module elliptic (
	PCLK, PRESET, Preset_0_0_, Pinp_0_0_, Pinp_1_1_, Pinp_2_2_, Pinp_3_3_, Pinp_4_4_, 
	Pinp_5_5_, Pinp_6_6_, Pinp_7_7_, Pinp_8_8_, Pinp_9_9_, Pinp_10_10_, Pinp_11_11_, Pinp_12_12_, Pinp_13_13_, Pinp_14_14_, 
	Pinp_15_15_, PDN, Pover_0_0_);

input PCLK, PRESET, Preset_0_0_, Pinp_0_0_, Pinp_1_1_, Pinp_2_2_, Pinp_3_3_, Pinp_4_4_, Pinp_5_5_, Pinp_6_6_, Pinp_7_7_, Pinp_8_8_, Pinp_9_9_, Pinp_10_10_, Pinp_11_11_, Pinp_12_12_, Pinp_13_13_, Pinp_14_14_, Pinp_15_15_;

output PDN, Pover_0_0_;

wire N_N9620, n16, N_N9577, n22, N_N9551, N_N9549, N_N9543, N_N9538, N_N9509, n41, N_N9461, N_N9443, N_N9425, N_N9409, N_N9330, N_N9328, N_N9297, N_N9295, N_N9293, N_N9279, N_N9274, N_N9243, N_N9241, N_N9149, n103, N_N9111, n126, N_N9039, N_N9012, N_N8971, N_N8969, N_N8967, N_N8952, N_N8934, n156, N_N8926, n157, N_N8922, N_N8874, n191, N_N8829, n193, N_N8825, n196, N_N8814, N_N8802, N_N8795, N_N8755, N_N8737, n227, N_N8722, N_N8709, N_N8690, N_N8684, N_N8614, N_N8612, N_N8576, N_N8565, N_N8540, N_N8527, N_N8507, N_N8478, n315, N_N8451, N_N8446, N_N8399, n338, N_N8385, N_N8365, N_N8364, N_N8363, n349, N_N8356, N_N8347, N_N8345, n360, N_N8317, N_N8311, n365, N_N8299, N_N8293, n370, N_N8286, n371, N_N8283, N_N8217, N_N8190, n404, N_N8181, N_N8178, N_N8172, N_N8170, N_N8169, n413, N_N8147, N_N8140, N_N8137, N_N8136, N_N8122, N_N8117, N_N8036, N_N8025, N_N8015, N_N7998, N_N7984, N_N7982, N_N7981, N_N7960, N_N7957, N_N7894, N_N7893, n486, N_N7891, N_N7883, N_N7870, n501, N_N7828, N_N7799, N_N7796, N_N7795, N_N7785, n515, N_N7750, n516, N_N7747, N_N7690, N_N7633, N_N7608, n571, N_N7574, N_N7548, N_N7547, n584, N_N7538, n585, N_N7535, n590, N_N7529, N_N7528, N_N7515, n625, N_N7477, n626, N_N7475, N_N7470, N_N7465, N_N7460, N_N7451, N_N7450, N_N7449, N_N7448, N_N7447, N_N7446, n640, N_N7439, N_N7397, N_N7382, N_N7379, N_N7377, N_N7371, N_N7357, N_N7318, N_N7313, N_N7312, N_N7305, N_N7301, N_N7294, N_N7280, N_N7266, N_N7238, N_N7232, N_N7194, n778, N_N7193, N_N7188, N_N7163, N_N7162, N_N7158, N_N7137, N_N7132, N_N7131, N_N7126, N_N7096, n834, N_N7095, n835, N_N7094, N_N7087, N_N7077, N_N7063, n861, N_N7059, N_N7048, N_N7047, N_N7042, n874, N_N7038, n880, N_N7030, N_N7015, N_N7007, N_N7006, N_N7001, N_N7000, N_N6995, N_N6982, N_N6971, N_N6958, N_N6957, N_N6942, N_N6941, n942, N_N6928, N_N6927, N_N6926, N_N6924, N_N6917, n955, N_N11, n956, N_N10, n957, N_N9, n958, N_N8, n959, N_N7, n960, N_N6, n961, N_N5, n962, N_N4, n963, N_N3, n964, N_N2, n965, N_N1, n966, N_N0, n1323, n1347, n1348, n1349, n1350, n1346, n1352, n1353, n1354, n1355, n1351, n1357, n1358, n1359, n1360, n1356, n1362, n1363, n1364, n1365, n1361, n1367, n1368, n1369, n1370, n1366, n1372, n1373, n1374, n1375, n1371, n1377, n1378, n1379, n1380, n1376, n1382, n1383, n1384, n1385, n1381, n1387, n1388, n1389, n1390, n1386, n1392, n1393, n1394, n1395, n1391, n1397, n1398, n1399, n1400, n1396, n1402, n1403, n1404, n1405, n1401, n1407, n1408, n1409, n1410, n1406, n1412, n1413, n1414, n1415, n1411, n1417, n1418, n1419, n1420, n1416, n1422, n1423, n1424, n1425, n1421, n1503, n1500, n1507, n1504, n1511, n1508, n1515, n1512, n1519, n1516, n1522, n1520, n1526, n1523, n1530, n1527, n1534, n1531, n1538, n1535, n1542, n1539, n1546, n1543, n1550, n1547, n1608, n1607, n1799, n1800, n1798, n1802, n1801, n1806, n1805, n1804, n1807, n1809, n1808, n1826, n1855, n2066, n2065, n2064, n2080, n2079, n2093, n2099, n2106, n2105, n2104, n2109, n2108, n2143, n2142, n2247, n2269, n2268, n2283, n2282, n2285, n2284, n2364, n2363, n2366, n2365, n2373, n2419, n2434, n2433, n2649, n2648, n2651, n2650, n2693, n2782, N_N7729, n2787, N_N7199, n2789, n2819, N_N7098, n2838, n2845, n2847, n2849, n2851, n2853, n2855, n2857, n2858, n2977, n2979, n3007, n3008, n3010, n3011, n3111, n3112, n3115, n3118, n3132, n3133, n3136;

reg N_N8199, N_N9280, N_N8803, N_N8240, N_N8274, N_N8198, N_N8239, N_N8615, N_N7703, N_N8273, N_N8366, N_N8272, N_N8238, N_N8531, N_N7983, N_N8575, N_N7854, N_N8237, N_N8197, N_N8271, N_N8530, N_N8650, N_N7985, N_N8710, N_N8574, N_N8312, N_N8270, N_N8573, N_N8935, N_N8649, N_N8196, N_N8236, N_N9244, N_N8348, N_N9150, N_N8648, N_N8269, N_N8235, N_N9275, N_N8970, N_N9554, N_N9013, N_N8508, N_N8529, N_N9242, N_N8572, N_N8571, N_N9436, N_N8528, N_N8796, N_N7770, N_N9357, N_N8685, N_N9296, N_N9555, N_N7628, N_N9510, N_N9578, N_N8447, N_N9437, N_N7771, N_N8570, N_N8647, N_N7704, N_N8646, N_N7629, NDN3_11, NDN3_12, N_N8037, NDN3_16, NDN3_17, NDN3_19, NDN3_22, NDN3_25, NDN3_26, N_N7584, NDN3_28, NDN3_29, NDN3_40, NDN3_39, NDN3_42, NDN3_44, NDN3_46, N_N9358, N_N9539, N_N9556, N_N7306, NEN3_16, N_N9160, NEN3_19, NEN3_22, N_N8930, NEN3_28, N_N9438, NEN3_34, NEN3_36, NEN3_39, N_N7961, NLC1_2, N_N9359, N_N7476, N_N8577, N_N9289, N_N9557, N_N7630, N_N9161, N_N8691, N_N9439, N_N8798, N_N8869, N_N9360, N_N8911, N_N9290, N_N9558, N_N8993, N_N9162, N_N9034, N_N9440, N_N9361, N_N9298, N_N9559, N_N9163, N_N9550, PDN, N_N8171, N_N8173, N_N9011, N_N9552, N_N7701, N_N8964, N_N9291, N_N9560, N_N7627, N_N8913, N_N8756, N_N9164, N_N8016, N_N9441, N_N8847, N_N8631, N_N9362, Pover_0_0_, NDN1_4, N_N8561, N_N9292, N_N9561, NGFDN_3, N_N9165, N_N9442, N_N7768, N_N8118, NDN2_2, N_N8875, N_N7852, N_N7582, N_N9331, N_N9363, N_N9294, NDN3_2, NDN3_4, NDN3_7, NDN3_9, N_N9410, N_N8613, N_N8972, N_N9247, N_N9166, N_N8968, NAK3_13, N_N8668, N_N8923, N_N7769, N_N8933, N_N7702, N_N8978, N_N8141, N_N8200, N_N8929, N_N7853, N_N9031, N_N8241, N_N7583, NSr3_13, N_N9248, NSr3_14, NSr3_20, N_N9198, NSr3_23, NSr3_30, NSr3_35, NSr3_37, NSr3_38, NSr1_2, N_N8603;

always  @(posedge PCLK)
	N_N8199<=N_N8025;

 always  @(posedge PCLK)
	N_N9280<=N_N9279;

 always  @(posedge PCLK)
	N_N8803<=N_N8802;

 always  @(posedge PCLK)
	N_N8240<=N_N7548;

 always  @(posedge PCLK)
	N_N8274<=N_N6924;

 always  @(posedge PCLK)
	N_N8198<=N_N7048;

 always  @(posedge PCLK)
	N_N8239<=N_N7371;

 always  @(posedge PCLK)
	N_N8615<=N_N8614;

 always  @(posedge PCLK)
	N_N7703<=N_N7294;

 always  @(posedge PCLK)
	N_N8273<=N_N7007;

 always  @(posedge PCLK)
	N_N8366<=N_N8365;

 always  @(posedge PCLK)
	N_N8272<=N_N7894;

 always  @(posedge PCLK)
	N_N8238<=N_N6941;

 always  @(posedge PCLK)
	N_N8531<=N_N7547;

 always  @(posedge PCLK)
	N_N7983<=N_N7982;

 always  @(posedge PCLK)
	N_N8575<=N_N7131;

 always  @(posedge PCLK)
	N_N7854<=N_N7000;

 always  @(posedge PCLK)
	N_N8237<=N_N7633;

 always  @(posedge PCLK)
	N_N8197<=N_N7447;

 always  @(posedge PCLK)
	N_N8271<=N_N7047;

 always  @(posedge PCLK)
	N_N8530<=N_N6982;

 always  @(posedge PCLK)
	N_N8650<=N_N7785;

 always  @(posedge PCLK)
	N_N7985<=N_N7984;

 always  @(posedge PCLK)
	N_N8710<=N_N8709;

 always  @(posedge PCLK)
	N_N8574<=N_N7006;

 always  @(posedge PCLK)
	N_N8312<=N_N8311;

 always  @(posedge PCLK)
	N_N8270<=N_N8190;

 always  @(posedge PCLK)
	N_N8573<=N_N7063;

 always  @(posedge PCLK)
	N_N8935<=N_N8934;

 always  @(posedge PCLK)
	N_N8649<=N_N7280;

 always  @(posedge PCLK)
	N_N8196<=N_N7893;

 always  @(posedge PCLK)
	N_N8236<=N_N8137;

 always  @(posedge PCLK)
	N_N9244<=N_N9243;

 always  @(posedge PCLK)
	N_N8348<=N_N8347;

 always  @(posedge PCLK)
	N_N9150<=N_N9149;

 always  @(posedge PCLK)
	N_N8648<=N_N7194;

 always  @(posedge PCLK)
	N_N8269<=N_N7313;

 always  @(posedge PCLK)
	N_N8235<=N_N7465;

 always  @(posedge PCLK)
	N_N9275<=N_N9274;

 always  @(posedge PCLK)
	N_N8970<=N_N8969;

 always  @(posedge PCLK)
	N_N9554<=N_N7266;

 always  @(posedge PCLK)
	N_N9013<=N_N9012;

 always  @(posedge PCLK)
	N_N8508<=N_N8507;

 always  @(posedge PCLK)
	N_N8529<=N_N8136;

 always  @(posedge PCLK)
	N_N9242<=N_N9241;

 always  @(posedge PCLK)
	N_N8572<=N_N8169;

 always  @(posedge PCLK)
	N_N8571<=N_N7312;

 always  @(posedge PCLK)
	N_N9436<=N_N8363;

 always  @(posedge PCLK)
	N_N8528<=N_N7377;

 always  @(posedge PCLK)
	N_N8796<=N_N8795;

 always  @(posedge PCLK)
	N_N7770<=N_N7001;

 always  @(posedge PCLK)
	N_N9357<=N_N8364;

 always  @(posedge PCLK)
	N_N8685<=N_N8684;

 always  @(posedge PCLK)
	N_N9296<=N_N9295;

 always  @(posedge PCLK)
	N_N9555<=N_N6995;

 always  @(posedge PCLK)
	N_N7628<=N_N6971;

 always  @(posedge PCLK)
	N_N9510<=N_N9509;

 always  @(posedge PCLK)
	N_N9578<=N_N9577;

 always  @(posedge PCLK)
	N_N8447<=N_N8446;

 always  @(posedge PCLK)
	N_N9437<=N_N7137;

 always  @(posedge PCLK)
	N_N7771<=N_N7042;

 always  @(posedge PCLK)
	N_N8570<=N_N7305;

 always  @(posedge PCLK)
	N_N8647<=N_N8527;

 always  @(posedge PCLK)
	N_N7704<=N_N6957;

 always  @(posedge PCLK)
	N_N8646<=N_N6926;

 always  @(posedge PCLK)
	N_N7629<=N_N6958;

 always  @(posedge PCLK)
	NDN3_11<=N_N7096;

 always  @(posedge PCLK)
	NDN3_12<=N_N7460;

 always  @(posedge PCLK)
	N_N8037<=N_N8036;

 always  @(posedge PCLK)
	NDN3_16<=N_N8540;

 always  @(posedge PCLK)
	NDN3_17<=N_N7087;

 always  @(posedge PCLK)
	NDN3_19<=N_N9543;

 always  @(posedge PCLK)
	NDN3_22<=N_N7883;

 always  @(posedge PCLK)
	NDN3_25<=N_N8293;

 always  @(posedge PCLK)
	NDN3_26<=N_N9328;

 always  @(posedge PCLK)
	N_N7584<=N_N7301;

 always  @(posedge PCLK)
	NDN3_28<=N_N9620;

 always  @(posedge PCLK)
	NDN3_29<=N_N8217;

 always  @(posedge PCLK)
	NDN3_40<=N_N7158;

 always  @(posedge PCLK)
	NDN3_39<=N_N9425;

 always  @(posedge PCLK)
	NDN3_42<=N_N7690;

 always  @(posedge PCLK)
	NDN3_44<=N_N7232;

 always  @(posedge PCLK)
	NDN3_46<=N_N7574;

 always  @(posedge PCLK)
	N_N9358<=N_N7608;

 always  @(posedge PCLK)
	N_N9539<=N_N9538;

 always  @(posedge PCLK)
	N_N9556<=N_N7795;

 always  @(posedge PCLK)
	N_N7306<=N_N8147;

 always  @(posedge PCLK)
	NEN3_16<=N_N7038;

 always  @(posedge PCLK)
	N_N9160<=N_N9111;

 always  @(posedge PCLK)
	NEN3_19<=N_N7477;

 always  @(posedge PCLK)
	NEN3_22<=N_N8299;

 always  @(posedge PCLK)
	N_N8930<=N_N7077;

 always  @(posedge PCLK)
	NEN3_28<=N_N7529;

 always  @(posedge PCLK)
	N_N9438<=N_N7796;

 always  @(posedge PCLK)
	NEN3_34<=N_N8825;

 always  @(posedge PCLK)
	NEN3_36<=N_N7891;

 always  @(posedge PCLK)
	NEN3_39<=N_N8317;

 always  @(posedge PCLK)
	N_N7961<=N_N7960;

 always  @(posedge PCLK)
	NLC1_2<=N_N8814;

 always  @(posedge PCLK)
	N_N9359<=N_N7126;

 always  @(posedge PCLK)
	N_N7476<=N_N7475;

 always  @(posedge PCLK)
	N_N8577<=N_N8576;

 always  @(posedge PCLK)
	N_N9289<=N_N8178;

 always  @(posedge PCLK)
	N_N9557<=N_N7397;

 always  @(posedge PCLK)
	N_N7630<=N_N7238;

 always  @(posedge PCLK)
	N_N9161<=N_N8829;

 always  @(posedge PCLK)
	N_N8691<=N_N8690;

 always  @(posedge PCLK)
	N_N9439<=N_N7449;

 always  @(posedge PCLK)
	N_N8798<=N_N7747;

 always  @(posedge PCLK)
	N_N8869<=N_N7750;

 always  @(posedge PCLK)
	N_N9360<=N_N7450;

 always  @(posedge PCLK)
	N_N8911<=N_N7535;

 always  @(posedge PCLK)
	N_N9290<=N_N7451;

 always  @(posedge PCLK)
	N_N9558<=N_N6942;

 always  @(posedge PCLK)
	N_N8993<=N_N8181;

 always  @(posedge PCLK)
	N_N9162<=N_N9039;

 always  @(posedge PCLK)
	N_N9034<=N_N7538;

 always  @(posedge PCLK)
	N_N9440<=N_N7998;

 always  @(posedge PCLK)
	N_N9361<=N_N7799;

 always  @(posedge PCLK)
	N_N9298<=N_N9297;

 always  @(posedge PCLK)
	N_N9559<=N_N8737;

 always  @(posedge PCLK)
	N_N9163<=N_N7193;

 always  @(posedge PCLK)
	N_N9550<=N_N9549;

 always  @(posedge PCLK)
	PDN<=N_N7729;

 always  @(posedge PCLK)
	N_N8171<=N_N8170;

 always  @(posedge PCLK)
	N_N8173<=N_N8172;

 always  @(posedge PCLK)
	N_N9011<=N_N8385;

 always  @(posedge PCLK)
	N_N9552<=N_N9551;

 always  @(posedge PCLK)
	N_N7701<=N_N7515;

 always  @(posedge PCLK)
	N_N8964<=N_N8286;

 always  @(posedge PCLK)
	N_N9291<=N_N7957;

 always  @(posedge PCLK)
	N_N9560<=N_N8345;

 always  @(posedge PCLK)
	N_N7627<=N_N6917;

 always  @(posedge PCLK)
	N_N8913<=N_N7095;

 always  @(posedge PCLK)
	N_N8756<=N_N8755;

 always  @(posedge PCLK)
	N_N9164<=N_N7059;

 always  @(posedge PCLK)
	N_N8016<=N_N8015;

 always  @(posedge PCLK)
	N_N9441<=N_N8952;

 always  @(posedge PCLK)
	N_N8847<=N_N8283;

 always  @(posedge PCLK)
	N_N8631<=N_N7094;

 always  @(posedge PCLK)
	N_N9362<=N_N7870;

 always  @(posedge PCLK)
	Pover_0_0_<=N_N7199;

 always  @(posedge PCLK)
	NDN1_4<=N_N7015;

 always  @(posedge PCLK)
	N_N8561<=N_N7439;

 always  @(posedge PCLK)
	N_N9292<=N_N6927;

 always  @(posedge PCLK)
	N_N9561<=N_N7470;

 always  @(posedge PCLK)
	NGFDN_3<=N_N7098;

 always  @(posedge PCLK)
	N_N9165<=N_N6928;

 always  @(posedge PCLK)
	N_N9442<=N_N7382;

 always  @(posedge PCLK)
	N_N7768<=N_N7528;

 always  @(posedge PCLK)
	N_N8118<=N_N8117;

 always  @(posedge PCLK)
	NDN2_2<=N_N8122;

 always  @(posedge PCLK)
	N_N8875<=N_N8874;

 always  @(posedge PCLK)
	N_N7852<=N_N7448;

 always  @(posedge PCLK)
	N_N7582<=N_N7318;

 always  @(posedge PCLK)
	N_N9331<=N_N9330;

 always  @(posedge PCLK)
	N_N9363<=N_N7981;

 always  @(posedge PCLK)
	N_N9294<=N_N9293;

 always  @(posedge PCLK)
	NDN3_2<=N_N9443;

 always  @(posedge PCLK)
	NDN3_4<=N_N8565;

 always  @(posedge PCLK)
	NDN3_7<=N_N8399;

 always  @(posedge PCLK)
	NDN3_9<=N_N7188;

 always  @(posedge PCLK)
	N_N9410<=N_N9409;

 always  @(posedge PCLK)
	N_N8613<=N_N8612;

 always  @(posedge PCLK)
	N_N8972<=N_N8971;

 always  @(posedge PCLK)
	N_N9247<=N_N9461;

 always  @(posedge PCLK)
	N_N9166<=N_N7030;

 always  @(posedge PCLK)
	N_N8968<=N_N8967;

 always  @(posedge PCLK)
	NAK3_13<=N_N8478;

 always  @(posedge PCLK)
	N_N8668<=N_N8451;

 always  @(posedge PCLK)
	N_N8923<=N_N8922;

 always  @(posedge PCLK)
	N_N7769<=N_N7162;

 always  @(posedge PCLK)
	N_N8933<=N_N8926;

 always  @(posedge PCLK)
	N_N7702<=N_N7163;

 always  @(posedge PCLK)
	N_N8978<=N_N7828;

 always  @(posedge PCLK)
	N_N8141<=N_N8140;

 always  @(posedge PCLK)
	N_N8200<=N_N7132;

 always  @(posedge PCLK)
	N_N8929<=N_N8722;

 always  @(posedge PCLK)
	N_N7853<=N_N7446;

 always  @(posedge PCLK)
	N_N9031<=N_N8356;

 always  @(posedge PCLK)
	N_N8241<=N_N7379;

 always  @(posedge PCLK)
	N_N7583<=N_N7357;

 always  @(posedge PCLK)
	NSr3_13<=N_N11;

 always  @(posedge PCLK)
	N_N9248<=N_N10;

 always  @(posedge PCLK)
	NSr3_14<=N_N9;

 always  @(posedge PCLK)
	NSr3_20<=N_N8;

 always  @(posedge PCLK)
	N_N9198<=N_N7;

 always  @(posedge PCLK)
	NSr3_23<=N_N6;

 always  @(posedge PCLK)
	NSr3_30<=N_N5;

 always  @(posedge PCLK)
	NSr3_35<=N_N4;

 always  @(posedge PCLK)
	NSr3_37<=N_N3;

 always  @(posedge PCLK)
	NSr3_38<=N_N2;

 always  @(posedge PCLK)
	NSr1_2<=N_N1;

 always  @(posedge PCLK)
	N_N8603<=N_N0;

 assign N_N9620 = ( NEN3_28  &  (~ n1826) ) | ( NDN3_28  &  (~ n1826) ) ;
 assign n16 = ( PRESET  &  n1323 ) | ( n1323  &  (~ N_N9578) ) ;
 assign N_N9577 = ( (~ n16) ) ;
 assign n22 = ( (~ PRESET)  &  n2838 ) ;
 assign N_N9551 = ( N_N9552  &  n22 ) ;
 assign N_N9549 = ( N_N9550  &  n22 ) ;
 assign N_N9543 = ( NDN3_19  &  (~ n1826) ) | ( NEN3_19  &  (~ n1826) ) ;
 assign N_N9538 = ( N_N9539  &  n22 ) ;
 assign N_N9509 = ( N_N9510  &  n22 ) ;
 assign n41 = ( (~ PRESET)  &  n3115 ) | ( (~ PRESET)  &  (~ n413)  &  N_N9247 ) ;
 assign N_N9461 = ( n41  &  N_N9248 ) ;
 assign N_N9443 = ( NDN3_2  &  (~ n1826) ) | ( (~ n1607)  &  (~ n1826) ) ;
 assign N_N9425 = ( NDN3_39  &  (~ n1826) ) | ( NEN3_39  &  (~ n1826) ) ;
 assign N_N9409 = ( N_N9410  &  n22 ) ;
 assign N_N9330 = ( N_N9331  &  n22 ) ;
 assign N_N9328 = ( NDN3_26  &  (~ n1826) ) | ( NDN3_25  &  (~ n1826) ) ;
 assign N_N9297 = ( N_N9298  &  n22 ) ;
 assign N_N9295 = ( N_N9296  &  n22 ) ;
 assign N_N9293 = ( N_N9294  &  n22 ) ;
 assign N_N9279 = ( N_N9280  &  n22 ) ;
 assign N_N9274 = ( N_N9275  &  n22 ) ;
 assign N_N9243 = ( N_N9244  &  n22 ) ;
 assign N_N9241 = ( N_N9242  &  n22 ) ;
 assign N_N9149 = ( N_N9150  &  n22 ) ;
 assign n103 = ( PRESET  &  n1323 ) | ( n1323  &  (~ N_N9160) ) ;
 assign N_N9111 = ( (~ n103) ) ;
 assign n126 = ( PRESET  &  n1323 ) | ( n1323  &  (~ N_N9162) ) ;
 assign N_N9039 = ( (~ n126) ) ;
 assign N_N9012 = ( N_N9013  &  n22 ) ;
 assign N_N8971 = ( N_N8972  &  n22 ) ;
 assign N_N8969 = ( N_N8970  &  n22 ) ;
 assign N_N8967 = ( N_N8968  &  n22 ) ;
 assign N_N8952 = ( N_N9441  &  n22 ) ;
 assign N_N8934 = ( N_N8935  &  n22 ) ;
 assign n156 = ( PRESET  &  n1807 ) | ( n1804  &  n1807 ) | ( PRESET  &  (~ N_N8933) ) | ( n1804  &  (~ N_N8933) ) ;
 assign N_N8926 = ( (~ n156) ) ;
 assign n157 = ( PRESET  &  n1807 ) | ( n1807  &  n1808 ) | ( PRESET  &  (~ N_N8923) ) | ( n1808  &  (~ N_N8923) ) ;
 assign N_N8922 = ( (~ n157) ) ;
 assign N_N8874 = ( N_N8875  &  n22 ) ;
 assign n191 = ( PRESET  &  n1323 ) | ( n1323  &  (~ N_N9161) ) ;
 assign N_N8829 = ( (~ n191) ) ;
 assign n193 = ( (~ NEN3_34)  &  NGFDN_3 ) | ( n1826  &  NGFDN_3 ) | ( (~ NEN3_34)  &  n1855 ) | ( n1826  &  n1855 ) ;
 assign N_N8825 = ( (~ n193) ) ;
 assign n196 = ( (~ PRESET)  &  (~ PDN) ) ;
 assign N_N8814 = ( n196  &  NLC1_2 ) | ( n196  &  NSr1_2 ) ;
 assign N_N8802 = ( N_N8803  &  n22 ) ;
 assign N_N8795 = ( N_N8796  &  n22 ) ;
 assign N_N8755 = ( N_N8756  &  n22 ) ;
 assign N_N8737 = ( N_N9559  &  n22 ) ;
 assign n227 = ( N_N9198  &  (~ n1799)  &  n1800 ) ;
 assign N_N8722 = ( (~ PRESET)  &  N_N8929 ) | ( (~ PRESET)  &  n227 ) ;
 assign N_N8709 = ( N_N8710  &  n22 ) ;
 assign N_N8690 = ( N_N8691  &  n22 ) ;
 assign N_N8684 = ( N_N8685  &  n22 ) ;
 assign N_N8614 = ( N_N8615  &  n22 ) ;
 assign N_N8612 = ( N_N8613  &  n22 ) ;
 assign N_N8576 = ( N_N8577  &  n22 ) ;
 assign N_N8565 = ( NDN3_2  &  (~ n1826) ) | ( NDN3_4  &  (~ n1826) ) ;
 assign N_N8540 = ( NDN3_16  &  (~ n1826) ) | ( NEN3_16  &  (~ n1826) ) ;
 assign N_N8527 = ( N_N8647  &  n22 ) ;
 assign N_N8507 = ( N_N8508  &  n22 ) ;
 assign N_N8478 = ( (~ PRESET)  &  (~ n1798) ) ;
 assign n315 = ( (~ PRESET)  &  n1798 ) ;
 assign N_N8451 = ( N_N8668  &  n315 ) ;
 assign N_N8446 = ( N_N8447  &  n22 ) ;
 assign N_N8399 = ( NDN3_4  &  (~ n1826) ) | ( NDN3_7  &  (~ n1826) ) ;
 assign n338 = ( PRESET  &  n1807 ) | ( n1807  &  n2064 ) | ( PRESET  &  (~ N_N9011) ) | ( n2064  &  (~ N_N9011) ) ;
 assign N_N8385 = ( (~ n338) ) ;
 assign N_N8365 = ( N_N8366  &  n22 ) ;
 assign N_N8364 = ( N_N9357  &  n22 ) ;
 assign N_N8363 = ( N_N9436  &  n22 ) ;
 assign n349 = ( PRESET  &  n1807 ) | ( n1807  &  n2079 ) | ( PRESET  &  (~ N_N9031) ) | ( n2079  &  (~ N_N9031) ) ;
 assign N_N8356 = ( (~ n349) ) ;
 assign N_N8347 = ( N_N8348  &  n22 ) ;
 assign N_N8345 = ( N_N9560  &  n22 ) ;
 assign n360 = ( (~ NEN3_39)  &  NGFDN_3 ) | ( n1826  &  NGFDN_3 ) | ( (~ NEN3_39)  &  n2093 ) | ( n1826  &  n2093 ) ;
 assign N_N8317 = ( (~ n360) ) ;
 assign N_N8311 = ( N_N8312  &  n22 ) ;
 assign n365 = ( (~ NEN3_22)  &  NGFDN_3 ) | ( n1826  &  NGFDN_3 ) | ( (~ NEN3_22)  &  n2099 ) | ( n1826  &  n2099 ) ;
 assign N_N8299 = ( (~ n365) ) ;
 assign N_N8293 = ( NDN3_25  &  (~ n1826) ) | ( NDN3_22  &  (~ n1826) ) ;
 assign n370 = ( PRESET  &  n1807 ) | ( n1807  &  n2104 ) | ( PRESET  &  (~ N_N8964) ) | ( n2104  &  (~ N_N8964) ) ;
 assign N_N8286 = ( (~ n370) ) ;
 assign n371 = ( PRESET  &  n1807 ) | ( n1807  &  n2108 ) | ( PRESET  &  (~ N_N8847) ) | ( n2108  &  (~ N_N8847) ) ;
 assign N_N8283 = ( (~ n371) ) ;
 assign N_N8217 = ( NDN3_28  &  (~ n1826) ) | ( NDN3_29  &  (~ n1826) ) ;
 assign N_N8190 = ( N_N8270  &  n22 ) ;
 assign n404 = ( PRESET  &  n1807 ) | ( n1807  &  n2142 ) | ( PRESET  &  (~ N_N8993) ) | ( n2142  &  (~ N_N8993) ) ;
 assign N_N8181 = ( (~ n404) ) ;
 assign N_N8178 = ( N_N9289  &  n22 ) ;
 assign N_N8172 = ( N_N8173  &  n22 ) ;
 assign N_N8170 = ( N_N8171  &  n22 ) ;
 assign N_N8169 = ( N_N8572  &  n22 ) ;
 assign n413 = ( n1500  &  n2105  &  n1508  &  n1504  &  n1516  &  n1512  &  n3010  &  n3011 ) ;
 assign N_N8147 = ( (~ PRESET)  &  n413 ) ;
 assign N_N8140 = ( N_N8141  &  n22 ) ;
 assign N_N8137 = ( N_N8236  &  n22 ) ;
 assign N_N8136 = ( N_N8529  &  n22 ) ;
 assign N_N8122 = ( (~ PRESET)  &  NDN2_2  &  (~ n2782) ) ;
 assign N_N8117 = ( N_N8118  &  n22 ) ;
 assign N_N8036 = ( N_N8037  &  n22 ) ;
 assign N_N8025 = ( N_N8199  &  n22 ) ;
 assign N_N8015 = ( N_N8016  &  n22 ) ;
 assign N_N7998 = ( N_N9440  &  n22 ) ;
 assign N_N7984 = ( N_N7985  &  n22 ) ;
 assign N_N7982 = ( N_N7983  &  n22 ) ;
 assign N_N7981 = ( N_N9363  &  n22 ) ;
 assign N_N7960 = ( N_N7961  &  n22 ) ;
 assign N_N7957 = ( N_N9291  &  n22 ) ;
 assign N_N7894 = ( N_N8272  &  n22 ) ;
 assign N_N7893 = ( N_N8196  &  n22 ) ;
 assign n486 = ( (~ NEN3_36)  &  NGFDN_3 ) | ( n1826  &  NGFDN_3 ) | ( (~ NEN3_36)  &  n2247 ) | ( n1826  &  n2247 ) ;
 assign N_N7891 = ( (~ n486) ) ;
 assign N_N7883 = ( NDN3_22  &  (~ n1826) ) | ( NEN3_22  &  (~ n1826) ) ;
 assign N_N7870 = ( N_N9362  &  n22 ) ;
 assign n501 = ( PRESET  &  n1807 ) | ( n1807  &  n2268 ) | ( PRESET  &  (~ N_N8978) ) | ( n2268  &  (~ N_N8978) ) ;
 assign N_N7828 = ( (~ n501) ) ;
 assign N_N7799 = ( N_N9361  &  n22 ) ;
 assign N_N7796 = ( N_N9438  &  n22 ) ;
 assign N_N7795 = ( N_N9556  &  n22 ) ;
 assign N_N7785 = ( N_N8650  &  n22 ) ;
 assign n515 = ( PRESET  &  n1807 ) | ( n1807  &  n2282 ) | ( PRESET  &  (~ N_N8869) ) | ( n2282  &  (~ N_N8869) ) ;
 assign N_N7750 = ( (~ n515) ) ;
 assign n516 = ( PRESET  &  n1807 ) | ( n1807  &  n2284 ) | ( PRESET  &  (~ N_N8798) ) | ( n2284  &  (~ N_N8798) ) ;
 assign N_N7747 = ( (~ n516) ) ;
 assign N_N7690 = ( NDN3_42  &  (~ n1826) ) | ( NDN3_40  &  (~ n1826) ) ;
 assign N_N7633 = ( N_N8237  &  n22 ) ;
 assign N_N7608 = ( N_N9358  &  n22 ) ;
 assign n571 = ( (~ NDN3_44)  &  (~ N_N7098) ) | ( n1826  &  (~ N_N7098) ) ;
 assign N_N7574 = ( (~ n571) ) ;
 assign N_N7548 = ( N_N8240  &  n22 ) ;
 assign N_N7547 = ( N_N8531  &  n22 ) ;
 assign n584 = ( PRESET  &  n1807 ) | ( n1807  &  n2363 ) | ( PRESET  &  (~ N_N9034) ) | ( n2363  &  (~ N_N9034) ) ;
 assign N_N7538 = ( (~ n584) ) ;
 assign n585 = ( PRESET  &  n1807 ) | ( n1807  &  n2365 ) | ( PRESET  &  (~ N_N8911) ) | ( n2365  &  (~ N_N8911) ) ;
 assign N_N7535 = ( (~ n585) ) ;
 assign n590 = ( (~ NEN3_28)  &  NGFDN_3 ) | ( n1826  &  NGFDN_3 ) | ( (~ NEN3_28)  &  n2373 ) | ( n1826  &  n2373 ) ;
 assign N_N7529 = ( (~ n590) ) ;
 assign N_N7528 = ( N_N7768  &  n22 ) ;
 assign N_N7515 = ( N_N7701  &  n22 ) ;
 assign n625 = ( (~ NEN3_19)  &  NGFDN_3 ) | ( n1826  &  NGFDN_3 ) | ( (~ NEN3_19)  &  n2419 ) | ( n1826  &  n2419 ) ;
 assign N_N7477 = ( (~ n625) ) ;
 assign n626 = ( (~ Preset_0_0_)  &  (~ n1608) ) | ( (~ Preset_0_0_)  &  N_N7476 ) | ( n1608  &  N_N7476 ) ;
 assign N_N7475 = ( (~ PRESET)  &  n626 ) ;
 assign N_N7470 = ( N_N9561  &  n22 ) ;
 assign N_N7465 = ( N_N8235  &  n22 ) ;
 assign N_N7460 = ( NDN3_11  &  (~ n1826) ) | ( NDN3_12  &  (~ n1826) ) ;
 assign N_N7451 = ( N_N9290  &  n22 ) ;
 assign N_N7450 = ( N_N9360  &  n22 ) ;
 assign N_N7449 = ( N_N9439  &  n22 ) ;
 assign N_N7448 = ( N_N7852  &  n22 ) ;
 assign N_N7447 = ( N_N8197  &  n22 ) ;
 assign N_N7446 = ( N_N7853  &  n22 ) ;
 assign n640 = ( PRESET  &  n1807 ) | ( n1807  &  n2433 ) | ( PRESET  &  (~ N_N8561) ) | ( n2433  &  (~ N_N8561) ) ;
 assign N_N7439 = ( (~ n640) ) ;
 assign N_N7397 = ( N_N9557  &  n22 ) ;
 assign N_N7382 = ( N_N9442  &  n22 ) ;
 assign N_N7379 = ( N_N8241  &  n22 ) ;
 assign N_N7377 = ( N_N8528  &  n22 ) ;
 assign N_N7371 = ( N_N8239  &  n22 ) ;
 assign N_N7357 = ( N_N7583  &  n22 ) ;
 assign N_N7318 = ( N_N7582  &  n22 ) ;
 assign N_N7313 = ( N_N8269  &  n22 ) ;
 assign N_N7312 = ( N_N8571  &  n22 ) ;
 assign N_N7305 = ( N_N8570  &  n22 ) ;
 assign N_N7301 = ( N_N7584  &  n22 ) ;
 assign N_N7294 = ( N_N7703  &  n22 ) ;
 assign N_N7280 = ( N_N8649  &  n22 ) ;
 assign N_N7266 = ( N_N9554  &  n22 ) ;
 assign N_N7238 = ( N_N7630  &  n22 ) ;
 assign N_N7232 = ( NDN3_42  &  (~ n1826) ) | ( NDN3_44  &  (~ n1826) ) ;
 assign N_N7194 = ( N_N8648  &  n22 ) ;
 assign n778 = ( PRESET  &  n1323 ) | ( n1323  &  (~ N_N9163) ) ;
 assign N_N7193 = ( (~ n778) ) ;
 assign N_N7188 = ( NDN3_7  &  (~ n1826) ) | ( NDN3_9  &  (~ n1826) ) ;
 assign N_N7163 = ( N_N7702  &  n22 ) ;
 assign N_N7162 = ( N_N7769  &  n22 ) ;
 assign N_N7158 = ( NDN3_39  &  (~ n1826) ) | ( NDN3_40  &  (~ n1826) ) ;
 assign N_N7137 = ( N_N9437  &  n22 ) ;
 assign N_N7132 = ( N_N8200  &  n22 ) ;
 assign N_N7131 = ( N_N8575  &  n22 ) ;
 assign N_N7126 = ( N_N9359  &  n22 ) ;
 assign N_N7096 = ( NDN3_11  &  (~ n1826) ) | ( NDN3_9  &  (~ n1826) ) ;
 assign n834 = ( PRESET  &  n1807 ) | ( n1807  &  n2648 ) | ( PRESET  &  (~ N_N8913) ) | ( n2648  &  (~ N_N8913) ) ;
 assign N_N7095 = ( (~ n834) ) ;
 assign n835 = ( PRESET  &  n1807 ) | ( n1807  &  n2650 ) | ( PRESET  &  (~ N_N8631) ) | ( n2650  &  (~ N_N8631) ) ;
 assign N_N7094 = ( (~ n835) ) ;
 assign N_N7087 = ( NDN3_16  &  (~ n1826) ) | ( NDN3_17  &  (~ n1826) ) ;
 assign N_N7077 = ( n315  &  n227 ) | ( n315  &  N_N8930 ) ;
 assign N_N7063 = ( N_N8573  &  n22 ) ;
 assign n861 = ( PRESET  &  n1323 ) | ( n1323  &  (~ N_N9164) ) ;
 assign N_N7059 = ( (~ n861) ) ;
 assign N_N7048 = ( N_N8198  &  n22 ) ;
 assign N_N7047 = ( N_N8271  &  n22 ) ;
 assign N_N7042 = ( N_N7771  &  n22 ) ;
 assign n874 = ( (~ NEN3_16)  &  NGFDN_3 ) | ( n1826  &  NGFDN_3 ) | ( (~ NEN3_16)  &  n2693 ) | ( n1826  &  n2693 ) ;
 assign N_N7038 = ( (~ n874) ) ;
 assign n880 = ( PRESET  &  n1323 ) | ( n1323  &  (~ N_N9166) ) ;
 assign N_N7030 = ( (~ n880) ) ;
 assign N_N7015 = ( NDN1_4  &  n196 ) ;
 assign N_N7007 = ( N_N8273  &  n22 ) ;
 assign N_N7006 = ( N_N8574  &  n22 ) ;
 assign N_N7001 = ( N_N7770  &  n22 ) ;
 assign N_N7000 = ( N_N7854  &  n22 ) ;
 assign N_N6995 = ( N_N9555  &  n22 ) ;
 assign N_N6982 = ( N_N8530  &  n22 ) ;
 assign N_N6971 = ( N_N7628  &  n22 ) ;
 assign N_N6958 = ( N_N7629  &  n22 ) ;
 assign N_N6957 = ( N_N7704  &  n22 ) ;
 assign N_N6942 = ( N_N9558  &  n22 ) ;
 assign N_N6941 = ( N_N8238  &  n22 ) ;
 assign n942 = ( PRESET  &  n1323 ) | ( n1323  &  (~ N_N9165) ) ;
 assign N_N6928 = ( (~ n942) ) ;
 assign N_N6927 = ( N_N9292  &  n22 ) ;
 assign N_N6926 = ( N_N8646  &  n22 ) ;
 assign N_N6924 = ( N_N8274  &  n22 ) ;
 assign N_N6917 = ( N_N7627  &  n22 ) ;
 assign n955 = ( n196  &  (~ NSr3_13) ) | ( n196  &  NDN3_12  &  NAK3_13 ) ;
 assign N_N11 = ( (~ n955) ) ;
 assign n956 = ( (~ N_N9248)  &  n315 ) | ( n315  &  n413 ) ;
 assign N_N10 = ( (~ n956) ) ;
 assign n957 = ( n196  &  (~ NSr3_14) ) | ( n196  &  NAK3_13  &  (~ NSr3_13) ) ;
 assign N_N9 = ( (~ n957) ) ;
 assign n958 = ( n196  &  (~ NSr3_20) ) | ( n196  &  NDN3_17  &  NAK3_13 ) ;
 assign N_N8 = ( (~ n958) ) ;
 assign n959 = ( (~ N_N9248)  &  n315  &  (~ n1799) ) | ( n315  &  n413  &  (~ n1799) ) ;
 assign N_N7 = ( (~ n959) ) ;
 assign n960 = ( n196  &  (~ NSr3_23) ) | ( NDN3_19  &  n196  &  NAK3_13 ) ;
 assign N_N6 = ( (~ n960) ) ;
 assign n961 = ( n196  &  (~ NSr3_30) ) | ( NDN3_26  &  n196  &  NAK3_13 ) ;
 assign N_N5 = ( (~ n961) ) ;
 assign n962 = ( n196  &  (~ NSr3_35) ) | ( n196  &  NDN3_29  &  NAK3_13 ) ;
 assign N_N4 = ( (~ n962) ) ;
 assign n963 = ( n196  &  (~ NSr3_37) ) | ( NEN3_34  &  n196  &  NAK3_13 ) ;
 assign N_N3 = ( (~ n963) ) ;
 assign n964 = ( n196  &  (~ NSr3_38) ) | ( NEN3_36  &  n196  &  NAK3_13 ) ;
 assign N_N2 = ( (~ n964) ) ;
 assign n965 = ( n196  &  (~ NSr1_2) ) | ( n196  &  NGFDN_3 ) | ( n196  &  n2782 ) ;
 assign N_N1 = ( (~ n965) ) ;
 assign n966 = ( (~ PRESET)  &  (~ N_N8603)  &  (~ n3133) ) | ( (~ PRESET)  &  (~ n3007)  &  (~ n3133) ) ;
 assign N_N0 = ( (~ n966) ) ;
 assign n1323 = ( PRESET ) | ( n2838 ) ;
 assign n1347 = ( (~ N_N9552)  &  (~ N_N9363) ) | ( (~ N_N9552)  &  (~ n2857) ) | ( (~ N_N9363)  &  n2858 ) | ( (~ n2857)  &  n2858 ) ;
 assign n1348 = ( (~ N_N9362)  &  (~ N_N9361) ) | ( (~ N_N9362)  &  n2853 ) | ( (~ N_N9361)  &  n2855 ) | ( n2853  &  n2855 ) ;
 assign n1349 = ( (~ N_N9360)  &  (~ N_N9359) ) | ( (~ N_N9360)  &  n2849 ) | ( (~ N_N9359)  &  n2851 ) | ( n2849  &  n2851 ) ;
 assign n1350 = ( (~ N_N9357)  &  (~ N_N9358) ) | ( (~ N_N9358)  &  n2845 ) | ( (~ N_N9357)  &  n2847 ) | ( n2845  &  n2847 ) ;
 assign n1346 = ( n1347  &  n1348  &  n1349  &  n1350 ) ;
 assign n1352 = ( (~ N_N9539)  &  (~ N_N9410) ) | ( (~ N_N9410)  &  n2847 ) | ( (~ N_N9539)  &  (~ n2857) ) | ( n2847  &  (~ n2857) ) ;
 assign n1353 = ( (~ N_N9298)  &  (~ N_N9296) ) | ( (~ N_N9298)  &  n2845 ) | ( (~ N_N9296)  &  n2853 ) | ( n2845  &  n2853 ) ;
 assign n1354 = ( (~ N_N9291)  &  (~ N_N9292) ) | ( (~ N_N9291)  &  n2855 ) | ( (~ N_N9292)  &  n2858 ) | ( n2855  &  n2858 ) ;
 assign n1355 = ( (~ N_N9289)  &  (~ N_N9290) ) | ( (~ N_N9290)  &  n2849 ) | ( (~ N_N9289)  &  n2851 ) | ( n2849  &  n2851 ) ;
 assign n1351 = ( n1352  &  n1353  &  n1354  &  n1355 ) ;
 assign n1357 = ( (~ N_N9578)  &  (~ n2857) ) | ( n2845  &  (~ n2857) ) | ( (~ N_N9578)  &  (~ N_N9166) ) | ( n2845  &  (~ N_N9166) ) ;
 assign n1358 = ( n2855  &  n2858 ) | ( n2855  &  (~ N_N9164) ) | ( n2858  &  (~ N_N9165) ) | ( (~ N_N9164)  &  (~ N_N9165) ) ;
 assign n1359 = ( n2851  &  n2853 ) | ( n2853  &  (~ N_N9162) ) | ( n2851  &  (~ N_N9163) ) | ( (~ N_N9162)  &  (~ N_N9163) ) ;
 assign n1360 = ( n2847  &  n2849 ) | ( n2849  &  (~ N_N9160) ) | ( n2847  &  (~ N_N9161) ) | ( (~ N_N9160)  &  (~ N_N9161) ) ;
 assign n1356 = ( n1357  &  n1358  &  n1359  &  n1360 ) ;
 assign n1362 = ( (~ N_N8875)  &  (~ N_N8613) ) | ( (~ N_N8613)  &  n2847 ) | ( (~ N_N8875)  &  n2849 ) | ( n2847  &  n2849 ) ;
 assign n1363 = ( (~ N_N8141)  &  (~ N_N7983) ) | ( (~ N_N7983)  &  n2851 ) | ( (~ N_N8141)  &  n2853 ) | ( n2851  &  n2853 ) ;
 assign n1364 = ( (~ N_N7630)  &  (~ N_N7629) ) | ( (~ N_N7630)  &  n2855 ) | ( (~ N_N7629)  &  (~ n2857) ) | ( n2855  &  (~ n2857) ) ;
 assign n1365 = ( (~ N_N7628)  &  (~ N_N7627) ) | ( (~ N_N7628)  &  n2845 ) | ( (~ N_N7627)  &  n2858 ) | ( n2845  &  n2858 ) ;
 assign n1361 = ( n1362  &  n1363  &  n1364  &  n1365 ) ;
 assign n1367 = ( (~ N_N8968)  &  (~ N_N8691) ) | ( (~ N_N8691)  &  n2849 ) | ( (~ N_N8968)  &  (~ n2857) ) | ( n2849  &  (~ n2857) ) ;
 assign n1368 = ( (~ N_N8447)  &  (~ N_N8016) ) | ( (~ N_N8447)  &  n2845 ) | ( (~ N_N8016)  &  n2858 ) | ( n2845  &  n2858 ) ;
 assign n1369 = ( (~ N_N7985)  &  (~ N_N7584) ) | ( (~ N_N7584)  &  n2853 ) | ( (~ N_N7985)  &  n2855 ) | ( n2853  &  n2855 ) ;
 assign n1370 = ( (~ N_N7583)  &  (~ N_N7582) ) | ( (~ N_N7583)  &  n2847 ) | ( (~ N_N7582)  &  n2851 ) | ( n2847  &  n2851 ) ;
 assign n1366 = ( n1367  &  n1368  &  n1369  &  n1370 ) ;
 assign n1372 = ( (~ N_N9294)  &  (~ N_N8685) ) | ( (~ N_N8685)  &  n2849 ) | ( (~ N_N9294)  &  n2858 ) | ( n2849  &  n2858 ) ;
 assign n1373 = ( (~ N_N8577)  &  (~ N_N8118) ) | ( (~ N_N8577)  &  n2847 ) | ( (~ N_N8118)  &  (~ n2857) ) | ( n2847  &  (~ n2857) ) ;
 assign n1374 = ( (~ N_N7703)  &  (~ N_N7704) ) | ( (~ N_N7704)  &  n2853 ) | ( (~ N_N7703)  &  n2855 ) | ( n2853  &  n2855 ) ;
 assign n1375 = ( (~ N_N7701)  &  (~ N_N7702) ) | ( (~ N_N7702)  &  n2845 ) | ( (~ N_N7701)  &  n2851 ) | ( n2845  &  n2851 ) ;
 assign n1371 = ( n1372  &  n1373  &  n1374  &  n1375 ) ;
 assign n1377 = ( (~ N_N9331)  &  (~ N_N8803) ) | ( (~ N_N8803)  &  n2849 ) | ( (~ N_N9331)  &  n2853 ) | ( n2849  &  n2853 ) ;
 assign n1378 = ( (~ N_N8173)  &  (~ N_N7961) ) | ( (~ N_N7961)  &  n2845 ) | ( (~ N_N8173)  &  (~ n2857) ) | ( n2845  &  (~ n2857) ) ;
 assign n1379 = ( (~ N_N7771)  &  (~ N_N7770) ) | ( (~ N_N7770)  &  n2855 ) | ( (~ N_N7771)  &  n2858 ) | ( n2855  &  n2858 ) ;
 assign n1380 = ( (~ N_N7768)  &  (~ N_N7769) ) | ( (~ N_N7769)  &  n2847 ) | ( (~ N_N7768)  &  n2851 ) | ( n2847  &  n2851 ) ;
 assign n1376 = ( n1377  &  n1378  &  n1379  &  n1380 ) ;
 assign n1382 = ( (~ N_N9560)  &  (~ N_N9561) ) | ( (~ N_N9561)  &  n2855 ) | ( (~ N_N9560)  &  (~ n2857) ) | ( n2855  &  (~ n2857) ) ;
 assign n1383 = ( (~ N_N9559)  &  (~ N_N9558) ) | ( (~ N_N9559)  &  n2853 ) | ( (~ N_N9558)  &  n2858 ) | ( n2853  &  n2858 ) ;
 assign n1384 = ( (~ N_N9556)  &  (~ N_N9557) ) | ( (~ N_N9557)  &  n2849 ) | ( (~ N_N9556)  &  n2851 ) | ( n2849  &  n2851 ) ;
 assign n1385 = ( (~ N_N9554)  &  (~ N_N9555) ) | ( (~ N_N9555)  &  n2845 ) | ( (~ N_N9554)  &  n2847 ) | ( n2845  &  n2847 ) ;
 assign n1381 = ( n1382  &  n1383  &  n1384  &  n1385 ) ;
 assign n1387 = ( (~ N_N9550)  &  (~ N_N9442) ) | ( (~ N_N9550)  &  (~ n2857) ) | ( (~ N_N9442)  &  n2858 ) | ( (~ n2857)  &  n2858 ) ;
 assign n1388 = ( (~ N_N9441)  &  (~ N_N9440) ) | ( (~ N_N9441)  &  n2853 ) | ( (~ N_N9440)  &  n2855 ) | ( n2853  &  n2855 ) ;
 assign n1389 = ( (~ N_N9438)  &  (~ N_N9439) ) | ( (~ N_N9439)  &  n2849 ) | ( (~ N_N9438)  &  n2851 ) | ( n2849  &  n2851 ) ;
 assign n1390 = ( (~ N_N9436)  &  (~ N_N9437) ) | ( (~ N_N9437)  &  n2845 ) | ( (~ N_N9436)  &  n2847 ) | ( n2845  &  n2847 ) ;
 assign n1386 = ( n1387  &  n1388  &  n1389  &  n1390 ) ;
 assign n1392 = ( (~ N_N8508)  &  (~ N_N8348) ) | ( (~ N_N8348)  &  n2845 ) | ( (~ N_N8508)  &  n2849 ) | ( n2845  &  n2849 ) ;
 assign n1393 = ( (~ N_N8273)  &  (~ N_N8274) ) | ( (~ N_N8274)  &  n2855 ) | ( (~ N_N8273)  &  (~ n2857) ) | ( n2855  &  (~ n2857) ) ;
 assign n1394 = ( (~ N_N8272)  &  (~ N_N8271) ) | ( (~ N_N8272)  &  n2853 ) | ( (~ N_N8271)  &  n2858 ) | ( n2853  &  n2858 ) ;
 assign n1395 = ( (~ N_N8270)  &  (~ N_N8269) ) | ( (~ N_N8270)  &  n2847 ) | ( (~ N_N8269)  &  n2851 ) | ( n2847  &  n2851 ) ;
 assign n1391 = ( n1392  &  n1393  &  n1394  &  n1395 ) ;
 assign n1397 = ( (~ N_N9280)  &  (~ N_N8710) ) | ( (~ N_N9280)  &  n2847 ) | ( (~ N_N8710)  &  n2858 ) | ( n2847  &  n2858 ) ;
 assign n1398 = ( (~ N_N8366)  &  (~ N_N8200) ) | ( (~ N_N8200)  &  n2851 ) | ( (~ N_N8366)  &  (~ n2857) ) | ( n2851  &  (~ n2857) ) ;
 assign n1399 = ( (~ N_N8199)  &  (~ N_N8198) ) | ( (~ N_N8199)  &  n2853 ) | ( (~ N_N8198)  &  n2855 ) | ( n2853  &  n2855 ) ;
 assign n1400 = ( (~ N_N8196)  &  (~ N_N8197) ) | ( (~ N_N8197)  &  n2845 ) | ( (~ N_N8196)  &  n2849 ) | ( n2845  &  n2849 ) ;
 assign n1396 = ( n1397  &  n1398  &  n1399  &  n1400 ) ;
 assign n1402 = ( (~ N_N8312)  &  (~ N_N8241) ) | ( (~ N_N8241)  &  n2849 ) | ( (~ N_N8312)  &  (~ n2857) ) | ( n2849  &  (~ n2857) ) ;
 assign n1403 = ( (~ N_N8240)  &  (~ N_N8239) ) | ( (~ N_N8239)  &  n2855 ) | ( (~ N_N8240)  &  n2858 ) | ( n2855  &  n2858 ) ;
 assign n1404 = ( (~ N_N8237)  &  (~ N_N8238) ) | ( (~ N_N8238)  &  n2851 ) | ( (~ N_N8237)  &  n2853 ) | ( n2851  &  n2853 ) ;
 assign n1405 = ( (~ N_N8236)  &  (~ N_N8235) ) | ( (~ N_N8236)  &  n2845 ) | ( (~ N_N8235)  &  n2847 ) | ( n2845  &  n2847 ) ;
 assign n1401 = ( n1402  &  n1403  &  n1404  &  n1405 ) ;
 assign n1407 = ( (~ N_N9510)  &  (~ N_N8972) ) | ( (~ N_N9510)  &  n2851 ) | ( (~ N_N8972)  &  n2855 ) | ( n2851  &  n2855 ) ;
 assign n1408 = ( (~ N_N8756)  &  (~ N_N8171) ) | ( (~ N_N8756)  &  n2845 ) | ( (~ N_N8171)  &  n2847 ) | ( n2845  &  n2847 ) ;
 assign n1409 = ( (~ N_N8037)  &  (~ N_N7854) ) | ( (~ N_N7854)  &  (~ n2857) ) | ( (~ N_N8037)  &  n2858 ) | ( (~ n2857)  &  n2858 ) ;
 assign n1410 = ( (~ N_N7852)  &  (~ N_N7853) ) | ( (~ N_N7853)  &  n2849 ) | ( (~ N_N7852)  &  n2853 ) | ( n2849  &  n2853 ) ;
 assign n1406 = ( n1407  &  n1408  &  n1409  &  n1410 ) ;
 assign n1412 = ( (~ N_N9242)  &  (~ N_N9013) ) | ( (~ N_N9013)  &  n2851 ) | ( (~ N_N9242)  &  n2853 ) | ( n2851  &  n2853 ) ;
 assign n1413 = ( (~ N_N8796)  &  (~ N_N8650) ) | ( (~ N_N8650)  &  n2849 ) | ( (~ N_N8796)  &  (~ n2857) ) | ( n2849  &  (~ n2857) ) ;
 assign n1414 = ( (~ N_N8649)  &  (~ N_N8648) ) | ( (~ N_N8648)  &  n2855 ) | ( (~ N_N8649)  &  n2858 ) | ( n2855  &  n2858 ) ;
 assign n1415 = ( (~ N_N8647)  &  (~ N_N8646) ) | ( (~ N_N8647)  &  n2845 ) | ( (~ N_N8646)  &  n2847 ) | ( n2845  &  n2847 ) ;
 assign n1411 = ( n1412  &  n1413  &  n1414  &  n1415 ) ;
 assign n1417 = ( (~ N_N9150)  &  (~ N_N8970) ) | ( (~ N_N9150)  &  n2851 ) | ( (~ N_N8970)  &  n2853 ) | ( n2851  &  n2853 ) ;
 assign n1418 = ( (~ N_N8575)  &  (~ N_N8574) ) | ( (~ N_N8575)  &  n2855 ) | ( (~ N_N8574)  &  (~ n2857) ) | ( n2855  &  (~ n2857) ) ;
 assign n1419 = ( (~ N_N8572)  &  (~ N_N8573) ) | ( (~ N_N8573)  &  n2849 ) | ( (~ N_N8572)  &  n2858 ) | ( n2849  &  n2858 ) ;
 assign n1420 = ( (~ N_N8571)  &  (~ N_N8570) ) | ( (~ N_N8571)  &  n2845 ) | ( (~ N_N8570)  &  n2847 ) | ( n2845  &  n2847 ) ;
 assign n1416 = ( n1417  &  n1418  &  n1419  &  n1420 ) ;
 assign n1422 = ( (~ N_N9275)  &  (~ N_N9244) ) | ( (~ N_N9244)  &  n2849 ) | ( (~ N_N9275)  &  n2851 ) | ( n2849  &  n2851 ) ;
 assign n1423 = ( (~ N_N8935)  &  (~ N_N8615) ) | ( (~ N_N8615)  &  n2853 ) | ( (~ N_N8935)  &  (~ n2857) ) | ( n2853  &  (~ n2857) ) ;
 assign n1424 = ( (~ N_N8531)  &  (~ N_N8530) ) | ( (~ N_N8530)  &  n2855 ) | ( (~ N_N8531)  &  n2858 ) | ( n2855  &  n2858 ) ;
 assign n1425 = ( (~ N_N8529)  &  (~ N_N8528) ) | ( (~ N_N8529)  &  n2845 ) | ( (~ N_N8528)  &  n2847 ) | ( n2845  &  n2847 ) ;
 assign n1421 = ( n1422  &  n1423  &  n1424  &  n1425 ) ;
 assign n1503 = ( N_N8869 ) | ( n1515 ) ;
 assign n1500 = ( n1503  &  (~ n1515) ) | ( n1503  &  (~ N_N8869) ) ;
 assign n1507 = ( N_N8978 ) | ( n1519 ) ;
 assign n1504 = ( n1507  &  (~ n1519) ) | ( n1507  &  (~ N_N8978) ) ;
 assign n1511 = ( N_N8933 ) | ( n1503 ) ;
 assign n1508 = ( (~ n1503)  &  n1511 ) | ( n1511  &  (~ N_N8933) ) ;
 assign n1515 = ( N_N8923 ) | ( n1522 ) ;
 assign n1512 = ( n1515  &  (~ n1522) ) | ( n1515  &  (~ N_N8923) ) ;
 assign n1519 = ( N_N8911 ) | ( n1511 ) ;
 assign n1516 = ( (~ n1511)  &  n1519 ) | ( n1519  &  (~ N_N8911) ) ;
 assign n1522 = ( (~ N_N8603) ) | ( N_N8798 ) ;
 assign n1520 = ( n1522  &  N_N8603 ) | ( n1522  &  (~ N_N8798) ) ;
 assign n1526 = ( N_N8913 ) | ( n1534 ) ;
 assign n1523 = ( n1526  &  (~ n1534) ) | ( n1526  &  (~ N_N8913) ) ;
 assign n1530 = ( N_N9031 ) | ( n1546 ) ;
 assign n1527 = ( n1530  &  (~ n1546) ) | ( n1530  &  (~ N_N9031) ) ;
 assign n1534 = ( N_N8847 ) | ( n1538 ) ;
 assign n1531 = ( n1534  &  (~ n1538) ) | ( n1534  &  (~ N_N8847) ) ;
 assign n1538 = ( N_N8631 ) | ( n1542 ) ;
 assign n1535 = ( n1538  &  (~ n1542) ) | ( n1538  &  (~ N_N8631) ) ;
 assign n1542 = ( N_N8561 ) | ( n1550 ) ;
 assign n1539 = ( n1542  &  (~ n1550) ) | ( n1542  &  (~ N_N8561) ) ;
 assign n1546 = ( N_N8993 ) | ( n1507 ) ;
 assign n1543 = ( (~ n1507)  &  n1546 ) | ( n1546  &  (~ N_N8993) ) ;
 assign n1550 = ( N_N9034 ) | ( n1530 ) ;
 assign n1547 = ( (~ n1530)  &  n1550 ) | ( n1550  &  (~ N_N9034) ) ;
 assign n1608 = ( NLC1_2 ) | ( (~ NSr1_2) ) ;
 assign n1607 = ( Preset_0_0_  &  (~ n3136) ) | ( n1608  &  (~ n3136) ) ;
 assign n1799 = ( n2851  &  n2849  &  n2858  &  n2853  &  n2847  &  n2845  &  n2977 ) ;
 assign n1800 = ( N_N8930  &  n3118 ) | ( (~ n3111)  &  n3118 ) | ( (~ n3112)  &  n3118 ) ;
 assign n1798 = ( N_N9198  &  n1799 ) | ( N_N9198  &  n1800 ) ;
 assign n1802 = ( N_N8668 ) | ( n1798 ) ;
 assign n1801 = ( n1800  &  (~ n3115) ) | ( n1802  &  (~ n3115) ) ;
 assign n1806 = ( n1371  &  (~ N_N8933) ) | ( n1801  &  (~ N_N8933) ) | ( n1371  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n1805 = ( (~ N_N9248) ) | ( N_N7306 ) | ( (~ N_N9247) ) ;
 assign n1804 = ( n1806  &  n1508 ) | ( n1806  &  n1805 ) ;
 assign n1807 = ( PRESET ) | ( (~ n3007) ) ;
 assign n1809 = ( n1361  &  (~ N_N8923) ) | ( n1801  &  (~ N_N8923) ) | ( n1361  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n1808 = ( n1809  &  n1512 ) | ( n1809  &  n1805 ) ;
 assign n1826 = ( NGFDN_3 ) | ( PRESET ) ;
 assign n1855 = ( NSr3_35 ) | ( PRESET ) ;
 assign n2066 = ( n1411  &  (~ N_N9011) ) | ( n1801  &  (~ N_N9011) ) | ( n1411  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2065 = ( (~ N_N9011)  &  n2789 ) | ( N_N9011  &  (~ n2789) ) ;
 assign n2064 = ( n2066  &  n2065 ) | ( n2066  &  n1805 ) ;
 assign n2080 = ( n1406  &  (~ N_N9031) ) | ( n1801  &  (~ N_N9031) ) | ( n1406  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2079 = ( n2080  &  n1527 ) | ( n2080  &  n1805 ) ;
 assign n2093 = ( NSr3_38 ) | ( PRESET ) ;
 assign n2099 = ( NSr3_23 ) | ( PRESET ) ;
 assign n2106 = ( n1416  &  (~ N_N8964) ) | ( n1801  &  (~ N_N8964) ) | ( n1416  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2105 = ( (~ N_N8964)  &  n1526 ) | ( N_N8964  &  (~ n1526) ) ;
 assign n2104 = ( n2106  &  n2105 ) | ( n2106  &  n1805 ) ;
 assign n2109 = ( n1391  &  (~ N_N8847) ) | ( n1801  &  (~ N_N8847) ) | ( n1391  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2108 = ( n2109  &  n1531 ) | ( n2109  &  n1805 ) ;
 assign n2143 = ( n1386  &  (~ N_N8993) ) | ( n1801  &  (~ N_N8993) ) | ( n1386  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2142 = ( n2143  &  n1543 ) | ( n2143  &  n1805 ) ;
 assign n2247 = ( NSr3_37 ) | ( PRESET ) ;
 assign n2269 = ( n1376  &  (~ N_N8978) ) | ( n1801  &  (~ N_N8978) ) | ( n1376  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2268 = ( n2269  &  n1504 ) | ( n2269  &  n1805 ) ;
 assign n2283 = ( n1351  &  (~ N_N8869) ) | ( n1801  &  (~ N_N8869) ) | ( n1351  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2282 = ( n2283  &  n1500 ) | ( n2283  &  n1805 ) ;
 assign n2285 = ( n1356  &  (~ N_N8798) ) | ( n1801  &  (~ N_N8798) ) | ( n1356  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2284 = ( n2285  &  n1520 ) | ( n2285  &  n1805 ) ;
 assign n2364 = ( n1381  &  (~ N_N9034) ) | ( n1801  &  (~ N_N9034) ) | ( n1381  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2363 = ( n2364  &  n1547 ) | ( n2364  &  n1805 ) ;
 assign n2366 = ( n1346  &  (~ N_N8911) ) | ( n1801  &  (~ N_N8911) ) | ( n1346  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2365 = ( n2366  &  n1516 ) | ( n2366  &  n1805 ) ;
 assign n2373 = ( NSr3_30 ) | ( PRESET ) ;
 assign n2419 = ( NSr3_20 ) | ( PRESET ) ;
 assign n2434 = ( n1396  &  (~ N_N8561) ) | ( n1801  &  (~ N_N8561) ) | ( n1396  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2433 = ( n2434  &  n1539 ) | ( n2434  &  n1805 ) ;
 assign n2649 = ( n1421  &  (~ N_N8913) ) | ( n1801  &  (~ N_N8913) ) | ( n1421  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2648 = ( n2649  &  n1523 ) | ( n2649  &  n1805 ) ;
 assign n2651 = ( n1401  &  (~ N_N8631) ) | ( n1801  &  (~ N_N8631) ) | ( n1401  &  n3008 ) | ( n1801  &  n3008 ) ;
 assign n2650 = ( n2651  &  n1535 ) | ( n2651  &  n1805 ) ;
 assign n2693 = ( NSr3_14 ) | ( PRESET ) ;
 assign n2782 = ( Preset_0_0_  &  (~ n1608) ) ;
 assign N_N7729 = ( n196  &  (~ NSr1_2) ) ;
 assign n2787 = ( (~ PRESET)  &  (~ PDN)  &  Pover_0_0_ ) | ( (~ PRESET)  &  Pover_0_0_  &  NDN1_4 ) ;
 assign N_N7199 = ( N_N7729 ) | ( n2787 ) ;
 assign n2789 = ( N_N8964 ) | ( n1526 ) ;
 assign n2819 = ( (~ NGFDN_3)  &  NDN3_46 ) ;
 assign N_N7098 = ( (~ PRESET)  &  n2819 ) ;
 assign n2838 = ( NDN2_2 ) | ( (~ n2782) ) ;
 assign n2845 = ( (~ NEN3_36) ) | ( (~ NSr3_38) ) ;
 assign n2847 = ( (~ NEN3_34) ) | ( (~ NSr3_37) ) ;
 assign n2849 = ( (~ NDN3_29) ) | ( (~ NSr3_35) ) ;
 assign n2851 = ( (~ NDN3_26) ) | ( (~ NSr3_30) ) ;
 assign n2853 = ( (~ NDN3_19) ) | ( (~ NSr3_23) ) ;
 assign n2855 = ( NSr3_13 ) | ( (~ NSr3_14) ) ;
 assign n2857 = ( NSr3_13  &  NDN3_12 ) ;
 assign n2858 = ( (~ NDN3_17) ) | ( (~ NSr3_20) ) ;
 assign n2977 = ( n2855  &  (~ n2857) ) ;
 assign n2979 = ( n1805  &  (~ n3115) ) ;
 assign n3007 = ( n1802  &  n2979 ) ;
 assign n3008 = ( (~ n1800) ) | ( n1802 ) ;
 assign n3010 = ( (~ N_N8603)  &  n1520  &  (~ n1805) ) ;
 assign n3011 = ( n1531  &  n1527  &  n1539  &  n1535  &  n1547  &  n1543  &  n1523  &  n2065 ) ;
 assign n3111 = ( n1346  &  n1406  &  n1356  &  n1351  &  n1366  &  n1361  &  n1376  &  n1371 ) ;
 assign n3112 = ( n1416  &  n1411  &  n1381  &  n1421  &  n1391  &  n1386  &  n1401  &  n1396 ) ;
 assign n3115 = ( n227  &  (~ N_N9247) ) ;
 assign n3118 = ( N_N8929 ) | ( (~ N_N8930) ) ;
 assign n3132 = ( N_N8603  &  n1805 ) | ( (~ N_N8603)  &  n3008 ) | ( n1805  &  n3008 ) ;
 assign n3133 = ( n1366  &  (~ n3007)  &  n3132 ) | ( n1801  &  (~ n3007)  &  n3132 ) ;
 assign n3136 = ( NSr1_2  &  N_N7476  &  NLC1_2 ) ;


endmodule

