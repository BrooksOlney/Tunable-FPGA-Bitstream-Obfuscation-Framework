module ex1010x5_map (i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_, o_1_, o_2_, o_0_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

	input i_9_;
	input i_7_;
	input i_8_;
	input i_5_;
	input i_6_;
	input i_3_;
	input i_4_;
	input i_1_;
	input i_2_;
	input i_0_;
	output o_1_;
	output o_2_;
	output o_0_;
	output o_9_;
	output o_7_;
	output o_8_;
	output o_5_;
	output o_6_;
	output o_3_;
	output o_4_;



	wire x12042x, x12038x, n_n1007, n_n1009, x12041x, x12589x, x12151x, x12152x, n_n1398, n_n1392, x13147x, x13136x, x13137x, x13684x, x13573x, x13574x, x14222x, x14216x, n_n3251, n_n3253, x14780x;
	wire n_n3623, n_n3624, x14775x, x14778x, x15301x, n_n2523, x15300x, x15817x, n_n2898, x15816x, x16324x, n_n1706, x15943x, n_n1784, x16320x, x16831x, x16832x, n_n1014, n_n1013, x11894x, n_n1010;
	wire n_n1012, n_n1020, n_n1052, n_n1054, x11977x, x12036x, n_n1017, n_n1045, x11953x, x11960x, x11961x, n_n1023, n_n1061, n_n1062, x12020x, x12028x, n_n1015, x11747x, n_n942, n_n941, n_n1396;
	wire n_n1397, x12391x, n_n1394, n_n1393, x12062x, x12063x, x12083x, x12084x, n_n1323, x12129x, x12130x, x12150x, x12440x, n_n1480, n_n1418, x12431x, n_n1481, x12585x, n_n1425, n_n1423, x12517x;
	wire n_n1399, x12693x, n_n539, n_n540, x13146x, n_n630, n_n657, n_n656, x13088x, n_n629, n_n627, n_n628, x12867x, x13001x, x13002x, x13645x, x13646x, n_n3921, x13683x, n_n3990, n_n3992;
	wire n_n3988, n_n3987, n_n3989, n_n3993, n_n3995, x13555x, x13569x, n_n3192, x13782x, x13783x, x14221x, n_n3257, n_n3259, x14214x, n_n3254, n_n3256, x14067x, n_n3260, n_n3262, x14211x, x14540x;
	wire n_n3625, n_n3627, n_n3629, n_n3631, x14591x, n_n3661, n_n3660, x14566x, n_n3634, x14638x, x14613x, n_n3635, n_n3676, x14612x, x14388x, n_n659, n_n3649, x22190x, n_n3543, x14343x, n_n3626;
	wire n_n2530, n_n2529, x15169x, n_n2533, n_n2532, x15297x, n_n2526, n_n2542, n_n2541, x15264x, n_n2449, n_n2531, x14890x, x14891x, n_n2906, n_n2908, n_n2902, x15677x, n_n2921, n_n2903, n_n2905;
	wire n_n2922, x15806x, n_n2827, n_n2821, n_n2826, n_n2907, x15811x, n_n1793, n_n1792, n_n1794, n_n1787, n_n1709, x15899x, x15900x, x15901x, n_n1712, n_n1711, x15939x, x15940x, x16242x, n_n1789;
	wire n_n1790, x15991x, x16318x, x16319x, n_n1801, n_n1800, x16470x, n_n2165, n_n2164, n_n2162, n_n2163, n_n2166, n_n2160, x16764x, x16826x, x16827x, x11530x, n_n1107, x11501x, n_n1038, x11500x;
	wire x11581x, n_n1034, n_n1035, n_n1083, n_n1082, x11766x, n_n1028, x11892x, n_n1026, n_n1071, n_n1072, x11815x, x11832x, n_n1088, x11851x, n_n1032, x11884x, x11850x, x12199x, n_n1412, n_n1413;
	wire x12247x, n_n1466, x12223x, n_n1415, x12222x, n_n1450, n_n1451, x12324x, n_n1408, x12389x, n_n1442, n_n1405, x12296x, x12305x, x12295x, n_n1404, x12381x, x12380x, n_n553, x12683x, x12684x;
	wire x12689x, x12690x, n_n546, x12640x, x12641x, x12647x, x12648x, x12656x, x12657x, n_n551, x12670x, x12671x, n_n543, n_n542, x13142x, x13143x, n_n4748, n_n4725, n_n4788, n_n4802, x13644x;
	wire x13630x, x13631x, x13636x, x13637x, x13650x, x13651x, n_n3932, x13663x, x13664x, x13616x, n_n3926, n_n3924, x13615x, x13681x, x13761x, x13747x, x13748x, x13753x, x13754x, n_n4853, n_n4847;
	wire n_n4864, n_n4912, x13781x, x13767x, x13768x, x13773x, x13774x, n_n3189, n_n3205, x13728x, x13729x, x14218x, n_n3653, x14530x, n_n3729, n_n3731, x14538x, n_n3638, n_n3639, n_n3685, n_n3686;
	wire x14682x, x14730x, n_n3645, n_n3702, x14722x, x14721x, n_n3650, n_n3652, x14436x, x14513x, n_n3658, x14507x, n_n3732, n_n3734, n_n2548, n_n2598, n_n2597, n_n2549, x14933x, n_n2589, n_n2588;
	wire n_n2546, n_n2545, x14979x, n_n2560, n_n2559, x15167x, n_n2558, n_n2557, x15103x, n_n2554, n_n2553, x15150x, x15503x, n_n2990, n_n2991, n_n2926, x15494x, x15549x, n_n2934, n_n3004, n_n3005;
	wire x15543x, n_n2915, n_n2952, x15633x, x15642x, x15632x, n_n2912, n_n2911, x15594x, x15674x, x15675x, x16027x, n_n1882, n_n1817, x16018x, x16017x, x16072x, n_n1877, x16048x, n_n1812, n_n1876;
	wire x16114x, n_n1896, x16086x, n_n1818, x16085x, x16289x, n_n1832, x16262x, n_n1797, x16261x, n_n2175, x16456x, n_n2223, n_n2225, x16468x, x16598x, n_n2189, x16590x, n_n2253, x16589x, x16645x;
	wire n_n2185, n_n2184, n_n2178, x16365x, x16376x, x16362x, x16363x, n_n2236, n_n2237, n_n2182, n_n2183, x16423x, x16557x, n_n2190, n_n2268, x16545x, x16544x, x467x, n_n2173, n_n2172, n_n2214;
	wire x16742x, n_n2170, n_n2169, x16705x, n_n2168, x16762x, n_n2087, x16516x, x16517x, n_n2103, n_n2084, x16821x, x16822x, x16824x, n_n4440, n_n4434, n_n4442, n_n4443, x22164x, n_n1113, n_n4448;
	wire n_n4450, x368x, n_n3889, x32x, n_n1112, x37x, x84x, n_n4428, x79x, x11524x, x11528x, x13x, x572x, x129x, x308x, x22163x, x130x, n_n4524, x170x, n_n4492, x22162x;
	wire n_n1111, x206x, x11516x, x11517x, n_n4498, n_n4499, x307x, x162x, x347x, n_n455, n_n473, n_n532, n_n534, n_n4243, n_n4542, x201x, n_n4549, n_n4551, x22161x, n_n1104, n_n4557;
	wire n_n4561, x213x, x11542x, n_n1103, n_n482, n_n520, x20x, n_n3875, n_n526, n_n530, x11577x, n_n1099, x11555x, x11556x, x11557x, n_n1100, x224x, x11572x, x11573x, n_n4317, n_n4318;
	wire n_n4320, n_n4316, x11587x, n_n1123, n_n1117, n_n1115, x11604x, n_n1040, x300x, n_n1120, n_n3176, x11618x, x161x, n_n1041, n_n4337, n_n4344, n_n4335, x11620x, x22150x, n_n1121, n_n4327;
	wire n_n4331, x410x, x11631x, x11632x, x11719x, x11720x, x11726x, x11727x, x11736x, x11698x, x11699x, x11732x, x22198x, x11734x, x11705x, x11706x, n_n947, x11735x, x11660x, x11661x, x11667x;
	wire x11668x, x11743x, x11745x, n_n4800, x11757x, n_n4798, x439x, x24x, x530x, n_n4812, x11762x, x151x, n_n4787, x313x, n_n4792, n_n2003, x292x, n_n3460, x177x, n_n4838, x11782x;
	wire x11778x, n_n1086, n_n1087, x315x, x191x, x11889x, n_n1057, x11908x, x11907x, n_n5223, n_n5221, n_n5215, x181x, x22157x, n_n5200, n_n5188, n_n1927, x188x, x452x, n_n5207, n_n5203;
	wire x36x, x11976x, n_n1059, n_n1060, x211x, x422x, x12033x, n_n4506, n_n4546, n_n4555, n_n4562, x12061x, x12048x, x12049x, x12053x, x12054x, n_n4774, n_n4845, n_n4796, n_n4822, x12082x;
	wire x12068x, x12069x, x12074x, x12075x, n_n1330, n_n1331, x12110x, x12089x, x12090x, x12128x, x12117x, x12118x, n_n1333, n_n1341, x12141x, x12142x, x12146x, x12147x, n_n524, n_n518, n_n195;
	wire n_n4979, n_n4978, n_n4982, n_n4988, n_n4989, n_n4985, n_n4986, x12156x, n_n4991, n_n5000, n_n1576, x247x, x104x, n_n1455, n_n4983, n_n4984, x228x, x362x, x12196x, x22195x, x12164x;
	wire x12165x, x142x, x12176x, n_n3810, n_n1592, n_n1463, x12188x, x12190x, n_n325, n_n528, x402x, n_n4793, x179x, n_n4799, x22147x, n_n1471, n_n4779, n_n4780, n_n4783, n_n4778, n_n4775;
	wire x12209x, n_n4805, x71x, n_n4197, x440x, x12245x, n_n4865, x245x, n_n4852, x22146x, n_n4870, n_n4877, n_n1985, n_n3815, x12217x, n_n1468, x12235x, x12236x, x12240x, n_n4868, n_n4880;
	wire x330x, x263x, x324x, n_n5060, n_n5055, n_n5059, n_n5056, x12311x, n_n5054, n_n5042, x97x, x12316x, n_n5075, n_n5068, x12321x, x12322x, n_n1446, x12333x, x12334x, x12338x, x12339x;
	wire n_n1453, n_n1454, x12385x, x12386x, n_n4762, n_n4765, n_n4766, n_n4205, x12394x, n_n1473, x483x, n_n4740, n_n3475, x22143x, n_n1475, n_n4754, n_n4757, n_n4749, n_n4760, x12436x, n_n4747;
	wire n_n4755, n_n4761, n_n4752, x12437x, n_n4674, n_n4671, n_n1636, x417x, x12418x, x12416x, x12404x, x12405x, n_n1476, x10x, n_n464, n_n4689, x22206x, n_n4667, n_n4662, n_n4660, x72x;
	wire x12425x, n_n3903, n_n1504, n_n1693, x12452x, x12454x, n_n1427, x83x, x12460x, x12469x, x12468x, n_n1426, n_n4341, x67x, x53x, x448x, n_n1506, x283x, x364x, x12575x, n_n1508;
	wire n_n4332, n_n4328, x106x, n_n1703, x12581x, x12476x, x12485x, x12481x, x22141x, n_n1491, x12504x, x12505x, x12506x, n_n1496, x12513x, x12514x, x22140x, n_n1422, n_n1485, n_n1487, n_n1420;
	wire x12565x, x25x, n_n65, n_n5305, x15x, x592x, n_n5293, x19x, n_n5296, n_n491, x492x, n_n5284, n_n4578, n_n4611, n_n4633, n_n4581, x12597x, n_n559, n_n4641, n_n4643, n_n4646;
	wire n_n4647, x12600x, n_n4648, n_n4645, n_n4635, x140x, x12601x, n_n4572, n_n4531, x12607x, n_n4523, n_n4539, n_n4559, n_n4528, x12608x, n_n4718, x23x, n_n4727, n_n509, n_n4730, n_n4733;
	wire n_n4735, n_n4750, n_n4736, x12628x, x12629x, x165x, n_n522, n_n500, x258x, x131x, n_n4764, n_n4763, x12614x, n_n4656, n_n4676, n_n4703, n_n4698, x12621x, n_n557, n_n4885, n_n4911;
	wire n_n4903, n_n4895, x12679x, n_n260, n_n535, x38x, x11x, n_n4819, x395x, n_n4928, n_n4950, n_n4956, n_n4936, n_n4918, n_n4917, n_n4931, n_n4948, n_n4954, x496x, n_n4441, n_n536;
	wire n_n4404, n_n4384, x12700x, n_n4379, n_n4371, n_n4399, n_n4417, x12701x, n_n4460, n_n4473, x12707x, n_n4512, n_n4453, n_n4471, n_n4488, n_n4458, x12708x, n_n4363, n_n4347, n_n4315, x12714x;
	wire n_n4338, n_n4326, n_n4350, x12715x, n_n727, x13016x, n_n653, x13046x, x13015x, x74x, x398x, x13060x, x13065x, x13064x, n_n730, x13074x, x13075x, x13080x, x337x, x124x, n_n738;
	wire n_n737, x13085x, n_n719, n_n651, n_n650, x13130x, x13131x, n_n698, x12752x, n_n646, x12775x, x12751x, n_n648, n_n649, x12827x, n_n642, n_n641, x12865x, n_n634, x12984x, x12999x;
	wire n_n635, n_n637, n_n639, n_n638, x12947x, n_n5297, n_n4007, x13235x, x13234x, n_n4072, n_n4013, n_n4014, x13276x, x13303x, n_n4002, x13326x, n_n4036, n_n4037, n_n3998, n_n3999, x13374x;
	wire n_n4051, n_n4050, n_n4003, n_n4004, x13421x, x13482x, n_n4016, n_n4015, n_n4023, n_n4100, n_n4102, n_n4021, x13545x, n_n4020, x13501x, n_n4090, x13500x, x13553x, n_n4010, n_n4009, x13188x;
	wire n_n3996, n_n5017, n_n5015, n_n5037, x13606x, n_n5032, n_n5036, n_n5021, n_n5020, n_n5047, x13607x, n_n5156, n_n5191, n_n5175, n_n5177, x13611x, n_n5171, n_n5190, n_n5170, n_n5194, n_n5213;
	wire x13612x, n_n4392, n_n4391, x13623x, n_n4378, n_n4388, n_n4407, n_n4402, n_n4408, x13624x, n_n4781, n_n4742, n_n4808, n_n4663, n_n4665, n_n4672, n_n4707, n_n4724, n_n4679, n_n4701, n_n4692;
	wire n_n4686, n_n4913, n_n4905, n_n4846, n_n4901, n_n4904, n_n4842, n_n4841, n_n4867, n_n4570, x523x, x214x, n_n4576, n_n4552, n_n4580, n_n4617, n_n4637, n_n4613, n_n4602, x13657x, n_n4504;
	wire n_n4535, n_n4507, n_n4509, n_n4521, n_n4544, n_n4540, n_n4520, n_n4470, n_n4413, n_n4457, x13672x, n_n4459, n_n4420, n_n4472, n_n4480, n_n4410, x13673x, n_n4340, n_n4368, n_n4358, n_n4354;
	wire x13679x, n_n4325, n_n4362, n_n4312, n_n3937, n_n4339, n_n4401, n_n4314, n_n4389, x13689x, n_n4369, n_n4381, x13690x, n_n5182, n_n5173, n_n5165, n_n5230, x13703x, n_n5239, n_n5238, n_n5166;
	wire n_n5163, n_n5214, x13704x, n_n5274, n_n5300, n_n5254, n_n5287, x13710x, n_n5240, n_n5281, n_n5268, n_n5261, x13711x, n_n5302, x13713x, n_n4487, n_n4409, x13735x, n_n4456, n_n4484, n_n4462;
	wire x13736x, n_n4533, x13741x, n_n4532, n_n4545, x471x, n_n390, n_n4638, n_n4640, n_n4683, n_n4685, n_n3125, x13760x, n_n4786, n_n4767, n_n4723, n_n4571, n_n4594, n_n4629, n_n4583, n_n4630;
	wire n_n4900, n_n4849, n_n4908, n_n4891, n_n4896, n_n4977, n_n4920, n_n4922, n_n4959, n_n4980, n_n4953, x351x, n_n4972, n_n4816, n_n4828, x552x, n_n4844, n_n4818, n_n3272, n_n3274, n_n3322;
	wire x13875x, x13876x, n_n3336, n_n3280, n_n3279, x13916x, x13917x, n_n5331, n_n3277, n_n3275, x13827x, x14240x, x14226x, x14227x, x14232x, x14233x, n_n3546, n_n5307, n_n5266, x14256x, x14246x;
	wire x63x, n_n3545, n_n5057, n_n4994, n_n4974, x275x, x14273x, x14275x, x14261x, x14262x, x14267x, x14268x, x14276x, n_n3562, x14301x, x14302x, x14308x, x14309x, n_n3549, n_n4759, n_n4811;
	wire x14331x, x14332x, x14317x, x14318x, x14323x, x14324x, x14333x, n_n3565, x14290x, x14291x, x14339x, x14341x, x350x, n_n4758, x370x, x14376x, x95x, n_n4728, x22104x, n_n3707, x109x;
	wire n_n4743, n_n4745, n_n4210, x14382x, x14386x, x14448x, x14449x, x14455x, x14456x, x14457x, n_n4444, n_n4445, x22165x, x321x, x98x, n_n4426, n_n2802, x215x, x194x, n_n3727, n_n3726;
	wire x322x, x14535x, n_n5278, n_n5275, n_n5279, n_n5280, x22186x, n_n3664, n_n5267, n_n5262, x409x, x205x, x14548x, n_n3665, n_n5289, n_n5285, n_n5282, x14542x, x22107x, x14589x, n_n5312;
	wire n_n5313, x325x, n_n5315, x22106x, n_n5318, n_n5326, n_n5329, n_n5327, x14561x, n_n5292, x197x, x200x, x60x, x14562x, x14572x, x14573x, x14579x, x14580x, x14581x, x76x, x126x;
	wire n_n5144, n_n5143, n_n777, n_n3674, n_n5155, n_n5154, x195x, x14598x, n_n3673, x33x, x14635x, x14636x, n_n5113, n_n5114, n_n3412, n_n3771, n_n3772, n_n3670, x14629x, x14625x, n_n5121;
	wire n_n5119, x14604x, x22105x, n_n5111, n_n5112, n_n5107, n_n5108, n_n3051, x14644x, x14645x, x14648x, x14649x, x14654x, x14659x, x14660x, x14665x, x14666x, x136x, n_n5003, n_n5002, x299x;
	wire x14670x, n_n4995, n_n4999, x41x, n_n5018, n_n5014, x14681x, x40x, x295x, n_n4871, x14687x, n_n3696, x375x, x22111x, n_n3698, n_n4857, n_n4856, n_n4854, n_n4855, x14727x, x14728x;
	wire n_n3701, x14708x, x14709x, x22110x, x380x, x381x, x14712x, n_n4204, n_n4782, n_n4790, x14718x, n_n4890, x264x, x261x, n_n3694, n_n4899, x14739x, n_n3693, n_n3691, x14748x, x14749x;
	wire n_n3642, n_n3803, n_n3802, x14754x, x14764x, x14763x, n_n3641, n_n4882, n_n4881, n_n4878, x14769x, x14770x, n_n5330, x371x, x14793x, x14796x, x155x, x143x, x14785x, x14790x, x14791x;
	wire x14797x, x14807x, x14803x, x14804x, x14825x, x14826x, x14829x, x14813x, x14814x, x14820x, x14821x, x14828x, n_n1217, n_n4848, x14907x, x14904x, n_n3451, x174x, n_n4876, n_n4874, x14908x;
	wire n_n3450, n_n4894, n_n4889, x12179x, x49x, x14927x, x14918x, x14919x, x14926x, n_n4862, n_n4872, x14932x, n_n4987, n_n4993, x134x, x252x, x393x, x14940x, x14960x, x14948x, x14949x;
	wire n_n2596, n_n4939, x382x, x14974x, n_n2591, x14970x, x29x, n_n4965, x68x, x21x, x47x, x14986x, n_n2608, x164x, x22092x, n_n2607, n_n4776, n_n4777, x15021x, n_n4773, x15022x;
	wire x15025x, n_n2614, x15002x, x15003x, x15004x, n_n2552, n_n2611, x15013x, x15014x, x15015x, n_n2551, n_n2637, x15033x, x15034x, x15040x, n_n2634, x15049x, x15050x, x15055x, x156x, n_n2640;
	wire n_n2641, x15164x, n_n2570, x15221x, x15220x, n_n2538, x15269x, x15270x, x15278x, x15277x, n_n2539, n_n5167, n_n5164, n_n5162, x15284x, n_n2576, n_n5149, n_n5152, n_n5153, x407x, x22204x;
	wire n_n2577, n_n5138, n_n2304, x22184x, x15293x, n_n2568, n_n2569, x15184x, x15206x, x15205x, x90x, n_n2584, x15232x, x22093x, x15239x, x15240x, x15249x, x15248x, x15254x, x15255x, n_n2586;
	wire x15262x, n_n4359, n_n4397, x15308x, n_n4431, n_n4436, n_n4424, x15309x, n_n4451, n_n4476, x15316x, n_n4478, n_n2844, n_n4345, n_n4319, n_n4355, x15323x, n_n4357, n_n4348, n_n2846, n_n4514;
	wire n_n4511, n_n4525, n_n4543, n_n4527, n_n4534, x15341x, x15342x, n_n4598, n_n4612, x15329x, n_n2842, n_n4659, x75x, x15334x, n_n4634, n_n4631, n_n4691, n_n4687, x15335x, n_n5090, n_n5080;
	wire x279x, x15367x, x15369x, x15355x, x15356x, x15361x, x15362x, x15370x, x15374x, x15375x, x15381x, x15382x, x15383x, n_n2823, n_n4957, x141x, x15396x, x15398x, x15348x, x15349x, n_n2835;
	wire x15399x, x73x, n_n4700, x14x, n_n1760, n_n4711, x15414x, x15418x, n_n4769, n_n4794, n_n4797, x15406x, n_n4815, x15407x, n_n4817, n_n4843, n_n4823, x15413x, n_n2838, n_n4466, x412x;
	wire n_n4469, x22082x, n_n3001, x323x, n_n4449, x470x, x421x, n_n3003, n_n4463, n_n4455, n_n4452, x15459x, n_n4461, n_n4454, n_n4465, x15460x, x15463x, n_n4496, x163x, x22081x, n_n2999;
	wire n_n4489, x70x, n_n3515, n_n4486, x189x, n_n4490, n_n3509, x15433x, x15437x, n_n2997, x15445x, x15446x, x15453x, n_n2929, x100x, x237x, n_n4574, n_n4573, n_n3870, x276x, x222x;
	wire n_n2993, n_n4587, x365x, n_n4585, x15479x, n_n4554, x22090x, x15501x, n_n4618, n_n4232, n_n4620, x22226x, n_n4593, n_n4601, n_n4590, x15489x, n_n2987, x15471x, x15470x, n_n4628, x190x;
	wire x15493x, n_n4383, n_n4385, n_n4390, x15508x, n_n3007, n_n4366, x64x, x15512x, n_n4365, n_n4356, n_n4353, x15513x, n_n4373, n_n4374, x27x, x15547x, n_n3010, n_n3012, x15527x, n_n4433;
	wire n_n4438, x15531x, x22200x, n_n4416, n_n4414, x15536x, n_n4403, x15542x, x15607x, x15611x, x15618x, x22087x, n_n5106, x127x, x22086x, n_n5134, x15626x, n_n2957, x15602x, x15603x, x15638x;
	wire x15639x, n_n5136, n_n5124, x335x, x35x, x286x, x15554x, x15555x, x15564x, x15563x, n_n3031, n_n2943, n_n3385, x15575x, x15577x, n_n5179, n_n2948, n_n2949, x22180x, n_n5288, n_n5286;
	wire n_n2937, x15668x, x15649x, x15650x, n_n2939, n_n2940, x15671x, n_n3820, n_n2973, x15693x, x15695x, n_n2966, n_n2917, n_n2918, n_n2965, x15740x, n_n2977, n_n2979, x15766x, n_n2925, x15786x;
	wire x158x, x15791x, x15798x, x15797x, n_n2970, n_n2968, x15802x, x15803x, x15887x, x15871x, x15872x, n_n1717, x15845x, x15846x, x15898x, x15852x, x15853x, x15859x, x15860x, n_n1720, x15894x;
	wire x15895x, x15838x, x15823x, x15824x, x15829x, x15830x, x15932x, x15920x, x15921x, x15924x, x15925x, x15938x, x15909x, x15910x, x15915x, x15916x, x18x, x15978x, n_n5048, n_n5044, n_n5045;
	wire n_n5053, x15979x, n_n5025, n_n5023, n_n5024, x15983x, n_n1844, n_n5027, n_n5028, x50x, n_n5029, x22069x, x15989x, n_n3883, x65x, n_n1885, x78x, n_n4477, x184x, n_n4479, x376x;
	wire n_n1886, n_n4503, x16023x, n_n4500, x16024x, n_n4537, x11532x, n_n4529, x22223x, x16007x, n_n1889, n_n4526, n_n3504, x14108x, x14109x, n_n4517, n_n4584, n_n2401, n_n1878, x121x, x16036x;
	wire n_n4560, x430x, n_n4239, x16070x, n_n4575, n_n4577, x22201x, n_n4595, x172x, n_n4588, x45x, n_n2037, n_n4621, x16047x, x16065x, x16053x, x16054x, n_n1873, n_n4609, n_n4608, x51x;
	wire n_n2036, n_n4275, x16089x, n_n1894, n_n4380, x280x, x14460x, n_n4377, n_n1893, n_n4361, x16110x, x16111x, x22078x, n_n4279, x16080x, n_n1890, x16099x, x16100x, x16105x, n_n4321, x443x;
	wire n_n4744, x374x, x22073x, n_n1867, n_n4751, x22072x, n_n1866, n_n4722, x242x, x22177x, x16130x, x16135x, x16144x, x16141x, x22071x, n_n1811, n_n1863, x16233x, x16234x, x16238x, x16240x;
	wire n_n1846, x16157x, n_n1805, x16180x, x16156x, n_n1854, n_n1808, n_n1807, n_n1856, x16222x, n_n5157, n_n5160, x466x, n_n130, x16245x, n_n5174, x254x, x16248x, n_n1833, n_n5142, n_n5148;
	wire x196x, x22077x, x16287x, n_n5186, n_n5187, x152x, x22076x, n_n5212, n_n5189, x453x, x22218x, x16267x, x16268x, n_n1829, x16278x, x16279x, x220x, x454x, n_n5192, n_n5308, n_n5319;
	wire n_n5332, x117x, x16315x, n_n5310, n_n5311, n_n5309, n_n5304, x22068x, x218x, x22067x, n_n1825, n_n5298, x16301x, n_n1824, n_n5264, x77x, x334x, x203x, x16302x, n_n1826, x516x;
	wire x506x, n_n5320, n_n1900, x16314x, n_n2218, x16435x, x16436x, x16440x, x16441x, n_n4915, x22064x, x31x, n_n4937, n_n4933, n_n4935, x249x, x226x, x16447x, n_n3805, x16327x, n_n2220;
	wire x16466x, n_n4400, x16476x, n_n4405, n_n4406, x16477x, n_n4513, x16483x, n_n4518, n_n2102, x16487x, x256x, n_n4623, x16488x, n_n4547, x16494x, n_n4553, x16495x, n_n2130, n_n4803, x16514x;
	wire n_n4710, n_n4719, n_n4708, x16503x, n_n4772, n_n4706, n_n4699, x16504x, n_n4675, x16509x, n_n4661, x16510x, x345x, n_n2267, n_n4382, x423x, x16554x, n_n4386, n_n2435, x282x, x12447x;
	wire x16555x, n_n2263, x16526x, x16527x, x16533x, n_n4343, n_n4352, x399x, x22197x, n_n2446, n_n2443, n_n2445, n_n4336, x198x, n_n4491, n_n4497, x66x, n_n2257, n_n4254, n_n2258, n_n4505;
	wire x16595x, x16596x, n_n2261, x16568x, x16569x, n_n4247, n_n4510, x22063x, x22208x, x178x, x378x, n_n4568, x455x, n_n2251, x16606x, n_n4548, x16642x, x238x, x22062x, x16622x, x16611x;
	wire x16612x, x16617x, x16618x, x16628x, n_n2246, x16636x, x22061x, x16651x, n_n4367, x16652x, n_n5031, x13400x, x111x, x253x, x16715x, x16711x, x16713x, n_n2210, n_n2209, x16728x, x16729x;
	wire n_n5052, x22221x, n_n5040, x16741x, x16682x, n_n2204, x16681x, n_n5251, x435x, n_n1139, x16697x, x16693x, x358x, x16666x, n_n2205, x125x, x16703x, x16758x, n_n2196, x16757x, x462x;
	wire x16659x, x16660x, x16761x, n_n4432, n_n4421, x16769x, n_n4429, n_n5034, n_n5099, n_n5019, n_n5097, x16790x, n_n5104, n_n5117, n_n5122, x16791x, n_n5123, n_n5131, n_n5137, n_n5146, x16796x;
	wire n_n5193, n_n5168, x16797x, n_n4996, n_n4992, n_n4981, n_n5005, x16804x, x16805x, n_n4464, n_n4467, n_n4666, n_n4664, n_n4737, n_n4738, n_n4784, x17x, n_n4830, n_n4831, n_n4902, n_n4898;
	wire n_n4976, n_n4975, n_n5038, x12x, n_n5092, n_n5093, n_n5091, n_n4148, x233x, x236x, x13428x, n_n4095, n_n4720, n_n4717, x241x, n_n4863, x102x, n_n4859, n_n4858, x13171x, n_n4990;
	wire n_n4998, n_n5001, x103x, x13381x, n_n4927, n_n4958, n_n4324, n_n4923, n_n4924, n_n4921, n_n5035, n_n5109, x583x, n_n4597, n_n4605, x108x, n_n4596, x257x, x22114x, n_n3347, n_n4756;
	wire x22117x, n_n4887, n_n4888, n_n4883, x262x, n_n5026, n_n3424, n_n5178, n_n3399, n_n5181, n_n5184, n_n5185, n_n5183, x112x, x14026x, n_n3303, n_n5316, x502x, n_n5321, x268x, x459x;
	wire x13935x, n_n3292, n_n4615, n_n4616, n_n4607, n_n4606, x14072x, x14073x, n_n4625, n_n1649, x26x, n_n4619, x118x, x309x, n_n4639, n_n4642, x348x, n_n4632, x349x, x14080x, x14082x;
	wire x14081x, n_n3281, n_n5050, n_n5064, x120x, n_n5058, x13982x, x13983x, x13984x, x231x, n_n5046, x356x, x13991x, x13990x, x22222x, n_n3270, n_n5096, n_n5085, n_n5101, n_n5110, n_n5130;
	wire n_n5129, n_n5145, x13696x, x13697x, n_n4515, n_n4791, n_n4860, n_n4926, n_n4925, n_n5041, n_n5100, n_n4734, n_n4726, x101x, x244x, x15745x, n_n2981, n_n4861, x246x, n_n4869, x294x;
	wire x15678x, n_n5022, x296x, x298x, x15705x, n_n5004, n_n5006, n_n5007, n_n4907, n_n5132, n_n5088, n_n5081, n_n5098, n_n5095, n_n5172, n_n5234, x385x, n_n4934, n_n5324, n_n5335, x531x;
	wire n_n5010, n_n4967, n_n4962, n_n4897, n_n4886, n_n4929, x353x, n_n5245, n_n5235, n_n5248, x14834x, n_n4494, x14839x, n_n4475, x14840x, x14849x, n_n4770, n_n4771, n_n4826, x14869x, x14870x;
	wire n_n4697, n_n4681, x14855x, n_n4673, n_n4690, x14856x, x14861x, n_n4714, x14862x, x14871x, x14876x, n_n4396, n_n4375, x14877x, x14882x, n_n4330, n_n4351, n_n4313, x14883x, x234x, n_n4447;
	wire n_n4415, n_n4372, n_n4430, n_n4495, n_n4834, n_n4835, n_n4832, n_n4909, n_n5049, n_n4644, n_n4651, n_n4649, n_n4652, x311x, n_n4952, n_n4942, n_n4945, n_n4946, n_n4949, n_n5244, n_n5241;
	wire n_n5242, n_n5247, n_n5246, x319x, x16687x, x16563x, x147x, n_n4468, x260x, x16330x, n_n2226, n_n4850, x277x, x16336x, n_n2228, n_n4875, n_n4873, x16340x, x16341x, n_n5322, n_n2274;
	wire n_n5325, x115x, x16292x, n_n5303, n_n5306, n_n4804, n_n4795, x16349x, n_n4801, x16350x, n_n4840, x185x, x388x, n_n2230, n_n4837, x16357x, n_n3469, n_n2234, n_n4789, x22060x, x16374x;
	wire n_n4824, n_n4806, n_n4821, n_n4820, n_n4810, x16383x, n_n4753, x293x, n_n4702, n_n2378, n_n4709, x22219x, x16399x, n_n4696, n_n4695, n_n4712, x16395x, x39x, n_n4715, x16390x, x22176x;
	wire n_n1764, n_n4688, n_n3849, n_n3848, x16415x, x16406x, n_n2242, n_n4657, x431x, x16408x, x16414x, x69x, x16421x, n_n4963, n_n4960, n_n4964, x22065x, n_n5012, n_n5016, n_n5009, n_n5013;
	wire n_n4919, x341x, x16458x, x250x, n_n4827, n_n4474, x199x, n_n4825, n_n4879, n_n4938, n_n5043, n_n5294, n_n4916, n_n4930, n_n4947, x96x, n_n5206, n_n5204, x12091x, x12097x, n_n5089;
	wire n_n5116, n_n5063, x344x, x12099x, x12100x, n_n5258, n_n5232, n_n5255, n_n5216, n_n5222, x12109x, n_n4393, n_n4669, n_n4668, n_n4966, n_n4968, n_n5067, n_n5069, n_n5243, n_n5299, n_n4364;
	wire n_n3533, n_n1308, x316x, x11749x, x306x, n_n4914, x352x, x11786x, n_n1075, x166x, x22155x, n_n1064, n_n4807, x85x, n_n4851, n_n4836, x11773x, x372x, x11780x, n_n5161, n_n4482;
	wire n_n4704, n_n5105, n_n5120, n_n5127, n_n5273, n_n4398, n_n4522, n_n4246, n_n4670, n_n4732, n_n5086, n_n5087, n_n881, n_n4591, n_n4592, n_n4083, n_n3520, n_n4582, n_n4586, x14093x, n_n3348;
	wire x461x, x22120x, n_n3326, n_n2643, n_n5323, n_n4569, n_n4579, x14100x, x14101x, n_n4538, n_n3871, n_n4556, x14103x, n_n3350, x212x, n_n4536, x14112x, x14115x, x14117x, n_n5033, n_n5051;
	wire n_n5072, n_n5082, x13719x, n_n5079, n_n5065, x13720x, n_n3152, n_n5039, n_n5103, n_n5102, n_n4395, x281x, n_n4394, x216x, n_n4387, x425x, x22099x, x15045x, n_n4419, n_n4411, n_n4412;
	wire x15051x, n_n4360, n_n4483, n_n5115, x290x, n_n4144, x34x, x289x, x428x, x176x, x186x, x16522x, x16532x, n_n4349, x171x, n_n4376, n_n4502, x387x, n_n4610, n_n4614, n_n4600;
	wire n_n4603, x16632x, x119x, x271x, n_n5328, n_n5249, n_n5233, n_n5236, n_n5290, x392x, n_n5217, x449x, x16778x, x16777x, x16779x, n_n4833, n_n4940, x373x, n_n5128, x12253x, n_n4129;
	wire n_n3019, n_n4655, n_n4658, n_n4342, x22196x, n_n4622, n_n5073, n_n4152, x11790x, x11791x, n_n4932, x411x, x22175x, x11796x, n_n4971, x11802x, x11806x, x22160x, n_n4973, x11814x, n_n1077;
	wire x11824x, n_n4892, x11828x, x11830x, n_n1002, n_n5011, n_n5061, n_n5070, n_n5076, n_n5135, n_n5201, n_n5237, n_n5252, n_n4161, n_n5084, n_n5276, x22215x, n_n4082, x13149x, x22121x, n_n4068;
	wire n_n4196, x390x, x13166x, x389x, x326x, n_n4065, x13163x, x13178x, x13180x, n_n834, n_n4063, x13182x, x13186x, x22127x, n_n4060, x13199x, x42x, x13213x, x154x, x13204x, n_n4058;
	wire x331x, x13208x, n_n4944, x13209x, x210x, n_n814, x13226x, x317x, x13224x, x13227x, x13232x, n_n4172, n_n1970, x137x, x22128x, x94x, x13237x, x221x, x13244x, n_n4219, x13245x;
	wire n_n4716, n_n4713, x13251x, x13252x, x367x, x30x, x13253x, n_n4693, x81x, x426x, x22220x, x13269x, x312x, x22126x, n_n4078, x157x, x339x, n_n4680, x80x, x13264x, x22125x;
	wire n_n5078, n_n5083, x123x, x122x, x232x, x160x, x14653x, n_n5077, x159x, x22100x, n_n5169, n_n5197, n_n5176, n_n5205, n_n5211, x14253x, n_n5226, n_n5218, x14254x, n_n5295, n_n5256;
	wire n_n5257, n_n5283, n_n4370, n_n4435, n_n4493, x14284x, n_n4626, x14296x, n_n4721, n_n4678, n_n5158, n_n3427, n_n5150, n_n5147, x22115x, n_n3305, x13834x, n_n3318, x229x, x13841x, x13842x;
	wire n_n901, x14122x, n_n3358, x14128x, x14130x, n_n3285, n_n2059, n_n4423, x14138x, x14139x, x14147x, x14143x, x14146x, n_n3286, n_n3162, x153x, n_n3461, x304x, n_n2601, x14900x, n_n2727;
	wire x14920x, n_n2718, x22210x, x14955x, n_n1973, n_n2710, x58x, x22091x, n_n4684, x86x, n_n4694, x219x, x442x, n_n4705, x464x, n_n856, n_n5118, n_n5229, n_n5228, n_n889, n_n4541;
	wire n_n4677, x338x, x414x, x16724x, n_n4893, x16785x, n_n2095, x14962x, n_n5159, n_n5151, x406x, x12261x, n_n1443, x208x, x22205x, n_n1432, x12124x, n_n4627, n_n4955, n_n1128, x420x;
	wire x11592x, x11505x, x22169x, x458x, n_n1066, x11842x, x457x, x22159x, x11900x, x113x, x22182x, n_n5199, n_n5260, n_n5272, n_n4501, n_n5220, n_n5125, n_n5140, x13284x, n_n4039, x22202x;
	wire n_n4038, n_n5196, n_n5195, n_n2670, x13302x, x13306x, x144x, x13317x, x11915x, n_n4041, x13314x, n_n5126, x13322x, x13323x, x13293x, x13296x, n_n4026, x217x, x333x, x13332x, n_n4028;
	wire n_n5271, x22187x, x13348x, n_n5253, x13338x, n_n5259, x13339x, x13343x, n_n4031, n_n1530, n_n2290, x13351x, x13353x, n_n4032, x13361x, x223x, x384x, x450x, x13363x, x441x, x13370x;
	wire x13371x, x343x, x13383x, x404x, x13396x, x13398x, n_n1952, n_n789, x13394x, x13414x, x13405x, n_n4047, x22124x, n_n4048, x13420x, n_n4650, n_n5071, n_n5250, x13789x, n_n3333, x13994x;
	wire n_n3315, n_n4654, x13887x, x11854x, x192x, x193x, x13893x, x13894x, x248x, n_n3317, n_n4273, x22113x, n_n3367, x301x, x14163x, x14159x, n_n3288, x14170x, n_n3363, x14175x, n_n3362;
	wire x14179x, x14180x, n_n3287, n_n3369, x14186x, n_n4322, n_n4323, x363x, n_n3370, x22112x, x14193x, x227x, x427x, x332x, x22179x, n_n5208, x22217x, x22199x, x451x, x62x, x183x;
	wire x16695x, x22059x, x22225x, x16750x, x419x, x438x, n_n5334, n_n5333, n_n4813, x16812x, x16813x, n_n5225, n_n5224, x12287x, n_n3382, n_n1162, x11563x, x11913x, x28x, n_n4446, n_n4961;
	wire n_n5265, n_n1648, x22123x, x13438x, n_n4094, x91x, x13471x, x13091x, x22207x, n_n4086, x379x, x13477x, x13480x, x13450x, x13451x, n_n4079, x13464x, x13466x, x13487x, x13488x, x13503x;
	wire n_n4092, n_n4103, x13519x, n_n4097, x13533x, x13539x, x13544x, x55x, x22122x, x13551x, x14393x, x14394x, n_n2761, n_n3714, x14403x, x14404x, n_n4550, x22214x, n_n3722, x14416x, x14418x;
	wire x14424x, x14429x, n_n3719, x46x, x22168x, x14434x, n_n3329, x13924x, x13925x, x13793x, x13795x, x13799x, n_n3332, x13805x, x22116x, x13820x, n_n1988, n_n3327, x13825x, x13857x, x22119x;
	wire x22118x, n_n4910, x13868x, x138x, n_n3124, x13910x, x13903x, x13899x, x13909x, x456x, x357x, n_n5008, x13454x, x15754x, x15757x, x22172x, n_n5317, n_n2803, x22216x, x146x, x320x;
	wire x15177x, x22185x, x267x, x15191x, x22188x, x15192x, x15196x, n_n2651, n_n2566, x207x, x15203x, n_n5227, n_n5219, n_n1521, x328x, x22151x, n_n1093, x11980x, n_n1068, x11925x, x22193x;
	wire n_n1049, n_n1047, n_n1048, x22156x, x11940x, x175x, x11950x, x22189x, x11959x, x22192x, x22136x, n_n5210, x13568x, x13565x, x13457x, x22103x, n_n3708, n_n3710, x22102x, x14357x, x14362x;
	wire n_n3711, x22101x, x14371x, x14442x, x14467x, n_n3737, x14472x, n_n3736, x14511x, n_n3740, x14486x, x14488x, x14506x, x14494x, x22108x, x360x, x14527x, x13929x, x13930x, x13947x, x13950x;
	wire n_n3299, x446x, x434x, n_n3297, x13959x, x13960x, n_n3265, x13963x, x13965x, n_n3296, x12372x, x204x, x13973x, x13974x, x13976x, x13943x, n_n3293, n_n1167, n_n783, x14015x, x14006x;
	wire x14007x, x14014x, n_n3269, x14021x, x14022x, x14040x, x14041x, n_n3267, x14054x, x14056x, x14057x, n_n2665, n_n3300, x14047x, n_n3301, x14063x, x14065x, n_n4334, n_n1646, x48x, x383x;
	wire x15208x, x15210x, n_n5209, x22095x, x15061x, x15062x, n_n910, x15074x, x15075x, x128x, x291x, x15066x, x22224x, n_n2630, x15080x, x15081x, n_n1677, x15082x, n_n2629, x15091x, x15093x;
	wire x15096x, x15098x, x15101x, x22097x, n_n2619, x22167x, n_n2618, x15119x, x15120x, x15126x, n_n2621, x22096x, n_n2615, n_n2030, x15137x, x15139x, x82x, x15146x, x15147x, x469x, x15152x;
	wire x22098x, x133x, n_n1532, x12265x, n_n1444, x12349x, n_n1435, x22152x, n_n1067, x22166x, x11571x, x284x, x11603x, n_n897, n_n3355, n_n3354, x14207x, x15758x, n_n3037, x15562x, x22085x;
	wire x22183x, x14953x, x22094x, x88x, x15246x, x265x, x297x, x394x, x361x, n_n801, x405x, x12354x, n_n1436, x225x, x432x, x11859x, x22154x, x12003x, x22194x, x22153x, x12019x;
	wire x12025x, x13003x, x13010x, x12729x, x12730x, x12736x, n_n696, x15268x, x15271x, x139x, x22149x, n_n954, x11647x, x11648x, x11653x, x11654x, n_n725, x13025x, x13026x, x12741x, x22171x;
	wire x52x, x150x, x12745x, x13513x, x12497x, x12446x, x12269x, x12270x, n_n1439, x12278x, x12280x, x22145x, x22181x, x12301x, x12302x, x22144x, x11675x, x11676x, x12873x, n_n667, n_n761;
	wire x12878x, x12879x, x12880x, x12884x, x12889x, x12897x, x12896x, x22203x, x22211x, x303x, x13580x, x13587x, x13592x, x13593x, x13599x, x13600x, x22142x, x12357x, x12358x, x12952x, n_n664;
	wire x12958x, x12960x, x12902x, x12903x, x22130x, n_n681, x209x, x12913x, x12914x, x12921x, x12920x, x12922x, x12929x, x12928x, n_n684, x12939x, n_n683, x22129x, x12945x, x13538x, n_n2058;
	wire x22148x, x305x, x12662x, x22135x, x12669x, x13449x, x401x, x12492x, x12231x, x11867x, x11868x, x22089x, x12369x, x12364x, n_n1429, x12368x, x12379x, x11682x, n_n951, x11688x, x11689x;
	wire x22139x, n_n1489, x12531x, x12533x, x12415x, x12410x, x13027x, x22137x, n_n1482, x270x, x22138x, x22209x, x12559x, x12558x, x22170x, x617x, x15837x, x22074x, x22178x, n_n2982, x22088x;
	wire x16182x, n_n1840, x22066x, n_n1839, x15956x, x15957x, x15962x, x15963x, x15967x, x15968x, x15972x, x15973x, x12784x, x12785x, n_n691, x12724x, x12725x, x22191x, n_n632, x12767x, x12757x;
	wire x12758x, x12763x, n_n702, x12772x, x12773x, x12791x, n_n706, x12794x, x12795x, n_n709, x12804x, n_n710, x12811x, x12812x, x22132x, n_n704, x12824x, x12834x, n_n689, x12840x, x12841x;
	wire x12842x, x22131x, n_n686, x12854x, x12856x, x12863x, x15763x, x16146x, x16155x, n_n1852, x16166x, x16167x, n_n1850, x16177x, x16178x, x22212x, n_n662, x12975x, n_n661, x12980x, x12981x;
	wire x12989x, n_n670, n_n671, x12995x, x12996x, x13056x, x16189x, x16190x, x16192x, x16198x, x16197x, x22070x, n_n1858, n_n1857, x16211x, x16212x, x16215x, x22075x, x15886x, x15879x, x13029x;
	wire n_n722, x346x, x13036x, x13037x, x13038x, x13044x, x22173x, x15519x, x22213x, x15771x, x15778x, x15775x, x15777x, x22083x, x16095x, x16104x, x16227x, x11713x, x13051x, x22134x, x13079x;
	wire x13102x, n_n715, x13108x, x13109x, x22133x, n_n714, x13120x, x13121x, x13122x, x13126x, x15655x, x15712x, x15714x, x15713x, x22158x, x11875x, x22109x, x14485x, x15657x, x15719x, n_n2962;
	wire x15728x, x15725x, x14620x, x22084x, x15734x, x22080x, x15876x, x14504x, x16002x, x16064x, x22079x, x11881x, x11882x, x14703x, x16273x, x14761x, x15735x, x15737x, x15783x, x11742x, x22174x;
	wire x13141x, x13727x, x14059x, x14338x, x14846x, x14847x, x14887x, x14889x, x16462x, x22058x, x16818x, x16819x;

	assign o_1_ = (((!x12042x) & (!x12038x) & (!n_n1007) & (!n_n1009) & (x12041x)) + ((!x12042x) & (!x12038x) & (!n_n1007) & (n_n1009) & (!x12041x)) + ((!x12042x) & (!x12038x) & (!n_n1007) & (n_n1009) & (x12041x)) + ((!x12042x) & (!x12038x) & (n_n1007) & (!n_n1009) & (!x12041x)) + ((!x12042x) & (!x12038x) & (n_n1007) & (!n_n1009) & (x12041x)) + ((!x12042x) & (!x12038x) & (n_n1007) & (n_n1009) & (!x12041x)) + ((!x12042x) & (!x12038x) & (n_n1007) & (n_n1009) & (x12041x)) + ((!x12042x) & (x12038x) & (!n_n1007) & (!n_n1009) & (!x12041x)) + ((!x12042x) & (x12038x) & (!n_n1007) & (!n_n1009) & (x12041x)) + ((!x12042x) & (x12038x) & (!n_n1007) & (n_n1009) & (!x12041x)) + ((!x12042x) & (x12038x) & (!n_n1007) & (n_n1009) & (x12041x)) + ((!x12042x) & (x12038x) & (n_n1007) & (!n_n1009) & (!x12041x)) + ((!x12042x) & (x12038x) & (n_n1007) & (!n_n1009) & (x12041x)) + ((!x12042x) & (x12038x) & (n_n1007) & (n_n1009) & (!x12041x)) + ((!x12042x) & (x12038x) & (n_n1007) & (n_n1009) & (x12041x)) + ((x12042x) & (!x12038x) & (!n_n1007) & (!n_n1009) & (!x12041x)) + ((x12042x) & (!x12038x) & (!n_n1007) & (!n_n1009) & (x12041x)) + ((x12042x) & (!x12038x) & (!n_n1007) & (n_n1009) & (!x12041x)) + ((x12042x) & (!x12038x) & (!n_n1007) & (n_n1009) & (x12041x)) + ((x12042x) & (!x12038x) & (n_n1007) & (!n_n1009) & (!x12041x)) + ((x12042x) & (!x12038x) & (n_n1007) & (!n_n1009) & (x12041x)) + ((x12042x) & (!x12038x) & (n_n1007) & (n_n1009) & (!x12041x)) + ((x12042x) & (!x12038x) & (n_n1007) & (n_n1009) & (x12041x)) + ((x12042x) & (x12038x) & (!n_n1007) & (!n_n1009) & (!x12041x)) + ((x12042x) & (x12038x) & (!n_n1007) & (!n_n1009) & (x12041x)) + ((x12042x) & (x12038x) & (!n_n1007) & (n_n1009) & (!x12041x)) + ((x12042x) & (x12038x) & (!n_n1007) & (n_n1009) & (x12041x)) + ((x12042x) & (x12038x) & (n_n1007) & (!n_n1009) & (!x12041x)) + ((x12042x) & (x12038x) & (n_n1007) & (!n_n1009) & (x12041x)) + ((x12042x) & (x12038x) & (n_n1007) & (n_n1009) & (!x12041x)) + ((x12042x) & (x12038x) & (n_n1007) & (n_n1009) & (x12041x)));
	assign o_2_ = (((!x12589x) & (!x12151x) & (!x12152x) & (!n_n1398) & (n_n1392)) + ((!x12589x) & (!x12151x) & (!x12152x) & (n_n1398) & (!n_n1392)) + ((!x12589x) & (!x12151x) & (!x12152x) & (n_n1398) & (n_n1392)) + ((!x12589x) & (!x12151x) & (x12152x) & (!n_n1398) & (!n_n1392)) + ((!x12589x) & (!x12151x) & (x12152x) & (!n_n1398) & (n_n1392)) + ((!x12589x) & (!x12151x) & (x12152x) & (n_n1398) & (!n_n1392)) + ((!x12589x) & (!x12151x) & (x12152x) & (n_n1398) & (n_n1392)) + ((!x12589x) & (x12151x) & (!x12152x) & (!n_n1398) & (!n_n1392)) + ((!x12589x) & (x12151x) & (!x12152x) & (!n_n1398) & (n_n1392)) + ((!x12589x) & (x12151x) & (!x12152x) & (n_n1398) & (!n_n1392)) + ((!x12589x) & (x12151x) & (!x12152x) & (n_n1398) & (n_n1392)) + ((!x12589x) & (x12151x) & (x12152x) & (!n_n1398) & (!n_n1392)) + ((!x12589x) & (x12151x) & (x12152x) & (!n_n1398) & (n_n1392)) + ((!x12589x) & (x12151x) & (x12152x) & (n_n1398) & (!n_n1392)) + ((!x12589x) & (x12151x) & (x12152x) & (n_n1398) & (n_n1392)) + ((x12589x) & (!x12151x) & (!x12152x) & (!n_n1398) & (!n_n1392)) + ((x12589x) & (!x12151x) & (!x12152x) & (!n_n1398) & (n_n1392)) + ((x12589x) & (!x12151x) & (!x12152x) & (n_n1398) & (!n_n1392)) + ((x12589x) & (!x12151x) & (!x12152x) & (n_n1398) & (n_n1392)) + ((x12589x) & (!x12151x) & (x12152x) & (!n_n1398) & (!n_n1392)) + ((x12589x) & (!x12151x) & (x12152x) & (!n_n1398) & (n_n1392)) + ((x12589x) & (!x12151x) & (x12152x) & (n_n1398) & (!n_n1392)) + ((x12589x) & (!x12151x) & (x12152x) & (n_n1398) & (n_n1392)) + ((x12589x) & (x12151x) & (!x12152x) & (!n_n1398) & (!n_n1392)) + ((x12589x) & (x12151x) & (!x12152x) & (!n_n1398) & (n_n1392)) + ((x12589x) & (x12151x) & (!x12152x) & (n_n1398) & (!n_n1392)) + ((x12589x) & (x12151x) & (!x12152x) & (n_n1398) & (n_n1392)) + ((x12589x) & (x12151x) & (x12152x) & (!n_n1398) & (!n_n1392)) + ((x12589x) & (x12151x) & (x12152x) & (!n_n1398) & (n_n1392)) + ((x12589x) & (x12151x) & (x12152x) & (n_n1398) & (!n_n1392)) + ((x12589x) & (x12151x) & (x12152x) & (n_n1398) & (n_n1392)));
	assign o_0_ = (((!x13147x) & (!x13136x) & (x13137x)) + ((!x13147x) & (x13136x) & (!x13137x)) + ((!x13147x) & (x13136x) & (x13137x)) + ((x13147x) & (!x13136x) & (!x13137x)) + ((x13147x) & (!x13136x) & (x13137x)) + ((x13147x) & (x13136x) & (!x13137x)) + ((x13147x) & (x13136x) & (x13137x)));
	assign o_9_ = (((!x13684x) & (!x13573x) & (x13574x)) + ((!x13684x) & (x13573x) & (!x13574x)) + ((!x13684x) & (x13573x) & (x13574x)) + ((x13684x) & (!x13573x) & (!x13574x)) + ((x13684x) & (!x13573x) & (x13574x)) + ((x13684x) & (x13573x) & (!x13574x)) + ((x13684x) & (x13573x) & (x13574x)));
	assign o_7_ = (((!x14222x) & (!x14216x) & (!n_n3251) & (n_n3253)) + ((!x14222x) & (!x14216x) & (n_n3251) & (!n_n3253)) + ((!x14222x) & (!x14216x) & (n_n3251) & (n_n3253)) + ((!x14222x) & (x14216x) & (!n_n3251) & (!n_n3253)) + ((!x14222x) & (x14216x) & (!n_n3251) & (n_n3253)) + ((!x14222x) & (x14216x) & (n_n3251) & (!n_n3253)) + ((!x14222x) & (x14216x) & (n_n3251) & (n_n3253)) + ((x14222x) & (!x14216x) & (!n_n3251) & (!n_n3253)) + ((x14222x) & (!x14216x) & (!n_n3251) & (n_n3253)) + ((x14222x) & (!x14216x) & (n_n3251) & (!n_n3253)) + ((x14222x) & (!x14216x) & (n_n3251) & (n_n3253)) + ((x14222x) & (x14216x) & (!n_n3251) & (!n_n3253)) + ((x14222x) & (x14216x) & (!n_n3251) & (n_n3253)) + ((x14222x) & (x14216x) & (n_n3251) & (!n_n3253)) + ((x14222x) & (x14216x) & (n_n3251) & (n_n3253)));
	assign o_8_ = (((!x14780x) & (!n_n3623) & (!n_n3624) & (!x14775x) & (x14778x)) + ((!x14780x) & (!n_n3623) & (!n_n3624) & (x14775x) & (!x14778x)) + ((!x14780x) & (!n_n3623) & (!n_n3624) & (x14775x) & (x14778x)) + ((!x14780x) & (!n_n3623) & (n_n3624) & (!x14775x) & (!x14778x)) + ((!x14780x) & (!n_n3623) & (n_n3624) & (!x14775x) & (x14778x)) + ((!x14780x) & (!n_n3623) & (n_n3624) & (x14775x) & (!x14778x)) + ((!x14780x) & (!n_n3623) & (n_n3624) & (x14775x) & (x14778x)) + ((!x14780x) & (n_n3623) & (!n_n3624) & (!x14775x) & (!x14778x)) + ((!x14780x) & (n_n3623) & (!n_n3624) & (!x14775x) & (x14778x)) + ((!x14780x) & (n_n3623) & (!n_n3624) & (x14775x) & (!x14778x)) + ((!x14780x) & (n_n3623) & (!n_n3624) & (x14775x) & (x14778x)) + ((!x14780x) & (n_n3623) & (n_n3624) & (!x14775x) & (!x14778x)) + ((!x14780x) & (n_n3623) & (n_n3624) & (!x14775x) & (x14778x)) + ((!x14780x) & (n_n3623) & (n_n3624) & (x14775x) & (!x14778x)) + ((!x14780x) & (n_n3623) & (n_n3624) & (x14775x) & (x14778x)) + ((x14780x) & (!n_n3623) & (!n_n3624) & (!x14775x) & (!x14778x)) + ((x14780x) & (!n_n3623) & (!n_n3624) & (!x14775x) & (x14778x)) + ((x14780x) & (!n_n3623) & (!n_n3624) & (x14775x) & (!x14778x)) + ((x14780x) & (!n_n3623) & (!n_n3624) & (x14775x) & (x14778x)) + ((x14780x) & (!n_n3623) & (n_n3624) & (!x14775x) & (!x14778x)) + ((x14780x) & (!n_n3623) & (n_n3624) & (!x14775x) & (x14778x)) + ((x14780x) & (!n_n3623) & (n_n3624) & (x14775x) & (!x14778x)) + ((x14780x) & (!n_n3623) & (n_n3624) & (x14775x) & (x14778x)) + ((x14780x) & (n_n3623) & (!n_n3624) & (!x14775x) & (!x14778x)) + ((x14780x) & (n_n3623) & (!n_n3624) & (!x14775x) & (x14778x)) + ((x14780x) & (n_n3623) & (!n_n3624) & (x14775x) & (!x14778x)) + ((x14780x) & (n_n3623) & (!n_n3624) & (x14775x) & (x14778x)) + ((x14780x) & (n_n3623) & (n_n3624) & (!x14775x) & (!x14778x)) + ((x14780x) & (n_n3623) & (n_n3624) & (!x14775x) & (x14778x)) + ((x14780x) & (n_n3623) & (n_n3624) & (x14775x) & (!x14778x)) + ((x14780x) & (n_n3623) & (n_n3624) & (x14775x) & (x14778x)));
	assign o_5_ = (((!x15301x) & (!n_n2523) & (x15300x)) + ((!x15301x) & (n_n2523) & (!x15300x)) + ((!x15301x) & (n_n2523) & (x15300x)) + ((x15301x) & (!n_n2523) & (!x15300x)) + ((x15301x) & (!n_n2523) & (x15300x)) + ((x15301x) & (n_n2523) & (!x15300x)) + ((x15301x) & (n_n2523) & (x15300x)));
	assign o_6_ = (((!x15817x) & (!n_n2898) & (x15816x)) + ((!x15817x) & (n_n2898) & (!x15816x)) + ((!x15817x) & (n_n2898) & (x15816x)) + ((x15817x) & (!n_n2898) & (!x15816x)) + ((x15817x) & (!n_n2898) & (x15816x)) + ((x15817x) & (n_n2898) & (!x15816x)) + ((x15817x) & (n_n2898) & (x15816x)));
	assign o_3_ = (((!x16324x) & (!n_n1706) & (!x15943x) & (!n_n1784) & (x16320x)) + ((!x16324x) & (!n_n1706) & (!x15943x) & (n_n1784) & (!x16320x)) + ((!x16324x) & (!n_n1706) & (!x15943x) & (n_n1784) & (x16320x)) + ((!x16324x) & (!n_n1706) & (x15943x) & (!n_n1784) & (!x16320x)) + ((!x16324x) & (!n_n1706) & (x15943x) & (!n_n1784) & (x16320x)) + ((!x16324x) & (!n_n1706) & (x15943x) & (n_n1784) & (!x16320x)) + ((!x16324x) & (!n_n1706) & (x15943x) & (n_n1784) & (x16320x)) + ((!x16324x) & (n_n1706) & (!x15943x) & (!n_n1784) & (!x16320x)) + ((!x16324x) & (n_n1706) & (!x15943x) & (!n_n1784) & (x16320x)) + ((!x16324x) & (n_n1706) & (!x15943x) & (n_n1784) & (!x16320x)) + ((!x16324x) & (n_n1706) & (!x15943x) & (n_n1784) & (x16320x)) + ((!x16324x) & (n_n1706) & (x15943x) & (!n_n1784) & (!x16320x)) + ((!x16324x) & (n_n1706) & (x15943x) & (!n_n1784) & (x16320x)) + ((!x16324x) & (n_n1706) & (x15943x) & (n_n1784) & (!x16320x)) + ((!x16324x) & (n_n1706) & (x15943x) & (n_n1784) & (x16320x)) + ((x16324x) & (!n_n1706) & (!x15943x) & (!n_n1784) & (!x16320x)) + ((x16324x) & (!n_n1706) & (!x15943x) & (!n_n1784) & (x16320x)) + ((x16324x) & (!n_n1706) & (!x15943x) & (n_n1784) & (!x16320x)) + ((x16324x) & (!n_n1706) & (!x15943x) & (n_n1784) & (x16320x)) + ((x16324x) & (!n_n1706) & (x15943x) & (!n_n1784) & (!x16320x)) + ((x16324x) & (!n_n1706) & (x15943x) & (!n_n1784) & (x16320x)) + ((x16324x) & (!n_n1706) & (x15943x) & (n_n1784) & (!x16320x)) + ((x16324x) & (!n_n1706) & (x15943x) & (n_n1784) & (x16320x)) + ((x16324x) & (n_n1706) & (!x15943x) & (!n_n1784) & (!x16320x)) + ((x16324x) & (n_n1706) & (!x15943x) & (!n_n1784) & (x16320x)) + ((x16324x) & (n_n1706) & (!x15943x) & (n_n1784) & (!x16320x)) + ((x16324x) & (n_n1706) & (!x15943x) & (n_n1784) & (x16320x)) + ((x16324x) & (n_n1706) & (x15943x) & (!n_n1784) & (!x16320x)) + ((x16324x) & (n_n1706) & (x15943x) & (!n_n1784) & (x16320x)) + ((x16324x) & (n_n1706) & (x15943x) & (n_n1784) & (!x16320x)) + ((x16324x) & (n_n1706) & (x15943x) & (n_n1784) & (x16320x)));
	assign o_4_ = (((!x16831x) & (x16832x)) + ((x16831x) & (!x16832x)) + ((x16831x) & (x16832x)));
	assign x12042x = (((!n_n1014) & (!n_n1013) & (!x11894x) & (!n_n1010) & (n_n1012)) + ((!n_n1014) & (!n_n1013) & (!x11894x) & (n_n1010) & (!n_n1012)) + ((!n_n1014) & (!n_n1013) & (!x11894x) & (n_n1010) & (n_n1012)) + ((!n_n1014) & (!n_n1013) & (x11894x) & (!n_n1010) & (!n_n1012)) + ((!n_n1014) & (!n_n1013) & (x11894x) & (!n_n1010) & (n_n1012)) + ((!n_n1014) & (!n_n1013) & (x11894x) & (n_n1010) & (!n_n1012)) + ((!n_n1014) & (!n_n1013) & (x11894x) & (n_n1010) & (n_n1012)) + ((!n_n1014) & (n_n1013) & (!x11894x) & (!n_n1010) & (!n_n1012)) + ((!n_n1014) & (n_n1013) & (!x11894x) & (!n_n1010) & (n_n1012)) + ((!n_n1014) & (n_n1013) & (!x11894x) & (n_n1010) & (!n_n1012)) + ((!n_n1014) & (n_n1013) & (!x11894x) & (n_n1010) & (n_n1012)) + ((!n_n1014) & (n_n1013) & (x11894x) & (!n_n1010) & (!n_n1012)) + ((!n_n1014) & (n_n1013) & (x11894x) & (!n_n1010) & (n_n1012)) + ((!n_n1014) & (n_n1013) & (x11894x) & (n_n1010) & (!n_n1012)) + ((!n_n1014) & (n_n1013) & (x11894x) & (n_n1010) & (n_n1012)) + ((n_n1014) & (!n_n1013) & (!x11894x) & (!n_n1010) & (!n_n1012)) + ((n_n1014) & (!n_n1013) & (!x11894x) & (!n_n1010) & (n_n1012)) + ((n_n1014) & (!n_n1013) & (!x11894x) & (n_n1010) & (!n_n1012)) + ((n_n1014) & (!n_n1013) & (!x11894x) & (n_n1010) & (n_n1012)) + ((n_n1014) & (!n_n1013) & (x11894x) & (!n_n1010) & (!n_n1012)) + ((n_n1014) & (!n_n1013) & (x11894x) & (!n_n1010) & (n_n1012)) + ((n_n1014) & (!n_n1013) & (x11894x) & (n_n1010) & (!n_n1012)) + ((n_n1014) & (!n_n1013) & (x11894x) & (n_n1010) & (n_n1012)) + ((n_n1014) & (n_n1013) & (!x11894x) & (!n_n1010) & (!n_n1012)) + ((n_n1014) & (n_n1013) & (!x11894x) & (!n_n1010) & (n_n1012)) + ((n_n1014) & (n_n1013) & (!x11894x) & (n_n1010) & (!n_n1012)) + ((n_n1014) & (n_n1013) & (!x11894x) & (n_n1010) & (n_n1012)) + ((n_n1014) & (n_n1013) & (x11894x) & (!n_n1010) & (!n_n1012)) + ((n_n1014) & (n_n1013) & (x11894x) & (!n_n1010) & (n_n1012)) + ((n_n1014) & (n_n1013) & (x11894x) & (n_n1010) & (!n_n1012)) + ((n_n1014) & (n_n1013) & (x11894x) & (n_n1010) & (n_n1012)));
	assign x12038x = (((!n_n1020) & (!n_n1052) & (!n_n1054) & (!x11977x) & (x12036x)) + ((!n_n1020) & (!n_n1052) & (!n_n1054) & (x11977x) & (!x12036x)) + ((!n_n1020) & (!n_n1052) & (!n_n1054) & (x11977x) & (x12036x)) + ((!n_n1020) & (!n_n1052) & (n_n1054) & (!x11977x) & (!x12036x)) + ((!n_n1020) & (!n_n1052) & (n_n1054) & (!x11977x) & (x12036x)) + ((!n_n1020) & (!n_n1052) & (n_n1054) & (x11977x) & (!x12036x)) + ((!n_n1020) & (!n_n1052) & (n_n1054) & (x11977x) & (x12036x)) + ((!n_n1020) & (n_n1052) & (!n_n1054) & (!x11977x) & (!x12036x)) + ((!n_n1020) & (n_n1052) & (!n_n1054) & (!x11977x) & (x12036x)) + ((!n_n1020) & (n_n1052) & (!n_n1054) & (x11977x) & (!x12036x)) + ((!n_n1020) & (n_n1052) & (!n_n1054) & (x11977x) & (x12036x)) + ((!n_n1020) & (n_n1052) & (n_n1054) & (!x11977x) & (!x12036x)) + ((!n_n1020) & (n_n1052) & (n_n1054) & (!x11977x) & (x12036x)) + ((!n_n1020) & (n_n1052) & (n_n1054) & (x11977x) & (!x12036x)) + ((!n_n1020) & (n_n1052) & (n_n1054) & (x11977x) & (x12036x)) + ((n_n1020) & (!n_n1052) & (!n_n1054) & (!x11977x) & (!x12036x)) + ((n_n1020) & (!n_n1052) & (!n_n1054) & (!x11977x) & (x12036x)) + ((n_n1020) & (!n_n1052) & (!n_n1054) & (x11977x) & (!x12036x)) + ((n_n1020) & (!n_n1052) & (!n_n1054) & (x11977x) & (x12036x)) + ((n_n1020) & (!n_n1052) & (n_n1054) & (!x11977x) & (!x12036x)) + ((n_n1020) & (!n_n1052) & (n_n1054) & (!x11977x) & (x12036x)) + ((n_n1020) & (!n_n1052) & (n_n1054) & (x11977x) & (!x12036x)) + ((n_n1020) & (!n_n1052) & (n_n1054) & (x11977x) & (x12036x)) + ((n_n1020) & (n_n1052) & (!n_n1054) & (!x11977x) & (!x12036x)) + ((n_n1020) & (n_n1052) & (!n_n1054) & (!x11977x) & (x12036x)) + ((n_n1020) & (n_n1052) & (!n_n1054) & (x11977x) & (!x12036x)) + ((n_n1020) & (n_n1052) & (!n_n1054) & (x11977x) & (x12036x)) + ((n_n1020) & (n_n1052) & (n_n1054) & (!x11977x) & (!x12036x)) + ((n_n1020) & (n_n1052) & (n_n1054) & (!x11977x) & (x12036x)) + ((n_n1020) & (n_n1052) & (n_n1054) & (x11977x) & (!x12036x)) + ((n_n1020) & (n_n1052) & (n_n1054) & (x11977x) & (x12036x)));
	assign n_n1007 = (((!n_n1017) & (!n_n1045) & (!x11953x) & (!x11960x) & (x11961x)) + ((!n_n1017) & (!n_n1045) & (!x11953x) & (x11960x) & (!x11961x)) + ((!n_n1017) & (!n_n1045) & (!x11953x) & (x11960x) & (x11961x)) + ((!n_n1017) & (!n_n1045) & (x11953x) & (!x11960x) & (!x11961x)) + ((!n_n1017) & (!n_n1045) & (x11953x) & (!x11960x) & (x11961x)) + ((!n_n1017) & (!n_n1045) & (x11953x) & (x11960x) & (!x11961x)) + ((!n_n1017) & (!n_n1045) & (x11953x) & (x11960x) & (x11961x)) + ((!n_n1017) & (n_n1045) & (!x11953x) & (!x11960x) & (!x11961x)) + ((!n_n1017) & (n_n1045) & (!x11953x) & (!x11960x) & (x11961x)) + ((!n_n1017) & (n_n1045) & (!x11953x) & (x11960x) & (!x11961x)) + ((!n_n1017) & (n_n1045) & (!x11953x) & (x11960x) & (x11961x)) + ((!n_n1017) & (n_n1045) & (x11953x) & (!x11960x) & (!x11961x)) + ((!n_n1017) & (n_n1045) & (x11953x) & (!x11960x) & (x11961x)) + ((!n_n1017) & (n_n1045) & (x11953x) & (x11960x) & (!x11961x)) + ((!n_n1017) & (n_n1045) & (x11953x) & (x11960x) & (x11961x)) + ((n_n1017) & (!n_n1045) & (!x11953x) & (!x11960x) & (!x11961x)) + ((n_n1017) & (!n_n1045) & (!x11953x) & (!x11960x) & (x11961x)) + ((n_n1017) & (!n_n1045) & (!x11953x) & (x11960x) & (!x11961x)) + ((n_n1017) & (!n_n1045) & (!x11953x) & (x11960x) & (x11961x)) + ((n_n1017) & (!n_n1045) & (x11953x) & (!x11960x) & (!x11961x)) + ((n_n1017) & (!n_n1045) & (x11953x) & (!x11960x) & (x11961x)) + ((n_n1017) & (!n_n1045) & (x11953x) & (x11960x) & (!x11961x)) + ((n_n1017) & (!n_n1045) & (x11953x) & (x11960x) & (x11961x)) + ((n_n1017) & (n_n1045) & (!x11953x) & (!x11960x) & (!x11961x)) + ((n_n1017) & (n_n1045) & (!x11953x) & (!x11960x) & (x11961x)) + ((n_n1017) & (n_n1045) & (!x11953x) & (x11960x) & (!x11961x)) + ((n_n1017) & (n_n1045) & (!x11953x) & (x11960x) & (x11961x)) + ((n_n1017) & (n_n1045) & (x11953x) & (!x11960x) & (!x11961x)) + ((n_n1017) & (n_n1045) & (x11953x) & (!x11960x) & (x11961x)) + ((n_n1017) & (n_n1045) & (x11953x) & (x11960x) & (!x11961x)) + ((n_n1017) & (n_n1045) & (x11953x) & (x11960x) & (x11961x)));
	assign n_n1009 = (((!n_n1023) & (!n_n1061) & (!n_n1062) & (!x12020x) & (x12028x)) + ((!n_n1023) & (!n_n1061) & (!n_n1062) & (x12020x) & (!x12028x)) + ((!n_n1023) & (!n_n1061) & (!n_n1062) & (x12020x) & (x12028x)) + ((!n_n1023) & (!n_n1061) & (n_n1062) & (!x12020x) & (!x12028x)) + ((!n_n1023) & (!n_n1061) & (n_n1062) & (!x12020x) & (x12028x)) + ((!n_n1023) & (!n_n1061) & (n_n1062) & (x12020x) & (!x12028x)) + ((!n_n1023) & (!n_n1061) & (n_n1062) & (x12020x) & (x12028x)) + ((!n_n1023) & (n_n1061) & (!n_n1062) & (!x12020x) & (!x12028x)) + ((!n_n1023) & (n_n1061) & (!n_n1062) & (!x12020x) & (x12028x)) + ((!n_n1023) & (n_n1061) & (!n_n1062) & (x12020x) & (!x12028x)) + ((!n_n1023) & (n_n1061) & (!n_n1062) & (x12020x) & (x12028x)) + ((!n_n1023) & (n_n1061) & (n_n1062) & (!x12020x) & (!x12028x)) + ((!n_n1023) & (n_n1061) & (n_n1062) & (!x12020x) & (x12028x)) + ((!n_n1023) & (n_n1061) & (n_n1062) & (x12020x) & (!x12028x)) + ((!n_n1023) & (n_n1061) & (n_n1062) & (x12020x) & (x12028x)) + ((n_n1023) & (!n_n1061) & (!n_n1062) & (!x12020x) & (!x12028x)) + ((n_n1023) & (!n_n1061) & (!n_n1062) & (!x12020x) & (x12028x)) + ((n_n1023) & (!n_n1061) & (!n_n1062) & (x12020x) & (!x12028x)) + ((n_n1023) & (!n_n1061) & (!n_n1062) & (x12020x) & (x12028x)) + ((n_n1023) & (!n_n1061) & (n_n1062) & (!x12020x) & (!x12028x)) + ((n_n1023) & (!n_n1061) & (n_n1062) & (!x12020x) & (x12028x)) + ((n_n1023) & (!n_n1061) & (n_n1062) & (x12020x) & (!x12028x)) + ((n_n1023) & (!n_n1061) & (n_n1062) & (x12020x) & (x12028x)) + ((n_n1023) & (n_n1061) & (!n_n1062) & (!x12020x) & (!x12028x)) + ((n_n1023) & (n_n1061) & (!n_n1062) & (!x12020x) & (x12028x)) + ((n_n1023) & (n_n1061) & (!n_n1062) & (x12020x) & (!x12028x)) + ((n_n1023) & (n_n1061) & (!n_n1062) & (x12020x) & (x12028x)) + ((n_n1023) & (n_n1061) & (n_n1062) & (!x12020x) & (!x12028x)) + ((n_n1023) & (n_n1061) & (n_n1062) & (!x12020x) & (x12028x)) + ((n_n1023) & (n_n1061) & (n_n1062) & (x12020x) & (!x12028x)) + ((n_n1023) & (n_n1061) & (n_n1062) & (x12020x) & (x12028x)));
	assign x12041x = (((!n_n1015) & (!x11747x) & (!n_n942) & (n_n941)) + ((!n_n1015) & (!x11747x) & (n_n942) & (!n_n941)) + ((!n_n1015) & (!x11747x) & (n_n942) & (n_n941)) + ((!n_n1015) & (x11747x) & (!n_n942) & (!n_n941)) + ((!n_n1015) & (x11747x) & (!n_n942) & (n_n941)) + ((!n_n1015) & (x11747x) & (n_n942) & (!n_n941)) + ((!n_n1015) & (x11747x) & (n_n942) & (n_n941)) + ((n_n1015) & (!x11747x) & (!n_n942) & (!n_n941)) + ((n_n1015) & (!x11747x) & (!n_n942) & (n_n941)) + ((n_n1015) & (!x11747x) & (n_n942) & (!n_n941)) + ((n_n1015) & (!x11747x) & (n_n942) & (n_n941)) + ((n_n1015) & (x11747x) & (!n_n942) & (!n_n941)) + ((n_n1015) & (x11747x) & (!n_n942) & (n_n941)) + ((n_n1015) & (x11747x) & (n_n942) & (!n_n941)) + ((n_n1015) & (x11747x) & (n_n942) & (n_n941)));
	assign x12589x = (((!n_n1396) & (!n_n1397) & (!x12391x) & (!n_n1394) & (n_n1393)) + ((!n_n1396) & (!n_n1397) & (!x12391x) & (n_n1394) & (!n_n1393)) + ((!n_n1396) & (!n_n1397) & (!x12391x) & (n_n1394) & (n_n1393)) + ((!n_n1396) & (!n_n1397) & (x12391x) & (!n_n1394) & (!n_n1393)) + ((!n_n1396) & (!n_n1397) & (x12391x) & (!n_n1394) & (n_n1393)) + ((!n_n1396) & (!n_n1397) & (x12391x) & (n_n1394) & (!n_n1393)) + ((!n_n1396) & (!n_n1397) & (x12391x) & (n_n1394) & (n_n1393)) + ((!n_n1396) & (n_n1397) & (!x12391x) & (!n_n1394) & (!n_n1393)) + ((!n_n1396) & (n_n1397) & (!x12391x) & (!n_n1394) & (n_n1393)) + ((!n_n1396) & (n_n1397) & (!x12391x) & (n_n1394) & (!n_n1393)) + ((!n_n1396) & (n_n1397) & (!x12391x) & (n_n1394) & (n_n1393)) + ((!n_n1396) & (n_n1397) & (x12391x) & (!n_n1394) & (!n_n1393)) + ((!n_n1396) & (n_n1397) & (x12391x) & (!n_n1394) & (n_n1393)) + ((!n_n1396) & (n_n1397) & (x12391x) & (n_n1394) & (!n_n1393)) + ((!n_n1396) & (n_n1397) & (x12391x) & (n_n1394) & (n_n1393)) + ((n_n1396) & (!n_n1397) & (!x12391x) & (!n_n1394) & (!n_n1393)) + ((n_n1396) & (!n_n1397) & (!x12391x) & (!n_n1394) & (n_n1393)) + ((n_n1396) & (!n_n1397) & (!x12391x) & (n_n1394) & (!n_n1393)) + ((n_n1396) & (!n_n1397) & (!x12391x) & (n_n1394) & (n_n1393)) + ((n_n1396) & (!n_n1397) & (x12391x) & (!n_n1394) & (!n_n1393)) + ((n_n1396) & (!n_n1397) & (x12391x) & (!n_n1394) & (n_n1393)) + ((n_n1396) & (!n_n1397) & (x12391x) & (n_n1394) & (!n_n1393)) + ((n_n1396) & (!n_n1397) & (x12391x) & (n_n1394) & (n_n1393)) + ((n_n1396) & (n_n1397) & (!x12391x) & (!n_n1394) & (!n_n1393)) + ((n_n1396) & (n_n1397) & (!x12391x) & (!n_n1394) & (n_n1393)) + ((n_n1396) & (n_n1397) & (!x12391x) & (n_n1394) & (!n_n1393)) + ((n_n1396) & (n_n1397) & (!x12391x) & (n_n1394) & (n_n1393)) + ((n_n1396) & (n_n1397) & (x12391x) & (!n_n1394) & (!n_n1393)) + ((n_n1396) & (n_n1397) & (x12391x) & (!n_n1394) & (n_n1393)) + ((n_n1396) & (n_n1397) & (x12391x) & (n_n1394) & (!n_n1393)) + ((n_n1396) & (n_n1397) & (x12391x) & (n_n1394) & (n_n1393)));
	assign x12151x = (((!x12062x) & (!x12063x) & (!x12083x) & (x12084x)) + ((!x12062x) & (!x12063x) & (x12083x) & (!x12084x)) + ((!x12062x) & (!x12063x) & (x12083x) & (x12084x)) + ((!x12062x) & (x12063x) & (!x12083x) & (!x12084x)) + ((!x12062x) & (x12063x) & (!x12083x) & (x12084x)) + ((!x12062x) & (x12063x) & (x12083x) & (!x12084x)) + ((!x12062x) & (x12063x) & (x12083x) & (x12084x)) + ((x12062x) & (!x12063x) & (!x12083x) & (!x12084x)) + ((x12062x) & (!x12063x) & (!x12083x) & (x12084x)) + ((x12062x) & (!x12063x) & (x12083x) & (!x12084x)) + ((x12062x) & (!x12063x) & (x12083x) & (x12084x)) + ((x12062x) & (x12063x) & (!x12083x) & (!x12084x)) + ((x12062x) & (x12063x) & (!x12083x) & (x12084x)) + ((x12062x) & (x12063x) & (x12083x) & (!x12084x)) + ((x12062x) & (x12063x) & (x12083x) & (x12084x)));
	assign x12152x = (((!n_n1323) & (!x12129x) & (!x12130x) & (x12150x)) + ((!n_n1323) & (!x12129x) & (x12130x) & (!x12150x)) + ((!n_n1323) & (!x12129x) & (x12130x) & (x12150x)) + ((!n_n1323) & (x12129x) & (!x12130x) & (!x12150x)) + ((!n_n1323) & (x12129x) & (!x12130x) & (x12150x)) + ((!n_n1323) & (x12129x) & (x12130x) & (!x12150x)) + ((!n_n1323) & (x12129x) & (x12130x) & (x12150x)) + ((n_n1323) & (!x12129x) & (!x12130x) & (!x12150x)) + ((n_n1323) & (!x12129x) & (!x12130x) & (x12150x)) + ((n_n1323) & (!x12129x) & (x12130x) & (!x12150x)) + ((n_n1323) & (!x12129x) & (x12130x) & (x12150x)) + ((n_n1323) & (x12129x) & (!x12130x) & (!x12150x)) + ((n_n1323) & (x12129x) & (!x12130x) & (x12150x)) + ((n_n1323) & (x12129x) & (x12130x) & (!x12150x)) + ((n_n1323) & (x12129x) & (x12130x) & (x12150x)));
	assign n_n1398 = (((!x12440x) & (!n_n1480) & (!n_n1418) & (!x12431x) & (n_n1481)) + ((!x12440x) & (!n_n1480) & (!n_n1418) & (x12431x) & (!n_n1481)) + ((!x12440x) & (!n_n1480) & (!n_n1418) & (x12431x) & (n_n1481)) + ((!x12440x) & (!n_n1480) & (n_n1418) & (!x12431x) & (!n_n1481)) + ((!x12440x) & (!n_n1480) & (n_n1418) & (!x12431x) & (n_n1481)) + ((!x12440x) & (!n_n1480) & (n_n1418) & (x12431x) & (!n_n1481)) + ((!x12440x) & (!n_n1480) & (n_n1418) & (x12431x) & (n_n1481)) + ((!x12440x) & (n_n1480) & (!n_n1418) & (!x12431x) & (!n_n1481)) + ((!x12440x) & (n_n1480) & (!n_n1418) & (!x12431x) & (n_n1481)) + ((!x12440x) & (n_n1480) & (!n_n1418) & (x12431x) & (!n_n1481)) + ((!x12440x) & (n_n1480) & (!n_n1418) & (x12431x) & (n_n1481)) + ((!x12440x) & (n_n1480) & (n_n1418) & (!x12431x) & (!n_n1481)) + ((!x12440x) & (n_n1480) & (n_n1418) & (!x12431x) & (n_n1481)) + ((!x12440x) & (n_n1480) & (n_n1418) & (x12431x) & (!n_n1481)) + ((!x12440x) & (n_n1480) & (n_n1418) & (x12431x) & (n_n1481)) + ((x12440x) & (!n_n1480) & (!n_n1418) & (!x12431x) & (!n_n1481)) + ((x12440x) & (!n_n1480) & (!n_n1418) & (!x12431x) & (n_n1481)) + ((x12440x) & (!n_n1480) & (!n_n1418) & (x12431x) & (!n_n1481)) + ((x12440x) & (!n_n1480) & (!n_n1418) & (x12431x) & (n_n1481)) + ((x12440x) & (!n_n1480) & (n_n1418) & (!x12431x) & (!n_n1481)) + ((x12440x) & (!n_n1480) & (n_n1418) & (!x12431x) & (n_n1481)) + ((x12440x) & (!n_n1480) & (n_n1418) & (x12431x) & (!n_n1481)) + ((x12440x) & (!n_n1480) & (n_n1418) & (x12431x) & (n_n1481)) + ((x12440x) & (n_n1480) & (!n_n1418) & (!x12431x) & (!n_n1481)) + ((x12440x) & (n_n1480) & (!n_n1418) & (!x12431x) & (n_n1481)) + ((x12440x) & (n_n1480) & (!n_n1418) & (x12431x) & (!n_n1481)) + ((x12440x) & (n_n1480) & (!n_n1418) & (x12431x) & (n_n1481)) + ((x12440x) & (n_n1480) & (n_n1418) & (!x12431x) & (!n_n1481)) + ((x12440x) & (n_n1480) & (n_n1418) & (!x12431x) & (n_n1481)) + ((x12440x) & (n_n1480) & (n_n1418) & (x12431x) & (!n_n1481)) + ((x12440x) & (n_n1480) & (n_n1418) & (x12431x) & (n_n1481)));
	assign n_n1392 = (((!x12585x) & (!n_n1425) & (!n_n1423) & (!x12517x) & (n_n1399)) + ((!x12585x) & (!n_n1425) & (!n_n1423) & (x12517x) & (!n_n1399)) + ((!x12585x) & (!n_n1425) & (!n_n1423) & (x12517x) & (n_n1399)) + ((!x12585x) & (!n_n1425) & (n_n1423) & (!x12517x) & (!n_n1399)) + ((!x12585x) & (!n_n1425) & (n_n1423) & (!x12517x) & (n_n1399)) + ((!x12585x) & (!n_n1425) & (n_n1423) & (x12517x) & (!n_n1399)) + ((!x12585x) & (!n_n1425) & (n_n1423) & (x12517x) & (n_n1399)) + ((!x12585x) & (n_n1425) & (!n_n1423) & (!x12517x) & (!n_n1399)) + ((!x12585x) & (n_n1425) & (!n_n1423) & (!x12517x) & (n_n1399)) + ((!x12585x) & (n_n1425) & (!n_n1423) & (x12517x) & (!n_n1399)) + ((!x12585x) & (n_n1425) & (!n_n1423) & (x12517x) & (n_n1399)) + ((!x12585x) & (n_n1425) & (n_n1423) & (!x12517x) & (!n_n1399)) + ((!x12585x) & (n_n1425) & (n_n1423) & (!x12517x) & (n_n1399)) + ((!x12585x) & (n_n1425) & (n_n1423) & (x12517x) & (!n_n1399)) + ((!x12585x) & (n_n1425) & (n_n1423) & (x12517x) & (n_n1399)) + ((x12585x) & (!n_n1425) & (!n_n1423) & (!x12517x) & (!n_n1399)) + ((x12585x) & (!n_n1425) & (!n_n1423) & (!x12517x) & (n_n1399)) + ((x12585x) & (!n_n1425) & (!n_n1423) & (x12517x) & (!n_n1399)) + ((x12585x) & (!n_n1425) & (!n_n1423) & (x12517x) & (n_n1399)) + ((x12585x) & (!n_n1425) & (n_n1423) & (!x12517x) & (!n_n1399)) + ((x12585x) & (!n_n1425) & (n_n1423) & (!x12517x) & (n_n1399)) + ((x12585x) & (!n_n1425) & (n_n1423) & (x12517x) & (!n_n1399)) + ((x12585x) & (!n_n1425) & (n_n1423) & (x12517x) & (n_n1399)) + ((x12585x) & (n_n1425) & (!n_n1423) & (!x12517x) & (!n_n1399)) + ((x12585x) & (n_n1425) & (!n_n1423) & (!x12517x) & (n_n1399)) + ((x12585x) & (n_n1425) & (!n_n1423) & (x12517x) & (!n_n1399)) + ((x12585x) & (n_n1425) & (!n_n1423) & (x12517x) & (n_n1399)) + ((x12585x) & (n_n1425) & (n_n1423) & (!x12517x) & (!n_n1399)) + ((x12585x) & (n_n1425) & (n_n1423) & (!x12517x) & (n_n1399)) + ((x12585x) & (n_n1425) & (n_n1423) & (x12517x) & (!n_n1399)) + ((x12585x) & (n_n1425) & (n_n1423) & (x12517x) & (n_n1399)));
	assign x13147x = (((!x12693x) & (!n_n539) & (!n_n540) & (x13146x)) + ((!x12693x) & (!n_n539) & (n_n540) & (!x13146x)) + ((!x12693x) & (!n_n539) & (n_n540) & (x13146x)) + ((!x12693x) & (n_n539) & (!n_n540) & (!x13146x)) + ((!x12693x) & (n_n539) & (!n_n540) & (x13146x)) + ((!x12693x) & (n_n539) & (n_n540) & (!x13146x)) + ((!x12693x) & (n_n539) & (n_n540) & (x13146x)) + ((x12693x) & (!n_n539) & (!n_n540) & (!x13146x)) + ((x12693x) & (!n_n539) & (!n_n540) & (x13146x)) + ((x12693x) & (!n_n539) & (n_n540) & (!x13146x)) + ((x12693x) & (!n_n539) & (n_n540) & (x13146x)) + ((x12693x) & (n_n539) & (!n_n540) & (!x13146x)) + ((x12693x) & (n_n539) & (!n_n540) & (x13146x)) + ((x12693x) & (n_n539) & (n_n540) & (!x13146x)) + ((x12693x) & (n_n539) & (n_n540) & (x13146x)));
	assign x13136x = (((!n_n630) & (!n_n657) & (!n_n656) & (!x13088x) & (n_n629)) + ((!n_n630) & (!n_n657) & (!n_n656) & (x13088x) & (!n_n629)) + ((!n_n630) & (!n_n657) & (!n_n656) & (x13088x) & (n_n629)) + ((!n_n630) & (!n_n657) & (n_n656) & (!x13088x) & (!n_n629)) + ((!n_n630) & (!n_n657) & (n_n656) & (!x13088x) & (n_n629)) + ((!n_n630) & (!n_n657) & (n_n656) & (x13088x) & (!n_n629)) + ((!n_n630) & (!n_n657) & (n_n656) & (x13088x) & (n_n629)) + ((!n_n630) & (n_n657) & (!n_n656) & (!x13088x) & (!n_n629)) + ((!n_n630) & (n_n657) & (!n_n656) & (!x13088x) & (n_n629)) + ((!n_n630) & (n_n657) & (!n_n656) & (x13088x) & (!n_n629)) + ((!n_n630) & (n_n657) & (!n_n656) & (x13088x) & (n_n629)) + ((!n_n630) & (n_n657) & (n_n656) & (!x13088x) & (!n_n629)) + ((!n_n630) & (n_n657) & (n_n656) & (!x13088x) & (n_n629)) + ((!n_n630) & (n_n657) & (n_n656) & (x13088x) & (!n_n629)) + ((!n_n630) & (n_n657) & (n_n656) & (x13088x) & (n_n629)) + ((n_n630) & (!n_n657) & (!n_n656) & (!x13088x) & (!n_n629)) + ((n_n630) & (!n_n657) & (!n_n656) & (!x13088x) & (n_n629)) + ((n_n630) & (!n_n657) & (!n_n656) & (x13088x) & (!n_n629)) + ((n_n630) & (!n_n657) & (!n_n656) & (x13088x) & (n_n629)) + ((n_n630) & (!n_n657) & (n_n656) & (!x13088x) & (!n_n629)) + ((n_n630) & (!n_n657) & (n_n656) & (!x13088x) & (n_n629)) + ((n_n630) & (!n_n657) & (n_n656) & (x13088x) & (!n_n629)) + ((n_n630) & (!n_n657) & (n_n656) & (x13088x) & (n_n629)) + ((n_n630) & (n_n657) & (!n_n656) & (!x13088x) & (!n_n629)) + ((n_n630) & (n_n657) & (!n_n656) & (!x13088x) & (n_n629)) + ((n_n630) & (n_n657) & (!n_n656) & (x13088x) & (!n_n629)) + ((n_n630) & (n_n657) & (!n_n656) & (x13088x) & (n_n629)) + ((n_n630) & (n_n657) & (n_n656) & (!x13088x) & (!n_n629)) + ((n_n630) & (n_n657) & (n_n656) & (!x13088x) & (n_n629)) + ((n_n630) & (n_n657) & (n_n656) & (x13088x) & (!n_n629)) + ((n_n630) & (n_n657) & (n_n656) & (x13088x) & (n_n629)));
	assign x13137x = (((!n_n627) & (!n_n628) & (!x12867x) & (!x13001x) & (x13002x)) + ((!n_n627) & (!n_n628) & (!x12867x) & (x13001x) & (!x13002x)) + ((!n_n627) & (!n_n628) & (!x12867x) & (x13001x) & (x13002x)) + ((!n_n627) & (!n_n628) & (x12867x) & (!x13001x) & (!x13002x)) + ((!n_n627) & (!n_n628) & (x12867x) & (!x13001x) & (x13002x)) + ((!n_n627) & (!n_n628) & (x12867x) & (x13001x) & (!x13002x)) + ((!n_n627) & (!n_n628) & (x12867x) & (x13001x) & (x13002x)) + ((!n_n627) & (n_n628) & (!x12867x) & (!x13001x) & (!x13002x)) + ((!n_n627) & (n_n628) & (!x12867x) & (!x13001x) & (x13002x)) + ((!n_n627) & (n_n628) & (!x12867x) & (x13001x) & (!x13002x)) + ((!n_n627) & (n_n628) & (!x12867x) & (x13001x) & (x13002x)) + ((!n_n627) & (n_n628) & (x12867x) & (!x13001x) & (!x13002x)) + ((!n_n627) & (n_n628) & (x12867x) & (!x13001x) & (x13002x)) + ((!n_n627) & (n_n628) & (x12867x) & (x13001x) & (!x13002x)) + ((!n_n627) & (n_n628) & (x12867x) & (x13001x) & (x13002x)) + ((n_n627) & (!n_n628) & (!x12867x) & (!x13001x) & (!x13002x)) + ((n_n627) & (!n_n628) & (!x12867x) & (!x13001x) & (x13002x)) + ((n_n627) & (!n_n628) & (!x12867x) & (x13001x) & (!x13002x)) + ((n_n627) & (!n_n628) & (!x12867x) & (x13001x) & (x13002x)) + ((n_n627) & (!n_n628) & (x12867x) & (!x13001x) & (!x13002x)) + ((n_n627) & (!n_n628) & (x12867x) & (!x13001x) & (x13002x)) + ((n_n627) & (!n_n628) & (x12867x) & (x13001x) & (!x13002x)) + ((n_n627) & (!n_n628) & (x12867x) & (x13001x) & (x13002x)) + ((n_n627) & (n_n628) & (!x12867x) & (!x13001x) & (!x13002x)) + ((n_n627) & (n_n628) & (!x12867x) & (!x13001x) & (x13002x)) + ((n_n627) & (n_n628) & (!x12867x) & (x13001x) & (!x13002x)) + ((n_n627) & (n_n628) & (!x12867x) & (x13001x) & (x13002x)) + ((n_n627) & (n_n628) & (x12867x) & (!x13001x) & (!x13002x)) + ((n_n627) & (n_n628) & (x12867x) & (!x13001x) & (x13002x)) + ((n_n627) & (n_n628) & (x12867x) & (x13001x) & (!x13002x)) + ((n_n627) & (n_n628) & (x12867x) & (x13001x) & (x13002x)));
	assign x13684x = (((!x13645x) & (!x13646x) & (!n_n3921) & (x13683x)) + ((!x13645x) & (!x13646x) & (n_n3921) & (!x13683x)) + ((!x13645x) & (!x13646x) & (n_n3921) & (x13683x)) + ((!x13645x) & (x13646x) & (!n_n3921) & (!x13683x)) + ((!x13645x) & (x13646x) & (!n_n3921) & (x13683x)) + ((!x13645x) & (x13646x) & (n_n3921) & (!x13683x)) + ((!x13645x) & (x13646x) & (n_n3921) & (x13683x)) + ((x13645x) & (!x13646x) & (!n_n3921) & (!x13683x)) + ((x13645x) & (!x13646x) & (!n_n3921) & (x13683x)) + ((x13645x) & (!x13646x) & (n_n3921) & (!x13683x)) + ((x13645x) & (!x13646x) & (n_n3921) & (x13683x)) + ((x13645x) & (x13646x) & (!n_n3921) & (!x13683x)) + ((x13645x) & (x13646x) & (!n_n3921) & (x13683x)) + ((x13645x) & (x13646x) & (n_n3921) & (!x13683x)) + ((x13645x) & (x13646x) & (n_n3921) & (x13683x)));
	assign x13573x = (((!n_n3990) & (!n_n3992) & (!n_n3988) & (n_n3987)) + ((!n_n3990) & (!n_n3992) & (n_n3988) & (!n_n3987)) + ((!n_n3990) & (!n_n3992) & (n_n3988) & (n_n3987)) + ((!n_n3990) & (n_n3992) & (!n_n3988) & (!n_n3987)) + ((!n_n3990) & (n_n3992) & (!n_n3988) & (n_n3987)) + ((!n_n3990) & (n_n3992) & (n_n3988) & (!n_n3987)) + ((!n_n3990) & (n_n3992) & (n_n3988) & (n_n3987)) + ((n_n3990) & (!n_n3992) & (!n_n3988) & (!n_n3987)) + ((n_n3990) & (!n_n3992) & (!n_n3988) & (n_n3987)) + ((n_n3990) & (!n_n3992) & (n_n3988) & (!n_n3987)) + ((n_n3990) & (!n_n3992) & (n_n3988) & (n_n3987)) + ((n_n3990) & (n_n3992) & (!n_n3988) & (!n_n3987)) + ((n_n3990) & (n_n3992) & (!n_n3988) & (n_n3987)) + ((n_n3990) & (n_n3992) & (n_n3988) & (!n_n3987)) + ((n_n3990) & (n_n3992) & (n_n3988) & (n_n3987)));
	assign x13574x = (((!n_n3989) & (!n_n3993) & (!n_n3995) & (!x13555x) & (x13569x)) + ((!n_n3989) & (!n_n3993) & (!n_n3995) & (x13555x) & (!x13569x)) + ((!n_n3989) & (!n_n3993) & (!n_n3995) & (x13555x) & (x13569x)) + ((!n_n3989) & (!n_n3993) & (n_n3995) & (!x13555x) & (!x13569x)) + ((!n_n3989) & (!n_n3993) & (n_n3995) & (!x13555x) & (x13569x)) + ((!n_n3989) & (!n_n3993) & (n_n3995) & (x13555x) & (!x13569x)) + ((!n_n3989) & (!n_n3993) & (n_n3995) & (x13555x) & (x13569x)) + ((!n_n3989) & (n_n3993) & (!n_n3995) & (!x13555x) & (!x13569x)) + ((!n_n3989) & (n_n3993) & (!n_n3995) & (!x13555x) & (x13569x)) + ((!n_n3989) & (n_n3993) & (!n_n3995) & (x13555x) & (!x13569x)) + ((!n_n3989) & (n_n3993) & (!n_n3995) & (x13555x) & (x13569x)) + ((!n_n3989) & (n_n3993) & (n_n3995) & (!x13555x) & (!x13569x)) + ((!n_n3989) & (n_n3993) & (n_n3995) & (!x13555x) & (x13569x)) + ((!n_n3989) & (n_n3993) & (n_n3995) & (x13555x) & (!x13569x)) + ((!n_n3989) & (n_n3993) & (n_n3995) & (x13555x) & (x13569x)) + ((n_n3989) & (!n_n3993) & (!n_n3995) & (!x13555x) & (!x13569x)) + ((n_n3989) & (!n_n3993) & (!n_n3995) & (!x13555x) & (x13569x)) + ((n_n3989) & (!n_n3993) & (!n_n3995) & (x13555x) & (!x13569x)) + ((n_n3989) & (!n_n3993) & (!n_n3995) & (x13555x) & (x13569x)) + ((n_n3989) & (!n_n3993) & (n_n3995) & (!x13555x) & (!x13569x)) + ((n_n3989) & (!n_n3993) & (n_n3995) & (!x13555x) & (x13569x)) + ((n_n3989) & (!n_n3993) & (n_n3995) & (x13555x) & (!x13569x)) + ((n_n3989) & (!n_n3993) & (n_n3995) & (x13555x) & (x13569x)) + ((n_n3989) & (n_n3993) & (!n_n3995) & (!x13555x) & (!x13569x)) + ((n_n3989) & (n_n3993) & (!n_n3995) & (!x13555x) & (x13569x)) + ((n_n3989) & (n_n3993) & (!n_n3995) & (x13555x) & (!x13569x)) + ((n_n3989) & (n_n3993) & (!n_n3995) & (x13555x) & (x13569x)) + ((n_n3989) & (n_n3993) & (n_n3995) & (!x13555x) & (!x13569x)) + ((n_n3989) & (n_n3993) & (n_n3995) & (!x13555x) & (x13569x)) + ((n_n3989) & (n_n3993) & (n_n3995) & (x13555x) & (!x13569x)) + ((n_n3989) & (n_n3993) & (n_n3995) & (x13555x) & (x13569x)));
	assign x14222x = (((!n_n3192) & (!x13782x) & (!x13783x) & (x14221x)) + ((!n_n3192) & (!x13782x) & (x13783x) & (!x14221x)) + ((!n_n3192) & (!x13782x) & (x13783x) & (x14221x)) + ((!n_n3192) & (x13782x) & (!x13783x) & (!x14221x)) + ((!n_n3192) & (x13782x) & (!x13783x) & (x14221x)) + ((!n_n3192) & (x13782x) & (x13783x) & (!x14221x)) + ((!n_n3192) & (x13782x) & (x13783x) & (x14221x)) + ((n_n3192) & (!x13782x) & (!x13783x) & (!x14221x)) + ((n_n3192) & (!x13782x) & (!x13783x) & (x14221x)) + ((n_n3192) & (!x13782x) & (x13783x) & (!x14221x)) + ((n_n3192) & (!x13782x) & (x13783x) & (x14221x)) + ((n_n3192) & (x13782x) & (!x13783x) & (!x14221x)) + ((n_n3192) & (x13782x) & (!x13783x) & (x14221x)) + ((n_n3192) & (x13782x) & (x13783x) & (!x14221x)) + ((n_n3192) & (x13782x) & (x13783x) & (x14221x)));
	assign x14216x = (((!n_n3257) & (!n_n3259) & (x14214x)) + ((!n_n3257) & (n_n3259) & (!x14214x)) + ((!n_n3257) & (n_n3259) & (x14214x)) + ((n_n3257) & (!n_n3259) & (!x14214x)) + ((n_n3257) & (!n_n3259) & (x14214x)) + ((n_n3257) & (n_n3259) & (!x14214x)) + ((n_n3257) & (n_n3259) & (x14214x)));
	assign n_n3251 = (((!n_n3254) & (!n_n3256) & (x14067x)) + ((!n_n3254) & (n_n3256) & (!x14067x)) + ((!n_n3254) & (n_n3256) & (x14067x)) + ((n_n3254) & (!n_n3256) & (!x14067x)) + ((n_n3254) & (!n_n3256) & (x14067x)) + ((n_n3254) & (n_n3256) & (!x14067x)) + ((n_n3254) & (n_n3256) & (x14067x)));
	assign n_n3253 = (((!n_n3260) & (!n_n3262) & (x14211x)) + ((!n_n3260) & (n_n3262) & (!x14211x)) + ((!n_n3260) & (n_n3262) & (x14211x)) + ((n_n3260) & (!n_n3262) & (!x14211x)) + ((n_n3260) & (!n_n3262) & (x14211x)) + ((n_n3260) & (n_n3262) & (!x14211x)) + ((n_n3260) & (n_n3262) & (x14211x)));
	assign x14780x = (((!x14540x) & (!n_n3625) & (!n_n3627) & (!n_n3629) & (n_n3631)) + ((!x14540x) & (!n_n3625) & (!n_n3627) & (n_n3629) & (!n_n3631)) + ((!x14540x) & (!n_n3625) & (!n_n3627) & (n_n3629) & (n_n3631)) + ((!x14540x) & (!n_n3625) & (n_n3627) & (!n_n3629) & (!n_n3631)) + ((!x14540x) & (!n_n3625) & (n_n3627) & (!n_n3629) & (n_n3631)) + ((!x14540x) & (!n_n3625) & (n_n3627) & (n_n3629) & (!n_n3631)) + ((!x14540x) & (!n_n3625) & (n_n3627) & (n_n3629) & (n_n3631)) + ((!x14540x) & (n_n3625) & (!n_n3627) & (!n_n3629) & (!n_n3631)) + ((!x14540x) & (n_n3625) & (!n_n3627) & (!n_n3629) & (n_n3631)) + ((!x14540x) & (n_n3625) & (!n_n3627) & (n_n3629) & (!n_n3631)) + ((!x14540x) & (n_n3625) & (!n_n3627) & (n_n3629) & (n_n3631)) + ((!x14540x) & (n_n3625) & (n_n3627) & (!n_n3629) & (!n_n3631)) + ((!x14540x) & (n_n3625) & (n_n3627) & (!n_n3629) & (n_n3631)) + ((!x14540x) & (n_n3625) & (n_n3627) & (n_n3629) & (!n_n3631)) + ((!x14540x) & (n_n3625) & (n_n3627) & (n_n3629) & (n_n3631)) + ((x14540x) & (!n_n3625) & (!n_n3627) & (!n_n3629) & (!n_n3631)) + ((x14540x) & (!n_n3625) & (!n_n3627) & (!n_n3629) & (n_n3631)) + ((x14540x) & (!n_n3625) & (!n_n3627) & (n_n3629) & (!n_n3631)) + ((x14540x) & (!n_n3625) & (!n_n3627) & (n_n3629) & (n_n3631)) + ((x14540x) & (!n_n3625) & (n_n3627) & (!n_n3629) & (!n_n3631)) + ((x14540x) & (!n_n3625) & (n_n3627) & (!n_n3629) & (n_n3631)) + ((x14540x) & (!n_n3625) & (n_n3627) & (n_n3629) & (!n_n3631)) + ((x14540x) & (!n_n3625) & (n_n3627) & (n_n3629) & (n_n3631)) + ((x14540x) & (n_n3625) & (!n_n3627) & (!n_n3629) & (!n_n3631)) + ((x14540x) & (n_n3625) & (!n_n3627) & (!n_n3629) & (n_n3631)) + ((x14540x) & (n_n3625) & (!n_n3627) & (n_n3629) & (!n_n3631)) + ((x14540x) & (n_n3625) & (!n_n3627) & (n_n3629) & (n_n3631)) + ((x14540x) & (n_n3625) & (n_n3627) & (!n_n3629) & (!n_n3631)) + ((x14540x) & (n_n3625) & (n_n3627) & (!n_n3629) & (n_n3631)) + ((x14540x) & (n_n3625) & (n_n3627) & (n_n3629) & (!n_n3631)) + ((x14540x) & (n_n3625) & (n_n3627) & (n_n3629) & (n_n3631)));
	assign n_n3623 = (((!x14591x) & (!n_n3661) & (!n_n3660) & (!x14566x) & (n_n3634)) + ((!x14591x) & (!n_n3661) & (!n_n3660) & (x14566x) & (!n_n3634)) + ((!x14591x) & (!n_n3661) & (!n_n3660) & (x14566x) & (n_n3634)) + ((!x14591x) & (!n_n3661) & (n_n3660) & (!x14566x) & (!n_n3634)) + ((!x14591x) & (!n_n3661) & (n_n3660) & (!x14566x) & (n_n3634)) + ((!x14591x) & (!n_n3661) & (n_n3660) & (x14566x) & (!n_n3634)) + ((!x14591x) & (!n_n3661) & (n_n3660) & (x14566x) & (n_n3634)) + ((!x14591x) & (n_n3661) & (!n_n3660) & (!x14566x) & (!n_n3634)) + ((!x14591x) & (n_n3661) & (!n_n3660) & (!x14566x) & (n_n3634)) + ((!x14591x) & (n_n3661) & (!n_n3660) & (x14566x) & (!n_n3634)) + ((!x14591x) & (n_n3661) & (!n_n3660) & (x14566x) & (n_n3634)) + ((!x14591x) & (n_n3661) & (n_n3660) & (!x14566x) & (!n_n3634)) + ((!x14591x) & (n_n3661) & (n_n3660) & (!x14566x) & (n_n3634)) + ((!x14591x) & (n_n3661) & (n_n3660) & (x14566x) & (!n_n3634)) + ((!x14591x) & (n_n3661) & (n_n3660) & (x14566x) & (n_n3634)) + ((x14591x) & (!n_n3661) & (!n_n3660) & (!x14566x) & (!n_n3634)) + ((x14591x) & (!n_n3661) & (!n_n3660) & (!x14566x) & (n_n3634)) + ((x14591x) & (!n_n3661) & (!n_n3660) & (x14566x) & (!n_n3634)) + ((x14591x) & (!n_n3661) & (!n_n3660) & (x14566x) & (n_n3634)) + ((x14591x) & (!n_n3661) & (n_n3660) & (!x14566x) & (!n_n3634)) + ((x14591x) & (!n_n3661) & (n_n3660) & (!x14566x) & (n_n3634)) + ((x14591x) & (!n_n3661) & (n_n3660) & (x14566x) & (!n_n3634)) + ((x14591x) & (!n_n3661) & (n_n3660) & (x14566x) & (n_n3634)) + ((x14591x) & (n_n3661) & (!n_n3660) & (!x14566x) & (!n_n3634)) + ((x14591x) & (n_n3661) & (!n_n3660) & (!x14566x) & (n_n3634)) + ((x14591x) & (n_n3661) & (!n_n3660) & (x14566x) & (!n_n3634)) + ((x14591x) & (n_n3661) & (!n_n3660) & (x14566x) & (n_n3634)) + ((x14591x) & (n_n3661) & (n_n3660) & (!x14566x) & (!n_n3634)) + ((x14591x) & (n_n3661) & (n_n3660) & (!x14566x) & (n_n3634)) + ((x14591x) & (n_n3661) & (n_n3660) & (x14566x) & (!n_n3634)) + ((x14591x) & (n_n3661) & (n_n3660) & (x14566x) & (n_n3634)));
	assign n_n3624 = (((!x14638x) & (!x14613x) & (!n_n3635) & (!n_n3676) & (x14612x)) + ((!x14638x) & (!x14613x) & (!n_n3635) & (n_n3676) & (!x14612x)) + ((!x14638x) & (!x14613x) & (!n_n3635) & (n_n3676) & (x14612x)) + ((!x14638x) & (!x14613x) & (n_n3635) & (!n_n3676) & (!x14612x)) + ((!x14638x) & (!x14613x) & (n_n3635) & (!n_n3676) & (x14612x)) + ((!x14638x) & (!x14613x) & (n_n3635) & (n_n3676) & (!x14612x)) + ((!x14638x) & (!x14613x) & (n_n3635) & (n_n3676) & (x14612x)) + ((!x14638x) & (x14613x) & (!n_n3635) & (!n_n3676) & (!x14612x)) + ((!x14638x) & (x14613x) & (!n_n3635) & (!n_n3676) & (x14612x)) + ((!x14638x) & (x14613x) & (!n_n3635) & (n_n3676) & (!x14612x)) + ((!x14638x) & (x14613x) & (!n_n3635) & (n_n3676) & (x14612x)) + ((!x14638x) & (x14613x) & (n_n3635) & (!n_n3676) & (!x14612x)) + ((!x14638x) & (x14613x) & (n_n3635) & (!n_n3676) & (x14612x)) + ((!x14638x) & (x14613x) & (n_n3635) & (n_n3676) & (!x14612x)) + ((!x14638x) & (x14613x) & (n_n3635) & (n_n3676) & (x14612x)) + ((x14638x) & (!x14613x) & (!n_n3635) & (!n_n3676) & (!x14612x)) + ((x14638x) & (!x14613x) & (!n_n3635) & (!n_n3676) & (x14612x)) + ((x14638x) & (!x14613x) & (!n_n3635) & (n_n3676) & (!x14612x)) + ((x14638x) & (!x14613x) & (!n_n3635) & (n_n3676) & (x14612x)) + ((x14638x) & (!x14613x) & (n_n3635) & (!n_n3676) & (!x14612x)) + ((x14638x) & (!x14613x) & (n_n3635) & (!n_n3676) & (x14612x)) + ((x14638x) & (!x14613x) & (n_n3635) & (n_n3676) & (!x14612x)) + ((x14638x) & (!x14613x) & (n_n3635) & (n_n3676) & (x14612x)) + ((x14638x) & (x14613x) & (!n_n3635) & (!n_n3676) & (!x14612x)) + ((x14638x) & (x14613x) & (!n_n3635) & (!n_n3676) & (x14612x)) + ((x14638x) & (x14613x) & (!n_n3635) & (n_n3676) & (!x14612x)) + ((x14638x) & (x14613x) & (!n_n3635) & (n_n3676) & (x14612x)) + ((x14638x) & (x14613x) & (n_n3635) & (!n_n3676) & (!x14612x)) + ((x14638x) & (x14613x) & (n_n3635) & (!n_n3676) & (x14612x)) + ((x14638x) & (x14613x) & (n_n3635) & (n_n3676) & (!x14612x)) + ((x14638x) & (x14613x) & (n_n3635) & (n_n3676) & (x14612x)));
	assign x14775x = (((!x14388x) & (!n_n659) & (!n_n3649) & (!x22190x)) + ((!x14388x) & (!n_n659) & (n_n3649) & (!x22190x)) + ((!x14388x) & (!n_n659) & (n_n3649) & (x22190x)) + ((!x14388x) & (n_n659) & (!n_n3649) & (!x22190x)) + ((!x14388x) & (n_n659) & (!n_n3649) & (x22190x)) + ((!x14388x) & (n_n659) & (n_n3649) & (!x22190x)) + ((!x14388x) & (n_n659) & (n_n3649) & (x22190x)) + ((x14388x) & (!n_n659) & (!n_n3649) & (!x22190x)) + ((x14388x) & (!n_n659) & (!n_n3649) & (x22190x)) + ((x14388x) & (!n_n659) & (n_n3649) & (!x22190x)) + ((x14388x) & (!n_n659) & (n_n3649) & (x22190x)) + ((x14388x) & (n_n659) & (!n_n3649) & (!x22190x)) + ((x14388x) & (n_n659) & (!n_n3649) & (x22190x)) + ((x14388x) & (n_n659) & (n_n3649) & (!x22190x)) + ((x14388x) & (n_n659) & (n_n3649) & (x22190x)));
	assign x14778x = (((!n_n3543) & (!x14343x) & (n_n3626)) + ((!n_n3543) & (x14343x) & (!n_n3626)) + ((!n_n3543) & (x14343x) & (n_n3626)) + ((n_n3543) & (!x14343x) & (!n_n3626)) + ((n_n3543) & (!x14343x) & (n_n3626)) + ((n_n3543) & (x14343x) & (!n_n3626)) + ((n_n3543) & (x14343x) & (n_n3626)));
	assign x15301x = (((!n_n2530) & (!n_n2529) & (!x15169x) & (!n_n2533) & (n_n2532)) + ((!n_n2530) & (!n_n2529) & (!x15169x) & (n_n2533) & (!n_n2532)) + ((!n_n2530) & (!n_n2529) & (!x15169x) & (n_n2533) & (n_n2532)) + ((!n_n2530) & (!n_n2529) & (x15169x) & (!n_n2533) & (!n_n2532)) + ((!n_n2530) & (!n_n2529) & (x15169x) & (!n_n2533) & (n_n2532)) + ((!n_n2530) & (!n_n2529) & (x15169x) & (n_n2533) & (!n_n2532)) + ((!n_n2530) & (!n_n2529) & (x15169x) & (n_n2533) & (n_n2532)) + ((!n_n2530) & (n_n2529) & (!x15169x) & (!n_n2533) & (!n_n2532)) + ((!n_n2530) & (n_n2529) & (!x15169x) & (!n_n2533) & (n_n2532)) + ((!n_n2530) & (n_n2529) & (!x15169x) & (n_n2533) & (!n_n2532)) + ((!n_n2530) & (n_n2529) & (!x15169x) & (n_n2533) & (n_n2532)) + ((!n_n2530) & (n_n2529) & (x15169x) & (!n_n2533) & (!n_n2532)) + ((!n_n2530) & (n_n2529) & (x15169x) & (!n_n2533) & (n_n2532)) + ((!n_n2530) & (n_n2529) & (x15169x) & (n_n2533) & (!n_n2532)) + ((!n_n2530) & (n_n2529) & (x15169x) & (n_n2533) & (n_n2532)) + ((n_n2530) & (!n_n2529) & (!x15169x) & (!n_n2533) & (!n_n2532)) + ((n_n2530) & (!n_n2529) & (!x15169x) & (!n_n2533) & (n_n2532)) + ((n_n2530) & (!n_n2529) & (!x15169x) & (n_n2533) & (!n_n2532)) + ((n_n2530) & (!n_n2529) & (!x15169x) & (n_n2533) & (n_n2532)) + ((n_n2530) & (!n_n2529) & (x15169x) & (!n_n2533) & (!n_n2532)) + ((n_n2530) & (!n_n2529) & (x15169x) & (!n_n2533) & (n_n2532)) + ((n_n2530) & (!n_n2529) & (x15169x) & (n_n2533) & (!n_n2532)) + ((n_n2530) & (!n_n2529) & (x15169x) & (n_n2533) & (n_n2532)) + ((n_n2530) & (n_n2529) & (!x15169x) & (!n_n2533) & (!n_n2532)) + ((n_n2530) & (n_n2529) & (!x15169x) & (!n_n2533) & (n_n2532)) + ((n_n2530) & (n_n2529) & (!x15169x) & (n_n2533) & (!n_n2532)) + ((n_n2530) & (n_n2529) & (!x15169x) & (n_n2533) & (n_n2532)) + ((n_n2530) & (n_n2529) & (x15169x) & (!n_n2533) & (!n_n2532)) + ((n_n2530) & (n_n2529) & (x15169x) & (!n_n2533) & (n_n2532)) + ((n_n2530) & (n_n2529) & (x15169x) & (n_n2533) & (!n_n2532)) + ((n_n2530) & (n_n2529) & (x15169x) & (n_n2533) & (n_n2532)));
	assign n_n2523 = (((!x15297x) & (!n_n2526) & (!n_n2542) & (!n_n2541) & (x15264x)) + ((!x15297x) & (!n_n2526) & (!n_n2542) & (n_n2541) & (!x15264x)) + ((!x15297x) & (!n_n2526) & (!n_n2542) & (n_n2541) & (x15264x)) + ((!x15297x) & (!n_n2526) & (n_n2542) & (!n_n2541) & (!x15264x)) + ((!x15297x) & (!n_n2526) & (n_n2542) & (!n_n2541) & (x15264x)) + ((!x15297x) & (!n_n2526) & (n_n2542) & (n_n2541) & (!x15264x)) + ((!x15297x) & (!n_n2526) & (n_n2542) & (n_n2541) & (x15264x)) + ((!x15297x) & (n_n2526) & (!n_n2542) & (!n_n2541) & (!x15264x)) + ((!x15297x) & (n_n2526) & (!n_n2542) & (!n_n2541) & (x15264x)) + ((!x15297x) & (n_n2526) & (!n_n2542) & (n_n2541) & (!x15264x)) + ((!x15297x) & (n_n2526) & (!n_n2542) & (n_n2541) & (x15264x)) + ((!x15297x) & (n_n2526) & (n_n2542) & (!n_n2541) & (!x15264x)) + ((!x15297x) & (n_n2526) & (n_n2542) & (!n_n2541) & (x15264x)) + ((!x15297x) & (n_n2526) & (n_n2542) & (n_n2541) & (!x15264x)) + ((!x15297x) & (n_n2526) & (n_n2542) & (n_n2541) & (x15264x)) + ((x15297x) & (!n_n2526) & (!n_n2542) & (!n_n2541) & (!x15264x)) + ((x15297x) & (!n_n2526) & (!n_n2542) & (!n_n2541) & (x15264x)) + ((x15297x) & (!n_n2526) & (!n_n2542) & (n_n2541) & (!x15264x)) + ((x15297x) & (!n_n2526) & (!n_n2542) & (n_n2541) & (x15264x)) + ((x15297x) & (!n_n2526) & (n_n2542) & (!n_n2541) & (!x15264x)) + ((x15297x) & (!n_n2526) & (n_n2542) & (!n_n2541) & (x15264x)) + ((x15297x) & (!n_n2526) & (n_n2542) & (n_n2541) & (!x15264x)) + ((x15297x) & (!n_n2526) & (n_n2542) & (n_n2541) & (x15264x)) + ((x15297x) & (n_n2526) & (!n_n2542) & (!n_n2541) & (!x15264x)) + ((x15297x) & (n_n2526) & (!n_n2542) & (!n_n2541) & (x15264x)) + ((x15297x) & (n_n2526) & (!n_n2542) & (n_n2541) & (!x15264x)) + ((x15297x) & (n_n2526) & (!n_n2542) & (n_n2541) & (x15264x)) + ((x15297x) & (n_n2526) & (n_n2542) & (!n_n2541) & (!x15264x)) + ((x15297x) & (n_n2526) & (n_n2542) & (!n_n2541) & (x15264x)) + ((x15297x) & (n_n2526) & (n_n2542) & (n_n2541) & (!x15264x)) + ((x15297x) & (n_n2526) & (n_n2542) & (n_n2541) & (x15264x)));
	assign x15300x = (((!n_n2449) & (!n_n2531) & (!x14890x) & (x14891x)) + ((!n_n2449) & (!n_n2531) & (x14890x) & (!x14891x)) + ((!n_n2449) & (!n_n2531) & (x14890x) & (x14891x)) + ((!n_n2449) & (n_n2531) & (!x14890x) & (!x14891x)) + ((!n_n2449) & (n_n2531) & (!x14890x) & (x14891x)) + ((!n_n2449) & (n_n2531) & (x14890x) & (!x14891x)) + ((!n_n2449) & (n_n2531) & (x14890x) & (x14891x)) + ((n_n2449) & (!n_n2531) & (!x14890x) & (!x14891x)) + ((n_n2449) & (!n_n2531) & (!x14890x) & (x14891x)) + ((n_n2449) & (!n_n2531) & (x14890x) & (!x14891x)) + ((n_n2449) & (!n_n2531) & (x14890x) & (x14891x)) + ((n_n2449) & (n_n2531) & (!x14890x) & (!x14891x)) + ((n_n2449) & (n_n2531) & (!x14890x) & (x14891x)) + ((n_n2449) & (n_n2531) & (x14890x) & (!x14891x)) + ((n_n2449) & (n_n2531) & (x14890x) & (x14891x)));
	assign x15817x = (((!n_n2906) & (!n_n2908) & (!n_n2902) & (x15677x)) + ((!n_n2906) & (!n_n2908) & (n_n2902) & (!x15677x)) + ((!n_n2906) & (!n_n2908) & (n_n2902) & (x15677x)) + ((!n_n2906) & (n_n2908) & (!n_n2902) & (!x15677x)) + ((!n_n2906) & (n_n2908) & (!n_n2902) & (x15677x)) + ((!n_n2906) & (n_n2908) & (n_n2902) & (!x15677x)) + ((!n_n2906) & (n_n2908) & (n_n2902) & (x15677x)) + ((n_n2906) & (!n_n2908) & (!n_n2902) & (!x15677x)) + ((n_n2906) & (!n_n2908) & (!n_n2902) & (x15677x)) + ((n_n2906) & (!n_n2908) & (n_n2902) & (!x15677x)) + ((n_n2906) & (!n_n2908) & (n_n2902) & (x15677x)) + ((n_n2906) & (n_n2908) & (!n_n2902) & (!x15677x)) + ((n_n2906) & (n_n2908) & (!n_n2902) & (x15677x)) + ((n_n2906) & (n_n2908) & (n_n2902) & (!x15677x)) + ((n_n2906) & (n_n2908) & (n_n2902) & (x15677x)));
	assign n_n2898 = (((!n_n2921) & (!n_n2903) & (!n_n2905) & (!n_n2922) & (x15806x)) + ((!n_n2921) & (!n_n2903) & (!n_n2905) & (n_n2922) & (!x15806x)) + ((!n_n2921) & (!n_n2903) & (!n_n2905) & (n_n2922) & (x15806x)) + ((!n_n2921) & (!n_n2903) & (n_n2905) & (!n_n2922) & (!x15806x)) + ((!n_n2921) & (!n_n2903) & (n_n2905) & (!n_n2922) & (x15806x)) + ((!n_n2921) & (!n_n2903) & (n_n2905) & (n_n2922) & (!x15806x)) + ((!n_n2921) & (!n_n2903) & (n_n2905) & (n_n2922) & (x15806x)) + ((!n_n2921) & (n_n2903) & (!n_n2905) & (!n_n2922) & (!x15806x)) + ((!n_n2921) & (n_n2903) & (!n_n2905) & (!n_n2922) & (x15806x)) + ((!n_n2921) & (n_n2903) & (!n_n2905) & (n_n2922) & (!x15806x)) + ((!n_n2921) & (n_n2903) & (!n_n2905) & (n_n2922) & (x15806x)) + ((!n_n2921) & (n_n2903) & (n_n2905) & (!n_n2922) & (!x15806x)) + ((!n_n2921) & (n_n2903) & (n_n2905) & (!n_n2922) & (x15806x)) + ((!n_n2921) & (n_n2903) & (n_n2905) & (n_n2922) & (!x15806x)) + ((!n_n2921) & (n_n2903) & (n_n2905) & (n_n2922) & (x15806x)) + ((n_n2921) & (!n_n2903) & (!n_n2905) & (!n_n2922) & (!x15806x)) + ((n_n2921) & (!n_n2903) & (!n_n2905) & (!n_n2922) & (x15806x)) + ((n_n2921) & (!n_n2903) & (!n_n2905) & (n_n2922) & (!x15806x)) + ((n_n2921) & (!n_n2903) & (!n_n2905) & (n_n2922) & (x15806x)) + ((n_n2921) & (!n_n2903) & (n_n2905) & (!n_n2922) & (!x15806x)) + ((n_n2921) & (!n_n2903) & (n_n2905) & (!n_n2922) & (x15806x)) + ((n_n2921) & (!n_n2903) & (n_n2905) & (n_n2922) & (!x15806x)) + ((n_n2921) & (!n_n2903) & (n_n2905) & (n_n2922) & (x15806x)) + ((n_n2921) & (n_n2903) & (!n_n2905) & (!n_n2922) & (!x15806x)) + ((n_n2921) & (n_n2903) & (!n_n2905) & (!n_n2922) & (x15806x)) + ((n_n2921) & (n_n2903) & (!n_n2905) & (n_n2922) & (!x15806x)) + ((n_n2921) & (n_n2903) & (!n_n2905) & (n_n2922) & (x15806x)) + ((n_n2921) & (n_n2903) & (n_n2905) & (!n_n2922) & (!x15806x)) + ((n_n2921) & (n_n2903) & (n_n2905) & (!n_n2922) & (x15806x)) + ((n_n2921) & (n_n2903) & (n_n2905) & (n_n2922) & (!x15806x)) + ((n_n2921) & (n_n2903) & (n_n2905) & (n_n2922) & (x15806x)));
	assign x15816x = (((!n_n2827) & (!n_n2821) & (!n_n2826) & (!n_n2907) & (x15811x)) + ((!n_n2827) & (!n_n2821) & (!n_n2826) & (n_n2907) & (!x15811x)) + ((!n_n2827) & (!n_n2821) & (!n_n2826) & (n_n2907) & (x15811x)) + ((!n_n2827) & (!n_n2821) & (n_n2826) & (!n_n2907) & (!x15811x)) + ((!n_n2827) & (!n_n2821) & (n_n2826) & (!n_n2907) & (x15811x)) + ((!n_n2827) & (!n_n2821) & (n_n2826) & (n_n2907) & (!x15811x)) + ((!n_n2827) & (!n_n2821) & (n_n2826) & (n_n2907) & (x15811x)) + ((!n_n2827) & (n_n2821) & (!n_n2826) & (!n_n2907) & (!x15811x)) + ((!n_n2827) & (n_n2821) & (!n_n2826) & (!n_n2907) & (x15811x)) + ((!n_n2827) & (n_n2821) & (!n_n2826) & (n_n2907) & (!x15811x)) + ((!n_n2827) & (n_n2821) & (!n_n2826) & (n_n2907) & (x15811x)) + ((!n_n2827) & (n_n2821) & (n_n2826) & (!n_n2907) & (!x15811x)) + ((!n_n2827) & (n_n2821) & (n_n2826) & (!n_n2907) & (x15811x)) + ((!n_n2827) & (n_n2821) & (n_n2826) & (n_n2907) & (!x15811x)) + ((!n_n2827) & (n_n2821) & (n_n2826) & (n_n2907) & (x15811x)) + ((n_n2827) & (!n_n2821) & (!n_n2826) & (!n_n2907) & (!x15811x)) + ((n_n2827) & (!n_n2821) & (!n_n2826) & (!n_n2907) & (x15811x)) + ((n_n2827) & (!n_n2821) & (!n_n2826) & (n_n2907) & (!x15811x)) + ((n_n2827) & (!n_n2821) & (!n_n2826) & (n_n2907) & (x15811x)) + ((n_n2827) & (!n_n2821) & (n_n2826) & (!n_n2907) & (!x15811x)) + ((n_n2827) & (!n_n2821) & (n_n2826) & (!n_n2907) & (x15811x)) + ((n_n2827) & (!n_n2821) & (n_n2826) & (n_n2907) & (!x15811x)) + ((n_n2827) & (!n_n2821) & (n_n2826) & (n_n2907) & (x15811x)) + ((n_n2827) & (n_n2821) & (!n_n2826) & (!n_n2907) & (!x15811x)) + ((n_n2827) & (n_n2821) & (!n_n2826) & (!n_n2907) & (x15811x)) + ((n_n2827) & (n_n2821) & (!n_n2826) & (n_n2907) & (!x15811x)) + ((n_n2827) & (n_n2821) & (!n_n2826) & (n_n2907) & (x15811x)) + ((n_n2827) & (n_n2821) & (n_n2826) & (!n_n2907) & (!x15811x)) + ((n_n2827) & (n_n2821) & (n_n2826) & (!n_n2907) & (x15811x)) + ((n_n2827) & (n_n2821) & (n_n2826) & (n_n2907) & (!x15811x)) + ((n_n2827) & (n_n2821) & (n_n2826) & (n_n2907) & (x15811x)));
	assign x16324x = (((!n_n1793) & (!n_n1792) & (!n_n1794) & (n_n1787)) + ((!n_n1793) & (!n_n1792) & (n_n1794) & (!n_n1787)) + ((!n_n1793) & (!n_n1792) & (n_n1794) & (n_n1787)) + ((!n_n1793) & (n_n1792) & (!n_n1794) & (!n_n1787)) + ((!n_n1793) & (n_n1792) & (!n_n1794) & (n_n1787)) + ((!n_n1793) & (n_n1792) & (n_n1794) & (!n_n1787)) + ((!n_n1793) & (n_n1792) & (n_n1794) & (n_n1787)) + ((n_n1793) & (!n_n1792) & (!n_n1794) & (!n_n1787)) + ((n_n1793) & (!n_n1792) & (!n_n1794) & (n_n1787)) + ((n_n1793) & (!n_n1792) & (n_n1794) & (!n_n1787)) + ((n_n1793) & (!n_n1792) & (n_n1794) & (n_n1787)) + ((n_n1793) & (n_n1792) & (!n_n1794) & (!n_n1787)) + ((n_n1793) & (n_n1792) & (!n_n1794) & (n_n1787)) + ((n_n1793) & (n_n1792) & (n_n1794) & (!n_n1787)) + ((n_n1793) & (n_n1792) & (n_n1794) & (n_n1787)));
	assign n_n1706 = (((!n_n1709) & (!x15899x) & (!x15900x) & (x15901x)) + ((!n_n1709) & (!x15899x) & (x15900x) & (!x15901x)) + ((!n_n1709) & (!x15899x) & (x15900x) & (x15901x)) + ((!n_n1709) & (x15899x) & (!x15900x) & (!x15901x)) + ((!n_n1709) & (x15899x) & (!x15900x) & (x15901x)) + ((!n_n1709) & (x15899x) & (x15900x) & (!x15901x)) + ((!n_n1709) & (x15899x) & (x15900x) & (x15901x)) + ((n_n1709) & (!x15899x) & (!x15900x) & (!x15901x)) + ((n_n1709) & (!x15899x) & (!x15900x) & (x15901x)) + ((n_n1709) & (!x15899x) & (x15900x) & (!x15901x)) + ((n_n1709) & (!x15899x) & (x15900x) & (x15901x)) + ((n_n1709) & (x15899x) & (!x15900x) & (!x15901x)) + ((n_n1709) & (x15899x) & (!x15900x) & (x15901x)) + ((n_n1709) & (x15899x) & (x15900x) & (!x15901x)) + ((n_n1709) & (x15899x) & (x15900x) & (x15901x)));
	assign x15943x = (((!n_n1712) & (!n_n1711) & (!x15939x) & (x15940x)) + ((!n_n1712) & (!n_n1711) & (x15939x) & (!x15940x)) + ((!n_n1712) & (!n_n1711) & (x15939x) & (x15940x)) + ((!n_n1712) & (n_n1711) & (!x15939x) & (!x15940x)) + ((!n_n1712) & (n_n1711) & (!x15939x) & (x15940x)) + ((!n_n1712) & (n_n1711) & (x15939x) & (!x15940x)) + ((!n_n1712) & (n_n1711) & (x15939x) & (x15940x)) + ((n_n1712) & (!n_n1711) & (!x15939x) & (!x15940x)) + ((n_n1712) & (!n_n1711) & (!x15939x) & (x15940x)) + ((n_n1712) & (!n_n1711) & (x15939x) & (!x15940x)) + ((n_n1712) & (!n_n1711) & (x15939x) & (x15940x)) + ((n_n1712) & (n_n1711) & (!x15939x) & (!x15940x)) + ((n_n1712) & (n_n1711) & (!x15939x) & (x15940x)) + ((n_n1712) & (n_n1711) & (x15939x) & (!x15940x)) + ((n_n1712) & (n_n1711) & (x15939x) & (x15940x)));
	assign n_n1784 = (((!x16242x) & (!n_n1789) & (n_n1790)) + ((!x16242x) & (n_n1789) & (!n_n1790)) + ((!x16242x) & (n_n1789) & (n_n1790)) + ((x16242x) & (!n_n1789) & (!n_n1790)) + ((x16242x) & (!n_n1789) & (n_n1790)) + ((x16242x) & (n_n1789) & (!n_n1790)) + ((x16242x) & (n_n1789) & (n_n1790)));
	assign x16320x = (((!x15991x) & (!x16318x) & (!x16319x) & (!n_n1801) & (n_n1800)) + ((!x15991x) & (!x16318x) & (!x16319x) & (n_n1801) & (!n_n1800)) + ((!x15991x) & (!x16318x) & (!x16319x) & (n_n1801) & (n_n1800)) + ((!x15991x) & (!x16318x) & (x16319x) & (!n_n1801) & (!n_n1800)) + ((!x15991x) & (!x16318x) & (x16319x) & (!n_n1801) & (n_n1800)) + ((!x15991x) & (!x16318x) & (x16319x) & (n_n1801) & (!n_n1800)) + ((!x15991x) & (!x16318x) & (x16319x) & (n_n1801) & (n_n1800)) + ((!x15991x) & (x16318x) & (!x16319x) & (!n_n1801) & (!n_n1800)) + ((!x15991x) & (x16318x) & (!x16319x) & (!n_n1801) & (n_n1800)) + ((!x15991x) & (x16318x) & (!x16319x) & (n_n1801) & (!n_n1800)) + ((!x15991x) & (x16318x) & (!x16319x) & (n_n1801) & (n_n1800)) + ((!x15991x) & (x16318x) & (x16319x) & (!n_n1801) & (!n_n1800)) + ((!x15991x) & (x16318x) & (x16319x) & (!n_n1801) & (n_n1800)) + ((!x15991x) & (x16318x) & (x16319x) & (n_n1801) & (!n_n1800)) + ((!x15991x) & (x16318x) & (x16319x) & (n_n1801) & (n_n1800)) + ((x15991x) & (!x16318x) & (!x16319x) & (!n_n1801) & (!n_n1800)) + ((x15991x) & (!x16318x) & (!x16319x) & (!n_n1801) & (n_n1800)) + ((x15991x) & (!x16318x) & (!x16319x) & (n_n1801) & (!n_n1800)) + ((x15991x) & (!x16318x) & (!x16319x) & (n_n1801) & (n_n1800)) + ((x15991x) & (!x16318x) & (x16319x) & (!n_n1801) & (!n_n1800)) + ((x15991x) & (!x16318x) & (x16319x) & (!n_n1801) & (n_n1800)) + ((x15991x) & (!x16318x) & (x16319x) & (n_n1801) & (!n_n1800)) + ((x15991x) & (!x16318x) & (x16319x) & (n_n1801) & (n_n1800)) + ((x15991x) & (x16318x) & (!x16319x) & (!n_n1801) & (!n_n1800)) + ((x15991x) & (x16318x) & (!x16319x) & (!n_n1801) & (n_n1800)) + ((x15991x) & (x16318x) & (!x16319x) & (n_n1801) & (!n_n1800)) + ((x15991x) & (x16318x) & (!x16319x) & (n_n1801) & (n_n1800)) + ((x15991x) & (x16318x) & (x16319x) & (!n_n1801) & (!n_n1800)) + ((x15991x) & (x16318x) & (x16319x) & (!n_n1801) & (n_n1800)) + ((x15991x) & (x16318x) & (x16319x) & (n_n1801) & (!n_n1800)) + ((x15991x) & (x16318x) & (x16319x) & (n_n1801) & (n_n1800)));
	assign x16831x = (((!x16470x) & (!n_n2165) & (!n_n2164) & (!n_n2162) & (n_n2163)) + ((!x16470x) & (!n_n2165) & (!n_n2164) & (n_n2162) & (!n_n2163)) + ((!x16470x) & (!n_n2165) & (!n_n2164) & (n_n2162) & (n_n2163)) + ((!x16470x) & (!n_n2165) & (n_n2164) & (!n_n2162) & (!n_n2163)) + ((!x16470x) & (!n_n2165) & (n_n2164) & (!n_n2162) & (n_n2163)) + ((!x16470x) & (!n_n2165) & (n_n2164) & (n_n2162) & (!n_n2163)) + ((!x16470x) & (!n_n2165) & (n_n2164) & (n_n2162) & (n_n2163)) + ((!x16470x) & (n_n2165) & (!n_n2164) & (!n_n2162) & (!n_n2163)) + ((!x16470x) & (n_n2165) & (!n_n2164) & (!n_n2162) & (n_n2163)) + ((!x16470x) & (n_n2165) & (!n_n2164) & (n_n2162) & (!n_n2163)) + ((!x16470x) & (n_n2165) & (!n_n2164) & (n_n2162) & (n_n2163)) + ((!x16470x) & (n_n2165) & (n_n2164) & (!n_n2162) & (!n_n2163)) + ((!x16470x) & (n_n2165) & (n_n2164) & (!n_n2162) & (n_n2163)) + ((!x16470x) & (n_n2165) & (n_n2164) & (n_n2162) & (!n_n2163)) + ((!x16470x) & (n_n2165) & (n_n2164) & (n_n2162) & (n_n2163)) + ((x16470x) & (!n_n2165) & (!n_n2164) & (!n_n2162) & (!n_n2163)) + ((x16470x) & (!n_n2165) & (!n_n2164) & (!n_n2162) & (n_n2163)) + ((x16470x) & (!n_n2165) & (!n_n2164) & (n_n2162) & (!n_n2163)) + ((x16470x) & (!n_n2165) & (!n_n2164) & (n_n2162) & (n_n2163)) + ((x16470x) & (!n_n2165) & (n_n2164) & (!n_n2162) & (!n_n2163)) + ((x16470x) & (!n_n2165) & (n_n2164) & (!n_n2162) & (n_n2163)) + ((x16470x) & (!n_n2165) & (n_n2164) & (n_n2162) & (!n_n2163)) + ((x16470x) & (!n_n2165) & (n_n2164) & (n_n2162) & (n_n2163)) + ((x16470x) & (n_n2165) & (!n_n2164) & (!n_n2162) & (!n_n2163)) + ((x16470x) & (n_n2165) & (!n_n2164) & (!n_n2162) & (n_n2163)) + ((x16470x) & (n_n2165) & (!n_n2164) & (n_n2162) & (!n_n2163)) + ((x16470x) & (n_n2165) & (!n_n2164) & (n_n2162) & (n_n2163)) + ((x16470x) & (n_n2165) & (n_n2164) & (!n_n2162) & (!n_n2163)) + ((x16470x) & (n_n2165) & (n_n2164) & (!n_n2162) & (n_n2163)) + ((x16470x) & (n_n2165) & (n_n2164) & (n_n2162) & (!n_n2163)) + ((x16470x) & (n_n2165) & (n_n2164) & (n_n2162) & (n_n2163)));
	assign x16832x = (((!n_n2166) & (!n_n2160) & (!x16764x) & (!x16826x) & (x16827x)) + ((!n_n2166) & (!n_n2160) & (!x16764x) & (x16826x) & (!x16827x)) + ((!n_n2166) & (!n_n2160) & (!x16764x) & (x16826x) & (x16827x)) + ((!n_n2166) & (!n_n2160) & (x16764x) & (!x16826x) & (!x16827x)) + ((!n_n2166) & (!n_n2160) & (x16764x) & (!x16826x) & (x16827x)) + ((!n_n2166) & (!n_n2160) & (x16764x) & (x16826x) & (!x16827x)) + ((!n_n2166) & (!n_n2160) & (x16764x) & (x16826x) & (x16827x)) + ((!n_n2166) & (n_n2160) & (!x16764x) & (!x16826x) & (!x16827x)) + ((!n_n2166) & (n_n2160) & (!x16764x) & (!x16826x) & (x16827x)) + ((!n_n2166) & (n_n2160) & (!x16764x) & (x16826x) & (!x16827x)) + ((!n_n2166) & (n_n2160) & (!x16764x) & (x16826x) & (x16827x)) + ((!n_n2166) & (n_n2160) & (x16764x) & (!x16826x) & (!x16827x)) + ((!n_n2166) & (n_n2160) & (x16764x) & (!x16826x) & (x16827x)) + ((!n_n2166) & (n_n2160) & (x16764x) & (x16826x) & (!x16827x)) + ((!n_n2166) & (n_n2160) & (x16764x) & (x16826x) & (x16827x)) + ((n_n2166) & (!n_n2160) & (!x16764x) & (!x16826x) & (!x16827x)) + ((n_n2166) & (!n_n2160) & (!x16764x) & (!x16826x) & (x16827x)) + ((n_n2166) & (!n_n2160) & (!x16764x) & (x16826x) & (!x16827x)) + ((n_n2166) & (!n_n2160) & (!x16764x) & (x16826x) & (x16827x)) + ((n_n2166) & (!n_n2160) & (x16764x) & (!x16826x) & (!x16827x)) + ((n_n2166) & (!n_n2160) & (x16764x) & (!x16826x) & (x16827x)) + ((n_n2166) & (!n_n2160) & (x16764x) & (x16826x) & (!x16827x)) + ((n_n2166) & (!n_n2160) & (x16764x) & (x16826x) & (x16827x)) + ((n_n2166) & (n_n2160) & (!x16764x) & (!x16826x) & (!x16827x)) + ((n_n2166) & (n_n2160) & (!x16764x) & (!x16826x) & (x16827x)) + ((n_n2166) & (n_n2160) & (!x16764x) & (x16826x) & (!x16827x)) + ((n_n2166) & (n_n2160) & (!x16764x) & (x16826x) & (x16827x)) + ((n_n2166) & (n_n2160) & (x16764x) & (!x16826x) & (!x16827x)) + ((n_n2166) & (n_n2160) & (x16764x) & (!x16826x) & (x16827x)) + ((n_n2166) & (n_n2160) & (x16764x) & (x16826x) & (!x16827x)) + ((n_n2166) & (n_n2160) & (x16764x) & (x16826x) & (x16827x)));
	assign n_n1014 = (((!x11530x) & (!n_n1107) & (!x11501x) & (!n_n1038) & (x11500x)) + ((!x11530x) & (!n_n1107) & (!x11501x) & (n_n1038) & (!x11500x)) + ((!x11530x) & (!n_n1107) & (!x11501x) & (n_n1038) & (x11500x)) + ((!x11530x) & (!n_n1107) & (x11501x) & (!n_n1038) & (!x11500x)) + ((!x11530x) & (!n_n1107) & (x11501x) & (!n_n1038) & (x11500x)) + ((!x11530x) & (!n_n1107) & (x11501x) & (n_n1038) & (!x11500x)) + ((!x11530x) & (!n_n1107) & (x11501x) & (n_n1038) & (x11500x)) + ((!x11530x) & (n_n1107) & (!x11501x) & (!n_n1038) & (!x11500x)) + ((!x11530x) & (n_n1107) & (!x11501x) & (!n_n1038) & (x11500x)) + ((!x11530x) & (n_n1107) & (!x11501x) & (n_n1038) & (!x11500x)) + ((!x11530x) & (n_n1107) & (!x11501x) & (n_n1038) & (x11500x)) + ((!x11530x) & (n_n1107) & (x11501x) & (!n_n1038) & (!x11500x)) + ((!x11530x) & (n_n1107) & (x11501x) & (!n_n1038) & (x11500x)) + ((!x11530x) & (n_n1107) & (x11501x) & (n_n1038) & (!x11500x)) + ((!x11530x) & (n_n1107) & (x11501x) & (n_n1038) & (x11500x)) + ((x11530x) & (!n_n1107) & (!x11501x) & (!n_n1038) & (!x11500x)) + ((x11530x) & (!n_n1107) & (!x11501x) & (!n_n1038) & (x11500x)) + ((x11530x) & (!n_n1107) & (!x11501x) & (n_n1038) & (!x11500x)) + ((x11530x) & (!n_n1107) & (!x11501x) & (n_n1038) & (x11500x)) + ((x11530x) & (!n_n1107) & (x11501x) & (!n_n1038) & (!x11500x)) + ((x11530x) & (!n_n1107) & (x11501x) & (!n_n1038) & (x11500x)) + ((x11530x) & (!n_n1107) & (x11501x) & (n_n1038) & (!x11500x)) + ((x11530x) & (!n_n1107) & (x11501x) & (n_n1038) & (x11500x)) + ((x11530x) & (n_n1107) & (!x11501x) & (!n_n1038) & (!x11500x)) + ((x11530x) & (n_n1107) & (!x11501x) & (!n_n1038) & (x11500x)) + ((x11530x) & (n_n1107) & (!x11501x) & (n_n1038) & (!x11500x)) + ((x11530x) & (n_n1107) & (!x11501x) & (n_n1038) & (x11500x)) + ((x11530x) & (n_n1107) & (x11501x) & (!n_n1038) & (!x11500x)) + ((x11530x) & (n_n1107) & (x11501x) & (!n_n1038) & (x11500x)) + ((x11530x) & (n_n1107) & (x11501x) & (n_n1038) & (!x11500x)) + ((x11530x) & (n_n1107) & (x11501x) & (n_n1038) & (x11500x)));
	assign n_n1013 = (((!x11581x) & (!n_n1034) & (n_n1035)) + ((!x11581x) & (n_n1034) & (!n_n1035)) + ((!x11581x) & (n_n1034) & (n_n1035)) + ((x11581x) & (!n_n1034) & (!n_n1035)) + ((x11581x) & (!n_n1034) & (n_n1035)) + ((x11581x) & (n_n1034) & (!n_n1035)) + ((x11581x) & (n_n1034) & (n_n1035)));
	assign x11894x = (((!n_n1083) & (!n_n1082) & (!x11766x) & (!n_n1028) & (x11892x)) + ((!n_n1083) & (!n_n1082) & (!x11766x) & (n_n1028) & (!x11892x)) + ((!n_n1083) & (!n_n1082) & (!x11766x) & (n_n1028) & (x11892x)) + ((!n_n1083) & (!n_n1082) & (x11766x) & (!n_n1028) & (!x11892x)) + ((!n_n1083) & (!n_n1082) & (x11766x) & (!n_n1028) & (x11892x)) + ((!n_n1083) & (!n_n1082) & (x11766x) & (n_n1028) & (!x11892x)) + ((!n_n1083) & (!n_n1082) & (x11766x) & (n_n1028) & (x11892x)) + ((!n_n1083) & (n_n1082) & (!x11766x) & (!n_n1028) & (!x11892x)) + ((!n_n1083) & (n_n1082) & (!x11766x) & (!n_n1028) & (x11892x)) + ((!n_n1083) & (n_n1082) & (!x11766x) & (n_n1028) & (!x11892x)) + ((!n_n1083) & (n_n1082) & (!x11766x) & (n_n1028) & (x11892x)) + ((!n_n1083) & (n_n1082) & (x11766x) & (!n_n1028) & (!x11892x)) + ((!n_n1083) & (n_n1082) & (x11766x) & (!n_n1028) & (x11892x)) + ((!n_n1083) & (n_n1082) & (x11766x) & (n_n1028) & (!x11892x)) + ((!n_n1083) & (n_n1082) & (x11766x) & (n_n1028) & (x11892x)) + ((n_n1083) & (!n_n1082) & (!x11766x) & (!n_n1028) & (!x11892x)) + ((n_n1083) & (!n_n1082) & (!x11766x) & (!n_n1028) & (x11892x)) + ((n_n1083) & (!n_n1082) & (!x11766x) & (n_n1028) & (!x11892x)) + ((n_n1083) & (!n_n1082) & (!x11766x) & (n_n1028) & (x11892x)) + ((n_n1083) & (!n_n1082) & (x11766x) & (!n_n1028) & (!x11892x)) + ((n_n1083) & (!n_n1082) & (x11766x) & (!n_n1028) & (x11892x)) + ((n_n1083) & (!n_n1082) & (x11766x) & (n_n1028) & (!x11892x)) + ((n_n1083) & (!n_n1082) & (x11766x) & (n_n1028) & (x11892x)) + ((n_n1083) & (n_n1082) & (!x11766x) & (!n_n1028) & (!x11892x)) + ((n_n1083) & (n_n1082) & (!x11766x) & (!n_n1028) & (x11892x)) + ((n_n1083) & (n_n1082) & (!x11766x) & (n_n1028) & (!x11892x)) + ((n_n1083) & (n_n1082) & (!x11766x) & (n_n1028) & (x11892x)) + ((n_n1083) & (n_n1082) & (x11766x) & (!n_n1028) & (!x11892x)) + ((n_n1083) & (n_n1082) & (x11766x) & (!n_n1028) & (x11892x)) + ((n_n1083) & (n_n1082) & (x11766x) & (n_n1028) & (!x11892x)) + ((n_n1083) & (n_n1082) & (x11766x) & (n_n1028) & (x11892x)));
	assign n_n1010 = (((!n_n1026) & (!n_n1071) & (!n_n1072) & (!x11815x) & (x11832x)) + ((!n_n1026) & (!n_n1071) & (!n_n1072) & (x11815x) & (!x11832x)) + ((!n_n1026) & (!n_n1071) & (!n_n1072) & (x11815x) & (x11832x)) + ((!n_n1026) & (!n_n1071) & (n_n1072) & (!x11815x) & (!x11832x)) + ((!n_n1026) & (!n_n1071) & (n_n1072) & (!x11815x) & (x11832x)) + ((!n_n1026) & (!n_n1071) & (n_n1072) & (x11815x) & (!x11832x)) + ((!n_n1026) & (!n_n1071) & (n_n1072) & (x11815x) & (x11832x)) + ((!n_n1026) & (n_n1071) & (!n_n1072) & (!x11815x) & (!x11832x)) + ((!n_n1026) & (n_n1071) & (!n_n1072) & (!x11815x) & (x11832x)) + ((!n_n1026) & (n_n1071) & (!n_n1072) & (x11815x) & (!x11832x)) + ((!n_n1026) & (n_n1071) & (!n_n1072) & (x11815x) & (x11832x)) + ((!n_n1026) & (n_n1071) & (n_n1072) & (!x11815x) & (!x11832x)) + ((!n_n1026) & (n_n1071) & (n_n1072) & (!x11815x) & (x11832x)) + ((!n_n1026) & (n_n1071) & (n_n1072) & (x11815x) & (!x11832x)) + ((!n_n1026) & (n_n1071) & (n_n1072) & (x11815x) & (x11832x)) + ((n_n1026) & (!n_n1071) & (!n_n1072) & (!x11815x) & (!x11832x)) + ((n_n1026) & (!n_n1071) & (!n_n1072) & (!x11815x) & (x11832x)) + ((n_n1026) & (!n_n1071) & (!n_n1072) & (x11815x) & (!x11832x)) + ((n_n1026) & (!n_n1071) & (!n_n1072) & (x11815x) & (x11832x)) + ((n_n1026) & (!n_n1071) & (n_n1072) & (!x11815x) & (!x11832x)) + ((n_n1026) & (!n_n1071) & (n_n1072) & (!x11815x) & (x11832x)) + ((n_n1026) & (!n_n1071) & (n_n1072) & (x11815x) & (!x11832x)) + ((n_n1026) & (!n_n1071) & (n_n1072) & (x11815x) & (x11832x)) + ((n_n1026) & (n_n1071) & (!n_n1072) & (!x11815x) & (!x11832x)) + ((n_n1026) & (n_n1071) & (!n_n1072) & (!x11815x) & (x11832x)) + ((n_n1026) & (n_n1071) & (!n_n1072) & (x11815x) & (!x11832x)) + ((n_n1026) & (n_n1071) & (!n_n1072) & (x11815x) & (x11832x)) + ((n_n1026) & (n_n1071) & (n_n1072) & (!x11815x) & (!x11832x)) + ((n_n1026) & (n_n1071) & (n_n1072) & (!x11815x) & (x11832x)) + ((n_n1026) & (n_n1071) & (n_n1072) & (x11815x) & (!x11832x)) + ((n_n1026) & (n_n1071) & (n_n1072) & (x11815x) & (x11832x)));
	assign n_n1012 = (((!n_n1088) & (!x11851x) & (!n_n1032) & (!x11884x) & (x11850x)) + ((!n_n1088) & (!x11851x) & (!n_n1032) & (x11884x) & (!x11850x)) + ((!n_n1088) & (!x11851x) & (!n_n1032) & (x11884x) & (x11850x)) + ((!n_n1088) & (!x11851x) & (n_n1032) & (!x11884x) & (!x11850x)) + ((!n_n1088) & (!x11851x) & (n_n1032) & (!x11884x) & (x11850x)) + ((!n_n1088) & (!x11851x) & (n_n1032) & (x11884x) & (!x11850x)) + ((!n_n1088) & (!x11851x) & (n_n1032) & (x11884x) & (x11850x)) + ((!n_n1088) & (x11851x) & (!n_n1032) & (!x11884x) & (!x11850x)) + ((!n_n1088) & (x11851x) & (!n_n1032) & (!x11884x) & (x11850x)) + ((!n_n1088) & (x11851x) & (!n_n1032) & (x11884x) & (!x11850x)) + ((!n_n1088) & (x11851x) & (!n_n1032) & (x11884x) & (x11850x)) + ((!n_n1088) & (x11851x) & (n_n1032) & (!x11884x) & (!x11850x)) + ((!n_n1088) & (x11851x) & (n_n1032) & (!x11884x) & (x11850x)) + ((!n_n1088) & (x11851x) & (n_n1032) & (x11884x) & (!x11850x)) + ((!n_n1088) & (x11851x) & (n_n1032) & (x11884x) & (x11850x)) + ((n_n1088) & (!x11851x) & (!n_n1032) & (!x11884x) & (!x11850x)) + ((n_n1088) & (!x11851x) & (!n_n1032) & (!x11884x) & (x11850x)) + ((n_n1088) & (!x11851x) & (!n_n1032) & (x11884x) & (!x11850x)) + ((n_n1088) & (!x11851x) & (!n_n1032) & (x11884x) & (x11850x)) + ((n_n1088) & (!x11851x) & (n_n1032) & (!x11884x) & (!x11850x)) + ((n_n1088) & (!x11851x) & (n_n1032) & (!x11884x) & (x11850x)) + ((n_n1088) & (!x11851x) & (n_n1032) & (x11884x) & (!x11850x)) + ((n_n1088) & (!x11851x) & (n_n1032) & (x11884x) & (x11850x)) + ((n_n1088) & (x11851x) & (!n_n1032) & (!x11884x) & (!x11850x)) + ((n_n1088) & (x11851x) & (!n_n1032) & (!x11884x) & (x11850x)) + ((n_n1088) & (x11851x) & (!n_n1032) & (x11884x) & (!x11850x)) + ((n_n1088) & (x11851x) & (!n_n1032) & (x11884x) & (x11850x)) + ((n_n1088) & (x11851x) & (n_n1032) & (!x11884x) & (!x11850x)) + ((n_n1088) & (x11851x) & (n_n1032) & (!x11884x) & (x11850x)) + ((n_n1088) & (x11851x) & (n_n1032) & (x11884x) & (!x11850x)) + ((n_n1088) & (x11851x) & (n_n1032) & (x11884x) & (x11850x)));
	assign n_n1396 = (((!x12199x) & (!n_n1412) & (n_n1413)) + ((!x12199x) & (n_n1412) & (!n_n1413)) + ((!x12199x) & (n_n1412) & (n_n1413)) + ((x12199x) & (!n_n1412) & (!n_n1413)) + ((x12199x) & (!n_n1412) & (n_n1413)) + ((x12199x) & (n_n1412) & (!n_n1413)) + ((x12199x) & (n_n1412) & (n_n1413)));
	assign n_n1397 = (((!x12247x) & (!n_n1466) & (!x12223x) & (!n_n1415) & (x12222x)) + ((!x12247x) & (!n_n1466) & (!x12223x) & (n_n1415) & (!x12222x)) + ((!x12247x) & (!n_n1466) & (!x12223x) & (n_n1415) & (x12222x)) + ((!x12247x) & (!n_n1466) & (x12223x) & (!n_n1415) & (!x12222x)) + ((!x12247x) & (!n_n1466) & (x12223x) & (!n_n1415) & (x12222x)) + ((!x12247x) & (!n_n1466) & (x12223x) & (n_n1415) & (!x12222x)) + ((!x12247x) & (!n_n1466) & (x12223x) & (n_n1415) & (x12222x)) + ((!x12247x) & (n_n1466) & (!x12223x) & (!n_n1415) & (!x12222x)) + ((!x12247x) & (n_n1466) & (!x12223x) & (!n_n1415) & (x12222x)) + ((!x12247x) & (n_n1466) & (!x12223x) & (n_n1415) & (!x12222x)) + ((!x12247x) & (n_n1466) & (!x12223x) & (n_n1415) & (x12222x)) + ((!x12247x) & (n_n1466) & (x12223x) & (!n_n1415) & (!x12222x)) + ((!x12247x) & (n_n1466) & (x12223x) & (!n_n1415) & (x12222x)) + ((!x12247x) & (n_n1466) & (x12223x) & (n_n1415) & (!x12222x)) + ((!x12247x) & (n_n1466) & (x12223x) & (n_n1415) & (x12222x)) + ((x12247x) & (!n_n1466) & (!x12223x) & (!n_n1415) & (!x12222x)) + ((x12247x) & (!n_n1466) & (!x12223x) & (!n_n1415) & (x12222x)) + ((x12247x) & (!n_n1466) & (!x12223x) & (n_n1415) & (!x12222x)) + ((x12247x) & (!n_n1466) & (!x12223x) & (n_n1415) & (x12222x)) + ((x12247x) & (!n_n1466) & (x12223x) & (!n_n1415) & (!x12222x)) + ((x12247x) & (!n_n1466) & (x12223x) & (!n_n1415) & (x12222x)) + ((x12247x) & (!n_n1466) & (x12223x) & (n_n1415) & (!x12222x)) + ((x12247x) & (!n_n1466) & (x12223x) & (n_n1415) & (x12222x)) + ((x12247x) & (n_n1466) & (!x12223x) & (!n_n1415) & (!x12222x)) + ((x12247x) & (n_n1466) & (!x12223x) & (!n_n1415) & (x12222x)) + ((x12247x) & (n_n1466) & (!x12223x) & (n_n1415) & (!x12222x)) + ((x12247x) & (n_n1466) & (!x12223x) & (n_n1415) & (x12222x)) + ((x12247x) & (n_n1466) & (x12223x) & (!n_n1415) & (!x12222x)) + ((x12247x) & (n_n1466) & (x12223x) & (!n_n1415) & (x12222x)) + ((x12247x) & (n_n1466) & (x12223x) & (n_n1415) & (!x12222x)) + ((x12247x) & (n_n1466) & (x12223x) & (n_n1415) & (x12222x)));
	assign x12391x = (((!n_n1450) & (!n_n1451) & (!x12324x) & (!n_n1408) & (x12389x)) + ((!n_n1450) & (!n_n1451) & (!x12324x) & (n_n1408) & (!x12389x)) + ((!n_n1450) & (!n_n1451) & (!x12324x) & (n_n1408) & (x12389x)) + ((!n_n1450) & (!n_n1451) & (x12324x) & (!n_n1408) & (!x12389x)) + ((!n_n1450) & (!n_n1451) & (x12324x) & (!n_n1408) & (x12389x)) + ((!n_n1450) & (!n_n1451) & (x12324x) & (n_n1408) & (!x12389x)) + ((!n_n1450) & (!n_n1451) & (x12324x) & (n_n1408) & (x12389x)) + ((!n_n1450) & (n_n1451) & (!x12324x) & (!n_n1408) & (!x12389x)) + ((!n_n1450) & (n_n1451) & (!x12324x) & (!n_n1408) & (x12389x)) + ((!n_n1450) & (n_n1451) & (!x12324x) & (n_n1408) & (!x12389x)) + ((!n_n1450) & (n_n1451) & (!x12324x) & (n_n1408) & (x12389x)) + ((!n_n1450) & (n_n1451) & (x12324x) & (!n_n1408) & (!x12389x)) + ((!n_n1450) & (n_n1451) & (x12324x) & (!n_n1408) & (x12389x)) + ((!n_n1450) & (n_n1451) & (x12324x) & (n_n1408) & (!x12389x)) + ((!n_n1450) & (n_n1451) & (x12324x) & (n_n1408) & (x12389x)) + ((n_n1450) & (!n_n1451) & (!x12324x) & (!n_n1408) & (!x12389x)) + ((n_n1450) & (!n_n1451) & (!x12324x) & (!n_n1408) & (x12389x)) + ((n_n1450) & (!n_n1451) & (!x12324x) & (n_n1408) & (!x12389x)) + ((n_n1450) & (!n_n1451) & (!x12324x) & (n_n1408) & (x12389x)) + ((n_n1450) & (!n_n1451) & (x12324x) & (!n_n1408) & (!x12389x)) + ((n_n1450) & (!n_n1451) & (x12324x) & (!n_n1408) & (x12389x)) + ((n_n1450) & (!n_n1451) & (x12324x) & (n_n1408) & (!x12389x)) + ((n_n1450) & (!n_n1451) & (x12324x) & (n_n1408) & (x12389x)) + ((n_n1450) & (n_n1451) & (!x12324x) & (!n_n1408) & (!x12389x)) + ((n_n1450) & (n_n1451) & (!x12324x) & (!n_n1408) & (x12389x)) + ((n_n1450) & (n_n1451) & (!x12324x) & (n_n1408) & (!x12389x)) + ((n_n1450) & (n_n1451) & (!x12324x) & (n_n1408) & (x12389x)) + ((n_n1450) & (n_n1451) & (x12324x) & (!n_n1408) & (!x12389x)) + ((n_n1450) & (n_n1451) & (x12324x) & (!n_n1408) & (x12389x)) + ((n_n1450) & (n_n1451) & (x12324x) & (n_n1408) & (!x12389x)) + ((n_n1450) & (n_n1451) & (x12324x) & (n_n1408) & (x12389x)));
	assign n_n1394 = (((!n_n1442) & (!n_n1405) & (!x12296x) & (!x12305x) & (x12295x)) + ((!n_n1442) & (!n_n1405) & (!x12296x) & (x12305x) & (!x12295x)) + ((!n_n1442) & (!n_n1405) & (!x12296x) & (x12305x) & (x12295x)) + ((!n_n1442) & (!n_n1405) & (x12296x) & (!x12305x) & (!x12295x)) + ((!n_n1442) & (!n_n1405) & (x12296x) & (!x12305x) & (x12295x)) + ((!n_n1442) & (!n_n1405) & (x12296x) & (x12305x) & (!x12295x)) + ((!n_n1442) & (!n_n1405) & (x12296x) & (x12305x) & (x12295x)) + ((!n_n1442) & (n_n1405) & (!x12296x) & (!x12305x) & (!x12295x)) + ((!n_n1442) & (n_n1405) & (!x12296x) & (!x12305x) & (x12295x)) + ((!n_n1442) & (n_n1405) & (!x12296x) & (x12305x) & (!x12295x)) + ((!n_n1442) & (n_n1405) & (!x12296x) & (x12305x) & (x12295x)) + ((!n_n1442) & (n_n1405) & (x12296x) & (!x12305x) & (!x12295x)) + ((!n_n1442) & (n_n1405) & (x12296x) & (!x12305x) & (x12295x)) + ((!n_n1442) & (n_n1405) & (x12296x) & (x12305x) & (!x12295x)) + ((!n_n1442) & (n_n1405) & (x12296x) & (x12305x) & (x12295x)) + ((n_n1442) & (!n_n1405) & (!x12296x) & (!x12305x) & (!x12295x)) + ((n_n1442) & (!n_n1405) & (!x12296x) & (!x12305x) & (x12295x)) + ((n_n1442) & (!n_n1405) & (!x12296x) & (x12305x) & (!x12295x)) + ((n_n1442) & (!n_n1405) & (!x12296x) & (x12305x) & (x12295x)) + ((n_n1442) & (!n_n1405) & (x12296x) & (!x12305x) & (!x12295x)) + ((n_n1442) & (!n_n1405) & (x12296x) & (!x12305x) & (x12295x)) + ((n_n1442) & (!n_n1405) & (x12296x) & (x12305x) & (!x12295x)) + ((n_n1442) & (!n_n1405) & (x12296x) & (x12305x) & (x12295x)) + ((n_n1442) & (n_n1405) & (!x12296x) & (!x12305x) & (!x12295x)) + ((n_n1442) & (n_n1405) & (!x12296x) & (!x12305x) & (x12295x)) + ((n_n1442) & (n_n1405) & (!x12296x) & (x12305x) & (!x12295x)) + ((n_n1442) & (n_n1405) & (!x12296x) & (x12305x) & (x12295x)) + ((n_n1442) & (n_n1405) & (x12296x) & (!x12305x) & (!x12295x)) + ((n_n1442) & (n_n1405) & (x12296x) & (!x12305x) & (x12295x)) + ((n_n1442) & (n_n1405) & (x12296x) & (x12305x) & (!x12295x)) + ((n_n1442) & (n_n1405) & (x12296x) & (x12305x) & (x12295x)));
	assign n_n1393 = (((!n_n1404) & (!x12381x) & (x12380x)) + ((!n_n1404) & (x12381x) & (!x12380x)) + ((!n_n1404) & (x12381x) & (x12380x)) + ((n_n1404) & (!x12381x) & (!x12380x)) + ((n_n1404) & (!x12381x) & (x12380x)) + ((n_n1404) & (x12381x) & (!x12380x)) + ((n_n1404) & (x12381x) & (x12380x)));
	assign x12693x = (((!n_n553) & (!x12683x) & (!x12684x) & (!x12689x) & (x12690x)) + ((!n_n553) & (!x12683x) & (!x12684x) & (x12689x) & (!x12690x)) + ((!n_n553) & (!x12683x) & (!x12684x) & (x12689x) & (x12690x)) + ((!n_n553) & (!x12683x) & (x12684x) & (!x12689x) & (!x12690x)) + ((!n_n553) & (!x12683x) & (x12684x) & (!x12689x) & (x12690x)) + ((!n_n553) & (!x12683x) & (x12684x) & (x12689x) & (!x12690x)) + ((!n_n553) & (!x12683x) & (x12684x) & (x12689x) & (x12690x)) + ((!n_n553) & (x12683x) & (!x12684x) & (!x12689x) & (!x12690x)) + ((!n_n553) & (x12683x) & (!x12684x) & (!x12689x) & (x12690x)) + ((!n_n553) & (x12683x) & (!x12684x) & (x12689x) & (!x12690x)) + ((!n_n553) & (x12683x) & (!x12684x) & (x12689x) & (x12690x)) + ((!n_n553) & (x12683x) & (x12684x) & (!x12689x) & (!x12690x)) + ((!n_n553) & (x12683x) & (x12684x) & (!x12689x) & (x12690x)) + ((!n_n553) & (x12683x) & (x12684x) & (x12689x) & (!x12690x)) + ((!n_n553) & (x12683x) & (x12684x) & (x12689x) & (x12690x)) + ((n_n553) & (!x12683x) & (!x12684x) & (!x12689x) & (!x12690x)) + ((n_n553) & (!x12683x) & (!x12684x) & (!x12689x) & (x12690x)) + ((n_n553) & (!x12683x) & (!x12684x) & (x12689x) & (!x12690x)) + ((n_n553) & (!x12683x) & (!x12684x) & (x12689x) & (x12690x)) + ((n_n553) & (!x12683x) & (x12684x) & (!x12689x) & (!x12690x)) + ((n_n553) & (!x12683x) & (x12684x) & (!x12689x) & (x12690x)) + ((n_n553) & (!x12683x) & (x12684x) & (x12689x) & (!x12690x)) + ((n_n553) & (!x12683x) & (x12684x) & (x12689x) & (x12690x)) + ((n_n553) & (x12683x) & (!x12684x) & (!x12689x) & (!x12690x)) + ((n_n553) & (x12683x) & (!x12684x) & (!x12689x) & (x12690x)) + ((n_n553) & (x12683x) & (!x12684x) & (x12689x) & (!x12690x)) + ((n_n553) & (x12683x) & (!x12684x) & (x12689x) & (x12690x)) + ((n_n553) & (x12683x) & (x12684x) & (!x12689x) & (!x12690x)) + ((n_n553) & (x12683x) & (x12684x) & (!x12689x) & (x12690x)) + ((n_n553) & (x12683x) & (x12684x) & (x12689x) & (!x12690x)) + ((n_n553) & (x12683x) & (x12684x) & (x12689x) & (x12690x)));
	assign n_n539 = (((!n_n546) & (!x12640x) & (!x12641x) & (!x12647x) & (x12648x)) + ((!n_n546) & (!x12640x) & (!x12641x) & (x12647x) & (!x12648x)) + ((!n_n546) & (!x12640x) & (!x12641x) & (x12647x) & (x12648x)) + ((!n_n546) & (!x12640x) & (x12641x) & (!x12647x) & (!x12648x)) + ((!n_n546) & (!x12640x) & (x12641x) & (!x12647x) & (x12648x)) + ((!n_n546) & (!x12640x) & (x12641x) & (x12647x) & (!x12648x)) + ((!n_n546) & (!x12640x) & (x12641x) & (x12647x) & (x12648x)) + ((!n_n546) & (x12640x) & (!x12641x) & (!x12647x) & (!x12648x)) + ((!n_n546) & (x12640x) & (!x12641x) & (!x12647x) & (x12648x)) + ((!n_n546) & (x12640x) & (!x12641x) & (x12647x) & (!x12648x)) + ((!n_n546) & (x12640x) & (!x12641x) & (x12647x) & (x12648x)) + ((!n_n546) & (x12640x) & (x12641x) & (!x12647x) & (!x12648x)) + ((!n_n546) & (x12640x) & (x12641x) & (!x12647x) & (x12648x)) + ((!n_n546) & (x12640x) & (x12641x) & (x12647x) & (!x12648x)) + ((!n_n546) & (x12640x) & (x12641x) & (x12647x) & (x12648x)) + ((n_n546) & (!x12640x) & (!x12641x) & (!x12647x) & (!x12648x)) + ((n_n546) & (!x12640x) & (!x12641x) & (!x12647x) & (x12648x)) + ((n_n546) & (!x12640x) & (!x12641x) & (x12647x) & (!x12648x)) + ((n_n546) & (!x12640x) & (!x12641x) & (x12647x) & (x12648x)) + ((n_n546) & (!x12640x) & (x12641x) & (!x12647x) & (!x12648x)) + ((n_n546) & (!x12640x) & (x12641x) & (!x12647x) & (x12648x)) + ((n_n546) & (!x12640x) & (x12641x) & (x12647x) & (!x12648x)) + ((n_n546) & (!x12640x) & (x12641x) & (x12647x) & (x12648x)) + ((n_n546) & (x12640x) & (!x12641x) & (!x12647x) & (!x12648x)) + ((n_n546) & (x12640x) & (!x12641x) & (!x12647x) & (x12648x)) + ((n_n546) & (x12640x) & (!x12641x) & (x12647x) & (!x12648x)) + ((n_n546) & (x12640x) & (!x12641x) & (x12647x) & (x12648x)) + ((n_n546) & (x12640x) & (x12641x) & (!x12647x) & (!x12648x)) + ((n_n546) & (x12640x) & (x12641x) & (!x12647x) & (x12648x)) + ((n_n546) & (x12640x) & (x12641x) & (x12647x) & (!x12648x)) + ((n_n546) & (x12640x) & (x12641x) & (x12647x) & (x12648x)));
	assign n_n540 = (((!x12656x) & (!x12657x) & (!n_n551) & (!x12670x) & (x12671x)) + ((!x12656x) & (!x12657x) & (!n_n551) & (x12670x) & (!x12671x)) + ((!x12656x) & (!x12657x) & (!n_n551) & (x12670x) & (x12671x)) + ((!x12656x) & (!x12657x) & (n_n551) & (!x12670x) & (!x12671x)) + ((!x12656x) & (!x12657x) & (n_n551) & (!x12670x) & (x12671x)) + ((!x12656x) & (!x12657x) & (n_n551) & (x12670x) & (!x12671x)) + ((!x12656x) & (!x12657x) & (n_n551) & (x12670x) & (x12671x)) + ((!x12656x) & (x12657x) & (!n_n551) & (!x12670x) & (!x12671x)) + ((!x12656x) & (x12657x) & (!n_n551) & (!x12670x) & (x12671x)) + ((!x12656x) & (x12657x) & (!n_n551) & (x12670x) & (!x12671x)) + ((!x12656x) & (x12657x) & (!n_n551) & (x12670x) & (x12671x)) + ((!x12656x) & (x12657x) & (n_n551) & (!x12670x) & (!x12671x)) + ((!x12656x) & (x12657x) & (n_n551) & (!x12670x) & (x12671x)) + ((!x12656x) & (x12657x) & (n_n551) & (x12670x) & (!x12671x)) + ((!x12656x) & (x12657x) & (n_n551) & (x12670x) & (x12671x)) + ((x12656x) & (!x12657x) & (!n_n551) & (!x12670x) & (!x12671x)) + ((x12656x) & (!x12657x) & (!n_n551) & (!x12670x) & (x12671x)) + ((x12656x) & (!x12657x) & (!n_n551) & (x12670x) & (!x12671x)) + ((x12656x) & (!x12657x) & (!n_n551) & (x12670x) & (x12671x)) + ((x12656x) & (!x12657x) & (n_n551) & (!x12670x) & (!x12671x)) + ((x12656x) & (!x12657x) & (n_n551) & (!x12670x) & (x12671x)) + ((x12656x) & (!x12657x) & (n_n551) & (x12670x) & (!x12671x)) + ((x12656x) & (!x12657x) & (n_n551) & (x12670x) & (x12671x)) + ((x12656x) & (x12657x) & (!n_n551) & (!x12670x) & (!x12671x)) + ((x12656x) & (x12657x) & (!n_n551) & (!x12670x) & (x12671x)) + ((x12656x) & (x12657x) & (!n_n551) & (x12670x) & (!x12671x)) + ((x12656x) & (x12657x) & (!n_n551) & (x12670x) & (x12671x)) + ((x12656x) & (x12657x) & (n_n551) & (!x12670x) & (!x12671x)) + ((x12656x) & (x12657x) & (n_n551) & (!x12670x) & (x12671x)) + ((x12656x) & (x12657x) & (n_n551) & (x12670x) & (!x12671x)) + ((x12656x) & (x12657x) & (n_n551) & (x12670x) & (x12671x)));
	assign x13146x = (((!n_n543) & (!n_n542) & (!x13142x) & (x13143x)) + ((!n_n543) & (!n_n542) & (x13142x) & (!x13143x)) + ((!n_n543) & (!n_n542) & (x13142x) & (x13143x)) + ((!n_n543) & (n_n542) & (!x13142x) & (!x13143x)) + ((!n_n543) & (n_n542) & (!x13142x) & (x13143x)) + ((!n_n543) & (n_n542) & (x13142x) & (!x13143x)) + ((!n_n543) & (n_n542) & (x13142x) & (x13143x)) + ((n_n543) & (!n_n542) & (!x13142x) & (!x13143x)) + ((n_n543) & (!n_n542) & (!x13142x) & (x13143x)) + ((n_n543) & (!n_n542) & (x13142x) & (!x13143x)) + ((n_n543) & (!n_n542) & (x13142x) & (x13143x)) + ((n_n543) & (n_n542) & (!x13142x) & (!x13143x)) + ((n_n543) & (n_n542) & (!x13142x) & (x13143x)) + ((n_n543) & (n_n542) & (x13142x) & (!x13143x)) + ((n_n543) & (n_n542) & (x13142x) & (x13143x)));
	assign x13645x = (((!n_n4748) & (!n_n4725) & (!n_n4788) & (!n_n4802) & (x13644x)) + ((!n_n4748) & (!n_n4725) & (!n_n4788) & (n_n4802) & (!x13644x)) + ((!n_n4748) & (!n_n4725) & (!n_n4788) & (n_n4802) & (x13644x)) + ((!n_n4748) & (!n_n4725) & (n_n4788) & (!n_n4802) & (!x13644x)) + ((!n_n4748) & (!n_n4725) & (n_n4788) & (!n_n4802) & (x13644x)) + ((!n_n4748) & (!n_n4725) & (n_n4788) & (n_n4802) & (!x13644x)) + ((!n_n4748) & (!n_n4725) & (n_n4788) & (n_n4802) & (x13644x)) + ((!n_n4748) & (n_n4725) & (!n_n4788) & (!n_n4802) & (!x13644x)) + ((!n_n4748) & (n_n4725) & (!n_n4788) & (!n_n4802) & (x13644x)) + ((!n_n4748) & (n_n4725) & (!n_n4788) & (n_n4802) & (!x13644x)) + ((!n_n4748) & (n_n4725) & (!n_n4788) & (n_n4802) & (x13644x)) + ((!n_n4748) & (n_n4725) & (n_n4788) & (!n_n4802) & (!x13644x)) + ((!n_n4748) & (n_n4725) & (n_n4788) & (!n_n4802) & (x13644x)) + ((!n_n4748) & (n_n4725) & (n_n4788) & (n_n4802) & (!x13644x)) + ((!n_n4748) & (n_n4725) & (n_n4788) & (n_n4802) & (x13644x)) + ((n_n4748) & (!n_n4725) & (!n_n4788) & (!n_n4802) & (!x13644x)) + ((n_n4748) & (!n_n4725) & (!n_n4788) & (!n_n4802) & (x13644x)) + ((n_n4748) & (!n_n4725) & (!n_n4788) & (n_n4802) & (!x13644x)) + ((n_n4748) & (!n_n4725) & (!n_n4788) & (n_n4802) & (x13644x)) + ((n_n4748) & (!n_n4725) & (n_n4788) & (!n_n4802) & (!x13644x)) + ((n_n4748) & (!n_n4725) & (n_n4788) & (!n_n4802) & (x13644x)) + ((n_n4748) & (!n_n4725) & (n_n4788) & (n_n4802) & (!x13644x)) + ((n_n4748) & (!n_n4725) & (n_n4788) & (n_n4802) & (x13644x)) + ((n_n4748) & (n_n4725) & (!n_n4788) & (!n_n4802) & (!x13644x)) + ((n_n4748) & (n_n4725) & (!n_n4788) & (!n_n4802) & (x13644x)) + ((n_n4748) & (n_n4725) & (!n_n4788) & (n_n4802) & (!x13644x)) + ((n_n4748) & (n_n4725) & (!n_n4788) & (n_n4802) & (x13644x)) + ((n_n4748) & (n_n4725) & (n_n4788) & (!n_n4802) & (!x13644x)) + ((n_n4748) & (n_n4725) & (n_n4788) & (!n_n4802) & (x13644x)) + ((n_n4748) & (n_n4725) & (n_n4788) & (n_n4802) & (!x13644x)) + ((n_n4748) & (n_n4725) & (n_n4788) & (n_n4802) & (x13644x)));
	assign x13646x = (((!x13630x) & (!x13631x) & (!x13636x) & (x13637x)) + ((!x13630x) & (!x13631x) & (x13636x) & (!x13637x)) + ((!x13630x) & (!x13631x) & (x13636x) & (x13637x)) + ((!x13630x) & (x13631x) & (!x13636x) & (!x13637x)) + ((!x13630x) & (x13631x) & (!x13636x) & (x13637x)) + ((!x13630x) & (x13631x) & (x13636x) & (!x13637x)) + ((!x13630x) & (x13631x) & (x13636x) & (x13637x)) + ((x13630x) & (!x13631x) & (!x13636x) & (!x13637x)) + ((x13630x) & (!x13631x) & (!x13636x) & (x13637x)) + ((x13630x) & (!x13631x) & (x13636x) & (!x13637x)) + ((x13630x) & (!x13631x) & (x13636x) & (x13637x)) + ((x13630x) & (x13631x) & (!x13636x) & (!x13637x)) + ((x13630x) & (x13631x) & (!x13636x) & (x13637x)) + ((x13630x) & (x13631x) & (x13636x) & (!x13637x)) + ((x13630x) & (x13631x) & (x13636x) & (x13637x)));
	assign n_n3921 = (((!x13650x) & (!x13651x) & (!n_n3932) & (!x13663x) & (x13664x)) + ((!x13650x) & (!x13651x) & (!n_n3932) & (x13663x) & (!x13664x)) + ((!x13650x) & (!x13651x) & (!n_n3932) & (x13663x) & (x13664x)) + ((!x13650x) & (!x13651x) & (n_n3932) & (!x13663x) & (!x13664x)) + ((!x13650x) & (!x13651x) & (n_n3932) & (!x13663x) & (x13664x)) + ((!x13650x) & (!x13651x) & (n_n3932) & (x13663x) & (!x13664x)) + ((!x13650x) & (!x13651x) & (n_n3932) & (x13663x) & (x13664x)) + ((!x13650x) & (x13651x) & (!n_n3932) & (!x13663x) & (!x13664x)) + ((!x13650x) & (x13651x) & (!n_n3932) & (!x13663x) & (x13664x)) + ((!x13650x) & (x13651x) & (!n_n3932) & (x13663x) & (!x13664x)) + ((!x13650x) & (x13651x) & (!n_n3932) & (x13663x) & (x13664x)) + ((!x13650x) & (x13651x) & (n_n3932) & (!x13663x) & (!x13664x)) + ((!x13650x) & (x13651x) & (n_n3932) & (!x13663x) & (x13664x)) + ((!x13650x) & (x13651x) & (n_n3932) & (x13663x) & (!x13664x)) + ((!x13650x) & (x13651x) & (n_n3932) & (x13663x) & (x13664x)) + ((x13650x) & (!x13651x) & (!n_n3932) & (!x13663x) & (!x13664x)) + ((x13650x) & (!x13651x) & (!n_n3932) & (!x13663x) & (x13664x)) + ((x13650x) & (!x13651x) & (!n_n3932) & (x13663x) & (!x13664x)) + ((x13650x) & (!x13651x) & (!n_n3932) & (x13663x) & (x13664x)) + ((x13650x) & (!x13651x) & (n_n3932) & (!x13663x) & (!x13664x)) + ((x13650x) & (!x13651x) & (n_n3932) & (!x13663x) & (x13664x)) + ((x13650x) & (!x13651x) & (n_n3932) & (x13663x) & (!x13664x)) + ((x13650x) & (!x13651x) & (n_n3932) & (x13663x) & (x13664x)) + ((x13650x) & (x13651x) & (!n_n3932) & (!x13663x) & (!x13664x)) + ((x13650x) & (x13651x) & (!n_n3932) & (!x13663x) & (x13664x)) + ((x13650x) & (x13651x) & (!n_n3932) & (x13663x) & (!x13664x)) + ((x13650x) & (x13651x) & (!n_n3932) & (x13663x) & (x13664x)) + ((x13650x) & (x13651x) & (n_n3932) & (!x13663x) & (!x13664x)) + ((x13650x) & (x13651x) & (n_n3932) & (!x13663x) & (x13664x)) + ((x13650x) & (x13651x) & (n_n3932) & (x13663x) & (!x13664x)) + ((x13650x) & (x13651x) & (n_n3932) & (x13663x) & (x13664x)));
	assign x13683x = (((!x13616x) & (!n_n3926) & (!n_n3924) & (!x13615x) & (x13681x)) + ((!x13616x) & (!n_n3926) & (!n_n3924) & (x13615x) & (!x13681x)) + ((!x13616x) & (!n_n3926) & (!n_n3924) & (x13615x) & (x13681x)) + ((!x13616x) & (!n_n3926) & (n_n3924) & (!x13615x) & (!x13681x)) + ((!x13616x) & (!n_n3926) & (n_n3924) & (!x13615x) & (x13681x)) + ((!x13616x) & (!n_n3926) & (n_n3924) & (x13615x) & (!x13681x)) + ((!x13616x) & (!n_n3926) & (n_n3924) & (x13615x) & (x13681x)) + ((!x13616x) & (n_n3926) & (!n_n3924) & (!x13615x) & (!x13681x)) + ((!x13616x) & (n_n3926) & (!n_n3924) & (!x13615x) & (x13681x)) + ((!x13616x) & (n_n3926) & (!n_n3924) & (x13615x) & (!x13681x)) + ((!x13616x) & (n_n3926) & (!n_n3924) & (x13615x) & (x13681x)) + ((!x13616x) & (n_n3926) & (n_n3924) & (!x13615x) & (!x13681x)) + ((!x13616x) & (n_n3926) & (n_n3924) & (!x13615x) & (x13681x)) + ((!x13616x) & (n_n3926) & (n_n3924) & (x13615x) & (!x13681x)) + ((!x13616x) & (n_n3926) & (n_n3924) & (x13615x) & (x13681x)) + ((x13616x) & (!n_n3926) & (!n_n3924) & (!x13615x) & (!x13681x)) + ((x13616x) & (!n_n3926) & (!n_n3924) & (!x13615x) & (x13681x)) + ((x13616x) & (!n_n3926) & (!n_n3924) & (x13615x) & (!x13681x)) + ((x13616x) & (!n_n3926) & (!n_n3924) & (x13615x) & (x13681x)) + ((x13616x) & (!n_n3926) & (n_n3924) & (!x13615x) & (!x13681x)) + ((x13616x) & (!n_n3926) & (n_n3924) & (!x13615x) & (x13681x)) + ((x13616x) & (!n_n3926) & (n_n3924) & (x13615x) & (!x13681x)) + ((x13616x) & (!n_n3926) & (n_n3924) & (x13615x) & (x13681x)) + ((x13616x) & (n_n3926) & (!n_n3924) & (!x13615x) & (!x13681x)) + ((x13616x) & (n_n3926) & (!n_n3924) & (!x13615x) & (x13681x)) + ((x13616x) & (n_n3926) & (!n_n3924) & (x13615x) & (!x13681x)) + ((x13616x) & (n_n3926) & (!n_n3924) & (x13615x) & (x13681x)) + ((x13616x) & (n_n3926) & (n_n3924) & (!x13615x) & (!x13681x)) + ((x13616x) & (n_n3926) & (n_n3924) & (!x13615x) & (x13681x)) + ((x13616x) & (n_n3926) & (n_n3924) & (x13615x) & (!x13681x)) + ((x13616x) & (n_n3926) & (n_n3924) & (x13615x) & (x13681x)));
	assign n_n3192 = (((!x13761x) & (!x13747x) & (!x13748x) & (!x13753x) & (x13754x)) + ((!x13761x) & (!x13747x) & (!x13748x) & (x13753x) & (!x13754x)) + ((!x13761x) & (!x13747x) & (!x13748x) & (x13753x) & (x13754x)) + ((!x13761x) & (!x13747x) & (x13748x) & (!x13753x) & (!x13754x)) + ((!x13761x) & (!x13747x) & (x13748x) & (!x13753x) & (x13754x)) + ((!x13761x) & (!x13747x) & (x13748x) & (x13753x) & (!x13754x)) + ((!x13761x) & (!x13747x) & (x13748x) & (x13753x) & (x13754x)) + ((!x13761x) & (x13747x) & (!x13748x) & (!x13753x) & (!x13754x)) + ((!x13761x) & (x13747x) & (!x13748x) & (!x13753x) & (x13754x)) + ((!x13761x) & (x13747x) & (!x13748x) & (x13753x) & (!x13754x)) + ((!x13761x) & (x13747x) & (!x13748x) & (x13753x) & (x13754x)) + ((!x13761x) & (x13747x) & (x13748x) & (!x13753x) & (!x13754x)) + ((!x13761x) & (x13747x) & (x13748x) & (!x13753x) & (x13754x)) + ((!x13761x) & (x13747x) & (x13748x) & (x13753x) & (!x13754x)) + ((!x13761x) & (x13747x) & (x13748x) & (x13753x) & (x13754x)) + ((x13761x) & (!x13747x) & (!x13748x) & (!x13753x) & (!x13754x)) + ((x13761x) & (!x13747x) & (!x13748x) & (!x13753x) & (x13754x)) + ((x13761x) & (!x13747x) & (!x13748x) & (x13753x) & (!x13754x)) + ((x13761x) & (!x13747x) & (!x13748x) & (x13753x) & (x13754x)) + ((x13761x) & (!x13747x) & (x13748x) & (!x13753x) & (!x13754x)) + ((x13761x) & (!x13747x) & (x13748x) & (!x13753x) & (x13754x)) + ((x13761x) & (!x13747x) & (x13748x) & (x13753x) & (!x13754x)) + ((x13761x) & (!x13747x) & (x13748x) & (x13753x) & (x13754x)) + ((x13761x) & (x13747x) & (!x13748x) & (!x13753x) & (!x13754x)) + ((x13761x) & (x13747x) & (!x13748x) & (!x13753x) & (x13754x)) + ((x13761x) & (x13747x) & (!x13748x) & (x13753x) & (!x13754x)) + ((x13761x) & (x13747x) & (!x13748x) & (x13753x) & (x13754x)) + ((x13761x) & (x13747x) & (x13748x) & (!x13753x) & (!x13754x)) + ((x13761x) & (x13747x) & (x13748x) & (!x13753x) & (x13754x)) + ((x13761x) & (x13747x) & (x13748x) & (x13753x) & (!x13754x)) + ((x13761x) & (x13747x) & (x13748x) & (x13753x) & (x13754x)));
	assign x13782x = (((!n_n4853) & (!n_n4847) & (!n_n4864) & (!n_n4912) & (x13781x)) + ((!n_n4853) & (!n_n4847) & (!n_n4864) & (n_n4912) & (!x13781x)) + ((!n_n4853) & (!n_n4847) & (!n_n4864) & (n_n4912) & (x13781x)) + ((!n_n4853) & (!n_n4847) & (n_n4864) & (!n_n4912) & (!x13781x)) + ((!n_n4853) & (!n_n4847) & (n_n4864) & (!n_n4912) & (x13781x)) + ((!n_n4853) & (!n_n4847) & (n_n4864) & (n_n4912) & (!x13781x)) + ((!n_n4853) & (!n_n4847) & (n_n4864) & (n_n4912) & (x13781x)) + ((!n_n4853) & (n_n4847) & (!n_n4864) & (!n_n4912) & (!x13781x)) + ((!n_n4853) & (n_n4847) & (!n_n4864) & (!n_n4912) & (x13781x)) + ((!n_n4853) & (n_n4847) & (!n_n4864) & (n_n4912) & (!x13781x)) + ((!n_n4853) & (n_n4847) & (!n_n4864) & (n_n4912) & (x13781x)) + ((!n_n4853) & (n_n4847) & (n_n4864) & (!n_n4912) & (!x13781x)) + ((!n_n4853) & (n_n4847) & (n_n4864) & (!n_n4912) & (x13781x)) + ((!n_n4853) & (n_n4847) & (n_n4864) & (n_n4912) & (!x13781x)) + ((!n_n4853) & (n_n4847) & (n_n4864) & (n_n4912) & (x13781x)) + ((n_n4853) & (!n_n4847) & (!n_n4864) & (!n_n4912) & (!x13781x)) + ((n_n4853) & (!n_n4847) & (!n_n4864) & (!n_n4912) & (x13781x)) + ((n_n4853) & (!n_n4847) & (!n_n4864) & (n_n4912) & (!x13781x)) + ((n_n4853) & (!n_n4847) & (!n_n4864) & (n_n4912) & (x13781x)) + ((n_n4853) & (!n_n4847) & (n_n4864) & (!n_n4912) & (!x13781x)) + ((n_n4853) & (!n_n4847) & (n_n4864) & (!n_n4912) & (x13781x)) + ((n_n4853) & (!n_n4847) & (n_n4864) & (n_n4912) & (!x13781x)) + ((n_n4853) & (!n_n4847) & (n_n4864) & (n_n4912) & (x13781x)) + ((n_n4853) & (n_n4847) & (!n_n4864) & (!n_n4912) & (!x13781x)) + ((n_n4853) & (n_n4847) & (!n_n4864) & (!n_n4912) & (x13781x)) + ((n_n4853) & (n_n4847) & (!n_n4864) & (n_n4912) & (!x13781x)) + ((n_n4853) & (n_n4847) & (!n_n4864) & (n_n4912) & (x13781x)) + ((n_n4853) & (n_n4847) & (n_n4864) & (!n_n4912) & (!x13781x)) + ((n_n4853) & (n_n4847) & (n_n4864) & (!n_n4912) & (x13781x)) + ((n_n4853) & (n_n4847) & (n_n4864) & (n_n4912) & (!x13781x)) + ((n_n4853) & (n_n4847) & (n_n4864) & (n_n4912) & (x13781x)));
	assign x13783x = (((!x13767x) & (!x13768x) & (!x13773x) & (x13774x)) + ((!x13767x) & (!x13768x) & (x13773x) & (!x13774x)) + ((!x13767x) & (!x13768x) & (x13773x) & (x13774x)) + ((!x13767x) & (x13768x) & (!x13773x) & (!x13774x)) + ((!x13767x) & (x13768x) & (!x13773x) & (x13774x)) + ((!x13767x) & (x13768x) & (x13773x) & (!x13774x)) + ((!x13767x) & (x13768x) & (x13773x) & (x13774x)) + ((x13767x) & (!x13768x) & (!x13773x) & (!x13774x)) + ((x13767x) & (!x13768x) & (!x13773x) & (x13774x)) + ((x13767x) & (!x13768x) & (x13773x) & (!x13774x)) + ((x13767x) & (!x13768x) & (x13773x) & (x13774x)) + ((x13767x) & (x13768x) & (!x13773x) & (!x13774x)) + ((x13767x) & (x13768x) & (!x13773x) & (x13774x)) + ((x13767x) & (x13768x) & (x13773x) & (!x13774x)) + ((x13767x) & (x13768x) & (x13773x) & (x13774x)));
	assign x14221x = (((!n_n3189) & (!n_n3205) & (!x13728x) & (!x13729x) & (x14218x)) + ((!n_n3189) & (!n_n3205) & (!x13728x) & (x13729x) & (!x14218x)) + ((!n_n3189) & (!n_n3205) & (!x13728x) & (x13729x) & (x14218x)) + ((!n_n3189) & (!n_n3205) & (x13728x) & (!x13729x) & (!x14218x)) + ((!n_n3189) & (!n_n3205) & (x13728x) & (!x13729x) & (x14218x)) + ((!n_n3189) & (!n_n3205) & (x13728x) & (x13729x) & (!x14218x)) + ((!n_n3189) & (!n_n3205) & (x13728x) & (x13729x) & (x14218x)) + ((!n_n3189) & (n_n3205) & (!x13728x) & (!x13729x) & (!x14218x)) + ((!n_n3189) & (n_n3205) & (!x13728x) & (!x13729x) & (x14218x)) + ((!n_n3189) & (n_n3205) & (!x13728x) & (x13729x) & (!x14218x)) + ((!n_n3189) & (n_n3205) & (!x13728x) & (x13729x) & (x14218x)) + ((!n_n3189) & (n_n3205) & (x13728x) & (!x13729x) & (!x14218x)) + ((!n_n3189) & (n_n3205) & (x13728x) & (!x13729x) & (x14218x)) + ((!n_n3189) & (n_n3205) & (x13728x) & (x13729x) & (!x14218x)) + ((!n_n3189) & (n_n3205) & (x13728x) & (x13729x) & (x14218x)) + ((n_n3189) & (!n_n3205) & (!x13728x) & (!x13729x) & (!x14218x)) + ((n_n3189) & (!n_n3205) & (!x13728x) & (!x13729x) & (x14218x)) + ((n_n3189) & (!n_n3205) & (!x13728x) & (x13729x) & (!x14218x)) + ((n_n3189) & (!n_n3205) & (!x13728x) & (x13729x) & (x14218x)) + ((n_n3189) & (!n_n3205) & (x13728x) & (!x13729x) & (!x14218x)) + ((n_n3189) & (!n_n3205) & (x13728x) & (!x13729x) & (x14218x)) + ((n_n3189) & (!n_n3205) & (x13728x) & (x13729x) & (!x14218x)) + ((n_n3189) & (!n_n3205) & (x13728x) & (x13729x) & (x14218x)) + ((n_n3189) & (n_n3205) & (!x13728x) & (!x13729x) & (!x14218x)) + ((n_n3189) & (n_n3205) & (!x13728x) & (!x13729x) & (x14218x)) + ((n_n3189) & (n_n3205) & (!x13728x) & (x13729x) & (!x14218x)) + ((n_n3189) & (n_n3205) & (!x13728x) & (x13729x) & (x14218x)) + ((n_n3189) & (n_n3205) & (x13728x) & (!x13729x) & (!x14218x)) + ((n_n3189) & (n_n3205) & (x13728x) & (!x13729x) & (x14218x)) + ((n_n3189) & (n_n3205) & (x13728x) & (x13729x) & (!x14218x)) + ((n_n3189) & (n_n3205) & (x13728x) & (x13729x) & (x14218x)));
	assign x14540x = (((!n_n3653) & (!x14530x) & (!n_n3729) & (!n_n3731) & (x14538x)) + ((!n_n3653) & (!x14530x) & (!n_n3729) & (n_n3731) & (!x14538x)) + ((!n_n3653) & (!x14530x) & (!n_n3729) & (n_n3731) & (x14538x)) + ((!n_n3653) & (!x14530x) & (n_n3729) & (!n_n3731) & (!x14538x)) + ((!n_n3653) & (!x14530x) & (n_n3729) & (!n_n3731) & (x14538x)) + ((!n_n3653) & (!x14530x) & (n_n3729) & (n_n3731) & (!x14538x)) + ((!n_n3653) & (!x14530x) & (n_n3729) & (n_n3731) & (x14538x)) + ((!n_n3653) & (x14530x) & (!n_n3729) & (!n_n3731) & (!x14538x)) + ((!n_n3653) & (x14530x) & (!n_n3729) & (!n_n3731) & (x14538x)) + ((!n_n3653) & (x14530x) & (!n_n3729) & (n_n3731) & (!x14538x)) + ((!n_n3653) & (x14530x) & (!n_n3729) & (n_n3731) & (x14538x)) + ((!n_n3653) & (x14530x) & (n_n3729) & (!n_n3731) & (!x14538x)) + ((!n_n3653) & (x14530x) & (n_n3729) & (!n_n3731) & (x14538x)) + ((!n_n3653) & (x14530x) & (n_n3729) & (n_n3731) & (!x14538x)) + ((!n_n3653) & (x14530x) & (n_n3729) & (n_n3731) & (x14538x)) + ((n_n3653) & (!x14530x) & (!n_n3729) & (!n_n3731) & (!x14538x)) + ((n_n3653) & (!x14530x) & (!n_n3729) & (!n_n3731) & (x14538x)) + ((n_n3653) & (!x14530x) & (!n_n3729) & (n_n3731) & (!x14538x)) + ((n_n3653) & (!x14530x) & (!n_n3729) & (n_n3731) & (x14538x)) + ((n_n3653) & (!x14530x) & (n_n3729) & (!n_n3731) & (!x14538x)) + ((n_n3653) & (!x14530x) & (n_n3729) & (!n_n3731) & (x14538x)) + ((n_n3653) & (!x14530x) & (n_n3729) & (n_n3731) & (!x14538x)) + ((n_n3653) & (!x14530x) & (n_n3729) & (n_n3731) & (x14538x)) + ((n_n3653) & (x14530x) & (!n_n3729) & (!n_n3731) & (!x14538x)) + ((n_n3653) & (x14530x) & (!n_n3729) & (!n_n3731) & (x14538x)) + ((n_n3653) & (x14530x) & (!n_n3729) & (n_n3731) & (!x14538x)) + ((n_n3653) & (x14530x) & (!n_n3729) & (n_n3731) & (x14538x)) + ((n_n3653) & (x14530x) & (n_n3729) & (!n_n3731) & (!x14538x)) + ((n_n3653) & (x14530x) & (n_n3729) & (!n_n3731) & (x14538x)) + ((n_n3653) & (x14530x) & (n_n3729) & (n_n3731) & (!x14538x)) + ((n_n3653) & (x14530x) & (n_n3729) & (n_n3731) & (x14538x)));
	assign n_n3625 = (((!n_n3638) & (!n_n3639) & (!n_n3685) & (!n_n3686) & (x14682x)) + ((!n_n3638) & (!n_n3639) & (!n_n3685) & (n_n3686) & (!x14682x)) + ((!n_n3638) & (!n_n3639) & (!n_n3685) & (n_n3686) & (x14682x)) + ((!n_n3638) & (!n_n3639) & (n_n3685) & (!n_n3686) & (!x14682x)) + ((!n_n3638) & (!n_n3639) & (n_n3685) & (!n_n3686) & (x14682x)) + ((!n_n3638) & (!n_n3639) & (n_n3685) & (n_n3686) & (!x14682x)) + ((!n_n3638) & (!n_n3639) & (n_n3685) & (n_n3686) & (x14682x)) + ((!n_n3638) & (n_n3639) & (!n_n3685) & (!n_n3686) & (!x14682x)) + ((!n_n3638) & (n_n3639) & (!n_n3685) & (!n_n3686) & (x14682x)) + ((!n_n3638) & (n_n3639) & (!n_n3685) & (n_n3686) & (!x14682x)) + ((!n_n3638) & (n_n3639) & (!n_n3685) & (n_n3686) & (x14682x)) + ((!n_n3638) & (n_n3639) & (n_n3685) & (!n_n3686) & (!x14682x)) + ((!n_n3638) & (n_n3639) & (n_n3685) & (!n_n3686) & (x14682x)) + ((!n_n3638) & (n_n3639) & (n_n3685) & (n_n3686) & (!x14682x)) + ((!n_n3638) & (n_n3639) & (n_n3685) & (n_n3686) & (x14682x)) + ((n_n3638) & (!n_n3639) & (!n_n3685) & (!n_n3686) & (!x14682x)) + ((n_n3638) & (!n_n3639) & (!n_n3685) & (!n_n3686) & (x14682x)) + ((n_n3638) & (!n_n3639) & (!n_n3685) & (n_n3686) & (!x14682x)) + ((n_n3638) & (!n_n3639) & (!n_n3685) & (n_n3686) & (x14682x)) + ((n_n3638) & (!n_n3639) & (n_n3685) & (!n_n3686) & (!x14682x)) + ((n_n3638) & (!n_n3639) & (n_n3685) & (!n_n3686) & (x14682x)) + ((n_n3638) & (!n_n3639) & (n_n3685) & (n_n3686) & (!x14682x)) + ((n_n3638) & (!n_n3639) & (n_n3685) & (n_n3686) & (x14682x)) + ((n_n3638) & (n_n3639) & (!n_n3685) & (!n_n3686) & (!x14682x)) + ((n_n3638) & (n_n3639) & (!n_n3685) & (!n_n3686) & (x14682x)) + ((n_n3638) & (n_n3639) & (!n_n3685) & (n_n3686) & (!x14682x)) + ((n_n3638) & (n_n3639) & (!n_n3685) & (n_n3686) & (x14682x)) + ((n_n3638) & (n_n3639) & (n_n3685) & (!n_n3686) & (!x14682x)) + ((n_n3638) & (n_n3639) & (n_n3685) & (!n_n3686) & (x14682x)) + ((n_n3638) & (n_n3639) & (n_n3685) & (n_n3686) & (!x14682x)) + ((n_n3638) & (n_n3639) & (n_n3685) & (n_n3686) & (x14682x)));
	assign n_n3627 = (((!x14730x) & (!n_n3645) & (!n_n3702) & (!x14722x) & (x14721x)) + ((!x14730x) & (!n_n3645) & (!n_n3702) & (x14722x) & (!x14721x)) + ((!x14730x) & (!n_n3645) & (!n_n3702) & (x14722x) & (x14721x)) + ((!x14730x) & (!n_n3645) & (n_n3702) & (!x14722x) & (!x14721x)) + ((!x14730x) & (!n_n3645) & (n_n3702) & (!x14722x) & (x14721x)) + ((!x14730x) & (!n_n3645) & (n_n3702) & (x14722x) & (!x14721x)) + ((!x14730x) & (!n_n3645) & (n_n3702) & (x14722x) & (x14721x)) + ((!x14730x) & (n_n3645) & (!n_n3702) & (!x14722x) & (!x14721x)) + ((!x14730x) & (n_n3645) & (!n_n3702) & (!x14722x) & (x14721x)) + ((!x14730x) & (n_n3645) & (!n_n3702) & (x14722x) & (!x14721x)) + ((!x14730x) & (n_n3645) & (!n_n3702) & (x14722x) & (x14721x)) + ((!x14730x) & (n_n3645) & (n_n3702) & (!x14722x) & (!x14721x)) + ((!x14730x) & (n_n3645) & (n_n3702) & (!x14722x) & (x14721x)) + ((!x14730x) & (n_n3645) & (n_n3702) & (x14722x) & (!x14721x)) + ((!x14730x) & (n_n3645) & (n_n3702) & (x14722x) & (x14721x)) + ((x14730x) & (!n_n3645) & (!n_n3702) & (!x14722x) & (!x14721x)) + ((x14730x) & (!n_n3645) & (!n_n3702) & (!x14722x) & (x14721x)) + ((x14730x) & (!n_n3645) & (!n_n3702) & (x14722x) & (!x14721x)) + ((x14730x) & (!n_n3645) & (!n_n3702) & (x14722x) & (x14721x)) + ((x14730x) & (!n_n3645) & (n_n3702) & (!x14722x) & (!x14721x)) + ((x14730x) & (!n_n3645) & (n_n3702) & (!x14722x) & (x14721x)) + ((x14730x) & (!n_n3645) & (n_n3702) & (x14722x) & (!x14721x)) + ((x14730x) & (!n_n3645) & (n_n3702) & (x14722x) & (x14721x)) + ((x14730x) & (n_n3645) & (!n_n3702) & (!x14722x) & (!x14721x)) + ((x14730x) & (n_n3645) & (!n_n3702) & (!x14722x) & (x14721x)) + ((x14730x) & (n_n3645) & (!n_n3702) & (x14722x) & (!x14721x)) + ((x14730x) & (n_n3645) & (!n_n3702) & (x14722x) & (x14721x)) + ((x14730x) & (n_n3645) & (n_n3702) & (!x14722x) & (!x14721x)) + ((x14730x) & (n_n3645) & (n_n3702) & (!x14722x) & (x14721x)) + ((x14730x) & (n_n3645) & (n_n3702) & (x14722x) & (!x14721x)) + ((x14730x) & (n_n3645) & (n_n3702) & (x14722x) & (x14721x)));
	assign n_n3629 = (((!n_n3650) & (!n_n3652) & (x14436x)) + ((!n_n3650) & (n_n3652) & (!x14436x)) + ((!n_n3650) & (n_n3652) & (x14436x)) + ((n_n3650) & (!n_n3652) & (!x14436x)) + ((n_n3650) & (!n_n3652) & (x14436x)) + ((n_n3650) & (n_n3652) & (!x14436x)) + ((n_n3650) & (n_n3652) & (x14436x)));
	assign n_n3631 = (((!x14513x) & (!n_n3658) & (!x14507x) & (!n_n3732) & (n_n3734)) + ((!x14513x) & (!n_n3658) & (!x14507x) & (n_n3732) & (!n_n3734)) + ((!x14513x) & (!n_n3658) & (!x14507x) & (n_n3732) & (n_n3734)) + ((!x14513x) & (!n_n3658) & (x14507x) & (!n_n3732) & (!n_n3734)) + ((!x14513x) & (!n_n3658) & (x14507x) & (!n_n3732) & (n_n3734)) + ((!x14513x) & (!n_n3658) & (x14507x) & (n_n3732) & (!n_n3734)) + ((!x14513x) & (!n_n3658) & (x14507x) & (n_n3732) & (n_n3734)) + ((!x14513x) & (n_n3658) & (!x14507x) & (!n_n3732) & (!n_n3734)) + ((!x14513x) & (n_n3658) & (!x14507x) & (!n_n3732) & (n_n3734)) + ((!x14513x) & (n_n3658) & (!x14507x) & (n_n3732) & (!n_n3734)) + ((!x14513x) & (n_n3658) & (!x14507x) & (n_n3732) & (n_n3734)) + ((!x14513x) & (n_n3658) & (x14507x) & (!n_n3732) & (!n_n3734)) + ((!x14513x) & (n_n3658) & (x14507x) & (!n_n3732) & (n_n3734)) + ((!x14513x) & (n_n3658) & (x14507x) & (n_n3732) & (!n_n3734)) + ((!x14513x) & (n_n3658) & (x14507x) & (n_n3732) & (n_n3734)) + ((x14513x) & (!n_n3658) & (!x14507x) & (!n_n3732) & (!n_n3734)) + ((x14513x) & (!n_n3658) & (!x14507x) & (!n_n3732) & (n_n3734)) + ((x14513x) & (!n_n3658) & (!x14507x) & (n_n3732) & (!n_n3734)) + ((x14513x) & (!n_n3658) & (!x14507x) & (n_n3732) & (n_n3734)) + ((x14513x) & (!n_n3658) & (x14507x) & (!n_n3732) & (!n_n3734)) + ((x14513x) & (!n_n3658) & (x14507x) & (!n_n3732) & (n_n3734)) + ((x14513x) & (!n_n3658) & (x14507x) & (n_n3732) & (!n_n3734)) + ((x14513x) & (!n_n3658) & (x14507x) & (n_n3732) & (n_n3734)) + ((x14513x) & (n_n3658) & (!x14507x) & (!n_n3732) & (!n_n3734)) + ((x14513x) & (n_n3658) & (!x14507x) & (!n_n3732) & (n_n3734)) + ((x14513x) & (n_n3658) & (!x14507x) & (n_n3732) & (!n_n3734)) + ((x14513x) & (n_n3658) & (!x14507x) & (n_n3732) & (n_n3734)) + ((x14513x) & (n_n3658) & (x14507x) & (!n_n3732) & (!n_n3734)) + ((x14513x) & (n_n3658) & (x14507x) & (!n_n3732) & (n_n3734)) + ((x14513x) & (n_n3658) & (x14507x) & (n_n3732) & (!n_n3734)) + ((x14513x) & (n_n3658) & (x14507x) & (n_n3732) & (n_n3734)));
	assign n_n2530 = (((!n_n2548) & (!n_n2598) & (!n_n2597) & (!n_n2549) & (x14933x)) + ((!n_n2548) & (!n_n2598) & (!n_n2597) & (n_n2549) & (!x14933x)) + ((!n_n2548) & (!n_n2598) & (!n_n2597) & (n_n2549) & (x14933x)) + ((!n_n2548) & (!n_n2598) & (n_n2597) & (!n_n2549) & (!x14933x)) + ((!n_n2548) & (!n_n2598) & (n_n2597) & (!n_n2549) & (x14933x)) + ((!n_n2548) & (!n_n2598) & (n_n2597) & (n_n2549) & (!x14933x)) + ((!n_n2548) & (!n_n2598) & (n_n2597) & (n_n2549) & (x14933x)) + ((!n_n2548) & (n_n2598) & (!n_n2597) & (!n_n2549) & (!x14933x)) + ((!n_n2548) & (n_n2598) & (!n_n2597) & (!n_n2549) & (x14933x)) + ((!n_n2548) & (n_n2598) & (!n_n2597) & (n_n2549) & (!x14933x)) + ((!n_n2548) & (n_n2598) & (!n_n2597) & (n_n2549) & (x14933x)) + ((!n_n2548) & (n_n2598) & (n_n2597) & (!n_n2549) & (!x14933x)) + ((!n_n2548) & (n_n2598) & (n_n2597) & (!n_n2549) & (x14933x)) + ((!n_n2548) & (n_n2598) & (n_n2597) & (n_n2549) & (!x14933x)) + ((!n_n2548) & (n_n2598) & (n_n2597) & (n_n2549) & (x14933x)) + ((n_n2548) & (!n_n2598) & (!n_n2597) & (!n_n2549) & (!x14933x)) + ((n_n2548) & (!n_n2598) & (!n_n2597) & (!n_n2549) & (x14933x)) + ((n_n2548) & (!n_n2598) & (!n_n2597) & (n_n2549) & (!x14933x)) + ((n_n2548) & (!n_n2598) & (!n_n2597) & (n_n2549) & (x14933x)) + ((n_n2548) & (!n_n2598) & (n_n2597) & (!n_n2549) & (!x14933x)) + ((n_n2548) & (!n_n2598) & (n_n2597) & (!n_n2549) & (x14933x)) + ((n_n2548) & (!n_n2598) & (n_n2597) & (n_n2549) & (!x14933x)) + ((n_n2548) & (!n_n2598) & (n_n2597) & (n_n2549) & (x14933x)) + ((n_n2548) & (n_n2598) & (!n_n2597) & (!n_n2549) & (!x14933x)) + ((n_n2548) & (n_n2598) & (!n_n2597) & (!n_n2549) & (x14933x)) + ((n_n2548) & (n_n2598) & (!n_n2597) & (n_n2549) & (!x14933x)) + ((n_n2548) & (n_n2598) & (!n_n2597) & (n_n2549) & (x14933x)) + ((n_n2548) & (n_n2598) & (n_n2597) & (!n_n2549) & (!x14933x)) + ((n_n2548) & (n_n2598) & (n_n2597) & (!n_n2549) & (x14933x)) + ((n_n2548) & (n_n2598) & (n_n2597) & (n_n2549) & (!x14933x)) + ((n_n2548) & (n_n2598) & (n_n2597) & (n_n2549) & (x14933x)));
	assign n_n2529 = (((!n_n2589) & (!n_n2588) & (!n_n2546) & (!n_n2545) & (x14979x)) + ((!n_n2589) & (!n_n2588) & (!n_n2546) & (n_n2545) & (!x14979x)) + ((!n_n2589) & (!n_n2588) & (!n_n2546) & (n_n2545) & (x14979x)) + ((!n_n2589) & (!n_n2588) & (n_n2546) & (!n_n2545) & (!x14979x)) + ((!n_n2589) & (!n_n2588) & (n_n2546) & (!n_n2545) & (x14979x)) + ((!n_n2589) & (!n_n2588) & (n_n2546) & (n_n2545) & (!x14979x)) + ((!n_n2589) & (!n_n2588) & (n_n2546) & (n_n2545) & (x14979x)) + ((!n_n2589) & (n_n2588) & (!n_n2546) & (!n_n2545) & (!x14979x)) + ((!n_n2589) & (n_n2588) & (!n_n2546) & (!n_n2545) & (x14979x)) + ((!n_n2589) & (n_n2588) & (!n_n2546) & (n_n2545) & (!x14979x)) + ((!n_n2589) & (n_n2588) & (!n_n2546) & (n_n2545) & (x14979x)) + ((!n_n2589) & (n_n2588) & (n_n2546) & (!n_n2545) & (!x14979x)) + ((!n_n2589) & (n_n2588) & (n_n2546) & (!n_n2545) & (x14979x)) + ((!n_n2589) & (n_n2588) & (n_n2546) & (n_n2545) & (!x14979x)) + ((!n_n2589) & (n_n2588) & (n_n2546) & (n_n2545) & (x14979x)) + ((n_n2589) & (!n_n2588) & (!n_n2546) & (!n_n2545) & (!x14979x)) + ((n_n2589) & (!n_n2588) & (!n_n2546) & (!n_n2545) & (x14979x)) + ((n_n2589) & (!n_n2588) & (!n_n2546) & (n_n2545) & (!x14979x)) + ((n_n2589) & (!n_n2588) & (!n_n2546) & (n_n2545) & (x14979x)) + ((n_n2589) & (!n_n2588) & (n_n2546) & (!n_n2545) & (!x14979x)) + ((n_n2589) & (!n_n2588) & (n_n2546) & (!n_n2545) & (x14979x)) + ((n_n2589) & (!n_n2588) & (n_n2546) & (n_n2545) & (!x14979x)) + ((n_n2589) & (!n_n2588) & (n_n2546) & (n_n2545) & (x14979x)) + ((n_n2589) & (n_n2588) & (!n_n2546) & (!n_n2545) & (!x14979x)) + ((n_n2589) & (n_n2588) & (!n_n2546) & (!n_n2545) & (x14979x)) + ((n_n2589) & (n_n2588) & (!n_n2546) & (n_n2545) & (!x14979x)) + ((n_n2589) & (n_n2588) & (!n_n2546) & (n_n2545) & (x14979x)) + ((n_n2589) & (n_n2588) & (n_n2546) & (!n_n2545) & (!x14979x)) + ((n_n2589) & (n_n2588) & (n_n2546) & (!n_n2545) & (x14979x)) + ((n_n2589) & (n_n2588) & (n_n2546) & (n_n2545) & (!x14979x)) + ((n_n2589) & (n_n2588) & (n_n2546) & (n_n2545) & (x14979x)));
	assign x15169x = (((!n_n2560) & (!n_n2559) & (x15167x)) + ((!n_n2560) & (n_n2559) & (!x15167x)) + ((!n_n2560) & (n_n2559) & (x15167x)) + ((n_n2560) & (!n_n2559) & (!x15167x)) + ((n_n2560) & (!n_n2559) & (x15167x)) + ((n_n2560) & (n_n2559) & (!x15167x)) + ((n_n2560) & (n_n2559) & (x15167x)));
	assign n_n2533 = (((!n_n2558) & (!n_n2557) & (x15103x)) + ((!n_n2558) & (n_n2557) & (!x15103x)) + ((!n_n2558) & (n_n2557) & (x15103x)) + ((n_n2558) & (!n_n2557) & (!x15103x)) + ((n_n2558) & (!n_n2557) & (x15103x)) + ((n_n2558) & (n_n2557) & (!x15103x)) + ((n_n2558) & (n_n2557) & (x15103x)));
	assign n_n2532 = (((!n_n2554) & (!n_n2553) & (x15150x)) + ((!n_n2554) & (n_n2553) & (!x15150x)) + ((!n_n2554) & (n_n2553) & (x15150x)) + ((n_n2554) & (!n_n2553) & (!x15150x)) + ((n_n2554) & (!n_n2553) & (x15150x)) + ((n_n2554) & (n_n2553) & (!x15150x)) + ((n_n2554) & (n_n2553) & (x15150x)));
	assign n_n2906 = (((!x15503x) & (!n_n2990) & (!n_n2991) & (!n_n2926) & (x15494x)) + ((!x15503x) & (!n_n2990) & (!n_n2991) & (n_n2926) & (!x15494x)) + ((!x15503x) & (!n_n2990) & (!n_n2991) & (n_n2926) & (x15494x)) + ((!x15503x) & (!n_n2990) & (n_n2991) & (!n_n2926) & (!x15494x)) + ((!x15503x) & (!n_n2990) & (n_n2991) & (!n_n2926) & (x15494x)) + ((!x15503x) & (!n_n2990) & (n_n2991) & (n_n2926) & (!x15494x)) + ((!x15503x) & (!n_n2990) & (n_n2991) & (n_n2926) & (x15494x)) + ((!x15503x) & (n_n2990) & (!n_n2991) & (!n_n2926) & (!x15494x)) + ((!x15503x) & (n_n2990) & (!n_n2991) & (!n_n2926) & (x15494x)) + ((!x15503x) & (n_n2990) & (!n_n2991) & (n_n2926) & (!x15494x)) + ((!x15503x) & (n_n2990) & (!n_n2991) & (n_n2926) & (x15494x)) + ((!x15503x) & (n_n2990) & (n_n2991) & (!n_n2926) & (!x15494x)) + ((!x15503x) & (n_n2990) & (n_n2991) & (!n_n2926) & (x15494x)) + ((!x15503x) & (n_n2990) & (n_n2991) & (n_n2926) & (!x15494x)) + ((!x15503x) & (n_n2990) & (n_n2991) & (n_n2926) & (x15494x)) + ((x15503x) & (!n_n2990) & (!n_n2991) & (!n_n2926) & (!x15494x)) + ((x15503x) & (!n_n2990) & (!n_n2991) & (!n_n2926) & (x15494x)) + ((x15503x) & (!n_n2990) & (!n_n2991) & (n_n2926) & (!x15494x)) + ((x15503x) & (!n_n2990) & (!n_n2991) & (n_n2926) & (x15494x)) + ((x15503x) & (!n_n2990) & (n_n2991) & (!n_n2926) & (!x15494x)) + ((x15503x) & (!n_n2990) & (n_n2991) & (!n_n2926) & (x15494x)) + ((x15503x) & (!n_n2990) & (n_n2991) & (n_n2926) & (!x15494x)) + ((x15503x) & (!n_n2990) & (n_n2991) & (n_n2926) & (x15494x)) + ((x15503x) & (n_n2990) & (!n_n2991) & (!n_n2926) & (!x15494x)) + ((x15503x) & (n_n2990) & (!n_n2991) & (!n_n2926) & (x15494x)) + ((x15503x) & (n_n2990) & (!n_n2991) & (n_n2926) & (!x15494x)) + ((x15503x) & (n_n2990) & (!n_n2991) & (n_n2926) & (x15494x)) + ((x15503x) & (n_n2990) & (n_n2991) & (!n_n2926) & (!x15494x)) + ((x15503x) & (n_n2990) & (n_n2991) & (!n_n2926) & (x15494x)) + ((x15503x) & (n_n2990) & (n_n2991) & (n_n2926) & (!x15494x)) + ((x15503x) & (n_n2990) & (n_n2991) & (n_n2926) & (x15494x)));
	assign n_n2908 = (((!x15549x) & (!n_n2934) & (!n_n3004) & (!n_n3005) & (x15543x)) + ((!x15549x) & (!n_n2934) & (!n_n3004) & (n_n3005) & (!x15543x)) + ((!x15549x) & (!n_n2934) & (!n_n3004) & (n_n3005) & (x15543x)) + ((!x15549x) & (!n_n2934) & (n_n3004) & (!n_n3005) & (!x15543x)) + ((!x15549x) & (!n_n2934) & (n_n3004) & (!n_n3005) & (x15543x)) + ((!x15549x) & (!n_n2934) & (n_n3004) & (n_n3005) & (!x15543x)) + ((!x15549x) & (!n_n2934) & (n_n3004) & (n_n3005) & (x15543x)) + ((!x15549x) & (n_n2934) & (!n_n3004) & (!n_n3005) & (!x15543x)) + ((!x15549x) & (n_n2934) & (!n_n3004) & (!n_n3005) & (x15543x)) + ((!x15549x) & (n_n2934) & (!n_n3004) & (n_n3005) & (!x15543x)) + ((!x15549x) & (n_n2934) & (!n_n3004) & (n_n3005) & (x15543x)) + ((!x15549x) & (n_n2934) & (n_n3004) & (!n_n3005) & (!x15543x)) + ((!x15549x) & (n_n2934) & (n_n3004) & (!n_n3005) & (x15543x)) + ((!x15549x) & (n_n2934) & (n_n3004) & (n_n3005) & (!x15543x)) + ((!x15549x) & (n_n2934) & (n_n3004) & (n_n3005) & (x15543x)) + ((x15549x) & (!n_n2934) & (!n_n3004) & (!n_n3005) & (!x15543x)) + ((x15549x) & (!n_n2934) & (!n_n3004) & (!n_n3005) & (x15543x)) + ((x15549x) & (!n_n2934) & (!n_n3004) & (n_n3005) & (!x15543x)) + ((x15549x) & (!n_n2934) & (!n_n3004) & (n_n3005) & (x15543x)) + ((x15549x) & (!n_n2934) & (n_n3004) & (!n_n3005) & (!x15543x)) + ((x15549x) & (!n_n2934) & (n_n3004) & (!n_n3005) & (x15543x)) + ((x15549x) & (!n_n2934) & (n_n3004) & (n_n3005) & (!x15543x)) + ((x15549x) & (!n_n2934) & (n_n3004) & (n_n3005) & (x15543x)) + ((x15549x) & (n_n2934) & (!n_n3004) & (!n_n3005) & (!x15543x)) + ((x15549x) & (n_n2934) & (!n_n3004) & (!n_n3005) & (x15543x)) + ((x15549x) & (n_n2934) & (!n_n3004) & (n_n3005) & (!x15543x)) + ((x15549x) & (n_n2934) & (!n_n3004) & (n_n3005) & (x15543x)) + ((x15549x) & (n_n2934) & (n_n3004) & (!n_n3005) & (!x15543x)) + ((x15549x) & (n_n2934) & (n_n3004) & (!n_n3005) & (x15543x)) + ((x15549x) & (n_n2934) & (n_n3004) & (n_n3005) & (!x15543x)) + ((x15549x) & (n_n2934) & (n_n3004) & (n_n3005) & (x15543x)));
	assign n_n2902 = (((!n_n2915) & (!n_n2952) & (!x15633x) & (!x15642x) & (x15632x)) + ((!n_n2915) & (!n_n2952) & (!x15633x) & (x15642x) & (!x15632x)) + ((!n_n2915) & (!n_n2952) & (!x15633x) & (x15642x) & (x15632x)) + ((!n_n2915) & (!n_n2952) & (x15633x) & (!x15642x) & (!x15632x)) + ((!n_n2915) & (!n_n2952) & (x15633x) & (!x15642x) & (x15632x)) + ((!n_n2915) & (!n_n2952) & (x15633x) & (x15642x) & (!x15632x)) + ((!n_n2915) & (!n_n2952) & (x15633x) & (x15642x) & (x15632x)) + ((!n_n2915) & (n_n2952) & (!x15633x) & (!x15642x) & (!x15632x)) + ((!n_n2915) & (n_n2952) & (!x15633x) & (!x15642x) & (x15632x)) + ((!n_n2915) & (n_n2952) & (!x15633x) & (x15642x) & (!x15632x)) + ((!n_n2915) & (n_n2952) & (!x15633x) & (x15642x) & (x15632x)) + ((!n_n2915) & (n_n2952) & (x15633x) & (!x15642x) & (!x15632x)) + ((!n_n2915) & (n_n2952) & (x15633x) & (!x15642x) & (x15632x)) + ((!n_n2915) & (n_n2952) & (x15633x) & (x15642x) & (!x15632x)) + ((!n_n2915) & (n_n2952) & (x15633x) & (x15642x) & (x15632x)) + ((n_n2915) & (!n_n2952) & (!x15633x) & (!x15642x) & (!x15632x)) + ((n_n2915) & (!n_n2952) & (!x15633x) & (!x15642x) & (x15632x)) + ((n_n2915) & (!n_n2952) & (!x15633x) & (x15642x) & (!x15632x)) + ((n_n2915) & (!n_n2952) & (!x15633x) & (x15642x) & (x15632x)) + ((n_n2915) & (!n_n2952) & (x15633x) & (!x15642x) & (!x15632x)) + ((n_n2915) & (!n_n2952) & (x15633x) & (!x15642x) & (x15632x)) + ((n_n2915) & (!n_n2952) & (x15633x) & (x15642x) & (!x15632x)) + ((n_n2915) & (!n_n2952) & (x15633x) & (x15642x) & (x15632x)) + ((n_n2915) & (n_n2952) & (!x15633x) & (!x15642x) & (!x15632x)) + ((n_n2915) & (n_n2952) & (!x15633x) & (!x15642x) & (x15632x)) + ((n_n2915) & (n_n2952) & (!x15633x) & (x15642x) & (!x15632x)) + ((n_n2915) & (n_n2952) & (!x15633x) & (x15642x) & (x15632x)) + ((n_n2915) & (n_n2952) & (x15633x) & (!x15642x) & (!x15632x)) + ((n_n2915) & (n_n2952) & (x15633x) & (!x15642x) & (x15632x)) + ((n_n2915) & (n_n2952) & (x15633x) & (x15642x) & (!x15632x)) + ((n_n2915) & (n_n2952) & (x15633x) & (x15642x) & (x15632x)));
	assign x15677x = (((!n_n2912) & (!n_n2911) & (!x15594x) & (!x15674x) & (x15675x)) + ((!n_n2912) & (!n_n2911) & (!x15594x) & (x15674x) & (!x15675x)) + ((!n_n2912) & (!n_n2911) & (!x15594x) & (x15674x) & (x15675x)) + ((!n_n2912) & (!n_n2911) & (x15594x) & (!x15674x) & (!x15675x)) + ((!n_n2912) & (!n_n2911) & (x15594x) & (!x15674x) & (x15675x)) + ((!n_n2912) & (!n_n2911) & (x15594x) & (x15674x) & (!x15675x)) + ((!n_n2912) & (!n_n2911) & (x15594x) & (x15674x) & (x15675x)) + ((!n_n2912) & (n_n2911) & (!x15594x) & (!x15674x) & (!x15675x)) + ((!n_n2912) & (n_n2911) & (!x15594x) & (!x15674x) & (x15675x)) + ((!n_n2912) & (n_n2911) & (!x15594x) & (x15674x) & (!x15675x)) + ((!n_n2912) & (n_n2911) & (!x15594x) & (x15674x) & (x15675x)) + ((!n_n2912) & (n_n2911) & (x15594x) & (!x15674x) & (!x15675x)) + ((!n_n2912) & (n_n2911) & (x15594x) & (!x15674x) & (x15675x)) + ((!n_n2912) & (n_n2911) & (x15594x) & (x15674x) & (!x15675x)) + ((!n_n2912) & (n_n2911) & (x15594x) & (x15674x) & (x15675x)) + ((n_n2912) & (!n_n2911) & (!x15594x) & (!x15674x) & (!x15675x)) + ((n_n2912) & (!n_n2911) & (!x15594x) & (!x15674x) & (x15675x)) + ((n_n2912) & (!n_n2911) & (!x15594x) & (x15674x) & (!x15675x)) + ((n_n2912) & (!n_n2911) & (!x15594x) & (x15674x) & (x15675x)) + ((n_n2912) & (!n_n2911) & (x15594x) & (!x15674x) & (!x15675x)) + ((n_n2912) & (!n_n2911) & (x15594x) & (!x15674x) & (x15675x)) + ((n_n2912) & (!n_n2911) & (x15594x) & (x15674x) & (!x15675x)) + ((n_n2912) & (!n_n2911) & (x15594x) & (x15674x) & (x15675x)) + ((n_n2912) & (n_n2911) & (!x15594x) & (!x15674x) & (!x15675x)) + ((n_n2912) & (n_n2911) & (!x15594x) & (!x15674x) & (x15675x)) + ((n_n2912) & (n_n2911) & (!x15594x) & (x15674x) & (!x15675x)) + ((n_n2912) & (n_n2911) & (!x15594x) & (x15674x) & (x15675x)) + ((n_n2912) & (n_n2911) & (x15594x) & (!x15674x) & (!x15675x)) + ((n_n2912) & (n_n2911) & (x15594x) & (!x15674x) & (x15675x)) + ((n_n2912) & (n_n2911) & (x15594x) & (x15674x) & (!x15675x)) + ((n_n2912) & (n_n2911) & (x15594x) & (x15674x) & (x15675x)));
	assign n_n1793 = (((!x16027x) & (!n_n1882) & (!n_n1817) & (!x16018x) & (x16017x)) + ((!x16027x) & (!n_n1882) & (!n_n1817) & (x16018x) & (!x16017x)) + ((!x16027x) & (!n_n1882) & (!n_n1817) & (x16018x) & (x16017x)) + ((!x16027x) & (!n_n1882) & (n_n1817) & (!x16018x) & (!x16017x)) + ((!x16027x) & (!n_n1882) & (n_n1817) & (!x16018x) & (x16017x)) + ((!x16027x) & (!n_n1882) & (n_n1817) & (x16018x) & (!x16017x)) + ((!x16027x) & (!n_n1882) & (n_n1817) & (x16018x) & (x16017x)) + ((!x16027x) & (n_n1882) & (!n_n1817) & (!x16018x) & (!x16017x)) + ((!x16027x) & (n_n1882) & (!n_n1817) & (!x16018x) & (x16017x)) + ((!x16027x) & (n_n1882) & (!n_n1817) & (x16018x) & (!x16017x)) + ((!x16027x) & (n_n1882) & (!n_n1817) & (x16018x) & (x16017x)) + ((!x16027x) & (n_n1882) & (n_n1817) & (!x16018x) & (!x16017x)) + ((!x16027x) & (n_n1882) & (n_n1817) & (!x16018x) & (x16017x)) + ((!x16027x) & (n_n1882) & (n_n1817) & (x16018x) & (!x16017x)) + ((!x16027x) & (n_n1882) & (n_n1817) & (x16018x) & (x16017x)) + ((x16027x) & (!n_n1882) & (!n_n1817) & (!x16018x) & (!x16017x)) + ((x16027x) & (!n_n1882) & (!n_n1817) & (!x16018x) & (x16017x)) + ((x16027x) & (!n_n1882) & (!n_n1817) & (x16018x) & (!x16017x)) + ((x16027x) & (!n_n1882) & (!n_n1817) & (x16018x) & (x16017x)) + ((x16027x) & (!n_n1882) & (n_n1817) & (!x16018x) & (!x16017x)) + ((x16027x) & (!n_n1882) & (n_n1817) & (!x16018x) & (x16017x)) + ((x16027x) & (!n_n1882) & (n_n1817) & (x16018x) & (!x16017x)) + ((x16027x) & (!n_n1882) & (n_n1817) & (x16018x) & (x16017x)) + ((x16027x) & (n_n1882) & (!n_n1817) & (!x16018x) & (!x16017x)) + ((x16027x) & (n_n1882) & (!n_n1817) & (!x16018x) & (x16017x)) + ((x16027x) & (n_n1882) & (!n_n1817) & (x16018x) & (!x16017x)) + ((x16027x) & (n_n1882) & (!n_n1817) & (x16018x) & (x16017x)) + ((x16027x) & (n_n1882) & (n_n1817) & (!x16018x) & (!x16017x)) + ((x16027x) & (n_n1882) & (n_n1817) & (!x16018x) & (x16017x)) + ((x16027x) & (n_n1882) & (n_n1817) & (x16018x) & (!x16017x)) + ((x16027x) & (n_n1882) & (n_n1817) & (x16018x) & (x16017x)));
	assign n_n1792 = (((!x16072x) & (!n_n1877) & (!x16048x) & (!n_n1812) & (n_n1876)) + ((!x16072x) & (!n_n1877) & (!x16048x) & (n_n1812) & (!n_n1876)) + ((!x16072x) & (!n_n1877) & (!x16048x) & (n_n1812) & (n_n1876)) + ((!x16072x) & (!n_n1877) & (x16048x) & (!n_n1812) & (!n_n1876)) + ((!x16072x) & (!n_n1877) & (x16048x) & (!n_n1812) & (n_n1876)) + ((!x16072x) & (!n_n1877) & (x16048x) & (n_n1812) & (!n_n1876)) + ((!x16072x) & (!n_n1877) & (x16048x) & (n_n1812) & (n_n1876)) + ((!x16072x) & (n_n1877) & (!x16048x) & (!n_n1812) & (!n_n1876)) + ((!x16072x) & (n_n1877) & (!x16048x) & (!n_n1812) & (n_n1876)) + ((!x16072x) & (n_n1877) & (!x16048x) & (n_n1812) & (!n_n1876)) + ((!x16072x) & (n_n1877) & (!x16048x) & (n_n1812) & (n_n1876)) + ((!x16072x) & (n_n1877) & (x16048x) & (!n_n1812) & (!n_n1876)) + ((!x16072x) & (n_n1877) & (x16048x) & (!n_n1812) & (n_n1876)) + ((!x16072x) & (n_n1877) & (x16048x) & (n_n1812) & (!n_n1876)) + ((!x16072x) & (n_n1877) & (x16048x) & (n_n1812) & (n_n1876)) + ((x16072x) & (!n_n1877) & (!x16048x) & (!n_n1812) & (!n_n1876)) + ((x16072x) & (!n_n1877) & (!x16048x) & (!n_n1812) & (n_n1876)) + ((x16072x) & (!n_n1877) & (!x16048x) & (n_n1812) & (!n_n1876)) + ((x16072x) & (!n_n1877) & (!x16048x) & (n_n1812) & (n_n1876)) + ((x16072x) & (!n_n1877) & (x16048x) & (!n_n1812) & (!n_n1876)) + ((x16072x) & (!n_n1877) & (x16048x) & (!n_n1812) & (n_n1876)) + ((x16072x) & (!n_n1877) & (x16048x) & (n_n1812) & (!n_n1876)) + ((x16072x) & (!n_n1877) & (x16048x) & (n_n1812) & (n_n1876)) + ((x16072x) & (n_n1877) & (!x16048x) & (!n_n1812) & (!n_n1876)) + ((x16072x) & (n_n1877) & (!x16048x) & (!n_n1812) & (n_n1876)) + ((x16072x) & (n_n1877) & (!x16048x) & (n_n1812) & (!n_n1876)) + ((x16072x) & (n_n1877) & (!x16048x) & (n_n1812) & (n_n1876)) + ((x16072x) & (n_n1877) & (x16048x) & (!n_n1812) & (!n_n1876)) + ((x16072x) & (n_n1877) & (x16048x) & (!n_n1812) & (n_n1876)) + ((x16072x) & (n_n1877) & (x16048x) & (n_n1812) & (!n_n1876)) + ((x16072x) & (n_n1877) & (x16048x) & (n_n1812) & (n_n1876)));
	assign n_n1794 = (((!x16114x) & (!n_n1896) & (!x16086x) & (!n_n1818) & (x16085x)) + ((!x16114x) & (!n_n1896) & (!x16086x) & (n_n1818) & (!x16085x)) + ((!x16114x) & (!n_n1896) & (!x16086x) & (n_n1818) & (x16085x)) + ((!x16114x) & (!n_n1896) & (x16086x) & (!n_n1818) & (!x16085x)) + ((!x16114x) & (!n_n1896) & (x16086x) & (!n_n1818) & (x16085x)) + ((!x16114x) & (!n_n1896) & (x16086x) & (n_n1818) & (!x16085x)) + ((!x16114x) & (!n_n1896) & (x16086x) & (n_n1818) & (x16085x)) + ((!x16114x) & (n_n1896) & (!x16086x) & (!n_n1818) & (!x16085x)) + ((!x16114x) & (n_n1896) & (!x16086x) & (!n_n1818) & (x16085x)) + ((!x16114x) & (n_n1896) & (!x16086x) & (n_n1818) & (!x16085x)) + ((!x16114x) & (n_n1896) & (!x16086x) & (n_n1818) & (x16085x)) + ((!x16114x) & (n_n1896) & (x16086x) & (!n_n1818) & (!x16085x)) + ((!x16114x) & (n_n1896) & (x16086x) & (!n_n1818) & (x16085x)) + ((!x16114x) & (n_n1896) & (x16086x) & (n_n1818) & (!x16085x)) + ((!x16114x) & (n_n1896) & (x16086x) & (n_n1818) & (x16085x)) + ((x16114x) & (!n_n1896) & (!x16086x) & (!n_n1818) & (!x16085x)) + ((x16114x) & (!n_n1896) & (!x16086x) & (!n_n1818) & (x16085x)) + ((x16114x) & (!n_n1896) & (!x16086x) & (n_n1818) & (!x16085x)) + ((x16114x) & (!n_n1896) & (!x16086x) & (n_n1818) & (x16085x)) + ((x16114x) & (!n_n1896) & (x16086x) & (!n_n1818) & (!x16085x)) + ((x16114x) & (!n_n1896) & (x16086x) & (!n_n1818) & (x16085x)) + ((x16114x) & (!n_n1896) & (x16086x) & (n_n1818) & (!x16085x)) + ((x16114x) & (!n_n1896) & (x16086x) & (n_n1818) & (x16085x)) + ((x16114x) & (n_n1896) & (!x16086x) & (!n_n1818) & (!x16085x)) + ((x16114x) & (n_n1896) & (!x16086x) & (!n_n1818) & (x16085x)) + ((x16114x) & (n_n1896) & (!x16086x) & (n_n1818) & (!x16085x)) + ((x16114x) & (n_n1896) & (!x16086x) & (n_n1818) & (x16085x)) + ((x16114x) & (n_n1896) & (x16086x) & (!n_n1818) & (!x16085x)) + ((x16114x) & (n_n1896) & (x16086x) & (!n_n1818) & (x16085x)) + ((x16114x) & (n_n1896) & (x16086x) & (n_n1818) & (!x16085x)) + ((x16114x) & (n_n1896) & (x16086x) & (n_n1818) & (x16085x)));
	assign n_n1787 = (((!x16289x) & (!n_n1832) & (!x16262x) & (!n_n1797) & (x16261x)) + ((!x16289x) & (!n_n1832) & (!x16262x) & (n_n1797) & (!x16261x)) + ((!x16289x) & (!n_n1832) & (!x16262x) & (n_n1797) & (x16261x)) + ((!x16289x) & (!n_n1832) & (x16262x) & (!n_n1797) & (!x16261x)) + ((!x16289x) & (!n_n1832) & (x16262x) & (!n_n1797) & (x16261x)) + ((!x16289x) & (!n_n1832) & (x16262x) & (n_n1797) & (!x16261x)) + ((!x16289x) & (!n_n1832) & (x16262x) & (n_n1797) & (x16261x)) + ((!x16289x) & (n_n1832) & (!x16262x) & (!n_n1797) & (!x16261x)) + ((!x16289x) & (n_n1832) & (!x16262x) & (!n_n1797) & (x16261x)) + ((!x16289x) & (n_n1832) & (!x16262x) & (n_n1797) & (!x16261x)) + ((!x16289x) & (n_n1832) & (!x16262x) & (n_n1797) & (x16261x)) + ((!x16289x) & (n_n1832) & (x16262x) & (!n_n1797) & (!x16261x)) + ((!x16289x) & (n_n1832) & (x16262x) & (!n_n1797) & (x16261x)) + ((!x16289x) & (n_n1832) & (x16262x) & (n_n1797) & (!x16261x)) + ((!x16289x) & (n_n1832) & (x16262x) & (n_n1797) & (x16261x)) + ((x16289x) & (!n_n1832) & (!x16262x) & (!n_n1797) & (!x16261x)) + ((x16289x) & (!n_n1832) & (!x16262x) & (!n_n1797) & (x16261x)) + ((x16289x) & (!n_n1832) & (!x16262x) & (n_n1797) & (!x16261x)) + ((x16289x) & (!n_n1832) & (!x16262x) & (n_n1797) & (x16261x)) + ((x16289x) & (!n_n1832) & (x16262x) & (!n_n1797) & (!x16261x)) + ((x16289x) & (!n_n1832) & (x16262x) & (!n_n1797) & (x16261x)) + ((x16289x) & (!n_n1832) & (x16262x) & (n_n1797) & (!x16261x)) + ((x16289x) & (!n_n1832) & (x16262x) & (n_n1797) & (x16261x)) + ((x16289x) & (n_n1832) & (!x16262x) & (!n_n1797) & (!x16261x)) + ((x16289x) & (n_n1832) & (!x16262x) & (!n_n1797) & (x16261x)) + ((x16289x) & (n_n1832) & (!x16262x) & (n_n1797) & (!x16261x)) + ((x16289x) & (n_n1832) & (!x16262x) & (n_n1797) & (x16261x)) + ((x16289x) & (n_n1832) & (x16262x) & (!n_n1797) & (!x16261x)) + ((x16289x) & (n_n1832) & (x16262x) & (!n_n1797) & (x16261x)) + ((x16289x) & (n_n1832) & (x16262x) & (n_n1797) & (!x16261x)) + ((x16289x) & (n_n1832) & (x16262x) & (n_n1797) & (x16261x)));
	assign x16470x = (((!n_n2175) & (!x16456x) & (!n_n2223) & (!n_n2225) & (x16468x)) + ((!n_n2175) & (!x16456x) & (!n_n2223) & (n_n2225) & (!x16468x)) + ((!n_n2175) & (!x16456x) & (!n_n2223) & (n_n2225) & (x16468x)) + ((!n_n2175) & (!x16456x) & (n_n2223) & (!n_n2225) & (!x16468x)) + ((!n_n2175) & (!x16456x) & (n_n2223) & (!n_n2225) & (x16468x)) + ((!n_n2175) & (!x16456x) & (n_n2223) & (n_n2225) & (!x16468x)) + ((!n_n2175) & (!x16456x) & (n_n2223) & (n_n2225) & (x16468x)) + ((!n_n2175) & (x16456x) & (!n_n2223) & (!n_n2225) & (!x16468x)) + ((!n_n2175) & (x16456x) & (!n_n2223) & (!n_n2225) & (x16468x)) + ((!n_n2175) & (x16456x) & (!n_n2223) & (n_n2225) & (!x16468x)) + ((!n_n2175) & (x16456x) & (!n_n2223) & (n_n2225) & (x16468x)) + ((!n_n2175) & (x16456x) & (n_n2223) & (!n_n2225) & (!x16468x)) + ((!n_n2175) & (x16456x) & (n_n2223) & (!n_n2225) & (x16468x)) + ((!n_n2175) & (x16456x) & (n_n2223) & (n_n2225) & (!x16468x)) + ((!n_n2175) & (x16456x) & (n_n2223) & (n_n2225) & (x16468x)) + ((n_n2175) & (!x16456x) & (!n_n2223) & (!n_n2225) & (!x16468x)) + ((n_n2175) & (!x16456x) & (!n_n2223) & (!n_n2225) & (x16468x)) + ((n_n2175) & (!x16456x) & (!n_n2223) & (n_n2225) & (!x16468x)) + ((n_n2175) & (!x16456x) & (!n_n2223) & (n_n2225) & (x16468x)) + ((n_n2175) & (!x16456x) & (n_n2223) & (!n_n2225) & (!x16468x)) + ((n_n2175) & (!x16456x) & (n_n2223) & (!n_n2225) & (x16468x)) + ((n_n2175) & (!x16456x) & (n_n2223) & (n_n2225) & (!x16468x)) + ((n_n2175) & (!x16456x) & (n_n2223) & (n_n2225) & (x16468x)) + ((n_n2175) & (x16456x) & (!n_n2223) & (!n_n2225) & (!x16468x)) + ((n_n2175) & (x16456x) & (!n_n2223) & (!n_n2225) & (x16468x)) + ((n_n2175) & (x16456x) & (!n_n2223) & (n_n2225) & (!x16468x)) + ((n_n2175) & (x16456x) & (!n_n2223) & (n_n2225) & (x16468x)) + ((n_n2175) & (x16456x) & (n_n2223) & (!n_n2225) & (!x16468x)) + ((n_n2175) & (x16456x) & (n_n2223) & (!n_n2225) & (x16468x)) + ((n_n2175) & (x16456x) & (n_n2223) & (n_n2225) & (!x16468x)) + ((n_n2175) & (x16456x) & (n_n2223) & (n_n2225) & (x16468x)));
	assign n_n2165 = (((!x16598x) & (!n_n2189) & (!x16590x) & (!n_n2253) & (x16589x)) + ((!x16598x) & (!n_n2189) & (!x16590x) & (n_n2253) & (!x16589x)) + ((!x16598x) & (!n_n2189) & (!x16590x) & (n_n2253) & (x16589x)) + ((!x16598x) & (!n_n2189) & (x16590x) & (!n_n2253) & (!x16589x)) + ((!x16598x) & (!n_n2189) & (x16590x) & (!n_n2253) & (x16589x)) + ((!x16598x) & (!n_n2189) & (x16590x) & (n_n2253) & (!x16589x)) + ((!x16598x) & (!n_n2189) & (x16590x) & (n_n2253) & (x16589x)) + ((!x16598x) & (n_n2189) & (!x16590x) & (!n_n2253) & (!x16589x)) + ((!x16598x) & (n_n2189) & (!x16590x) & (!n_n2253) & (x16589x)) + ((!x16598x) & (n_n2189) & (!x16590x) & (n_n2253) & (!x16589x)) + ((!x16598x) & (n_n2189) & (!x16590x) & (n_n2253) & (x16589x)) + ((!x16598x) & (n_n2189) & (x16590x) & (!n_n2253) & (!x16589x)) + ((!x16598x) & (n_n2189) & (x16590x) & (!n_n2253) & (x16589x)) + ((!x16598x) & (n_n2189) & (x16590x) & (n_n2253) & (!x16589x)) + ((!x16598x) & (n_n2189) & (x16590x) & (n_n2253) & (x16589x)) + ((x16598x) & (!n_n2189) & (!x16590x) & (!n_n2253) & (!x16589x)) + ((x16598x) & (!n_n2189) & (!x16590x) & (!n_n2253) & (x16589x)) + ((x16598x) & (!n_n2189) & (!x16590x) & (n_n2253) & (!x16589x)) + ((x16598x) & (!n_n2189) & (!x16590x) & (n_n2253) & (x16589x)) + ((x16598x) & (!n_n2189) & (x16590x) & (!n_n2253) & (!x16589x)) + ((x16598x) & (!n_n2189) & (x16590x) & (!n_n2253) & (x16589x)) + ((x16598x) & (!n_n2189) & (x16590x) & (n_n2253) & (!x16589x)) + ((x16598x) & (!n_n2189) & (x16590x) & (n_n2253) & (x16589x)) + ((x16598x) & (n_n2189) & (!x16590x) & (!n_n2253) & (!x16589x)) + ((x16598x) & (n_n2189) & (!x16590x) & (!n_n2253) & (x16589x)) + ((x16598x) & (n_n2189) & (!x16590x) & (n_n2253) & (!x16589x)) + ((x16598x) & (n_n2189) & (!x16590x) & (n_n2253) & (x16589x)) + ((x16598x) & (n_n2189) & (x16590x) & (!n_n2253) & (!x16589x)) + ((x16598x) & (n_n2189) & (x16590x) & (!n_n2253) & (x16589x)) + ((x16598x) & (n_n2189) & (x16590x) & (n_n2253) & (!x16589x)) + ((x16598x) & (n_n2189) & (x16590x) & (n_n2253) & (x16589x)));
	assign n_n2164 = (((!x16645x) & (!n_n2185) & (n_n2184)) + ((!x16645x) & (n_n2185) & (!n_n2184)) + ((!x16645x) & (n_n2185) & (n_n2184)) + ((x16645x) & (!n_n2185) & (!n_n2184)) + ((x16645x) & (!n_n2185) & (n_n2184)) + ((x16645x) & (n_n2185) & (!n_n2184)) + ((x16645x) & (n_n2185) & (n_n2184)));
	assign n_n2162 = (((!n_n2178) & (!x16365x) & (!x16376x) & (!x16362x) & (x16363x)) + ((!n_n2178) & (!x16365x) & (!x16376x) & (x16362x) & (!x16363x)) + ((!n_n2178) & (!x16365x) & (!x16376x) & (x16362x) & (x16363x)) + ((!n_n2178) & (!x16365x) & (x16376x) & (!x16362x) & (!x16363x)) + ((!n_n2178) & (!x16365x) & (x16376x) & (!x16362x) & (x16363x)) + ((!n_n2178) & (!x16365x) & (x16376x) & (x16362x) & (!x16363x)) + ((!n_n2178) & (!x16365x) & (x16376x) & (x16362x) & (x16363x)) + ((!n_n2178) & (x16365x) & (!x16376x) & (!x16362x) & (!x16363x)) + ((!n_n2178) & (x16365x) & (!x16376x) & (!x16362x) & (x16363x)) + ((!n_n2178) & (x16365x) & (!x16376x) & (x16362x) & (!x16363x)) + ((!n_n2178) & (x16365x) & (!x16376x) & (x16362x) & (x16363x)) + ((!n_n2178) & (x16365x) & (x16376x) & (!x16362x) & (!x16363x)) + ((!n_n2178) & (x16365x) & (x16376x) & (!x16362x) & (x16363x)) + ((!n_n2178) & (x16365x) & (x16376x) & (x16362x) & (!x16363x)) + ((!n_n2178) & (x16365x) & (x16376x) & (x16362x) & (x16363x)) + ((n_n2178) & (!x16365x) & (!x16376x) & (!x16362x) & (!x16363x)) + ((n_n2178) & (!x16365x) & (!x16376x) & (!x16362x) & (x16363x)) + ((n_n2178) & (!x16365x) & (!x16376x) & (x16362x) & (!x16363x)) + ((n_n2178) & (!x16365x) & (!x16376x) & (x16362x) & (x16363x)) + ((n_n2178) & (!x16365x) & (x16376x) & (!x16362x) & (!x16363x)) + ((n_n2178) & (!x16365x) & (x16376x) & (!x16362x) & (x16363x)) + ((n_n2178) & (!x16365x) & (x16376x) & (x16362x) & (!x16363x)) + ((n_n2178) & (!x16365x) & (x16376x) & (x16362x) & (x16363x)) + ((n_n2178) & (x16365x) & (!x16376x) & (!x16362x) & (!x16363x)) + ((n_n2178) & (x16365x) & (!x16376x) & (!x16362x) & (x16363x)) + ((n_n2178) & (x16365x) & (!x16376x) & (x16362x) & (!x16363x)) + ((n_n2178) & (x16365x) & (!x16376x) & (x16362x) & (x16363x)) + ((n_n2178) & (x16365x) & (x16376x) & (!x16362x) & (!x16363x)) + ((n_n2178) & (x16365x) & (x16376x) & (!x16362x) & (x16363x)) + ((n_n2178) & (x16365x) & (x16376x) & (x16362x) & (!x16363x)) + ((n_n2178) & (x16365x) & (x16376x) & (x16362x) & (x16363x)));
	assign n_n2163 = (((!n_n2236) & (!n_n2237) & (!n_n2182) & (!n_n2183) & (x16423x)) + ((!n_n2236) & (!n_n2237) & (!n_n2182) & (n_n2183) & (!x16423x)) + ((!n_n2236) & (!n_n2237) & (!n_n2182) & (n_n2183) & (x16423x)) + ((!n_n2236) & (!n_n2237) & (n_n2182) & (!n_n2183) & (!x16423x)) + ((!n_n2236) & (!n_n2237) & (n_n2182) & (!n_n2183) & (x16423x)) + ((!n_n2236) & (!n_n2237) & (n_n2182) & (n_n2183) & (!x16423x)) + ((!n_n2236) & (!n_n2237) & (n_n2182) & (n_n2183) & (x16423x)) + ((!n_n2236) & (n_n2237) & (!n_n2182) & (!n_n2183) & (!x16423x)) + ((!n_n2236) & (n_n2237) & (!n_n2182) & (!n_n2183) & (x16423x)) + ((!n_n2236) & (n_n2237) & (!n_n2182) & (n_n2183) & (!x16423x)) + ((!n_n2236) & (n_n2237) & (!n_n2182) & (n_n2183) & (x16423x)) + ((!n_n2236) & (n_n2237) & (n_n2182) & (!n_n2183) & (!x16423x)) + ((!n_n2236) & (n_n2237) & (n_n2182) & (!n_n2183) & (x16423x)) + ((!n_n2236) & (n_n2237) & (n_n2182) & (n_n2183) & (!x16423x)) + ((!n_n2236) & (n_n2237) & (n_n2182) & (n_n2183) & (x16423x)) + ((n_n2236) & (!n_n2237) & (!n_n2182) & (!n_n2183) & (!x16423x)) + ((n_n2236) & (!n_n2237) & (!n_n2182) & (!n_n2183) & (x16423x)) + ((n_n2236) & (!n_n2237) & (!n_n2182) & (n_n2183) & (!x16423x)) + ((n_n2236) & (!n_n2237) & (!n_n2182) & (n_n2183) & (x16423x)) + ((n_n2236) & (!n_n2237) & (n_n2182) & (!n_n2183) & (!x16423x)) + ((n_n2236) & (!n_n2237) & (n_n2182) & (!n_n2183) & (x16423x)) + ((n_n2236) & (!n_n2237) & (n_n2182) & (n_n2183) & (!x16423x)) + ((n_n2236) & (!n_n2237) & (n_n2182) & (n_n2183) & (x16423x)) + ((n_n2236) & (n_n2237) & (!n_n2182) & (!n_n2183) & (!x16423x)) + ((n_n2236) & (n_n2237) & (!n_n2182) & (!n_n2183) & (x16423x)) + ((n_n2236) & (n_n2237) & (!n_n2182) & (n_n2183) & (!x16423x)) + ((n_n2236) & (n_n2237) & (!n_n2182) & (n_n2183) & (x16423x)) + ((n_n2236) & (n_n2237) & (n_n2182) & (!n_n2183) & (!x16423x)) + ((n_n2236) & (n_n2237) & (n_n2182) & (!n_n2183) & (x16423x)) + ((n_n2236) & (n_n2237) & (n_n2182) & (n_n2183) & (!x16423x)) + ((n_n2236) & (n_n2237) & (n_n2182) & (n_n2183) & (x16423x)));
	assign n_n2166 = (((!x16557x) & (!n_n2190) & (!n_n2268) & (!x16545x) & (x16544x)) + ((!x16557x) & (!n_n2190) & (!n_n2268) & (x16545x) & (!x16544x)) + ((!x16557x) & (!n_n2190) & (!n_n2268) & (x16545x) & (x16544x)) + ((!x16557x) & (!n_n2190) & (n_n2268) & (!x16545x) & (!x16544x)) + ((!x16557x) & (!n_n2190) & (n_n2268) & (!x16545x) & (x16544x)) + ((!x16557x) & (!n_n2190) & (n_n2268) & (x16545x) & (!x16544x)) + ((!x16557x) & (!n_n2190) & (n_n2268) & (x16545x) & (x16544x)) + ((!x16557x) & (n_n2190) & (!n_n2268) & (!x16545x) & (!x16544x)) + ((!x16557x) & (n_n2190) & (!n_n2268) & (!x16545x) & (x16544x)) + ((!x16557x) & (n_n2190) & (!n_n2268) & (x16545x) & (!x16544x)) + ((!x16557x) & (n_n2190) & (!n_n2268) & (x16545x) & (x16544x)) + ((!x16557x) & (n_n2190) & (n_n2268) & (!x16545x) & (!x16544x)) + ((!x16557x) & (n_n2190) & (n_n2268) & (!x16545x) & (x16544x)) + ((!x16557x) & (n_n2190) & (n_n2268) & (x16545x) & (!x16544x)) + ((!x16557x) & (n_n2190) & (n_n2268) & (x16545x) & (x16544x)) + ((x16557x) & (!n_n2190) & (!n_n2268) & (!x16545x) & (!x16544x)) + ((x16557x) & (!n_n2190) & (!n_n2268) & (!x16545x) & (x16544x)) + ((x16557x) & (!n_n2190) & (!n_n2268) & (x16545x) & (!x16544x)) + ((x16557x) & (!n_n2190) & (!n_n2268) & (x16545x) & (x16544x)) + ((x16557x) & (!n_n2190) & (n_n2268) & (!x16545x) & (!x16544x)) + ((x16557x) & (!n_n2190) & (n_n2268) & (!x16545x) & (x16544x)) + ((x16557x) & (!n_n2190) & (n_n2268) & (x16545x) & (!x16544x)) + ((x16557x) & (!n_n2190) & (n_n2268) & (x16545x) & (x16544x)) + ((x16557x) & (n_n2190) & (!n_n2268) & (!x16545x) & (!x16544x)) + ((x16557x) & (n_n2190) & (!n_n2268) & (!x16545x) & (x16544x)) + ((x16557x) & (n_n2190) & (!n_n2268) & (x16545x) & (!x16544x)) + ((x16557x) & (n_n2190) & (!n_n2268) & (x16545x) & (x16544x)) + ((x16557x) & (n_n2190) & (n_n2268) & (!x16545x) & (!x16544x)) + ((x16557x) & (n_n2190) & (n_n2268) & (!x16545x) & (x16544x)) + ((x16557x) & (n_n2190) & (n_n2268) & (x16545x) & (!x16544x)) + ((x16557x) & (n_n2190) & (n_n2268) & (x16545x) & (x16544x)));
	assign n_n2160 = (((!x467x) & (!n_n2173) & (!n_n2172) & (!n_n2214) & (x16742x)) + ((!x467x) & (!n_n2173) & (!n_n2172) & (n_n2214) & (!x16742x)) + ((!x467x) & (!n_n2173) & (!n_n2172) & (n_n2214) & (x16742x)) + ((!x467x) & (!n_n2173) & (n_n2172) & (!n_n2214) & (!x16742x)) + ((!x467x) & (!n_n2173) & (n_n2172) & (!n_n2214) & (x16742x)) + ((!x467x) & (!n_n2173) & (n_n2172) & (n_n2214) & (!x16742x)) + ((!x467x) & (!n_n2173) & (n_n2172) & (n_n2214) & (x16742x)) + ((!x467x) & (n_n2173) & (!n_n2172) & (!n_n2214) & (!x16742x)) + ((!x467x) & (n_n2173) & (!n_n2172) & (!n_n2214) & (x16742x)) + ((!x467x) & (n_n2173) & (!n_n2172) & (n_n2214) & (!x16742x)) + ((!x467x) & (n_n2173) & (!n_n2172) & (n_n2214) & (x16742x)) + ((!x467x) & (n_n2173) & (n_n2172) & (!n_n2214) & (!x16742x)) + ((!x467x) & (n_n2173) & (n_n2172) & (!n_n2214) & (x16742x)) + ((!x467x) & (n_n2173) & (n_n2172) & (n_n2214) & (!x16742x)) + ((!x467x) & (n_n2173) & (n_n2172) & (n_n2214) & (x16742x)) + ((x467x) & (!n_n2173) & (!n_n2172) & (!n_n2214) & (!x16742x)) + ((x467x) & (!n_n2173) & (!n_n2172) & (!n_n2214) & (x16742x)) + ((x467x) & (!n_n2173) & (!n_n2172) & (n_n2214) & (!x16742x)) + ((x467x) & (!n_n2173) & (!n_n2172) & (n_n2214) & (x16742x)) + ((x467x) & (!n_n2173) & (n_n2172) & (!n_n2214) & (!x16742x)) + ((x467x) & (!n_n2173) & (n_n2172) & (!n_n2214) & (x16742x)) + ((x467x) & (!n_n2173) & (n_n2172) & (n_n2214) & (!x16742x)) + ((x467x) & (!n_n2173) & (n_n2172) & (n_n2214) & (x16742x)) + ((x467x) & (n_n2173) & (!n_n2172) & (!n_n2214) & (!x16742x)) + ((x467x) & (n_n2173) & (!n_n2172) & (!n_n2214) & (x16742x)) + ((x467x) & (n_n2173) & (!n_n2172) & (n_n2214) & (!x16742x)) + ((x467x) & (n_n2173) & (!n_n2172) & (n_n2214) & (x16742x)) + ((x467x) & (n_n2173) & (n_n2172) & (!n_n2214) & (!x16742x)) + ((x467x) & (n_n2173) & (n_n2172) & (!n_n2214) & (x16742x)) + ((x467x) & (n_n2173) & (n_n2172) & (n_n2214) & (!x16742x)) + ((x467x) & (n_n2173) & (n_n2172) & (n_n2214) & (x16742x)));
	assign x16764x = (((!n_n2170) & (!n_n2169) & (!x16705x) & (!n_n2168) & (x16762x)) + ((!n_n2170) & (!n_n2169) & (!x16705x) & (n_n2168) & (!x16762x)) + ((!n_n2170) & (!n_n2169) & (!x16705x) & (n_n2168) & (x16762x)) + ((!n_n2170) & (!n_n2169) & (x16705x) & (!n_n2168) & (!x16762x)) + ((!n_n2170) & (!n_n2169) & (x16705x) & (!n_n2168) & (x16762x)) + ((!n_n2170) & (!n_n2169) & (x16705x) & (n_n2168) & (!x16762x)) + ((!n_n2170) & (!n_n2169) & (x16705x) & (n_n2168) & (x16762x)) + ((!n_n2170) & (n_n2169) & (!x16705x) & (!n_n2168) & (!x16762x)) + ((!n_n2170) & (n_n2169) & (!x16705x) & (!n_n2168) & (x16762x)) + ((!n_n2170) & (n_n2169) & (!x16705x) & (n_n2168) & (!x16762x)) + ((!n_n2170) & (n_n2169) & (!x16705x) & (n_n2168) & (x16762x)) + ((!n_n2170) & (n_n2169) & (x16705x) & (!n_n2168) & (!x16762x)) + ((!n_n2170) & (n_n2169) & (x16705x) & (!n_n2168) & (x16762x)) + ((!n_n2170) & (n_n2169) & (x16705x) & (n_n2168) & (!x16762x)) + ((!n_n2170) & (n_n2169) & (x16705x) & (n_n2168) & (x16762x)) + ((n_n2170) & (!n_n2169) & (!x16705x) & (!n_n2168) & (!x16762x)) + ((n_n2170) & (!n_n2169) & (!x16705x) & (!n_n2168) & (x16762x)) + ((n_n2170) & (!n_n2169) & (!x16705x) & (n_n2168) & (!x16762x)) + ((n_n2170) & (!n_n2169) & (!x16705x) & (n_n2168) & (x16762x)) + ((n_n2170) & (!n_n2169) & (x16705x) & (!n_n2168) & (!x16762x)) + ((n_n2170) & (!n_n2169) & (x16705x) & (!n_n2168) & (x16762x)) + ((n_n2170) & (!n_n2169) & (x16705x) & (n_n2168) & (!x16762x)) + ((n_n2170) & (!n_n2169) & (x16705x) & (n_n2168) & (x16762x)) + ((n_n2170) & (n_n2169) & (!x16705x) & (!n_n2168) & (!x16762x)) + ((n_n2170) & (n_n2169) & (!x16705x) & (!n_n2168) & (x16762x)) + ((n_n2170) & (n_n2169) & (!x16705x) & (n_n2168) & (!x16762x)) + ((n_n2170) & (n_n2169) & (!x16705x) & (n_n2168) & (x16762x)) + ((n_n2170) & (n_n2169) & (x16705x) & (!n_n2168) & (!x16762x)) + ((n_n2170) & (n_n2169) & (x16705x) & (!n_n2168) & (x16762x)) + ((n_n2170) & (n_n2169) & (x16705x) & (n_n2168) & (!x16762x)) + ((n_n2170) & (n_n2169) & (x16705x) & (n_n2168) & (x16762x)));
	assign x16826x = (((!n_n2087) & (!x16516x) & (x16517x)) + ((!n_n2087) & (x16516x) & (!x16517x)) + ((!n_n2087) & (x16516x) & (x16517x)) + ((n_n2087) & (!x16516x) & (!x16517x)) + ((n_n2087) & (!x16516x) & (x16517x)) + ((n_n2087) & (x16516x) & (!x16517x)) + ((n_n2087) & (x16516x) & (x16517x)));
	assign x16827x = (((!n_n2103) & (!n_n2084) & (!x16821x) & (!x16822x) & (x16824x)) + ((!n_n2103) & (!n_n2084) & (!x16821x) & (x16822x) & (!x16824x)) + ((!n_n2103) & (!n_n2084) & (!x16821x) & (x16822x) & (x16824x)) + ((!n_n2103) & (!n_n2084) & (x16821x) & (!x16822x) & (!x16824x)) + ((!n_n2103) & (!n_n2084) & (x16821x) & (!x16822x) & (x16824x)) + ((!n_n2103) & (!n_n2084) & (x16821x) & (x16822x) & (!x16824x)) + ((!n_n2103) & (!n_n2084) & (x16821x) & (x16822x) & (x16824x)) + ((!n_n2103) & (n_n2084) & (!x16821x) & (!x16822x) & (!x16824x)) + ((!n_n2103) & (n_n2084) & (!x16821x) & (!x16822x) & (x16824x)) + ((!n_n2103) & (n_n2084) & (!x16821x) & (x16822x) & (!x16824x)) + ((!n_n2103) & (n_n2084) & (!x16821x) & (x16822x) & (x16824x)) + ((!n_n2103) & (n_n2084) & (x16821x) & (!x16822x) & (!x16824x)) + ((!n_n2103) & (n_n2084) & (x16821x) & (!x16822x) & (x16824x)) + ((!n_n2103) & (n_n2084) & (x16821x) & (x16822x) & (!x16824x)) + ((!n_n2103) & (n_n2084) & (x16821x) & (x16822x) & (x16824x)) + ((n_n2103) & (!n_n2084) & (!x16821x) & (!x16822x) & (!x16824x)) + ((n_n2103) & (!n_n2084) & (!x16821x) & (!x16822x) & (x16824x)) + ((n_n2103) & (!n_n2084) & (!x16821x) & (x16822x) & (!x16824x)) + ((n_n2103) & (!n_n2084) & (!x16821x) & (x16822x) & (x16824x)) + ((n_n2103) & (!n_n2084) & (x16821x) & (!x16822x) & (!x16824x)) + ((n_n2103) & (!n_n2084) & (x16821x) & (!x16822x) & (x16824x)) + ((n_n2103) & (!n_n2084) & (x16821x) & (x16822x) & (!x16824x)) + ((n_n2103) & (!n_n2084) & (x16821x) & (x16822x) & (x16824x)) + ((n_n2103) & (n_n2084) & (!x16821x) & (!x16822x) & (!x16824x)) + ((n_n2103) & (n_n2084) & (!x16821x) & (!x16822x) & (x16824x)) + ((n_n2103) & (n_n2084) & (!x16821x) & (x16822x) & (!x16824x)) + ((n_n2103) & (n_n2084) & (!x16821x) & (x16822x) & (x16824x)) + ((n_n2103) & (n_n2084) & (x16821x) & (!x16822x) & (!x16824x)) + ((n_n2103) & (n_n2084) & (x16821x) & (!x16822x) & (x16824x)) + ((n_n2103) & (n_n2084) & (x16821x) & (x16822x) & (!x16824x)) + ((n_n2103) & (n_n2084) & (x16821x) & (x16822x) & (x16824x)));
	assign n_n1113 = (((!n_n4440) & (!n_n4434) & (!n_n4442) & (!n_n4443) & (!x22164x)) + ((!n_n4440) & (!n_n4434) & (!n_n4442) & (n_n4443) & (!x22164x)) + ((!n_n4440) & (!n_n4434) & (!n_n4442) & (n_n4443) & (x22164x)) + ((!n_n4440) & (!n_n4434) & (n_n4442) & (!n_n4443) & (!x22164x)) + ((!n_n4440) & (!n_n4434) & (n_n4442) & (!n_n4443) & (x22164x)) + ((!n_n4440) & (!n_n4434) & (n_n4442) & (n_n4443) & (!x22164x)) + ((!n_n4440) & (!n_n4434) & (n_n4442) & (n_n4443) & (x22164x)) + ((!n_n4440) & (n_n4434) & (!n_n4442) & (!n_n4443) & (!x22164x)) + ((!n_n4440) & (n_n4434) & (!n_n4442) & (!n_n4443) & (x22164x)) + ((!n_n4440) & (n_n4434) & (!n_n4442) & (n_n4443) & (!x22164x)) + ((!n_n4440) & (n_n4434) & (!n_n4442) & (n_n4443) & (x22164x)) + ((!n_n4440) & (n_n4434) & (n_n4442) & (!n_n4443) & (!x22164x)) + ((!n_n4440) & (n_n4434) & (n_n4442) & (!n_n4443) & (x22164x)) + ((!n_n4440) & (n_n4434) & (n_n4442) & (n_n4443) & (!x22164x)) + ((!n_n4440) & (n_n4434) & (n_n4442) & (n_n4443) & (x22164x)) + ((n_n4440) & (!n_n4434) & (!n_n4442) & (!n_n4443) & (!x22164x)) + ((n_n4440) & (!n_n4434) & (!n_n4442) & (!n_n4443) & (x22164x)) + ((n_n4440) & (!n_n4434) & (!n_n4442) & (n_n4443) & (!x22164x)) + ((n_n4440) & (!n_n4434) & (!n_n4442) & (n_n4443) & (x22164x)) + ((n_n4440) & (!n_n4434) & (n_n4442) & (!n_n4443) & (!x22164x)) + ((n_n4440) & (!n_n4434) & (n_n4442) & (!n_n4443) & (x22164x)) + ((n_n4440) & (!n_n4434) & (n_n4442) & (n_n4443) & (!x22164x)) + ((n_n4440) & (!n_n4434) & (n_n4442) & (n_n4443) & (x22164x)) + ((n_n4440) & (n_n4434) & (!n_n4442) & (!n_n4443) & (!x22164x)) + ((n_n4440) & (n_n4434) & (!n_n4442) & (!n_n4443) & (x22164x)) + ((n_n4440) & (n_n4434) & (!n_n4442) & (n_n4443) & (!x22164x)) + ((n_n4440) & (n_n4434) & (!n_n4442) & (n_n4443) & (x22164x)) + ((n_n4440) & (n_n4434) & (n_n4442) & (!n_n4443) & (!x22164x)) + ((n_n4440) & (n_n4434) & (n_n4442) & (!n_n4443) & (x22164x)) + ((n_n4440) & (n_n4434) & (n_n4442) & (n_n4443) & (!x22164x)) + ((n_n4440) & (n_n4434) & (n_n4442) & (n_n4443) & (x22164x)));
	assign n_n1112 = (((!n_n4448) & (!n_n4450) & (!x368x) & (!n_n3889) & (x32x)) + ((!n_n4448) & (!n_n4450) & (!x368x) & (n_n3889) & (!x32x)) + ((!n_n4448) & (!n_n4450) & (!x368x) & (n_n3889) & (x32x)) + ((!n_n4448) & (!n_n4450) & (x368x) & (!n_n3889) & (!x32x)) + ((!n_n4448) & (!n_n4450) & (x368x) & (!n_n3889) & (x32x)) + ((!n_n4448) & (!n_n4450) & (x368x) & (n_n3889) & (!x32x)) + ((!n_n4448) & (!n_n4450) & (x368x) & (n_n3889) & (x32x)) + ((!n_n4448) & (n_n4450) & (!x368x) & (!n_n3889) & (!x32x)) + ((!n_n4448) & (n_n4450) & (!x368x) & (!n_n3889) & (x32x)) + ((!n_n4448) & (n_n4450) & (!x368x) & (n_n3889) & (!x32x)) + ((!n_n4448) & (n_n4450) & (!x368x) & (n_n3889) & (x32x)) + ((!n_n4448) & (n_n4450) & (x368x) & (!n_n3889) & (!x32x)) + ((!n_n4448) & (n_n4450) & (x368x) & (!n_n3889) & (x32x)) + ((!n_n4448) & (n_n4450) & (x368x) & (n_n3889) & (!x32x)) + ((!n_n4448) & (n_n4450) & (x368x) & (n_n3889) & (x32x)) + ((n_n4448) & (!n_n4450) & (!x368x) & (!n_n3889) & (!x32x)) + ((n_n4448) & (!n_n4450) & (!x368x) & (!n_n3889) & (x32x)) + ((n_n4448) & (!n_n4450) & (!x368x) & (n_n3889) & (!x32x)) + ((n_n4448) & (!n_n4450) & (!x368x) & (n_n3889) & (x32x)) + ((n_n4448) & (!n_n4450) & (x368x) & (!n_n3889) & (!x32x)) + ((n_n4448) & (!n_n4450) & (x368x) & (!n_n3889) & (x32x)) + ((n_n4448) & (!n_n4450) & (x368x) & (n_n3889) & (!x32x)) + ((n_n4448) & (!n_n4450) & (x368x) & (n_n3889) & (x32x)) + ((n_n4448) & (n_n4450) & (!x368x) & (!n_n3889) & (!x32x)) + ((n_n4448) & (n_n4450) & (!x368x) & (!n_n3889) & (x32x)) + ((n_n4448) & (n_n4450) & (!x368x) & (n_n3889) & (!x32x)) + ((n_n4448) & (n_n4450) & (!x368x) & (n_n3889) & (x32x)) + ((n_n4448) & (n_n4450) & (x368x) & (!n_n3889) & (!x32x)) + ((n_n4448) & (n_n4450) & (x368x) & (!n_n3889) & (x32x)) + ((n_n4448) & (n_n4450) & (x368x) & (n_n3889) & (!x32x)) + ((n_n4448) & (n_n4450) & (x368x) & (n_n3889) & (x32x)));
	assign x11528x = (((!x37x) & (!x84x) & (!n_n4428) & (!x79x) & (x11524x)) + ((!x37x) & (!x84x) & (!n_n4428) & (x79x) & (!x11524x)) + ((!x37x) & (!x84x) & (!n_n4428) & (x79x) & (x11524x)) + ((!x37x) & (!x84x) & (n_n4428) & (!x79x) & (!x11524x)) + ((!x37x) & (!x84x) & (n_n4428) & (!x79x) & (x11524x)) + ((!x37x) & (!x84x) & (n_n4428) & (x79x) & (!x11524x)) + ((!x37x) & (!x84x) & (n_n4428) & (x79x) & (x11524x)) + ((!x37x) & (x84x) & (!n_n4428) & (!x79x) & (!x11524x)) + ((!x37x) & (x84x) & (!n_n4428) & (!x79x) & (x11524x)) + ((!x37x) & (x84x) & (!n_n4428) & (x79x) & (!x11524x)) + ((!x37x) & (x84x) & (!n_n4428) & (x79x) & (x11524x)) + ((!x37x) & (x84x) & (n_n4428) & (!x79x) & (!x11524x)) + ((!x37x) & (x84x) & (n_n4428) & (!x79x) & (x11524x)) + ((!x37x) & (x84x) & (n_n4428) & (x79x) & (!x11524x)) + ((!x37x) & (x84x) & (n_n4428) & (x79x) & (x11524x)) + ((x37x) & (!x84x) & (!n_n4428) & (!x79x) & (!x11524x)) + ((x37x) & (!x84x) & (!n_n4428) & (!x79x) & (x11524x)) + ((x37x) & (!x84x) & (!n_n4428) & (x79x) & (!x11524x)) + ((x37x) & (!x84x) & (!n_n4428) & (x79x) & (x11524x)) + ((x37x) & (!x84x) & (n_n4428) & (!x79x) & (!x11524x)) + ((x37x) & (!x84x) & (n_n4428) & (!x79x) & (x11524x)) + ((x37x) & (!x84x) & (n_n4428) & (x79x) & (!x11524x)) + ((x37x) & (!x84x) & (n_n4428) & (x79x) & (x11524x)) + ((x37x) & (x84x) & (!n_n4428) & (!x79x) & (!x11524x)) + ((x37x) & (x84x) & (!n_n4428) & (!x79x) & (x11524x)) + ((x37x) & (x84x) & (!n_n4428) & (x79x) & (!x11524x)) + ((x37x) & (x84x) & (!n_n4428) & (x79x) & (x11524x)) + ((x37x) & (x84x) & (n_n4428) & (!x79x) & (!x11524x)) + ((x37x) & (x84x) & (n_n4428) & (!x79x) & (x11524x)) + ((x37x) & (x84x) & (n_n4428) & (x79x) & (!x11524x)) + ((x37x) & (x84x) & (n_n4428) & (x79x) & (x11524x)));
	assign x11530x = (((!n_n1113) & (!n_n1112) & (x11528x)) + ((!n_n1113) & (n_n1112) & (!x11528x)) + ((!n_n1113) & (n_n1112) & (x11528x)) + ((n_n1113) & (!n_n1112) & (!x11528x)) + ((n_n1113) & (!n_n1112) & (x11528x)) + ((n_n1113) & (n_n1112) & (!x11528x)) + ((n_n1113) & (n_n1112) & (x11528x)));
	assign n_n1107 = (((!x13x) & (!x572x) & (!x129x) & (!x308x) & (!x22163x)) + ((!x13x) & (!x572x) & (!x129x) & (x308x) & (!x22163x)) + ((!x13x) & (!x572x) & (!x129x) & (x308x) & (x22163x)) + ((!x13x) & (!x572x) & (x129x) & (!x308x) & (!x22163x)) + ((!x13x) & (!x572x) & (x129x) & (!x308x) & (x22163x)) + ((!x13x) & (!x572x) & (x129x) & (x308x) & (!x22163x)) + ((!x13x) & (!x572x) & (x129x) & (x308x) & (x22163x)) + ((!x13x) & (x572x) & (!x129x) & (!x308x) & (!x22163x)) + ((!x13x) & (x572x) & (!x129x) & (x308x) & (!x22163x)) + ((!x13x) & (x572x) & (!x129x) & (x308x) & (x22163x)) + ((!x13x) & (x572x) & (x129x) & (!x308x) & (!x22163x)) + ((!x13x) & (x572x) & (x129x) & (!x308x) & (x22163x)) + ((!x13x) & (x572x) & (x129x) & (x308x) & (!x22163x)) + ((!x13x) & (x572x) & (x129x) & (x308x) & (x22163x)) + ((x13x) & (!x572x) & (!x129x) & (!x308x) & (!x22163x)) + ((x13x) & (!x572x) & (!x129x) & (x308x) & (!x22163x)) + ((x13x) & (!x572x) & (!x129x) & (x308x) & (x22163x)) + ((x13x) & (!x572x) & (x129x) & (!x308x) & (!x22163x)) + ((x13x) & (!x572x) & (x129x) & (!x308x) & (x22163x)) + ((x13x) & (!x572x) & (x129x) & (x308x) & (!x22163x)) + ((x13x) & (!x572x) & (x129x) & (x308x) & (x22163x)) + ((x13x) & (x572x) & (!x129x) & (!x308x) & (!x22163x)) + ((x13x) & (x572x) & (!x129x) & (!x308x) & (x22163x)) + ((x13x) & (x572x) & (!x129x) & (x308x) & (!x22163x)) + ((x13x) & (x572x) & (!x129x) & (x308x) & (x22163x)) + ((x13x) & (x572x) & (x129x) & (!x308x) & (!x22163x)) + ((x13x) & (x572x) & (x129x) & (!x308x) & (x22163x)) + ((x13x) & (x572x) & (x129x) & (x308x) & (!x22163x)) + ((x13x) & (x572x) & (x129x) & (x308x) & (x22163x)));
	assign x11501x = (((!x130x) & (!n_n4524) & (!x170x) & (!n_n4492) & (!x22162x)) + ((!x130x) & (!n_n4524) & (!x170x) & (n_n4492) & (!x22162x)) + ((!x130x) & (!n_n4524) & (!x170x) & (n_n4492) & (x22162x)) + ((!x130x) & (!n_n4524) & (x170x) & (!n_n4492) & (!x22162x)) + ((!x130x) & (!n_n4524) & (x170x) & (!n_n4492) & (x22162x)) + ((!x130x) & (!n_n4524) & (x170x) & (n_n4492) & (!x22162x)) + ((!x130x) & (!n_n4524) & (x170x) & (n_n4492) & (x22162x)) + ((!x130x) & (n_n4524) & (!x170x) & (!n_n4492) & (!x22162x)) + ((!x130x) & (n_n4524) & (!x170x) & (!n_n4492) & (x22162x)) + ((!x130x) & (n_n4524) & (!x170x) & (n_n4492) & (!x22162x)) + ((!x130x) & (n_n4524) & (!x170x) & (n_n4492) & (x22162x)) + ((!x130x) & (n_n4524) & (x170x) & (!n_n4492) & (!x22162x)) + ((!x130x) & (n_n4524) & (x170x) & (!n_n4492) & (x22162x)) + ((!x130x) & (n_n4524) & (x170x) & (n_n4492) & (!x22162x)) + ((!x130x) & (n_n4524) & (x170x) & (n_n4492) & (x22162x)) + ((x130x) & (!n_n4524) & (!x170x) & (!n_n4492) & (!x22162x)) + ((x130x) & (!n_n4524) & (!x170x) & (!n_n4492) & (x22162x)) + ((x130x) & (!n_n4524) & (!x170x) & (n_n4492) & (!x22162x)) + ((x130x) & (!n_n4524) & (!x170x) & (n_n4492) & (x22162x)) + ((x130x) & (!n_n4524) & (x170x) & (!n_n4492) & (!x22162x)) + ((x130x) & (!n_n4524) & (x170x) & (!n_n4492) & (x22162x)) + ((x130x) & (!n_n4524) & (x170x) & (n_n4492) & (!x22162x)) + ((x130x) & (!n_n4524) & (x170x) & (n_n4492) & (x22162x)) + ((x130x) & (n_n4524) & (!x170x) & (!n_n4492) & (!x22162x)) + ((x130x) & (n_n4524) & (!x170x) & (!n_n4492) & (x22162x)) + ((x130x) & (n_n4524) & (!x170x) & (n_n4492) & (!x22162x)) + ((x130x) & (n_n4524) & (!x170x) & (n_n4492) & (x22162x)) + ((x130x) & (n_n4524) & (x170x) & (!n_n4492) & (!x22162x)) + ((x130x) & (n_n4524) & (x170x) & (!n_n4492) & (x22162x)) + ((x130x) & (n_n4524) & (x170x) & (n_n4492) & (!x22162x)) + ((x130x) & (n_n4524) & (x170x) & (n_n4492) & (x22162x)));
	assign n_n1038 = (((!n_n1111) & (!x206x) & (!x11516x) & (x11517x)) + ((!n_n1111) & (!x206x) & (x11516x) & (!x11517x)) + ((!n_n1111) & (!x206x) & (x11516x) & (x11517x)) + ((!n_n1111) & (x206x) & (!x11516x) & (!x11517x)) + ((!n_n1111) & (x206x) & (!x11516x) & (x11517x)) + ((!n_n1111) & (x206x) & (x11516x) & (!x11517x)) + ((!n_n1111) & (x206x) & (x11516x) & (x11517x)) + ((n_n1111) & (!x206x) & (!x11516x) & (!x11517x)) + ((n_n1111) & (!x206x) & (!x11516x) & (x11517x)) + ((n_n1111) & (!x206x) & (x11516x) & (!x11517x)) + ((n_n1111) & (!x206x) & (x11516x) & (x11517x)) + ((n_n1111) & (x206x) & (!x11516x) & (!x11517x)) + ((n_n1111) & (x206x) & (!x11516x) & (x11517x)) + ((n_n1111) & (x206x) & (x11516x) & (!x11517x)) + ((n_n1111) & (x206x) & (x11516x) & (x11517x)));
	assign x11500x = (((!n_n4498) & (!n_n4499) & (!x307x) & (!x162x) & (x347x)) + ((!n_n4498) & (!n_n4499) & (!x307x) & (x162x) & (!x347x)) + ((!n_n4498) & (!n_n4499) & (!x307x) & (x162x) & (x347x)) + ((!n_n4498) & (!n_n4499) & (x307x) & (!x162x) & (!x347x)) + ((!n_n4498) & (!n_n4499) & (x307x) & (!x162x) & (x347x)) + ((!n_n4498) & (!n_n4499) & (x307x) & (x162x) & (!x347x)) + ((!n_n4498) & (!n_n4499) & (x307x) & (x162x) & (x347x)) + ((!n_n4498) & (n_n4499) & (!x307x) & (!x162x) & (!x347x)) + ((!n_n4498) & (n_n4499) & (!x307x) & (!x162x) & (x347x)) + ((!n_n4498) & (n_n4499) & (!x307x) & (x162x) & (!x347x)) + ((!n_n4498) & (n_n4499) & (!x307x) & (x162x) & (x347x)) + ((!n_n4498) & (n_n4499) & (x307x) & (!x162x) & (!x347x)) + ((!n_n4498) & (n_n4499) & (x307x) & (!x162x) & (x347x)) + ((!n_n4498) & (n_n4499) & (x307x) & (x162x) & (!x347x)) + ((!n_n4498) & (n_n4499) & (x307x) & (x162x) & (x347x)) + ((n_n4498) & (!n_n4499) & (!x307x) & (!x162x) & (!x347x)) + ((n_n4498) & (!n_n4499) & (!x307x) & (!x162x) & (x347x)) + ((n_n4498) & (!n_n4499) & (!x307x) & (x162x) & (!x347x)) + ((n_n4498) & (!n_n4499) & (!x307x) & (x162x) & (x347x)) + ((n_n4498) & (!n_n4499) & (x307x) & (!x162x) & (!x347x)) + ((n_n4498) & (!n_n4499) & (x307x) & (!x162x) & (x347x)) + ((n_n4498) & (!n_n4499) & (x307x) & (x162x) & (!x347x)) + ((n_n4498) & (!n_n4499) & (x307x) & (x162x) & (x347x)) + ((n_n4498) & (n_n4499) & (!x307x) & (!x162x) & (!x347x)) + ((n_n4498) & (n_n4499) & (!x307x) & (!x162x) & (x347x)) + ((n_n4498) & (n_n4499) & (!x307x) & (x162x) & (!x347x)) + ((n_n4498) & (n_n4499) & (!x307x) & (x162x) & (x347x)) + ((n_n4498) & (n_n4499) & (x307x) & (!x162x) & (!x347x)) + ((n_n4498) & (n_n4499) & (x307x) & (!x162x) & (x347x)) + ((n_n4498) & (n_n4499) & (x307x) & (x162x) & (!x347x)) + ((n_n4498) & (n_n4499) & (x307x) & (x162x) & (x347x)));
	assign n_n4243 = (((!i_9_) & (n_n455) & (n_n473) & (!n_n532) & (n_n534)) + ((!i_9_) & (n_n455) & (n_n473) & (n_n532) & (!n_n534)) + ((!i_9_) & (n_n455) & (n_n473) & (n_n532) & (n_n534)) + ((i_9_) & (n_n455) & (n_n473) & (n_n532) & (!n_n534)) + ((i_9_) & (n_n455) & (n_n473) & (n_n532) & (n_n534)));
	assign n_n1104 = (((!n_n4542) & (!x201x) & (!n_n4549) & (!n_n4551) & (!x22161x)) + ((!n_n4542) & (!x201x) & (!n_n4549) & (n_n4551) & (!x22161x)) + ((!n_n4542) & (!x201x) & (!n_n4549) & (n_n4551) & (x22161x)) + ((!n_n4542) & (!x201x) & (n_n4549) & (!n_n4551) & (!x22161x)) + ((!n_n4542) & (!x201x) & (n_n4549) & (!n_n4551) & (x22161x)) + ((!n_n4542) & (!x201x) & (n_n4549) & (n_n4551) & (!x22161x)) + ((!n_n4542) & (!x201x) & (n_n4549) & (n_n4551) & (x22161x)) + ((!n_n4542) & (x201x) & (!n_n4549) & (!n_n4551) & (!x22161x)) + ((!n_n4542) & (x201x) & (!n_n4549) & (!n_n4551) & (x22161x)) + ((!n_n4542) & (x201x) & (!n_n4549) & (n_n4551) & (!x22161x)) + ((!n_n4542) & (x201x) & (!n_n4549) & (n_n4551) & (x22161x)) + ((!n_n4542) & (x201x) & (n_n4549) & (!n_n4551) & (!x22161x)) + ((!n_n4542) & (x201x) & (n_n4549) & (!n_n4551) & (x22161x)) + ((!n_n4542) & (x201x) & (n_n4549) & (n_n4551) & (!x22161x)) + ((!n_n4542) & (x201x) & (n_n4549) & (n_n4551) & (x22161x)) + ((n_n4542) & (!x201x) & (!n_n4549) & (!n_n4551) & (!x22161x)) + ((n_n4542) & (!x201x) & (!n_n4549) & (!n_n4551) & (x22161x)) + ((n_n4542) & (!x201x) & (!n_n4549) & (n_n4551) & (!x22161x)) + ((n_n4542) & (!x201x) & (!n_n4549) & (n_n4551) & (x22161x)) + ((n_n4542) & (!x201x) & (n_n4549) & (!n_n4551) & (!x22161x)) + ((n_n4542) & (!x201x) & (n_n4549) & (!n_n4551) & (x22161x)) + ((n_n4542) & (!x201x) & (n_n4549) & (n_n4551) & (!x22161x)) + ((n_n4542) & (!x201x) & (n_n4549) & (n_n4551) & (x22161x)) + ((n_n4542) & (x201x) & (!n_n4549) & (!n_n4551) & (!x22161x)) + ((n_n4542) & (x201x) & (!n_n4549) & (!n_n4551) & (x22161x)) + ((n_n4542) & (x201x) & (!n_n4549) & (n_n4551) & (!x22161x)) + ((n_n4542) & (x201x) & (!n_n4549) & (n_n4551) & (x22161x)) + ((n_n4542) & (x201x) & (n_n4549) & (!n_n4551) & (!x22161x)) + ((n_n4542) & (x201x) & (n_n4549) & (!n_n4551) & (x22161x)) + ((n_n4542) & (x201x) & (n_n4549) & (n_n4551) & (!x22161x)) + ((n_n4542) & (x201x) & (n_n4549) & (n_n4551) & (x22161x)));
	assign n_n1103 = (((!n_n4557) & (!n_n4561) & (!x213x) & (x11542x)) + ((!n_n4557) & (!n_n4561) & (x213x) & (!x11542x)) + ((!n_n4557) & (!n_n4561) & (x213x) & (x11542x)) + ((!n_n4557) & (n_n4561) & (!x213x) & (!x11542x)) + ((!n_n4557) & (n_n4561) & (!x213x) & (x11542x)) + ((!n_n4557) & (n_n4561) & (x213x) & (!x11542x)) + ((!n_n4557) & (n_n4561) & (x213x) & (x11542x)) + ((n_n4557) & (!n_n4561) & (!x213x) & (!x11542x)) + ((n_n4557) & (!n_n4561) & (!x213x) & (x11542x)) + ((n_n4557) & (!n_n4561) & (x213x) & (!x11542x)) + ((n_n4557) & (!n_n4561) & (x213x) & (x11542x)) + ((n_n4557) & (n_n4561) & (!x213x) & (!x11542x)) + ((n_n4557) & (n_n4561) & (!x213x) & (x11542x)) + ((n_n4557) & (n_n4561) & (x213x) & (!x11542x)) + ((n_n4557) & (n_n4561) & (x213x) & (x11542x)));
	assign n_n3875 = (((!i_9_) & (n_n482) & (n_n455) & (!n_n520) & (x20x)) + ((!i_9_) & (n_n482) & (n_n455) & (n_n520) & (!x20x)) + ((!i_9_) & (n_n482) & (n_n455) & (n_n520) & (x20x)) + ((i_9_) & (n_n482) & (n_n455) & (!n_n520) & (x20x)) + ((i_9_) & (n_n482) & (n_n455) & (n_n520) & (!x20x)) + ((i_9_) & (n_n482) & (n_n455) & (n_n520) & (x20x)));
	assign x11577x = (((!i_9_) & (!n_n526) & (n_n482) & (n_n455) & (n_n530)) + ((!i_9_) & (n_n526) & (n_n482) & (n_n455) & (!n_n530)) + ((!i_9_) & (n_n526) & (n_n482) & (n_n455) & (n_n530)) + ((i_9_) & (n_n526) & (n_n482) & (n_n455) & (!n_n530)) + ((i_9_) & (n_n526) & (n_n482) & (n_n455) & (n_n530)));
	assign x11581x = (((!n_n4243) & (!n_n1104) & (!n_n1103) & (!n_n3875) & (x11577x)) + ((!n_n4243) & (!n_n1104) & (!n_n1103) & (n_n3875) & (!x11577x)) + ((!n_n4243) & (!n_n1104) & (!n_n1103) & (n_n3875) & (x11577x)) + ((!n_n4243) & (!n_n1104) & (n_n1103) & (!n_n3875) & (!x11577x)) + ((!n_n4243) & (!n_n1104) & (n_n1103) & (!n_n3875) & (x11577x)) + ((!n_n4243) & (!n_n1104) & (n_n1103) & (n_n3875) & (!x11577x)) + ((!n_n4243) & (!n_n1104) & (n_n1103) & (n_n3875) & (x11577x)) + ((!n_n4243) & (n_n1104) & (!n_n1103) & (!n_n3875) & (!x11577x)) + ((!n_n4243) & (n_n1104) & (!n_n1103) & (!n_n3875) & (x11577x)) + ((!n_n4243) & (n_n1104) & (!n_n1103) & (n_n3875) & (!x11577x)) + ((!n_n4243) & (n_n1104) & (!n_n1103) & (n_n3875) & (x11577x)) + ((!n_n4243) & (n_n1104) & (n_n1103) & (!n_n3875) & (!x11577x)) + ((!n_n4243) & (n_n1104) & (n_n1103) & (!n_n3875) & (x11577x)) + ((!n_n4243) & (n_n1104) & (n_n1103) & (n_n3875) & (!x11577x)) + ((!n_n4243) & (n_n1104) & (n_n1103) & (n_n3875) & (x11577x)) + ((n_n4243) & (!n_n1104) & (!n_n1103) & (!n_n3875) & (!x11577x)) + ((n_n4243) & (!n_n1104) & (!n_n1103) & (!n_n3875) & (x11577x)) + ((n_n4243) & (!n_n1104) & (!n_n1103) & (n_n3875) & (!x11577x)) + ((n_n4243) & (!n_n1104) & (!n_n1103) & (n_n3875) & (x11577x)) + ((n_n4243) & (!n_n1104) & (n_n1103) & (!n_n3875) & (!x11577x)) + ((n_n4243) & (!n_n1104) & (n_n1103) & (!n_n3875) & (x11577x)) + ((n_n4243) & (!n_n1104) & (n_n1103) & (n_n3875) & (!x11577x)) + ((n_n4243) & (!n_n1104) & (n_n1103) & (n_n3875) & (x11577x)) + ((n_n4243) & (n_n1104) & (!n_n1103) & (!n_n3875) & (!x11577x)) + ((n_n4243) & (n_n1104) & (!n_n1103) & (!n_n3875) & (x11577x)) + ((n_n4243) & (n_n1104) & (!n_n1103) & (n_n3875) & (!x11577x)) + ((n_n4243) & (n_n1104) & (!n_n1103) & (n_n3875) & (x11577x)) + ((n_n4243) & (n_n1104) & (n_n1103) & (!n_n3875) & (!x11577x)) + ((n_n4243) & (n_n1104) & (n_n1103) & (!n_n3875) & (x11577x)) + ((n_n4243) & (n_n1104) & (n_n1103) & (n_n3875) & (!x11577x)) + ((n_n4243) & (n_n1104) & (n_n1103) & (n_n3875) & (x11577x)));
	assign n_n1034 = (((!n_n1099) & (!x11555x) & (!x11556x) & (x11557x)) + ((!n_n1099) & (!x11555x) & (x11556x) & (!x11557x)) + ((!n_n1099) & (!x11555x) & (x11556x) & (x11557x)) + ((!n_n1099) & (x11555x) & (!x11556x) & (!x11557x)) + ((!n_n1099) & (x11555x) & (!x11556x) & (x11557x)) + ((!n_n1099) & (x11555x) & (x11556x) & (!x11557x)) + ((!n_n1099) & (x11555x) & (x11556x) & (x11557x)) + ((n_n1099) & (!x11555x) & (!x11556x) & (!x11557x)) + ((n_n1099) & (!x11555x) & (!x11556x) & (x11557x)) + ((n_n1099) & (!x11555x) & (x11556x) & (!x11557x)) + ((n_n1099) & (!x11555x) & (x11556x) & (x11557x)) + ((n_n1099) & (x11555x) & (!x11556x) & (!x11557x)) + ((n_n1099) & (x11555x) & (!x11556x) & (x11557x)) + ((n_n1099) & (x11555x) & (x11556x) & (!x11557x)) + ((n_n1099) & (x11555x) & (x11556x) & (x11557x)));
	assign n_n1035 = (((!n_n1100) & (!x224x) & (!x11572x) & (x11573x)) + ((!n_n1100) & (!x224x) & (x11572x) & (!x11573x)) + ((!n_n1100) & (!x224x) & (x11572x) & (x11573x)) + ((!n_n1100) & (x224x) & (!x11572x) & (!x11573x)) + ((!n_n1100) & (x224x) & (!x11572x) & (x11573x)) + ((!n_n1100) & (x224x) & (x11572x) & (!x11573x)) + ((!n_n1100) & (x224x) & (x11572x) & (x11573x)) + ((n_n1100) & (!x224x) & (!x11572x) & (!x11573x)) + ((n_n1100) & (!x224x) & (!x11572x) & (x11573x)) + ((n_n1100) & (!x224x) & (x11572x) & (!x11573x)) + ((n_n1100) & (!x224x) & (x11572x) & (x11573x)) + ((n_n1100) & (x224x) & (!x11572x) & (!x11573x)) + ((n_n1100) & (x224x) & (!x11572x) & (x11573x)) + ((n_n1100) & (x224x) & (x11572x) & (!x11573x)) + ((n_n1100) & (x224x) & (x11572x) & (x11573x)));
	assign n_n1123 = (((!n_n4317) & (!n_n4318) & (!n_n4320) & (!n_n4316) & (x11587x)) + ((!n_n4317) & (!n_n4318) & (!n_n4320) & (n_n4316) & (!x11587x)) + ((!n_n4317) & (!n_n4318) & (!n_n4320) & (n_n4316) & (x11587x)) + ((!n_n4317) & (!n_n4318) & (n_n4320) & (!n_n4316) & (!x11587x)) + ((!n_n4317) & (!n_n4318) & (n_n4320) & (!n_n4316) & (x11587x)) + ((!n_n4317) & (!n_n4318) & (n_n4320) & (n_n4316) & (!x11587x)) + ((!n_n4317) & (!n_n4318) & (n_n4320) & (n_n4316) & (x11587x)) + ((!n_n4317) & (n_n4318) & (!n_n4320) & (!n_n4316) & (!x11587x)) + ((!n_n4317) & (n_n4318) & (!n_n4320) & (!n_n4316) & (x11587x)) + ((!n_n4317) & (n_n4318) & (!n_n4320) & (n_n4316) & (!x11587x)) + ((!n_n4317) & (n_n4318) & (!n_n4320) & (n_n4316) & (x11587x)) + ((!n_n4317) & (n_n4318) & (n_n4320) & (!n_n4316) & (!x11587x)) + ((!n_n4317) & (n_n4318) & (n_n4320) & (!n_n4316) & (x11587x)) + ((!n_n4317) & (n_n4318) & (n_n4320) & (n_n4316) & (!x11587x)) + ((!n_n4317) & (n_n4318) & (n_n4320) & (n_n4316) & (x11587x)) + ((n_n4317) & (!n_n4318) & (!n_n4320) & (!n_n4316) & (!x11587x)) + ((n_n4317) & (!n_n4318) & (!n_n4320) & (!n_n4316) & (x11587x)) + ((n_n4317) & (!n_n4318) & (!n_n4320) & (n_n4316) & (!x11587x)) + ((n_n4317) & (!n_n4318) & (!n_n4320) & (n_n4316) & (x11587x)) + ((n_n4317) & (!n_n4318) & (n_n4320) & (!n_n4316) & (!x11587x)) + ((n_n4317) & (!n_n4318) & (n_n4320) & (!n_n4316) & (x11587x)) + ((n_n4317) & (!n_n4318) & (n_n4320) & (n_n4316) & (!x11587x)) + ((n_n4317) & (!n_n4318) & (n_n4320) & (n_n4316) & (x11587x)) + ((n_n4317) & (n_n4318) & (!n_n4320) & (!n_n4316) & (!x11587x)) + ((n_n4317) & (n_n4318) & (!n_n4320) & (!n_n4316) & (x11587x)) + ((n_n4317) & (n_n4318) & (!n_n4320) & (n_n4316) & (!x11587x)) + ((n_n4317) & (n_n4318) & (!n_n4320) & (n_n4316) & (x11587x)) + ((n_n4317) & (n_n4318) & (n_n4320) & (!n_n4316) & (!x11587x)) + ((n_n4317) & (n_n4318) & (n_n4320) & (!n_n4316) & (x11587x)) + ((n_n4317) & (n_n4318) & (n_n4320) & (n_n4316) & (!x11587x)) + ((n_n4317) & (n_n4318) & (n_n4320) & (n_n4316) & (x11587x)));
	assign n_n1040 = (((!n_n1117) & (!n_n1115) & (x11604x)) + ((!n_n1117) & (n_n1115) & (!x11604x)) + ((!n_n1117) & (n_n1115) & (x11604x)) + ((n_n1117) & (!n_n1115) & (!x11604x)) + ((n_n1117) & (!n_n1115) & (x11604x)) + ((n_n1117) & (n_n1115) & (!x11604x)) + ((n_n1117) & (n_n1115) & (x11604x)));
	assign n_n1041 = (((!x300x) & (!n_n1120) & (!n_n3176) & (!x11618x) & (x161x)) + ((!x300x) & (!n_n1120) & (!n_n3176) & (x11618x) & (!x161x)) + ((!x300x) & (!n_n1120) & (!n_n3176) & (x11618x) & (x161x)) + ((!x300x) & (!n_n1120) & (n_n3176) & (!x11618x) & (!x161x)) + ((!x300x) & (!n_n1120) & (n_n3176) & (!x11618x) & (x161x)) + ((!x300x) & (!n_n1120) & (n_n3176) & (x11618x) & (!x161x)) + ((!x300x) & (!n_n1120) & (n_n3176) & (x11618x) & (x161x)) + ((!x300x) & (n_n1120) & (!n_n3176) & (!x11618x) & (!x161x)) + ((!x300x) & (n_n1120) & (!n_n3176) & (!x11618x) & (x161x)) + ((!x300x) & (n_n1120) & (!n_n3176) & (x11618x) & (!x161x)) + ((!x300x) & (n_n1120) & (!n_n3176) & (x11618x) & (x161x)) + ((!x300x) & (n_n1120) & (n_n3176) & (!x11618x) & (!x161x)) + ((!x300x) & (n_n1120) & (n_n3176) & (!x11618x) & (x161x)) + ((!x300x) & (n_n1120) & (n_n3176) & (x11618x) & (!x161x)) + ((!x300x) & (n_n1120) & (n_n3176) & (x11618x) & (x161x)) + ((x300x) & (!n_n1120) & (!n_n3176) & (!x11618x) & (!x161x)) + ((x300x) & (!n_n1120) & (!n_n3176) & (!x11618x) & (x161x)) + ((x300x) & (!n_n1120) & (!n_n3176) & (x11618x) & (!x161x)) + ((x300x) & (!n_n1120) & (!n_n3176) & (x11618x) & (x161x)) + ((x300x) & (!n_n1120) & (n_n3176) & (!x11618x) & (!x161x)) + ((x300x) & (!n_n1120) & (n_n3176) & (!x11618x) & (x161x)) + ((x300x) & (!n_n1120) & (n_n3176) & (x11618x) & (!x161x)) + ((x300x) & (!n_n1120) & (n_n3176) & (x11618x) & (x161x)) + ((x300x) & (n_n1120) & (!n_n3176) & (!x11618x) & (!x161x)) + ((x300x) & (n_n1120) & (!n_n3176) & (!x11618x) & (x161x)) + ((x300x) & (n_n1120) & (!n_n3176) & (x11618x) & (!x161x)) + ((x300x) & (n_n1120) & (!n_n3176) & (x11618x) & (x161x)) + ((x300x) & (n_n1120) & (n_n3176) & (!x11618x) & (!x161x)) + ((x300x) & (n_n1120) & (n_n3176) & (!x11618x) & (x161x)) + ((x300x) & (n_n1120) & (n_n3176) & (x11618x) & (!x161x)) + ((x300x) & (n_n1120) & (n_n3176) & (x11618x) & (x161x)));
	assign n_n1121 = (((!n_n4337) & (!n_n4344) & (!n_n4335) & (!x11620x) & (!x22150x)) + ((!n_n4337) & (!n_n4344) & (!n_n4335) & (x11620x) & (!x22150x)) + ((!n_n4337) & (!n_n4344) & (!n_n4335) & (x11620x) & (x22150x)) + ((!n_n4337) & (!n_n4344) & (n_n4335) & (!x11620x) & (!x22150x)) + ((!n_n4337) & (!n_n4344) & (n_n4335) & (!x11620x) & (x22150x)) + ((!n_n4337) & (!n_n4344) & (n_n4335) & (x11620x) & (!x22150x)) + ((!n_n4337) & (!n_n4344) & (n_n4335) & (x11620x) & (x22150x)) + ((!n_n4337) & (n_n4344) & (!n_n4335) & (!x11620x) & (!x22150x)) + ((!n_n4337) & (n_n4344) & (!n_n4335) & (!x11620x) & (x22150x)) + ((!n_n4337) & (n_n4344) & (!n_n4335) & (x11620x) & (!x22150x)) + ((!n_n4337) & (n_n4344) & (!n_n4335) & (x11620x) & (x22150x)) + ((!n_n4337) & (n_n4344) & (n_n4335) & (!x11620x) & (!x22150x)) + ((!n_n4337) & (n_n4344) & (n_n4335) & (!x11620x) & (x22150x)) + ((!n_n4337) & (n_n4344) & (n_n4335) & (x11620x) & (!x22150x)) + ((!n_n4337) & (n_n4344) & (n_n4335) & (x11620x) & (x22150x)) + ((n_n4337) & (!n_n4344) & (!n_n4335) & (!x11620x) & (!x22150x)) + ((n_n4337) & (!n_n4344) & (!n_n4335) & (!x11620x) & (x22150x)) + ((n_n4337) & (!n_n4344) & (!n_n4335) & (x11620x) & (!x22150x)) + ((n_n4337) & (!n_n4344) & (!n_n4335) & (x11620x) & (x22150x)) + ((n_n4337) & (!n_n4344) & (n_n4335) & (!x11620x) & (!x22150x)) + ((n_n4337) & (!n_n4344) & (n_n4335) & (!x11620x) & (x22150x)) + ((n_n4337) & (!n_n4344) & (n_n4335) & (x11620x) & (!x22150x)) + ((n_n4337) & (!n_n4344) & (n_n4335) & (x11620x) & (x22150x)) + ((n_n4337) & (n_n4344) & (!n_n4335) & (!x11620x) & (!x22150x)) + ((n_n4337) & (n_n4344) & (!n_n4335) & (!x11620x) & (x22150x)) + ((n_n4337) & (n_n4344) & (!n_n4335) & (x11620x) & (!x22150x)) + ((n_n4337) & (n_n4344) & (!n_n4335) & (x11620x) & (x22150x)) + ((n_n4337) & (n_n4344) & (n_n4335) & (!x11620x) & (!x22150x)) + ((n_n4337) & (n_n4344) & (n_n4335) & (!x11620x) & (x22150x)) + ((n_n4337) & (n_n4344) & (n_n4335) & (x11620x) & (!x22150x)) + ((n_n4337) & (n_n4344) & (n_n4335) & (x11620x) & (x22150x)));
	assign x11632x = (((!n_n4327) & (!n_n4331) & (!x410x) & (x11631x)) + ((!n_n4327) & (!n_n4331) & (x410x) & (!x11631x)) + ((!n_n4327) & (!n_n4331) & (x410x) & (x11631x)) + ((!n_n4327) & (n_n4331) & (!x410x) & (!x11631x)) + ((!n_n4327) & (n_n4331) & (!x410x) & (x11631x)) + ((!n_n4327) & (n_n4331) & (x410x) & (!x11631x)) + ((!n_n4327) & (n_n4331) & (x410x) & (x11631x)) + ((n_n4327) & (!n_n4331) & (!x410x) & (!x11631x)) + ((n_n4327) & (!n_n4331) & (!x410x) & (x11631x)) + ((n_n4327) & (!n_n4331) & (x410x) & (!x11631x)) + ((n_n4327) & (!n_n4331) & (x410x) & (x11631x)) + ((n_n4327) & (n_n4331) & (!x410x) & (!x11631x)) + ((n_n4327) & (n_n4331) & (!x410x) & (x11631x)) + ((n_n4327) & (n_n4331) & (x410x) & (!x11631x)) + ((n_n4327) & (n_n4331) & (x410x) & (x11631x)));
	assign n_n1015 = (((!n_n1123) & (!n_n1040) & (!n_n1041) & (!n_n1121) & (x11632x)) + ((!n_n1123) & (!n_n1040) & (!n_n1041) & (n_n1121) & (!x11632x)) + ((!n_n1123) & (!n_n1040) & (!n_n1041) & (n_n1121) & (x11632x)) + ((!n_n1123) & (!n_n1040) & (n_n1041) & (!n_n1121) & (!x11632x)) + ((!n_n1123) & (!n_n1040) & (n_n1041) & (!n_n1121) & (x11632x)) + ((!n_n1123) & (!n_n1040) & (n_n1041) & (n_n1121) & (!x11632x)) + ((!n_n1123) & (!n_n1040) & (n_n1041) & (n_n1121) & (x11632x)) + ((!n_n1123) & (n_n1040) & (!n_n1041) & (!n_n1121) & (!x11632x)) + ((!n_n1123) & (n_n1040) & (!n_n1041) & (!n_n1121) & (x11632x)) + ((!n_n1123) & (n_n1040) & (!n_n1041) & (n_n1121) & (!x11632x)) + ((!n_n1123) & (n_n1040) & (!n_n1041) & (n_n1121) & (x11632x)) + ((!n_n1123) & (n_n1040) & (n_n1041) & (!n_n1121) & (!x11632x)) + ((!n_n1123) & (n_n1040) & (n_n1041) & (!n_n1121) & (x11632x)) + ((!n_n1123) & (n_n1040) & (n_n1041) & (n_n1121) & (!x11632x)) + ((!n_n1123) & (n_n1040) & (n_n1041) & (n_n1121) & (x11632x)) + ((n_n1123) & (!n_n1040) & (!n_n1041) & (!n_n1121) & (!x11632x)) + ((n_n1123) & (!n_n1040) & (!n_n1041) & (!n_n1121) & (x11632x)) + ((n_n1123) & (!n_n1040) & (!n_n1041) & (n_n1121) & (!x11632x)) + ((n_n1123) & (!n_n1040) & (!n_n1041) & (n_n1121) & (x11632x)) + ((n_n1123) & (!n_n1040) & (n_n1041) & (!n_n1121) & (!x11632x)) + ((n_n1123) & (!n_n1040) & (n_n1041) & (!n_n1121) & (x11632x)) + ((n_n1123) & (!n_n1040) & (n_n1041) & (n_n1121) & (!x11632x)) + ((n_n1123) & (!n_n1040) & (n_n1041) & (n_n1121) & (x11632x)) + ((n_n1123) & (n_n1040) & (!n_n1041) & (!n_n1121) & (!x11632x)) + ((n_n1123) & (n_n1040) & (!n_n1041) & (!n_n1121) & (x11632x)) + ((n_n1123) & (n_n1040) & (!n_n1041) & (n_n1121) & (!x11632x)) + ((n_n1123) & (n_n1040) & (!n_n1041) & (n_n1121) & (x11632x)) + ((n_n1123) & (n_n1040) & (n_n1041) & (!n_n1121) & (!x11632x)) + ((n_n1123) & (n_n1040) & (n_n1041) & (!n_n1121) & (x11632x)) + ((n_n1123) & (n_n1040) & (n_n1041) & (n_n1121) & (!x11632x)) + ((n_n1123) & (n_n1040) & (n_n1041) & (n_n1121) & (x11632x)));
	assign x11736x = (((!x11719x) & (!x11720x) & (!x11726x) & (x11727x)) + ((!x11719x) & (!x11720x) & (x11726x) & (!x11727x)) + ((!x11719x) & (!x11720x) & (x11726x) & (x11727x)) + ((!x11719x) & (x11720x) & (!x11726x) & (!x11727x)) + ((!x11719x) & (x11720x) & (!x11726x) & (x11727x)) + ((!x11719x) & (x11720x) & (x11726x) & (!x11727x)) + ((!x11719x) & (x11720x) & (x11726x) & (x11727x)) + ((x11719x) & (!x11720x) & (!x11726x) & (!x11727x)) + ((x11719x) & (!x11720x) & (!x11726x) & (x11727x)) + ((x11719x) & (!x11720x) & (x11726x) & (!x11727x)) + ((x11719x) & (!x11720x) & (x11726x) & (x11727x)) + ((x11719x) & (x11720x) & (!x11726x) & (!x11727x)) + ((x11719x) & (x11720x) & (!x11726x) & (x11727x)) + ((x11719x) & (x11720x) & (x11726x) & (!x11727x)) + ((x11719x) & (x11720x) & (x11726x) & (x11727x)));
	assign x11734x = (((!x11698x) & (!x11699x) & (!x11732x) & (!x22198x)) + ((!x11698x) & (!x11699x) & (x11732x) & (!x22198x)) + ((!x11698x) & (!x11699x) & (x11732x) & (x22198x)) + ((!x11698x) & (x11699x) & (!x11732x) & (!x22198x)) + ((!x11698x) & (x11699x) & (!x11732x) & (x22198x)) + ((!x11698x) & (x11699x) & (x11732x) & (!x22198x)) + ((!x11698x) & (x11699x) & (x11732x) & (x22198x)) + ((x11698x) & (!x11699x) & (!x11732x) & (!x22198x)) + ((x11698x) & (!x11699x) & (!x11732x) & (x22198x)) + ((x11698x) & (!x11699x) & (x11732x) & (!x22198x)) + ((x11698x) & (!x11699x) & (x11732x) & (x22198x)) + ((x11698x) & (x11699x) & (!x11732x) & (!x22198x)) + ((x11698x) & (x11699x) & (!x11732x) & (x22198x)) + ((x11698x) & (x11699x) & (x11732x) & (!x22198x)) + ((x11698x) & (x11699x) & (x11732x) & (x22198x)));
	assign x11735x = (((!x11705x) & (!x11706x) & (n_n947)) + ((!x11705x) & (x11706x) & (!n_n947)) + ((!x11705x) & (x11706x) & (n_n947)) + ((x11705x) & (!x11706x) & (!n_n947)) + ((x11705x) & (!x11706x) & (n_n947)) + ((x11705x) & (x11706x) & (!n_n947)) + ((x11705x) & (x11706x) & (n_n947)));
	assign x11745x = (((!x11660x) & (!x11661x) & (!x11667x) & (!x11668x) & (x11743x)) + ((!x11660x) & (!x11661x) & (!x11667x) & (x11668x) & (!x11743x)) + ((!x11660x) & (!x11661x) & (!x11667x) & (x11668x) & (x11743x)) + ((!x11660x) & (!x11661x) & (x11667x) & (!x11668x) & (!x11743x)) + ((!x11660x) & (!x11661x) & (x11667x) & (!x11668x) & (x11743x)) + ((!x11660x) & (!x11661x) & (x11667x) & (x11668x) & (!x11743x)) + ((!x11660x) & (!x11661x) & (x11667x) & (x11668x) & (x11743x)) + ((!x11660x) & (x11661x) & (!x11667x) & (!x11668x) & (!x11743x)) + ((!x11660x) & (x11661x) & (!x11667x) & (!x11668x) & (x11743x)) + ((!x11660x) & (x11661x) & (!x11667x) & (x11668x) & (!x11743x)) + ((!x11660x) & (x11661x) & (!x11667x) & (x11668x) & (x11743x)) + ((!x11660x) & (x11661x) & (x11667x) & (!x11668x) & (!x11743x)) + ((!x11660x) & (x11661x) & (x11667x) & (!x11668x) & (x11743x)) + ((!x11660x) & (x11661x) & (x11667x) & (x11668x) & (!x11743x)) + ((!x11660x) & (x11661x) & (x11667x) & (x11668x) & (x11743x)) + ((x11660x) & (!x11661x) & (!x11667x) & (!x11668x) & (!x11743x)) + ((x11660x) & (!x11661x) & (!x11667x) & (!x11668x) & (x11743x)) + ((x11660x) & (!x11661x) & (!x11667x) & (x11668x) & (!x11743x)) + ((x11660x) & (!x11661x) & (!x11667x) & (x11668x) & (x11743x)) + ((x11660x) & (!x11661x) & (x11667x) & (!x11668x) & (!x11743x)) + ((x11660x) & (!x11661x) & (x11667x) & (!x11668x) & (x11743x)) + ((x11660x) & (!x11661x) & (x11667x) & (x11668x) & (!x11743x)) + ((x11660x) & (!x11661x) & (x11667x) & (x11668x) & (x11743x)) + ((x11660x) & (x11661x) & (!x11667x) & (!x11668x) & (!x11743x)) + ((x11660x) & (x11661x) & (!x11667x) & (!x11668x) & (x11743x)) + ((x11660x) & (x11661x) & (!x11667x) & (x11668x) & (!x11743x)) + ((x11660x) & (x11661x) & (!x11667x) & (x11668x) & (x11743x)) + ((x11660x) & (x11661x) & (x11667x) & (!x11668x) & (!x11743x)) + ((x11660x) & (x11661x) & (x11667x) & (!x11668x) & (x11743x)) + ((x11660x) & (x11661x) & (x11667x) & (x11668x) & (!x11743x)) + ((x11660x) & (x11661x) & (x11667x) & (x11668x) & (x11743x)));
	assign x11747x = (((!x11736x) & (!x11734x) & (!x11735x) & (x11745x)) + ((!x11736x) & (!x11734x) & (x11735x) & (!x11745x)) + ((!x11736x) & (!x11734x) & (x11735x) & (x11745x)) + ((!x11736x) & (x11734x) & (!x11735x) & (!x11745x)) + ((!x11736x) & (x11734x) & (!x11735x) & (x11745x)) + ((!x11736x) & (x11734x) & (x11735x) & (!x11745x)) + ((!x11736x) & (x11734x) & (x11735x) & (x11745x)) + ((x11736x) & (!x11734x) & (!x11735x) & (!x11745x)) + ((x11736x) & (!x11734x) & (!x11735x) & (x11745x)) + ((x11736x) & (!x11734x) & (x11735x) & (!x11745x)) + ((x11736x) & (!x11734x) & (x11735x) & (x11745x)) + ((x11736x) & (x11734x) & (!x11735x) & (!x11745x)) + ((x11736x) & (x11734x) & (!x11735x) & (x11745x)) + ((x11736x) & (x11734x) & (x11735x) & (!x11745x)) + ((x11736x) & (x11734x) & (x11735x) & (x11745x)));
	assign n_n1083 = (((!n_n4800) & (!x11757x) & (!n_n4798) & (x439x)) + ((!n_n4800) & (!x11757x) & (n_n4798) & (!x439x)) + ((!n_n4800) & (!x11757x) & (n_n4798) & (x439x)) + ((!n_n4800) & (x11757x) & (!n_n4798) & (!x439x)) + ((!n_n4800) & (x11757x) & (!n_n4798) & (x439x)) + ((!n_n4800) & (x11757x) & (n_n4798) & (!x439x)) + ((!n_n4800) & (x11757x) & (n_n4798) & (x439x)) + ((n_n4800) & (!x11757x) & (!n_n4798) & (!x439x)) + ((n_n4800) & (!x11757x) & (!n_n4798) & (x439x)) + ((n_n4800) & (!x11757x) & (n_n4798) & (!x439x)) + ((n_n4800) & (!x11757x) & (n_n4798) & (x439x)) + ((n_n4800) & (x11757x) & (!n_n4798) & (!x439x)) + ((n_n4800) & (x11757x) & (!n_n4798) & (x439x)) + ((n_n4800) & (x11757x) & (n_n4798) & (!x439x)) + ((n_n4800) & (x11757x) & (n_n4798) & (x439x)));
	assign n_n1082 = (((!x24x) & (!x530x) & (!n_n4812) & (!x11762x) & (x151x)) + ((!x24x) & (!x530x) & (!n_n4812) & (x11762x) & (!x151x)) + ((!x24x) & (!x530x) & (!n_n4812) & (x11762x) & (x151x)) + ((!x24x) & (!x530x) & (n_n4812) & (!x11762x) & (!x151x)) + ((!x24x) & (!x530x) & (n_n4812) & (!x11762x) & (x151x)) + ((!x24x) & (!x530x) & (n_n4812) & (x11762x) & (!x151x)) + ((!x24x) & (!x530x) & (n_n4812) & (x11762x) & (x151x)) + ((!x24x) & (x530x) & (!n_n4812) & (!x11762x) & (x151x)) + ((!x24x) & (x530x) & (!n_n4812) & (x11762x) & (!x151x)) + ((!x24x) & (x530x) & (!n_n4812) & (x11762x) & (x151x)) + ((!x24x) & (x530x) & (n_n4812) & (!x11762x) & (!x151x)) + ((!x24x) & (x530x) & (n_n4812) & (!x11762x) & (x151x)) + ((!x24x) & (x530x) & (n_n4812) & (x11762x) & (!x151x)) + ((!x24x) & (x530x) & (n_n4812) & (x11762x) & (x151x)) + ((x24x) & (!x530x) & (!n_n4812) & (!x11762x) & (x151x)) + ((x24x) & (!x530x) & (!n_n4812) & (x11762x) & (!x151x)) + ((x24x) & (!x530x) & (!n_n4812) & (x11762x) & (x151x)) + ((x24x) & (!x530x) & (n_n4812) & (!x11762x) & (!x151x)) + ((x24x) & (!x530x) & (n_n4812) & (!x11762x) & (x151x)) + ((x24x) & (!x530x) & (n_n4812) & (x11762x) & (!x151x)) + ((x24x) & (!x530x) & (n_n4812) & (x11762x) & (x151x)) + ((x24x) & (x530x) & (!n_n4812) & (!x11762x) & (!x151x)) + ((x24x) & (x530x) & (!n_n4812) & (!x11762x) & (x151x)) + ((x24x) & (x530x) & (!n_n4812) & (x11762x) & (!x151x)) + ((x24x) & (x530x) & (!n_n4812) & (x11762x) & (x151x)) + ((x24x) & (x530x) & (n_n4812) & (!x11762x) & (!x151x)) + ((x24x) & (x530x) & (n_n4812) & (!x11762x) & (x151x)) + ((x24x) & (x530x) & (n_n4812) & (x11762x) & (!x151x)) + ((x24x) & (x530x) & (n_n4812) & (x11762x) & (x151x)));
	assign x11766x = (((!n_n4787) & (!x313x) & (!n_n4792) & (!n_n2003) & (x292x)) + ((!n_n4787) & (!x313x) & (!n_n4792) & (n_n2003) & (!x292x)) + ((!n_n4787) & (!x313x) & (!n_n4792) & (n_n2003) & (x292x)) + ((!n_n4787) & (!x313x) & (n_n4792) & (!n_n2003) & (!x292x)) + ((!n_n4787) & (!x313x) & (n_n4792) & (!n_n2003) & (x292x)) + ((!n_n4787) & (!x313x) & (n_n4792) & (n_n2003) & (!x292x)) + ((!n_n4787) & (!x313x) & (n_n4792) & (n_n2003) & (x292x)) + ((!n_n4787) & (x313x) & (!n_n4792) & (!n_n2003) & (!x292x)) + ((!n_n4787) & (x313x) & (!n_n4792) & (!n_n2003) & (x292x)) + ((!n_n4787) & (x313x) & (!n_n4792) & (n_n2003) & (!x292x)) + ((!n_n4787) & (x313x) & (!n_n4792) & (n_n2003) & (x292x)) + ((!n_n4787) & (x313x) & (n_n4792) & (!n_n2003) & (!x292x)) + ((!n_n4787) & (x313x) & (n_n4792) & (!n_n2003) & (x292x)) + ((!n_n4787) & (x313x) & (n_n4792) & (n_n2003) & (!x292x)) + ((!n_n4787) & (x313x) & (n_n4792) & (n_n2003) & (x292x)) + ((n_n4787) & (!x313x) & (!n_n4792) & (!n_n2003) & (!x292x)) + ((n_n4787) & (!x313x) & (!n_n4792) & (!n_n2003) & (x292x)) + ((n_n4787) & (!x313x) & (!n_n4792) & (n_n2003) & (!x292x)) + ((n_n4787) & (!x313x) & (!n_n4792) & (n_n2003) & (x292x)) + ((n_n4787) & (!x313x) & (n_n4792) & (!n_n2003) & (!x292x)) + ((n_n4787) & (!x313x) & (n_n4792) & (!n_n2003) & (x292x)) + ((n_n4787) & (!x313x) & (n_n4792) & (n_n2003) & (!x292x)) + ((n_n4787) & (!x313x) & (n_n4792) & (n_n2003) & (x292x)) + ((n_n4787) & (x313x) & (!n_n4792) & (!n_n2003) & (!x292x)) + ((n_n4787) & (x313x) & (!n_n4792) & (!n_n2003) & (x292x)) + ((n_n4787) & (x313x) & (!n_n4792) & (n_n2003) & (!x292x)) + ((n_n4787) & (x313x) & (!n_n4792) & (n_n2003) & (x292x)) + ((n_n4787) & (x313x) & (n_n4792) & (!n_n2003) & (!x292x)) + ((n_n4787) & (x313x) & (n_n4792) & (!n_n2003) & (x292x)) + ((n_n4787) & (x313x) & (n_n4792) & (n_n2003) & (!x292x)) + ((n_n4787) & (x313x) & (n_n4792) & (n_n2003) & (x292x)));
	assign n_n1028 = (((!n_n3460) & (!x177x) & (!n_n4838) & (!x11782x) & (x11778x)) + ((!n_n3460) & (!x177x) & (!n_n4838) & (x11782x) & (!x11778x)) + ((!n_n3460) & (!x177x) & (!n_n4838) & (x11782x) & (x11778x)) + ((!n_n3460) & (!x177x) & (n_n4838) & (!x11782x) & (!x11778x)) + ((!n_n3460) & (!x177x) & (n_n4838) & (!x11782x) & (x11778x)) + ((!n_n3460) & (!x177x) & (n_n4838) & (x11782x) & (!x11778x)) + ((!n_n3460) & (!x177x) & (n_n4838) & (x11782x) & (x11778x)) + ((!n_n3460) & (x177x) & (!n_n4838) & (!x11782x) & (!x11778x)) + ((!n_n3460) & (x177x) & (!n_n4838) & (!x11782x) & (x11778x)) + ((!n_n3460) & (x177x) & (!n_n4838) & (x11782x) & (!x11778x)) + ((!n_n3460) & (x177x) & (!n_n4838) & (x11782x) & (x11778x)) + ((!n_n3460) & (x177x) & (n_n4838) & (!x11782x) & (!x11778x)) + ((!n_n3460) & (x177x) & (n_n4838) & (!x11782x) & (x11778x)) + ((!n_n3460) & (x177x) & (n_n4838) & (x11782x) & (!x11778x)) + ((!n_n3460) & (x177x) & (n_n4838) & (x11782x) & (x11778x)) + ((n_n3460) & (!x177x) & (!n_n4838) & (!x11782x) & (!x11778x)) + ((n_n3460) & (!x177x) & (!n_n4838) & (!x11782x) & (x11778x)) + ((n_n3460) & (!x177x) & (!n_n4838) & (x11782x) & (!x11778x)) + ((n_n3460) & (!x177x) & (!n_n4838) & (x11782x) & (x11778x)) + ((n_n3460) & (!x177x) & (n_n4838) & (!x11782x) & (!x11778x)) + ((n_n3460) & (!x177x) & (n_n4838) & (!x11782x) & (x11778x)) + ((n_n3460) & (!x177x) & (n_n4838) & (x11782x) & (!x11778x)) + ((n_n3460) & (!x177x) & (n_n4838) & (x11782x) & (x11778x)) + ((n_n3460) & (x177x) & (!n_n4838) & (!x11782x) & (!x11778x)) + ((n_n3460) & (x177x) & (!n_n4838) & (!x11782x) & (x11778x)) + ((n_n3460) & (x177x) & (!n_n4838) & (x11782x) & (!x11778x)) + ((n_n3460) & (x177x) & (!n_n4838) & (x11782x) & (x11778x)) + ((n_n3460) & (x177x) & (n_n4838) & (!x11782x) & (!x11778x)) + ((n_n3460) & (x177x) & (n_n4838) & (!x11782x) & (x11778x)) + ((n_n3460) & (x177x) & (n_n4838) & (x11782x) & (!x11778x)) + ((n_n3460) & (x177x) & (n_n4838) & (x11782x) & (x11778x)));
	assign x11892x = (((!n_n1086) & (!n_n1087) & (!x315x) & (!x191x) & (x11889x)) + ((!n_n1086) & (!n_n1087) & (!x315x) & (x191x) & (!x11889x)) + ((!n_n1086) & (!n_n1087) & (!x315x) & (x191x) & (x11889x)) + ((!n_n1086) & (!n_n1087) & (x315x) & (!x191x) & (!x11889x)) + ((!n_n1086) & (!n_n1087) & (x315x) & (!x191x) & (x11889x)) + ((!n_n1086) & (!n_n1087) & (x315x) & (x191x) & (!x11889x)) + ((!n_n1086) & (!n_n1087) & (x315x) & (x191x) & (x11889x)) + ((!n_n1086) & (n_n1087) & (!x315x) & (!x191x) & (!x11889x)) + ((!n_n1086) & (n_n1087) & (!x315x) & (!x191x) & (x11889x)) + ((!n_n1086) & (n_n1087) & (!x315x) & (x191x) & (!x11889x)) + ((!n_n1086) & (n_n1087) & (!x315x) & (x191x) & (x11889x)) + ((!n_n1086) & (n_n1087) & (x315x) & (!x191x) & (!x11889x)) + ((!n_n1086) & (n_n1087) & (x315x) & (!x191x) & (x11889x)) + ((!n_n1086) & (n_n1087) & (x315x) & (x191x) & (!x11889x)) + ((!n_n1086) & (n_n1087) & (x315x) & (x191x) & (x11889x)) + ((n_n1086) & (!n_n1087) & (!x315x) & (!x191x) & (!x11889x)) + ((n_n1086) & (!n_n1087) & (!x315x) & (!x191x) & (x11889x)) + ((n_n1086) & (!n_n1087) & (!x315x) & (x191x) & (!x11889x)) + ((n_n1086) & (!n_n1087) & (!x315x) & (x191x) & (x11889x)) + ((n_n1086) & (!n_n1087) & (x315x) & (!x191x) & (!x11889x)) + ((n_n1086) & (!n_n1087) & (x315x) & (!x191x) & (x11889x)) + ((n_n1086) & (!n_n1087) & (x315x) & (x191x) & (!x11889x)) + ((n_n1086) & (!n_n1087) & (x315x) & (x191x) & (x11889x)) + ((n_n1086) & (n_n1087) & (!x315x) & (!x191x) & (!x11889x)) + ((n_n1086) & (n_n1087) & (!x315x) & (!x191x) & (x11889x)) + ((n_n1086) & (n_n1087) & (!x315x) & (x191x) & (!x11889x)) + ((n_n1086) & (n_n1087) & (!x315x) & (x191x) & (x11889x)) + ((n_n1086) & (n_n1087) & (x315x) & (!x191x) & (!x11889x)) + ((n_n1086) & (n_n1087) & (x315x) & (!x191x) & (x11889x)) + ((n_n1086) & (n_n1087) & (x315x) & (x191x) & (!x11889x)) + ((n_n1086) & (n_n1087) & (x315x) & (x191x) & (x11889x)));
	assign n_n1020 = (((!n_n1057) & (!x11908x) & (x11907x)) + ((!n_n1057) & (x11908x) & (!x11907x)) + ((!n_n1057) & (x11908x) & (x11907x)) + ((n_n1057) & (!x11908x) & (!x11907x)) + ((n_n1057) & (!x11908x) & (x11907x)) + ((n_n1057) & (x11908x) & (!x11907x)) + ((n_n1057) & (x11908x) & (x11907x)));
	assign n_n1052 = (((!n_n5223) & (!n_n5221) & (!n_n5215) & (!x181x) & (!x22157x)) + ((!n_n5223) & (!n_n5221) & (!n_n5215) & (x181x) & (!x22157x)) + ((!n_n5223) & (!n_n5221) & (!n_n5215) & (x181x) & (x22157x)) + ((!n_n5223) & (!n_n5221) & (n_n5215) & (!x181x) & (!x22157x)) + ((!n_n5223) & (!n_n5221) & (n_n5215) & (!x181x) & (x22157x)) + ((!n_n5223) & (!n_n5221) & (n_n5215) & (x181x) & (!x22157x)) + ((!n_n5223) & (!n_n5221) & (n_n5215) & (x181x) & (x22157x)) + ((!n_n5223) & (n_n5221) & (!n_n5215) & (!x181x) & (!x22157x)) + ((!n_n5223) & (n_n5221) & (!n_n5215) & (!x181x) & (x22157x)) + ((!n_n5223) & (n_n5221) & (!n_n5215) & (x181x) & (!x22157x)) + ((!n_n5223) & (n_n5221) & (!n_n5215) & (x181x) & (x22157x)) + ((!n_n5223) & (n_n5221) & (n_n5215) & (!x181x) & (!x22157x)) + ((!n_n5223) & (n_n5221) & (n_n5215) & (!x181x) & (x22157x)) + ((!n_n5223) & (n_n5221) & (n_n5215) & (x181x) & (!x22157x)) + ((!n_n5223) & (n_n5221) & (n_n5215) & (x181x) & (x22157x)) + ((n_n5223) & (!n_n5221) & (!n_n5215) & (!x181x) & (!x22157x)) + ((n_n5223) & (!n_n5221) & (!n_n5215) & (!x181x) & (x22157x)) + ((n_n5223) & (!n_n5221) & (!n_n5215) & (x181x) & (!x22157x)) + ((n_n5223) & (!n_n5221) & (!n_n5215) & (x181x) & (x22157x)) + ((n_n5223) & (!n_n5221) & (n_n5215) & (!x181x) & (!x22157x)) + ((n_n5223) & (!n_n5221) & (n_n5215) & (!x181x) & (x22157x)) + ((n_n5223) & (!n_n5221) & (n_n5215) & (x181x) & (!x22157x)) + ((n_n5223) & (!n_n5221) & (n_n5215) & (x181x) & (x22157x)) + ((n_n5223) & (n_n5221) & (!n_n5215) & (!x181x) & (!x22157x)) + ((n_n5223) & (n_n5221) & (!n_n5215) & (!x181x) & (x22157x)) + ((n_n5223) & (n_n5221) & (!n_n5215) & (x181x) & (!x22157x)) + ((n_n5223) & (n_n5221) & (!n_n5215) & (x181x) & (x22157x)) + ((n_n5223) & (n_n5221) & (n_n5215) & (!x181x) & (!x22157x)) + ((n_n5223) & (n_n5221) & (n_n5215) & (!x181x) & (x22157x)) + ((n_n5223) & (n_n5221) & (n_n5215) & (x181x) & (!x22157x)) + ((n_n5223) & (n_n5221) & (n_n5215) & (x181x) & (x22157x)));
	assign n_n1054 = (((!n_n5200) & (!n_n5188) & (!n_n1927) & (!x188x) & (x452x)) + ((!n_n5200) & (!n_n5188) & (!n_n1927) & (x188x) & (!x452x)) + ((!n_n5200) & (!n_n5188) & (!n_n1927) & (x188x) & (x452x)) + ((!n_n5200) & (!n_n5188) & (n_n1927) & (!x188x) & (!x452x)) + ((!n_n5200) & (!n_n5188) & (n_n1927) & (!x188x) & (x452x)) + ((!n_n5200) & (!n_n5188) & (n_n1927) & (x188x) & (!x452x)) + ((!n_n5200) & (!n_n5188) & (n_n1927) & (x188x) & (x452x)) + ((!n_n5200) & (n_n5188) & (!n_n1927) & (!x188x) & (!x452x)) + ((!n_n5200) & (n_n5188) & (!n_n1927) & (!x188x) & (x452x)) + ((!n_n5200) & (n_n5188) & (!n_n1927) & (x188x) & (!x452x)) + ((!n_n5200) & (n_n5188) & (!n_n1927) & (x188x) & (x452x)) + ((!n_n5200) & (n_n5188) & (n_n1927) & (!x188x) & (!x452x)) + ((!n_n5200) & (n_n5188) & (n_n1927) & (!x188x) & (x452x)) + ((!n_n5200) & (n_n5188) & (n_n1927) & (x188x) & (!x452x)) + ((!n_n5200) & (n_n5188) & (n_n1927) & (x188x) & (x452x)) + ((n_n5200) & (!n_n5188) & (!n_n1927) & (!x188x) & (!x452x)) + ((n_n5200) & (!n_n5188) & (!n_n1927) & (!x188x) & (x452x)) + ((n_n5200) & (!n_n5188) & (!n_n1927) & (x188x) & (!x452x)) + ((n_n5200) & (!n_n5188) & (!n_n1927) & (x188x) & (x452x)) + ((n_n5200) & (!n_n5188) & (n_n1927) & (!x188x) & (!x452x)) + ((n_n5200) & (!n_n5188) & (n_n1927) & (!x188x) & (x452x)) + ((n_n5200) & (!n_n5188) & (n_n1927) & (x188x) & (!x452x)) + ((n_n5200) & (!n_n5188) & (n_n1927) & (x188x) & (x452x)) + ((n_n5200) & (n_n5188) & (!n_n1927) & (!x188x) & (!x452x)) + ((n_n5200) & (n_n5188) & (!n_n1927) & (!x188x) & (x452x)) + ((n_n5200) & (n_n5188) & (!n_n1927) & (x188x) & (!x452x)) + ((n_n5200) & (n_n5188) & (!n_n1927) & (x188x) & (x452x)) + ((n_n5200) & (n_n5188) & (n_n1927) & (!x188x) & (!x452x)) + ((n_n5200) & (n_n5188) & (n_n1927) & (!x188x) & (x452x)) + ((n_n5200) & (n_n5188) & (n_n1927) & (x188x) & (!x452x)) + ((n_n5200) & (n_n5188) & (n_n1927) & (x188x) & (x452x)));
	assign x11977x = (((!n_n5207) & (!n_n5203) & (!x36x) & (x11976x)) + ((!n_n5207) & (!n_n5203) & (x36x) & (!x11976x)) + ((!n_n5207) & (!n_n5203) & (x36x) & (x11976x)) + ((!n_n5207) & (n_n5203) & (!x36x) & (!x11976x)) + ((!n_n5207) & (n_n5203) & (!x36x) & (x11976x)) + ((!n_n5207) & (n_n5203) & (x36x) & (!x11976x)) + ((!n_n5207) & (n_n5203) & (x36x) & (x11976x)) + ((n_n5207) & (!n_n5203) & (!x36x) & (!x11976x)) + ((n_n5207) & (!n_n5203) & (!x36x) & (x11976x)) + ((n_n5207) & (!n_n5203) & (x36x) & (!x11976x)) + ((n_n5207) & (!n_n5203) & (x36x) & (x11976x)) + ((n_n5207) & (n_n5203) & (!x36x) & (!x11976x)) + ((n_n5207) & (n_n5203) & (!x36x) & (x11976x)) + ((n_n5207) & (n_n5203) & (x36x) & (!x11976x)) + ((n_n5207) & (n_n5203) & (x36x) & (x11976x)));
	assign x12036x = (((!n_n1059) & (!n_n1060) & (!x211x) & (!x422x) & (x12033x)) + ((!n_n1059) & (!n_n1060) & (!x211x) & (x422x) & (!x12033x)) + ((!n_n1059) & (!n_n1060) & (!x211x) & (x422x) & (x12033x)) + ((!n_n1059) & (!n_n1060) & (x211x) & (!x422x) & (!x12033x)) + ((!n_n1059) & (!n_n1060) & (x211x) & (!x422x) & (x12033x)) + ((!n_n1059) & (!n_n1060) & (x211x) & (x422x) & (!x12033x)) + ((!n_n1059) & (!n_n1060) & (x211x) & (x422x) & (x12033x)) + ((!n_n1059) & (n_n1060) & (!x211x) & (!x422x) & (!x12033x)) + ((!n_n1059) & (n_n1060) & (!x211x) & (!x422x) & (x12033x)) + ((!n_n1059) & (n_n1060) & (!x211x) & (x422x) & (!x12033x)) + ((!n_n1059) & (n_n1060) & (!x211x) & (x422x) & (x12033x)) + ((!n_n1059) & (n_n1060) & (x211x) & (!x422x) & (!x12033x)) + ((!n_n1059) & (n_n1060) & (x211x) & (!x422x) & (x12033x)) + ((!n_n1059) & (n_n1060) & (x211x) & (x422x) & (!x12033x)) + ((!n_n1059) & (n_n1060) & (x211x) & (x422x) & (x12033x)) + ((n_n1059) & (!n_n1060) & (!x211x) & (!x422x) & (!x12033x)) + ((n_n1059) & (!n_n1060) & (!x211x) & (!x422x) & (x12033x)) + ((n_n1059) & (!n_n1060) & (!x211x) & (x422x) & (!x12033x)) + ((n_n1059) & (!n_n1060) & (!x211x) & (x422x) & (x12033x)) + ((n_n1059) & (!n_n1060) & (x211x) & (!x422x) & (!x12033x)) + ((n_n1059) & (!n_n1060) & (x211x) & (!x422x) & (x12033x)) + ((n_n1059) & (!n_n1060) & (x211x) & (x422x) & (!x12033x)) + ((n_n1059) & (!n_n1060) & (x211x) & (x422x) & (x12033x)) + ((n_n1059) & (n_n1060) & (!x211x) & (!x422x) & (!x12033x)) + ((n_n1059) & (n_n1060) & (!x211x) & (!x422x) & (x12033x)) + ((n_n1059) & (n_n1060) & (!x211x) & (x422x) & (!x12033x)) + ((n_n1059) & (n_n1060) & (!x211x) & (x422x) & (x12033x)) + ((n_n1059) & (n_n1060) & (x211x) & (!x422x) & (!x12033x)) + ((n_n1059) & (n_n1060) & (x211x) & (!x422x) & (x12033x)) + ((n_n1059) & (n_n1060) & (x211x) & (x422x) & (!x12033x)) + ((n_n1059) & (n_n1060) & (x211x) & (x422x) & (x12033x)));
	assign x12062x = (((!n_n4506) & (!n_n4546) & (!n_n4555) & (!n_n4562) & (x12061x)) + ((!n_n4506) & (!n_n4546) & (!n_n4555) & (n_n4562) & (!x12061x)) + ((!n_n4506) & (!n_n4546) & (!n_n4555) & (n_n4562) & (x12061x)) + ((!n_n4506) & (!n_n4546) & (n_n4555) & (!n_n4562) & (!x12061x)) + ((!n_n4506) & (!n_n4546) & (n_n4555) & (!n_n4562) & (x12061x)) + ((!n_n4506) & (!n_n4546) & (n_n4555) & (n_n4562) & (!x12061x)) + ((!n_n4506) & (!n_n4546) & (n_n4555) & (n_n4562) & (x12061x)) + ((!n_n4506) & (n_n4546) & (!n_n4555) & (!n_n4562) & (!x12061x)) + ((!n_n4506) & (n_n4546) & (!n_n4555) & (!n_n4562) & (x12061x)) + ((!n_n4506) & (n_n4546) & (!n_n4555) & (n_n4562) & (!x12061x)) + ((!n_n4506) & (n_n4546) & (!n_n4555) & (n_n4562) & (x12061x)) + ((!n_n4506) & (n_n4546) & (n_n4555) & (!n_n4562) & (!x12061x)) + ((!n_n4506) & (n_n4546) & (n_n4555) & (!n_n4562) & (x12061x)) + ((!n_n4506) & (n_n4546) & (n_n4555) & (n_n4562) & (!x12061x)) + ((!n_n4506) & (n_n4546) & (n_n4555) & (n_n4562) & (x12061x)) + ((n_n4506) & (!n_n4546) & (!n_n4555) & (!n_n4562) & (!x12061x)) + ((n_n4506) & (!n_n4546) & (!n_n4555) & (!n_n4562) & (x12061x)) + ((n_n4506) & (!n_n4546) & (!n_n4555) & (n_n4562) & (!x12061x)) + ((n_n4506) & (!n_n4546) & (!n_n4555) & (n_n4562) & (x12061x)) + ((n_n4506) & (!n_n4546) & (n_n4555) & (!n_n4562) & (!x12061x)) + ((n_n4506) & (!n_n4546) & (n_n4555) & (!n_n4562) & (x12061x)) + ((n_n4506) & (!n_n4546) & (n_n4555) & (n_n4562) & (!x12061x)) + ((n_n4506) & (!n_n4546) & (n_n4555) & (n_n4562) & (x12061x)) + ((n_n4506) & (n_n4546) & (!n_n4555) & (!n_n4562) & (!x12061x)) + ((n_n4506) & (n_n4546) & (!n_n4555) & (!n_n4562) & (x12061x)) + ((n_n4506) & (n_n4546) & (!n_n4555) & (n_n4562) & (!x12061x)) + ((n_n4506) & (n_n4546) & (!n_n4555) & (n_n4562) & (x12061x)) + ((n_n4506) & (n_n4546) & (n_n4555) & (!n_n4562) & (!x12061x)) + ((n_n4506) & (n_n4546) & (n_n4555) & (!n_n4562) & (x12061x)) + ((n_n4506) & (n_n4546) & (n_n4555) & (n_n4562) & (!x12061x)) + ((n_n4506) & (n_n4546) & (n_n4555) & (n_n4562) & (x12061x)));
	assign x12063x = (((!x12048x) & (!x12049x) & (!x12053x) & (x12054x)) + ((!x12048x) & (!x12049x) & (x12053x) & (!x12054x)) + ((!x12048x) & (!x12049x) & (x12053x) & (x12054x)) + ((!x12048x) & (x12049x) & (!x12053x) & (!x12054x)) + ((!x12048x) & (x12049x) & (!x12053x) & (x12054x)) + ((!x12048x) & (x12049x) & (x12053x) & (!x12054x)) + ((!x12048x) & (x12049x) & (x12053x) & (x12054x)) + ((x12048x) & (!x12049x) & (!x12053x) & (!x12054x)) + ((x12048x) & (!x12049x) & (!x12053x) & (x12054x)) + ((x12048x) & (!x12049x) & (x12053x) & (!x12054x)) + ((x12048x) & (!x12049x) & (x12053x) & (x12054x)) + ((x12048x) & (x12049x) & (!x12053x) & (!x12054x)) + ((x12048x) & (x12049x) & (!x12053x) & (x12054x)) + ((x12048x) & (x12049x) & (x12053x) & (!x12054x)) + ((x12048x) & (x12049x) & (x12053x) & (x12054x)));
	assign x12083x = (((!n_n4774) & (!n_n4845) & (!n_n4796) & (!n_n4822) & (x12082x)) + ((!n_n4774) & (!n_n4845) & (!n_n4796) & (n_n4822) & (!x12082x)) + ((!n_n4774) & (!n_n4845) & (!n_n4796) & (n_n4822) & (x12082x)) + ((!n_n4774) & (!n_n4845) & (n_n4796) & (!n_n4822) & (!x12082x)) + ((!n_n4774) & (!n_n4845) & (n_n4796) & (!n_n4822) & (x12082x)) + ((!n_n4774) & (!n_n4845) & (n_n4796) & (n_n4822) & (!x12082x)) + ((!n_n4774) & (!n_n4845) & (n_n4796) & (n_n4822) & (x12082x)) + ((!n_n4774) & (n_n4845) & (!n_n4796) & (!n_n4822) & (!x12082x)) + ((!n_n4774) & (n_n4845) & (!n_n4796) & (!n_n4822) & (x12082x)) + ((!n_n4774) & (n_n4845) & (!n_n4796) & (n_n4822) & (!x12082x)) + ((!n_n4774) & (n_n4845) & (!n_n4796) & (n_n4822) & (x12082x)) + ((!n_n4774) & (n_n4845) & (n_n4796) & (!n_n4822) & (!x12082x)) + ((!n_n4774) & (n_n4845) & (n_n4796) & (!n_n4822) & (x12082x)) + ((!n_n4774) & (n_n4845) & (n_n4796) & (n_n4822) & (!x12082x)) + ((!n_n4774) & (n_n4845) & (n_n4796) & (n_n4822) & (x12082x)) + ((n_n4774) & (!n_n4845) & (!n_n4796) & (!n_n4822) & (!x12082x)) + ((n_n4774) & (!n_n4845) & (!n_n4796) & (!n_n4822) & (x12082x)) + ((n_n4774) & (!n_n4845) & (!n_n4796) & (n_n4822) & (!x12082x)) + ((n_n4774) & (!n_n4845) & (!n_n4796) & (n_n4822) & (x12082x)) + ((n_n4774) & (!n_n4845) & (n_n4796) & (!n_n4822) & (!x12082x)) + ((n_n4774) & (!n_n4845) & (n_n4796) & (!n_n4822) & (x12082x)) + ((n_n4774) & (!n_n4845) & (n_n4796) & (n_n4822) & (!x12082x)) + ((n_n4774) & (!n_n4845) & (n_n4796) & (n_n4822) & (x12082x)) + ((n_n4774) & (n_n4845) & (!n_n4796) & (!n_n4822) & (!x12082x)) + ((n_n4774) & (n_n4845) & (!n_n4796) & (!n_n4822) & (x12082x)) + ((n_n4774) & (n_n4845) & (!n_n4796) & (n_n4822) & (!x12082x)) + ((n_n4774) & (n_n4845) & (!n_n4796) & (n_n4822) & (x12082x)) + ((n_n4774) & (n_n4845) & (n_n4796) & (!n_n4822) & (!x12082x)) + ((n_n4774) & (n_n4845) & (n_n4796) & (!n_n4822) & (x12082x)) + ((n_n4774) & (n_n4845) & (n_n4796) & (n_n4822) & (!x12082x)) + ((n_n4774) & (n_n4845) & (n_n4796) & (n_n4822) & (x12082x)));
	assign x12084x = (((!x12068x) & (!x12069x) & (!x12074x) & (x12075x)) + ((!x12068x) & (!x12069x) & (x12074x) & (!x12075x)) + ((!x12068x) & (!x12069x) & (x12074x) & (x12075x)) + ((!x12068x) & (x12069x) & (!x12074x) & (!x12075x)) + ((!x12068x) & (x12069x) & (!x12074x) & (x12075x)) + ((!x12068x) & (x12069x) & (x12074x) & (!x12075x)) + ((!x12068x) & (x12069x) & (x12074x) & (x12075x)) + ((x12068x) & (!x12069x) & (!x12074x) & (!x12075x)) + ((x12068x) & (!x12069x) & (!x12074x) & (x12075x)) + ((x12068x) & (!x12069x) & (x12074x) & (!x12075x)) + ((x12068x) & (!x12069x) & (x12074x) & (x12075x)) + ((x12068x) & (x12069x) & (!x12074x) & (!x12075x)) + ((x12068x) & (x12069x) & (!x12074x) & (x12075x)) + ((x12068x) & (x12069x) & (x12074x) & (!x12075x)) + ((x12068x) & (x12069x) & (x12074x) & (x12075x)));
	assign n_n1323 = (((!n_n1330) & (!n_n1331) & (x12110x)) + ((!n_n1330) & (n_n1331) & (!x12110x)) + ((!n_n1330) & (n_n1331) & (x12110x)) + ((n_n1330) & (!n_n1331) & (!x12110x)) + ((n_n1330) & (!n_n1331) & (x12110x)) + ((n_n1330) & (n_n1331) & (!x12110x)) + ((n_n1330) & (n_n1331) & (x12110x)));
	assign x12129x = (((!x12089x) & (!x12090x) & (x12128x)) + ((!x12089x) & (x12090x) & (!x12128x)) + ((!x12089x) & (x12090x) & (x12128x)) + ((x12089x) & (!x12090x) & (!x12128x)) + ((x12089x) & (!x12090x) & (x12128x)) + ((x12089x) & (x12090x) & (!x12128x)) + ((x12089x) & (x12090x) & (x12128x)));
	assign x12130x = (((!x12117x) & (!x12118x) & (n_n1333)) + ((!x12117x) & (x12118x) & (!n_n1333)) + ((!x12117x) & (x12118x) & (n_n1333)) + ((x12117x) & (!x12118x) & (!n_n1333)) + ((x12117x) & (!x12118x) & (n_n1333)) + ((x12117x) & (x12118x) & (!n_n1333)) + ((x12117x) & (x12118x) & (n_n1333)));
	assign x12150x = (((!n_n1341) & (!x12141x) & (!x12142x) & (!x12146x) & (x12147x)) + ((!n_n1341) & (!x12141x) & (!x12142x) & (x12146x) & (!x12147x)) + ((!n_n1341) & (!x12141x) & (!x12142x) & (x12146x) & (x12147x)) + ((!n_n1341) & (!x12141x) & (x12142x) & (!x12146x) & (!x12147x)) + ((!n_n1341) & (!x12141x) & (x12142x) & (!x12146x) & (x12147x)) + ((!n_n1341) & (!x12141x) & (x12142x) & (x12146x) & (!x12147x)) + ((!n_n1341) & (!x12141x) & (x12142x) & (x12146x) & (x12147x)) + ((!n_n1341) & (x12141x) & (!x12142x) & (!x12146x) & (!x12147x)) + ((!n_n1341) & (x12141x) & (!x12142x) & (!x12146x) & (x12147x)) + ((!n_n1341) & (x12141x) & (!x12142x) & (x12146x) & (!x12147x)) + ((!n_n1341) & (x12141x) & (!x12142x) & (x12146x) & (x12147x)) + ((!n_n1341) & (x12141x) & (x12142x) & (!x12146x) & (!x12147x)) + ((!n_n1341) & (x12141x) & (x12142x) & (!x12146x) & (x12147x)) + ((!n_n1341) & (x12141x) & (x12142x) & (x12146x) & (!x12147x)) + ((!n_n1341) & (x12141x) & (x12142x) & (x12146x) & (x12147x)) + ((n_n1341) & (!x12141x) & (!x12142x) & (!x12146x) & (!x12147x)) + ((n_n1341) & (!x12141x) & (!x12142x) & (!x12146x) & (x12147x)) + ((n_n1341) & (!x12141x) & (!x12142x) & (x12146x) & (!x12147x)) + ((n_n1341) & (!x12141x) & (!x12142x) & (x12146x) & (x12147x)) + ((n_n1341) & (!x12141x) & (x12142x) & (!x12146x) & (!x12147x)) + ((n_n1341) & (!x12141x) & (x12142x) & (!x12146x) & (x12147x)) + ((n_n1341) & (!x12141x) & (x12142x) & (x12146x) & (!x12147x)) + ((n_n1341) & (!x12141x) & (x12142x) & (x12146x) & (x12147x)) + ((n_n1341) & (x12141x) & (!x12142x) & (!x12146x) & (!x12147x)) + ((n_n1341) & (x12141x) & (!x12142x) & (!x12146x) & (x12147x)) + ((n_n1341) & (x12141x) & (!x12142x) & (x12146x) & (!x12147x)) + ((n_n1341) & (x12141x) & (!x12142x) & (x12146x) & (x12147x)) + ((n_n1341) & (x12141x) & (x12142x) & (!x12146x) & (!x12147x)) + ((n_n1341) & (x12141x) & (x12142x) & (!x12146x) & (x12147x)) + ((n_n1341) & (x12141x) & (x12142x) & (x12146x) & (!x12147x)) + ((n_n1341) & (x12141x) & (x12142x) & (x12146x) & (x12147x)));
	assign n_n4979 = (((!i_9_) & (n_n524) & (n_n518) & (n_n195)));
	assign n_n4978 = (((i_9_) & (n_n524) & (n_n518) & (n_n195)));
	assign x12156x = (((!n_n4982) & (!n_n4988) & (!n_n4989) & (!n_n4985) & (n_n4986)) + ((!n_n4982) & (!n_n4988) & (!n_n4989) & (n_n4985) & (!n_n4986)) + ((!n_n4982) & (!n_n4988) & (!n_n4989) & (n_n4985) & (n_n4986)) + ((!n_n4982) & (!n_n4988) & (n_n4989) & (!n_n4985) & (!n_n4986)) + ((!n_n4982) & (!n_n4988) & (n_n4989) & (!n_n4985) & (n_n4986)) + ((!n_n4982) & (!n_n4988) & (n_n4989) & (n_n4985) & (!n_n4986)) + ((!n_n4982) & (!n_n4988) & (n_n4989) & (n_n4985) & (n_n4986)) + ((!n_n4982) & (n_n4988) & (!n_n4989) & (!n_n4985) & (!n_n4986)) + ((!n_n4982) & (n_n4988) & (!n_n4989) & (!n_n4985) & (n_n4986)) + ((!n_n4982) & (n_n4988) & (!n_n4989) & (n_n4985) & (!n_n4986)) + ((!n_n4982) & (n_n4988) & (!n_n4989) & (n_n4985) & (n_n4986)) + ((!n_n4982) & (n_n4988) & (n_n4989) & (!n_n4985) & (!n_n4986)) + ((!n_n4982) & (n_n4988) & (n_n4989) & (!n_n4985) & (n_n4986)) + ((!n_n4982) & (n_n4988) & (n_n4989) & (n_n4985) & (!n_n4986)) + ((!n_n4982) & (n_n4988) & (n_n4989) & (n_n4985) & (n_n4986)) + ((n_n4982) & (!n_n4988) & (!n_n4989) & (!n_n4985) & (!n_n4986)) + ((n_n4982) & (!n_n4988) & (!n_n4989) & (!n_n4985) & (n_n4986)) + ((n_n4982) & (!n_n4988) & (!n_n4989) & (n_n4985) & (!n_n4986)) + ((n_n4982) & (!n_n4988) & (!n_n4989) & (n_n4985) & (n_n4986)) + ((n_n4982) & (!n_n4988) & (n_n4989) & (!n_n4985) & (!n_n4986)) + ((n_n4982) & (!n_n4988) & (n_n4989) & (!n_n4985) & (n_n4986)) + ((n_n4982) & (!n_n4988) & (n_n4989) & (n_n4985) & (!n_n4986)) + ((n_n4982) & (!n_n4988) & (n_n4989) & (n_n4985) & (n_n4986)) + ((n_n4982) & (n_n4988) & (!n_n4989) & (!n_n4985) & (!n_n4986)) + ((n_n4982) & (n_n4988) & (!n_n4989) & (!n_n4985) & (n_n4986)) + ((n_n4982) & (n_n4988) & (!n_n4989) & (n_n4985) & (!n_n4986)) + ((n_n4982) & (n_n4988) & (!n_n4989) & (n_n4985) & (n_n4986)) + ((n_n4982) & (n_n4988) & (n_n4989) & (!n_n4985) & (!n_n4986)) + ((n_n4982) & (n_n4988) & (n_n4989) & (!n_n4985) & (n_n4986)) + ((n_n4982) & (n_n4988) & (n_n4989) & (n_n4985) & (!n_n4986)) + ((n_n4982) & (n_n4988) & (n_n4989) & (n_n4985) & (n_n4986)));
	assign n_n1455 = (((!n_n4991) & (!n_n5000) & (!n_n1576) & (!x247x) & (x104x)) + ((!n_n4991) & (!n_n5000) & (!n_n1576) & (x247x) & (!x104x)) + ((!n_n4991) & (!n_n5000) & (!n_n1576) & (x247x) & (x104x)) + ((!n_n4991) & (!n_n5000) & (n_n1576) & (!x247x) & (!x104x)) + ((!n_n4991) & (!n_n5000) & (n_n1576) & (!x247x) & (x104x)) + ((!n_n4991) & (!n_n5000) & (n_n1576) & (x247x) & (!x104x)) + ((!n_n4991) & (!n_n5000) & (n_n1576) & (x247x) & (x104x)) + ((!n_n4991) & (n_n5000) & (!n_n1576) & (!x247x) & (!x104x)) + ((!n_n4991) & (n_n5000) & (!n_n1576) & (!x247x) & (x104x)) + ((!n_n4991) & (n_n5000) & (!n_n1576) & (x247x) & (!x104x)) + ((!n_n4991) & (n_n5000) & (!n_n1576) & (x247x) & (x104x)) + ((!n_n4991) & (n_n5000) & (n_n1576) & (!x247x) & (!x104x)) + ((!n_n4991) & (n_n5000) & (n_n1576) & (!x247x) & (x104x)) + ((!n_n4991) & (n_n5000) & (n_n1576) & (x247x) & (!x104x)) + ((!n_n4991) & (n_n5000) & (n_n1576) & (x247x) & (x104x)) + ((n_n4991) & (!n_n5000) & (!n_n1576) & (!x247x) & (!x104x)) + ((n_n4991) & (!n_n5000) & (!n_n1576) & (!x247x) & (x104x)) + ((n_n4991) & (!n_n5000) & (!n_n1576) & (x247x) & (!x104x)) + ((n_n4991) & (!n_n5000) & (!n_n1576) & (x247x) & (x104x)) + ((n_n4991) & (!n_n5000) & (n_n1576) & (!x247x) & (!x104x)) + ((n_n4991) & (!n_n5000) & (n_n1576) & (!x247x) & (x104x)) + ((n_n4991) & (!n_n5000) & (n_n1576) & (x247x) & (!x104x)) + ((n_n4991) & (!n_n5000) & (n_n1576) & (x247x) & (x104x)) + ((n_n4991) & (n_n5000) & (!n_n1576) & (!x247x) & (!x104x)) + ((n_n4991) & (n_n5000) & (!n_n1576) & (!x247x) & (x104x)) + ((n_n4991) & (n_n5000) & (!n_n1576) & (x247x) & (!x104x)) + ((n_n4991) & (n_n5000) & (!n_n1576) & (x247x) & (x104x)) + ((n_n4991) & (n_n5000) & (n_n1576) & (!x247x) & (!x104x)) + ((n_n4991) & (n_n5000) & (n_n1576) & (!x247x) & (x104x)) + ((n_n4991) & (n_n5000) & (n_n1576) & (x247x) & (!x104x)) + ((n_n4991) & (n_n5000) & (n_n1576) & (x247x) & (x104x)));
	assign x22195x = (((!n_n4983) & (!n_n4984) & (!x228x) & (!x362x) & (!x12196x)));
	assign x12199x = (((!n_n4979) & (!n_n4978) & (!x12156x) & (!n_n1455) & (!x22195x)) + ((!n_n4979) & (!n_n4978) & (!x12156x) & (n_n1455) & (!x22195x)) + ((!n_n4979) & (!n_n4978) & (!x12156x) & (n_n1455) & (x22195x)) + ((!n_n4979) & (!n_n4978) & (x12156x) & (!n_n1455) & (!x22195x)) + ((!n_n4979) & (!n_n4978) & (x12156x) & (!n_n1455) & (x22195x)) + ((!n_n4979) & (!n_n4978) & (x12156x) & (n_n1455) & (!x22195x)) + ((!n_n4979) & (!n_n4978) & (x12156x) & (n_n1455) & (x22195x)) + ((!n_n4979) & (n_n4978) & (!x12156x) & (!n_n1455) & (!x22195x)) + ((!n_n4979) & (n_n4978) & (!x12156x) & (!n_n1455) & (x22195x)) + ((!n_n4979) & (n_n4978) & (!x12156x) & (n_n1455) & (!x22195x)) + ((!n_n4979) & (n_n4978) & (!x12156x) & (n_n1455) & (x22195x)) + ((!n_n4979) & (n_n4978) & (x12156x) & (!n_n1455) & (!x22195x)) + ((!n_n4979) & (n_n4978) & (x12156x) & (!n_n1455) & (x22195x)) + ((!n_n4979) & (n_n4978) & (x12156x) & (n_n1455) & (!x22195x)) + ((!n_n4979) & (n_n4978) & (x12156x) & (n_n1455) & (x22195x)) + ((n_n4979) & (!n_n4978) & (!x12156x) & (!n_n1455) & (!x22195x)) + ((n_n4979) & (!n_n4978) & (!x12156x) & (!n_n1455) & (x22195x)) + ((n_n4979) & (!n_n4978) & (!x12156x) & (n_n1455) & (!x22195x)) + ((n_n4979) & (!n_n4978) & (!x12156x) & (n_n1455) & (x22195x)) + ((n_n4979) & (!n_n4978) & (x12156x) & (!n_n1455) & (!x22195x)) + ((n_n4979) & (!n_n4978) & (x12156x) & (!n_n1455) & (x22195x)) + ((n_n4979) & (!n_n4978) & (x12156x) & (n_n1455) & (!x22195x)) + ((n_n4979) & (!n_n4978) & (x12156x) & (n_n1455) & (x22195x)) + ((n_n4979) & (n_n4978) & (!x12156x) & (!n_n1455) & (!x22195x)) + ((n_n4979) & (n_n4978) & (!x12156x) & (!n_n1455) & (x22195x)) + ((n_n4979) & (n_n4978) & (!x12156x) & (n_n1455) & (!x22195x)) + ((n_n4979) & (n_n4978) & (!x12156x) & (n_n1455) & (x22195x)) + ((n_n4979) & (n_n4978) & (x12156x) & (!n_n1455) & (!x22195x)) + ((n_n4979) & (n_n4978) & (x12156x) & (!n_n1455) & (x22195x)) + ((n_n4979) & (n_n4978) & (x12156x) & (n_n1455) & (!x22195x)) + ((n_n4979) & (n_n4978) & (x12156x) & (n_n1455) & (x22195x)));
	assign n_n1412 = (((!x12164x) & (!x12165x) & (!x142x) & (x12176x)) + ((!x12164x) & (!x12165x) & (x142x) & (!x12176x)) + ((!x12164x) & (!x12165x) & (x142x) & (x12176x)) + ((!x12164x) & (x12165x) & (!x142x) & (!x12176x)) + ((!x12164x) & (x12165x) & (!x142x) & (x12176x)) + ((!x12164x) & (x12165x) & (x142x) & (!x12176x)) + ((!x12164x) & (x12165x) & (x142x) & (x12176x)) + ((x12164x) & (!x12165x) & (!x142x) & (!x12176x)) + ((x12164x) & (!x12165x) & (!x142x) & (x12176x)) + ((x12164x) & (!x12165x) & (x142x) & (!x12176x)) + ((x12164x) & (!x12165x) & (x142x) & (x12176x)) + ((x12164x) & (x12165x) & (!x142x) & (!x12176x)) + ((x12164x) & (x12165x) & (!x142x) & (x12176x)) + ((x12164x) & (x12165x) & (x142x) & (!x12176x)) + ((x12164x) & (x12165x) & (x142x) & (x12176x)));
	assign n_n1413 = (((!n_n3810) & (!n_n1592) & (!n_n1463) & (!x12188x) & (x12190x)) + ((!n_n3810) & (!n_n1592) & (!n_n1463) & (x12188x) & (!x12190x)) + ((!n_n3810) & (!n_n1592) & (!n_n1463) & (x12188x) & (x12190x)) + ((!n_n3810) & (!n_n1592) & (n_n1463) & (!x12188x) & (!x12190x)) + ((!n_n3810) & (!n_n1592) & (n_n1463) & (!x12188x) & (x12190x)) + ((!n_n3810) & (!n_n1592) & (n_n1463) & (x12188x) & (!x12190x)) + ((!n_n3810) & (!n_n1592) & (n_n1463) & (x12188x) & (x12190x)) + ((!n_n3810) & (n_n1592) & (!n_n1463) & (!x12188x) & (!x12190x)) + ((!n_n3810) & (n_n1592) & (!n_n1463) & (!x12188x) & (x12190x)) + ((!n_n3810) & (n_n1592) & (!n_n1463) & (x12188x) & (!x12190x)) + ((!n_n3810) & (n_n1592) & (!n_n1463) & (x12188x) & (x12190x)) + ((!n_n3810) & (n_n1592) & (n_n1463) & (!x12188x) & (!x12190x)) + ((!n_n3810) & (n_n1592) & (n_n1463) & (!x12188x) & (x12190x)) + ((!n_n3810) & (n_n1592) & (n_n1463) & (x12188x) & (!x12190x)) + ((!n_n3810) & (n_n1592) & (n_n1463) & (x12188x) & (x12190x)) + ((n_n3810) & (!n_n1592) & (!n_n1463) & (!x12188x) & (!x12190x)) + ((n_n3810) & (!n_n1592) & (!n_n1463) & (!x12188x) & (x12190x)) + ((n_n3810) & (!n_n1592) & (!n_n1463) & (x12188x) & (!x12190x)) + ((n_n3810) & (!n_n1592) & (!n_n1463) & (x12188x) & (x12190x)) + ((n_n3810) & (!n_n1592) & (n_n1463) & (!x12188x) & (!x12190x)) + ((n_n3810) & (!n_n1592) & (n_n1463) & (!x12188x) & (x12190x)) + ((n_n3810) & (!n_n1592) & (n_n1463) & (x12188x) & (!x12190x)) + ((n_n3810) & (!n_n1592) & (n_n1463) & (x12188x) & (x12190x)) + ((n_n3810) & (n_n1592) & (!n_n1463) & (!x12188x) & (!x12190x)) + ((n_n3810) & (n_n1592) & (!n_n1463) & (!x12188x) & (x12190x)) + ((n_n3810) & (n_n1592) & (!n_n1463) & (x12188x) & (!x12190x)) + ((n_n3810) & (n_n1592) & (!n_n1463) & (x12188x) & (x12190x)) + ((n_n3810) & (n_n1592) & (n_n1463) & (!x12188x) & (!x12190x)) + ((n_n3810) & (n_n1592) & (n_n1463) & (!x12188x) & (x12190x)) + ((n_n3810) & (n_n1592) & (n_n1463) & (x12188x) & (!x12190x)) + ((n_n3810) & (n_n1592) & (n_n1463) & (x12188x) & (x12190x)));
	assign x315x = (((!i_9_) & (n_n482) & (n_n534) & (n_n325)) + ((i_9_) & (n_n482) & (n_n534) & (n_n325)));
	assign x402x = (((!i_9_) & (n_n482) & (!n_n528) & (n_n325) & (n_n530)) + ((!i_9_) & (n_n482) & (n_n528) & (n_n325) & (n_n530)) + ((i_9_) & (n_n482) & (n_n528) & (n_n325) & (!n_n530)) + ((i_9_) & (n_n482) & (n_n528) & (n_n325) & (n_n530)));
	assign n_n1471 = (((!n_n4792) & (!n_n4793) & (!x179x) & (!n_n4799) & (!x22147x)) + ((!n_n4792) & (!n_n4793) & (!x179x) & (n_n4799) & (!x22147x)) + ((!n_n4792) & (!n_n4793) & (!x179x) & (n_n4799) & (x22147x)) + ((!n_n4792) & (!n_n4793) & (x179x) & (!n_n4799) & (!x22147x)) + ((!n_n4792) & (!n_n4793) & (x179x) & (!n_n4799) & (x22147x)) + ((!n_n4792) & (!n_n4793) & (x179x) & (n_n4799) & (!x22147x)) + ((!n_n4792) & (!n_n4793) & (x179x) & (n_n4799) & (x22147x)) + ((!n_n4792) & (n_n4793) & (!x179x) & (!n_n4799) & (!x22147x)) + ((!n_n4792) & (n_n4793) & (!x179x) & (!n_n4799) & (x22147x)) + ((!n_n4792) & (n_n4793) & (!x179x) & (n_n4799) & (!x22147x)) + ((!n_n4792) & (n_n4793) & (!x179x) & (n_n4799) & (x22147x)) + ((!n_n4792) & (n_n4793) & (x179x) & (!n_n4799) & (!x22147x)) + ((!n_n4792) & (n_n4793) & (x179x) & (!n_n4799) & (x22147x)) + ((!n_n4792) & (n_n4793) & (x179x) & (n_n4799) & (!x22147x)) + ((!n_n4792) & (n_n4793) & (x179x) & (n_n4799) & (x22147x)) + ((n_n4792) & (!n_n4793) & (!x179x) & (!n_n4799) & (!x22147x)) + ((n_n4792) & (!n_n4793) & (!x179x) & (!n_n4799) & (x22147x)) + ((n_n4792) & (!n_n4793) & (!x179x) & (n_n4799) & (!x22147x)) + ((n_n4792) & (!n_n4793) & (!x179x) & (n_n4799) & (x22147x)) + ((n_n4792) & (!n_n4793) & (x179x) & (!n_n4799) & (!x22147x)) + ((n_n4792) & (!n_n4793) & (x179x) & (!n_n4799) & (x22147x)) + ((n_n4792) & (!n_n4793) & (x179x) & (n_n4799) & (!x22147x)) + ((n_n4792) & (!n_n4793) & (x179x) & (n_n4799) & (x22147x)) + ((n_n4792) & (n_n4793) & (!x179x) & (!n_n4799) & (!x22147x)) + ((n_n4792) & (n_n4793) & (!x179x) & (!n_n4799) & (x22147x)) + ((n_n4792) & (n_n4793) & (!x179x) & (n_n4799) & (!x22147x)) + ((n_n4792) & (n_n4793) & (!x179x) & (n_n4799) & (x22147x)) + ((n_n4792) & (n_n4793) & (x179x) & (!n_n4799) & (!x22147x)) + ((n_n4792) & (n_n4793) & (x179x) & (!n_n4799) & (x22147x)) + ((n_n4792) & (n_n4793) & (x179x) & (n_n4799) & (!x22147x)) + ((n_n4792) & (n_n4793) & (x179x) & (n_n4799) & (x22147x)));
	assign x12209x = (((!n_n4779) & (!n_n4780) & (!n_n4783) & (!n_n4778) & (n_n4775)) + ((!n_n4779) & (!n_n4780) & (!n_n4783) & (n_n4778) & (!n_n4775)) + ((!n_n4779) & (!n_n4780) & (!n_n4783) & (n_n4778) & (n_n4775)) + ((!n_n4779) & (!n_n4780) & (n_n4783) & (!n_n4778) & (!n_n4775)) + ((!n_n4779) & (!n_n4780) & (n_n4783) & (!n_n4778) & (n_n4775)) + ((!n_n4779) & (!n_n4780) & (n_n4783) & (n_n4778) & (!n_n4775)) + ((!n_n4779) & (!n_n4780) & (n_n4783) & (n_n4778) & (n_n4775)) + ((!n_n4779) & (n_n4780) & (!n_n4783) & (!n_n4778) & (!n_n4775)) + ((!n_n4779) & (n_n4780) & (!n_n4783) & (!n_n4778) & (n_n4775)) + ((!n_n4779) & (n_n4780) & (!n_n4783) & (n_n4778) & (!n_n4775)) + ((!n_n4779) & (n_n4780) & (!n_n4783) & (n_n4778) & (n_n4775)) + ((!n_n4779) & (n_n4780) & (n_n4783) & (!n_n4778) & (!n_n4775)) + ((!n_n4779) & (n_n4780) & (n_n4783) & (!n_n4778) & (n_n4775)) + ((!n_n4779) & (n_n4780) & (n_n4783) & (n_n4778) & (!n_n4775)) + ((!n_n4779) & (n_n4780) & (n_n4783) & (n_n4778) & (n_n4775)) + ((n_n4779) & (!n_n4780) & (!n_n4783) & (!n_n4778) & (!n_n4775)) + ((n_n4779) & (!n_n4780) & (!n_n4783) & (!n_n4778) & (n_n4775)) + ((n_n4779) & (!n_n4780) & (!n_n4783) & (n_n4778) & (!n_n4775)) + ((n_n4779) & (!n_n4780) & (!n_n4783) & (n_n4778) & (n_n4775)) + ((n_n4779) & (!n_n4780) & (n_n4783) & (!n_n4778) & (!n_n4775)) + ((n_n4779) & (!n_n4780) & (n_n4783) & (!n_n4778) & (n_n4775)) + ((n_n4779) & (!n_n4780) & (n_n4783) & (n_n4778) & (!n_n4775)) + ((n_n4779) & (!n_n4780) & (n_n4783) & (n_n4778) & (n_n4775)) + ((n_n4779) & (n_n4780) & (!n_n4783) & (!n_n4778) & (!n_n4775)) + ((n_n4779) & (n_n4780) & (!n_n4783) & (!n_n4778) & (n_n4775)) + ((n_n4779) & (n_n4780) & (!n_n4783) & (n_n4778) & (!n_n4775)) + ((n_n4779) & (n_n4780) & (!n_n4783) & (n_n4778) & (n_n4775)) + ((n_n4779) & (n_n4780) & (n_n4783) & (!n_n4778) & (!n_n4775)) + ((n_n4779) & (n_n4780) & (n_n4783) & (!n_n4778) & (n_n4775)) + ((n_n4779) & (n_n4780) & (n_n4783) & (n_n4778) & (!n_n4775)) + ((n_n4779) & (n_n4780) & (n_n4783) & (n_n4778) & (n_n4775)));
	assign x12245x = (((!n_n4802) & (!n_n4805) & (!x71x) & (!n_n4197) & (x440x)) + ((!n_n4802) & (!n_n4805) & (!x71x) & (n_n4197) & (!x440x)) + ((!n_n4802) & (!n_n4805) & (!x71x) & (n_n4197) & (x440x)) + ((!n_n4802) & (!n_n4805) & (x71x) & (!n_n4197) & (!x440x)) + ((!n_n4802) & (!n_n4805) & (x71x) & (!n_n4197) & (x440x)) + ((!n_n4802) & (!n_n4805) & (x71x) & (n_n4197) & (!x440x)) + ((!n_n4802) & (!n_n4805) & (x71x) & (n_n4197) & (x440x)) + ((!n_n4802) & (n_n4805) & (!x71x) & (!n_n4197) & (!x440x)) + ((!n_n4802) & (n_n4805) & (!x71x) & (!n_n4197) & (x440x)) + ((!n_n4802) & (n_n4805) & (!x71x) & (n_n4197) & (!x440x)) + ((!n_n4802) & (n_n4805) & (!x71x) & (n_n4197) & (x440x)) + ((!n_n4802) & (n_n4805) & (x71x) & (!n_n4197) & (!x440x)) + ((!n_n4802) & (n_n4805) & (x71x) & (!n_n4197) & (x440x)) + ((!n_n4802) & (n_n4805) & (x71x) & (n_n4197) & (!x440x)) + ((!n_n4802) & (n_n4805) & (x71x) & (n_n4197) & (x440x)) + ((n_n4802) & (!n_n4805) & (!x71x) & (!n_n4197) & (!x440x)) + ((n_n4802) & (!n_n4805) & (!x71x) & (!n_n4197) & (x440x)) + ((n_n4802) & (!n_n4805) & (!x71x) & (n_n4197) & (!x440x)) + ((n_n4802) & (!n_n4805) & (!x71x) & (n_n4197) & (x440x)) + ((n_n4802) & (!n_n4805) & (x71x) & (!n_n4197) & (!x440x)) + ((n_n4802) & (!n_n4805) & (x71x) & (!n_n4197) & (x440x)) + ((n_n4802) & (!n_n4805) & (x71x) & (n_n4197) & (!x440x)) + ((n_n4802) & (!n_n4805) & (x71x) & (n_n4197) & (x440x)) + ((n_n4802) & (n_n4805) & (!x71x) & (!n_n4197) & (!x440x)) + ((n_n4802) & (n_n4805) & (!x71x) & (!n_n4197) & (x440x)) + ((n_n4802) & (n_n4805) & (!x71x) & (n_n4197) & (!x440x)) + ((n_n4802) & (n_n4805) & (!x71x) & (n_n4197) & (x440x)) + ((n_n4802) & (n_n4805) & (x71x) & (!n_n4197) & (!x440x)) + ((n_n4802) & (n_n4805) & (x71x) & (!n_n4197) & (x440x)) + ((n_n4802) & (n_n4805) & (x71x) & (n_n4197) & (!x440x)) + ((n_n4802) & (n_n4805) & (x71x) & (n_n4197) & (x440x)));
	assign x12247x = (((!x315x) & (!x402x) & (!n_n1471) & (!x12209x) & (x12245x)) + ((!x315x) & (!x402x) & (!n_n1471) & (x12209x) & (!x12245x)) + ((!x315x) & (!x402x) & (!n_n1471) & (x12209x) & (x12245x)) + ((!x315x) & (!x402x) & (n_n1471) & (!x12209x) & (!x12245x)) + ((!x315x) & (!x402x) & (n_n1471) & (!x12209x) & (x12245x)) + ((!x315x) & (!x402x) & (n_n1471) & (x12209x) & (!x12245x)) + ((!x315x) & (!x402x) & (n_n1471) & (x12209x) & (x12245x)) + ((!x315x) & (x402x) & (!n_n1471) & (!x12209x) & (!x12245x)) + ((!x315x) & (x402x) & (!n_n1471) & (!x12209x) & (x12245x)) + ((!x315x) & (x402x) & (!n_n1471) & (x12209x) & (!x12245x)) + ((!x315x) & (x402x) & (!n_n1471) & (x12209x) & (x12245x)) + ((!x315x) & (x402x) & (n_n1471) & (!x12209x) & (!x12245x)) + ((!x315x) & (x402x) & (n_n1471) & (!x12209x) & (x12245x)) + ((!x315x) & (x402x) & (n_n1471) & (x12209x) & (!x12245x)) + ((!x315x) & (x402x) & (n_n1471) & (x12209x) & (x12245x)) + ((x315x) & (!x402x) & (!n_n1471) & (!x12209x) & (!x12245x)) + ((x315x) & (!x402x) & (!n_n1471) & (!x12209x) & (x12245x)) + ((x315x) & (!x402x) & (!n_n1471) & (x12209x) & (!x12245x)) + ((x315x) & (!x402x) & (!n_n1471) & (x12209x) & (x12245x)) + ((x315x) & (!x402x) & (n_n1471) & (!x12209x) & (!x12245x)) + ((x315x) & (!x402x) & (n_n1471) & (!x12209x) & (x12245x)) + ((x315x) & (!x402x) & (n_n1471) & (x12209x) & (!x12245x)) + ((x315x) & (!x402x) & (n_n1471) & (x12209x) & (x12245x)) + ((x315x) & (x402x) & (!n_n1471) & (!x12209x) & (!x12245x)) + ((x315x) & (x402x) & (!n_n1471) & (!x12209x) & (x12245x)) + ((x315x) & (x402x) & (!n_n1471) & (x12209x) & (!x12245x)) + ((x315x) & (x402x) & (!n_n1471) & (x12209x) & (x12245x)) + ((x315x) & (x402x) & (n_n1471) & (!x12209x) & (!x12245x)) + ((x315x) & (x402x) & (n_n1471) & (!x12209x) & (x12245x)) + ((x315x) & (x402x) & (n_n1471) & (x12209x) & (!x12245x)) + ((x315x) & (x402x) & (n_n1471) & (x12209x) & (x12245x)));
	assign n_n1466 = (((!n_n4865) & (!x245x) & (!n_n4853) & (!n_n4852) & (!x22146x)) + ((!n_n4865) & (!x245x) & (!n_n4853) & (n_n4852) & (!x22146x)) + ((!n_n4865) & (!x245x) & (!n_n4853) & (n_n4852) & (x22146x)) + ((!n_n4865) & (!x245x) & (n_n4853) & (!n_n4852) & (!x22146x)) + ((!n_n4865) & (!x245x) & (n_n4853) & (!n_n4852) & (x22146x)) + ((!n_n4865) & (!x245x) & (n_n4853) & (n_n4852) & (!x22146x)) + ((!n_n4865) & (!x245x) & (n_n4853) & (n_n4852) & (x22146x)) + ((!n_n4865) & (x245x) & (!n_n4853) & (!n_n4852) & (!x22146x)) + ((!n_n4865) & (x245x) & (!n_n4853) & (!n_n4852) & (x22146x)) + ((!n_n4865) & (x245x) & (!n_n4853) & (n_n4852) & (!x22146x)) + ((!n_n4865) & (x245x) & (!n_n4853) & (n_n4852) & (x22146x)) + ((!n_n4865) & (x245x) & (n_n4853) & (!n_n4852) & (!x22146x)) + ((!n_n4865) & (x245x) & (n_n4853) & (!n_n4852) & (x22146x)) + ((!n_n4865) & (x245x) & (n_n4853) & (n_n4852) & (!x22146x)) + ((!n_n4865) & (x245x) & (n_n4853) & (n_n4852) & (x22146x)) + ((n_n4865) & (!x245x) & (!n_n4853) & (!n_n4852) & (!x22146x)) + ((n_n4865) & (!x245x) & (!n_n4853) & (!n_n4852) & (x22146x)) + ((n_n4865) & (!x245x) & (!n_n4853) & (n_n4852) & (!x22146x)) + ((n_n4865) & (!x245x) & (!n_n4853) & (n_n4852) & (x22146x)) + ((n_n4865) & (!x245x) & (n_n4853) & (!n_n4852) & (!x22146x)) + ((n_n4865) & (!x245x) & (n_n4853) & (!n_n4852) & (x22146x)) + ((n_n4865) & (!x245x) & (n_n4853) & (n_n4852) & (!x22146x)) + ((n_n4865) & (!x245x) & (n_n4853) & (n_n4852) & (x22146x)) + ((n_n4865) & (x245x) & (!n_n4853) & (!n_n4852) & (!x22146x)) + ((n_n4865) & (x245x) & (!n_n4853) & (!n_n4852) & (x22146x)) + ((n_n4865) & (x245x) & (!n_n4853) & (n_n4852) & (!x22146x)) + ((n_n4865) & (x245x) & (!n_n4853) & (n_n4852) & (x22146x)) + ((n_n4865) & (x245x) & (n_n4853) & (!n_n4852) & (!x22146x)) + ((n_n4865) & (x245x) & (n_n4853) & (!n_n4852) & (x22146x)) + ((n_n4865) & (x245x) & (n_n4853) & (n_n4852) & (!x22146x)) + ((n_n4865) & (x245x) & (n_n4853) & (n_n4852) & (x22146x)));
	assign x12223x = (((!n_n4870) & (!n_n4877) & (!n_n1985) & (!n_n3815) & (x12217x)) + ((!n_n4870) & (!n_n4877) & (!n_n1985) & (n_n3815) & (!x12217x)) + ((!n_n4870) & (!n_n4877) & (!n_n1985) & (n_n3815) & (x12217x)) + ((!n_n4870) & (!n_n4877) & (n_n1985) & (!n_n3815) & (!x12217x)) + ((!n_n4870) & (!n_n4877) & (n_n1985) & (!n_n3815) & (x12217x)) + ((!n_n4870) & (!n_n4877) & (n_n1985) & (n_n3815) & (!x12217x)) + ((!n_n4870) & (!n_n4877) & (n_n1985) & (n_n3815) & (x12217x)) + ((!n_n4870) & (n_n4877) & (!n_n1985) & (!n_n3815) & (!x12217x)) + ((!n_n4870) & (n_n4877) & (!n_n1985) & (!n_n3815) & (x12217x)) + ((!n_n4870) & (n_n4877) & (!n_n1985) & (n_n3815) & (!x12217x)) + ((!n_n4870) & (n_n4877) & (!n_n1985) & (n_n3815) & (x12217x)) + ((!n_n4870) & (n_n4877) & (n_n1985) & (!n_n3815) & (!x12217x)) + ((!n_n4870) & (n_n4877) & (n_n1985) & (!n_n3815) & (x12217x)) + ((!n_n4870) & (n_n4877) & (n_n1985) & (n_n3815) & (!x12217x)) + ((!n_n4870) & (n_n4877) & (n_n1985) & (n_n3815) & (x12217x)) + ((n_n4870) & (!n_n4877) & (!n_n1985) & (!n_n3815) & (!x12217x)) + ((n_n4870) & (!n_n4877) & (!n_n1985) & (!n_n3815) & (x12217x)) + ((n_n4870) & (!n_n4877) & (!n_n1985) & (n_n3815) & (!x12217x)) + ((n_n4870) & (!n_n4877) & (!n_n1985) & (n_n3815) & (x12217x)) + ((n_n4870) & (!n_n4877) & (n_n1985) & (!n_n3815) & (!x12217x)) + ((n_n4870) & (!n_n4877) & (n_n1985) & (!n_n3815) & (x12217x)) + ((n_n4870) & (!n_n4877) & (n_n1985) & (n_n3815) & (!x12217x)) + ((n_n4870) & (!n_n4877) & (n_n1985) & (n_n3815) & (x12217x)) + ((n_n4870) & (n_n4877) & (!n_n1985) & (!n_n3815) & (!x12217x)) + ((n_n4870) & (n_n4877) & (!n_n1985) & (!n_n3815) & (x12217x)) + ((n_n4870) & (n_n4877) & (!n_n1985) & (n_n3815) & (!x12217x)) + ((n_n4870) & (n_n4877) & (!n_n1985) & (n_n3815) & (x12217x)) + ((n_n4870) & (n_n4877) & (n_n1985) & (!n_n3815) & (!x12217x)) + ((n_n4870) & (n_n4877) & (n_n1985) & (!n_n3815) & (x12217x)) + ((n_n4870) & (n_n4877) & (n_n1985) & (n_n3815) & (!x12217x)) + ((n_n4870) & (n_n4877) & (n_n1985) & (n_n3815) & (x12217x)));
	assign n_n1415 = (((!n_n1468) & (!x12235x) & (!x12236x) & (x12240x)) + ((!n_n1468) & (!x12235x) & (x12236x) & (!x12240x)) + ((!n_n1468) & (!x12235x) & (x12236x) & (x12240x)) + ((!n_n1468) & (x12235x) & (!x12236x) & (!x12240x)) + ((!n_n1468) & (x12235x) & (!x12236x) & (x12240x)) + ((!n_n1468) & (x12235x) & (x12236x) & (!x12240x)) + ((!n_n1468) & (x12235x) & (x12236x) & (x12240x)) + ((n_n1468) & (!x12235x) & (!x12236x) & (!x12240x)) + ((n_n1468) & (!x12235x) & (!x12236x) & (x12240x)) + ((n_n1468) & (!x12235x) & (x12236x) & (!x12240x)) + ((n_n1468) & (!x12235x) & (x12236x) & (x12240x)) + ((n_n1468) & (x12235x) & (!x12236x) & (!x12240x)) + ((n_n1468) & (x12235x) & (!x12236x) & (x12240x)) + ((n_n1468) & (x12235x) & (x12236x) & (!x12240x)) + ((n_n1468) & (x12235x) & (x12236x) & (x12240x)));
	assign x12222x = (((!n_n4868) & (!n_n4880) & (!x330x) & (!x263x) & (x324x)) + ((!n_n4868) & (!n_n4880) & (!x330x) & (x263x) & (!x324x)) + ((!n_n4868) & (!n_n4880) & (!x330x) & (x263x) & (x324x)) + ((!n_n4868) & (!n_n4880) & (x330x) & (!x263x) & (!x324x)) + ((!n_n4868) & (!n_n4880) & (x330x) & (!x263x) & (x324x)) + ((!n_n4868) & (!n_n4880) & (x330x) & (x263x) & (!x324x)) + ((!n_n4868) & (!n_n4880) & (x330x) & (x263x) & (x324x)) + ((!n_n4868) & (n_n4880) & (!x330x) & (!x263x) & (!x324x)) + ((!n_n4868) & (n_n4880) & (!x330x) & (!x263x) & (x324x)) + ((!n_n4868) & (n_n4880) & (!x330x) & (x263x) & (!x324x)) + ((!n_n4868) & (n_n4880) & (!x330x) & (x263x) & (x324x)) + ((!n_n4868) & (n_n4880) & (x330x) & (!x263x) & (!x324x)) + ((!n_n4868) & (n_n4880) & (x330x) & (!x263x) & (x324x)) + ((!n_n4868) & (n_n4880) & (x330x) & (x263x) & (!x324x)) + ((!n_n4868) & (n_n4880) & (x330x) & (x263x) & (x324x)) + ((n_n4868) & (!n_n4880) & (!x330x) & (!x263x) & (!x324x)) + ((n_n4868) & (!n_n4880) & (!x330x) & (!x263x) & (x324x)) + ((n_n4868) & (!n_n4880) & (!x330x) & (x263x) & (!x324x)) + ((n_n4868) & (!n_n4880) & (!x330x) & (x263x) & (x324x)) + ((n_n4868) & (!n_n4880) & (x330x) & (!x263x) & (!x324x)) + ((n_n4868) & (!n_n4880) & (x330x) & (!x263x) & (x324x)) + ((n_n4868) & (!n_n4880) & (x330x) & (x263x) & (!x324x)) + ((n_n4868) & (!n_n4880) & (x330x) & (x263x) & (x324x)) + ((n_n4868) & (n_n4880) & (!x330x) & (!x263x) & (!x324x)) + ((n_n4868) & (n_n4880) & (!x330x) & (!x263x) & (x324x)) + ((n_n4868) & (n_n4880) & (!x330x) & (x263x) & (!x324x)) + ((n_n4868) & (n_n4880) & (!x330x) & (x263x) & (x324x)) + ((n_n4868) & (n_n4880) & (x330x) & (!x263x) & (!x324x)) + ((n_n4868) & (n_n4880) & (x330x) & (!x263x) & (x324x)) + ((n_n4868) & (n_n4880) & (x330x) & (x263x) & (!x324x)) + ((n_n4868) & (n_n4880) & (x330x) & (x263x) & (x324x)));
	assign n_n1450 = (((!n_n5060) & (!n_n5055) & (!n_n5059) & (!n_n5056) & (x12311x)) + ((!n_n5060) & (!n_n5055) & (!n_n5059) & (n_n5056) & (!x12311x)) + ((!n_n5060) & (!n_n5055) & (!n_n5059) & (n_n5056) & (x12311x)) + ((!n_n5060) & (!n_n5055) & (n_n5059) & (!n_n5056) & (!x12311x)) + ((!n_n5060) & (!n_n5055) & (n_n5059) & (!n_n5056) & (x12311x)) + ((!n_n5060) & (!n_n5055) & (n_n5059) & (n_n5056) & (!x12311x)) + ((!n_n5060) & (!n_n5055) & (n_n5059) & (n_n5056) & (x12311x)) + ((!n_n5060) & (n_n5055) & (!n_n5059) & (!n_n5056) & (!x12311x)) + ((!n_n5060) & (n_n5055) & (!n_n5059) & (!n_n5056) & (x12311x)) + ((!n_n5060) & (n_n5055) & (!n_n5059) & (n_n5056) & (!x12311x)) + ((!n_n5060) & (n_n5055) & (!n_n5059) & (n_n5056) & (x12311x)) + ((!n_n5060) & (n_n5055) & (n_n5059) & (!n_n5056) & (!x12311x)) + ((!n_n5060) & (n_n5055) & (n_n5059) & (!n_n5056) & (x12311x)) + ((!n_n5060) & (n_n5055) & (n_n5059) & (n_n5056) & (!x12311x)) + ((!n_n5060) & (n_n5055) & (n_n5059) & (n_n5056) & (x12311x)) + ((n_n5060) & (!n_n5055) & (!n_n5059) & (!n_n5056) & (!x12311x)) + ((n_n5060) & (!n_n5055) & (!n_n5059) & (!n_n5056) & (x12311x)) + ((n_n5060) & (!n_n5055) & (!n_n5059) & (n_n5056) & (!x12311x)) + ((n_n5060) & (!n_n5055) & (!n_n5059) & (n_n5056) & (x12311x)) + ((n_n5060) & (!n_n5055) & (n_n5059) & (!n_n5056) & (!x12311x)) + ((n_n5060) & (!n_n5055) & (n_n5059) & (!n_n5056) & (x12311x)) + ((n_n5060) & (!n_n5055) & (n_n5059) & (n_n5056) & (!x12311x)) + ((n_n5060) & (!n_n5055) & (n_n5059) & (n_n5056) & (x12311x)) + ((n_n5060) & (n_n5055) & (!n_n5059) & (!n_n5056) & (!x12311x)) + ((n_n5060) & (n_n5055) & (!n_n5059) & (!n_n5056) & (x12311x)) + ((n_n5060) & (n_n5055) & (!n_n5059) & (n_n5056) & (!x12311x)) + ((n_n5060) & (n_n5055) & (!n_n5059) & (n_n5056) & (x12311x)) + ((n_n5060) & (n_n5055) & (n_n5059) & (!n_n5056) & (!x12311x)) + ((n_n5060) & (n_n5055) & (n_n5059) & (!n_n5056) & (x12311x)) + ((n_n5060) & (n_n5055) & (n_n5059) & (n_n5056) & (!x12311x)) + ((n_n5060) & (n_n5055) & (n_n5059) & (n_n5056) & (x12311x)));
	assign n_n1451 = (((!n_n5054) & (!n_n5042) & (!x97x) & (x12316x)) + ((!n_n5054) & (!n_n5042) & (x97x) & (!x12316x)) + ((!n_n5054) & (!n_n5042) & (x97x) & (x12316x)) + ((!n_n5054) & (n_n5042) & (!x97x) & (!x12316x)) + ((!n_n5054) & (n_n5042) & (!x97x) & (x12316x)) + ((!n_n5054) & (n_n5042) & (x97x) & (!x12316x)) + ((!n_n5054) & (n_n5042) & (x97x) & (x12316x)) + ((n_n5054) & (!n_n5042) & (!x97x) & (!x12316x)) + ((n_n5054) & (!n_n5042) & (!x97x) & (x12316x)) + ((n_n5054) & (!n_n5042) & (x97x) & (!x12316x)) + ((n_n5054) & (!n_n5042) & (x97x) & (x12316x)) + ((n_n5054) & (n_n5042) & (!x97x) & (!x12316x)) + ((n_n5054) & (n_n5042) & (!x97x) & (x12316x)) + ((n_n5054) & (n_n5042) & (x97x) & (!x12316x)) + ((n_n5054) & (n_n5042) & (x97x) & (x12316x)));
	assign x12324x = (((!n_n5075) & (!n_n5068) & (!x12321x) & (x12322x)) + ((!n_n5075) & (!n_n5068) & (x12321x) & (!x12322x)) + ((!n_n5075) & (!n_n5068) & (x12321x) & (x12322x)) + ((!n_n5075) & (n_n5068) & (!x12321x) & (!x12322x)) + ((!n_n5075) & (n_n5068) & (!x12321x) & (x12322x)) + ((!n_n5075) & (n_n5068) & (x12321x) & (!x12322x)) + ((!n_n5075) & (n_n5068) & (x12321x) & (x12322x)) + ((n_n5075) & (!n_n5068) & (!x12321x) & (!x12322x)) + ((n_n5075) & (!n_n5068) & (!x12321x) & (x12322x)) + ((n_n5075) & (!n_n5068) & (x12321x) & (!x12322x)) + ((n_n5075) & (!n_n5068) & (x12321x) & (x12322x)) + ((n_n5075) & (n_n5068) & (!x12321x) & (!x12322x)) + ((n_n5075) & (n_n5068) & (!x12321x) & (x12322x)) + ((n_n5075) & (n_n5068) & (x12321x) & (!x12322x)) + ((n_n5075) & (n_n5068) & (x12321x) & (x12322x)));
	assign n_n1408 = (((!n_n1446) & (!x12333x) & (!x12334x) & (!x12338x) & (x12339x)) + ((!n_n1446) & (!x12333x) & (!x12334x) & (x12338x) & (!x12339x)) + ((!n_n1446) & (!x12333x) & (!x12334x) & (x12338x) & (x12339x)) + ((!n_n1446) & (!x12333x) & (x12334x) & (!x12338x) & (!x12339x)) + ((!n_n1446) & (!x12333x) & (x12334x) & (!x12338x) & (x12339x)) + ((!n_n1446) & (!x12333x) & (x12334x) & (x12338x) & (!x12339x)) + ((!n_n1446) & (!x12333x) & (x12334x) & (x12338x) & (x12339x)) + ((!n_n1446) & (x12333x) & (!x12334x) & (!x12338x) & (!x12339x)) + ((!n_n1446) & (x12333x) & (!x12334x) & (!x12338x) & (x12339x)) + ((!n_n1446) & (x12333x) & (!x12334x) & (x12338x) & (!x12339x)) + ((!n_n1446) & (x12333x) & (!x12334x) & (x12338x) & (x12339x)) + ((!n_n1446) & (x12333x) & (x12334x) & (!x12338x) & (!x12339x)) + ((!n_n1446) & (x12333x) & (x12334x) & (!x12338x) & (x12339x)) + ((!n_n1446) & (x12333x) & (x12334x) & (x12338x) & (!x12339x)) + ((!n_n1446) & (x12333x) & (x12334x) & (x12338x) & (x12339x)) + ((n_n1446) & (!x12333x) & (!x12334x) & (!x12338x) & (!x12339x)) + ((n_n1446) & (!x12333x) & (!x12334x) & (!x12338x) & (x12339x)) + ((n_n1446) & (!x12333x) & (!x12334x) & (x12338x) & (!x12339x)) + ((n_n1446) & (!x12333x) & (!x12334x) & (x12338x) & (x12339x)) + ((n_n1446) & (!x12333x) & (x12334x) & (!x12338x) & (!x12339x)) + ((n_n1446) & (!x12333x) & (x12334x) & (!x12338x) & (x12339x)) + ((n_n1446) & (!x12333x) & (x12334x) & (x12338x) & (!x12339x)) + ((n_n1446) & (!x12333x) & (x12334x) & (x12338x) & (x12339x)) + ((n_n1446) & (x12333x) & (!x12334x) & (!x12338x) & (!x12339x)) + ((n_n1446) & (x12333x) & (!x12334x) & (!x12338x) & (x12339x)) + ((n_n1446) & (x12333x) & (!x12334x) & (x12338x) & (!x12339x)) + ((n_n1446) & (x12333x) & (!x12334x) & (x12338x) & (x12339x)) + ((n_n1446) & (x12333x) & (x12334x) & (!x12338x) & (!x12339x)) + ((n_n1446) & (x12333x) & (x12334x) & (!x12338x) & (x12339x)) + ((n_n1446) & (x12333x) & (x12334x) & (x12338x) & (!x12339x)) + ((n_n1446) & (x12333x) & (x12334x) & (x12338x) & (x12339x)));
	assign x12389x = (((!n_n1453) & (!n_n1454) & (!x12385x) & (x12386x)) + ((!n_n1453) & (!n_n1454) & (x12385x) & (!x12386x)) + ((!n_n1453) & (!n_n1454) & (x12385x) & (x12386x)) + ((!n_n1453) & (n_n1454) & (!x12385x) & (!x12386x)) + ((!n_n1453) & (n_n1454) & (!x12385x) & (x12386x)) + ((!n_n1453) & (n_n1454) & (x12385x) & (!x12386x)) + ((!n_n1453) & (n_n1454) & (x12385x) & (x12386x)) + ((n_n1453) & (!n_n1454) & (!x12385x) & (!x12386x)) + ((n_n1453) & (!n_n1454) & (!x12385x) & (x12386x)) + ((n_n1453) & (!n_n1454) & (x12385x) & (!x12386x)) + ((n_n1453) & (!n_n1454) & (x12385x) & (x12386x)) + ((n_n1453) & (n_n1454) & (!x12385x) & (!x12386x)) + ((n_n1453) & (n_n1454) & (!x12385x) & (x12386x)) + ((n_n1453) & (n_n1454) & (x12385x) & (!x12386x)) + ((n_n1453) & (n_n1454) & (x12385x) & (x12386x)));
	assign n_n1473 = (((!n_n4762) & (!n_n4765) & (!n_n4766) & (!n_n4205) & (x12394x)) + ((!n_n4762) & (!n_n4765) & (!n_n4766) & (n_n4205) & (!x12394x)) + ((!n_n4762) & (!n_n4765) & (!n_n4766) & (n_n4205) & (x12394x)) + ((!n_n4762) & (!n_n4765) & (n_n4766) & (!n_n4205) & (!x12394x)) + ((!n_n4762) & (!n_n4765) & (n_n4766) & (!n_n4205) & (x12394x)) + ((!n_n4762) & (!n_n4765) & (n_n4766) & (n_n4205) & (!x12394x)) + ((!n_n4762) & (!n_n4765) & (n_n4766) & (n_n4205) & (x12394x)) + ((!n_n4762) & (n_n4765) & (!n_n4766) & (!n_n4205) & (!x12394x)) + ((!n_n4762) & (n_n4765) & (!n_n4766) & (!n_n4205) & (x12394x)) + ((!n_n4762) & (n_n4765) & (!n_n4766) & (n_n4205) & (!x12394x)) + ((!n_n4762) & (n_n4765) & (!n_n4766) & (n_n4205) & (x12394x)) + ((!n_n4762) & (n_n4765) & (n_n4766) & (!n_n4205) & (!x12394x)) + ((!n_n4762) & (n_n4765) & (n_n4766) & (!n_n4205) & (x12394x)) + ((!n_n4762) & (n_n4765) & (n_n4766) & (n_n4205) & (!x12394x)) + ((!n_n4762) & (n_n4765) & (n_n4766) & (n_n4205) & (x12394x)) + ((n_n4762) & (!n_n4765) & (!n_n4766) & (!n_n4205) & (!x12394x)) + ((n_n4762) & (!n_n4765) & (!n_n4766) & (!n_n4205) & (x12394x)) + ((n_n4762) & (!n_n4765) & (!n_n4766) & (n_n4205) & (!x12394x)) + ((n_n4762) & (!n_n4765) & (!n_n4766) & (n_n4205) & (x12394x)) + ((n_n4762) & (!n_n4765) & (n_n4766) & (!n_n4205) & (!x12394x)) + ((n_n4762) & (!n_n4765) & (n_n4766) & (!n_n4205) & (x12394x)) + ((n_n4762) & (!n_n4765) & (n_n4766) & (n_n4205) & (!x12394x)) + ((n_n4762) & (!n_n4765) & (n_n4766) & (n_n4205) & (x12394x)) + ((n_n4762) & (n_n4765) & (!n_n4766) & (!n_n4205) & (!x12394x)) + ((n_n4762) & (n_n4765) & (!n_n4766) & (!n_n4205) & (x12394x)) + ((n_n4762) & (n_n4765) & (!n_n4766) & (n_n4205) & (!x12394x)) + ((n_n4762) & (n_n4765) & (!n_n4766) & (n_n4205) & (x12394x)) + ((n_n4762) & (n_n4765) & (n_n4766) & (!n_n4205) & (!x12394x)) + ((n_n4762) & (n_n4765) & (n_n4766) & (!n_n4205) & (x12394x)) + ((n_n4762) & (n_n4765) & (n_n4766) & (n_n4205) & (!x12394x)) + ((n_n4762) & (n_n4765) & (n_n4766) & (n_n4205) & (x12394x)));
	assign n_n1475 = (((!x483x) & (!x20x) & (!n_n4740) & (!n_n3475) & (!x22143x)) + ((!x483x) & (!x20x) & (!n_n4740) & (n_n3475) & (!x22143x)) + ((!x483x) & (!x20x) & (!n_n4740) & (n_n3475) & (x22143x)) + ((!x483x) & (!x20x) & (n_n4740) & (!n_n3475) & (!x22143x)) + ((!x483x) & (!x20x) & (n_n4740) & (!n_n3475) & (x22143x)) + ((!x483x) & (!x20x) & (n_n4740) & (n_n3475) & (!x22143x)) + ((!x483x) & (!x20x) & (n_n4740) & (n_n3475) & (x22143x)) + ((!x483x) & (x20x) & (!n_n4740) & (!n_n3475) & (!x22143x)) + ((!x483x) & (x20x) & (!n_n4740) & (n_n3475) & (!x22143x)) + ((!x483x) & (x20x) & (!n_n4740) & (n_n3475) & (x22143x)) + ((!x483x) & (x20x) & (n_n4740) & (!n_n3475) & (!x22143x)) + ((!x483x) & (x20x) & (n_n4740) & (!n_n3475) & (x22143x)) + ((!x483x) & (x20x) & (n_n4740) & (n_n3475) & (!x22143x)) + ((!x483x) & (x20x) & (n_n4740) & (n_n3475) & (x22143x)) + ((x483x) & (!x20x) & (!n_n4740) & (!n_n3475) & (!x22143x)) + ((x483x) & (!x20x) & (!n_n4740) & (n_n3475) & (!x22143x)) + ((x483x) & (!x20x) & (!n_n4740) & (n_n3475) & (x22143x)) + ((x483x) & (!x20x) & (n_n4740) & (!n_n3475) & (!x22143x)) + ((x483x) & (!x20x) & (n_n4740) & (!n_n3475) & (x22143x)) + ((x483x) & (!x20x) & (n_n4740) & (n_n3475) & (!x22143x)) + ((x483x) & (!x20x) & (n_n4740) & (n_n3475) & (x22143x)) + ((x483x) & (x20x) & (!n_n4740) & (!n_n3475) & (!x22143x)) + ((x483x) & (x20x) & (!n_n4740) & (!n_n3475) & (x22143x)) + ((x483x) & (x20x) & (!n_n4740) & (n_n3475) & (!x22143x)) + ((x483x) & (x20x) & (!n_n4740) & (n_n3475) & (x22143x)) + ((x483x) & (x20x) & (n_n4740) & (!n_n3475) & (!x22143x)) + ((x483x) & (x20x) & (n_n4740) & (!n_n3475) & (x22143x)) + ((x483x) & (x20x) & (n_n4740) & (n_n3475) & (!x22143x)) + ((x483x) & (x20x) & (n_n4740) & (n_n3475) & (x22143x)));
	assign x12436x = (((!n_n4754) & (!n_n4757) & (!n_n4749) & (n_n4760)) + ((!n_n4754) & (!n_n4757) & (n_n4749) & (!n_n4760)) + ((!n_n4754) & (!n_n4757) & (n_n4749) & (n_n4760)) + ((!n_n4754) & (n_n4757) & (!n_n4749) & (!n_n4760)) + ((!n_n4754) & (n_n4757) & (!n_n4749) & (n_n4760)) + ((!n_n4754) & (n_n4757) & (n_n4749) & (!n_n4760)) + ((!n_n4754) & (n_n4757) & (n_n4749) & (n_n4760)) + ((n_n4754) & (!n_n4757) & (!n_n4749) & (!n_n4760)) + ((n_n4754) & (!n_n4757) & (!n_n4749) & (n_n4760)) + ((n_n4754) & (!n_n4757) & (n_n4749) & (!n_n4760)) + ((n_n4754) & (!n_n4757) & (n_n4749) & (n_n4760)) + ((n_n4754) & (n_n4757) & (!n_n4749) & (!n_n4760)) + ((n_n4754) & (n_n4757) & (!n_n4749) & (n_n4760)) + ((n_n4754) & (n_n4757) & (n_n4749) & (!n_n4760)) + ((n_n4754) & (n_n4757) & (n_n4749) & (n_n4760)));
	assign x12437x = (((!n_n4748) & (!n_n4747) & (!n_n4755) & (!n_n4761) & (n_n4752)) + ((!n_n4748) & (!n_n4747) & (!n_n4755) & (n_n4761) & (!n_n4752)) + ((!n_n4748) & (!n_n4747) & (!n_n4755) & (n_n4761) & (n_n4752)) + ((!n_n4748) & (!n_n4747) & (n_n4755) & (!n_n4761) & (!n_n4752)) + ((!n_n4748) & (!n_n4747) & (n_n4755) & (!n_n4761) & (n_n4752)) + ((!n_n4748) & (!n_n4747) & (n_n4755) & (n_n4761) & (!n_n4752)) + ((!n_n4748) & (!n_n4747) & (n_n4755) & (n_n4761) & (n_n4752)) + ((!n_n4748) & (n_n4747) & (!n_n4755) & (!n_n4761) & (!n_n4752)) + ((!n_n4748) & (n_n4747) & (!n_n4755) & (!n_n4761) & (n_n4752)) + ((!n_n4748) & (n_n4747) & (!n_n4755) & (n_n4761) & (!n_n4752)) + ((!n_n4748) & (n_n4747) & (!n_n4755) & (n_n4761) & (n_n4752)) + ((!n_n4748) & (n_n4747) & (n_n4755) & (!n_n4761) & (!n_n4752)) + ((!n_n4748) & (n_n4747) & (n_n4755) & (!n_n4761) & (n_n4752)) + ((!n_n4748) & (n_n4747) & (n_n4755) & (n_n4761) & (!n_n4752)) + ((!n_n4748) & (n_n4747) & (n_n4755) & (n_n4761) & (n_n4752)) + ((n_n4748) & (!n_n4747) & (!n_n4755) & (!n_n4761) & (!n_n4752)) + ((n_n4748) & (!n_n4747) & (!n_n4755) & (!n_n4761) & (n_n4752)) + ((n_n4748) & (!n_n4747) & (!n_n4755) & (n_n4761) & (!n_n4752)) + ((n_n4748) & (!n_n4747) & (!n_n4755) & (n_n4761) & (n_n4752)) + ((n_n4748) & (!n_n4747) & (n_n4755) & (!n_n4761) & (!n_n4752)) + ((n_n4748) & (!n_n4747) & (n_n4755) & (!n_n4761) & (n_n4752)) + ((n_n4748) & (!n_n4747) & (n_n4755) & (n_n4761) & (!n_n4752)) + ((n_n4748) & (!n_n4747) & (n_n4755) & (n_n4761) & (n_n4752)) + ((n_n4748) & (n_n4747) & (!n_n4755) & (!n_n4761) & (!n_n4752)) + ((n_n4748) & (n_n4747) & (!n_n4755) & (!n_n4761) & (n_n4752)) + ((n_n4748) & (n_n4747) & (!n_n4755) & (n_n4761) & (!n_n4752)) + ((n_n4748) & (n_n4747) & (!n_n4755) & (n_n4761) & (n_n4752)) + ((n_n4748) & (n_n4747) & (n_n4755) & (!n_n4761) & (!n_n4752)) + ((n_n4748) & (n_n4747) & (n_n4755) & (!n_n4761) & (n_n4752)) + ((n_n4748) & (n_n4747) & (n_n4755) & (n_n4761) & (!n_n4752)) + ((n_n4748) & (n_n4747) & (n_n4755) & (n_n4761) & (n_n4752)));
	assign x12440x = (((!n_n1473) & (!n_n1475) & (!x12436x) & (x12437x)) + ((!n_n1473) & (!n_n1475) & (x12436x) & (!x12437x)) + ((!n_n1473) & (!n_n1475) & (x12436x) & (x12437x)) + ((!n_n1473) & (n_n1475) & (!x12436x) & (!x12437x)) + ((!n_n1473) & (n_n1475) & (!x12436x) & (x12437x)) + ((!n_n1473) & (n_n1475) & (x12436x) & (!x12437x)) + ((!n_n1473) & (n_n1475) & (x12436x) & (x12437x)) + ((n_n1473) & (!n_n1475) & (!x12436x) & (!x12437x)) + ((n_n1473) & (!n_n1475) & (!x12436x) & (x12437x)) + ((n_n1473) & (!n_n1475) & (x12436x) & (!x12437x)) + ((n_n1473) & (!n_n1475) & (x12436x) & (x12437x)) + ((n_n1473) & (n_n1475) & (!x12436x) & (!x12437x)) + ((n_n1473) & (n_n1475) & (!x12436x) & (x12437x)) + ((n_n1473) & (n_n1475) & (x12436x) & (!x12437x)) + ((n_n1473) & (n_n1475) & (x12436x) & (x12437x)));
	assign n_n1480 = (((!n_n4674) & (!n_n4671) & (!n_n1636) & (!x417x) & (x12418x)) + ((!n_n4674) & (!n_n4671) & (!n_n1636) & (x417x) & (!x12418x)) + ((!n_n4674) & (!n_n4671) & (!n_n1636) & (x417x) & (x12418x)) + ((!n_n4674) & (!n_n4671) & (n_n1636) & (!x417x) & (!x12418x)) + ((!n_n4674) & (!n_n4671) & (n_n1636) & (!x417x) & (x12418x)) + ((!n_n4674) & (!n_n4671) & (n_n1636) & (x417x) & (!x12418x)) + ((!n_n4674) & (!n_n4671) & (n_n1636) & (x417x) & (x12418x)) + ((!n_n4674) & (n_n4671) & (!n_n1636) & (!x417x) & (!x12418x)) + ((!n_n4674) & (n_n4671) & (!n_n1636) & (!x417x) & (x12418x)) + ((!n_n4674) & (n_n4671) & (!n_n1636) & (x417x) & (!x12418x)) + ((!n_n4674) & (n_n4671) & (!n_n1636) & (x417x) & (x12418x)) + ((!n_n4674) & (n_n4671) & (n_n1636) & (!x417x) & (!x12418x)) + ((!n_n4674) & (n_n4671) & (n_n1636) & (!x417x) & (x12418x)) + ((!n_n4674) & (n_n4671) & (n_n1636) & (x417x) & (!x12418x)) + ((!n_n4674) & (n_n4671) & (n_n1636) & (x417x) & (x12418x)) + ((n_n4674) & (!n_n4671) & (!n_n1636) & (!x417x) & (!x12418x)) + ((n_n4674) & (!n_n4671) & (!n_n1636) & (!x417x) & (x12418x)) + ((n_n4674) & (!n_n4671) & (!n_n1636) & (x417x) & (!x12418x)) + ((n_n4674) & (!n_n4671) & (!n_n1636) & (x417x) & (x12418x)) + ((n_n4674) & (!n_n4671) & (n_n1636) & (!x417x) & (!x12418x)) + ((n_n4674) & (!n_n4671) & (n_n1636) & (!x417x) & (x12418x)) + ((n_n4674) & (!n_n4671) & (n_n1636) & (x417x) & (!x12418x)) + ((n_n4674) & (!n_n4671) & (n_n1636) & (x417x) & (x12418x)) + ((n_n4674) & (n_n4671) & (!n_n1636) & (!x417x) & (!x12418x)) + ((n_n4674) & (n_n4671) & (!n_n1636) & (!x417x) & (x12418x)) + ((n_n4674) & (n_n4671) & (!n_n1636) & (x417x) & (!x12418x)) + ((n_n4674) & (n_n4671) & (!n_n1636) & (x417x) & (x12418x)) + ((n_n4674) & (n_n4671) & (n_n1636) & (!x417x) & (!x12418x)) + ((n_n4674) & (n_n4671) & (n_n1636) & (!x417x) & (x12418x)) + ((n_n4674) & (n_n4671) & (n_n1636) & (x417x) & (!x12418x)) + ((n_n4674) & (n_n4671) & (n_n1636) & (x417x) & (x12418x)));
	assign n_n1418 = (((!x12416x) & (!x12404x) & (!x12405x) & (n_n1476)) + ((!x12416x) & (!x12404x) & (x12405x) & (!n_n1476)) + ((!x12416x) & (!x12404x) & (x12405x) & (n_n1476)) + ((!x12416x) & (x12404x) & (!x12405x) & (!n_n1476)) + ((!x12416x) & (x12404x) & (!x12405x) & (n_n1476)) + ((!x12416x) & (x12404x) & (x12405x) & (!n_n1476)) + ((!x12416x) & (x12404x) & (x12405x) & (n_n1476)) + ((x12416x) & (!x12404x) & (!x12405x) & (!n_n1476)) + ((x12416x) & (!x12404x) & (!x12405x) & (n_n1476)) + ((x12416x) & (!x12404x) & (x12405x) & (!n_n1476)) + ((x12416x) & (!x12404x) & (x12405x) & (n_n1476)) + ((x12416x) & (x12404x) & (!x12405x) & (!n_n1476)) + ((x12416x) & (x12404x) & (!x12405x) & (n_n1476)) + ((x12416x) & (x12404x) & (x12405x) & (!n_n1476)) + ((x12416x) & (x12404x) & (x12405x) & (n_n1476)));
	assign x12431x = (((!x10x) & (!n_n530) & (!n_n464) & (!n_n4689) & (!x22206x)) + ((!x10x) & (!n_n530) & (!n_n464) & (n_n4689) & (!x22206x)) + ((!x10x) & (!n_n530) & (!n_n464) & (n_n4689) & (x22206x)) + ((!x10x) & (!n_n530) & (n_n464) & (!n_n4689) & (!x22206x)) + ((!x10x) & (!n_n530) & (n_n464) & (n_n4689) & (!x22206x)) + ((!x10x) & (!n_n530) & (n_n464) & (n_n4689) & (x22206x)) + ((!x10x) & (n_n530) & (!n_n464) & (!n_n4689) & (!x22206x)) + ((!x10x) & (n_n530) & (!n_n464) & (n_n4689) & (!x22206x)) + ((!x10x) & (n_n530) & (!n_n464) & (n_n4689) & (x22206x)) + ((!x10x) & (n_n530) & (n_n464) & (!n_n4689) & (!x22206x)) + ((!x10x) & (n_n530) & (n_n464) & (n_n4689) & (!x22206x)) + ((!x10x) & (n_n530) & (n_n464) & (n_n4689) & (x22206x)) + ((x10x) & (!n_n530) & (!n_n464) & (!n_n4689) & (!x22206x)) + ((x10x) & (!n_n530) & (!n_n464) & (n_n4689) & (!x22206x)) + ((x10x) & (!n_n530) & (!n_n464) & (n_n4689) & (x22206x)) + ((x10x) & (!n_n530) & (n_n464) & (!n_n4689) & (!x22206x)) + ((x10x) & (!n_n530) & (n_n464) & (n_n4689) & (!x22206x)) + ((x10x) & (!n_n530) & (n_n464) & (n_n4689) & (x22206x)) + ((x10x) & (n_n530) & (!n_n464) & (!n_n4689) & (!x22206x)) + ((x10x) & (n_n530) & (!n_n464) & (n_n4689) & (!x22206x)) + ((x10x) & (n_n530) & (!n_n464) & (n_n4689) & (x22206x)) + ((x10x) & (n_n530) & (n_n464) & (!n_n4689) & (!x22206x)) + ((x10x) & (n_n530) & (n_n464) & (!n_n4689) & (x22206x)) + ((x10x) & (n_n530) & (n_n464) & (n_n4689) & (!x22206x)) + ((x10x) & (n_n530) & (n_n464) & (n_n4689) & (x22206x)));
	assign n_n1481 = (((!n_n4667) & (!n_n4662) & (!n_n4660) & (!x72x) & (x12425x)) + ((!n_n4667) & (!n_n4662) & (!n_n4660) & (x72x) & (!x12425x)) + ((!n_n4667) & (!n_n4662) & (!n_n4660) & (x72x) & (x12425x)) + ((!n_n4667) & (!n_n4662) & (n_n4660) & (!x72x) & (!x12425x)) + ((!n_n4667) & (!n_n4662) & (n_n4660) & (!x72x) & (x12425x)) + ((!n_n4667) & (!n_n4662) & (n_n4660) & (x72x) & (!x12425x)) + ((!n_n4667) & (!n_n4662) & (n_n4660) & (x72x) & (x12425x)) + ((!n_n4667) & (n_n4662) & (!n_n4660) & (!x72x) & (!x12425x)) + ((!n_n4667) & (n_n4662) & (!n_n4660) & (!x72x) & (x12425x)) + ((!n_n4667) & (n_n4662) & (!n_n4660) & (x72x) & (!x12425x)) + ((!n_n4667) & (n_n4662) & (!n_n4660) & (x72x) & (x12425x)) + ((!n_n4667) & (n_n4662) & (n_n4660) & (!x72x) & (!x12425x)) + ((!n_n4667) & (n_n4662) & (n_n4660) & (!x72x) & (x12425x)) + ((!n_n4667) & (n_n4662) & (n_n4660) & (x72x) & (!x12425x)) + ((!n_n4667) & (n_n4662) & (n_n4660) & (x72x) & (x12425x)) + ((n_n4667) & (!n_n4662) & (!n_n4660) & (!x72x) & (!x12425x)) + ((n_n4667) & (!n_n4662) & (!n_n4660) & (!x72x) & (x12425x)) + ((n_n4667) & (!n_n4662) & (!n_n4660) & (x72x) & (!x12425x)) + ((n_n4667) & (!n_n4662) & (!n_n4660) & (x72x) & (x12425x)) + ((n_n4667) & (!n_n4662) & (n_n4660) & (!x72x) & (!x12425x)) + ((n_n4667) & (!n_n4662) & (n_n4660) & (!x72x) & (x12425x)) + ((n_n4667) & (!n_n4662) & (n_n4660) & (x72x) & (!x12425x)) + ((n_n4667) & (!n_n4662) & (n_n4660) & (x72x) & (x12425x)) + ((n_n4667) & (n_n4662) & (!n_n4660) & (!x72x) & (!x12425x)) + ((n_n4667) & (n_n4662) & (!n_n4660) & (!x72x) & (x12425x)) + ((n_n4667) & (n_n4662) & (!n_n4660) & (x72x) & (!x12425x)) + ((n_n4667) & (n_n4662) & (!n_n4660) & (x72x) & (x12425x)) + ((n_n4667) & (n_n4662) & (n_n4660) & (!x72x) & (!x12425x)) + ((n_n4667) & (n_n4662) & (n_n4660) & (!x72x) & (x12425x)) + ((n_n4667) & (n_n4662) & (n_n4660) & (x72x) & (!x12425x)) + ((n_n4667) & (n_n4662) & (n_n4660) & (x72x) & (x12425x)));
	assign n_n1427 = (((!n_n3903) & (!n_n1504) & (!n_n1693) & (!x12452x) & (x12454x)) + ((!n_n3903) & (!n_n1504) & (!n_n1693) & (x12452x) & (!x12454x)) + ((!n_n3903) & (!n_n1504) & (!n_n1693) & (x12452x) & (x12454x)) + ((!n_n3903) & (!n_n1504) & (n_n1693) & (!x12452x) & (!x12454x)) + ((!n_n3903) & (!n_n1504) & (n_n1693) & (!x12452x) & (x12454x)) + ((!n_n3903) & (!n_n1504) & (n_n1693) & (x12452x) & (!x12454x)) + ((!n_n3903) & (!n_n1504) & (n_n1693) & (x12452x) & (x12454x)) + ((!n_n3903) & (n_n1504) & (!n_n1693) & (!x12452x) & (!x12454x)) + ((!n_n3903) & (n_n1504) & (!n_n1693) & (!x12452x) & (x12454x)) + ((!n_n3903) & (n_n1504) & (!n_n1693) & (x12452x) & (!x12454x)) + ((!n_n3903) & (n_n1504) & (!n_n1693) & (x12452x) & (x12454x)) + ((!n_n3903) & (n_n1504) & (n_n1693) & (!x12452x) & (!x12454x)) + ((!n_n3903) & (n_n1504) & (n_n1693) & (!x12452x) & (x12454x)) + ((!n_n3903) & (n_n1504) & (n_n1693) & (x12452x) & (!x12454x)) + ((!n_n3903) & (n_n1504) & (n_n1693) & (x12452x) & (x12454x)) + ((n_n3903) & (!n_n1504) & (!n_n1693) & (!x12452x) & (!x12454x)) + ((n_n3903) & (!n_n1504) & (!n_n1693) & (!x12452x) & (x12454x)) + ((n_n3903) & (!n_n1504) & (!n_n1693) & (x12452x) & (!x12454x)) + ((n_n3903) & (!n_n1504) & (!n_n1693) & (x12452x) & (x12454x)) + ((n_n3903) & (!n_n1504) & (n_n1693) & (!x12452x) & (!x12454x)) + ((n_n3903) & (!n_n1504) & (n_n1693) & (!x12452x) & (x12454x)) + ((n_n3903) & (!n_n1504) & (n_n1693) & (x12452x) & (!x12454x)) + ((n_n3903) & (!n_n1504) & (n_n1693) & (x12452x) & (x12454x)) + ((n_n3903) & (n_n1504) & (!n_n1693) & (!x12452x) & (!x12454x)) + ((n_n3903) & (n_n1504) & (!n_n1693) & (!x12452x) & (x12454x)) + ((n_n3903) & (n_n1504) & (!n_n1693) & (x12452x) & (!x12454x)) + ((n_n3903) & (n_n1504) & (!n_n1693) & (x12452x) & (x12454x)) + ((n_n3903) & (n_n1504) & (n_n1693) & (!x12452x) & (!x12454x)) + ((n_n3903) & (n_n1504) & (n_n1693) & (!x12452x) & (x12454x)) + ((n_n3903) & (n_n1504) & (n_n1693) & (x12452x) & (!x12454x)) + ((n_n3903) & (n_n1504) & (n_n1693) & (x12452x) & (x12454x)));
	assign n_n1426 = (((!x83x) & (!x79x) & (!x12460x) & (!x12469x) & (x12468x)) + ((!x83x) & (!x79x) & (!x12460x) & (x12469x) & (!x12468x)) + ((!x83x) & (!x79x) & (!x12460x) & (x12469x) & (x12468x)) + ((!x83x) & (!x79x) & (x12460x) & (!x12469x) & (!x12468x)) + ((!x83x) & (!x79x) & (x12460x) & (!x12469x) & (x12468x)) + ((!x83x) & (!x79x) & (x12460x) & (x12469x) & (!x12468x)) + ((!x83x) & (!x79x) & (x12460x) & (x12469x) & (x12468x)) + ((!x83x) & (x79x) & (!x12460x) & (!x12469x) & (!x12468x)) + ((!x83x) & (x79x) & (!x12460x) & (!x12469x) & (x12468x)) + ((!x83x) & (x79x) & (!x12460x) & (x12469x) & (!x12468x)) + ((!x83x) & (x79x) & (!x12460x) & (x12469x) & (x12468x)) + ((!x83x) & (x79x) & (x12460x) & (!x12469x) & (!x12468x)) + ((!x83x) & (x79x) & (x12460x) & (!x12469x) & (x12468x)) + ((!x83x) & (x79x) & (x12460x) & (x12469x) & (!x12468x)) + ((!x83x) & (x79x) & (x12460x) & (x12469x) & (x12468x)) + ((x83x) & (!x79x) & (!x12460x) & (!x12469x) & (!x12468x)) + ((x83x) & (!x79x) & (!x12460x) & (!x12469x) & (x12468x)) + ((x83x) & (!x79x) & (!x12460x) & (x12469x) & (!x12468x)) + ((x83x) & (!x79x) & (!x12460x) & (x12469x) & (x12468x)) + ((x83x) & (!x79x) & (x12460x) & (!x12469x) & (!x12468x)) + ((x83x) & (!x79x) & (x12460x) & (!x12469x) & (x12468x)) + ((x83x) & (!x79x) & (x12460x) & (x12469x) & (!x12468x)) + ((x83x) & (!x79x) & (x12460x) & (x12469x) & (x12468x)) + ((x83x) & (x79x) & (!x12460x) & (!x12469x) & (!x12468x)) + ((x83x) & (x79x) & (!x12460x) & (!x12469x) & (x12468x)) + ((x83x) & (x79x) & (!x12460x) & (x12469x) & (!x12468x)) + ((x83x) & (x79x) & (!x12460x) & (x12469x) & (x12468x)) + ((x83x) & (x79x) & (x12460x) & (!x12469x) & (!x12468x)) + ((x83x) & (x79x) & (x12460x) & (!x12469x) & (x12468x)) + ((x83x) & (x79x) & (x12460x) & (x12469x) & (!x12468x)) + ((x83x) & (x79x) & (x12460x) & (x12469x) & (x12468x)));
	assign n_n1506 = (((!n_n4344) & (!n_n4341) & (!x67x) & (!x53x) & (x448x)) + ((!n_n4344) & (!n_n4341) & (!x67x) & (x53x) & (!x448x)) + ((!n_n4344) & (!n_n4341) & (!x67x) & (x53x) & (x448x)) + ((!n_n4344) & (!n_n4341) & (x67x) & (!x53x) & (!x448x)) + ((!n_n4344) & (!n_n4341) & (x67x) & (!x53x) & (x448x)) + ((!n_n4344) & (!n_n4341) & (x67x) & (x53x) & (!x448x)) + ((!n_n4344) & (!n_n4341) & (x67x) & (x53x) & (x448x)) + ((!n_n4344) & (n_n4341) & (!x67x) & (!x53x) & (!x448x)) + ((!n_n4344) & (n_n4341) & (!x67x) & (!x53x) & (x448x)) + ((!n_n4344) & (n_n4341) & (!x67x) & (x53x) & (!x448x)) + ((!n_n4344) & (n_n4341) & (!x67x) & (x53x) & (x448x)) + ((!n_n4344) & (n_n4341) & (x67x) & (!x53x) & (!x448x)) + ((!n_n4344) & (n_n4341) & (x67x) & (!x53x) & (x448x)) + ((!n_n4344) & (n_n4341) & (x67x) & (x53x) & (!x448x)) + ((!n_n4344) & (n_n4341) & (x67x) & (x53x) & (x448x)) + ((n_n4344) & (!n_n4341) & (!x67x) & (!x53x) & (!x448x)) + ((n_n4344) & (!n_n4341) & (!x67x) & (!x53x) & (x448x)) + ((n_n4344) & (!n_n4341) & (!x67x) & (x53x) & (!x448x)) + ((n_n4344) & (!n_n4341) & (!x67x) & (x53x) & (x448x)) + ((n_n4344) & (!n_n4341) & (x67x) & (!x53x) & (!x448x)) + ((n_n4344) & (!n_n4341) & (x67x) & (!x53x) & (x448x)) + ((n_n4344) & (!n_n4341) & (x67x) & (x53x) & (!x448x)) + ((n_n4344) & (!n_n4341) & (x67x) & (x53x) & (x448x)) + ((n_n4344) & (n_n4341) & (!x67x) & (!x53x) & (!x448x)) + ((n_n4344) & (n_n4341) & (!x67x) & (!x53x) & (x448x)) + ((n_n4344) & (n_n4341) & (!x67x) & (x53x) & (!x448x)) + ((n_n4344) & (n_n4341) & (!x67x) & (x53x) & (x448x)) + ((n_n4344) & (n_n4341) & (x67x) & (!x53x) & (!x448x)) + ((n_n4344) & (n_n4341) & (x67x) & (!x53x) & (x448x)) + ((n_n4344) & (n_n4341) & (x67x) & (x53x) & (!x448x)) + ((n_n4344) & (n_n4341) & (x67x) & (x53x) & (x448x)));
	assign n_n1508 = (((!n_n4318) & (!n_n4320) & (!x283x) & (!x364x) & (x12575x)) + ((!n_n4318) & (!n_n4320) & (!x283x) & (x364x) & (!x12575x)) + ((!n_n4318) & (!n_n4320) & (!x283x) & (x364x) & (x12575x)) + ((!n_n4318) & (!n_n4320) & (x283x) & (!x364x) & (!x12575x)) + ((!n_n4318) & (!n_n4320) & (x283x) & (!x364x) & (x12575x)) + ((!n_n4318) & (!n_n4320) & (x283x) & (x364x) & (!x12575x)) + ((!n_n4318) & (!n_n4320) & (x283x) & (x364x) & (x12575x)) + ((!n_n4318) & (n_n4320) & (!x283x) & (!x364x) & (!x12575x)) + ((!n_n4318) & (n_n4320) & (!x283x) & (!x364x) & (x12575x)) + ((!n_n4318) & (n_n4320) & (!x283x) & (x364x) & (!x12575x)) + ((!n_n4318) & (n_n4320) & (!x283x) & (x364x) & (x12575x)) + ((!n_n4318) & (n_n4320) & (x283x) & (!x364x) & (!x12575x)) + ((!n_n4318) & (n_n4320) & (x283x) & (!x364x) & (x12575x)) + ((!n_n4318) & (n_n4320) & (x283x) & (x364x) & (!x12575x)) + ((!n_n4318) & (n_n4320) & (x283x) & (x364x) & (x12575x)) + ((n_n4318) & (!n_n4320) & (!x283x) & (!x364x) & (!x12575x)) + ((n_n4318) & (!n_n4320) & (!x283x) & (!x364x) & (x12575x)) + ((n_n4318) & (!n_n4320) & (!x283x) & (x364x) & (!x12575x)) + ((n_n4318) & (!n_n4320) & (!x283x) & (x364x) & (x12575x)) + ((n_n4318) & (!n_n4320) & (x283x) & (!x364x) & (!x12575x)) + ((n_n4318) & (!n_n4320) & (x283x) & (!x364x) & (x12575x)) + ((n_n4318) & (!n_n4320) & (x283x) & (x364x) & (!x12575x)) + ((n_n4318) & (!n_n4320) & (x283x) & (x364x) & (x12575x)) + ((n_n4318) & (n_n4320) & (!x283x) & (!x364x) & (!x12575x)) + ((n_n4318) & (n_n4320) & (!x283x) & (!x364x) & (x12575x)) + ((n_n4318) & (n_n4320) & (!x283x) & (x364x) & (!x12575x)) + ((n_n4318) & (n_n4320) & (!x283x) & (x364x) & (x12575x)) + ((n_n4318) & (n_n4320) & (x283x) & (!x364x) & (!x12575x)) + ((n_n4318) & (n_n4320) & (x283x) & (!x364x) & (x12575x)) + ((n_n4318) & (n_n4320) & (x283x) & (x364x) & (!x12575x)) + ((n_n4318) & (n_n4320) & (x283x) & (x364x) & (x12575x)));
	assign x12581x = (((!n_n4332) & (!n_n4328) & (!x410x) & (!x106x) & (n_n1703)) + ((!n_n4332) & (!n_n4328) & (!x410x) & (x106x) & (!n_n1703)) + ((!n_n4332) & (!n_n4328) & (!x410x) & (x106x) & (n_n1703)) + ((!n_n4332) & (!n_n4328) & (x410x) & (!x106x) & (!n_n1703)) + ((!n_n4332) & (!n_n4328) & (x410x) & (!x106x) & (n_n1703)) + ((!n_n4332) & (!n_n4328) & (x410x) & (x106x) & (!n_n1703)) + ((!n_n4332) & (!n_n4328) & (x410x) & (x106x) & (n_n1703)) + ((!n_n4332) & (n_n4328) & (!x410x) & (!x106x) & (!n_n1703)) + ((!n_n4332) & (n_n4328) & (!x410x) & (!x106x) & (n_n1703)) + ((!n_n4332) & (n_n4328) & (!x410x) & (x106x) & (!n_n1703)) + ((!n_n4332) & (n_n4328) & (!x410x) & (x106x) & (n_n1703)) + ((!n_n4332) & (n_n4328) & (x410x) & (!x106x) & (!n_n1703)) + ((!n_n4332) & (n_n4328) & (x410x) & (!x106x) & (n_n1703)) + ((!n_n4332) & (n_n4328) & (x410x) & (x106x) & (!n_n1703)) + ((!n_n4332) & (n_n4328) & (x410x) & (x106x) & (n_n1703)) + ((n_n4332) & (!n_n4328) & (!x410x) & (!x106x) & (!n_n1703)) + ((n_n4332) & (!n_n4328) & (!x410x) & (!x106x) & (n_n1703)) + ((n_n4332) & (!n_n4328) & (!x410x) & (x106x) & (!n_n1703)) + ((n_n4332) & (!n_n4328) & (!x410x) & (x106x) & (n_n1703)) + ((n_n4332) & (!n_n4328) & (x410x) & (!x106x) & (!n_n1703)) + ((n_n4332) & (!n_n4328) & (x410x) & (!x106x) & (n_n1703)) + ((n_n4332) & (!n_n4328) & (x410x) & (x106x) & (!n_n1703)) + ((n_n4332) & (!n_n4328) & (x410x) & (x106x) & (n_n1703)) + ((n_n4332) & (n_n4328) & (!x410x) & (!x106x) & (!n_n1703)) + ((n_n4332) & (n_n4328) & (!x410x) & (!x106x) & (n_n1703)) + ((n_n4332) & (n_n4328) & (!x410x) & (x106x) & (!n_n1703)) + ((n_n4332) & (n_n4328) & (!x410x) & (x106x) & (n_n1703)) + ((n_n4332) & (n_n4328) & (x410x) & (!x106x) & (!n_n1703)) + ((n_n4332) & (n_n4328) & (x410x) & (!x106x) & (n_n1703)) + ((n_n4332) & (n_n4328) & (x410x) & (x106x) & (!n_n1703)) + ((n_n4332) & (n_n4328) & (x410x) & (x106x) & (n_n1703)));
	assign x12585x = (((!n_n1427) & (!n_n1426) & (!n_n1506) & (!n_n1508) & (x12581x)) + ((!n_n1427) & (!n_n1426) & (!n_n1506) & (n_n1508) & (!x12581x)) + ((!n_n1427) & (!n_n1426) & (!n_n1506) & (n_n1508) & (x12581x)) + ((!n_n1427) & (!n_n1426) & (n_n1506) & (!n_n1508) & (!x12581x)) + ((!n_n1427) & (!n_n1426) & (n_n1506) & (!n_n1508) & (x12581x)) + ((!n_n1427) & (!n_n1426) & (n_n1506) & (n_n1508) & (!x12581x)) + ((!n_n1427) & (!n_n1426) & (n_n1506) & (n_n1508) & (x12581x)) + ((!n_n1427) & (n_n1426) & (!n_n1506) & (!n_n1508) & (!x12581x)) + ((!n_n1427) & (n_n1426) & (!n_n1506) & (!n_n1508) & (x12581x)) + ((!n_n1427) & (n_n1426) & (!n_n1506) & (n_n1508) & (!x12581x)) + ((!n_n1427) & (n_n1426) & (!n_n1506) & (n_n1508) & (x12581x)) + ((!n_n1427) & (n_n1426) & (n_n1506) & (!n_n1508) & (!x12581x)) + ((!n_n1427) & (n_n1426) & (n_n1506) & (!n_n1508) & (x12581x)) + ((!n_n1427) & (n_n1426) & (n_n1506) & (n_n1508) & (!x12581x)) + ((!n_n1427) & (n_n1426) & (n_n1506) & (n_n1508) & (x12581x)) + ((n_n1427) & (!n_n1426) & (!n_n1506) & (!n_n1508) & (!x12581x)) + ((n_n1427) & (!n_n1426) & (!n_n1506) & (!n_n1508) & (x12581x)) + ((n_n1427) & (!n_n1426) & (!n_n1506) & (n_n1508) & (!x12581x)) + ((n_n1427) & (!n_n1426) & (!n_n1506) & (n_n1508) & (x12581x)) + ((n_n1427) & (!n_n1426) & (n_n1506) & (!n_n1508) & (!x12581x)) + ((n_n1427) & (!n_n1426) & (n_n1506) & (!n_n1508) & (x12581x)) + ((n_n1427) & (!n_n1426) & (n_n1506) & (n_n1508) & (!x12581x)) + ((n_n1427) & (!n_n1426) & (n_n1506) & (n_n1508) & (x12581x)) + ((n_n1427) & (n_n1426) & (!n_n1506) & (!n_n1508) & (!x12581x)) + ((n_n1427) & (n_n1426) & (!n_n1506) & (!n_n1508) & (x12581x)) + ((n_n1427) & (n_n1426) & (!n_n1506) & (n_n1508) & (!x12581x)) + ((n_n1427) & (n_n1426) & (!n_n1506) & (n_n1508) & (x12581x)) + ((n_n1427) & (n_n1426) & (n_n1506) & (!n_n1508) & (!x12581x)) + ((n_n1427) & (n_n1426) & (n_n1506) & (!n_n1508) & (x12581x)) + ((n_n1427) & (n_n1426) & (n_n1506) & (n_n1508) & (!x12581x)) + ((n_n1427) & (n_n1426) & (n_n1506) & (n_n1508) & (x12581x)));
	assign n_n1425 = (((!x12476x) & (!x12485x) & (!x12481x) & (!x22141x)) + ((!x12476x) & (!x12485x) & (x12481x) & (!x22141x)) + ((!x12476x) & (!x12485x) & (x12481x) & (x22141x)) + ((!x12476x) & (x12485x) & (!x12481x) & (!x22141x)) + ((!x12476x) & (x12485x) & (!x12481x) & (x22141x)) + ((!x12476x) & (x12485x) & (x12481x) & (!x22141x)) + ((!x12476x) & (x12485x) & (x12481x) & (x22141x)) + ((x12476x) & (!x12485x) & (!x12481x) & (!x22141x)) + ((x12476x) & (!x12485x) & (!x12481x) & (x22141x)) + ((x12476x) & (!x12485x) & (x12481x) & (!x22141x)) + ((x12476x) & (!x12485x) & (x12481x) & (x22141x)) + ((x12476x) & (x12485x) & (!x12481x) & (!x22141x)) + ((x12476x) & (x12485x) & (!x12481x) & (x22141x)) + ((x12476x) & (x12485x) & (x12481x) & (!x22141x)) + ((x12476x) & (x12485x) & (x12481x) & (x22141x)));
	assign n_n1423 = (((!n_n1491) & (!x12504x) & (!x12505x) & (x12506x)) + ((!n_n1491) & (!x12504x) & (x12505x) & (!x12506x)) + ((!n_n1491) & (!x12504x) & (x12505x) & (x12506x)) + ((!n_n1491) & (x12504x) & (!x12505x) & (!x12506x)) + ((!n_n1491) & (x12504x) & (!x12505x) & (x12506x)) + ((!n_n1491) & (x12504x) & (x12505x) & (!x12506x)) + ((!n_n1491) & (x12504x) & (x12505x) & (x12506x)) + ((n_n1491) & (!x12504x) & (!x12505x) & (!x12506x)) + ((n_n1491) & (!x12504x) & (!x12505x) & (x12506x)) + ((n_n1491) & (!x12504x) & (x12505x) & (!x12506x)) + ((n_n1491) & (!x12504x) & (x12505x) & (x12506x)) + ((n_n1491) & (x12504x) & (!x12505x) & (!x12506x)) + ((n_n1491) & (x12504x) & (!x12505x) & (x12506x)) + ((n_n1491) & (x12504x) & (x12505x) & (!x12506x)) + ((n_n1491) & (x12504x) & (x12505x) & (x12506x)));
	assign x12517x = (((!n_n1496) & (!x12513x) & (!x12514x) & (!x22140x)) + ((!n_n1496) & (!x12513x) & (x12514x) & (!x22140x)) + ((!n_n1496) & (!x12513x) & (x12514x) & (x22140x)) + ((!n_n1496) & (x12513x) & (!x12514x) & (!x22140x)) + ((!n_n1496) & (x12513x) & (!x12514x) & (x22140x)) + ((!n_n1496) & (x12513x) & (x12514x) & (!x22140x)) + ((!n_n1496) & (x12513x) & (x12514x) & (x22140x)) + ((n_n1496) & (!x12513x) & (!x12514x) & (!x22140x)) + ((n_n1496) & (!x12513x) & (!x12514x) & (x22140x)) + ((n_n1496) & (!x12513x) & (x12514x) & (!x22140x)) + ((n_n1496) & (!x12513x) & (x12514x) & (x22140x)) + ((n_n1496) & (x12513x) & (!x12514x) & (!x22140x)) + ((n_n1496) & (x12513x) & (!x12514x) & (x22140x)) + ((n_n1496) & (x12513x) & (x12514x) & (!x22140x)) + ((n_n1496) & (x12513x) & (x12514x) & (x22140x)));
	assign n_n1399 = (((!n_n1422) & (!n_n1485) & (!n_n1487) & (!n_n1420) & (x12565x)) + ((!n_n1422) & (!n_n1485) & (!n_n1487) & (n_n1420) & (!x12565x)) + ((!n_n1422) & (!n_n1485) & (!n_n1487) & (n_n1420) & (x12565x)) + ((!n_n1422) & (!n_n1485) & (n_n1487) & (!n_n1420) & (!x12565x)) + ((!n_n1422) & (!n_n1485) & (n_n1487) & (!n_n1420) & (x12565x)) + ((!n_n1422) & (!n_n1485) & (n_n1487) & (n_n1420) & (!x12565x)) + ((!n_n1422) & (!n_n1485) & (n_n1487) & (n_n1420) & (x12565x)) + ((!n_n1422) & (n_n1485) & (!n_n1487) & (!n_n1420) & (!x12565x)) + ((!n_n1422) & (n_n1485) & (!n_n1487) & (!n_n1420) & (x12565x)) + ((!n_n1422) & (n_n1485) & (!n_n1487) & (n_n1420) & (!x12565x)) + ((!n_n1422) & (n_n1485) & (!n_n1487) & (n_n1420) & (x12565x)) + ((!n_n1422) & (n_n1485) & (n_n1487) & (!n_n1420) & (!x12565x)) + ((!n_n1422) & (n_n1485) & (n_n1487) & (!n_n1420) & (x12565x)) + ((!n_n1422) & (n_n1485) & (n_n1487) & (n_n1420) & (!x12565x)) + ((!n_n1422) & (n_n1485) & (n_n1487) & (n_n1420) & (x12565x)) + ((n_n1422) & (!n_n1485) & (!n_n1487) & (!n_n1420) & (!x12565x)) + ((n_n1422) & (!n_n1485) & (!n_n1487) & (!n_n1420) & (x12565x)) + ((n_n1422) & (!n_n1485) & (!n_n1487) & (n_n1420) & (!x12565x)) + ((n_n1422) & (!n_n1485) & (!n_n1487) & (n_n1420) & (x12565x)) + ((n_n1422) & (!n_n1485) & (n_n1487) & (!n_n1420) & (!x12565x)) + ((n_n1422) & (!n_n1485) & (n_n1487) & (!n_n1420) & (x12565x)) + ((n_n1422) & (!n_n1485) & (n_n1487) & (n_n1420) & (!x12565x)) + ((n_n1422) & (!n_n1485) & (n_n1487) & (n_n1420) & (x12565x)) + ((n_n1422) & (n_n1485) & (!n_n1487) & (!n_n1420) & (!x12565x)) + ((n_n1422) & (n_n1485) & (!n_n1487) & (!n_n1420) & (x12565x)) + ((n_n1422) & (n_n1485) & (!n_n1487) & (n_n1420) & (!x12565x)) + ((n_n1422) & (n_n1485) & (!n_n1487) & (n_n1420) & (x12565x)) + ((n_n1422) & (n_n1485) & (n_n1487) & (!n_n1420) & (!x12565x)) + ((n_n1422) & (n_n1485) & (n_n1487) & (!n_n1420) & (x12565x)) + ((n_n1422) & (n_n1485) & (n_n1487) & (n_n1420) & (!x12565x)) + ((n_n1422) & (n_n1485) & (n_n1487) & (n_n1420) & (x12565x)));
	assign x25x = (((!i_9_) & (i_7_) & (i_8_) & (i_6_)));
	assign n_n473 = (((i_5_) & (!i_3_) & (!i_4_)));
	assign n_n534 = (((i_7_) & (i_8_) & (i_6_)));
	assign n_n65 = (((!i_1_) & (!i_2_) & (!i_0_)));
	assign n_n5305 = (((!i_9_) & (n_n473) & (n_n534) & (n_n65)));
	assign x15x = (((!i_9_) & (!i_7_) & (i_8_) & (i_6_)));
	assign x592x = (((!i_5_) & (!i_3_) & (i_4_) & (n_n65)));
	assign n_n482 = (((!i_5_) & (!i_3_) & (i_4_)));
	assign n_n530 = (((!i_7_) & (i_8_) & (i_6_)));
	assign n_n5293 = (((!i_9_) & (n_n482) & (n_n530) & (n_n65)));
	assign x19x = (((i_9_) & (!i_1_) & (!i_2_) & (!i_0_)));
	assign n_n5296 = (((i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n482)));
	assign n_n491 = (((i_5_) & (!i_3_) & (i_4_)));
	assign x492x = (((!i_7_) & (i_8_) & (!i_6_) & (n_n491)));
	assign n_n5284 = (((!i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n491)));
	assign n_n559 = (((!n_n4578) & (!n_n4611) & (!n_n4633) & (!n_n4581) & (x12597x)) + ((!n_n4578) & (!n_n4611) & (!n_n4633) & (n_n4581) & (!x12597x)) + ((!n_n4578) & (!n_n4611) & (!n_n4633) & (n_n4581) & (x12597x)) + ((!n_n4578) & (!n_n4611) & (n_n4633) & (!n_n4581) & (!x12597x)) + ((!n_n4578) & (!n_n4611) & (n_n4633) & (!n_n4581) & (x12597x)) + ((!n_n4578) & (!n_n4611) & (n_n4633) & (n_n4581) & (!x12597x)) + ((!n_n4578) & (!n_n4611) & (n_n4633) & (n_n4581) & (x12597x)) + ((!n_n4578) & (n_n4611) & (!n_n4633) & (!n_n4581) & (!x12597x)) + ((!n_n4578) & (n_n4611) & (!n_n4633) & (!n_n4581) & (x12597x)) + ((!n_n4578) & (n_n4611) & (!n_n4633) & (n_n4581) & (!x12597x)) + ((!n_n4578) & (n_n4611) & (!n_n4633) & (n_n4581) & (x12597x)) + ((!n_n4578) & (n_n4611) & (n_n4633) & (!n_n4581) & (!x12597x)) + ((!n_n4578) & (n_n4611) & (n_n4633) & (!n_n4581) & (x12597x)) + ((!n_n4578) & (n_n4611) & (n_n4633) & (n_n4581) & (!x12597x)) + ((!n_n4578) & (n_n4611) & (n_n4633) & (n_n4581) & (x12597x)) + ((n_n4578) & (!n_n4611) & (!n_n4633) & (!n_n4581) & (!x12597x)) + ((n_n4578) & (!n_n4611) & (!n_n4633) & (!n_n4581) & (x12597x)) + ((n_n4578) & (!n_n4611) & (!n_n4633) & (n_n4581) & (!x12597x)) + ((n_n4578) & (!n_n4611) & (!n_n4633) & (n_n4581) & (x12597x)) + ((n_n4578) & (!n_n4611) & (n_n4633) & (!n_n4581) & (!x12597x)) + ((n_n4578) & (!n_n4611) & (n_n4633) & (!n_n4581) & (x12597x)) + ((n_n4578) & (!n_n4611) & (n_n4633) & (n_n4581) & (!x12597x)) + ((n_n4578) & (!n_n4611) & (n_n4633) & (n_n4581) & (x12597x)) + ((n_n4578) & (n_n4611) & (!n_n4633) & (!n_n4581) & (!x12597x)) + ((n_n4578) & (n_n4611) & (!n_n4633) & (!n_n4581) & (x12597x)) + ((n_n4578) & (n_n4611) & (!n_n4633) & (n_n4581) & (!x12597x)) + ((n_n4578) & (n_n4611) & (!n_n4633) & (n_n4581) & (x12597x)) + ((n_n4578) & (n_n4611) & (n_n4633) & (!n_n4581) & (!x12597x)) + ((n_n4578) & (n_n4611) & (n_n4633) & (!n_n4581) & (x12597x)) + ((n_n4578) & (n_n4611) & (n_n4633) & (n_n4581) & (!x12597x)) + ((n_n4578) & (n_n4611) & (n_n4633) & (n_n4581) & (x12597x)));
	assign x12600x = (((!n_n4641) & (!n_n4643) & (!n_n4646) & (n_n4647)) + ((!n_n4641) & (!n_n4643) & (n_n4646) & (!n_n4647)) + ((!n_n4641) & (!n_n4643) & (n_n4646) & (n_n4647)) + ((!n_n4641) & (n_n4643) & (!n_n4646) & (!n_n4647)) + ((!n_n4641) & (n_n4643) & (!n_n4646) & (n_n4647)) + ((!n_n4641) & (n_n4643) & (n_n4646) & (!n_n4647)) + ((!n_n4641) & (n_n4643) & (n_n4646) & (n_n4647)) + ((n_n4641) & (!n_n4643) & (!n_n4646) & (!n_n4647)) + ((n_n4641) & (!n_n4643) & (!n_n4646) & (n_n4647)) + ((n_n4641) & (!n_n4643) & (n_n4646) & (!n_n4647)) + ((n_n4641) & (!n_n4643) & (n_n4646) & (n_n4647)) + ((n_n4641) & (n_n4643) & (!n_n4646) & (!n_n4647)) + ((n_n4641) & (n_n4643) & (!n_n4646) & (n_n4647)) + ((n_n4641) & (n_n4643) & (n_n4646) & (!n_n4647)) + ((n_n4641) & (n_n4643) & (n_n4646) & (n_n4647)));
	assign x12601x = (((!n_n4648) & (!n_n4645) & (!n_n4635) & (x140x)) + ((!n_n4648) & (!n_n4645) & (n_n4635) & (!x140x)) + ((!n_n4648) & (!n_n4645) & (n_n4635) & (x140x)) + ((!n_n4648) & (n_n4645) & (!n_n4635) & (!x140x)) + ((!n_n4648) & (n_n4645) & (!n_n4635) & (x140x)) + ((!n_n4648) & (n_n4645) & (n_n4635) & (!x140x)) + ((!n_n4648) & (n_n4645) & (n_n4635) & (x140x)) + ((n_n4648) & (!n_n4645) & (!n_n4635) & (!x140x)) + ((n_n4648) & (!n_n4645) & (!n_n4635) & (x140x)) + ((n_n4648) & (!n_n4645) & (n_n4635) & (!x140x)) + ((n_n4648) & (!n_n4645) & (n_n4635) & (x140x)) + ((n_n4648) & (n_n4645) & (!n_n4635) & (!x140x)) + ((n_n4648) & (n_n4645) & (!n_n4635) & (x140x)) + ((n_n4648) & (n_n4645) & (n_n4635) & (!x140x)) + ((n_n4648) & (n_n4645) & (n_n4635) & (x140x)));
	assign x12607x = (((!n_n4557) & (!n_n4572) & (!n_n4531) & (n_n4555)) + ((!n_n4557) & (!n_n4572) & (n_n4531) & (!n_n4555)) + ((!n_n4557) & (!n_n4572) & (n_n4531) & (n_n4555)) + ((!n_n4557) & (n_n4572) & (!n_n4531) & (!n_n4555)) + ((!n_n4557) & (n_n4572) & (!n_n4531) & (n_n4555)) + ((!n_n4557) & (n_n4572) & (n_n4531) & (!n_n4555)) + ((!n_n4557) & (n_n4572) & (n_n4531) & (n_n4555)) + ((n_n4557) & (!n_n4572) & (!n_n4531) & (!n_n4555)) + ((n_n4557) & (!n_n4572) & (!n_n4531) & (n_n4555)) + ((n_n4557) & (!n_n4572) & (n_n4531) & (!n_n4555)) + ((n_n4557) & (!n_n4572) & (n_n4531) & (n_n4555)) + ((n_n4557) & (n_n4572) & (!n_n4531) & (!n_n4555)) + ((n_n4557) & (n_n4572) & (!n_n4531) & (n_n4555)) + ((n_n4557) & (n_n4572) & (n_n4531) & (!n_n4555)) + ((n_n4557) & (n_n4572) & (n_n4531) & (n_n4555)));
	assign x12608x = (((!n_n4523) & (!n_n4539) & (!n_n4549) & (!n_n4559) & (n_n4528)) + ((!n_n4523) & (!n_n4539) & (!n_n4549) & (n_n4559) & (!n_n4528)) + ((!n_n4523) & (!n_n4539) & (!n_n4549) & (n_n4559) & (n_n4528)) + ((!n_n4523) & (!n_n4539) & (n_n4549) & (!n_n4559) & (!n_n4528)) + ((!n_n4523) & (!n_n4539) & (n_n4549) & (!n_n4559) & (n_n4528)) + ((!n_n4523) & (!n_n4539) & (n_n4549) & (n_n4559) & (!n_n4528)) + ((!n_n4523) & (!n_n4539) & (n_n4549) & (n_n4559) & (n_n4528)) + ((!n_n4523) & (n_n4539) & (!n_n4549) & (!n_n4559) & (!n_n4528)) + ((!n_n4523) & (n_n4539) & (!n_n4549) & (!n_n4559) & (n_n4528)) + ((!n_n4523) & (n_n4539) & (!n_n4549) & (n_n4559) & (!n_n4528)) + ((!n_n4523) & (n_n4539) & (!n_n4549) & (n_n4559) & (n_n4528)) + ((!n_n4523) & (n_n4539) & (n_n4549) & (!n_n4559) & (!n_n4528)) + ((!n_n4523) & (n_n4539) & (n_n4549) & (!n_n4559) & (n_n4528)) + ((!n_n4523) & (n_n4539) & (n_n4549) & (n_n4559) & (!n_n4528)) + ((!n_n4523) & (n_n4539) & (n_n4549) & (n_n4559) & (n_n4528)) + ((n_n4523) & (!n_n4539) & (!n_n4549) & (!n_n4559) & (!n_n4528)) + ((n_n4523) & (!n_n4539) & (!n_n4549) & (!n_n4559) & (n_n4528)) + ((n_n4523) & (!n_n4539) & (!n_n4549) & (n_n4559) & (!n_n4528)) + ((n_n4523) & (!n_n4539) & (!n_n4549) & (n_n4559) & (n_n4528)) + ((n_n4523) & (!n_n4539) & (n_n4549) & (!n_n4559) & (!n_n4528)) + ((n_n4523) & (!n_n4539) & (n_n4549) & (!n_n4559) & (n_n4528)) + ((n_n4523) & (!n_n4539) & (n_n4549) & (n_n4559) & (!n_n4528)) + ((n_n4523) & (!n_n4539) & (n_n4549) & (n_n4559) & (n_n4528)) + ((n_n4523) & (n_n4539) & (!n_n4549) & (!n_n4559) & (!n_n4528)) + ((n_n4523) & (n_n4539) & (!n_n4549) & (!n_n4559) & (n_n4528)) + ((n_n4523) & (n_n4539) & (!n_n4549) & (n_n4559) & (!n_n4528)) + ((n_n4523) & (n_n4539) & (!n_n4549) & (n_n4559) & (n_n4528)) + ((n_n4523) & (n_n4539) & (n_n4549) & (!n_n4559) & (!n_n4528)) + ((n_n4523) & (n_n4539) & (n_n4549) & (!n_n4559) & (n_n4528)) + ((n_n4523) & (n_n4539) & (n_n4549) & (n_n4559) & (!n_n4528)) + ((n_n4523) & (n_n4539) & (n_n4549) & (n_n4559) & (n_n4528)));
	assign n_n543 = (((!n_n559) & (!x12600x) & (!x12601x) & (!x12607x) & (x12608x)) + ((!n_n559) & (!x12600x) & (!x12601x) & (x12607x) & (!x12608x)) + ((!n_n559) & (!x12600x) & (!x12601x) & (x12607x) & (x12608x)) + ((!n_n559) & (!x12600x) & (x12601x) & (!x12607x) & (!x12608x)) + ((!n_n559) & (!x12600x) & (x12601x) & (!x12607x) & (x12608x)) + ((!n_n559) & (!x12600x) & (x12601x) & (x12607x) & (!x12608x)) + ((!n_n559) & (!x12600x) & (x12601x) & (x12607x) & (x12608x)) + ((!n_n559) & (x12600x) & (!x12601x) & (!x12607x) & (!x12608x)) + ((!n_n559) & (x12600x) & (!x12601x) & (!x12607x) & (x12608x)) + ((!n_n559) & (x12600x) & (!x12601x) & (x12607x) & (!x12608x)) + ((!n_n559) & (x12600x) & (!x12601x) & (x12607x) & (x12608x)) + ((!n_n559) & (x12600x) & (x12601x) & (!x12607x) & (!x12608x)) + ((!n_n559) & (x12600x) & (x12601x) & (!x12607x) & (x12608x)) + ((!n_n559) & (x12600x) & (x12601x) & (x12607x) & (!x12608x)) + ((!n_n559) & (x12600x) & (x12601x) & (x12607x) & (x12608x)) + ((n_n559) & (!x12600x) & (!x12601x) & (!x12607x) & (!x12608x)) + ((n_n559) & (!x12600x) & (!x12601x) & (!x12607x) & (x12608x)) + ((n_n559) & (!x12600x) & (!x12601x) & (x12607x) & (!x12608x)) + ((n_n559) & (!x12600x) & (!x12601x) & (x12607x) & (x12608x)) + ((n_n559) & (!x12600x) & (x12601x) & (!x12607x) & (!x12608x)) + ((n_n559) & (!x12600x) & (x12601x) & (!x12607x) & (x12608x)) + ((n_n559) & (!x12600x) & (x12601x) & (x12607x) & (!x12608x)) + ((n_n559) & (!x12600x) & (x12601x) & (x12607x) & (x12608x)) + ((n_n559) & (x12600x) & (!x12601x) & (!x12607x) & (!x12608x)) + ((n_n559) & (x12600x) & (!x12601x) & (!x12607x) & (x12608x)) + ((n_n559) & (x12600x) & (!x12601x) & (x12607x) & (!x12608x)) + ((n_n559) & (x12600x) & (!x12601x) & (x12607x) & (x12608x)) + ((n_n559) & (x12600x) & (x12601x) & (!x12607x) & (!x12608x)) + ((n_n559) & (x12600x) & (x12601x) & (!x12607x) & (x12608x)) + ((n_n559) & (x12600x) & (x12601x) & (x12607x) & (!x12608x)) + ((n_n559) & (x12600x) & (x12601x) & (x12607x) & (x12608x)));
	assign n_n4718 = (((i_9_) & (n_n518) & (n_n528) & (n_n325)));
	assign n_n4727 = (((!i_5_) & (i_3_) & (i_4_) & (n_n325) & (x23x)));
	assign n_n4730 = (((i_9_) & (n_n532) & (n_n509) & (n_n325)));
	assign n_n4733 = (((!i_9_) & (n_n509) & (n_n325) & (n_n530)));
	assign x12628x = (((!n_n4735) & (!n_n4749) & (!n_n4750) & (!n_n4740) & (n_n4736)) + ((!n_n4735) & (!n_n4749) & (!n_n4750) & (n_n4740) & (!n_n4736)) + ((!n_n4735) & (!n_n4749) & (!n_n4750) & (n_n4740) & (n_n4736)) + ((!n_n4735) & (!n_n4749) & (n_n4750) & (!n_n4740) & (!n_n4736)) + ((!n_n4735) & (!n_n4749) & (n_n4750) & (!n_n4740) & (n_n4736)) + ((!n_n4735) & (!n_n4749) & (n_n4750) & (n_n4740) & (!n_n4736)) + ((!n_n4735) & (!n_n4749) & (n_n4750) & (n_n4740) & (n_n4736)) + ((!n_n4735) & (n_n4749) & (!n_n4750) & (!n_n4740) & (!n_n4736)) + ((!n_n4735) & (n_n4749) & (!n_n4750) & (!n_n4740) & (n_n4736)) + ((!n_n4735) & (n_n4749) & (!n_n4750) & (n_n4740) & (!n_n4736)) + ((!n_n4735) & (n_n4749) & (!n_n4750) & (n_n4740) & (n_n4736)) + ((!n_n4735) & (n_n4749) & (n_n4750) & (!n_n4740) & (!n_n4736)) + ((!n_n4735) & (n_n4749) & (n_n4750) & (!n_n4740) & (n_n4736)) + ((!n_n4735) & (n_n4749) & (n_n4750) & (n_n4740) & (!n_n4736)) + ((!n_n4735) & (n_n4749) & (n_n4750) & (n_n4740) & (n_n4736)) + ((n_n4735) & (!n_n4749) & (!n_n4750) & (!n_n4740) & (!n_n4736)) + ((n_n4735) & (!n_n4749) & (!n_n4750) & (!n_n4740) & (n_n4736)) + ((n_n4735) & (!n_n4749) & (!n_n4750) & (n_n4740) & (!n_n4736)) + ((n_n4735) & (!n_n4749) & (!n_n4750) & (n_n4740) & (n_n4736)) + ((n_n4735) & (!n_n4749) & (n_n4750) & (!n_n4740) & (!n_n4736)) + ((n_n4735) & (!n_n4749) & (n_n4750) & (!n_n4740) & (n_n4736)) + ((n_n4735) & (!n_n4749) & (n_n4750) & (n_n4740) & (!n_n4736)) + ((n_n4735) & (!n_n4749) & (n_n4750) & (n_n4740) & (n_n4736)) + ((n_n4735) & (n_n4749) & (!n_n4750) & (!n_n4740) & (!n_n4736)) + ((n_n4735) & (n_n4749) & (!n_n4750) & (!n_n4740) & (n_n4736)) + ((n_n4735) & (n_n4749) & (!n_n4750) & (n_n4740) & (!n_n4736)) + ((n_n4735) & (n_n4749) & (!n_n4750) & (n_n4740) & (n_n4736)) + ((n_n4735) & (n_n4749) & (n_n4750) & (!n_n4740) & (!n_n4736)) + ((n_n4735) & (n_n4749) & (n_n4750) & (!n_n4740) & (n_n4736)) + ((n_n4735) & (n_n4749) & (n_n4750) & (n_n4740) & (!n_n4736)) + ((n_n4735) & (n_n4749) & (n_n4750) & (n_n4740) & (n_n4736)));
	assign x12629x = (((!n_n4718) & (!n_n4727) & (!n_n4730) & (!n_n4733) & (x12628x)) + ((!n_n4718) & (!n_n4727) & (!n_n4730) & (n_n4733) & (!x12628x)) + ((!n_n4718) & (!n_n4727) & (!n_n4730) & (n_n4733) & (x12628x)) + ((!n_n4718) & (!n_n4727) & (n_n4730) & (!n_n4733) & (!x12628x)) + ((!n_n4718) & (!n_n4727) & (n_n4730) & (!n_n4733) & (x12628x)) + ((!n_n4718) & (!n_n4727) & (n_n4730) & (n_n4733) & (!x12628x)) + ((!n_n4718) & (!n_n4727) & (n_n4730) & (n_n4733) & (x12628x)) + ((!n_n4718) & (n_n4727) & (!n_n4730) & (!n_n4733) & (!x12628x)) + ((!n_n4718) & (n_n4727) & (!n_n4730) & (!n_n4733) & (x12628x)) + ((!n_n4718) & (n_n4727) & (!n_n4730) & (n_n4733) & (!x12628x)) + ((!n_n4718) & (n_n4727) & (!n_n4730) & (n_n4733) & (x12628x)) + ((!n_n4718) & (n_n4727) & (n_n4730) & (!n_n4733) & (!x12628x)) + ((!n_n4718) & (n_n4727) & (n_n4730) & (!n_n4733) & (x12628x)) + ((!n_n4718) & (n_n4727) & (n_n4730) & (n_n4733) & (!x12628x)) + ((!n_n4718) & (n_n4727) & (n_n4730) & (n_n4733) & (x12628x)) + ((n_n4718) & (!n_n4727) & (!n_n4730) & (!n_n4733) & (!x12628x)) + ((n_n4718) & (!n_n4727) & (!n_n4730) & (!n_n4733) & (x12628x)) + ((n_n4718) & (!n_n4727) & (!n_n4730) & (n_n4733) & (!x12628x)) + ((n_n4718) & (!n_n4727) & (!n_n4730) & (n_n4733) & (x12628x)) + ((n_n4718) & (!n_n4727) & (n_n4730) & (!n_n4733) & (!x12628x)) + ((n_n4718) & (!n_n4727) & (n_n4730) & (!n_n4733) & (x12628x)) + ((n_n4718) & (!n_n4727) & (n_n4730) & (n_n4733) & (!x12628x)) + ((n_n4718) & (!n_n4727) & (n_n4730) & (n_n4733) & (x12628x)) + ((n_n4718) & (n_n4727) & (!n_n4730) & (!n_n4733) & (!x12628x)) + ((n_n4718) & (n_n4727) & (!n_n4730) & (!n_n4733) & (x12628x)) + ((n_n4718) & (n_n4727) & (!n_n4730) & (n_n4733) & (!x12628x)) + ((n_n4718) & (n_n4727) & (!n_n4730) & (n_n4733) & (x12628x)) + ((n_n4718) & (n_n4727) & (n_n4730) & (!n_n4733) & (!x12628x)) + ((n_n4718) & (n_n4727) & (n_n4730) & (!n_n4733) & (x12628x)) + ((n_n4718) & (n_n4727) & (n_n4730) & (n_n4733) & (!x12628x)) + ((n_n4718) & (n_n4727) & (n_n4730) & (n_n4733) & (x12628x)));
	assign x165x = (((!i_9_) & (!n_n528) & (n_n325) & (n_n491) & (n_n530)) + ((!i_9_) & (n_n528) & (n_n325) & (n_n491) & (n_n530)) + ((i_9_) & (n_n528) & (n_n325) & (n_n491) & (!n_n530)) + ((i_9_) & (n_n528) & (n_n325) & (n_n491) & (n_n530)));
	assign x258x = (((!i_9_) & (n_n526) & (n_n325) & (!n_n522) & (n_n500)) + ((!i_9_) & (n_n526) & (n_n325) & (n_n522) & (n_n500)) + ((i_9_) & (!n_n526) & (n_n325) & (n_n522) & (n_n500)) + ((i_9_) & (n_n526) & (n_n325) & (n_n522) & (n_n500)));
	assign x12614x = (((!x131x) & (!n_n4792) & (!n_n4764) & (n_n4763)) + ((!x131x) & (!n_n4792) & (n_n4764) & (!n_n4763)) + ((!x131x) & (!n_n4792) & (n_n4764) & (n_n4763)) + ((!x131x) & (n_n4792) & (!n_n4764) & (!n_n4763)) + ((!x131x) & (n_n4792) & (!n_n4764) & (n_n4763)) + ((!x131x) & (n_n4792) & (n_n4764) & (!n_n4763)) + ((!x131x) & (n_n4792) & (n_n4764) & (n_n4763)) + ((x131x) & (!n_n4792) & (!n_n4764) & (!n_n4763)) + ((x131x) & (!n_n4792) & (!n_n4764) & (n_n4763)) + ((x131x) & (!n_n4792) & (n_n4764) & (!n_n4763)) + ((x131x) & (!n_n4792) & (n_n4764) & (n_n4763)) + ((x131x) & (n_n4792) & (!n_n4764) & (!n_n4763)) + ((x131x) & (n_n4792) & (!n_n4764) & (n_n4763)) + ((x131x) & (n_n4792) & (n_n4764) & (!n_n4763)) + ((x131x) & (n_n4792) & (n_n4764) & (n_n4763)));
	assign n_n557 = (((!n_n4656) & (!n_n4676) & (!n_n4703) & (!n_n4698) & (x12621x)) + ((!n_n4656) & (!n_n4676) & (!n_n4703) & (n_n4698) & (!x12621x)) + ((!n_n4656) & (!n_n4676) & (!n_n4703) & (n_n4698) & (x12621x)) + ((!n_n4656) & (!n_n4676) & (n_n4703) & (!n_n4698) & (!x12621x)) + ((!n_n4656) & (!n_n4676) & (n_n4703) & (!n_n4698) & (x12621x)) + ((!n_n4656) & (!n_n4676) & (n_n4703) & (n_n4698) & (!x12621x)) + ((!n_n4656) & (!n_n4676) & (n_n4703) & (n_n4698) & (x12621x)) + ((!n_n4656) & (n_n4676) & (!n_n4703) & (!n_n4698) & (!x12621x)) + ((!n_n4656) & (n_n4676) & (!n_n4703) & (!n_n4698) & (x12621x)) + ((!n_n4656) & (n_n4676) & (!n_n4703) & (n_n4698) & (!x12621x)) + ((!n_n4656) & (n_n4676) & (!n_n4703) & (n_n4698) & (x12621x)) + ((!n_n4656) & (n_n4676) & (n_n4703) & (!n_n4698) & (!x12621x)) + ((!n_n4656) & (n_n4676) & (n_n4703) & (!n_n4698) & (x12621x)) + ((!n_n4656) & (n_n4676) & (n_n4703) & (n_n4698) & (!x12621x)) + ((!n_n4656) & (n_n4676) & (n_n4703) & (n_n4698) & (x12621x)) + ((n_n4656) & (!n_n4676) & (!n_n4703) & (!n_n4698) & (!x12621x)) + ((n_n4656) & (!n_n4676) & (!n_n4703) & (!n_n4698) & (x12621x)) + ((n_n4656) & (!n_n4676) & (!n_n4703) & (n_n4698) & (!x12621x)) + ((n_n4656) & (!n_n4676) & (!n_n4703) & (n_n4698) & (x12621x)) + ((n_n4656) & (!n_n4676) & (n_n4703) & (!n_n4698) & (!x12621x)) + ((n_n4656) & (!n_n4676) & (n_n4703) & (!n_n4698) & (x12621x)) + ((n_n4656) & (!n_n4676) & (n_n4703) & (n_n4698) & (!x12621x)) + ((n_n4656) & (!n_n4676) & (n_n4703) & (n_n4698) & (x12621x)) + ((n_n4656) & (n_n4676) & (!n_n4703) & (!n_n4698) & (!x12621x)) + ((n_n4656) & (n_n4676) & (!n_n4703) & (!n_n4698) & (x12621x)) + ((n_n4656) & (n_n4676) & (!n_n4703) & (n_n4698) & (!x12621x)) + ((n_n4656) & (n_n4676) & (!n_n4703) & (n_n4698) & (x12621x)) + ((n_n4656) & (n_n4676) & (n_n4703) & (!n_n4698) & (!x12621x)) + ((n_n4656) & (n_n4676) & (n_n4703) & (!n_n4698) & (x12621x)) + ((n_n4656) & (n_n4676) & (n_n4703) & (n_n4698) & (!x12621x)) + ((n_n4656) & (n_n4676) & (n_n4703) & (n_n4698) & (x12621x)));
	assign n_n542 = (((!x12629x) & (!x165x) & (!x258x) & (!x12614x) & (n_n557)) + ((!x12629x) & (!x165x) & (!x258x) & (x12614x) & (!n_n557)) + ((!x12629x) & (!x165x) & (!x258x) & (x12614x) & (n_n557)) + ((!x12629x) & (!x165x) & (x258x) & (!x12614x) & (!n_n557)) + ((!x12629x) & (!x165x) & (x258x) & (!x12614x) & (n_n557)) + ((!x12629x) & (!x165x) & (x258x) & (x12614x) & (!n_n557)) + ((!x12629x) & (!x165x) & (x258x) & (x12614x) & (n_n557)) + ((!x12629x) & (x165x) & (!x258x) & (!x12614x) & (!n_n557)) + ((!x12629x) & (x165x) & (!x258x) & (!x12614x) & (n_n557)) + ((!x12629x) & (x165x) & (!x258x) & (x12614x) & (!n_n557)) + ((!x12629x) & (x165x) & (!x258x) & (x12614x) & (n_n557)) + ((!x12629x) & (x165x) & (x258x) & (!x12614x) & (!n_n557)) + ((!x12629x) & (x165x) & (x258x) & (!x12614x) & (n_n557)) + ((!x12629x) & (x165x) & (x258x) & (x12614x) & (!n_n557)) + ((!x12629x) & (x165x) & (x258x) & (x12614x) & (n_n557)) + ((x12629x) & (!x165x) & (!x258x) & (!x12614x) & (!n_n557)) + ((x12629x) & (!x165x) & (!x258x) & (!x12614x) & (n_n557)) + ((x12629x) & (!x165x) & (!x258x) & (x12614x) & (!n_n557)) + ((x12629x) & (!x165x) & (!x258x) & (x12614x) & (n_n557)) + ((x12629x) & (!x165x) & (x258x) & (!x12614x) & (!n_n557)) + ((x12629x) & (!x165x) & (x258x) & (!x12614x) & (n_n557)) + ((x12629x) & (!x165x) & (x258x) & (x12614x) & (!n_n557)) + ((x12629x) & (!x165x) & (x258x) & (x12614x) & (n_n557)) + ((x12629x) & (x165x) & (!x258x) & (!x12614x) & (!n_n557)) + ((x12629x) & (x165x) & (!x258x) & (!x12614x) & (n_n557)) + ((x12629x) & (x165x) & (!x258x) & (x12614x) & (!n_n557)) + ((x12629x) & (x165x) & (!x258x) & (x12614x) & (n_n557)) + ((x12629x) & (x165x) & (x258x) & (!x12614x) & (!n_n557)) + ((x12629x) & (x165x) & (x258x) & (!x12614x) & (n_n557)) + ((x12629x) & (x165x) & (x258x) & (x12614x) & (!n_n557)) + ((x12629x) & (x165x) & (x258x) & (x12614x) & (n_n557)));
	assign n_n553 = (((!n_n4885) & (!n_n4911) & (!n_n4903) & (!n_n4895) & (x12679x)) + ((!n_n4885) & (!n_n4911) & (!n_n4903) & (n_n4895) & (!x12679x)) + ((!n_n4885) & (!n_n4911) & (!n_n4903) & (n_n4895) & (x12679x)) + ((!n_n4885) & (!n_n4911) & (n_n4903) & (!n_n4895) & (!x12679x)) + ((!n_n4885) & (!n_n4911) & (n_n4903) & (!n_n4895) & (x12679x)) + ((!n_n4885) & (!n_n4911) & (n_n4903) & (n_n4895) & (!x12679x)) + ((!n_n4885) & (!n_n4911) & (n_n4903) & (n_n4895) & (x12679x)) + ((!n_n4885) & (n_n4911) & (!n_n4903) & (!n_n4895) & (!x12679x)) + ((!n_n4885) & (n_n4911) & (!n_n4903) & (!n_n4895) & (x12679x)) + ((!n_n4885) & (n_n4911) & (!n_n4903) & (n_n4895) & (!x12679x)) + ((!n_n4885) & (n_n4911) & (!n_n4903) & (n_n4895) & (x12679x)) + ((!n_n4885) & (n_n4911) & (n_n4903) & (!n_n4895) & (!x12679x)) + ((!n_n4885) & (n_n4911) & (n_n4903) & (!n_n4895) & (x12679x)) + ((!n_n4885) & (n_n4911) & (n_n4903) & (n_n4895) & (!x12679x)) + ((!n_n4885) & (n_n4911) & (n_n4903) & (n_n4895) & (x12679x)) + ((n_n4885) & (!n_n4911) & (!n_n4903) & (!n_n4895) & (!x12679x)) + ((n_n4885) & (!n_n4911) & (!n_n4903) & (!n_n4895) & (x12679x)) + ((n_n4885) & (!n_n4911) & (!n_n4903) & (n_n4895) & (!x12679x)) + ((n_n4885) & (!n_n4911) & (!n_n4903) & (n_n4895) & (x12679x)) + ((n_n4885) & (!n_n4911) & (n_n4903) & (!n_n4895) & (!x12679x)) + ((n_n4885) & (!n_n4911) & (n_n4903) & (!n_n4895) & (x12679x)) + ((n_n4885) & (!n_n4911) & (n_n4903) & (n_n4895) & (!x12679x)) + ((n_n4885) & (!n_n4911) & (n_n4903) & (n_n4895) & (x12679x)) + ((n_n4885) & (n_n4911) & (!n_n4903) & (!n_n4895) & (!x12679x)) + ((n_n4885) & (n_n4911) & (!n_n4903) & (!n_n4895) & (x12679x)) + ((n_n4885) & (n_n4911) & (!n_n4903) & (n_n4895) & (!x12679x)) + ((n_n4885) & (n_n4911) & (!n_n4903) & (n_n4895) & (x12679x)) + ((n_n4885) & (n_n4911) & (n_n4903) & (!n_n4895) & (!x12679x)) + ((n_n4885) & (n_n4911) & (n_n4903) & (!n_n4895) & (x12679x)) + ((n_n4885) & (n_n4911) & (n_n4903) & (n_n4895) & (!x12679x)) + ((n_n4885) & (n_n4911) & (n_n4903) & (n_n4895) & (x12679x)));
	assign x12683x = (((!x25x) & (!n_n260) & (!n_n535) & (!n_n4800) & (x38x)) + ((!x25x) & (!n_n260) & (!n_n535) & (n_n4800) & (!x38x)) + ((!x25x) & (!n_n260) & (!n_n535) & (n_n4800) & (x38x)) + ((!x25x) & (!n_n260) & (n_n535) & (!n_n4800) & (x38x)) + ((!x25x) & (!n_n260) & (n_n535) & (n_n4800) & (!x38x)) + ((!x25x) & (!n_n260) & (n_n535) & (n_n4800) & (x38x)) + ((!x25x) & (n_n260) & (!n_n535) & (!n_n4800) & (x38x)) + ((!x25x) & (n_n260) & (!n_n535) & (n_n4800) & (!x38x)) + ((!x25x) & (n_n260) & (!n_n535) & (n_n4800) & (x38x)) + ((!x25x) & (n_n260) & (n_n535) & (!n_n4800) & (x38x)) + ((!x25x) & (n_n260) & (n_n535) & (n_n4800) & (!x38x)) + ((!x25x) & (n_n260) & (n_n535) & (n_n4800) & (x38x)) + ((x25x) & (!n_n260) & (!n_n535) & (!n_n4800) & (x38x)) + ((x25x) & (!n_n260) & (!n_n535) & (n_n4800) & (!x38x)) + ((x25x) & (!n_n260) & (!n_n535) & (n_n4800) & (x38x)) + ((x25x) & (!n_n260) & (n_n535) & (!n_n4800) & (x38x)) + ((x25x) & (!n_n260) & (n_n535) & (n_n4800) & (!x38x)) + ((x25x) & (!n_n260) & (n_n535) & (n_n4800) & (x38x)) + ((x25x) & (n_n260) & (!n_n535) & (!n_n4800) & (x38x)) + ((x25x) & (n_n260) & (!n_n535) & (n_n4800) & (!x38x)) + ((x25x) & (n_n260) & (!n_n535) & (n_n4800) & (x38x)) + ((x25x) & (n_n260) & (n_n535) & (!n_n4800) & (!x38x)) + ((x25x) & (n_n260) & (n_n535) & (!n_n4800) & (x38x)) + ((x25x) & (n_n260) & (n_n535) & (n_n4800) & (!x38x)) + ((x25x) & (n_n260) & (n_n535) & (n_n4800) & (x38x)));
	assign x12684x = (((!x11x) & (!n_n4870) & (!x530x) & (!n_n4819) & (x395x)) + ((!x11x) & (!n_n4870) & (!x530x) & (n_n4819) & (!x395x)) + ((!x11x) & (!n_n4870) & (!x530x) & (n_n4819) & (x395x)) + ((!x11x) & (!n_n4870) & (x530x) & (!n_n4819) & (x395x)) + ((!x11x) & (!n_n4870) & (x530x) & (n_n4819) & (!x395x)) + ((!x11x) & (!n_n4870) & (x530x) & (n_n4819) & (x395x)) + ((!x11x) & (n_n4870) & (!x530x) & (!n_n4819) & (!x395x)) + ((!x11x) & (n_n4870) & (!x530x) & (!n_n4819) & (x395x)) + ((!x11x) & (n_n4870) & (!x530x) & (n_n4819) & (!x395x)) + ((!x11x) & (n_n4870) & (!x530x) & (n_n4819) & (x395x)) + ((!x11x) & (n_n4870) & (x530x) & (!n_n4819) & (!x395x)) + ((!x11x) & (n_n4870) & (x530x) & (!n_n4819) & (x395x)) + ((!x11x) & (n_n4870) & (x530x) & (n_n4819) & (!x395x)) + ((!x11x) & (n_n4870) & (x530x) & (n_n4819) & (x395x)) + ((x11x) & (!n_n4870) & (!x530x) & (!n_n4819) & (x395x)) + ((x11x) & (!n_n4870) & (!x530x) & (n_n4819) & (!x395x)) + ((x11x) & (!n_n4870) & (!x530x) & (n_n4819) & (x395x)) + ((x11x) & (!n_n4870) & (x530x) & (!n_n4819) & (!x395x)) + ((x11x) & (!n_n4870) & (x530x) & (!n_n4819) & (x395x)) + ((x11x) & (!n_n4870) & (x530x) & (n_n4819) & (!x395x)) + ((x11x) & (!n_n4870) & (x530x) & (n_n4819) & (x395x)) + ((x11x) & (n_n4870) & (!x530x) & (!n_n4819) & (!x395x)) + ((x11x) & (n_n4870) & (!x530x) & (!n_n4819) & (x395x)) + ((x11x) & (n_n4870) & (!x530x) & (n_n4819) & (!x395x)) + ((x11x) & (n_n4870) & (!x530x) & (n_n4819) & (x395x)) + ((x11x) & (n_n4870) & (x530x) & (!n_n4819) & (!x395x)) + ((x11x) & (n_n4870) & (x530x) & (!n_n4819) & (x395x)) + ((x11x) & (n_n4870) & (x530x) & (n_n4819) & (!x395x)) + ((x11x) & (n_n4870) & (x530x) & (n_n4819) & (x395x)));
	assign x12689x = (((!n_n4928) & (!n_n4950) & (!n_n4956) & (n_n4936)) + ((!n_n4928) & (!n_n4950) & (n_n4956) & (!n_n4936)) + ((!n_n4928) & (!n_n4950) & (n_n4956) & (n_n4936)) + ((!n_n4928) & (n_n4950) & (!n_n4956) & (!n_n4936)) + ((!n_n4928) & (n_n4950) & (!n_n4956) & (n_n4936)) + ((!n_n4928) & (n_n4950) & (n_n4956) & (!n_n4936)) + ((!n_n4928) & (n_n4950) & (n_n4956) & (n_n4936)) + ((n_n4928) & (!n_n4950) & (!n_n4956) & (!n_n4936)) + ((n_n4928) & (!n_n4950) & (!n_n4956) & (n_n4936)) + ((n_n4928) & (!n_n4950) & (n_n4956) & (!n_n4936)) + ((n_n4928) & (!n_n4950) & (n_n4956) & (n_n4936)) + ((n_n4928) & (n_n4950) & (!n_n4956) & (!n_n4936)) + ((n_n4928) & (n_n4950) & (!n_n4956) & (n_n4936)) + ((n_n4928) & (n_n4950) & (n_n4956) & (!n_n4936)) + ((n_n4928) & (n_n4950) & (n_n4956) & (n_n4936)));
	assign x12690x = (((!n_n4918) & (!n_n4917) & (!n_n4931) & (!n_n4948) & (n_n4954)) + ((!n_n4918) & (!n_n4917) & (!n_n4931) & (n_n4948) & (!n_n4954)) + ((!n_n4918) & (!n_n4917) & (!n_n4931) & (n_n4948) & (n_n4954)) + ((!n_n4918) & (!n_n4917) & (n_n4931) & (!n_n4948) & (!n_n4954)) + ((!n_n4918) & (!n_n4917) & (n_n4931) & (!n_n4948) & (n_n4954)) + ((!n_n4918) & (!n_n4917) & (n_n4931) & (n_n4948) & (!n_n4954)) + ((!n_n4918) & (!n_n4917) & (n_n4931) & (n_n4948) & (n_n4954)) + ((!n_n4918) & (n_n4917) & (!n_n4931) & (!n_n4948) & (!n_n4954)) + ((!n_n4918) & (n_n4917) & (!n_n4931) & (!n_n4948) & (n_n4954)) + ((!n_n4918) & (n_n4917) & (!n_n4931) & (n_n4948) & (!n_n4954)) + ((!n_n4918) & (n_n4917) & (!n_n4931) & (n_n4948) & (n_n4954)) + ((!n_n4918) & (n_n4917) & (n_n4931) & (!n_n4948) & (!n_n4954)) + ((!n_n4918) & (n_n4917) & (n_n4931) & (!n_n4948) & (n_n4954)) + ((!n_n4918) & (n_n4917) & (n_n4931) & (n_n4948) & (!n_n4954)) + ((!n_n4918) & (n_n4917) & (n_n4931) & (n_n4948) & (n_n4954)) + ((n_n4918) & (!n_n4917) & (!n_n4931) & (!n_n4948) & (!n_n4954)) + ((n_n4918) & (!n_n4917) & (!n_n4931) & (!n_n4948) & (n_n4954)) + ((n_n4918) & (!n_n4917) & (!n_n4931) & (n_n4948) & (!n_n4954)) + ((n_n4918) & (!n_n4917) & (!n_n4931) & (n_n4948) & (n_n4954)) + ((n_n4918) & (!n_n4917) & (n_n4931) & (!n_n4948) & (!n_n4954)) + ((n_n4918) & (!n_n4917) & (n_n4931) & (!n_n4948) & (n_n4954)) + ((n_n4918) & (!n_n4917) & (n_n4931) & (n_n4948) & (!n_n4954)) + ((n_n4918) & (!n_n4917) & (n_n4931) & (n_n4948) & (n_n4954)) + ((n_n4918) & (n_n4917) & (!n_n4931) & (!n_n4948) & (!n_n4954)) + ((n_n4918) & (n_n4917) & (!n_n4931) & (!n_n4948) & (n_n4954)) + ((n_n4918) & (n_n4917) & (!n_n4931) & (n_n4948) & (!n_n4954)) + ((n_n4918) & (n_n4917) & (!n_n4931) & (n_n4948) & (n_n4954)) + ((n_n4918) & (n_n4917) & (n_n4931) & (!n_n4948) & (!n_n4954)) + ((n_n4918) & (n_n4917) & (n_n4931) & (!n_n4948) & (n_n4954)) + ((n_n4918) & (n_n4917) & (n_n4931) & (n_n4948) & (!n_n4954)) + ((n_n4918) & (n_n4917) & (n_n4931) & (n_n4948) & (n_n4954)));
	assign x20x = (((!i_9_) & (!i_7_) & (i_8_) & (!i_6_)));
	assign x496x = (((i_1_) & (i_2_) & (i_0_) & (n_n464)));
	assign n_n4441 = (((!i_9_) & (n_n455) & (n_n534) & (n_n535)));
	assign n_n4404 = (((i_9_) & (n_n536) & (n_n482) & (n_n522)));
	assign n_n4384 = (((i_9_) & (n_n536) & (n_n526) & (n_n491)));
	assign x12700x = (((!x20x) & (!x496x) & (!n_n4441) & (!n_n4404) & (n_n4384)) + ((!x20x) & (!x496x) & (!n_n4441) & (n_n4404) & (!n_n4384)) + ((!x20x) & (!x496x) & (!n_n4441) & (n_n4404) & (n_n4384)) + ((!x20x) & (!x496x) & (n_n4441) & (!n_n4404) & (!n_n4384)) + ((!x20x) & (!x496x) & (n_n4441) & (!n_n4404) & (n_n4384)) + ((!x20x) & (!x496x) & (n_n4441) & (n_n4404) & (!n_n4384)) + ((!x20x) & (!x496x) & (n_n4441) & (n_n4404) & (n_n4384)) + ((!x20x) & (x496x) & (!n_n4441) & (!n_n4404) & (n_n4384)) + ((!x20x) & (x496x) & (!n_n4441) & (n_n4404) & (!n_n4384)) + ((!x20x) & (x496x) & (!n_n4441) & (n_n4404) & (n_n4384)) + ((!x20x) & (x496x) & (n_n4441) & (!n_n4404) & (!n_n4384)) + ((!x20x) & (x496x) & (n_n4441) & (!n_n4404) & (n_n4384)) + ((!x20x) & (x496x) & (n_n4441) & (n_n4404) & (!n_n4384)) + ((!x20x) & (x496x) & (n_n4441) & (n_n4404) & (n_n4384)) + ((x20x) & (!x496x) & (!n_n4441) & (!n_n4404) & (n_n4384)) + ((x20x) & (!x496x) & (!n_n4441) & (n_n4404) & (!n_n4384)) + ((x20x) & (!x496x) & (!n_n4441) & (n_n4404) & (n_n4384)) + ((x20x) & (!x496x) & (n_n4441) & (!n_n4404) & (!n_n4384)) + ((x20x) & (!x496x) & (n_n4441) & (!n_n4404) & (n_n4384)) + ((x20x) & (!x496x) & (n_n4441) & (n_n4404) & (!n_n4384)) + ((x20x) & (!x496x) & (n_n4441) & (n_n4404) & (n_n4384)) + ((x20x) & (x496x) & (!n_n4441) & (!n_n4404) & (!n_n4384)) + ((x20x) & (x496x) & (!n_n4441) & (!n_n4404) & (n_n4384)) + ((x20x) & (x496x) & (!n_n4441) & (n_n4404) & (!n_n4384)) + ((x20x) & (x496x) & (!n_n4441) & (n_n4404) & (n_n4384)) + ((x20x) & (x496x) & (n_n4441) & (!n_n4404) & (!n_n4384)) + ((x20x) & (x496x) & (n_n4441) & (!n_n4404) & (n_n4384)) + ((x20x) & (x496x) & (n_n4441) & (n_n4404) & (!n_n4384)) + ((x20x) & (x496x) & (n_n4441) & (n_n4404) & (n_n4384)));
	assign n_n4379 = (((!i_9_) & (n_n536) & (n_n532) & (n_n491)));
	assign n_n4371 = (((!i_9_) & (n_n536) & (n_n524) & (n_n500)));
	assign n_n4442 = (((i_9_) & (n_n455) & (n_n532) & (n_n535)));
	assign n_n4399 = (((!i_9_) & (n_n536) & (n_n482) & (n_n528)));
	assign n_n4417 = (((!i_9_) & (n_n536) & (n_n526) & (n_n473)));
	assign x12701x = (((!n_n4379) & (!n_n4371) & (!n_n4442) & (!n_n4399) & (n_n4417)) + ((!n_n4379) & (!n_n4371) & (!n_n4442) & (n_n4399) & (!n_n4417)) + ((!n_n4379) & (!n_n4371) & (!n_n4442) & (n_n4399) & (n_n4417)) + ((!n_n4379) & (!n_n4371) & (n_n4442) & (!n_n4399) & (!n_n4417)) + ((!n_n4379) & (!n_n4371) & (n_n4442) & (!n_n4399) & (n_n4417)) + ((!n_n4379) & (!n_n4371) & (n_n4442) & (n_n4399) & (!n_n4417)) + ((!n_n4379) & (!n_n4371) & (n_n4442) & (n_n4399) & (n_n4417)) + ((!n_n4379) & (n_n4371) & (!n_n4442) & (!n_n4399) & (!n_n4417)) + ((!n_n4379) & (n_n4371) & (!n_n4442) & (!n_n4399) & (n_n4417)) + ((!n_n4379) & (n_n4371) & (!n_n4442) & (n_n4399) & (!n_n4417)) + ((!n_n4379) & (n_n4371) & (!n_n4442) & (n_n4399) & (n_n4417)) + ((!n_n4379) & (n_n4371) & (n_n4442) & (!n_n4399) & (!n_n4417)) + ((!n_n4379) & (n_n4371) & (n_n4442) & (!n_n4399) & (n_n4417)) + ((!n_n4379) & (n_n4371) & (n_n4442) & (n_n4399) & (!n_n4417)) + ((!n_n4379) & (n_n4371) & (n_n4442) & (n_n4399) & (n_n4417)) + ((n_n4379) & (!n_n4371) & (!n_n4442) & (!n_n4399) & (!n_n4417)) + ((n_n4379) & (!n_n4371) & (!n_n4442) & (!n_n4399) & (n_n4417)) + ((n_n4379) & (!n_n4371) & (!n_n4442) & (n_n4399) & (!n_n4417)) + ((n_n4379) & (!n_n4371) & (!n_n4442) & (n_n4399) & (n_n4417)) + ((n_n4379) & (!n_n4371) & (n_n4442) & (!n_n4399) & (!n_n4417)) + ((n_n4379) & (!n_n4371) & (n_n4442) & (!n_n4399) & (n_n4417)) + ((n_n4379) & (!n_n4371) & (n_n4442) & (n_n4399) & (!n_n4417)) + ((n_n4379) & (!n_n4371) & (n_n4442) & (n_n4399) & (n_n4417)) + ((n_n4379) & (n_n4371) & (!n_n4442) & (!n_n4399) & (!n_n4417)) + ((n_n4379) & (n_n4371) & (!n_n4442) & (!n_n4399) & (n_n4417)) + ((n_n4379) & (n_n4371) & (!n_n4442) & (n_n4399) & (!n_n4417)) + ((n_n4379) & (n_n4371) & (!n_n4442) & (n_n4399) & (n_n4417)) + ((n_n4379) & (n_n4371) & (n_n4442) & (!n_n4399) & (!n_n4417)) + ((n_n4379) & (n_n4371) & (n_n4442) & (!n_n4399) & (n_n4417)) + ((n_n4379) & (n_n4371) & (n_n4442) & (n_n4399) & (!n_n4417)) + ((n_n4379) & (n_n4371) & (n_n4442) & (n_n4399) & (n_n4417)));
	assign n_n4450 = (((i_9_) & (n_n524) & (n_n455) & (n_n535)));
	assign n_n4460 = (((i_9_) & (n_n518) & (n_n455) & (n_n530)));
	assign n_n4473 = (((!i_9_) & (n_n455) & (n_n534) & (n_n509)));
	assign n_n4506 = (((i_9_) & (n_n455) & (n_n532) & (n_n491)));
	assign x12707x = (((!n_n4450) & (!n_n4460) & (!n_n4473) & (n_n4506)) + ((!n_n4450) & (!n_n4460) & (n_n4473) & (!n_n4506)) + ((!n_n4450) & (!n_n4460) & (n_n4473) & (n_n4506)) + ((!n_n4450) & (n_n4460) & (!n_n4473) & (!n_n4506)) + ((!n_n4450) & (n_n4460) & (!n_n4473) & (n_n4506)) + ((!n_n4450) & (n_n4460) & (n_n4473) & (!n_n4506)) + ((!n_n4450) & (n_n4460) & (n_n4473) & (n_n4506)) + ((n_n4450) & (!n_n4460) & (!n_n4473) & (!n_n4506)) + ((n_n4450) & (!n_n4460) & (!n_n4473) & (n_n4506)) + ((n_n4450) & (!n_n4460) & (n_n4473) & (!n_n4506)) + ((n_n4450) & (!n_n4460) & (n_n4473) & (n_n4506)) + ((n_n4450) & (n_n4460) & (!n_n4473) & (!n_n4506)) + ((n_n4450) & (n_n4460) & (!n_n4473) & (n_n4506)) + ((n_n4450) & (n_n4460) & (n_n4473) & (!n_n4506)) + ((n_n4450) & (n_n4460) & (n_n4473) & (n_n4506)));
	assign n_n4512 = (((i_9_) & (n_n526) & (n_n455) & (n_n491)));
	assign n_n4453 = (((i_1_) & (!i_2_) & (i_0_) & (n_n535) & (x20x)));
	assign n_n4471 = (((!i_5_) & (i_3_) & (i_4_) & (n_n455) & (x23x)));
	assign n_n4488 = (((i_9_) & (n_n455) & (n_n534) & (n_n500)));
	assign n_n4458 = (((i_9_) & (n_n518) & (n_n455) & (n_n532)));
	assign x12708x = (((!n_n4512) & (!n_n4453) & (!n_n4471) & (!n_n4488) & (n_n4458)) + ((!n_n4512) & (!n_n4453) & (!n_n4471) & (n_n4488) & (!n_n4458)) + ((!n_n4512) & (!n_n4453) & (!n_n4471) & (n_n4488) & (n_n4458)) + ((!n_n4512) & (!n_n4453) & (n_n4471) & (!n_n4488) & (!n_n4458)) + ((!n_n4512) & (!n_n4453) & (n_n4471) & (!n_n4488) & (n_n4458)) + ((!n_n4512) & (!n_n4453) & (n_n4471) & (n_n4488) & (!n_n4458)) + ((!n_n4512) & (!n_n4453) & (n_n4471) & (n_n4488) & (n_n4458)) + ((!n_n4512) & (n_n4453) & (!n_n4471) & (!n_n4488) & (!n_n4458)) + ((!n_n4512) & (n_n4453) & (!n_n4471) & (!n_n4488) & (n_n4458)) + ((!n_n4512) & (n_n4453) & (!n_n4471) & (n_n4488) & (!n_n4458)) + ((!n_n4512) & (n_n4453) & (!n_n4471) & (n_n4488) & (n_n4458)) + ((!n_n4512) & (n_n4453) & (n_n4471) & (!n_n4488) & (!n_n4458)) + ((!n_n4512) & (n_n4453) & (n_n4471) & (!n_n4488) & (n_n4458)) + ((!n_n4512) & (n_n4453) & (n_n4471) & (n_n4488) & (!n_n4458)) + ((!n_n4512) & (n_n4453) & (n_n4471) & (n_n4488) & (n_n4458)) + ((n_n4512) & (!n_n4453) & (!n_n4471) & (!n_n4488) & (!n_n4458)) + ((n_n4512) & (!n_n4453) & (!n_n4471) & (!n_n4488) & (n_n4458)) + ((n_n4512) & (!n_n4453) & (!n_n4471) & (n_n4488) & (!n_n4458)) + ((n_n4512) & (!n_n4453) & (!n_n4471) & (n_n4488) & (n_n4458)) + ((n_n4512) & (!n_n4453) & (n_n4471) & (!n_n4488) & (!n_n4458)) + ((n_n4512) & (!n_n4453) & (n_n4471) & (!n_n4488) & (n_n4458)) + ((n_n4512) & (!n_n4453) & (n_n4471) & (n_n4488) & (!n_n4458)) + ((n_n4512) & (!n_n4453) & (n_n4471) & (n_n4488) & (n_n4458)) + ((n_n4512) & (n_n4453) & (!n_n4471) & (!n_n4488) & (!n_n4458)) + ((n_n4512) & (n_n4453) & (!n_n4471) & (!n_n4488) & (n_n4458)) + ((n_n4512) & (n_n4453) & (!n_n4471) & (n_n4488) & (!n_n4458)) + ((n_n4512) & (n_n4453) & (!n_n4471) & (n_n4488) & (n_n4458)) + ((n_n4512) & (n_n4453) & (n_n4471) & (!n_n4488) & (!n_n4458)) + ((n_n4512) & (n_n4453) & (n_n4471) & (!n_n4488) & (n_n4458)) + ((n_n4512) & (n_n4453) & (n_n4471) & (n_n4488) & (!n_n4458)) + ((n_n4512) & (n_n4453) & (n_n4471) & (n_n4488) & (n_n4458)));
	assign n_n4363 = (((!i_9_) & (n_n536) & (n_n532) & (n_n500)));
	assign n_n4347 = (((!i_9_) & (n_n536) & (n_n532) & (n_n509)));
	assign n_n4320 = (((i_9_) & (n_n536) & (n_n526) & (n_n535)));
	assign n_n4315 = (((!i_9_) & (n_n536) & (n_n532) & (n_n535)));
	assign x12714x = (((!n_n4363) & (!n_n4347) & (!n_n4320) & (n_n4315)) + ((!n_n4363) & (!n_n4347) & (n_n4320) & (!n_n4315)) + ((!n_n4363) & (!n_n4347) & (n_n4320) & (n_n4315)) + ((!n_n4363) & (n_n4347) & (!n_n4320) & (!n_n4315)) + ((!n_n4363) & (n_n4347) & (!n_n4320) & (n_n4315)) + ((!n_n4363) & (n_n4347) & (n_n4320) & (!n_n4315)) + ((!n_n4363) & (n_n4347) & (n_n4320) & (n_n4315)) + ((n_n4363) & (!n_n4347) & (!n_n4320) & (!n_n4315)) + ((n_n4363) & (!n_n4347) & (!n_n4320) & (n_n4315)) + ((n_n4363) & (!n_n4347) & (n_n4320) & (!n_n4315)) + ((n_n4363) & (!n_n4347) & (n_n4320) & (n_n4315)) + ((n_n4363) & (n_n4347) & (!n_n4320) & (!n_n4315)) + ((n_n4363) & (n_n4347) & (!n_n4320) & (n_n4315)) + ((n_n4363) & (n_n4347) & (n_n4320) & (!n_n4315)) + ((n_n4363) & (n_n4347) & (n_n4320) & (n_n4315)));
	assign n_n4338 = (((i_9_) & (n_n536) & (n_n524) & (n_n518)));
	assign n_n4327 = (((i_1_) & (i_2_) & (i_0_) & (n_n535) & (x23x)));
	assign n_n4326 = (((i_9_) & (n_n536) & (n_n535) & (n_n520)));
	assign n_n4350 = (((i_9_) & (n_n536) & (n_n528) & (n_n509)));
	assign n_n4331 = (((!i_9_) & (n_n536) & (n_n518) & (n_n532)));
	assign x12715x = (((!n_n4338) & (!n_n4327) & (!n_n4326) & (!n_n4350) & (n_n4331)) + ((!n_n4338) & (!n_n4327) & (!n_n4326) & (n_n4350) & (!n_n4331)) + ((!n_n4338) & (!n_n4327) & (!n_n4326) & (n_n4350) & (n_n4331)) + ((!n_n4338) & (!n_n4327) & (n_n4326) & (!n_n4350) & (!n_n4331)) + ((!n_n4338) & (!n_n4327) & (n_n4326) & (!n_n4350) & (n_n4331)) + ((!n_n4338) & (!n_n4327) & (n_n4326) & (n_n4350) & (!n_n4331)) + ((!n_n4338) & (!n_n4327) & (n_n4326) & (n_n4350) & (n_n4331)) + ((!n_n4338) & (n_n4327) & (!n_n4326) & (!n_n4350) & (!n_n4331)) + ((!n_n4338) & (n_n4327) & (!n_n4326) & (!n_n4350) & (n_n4331)) + ((!n_n4338) & (n_n4327) & (!n_n4326) & (n_n4350) & (!n_n4331)) + ((!n_n4338) & (n_n4327) & (!n_n4326) & (n_n4350) & (n_n4331)) + ((!n_n4338) & (n_n4327) & (n_n4326) & (!n_n4350) & (!n_n4331)) + ((!n_n4338) & (n_n4327) & (n_n4326) & (!n_n4350) & (n_n4331)) + ((!n_n4338) & (n_n4327) & (n_n4326) & (n_n4350) & (!n_n4331)) + ((!n_n4338) & (n_n4327) & (n_n4326) & (n_n4350) & (n_n4331)) + ((n_n4338) & (!n_n4327) & (!n_n4326) & (!n_n4350) & (!n_n4331)) + ((n_n4338) & (!n_n4327) & (!n_n4326) & (!n_n4350) & (n_n4331)) + ((n_n4338) & (!n_n4327) & (!n_n4326) & (n_n4350) & (!n_n4331)) + ((n_n4338) & (!n_n4327) & (!n_n4326) & (n_n4350) & (n_n4331)) + ((n_n4338) & (!n_n4327) & (n_n4326) & (!n_n4350) & (!n_n4331)) + ((n_n4338) & (!n_n4327) & (n_n4326) & (!n_n4350) & (n_n4331)) + ((n_n4338) & (!n_n4327) & (n_n4326) & (n_n4350) & (!n_n4331)) + ((n_n4338) & (!n_n4327) & (n_n4326) & (n_n4350) & (n_n4331)) + ((n_n4338) & (n_n4327) & (!n_n4326) & (!n_n4350) & (!n_n4331)) + ((n_n4338) & (n_n4327) & (!n_n4326) & (!n_n4350) & (n_n4331)) + ((n_n4338) & (n_n4327) & (!n_n4326) & (n_n4350) & (!n_n4331)) + ((n_n4338) & (n_n4327) & (!n_n4326) & (n_n4350) & (n_n4331)) + ((n_n4338) & (n_n4327) & (n_n4326) & (!n_n4350) & (!n_n4331)) + ((n_n4338) & (n_n4327) & (n_n4326) & (!n_n4350) & (n_n4331)) + ((n_n4338) & (n_n4327) & (n_n4326) & (n_n4350) & (!n_n4331)) + ((n_n4338) & (n_n4327) & (n_n4326) & (n_n4350) & (n_n4331)));
	assign n_n630 = (((!n_n727) & (!x13016x) & (!n_n653) & (!x13046x) & (x13015x)) + ((!n_n727) & (!x13016x) & (!n_n653) & (x13046x) & (!x13015x)) + ((!n_n727) & (!x13016x) & (!n_n653) & (x13046x) & (x13015x)) + ((!n_n727) & (!x13016x) & (n_n653) & (!x13046x) & (!x13015x)) + ((!n_n727) & (!x13016x) & (n_n653) & (!x13046x) & (x13015x)) + ((!n_n727) & (!x13016x) & (n_n653) & (x13046x) & (!x13015x)) + ((!n_n727) & (!x13016x) & (n_n653) & (x13046x) & (x13015x)) + ((!n_n727) & (x13016x) & (!n_n653) & (!x13046x) & (!x13015x)) + ((!n_n727) & (x13016x) & (!n_n653) & (!x13046x) & (x13015x)) + ((!n_n727) & (x13016x) & (!n_n653) & (x13046x) & (!x13015x)) + ((!n_n727) & (x13016x) & (!n_n653) & (x13046x) & (x13015x)) + ((!n_n727) & (x13016x) & (n_n653) & (!x13046x) & (!x13015x)) + ((!n_n727) & (x13016x) & (n_n653) & (!x13046x) & (x13015x)) + ((!n_n727) & (x13016x) & (n_n653) & (x13046x) & (!x13015x)) + ((!n_n727) & (x13016x) & (n_n653) & (x13046x) & (x13015x)) + ((n_n727) & (!x13016x) & (!n_n653) & (!x13046x) & (!x13015x)) + ((n_n727) & (!x13016x) & (!n_n653) & (!x13046x) & (x13015x)) + ((n_n727) & (!x13016x) & (!n_n653) & (x13046x) & (!x13015x)) + ((n_n727) & (!x13016x) & (!n_n653) & (x13046x) & (x13015x)) + ((n_n727) & (!x13016x) & (n_n653) & (!x13046x) & (!x13015x)) + ((n_n727) & (!x13016x) & (n_n653) & (!x13046x) & (x13015x)) + ((n_n727) & (!x13016x) & (n_n653) & (x13046x) & (!x13015x)) + ((n_n727) & (!x13016x) & (n_n653) & (x13046x) & (x13015x)) + ((n_n727) & (x13016x) & (!n_n653) & (!x13046x) & (!x13015x)) + ((n_n727) & (x13016x) & (!n_n653) & (!x13046x) & (x13015x)) + ((n_n727) & (x13016x) & (!n_n653) & (x13046x) & (!x13015x)) + ((n_n727) & (x13016x) & (!n_n653) & (x13046x) & (x13015x)) + ((n_n727) & (x13016x) & (n_n653) & (!x13046x) & (!x13015x)) + ((n_n727) & (x13016x) & (n_n653) & (!x13046x) & (x13015x)) + ((n_n727) & (x13016x) & (n_n653) & (x13046x) & (!x13015x)) + ((n_n727) & (x13016x) & (n_n653) & (x13046x) & (x13015x)));
	assign n_n657 = (((!x74x) & (!x398x) & (!x13060x) & (!x13065x) & (x13064x)) + ((!x74x) & (!x398x) & (!x13060x) & (x13065x) & (!x13064x)) + ((!x74x) & (!x398x) & (!x13060x) & (x13065x) & (x13064x)) + ((!x74x) & (!x398x) & (x13060x) & (!x13065x) & (!x13064x)) + ((!x74x) & (!x398x) & (x13060x) & (!x13065x) & (x13064x)) + ((!x74x) & (!x398x) & (x13060x) & (x13065x) & (!x13064x)) + ((!x74x) & (!x398x) & (x13060x) & (x13065x) & (x13064x)) + ((!x74x) & (x398x) & (!x13060x) & (!x13065x) & (!x13064x)) + ((!x74x) & (x398x) & (!x13060x) & (!x13065x) & (x13064x)) + ((!x74x) & (x398x) & (!x13060x) & (x13065x) & (!x13064x)) + ((!x74x) & (x398x) & (!x13060x) & (x13065x) & (x13064x)) + ((!x74x) & (x398x) & (x13060x) & (!x13065x) & (!x13064x)) + ((!x74x) & (x398x) & (x13060x) & (!x13065x) & (x13064x)) + ((!x74x) & (x398x) & (x13060x) & (x13065x) & (!x13064x)) + ((!x74x) & (x398x) & (x13060x) & (x13065x) & (x13064x)) + ((x74x) & (!x398x) & (!x13060x) & (!x13065x) & (!x13064x)) + ((x74x) & (!x398x) & (!x13060x) & (!x13065x) & (x13064x)) + ((x74x) & (!x398x) & (!x13060x) & (x13065x) & (!x13064x)) + ((x74x) & (!x398x) & (!x13060x) & (x13065x) & (x13064x)) + ((x74x) & (!x398x) & (x13060x) & (!x13065x) & (!x13064x)) + ((x74x) & (!x398x) & (x13060x) & (!x13065x) & (x13064x)) + ((x74x) & (!x398x) & (x13060x) & (x13065x) & (!x13064x)) + ((x74x) & (!x398x) & (x13060x) & (x13065x) & (x13064x)) + ((x74x) & (x398x) & (!x13060x) & (!x13065x) & (!x13064x)) + ((x74x) & (x398x) & (!x13060x) & (!x13065x) & (x13064x)) + ((x74x) & (x398x) & (!x13060x) & (x13065x) & (!x13064x)) + ((x74x) & (x398x) & (!x13060x) & (x13065x) & (x13064x)) + ((x74x) & (x398x) & (x13060x) & (!x13065x) & (!x13064x)) + ((x74x) & (x398x) & (x13060x) & (!x13065x) & (x13064x)) + ((x74x) & (x398x) & (x13060x) & (x13065x) & (!x13064x)) + ((x74x) & (x398x) & (x13060x) & (x13065x) & (x13064x)));
	assign n_n656 = (((!n_n730) & (!x13074x) & (!x13075x) & (x13080x)) + ((!n_n730) & (!x13074x) & (x13075x) & (!x13080x)) + ((!n_n730) & (!x13074x) & (x13075x) & (x13080x)) + ((!n_n730) & (x13074x) & (!x13075x) & (!x13080x)) + ((!n_n730) & (x13074x) & (!x13075x) & (x13080x)) + ((!n_n730) & (x13074x) & (x13075x) & (!x13080x)) + ((!n_n730) & (x13074x) & (x13075x) & (x13080x)) + ((n_n730) & (!x13074x) & (!x13075x) & (!x13080x)) + ((n_n730) & (!x13074x) & (!x13075x) & (x13080x)) + ((n_n730) & (!x13074x) & (x13075x) & (!x13080x)) + ((n_n730) & (!x13074x) & (x13075x) & (x13080x)) + ((n_n730) & (x13074x) & (!x13075x) & (!x13080x)) + ((n_n730) & (x13074x) & (!x13075x) & (x13080x)) + ((n_n730) & (x13074x) & (x13075x) & (!x13080x)) + ((n_n730) & (x13074x) & (x13075x) & (x13080x)));
	assign x13088x = (((!x337x) & (!x124x) & (!n_n738) & (!n_n737) & (x13085x)) + ((!x337x) & (!x124x) & (!n_n738) & (n_n737) & (!x13085x)) + ((!x337x) & (!x124x) & (!n_n738) & (n_n737) & (x13085x)) + ((!x337x) & (!x124x) & (n_n738) & (!n_n737) & (!x13085x)) + ((!x337x) & (!x124x) & (n_n738) & (!n_n737) & (x13085x)) + ((!x337x) & (!x124x) & (n_n738) & (n_n737) & (!x13085x)) + ((!x337x) & (!x124x) & (n_n738) & (n_n737) & (x13085x)) + ((!x337x) & (x124x) & (!n_n738) & (!n_n737) & (!x13085x)) + ((!x337x) & (x124x) & (!n_n738) & (!n_n737) & (x13085x)) + ((!x337x) & (x124x) & (!n_n738) & (n_n737) & (!x13085x)) + ((!x337x) & (x124x) & (!n_n738) & (n_n737) & (x13085x)) + ((!x337x) & (x124x) & (n_n738) & (!n_n737) & (!x13085x)) + ((!x337x) & (x124x) & (n_n738) & (!n_n737) & (x13085x)) + ((!x337x) & (x124x) & (n_n738) & (n_n737) & (!x13085x)) + ((!x337x) & (x124x) & (n_n738) & (n_n737) & (x13085x)) + ((x337x) & (!x124x) & (!n_n738) & (!n_n737) & (!x13085x)) + ((x337x) & (!x124x) & (!n_n738) & (!n_n737) & (x13085x)) + ((x337x) & (!x124x) & (!n_n738) & (n_n737) & (!x13085x)) + ((x337x) & (!x124x) & (!n_n738) & (n_n737) & (x13085x)) + ((x337x) & (!x124x) & (n_n738) & (!n_n737) & (!x13085x)) + ((x337x) & (!x124x) & (n_n738) & (!n_n737) & (x13085x)) + ((x337x) & (!x124x) & (n_n738) & (n_n737) & (!x13085x)) + ((x337x) & (!x124x) & (n_n738) & (n_n737) & (x13085x)) + ((x337x) & (x124x) & (!n_n738) & (!n_n737) & (!x13085x)) + ((x337x) & (x124x) & (!n_n738) & (!n_n737) & (x13085x)) + ((x337x) & (x124x) & (!n_n738) & (n_n737) & (!x13085x)) + ((x337x) & (x124x) & (!n_n738) & (n_n737) & (x13085x)) + ((x337x) & (x124x) & (n_n738) & (!n_n737) & (!x13085x)) + ((x337x) & (x124x) & (n_n738) & (!n_n737) & (x13085x)) + ((x337x) & (x124x) & (n_n738) & (n_n737) & (!x13085x)) + ((x337x) & (x124x) & (n_n738) & (n_n737) & (x13085x)));
	assign n_n629 = (((!n_n719) & (!n_n651) & (!n_n650) & (!x13130x) & (x13131x)) + ((!n_n719) & (!n_n651) & (!n_n650) & (x13130x) & (!x13131x)) + ((!n_n719) & (!n_n651) & (!n_n650) & (x13130x) & (x13131x)) + ((!n_n719) & (!n_n651) & (n_n650) & (!x13130x) & (!x13131x)) + ((!n_n719) & (!n_n651) & (n_n650) & (!x13130x) & (x13131x)) + ((!n_n719) & (!n_n651) & (n_n650) & (x13130x) & (!x13131x)) + ((!n_n719) & (!n_n651) & (n_n650) & (x13130x) & (x13131x)) + ((!n_n719) & (n_n651) & (!n_n650) & (!x13130x) & (!x13131x)) + ((!n_n719) & (n_n651) & (!n_n650) & (!x13130x) & (x13131x)) + ((!n_n719) & (n_n651) & (!n_n650) & (x13130x) & (!x13131x)) + ((!n_n719) & (n_n651) & (!n_n650) & (x13130x) & (x13131x)) + ((!n_n719) & (n_n651) & (n_n650) & (!x13130x) & (!x13131x)) + ((!n_n719) & (n_n651) & (n_n650) & (!x13130x) & (x13131x)) + ((!n_n719) & (n_n651) & (n_n650) & (x13130x) & (!x13131x)) + ((!n_n719) & (n_n651) & (n_n650) & (x13130x) & (x13131x)) + ((n_n719) & (!n_n651) & (!n_n650) & (!x13130x) & (!x13131x)) + ((n_n719) & (!n_n651) & (!n_n650) & (!x13130x) & (x13131x)) + ((n_n719) & (!n_n651) & (!n_n650) & (x13130x) & (!x13131x)) + ((n_n719) & (!n_n651) & (!n_n650) & (x13130x) & (x13131x)) + ((n_n719) & (!n_n651) & (n_n650) & (!x13130x) & (!x13131x)) + ((n_n719) & (!n_n651) & (n_n650) & (!x13130x) & (x13131x)) + ((n_n719) & (!n_n651) & (n_n650) & (x13130x) & (!x13131x)) + ((n_n719) & (!n_n651) & (n_n650) & (x13130x) & (x13131x)) + ((n_n719) & (n_n651) & (!n_n650) & (!x13130x) & (!x13131x)) + ((n_n719) & (n_n651) & (!n_n650) & (!x13130x) & (x13131x)) + ((n_n719) & (n_n651) & (!n_n650) & (x13130x) & (!x13131x)) + ((n_n719) & (n_n651) & (!n_n650) & (x13130x) & (x13131x)) + ((n_n719) & (n_n651) & (n_n650) & (!x13130x) & (!x13131x)) + ((n_n719) & (n_n651) & (n_n650) & (!x13130x) & (x13131x)) + ((n_n719) & (n_n651) & (n_n650) & (x13130x) & (!x13131x)) + ((n_n719) & (n_n651) & (n_n650) & (x13130x) & (x13131x)));
	assign n_n627 = (((!n_n698) & (!x12752x) & (!n_n646) & (!x12775x) & (x12751x)) + ((!n_n698) & (!x12752x) & (!n_n646) & (x12775x) & (!x12751x)) + ((!n_n698) & (!x12752x) & (!n_n646) & (x12775x) & (x12751x)) + ((!n_n698) & (!x12752x) & (n_n646) & (!x12775x) & (!x12751x)) + ((!n_n698) & (!x12752x) & (n_n646) & (!x12775x) & (x12751x)) + ((!n_n698) & (!x12752x) & (n_n646) & (x12775x) & (!x12751x)) + ((!n_n698) & (!x12752x) & (n_n646) & (x12775x) & (x12751x)) + ((!n_n698) & (x12752x) & (!n_n646) & (!x12775x) & (!x12751x)) + ((!n_n698) & (x12752x) & (!n_n646) & (!x12775x) & (x12751x)) + ((!n_n698) & (x12752x) & (!n_n646) & (x12775x) & (!x12751x)) + ((!n_n698) & (x12752x) & (!n_n646) & (x12775x) & (x12751x)) + ((!n_n698) & (x12752x) & (n_n646) & (!x12775x) & (!x12751x)) + ((!n_n698) & (x12752x) & (n_n646) & (!x12775x) & (x12751x)) + ((!n_n698) & (x12752x) & (n_n646) & (x12775x) & (!x12751x)) + ((!n_n698) & (x12752x) & (n_n646) & (x12775x) & (x12751x)) + ((n_n698) & (!x12752x) & (!n_n646) & (!x12775x) & (!x12751x)) + ((n_n698) & (!x12752x) & (!n_n646) & (!x12775x) & (x12751x)) + ((n_n698) & (!x12752x) & (!n_n646) & (x12775x) & (!x12751x)) + ((n_n698) & (!x12752x) & (!n_n646) & (x12775x) & (x12751x)) + ((n_n698) & (!x12752x) & (n_n646) & (!x12775x) & (!x12751x)) + ((n_n698) & (!x12752x) & (n_n646) & (!x12775x) & (x12751x)) + ((n_n698) & (!x12752x) & (n_n646) & (x12775x) & (!x12751x)) + ((n_n698) & (!x12752x) & (n_n646) & (x12775x) & (x12751x)) + ((n_n698) & (x12752x) & (!n_n646) & (!x12775x) & (!x12751x)) + ((n_n698) & (x12752x) & (!n_n646) & (!x12775x) & (x12751x)) + ((n_n698) & (x12752x) & (!n_n646) & (x12775x) & (!x12751x)) + ((n_n698) & (x12752x) & (!n_n646) & (x12775x) & (x12751x)) + ((n_n698) & (x12752x) & (n_n646) & (!x12775x) & (!x12751x)) + ((n_n698) & (x12752x) & (n_n646) & (!x12775x) & (x12751x)) + ((n_n698) & (x12752x) & (n_n646) & (x12775x) & (!x12751x)) + ((n_n698) & (x12752x) & (n_n646) & (x12775x) & (x12751x)));
	assign n_n628 = (((!n_n648) & (!n_n649) & (x12827x)) + ((!n_n648) & (n_n649) & (!x12827x)) + ((!n_n648) & (n_n649) & (x12827x)) + ((n_n648) & (!n_n649) & (!x12827x)) + ((n_n648) & (!n_n649) & (x12827x)) + ((n_n648) & (n_n649) & (!x12827x)) + ((n_n648) & (n_n649) & (x12827x)));
	assign x12867x = (((!n_n642) & (!n_n641) & (x12865x)) + ((!n_n642) & (n_n641) & (!x12865x)) + ((!n_n642) & (n_n641) & (x12865x)) + ((n_n642) & (!n_n641) & (!x12865x)) + ((n_n642) & (!n_n641) & (x12865x)) + ((n_n642) & (n_n641) & (!x12865x)) + ((n_n642) & (n_n641) & (x12865x)));
	assign x13001x = (((!n_n634) & (!x12984x) & (x12999x)) + ((!n_n634) & (x12984x) & (!x12999x)) + ((!n_n634) & (x12984x) & (x12999x)) + ((n_n634) & (!x12984x) & (!x12999x)) + ((n_n634) & (!x12984x) & (x12999x)) + ((n_n634) & (x12984x) & (!x12999x)) + ((n_n634) & (x12984x) & (x12999x)));
	assign x13002x = (((!n_n635) & (!n_n637) & (!n_n639) & (!n_n638) & (x12947x)) + ((!n_n635) & (!n_n637) & (!n_n639) & (n_n638) & (!x12947x)) + ((!n_n635) & (!n_n637) & (!n_n639) & (n_n638) & (x12947x)) + ((!n_n635) & (!n_n637) & (n_n639) & (!n_n638) & (!x12947x)) + ((!n_n635) & (!n_n637) & (n_n639) & (!n_n638) & (x12947x)) + ((!n_n635) & (!n_n637) & (n_n639) & (n_n638) & (!x12947x)) + ((!n_n635) & (!n_n637) & (n_n639) & (n_n638) & (x12947x)) + ((!n_n635) & (n_n637) & (!n_n639) & (!n_n638) & (!x12947x)) + ((!n_n635) & (n_n637) & (!n_n639) & (!n_n638) & (x12947x)) + ((!n_n635) & (n_n637) & (!n_n639) & (n_n638) & (!x12947x)) + ((!n_n635) & (n_n637) & (!n_n639) & (n_n638) & (x12947x)) + ((!n_n635) & (n_n637) & (n_n639) & (!n_n638) & (!x12947x)) + ((!n_n635) & (n_n637) & (n_n639) & (!n_n638) & (x12947x)) + ((!n_n635) & (n_n637) & (n_n639) & (n_n638) & (!x12947x)) + ((!n_n635) & (n_n637) & (n_n639) & (n_n638) & (x12947x)) + ((n_n635) & (!n_n637) & (!n_n639) & (!n_n638) & (!x12947x)) + ((n_n635) & (!n_n637) & (!n_n639) & (!n_n638) & (x12947x)) + ((n_n635) & (!n_n637) & (!n_n639) & (n_n638) & (!x12947x)) + ((n_n635) & (!n_n637) & (!n_n639) & (n_n638) & (x12947x)) + ((n_n635) & (!n_n637) & (n_n639) & (!n_n638) & (!x12947x)) + ((n_n635) & (!n_n637) & (n_n639) & (!n_n638) & (x12947x)) + ((n_n635) & (!n_n637) & (n_n639) & (n_n638) & (!x12947x)) + ((n_n635) & (!n_n637) & (n_n639) & (n_n638) & (x12947x)) + ((n_n635) & (n_n637) & (!n_n639) & (!n_n638) & (!x12947x)) + ((n_n635) & (n_n637) & (!n_n639) & (!n_n638) & (x12947x)) + ((n_n635) & (n_n637) & (!n_n639) & (n_n638) & (!x12947x)) + ((n_n635) & (n_n637) & (!n_n639) & (n_n638) & (x12947x)) + ((n_n635) & (n_n637) & (n_n639) & (!n_n638) & (!x12947x)) + ((n_n635) & (n_n637) & (n_n639) & (!n_n638) & (x12947x)) + ((n_n635) & (n_n637) & (n_n639) & (n_n638) & (!x12947x)) + ((n_n635) & (n_n637) & (n_n639) & (n_n638) & (x12947x)));
	assign n_n526 = (((i_7_) & (i_8_) & (!i_6_)));
	assign n_n5297 = (((!i_9_) & (n_n526) & (n_n482) & (n_n65)));
	assign n_n3990 = (((!n_n4007) & (!x13235x) & (x13234x)) + ((!n_n4007) & (x13235x) & (!x13234x)) + ((!n_n4007) & (x13235x) & (x13234x)) + ((n_n4007) & (!x13235x) & (!x13234x)) + ((n_n4007) & (!x13235x) & (x13234x)) + ((n_n4007) & (x13235x) & (!x13234x)) + ((n_n4007) & (x13235x) & (x13234x)));
	assign n_n3992 = (((!n_n4072) & (!n_n1087) & (!n_n4013) & (!n_n4014) & (x13276x)) + ((!n_n4072) & (!n_n1087) & (!n_n4013) & (n_n4014) & (!x13276x)) + ((!n_n4072) & (!n_n1087) & (!n_n4013) & (n_n4014) & (x13276x)) + ((!n_n4072) & (!n_n1087) & (n_n4013) & (!n_n4014) & (!x13276x)) + ((!n_n4072) & (!n_n1087) & (n_n4013) & (!n_n4014) & (x13276x)) + ((!n_n4072) & (!n_n1087) & (n_n4013) & (n_n4014) & (!x13276x)) + ((!n_n4072) & (!n_n1087) & (n_n4013) & (n_n4014) & (x13276x)) + ((!n_n4072) & (n_n1087) & (!n_n4013) & (!n_n4014) & (!x13276x)) + ((!n_n4072) & (n_n1087) & (!n_n4013) & (!n_n4014) & (x13276x)) + ((!n_n4072) & (n_n1087) & (!n_n4013) & (n_n4014) & (!x13276x)) + ((!n_n4072) & (n_n1087) & (!n_n4013) & (n_n4014) & (x13276x)) + ((!n_n4072) & (n_n1087) & (n_n4013) & (!n_n4014) & (!x13276x)) + ((!n_n4072) & (n_n1087) & (n_n4013) & (!n_n4014) & (x13276x)) + ((!n_n4072) & (n_n1087) & (n_n4013) & (n_n4014) & (!x13276x)) + ((!n_n4072) & (n_n1087) & (n_n4013) & (n_n4014) & (x13276x)) + ((n_n4072) & (!n_n1087) & (!n_n4013) & (!n_n4014) & (!x13276x)) + ((n_n4072) & (!n_n1087) & (!n_n4013) & (!n_n4014) & (x13276x)) + ((n_n4072) & (!n_n1087) & (!n_n4013) & (n_n4014) & (!x13276x)) + ((n_n4072) & (!n_n1087) & (!n_n4013) & (n_n4014) & (x13276x)) + ((n_n4072) & (!n_n1087) & (n_n4013) & (!n_n4014) & (!x13276x)) + ((n_n4072) & (!n_n1087) & (n_n4013) & (!n_n4014) & (x13276x)) + ((n_n4072) & (!n_n1087) & (n_n4013) & (n_n4014) & (!x13276x)) + ((n_n4072) & (!n_n1087) & (n_n4013) & (n_n4014) & (x13276x)) + ((n_n4072) & (n_n1087) & (!n_n4013) & (!n_n4014) & (!x13276x)) + ((n_n4072) & (n_n1087) & (!n_n4013) & (!n_n4014) & (x13276x)) + ((n_n4072) & (n_n1087) & (!n_n4013) & (n_n4014) & (!x13276x)) + ((n_n4072) & (n_n1087) & (!n_n4013) & (n_n4014) & (x13276x)) + ((n_n4072) & (n_n1087) & (n_n4013) & (!n_n4014) & (!x13276x)) + ((n_n4072) & (n_n1087) & (n_n4013) & (!n_n4014) & (x13276x)) + ((n_n4072) & (n_n1087) & (n_n4013) & (n_n4014) & (!x13276x)) + ((n_n4072) & (n_n1087) & (n_n4013) & (n_n4014) & (x13276x)));
	assign n_n3988 = (((!x13303x) & (!n_n4002) & (!x13326x) & (!n_n4036) & (n_n4037)) + ((!x13303x) & (!n_n4002) & (!x13326x) & (n_n4036) & (!n_n4037)) + ((!x13303x) & (!n_n4002) & (!x13326x) & (n_n4036) & (n_n4037)) + ((!x13303x) & (!n_n4002) & (x13326x) & (!n_n4036) & (!n_n4037)) + ((!x13303x) & (!n_n4002) & (x13326x) & (!n_n4036) & (n_n4037)) + ((!x13303x) & (!n_n4002) & (x13326x) & (n_n4036) & (!n_n4037)) + ((!x13303x) & (!n_n4002) & (x13326x) & (n_n4036) & (n_n4037)) + ((!x13303x) & (n_n4002) & (!x13326x) & (!n_n4036) & (!n_n4037)) + ((!x13303x) & (n_n4002) & (!x13326x) & (!n_n4036) & (n_n4037)) + ((!x13303x) & (n_n4002) & (!x13326x) & (n_n4036) & (!n_n4037)) + ((!x13303x) & (n_n4002) & (!x13326x) & (n_n4036) & (n_n4037)) + ((!x13303x) & (n_n4002) & (x13326x) & (!n_n4036) & (!n_n4037)) + ((!x13303x) & (n_n4002) & (x13326x) & (!n_n4036) & (n_n4037)) + ((!x13303x) & (n_n4002) & (x13326x) & (n_n4036) & (!n_n4037)) + ((!x13303x) & (n_n4002) & (x13326x) & (n_n4036) & (n_n4037)) + ((x13303x) & (!n_n4002) & (!x13326x) & (!n_n4036) & (!n_n4037)) + ((x13303x) & (!n_n4002) & (!x13326x) & (!n_n4036) & (n_n4037)) + ((x13303x) & (!n_n4002) & (!x13326x) & (n_n4036) & (!n_n4037)) + ((x13303x) & (!n_n4002) & (!x13326x) & (n_n4036) & (n_n4037)) + ((x13303x) & (!n_n4002) & (x13326x) & (!n_n4036) & (!n_n4037)) + ((x13303x) & (!n_n4002) & (x13326x) & (!n_n4036) & (n_n4037)) + ((x13303x) & (!n_n4002) & (x13326x) & (n_n4036) & (!n_n4037)) + ((x13303x) & (!n_n4002) & (x13326x) & (n_n4036) & (n_n4037)) + ((x13303x) & (n_n4002) & (!x13326x) & (!n_n4036) & (!n_n4037)) + ((x13303x) & (n_n4002) & (!x13326x) & (!n_n4036) & (n_n4037)) + ((x13303x) & (n_n4002) & (!x13326x) & (n_n4036) & (!n_n4037)) + ((x13303x) & (n_n4002) & (!x13326x) & (n_n4036) & (n_n4037)) + ((x13303x) & (n_n4002) & (x13326x) & (!n_n4036) & (!n_n4037)) + ((x13303x) & (n_n4002) & (x13326x) & (!n_n4036) & (n_n4037)) + ((x13303x) & (n_n4002) & (x13326x) & (n_n4036) & (!n_n4037)) + ((x13303x) & (n_n4002) & (x13326x) & (n_n4036) & (n_n4037)));
	assign n_n3987 = (((!n_n3998) & (!n_n3999) & (x13374x)) + ((!n_n3998) & (n_n3999) & (!x13374x)) + ((!n_n3998) & (n_n3999) & (x13374x)) + ((n_n3998) & (!n_n3999) & (!x13374x)) + ((n_n3998) & (!n_n3999) & (x13374x)) + ((n_n3998) & (n_n3999) & (!x13374x)) + ((n_n3998) & (n_n3999) & (x13374x)));
	assign n_n3989 = (((!n_n4051) & (!n_n4050) & (!n_n4003) & (!n_n4004) & (x13421x)) + ((!n_n4051) & (!n_n4050) & (!n_n4003) & (n_n4004) & (!x13421x)) + ((!n_n4051) & (!n_n4050) & (!n_n4003) & (n_n4004) & (x13421x)) + ((!n_n4051) & (!n_n4050) & (n_n4003) & (!n_n4004) & (!x13421x)) + ((!n_n4051) & (!n_n4050) & (n_n4003) & (!n_n4004) & (x13421x)) + ((!n_n4051) & (!n_n4050) & (n_n4003) & (n_n4004) & (!x13421x)) + ((!n_n4051) & (!n_n4050) & (n_n4003) & (n_n4004) & (x13421x)) + ((!n_n4051) & (n_n4050) & (!n_n4003) & (!n_n4004) & (!x13421x)) + ((!n_n4051) & (n_n4050) & (!n_n4003) & (!n_n4004) & (x13421x)) + ((!n_n4051) & (n_n4050) & (!n_n4003) & (n_n4004) & (!x13421x)) + ((!n_n4051) & (n_n4050) & (!n_n4003) & (n_n4004) & (x13421x)) + ((!n_n4051) & (n_n4050) & (n_n4003) & (!n_n4004) & (!x13421x)) + ((!n_n4051) & (n_n4050) & (n_n4003) & (!n_n4004) & (x13421x)) + ((!n_n4051) & (n_n4050) & (n_n4003) & (n_n4004) & (!x13421x)) + ((!n_n4051) & (n_n4050) & (n_n4003) & (n_n4004) & (x13421x)) + ((n_n4051) & (!n_n4050) & (!n_n4003) & (!n_n4004) & (!x13421x)) + ((n_n4051) & (!n_n4050) & (!n_n4003) & (!n_n4004) & (x13421x)) + ((n_n4051) & (!n_n4050) & (!n_n4003) & (n_n4004) & (!x13421x)) + ((n_n4051) & (!n_n4050) & (!n_n4003) & (n_n4004) & (x13421x)) + ((n_n4051) & (!n_n4050) & (n_n4003) & (!n_n4004) & (!x13421x)) + ((n_n4051) & (!n_n4050) & (n_n4003) & (!n_n4004) & (x13421x)) + ((n_n4051) & (!n_n4050) & (n_n4003) & (n_n4004) & (!x13421x)) + ((n_n4051) & (!n_n4050) & (n_n4003) & (n_n4004) & (x13421x)) + ((n_n4051) & (n_n4050) & (!n_n4003) & (!n_n4004) & (!x13421x)) + ((n_n4051) & (n_n4050) & (!n_n4003) & (!n_n4004) & (x13421x)) + ((n_n4051) & (n_n4050) & (!n_n4003) & (n_n4004) & (!x13421x)) + ((n_n4051) & (n_n4050) & (!n_n4003) & (n_n4004) & (x13421x)) + ((n_n4051) & (n_n4050) & (n_n4003) & (!n_n4004) & (!x13421x)) + ((n_n4051) & (n_n4050) & (n_n4003) & (!n_n4004) & (x13421x)) + ((n_n4051) & (n_n4050) & (n_n4003) & (n_n4004) & (!x13421x)) + ((n_n4051) & (n_n4050) & (n_n4003) & (n_n4004) & (x13421x)));
	assign n_n3993 = (((!x13482x) & (!n_n4016) & (n_n4015)) + ((!x13482x) & (n_n4016) & (!n_n4015)) + ((!x13482x) & (n_n4016) & (n_n4015)) + ((x13482x) & (!n_n4016) & (!n_n4015)) + ((x13482x) & (!n_n4016) & (n_n4015)) + ((x13482x) & (n_n4016) & (!n_n4015)) + ((x13482x) & (n_n4016) & (n_n4015)));
	assign n_n3995 = (((!n_n4023) & (!n_n4100) & (!n_n4102) & (!n_n4021) & (x13545x)) + ((!n_n4023) & (!n_n4100) & (!n_n4102) & (n_n4021) & (!x13545x)) + ((!n_n4023) & (!n_n4100) & (!n_n4102) & (n_n4021) & (x13545x)) + ((!n_n4023) & (!n_n4100) & (n_n4102) & (!n_n4021) & (!x13545x)) + ((!n_n4023) & (!n_n4100) & (n_n4102) & (!n_n4021) & (x13545x)) + ((!n_n4023) & (!n_n4100) & (n_n4102) & (n_n4021) & (!x13545x)) + ((!n_n4023) & (!n_n4100) & (n_n4102) & (n_n4021) & (x13545x)) + ((!n_n4023) & (n_n4100) & (!n_n4102) & (!n_n4021) & (!x13545x)) + ((!n_n4023) & (n_n4100) & (!n_n4102) & (!n_n4021) & (x13545x)) + ((!n_n4023) & (n_n4100) & (!n_n4102) & (n_n4021) & (!x13545x)) + ((!n_n4023) & (n_n4100) & (!n_n4102) & (n_n4021) & (x13545x)) + ((!n_n4023) & (n_n4100) & (n_n4102) & (!n_n4021) & (!x13545x)) + ((!n_n4023) & (n_n4100) & (n_n4102) & (!n_n4021) & (x13545x)) + ((!n_n4023) & (n_n4100) & (n_n4102) & (n_n4021) & (!x13545x)) + ((!n_n4023) & (n_n4100) & (n_n4102) & (n_n4021) & (x13545x)) + ((n_n4023) & (!n_n4100) & (!n_n4102) & (!n_n4021) & (!x13545x)) + ((n_n4023) & (!n_n4100) & (!n_n4102) & (!n_n4021) & (x13545x)) + ((n_n4023) & (!n_n4100) & (!n_n4102) & (n_n4021) & (!x13545x)) + ((n_n4023) & (!n_n4100) & (!n_n4102) & (n_n4021) & (x13545x)) + ((n_n4023) & (!n_n4100) & (n_n4102) & (!n_n4021) & (!x13545x)) + ((n_n4023) & (!n_n4100) & (n_n4102) & (!n_n4021) & (x13545x)) + ((n_n4023) & (!n_n4100) & (n_n4102) & (n_n4021) & (!x13545x)) + ((n_n4023) & (!n_n4100) & (n_n4102) & (n_n4021) & (x13545x)) + ((n_n4023) & (n_n4100) & (!n_n4102) & (!n_n4021) & (!x13545x)) + ((n_n4023) & (n_n4100) & (!n_n4102) & (!n_n4021) & (x13545x)) + ((n_n4023) & (n_n4100) & (!n_n4102) & (n_n4021) & (!x13545x)) + ((n_n4023) & (n_n4100) & (!n_n4102) & (n_n4021) & (x13545x)) + ((n_n4023) & (n_n4100) & (n_n4102) & (!n_n4021) & (!x13545x)) + ((n_n4023) & (n_n4100) & (n_n4102) & (!n_n4021) & (x13545x)) + ((n_n4023) & (n_n4100) & (n_n4102) & (n_n4021) & (!x13545x)) + ((n_n4023) & (n_n4100) & (n_n4102) & (n_n4021) & (x13545x)));
	assign x13555x = (((!n_n4020) & (!x13501x) & (!n_n4090) & (!x13500x) & (x13553x)) + ((!n_n4020) & (!x13501x) & (!n_n4090) & (x13500x) & (!x13553x)) + ((!n_n4020) & (!x13501x) & (!n_n4090) & (x13500x) & (x13553x)) + ((!n_n4020) & (!x13501x) & (n_n4090) & (!x13500x) & (!x13553x)) + ((!n_n4020) & (!x13501x) & (n_n4090) & (!x13500x) & (x13553x)) + ((!n_n4020) & (!x13501x) & (n_n4090) & (x13500x) & (!x13553x)) + ((!n_n4020) & (!x13501x) & (n_n4090) & (x13500x) & (x13553x)) + ((!n_n4020) & (x13501x) & (!n_n4090) & (!x13500x) & (!x13553x)) + ((!n_n4020) & (x13501x) & (!n_n4090) & (!x13500x) & (x13553x)) + ((!n_n4020) & (x13501x) & (!n_n4090) & (x13500x) & (!x13553x)) + ((!n_n4020) & (x13501x) & (!n_n4090) & (x13500x) & (x13553x)) + ((!n_n4020) & (x13501x) & (n_n4090) & (!x13500x) & (!x13553x)) + ((!n_n4020) & (x13501x) & (n_n4090) & (!x13500x) & (x13553x)) + ((!n_n4020) & (x13501x) & (n_n4090) & (x13500x) & (!x13553x)) + ((!n_n4020) & (x13501x) & (n_n4090) & (x13500x) & (x13553x)) + ((n_n4020) & (!x13501x) & (!n_n4090) & (!x13500x) & (!x13553x)) + ((n_n4020) & (!x13501x) & (!n_n4090) & (!x13500x) & (x13553x)) + ((n_n4020) & (!x13501x) & (!n_n4090) & (x13500x) & (!x13553x)) + ((n_n4020) & (!x13501x) & (!n_n4090) & (x13500x) & (x13553x)) + ((n_n4020) & (!x13501x) & (n_n4090) & (!x13500x) & (!x13553x)) + ((n_n4020) & (!x13501x) & (n_n4090) & (!x13500x) & (x13553x)) + ((n_n4020) & (!x13501x) & (n_n4090) & (x13500x) & (!x13553x)) + ((n_n4020) & (!x13501x) & (n_n4090) & (x13500x) & (x13553x)) + ((n_n4020) & (x13501x) & (!n_n4090) & (!x13500x) & (!x13553x)) + ((n_n4020) & (x13501x) & (!n_n4090) & (!x13500x) & (x13553x)) + ((n_n4020) & (x13501x) & (!n_n4090) & (x13500x) & (!x13553x)) + ((n_n4020) & (x13501x) & (!n_n4090) & (x13500x) & (x13553x)) + ((n_n4020) & (x13501x) & (n_n4090) & (!x13500x) & (!x13553x)) + ((n_n4020) & (x13501x) & (n_n4090) & (!x13500x) & (x13553x)) + ((n_n4020) & (x13501x) & (n_n4090) & (x13500x) & (!x13553x)) + ((n_n4020) & (x13501x) & (n_n4090) & (x13500x) & (x13553x)));
	assign x13569x = (((!n_n4010) & (!n_n4009) & (!x13188x) & (n_n3996)) + ((!n_n4010) & (!n_n4009) & (x13188x) & (!n_n3996)) + ((!n_n4010) & (!n_n4009) & (x13188x) & (n_n3996)) + ((!n_n4010) & (n_n4009) & (!x13188x) & (!n_n3996)) + ((!n_n4010) & (n_n4009) & (!x13188x) & (n_n3996)) + ((!n_n4010) & (n_n4009) & (x13188x) & (!n_n3996)) + ((!n_n4010) & (n_n4009) & (x13188x) & (n_n3996)) + ((n_n4010) & (!n_n4009) & (!x13188x) & (!n_n3996)) + ((n_n4010) & (!n_n4009) & (!x13188x) & (n_n3996)) + ((n_n4010) & (!n_n4009) & (x13188x) & (!n_n3996)) + ((n_n4010) & (!n_n4009) & (x13188x) & (n_n3996)) + ((n_n4010) & (n_n4009) & (!x13188x) & (!n_n3996)) + ((n_n4010) & (n_n4009) & (!x13188x) & (n_n3996)) + ((n_n4010) & (n_n4009) & (x13188x) & (!n_n3996)) + ((n_n4010) & (n_n4009) & (x13188x) & (n_n3996)));
	assign x13606x = (((!n_n5017) & (!n_n5015) & (!n_n5037) & (n_n5056)) + ((!n_n5017) & (!n_n5015) & (n_n5037) & (!n_n5056)) + ((!n_n5017) & (!n_n5015) & (n_n5037) & (n_n5056)) + ((!n_n5017) & (n_n5015) & (!n_n5037) & (!n_n5056)) + ((!n_n5017) & (n_n5015) & (!n_n5037) & (n_n5056)) + ((!n_n5017) & (n_n5015) & (n_n5037) & (!n_n5056)) + ((!n_n5017) & (n_n5015) & (n_n5037) & (n_n5056)) + ((n_n5017) & (!n_n5015) & (!n_n5037) & (!n_n5056)) + ((n_n5017) & (!n_n5015) & (!n_n5037) & (n_n5056)) + ((n_n5017) & (!n_n5015) & (n_n5037) & (!n_n5056)) + ((n_n5017) & (!n_n5015) & (n_n5037) & (n_n5056)) + ((n_n5017) & (n_n5015) & (!n_n5037) & (!n_n5056)) + ((n_n5017) & (n_n5015) & (!n_n5037) & (n_n5056)) + ((n_n5017) & (n_n5015) & (n_n5037) & (!n_n5056)) + ((n_n5017) & (n_n5015) & (n_n5037) & (n_n5056)));
	assign x13607x = (((!n_n5032) & (!n_n5036) & (!n_n5021) & (!n_n5020) & (n_n5047)) + ((!n_n5032) & (!n_n5036) & (!n_n5021) & (n_n5020) & (!n_n5047)) + ((!n_n5032) & (!n_n5036) & (!n_n5021) & (n_n5020) & (n_n5047)) + ((!n_n5032) & (!n_n5036) & (n_n5021) & (!n_n5020) & (!n_n5047)) + ((!n_n5032) & (!n_n5036) & (n_n5021) & (!n_n5020) & (n_n5047)) + ((!n_n5032) & (!n_n5036) & (n_n5021) & (n_n5020) & (!n_n5047)) + ((!n_n5032) & (!n_n5036) & (n_n5021) & (n_n5020) & (n_n5047)) + ((!n_n5032) & (n_n5036) & (!n_n5021) & (!n_n5020) & (!n_n5047)) + ((!n_n5032) & (n_n5036) & (!n_n5021) & (!n_n5020) & (n_n5047)) + ((!n_n5032) & (n_n5036) & (!n_n5021) & (n_n5020) & (!n_n5047)) + ((!n_n5032) & (n_n5036) & (!n_n5021) & (n_n5020) & (n_n5047)) + ((!n_n5032) & (n_n5036) & (n_n5021) & (!n_n5020) & (!n_n5047)) + ((!n_n5032) & (n_n5036) & (n_n5021) & (!n_n5020) & (n_n5047)) + ((!n_n5032) & (n_n5036) & (n_n5021) & (n_n5020) & (!n_n5047)) + ((!n_n5032) & (n_n5036) & (n_n5021) & (n_n5020) & (n_n5047)) + ((n_n5032) & (!n_n5036) & (!n_n5021) & (!n_n5020) & (!n_n5047)) + ((n_n5032) & (!n_n5036) & (!n_n5021) & (!n_n5020) & (n_n5047)) + ((n_n5032) & (!n_n5036) & (!n_n5021) & (n_n5020) & (!n_n5047)) + ((n_n5032) & (!n_n5036) & (!n_n5021) & (n_n5020) & (n_n5047)) + ((n_n5032) & (!n_n5036) & (n_n5021) & (!n_n5020) & (!n_n5047)) + ((n_n5032) & (!n_n5036) & (n_n5021) & (!n_n5020) & (n_n5047)) + ((n_n5032) & (!n_n5036) & (n_n5021) & (n_n5020) & (!n_n5047)) + ((n_n5032) & (!n_n5036) & (n_n5021) & (n_n5020) & (n_n5047)) + ((n_n5032) & (n_n5036) & (!n_n5021) & (!n_n5020) & (!n_n5047)) + ((n_n5032) & (n_n5036) & (!n_n5021) & (!n_n5020) & (n_n5047)) + ((n_n5032) & (n_n5036) & (!n_n5021) & (n_n5020) & (!n_n5047)) + ((n_n5032) & (n_n5036) & (!n_n5021) & (n_n5020) & (n_n5047)) + ((n_n5032) & (n_n5036) & (n_n5021) & (!n_n5020) & (!n_n5047)) + ((n_n5032) & (n_n5036) & (n_n5021) & (!n_n5020) & (n_n5047)) + ((n_n5032) & (n_n5036) & (n_n5021) & (n_n5020) & (!n_n5047)) + ((n_n5032) & (n_n5036) & (n_n5021) & (n_n5020) & (n_n5047)));
	assign x13611x = (((!n_n5156) & (!n_n5191) & (!n_n5175) & (n_n5177)) + ((!n_n5156) & (!n_n5191) & (n_n5175) & (!n_n5177)) + ((!n_n5156) & (!n_n5191) & (n_n5175) & (n_n5177)) + ((!n_n5156) & (n_n5191) & (!n_n5175) & (!n_n5177)) + ((!n_n5156) & (n_n5191) & (!n_n5175) & (n_n5177)) + ((!n_n5156) & (n_n5191) & (n_n5175) & (!n_n5177)) + ((!n_n5156) & (n_n5191) & (n_n5175) & (n_n5177)) + ((n_n5156) & (!n_n5191) & (!n_n5175) & (!n_n5177)) + ((n_n5156) & (!n_n5191) & (!n_n5175) & (n_n5177)) + ((n_n5156) & (!n_n5191) & (n_n5175) & (!n_n5177)) + ((n_n5156) & (!n_n5191) & (n_n5175) & (n_n5177)) + ((n_n5156) & (n_n5191) & (!n_n5175) & (!n_n5177)) + ((n_n5156) & (n_n5191) & (!n_n5175) & (n_n5177)) + ((n_n5156) & (n_n5191) & (n_n5175) & (!n_n5177)) + ((n_n5156) & (n_n5191) & (n_n5175) & (n_n5177)));
	assign x13612x = (((!n_n5171) & (!n_n5190) & (!n_n5170) & (!n_n5194) & (n_n5213)) + ((!n_n5171) & (!n_n5190) & (!n_n5170) & (n_n5194) & (!n_n5213)) + ((!n_n5171) & (!n_n5190) & (!n_n5170) & (n_n5194) & (n_n5213)) + ((!n_n5171) & (!n_n5190) & (n_n5170) & (!n_n5194) & (!n_n5213)) + ((!n_n5171) & (!n_n5190) & (n_n5170) & (!n_n5194) & (n_n5213)) + ((!n_n5171) & (!n_n5190) & (n_n5170) & (n_n5194) & (!n_n5213)) + ((!n_n5171) & (!n_n5190) & (n_n5170) & (n_n5194) & (n_n5213)) + ((!n_n5171) & (n_n5190) & (!n_n5170) & (!n_n5194) & (!n_n5213)) + ((!n_n5171) & (n_n5190) & (!n_n5170) & (!n_n5194) & (n_n5213)) + ((!n_n5171) & (n_n5190) & (!n_n5170) & (n_n5194) & (!n_n5213)) + ((!n_n5171) & (n_n5190) & (!n_n5170) & (n_n5194) & (n_n5213)) + ((!n_n5171) & (n_n5190) & (n_n5170) & (!n_n5194) & (!n_n5213)) + ((!n_n5171) & (n_n5190) & (n_n5170) & (!n_n5194) & (n_n5213)) + ((!n_n5171) & (n_n5190) & (n_n5170) & (n_n5194) & (!n_n5213)) + ((!n_n5171) & (n_n5190) & (n_n5170) & (n_n5194) & (n_n5213)) + ((n_n5171) & (!n_n5190) & (!n_n5170) & (!n_n5194) & (!n_n5213)) + ((n_n5171) & (!n_n5190) & (!n_n5170) & (!n_n5194) & (n_n5213)) + ((n_n5171) & (!n_n5190) & (!n_n5170) & (n_n5194) & (!n_n5213)) + ((n_n5171) & (!n_n5190) & (!n_n5170) & (n_n5194) & (n_n5213)) + ((n_n5171) & (!n_n5190) & (n_n5170) & (!n_n5194) & (!n_n5213)) + ((n_n5171) & (!n_n5190) & (n_n5170) & (!n_n5194) & (n_n5213)) + ((n_n5171) & (!n_n5190) & (n_n5170) & (n_n5194) & (!n_n5213)) + ((n_n5171) & (!n_n5190) & (n_n5170) & (n_n5194) & (n_n5213)) + ((n_n5171) & (n_n5190) & (!n_n5170) & (!n_n5194) & (!n_n5213)) + ((n_n5171) & (n_n5190) & (!n_n5170) & (!n_n5194) & (n_n5213)) + ((n_n5171) & (n_n5190) & (!n_n5170) & (n_n5194) & (!n_n5213)) + ((n_n5171) & (n_n5190) & (!n_n5170) & (n_n5194) & (n_n5213)) + ((n_n5171) & (n_n5190) & (n_n5170) & (!n_n5194) & (!n_n5213)) + ((n_n5171) & (n_n5190) & (n_n5170) & (!n_n5194) & (n_n5213)) + ((n_n5171) & (n_n5190) & (n_n5170) & (n_n5194) & (!n_n5213)) + ((n_n5171) & (n_n5190) & (n_n5170) & (n_n5194) & (n_n5213)));
	assign x13616x = (((!x13606x) & (!x13607x) & (!x13611x) & (x13612x)) + ((!x13606x) & (!x13607x) & (x13611x) & (!x13612x)) + ((!x13606x) & (!x13607x) & (x13611x) & (x13612x)) + ((!x13606x) & (x13607x) & (!x13611x) & (!x13612x)) + ((!x13606x) & (x13607x) & (!x13611x) & (x13612x)) + ((!x13606x) & (x13607x) & (x13611x) & (!x13612x)) + ((!x13606x) & (x13607x) & (x13611x) & (x13612x)) + ((x13606x) & (!x13607x) & (!x13611x) & (!x13612x)) + ((x13606x) & (!x13607x) & (!x13611x) & (x13612x)) + ((x13606x) & (!x13607x) & (x13611x) & (!x13612x)) + ((x13606x) & (!x13607x) & (x13611x) & (x13612x)) + ((x13606x) & (x13607x) & (!x13611x) & (!x13612x)) + ((x13606x) & (x13607x) & (!x13611x) & (x13612x)) + ((x13606x) & (x13607x) & (x13611x) & (!x13612x)) + ((x13606x) & (x13607x) & (x13611x) & (x13612x)));
	assign n_n4392 = (((i_9_) & (n_n536) & (n_n482) & (n_n534)));
	assign n_n4391 = (((i_1_) & (i_2_) & (i_0_) & (n_n491) & (x23x)));
	assign x13623x = (((!n_n4371) & (!n_n4392) & (!n_n4391) & (n_n4399)) + ((!n_n4371) & (!n_n4392) & (n_n4391) & (!n_n4399)) + ((!n_n4371) & (!n_n4392) & (n_n4391) & (n_n4399)) + ((!n_n4371) & (n_n4392) & (!n_n4391) & (!n_n4399)) + ((!n_n4371) & (n_n4392) & (!n_n4391) & (n_n4399)) + ((!n_n4371) & (n_n4392) & (n_n4391) & (!n_n4399)) + ((!n_n4371) & (n_n4392) & (n_n4391) & (n_n4399)) + ((n_n4371) & (!n_n4392) & (!n_n4391) & (!n_n4399)) + ((n_n4371) & (!n_n4392) & (!n_n4391) & (n_n4399)) + ((n_n4371) & (!n_n4392) & (n_n4391) & (!n_n4399)) + ((n_n4371) & (!n_n4392) & (n_n4391) & (n_n4399)) + ((n_n4371) & (n_n4392) & (!n_n4391) & (!n_n4399)) + ((n_n4371) & (n_n4392) & (!n_n4391) & (n_n4399)) + ((n_n4371) & (n_n4392) & (n_n4391) & (!n_n4399)) + ((n_n4371) & (n_n4392) & (n_n4391) & (n_n4399)));
	assign n_n4378 = (((i_9_) & (n_n536) & (n_n532) & (n_n491)));
	assign n_n4388 = (((i_9_) & (n_n536) & (n_n522) & (n_n491)));
	assign n_n4407 = (((i_1_) & (i_2_) & (i_0_) & (n_n482) & (x23x)));
	assign n_n4402 = (((i_9_) & (n_n536) & (n_n524) & (n_n482)));
	assign n_n4408 = (((i_9_) & (n_n536) & (n_n473) & (n_n534)));
	assign x13624x = (((!n_n4378) & (!n_n4388) & (!n_n4407) & (!n_n4402) & (n_n4408)) + ((!n_n4378) & (!n_n4388) & (!n_n4407) & (n_n4402) & (!n_n4408)) + ((!n_n4378) & (!n_n4388) & (!n_n4407) & (n_n4402) & (n_n4408)) + ((!n_n4378) & (!n_n4388) & (n_n4407) & (!n_n4402) & (!n_n4408)) + ((!n_n4378) & (!n_n4388) & (n_n4407) & (!n_n4402) & (n_n4408)) + ((!n_n4378) & (!n_n4388) & (n_n4407) & (n_n4402) & (!n_n4408)) + ((!n_n4378) & (!n_n4388) & (n_n4407) & (n_n4402) & (n_n4408)) + ((!n_n4378) & (n_n4388) & (!n_n4407) & (!n_n4402) & (!n_n4408)) + ((!n_n4378) & (n_n4388) & (!n_n4407) & (!n_n4402) & (n_n4408)) + ((!n_n4378) & (n_n4388) & (!n_n4407) & (n_n4402) & (!n_n4408)) + ((!n_n4378) & (n_n4388) & (!n_n4407) & (n_n4402) & (n_n4408)) + ((!n_n4378) & (n_n4388) & (n_n4407) & (!n_n4402) & (!n_n4408)) + ((!n_n4378) & (n_n4388) & (n_n4407) & (!n_n4402) & (n_n4408)) + ((!n_n4378) & (n_n4388) & (n_n4407) & (n_n4402) & (!n_n4408)) + ((!n_n4378) & (n_n4388) & (n_n4407) & (n_n4402) & (n_n4408)) + ((n_n4378) & (!n_n4388) & (!n_n4407) & (!n_n4402) & (!n_n4408)) + ((n_n4378) & (!n_n4388) & (!n_n4407) & (!n_n4402) & (n_n4408)) + ((n_n4378) & (!n_n4388) & (!n_n4407) & (n_n4402) & (!n_n4408)) + ((n_n4378) & (!n_n4388) & (!n_n4407) & (n_n4402) & (n_n4408)) + ((n_n4378) & (!n_n4388) & (n_n4407) & (!n_n4402) & (!n_n4408)) + ((n_n4378) & (!n_n4388) & (n_n4407) & (!n_n4402) & (n_n4408)) + ((n_n4378) & (!n_n4388) & (n_n4407) & (n_n4402) & (!n_n4408)) + ((n_n4378) & (!n_n4388) & (n_n4407) & (n_n4402) & (n_n4408)) + ((n_n4378) & (n_n4388) & (!n_n4407) & (!n_n4402) & (!n_n4408)) + ((n_n4378) & (n_n4388) & (!n_n4407) & (!n_n4402) & (n_n4408)) + ((n_n4378) & (n_n4388) & (!n_n4407) & (n_n4402) & (!n_n4408)) + ((n_n4378) & (n_n4388) & (!n_n4407) & (n_n4402) & (n_n4408)) + ((n_n4378) & (n_n4388) & (n_n4407) & (!n_n4402) & (!n_n4408)) + ((n_n4378) & (n_n4388) & (n_n4407) & (!n_n4402) & (n_n4408)) + ((n_n4378) & (n_n4388) & (n_n4407) & (n_n4402) & (!n_n4408)) + ((n_n4378) & (n_n4388) & (n_n4407) & (n_n4402) & (n_n4408)));
	assign n_n4748 = (((i_9_) & (n_n325) & (n_n500) & (n_n530)));
	assign n_n4725 = (((!i_5_) & (i_3_) & (i_4_) & (n_n325) & (x20x)));
	assign n_n4788 = (((i_9_) & (n_n482) & (n_n325) & (n_n522)));
	assign n_n4802 = (((i_9_) & (n_n524) & (n_n473) & (n_n325)));
	assign x13644x = (((!n_n4781) & (!n_n4733) & (!n_n4765) & (!n_n4742) & (n_n4808)) + ((!n_n4781) & (!n_n4733) & (!n_n4765) & (n_n4742) & (!n_n4808)) + ((!n_n4781) & (!n_n4733) & (!n_n4765) & (n_n4742) & (n_n4808)) + ((!n_n4781) & (!n_n4733) & (n_n4765) & (!n_n4742) & (!n_n4808)) + ((!n_n4781) & (!n_n4733) & (n_n4765) & (!n_n4742) & (n_n4808)) + ((!n_n4781) & (!n_n4733) & (n_n4765) & (n_n4742) & (!n_n4808)) + ((!n_n4781) & (!n_n4733) & (n_n4765) & (n_n4742) & (n_n4808)) + ((!n_n4781) & (n_n4733) & (!n_n4765) & (!n_n4742) & (!n_n4808)) + ((!n_n4781) & (n_n4733) & (!n_n4765) & (!n_n4742) & (n_n4808)) + ((!n_n4781) & (n_n4733) & (!n_n4765) & (n_n4742) & (!n_n4808)) + ((!n_n4781) & (n_n4733) & (!n_n4765) & (n_n4742) & (n_n4808)) + ((!n_n4781) & (n_n4733) & (n_n4765) & (!n_n4742) & (!n_n4808)) + ((!n_n4781) & (n_n4733) & (n_n4765) & (!n_n4742) & (n_n4808)) + ((!n_n4781) & (n_n4733) & (n_n4765) & (n_n4742) & (!n_n4808)) + ((!n_n4781) & (n_n4733) & (n_n4765) & (n_n4742) & (n_n4808)) + ((n_n4781) & (!n_n4733) & (!n_n4765) & (!n_n4742) & (!n_n4808)) + ((n_n4781) & (!n_n4733) & (!n_n4765) & (!n_n4742) & (n_n4808)) + ((n_n4781) & (!n_n4733) & (!n_n4765) & (n_n4742) & (!n_n4808)) + ((n_n4781) & (!n_n4733) & (!n_n4765) & (n_n4742) & (n_n4808)) + ((n_n4781) & (!n_n4733) & (n_n4765) & (!n_n4742) & (!n_n4808)) + ((n_n4781) & (!n_n4733) & (n_n4765) & (!n_n4742) & (n_n4808)) + ((n_n4781) & (!n_n4733) & (n_n4765) & (n_n4742) & (!n_n4808)) + ((n_n4781) & (!n_n4733) & (n_n4765) & (n_n4742) & (n_n4808)) + ((n_n4781) & (n_n4733) & (!n_n4765) & (!n_n4742) & (!n_n4808)) + ((n_n4781) & (n_n4733) & (!n_n4765) & (!n_n4742) & (n_n4808)) + ((n_n4781) & (n_n4733) & (!n_n4765) & (n_n4742) & (!n_n4808)) + ((n_n4781) & (n_n4733) & (!n_n4765) & (n_n4742) & (n_n4808)) + ((n_n4781) & (n_n4733) & (n_n4765) & (!n_n4742) & (!n_n4808)) + ((n_n4781) & (n_n4733) & (n_n4765) & (!n_n4742) & (n_n4808)) + ((n_n4781) & (n_n4733) & (n_n4765) & (n_n4742) & (!n_n4808)) + ((n_n4781) & (n_n4733) & (n_n4765) & (n_n4742) & (n_n4808)));
	assign x13630x = (((!n_n4663) & (!n_n4665) & (!n_n4672) & (n_n4707)) + ((!n_n4663) & (!n_n4665) & (n_n4672) & (!n_n4707)) + ((!n_n4663) & (!n_n4665) & (n_n4672) & (n_n4707)) + ((!n_n4663) & (n_n4665) & (!n_n4672) & (!n_n4707)) + ((!n_n4663) & (n_n4665) & (!n_n4672) & (n_n4707)) + ((!n_n4663) & (n_n4665) & (n_n4672) & (!n_n4707)) + ((!n_n4663) & (n_n4665) & (n_n4672) & (n_n4707)) + ((n_n4663) & (!n_n4665) & (!n_n4672) & (!n_n4707)) + ((n_n4663) & (!n_n4665) & (!n_n4672) & (n_n4707)) + ((n_n4663) & (!n_n4665) & (n_n4672) & (!n_n4707)) + ((n_n4663) & (!n_n4665) & (n_n4672) & (n_n4707)) + ((n_n4663) & (n_n4665) & (!n_n4672) & (!n_n4707)) + ((n_n4663) & (n_n4665) & (!n_n4672) & (n_n4707)) + ((n_n4663) & (n_n4665) & (n_n4672) & (!n_n4707)) + ((n_n4663) & (n_n4665) & (n_n4672) & (n_n4707)));
	assign x13631x = (((!n_n4724) & (!n_n4679) & (!n_n4701) & (!n_n4692) & (n_n4686)) + ((!n_n4724) & (!n_n4679) & (!n_n4701) & (n_n4692) & (!n_n4686)) + ((!n_n4724) & (!n_n4679) & (!n_n4701) & (n_n4692) & (n_n4686)) + ((!n_n4724) & (!n_n4679) & (n_n4701) & (!n_n4692) & (!n_n4686)) + ((!n_n4724) & (!n_n4679) & (n_n4701) & (!n_n4692) & (n_n4686)) + ((!n_n4724) & (!n_n4679) & (n_n4701) & (n_n4692) & (!n_n4686)) + ((!n_n4724) & (!n_n4679) & (n_n4701) & (n_n4692) & (n_n4686)) + ((!n_n4724) & (n_n4679) & (!n_n4701) & (!n_n4692) & (!n_n4686)) + ((!n_n4724) & (n_n4679) & (!n_n4701) & (!n_n4692) & (n_n4686)) + ((!n_n4724) & (n_n4679) & (!n_n4701) & (n_n4692) & (!n_n4686)) + ((!n_n4724) & (n_n4679) & (!n_n4701) & (n_n4692) & (n_n4686)) + ((!n_n4724) & (n_n4679) & (n_n4701) & (!n_n4692) & (!n_n4686)) + ((!n_n4724) & (n_n4679) & (n_n4701) & (!n_n4692) & (n_n4686)) + ((!n_n4724) & (n_n4679) & (n_n4701) & (n_n4692) & (!n_n4686)) + ((!n_n4724) & (n_n4679) & (n_n4701) & (n_n4692) & (n_n4686)) + ((n_n4724) & (!n_n4679) & (!n_n4701) & (!n_n4692) & (!n_n4686)) + ((n_n4724) & (!n_n4679) & (!n_n4701) & (!n_n4692) & (n_n4686)) + ((n_n4724) & (!n_n4679) & (!n_n4701) & (n_n4692) & (!n_n4686)) + ((n_n4724) & (!n_n4679) & (!n_n4701) & (n_n4692) & (n_n4686)) + ((n_n4724) & (!n_n4679) & (n_n4701) & (!n_n4692) & (!n_n4686)) + ((n_n4724) & (!n_n4679) & (n_n4701) & (!n_n4692) & (n_n4686)) + ((n_n4724) & (!n_n4679) & (n_n4701) & (n_n4692) & (!n_n4686)) + ((n_n4724) & (!n_n4679) & (n_n4701) & (n_n4692) & (n_n4686)) + ((n_n4724) & (n_n4679) & (!n_n4701) & (!n_n4692) & (!n_n4686)) + ((n_n4724) & (n_n4679) & (!n_n4701) & (!n_n4692) & (n_n4686)) + ((n_n4724) & (n_n4679) & (!n_n4701) & (n_n4692) & (!n_n4686)) + ((n_n4724) & (n_n4679) & (!n_n4701) & (n_n4692) & (n_n4686)) + ((n_n4724) & (n_n4679) & (n_n4701) & (!n_n4692) & (!n_n4686)) + ((n_n4724) & (n_n4679) & (n_n4701) & (!n_n4692) & (n_n4686)) + ((n_n4724) & (n_n4679) & (n_n4701) & (n_n4692) & (!n_n4686)) + ((n_n4724) & (n_n4679) & (n_n4701) & (n_n4692) & (n_n4686)));
	assign x13636x = (((!n_n4913) & (!n_n4903) & (!n_n4905) & (n_n4846)) + ((!n_n4913) & (!n_n4903) & (n_n4905) & (!n_n4846)) + ((!n_n4913) & (!n_n4903) & (n_n4905) & (n_n4846)) + ((!n_n4913) & (n_n4903) & (!n_n4905) & (!n_n4846)) + ((!n_n4913) & (n_n4903) & (!n_n4905) & (n_n4846)) + ((!n_n4913) & (n_n4903) & (n_n4905) & (!n_n4846)) + ((!n_n4913) & (n_n4903) & (n_n4905) & (n_n4846)) + ((n_n4913) & (!n_n4903) & (!n_n4905) & (!n_n4846)) + ((n_n4913) & (!n_n4903) & (!n_n4905) & (n_n4846)) + ((n_n4913) & (!n_n4903) & (n_n4905) & (!n_n4846)) + ((n_n4913) & (!n_n4903) & (n_n4905) & (n_n4846)) + ((n_n4913) & (n_n4903) & (!n_n4905) & (!n_n4846)) + ((n_n4913) & (n_n4903) & (!n_n4905) & (n_n4846)) + ((n_n4913) & (n_n4903) & (n_n4905) & (!n_n4846)) + ((n_n4913) & (n_n4903) & (n_n4905) & (n_n4846)));
	assign x13637x = (((!n_n4901) & (!n_n4904) & (!n_n4842) & (!n_n4841) & (n_n4867)) + ((!n_n4901) & (!n_n4904) & (!n_n4842) & (n_n4841) & (!n_n4867)) + ((!n_n4901) & (!n_n4904) & (!n_n4842) & (n_n4841) & (n_n4867)) + ((!n_n4901) & (!n_n4904) & (n_n4842) & (!n_n4841) & (!n_n4867)) + ((!n_n4901) & (!n_n4904) & (n_n4842) & (!n_n4841) & (n_n4867)) + ((!n_n4901) & (!n_n4904) & (n_n4842) & (n_n4841) & (!n_n4867)) + ((!n_n4901) & (!n_n4904) & (n_n4842) & (n_n4841) & (n_n4867)) + ((!n_n4901) & (n_n4904) & (!n_n4842) & (!n_n4841) & (!n_n4867)) + ((!n_n4901) & (n_n4904) & (!n_n4842) & (!n_n4841) & (n_n4867)) + ((!n_n4901) & (n_n4904) & (!n_n4842) & (n_n4841) & (!n_n4867)) + ((!n_n4901) & (n_n4904) & (!n_n4842) & (n_n4841) & (n_n4867)) + ((!n_n4901) & (n_n4904) & (n_n4842) & (!n_n4841) & (!n_n4867)) + ((!n_n4901) & (n_n4904) & (n_n4842) & (!n_n4841) & (n_n4867)) + ((!n_n4901) & (n_n4904) & (n_n4842) & (n_n4841) & (!n_n4867)) + ((!n_n4901) & (n_n4904) & (n_n4842) & (n_n4841) & (n_n4867)) + ((n_n4901) & (!n_n4904) & (!n_n4842) & (!n_n4841) & (!n_n4867)) + ((n_n4901) & (!n_n4904) & (!n_n4842) & (!n_n4841) & (n_n4867)) + ((n_n4901) & (!n_n4904) & (!n_n4842) & (n_n4841) & (!n_n4867)) + ((n_n4901) & (!n_n4904) & (!n_n4842) & (n_n4841) & (n_n4867)) + ((n_n4901) & (!n_n4904) & (n_n4842) & (!n_n4841) & (!n_n4867)) + ((n_n4901) & (!n_n4904) & (n_n4842) & (!n_n4841) & (n_n4867)) + ((n_n4901) & (!n_n4904) & (n_n4842) & (n_n4841) & (!n_n4867)) + ((n_n4901) & (!n_n4904) & (n_n4842) & (n_n4841) & (n_n4867)) + ((n_n4901) & (n_n4904) & (!n_n4842) & (!n_n4841) & (!n_n4867)) + ((n_n4901) & (n_n4904) & (!n_n4842) & (!n_n4841) & (n_n4867)) + ((n_n4901) & (n_n4904) & (!n_n4842) & (n_n4841) & (!n_n4867)) + ((n_n4901) & (n_n4904) & (!n_n4842) & (n_n4841) & (n_n4867)) + ((n_n4901) & (n_n4904) & (n_n4842) & (!n_n4841) & (!n_n4867)) + ((n_n4901) & (n_n4904) & (n_n4842) & (!n_n4841) & (n_n4867)) + ((n_n4901) & (n_n4904) & (n_n4842) & (n_n4841) & (!n_n4867)) + ((n_n4901) & (n_n4904) & (n_n4842) & (n_n4841) & (n_n4867)));
	assign x13650x = (((!i_9_) & (!n_n534) & (!n_n4570) & (!x523x) & (x214x)) + ((!i_9_) & (!n_n534) & (!n_n4570) & (x523x) & (x214x)) + ((!i_9_) & (!n_n534) & (n_n4570) & (!x523x) & (!x214x)) + ((!i_9_) & (!n_n534) & (n_n4570) & (!x523x) & (x214x)) + ((!i_9_) & (!n_n534) & (n_n4570) & (x523x) & (!x214x)) + ((!i_9_) & (!n_n534) & (n_n4570) & (x523x) & (x214x)) + ((!i_9_) & (n_n534) & (!n_n4570) & (!x523x) & (x214x)) + ((!i_9_) & (n_n534) & (!n_n4570) & (x523x) & (!x214x)) + ((!i_9_) & (n_n534) & (!n_n4570) & (x523x) & (x214x)) + ((!i_9_) & (n_n534) & (n_n4570) & (!x523x) & (!x214x)) + ((!i_9_) & (n_n534) & (n_n4570) & (!x523x) & (x214x)) + ((!i_9_) & (n_n534) & (n_n4570) & (x523x) & (!x214x)) + ((!i_9_) & (n_n534) & (n_n4570) & (x523x) & (x214x)) + ((i_9_) & (!n_n534) & (!n_n4570) & (!x523x) & (x214x)) + ((i_9_) & (!n_n534) & (!n_n4570) & (x523x) & (x214x)) + ((i_9_) & (!n_n534) & (n_n4570) & (!x523x) & (!x214x)) + ((i_9_) & (!n_n534) & (n_n4570) & (!x523x) & (x214x)) + ((i_9_) & (!n_n534) & (n_n4570) & (x523x) & (!x214x)) + ((i_9_) & (!n_n534) & (n_n4570) & (x523x) & (x214x)) + ((i_9_) & (n_n534) & (!n_n4570) & (!x523x) & (x214x)) + ((i_9_) & (n_n534) & (!n_n4570) & (x523x) & (x214x)) + ((i_9_) & (n_n534) & (n_n4570) & (!x523x) & (!x214x)) + ((i_9_) & (n_n534) & (n_n4570) & (!x523x) & (x214x)) + ((i_9_) & (n_n534) & (n_n4570) & (x523x) & (!x214x)) + ((i_9_) & (n_n534) & (n_n4570) & (x523x) & (x214x)));
	assign x13651x = (((!n_n4576) & (!n_n4549) & (!n_n4551) & (!n_n4552) & (n_n4580)) + ((!n_n4576) & (!n_n4549) & (!n_n4551) & (n_n4552) & (!n_n4580)) + ((!n_n4576) & (!n_n4549) & (!n_n4551) & (n_n4552) & (n_n4580)) + ((!n_n4576) & (!n_n4549) & (n_n4551) & (!n_n4552) & (!n_n4580)) + ((!n_n4576) & (!n_n4549) & (n_n4551) & (!n_n4552) & (n_n4580)) + ((!n_n4576) & (!n_n4549) & (n_n4551) & (n_n4552) & (!n_n4580)) + ((!n_n4576) & (!n_n4549) & (n_n4551) & (n_n4552) & (n_n4580)) + ((!n_n4576) & (n_n4549) & (!n_n4551) & (!n_n4552) & (!n_n4580)) + ((!n_n4576) & (n_n4549) & (!n_n4551) & (!n_n4552) & (n_n4580)) + ((!n_n4576) & (n_n4549) & (!n_n4551) & (n_n4552) & (!n_n4580)) + ((!n_n4576) & (n_n4549) & (!n_n4551) & (n_n4552) & (n_n4580)) + ((!n_n4576) & (n_n4549) & (n_n4551) & (!n_n4552) & (!n_n4580)) + ((!n_n4576) & (n_n4549) & (n_n4551) & (!n_n4552) & (n_n4580)) + ((!n_n4576) & (n_n4549) & (n_n4551) & (n_n4552) & (!n_n4580)) + ((!n_n4576) & (n_n4549) & (n_n4551) & (n_n4552) & (n_n4580)) + ((n_n4576) & (!n_n4549) & (!n_n4551) & (!n_n4552) & (!n_n4580)) + ((n_n4576) & (!n_n4549) & (!n_n4551) & (!n_n4552) & (n_n4580)) + ((n_n4576) & (!n_n4549) & (!n_n4551) & (n_n4552) & (!n_n4580)) + ((n_n4576) & (!n_n4549) & (!n_n4551) & (n_n4552) & (n_n4580)) + ((n_n4576) & (!n_n4549) & (n_n4551) & (!n_n4552) & (!n_n4580)) + ((n_n4576) & (!n_n4549) & (n_n4551) & (!n_n4552) & (n_n4580)) + ((n_n4576) & (!n_n4549) & (n_n4551) & (n_n4552) & (!n_n4580)) + ((n_n4576) & (!n_n4549) & (n_n4551) & (n_n4552) & (n_n4580)) + ((n_n4576) & (n_n4549) & (!n_n4551) & (!n_n4552) & (!n_n4580)) + ((n_n4576) & (n_n4549) & (!n_n4551) & (!n_n4552) & (n_n4580)) + ((n_n4576) & (n_n4549) & (!n_n4551) & (n_n4552) & (!n_n4580)) + ((n_n4576) & (n_n4549) & (!n_n4551) & (n_n4552) & (n_n4580)) + ((n_n4576) & (n_n4549) & (n_n4551) & (!n_n4552) & (!n_n4580)) + ((n_n4576) & (n_n4549) & (n_n4551) & (!n_n4552) & (n_n4580)) + ((n_n4576) & (n_n4549) & (n_n4551) & (n_n4552) & (!n_n4580)) + ((n_n4576) & (n_n4549) & (n_n4551) & (n_n4552) & (n_n4580)));
	assign n_n3932 = (((!n_n4617) & (!n_n4637) & (!n_n4613) & (!n_n4602) & (x13657x)) + ((!n_n4617) & (!n_n4637) & (!n_n4613) & (n_n4602) & (!x13657x)) + ((!n_n4617) & (!n_n4637) & (!n_n4613) & (n_n4602) & (x13657x)) + ((!n_n4617) & (!n_n4637) & (n_n4613) & (!n_n4602) & (!x13657x)) + ((!n_n4617) & (!n_n4637) & (n_n4613) & (!n_n4602) & (x13657x)) + ((!n_n4617) & (!n_n4637) & (n_n4613) & (n_n4602) & (!x13657x)) + ((!n_n4617) & (!n_n4637) & (n_n4613) & (n_n4602) & (x13657x)) + ((!n_n4617) & (n_n4637) & (!n_n4613) & (!n_n4602) & (!x13657x)) + ((!n_n4617) & (n_n4637) & (!n_n4613) & (!n_n4602) & (x13657x)) + ((!n_n4617) & (n_n4637) & (!n_n4613) & (n_n4602) & (!x13657x)) + ((!n_n4617) & (n_n4637) & (!n_n4613) & (n_n4602) & (x13657x)) + ((!n_n4617) & (n_n4637) & (n_n4613) & (!n_n4602) & (!x13657x)) + ((!n_n4617) & (n_n4637) & (n_n4613) & (!n_n4602) & (x13657x)) + ((!n_n4617) & (n_n4637) & (n_n4613) & (n_n4602) & (!x13657x)) + ((!n_n4617) & (n_n4637) & (n_n4613) & (n_n4602) & (x13657x)) + ((n_n4617) & (!n_n4637) & (!n_n4613) & (!n_n4602) & (!x13657x)) + ((n_n4617) & (!n_n4637) & (!n_n4613) & (!n_n4602) & (x13657x)) + ((n_n4617) & (!n_n4637) & (!n_n4613) & (n_n4602) & (!x13657x)) + ((n_n4617) & (!n_n4637) & (!n_n4613) & (n_n4602) & (x13657x)) + ((n_n4617) & (!n_n4637) & (n_n4613) & (!n_n4602) & (!x13657x)) + ((n_n4617) & (!n_n4637) & (n_n4613) & (!n_n4602) & (x13657x)) + ((n_n4617) & (!n_n4637) & (n_n4613) & (n_n4602) & (!x13657x)) + ((n_n4617) & (!n_n4637) & (n_n4613) & (n_n4602) & (x13657x)) + ((n_n4617) & (n_n4637) & (!n_n4613) & (!n_n4602) & (!x13657x)) + ((n_n4617) & (n_n4637) & (!n_n4613) & (!n_n4602) & (x13657x)) + ((n_n4617) & (n_n4637) & (!n_n4613) & (n_n4602) & (!x13657x)) + ((n_n4617) & (n_n4637) & (!n_n4613) & (n_n4602) & (x13657x)) + ((n_n4617) & (n_n4637) & (n_n4613) & (!n_n4602) & (!x13657x)) + ((n_n4617) & (n_n4637) & (n_n4613) & (!n_n4602) & (x13657x)) + ((n_n4617) & (n_n4637) & (n_n4613) & (n_n4602) & (!x13657x)) + ((n_n4617) & (n_n4637) & (n_n4613) & (n_n4602) & (x13657x)));
	assign x13663x = (((!n_n4504) & (!n_n4535) & (!n_n4507) & (n_n4509)) + ((!n_n4504) & (!n_n4535) & (n_n4507) & (!n_n4509)) + ((!n_n4504) & (!n_n4535) & (n_n4507) & (n_n4509)) + ((!n_n4504) & (n_n4535) & (!n_n4507) & (!n_n4509)) + ((!n_n4504) & (n_n4535) & (!n_n4507) & (n_n4509)) + ((!n_n4504) & (n_n4535) & (n_n4507) & (!n_n4509)) + ((!n_n4504) & (n_n4535) & (n_n4507) & (n_n4509)) + ((n_n4504) & (!n_n4535) & (!n_n4507) & (!n_n4509)) + ((n_n4504) & (!n_n4535) & (!n_n4507) & (n_n4509)) + ((n_n4504) & (!n_n4535) & (n_n4507) & (!n_n4509)) + ((n_n4504) & (!n_n4535) & (n_n4507) & (n_n4509)) + ((n_n4504) & (n_n4535) & (!n_n4507) & (!n_n4509)) + ((n_n4504) & (n_n4535) & (!n_n4507) & (n_n4509)) + ((n_n4504) & (n_n4535) & (n_n4507) & (!n_n4509)) + ((n_n4504) & (n_n4535) & (n_n4507) & (n_n4509)));
	assign x13664x = (((!n_n4521) & (!n_n4544) & (!n_n4498) & (!n_n4540) & (n_n4520)) + ((!n_n4521) & (!n_n4544) & (!n_n4498) & (n_n4540) & (!n_n4520)) + ((!n_n4521) & (!n_n4544) & (!n_n4498) & (n_n4540) & (n_n4520)) + ((!n_n4521) & (!n_n4544) & (n_n4498) & (!n_n4540) & (!n_n4520)) + ((!n_n4521) & (!n_n4544) & (n_n4498) & (!n_n4540) & (n_n4520)) + ((!n_n4521) & (!n_n4544) & (n_n4498) & (n_n4540) & (!n_n4520)) + ((!n_n4521) & (!n_n4544) & (n_n4498) & (n_n4540) & (n_n4520)) + ((!n_n4521) & (n_n4544) & (!n_n4498) & (!n_n4540) & (!n_n4520)) + ((!n_n4521) & (n_n4544) & (!n_n4498) & (!n_n4540) & (n_n4520)) + ((!n_n4521) & (n_n4544) & (!n_n4498) & (n_n4540) & (!n_n4520)) + ((!n_n4521) & (n_n4544) & (!n_n4498) & (n_n4540) & (n_n4520)) + ((!n_n4521) & (n_n4544) & (n_n4498) & (!n_n4540) & (!n_n4520)) + ((!n_n4521) & (n_n4544) & (n_n4498) & (!n_n4540) & (n_n4520)) + ((!n_n4521) & (n_n4544) & (n_n4498) & (n_n4540) & (!n_n4520)) + ((!n_n4521) & (n_n4544) & (n_n4498) & (n_n4540) & (n_n4520)) + ((n_n4521) & (!n_n4544) & (!n_n4498) & (!n_n4540) & (!n_n4520)) + ((n_n4521) & (!n_n4544) & (!n_n4498) & (!n_n4540) & (n_n4520)) + ((n_n4521) & (!n_n4544) & (!n_n4498) & (n_n4540) & (!n_n4520)) + ((n_n4521) & (!n_n4544) & (!n_n4498) & (n_n4540) & (n_n4520)) + ((n_n4521) & (!n_n4544) & (n_n4498) & (!n_n4540) & (!n_n4520)) + ((n_n4521) & (!n_n4544) & (n_n4498) & (!n_n4540) & (n_n4520)) + ((n_n4521) & (!n_n4544) & (n_n4498) & (n_n4540) & (!n_n4520)) + ((n_n4521) & (!n_n4544) & (n_n4498) & (n_n4540) & (n_n4520)) + ((n_n4521) & (n_n4544) & (!n_n4498) & (!n_n4540) & (!n_n4520)) + ((n_n4521) & (n_n4544) & (!n_n4498) & (!n_n4540) & (n_n4520)) + ((n_n4521) & (n_n4544) & (!n_n4498) & (n_n4540) & (!n_n4520)) + ((n_n4521) & (n_n4544) & (!n_n4498) & (n_n4540) & (n_n4520)) + ((n_n4521) & (n_n4544) & (n_n4498) & (!n_n4540) & (!n_n4520)) + ((n_n4521) & (n_n4544) & (n_n4498) & (!n_n4540) & (n_n4520)) + ((n_n4521) & (n_n4544) & (n_n4498) & (n_n4540) & (!n_n4520)) + ((n_n4521) & (n_n4544) & (n_n4498) & (n_n4540) & (n_n4520)));
	assign n_n4470 = (((i_9_) & (n_n518) & (n_n455) & (n_n520)));
	assign n_n4413 = (((!i_9_) & (n_n536) & (n_n473) & (n_n530)));
	assign n_n4457 = (((!i_9_) & (n_n518) & (n_n455) & (n_n534)));
	assign x13672x = (((!n_n4470) & (!n_n4473) & (!n_n4413) & (n_n4457)) + ((!n_n4470) & (!n_n4473) & (n_n4413) & (!n_n4457)) + ((!n_n4470) & (!n_n4473) & (n_n4413) & (n_n4457)) + ((!n_n4470) & (n_n4473) & (!n_n4413) & (!n_n4457)) + ((!n_n4470) & (n_n4473) & (!n_n4413) & (n_n4457)) + ((!n_n4470) & (n_n4473) & (n_n4413) & (!n_n4457)) + ((!n_n4470) & (n_n4473) & (n_n4413) & (n_n4457)) + ((n_n4470) & (!n_n4473) & (!n_n4413) & (!n_n4457)) + ((n_n4470) & (!n_n4473) & (!n_n4413) & (n_n4457)) + ((n_n4470) & (!n_n4473) & (n_n4413) & (!n_n4457)) + ((n_n4470) & (!n_n4473) & (n_n4413) & (n_n4457)) + ((n_n4470) & (n_n4473) & (!n_n4413) & (!n_n4457)) + ((n_n4470) & (n_n4473) & (!n_n4413) & (n_n4457)) + ((n_n4470) & (n_n4473) & (n_n4413) & (!n_n4457)) + ((n_n4470) & (n_n4473) & (n_n4413) & (n_n4457)));
	assign n_n4459 = (((!i_9_) & (n_n518) & (n_n455) & (n_n532)));
	assign n_n4420 = (((i_9_) & (n_n536) & (n_n473) & (n_n522)));
	assign n_n4472 = (((i_9_) & (n_n455) & (n_n534) & (n_n509)));
	assign n_n4480 = (((i_9_) & (n_n526) & (n_n455) & (n_n509)));
	assign n_n4410 = (((i_9_) & (n_n536) & (n_n473) & (n_n532)));
	assign x13673x = (((!n_n4459) & (!n_n4420) & (!n_n4472) & (!n_n4480) & (n_n4410)) + ((!n_n4459) & (!n_n4420) & (!n_n4472) & (n_n4480) & (!n_n4410)) + ((!n_n4459) & (!n_n4420) & (!n_n4472) & (n_n4480) & (n_n4410)) + ((!n_n4459) & (!n_n4420) & (n_n4472) & (!n_n4480) & (!n_n4410)) + ((!n_n4459) & (!n_n4420) & (n_n4472) & (!n_n4480) & (n_n4410)) + ((!n_n4459) & (!n_n4420) & (n_n4472) & (n_n4480) & (!n_n4410)) + ((!n_n4459) & (!n_n4420) & (n_n4472) & (n_n4480) & (n_n4410)) + ((!n_n4459) & (n_n4420) & (!n_n4472) & (!n_n4480) & (!n_n4410)) + ((!n_n4459) & (n_n4420) & (!n_n4472) & (!n_n4480) & (n_n4410)) + ((!n_n4459) & (n_n4420) & (!n_n4472) & (n_n4480) & (!n_n4410)) + ((!n_n4459) & (n_n4420) & (!n_n4472) & (n_n4480) & (n_n4410)) + ((!n_n4459) & (n_n4420) & (n_n4472) & (!n_n4480) & (!n_n4410)) + ((!n_n4459) & (n_n4420) & (n_n4472) & (!n_n4480) & (n_n4410)) + ((!n_n4459) & (n_n4420) & (n_n4472) & (n_n4480) & (!n_n4410)) + ((!n_n4459) & (n_n4420) & (n_n4472) & (n_n4480) & (n_n4410)) + ((n_n4459) & (!n_n4420) & (!n_n4472) & (!n_n4480) & (!n_n4410)) + ((n_n4459) & (!n_n4420) & (!n_n4472) & (!n_n4480) & (n_n4410)) + ((n_n4459) & (!n_n4420) & (!n_n4472) & (n_n4480) & (!n_n4410)) + ((n_n4459) & (!n_n4420) & (!n_n4472) & (n_n4480) & (n_n4410)) + ((n_n4459) & (!n_n4420) & (n_n4472) & (!n_n4480) & (!n_n4410)) + ((n_n4459) & (!n_n4420) & (n_n4472) & (!n_n4480) & (n_n4410)) + ((n_n4459) & (!n_n4420) & (n_n4472) & (n_n4480) & (!n_n4410)) + ((n_n4459) & (!n_n4420) & (n_n4472) & (n_n4480) & (n_n4410)) + ((n_n4459) & (n_n4420) & (!n_n4472) & (!n_n4480) & (!n_n4410)) + ((n_n4459) & (n_n4420) & (!n_n4472) & (!n_n4480) & (n_n4410)) + ((n_n4459) & (n_n4420) & (!n_n4472) & (n_n4480) & (!n_n4410)) + ((n_n4459) & (n_n4420) & (!n_n4472) & (n_n4480) & (n_n4410)) + ((n_n4459) & (n_n4420) & (n_n4472) & (!n_n4480) & (!n_n4410)) + ((n_n4459) & (n_n4420) & (n_n4472) & (!n_n4480) & (n_n4410)) + ((n_n4459) & (n_n4420) & (n_n4472) & (n_n4480) & (!n_n4410)) + ((n_n4459) & (n_n4420) & (n_n4472) & (n_n4480) & (n_n4410)));
	assign n_n4340 = (((i_9_) & (n_n536) & (n_n518) & (n_n522)));
	assign n_n4368 = (((i_9_) & (n_n536) & (n_n526) & (n_n500)));
	assign n_n4341 = (((i_1_) & (i_2_) & (i_0_) & (n_n518) & (x20x)));
	assign n_n4358 = (((i_9_) & (n_n536) & (n_n509) & (n_n520)));
	assign n_n4354 = (((i_9_) & (n_n536) & (n_n524) & (n_n509)));
	assign x13679x = (((!n_n4340) & (!n_n4368) & (!n_n4341) & (!n_n4358) & (n_n4354)) + ((!n_n4340) & (!n_n4368) & (!n_n4341) & (n_n4358) & (!n_n4354)) + ((!n_n4340) & (!n_n4368) & (!n_n4341) & (n_n4358) & (n_n4354)) + ((!n_n4340) & (!n_n4368) & (n_n4341) & (!n_n4358) & (!n_n4354)) + ((!n_n4340) & (!n_n4368) & (n_n4341) & (!n_n4358) & (n_n4354)) + ((!n_n4340) & (!n_n4368) & (n_n4341) & (n_n4358) & (!n_n4354)) + ((!n_n4340) & (!n_n4368) & (n_n4341) & (n_n4358) & (n_n4354)) + ((!n_n4340) & (n_n4368) & (!n_n4341) & (!n_n4358) & (!n_n4354)) + ((!n_n4340) & (n_n4368) & (!n_n4341) & (!n_n4358) & (n_n4354)) + ((!n_n4340) & (n_n4368) & (!n_n4341) & (n_n4358) & (!n_n4354)) + ((!n_n4340) & (n_n4368) & (!n_n4341) & (n_n4358) & (n_n4354)) + ((!n_n4340) & (n_n4368) & (n_n4341) & (!n_n4358) & (!n_n4354)) + ((!n_n4340) & (n_n4368) & (n_n4341) & (!n_n4358) & (n_n4354)) + ((!n_n4340) & (n_n4368) & (n_n4341) & (n_n4358) & (!n_n4354)) + ((!n_n4340) & (n_n4368) & (n_n4341) & (n_n4358) & (n_n4354)) + ((n_n4340) & (!n_n4368) & (!n_n4341) & (!n_n4358) & (!n_n4354)) + ((n_n4340) & (!n_n4368) & (!n_n4341) & (!n_n4358) & (n_n4354)) + ((n_n4340) & (!n_n4368) & (!n_n4341) & (n_n4358) & (!n_n4354)) + ((n_n4340) & (!n_n4368) & (!n_n4341) & (n_n4358) & (n_n4354)) + ((n_n4340) & (!n_n4368) & (n_n4341) & (!n_n4358) & (!n_n4354)) + ((n_n4340) & (!n_n4368) & (n_n4341) & (!n_n4358) & (n_n4354)) + ((n_n4340) & (!n_n4368) & (n_n4341) & (n_n4358) & (!n_n4354)) + ((n_n4340) & (!n_n4368) & (n_n4341) & (n_n4358) & (n_n4354)) + ((n_n4340) & (n_n4368) & (!n_n4341) & (!n_n4358) & (!n_n4354)) + ((n_n4340) & (n_n4368) & (!n_n4341) & (!n_n4358) & (n_n4354)) + ((n_n4340) & (n_n4368) & (!n_n4341) & (n_n4358) & (!n_n4354)) + ((n_n4340) & (n_n4368) & (!n_n4341) & (n_n4358) & (n_n4354)) + ((n_n4340) & (n_n4368) & (n_n4341) & (!n_n4358) & (!n_n4354)) + ((n_n4340) & (n_n4368) & (n_n4341) & (!n_n4358) & (n_n4354)) + ((n_n4340) & (n_n4368) & (n_n4341) & (n_n4358) & (!n_n4354)) + ((n_n4340) & (n_n4368) & (n_n4341) & (n_n4358) & (n_n4354)));
	assign n_n4325 = (((i_1_) & (i_2_) & (i_0_) & (n_n535) & (x20x)));
	assign n_n4317 = (((!i_9_) & (n_n536) & (n_n535) & (n_n530)));
	assign n_n4362 = (((i_9_) & (n_n536) & (n_n532) & (n_n500)));
	assign n_n4312 = (((i_9_) & (n_n536) & (n_n534) & (n_n535)));
	assign n_n3937 = (((!x13679x) & (!n_n4325) & (!n_n4317) & (!n_n4362) & (n_n4312)) + ((!x13679x) & (!n_n4325) & (!n_n4317) & (n_n4362) & (!n_n4312)) + ((!x13679x) & (!n_n4325) & (!n_n4317) & (n_n4362) & (n_n4312)) + ((!x13679x) & (!n_n4325) & (n_n4317) & (!n_n4362) & (!n_n4312)) + ((!x13679x) & (!n_n4325) & (n_n4317) & (!n_n4362) & (n_n4312)) + ((!x13679x) & (!n_n4325) & (n_n4317) & (n_n4362) & (!n_n4312)) + ((!x13679x) & (!n_n4325) & (n_n4317) & (n_n4362) & (n_n4312)) + ((!x13679x) & (n_n4325) & (!n_n4317) & (!n_n4362) & (!n_n4312)) + ((!x13679x) & (n_n4325) & (!n_n4317) & (!n_n4362) & (n_n4312)) + ((!x13679x) & (n_n4325) & (!n_n4317) & (n_n4362) & (!n_n4312)) + ((!x13679x) & (n_n4325) & (!n_n4317) & (n_n4362) & (n_n4312)) + ((!x13679x) & (n_n4325) & (n_n4317) & (!n_n4362) & (!n_n4312)) + ((!x13679x) & (n_n4325) & (n_n4317) & (!n_n4362) & (n_n4312)) + ((!x13679x) & (n_n4325) & (n_n4317) & (n_n4362) & (!n_n4312)) + ((!x13679x) & (n_n4325) & (n_n4317) & (n_n4362) & (n_n4312)) + ((x13679x) & (!n_n4325) & (!n_n4317) & (!n_n4362) & (!n_n4312)) + ((x13679x) & (!n_n4325) & (!n_n4317) & (!n_n4362) & (n_n4312)) + ((x13679x) & (!n_n4325) & (!n_n4317) & (n_n4362) & (!n_n4312)) + ((x13679x) & (!n_n4325) & (!n_n4317) & (n_n4362) & (n_n4312)) + ((x13679x) & (!n_n4325) & (n_n4317) & (!n_n4362) & (!n_n4312)) + ((x13679x) & (!n_n4325) & (n_n4317) & (!n_n4362) & (n_n4312)) + ((x13679x) & (!n_n4325) & (n_n4317) & (n_n4362) & (!n_n4312)) + ((x13679x) & (!n_n4325) & (n_n4317) & (n_n4362) & (n_n4312)) + ((x13679x) & (n_n4325) & (!n_n4317) & (!n_n4362) & (!n_n4312)) + ((x13679x) & (n_n4325) & (!n_n4317) & (!n_n4362) & (n_n4312)) + ((x13679x) & (n_n4325) & (!n_n4317) & (n_n4362) & (!n_n4312)) + ((x13679x) & (n_n4325) & (!n_n4317) & (n_n4362) & (n_n4312)) + ((x13679x) & (n_n4325) & (n_n4317) & (!n_n4362) & (!n_n4312)) + ((x13679x) & (n_n4325) & (n_n4317) & (!n_n4362) & (n_n4312)) + ((x13679x) & (n_n4325) & (n_n4317) & (n_n4362) & (!n_n4312)) + ((x13679x) & (n_n4325) & (n_n4317) & (n_n4362) & (n_n4312)));
	assign n_n4339 = (((!i_9_) & (n_n536) & (n_n524) & (n_n518)));
	assign n_n4401 = (((!i_9_) & (n_n536) & (n_n526) & (n_n482)));
	assign n_n4314 = (((i_9_) & (n_n536) & (n_n532) & (n_n535)));
	assign n_n4389 = (((i_1_) & (i_2_) & (i_0_) & (n_n491) & (x20x)));
	assign x13689x = (((!n_n4339) & (!n_n4401) & (!n_n4314) & (n_n4389)) + ((!n_n4339) & (!n_n4401) & (n_n4314) & (!n_n4389)) + ((!n_n4339) & (!n_n4401) & (n_n4314) & (n_n4389)) + ((!n_n4339) & (n_n4401) & (!n_n4314) & (!n_n4389)) + ((!n_n4339) & (n_n4401) & (!n_n4314) & (n_n4389)) + ((!n_n4339) & (n_n4401) & (n_n4314) & (!n_n4389)) + ((!n_n4339) & (n_n4401) & (n_n4314) & (n_n4389)) + ((n_n4339) & (!n_n4401) & (!n_n4314) & (!n_n4389)) + ((n_n4339) & (!n_n4401) & (!n_n4314) & (n_n4389)) + ((n_n4339) & (!n_n4401) & (n_n4314) & (!n_n4389)) + ((n_n4339) & (!n_n4401) & (n_n4314) & (n_n4389)) + ((n_n4339) & (n_n4401) & (!n_n4314) & (!n_n4389)) + ((n_n4339) & (n_n4401) & (!n_n4314) & (n_n4389)) + ((n_n4339) & (n_n4401) & (n_n4314) & (!n_n4389)) + ((n_n4339) & (n_n4401) & (n_n4314) & (n_n4389)));
	assign n_n4369 = (((!i_9_) & (n_n536) & (n_n526) & (n_n500)));
	assign n_n4381 = (((!i_9_) & (n_n536) & (n_n491) & (n_n530)));
	assign x13690x = (((!n_n4369) & (!n_n4381) & (!n_n4340) & (!n_n4379) & (n_n4378)) + ((!n_n4369) & (!n_n4381) & (!n_n4340) & (n_n4379) & (!n_n4378)) + ((!n_n4369) & (!n_n4381) & (!n_n4340) & (n_n4379) & (n_n4378)) + ((!n_n4369) & (!n_n4381) & (n_n4340) & (!n_n4379) & (!n_n4378)) + ((!n_n4369) & (!n_n4381) & (n_n4340) & (!n_n4379) & (n_n4378)) + ((!n_n4369) & (!n_n4381) & (n_n4340) & (n_n4379) & (!n_n4378)) + ((!n_n4369) & (!n_n4381) & (n_n4340) & (n_n4379) & (n_n4378)) + ((!n_n4369) & (n_n4381) & (!n_n4340) & (!n_n4379) & (!n_n4378)) + ((!n_n4369) & (n_n4381) & (!n_n4340) & (!n_n4379) & (n_n4378)) + ((!n_n4369) & (n_n4381) & (!n_n4340) & (n_n4379) & (!n_n4378)) + ((!n_n4369) & (n_n4381) & (!n_n4340) & (n_n4379) & (n_n4378)) + ((!n_n4369) & (n_n4381) & (n_n4340) & (!n_n4379) & (!n_n4378)) + ((!n_n4369) & (n_n4381) & (n_n4340) & (!n_n4379) & (n_n4378)) + ((!n_n4369) & (n_n4381) & (n_n4340) & (n_n4379) & (!n_n4378)) + ((!n_n4369) & (n_n4381) & (n_n4340) & (n_n4379) & (n_n4378)) + ((n_n4369) & (!n_n4381) & (!n_n4340) & (!n_n4379) & (!n_n4378)) + ((n_n4369) & (!n_n4381) & (!n_n4340) & (!n_n4379) & (n_n4378)) + ((n_n4369) & (!n_n4381) & (!n_n4340) & (n_n4379) & (!n_n4378)) + ((n_n4369) & (!n_n4381) & (!n_n4340) & (n_n4379) & (n_n4378)) + ((n_n4369) & (!n_n4381) & (n_n4340) & (!n_n4379) & (!n_n4378)) + ((n_n4369) & (!n_n4381) & (n_n4340) & (!n_n4379) & (n_n4378)) + ((n_n4369) & (!n_n4381) & (n_n4340) & (n_n4379) & (!n_n4378)) + ((n_n4369) & (!n_n4381) & (n_n4340) & (n_n4379) & (n_n4378)) + ((n_n4369) & (n_n4381) & (!n_n4340) & (!n_n4379) & (!n_n4378)) + ((n_n4369) & (n_n4381) & (!n_n4340) & (!n_n4379) & (n_n4378)) + ((n_n4369) & (n_n4381) & (!n_n4340) & (n_n4379) & (!n_n4378)) + ((n_n4369) & (n_n4381) & (!n_n4340) & (n_n4379) & (n_n4378)) + ((n_n4369) & (n_n4381) & (n_n4340) & (!n_n4379) & (!n_n4378)) + ((n_n4369) & (n_n4381) & (n_n4340) & (!n_n4379) & (n_n4378)) + ((n_n4369) & (n_n4381) & (n_n4340) & (n_n4379) & (!n_n4378)) + ((n_n4369) & (n_n4381) & (n_n4340) & (n_n4379) & (n_n4378)));
	assign x13703x = (((!n_n5182) & (!n_n5173) & (!n_n5165) & (n_n5230)) + ((!n_n5182) & (!n_n5173) & (n_n5165) & (!n_n5230)) + ((!n_n5182) & (!n_n5173) & (n_n5165) & (n_n5230)) + ((!n_n5182) & (n_n5173) & (!n_n5165) & (!n_n5230)) + ((!n_n5182) & (n_n5173) & (!n_n5165) & (n_n5230)) + ((!n_n5182) & (n_n5173) & (n_n5165) & (!n_n5230)) + ((!n_n5182) & (n_n5173) & (n_n5165) & (n_n5230)) + ((n_n5182) & (!n_n5173) & (!n_n5165) & (!n_n5230)) + ((n_n5182) & (!n_n5173) & (!n_n5165) & (n_n5230)) + ((n_n5182) & (!n_n5173) & (n_n5165) & (!n_n5230)) + ((n_n5182) & (!n_n5173) & (n_n5165) & (n_n5230)) + ((n_n5182) & (n_n5173) & (!n_n5165) & (!n_n5230)) + ((n_n5182) & (n_n5173) & (!n_n5165) & (n_n5230)) + ((n_n5182) & (n_n5173) & (n_n5165) & (!n_n5230)) + ((n_n5182) & (n_n5173) & (n_n5165) & (n_n5230)));
	assign x13704x = (((!n_n5239) & (!n_n5238) & (!n_n5166) & (!n_n5163) & (n_n5214)) + ((!n_n5239) & (!n_n5238) & (!n_n5166) & (n_n5163) & (!n_n5214)) + ((!n_n5239) & (!n_n5238) & (!n_n5166) & (n_n5163) & (n_n5214)) + ((!n_n5239) & (!n_n5238) & (n_n5166) & (!n_n5163) & (!n_n5214)) + ((!n_n5239) & (!n_n5238) & (n_n5166) & (!n_n5163) & (n_n5214)) + ((!n_n5239) & (!n_n5238) & (n_n5166) & (n_n5163) & (!n_n5214)) + ((!n_n5239) & (!n_n5238) & (n_n5166) & (n_n5163) & (n_n5214)) + ((!n_n5239) & (n_n5238) & (!n_n5166) & (!n_n5163) & (!n_n5214)) + ((!n_n5239) & (n_n5238) & (!n_n5166) & (!n_n5163) & (n_n5214)) + ((!n_n5239) & (n_n5238) & (!n_n5166) & (n_n5163) & (!n_n5214)) + ((!n_n5239) & (n_n5238) & (!n_n5166) & (n_n5163) & (n_n5214)) + ((!n_n5239) & (n_n5238) & (n_n5166) & (!n_n5163) & (!n_n5214)) + ((!n_n5239) & (n_n5238) & (n_n5166) & (!n_n5163) & (n_n5214)) + ((!n_n5239) & (n_n5238) & (n_n5166) & (n_n5163) & (!n_n5214)) + ((!n_n5239) & (n_n5238) & (n_n5166) & (n_n5163) & (n_n5214)) + ((n_n5239) & (!n_n5238) & (!n_n5166) & (!n_n5163) & (!n_n5214)) + ((n_n5239) & (!n_n5238) & (!n_n5166) & (!n_n5163) & (n_n5214)) + ((n_n5239) & (!n_n5238) & (!n_n5166) & (n_n5163) & (!n_n5214)) + ((n_n5239) & (!n_n5238) & (!n_n5166) & (n_n5163) & (n_n5214)) + ((n_n5239) & (!n_n5238) & (n_n5166) & (!n_n5163) & (!n_n5214)) + ((n_n5239) & (!n_n5238) & (n_n5166) & (!n_n5163) & (n_n5214)) + ((n_n5239) & (!n_n5238) & (n_n5166) & (n_n5163) & (!n_n5214)) + ((n_n5239) & (!n_n5238) & (n_n5166) & (n_n5163) & (n_n5214)) + ((n_n5239) & (n_n5238) & (!n_n5166) & (!n_n5163) & (!n_n5214)) + ((n_n5239) & (n_n5238) & (!n_n5166) & (!n_n5163) & (n_n5214)) + ((n_n5239) & (n_n5238) & (!n_n5166) & (n_n5163) & (!n_n5214)) + ((n_n5239) & (n_n5238) & (!n_n5166) & (n_n5163) & (n_n5214)) + ((n_n5239) & (n_n5238) & (n_n5166) & (!n_n5163) & (!n_n5214)) + ((n_n5239) & (n_n5238) & (n_n5166) & (!n_n5163) & (n_n5214)) + ((n_n5239) & (n_n5238) & (n_n5166) & (n_n5163) & (!n_n5214)) + ((n_n5239) & (n_n5238) & (n_n5166) & (n_n5163) & (n_n5214)));
	assign x13710x = (((!n_n5274) & (!n_n5300) & (!n_n5254) & (n_n5287)) + ((!n_n5274) & (!n_n5300) & (n_n5254) & (!n_n5287)) + ((!n_n5274) & (!n_n5300) & (n_n5254) & (n_n5287)) + ((!n_n5274) & (n_n5300) & (!n_n5254) & (!n_n5287)) + ((!n_n5274) & (n_n5300) & (!n_n5254) & (n_n5287)) + ((!n_n5274) & (n_n5300) & (n_n5254) & (!n_n5287)) + ((!n_n5274) & (n_n5300) & (n_n5254) & (n_n5287)) + ((n_n5274) & (!n_n5300) & (!n_n5254) & (!n_n5287)) + ((n_n5274) & (!n_n5300) & (!n_n5254) & (n_n5287)) + ((n_n5274) & (!n_n5300) & (n_n5254) & (!n_n5287)) + ((n_n5274) & (!n_n5300) & (n_n5254) & (n_n5287)) + ((n_n5274) & (n_n5300) & (!n_n5254) & (!n_n5287)) + ((n_n5274) & (n_n5300) & (!n_n5254) & (n_n5287)) + ((n_n5274) & (n_n5300) & (n_n5254) & (!n_n5287)) + ((n_n5274) & (n_n5300) & (n_n5254) & (n_n5287)));
	assign x13711x = (((!n_n5293) & (!n_n5240) & (!n_n5281) & (!n_n5268) & (n_n5261)) + ((!n_n5293) & (!n_n5240) & (!n_n5281) & (n_n5268) & (!n_n5261)) + ((!n_n5293) & (!n_n5240) & (!n_n5281) & (n_n5268) & (n_n5261)) + ((!n_n5293) & (!n_n5240) & (n_n5281) & (!n_n5268) & (!n_n5261)) + ((!n_n5293) & (!n_n5240) & (n_n5281) & (!n_n5268) & (n_n5261)) + ((!n_n5293) & (!n_n5240) & (n_n5281) & (n_n5268) & (!n_n5261)) + ((!n_n5293) & (!n_n5240) & (n_n5281) & (n_n5268) & (n_n5261)) + ((!n_n5293) & (n_n5240) & (!n_n5281) & (!n_n5268) & (!n_n5261)) + ((!n_n5293) & (n_n5240) & (!n_n5281) & (!n_n5268) & (n_n5261)) + ((!n_n5293) & (n_n5240) & (!n_n5281) & (n_n5268) & (!n_n5261)) + ((!n_n5293) & (n_n5240) & (!n_n5281) & (n_n5268) & (n_n5261)) + ((!n_n5293) & (n_n5240) & (n_n5281) & (!n_n5268) & (!n_n5261)) + ((!n_n5293) & (n_n5240) & (n_n5281) & (!n_n5268) & (n_n5261)) + ((!n_n5293) & (n_n5240) & (n_n5281) & (n_n5268) & (!n_n5261)) + ((!n_n5293) & (n_n5240) & (n_n5281) & (n_n5268) & (n_n5261)) + ((n_n5293) & (!n_n5240) & (!n_n5281) & (!n_n5268) & (!n_n5261)) + ((n_n5293) & (!n_n5240) & (!n_n5281) & (!n_n5268) & (n_n5261)) + ((n_n5293) & (!n_n5240) & (!n_n5281) & (n_n5268) & (!n_n5261)) + ((n_n5293) & (!n_n5240) & (!n_n5281) & (n_n5268) & (n_n5261)) + ((n_n5293) & (!n_n5240) & (n_n5281) & (!n_n5268) & (!n_n5261)) + ((n_n5293) & (!n_n5240) & (n_n5281) & (!n_n5268) & (n_n5261)) + ((n_n5293) & (!n_n5240) & (n_n5281) & (n_n5268) & (!n_n5261)) + ((n_n5293) & (!n_n5240) & (n_n5281) & (n_n5268) & (n_n5261)) + ((n_n5293) & (n_n5240) & (!n_n5281) & (!n_n5268) & (!n_n5261)) + ((n_n5293) & (n_n5240) & (!n_n5281) & (!n_n5268) & (n_n5261)) + ((n_n5293) & (n_n5240) & (!n_n5281) & (n_n5268) & (!n_n5261)) + ((n_n5293) & (n_n5240) & (!n_n5281) & (n_n5268) & (n_n5261)) + ((n_n5293) & (n_n5240) & (n_n5281) & (!n_n5268) & (!n_n5261)) + ((n_n5293) & (n_n5240) & (n_n5281) & (!n_n5268) & (n_n5261)) + ((n_n5293) & (n_n5240) & (n_n5281) & (n_n5268) & (!n_n5261)) + ((n_n5293) & (n_n5240) & (n_n5281) & (n_n5268) & (n_n5261)));
	assign x13713x = (((!n_n5305) & (!n_n482) & (!x23x) & (!n_n65) & (n_n5302)) + ((!n_n5305) & (!n_n482) & (!x23x) & (n_n65) & (n_n5302)) + ((!n_n5305) & (!n_n482) & (x23x) & (!n_n65) & (n_n5302)) + ((!n_n5305) & (!n_n482) & (x23x) & (n_n65) & (n_n5302)) + ((!n_n5305) & (n_n482) & (!x23x) & (!n_n65) & (n_n5302)) + ((!n_n5305) & (n_n482) & (!x23x) & (n_n65) & (n_n5302)) + ((!n_n5305) & (n_n482) & (x23x) & (!n_n65) & (n_n5302)) + ((!n_n5305) & (n_n482) & (x23x) & (n_n65) & (!n_n5302)) + ((!n_n5305) & (n_n482) & (x23x) & (n_n65) & (n_n5302)) + ((n_n5305) & (!n_n482) & (!x23x) & (!n_n65) & (!n_n5302)) + ((n_n5305) & (!n_n482) & (!x23x) & (!n_n65) & (n_n5302)) + ((n_n5305) & (!n_n482) & (!x23x) & (n_n65) & (!n_n5302)) + ((n_n5305) & (!n_n482) & (!x23x) & (n_n65) & (n_n5302)) + ((n_n5305) & (!n_n482) & (x23x) & (!n_n65) & (!n_n5302)) + ((n_n5305) & (!n_n482) & (x23x) & (!n_n65) & (n_n5302)) + ((n_n5305) & (!n_n482) & (x23x) & (n_n65) & (!n_n5302)) + ((n_n5305) & (!n_n482) & (x23x) & (n_n65) & (n_n5302)) + ((n_n5305) & (n_n482) & (!x23x) & (!n_n65) & (!n_n5302)) + ((n_n5305) & (n_n482) & (!x23x) & (!n_n65) & (n_n5302)) + ((n_n5305) & (n_n482) & (!x23x) & (n_n65) & (!n_n5302)) + ((n_n5305) & (n_n482) & (!x23x) & (n_n65) & (n_n5302)) + ((n_n5305) & (n_n482) & (x23x) & (!n_n65) & (!n_n5302)) + ((n_n5305) & (n_n482) & (x23x) & (!n_n65) & (n_n5302)) + ((n_n5305) & (n_n482) & (x23x) & (n_n65) & (!n_n5302)) + ((n_n5305) & (n_n482) & (x23x) & (n_n65) & (n_n5302)));
	assign n_n3189 = (((!x13703x) & (!x13704x) & (!x13710x) & (!x13711x) & (x13713x)) + ((!x13703x) & (!x13704x) & (!x13710x) & (x13711x) & (!x13713x)) + ((!x13703x) & (!x13704x) & (!x13710x) & (x13711x) & (x13713x)) + ((!x13703x) & (!x13704x) & (x13710x) & (!x13711x) & (!x13713x)) + ((!x13703x) & (!x13704x) & (x13710x) & (!x13711x) & (x13713x)) + ((!x13703x) & (!x13704x) & (x13710x) & (x13711x) & (!x13713x)) + ((!x13703x) & (!x13704x) & (x13710x) & (x13711x) & (x13713x)) + ((!x13703x) & (x13704x) & (!x13710x) & (!x13711x) & (!x13713x)) + ((!x13703x) & (x13704x) & (!x13710x) & (!x13711x) & (x13713x)) + ((!x13703x) & (x13704x) & (!x13710x) & (x13711x) & (!x13713x)) + ((!x13703x) & (x13704x) & (!x13710x) & (x13711x) & (x13713x)) + ((!x13703x) & (x13704x) & (x13710x) & (!x13711x) & (!x13713x)) + ((!x13703x) & (x13704x) & (x13710x) & (!x13711x) & (x13713x)) + ((!x13703x) & (x13704x) & (x13710x) & (x13711x) & (!x13713x)) + ((!x13703x) & (x13704x) & (x13710x) & (x13711x) & (x13713x)) + ((x13703x) & (!x13704x) & (!x13710x) & (!x13711x) & (!x13713x)) + ((x13703x) & (!x13704x) & (!x13710x) & (!x13711x) & (x13713x)) + ((x13703x) & (!x13704x) & (!x13710x) & (x13711x) & (!x13713x)) + ((x13703x) & (!x13704x) & (!x13710x) & (x13711x) & (x13713x)) + ((x13703x) & (!x13704x) & (x13710x) & (!x13711x) & (!x13713x)) + ((x13703x) & (!x13704x) & (x13710x) & (!x13711x) & (x13713x)) + ((x13703x) & (!x13704x) & (x13710x) & (x13711x) & (!x13713x)) + ((x13703x) & (!x13704x) & (x13710x) & (x13711x) & (x13713x)) + ((x13703x) & (x13704x) & (!x13710x) & (!x13711x) & (!x13713x)) + ((x13703x) & (x13704x) & (!x13710x) & (!x13711x) & (x13713x)) + ((x13703x) & (x13704x) & (!x13710x) & (x13711x) & (!x13713x)) + ((x13703x) & (x13704x) & (!x13710x) & (x13711x) & (x13713x)) + ((x13703x) & (x13704x) & (x13710x) & (!x13711x) & (!x13713x)) + ((x13703x) & (x13704x) & (x13710x) & (!x13711x) & (x13713x)) + ((x13703x) & (x13704x) & (x13710x) & (x13711x) & (!x13713x)) + ((x13703x) & (x13704x) & (x13710x) & (x13711x) & (x13713x)));
	assign n_n4487 = (((i_1_) & (!i_2_) & (i_0_) & (n_n509) & (x23x)));
	assign n_n4409 = (((!i_9_) & (n_n536) & (n_n473) & (n_n534)));
	assign x13735x = (((!x20x) & (!x496x) & (!n_n4472) & (!n_n4487) & (n_n4409)) + ((!x20x) & (!x496x) & (!n_n4472) & (n_n4487) & (!n_n4409)) + ((!x20x) & (!x496x) & (!n_n4472) & (n_n4487) & (n_n4409)) + ((!x20x) & (!x496x) & (n_n4472) & (!n_n4487) & (!n_n4409)) + ((!x20x) & (!x496x) & (n_n4472) & (!n_n4487) & (n_n4409)) + ((!x20x) & (!x496x) & (n_n4472) & (n_n4487) & (!n_n4409)) + ((!x20x) & (!x496x) & (n_n4472) & (n_n4487) & (n_n4409)) + ((!x20x) & (x496x) & (!n_n4472) & (!n_n4487) & (n_n4409)) + ((!x20x) & (x496x) & (!n_n4472) & (n_n4487) & (!n_n4409)) + ((!x20x) & (x496x) & (!n_n4472) & (n_n4487) & (n_n4409)) + ((!x20x) & (x496x) & (n_n4472) & (!n_n4487) & (!n_n4409)) + ((!x20x) & (x496x) & (n_n4472) & (!n_n4487) & (n_n4409)) + ((!x20x) & (x496x) & (n_n4472) & (n_n4487) & (!n_n4409)) + ((!x20x) & (x496x) & (n_n4472) & (n_n4487) & (n_n4409)) + ((x20x) & (!x496x) & (!n_n4472) & (!n_n4487) & (n_n4409)) + ((x20x) & (!x496x) & (!n_n4472) & (n_n4487) & (!n_n4409)) + ((x20x) & (!x496x) & (!n_n4472) & (n_n4487) & (n_n4409)) + ((x20x) & (!x496x) & (n_n4472) & (!n_n4487) & (!n_n4409)) + ((x20x) & (!x496x) & (n_n4472) & (!n_n4487) & (n_n4409)) + ((x20x) & (!x496x) & (n_n4472) & (n_n4487) & (!n_n4409)) + ((x20x) & (!x496x) & (n_n4472) & (n_n4487) & (n_n4409)) + ((x20x) & (x496x) & (!n_n4472) & (!n_n4487) & (!n_n4409)) + ((x20x) & (x496x) & (!n_n4472) & (!n_n4487) & (n_n4409)) + ((x20x) & (x496x) & (!n_n4472) & (n_n4487) & (!n_n4409)) + ((x20x) & (x496x) & (!n_n4472) & (n_n4487) & (n_n4409)) + ((x20x) & (x496x) & (n_n4472) & (!n_n4487) & (!n_n4409)) + ((x20x) & (x496x) & (n_n4472) & (!n_n4487) & (n_n4409)) + ((x20x) & (x496x) & (n_n4472) & (n_n4487) & (!n_n4409)) + ((x20x) & (x496x) & (n_n4472) & (n_n4487) & (n_n4409)));
	assign n_n4456 = (((i_9_) & (n_n518) & (n_n455) & (n_n534)));
	assign n_n4484 = (((i_9_) & (n_n455) & (n_n509) & (n_n522)));
	assign n_n4462 = (((i_9_) & (n_n518) & (n_n455) & (n_n528)));
	assign n_n4428 = (((i_9_) & (n_n536) & (n_n530) & (n_n464)));
	assign x13736x = (((!n_n4456) & (!n_n4458) & (!n_n4484) & (!n_n4462) & (n_n4428)) + ((!n_n4456) & (!n_n4458) & (!n_n4484) & (n_n4462) & (!n_n4428)) + ((!n_n4456) & (!n_n4458) & (!n_n4484) & (n_n4462) & (n_n4428)) + ((!n_n4456) & (!n_n4458) & (n_n4484) & (!n_n4462) & (!n_n4428)) + ((!n_n4456) & (!n_n4458) & (n_n4484) & (!n_n4462) & (n_n4428)) + ((!n_n4456) & (!n_n4458) & (n_n4484) & (n_n4462) & (!n_n4428)) + ((!n_n4456) & (!n_n4458) & (n_n4484) & (n_n4462) & (n_n4428)) + ((!n_n4456) & (n_n4458) & (!n_n4484) & (!n_n4462) & (!n_n4428)) + ((!n_n4456) & (n_n4458) & (!n_n4484) & (!n_n4462) & (n_n4428)) + ((!n_n4456) & (n_n4458) & (!n_n4484) & (n_n4462) & (!n_n4428)) + ((!n_n4456) & (n_n4458) & (!n_n4484) & (n_n4462) & (n_n4428)) + ((!n_n4456) & (n_n4458) & (n_n4484) & (!n_n4462) & (!n_n4428)) + ((!n_n4456) & (n_n4458) & (n_n4484) & (!n_n4462) & (n_n4428)) + ((!n_n4456) & (n_n4458) & (n_n4484) & (n_n4462) & (!n_n4428)) + ((!n_n4456) & (n_n4458) & (n_n4484) & (n_n4462) & (n_n4428)) + ((n_n4456) & (!n_n4458) & (!n_n4484) & (!n_n4462) & (!n_n4428)) + ((n_n4456) & (!n_n4458) & (!n_n4484) & (!n_n4462) & (n_n4428)) + ((n_n4456) & (!n_n4458) & (!n_n4484) & (n_n4462) & (!n_n4428)) + ((n_n4456) & (!n_n4458) & (!n_n4484) & (n_n4462) & (n_n4428)) + ((n_n4456) & (!n_n4458) & (n_n4484) & (!n_n4462) & (!n_n4428)) + ((n_n4456) & (!n_n4458) & (n_n4484) & (!n_n4462) & (n_n4428)) + ((n_n4456) & (!n_n4458) & (n_n4484) & (n_n4462) & (!n_n4428)) + ((n_n4456) & (!n_n4458) & (n_n4484) & (n_n4462) & (n_n4428)) + ((n_n4456) & (n_n4458) & (!n_n4484) & (!n_n4462) & (!n_n4428)) + ((n_n4456) & (n_n4458) & (!n_n4484) & (!n_n4462) & (n_n4428)) + ((n_n4456) & (n_n4458) & (!n_n4484) & (n_n4462) & (!n_n4428)) + ((n_n4456) & (n_n4458) & (!n_n4484) & (n_n4462) & (n_n4428)) + ((n_n4456) & (n_n4458) & (n_n4484) & (!n_n4462) & (!n_n4428)) + ((n_n4456) & (n_n4458) & (n_n4484) & (!n_n4462) & (n_n4428)) + ((n_n4456) & (n_n4458) & (n_n4484) & (n_n4462) & (!n_n4428)) + ((n_n4456) & (n_n4458) & (n_n4484) & (n_n4462) & (n_n4428)));
	assign n_n4539 = (((!i_9_) & (n_n455) & (n_n473) & (n_n532)));
	assign n_n4544 = (((i_9_) & (n_n526) & (n_n455) & (n_n473)));
	assign n_n4533 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n455) & (x20x)));
	assign n_n4507 = (((!i_9_) & (n_n455) & (n_n532) & (n_n491)));
	assign x13741x = (((!n_n4539) & (!n_n4544) & (!n_n4533) & (n_n4507)) + ((!n_n4539) & (!n_n4544) & (n_n4533) & (!n_n4507)) + ((!n_n4539) & (!n_n4544) & (n_n4533) & (n_n4507)) + ((!n_n4539) & (n_n4544) & (!n_n4533) & (!n_n4507)) + ((!n_n4539) & (n_n4544) & (!n_n4533) & (n_n4507)) + ((!n_n4539) & (n_n4544) & (n_n4533) & (!n_n4507)) + ((!n_n4539) & (n_n4544) & (n_n4533) & (n_n4507)) + ((n_n4539) & (!n_n4544) & (!n_n4533) & (!n_n4507)) + ((n_n4539) & (!n_n4544) & (!n_n4533) & (n_n4507)) + ((n_n4539) & (!n_n4544) & (n_n4533) & (!n_n4507)) + ((n_n4539) & (!n_n4544) & (n_n4533) & (n_n4507)) + ((n_n4539) & (n_n4544) & (!n_n4533) & (!n_n4507)) + ((n_n4539) & (n_n4544) & (!n_n4533) & (n_n4507)) + ((n_n4539) & (n_n4544) & (n_n4533) & (!n_n4507)) + ((n_n4539) & (n_n4544) & (n_n4533) & (n_n4507)));
	assign n_n4499 = (((!i_9_) & (n_n524) & (n_n455) & (n_n500)));
	assign n_n4532 = (((i_9_) & (n_n482) & (n_n455) & (n_n522)));
	assign n_n4545 = (((!i_9_) & (n_n526) & (n_n455) & (n_n473)));
	assign x471x = (((!i_9_) & (n_n455) & (!n_n522) & (x20x) & (n_n464)) + ((!i_9_) & (n_n455) & (n_n522) & (x20x) & (n_n464)) + ((i_9_) & (n_n455) & (!n_n522) & (x20x) & (n_n464)) + ((i_9_) & (n_n455) & (n_n522) & (!x20x) & (n_n464)) + ((i_9_) & (n_n455) & (n_n522) & (x20x) & (n_n464)));
	assign n_n3205 = (((!x13741x) & (!n_n4499) & (!n_n4532) & (!n_n4545) & (x471x)) + ((!x13741x) & (!n_n4499) & (!n_n4532) & (n_n4545) & (!x471x)) + ((!x13741x) & (!n_n4499) & (!n_n4532) & (n_n4545) & (x471x)) + ((!x13741x) & (!n_n4499) & (n_n4532) & (!n_n4545) & (!x471x)) + ((!x13741x) & (!n_n4499) & (n_n4532) & (!n_n4545) & (x471x)) + ((!x13741x) & (!n_n4499) & (n_n4532) & (n_n4545) & (!x471x)) + ((!x13741x) & (!n_n4499) & (n_n4532) & (n_n4545) & (x471x)) + ((!x13741x) & (n_n4499) & (!n_n4532) & (!n_n4545) & (!x471x)) + ((!x13741x) & (n_n4499) & (!n_n4532) & (!n_n4545) & (x471x)) + ((!x13741x) & (n_n4499) & (!n_n4532) & (n_n4545) & (!x471x)) + ((!x13741x) & (n_n4499) & (!n_n4532) & (n_n4545) & (x471x)) + ((!x13741x) & (n_n4499) & (n_n4532) & (!n_n4545) & (!x471x)) + ((!x13741x) & (n_n4499) & (n_n4532) & (!n_n4545) & (x471x)) + ((!x13741x) & (n_n4499) & (n_n4532) & (n_n4545) & (!x471x)) + ((!x13741x) & (n_n4499) & (n_n4532) & (n_n4545) & (x471x)) + ((x13741x) & (!n_n4499) & (!n_n4532) & (!n_n4545) & (!x471x)) + ((x13741x) & (!n_n4499) & (!n_n4532) & (!n_n4545) & (x471x)) + ((x13741x) & (!n_n4499) & (!n_n4532) & (n_n4545) & (!x471x)) + ((x13741x) & (!n_n4499) & (!n_n4532) & (n_n4545) & (x471x)) + ((x13741x) & (!n_n4499) & (n_n4532) & (!n_n4545) & (!x471x)) + ((x13741x) & (!n_n4499) & (n_n4532) & (!n_n4545) & (x471x)) + ((x13741x) & (!n_n4499) & (n_n4532) & (n_n4545) & (!x471x)) + ((x13741x) & (!n_n4499) & (n_n4532) & (n_n4545) & (x471x)) + ((x13741x) & (n_n4499) & (!n_n4532) & (!n_n4545) & (!x471x)) + ((x13741x) & (n_n4499) & (!n_n4532) & (!n_n4545) & (x471x)) + ((x13741x) & (n_n4499) & (!n_n4532) & (n_n4545) & (!x471x)) + ((x13741x) & (n_n4499) & (!n_n4532) & (n_n4545) & (x471x)) + ((x13741x) & (n_n4499) & (n_n4532) & (!n_n4545) & (!x471x)) + ((x13741x) & (n_n4499) & (n_n4532) & (!n_n4545) & (x471x)) + ((x13741x) & (n_n4499) & (n_n4532) & (n_n4545) & (!x471x)) + ((x13741x) & (n_n4499) & (n_n4532) & (n_n4545) & (x471x)));
	assign n_n4638 = (((i_9_) & (n_n528) & (n_n390) & (n_n491)));
	assign n_n4640 = (((i_9_) & (n_n526) & (n_n390) & (n_n491)));
	assign n_n4662 = (((i_9_) & (n_n482) & (n_n390) & (n_n520)));
	assign n_n4683 = (((!i_9_) & (n_n390) & (n_n532) & (n_n464)));
	assign x13760x = (((!n_n482) & (!n_n390) & (!x23x) & (!n_n4685) & (n_n3125)) + ((!n_n482) & (!n_n390) & (!x23x) & (n_n4685) & (!n_n3125)) + ((!n_n482) & (!n_n390) & (!x23x) & (n_n4685) & (n_n3125)) + ((!n_n482) & (!n_n390) & (x23x) & (!n_n4685) & (n_n3125)) + ((!n_n482) & (!n_n390) & (x23x) & (n_n4685) & (!n_n3125)) + ((!n_n482) & (!n_n390) & (x23x) & (n_n4685) & (n_n3125)) + ((!n_n482) & (n_n390) & (!x23x) & (!n_n4685) & (n_n3125)) + ((!n_n482) & (n_n390) & (!x23x) & (n_n4685) & (!n_n3125)) + ((!n_n482) & (n_n390) & (!x23x) & (n_n4685) & (n_n3125)) + ((!n_n482) & (n_n390) & (x23x) & (!n_n4685) & (n_n3125)) + ((!n_n482) & (n_n390) & (x23x) & (n_n4685) & (!n_n3125)) + ((!n_n482) & (n_n390) & (x23x) & (n_n4685) & (n_n3125)) + ((n_n482) & (!n_n390) & (!x23x) & (!n_n4685) & (n_n3125)) + ((n_n482) & (!n_n390) & (!x23x) & (n_n4685) & (!n_n3125)) + ((n_n482) & (!n_n390) & (!x23x) & (n_n4685) & (n_n3125)) + ((n_n482) & (!n_n390) & (x23x) & (!n_n4685) & (n_n3125)) + ((n_n482) & (!n_n390) & (x23x) & (n_n4685) & (!n_n3125)) + ((n_n482) & (!n_n390) & (x23x) & (n_n4685) & (n_n3125)) + ((n_n482) & (n_n390) & (!x23x) & (!n_n4685) & (n_n3125)) + ((n_n482) & (n_n390) & (!x23x) & (n_n4685) & (!n_n3125)) + ((n_n482) & (n_n390) & (!x23x) & (n_n4685) & (n_n3125)) + ((n_n482) & (n_n390) & (x23x) & (!n_n4685) & (!n_n3125)) + ((n_n482) & (n_n390) & (x23x) & (!n_n4685) & (n_n3125)) + ((n_n482) & (n_n390) & (x23x) & (n_n4685) & (!n_n3125)) + ((n_n482) & (n_n390) & (x23x) & (n_n4685) & (n_n3125)));
	assign x13761x = (((!n_n4638) & (!n_n4640) & (!n_n4662) & (!n_n4683) & (x13760x)) + ((!n_n4638) & (!n_n4640) & (!n_n4662) & (n_n4683) & (!x13760x)) + ((!n_n4638) & (!n_n4640) & (!n_n4662) & (n_n4683) & (x13760x)) + ((!n_n4638) & (!n_n4640) & (n_n4662) & (!n_n4683) & (!x13760x)) + ((!n_n4638) & (!n_n4640) & (n_n4662) & (!n_n4683) & (x13760x)) + ((!n_n4638) & (!n_n4640) & (n_n4662) & (n_n4683) & (!x13760x)) + ((!n_n4638) & (!n_n4640) & (n_n4662) & (n_n4683) & (x13760x)) + ((!n_n4638) & (n_n4640) & (!n_n4662) & (!n_n4683) & (!x13760x)) + ((!n_n4638) & (n_n4640) & (!n_n4662) & (!n_n4683) & (x13760x)) + ((!n_n4638) & (n_n4640) & (!n_n4662) & (n_n4683) & (!x13760x)) + ((!n_n4638) & (n_n4640) & (!n_n4662) & (n_n4683) & (x13760x)) + ((!n_n4638) & (n_n4640) & (n_n4662) & (!n_n4683) & (!x13760x)) + ((!n_n4638) & (n_n4640) & (n_n4662) & (!n_n4683) & (x13760x)) + ((!n_n4638) & (n_n4640) & (n_n4662) & (n_n4683) & (!x13760x)) + ((!n_n4638) & (n_n4640) & (n_n4662) & (n_n4683) & (x13760x)) + ((n_n4638) & (!n_n4640) & (!n_n4662) & (!n_n4683) & (!x13760x)) + ((n_n4638) & (!n_n4640) & (!n_n4662) & (!n_n4683) & (x13760x)) + ((n_n4638) & (!n_n4640) & (!n_n4662) & (n_n4683) & (!x13760x)) + ((n_n4638) & (!n_n4640) & (!n_n4662) & (n_n4683) & (x13760x)) + ((n_n4638) & (!n_n4640) & (n_n4662) & (!n_n4683) & (!x13760x)) + ((n_n4638) & (!n_n4640) & (n_n4662) & (!n_n4683) & (x13760x)) + ((n_n4638) & (!n_n4640) & (n_n4662) & (n_n4683) & (!x13760x)) + ((n_n4638) & (!n_n4640) & (n_n4662) & (n_n4683) & (x13760x)) + ((n_n4638) & (n_n4640) & (!n_n4662) & (!n_n4683) & (!x13760x)) + ((n_n4638) & (n_n4640) & (!n_n4662) & (!n_n4683) & (x13760x)) + ((n_n4638) & (n_n4640) & (!n_n4662) & (n_n4683) & (!x13760x)) + ((n_n4638) & (n_n4640) & (!n_n4662) & (n_n4683) & (x13760x)) + ((n_n4638) & (n_n4640) & (n_n4662) & (!n_n4683) & (!x13760x)) + ((n_n4638) & (n_n4640) & (n_n4662) & (!n_n4683) & (x13760x)) + ((n_n4638) & (n_n4640) & (n_n4662) & (n_n4683) & (!x13760x)) + ((n_n4638) & (n_n4640) & (n_n4662) & (n_n4683) & (x13760x)));
	assign x13747x = (((!n_n4779) & (!n_n4786) & (!n_n4755) & (n_n4781)) + ((!n_n4779) & (!n_n4786) & (n_n4755) & (!n_n4781)) + ((!n_n4779) & (!n_n4786) & (n_n4755) & (n_n4781)) + ((!n_n4779) & (n_n4786) & (!n_n4755) & (!n_n4781)) + ((!n_n4779) & (n_n4786) & (!n_n4755) & (n_n4781)) + ((!n_n4779) & (n_n4786) & (n_n4755) & (!n_n4781)) + ((!n_n4779) & (n_n4786) & (n_n4755) & (n_n4781)) + ((n_n4779) & (!n_n4786) & (!n_n4755) & (!n_n4781)) + ((n_n4779) & (!n_n4786) & (!n_n4755) & (n_n4781)) + ((n_n4779) & (!n_n4786) & (n_n4755) & (!n_n4781)) + ((n_n4779) & (!n_n4786) & (n_n4755) & (n_n4781)) + ((n_n4779) & (n_n4786) & (!n_n4755) & (!n_n4781)) + ((n_n4779) & (n_n4786) & (!n_n4755) & (n_n4781)) + ((n_n4779) & (n_n4786) & (n_n4755) & (!n_n4781)) + ((n_n4779) & (n_n4786) & (n_n4755) & (n_n4781)));
	assign x13748x = (((!n_n4724) & (!n_n4767) & (!n_n4752) & (!n_n4799) & (n_n4723)) + ((!n_n4724) & (!n_n4767) & (!n_n4752) & (n_n4799) & (!n_n4723)) + ((!n_n4724) & (!n_n4767) & (!n_n4752) & (n_n4799) & (n_n4723)) + ((!n_n4724) & (!n_n4767) & (n_n4752) & (!n_n4799) & (!n_n4723)) + ((!n_n4724) & (!n_n4767) & (n_n4752) & (!n_n4799) & (n_n4723)) + ((!n_n4724) & (!n_n4767) & (n_n4752) & (n_n4799) & (!n_n4723)) + ((!n_n4724) & (!n_n4767) & (n_n4752) & (n_n4799) & (n_n4723)) + ((!n_n4724) & (n_n4767) & (!n_n4752) & (!n_n4799) & (!n_n4723)) + ((!n_n4724) & (n_n4767) & (!n_n4752) & (!n_n4799) & (n_n4723)) + ((!n_n4724) & (n_n4767) & (!n_n4752) & (n_n4799) & (!n_n4723)) + ((!n_n4724) & (n_n4767) & (!n_n4752) & (n_n4799) & (n_n4723)) + ((!n_n4724) & (n_n4767) & (n_n4752) & (!n_n4799) & (!n_n4723)) + ((!n_n4724) & (n_n4767) & (n_n4752) & (!n_n4799) & (n_n4723)) + ((!n_n4724) & (n_n4767) & (n_n4752) & (n_n4799) & (!n_n4723)) + ((!n_n4724) & (n_n4767) & (n_n4752) & (n_n4799) & (n_n4723)) + ((n_n4724) & (!n_n4767) & (!n_n4752) & (!n_n4799) & (!n_n4723)) + ((n_n4724) & (!n_n4767) & (!n_n4752) & (!n_n4799) & (n_n4723)) + ((n_n4724) & (!n_n4767) & (!n_n4752) & (n_n4799) & (!n_n4723)) + ((n_n4724) & (!n_n4767) & (!n_n4752) & (n_n4799) & (n_n4723)) + ((n_n4724) & (!n_n4767) & (n_n4752) & (!n_n4799) & (!n_n4723)) + ((n_n4724) & (!n_n4767) & (n_n4752) & (!n_n4799) & (n_n4723)) + ((n_n4724) & (!n_n4767) & (n_n4752) & (n_n4799) & (!n_n4723)) + ((n_n4724) & (!n_n4767) & (n_n4752) & (n_n4799) & (n_n4723)) + ((n_n4724) & (n_n4767) & (!n_n4752) & (!n_n4799) & (!n_n4723)) + ((n_n4724) & (n_n4767) & (!n_n4752) & (!n_n4799) & (n_n4723)) + ((n_n4724) & (n_n4767) & (!n_n4752) & (n_n4799) & (!n_n4723)) + ((n_n4724) & (n_n4767) & (!n_n4752) & (n_n4799) & (n_n4723)) + ((n_n4724) & (n_n4767) & (n_n4752) & (!n_n4799) & (!n_n4723)) + ((n_n4724) & (n_n4767) & (n_n4752) & (!n_n4799) & (n_n4723)) + ((n_n4724) & (n_n4767) & (n_n4752) & (n_n4799) & (!n_n4723)) + ((n_n4724) & (n_n4767) & (n_n4752) & (n_n4799) & (n_n4723)));
	assign x13753x = (((!n_n4571) & (!n_n4578) & (!n_n4570) & (n_n4594)) + ((!n_n4571) & (!n_n4578) & (n_n4570) & (!n_n4594)) + ((!n_n4571) & (!n_n4578) & (n_n4570) & (n_n4594)) + ((!n_n4571) & (n_n4578) & (!n_n4570) & (!n_n4594)) + ((!n_n4571) & (n_n4578) & (!n_n4570) & (n_n4594)) + ((!n_n4571) & (n_n4578) & (n_n4570) & (!n_n4594)) + ((!n_n4571) & (n_n4578) & (n_n4570) & (n_n4594)) + ((n_n4571) & (!n_n4578) & (!n_n4570) & (!n_n4594)) + ((n_n4571) & (!n_n4578) & (!n_n4570) & (n_n4594)) + ((n_n4571) & (!n_n4578) & (n_n4570) & (!n_n4594)) + ((n_n4571) & (!n_n4578) & (n_n4570) & (n_n4594)) + ((n_n4571) & (n_n4578) & (!n_n4570) & (!n_n4594)) + ((n_n4571) & (n_n4578) & (!n_n4570) & (n_n4594)) + ((n_n4571) & (n_n4578) & (n_n4570) & (!n_n4594)) + ((n_n4571) & (n_n4578) & (n_n4570) & (n_n4594)));
	assign x13754x = (((!n_n4633) & (!n_n4629) & (!n_n4583) & (!n_n4635) & (n_n4630)) + ((!n_n4633) & (!n_n4629) & (!n_n4583) & (n_n4635) & (!n_n4630)) + ((!n_n4633) & (!n_n4629) & (!n_n4583) & (n_n4635) & (n_n4630)) + ((!n_n4633) & (!n_n4629) & (n_n4583) & (!n_n4635) & (!n_n4630)) + ((!n_n4633) & (!n_n4629) & (n_n4583) & (!n_n4635) & (n_n4630)) + ((!n_n4633) & (!n_n4629) & (n_n4583) & (n_n4635) & (!n_n4630)) + ((!n_n4633) & (!n_n4629) & (n_n4583) & (n_n4635) & (n_n4630)) + ((!n_n4633) & (n_n4629) & (!n_n4583) & (!n_n4635) & (!n_n4630)) + ((!n_n4633) & (n_n4629) & (!n_n4583) & (!n_n4635) & (n_n4630)) + ((!n_n4633) & (n_n4629) & (!n_n4583) & (n_n4635) & (!n_n4630)) + ((!n_n4633) & (n_n4629) & (!n_n4583) & (n_n4635) & (n_n4630)) + ((!n_n4633) & (n_n4629) & (n_n4583) & (!n_n4635) & (!n_n4630)) + ((!n_n4633) & (n_n4629) & (n_n4583) & (!n_n4635) & (n_n4630)) + ((!n_n4633) & (n_n4629) & (n_n4583) & (n_n4635) & (!n_n4630)) + ((!n_n4633) & (n_n4629) & (n_n4583) & (n_n4635) & (n_n4630)) + ((n_n4633) & (!n_n4629) & (!n_n4583) & (!n_n4635) & (!n_n4630)) + ((n_n4633) & (!n_n4629) & (!n_n4583) & (!n_n4635) & (n_n4630)) + ((n_n4633) & (!n_n4629) & (!n_n4583) & (n_n4635) & (!n_n4630)) + ((n_n4633) & (!n_n4629) & (!n_n4583) & (n_n4635) & (n_n4630)) + ((n_n4633) & (!n_n4629) & (n_n4583) & (!n_n4635) & (!n_n4630)) + ((n_n4633) & (!n_n4629) & (n_n4583) & (!n_n4635) & (n_n4630)) + ((n_n4633) & (!n_n4629) & (n_n4583) & (n_n4635) & (!n_n4630)) + ((n_n4633) & (!n_n4629) & (n_n4583) & (n_n4635) & (n_n4630)) + ((n_n4633) & (n_n4629) & (!n_n4583) & (!n_n4635) & (!n_n4630)) + ((n_n4633) & (n_n4629) & (!n_n4583) & (!n_n4635) & (n_n4630)) + ((n_n4633) & (n_n4629) & (!n_n4583) & (n_n4635) & (!n_n4630)) + ((n_n4633) & (n_n4629) & (!n_n4583) & (n_n4635) & (n_n4630)) + ((n_n4633) & (n_n4629) & (n_n4583) & (!n_n4635) & (!n_n4630)) + ((n_n4633) & (n_n4629) & (n_n4583) & (!n_n4635) & (n_n4630)) + ((n_n4633) & (n_n4629) & (n_n4583) & (n_n4635) & (!n_n4630)) + ((n_n4633) & (n_n4629) & (n_n4583) & (n_n4635) & (n_n4630)));
	assign n_n4853 = (((!i_5_) & (i_3_) & (i_4_) & (n_n260) & (x20x)));
	assign n_n4847 = (((!i_9_) & (n_n518) & (n_n528) & (n_n260)));
	assign n_n4864 = (((i_9_) & (n_n526) & (n_n509) & (n_n260)));
	assign n_n4912 = (((i_9_) & (n_n526) & (n_n482) & (n_n260)));
	assign x13781x = (((!n_n4900) & (!n_n4849) & (!n_n4908) & (!n_n4891) & (n_n4896)) + ((!n_n4900) & (!n_n4849) & (!n_n4908) & (n_n4891) & (!n_n4896)) + ((!n_n4900) & (!n_n4849) & (!n_n4908) & (n_n4891) & (n_n4896)) + ((!n_n4900) & (!n_n4849) & (n_n4908) & (!n_n4891) & (!n_n4896)) + ((!n_n4900) & (!n_n4849) & (n_n4908) & (!n_n4891) & (n_n4896)) + ((!n_n4900) & (!n_n4849) & (n_n4908) & (n_n4891) & (!n_n4896)) + ((!n_n4900) & (!n_n4849) & (n_n4908) & (n_n4891) & (n_n4896)) + ((!n_n4900) & (n_n4849) & (!n_n4908) & (!n_n4891) & (!n_n4896)) + ((!n_n4900) & (n_n4849) & (!n_n4908) & (!n_n4891) & (n_n4896)) + ((!n_n4900) & (n_n4849) & (!n_n4908) & (n_n4891) & (!n_n4896)) + ((!n_n4900) & (n_n4849) & (!n_n4908) & (n_n4891) & (n_n4896)) + ((!n_n4900) & (n_n4849) & (n_n4908) & (!n_n4891) & (!n_n4896)) + ((!n_n4900) & (n_n4849) & (n_n4908) & (!n_n4891) & (n_n4896)) + ((!n_n4900) & (n_n4849) & (n_n4908) & (n_n4891) & (!n_n4896)) + ((!n_n4900) & (n_n4849) & (n_n4908) & (n_n4891) & (n_n4896)) + ((n_n4900) & (!n_n4849) & (!n_n4908) & (!n_n4891) & (!n_n4896)) + ((n_n4900) & (!n_n4849) & (!n_n4908) & (!n_n4891) & (n_n4896)) + ((n_n4900) & (!n_n4849) & (!n_n4908) & (n_n4891) & (!n_n4896)) + ((n_n4900) & (!n_n4849) & (!n_n4908) & (n_n4891) & (n_n4896)) + ((n_n4900) & (!n_n4849) & (n_n4908) & (!n_n4891) & (!n_n4896)) + ((n_n4900) & (!n_n4849) & (n_n4908) & (!n_n4891) & (n_n4896)) + ((n_n4900) & (!n_n4849) & (n_n4908) & (n_n4891) & (!n_n4896)) + ((n_n4900) & (!n_n4849) & (n_n4908) & (n_n4891) & (n_n4896)) + ((n_n4900) & (n_n4849) & (!n_n4908) & (!n_n4891) & (!n_n4896)) + ((n_n4900) & (n_n4849) & (!n_n4908) & (!n_n4891) & (n_n4896)) + ((n_n4900) & (n_n4849) & (!n_n4908) & (n_n4891) & (!n_n4896)) + ((n_n4900) & (n_n4849) & (!n_n4908) & (n_n4891) & (n_n4896)) + ((n_n4900) & (n_n4849) & (n_n4908) & (!n_n4891) & (!n_n4896)) + ((n_n4900) & (n_n4849) & (n_n4908) & (!n_n4891) & (n_n4896)) + ((n_n4900) & (n_n4849) & (n_n4908) & (n_n4891) & (!n_n4896)) + ((n_n4900) & (n_n4849) & (n_n4908) & (n_n4891) & (n_n4896)));
	assign x13767x = (((!n_n4977) & (!n_n4920) & (!n_n4922) & (n_n4959)) + ((!n_n4977) & (!n_n4920) & (n_n4922) & (!n_n4959)) + ((!n_n4977) & (!n_n4920) & (n_n4922) & (n_n4959)) + ((!n_n4977) & (n_n4920) & (!n_n4922) & (!n_n4959)) + ((!n_n4977) & (n_n4920) & (!n_n4922) & (n_n4959)) + ((!n_n4977) & (n_n4920) & (n_n4922) & (!n_n4959)) + ((!n_n4977) & (n_n4920) & (n_n4922) & (n_n4959)) + ((n_n4977) & (!n_n4920) & (!n_n4922) & (!n_n4959)) + ((n_n4977) & (!n_n4920) & (!n_n4922) & (n_n4959)) + ((n_n4977) & (!n_n4920) & (n_n4922) & (!n_n4959)) + ((n_n4977) & (!n_n4920) & (n_n4922) & (n_n4959)) + ((n_n4977) & (n_n4920) & (!n_n4922) & (!n_n4959)) + ((n_n4977) & (n_n4920) & (!n_n4922) & (n_n4959)) + ((n_n4977) & (n_n4920) & (n_n4922) & (!n_n4959)) + ((n_n4977) & (n_n4920) & (n_n4922) & (n_n4959)));
	assign x13768x = (((!n_n4980) & (!n_n4953) & (!x351x) & (n_n4972)) + ((!n_n4980) & (!n_n4953) & (x351x) & (!n_n4972)) + ((!n_n4980) & (!n_n4953) & (x351x) & (n_n4972)) + ((!n_n4980) & (n_n4953) & (!x351x) & (!n_n4972)) + ((!n_n4980) & (n_n4953) & (!x351x) & (n_n4972)) + ((!n_n4980) & (n_n4953) & (x351x) & (!n_n4972)) + ((!n_n4980) & (n_n4953) & (x351x) & (n_n4972)) + ((n_n4980) & (!n_n4953) & (!x351x) & (!n_n4972)) + ((n_n4980) & (!n_n4953) & (!x351x) & (n_n4972)) + ((n_n4980) & (!n_n4953) & (x351x) & (!n_n4972)) + ((n_n4980) & (!n_n4953) & (x351x) & (n_n4972)) + ((n_n4980) & (n_n4953) & (!x351x) & (!n_n4972)) + ((n_n4980) & (n_n4953) & (!x351x) & (n_n4972)) + ((n_n4980) & (n_n4953) & (x351x) & (!n_n4972)) + ((n_n4980) & (n_n4953) & (x351x) & (n_n4972)));
	assign x13773x = (((!x24x) & (!x530x) & (!n_n4816) & (!n_n4828) & (n_n4842)) + ((!x24x) & (!x530x) & (!n_n4816) & (n_n4828) & (!n_n4842)) + ((!x24x) & (!x530x) & (!n_n4816) & (n_n4828) & (n_n4842)) + ((!x24x) & (!x530x) & (n_n4816) & (!n_n4828) & (!n_n4842)) + ((!x24x) & (!x530x) & (n_n4816) & (!n_n4828) & (n_n4842)) + ((!x24x) & (!x530x) & (n_n4816) & (n_n4828) & (!n_n4842)) + ((!x24x) & (!x530x) & (n_n4816) & (n_n4828) & (n_n4842)) + ((!x24x) & (x530x) & (!n_n4816) & (!n_n4828) & (n_n4842)) + ((!x24x) & (x530x) & (!n_n4816) & (n_n4828) & (!n_n4842)) + ((!x24x) & (x530x) & (!n_n4816) & (n_n4828) & (n_n4842)) + ((!x24x) & (x530x) & (n_n4816) & (!n_n4828) & (!n_n4842)) + ((!x24x) & (x530x) & (n_n4816) & (!n_n4828) & (n_n4842)) + ((!x24x) & (x530x) & (n_n4816) & (n_n4828) & (!n_n4842)) + ((!x24x) & (x530x) & (n_n4816) & (n_n4828) & (n_n4842)) + ((x24x) & (!x530x) & (!n_n4816) & (!n_n4828) & (n_n4842)) + ((x24x) & (!x530x) & (!n_n4816) & (n_n4828) & (!n_n4842)) + ((x24x) & (!x530x) & (!n_n4816) & (n_n4828) & (n_n4842)) + ((x24x) & (!x530x) & (n_n4816) & (!n_n4828) & (!n_n4842)) + ((x24x) & (!x530x) & (n_n4816) & (!n_n4828) & (n_n4842)) + ((x24x) & (!x530x) & (n_n4816) & (n_n4828) & (!n_n4842)) + ((x24x) & (!x530x) & (n_n4816) & (n_n4828) & (n_n4842)) + ((x24x) & (x530x) & (!n_n4816) & (!n_n4828) & (!n_n4842)) + ((x24x) & (x530x) & (!n_n4816) & (!n_n4828) & (n_n4842)) + ((x24x) & (x530x) & (!n_n4816) & (n_n4828) & (!n_n4842)) + ((x24x) & (x530x) & (!n_n4816) & (n_n4828) & (n_n4842)) + ((x24x) & (x530x) & (n_n4816) & (!n_n4828) & (!n_n4842)) + ((x24x) & (x530x) & (n_n4816) & (!n_n4828) & (n_n4842)) + ((x24x) & (x530x) & (n_n4816) & (n_n4828) & (!n_n4842)) + ((x24x) & (x530x) & (n_n4816) & (n_n4828) & (n_n4842)));
	assign x13774x = (((!x552x) & (!x23x) & (!n_n4844) & (!n_n4818) & (x71x)) + ((!x552x) & (!x23x) & (!n_n4844) & (n_n4818) & (!x71x)) + ((!x552x) & (!x23x) & (!n_n4844) & (n_n4818) & (x71x)) + ((!x552x) & (!x23x) & (n_n4844) & (!n_n4818) & (!x71x)) + ((!x552x) & (!x23x) & (n_n4844) & (!n_n4818) & (x71x)) + ((!x552x) & (!x23x) & (n_n4844) & (n_n4818) & (!x71x)) + ((!x552x) & (!x23x) & (n_n4844) & (n_n4818) & (x71x)) + ((!x552x) & (x23x) & (!n_n4844) & (!n_n4818) & (x71x)) + ((!x552x) & (x23x) & (!n_n4844) & (n_n4818) & (!x71x)) + ((!x552x) & (x23x) & (!n_n4844) & (n_n4818) & (x71x)) + ((!x552x) & (x23x) & (n_n4844) & (!n_n4818) & (!x71x)) + ((!x552x) & (x23x) & (n_n4844) & (!n_n4818) & (x71x)) + ((!x552x) & (x23x) & (n_n4844) & (n_n4818) & (!x71x)) + ((!x552x) & (x23x) & (n_n4844) & (n_n4818) & (x71x)) + ((x552x) & (!x23x) & (!n_n4844) & (!n_n4818) & (x71x)) + ((x552x) & (!x23x) & (!n_n4844) & (n_n4818) & (!x71x)) + ((x552x) & (!x23x) & (!n_n4844) & (n_n4818) & (x71x)) + ((x552x) & (!x23x) & (n_n4844) & (!n_n4818) & (!x71x)) + ((x552x) & (!x23x) & (n_n4844) & (!n_n4818) & (x71x)) + ((x552x) & (!x23x) & (n_n4844) & (n_n4818) & (!x71x)) + ((x552x) & (!x23x) & (n_n4844) & (n_n4818) & (x71x)) + ((x552x) & (x23x) & (!n_n4844) & (!n_n4818) & (!x71x)) + ((x552x) & (x23x) & (!n_n4844) & (!n_n4818) & (x71x)) + ((x552x) & (x23x) & (!n_n4844) & (n_n4818) & (!x71x)) + ((x552x) & (x23x) & (!n_n4844) & (n_n4818) & (x71x)) + ((x552x) & (x23x) & (n_n4844) & (!n_n4818) & (!x71x)) + ((x552x) & (x23x) & (n_n4844) & (!n_n4818) & (x71x)) + ((x552x) & (x23x) & (n_n4844) & (n_n4818) & (!x71x)) + ((x552x) & (x23x) & (n_n4844) & (n_n4818) & (x71x)));
	assign n_n3257 = (((!n_n3272) & (!n_n3274) & (!n_n3322) & (!x13875x) & (x13876x)) + ((!n_n3272) & (!n_n3274) & (!n_n3322) & (x13875x) & (!x13876x)) + ((!n_n3272) & (!n_n3274) & (!n_n3322) & (x13875x) & (x13876x)) + ((!n_n3272) & (!n_n3274) & (n_n3322) & (!x13875x) & (!x13876x)) + ((!n_n3272) & (!n_n3274) & (n_n3322) & (!x13875x) & (x13876x)) + ((!n_n3272) & (!n_n3274) & (n_n3322) & (x13875x) & (!x13876x)) + ((!n_n3272) & (!n_n3274) & (n_n3322) & (x13875x) & (x13876x)) + ((!n_n3272) & (n_n3274) & (!n_n3322) & (!x13875x) & (!x13876x)) + ((!n_n3272) & (n_n3274) & (!n_n3322) & (!x13875x) & (x13876x)) + ((!n_n3272) & (n_n3274) & (!n_n3322) & (x13875x) & (!x13876x)) + ((!n_n3272) & (n_n3274) & (!n_n3322) & (x13875x) & (x13876x)) + ((!n_n3272) & (n_n3274) & (n_n3322) & (!x13875x) & (!x13876x)) + ((!n_n3272) & (n_n3274) & (n_n3322) & (!x13875x) & (x13876x)) + ((!n_n3272) & (n_n3274) & (n_n3322) & (x13875x) & (!x13876x)) + ((!n_n3272) & (n_n3274) & (n_n3322) & (x13875x) & (x13876x)) + ((n_n3272) & (!n_n3274) & (!n_n3322) & (!x13875x) & (!x13876x)) + ((n_n3272) & (!n_n3274) & (!n_n3322) & (!x13875x) & (x13876x)) + ((n_n3272) & (!n_n3274) & (!n_n3322) & (x13875x) & (!x13876x)) + ((n_n3272) & (!n_n3274) & (!n_n3322) & (x13875x) & (x13876x)) + ((n_n3272) & (!n_n3274) & (n_n3322) & (!x13875x) & (!x13876x)) + ((n_n3272) & (!n_n3274) & (n_n3322) & (!x13875x) & (x13876x)) + ((n_n3272) & (!n_n3274) & (n_n3322) & (x13875x) & (!x13876x)) + ((n_n3272) & (!n_n3274) & (n_n3322) & (x13875x) & (x13876x)) + ((n_n3272) & (n_n3274) & (!n_n3322) & (!x13875x) & (!x13876x)) + ((n_n3272) & (n_n3274) & (!n_n3322) & (!x13875x) & (x13876x)) + ((n_n3272) & (n_n3274) & (!n_n3322) & (x13875x) & (!x13876x)) + ((n_n3272) & (n_n3274) & (!n_n3322) & (x13875x) & (x13876x)) + ((n_n3272) & (n_n3274) & (n_n3322) & (!x13875x) & (!x13876x)) + ((n_n3272) & (n_n3274) & (n_n3322) & (!x13875x) & (x13876x)) + ((n_n3272) & (n_n3274) & (n_n3322) & (x13875x) & (!x13876x)) + ((n_n3272) & (n_n3274) & (n_n3322) & (x13875x) & (x13876x)));
	assign n_n3259 = (((!n_n3336) & (!n_n3280) & (!n_n3279) & (!x13916x) & (x13917x)) + ((!n_n3336) & (!n_n3280) & (!n_n3279) & (x13916x) & (!x13917x)) + ((!n_n3336) & (!n_n3280) & (!n_n3279) & (x13916x) & (x13917x)) + ((!n_n3336) & (!n_n3280) & (n_n3279) & (!x13916x) & (!x13917x)) + ((!n_n3336) & (!n_n3280) & (n_n3279) & (!x13916x) & (x13917x)) + ((!n_n3336) & (!n_n3280) & (n_n3279) & (x13916x) & (!x13917x)) + ((!n_n3336) & (!n_n3280) & (n_n3279) & (x13916x) & (x13917x)) + ((!n_n3336) & (n_n3280) & (!n_n3279) & (!x13916x) & (!x13917x)) + ((!n_n3336) & (n_n3280) & (!n_n3279) & (!x13916x) & (x13917x)) + ((!n_n3336) & (n_n3280) & (!n_n3279) & (x13916x) & (!x13917x)) + ((!n_n3336) & (n_n3280) & (!n_n3279) & (x13916x) & (x13917x)) + ((!n_n3336) & (n_n3280) & (n_n3279) & (!x13916x) & (!x13917x)) + ((!n_n3336) & (n_n3280) & (n_n3279) & (!x13916x) & (x13917x)) + ((!n_n3336) & (n_n3280) & (n_n3279) & (x13916x) & (!x13917x)) + ((!n_n3336) & (n_n3280) & (n_n3279) & (x13916x) & (x13917x)) + ((n_n3336) & (!n_n3280) & (!n_n3279) & (!x13916x) & (!x13917x)) + ((n_n3336) & (!n_n3280) & (!n_n3279) & (!x13916x) & (x13917x)) + ((n_n3336) & (!n_n3280) & (!n_n3279) & (x13916x) & (!x13917x)) + ((n_n3336) & (!n_n3280) & (!n_n3279) & (x13916x) & (x13917x)) + ((n_n3336) & (!n_n3280) & (n_n3279) & (!x13916x) & (!x13917x)) + ((n_n3336) & (!n_n3280) & (n_n3279) & (!x13916x) & (x13917x)) + ((n_n3336) & (!n_n3280) & (n_n3279) & (x13916x) & (!x13917x)) + ((n_n3336) & (!n_n3280) & (n_n3279) & (x13916x) & (x13917x)) + ((n_n3336) & (n_n3280) & (!n_n3279) & (!x13916x) & (!x13917x)) + ((n_n3336) & (n_n3280) & (!n_n3279) & (!x13916x) & (x13917x)) + ((n_n3336) & (n_n3280) & (!n_n3279) & (x13916x) & (!x13917x)) + ((n_n3336) & (n_n3280) & (!n_n3279) & (x13916x) & (x13917x)) + ((n_n3336) & (n_n3280) & (n_n3279) & (!x13916x) & (!x13917x)) + ((n_n3336) & (n_n3280) & (n_n3279) & (!x13916x) & (x13917x)) + ((n_n3336) & (n_n3280) & (n_n3279) & (x13916x) & (!x13917x)) + ((n_n3336) & (n_n3280) & (n_n3279) & (x13916x) & (x13917x)));
	assign x14214x = (((!n_n659) & (!n_n5331) & (!n_n3277) & (!n_n3275) & (x13827x)) + ((!n_n659) & (!n_n5331) & (!n_n3277) & (n_n3275) & (!x13827x)) + ((!n_n659) & (!n_n5331) & (!n_n3277) & (n_n3275) & (x13827x)) + ((!n_n659) & (!n_n5331) & (n_n3277) & (!n_n3275) & (!x13827x)) + ((!n_n659) & (!n_n5331) & (n_n3277) & (!n_n3275) & (x13827x)) + ((!n_n659) & (!n_n5331) & (n_n3277) & (n_n3275) & (!x13827x)) + ((!n_n659) & (!n_n5331) & (n_n3277) & (n_n3275) & (x13827x)) + ((!n_n659) & (n_n5331) & (!n_n3277) & (!n_n3275) & (!x13827x)) + ((!n_n659) & (n_n5331) & (!n_n3277) & (!n_n3275) & (x13827x)) + ((!n_n659) & (n_n5331) & (!n_n3277) & (n_n3275) & (!x13827x)) + ((!n_n659) & (n_n5331) & (!n_n3277) & (n_n3275) & (x13827x)) + ((!n_n659) & (n_n5331) & (n_n3277) & (!n_n3275) & (!x13827x)) + ((!n_n659) & (n_n5331) & (n_n3277) & (!n_n3275) & (x13827x)) + ((!n_n659) & (n_n5331) & (n_n3277) & (n_n3275) & (!x13827x)) + ((!n_n659) & (n_n5331) & (n_n3277) & (n_n3275) & (x13827x)) + ((n_n659) & (!n_n5331) & (!n_n3277) & (!n_n3275) & (!x13827x)) + ((n_n659) & (!n_n5331) & (!n_n3277) & (!n_n3275) & (x13827x)) + ((n_n659) & (!n_n5331) & (!n_n3277) & (n_n3275) & (!x13827x)) + ((n_n659) & (!n_n5331) & (!n_n3277) & (n_n3275) & (x13827x)) + ((n_n659) & (!n_n5331) & (n_n3277) & (!n_n3275) & (!x13827x)) + ((n_n659) & (!n_n5331) & (n_n3277) & (!n_n3275) & (x13827x)) + ((n_n659) & (!n_n5331) & (n_n3277) & (n_n3275) & (!x13827x)) + ((n_n659) & (!n_n5331) & (n_n3277) & (n_n3275) & (x13827x)) + ((n_n659) & (n_n5331) & (!n_n3277) & (!n_n3275) & (!x13827x)) + ((n_n659) & (n_n5331) & (!n_n3277) & (!n_n3275) & (x13827x)) + ((n_n659) & (n_n5331) & (!n_n3277) & (n_n3275) & (!x13827x)) + ((n_n659) & (n_n5331) & (!n_n3277) & (n_n3275) & (x13827x)) + ((n_n659) & (n_n5331) & (n_n3277) & (!n_n3275) & (!x13827x)) + ((n_n659) & (n_n5331) & (n_n3277) & (!n_n3275) & (x13827x)) + ((n_n659) & (n_n5331) & (n_n3277) & (n_n3275) & (!x13827x)) + ((n_n659) & (n_n5331) & (n_n3277) & (n_n3275) & (x13827x)));
	assign n_n3546 = (((!x14240x) & (!x14226x) & (!x14227x) & (!x14232x) & (x14233x)) + ((!x14240x) & (!x14226x) & (!x14227x) & (x14232x) & (!x14233x)) + ((!x14240x) & (!x14226x) & (!x14227x) & (x14232x) & (x14233x)) + ((!x14240x) & (!x14226x) & (x14227x) & (!x14232x) & (!x14233x)) + ((!x14240x) & (!x14226x) & (x14227x) & (!x14232x) & (x14233x)) + ((!x14240x) & (!x14226x) & (x14227x) & (x14232x) & (!x14233x)) + ((!x14240x) & (!x14226x) & (x14227x) & (x14232x) & (x14233x)) + ((!x14240x) & (x14226x) & (!x14227x) & (!x14232x) & (!x14233x)) + ((!x14240x) & (x14226x) & (!x14227x) & (!x14232x) & (x14233x)) + ((!x14240x) & (x14226x) & (!x14227x) & (x14232x) & (!x14233x)) + ((!x14240x) & (x14226x) & (!x14227x) & (x14232x) & (x14233x)) + ((!x14240x) & (x14226x) & (x14227x) & (!x14232x) & (!x14233x)) + ((!x14240x) & (x14226x) & (x14227x) & (!x14232x) & (x14233x)) + ((!x14240x) & (x14226x) & (x14227x) & (x14232x) & (!x14233x)) + ((!x14240x) & (x14226x) & (x14227x) & (x14232x) & (x14233x)) + ((x14240x) & (!x14226x) & (!x14227x) & (!x14232x) & (!x14233x)) + ((x14240x) & (!x14226x) & (!x14227x) & (!x14232x) & (x14233x)) + ((x14240x) & (!x14226x) & (!x14227x) & (x14232x) & (!x14233x)) + ((x14240x) & (!x14226x) & (!x14227x) & (x14232x) & (x14233x)) + ((x14240x) & (!x14226x) & (x14227x) & (!x14232x) & (!x14233x)) + ((x14240x) & (!x14226x) & (x14227x) & (!x14232x) & (x14233x)) + ((x14240x) & (!x14226x) & (x14227x) & (x14232x) & (!x14233x)) + ((x14240x) & (!x14226x) & (x14227x) & (x14232x) & (x14233x)) + ((x14240x) & (x14226x) & (!x14227x) & (!x14232x) & (!x14233x)) + ((x14240x) & (x14226x) & (!x14227x) & (!x14232x) & (x14233x)) + ((x14240x) & (x14226x) & (!x14227x) & (x14232x) & (!x14233x)) + ((x14240x) & (x14226x) & (!x14227x) & (x14232x) & (x14233x)) + ((x14240x) & (x14226x) & (x14227x) & (!x14232x) & (!x14233x)) + ((x14240x) & (x14226x) & (x14227x) & (!x14232x) & (x14233x)) + ((x14240x) & (x14226x) & (x14227x) & (x14232x) & (!x14233x)) + ((x14240x) & (x14226x) & (x14227x) & (x14232x) & (x14233x)));
	assign n_n3545 = (((!n_n5307) & (!n_n5266) & (!x14256x) & (!x14246x) & (x63x)) + ((!n_n5307) & (!n_n5266) & (!x14256x) & (x14246x) & (!x63x)) + ((!n_n5307) & (!n_n5266) & (!x14256x) & (x14246x) & (x63x)) + ((!n_n5307) & (!n_n5266) & (x14256x) & (!x14246x) & (!x63x)) + ((!n_n5307) & (!n_n5266) & (x14256x) & (!x14246x) & (x63x)) + ((!n_n5307) & (!n_n5266) & (x14256x) & (x14246x) & (!x63x)) + ((!n_n5307) & (!n_n5266) & (x14256x) & (x14246x) & (x63x)) + ((!n_n5307) & (n_n5266) & (!x14256x) & (!x14246x) & (!x63x)) + ((!n_n5307) & (n_n5266) & (!x14256x) & (!x14246x) & (x63x)) + ((!n_n5307) & (n_n5266) & (!x14256x) & (x14246x) & (!x63x)) + ((!n_n5307) & (n_n5266) & (!x14256x) & (x14246x) & (x63x)) + ((!n_n5307) & (n_n5266) & (x14256x) & (!x14246x) & (!x63x)) + ((!n_n5307) & (n_n5266) & (x14256x) & (!x14246x) & (x63x)) + ((!n_n5307) & (n_n5266) & (x14256x) & (x14246x) & (!x63x)) + ((!n_n5307) & (n_n5266) & (x14256x) & (x14246x) & (x63x)) + ((n_n5307) & (!n_n5266) & (!x14256x) & (!x14246x) & (!x63x)) + ((n_n5307) & (!n_n5266) & (!x14256x) & (!x14246x) & (x63x)) + ((n_n5307) & (!n_n5266) & (!x14256x) & (x14246x) & (!x63x)) + ((n_n5307) & (!n_n5266) & (!x14256x) & (x14246x) & (x63x)) + ((n_n5307) & (!n_n5266) & (x14256x) & (!x14246x) & (!x63x)) + ((n_n5307) & (!n_n5266) & (x14256x) & (!x14246x) & (x63x)) + ((n_n5307) & (!n_n5266) & (x14256x) & (x14246x) & (!x63x)) + ((n_n5307) & (!n_n5266) & (x14256x) & (x14246x) & (x63x)) + ((n_n5307) & (n_n5266) & (!x14256x) & (!x14246x) & (!x63x)) + ((n_n5307) & (n_n5266) & (!x14256x) & (!x14246x) & (x63x)) + ((n_n5307) & (n_n5266) & (!x14256x) & (x14246x) & (!x63x)) + ((n_n5307) & (n_n5266) & (!x14256x) & (x14246x) & (x63x)) + ((n_n5307) & (n_n5266) & (x14256x) & (!x14246x) & (!x63x)) + ((n_n5307) & (n_n5266) & (x14256x) & (!x14246x) & (x63x)) + ((n_n5307) & (n_n5266) & (x14256x) & (x14246x) & (!x63x)) + ((n_n5307) & (n_n5266) & (x14256x) & (x14246x) & (x63x)));
	assign x14275x = (((!n_n5057) & (!n_n4994) & (!n_n4974) & (!x275x) & (x14273x)) + ((!n_n5057) & (!n_n4994) & (!n_n4974) & (x275x) & (!x14273x)) + ((!n_n5057) & (!n_n4994) & (!n_n4974) & (x275x) & (x14273x)) + ((!n_n5057) & (!n_n4994) & (n_n4974) & (!x275x) & (!x14273x)) + ((!n_n5057) & (!n_n4994) & (n_n4974) & (!x275x) & (x14273x)) + ((!n_n5057) & (!n_n4994) & (n_n4974) & (x275x) & (!x14273x)) + ((!n_n5057) & (!n_n4994) & (n_n4974) & (x275x) & (x14273x)) + ((!n_n5057) & (n_n4994) & (!n_n4974) & (!x275x) & (!x14273x)) + ((!n_n5057) & (n_n4994) & (!n_n4974) & (!x275x) & (x14273x)) + ((!n_n5057) & (n_n4994) & (!n_n4974) & (x275x) & (!x14273x)) + ((!n_n5057) & (n_n4994) & (!n_n4974) & (x275x) & (x14273x)) + ((!n_n5057) & (n_n4994) & (n_n4974) & (!x275x) & (!x14273x)) + ((!n_n5057) & (n_n4994) & (n_n4974) & (!x275x) & (x14273x)) + ((!n_n5057) & (n_n4994) & (n_n4974) & (x275x) & (!x14273x)) + ((!n_n5057) & (n_n4994) & (n_n4974) & (x275x) & (x14273x)) + ((n_n5057) & (!n_n4994) & (!n_n4974) & (!x275x) & (!x14273x)) + ((n_n5057) & (!n_n4994) & (!n_n4974) & (!x275x) & (x14273x)) + ((n_n5057) & (!n_n4994) & (!n_n4974) & (x275x) & (!x14273x)) + ((n_n5057) & (!n_n4994) & (!n_n4974) & (x275x) & (x14273x)) + ((n_n5057) & (!n_n4994) & (n_n4974) & (!x275x) & (!x14273x)) + ((n_n5057) & (!n_n4994) & (n_n4974) & (!x275x) & (x14273x)) + ((n_n5057) & (!n_n4994) & (n_n4974) & (x275x) & (!x14273x)) + ((n_n5057) & (!n_n4994) & (n_n4974) & (x275x) & (x14273x)) + ((n_n5057) & (n_n4994) & (!n_n4974) & (!x275x) & (!x14273x)) + ((n_n5057) & (n_n4994) & (!n_n4974) & (!x275x) & (x14273x)) + ((n_n5057) & (n_n4994) & (!n_n4974) & (x275x) & (!x14273x)) + ((n_n5057) & (n_n4994) & (!n_n4974) & (x275x) & (x14273x)) + ((n_n5057) & (n_n4994) & (n_n4974) & (!x275x) & (!x14273x)) + ((n_n5057) & (n_n4994) & (n_n4974) & (!x275x) & (x14273x)) + ((n_n5057) & (n_n4994) & (n_n4974) & (x275x) & (!x14273x)) + ((n_n5057) & (n_n4994) & (n_n4974) & (x275x) & (x14273x)));
	assign x14276x = (((!x14261x) & (!x14262x) & (!x14267x) & (x14268x)) + ((!x14261x) & (!x14262x) & (x14267x) & (!x14268x)) + ((!x14261x) & (!x14262x) & (x14267x) & (x14268x)) + ((!x14261x) & (x14262x) & (!x14267x) & (!x14268x)) + ((!x14261x) & (x14262x) & (!x14267x) & (x14268x)) + ((!x14261x) & (x14262x) & (x14267x) & (!x14268x)) + ((!x14261x) & (x14262x) & (x14267x) & (x14268x)) + ((x14261x) & (!x14262x) & (!x14267x) & (!x14268x)) + ((x14261x) & (!x14262x) & (!x14267x) & (x14268x)) + ((x14261x) & (!x14262x) & (x14267x) & (!x14268x)) + ((x14261x) & (!x14262x) & (x14267x) & (x14268x)) + ((x14261x) & (x14262x) & (!x14267x) & (!x14268x)) + ((x14261x) & (x14262x) & (!x14267x) & (x14268x)) + ((x14261x) & (x14262x) & (x14267x) & (!x14268x)) + ((x14261x) & (x14262x) & (x14267x) & (x14268x)));
	assign n_n3543 = (((!n_n3546) & (!n_n3545) & (!x14275x) & (x14276x)) + ((!n_n3546) & (!n_n3545) & (x14275x) & (!x14276x)) + ((!n_n3546) & (!n_n3545) & (x14275x) & (x14276x)) + ((!n_n3546) & (n_n3545) & (!x14275x) & (!x14276x)) + ((!n_n3546) & (n_n3545) & (!x14275x) & (x14276x)) + ((!n_n3546) & (n_n3545) & (x14275x) & (!x14276x)) + ((!n_n3546) & (n_n3545) & (x14275x) & (x14276x)) + ((n_n3546) & (!n_n3545) & (!x14275x) & (!x14276x)) + ((n_n3546) & (!n_n3545) & (!x14275x) & (x14276x)) + ((n_n3546) & (!n_n3545) & (x14275x) & (!x14276x)) + ((n_n3546) & (!n_n3545) & (x14275x) & (x14276x)) + ((n_n3546) & (n_n3545) & (!x14275x) & (!x14276x)) + ((n_n3546) & (n_n3545) & (!x14275x) & (x14276x)) + ((n_n3546) & (n_n3545) & (x14275x) & (!x14276x)) + ((n_n3546) & (n_n3545) & (x14275x) & (x14276x)));
	assign n_n3549 = (((!n_n3562) & (!x14301x) & (!x14302x) & (!x14308x) & (x14309x)) + ((!n_n3562) & (!x14301x) & (!x14302x) & (x14308x) & (!x14309x)) + ((!n_n3562) & (!x14301x) & (!x14302x) & (x14308x) & (x14309x)) + ((!n_n3562) & (!x14301x) & (x14302x) & (!x14308x) & (!x14309x)) + ((!n_n3562) & (!x14301x) & (x14302x) & (!x14308x) & (x14309x)) + ((!n_n3562) & (!x14301x) & (x14302x) & (x14308x) & (!x14309x)) + ((!n_n3562) & (!x14301x) & (x14302x) & (x14308x) & (x14309x)) + ((!n_n3562) & (x14301x) & (!x14302x) & (!x14308x) & (!x14309x)) + ((!n_n3562) & (x14301x) & (!x14302x) & (!x14308x) & (x14309x)) + ((!n_n3562) & (x14301x) & (!x14302x) & (x14308x) & (!x14309x)) + ((!n_n3562) & (x14301x) & (!x14302x) & (x14308x) & (x14309x)) + ((!n_n3562) & (x14301x) & (x14302x) & (!x14308x) & (!x14309x)) + ((!n_n3562) & (x14301x) & (x14302x) & (!x14308x) & (x14309x)) + ((!n_n3562) & (x14301x) & (x14302x) & (x14308x) & (!x14309x)) + ((!n_n3562) & (x14301x) & (x14302x) & (x14308x) & (x14309x)) + ((n_n3562) & (!x14301x) & (!x14302x) & (!x14308x) & (!x14309x)) + ((n_n3562) & (!x14301x) & (!x14302x) & (!x14308x) & (x14309x)) + ((n_n3562) & (!x14301x) & (!x14302x) & (x14308x) & (!x14309x)) + ((n_n3562) & (!x14301x) & (!x14302x) & (x14308x) & (x14309x)) + ((n_n3562) & (!x14301x) & (x14302x) & (!x14308x) & (!x14309x)) + ((n_n3562) & (!x14301x) & (x14302x) & (!x14308x) & (x14309x)) + ((n_n3562) & (!x14301x) & (x14302x) & (x14308x) & (!x14309x)) + ((n_n3562) & (!x14301x) & (x14302x) & (x14308x) & (x14309x)) + ((n_n3562) & (x14301x) & (!x14302x) & (!x14308x) & (!x14309x)) + ((n_n3562) & (x14301x) & (!x14302x) & (!x14308x) & (x14309x)) + ((n_n3562) & (x14301x) & (!x14302x) & (x14308x) & (!x14309x)) + ((n_n3562) & (x14301x) & (!x14302x) & (x14308x) & (x14309x)) + ((n_n3562) & (x14301x) & (x14302x) & (!x14308x) & (!x14309x)) + ((n_n3562) & (x14301x) & (x14302x) & (!x14308x) & (x14309x)) + ((n_n3562) & (x14301x) & (x14302x) & (x14308x) & (!x14309x)) + ((n_n3562) & (x14301x) & (x14302x) & (x14308x) & (x14309x)));
	assign x14332x = (((!n_n4759) & (!n_n4811) & (!n_n4793) & (!n_n4778) & (x14331x)) + ((!n_n4759) & (!n_n4811) & (!n_n4793) & (n_n4778) & (!x14331x)) + ((!n_n4759) & (!n_n4811) & (!n_n4793) & (n_n4778) & (x14331x)) + ((!n_n4759) & (!n_n4811) & (n_n4793) & (!n_n4778) & (!x14331x)) + ((!n_n4759) & (!n_n4811) & (n_n4793) & (!n_n4778) & (x14331x)) + ((!n_n4759) & (!n_n4811) & (n_n4793) & (n_n4778) & (!x14331x)) + ((!n_n4759) & (!n_n4811) & (n_n4793) & (n_n4778) & (x14331x)) + ((!n_n4759) & (n_n4811) & (!n_n4793) & (!n_n4778) & (!x14331x)) + ((!n_n4759) & (n_n4811) & (!n_n4793) & (!n_n4778) & (x14331x)) + ((!n_n4759) & (n_n4811) & (!n_n4793) & (n_n4778) & (!x14331x)) + ((!n_n4759) & (n_n4811) & (!n_n4793) & (n_n4778) & (x14331x)) + ((!n_n4759) & (n_n4811) & (n_n4793) & (!n_n4778) & (!x14331x)) + ((!n_n4759) & (n_n4811) & (n_n4793) & (!n_n4778) & (x14331x)) + ((!n_n4759) & (n_n4811) & (n_n4793) & (n_n4778) & (!x14331x)) + ((!n_n4759) & (n_n4811) & (n_n4793) & (n_n4778) & (x14331x)) + ((n_n4759) & (!n_n4811) & (!n_n4793) & (!n_n4778) & (!x14331x)) + ((n_n4759) & (!n_n4811) & (!n_n4793) & (!n_n4778) & (x14331x)) + ((n_n4759) & (!n_n4811) & (!n_n4793) & (n_n4778) & (!x14331x)) + ((n_n4759) & (!n_n4811) & (!n_n4793) & (n_n4778) & (x14331x)) + ((n_n4759) & (!n_n4811) & (n_n4793) & (!n_n4778) & (!x14331x)) + ((n_n4759) & (!n_n4811) & (n_n4793) & (!n_n4778) & (x14331x)) + ((n_n4759) & (!n_n4811) & (n_n4793) & (n_n4778) & (!x14331x)) + ((n_n4759) & (!n_n4811) & (n_n4793) & (n_n4778) & (x14331x)) + ((n_n4759) & (n_n4811) & (!n_n4793) & (!n_n4778) & (!x14331x)) + ((n_n4759) & (n_n4811) & (!n_n4793) & (!n_n4778) & (x14331x)) + ((n_n4759) & (n_n4811) & (!n_n4793) & (n_n4778) & (!x14331x)) + ((n_n4759) & (n_n4811) & (!n_n4793) & (n_n4778) & (x14331x)) + ((n_n4759) & (n_n4811) & (n_n4793) & (!n_n4778) & (!x14331x)) + ((n_n4759) & (n_n4811) & (n_n4793) & (!n_n4778) & (x14331x)) + ((n_n4759) & (n_n4811) & (n_n4793) & (n_n4778) & (!x14331x)) + ((n_n4759) & (n_n4811) & (n_n4793) & (n_n4778) & (x14331x)));
	assign x14333x = (((!x14317x) & (!x14318x) & (!x14323x) & (x14324x)) + ((!x14317x) & (!x14318x) & (x14323x) & (!x14324x)) + ((!x14317x) & (!x14318x) & (x14323x) & (x14324x)) + ((!x14317x) & (x14318x) & (!x14323x) & (!x14324x)) + ((!x14317x) & (x14318x) & (!x14323x) & (x14324x)) + ((!x14317x) & (x14318x) & (x14323x) & (!x14324x)) + ((!x14317x) & (x14318x) & (x14323x) & (x14324x)) + ((x14317x) & (!x14318x) & (!x14323x) & (!x14324x)) + ((x14317x) & (!x14318x) & (!x14323x) & (x14324x)) + ((x14317x) & (!x14318x) & (x14323x) & (!x14324x)) + ((x14317x) & (!x14318x) & (x14323x) & (x14324x)) + ((x14317x) & (x14318x) & (!x14323x) & (!x14324x)) + ((x14317x) & (x14318x) & (!x14323x) & (x14324x)) + ((x14317x) & (x14318x) & (x14323x) & (!x14324x)) + ((x14317x) & (x14318x) & (x14323x) & (x14324x)));
	assign x14341x = (((!n_n3565) & (!x14290x) & (!x14291x) & (x14339x)) + ((!n_n3565) & (!x14290x) & (x14291x) & (!x14339x)) + ((!n_n3565) & (!x14290x) & (x14291x) & (x14339x)) + ((!n_n3565) & (x14290x) & (!x14291x) & (!x14339x)) + ((!n_n3565) & (x14290x) & (!x14291x) & (x14339x)) + ((!n_n3565) & (x14290x) & (x14291x) & (!x14339x)) + ((!n_n3565) & (x14290x) & (x14291x) & (x14339x)) + ((n_n3565) & (!x14290x) & (!x14291x) & (!x14339x)) + ((n_n3565) & (!x14290x) & (!x14291x) & (x14339x)) + ((n_n3565) & (!x14290x) & (x14291x) & (!x14339x)) + ((n_n3565) & (!x14290x) & (x14291x) & (x14339x)) + ((n_n3565) & (x14290x) & (!x14291x) & (!x14339x)) + ((n_n3565) & (x14290x) & (!x14291x) & (x14339x)) + ((n_n3565) & (x14290x) & (x14291x) & (!x14339x)) + ((n_n3565) & (x14290x) & (x14291x) & (x14339x)));
	assign x14343x = (((!n_n3549) & (!x14332x) & (!x14333x) & (x14341x)) + ((!n_n3549) & (!x14332x) & (x14333x) & (!x14341x)) + ((!n_n3549) & (!x14332x) & (x14333x) & (x14341x)) + ((!n_n3549) & (x14332x) & (!x14333x) & (!x14341x)) + ((!n_n3549) & (x14332x) & (!x14333x) & (x14341x)) + ((!n_n3549) & (x14332x) & (x14333x) & (!x14341x)) + ((!n_n3549) & (x14332x) & (x14333x) & (x14341x)) + ((n_n3549) & (!x14332x) & (!x14333x) & (!x14341x)) + ((n_n3549) & (!x14332x) & (!x14333x) & (x14341x)) + ((n_n3549) & (!x14332x) & (x14333x) & (!x14341x)) + ((n_n3549) & (!x14332x) & (x14333x) & (x14341x)) + ((n_n3549) & (x14332x) & (!x14333x) & (!x14341x)) + ((n_n3549) & (x14332x) & (!x14333x) & (x14341x)) + ((n_n3549) & (x14332x) & (x14333x) & (!x14341x)) + ((n_n3549) & (x14332x) & (x14333x) & (x14341x)));
	assign x350x = (((!i_9_) & (n_n532) & (n_n325) & (n_n491) & (!n_n530)) + ((!i_9_) & (n_n532) & (n_n325) & (n_n491) & (n_n530)) + ((i_9_) & (!n_n532) & (n_n325) & (n_n491) & (n_n530)) + ((i_9_) & (n_n532) & (n_n325) & (n_n491) & (n_n530)));
	assign x370x = (((!i_9_) & (!n_n534) & (!n_n325) & (!n_n491) & (n_n4758)) + ((!i_9_) & (!n_n534) & (!n_n325) & (n_n491) & (n_n4758)) + ((!i_9_) & (!n_n534) & (n_n325) & (!n_n491) & (n_n4758)) + ((!i_9_) & (!n_n534) & (n_n325) & (n_n491) & (n_n4758)) + ((!i_9_) & (n_n534) & (!n_n325) & (!n_n491) & (n_n4758)) + ((!i_9_) & (n_n534) & (!n_n325) & (n_n491) & (n_n4758)) + ((!i_9_) & (n_n534) & (n_n325) & (!n_n491) & (n_n4758)) + ((!i_9_) & (n_n534) & (n_n325) & (n_n491) & (n_n4758)) + ((i_9_) & (!n_n534) & (!n_n325) & (!n_n491) & (n_n4758)) + ((i_9_) & (!n_n534) & (!n_n325) & (n_n491) & (n_n4758)) + ((i_9_) & (!n_n534) & (n_n325) & (!n_n491) & (n_n4758)) + ((i_9_) & (!n_n534) & (n_n325) & (n_n491) & (n_n4758)) + ((i_9_) & (n_n534) & (!n_n325) & (!n_n491) & (n_n4758)) + ((i_9_) & (n_n534) & (!n_n325) & (n_n491) & (n_n4758)) + ((i_9_) & (n_n534) & (n_n325) & (!n_n491) & (n_n4758)) + ((i_9_) & (n_n534) & (n_n325) & (n_n491) & (!n_n4758)) + ((i_9_) & (n_n534) & (n_n325) & (n_n491) & (n_n4758)));
	assign x14376x = (((!n_n4761) & (!n_n4762) & (!n_n4767) & (!n_n4765) & (n_n4766)) + ((!n_n4761) & (!n_n4762) & (!n_n4767) & (n_n4765) & (!n_n4766)) + ((!n_n4761) & (!n_n4762) & (!n_n4767) & (n_n4765) & (n_n4766)) + ((!n_n4761) & (!n_n4762) & (n_n4767) & (!n_n4765) & (!n_n4766)) + ((!n_n4761) & (!n_n4762) & (n_n4767) & (!n_n4765) & (n_n4766)) + ((!n_n4761) & (!n_n4762) & (n_n4767) & (n_n4765) & (!n_n4766)) + ((!n_n4761) & (!n_n4762) & (n_n4767) & (n_n4765) & (n_n4766)) + ((!n_n4761) & (n_n4762) & (!n_n4767) & (!n_n4765) & (!n_n4766)) + ((!n_n4761) & (n_n4762) & (!n_n4767) & (!n_n4765) & (n_n4766)) + ((!n_n4761) & (n_n4762) & (!n_n4767) & (n_n4765) & (!n_n4766)) + ((!n_n4761) & (n_n4762) & (!n_n4767) & (n_n4765) & (n_n4766)) + ((!n_n4761) & (n_n4762) & (n_n4767) & (!n_n4765) & (!n_n4766)) + ((!n_n4761) & (n_n4762) & (n_n4767) & (!n_n4765) & (n_n4766)) + ((!n_n4761) & (n_n4762) & (n_n4767) & (n_n4765) & (!n_n4766)) + ((!n_n4761) & (n_n4762) & (n_n4767) & (n_n4765) & (n_n4766)) + ((n_n4761) & (!n_n4762) & (!n_n4767) & (!n_n4765) & (!n_n4766)) + ((n_n4761) & (!n_n4762) & (!n_n4767) & (!n_n4765) & (n_n4766)) + ((n_n4761) & (!n_n4762) & (!n_n4767) & (n_n4765) & (!n_n4766)) + ((n_n4761) & (!n_n4762) & (!n_n4767) & (n_n4765) & (n_n4766)) + ((n_n4761) & (!n_n4762) & (n_n4767) & (!n_n4765) & (!n_n4766)) + ((n_n4761) & (!n_n4762) & (n_n4767) & (!n_n4765) & (n_n4766)) + ((n_n4761) & (!n_n4762) & (n_n4767) & (n_n4765) & (!n_n4766)) + ((n_n4761) & (!n_n4762) & (n_n4767) & (n_n4765) & (n_n4766)) + ((n_n4761) & (n_n4762) & (!n_n4767) & (!n_n4765) & (!n_n4766)) + ((n_n4761) & (n_n4762) & (!n_n4767) & (!n_n4765) & (n_n4766)) + ((n_n4761) & (n_n4762) & (!n_n4767) & (n_n4765) & (!n_n4766)) + ((n_n4761) & (n_n4762) & (!n_n4767) & (n_n4765) & (n_n4766)) + ((n_n4761) & (n_n4762) & (n_n4767) & (!n_n4765) & (!n_n4766)) + ((n_n4761) & (n_n4762) & (n_n4767) & (!n_n4765) & (n_n4766)) + ((n_n4761) & (n_n4762) & (n_n4767) & (n_n4765) & (!n_n4766)) + ((n_n4761) & (n_n4762) & (n_n4767) & (n_n4765) & (n_n4766)));
	assign n_n3707 = (((!x95x) & (!n_n4728) & (!n_n4730) & (!n_n4742) & (!x22104x)) + ((!x95x) & (!n_n4728) & (!n_n4730) & (n_n4742) & (!x22104x)) + ((!x95x) & (!n_n4728) & (!n_n4730) & (n_n4742) & (x22104x)) + ((!x95x) & (!n_n4728) & (n_n4730) & (!n_n4742) & (!x22104x)) + ((!x95x) & (!n_n4728) & (n_n4730) & (!n_n4742) & (x22104x)) + ((!x95x) & (!n_n4728) & (n_n4730) & (n_n4742) & (!x22104x)) + ((!x95x) & (!n_n4728) & (n_n4730) & (n_n4742) & (x22104x)) + ((!x95x) & (n_n4728) & (!n_n4730) & (!n_n4742) & (!x22104x)) + ((!x95x) & (n_n4728) & (!n_n4730) & (!n_n4742) & (x22104x)) + ((!x95x) & (n_n4728) & (!n_n4730) & (n_n4742) & (!x22104x)) + ((!x95x) & (n_n4728) & (!n_n4730) & (n_n4742) & (x22104x)) + ((!x95x) & (n_n4728) & (n_n4730) & (!n_n4742) & (!x22104x)) + ((!x95x) & (n_n4728) & (n_n4730) & (!n_n4742) & (x22104x)) + ((!x95x) & (n_n4728) & (n_n4730) & (n_n4742) & (!x22104x)) + ((!x95x) & (n_n4728) & (n_n4730) & (n_n4742) & (x22104x)) + ((x95x) & (!n_n4728) & (!n_n4730) & (!n_n4742) & (!x22104x)) + ((x95x) & (!n_n4728) & (!n_n4730) & (!n_n4742) & (x22104x)) + ((x95x) & (!n_n4728) & (!n_n4730) & (n_n4742) & (!x22104x)) + ((x95x) & (!n_n4728) & (!n_n4730) & (n_n4742) & (x22104x)) + ((x95x) & (!n_n4728) & (n_n4730) & (!n_n4742) & (!x22104x)) + ((x95x) & (!n_n4728) & (n_n4730) & (!n_n4742) & (x22104x)) + ((x95x) & (!n_n4728) & (n_n4730) & (n_n4742) & (!x22104x)) + ((x95x) & (!n_n4728) & (n_n4730) & (n_n4742) & (x22104x)) + ((x95x) & (n_n4728) & (!n_n4730) & (!n_n4742) & (!x22104x)) + ((x95x) & (n_n4728) & (!n_n4730) & (!n_n4742) & (x22104x)) + ((x95x) & (n_n4728) & (!n_n4730) & (n_n4742) & (!x22104x)) + ((x95x) & (n_n4728) & (!n_n4730) & (n_n4742) & (x22104x)) + ((x95x) & (n_n4728) & (n_n4730) & (!n_n4742) & (!x22104x)) + ((x95x) & (n_n4728) & (n_n4730) & (!n_n4742) & (x22104x)) + ((x95x) & (n_n4728) & (n_n4730) & (n_n4742) & (!x22104x)) + ((x95x) & (n_n4728) & (n_n4730) & (n_n4742) & (x22104x)));
	assign x14386x = (((!x109x) & (!n_n4743) & (!n_n4745) & (!n_n4210) & (x14382x)) + ((!x109x) & (!n_n4743) & (!n_n4745) & (n_n4210) & (!x14382x)) + ((!x109x) & (!n_n4743) & (!n_n4745) & (n_n4210) & (x14382x)) + ((!x109x) & (!n_n4743) & (n_n4745) & (!n_n4210) & (!x14382x)) + ((!x109x) & (!n_n4743) & (n_n4745) & (!n_n4210) & (x14382x)) + ((!x109x) & (!n_n4743) & (n_n4745) & (n_n4210) & (!x14382x)) + ((!x109x) & (!n_n4743) & (n_n4745) & (n_n4210) & (x14382x)) + ((!x109x) & (n_n4743) & (!n_n4745) & (!n_n4210) & (!x14382x)) + ((!x109x) & (n_n4743) & (!n_n4745) & (!n_n4210) & (x14382x)) + ((!x109x) & (n_n4743) & (!n_n4745) & (n_n4210) & (!x14382x)) + ((!x109x) & (n_n4743) & (!n_n4745) & (n_n4210) & (x14382x)) + ((!x109x) & (n_n4743) & (n_n4745) & (!n_n4210) & (!x14382x)) + ((!x109x) & (n_n4743) & (n_n4745) & (!n_n4210) & (x14382x)) + ((!x109x) & (n_n4743) & (n_n4745) & (n_n4210) & (!x14382x)) + ((!x109x) & (n_n4743) & (n_n4745) & (n_n4210) & (x14382x)) + ((x109x) & (!n_n4743) & (!n_n4745) & (!n_n4210) & (!x14382x)) + ((x109x) & (!n_n4743) & (!n_n4745) & (!n_n4210) & (x14382x)) + ((x109x) & (!n_n4743) & (!n_n4745) & (n_n4210) & (!x14382x)) + ((x109x) & (!n_n4743) & (!n_n4745) & (n_n4210) & (x14382x)) + ((x109x) & (!n_n4743) & (n_n4745) & (!n_n4210) & (!x14382x)) + ((x109x) & (!n_n4743) & (n_n4745) & (!n_n4210) & (x14382x)) + ((x109x) & (!n_n4743) & (n_n4745) & (n_n4210) & (!x14382x)) + ((x109x) & (!n_n4743) & (n_n4745) & (n_n4210) & (x14382x)) + ((x109x) & (n_n4743) & (!n_n4745) & (!n_n4210) & (!x14382x)) + ((x109x) & (n_n4743) & (!n_n4745) & (!n_n4210) & (x14382x)) + ((x109x) & (n_n4743) & (!n_n4745) & (n_n4210) & (!x14382x)) + ((x109x) & (n_n4743) & (!n_n4745) & (n_n4210) & (x14382x)) + ((x109x) & (n_n4743) & (n_n4745) & (!n_n4210) & (!x14382x)) + ((x109x) & (n_n4743) & (n_n4745) & (!n_n4210) & (x14382x)) + ((x109x) & (n_n4743) & (n_n4745) & (n_n4210) & (!x14382x)) + ((x109x) & (n_n4743) & (n_n4745) & (n_n4210) & (x14382x)));
	assign x14388x = (((!x350x) & (!x370x) & (!x14376x) & (!n_n3707) & (x14386x)) + ((!x350x) & (!x370x) & (!x14376x) & (n_n3707) & (!x14386x)) + ((!x350x) & (!x370x) & (!x14376x) & (n_n3707) & (x14386x)) + ((!x350x) & (!x370x) & (x14376x) & (!n_n3707) & (!x14386x)) + ((!x350x) & (!x370x) & (x14376x) & (!n_n3707) & (x14386x)) + ((!x350x) & (!x370x) & (x14376x) & (n_n3707) & (!x14386x)) + ((!x350x) & (!x370x) & (x14376x) & (n_n3707) & (x14386x)) + ((!x350x) & (x370x) & (!x14376x) & (!n_n3707) & (!x14386x)) + ((!x350x) & (x370x) & (!x14376x) & (!n_n3707) & (x14386x)) + ((!x350x) & (x370x) & (!x14376x) & (n_n3707) & (!x14386x)) + ((!x350x) & (x370x) & (!x14376x) & (n_n3707) & (x14386x)) + ((!x350x) & (x370x) & (x14376x) & (!n_n3707) & (!x14386x)) + ((!x350x) & (x370x) & (x14376x) & (!n_n3707) & (x14386x)) + ((!x350x) & (x370x) & (x14376x) & (n_n3707) & (!x14386x)) + ((!x350x) & (x370x) & (x14376x) & (n_n3707) & (x14386x)) + ((x350x) & (!x370x) & (!x14376x) & (!n_n3707) & (!x14386x)) + ((x350x) & (!x370x) & (!x14376x) & (!n_n3707) & (x14386x)) + ((x350x) & (!x370x) & (!x14376x) & (n_n3707) & (!x14386x)) + ((x350x) & (!x370x) & (!x14376x) & (n_n3707) & (x14386x)) + ((x350x) & (!x370x) & (x14376x) & (!n_n3707) & (!x14386x)) + ((x350x) & (!x370x) & (x14376x) & (!n_n3707) & (x14386x)) + ((x350x) & (!x370x) & (x14376x) & (n_n3707) & (!x14386x)) + ((x350x) & (!x370x) & (x14376x) & (n_n3707) & (x14386x)) + ((x350x) & (x370x) & (!x14376x) & (!n_n3707) & (!x14386x)) + ((x350x) & (x370x) & (!x14376x) & (!n_n3707) & (x14386x)) + ((x350x) & (x370x) & (!x14376x) & (n_n3707) & (!x14386x)) + ((x350x) & (x370x) & (!x14376x) & (n_n3707) & (x14386x)) + ((x350x) & (x370x) & (x14376x) & (!n_n3707) & (!x14386x)) + ((x350x) & (x370x) & (x14376x) & (!n_n3707) & (x14386x)) + ((x350x) & (x370x) & (x14376x) & (n_n3707) & (!x14386x)) + ((x350x) & (x370x) & (x14376x) & (n_n3707) & (x14386x)));
	assign n_n3653 = (((!x14448x) & (!x14449x) & (!x14455x) & (!x14456x) & (x14457x)) + ((!x14448x) & (!x14449x) & (!x14455x) & (x14456x) & (!x14457x)) + ((!x14448x) & (!x14449x) & (!x14455x) & (x14456x) & (x14457x)) + ((!x14448x) & (!x14449x) & (x14455x) & (!x14456x) & (!x14457x)) + ((!x14448x) & (!x14449x) & (x14455x) & (!x14456x) & (x14457x)) + ((!x14448x) & (!x14449x) & (x14455x) & (x14456x) & (!x14457x)) + ((!x14448x) & (!x14449x) & (x14455x) & (x14456x) & (x14457x)) + ((!x14448x) & (x14449x) & (!x14455x) & (!x14456x) & (!x14457x)) + ((!x14448x) & (x14449x) & (!x14455x) & (!x14456x) & (x14457x)) + ((!x14448x) & (x14449x) & (!x14455x) & (x14456x) & (!x14457x)) + ((!x14448x) & (x14449x) & (!x14455x) & (x14456x) & (x14457x)) + ((!x14448x) & (x14449x) & (x14455x) & (!x14456x) & (!x14457x)) + ((!x14448x) & (x14449x) & (x14455x) & (!x14456x) & (x14457x)) + ((!x14448x) & (x14449x) & (x14455x) & (x14456x) & (!x14457x)) + ((!x14448x) & (x14449x) & (x14455x) & (x14456x) & (x14457x)) + ((x14448x) & (!x14449x) & (!x14455x) & (!x14456x) & (!x14457x)) + ((x14448x) & (!x14449x) & (!x14455x) & (!x14456x) & (x14457x)) + ((x14448x) & (!x14449x) & (!x14455x) & (x14456x) & (!x14457x)) + ((x14448x) & (!x14449x) & (!x14455x) & (x14456x) & (x14457x)) + ((x14448x) & (!x14449x) & (x14455x) & (!x14456x) & (!x14457x)) + ((x14448x) & (!x14449x) & (x14455x) & (!x14456x) & (x14457x)) + ((x14448x) & (!x14449x) & (x14455x) & (x14456x) & (!x14457x)) + ((x14448x) & (!x14449x) & (x14455x) & (x14456x) & (x14457x)) + ((x14448x) & (x14449x) & (!x14455x) & (!x14456x) & (!x14457x)) + ((x14448x) & (x14449x) & (!x14455x) & (!x14456x) & (x14457x)) + ((x14448x) & (x14449x) & (!x14455x) & (x14456x) & (!x14457x)) + ((x14448x) & (x14449x) & (!x14455x) & (x14456x) & (x14457x)) + ((x14448x) & (x14449x) & (x14455x) & (!x14456x) & (!x14457x)) + ((x14448x) & (x14449x) & (x14455x) & (!x14456x) & (x14457x)) + ((x14448x) & (x14449x) & (x14455x) & (x14456x) & (!x14457x)) + ((x14448x) & (x14449x) & (x14455x) & (x14456x) & (x14457x)));
	assign x14530x = (((!n_n4444) & (!n_n4445) & (!n_n4442) & (!x22165x)) + ((!n_n4444) & (!n_n4445) & (n_n4442) & (!x22165x)) + ((!n_n4444) & (!n_n4445) & (n_n4442) & (x22165x)) + ((!n_n4444) & (n_n4445) & (!n_n4442) & (!x22165x)) + ((!n_n4444) & (n_n4445) & (!n_n4442) & (x22165x)) + ((!n_n4444) & (n_n4445) & (n_n4442) & (!x22165x)) + ((!n_n4444) & (n_n4445) & (n_n4442) & (x22165x)) + ((n_n4444) & (!n_n4445) & (!n_n4442) & (!x22165x)) + ((n_n4444) & (!n_n4445) & (!n_n4442) & (x22165x)) + ((n_n4444) & (!n_n4445) & (n_n4442) & (!x22165x)) + ((n_n4444) & (!n_n4445) & (n_n4442) & (x22165x)) + ((n_n4444) & (n_n4445) & (!n_n4442) & (!x22165x)) + ((n_n4444) & (n_n4445) & (!n_n4442) & (x22165x)) + ((n_n4444) & (n_n4445) & (n_n4442) & (!x22165x)) + ((n_n4444) & (n_n4445) & (n_n4442) & (x22165x)));
	assign n_n3729 = (((!x15x) & (!n_n518) & (!n_n455) & (!x321x) & (n_n4458)) + ((!x15x) & (!n_n518) & (!n_n455) & (x321x) & (!n_n4458)) + ((!x15x) & (!n_n518) & (!n_n455) & (x321x) & (n_n4458)) + ((!x15x) & (!n_n518) & (n_n455) & (!x321x) & (n_n4458)) + ((!x15x) & (!n_n518) & (n_n455) & (x321x) & (!n_n4458)) + ((!x15x) & (!n_n518) & (n_n455) & (x321x) & (n_n4458)) + ((!x15x) & (n_n518) & (!n_n455) & (!x321x) & (n_n4458)) + ((!x15x) & (n_n518) & (!n_n455) & (x321x) & (!n_n4458)) + ((!x15x) & (n_n518) & (!n_n455) & (x321x) & (n_n4458)) + ((!x15x) & (n_n518) & (n_n455) & (!x321x) & (n_n4458)) + ((!x15x) & (n_n518) & (n_n455) & (x321x) & (!n_n4458)) + ((!x15x) & (n_n518) & (n_n455) & (x321x) & (n_n4458)) + ((x15x) & (!n_n518) & (!n_n455) & (!x321x) & (n_n4458)) + ((x15x) & (!n_n518) & (!n_n455) & (x321x) & (!n_n4458)) + ((x15x) & (!n_n518) & (!n_n455) & (x321x) & (n_n4458)) + ((x15x) & (!n_n518) & (n_n455) & (!x321x) & (n_n4458)) + ((x15x) & (!n_n518) & (n_n455) & (x321x) & (!n_n4458)) + ((x15x) & (!n_n518) & (n_n455) & (x321x) & (n_n4458)) + ((x15x) & (n_n518) & (!n_n455) & (!x321x) & (n_n4458)) + ((x15x) & (n_n518) & (!n_n455) & (x321x) & (!n_n4458)) + ((x15x) & (n_n518) & (!n_n455) & (x321x) & (n_n4458)) + ((x15x) & (n_n518) & (n_n455) & (!x321x) & (!n_n4458)) + ((x15x) & (n_n518) & (n_n455) & (!x321x) & (n_n4458)) + ((x15x) & (n_n518) & (n_n455) & (x321x) & (!n_n4458)) + ((x15x) & (n_n518) & (n_n455) & (x321x) & (n_n4458)));
	assign n_n3731 = (((!n_n4434) & (!x98x) & (!n_n4426) & (!n_n2802) & (x215x)) + ((!n_n4434) & (!x98x) & (!n_n4426) & (n_n2802) & (!x215x)) + ((!n_n4434) & (!x98x) & (!n_n4426) & (n_n2802) & (x215x)) + ((!n_n4434) & (!x98x) & (n_n4426) & (!n_n2802) & (!x215x)) + ((!n_n4434) & (!x98x) & (n_n4426) & (!n_n2802) & (x215x)) + ((!n_n4434) & (!x98x) & (n_n4426) & (n_n2802) & (!x215x)) + ((!n_n4434) & (!x98x) & (n_n4426) & (n_n2802) & (x215x)) + ((!n_n4434) & (x98x) & (!n_n4426) & (!n_n2802) & (!x215x)) + ((!n_n4434) & (x98x) & (!n_n4426) & (!n_n2802) & (x215x)) + ((!n_n4434) & (x98x) & (!n_n4426) & (n_n2802) & (!x215x)) + ((!n_n4434) & (x98x) & (!n_n4426) & (n_n2802) & (x215x)) + ((!n_n4434) & (x98x) & (n_n4426) & (!n_n2802) & (!x215x)) + ((!n_n4434) & (x98x) & (n_n4426) & (!n_n2802) & (x215x)) + ((!n_n4434) & (x98x) & (n_n4426) & (n_n2802) & (!x215x)) + ((!n_n4434) & (x98x) & (n_n4426) & (n_n2802) & (x215x)) + ((n_n4434) & (!x98x) & (!n_n4426) & (!n_n2802) & (!x215x)) + ((n_n4434) & (!x98x) & (!n_n4426) & (!n_n2802) & (x215x)) + ((n_n4434) & (!x98x) & (!n_n4426) & (n_n2802) & (!x215x)) + ((n_n4434) & (!x98x) & (!n_n4426) & (n_n2802) & (x215x)) + ((n_n4434) & (!x98x) & (n_n4426) & (!n_n2802) & (!x215x)) + ((n_n4434) & (!x98x) & (n_n4426) & (!n_n2802) & (x215x)) + ((n_n4434) & (!x98x) & (n_n4426) & (n_n2802) & (!x215x)) + ((n_n4434) & (!x98x) & (n_n4426) & (n_n2802) & (x215x)) + ((n_n4434) & (x98x) & (!n_n4426) & (!n_n2802) & (!x215x)) + ((n_n4434) & (x98x) & (!n_n4426) & (!n_n2802) & (x215x)) + ((n_n4434) & (x98x) & (!n_n4426) & (n_n2802) & (!x215x)) + ((n_n4434) & (x98x) & (!n_n4426) & (n_n2802) & (x215x)) + ((n_n4434) & (x98x) & (n_n4426) & (!n_n2802) & (!x215x)) + ((n_n4434) & (x98x) & (n_n4426) & (!n_n2802) & (x215x)) + ((n_n4434) & (x98x) & (n_n4426) & (n_n2802) & (!x215x)) + ((n_n4434) & (x98x) & (n_n4426) & (n_n2802) & (x215x)));
	assign x14538x = (((!x194x) & (!n_n3727) & (!n_n3726) & (!x322x) & (x14535x)) + ((!x194x) & (!n_n3727) & (!n_n3726) & (x322x) & (!x14535x)) + ((!x194x) & (!n_n3727) & (!n_n3726) & (x322x) & (x14535x)) + ((!x194x) & (!n_n3727) & (n_n3726) & (!x322x) & (!x14535x)) + ((!x194x) & (!n_n3727) & (n_n3726) & (!x322x) & (x14535x)) + ((!x194x) & (!n_n3727) & (n_n3726) & (x322x) & (!x14535x)) + ((!x194x) & (!n_n3727) & (n_n3726) & (x322x) & (x14535x)) + ((!x194x) & (n_n3727) & (!n_n3726) & (!x322x) & (!x14535x)) + ((!x194x) & (n_n3727) & (!n_n3726) & (!x322x) & (x14535x)) + ((!x194x) & (n_n3727) & (!n_n3726) & (x322x) & (!x14535x)) + ((!x194x) & (n_n3727) & (!n_n3726) & (x322x) & (x14535x)) + ((!x194x) & (n_n3727) & (n_n3726) & (!x322x) & (!x14535x)) + ((!x194x) & (n_n3727) & (n_n3726) & (!x322x) & (x14535x)) + ((!x194x) & (n_n3727) & (n_n3726) & (x322x) & (!x14535x)) + ((!x194x) & (n_n3727) & (n_n3726) & (x322x) & (x14535x)) + ((x194x) & (!n_n3727) & (!n_n3726) & (!x322x) & (!x14535x)) + ((x194x) & (!n_n3727) & (!n_n3726) & (!x322x) & (x14535x)) + ((x194x) & (!n_n3727) & (!n_n3726) & (x322x) & (!x14535x)) + ((x194x) & (!n_n3727) & (!n_n3726) & (x322x) & (x14535x)) + ((x194x) & (!n_n3727) & (n_n3726) & (!x322x) & (!x14535x)) + ((x194x) & (!n_n3727) & (n_n3726) & (!x322x) & (x14535x)) + ((x194x) & (!n_n3727) & (n_n3726) & (x322x) & (!x14535x)) + ((x194x) & (!n_n3727) & (n_n3726) & (x322x) & (x14535x)) + ((x194x) & (n_n3727) & (!n_n3726) & (!x322x) & (!x14535x)) + ((x194x) & (n_n3727) & (!n_n3726) & (!x322x) & (x14535x)) + ((x194x) & (n_n3727) & (!n_n3726) & (x322x) & (!x14535x)) + ((x194x) & (n_n3727) & (!n_n3726) & (x322x) & (x14535x)) + ((x194x) & (n_n3727) & (n_n3726) & (!x322x) & (!x14535x)) + ((x194x) & (n_n3727) & (n_n3726) & (!x322x) & (x14535x)) + ((x194x) & (n_n3727) & (n_n3726) & (x322x) & (!x14535x)) + ((x194x) & (n_n3727) & (n_n3726) & (x322x) & (x14535x)));
	assign n_n522 = (((!i_7_) & (i_8_) & (!i_6_)));
	assign n_n520 = (((!i_7_) & (!i_8_) & (!i_6_)));
	assign n_n464 = (((!i_5_) & (!i_3_) & (!i_4_)));
	assign n_n659 = (((!i_9_) & (!n_n522) & (n_n520) & (n_n464) & (n_n65)) + ((!i_9_) & (n_n522) & (!n_n520) & (n_n464) & (n_n65)) + ((!i_9_) & (n_n522) & (n_n520) & (n_n464) & (n_n65)) + ((i_9_) & (!n_n522) & (n_n520) & (n_n464) & (n_n65)) + ((i_9_) & (n_n522) & (!n_n520) & (n_n464) & (n_n65)) + ((i_9_) & (n_n522) & (n_n520) & (n_n464) & (n_n65)));
	assign n_n3664 = (((!n_n5278) & (!n_n5275) & (!n_n5279) & (!n_n5280) & (!x22186x)) + ((!n_n5278) & (!n_n5275) & (!n_n5279) & (n_n5280) & (!x22186x)) + ((!n_n5278) & (!n_n5275) & (!n_n5279) & (n_n5280) & (x22186x)) + ((!n_n5278) & (!n_n5275) & (n_n5279) & (!n_n5280) & (!x22186x)) + ((!n_n5278) & (!n_n5275) & (n_n5279) & (!n_n5280) & (x22186x)) + ((!n_n5278) & (!n_n5275) & (n_n5279) & (n_n5280) & (!x22186x)) + ((!n_n5278) & (!n_n5275) & (n_n5279) & (n_n5280) & (x22186x)) + ((!n_n5278) & (n_n5275) & (!n_n5279) & (!n_n5280) & (!x22186x)) + ((!n_n5278) & (n_n5275) & (!n_n5279) & (!n_n5280) & (x22186x)) + ((!n_n5278) & (n_n5275) & (!n_n5279) & (n_n5280) & (!x22186x)) + ((!n_n5278) & (n_n5275) & (!n_n5279) & (n_n5280) & (x22186x)) + ((!n_n5278) & (n_n5275) & (n_n5279) & (!n_n5280) & (!x22186x)) + ((!n_n5278) & (n_n5275) & (n_n5279) & (!n_n5280) & (x22186x)) + ((!n_n5278) & (n_n5275) & (n_n5279) & (n_n5280) & (!x22186x)) + ((!n_n5278) & (n_n5275) & (n_n5279) & (n_n5280) & (x22186x)) + ((n_n5278) & (!n_n5275) & (!n_n5279) & (!n_n5280) & (!x22186x)) + ((n_n5278) & (!n_n5275) & (!n_n5279) & (!n_n5280) & (x22186x)) + ((n_n5278) & (!n_n5275) & (!n_n5279) & (n_n5280) & (!x22186x)) + ((n_n5278) & (!n_n5275) & (!n_n5279) & (n_n5280) & (x22186x)) + ((n_n5278) & (!n_n5275) & (n_n5279) & (!n_n5280) & (!x22186x)) + ((n_n5278) & (!n_n5275) & (n_n5279) & (!n_n5280) & (x22186x)) + ((n_n5278) & (!n_n5275) & (n_n5279) & (n_n5280) & (!x22186x)) + ((n_n5278) & (!n_n5275) & (n_n5279) & (n_n5280) & (x22186x)) + ((n_n5278) & (n_n5275) & (!n_n5279) & (!n_n5280) & (!x22186x)) + ((n_n5278) & (n_n5275) & (!n_n5279) & (!n_n5280) & (x22186x)) + ((n_n5278) & (n_n5275) & (!n_n5279) & (n_n5280) & (!x22186x)) + ((n_n5278) & (n_n5275) & (!n_n5279) & (n_n5280) & (x22186x)) + ((n_n5278) & (n_n5275) & (n_n5279) & (!n_n5280) & (!x22186x)) + ((n_n5278) & (n_n5275) & (n_n5279) & (!n_n5280) & (x22186x)) + ((n_n5278) & (n_n5275) & (n_n5279) & (n_n5280) & (!x22186x)) + ((n_n5278) & (n_n5275) & (n_n5279) & (n_n5280) & (x22186x)));
	assign n_n3665 = (((!n_n5267) & (!n_n5262) & (!x409x) & (!x205x) & (x14548x)) + ((!n_n5267) & (!n_n5262) & (!x409x) & (x205x) & (!x14548x)) + ((!n_n5267) & (!n_n5262) & (!x409x) & (x205x) & (x14548x)) + ((!n_n5267) & (!n_n5262) & (x409x) & (!x205x) & (!x14548x)) + ((!n_n5267) & (!n_n5262) & (x409x) & (!x205x) & (x14548x)) + ((!n_n5267) & (!n_n5262) & (x409x) & (x205x) & (!x14548x)) + ((!n_n5267) & (!n_n5262) & (x409x) & (x205x) & (x14548x)) + ((!n_n5267) & (n_n5262) & (!x409x) & (!x205x) & (!x14548x)) + ((!n_n5267) & (n_n5262) & (!x409x) & (!x205x) & (x14548x)) + ((!n_n5267) & (n_n5262) & (!x409x) & (x205x) & (!x14548x)) + ((!n_n5267) & (n_n5262) & (!x409x) & (x205x) & (x14548x)) + ((!n_n5267) & (n_n5262) & (x409x) & (!x205x) & (!x14548x)) + ((!n_n5267) & (n_n5262) & (x409x) & (!x205x) & (x14548x)) + ((!n_n5267) & (n_n5262) & (x409x) & (x205x) & (!x14548x)) + ((!n_n5267) & (n_n5262) & (x409x) & (x205x) & (x14548x)) + ((n_n5267) & (!n_n5262) & (!x409x) & (!x205x) & (!x14548x)) + ((n_n5267) & (!n_n5262) & (!x409x) & (!x205x) & (x14548x)) + ((n_n5267) & (!n_n5262) & (!x409x) & (x205x) & (!x14548x)) + ((n_n5267) & (!n_n5262) & (!x409x) & (x205x) & (x14548x)) + ((n_n5267) & (!n_n5262) & (x409x) & (!x205x) & (!x14548x)) + ((n_n5267) & (!n_n5262) & (x409x) & (!x205x) & (x14548x)) + ((n_n5267) & (!n_n5262) & (x409x) & (x205x) & (!x14548x)) + ((n_n5267) & (!n_n5262) & (x409x) & (x205x) & (x14548x)) + ((n_n5267) & (n_n5262) & (!x409x) & (!x205x) & (!x14548x)) + ((n_n5267) & (n_n5262) & (!x409x) & (!x205x) & (x14548x)) + ((n_n5267) & (n_n5262) & (!x409x) & (x205x) & (!x14548x)) + ((n_n5267) & (n_n5262) & (!x409x) & (x205x) & (x14548x)) + ((n_n5267) & (n_n5262) & (x409x) & (!x205x) & (!x14548x)) + ((n_n5267) & (n_n5262) & (x409x) & (!x205x) & (x14548x)) + ((n_n5267) & (n_n5262) & (x409x) & (x205x) & (!x14548x)) + ((n_n5267) & (n_n5262) & (x409x) & (x205x) & (x14548x)));
	assign x14589x = (((!n_n5289) & (!n_n5285) & (!n_n5282) & (!x14542x) & (!x22107x)) + ((!n_n5289) & (!n_n5285) & (!n_n5282) & (x14542x) & (!x22107x)) + ((!n_n5289) & (!n_n5285) & (!n_n5282) & (x14542x) & (x22107x)) + ((!n_n5289) & (!n_n5285) & (n_n5282) & (!x14542x) & (!x22107x)) + ((!n_n5289) & (!n_n5285) & (n_n5282) & (!x14542x) & (x22107x)) + ((!n_n5289) & (!n_n5285) & (n_n5282) & (x14542x) & (!x22107x)) + ((!n_n5289) & (!n_n5285) & (n_n5282) & (x14542x) & (x22107x)) + ((!n_n5289) & (n_n5285) & (!n_n5282) & (!x14542x) & (!x22107x)) + ((!n_n5289) & (n_n5285) & (!n_n5282) & (!x14542x) & (x22107x)) + ((!n_n5289) & (n_n5285) & (!n_n5282) & (x14542x) & (!x22107x)) + ((!n_n5289) & (n_n5285) & (!n_n5282) & (x14542x) & (x22107x)) + ((!n_n5289) & (n_n5285) & (n_n5282) & (!x14542x) & (!x22107x)) + ((!n_n5289) & (n_n5285) & (n_n5282) & (!x14542x) & (x22107x)) + ((!n_n5289) & (n_n5285) & (n_n5282) & (x14542x) & (!x22107x)) + ((!n_n5289) & (n_n5285) & (n_n5282) & (x14542x) & (x22107x)) + ((n_n5289) & (!n_n5285) & (!n_n5282) & (!x14542x) & (!x22107x)) + ((n_n5289) & (!n_n5285) & (!n_n5282) & (!x14542x) & (x22107x)) + ((n_n5289) & (!n_n5285) & (!n_n5282) & (x14542x) & (!x22107x)) + ((n_n5289) & (!n_n5285) & (!n_n5282) & (x14542x) & (x22107x)) + ((n_n5289) & (!n_n5285) & (n_n5282) & (!x14542x) & (!x22107x)) + ((n_n5289) & (!n_n5285) & (n_n5282) & (!x14542x) & (x22107x)) + ((n_n5289) & (!n_n5285) & (n_n5282) & (x14542x) & (!x22107x)) + ((n_n5289) & (!n_n5285) & (n_n5282) & (x14542x) & (x22107x)) + ((n_n5289) & (n_n5285) & (!n_n5282) & (!x14542x) & (!x22107x)) + ((n_n5289) & (n_n5285) & (!n_n5282) & (!x14542x) & (x22107x)) + ((n_n5289) & (n_n5285) & (!n_n5282) & (x14542x) & (!x22107x)) + ((n_n5289) & (n_n5285) & (!n_n5282) & (x14542x) & (x22107x)) + ((n_n5289) & (n_n5285) & (n_n5282) & (!x14542x) & (!x22107x)) + ((n_n5289) & (n_n5285) & (n_n5282) & (!x14542x) & (x22107x)) + ((n_n5289) & (n_n5285) & (n_n5282) & (x14542x) & (!x22107x)) + ((n_n5289) & (n_n5285) & (n_n5282) & (x14542x) & (x22107x)));
	assign x14591x = (((!n_n3664) & (!n_n3665) & (x14589x)) + ((!n_n3664) & (n_n3665) & (!x14589x)) + ((!n_n3664) & (n_n3665) & (x14589x)) + ((n_n3664) & (!n_n3665) & (!x14589x)) + ((n_n3664) & (!n_n3665) & (x14589x)) + ((n_n3664) & (n_n3665) & (!x14589x)) + ((n_n3664) & (n_n3665) & (x14589x)));
	assign n_n3661 = (((!n_n5312) & (!n_n5313) & (!x325x) & (!n_n5315) & (!x22106x)) + ((!n_n5312) & (!n_n5313) & (!x325x) & (n_n5315) & (!x22106x)) + ((!n_n5312) & (!n_n5313) & (!x325x) & (n_n5315) & (x22106x)) + ((!n_n5312) & (!n_n5313) & (x325x) & (!n_n5315) & (!x22106x)) + ((!n_n5312) & (!n_n5313) & (x325x) & (!n_n5315) & (x22106x)) + ((!n_n5312) & (!n_n5313) & (x325x) & (n_n5315) & (!x22106x)) + ((!n_n5312) & (!n_n5313) & (x325x) & (n_n5315) & (x22106x)) + ((!n_n5312) & (n_n5313) & (!x325x) & (!n_n5315) & (!x22106x)) + ((!n_n5312) & (n_n5313) & (!x325x) & (!n_n5315) & (x22106x)) + ((!n_n5312) & (n_n5313) & (!x325x) & (n_n5315) & (!x22106x)) + ((!n_n5312) & (n_n5313) & (!x325x) & (n_n5315) & (x22106x)) + ((!n_n5312) & (n_n5313) & (x325x) & (!n_n5315) & (!x22106x)) + ((!n_n5312) & (n_n5313) & (x325x) & (!n_n5315) & (x22106x)) + ((!n_n5312) & (n_n5313) & (x325x) & (n_n5315) & (!x22106x)) + ((!n_n5312) & (n_n5313) & (x325x) & (n_n5315) & (x22106x)) + ((n_n5312) & (!n_n5313) & (!x325x) & (!n_n5315) & (!x22106x)) + ((n_n5312) & (!n_n5313) & (!x325x) & (!n_n5315) & (x22106x)) + ((n_n5312) & (!n_n5313) & (!x325x) & (n_n5315) & (!x22106x)) + ((n_n5312) & (!n_n5313) & (!x325x) & (n_n5315) & (x22106x)) + ((n_n5312) & (!n_n5313) & (x325x) & (!n_n5315) & (!x22106x)) + ((n_n5312) & (!n_n5313) & (x325x) & (!n_n5315) & (x22106x)) + ((n_n5312) & (!n_n5313) & (x325x) & (n_n5315) & (!x22106x)) + ((n_n5312) & (!n_n5313) & (x325x) & (n_n5315) & (x22106x)) + ((n_n5312) & (n_n5313) & (!x325x) & (!n_n5315) & (!x22106x)) + ((n_n5312) & (n_n5313) & (!x325x) & (!n_n5315) & (x22106x)) + ((n_n5312) & (n_n5313) & (!x325x) & (n_n5315) & (!x22106x)) + ((n_n5312) & (n_n5313) & (!x325x) & (n_n5315) & (x22106x)) + ((n_n5312) & (n_n5313) & (x325x) & (!n_n5315) & (!x22106x)) + ((n_n5312) & (n_n5313) & (x325x) & (!n_n5315) & (x22106x)) + ((n_n5312) & (n_n5313) & (x325x) & (n_n5315) & (!x22106x)) + ((n_n5312) & (n_n5313) & (x325x) & (n_n5315) & (x22106x)));
	assign n_n3660 = (((!n_n5318) & (!n_n5326) & (!n_n5329) & (!n_n5327) & (x14561x)) + ((!n_n5318) & (!n_n5326) & (!n_n5329) & (n_n5327) & (!x14561x)) + ((!n_n5318) & (!n_n5326) & (!n_n5329) & (n_n5327) & (x14561x)) + ((!n_n5318) & (!n_n5326) & (n_n5329) & (!n_n5327) & (!x14561x)) + ((!n_n5318) & (!n_n5326) & (n_n5329) & (!n_n5327) & (x14561x)) + ((!n_n5318) & (!n_n5326) & (n_n5329) & (n_n5327) & (!x14561x)) + ((!n_n5318) & (!n_n5326) & (n_n5329) & (n_n5327) & (x14561x)) + ((!n_n5318) & (n_n5326) & (!n_n5329) & (!n_n5327) & (!x14561x)) + ((!n_n5318) & (n_n5326) & (!n_n5329) & (!n_n5327) & (x14561x)) + ((!n_n5318) & (n_n5326) & (!n_n5329) & (n_n5327) & (!x14561x)) + ((!n_n5318) & (n_n5326) & (!n_n5329) & (n_n5327) & (x14561x)) + ((!n_n5318) & (n_n5326) & (n_n5329) & (!n_n5327) & (!x14561x)) + ((!n_n5318) & (n_n5326) & (n_n5329) & (!n_n5327) & (x14561x)) + ((!n_n5318) & (n_n5326) & (n_n5329) & (n_n5327) & (!x14561x)) + ((!n_n5318) & (n_n5326) & (n_n5329) & (n_n5327) & (x14561x)) + ((n_n5318) & (!n_n5326) & (!n_n5329) & (!n_n5327) & (!x14561x)) + ((n_n5318) & (!n_n5326) & (!n_n5329) & (!n_n5327) & (x14561x)) + ((n_n5318) & (!n_n5326) & (!n_n5329) & (n_n5327) & (!x14561x)) + ((n_n5318) & (!n_n5326) & (!n_n5329) & (n_n5327) & (x14561x)) + ((n_n5318) & (!n_n5326) & (n_n5329) & (!n_n5327) & (!x14561x)) + ((n_n5318) & (!n_n5326) & (n_n5329) & (!n_n5327) & (x14561x)) + ((n_n5318) & (!n_n5326) & (n_n5329) & (n_n5327) & (!x14561x)) + ((n_n5318) & (!n_n5326) & (n_n5329) & (n_n5327) & (x14561x)) + ((n_n5318) & (n_n5326) & (!n_n5329) & (!n_n5327) & (!x14561x)) + ((n_n5318) & (n_n5326) & (!n_n5329) & (!n_n5327) & (x14561x)) + ((n_n5318) & (n_n5326) & (!n_n5329) & (n_n5327) & (!x14561x)) + ((n_n5318) & (n_n5326) & (!n_n5329) & (n_n5327) & (x14561x)) + ((n_n5318) & (n_n5326) & (n_n5329) & (!n_n5327) & (!x14561x)) + ((n_n5318) & (n_n5326) & (n_n5329) & (!n_n5327) & (x14561x)) + ((n_n5318) & (n_n5326) & (n_n5329) & (n_n5327) & (!x14561x)) + ((n_n5318) & (n_n5326) & (n_n5329) & (n_n5327) & (x14561x)));
	assign x14566x = (((!n_n5292) & (!x197x) & (!x200x) & (!x60x) & (x14562x)) + ((!n_n5292) & (!x197x) & (!x200x) & (x60x) & (!x14562x)) + ((!n_n5292) & (!x197x) & (!x200x) & (x60x) & (x14562x)) + ((!n_n5292) & (!x197x) & (x200x) & (!x60x) & (!x14562x)) + ((!n_n5292) & (!x197x) & (x200x) & (!x60x) & (x14562x)) + ((!n_n5292) & (!x197x) & (x200x) & (x60x) & (!x14562x)) + ((!n_n5292) & (!x197x) & (x200x) & (x60x) & (x14562x)) + ((!n_n5292) & (x197x) & (!x200x) & (!x60x) & (!x14562x)) + ((!n_n5292) & (x197x) & (!x200x) & (!x60x) & (x14562x)) + ((!n_n5292) & (x197x) & (!x200x) & (x60x) & (!x14562x)) + ((!n_n5292) & (x197x) & (!x200x) & (x60x) & (x14562x)) + ((!n_n5292) & (x197x) & (x200x) & (!x60x) & (!x14562x)) + ((!n_n5292) & (x197x) & (x200x) & (!x60x) & (x14562x)) + ((!n_n5292) & (x197x) & (x200x) & (x60x) & (!x14562x)) + ((!n_n5292) & (x197x) & (x200x) & (x60x) & (x14562x)) + ((n_n5292) & (!x197x) & (!x200x) & (!x60x) & (!x14562x)) + ((n_n5292) & (!x197x) & (!x200x) & (!x60x) & (x14562x)) + ((n_n5292) & (!x197x) & (!x200x) & (x60x) & (!x14562x)) + ((n_n5292) & (!x197x) & (!x200x) & (x60x) & (x14562x)) + ((n_n5292) & (!x197x) & (x200x) & (!x60x) & (!x14562x)) + ((n_n5292) & (!x197x) & (x200x) & (!x60x) & (x14562x)) + ((n_n5292) & (!x197x) & (x200x) & (x60x) & (!x14562x)) + ((n_n5292) & (!x197x) & (x200x) & (x60x) & (x14562x)) + ((n_n5292) & (x197x) & (!x200x) & (!x60x) & (!x14562x)) + ((n_n5292) & (x197x) & (!x200x) & (!x60x) & (x14562x)) + ((n_n5292) & (x197x) & (!x200x) & (x60x) & (!x14562x)) + ((n_n5292) & (x197x) & (!x200x) & (x60x) & (x14562x)) + ((n_n5292) & (x197x) & (x200x) & (!x60x) & (!x14562x)) + ((n_n5292) & (x197x) & (x200x) & (!x60x) & (x14562x)) + ((n_n5292) & (x197x) & (x200x) & (x60x) & (!x14562x)) + ((n_n5292) & (x197x) & (x200x) & (x60x) & (x14562x)));
	assign n_n3634 = (((!x14572x) & (!x14573x) & (!x14579x) & (!x14580x) & (x14581x)) + ((!x14572x) & (!x14573x) & (!x14579x) & (x14580x) & (!x14581x)) + ((!x14572x) & (!x14573x) & (!x14579x) & (x14580x) & (x14581x)) + ((!x14572x) & (!x14573x) & (x14579x) & (!x14580x) & (!x14581x)) + ((!x14572x) & (!x14573x) & (x14579x) & (!x14580x) & (x14581x)) + ((!x14572x) & (!x14573x) & (x14579x) & (x14580x) & (!x14581x)) + ((!x14572x) & (!x14573x) & (x14579x) & (x14580x) & (x14581x)) + ((!x14572x) & (x14573x) & (!x14579x) & (!x14580x) & (!x14581x)) + ((!x14572x) & (x14573x) & (!x14579x) & (!x14580x) & (x14581x)) + ((!x14572x) & (x14573x) & (!x14579x) & (x14580x) & (!x14581x)) + ((!x14572x) & (x14573x) & (!x14579x) & (x14580x) & (x14581x)) + ((!x14572x) & (x14573x) & (x14579x) & (!x14580x) & (!x14581x)) + ((!x14572x) & (x14573x) & (x14579x) & (!x14580x) & (x14581x)) + ((!x14572x) & (x14573x) & (x14579x) & (x14580x) & (!x14581x)) + ((!x14572x) & (x14573x) & (x14579x) & (x14580x) & (x14581x)) + ((x14572x) & (!x14573x) & (!x14579x) & (!x14580x) & (!x14581x)) + ((x14572x) & (!x14573x) & (!x14579x) & (!x14580x) & (x14581x)) + ((x14572x) & (!x14573x) & (!x14579x) & (x14580x) & (!x14581x)) + ((x14572x) & (!x14573x) & (!x14579x) & (x14580x) & (x14581x)) + ((x14572x) & (!x14573x) & (x14579x) & (!x14580x) & (!x14581x)) + ((x14572x) & (!x14573x) & (x14579x) & (!x14580x) & (x14581x)) + ((x14572x) & (!x14573x) & (x14579x) & (x14580x) & (!x14581x)) + ((x14572x) & (!x14573x) & (x14579x) & (x14580x) & (x14581x)) + ((x14572x) & (x14573x) & (!x14579x) & (!x14580x) & (!x14581x)) + ((x14572x) & (x14573x) & (!x14579x) & (!x14580x) & (x14581x)) + ((x14572x) & (x14573x) & (!x14579x) & (x14580x) & (!x14581x)) + ((x14572x) & (x14573x) & (!x14579x) & (x14580x) & (x14581x)) + ((x14572x) & (x14573x) & (x14579x) & (!x14580x) & (!x14581x)) + ((x14572x) & (x14573x) & (x14579x) & (!x14580x) & (x14581x)) + ((x14572x) & (x14573x) & (x14579x) & (x14580x) & (!x14581x)) + ((x14572x) & (x14573x) & (x14579x) & (x14580x) & (x14581x)));
	assign n_n3674 = (((!x76x) & (!x126x) & (!n_n5144) & (!n_n5143) & (n_n777)) + ((!x76x) & (!x126x) & (!n_n5144) & (n_n5143) & (!n_n777)) + ((!x76x) & (!x126x) & (!n_n5144) & (n_n5143) & (n_n777)) + ((!x76x) & (!x126x) & (n_n5144) & (!n_n5143) & (!n_n777)) + ((!x76x) & (!x126x) & (n_n5144) & (!n_n5143) & (n_n777)) + ((!x76x) & (!x126x) & (n_n5144) & (n_n5143) & (!n_n777)) + ((!x76x) & (!x126x) & (n_n5144) & (n_n5143) & (n_n777)) + ((!x76x) & (x126x) & (!n_n5144) & (!n_n5143) & (!n_n777)) + ((!x76x) & (x126x) & (!n_n5144) & (!n_n5143) & (n_n777)) + ((!x76x) & (x126x) & (!n_n5144) & (n_n5143) & (!n_n777)) + ((!x76x) & (x126x) & (!n_n5144) & (n_n5143) & (n_n777)) + ((!x76x) & (x126x) & (n_n5144) & (!n_n5143) & (!n_n777)) + ((!x76x) & (x126x) & (n_n5144) & (!n_n5143) & (n_n777)) + ((!x76x) & (x126x) & (n_n5144) & (n_n5143) & (!n_n777)) + ((!x76x) & (x126x) & (n_n5144) & (n_n5143) & (n_n777)) + ((x76x) & (!x126x) & (!n_n5144) & (!n_n5143) & (!n_n777)) + ((x76x) & (!x126x) & (!n_n5144) & (!n_n5143) & (n_n777)) + ((x76x) & (!x126x) & (!n_n5144) & (n_n5143) & (!n_n777)) + ((x76x) & (!x126x) & (!n_n5144) & (n_n5143) & (n_n777)) + ((x76x) & (!x126x) & (n_n5144) & (!n_n5143) & (!n_n777)) + ((x76x) & (!x126x) & (n_n5144) & (!n_n5143) & (n_n777)) + ((x76x) & (!x126x) & (n_n5144) & (n_n5143) & (!n_n777)) + ((x76x) & (!x126x) & (n_n5144) & (n_n5143) & (n_n777)) + ((x76x) & (x126x) & (!n_n5144) & (!n_n5143) & (!n_n777)) + ((x76x) & (x126x) & (!n_n5144) & (!n_n5143) & (n_n777)) + ((x76x) & (x126x) & (!n_n5144) & (n_n5143) & (!n_n777)) + ((x76x) & (x126x) & (!n_n5144) & (n_n5143) & (n_n777)) + ((x76x) & (x126x) & (n_n5144) & (!n_n5143) & (!n_n777)) + ((x76x) & (x126x) & (n_n5144) & (!n_n5143) & (n_n777)) + ((x76x) & (x126x) & (n_n5144) & (n_n5143) & (!n_n777)) + ((x76x) & (x126x) & (n_n5144) & (n_n5143) & (n_n777)));
	assign n_n3673 = (((!n_n5155) & (!n_n5163) & (!n_n5154) & (!x195x) & (x14598x)) + ((!n_n5155) & (!n_n5163) & (!n_n5154) & (x195x) & (!x14598x)) + ((!n_n5155) & (!n_n5163) & (!n_n5154) & (x195x) & (x14598x)) + ((!n_n5155) & (!n_n5163) & (n_n5154) & (!x195x) & (!x14598x)) + ((!n_n5155) & (!n_n5163) & (n_n5154) & (!x195x) & (x14598x)) + ((!n_n5155) & (!n_n5163) & (n_n5154) & (x195x) & (!x14598x)) + ((!n_n5155) & (!n_n5163) & (n_n5154) & (x195x) & (x14598x)) + ((!n_n5155) & (n_n5163) & (!n_n5154) & (!x195x) & (!x14598x)) + ((!n_n5155) & (n_n5163) & (!n_n5154) & (!x195x) & (x14598x)) + ((!n_n5155) & (n_n5163) & (!n_n5154) & (x195x) & (!x14598x)) + ((!n_n5155) & (n_n5163) & (!n_n5154) & (x195x) & (x14598x)) + ((!n_n5155) & (n_n5163) & (n_n5154) & (!x195x) & (!x14598x)) + ((!n_n5155) & (n_n5163) & (n_n5154) & (!x195x) & (x14598x)) + ((!n_n5155) & (n_n5163) & (n_n5154) & (x195x) & (!x14598x)) + ((!n_n5155) & (n_n5163) & (n_n5154) & (x195x) & (x14598x)) + ((n_n5155) & (!n_n5163) & (!n_n5154) & (!x195x) & (!x14598x)) + ((n_n5155) & (!n_n5163) & (!n_n5154) & (!x195x) & (x14598x)) + ((n_n5155) & (!n_n5163) & (!n_n5154) & (x195x) & (!x14598x)) + ((n_n5155) & (!n_n5163) & (!n_n5154) & (x195x) & (x14598x)) + ((n_n5155) & (!n_n5163) & (n_n5154) & (!x195x) & (!x14598x)) + ((n_n5155) & (!n_n5163) & (n_n5154) & (!x195x) & (x14598x)) + ((n_n5155) & (!n_n5163) & (n_n5154) & (x195x) & (!x14598x)) + ((n_n5155) & (!n_n5163) & (n_n5154) & (x195x) & (x14598x)) + ((n_n5155) & (n_n5163) & (!n_n5154) & (!x195x) & (!x14598x)) + ((n_n5155) & (n_n5163) & (!n_n5154) & (!x195x) & (x14598x)) + ((n_n5155) & (n_n5163) & (!n_n5154) & (x195x) & (!x14598x)) + ((n_n5155) & (n_n5163) & (!n_n5154) & (x195x) & (x14598x)) + ((n_n5155) & (n_n5163) & (n_n5154) & (!x195x) & (!x14598x)) + ((n_n5155) & (n_n5163) & (n_n5154) & (!x195x) & (x14598x)) + ((n_n5155) & (n_n5163) & (n_n5154) & (x195x) & (!x14598x)) + ((n_n5155) & (n_n5163) & (n_n5154) & (x195x) & (x14598x)));
	assign x14636x = (((!n_n5171) & (!n_n5173) & (!x33x) & (x14635x)) + ((!n_n5171) & (!n_n5173) & (x33x) & (!x14635x)) + ((!n_n5171) & (!n_n5173) & (x33x) & (x14635x)) + ((!n_n5171) & (n_n5173) & (!x33x) & (!x14635x)) + ((!n_n5171) & (n_n5173) & (!x33x) & (x14635x)) + ((!n_n5171) & (n_n5173) & (x33x) & (!x14635x)) + ((!n_n5171) & (n_n5173) & (x33x) & (x14635x)) + ((n_n5171) & (!n_n5173) & (!x33x) & (!x14635x)) + ((n_n5171) & (!n_n5173) & (!x33x) & (x14635x)) + ((n_n5171) & (!n_n5173) & (x33x) & (!x14635x)) + ((n_n5171) & (!n_n5173) & (x33x) & (x14635x)) + ((n_n5171) & (n_n5173) & (!x33x) & (!x14635x)) + ((n_n5171) & (n_n5173) & (!x33x) & (x14635x)) + ((n_n5171) & (n_n5173) & (x33x) & (!x14635x)) + ((n_n5171) & (n_n5173) & (x33x) & (x14635x)));
	assign x14638x = (((!n_n3674) & (!n_n3673) & (x14636x)) + ((!n_n3674) & (n_n3673) & (!x14636x)) + ((!n_n3674) & (n_n3673) & (x14636x)) + ((n_n3674) & (!n_n3673) & (!x14636x)) + ((n_n3674) & (!n_n3673) & (x14636x)) + ((n_n3674) & (n_n3673) & (!x14636x)) + ((n_n3674) & (n_n3673) & (x14636x)));
	assign x14613x = (((!n_n5113) & (!n_n5114) & (!n_n3412) & (!n_n3771) & (n_n3772)) + ((!n_n5113) & (!n_n5114) & (!n_n3412) & (n_n3771) & (!n_n3772)) + ((!n_n5113) & (!n_n5114) & (!n_n3412) & (n_n3771) & (n_n3772)) + ((!n_n5113) & (!n_n5114) & (n_n3412) & (!n_n3771) & (!n_n3772)) + ((!n_n5113) & (!n_n5114) & (n_n3412) & (!n_n3771) & (n_n3772)) + ((!n_n5113) & (!n_n5114) & (n_n3412) & (n_n3771) & (!n_n3772)) + ((!n_n5113) & (!n_n5114) & (n_n3412) & (n_n3771) & (n_n3772)) + ((!n_n5113) & (n_n5114) & (!n_n3412) & (!n_n3771) & (!n_n3772)) + ((!n_n5113) & (n_n5114) & (!n_n3412) & (!n_n3771) & (n_n3772)) + ((!n_n5113) & (n_n5114) & (!n_n3412) & (n_n3771) & (!n_n3772)) + ((!n_n5113) & (n_n5114) & (!n_n3412) & (n_n3771) & (n_n3772)) + ((!n_n5113) & (n_n5114) & (n_n3412) & (!n_n3771) & (!n_n3772)) + ((!n_n5113) & (n_n5114) & (n_n3412) & (!n_n3771) & (n_n3772)) + ((!n_n5113) & (n_n5114) & (n_n3412) & (n_n3771) & (!n_n3772)) + ((!n_n5113) & (n_n5114) & (n_n3412) & (n_n3771) & (n_n3772)) + ((n_n5113) & (!n_n5114) & (!n_n3412) & (!n_n3771) & (!n_n3772)) + ((n_n5113) & (!n_n5114) & (!n_n3412) & (!n_n3771) & (n_n3772)) + ((n_n5113) & (!n_n5114) & (!n_n3412) & (n_n3771) & (!n_n3772)) + ((n_n5113) & (!n_n5114) & (!n_n3412) & (n_n3771) & (n_n3772)) + ((n_n5113) & (!n_n5114) & (n_n3412) & (!n_n3771) & (!n_n3772)) + ((n_n5113) & (!n_n5114) & (n_n3412) & (!n_n3771) & (n_n3772)) + ((n_n5113) & (!n_n5114) & (n_n3412) & (n_n3771) & (!n_n3772)) + ((n_n5113) & (!n_n5114) & (n_n3412) & (n_n3771) & (n_n3772)) + ((n_n5113) & (n_n5114) & (!n_n3412) & (!n_n3771) & (!n_n3772)) + ((n_n5113) & (n_n5114) & (!n_n3412) & (!n_n3771) & (n_n3772)) + ((n_n5113) & (n_n5114) & (!n_n3412) & (n_n3771) & (!n_n3772)) + ((n_n5113) & (n_n5114) & (!n_n3412) & (n_n3771) & (n_n3772)) + ((n_n5113) & (n_n5114) & (n_n3412) & (!n_n3771) & (!n_n3772)) + ((n_n5113) & (n_n5114) & (n_n3412) & (!n_n3771) & (n_n3772)) + ((n_n5113) & (n_n5114) & (n_n3412) & (n_n3771) & (!n_n3772)) + ((n_n5113) & (n_n5114) & (n_n3412) & (n_n3771) & (n_n3772)));
	assign n_n3635 = (((!n_n5203) & (!x188x) & (!n_n3670) & (!x14629x) & (x14625x)) + ((!n_n5203) & (!x188x) & (!n_n3670) & (x14629x) & (!x14625x)) + ((!n_n5203) & (!x188x) & (!n_n3670) & (x14629x) & (x14625x)) + ((!n_n5203) & (!x188x) & (n_n3670) & (!x14629x) & (!x14625x)) + ((!n_n5203) & (!x188x) & (n_n3670) & (!x14629x) & (x14625x)) + ((!n_n5203) & (!x188x) & (n_n3670) & (x14629x) & (!x14625x)) + ((!n_n5203) & (!x188x) & (n_n3670) & (x14629x) & (x14625x)) + ((!n_n5203) & (x188x) & (!n_n3670) & (!x14629x) & (!x14625x)) + ((!n_n5203) & (x188x) & (!n_n3670) & (!x14629x) & (x14625x)) + ((!n_n5203) & (x188x) & (!n_n3670) & (x14629x) & (!x14625x)) + ((!n_n5203) & (x188x) & (!n_n3670) & (x14629x) & (x14625x)) + ((!n_n5203) & (x188x) & (n_n3670) & (!x14629x) & (!x14625x)) + ((!n_n5203) & (x188x) & (n_n3670) & (!x14629x) & (x14625x)) + ((!n_n5203) & (x188x) & (n_n3670) & (x14629x) & (!x14625x)) + ((!n_n5203) & (x188x) & (n_n3670) & (x14629x) & (x14625x)) + ((n_n5203) & (!x188x) & (!n_n3670) & (!x14629x) & (!x14625x)) + ((n_n5203) & (!x188x) & (!n_n3670) & (!x14629x) & (x14625x)) + ((n_n5203) & (!x188x) & (!n_n3670) & (x14629x) & (!x14625x)) + ((n_n5203) & (!x188x) & (!n_n3670) & (x14629x) & (x14625x)) + ((n_n5203) & (!x188x) & (n_n3670) & (!x14629x) & (!x14625x)) + ((n_n5203) & (!x188x) & (n_n3670) & (!x14629x) & (x14625x)) + ((n_n5203) & (!x188x) & (n_n3670) & (x14629x) & (!x14625x)) + ((n_n5203) & (!x188x) & (n_n3670) & (x14629x) & (x14625x)) + ((n_n5203) & (x188x) & (!n_n3670) & (!x14629x) & (!x14625x)) + ((n_n5203) & (x188x) & (!n_n3670) & (!x14629x) & (x14625x)) + ((n_n5203) & (x188x) & (!n_n3670) & (x14629x) & (!x14625x)) + ((n_n5203) & (x188x) & (!n_n3670) & (x14629x) & (x14625x)) + ((n_n5203) & (x188x) & (n_n3670) & (!x14629x) & (!x14625x)) + ((n_n5203) & (x188x) & (n_n3670) & (!x14629x) & (x14625x)) + ((n_n5203) & (x188x) & (n_n3670) & (x14629x) & (!x14625x)) + ((n_n5203) & (x188x) & (n_n3670) & (x14629x) & (x14625x)));
	assign n_n3676 = (((!n_n5121) & (!n_n5119) & (!x14604x) & (!x22105x)) + ((!n_n5121) & (!n_n5119) & (x14604x) & (!x22105x)) + ((!n_n5121) & (!n_n5119) & (x14604x) & (x22105x)) + ((!n_n5121) & (n_n5119) & (!x14604x) & (!x22105x)) + ((!n_n5121) & (n_n5119) & (!x14604x) & (x22105x)) + ((!n_n5121) & (n_n5119) & (x14604x) & (!x22105x)) + ((!n_n5121) & (n_n5119) & (x14604x) & (x22105x)) + ((n_n5121) & (!n_n5119) & (!x14604x) & (!x22105x)) + ((n_n5121) & (!n_n5119) & (!x14604x) & (x22105x)) + ((n_n5121) & (!n_n5119) & (x14604x) & (!x22105x)) + ((n_n5121) & (!n_n5119) & (x14604x) & (x22105x)) + ((n_n5121) & (n_n5119) & (!x14604x) & (!x22105x)) + ((n_n5121) & (n_n5119) & (!x14604x) & (x22105x)) + ((n_n5121) & (n_n5119) & (x14604x) & (!x22105x)) + ((n_n5121) & (n_n5119) & (x14604x) & (x22105x)));
	assign x14612x = (((!n_n5111) & (!n_n5112) & (!n_n5107) & (!n_n5108) & (n_n3051)) + ((!n_n5111) & (!n_n5112) & (!n_n5107) & (n_n5108) & (!n_n3051)) + ((!n_n5111) & (!n_n5112) & (!n_n5107) & (n_n5108) & (n_n3051)) + ((!n_n5111) & (!n_n5112) & (n_n5107) & (!n_n5108) & (!n_n3051)) + ((!n_n5111) & (!n_n5112) & (n_n5107) & (!n_n5108) & (n_n3051)) + ((!n_n5111) & (!n_n5112) & (n_n5107) & (n_n5108) & (!n_n3051)) + ((!n_n5111) & (!n_n5112) & (n_n5107) & (n_n5108) & (n_n3051)) + ((!n_n5111) & (n_n5112) & (!n_n5107) & (!n_n5108) & (!n_n3051)) + ((!n_n5111) & (n_n5112) & (!n_n5107) & (!n_n5108) & (n_n3051)) + ((!n_n5111) & (n_n5112) & (!n_n5107) & (n_n5108) & (!n_n3051)) + ((!n_n5111) & (n_n5112) & (!n_n5107) & (n_n5108) & (n_n3051)) + ((!n_n5111) & (n_n5112) & (n_n5107) & (!n_n5108) & (!n_n3051)) + ((!n_n5111) & (n_n5112) & (n_n5107) & (!n_n5108) & (n_n3051)) + ((!n_n5111) & (n_n5112) & (n_n5107) & (n_n5108) & (!n_n3051)) + ((!n_n5111) & (n_n5112) & (n_n5107) & (n_n5108) & (n_n3051)) + ((n_n5111) & (!n_n5112) & (!n_n5107) & (!n_n5108) & (!n_n3051)) + ((n_n5111) & (!n_n5112) & (!n_n5107) & (!n_n5108) & (n_n3051)) + ((n_n5111) & (!n_n5112) & (!n_n5107) & (n_n5108) & (!n_n3051)) + ((n_n5111) & (!n_n5112) & (!n_n5107) & (n_n5108) & (n_n3051)) + ((n_n5111) & (!n_n5112) & (n_n5107) & (!n_n5108) & (!n_n3051)) + ((n_n5111) & (!n_n5112) & (n_n5107) & (!n_n5108) & (n_n3051)) + ((n_n5111) & (!n_n5112) & (n_n5107) & (n_n5108) & (!n_n3051)) + ((n_n5111) & (!n_n5112) & (n_n5107) & (n_n5108) & (n_n3051)) + ((n_n5111) & (n_n5112) & (!n_n5107) & (!n_n5108) & (!n_n3051)) + ((n_n5111) & (n_n5112) & (!n_n5107) & (!n_n5108) & (n_n3051)) + ((n_n5111) & (n_n5112) & (!n_n5107) & (n_n5108) & (!n_n3051)) + ((n_n5111) & (n_n5112) & (!n_n5107) & (n_n5108) & (n_n3051)) + ((n_n5111) & (n_n5112) & (n_n5107) & (!n_n5108) & (!n_n3051)) + ((n_n5111) & (n_n5112) & (n_n5107) & (!n_n5108) & (n_n3051)) + ((n_n5111) & (n_n5112) & (n_n5107) & (n_n5108) & (!n_n3051)) + ((n_n5111) & (n_n5112) & (n_n5107) & (n_n5108) & (n_n3051)));
	assign n_n3638 = (((!x14644x) & (!x14645x) & (!x14648x) & (!x14649x) & (x14654x)) + ((!x14644x) & (!x14645x) & (!x14648x) & (x14649x) & (!x14654x)) + ((!x14644x) & (!x14645x) & (!x14648x) & (x14649x) & (x14654x)) + ((!x14644x) & (!x14645x) & (x14648x) & (!x14649x) & (!x14654x)) + ((!x14644x) & (!x14645x) & (x14648x) & (!x14649x) & (x14654x)) + ((!x14644x) & (!x14645x) & (x14648x) & (x14649x) & (!x14654x)) + ((!x14644x) & (!x14645x) & (x14648x) & (x14649x) & (x14654x)) + ((!x14644x) & (x14645x) & (!x14648x) & (!x14649x) & (!x14654x)) + ((!x14644x) & (x14645x) & (!x14648x) & (!x14649x) & (x14654x)) + ((!x14644x) & (x14645x) & (!x14648x) & (x14649x) & (!x14654x)) + ((!x14644x) & (x14645x) & (!x14648x) & (x14649x) & (x14654x)) + ((!x14644x) & (x14645x) & (x14648x) & (!x14649x) & (!x14654x)) + ((!x14644x) & (x14645x) & (x14648x) & (!x14649x) & (x14654x)) + ((!x14644x) & (x14645x) & (x14648x) & (x14649x) & (!x14654x)) + ((!x14644x) & (x14645x) & (x14648x) & (x14649x) & (x14654x)) + ((x14644x) & (!x14645x) & (!x14648x) & (!x14649x) & (!x14654x)) + ((x14644x) & (!x14645x) & (!x14648x) & (!x14649x) & (x14654x)) + ((x14644x) & (!x14645x) & (!x14648x) & (x14649x) & (!x14654x)) + ((x14644x) & (!x14645x) & (!x14648x) & (x14649x) & (x14654x)) + ((x14644x) & (!x14645x) & (x14648x) & (!x14649x) & (!x14654x)) + ((x14644x) & (!x14645x) & (x14648x) & (!x14649x) & (x14654x)) + ((x14644x) & (!x14645x) & (x14648x) & (x14649x) & (!x14654x)) + ((x14644x) & (!x14645x) & (x14648x) & (x14649x) & (x14654x)) + ((x14644x) & (x14645x) & (!x14648x) & (!x14649x) & (!x14654x)) + ((x14644x) & (x14645x) & (!x14648x) & (!x14649x) & (x14654x)) + ((x14644x) & (x14645x) & (!x14648x) & (x14649x) & (!x14654x)) + ((x14644x) & (x14645x) & (!x14648x) & (x14649x) & (x14654x)) + ((x14644x) & (x14645x) & (x14648x) & (!x14649x) & (!x14654x)) + ((x14644x) & (x14645x) & (x14648x) & (!x14649x) & (x14654x)) + ((x14644x) & (x14645x) & (x14648x) & (x14649x) & (!x14654x)) + ((x14644x) & (x14645x) & (x14648x) & (x14649x) & (x14654x)));
	assign n_n3639 = (((!x14659x) & (!x14660x) & (!x467x) & (!x14665x) & (x14666x)) + ((!x14659x) & (!x14660x) & (!x467x) & (x14665x) & (!x14666x)) + ((!x14659x) & (!x14660x) & (!x467x) & (x14665x) & (x14666x)) + ((!x14659x) & (!x14660x) & (x467x) & (!x14665x) & (!x14666x)) + ((!x14659x) & (!x14660x) & (x467x) & (!x14665x) & (x14666x)) + ((!x14659x) & (!x14660x) & (x467x) & (x14665x) & (!x14666x)) + ((!x14659x) & (!x14660x) & (x467x) & (x14665x) & (x14666x)) + ((!x14659x) & (x14660x) & (!x467x) & (!x14665x) & (!x14666x)) + ((!x14659x) & (x14660x) & (!x467x) & (!x14665x) & (x14666x)) + ((!x14659x) & (x14660x) & (!x467x) & (x14665x) & (!x14666x)) + ((!x14659x) & (x14660x) & (!x467x) & (x14665x) & (x14666x)) + ((!x14659x) & (x14660x) & (x467x) & (!x14665x) & (!x14666x)) + ((!x14659x) & (x14660x) & (x467x) & (!x14665x) & (x14666x)) + ((!x14659x) & (x14660x) & (x467x) & (x14665x) & (!x14666x)) + ((!x14659x) & (x14660x) & (x467x) & (x14665x) & (x14666x)) + ((x14659x) & (!x14660x) & (!x467x) & (!x14665x) & (!x14666x)) + ((x14659x) & (!x14660x) & (!x467x) & (!x14665x) & (x14666x)) + ((x14659x) & (!x14660x) & (!x467x) & (x14665x) & (!x14666x)) + ((x14659x) & (!x14660x) & (!x467x) & (x14665x) & (x14666x)) + ((x14659x) & (!x14660x) & (x467x) & (!x14665x) & (!x14666x)) + ((x14659x) & (!x14660x) & (x467x) & (!x14665x) & (x14666x)) + ((x14659x) & (!x14660x) & (x467x) & (x14665x) & (!x14666x)) + ((x14659x) & (!x14660x) & (x467x) & (x14665x) & (x14666x)) + ((x14659x) & (x14660x) & (!x467x) & (!x14665x) & (!x14666x)) + ((x14659x) & (x14660x) & (!x467x) & (!x14665x) & (x14666x)) + ((x14659x) & (x14660x) & (!x467x) & (x14665x) & (!x14666x)) + ((x14659x) & (x14660x) & (!x467x) & (x14665x) & (x14666x)) + ((x14659x) & (x14660x) & (x467x) & (!x14665x) & (!x14666x)) + ((x14659x) & (x14660x) & (x467x) & (!x14665x) & (x14666x)) + ((x14659x) & (x14660x) & (x467x) & (x14665x) & (!x14666x)) + ((x14659x) & (x14660x) & (x467x) & (x14665x) & (x14666x)));
	assign n_n3685 = (((!x136x) & (!n_n5003) & (!n_n5002) & (!x299x) & (x14670x)) + ((!x136x) & (!n_n5003) & (!n_n5002) & (x299x) & (!x14670x)) + ((!x136x) & (!n_n5003) & (!n_n5002) & (x299x) & (x14670x)) + ((!x136x) & (!n_n5003) & (n_n5002) & (!x299x) & (!x14670x)) + ((!x136x) & (!n_n5003) & (n_n5002) & (!x299x) & (x14670x)) + ((!x136x) & (!n_n5003) & (n_n5002) & (x299x) & (!x14670x)) + ((!x136x) & (!n_n5003) & (n_n5002) & (x299x) & (x14670x)) + ((!x136x) & (n_n5003) & (!n_n5002) & (!x299x) & (!x14670x)) + ((!x136x) & (n_n5003) & (!n_n5002) & (!x299x) & (x14670x)) + ((!x136x) & (n_n5003) & (!n_n5002) & (x299x) & (!x14670x)) + ((!x136x) & (n_n5003) & (!n_n5002) & (x299x) & (x14670x)) + ((!x136x) & (n_n5003) & (n_n5002) & (!x299x) & (!x14670x)) + ((!x136x) & (n_n5003) & (n_n5002) & (!x299x) & (x14670x)) + ((!x136x) & (n_n5003) & (n_n5002) & (x299x) & (!x14670x)) + ((!x136x) & (n_n5003) & (n_n5002) & (x299x) & (x14670x)) + ((x136x) & (!n_n5003) & (!n_n5002) & (!x299x) & (!x14670x)) + ((x136x) & (!n_n5003) & (!n_n5002) & (!x299x) & (x14670x)) + ((x136x) & (!n_n5003) & (!n_n5002) & (x299x) & (!x14670x)) + ((x136x) & (!n_n5003) & (!n_n5002) & (x299x) & (x14670x)) + ((x136x) & (!n_n5003) & (n_n5002) & (!x299x) & (!x14670x)) + ((x136x) & (!n_n5003) & (n_n5002) & (!x299x) & (x14670x)) + ((x136x) & (!n_n5003) & (n_n5002) & (x299x) & (!x14670x)) + ((x136x) & (!n_n5003) & (n_n5002) & (x299x) & (x14670x)) + ((x136x) & (n_n5003) & (!n_n5002) & (!x299x) & (!x14670x)) + ((x136x) & (n_n5003) & (!n_n5002) & (!x299x) & (x14670x)) + ((x136x) & (n_n5003) & (!n_n5002) & (x299x) & (!x14670x)) + ((x136x) & (n_n5003) & (!n_n5002) & (x299x) & (x14670x)) + ((x136x) & (n_n5003) & (n_n5002) & (!x299x) & (!x14670x)) + ((x136x) & (n_n5003) & (n_n5002) & (!x299x) & (x14670x)) + ((x136x) & (n_n5003) & (n_n5002) & (x299x) & (!x14670x)) + ((x136x) & (n_n5003) & (n_n5002) & (x299x) & (x14670x)));
	assign n_n3686 = (((!n_n4995) & (!n_n4999) & (!x247x) & (!x41x) & (x104x)) + ((!n_n4995) & (!n_n4999) & (!x247x) & (x41x) & (!x104x)) + ((!n_n4995) & (!n_n4999) & (!x247x) & (x41x) & (x104x)) + ((!n_n4995) & (!n_n4999) & (x247x) & (!x41x) & (!x104x)) + ((!n_n4995) & (!n_n4999) & (x247x) & (!x41x) & (x104x)) + ((!n_n4995) & (!n_n4999) & (x247x) & (x41x) & (!x104x)) + ((!n_n4995) & (!n_n4999) & (x247x) & (x41x) & (x104x)) + ((!n_n4995) & (n_n4999) & (!x247x) & (!x41x) & (!x104x)) + ((!n_n4995) & (n_n4999) & (!x247x) & (!x41x) & (x104x)) + ((!n_n4995) & (n_n4999) & (!x247x) & (x41x) & (!x104x)) + ((!n_n4995) & (n_n4999) & (!x247x) & (x41x) & (x104x)) + ((!n_n4995) & (n_n4999) & (x247x) & (!x41x) & (!x104x)) + ((!n_n4995) & (n_n4999) & (x247x) & (!x41x) & (x104x)) + ((!n_n4995) & (n_n4999) & (x247x) & (x41x) & (!x104x)) + ((!n_n4995) & (n_n4999) & (x247x) & (x41x) & (x104x)) + ((n_n4995) & (!n_n4999) & (!x247x) & (!x41x) & (!x104x)) + ((n_n4995) & (!n_n4999) & (!x247x) & (!x41x) & (x104x)) + ((n_n4995) & (!n_n4999) & (!x247x) & (x41x) & (!x104x)) + ((n_n4995) & (!n_n4999) & (!x247x) & (x41x) & (x104x)) + ((n_n4995) & (!n_n4999) & (x247x) & (!x41x) & (!x104x)) + ((n_n4995) & (!n_n4999) & (x247x) & (!x41x) & (x104x)) + ((n_n4995) & (!n_n4999) & (x247x) & (x41x) & (!x104x)) + ((n_n4995) & (!n_n4999) & (x247x) & (x41x) & (x104x)) + ((n_n4995) & (n_n4999) & (!x247x) & (!x41x) & (!x104x)) + ((n_n4995) & (n_n4999) & (!x247x) & (!x41x) & (x104x)) + ((n_n4995) & (n_n4999) & (!x247x) & (x41x) & (!x104x)) + ((n_n4995) & (n_n4999) & (!x247x) & (x41x) & (x104x)) + ((n_n4995) & (n_n4999) & (x247x) & (!x41x) & (!x104x)) + ((n_n4995) & (n_n4999) & (x247x) & (!x41x) & (x104x)) + ((n_n4995) & (n_n4999) & (x247x) & (x41x) & (!x104x)) + ((n_n4995) & (n_n4999) & (x247x) & (x41x) & (x104x)));
	assign x14682x = (((!n_n5018) & (!n_n5017) & (!n_n5014) & (!n_n5020) & (x14681x)) + ((!n_n5018) & (!n_n5017) & (!n_n5014) & (n_n5020) & (!x14681x)) + ((!n_n5018) & (!n_n5017) & (!n_n5014) & (n_n5020) & (x14681x)) + ((!n_n5018) & (!n_n5017) & (n_n5014) & (!n_n5020) & (!x14681x)) + ((!n_n5018) & (!n_n5017) & (n_n5014) & (!n_n5020) & (x14681x)) + ((!n_n5018) & (!n_n5017) & (n_n5014) & (n_n5020) & (!x14681x)) + ((!n_n5018) & (!n_n5017) & (n_n5014) & (n_n5020) & (x14681x)) + ((!n_n5018) & (n_n5017) & (!n_n5014) & (!n_n5020) & (!x14681x)) + ((!n_n5018) & (n_n5017) & (!n_n5014) & (!n_n5020) & (x14681x)) + ((!n_n5018) & (n_n5017) & (!n_n5014) & (n_n5020) & (!x14681x)) + ((!n_n5018) & (n_n5017) & (!n_n5014) & (n_n5020) & (x14681x)) + ((!n_n5018) & (n_n5017) & (n_n5014) & (!n_n5020) & (!x14681x)) + ((!n_n5018) & (n_n5017) & (n_n5014) & (!n_n5020) & (x14681x)) + ((!n_n5018) & (n_n5017) & (n_n5014) & (n_n5020) & (!x14681x)) + ((!n_n5018) & (n_n5017) & (n_n5014) & (n_n5020) & (x14681x)) + ((n_n5018) & (!n_n5017) & (!n_n5014) & (!n_n5020) & (!x14681x)) + ((n_n5018) & (!n_n5017) & (!n_n5014) & (!n_n5020) & (x14681x)) + ((n_n5018) & (!n_n5017) & (!n_n5014) & (n_n5020) & (!x14681x)) + ((n_n5018) & (!n_n5017) & (!n_n5014) & (n_n5020) & (x14681x)) + ((n_n5018) & (!n_n5017) & (n_n5014) & (!n_n5020) & (!x14681x)) + ((n_n5018) & (!n_n5017) & (n_n5014) & (!n_n5020) & (x14681x)) + ((n_n5018) & (!n_n5017) & (n_n5014) & (n_n5020) & (!x14681x)) + ((n_n5018) & (!n_n5017) & (n_n5014) & (n_n5020) & (x14681x)) + ((n_n5018) & (n_n5017) & (!n_n5014) & (!n_n5020) & (!x14681x)) + ((n_n5018) & (n_n5017) & (!n_n5014) & (!n_n5020) & (x14681x)) + ((n_n5018) & (n_n5017) & (!n_n5014) & (n_n5020) & (!x14681x)) + ((n_n5018) & (n_n5017) & (!n_n5014) & (n_n5020) & (x14681x)) + ((n_n5018) & (n_n5017) & (n_n5014) & (!n_n5020) & (!x14681x)) + ((n_n5018) & (n_n5017) & (n_n5014) & (!n_n5020) & (x14681x)) + ((n_n5018) & (n_n5017) & (n_n5014) & (n_n5020) & (!x14681x)) + ((n_n5018) & (n_n5017) & (n_n5014) & (n_n5020) & (x14681x)));
	assign n_n3696 = (((!x40x) & (!x295x) & (!n_n4871) & (!x324x) & (x14687x)) + ((!x40x) & (!x295x) & (!n_n4871) & (x324x) & (!x14687x)) + ((!x40x) & (!x295x) & (!n_n4871) & (x324x) & (x14687x)) + ((!x40x) & (!x295x) & (n_n4871) & (!x324x) & (!x14687x)) + ((!x40x) & (!x295x) & (n_n4871) & (!x324x) & (x14687x)) + ((!x40x) & (!x295x) & (n_n4871) & (x324x) & (!x14687x)) + ((!x40x) & (!x295x) & (n_n4871) & (x324x) & (x14687x)) + ((!x40x) & (x295x) & (!n_n4871) & (!x324x) & (!x14687x)) + ((!x40x) & (x295x) & (!n_n4871) & (!x324x) & (x14687x)) + ((!x40x) & (x295x) & (!n_n4871) & (x324x) & (!x14687x)) + ((!x40x) & (x295x) & (!n_n4871) & (x324x) & (x14687x)) + ((!x40x) & (x295x) & (n_n4871) & (!x324x) & (!x14687x)) + ((!x40x) & (x295x) & (n_n4871) & (!x324x) & (x14687x)) + ((!x40x) & (x295x) & (n_n4871) & (x324x) & (!x14687x)) + ((!x40x) & (x295x) & (n_n4871) & (x324x) & (x14687x)) + ((x40x) & (!x295x) & (!n_n4871) & (!x324x) & (!x14687x)) + ((x40x) & (!x295x) & (!n_n4871) & (!x324x) & (x14687x)) + ((x40x) & (!x295x) & (!n_n4871) & (x324x) & (!x14687x)) + ((x40x) & (!x295x) & (!n_n4871) & (x324x) & (x14687x)) + ((x40x) & (!x295x) & (n_n4871) & (!x324x) & (!x14687x)) + ((x40x) & (!x295x) & (n_n4871) & (!x324x) & (x14687x)) + ((x40x) & (!x295x) & (n_n4871) & (x324x) & (!x14687x)) + ((x40x) & (!x295x) & (n_n4871) & (x324x) & (x14687x)) + ((x40x) & (x295x) & (!n_n4871) & (!x324x) & (!x14687x)) + ((x40x) & (x295x) & (!n_n4871) & (!x324x) & (x14687x)) + ((x40x) & (x295x) & (!n_n4871) & (x324x) & (!x14687x)) + ((x40x) & (x295x) & (!n_n4871) & (x324x) & (x14687x)) + ((x40x) & (x295x) & (n_n4871) & (!x324x) & (!x14687x)) + ((x40x) & (x295x) & (n_n4871) & (!x324x) & (x14687x)) + ((x40x) & (x295x) & (n_n4871) & (x324x) & (!x14687x)) + ((x40x) & (x295x) & (n_n4871) & (x324x) & (x14687x)));
	assign n_n3698 = (((!n_n4847) & (!n_n4846) & (!n_n4844) & (!x375x) & (!x22111x)) + ((!n_n4847) & (!n_n4846) & (!n_n4844) & (x375x) & (!x22111x)) + ((!n_n4847) & (!n_n4846) & (!n_n4844) & (x375x) & (x22111x)) + ((!n_n4847) & (!n_n4846) & (n_n4844) & (!x375x) & (!x22111x)) + ((!n_n4847) & (!n_n4846) & (n_n4844) & (!x375x) & (x22111x)) + ((!n_n4847) & (!n_n4846) & (n_n4844) & (x375x) & (!x22111x)) + ((!n_n4847) & (!n_n4846) & (n_n4844) & (x375x) & (x22111x)) + ((!n_n4847) & (n_n4846) & (!n_n4844) & (!x375x) & (!x22111x)) + ((!n_n4847) & (n_n4846) & (!n_n4844) & (!x375x) & (x22111x)) + ((!n_n4847) & (n_n4846) & (!n_n4844) & (x375x) & (!x22111x)) + ((!n_n4847) & (n_n4846) & (!n_n4844) & (x375x) & (x22111x)) + ((!n_n4847) & (n_n4846) & (n_n4844) & (!x375x) & (!x22111x)) + ((!n_n4847) & (n_n4846) & (n_n4844) & (!x375x) & (x22111x)) + ((!n_n4847) & (n_n4846) & (n_n4844) & (x375x) & (!x22111x)) + ((!n_n4847) & (n_n4846) & (n_n4844) & (x375x) & (x22111x)) + ((n_n4847) & (!n_n4846) & (!n_n4844) & (!x375x) & (!x22111x)) + ((n_n4847) & (!n_n4846) & (!n_n4844) & (!x375x) & (x22111x)) + ((n_n4847) & (!n_n4846) & (!n_n4844) & (x375x) & (!x22111x)) + ((n_n4847) & (!n_n4846) & (!n_n4844) & (x375x) & (x22111x)) + ((n_n4847) & (!n_n4846) & (n_n4844) & (!x375x) & (!x22111x)) + ((n_n4847) & (!n_n4846) & (n_n4844) & (!x375x) & (x22111x)) + ((n_n4847) & (!n_n4846) & (n_n4844) & (x375x) & (!x22111x)) + ((n_n4847) & (!n_n4846) & (n_n4844) & (x375x) & (x22111x)) + ((n_n4847) & (n_n4846) & (!n_n4844) & (!x375x) & (!x22111x)) + ((n_n4847) & (n_n4846) & (!n_n4844) & (!x375x) & (x22111x)) + ((n_n4847) & (n_n4846) & (!n_n4844) & (x375x) & (!x22111x)) + ((n_n4847) & (n_n4846) & (!n_n4844) & (x375x) & (x22111x)) + ((n_n4847) & (n_n4846) & (n_n4844) & (!x375x) & (!x22111x)) + ((n_n4847) & (n_n4846) & (n_n4844) & (!x375x) & (x22111x)) + ((n_n4847) & (n_n4846) & (n_n4844) & (x375x) & (!x22111x)) + ((n_n4847) & (n_n4846) & (n_n4844) & (x375x) & (x22111x)));
	assign x14728x = (((!n_n4857) & (!n_n4856) & (!n_n4854) & (!n_n4855) & (x14727x)) + ((!n_n4857) & (!n_n4856) & (!n_n4854) & (n_n4855) & (!x14727x)) + ((!n_n4857) & (!n_n4856) & (!n_n4854) & (n_n4855) & (x14727x)) + ((!n_n4857) & (!n_n4856) & (n_n4854) & (!n_n4855) & (!x14727x)) + ((!n_n4857) & (!n_n4856) & (n_n4854) & (!n_n4855) & (x14727x)) + ((!n_n4857) & (!n_n4856) & (n_n4854) & (n_n4855) & (!x14727x)) + ((!n_n4857) & (!n_n4856) & (n_n4854) & (n_n4855) & (x14727x)) + ((!n_n4857) & (n_n4856) & (!n_n4854) & (!n_n4855) & (!x14727x)) + ((!n_n4857) & (n_n4856) & (!n_n4854) & (!n_n4855) & (x14727x)) + ((!n_n4857) & (n_n4856) & (!n_n4854) & (n_n4855) & (!x14727x)) + ((!n_n4857) & (n_n4856) & (!n_n4854) & (n_n4855) & (x14727x)) + ((!n_n4857) & (n_n4856) & (n_n4854) & (!n_n4855) & (!x14727x)) + ((!n_n4857) & (n_n4856) & (n_n4854) & (!n_n4855) & (x14727x)) + ((!n_n4857) & (n_n4856) & (n_n4854) & (n_n4855) & (!x14727x)) + ((!n_n4857) & (n_n4856) & (n_n4854) & (n_n4855) & (x14727x)) + ((n_n4857) & (!n_n4856) & (!n_n4854) & (!n_n4855) & (!x14727x)) + ((n_n4857) & (!n_n4856) & (!n_n4854) & (!n_n4855) & (x14727x)) + ((n_n4857) & (!n_n4856) & (!n_n4854) & (n_n4855) & (!x14727x)) + ((n_n4857) & (!n_n4856) & (!n_n4854) & (n_n4855) & (x14727x)) + ((n_n4857) & (!n_n4856) & (n_n4854) & (!n_n4855) & (!x14727x)) + ((n_n4857) & (!n_n4856) & (n_n4854) & (!n_n4855) & (x14727x)) + ((n_n4857) & (!n_n4856) & (n_n4854) & (n_n4855) & (!x14727x)) + ((n_n4857) & (!n_n4856) & (n_n4854) & (n_n4855) & (x14727x)) + ((n_n4857) & (n_n4856) & (!n_n4854) & (!n_n4855) & (!x14727x)) + ((n_n4857) & (n_n4856) & (!n_n4854) & (!n_n4855) & (x14727x)) + ((n_n4857) & (n_n4856) & (!n_n4854) & (n_n4855) & (!x14727x)) + ((n_n4857) & (n_n4856) & (!n_n4854) & (n_n4855) & (x14727x)) + ((n_n4857) & (n_n4856) & (n_n4854) & (!n_n4855) & (!x14727x)) + ((n_n4857) & (n_n4856) & (n_n4854) & (!n_n4855) & (x14727x)) + ((n_n4857) & (n_n4856) & (n_n4854) & (n_n4855) & (!x14727x)) + ((n_n4857) & (n_n4856) & (n_n4854) & (n_n4855) & (x14727x)));
	assign x14730x = (((!n_n3696) & (!n_n3698) & (x14728x)) + ((!n_n3696) & (n_n3698) & (!x14728x)) + ((!n_n3696) & (n_n3698) & (x14728x)) + ((n_n3696) & (!n_n3698) & (!x14728x)) + ((n_n3696) & (!n_n3698) & (x14728x)) + ((n_n3696) & (n_n3698) & (!x14728x)) + ((n_n3696) & (n_n3698) & (x14728x)));
	assign n_n3645 = (((!n_n3701) & (!x14708x) & (!x14709x) & (!x22110x)) + ((!n_n3701) & (!x14708x) & (x14709x) & (!x22110x)) + ((!n_n3701) & (!x14708x) & (x14709x) & (x22110x)) + ((!n_n3701) & (x14708x) & (!x14709x) & (!x22110x)) + ((!n_n3701) & (x14708x) & (!x14709x) & (x22110x)) + ((!n_n3701) & (x14708x) & (x14709x) & (!x22110x)) + ((!n_n3701) & (x14708x) & (x14709x) & (x22110x)) + ((n_n3701) & (!x14708x) & (!x14709x) & (!x22110x)) + ((n_n3701) & (!x14708x) & (!x14709x) & (x22110x)) + ((n_n3701) & (!x14708x) & (x14709x) & (!x22110x)) + ((n_n3701) & (!x14708x) & (x14709x) & (x22110x)) + ((n_n3701) & (x14708x) & (!x14709x) & (!x22110x)) + ((n_n3701) & (x14708x) & (!x14709x) & (x22110x)) + ((n_n3701) & (x14708x) & (x14709x) & (!x22110x)) + ((n_n3701) & (x14708x) & (x14709x) & (x22110x)));
	assign n_n3702 = (((!x179x) & (!n_n4799) & (!x380x) & (!x381x) & (x14712x)) + ((!x179x) & (!n_n4799) & (!x380x) & (x381x) & (!x14712x)) + ((!x179x) & (!n_n4799) & (!x380x) & (x381x) & (x14712x)) + ((!x179x) & (!n_n4799) & (x380x) & (!x381x) & (!x14712x)) + ((!x179x) & (!n_n4799) & (x380x) & (!x381x) & (x14712x)) + ((!x179x) & (!n_n4799) & (x380x) & (x381x) & (!x14712x)) + ((!x179x) & (!n_n4799) & (x380x) & (x381x) & (x14712x)) + ((!x179x) & (n_n4799) & (!x380x) & (!x381x) & (!x14712x)) + ((!x179x) & (n_n4799) & (!x380x) & (!x381x) & (x14712x)) + ((!x179x) & (n_n4799) & (!x380x) & (x381x) & (!x14712x)) + ((!x179x) & (n_n4799) & (!x380x) & (x381x) & (x14712x)) + ((!x179x) & (n_n4799) & (x380x) & (!x381x) & (!x14712x)) + ((!x179x) & (n_n4799) & (x380x) & (!x381x) & (x14712x)) + ((!x179x) & (n_n4799) & (x380x) & (x381x) & (!x14712x)) + ((!x179x) & (n_n4799) & (x380x) & (x381x) & (x14712x)) + ((x179x) & (!n_n4799) & (!x380x) & (!x381x) & (!x14712x)) + ((x179x) & (!n_n4799) & (!x380x) & (!x381x) & (x14712x)) + ((x179x) & (!n_n4799) & (!x380x) & (x381x) & (!x14712x)) + ((x179x) & (!n_n4799) & (!x380x) & (x381x) & (x14712x)) + ((x179x) & (!n_n4799) & (x380x) & (!x381x) & (!x14712x)) + ((x179x) & (!n_n4799) & (x380x) & (!x381x) & (x14712x)) + ((x179x) & (!n_n4799) & (x380x) & (x381x) & (!x14712x)) + ((x179x) & (!n_n4799) & (x380x) & (x381x) & (x14712x)) + ((x179x) & (n_n4799) & (!x380x) & (!x381x) & (!x14712x)) + ((x179x) & (n_n4799) & (!x380x) & (!x381x) & (x14712x)) + ((x179x) & (n_n4799) & (!x380x) & (x381x) & (!x14712x)) + ((x179x) & (n_n4799) & (!x380x) & (x381x) & (x14712x)) + ((x179x) & (n_n4799) & (x380x) & (!x381x) & (!x14712x)) + ((x179x) & (n_n4799) & (x380x) & (!x381x) & (x14712x)) + ((x179x) & (n_n4799) & (x380x) & (x381x) & (!x14712x)) + ((x179x) & (n_n4799) & (x380x) & (x381x) & (x14712x)));
	assign x14722x = (((!n_n4786) & (!n_n4783) & (!n_n4205) & (!n_n4204) & (x12394x)) + ((!n_n4786) & (!n_n4783) & (!n_n4205) & (n_n4204) & (!x12394x)) + ((!n_n4786) & (!n_n4783) & (!n_n4205) & (n_n4204) & (x12394x)) + ((!n_n4786) & (!n_n4783) & (n_n4205) & (!n_n4204) & (!x12394x)) + ((!n_n4786) & (!n_n4783) & (n_n4205) & (!n_n4204) & (x12394x)) + ((!n_n4786) & (!n_n4783) & (n_n4205) & (n_n4204) & (!x12394x)) + ((!n_n4786) & (!n_n4783) & (n_n4205) & (n_n4204) & (x12394x)) + ((!n_n4786) & (n_n4783) & (!n_n4205) & (!n_n4204) & (!x12394x)) + ((!n_n4786) & (n_n4783) & (!n_n4205) & (!n_n4204) & (x12394x)) + ((!n_n4786) & (n_n4783) & (!n_n4205) & (n_n4204) & (!x12394x)) + ((!n_n4786) & (n_n4783) & (!n_n4205) & (n_n4204) & (x12394x)) + ((!n_n4786) & (n_n4783) & (n_n4205) & (!n_n4204) & (!x12394x)) + ((!n_n4786) & (n_n4783) & (n_n4205) & (!n_n4204) & (x12394x)) + ((!n_n4786) & (n_n4783) & (n_n4205) & (n_n4204) & (!x12394x)) + ((!n_n4786) & (n_n4783) & (n_n4205) & (n_n4204) & (x12394x)) + ((n_n4786) & (!n_n4783) & (!n_n4205) & (!n_n4204) & (!x12394x)) + ((n_n4786) & (!n_n4783) & (!n_n4205) & (!n_n4204) & (x12394x)) + ((n_n4786) & (!n_n4783) & (!n_n4205) & (n_n4204) & (!x12394x)) + ((n_n4786) & (!n_n4783) & (!n_n4205) & (n_n4204) & (x12394x)) + ((n_n4786) & (!n_n4783) & (n_n4205) & (!n_n4204) & (!x12394x)) + ((n_n4786) & (!n_n4783) & (n_n4205) & (!n_n4204) & (x12394x)) + ((n_n4786) & (!n_n4783) & (n_n4205) & (n_n4204) & (!x12394x)) + ((n_n4786) & (!n_n4783) & (n_n4205) & (n_n4204) & (x12394x)) + ((n_n4786) & (n_n4783) & (!n_n4205) & (!n_n4204) & (!x12394x)) + ((n_n4786) & (n_n4783) & (!n_n4205) & (!n_n4204) & (x12394x)) + ((n_n4786) & (n_n4783) & (!n_n4205) & (n_n4204) & (!x12394x)) + ((n_n4786) & (n_n4783) & (!n_n4205) & (n_n4204) & (x12394x)) + ((n_n4786) & (n_n4783) & (n_n4205) & (!n_n4204) & (!x12394x)) + ((n_n4786) & (n_n4783) & (n_n4205) & (!n_n4204) & (x12394x)) + ((n_n4786) & (n_n4783) & (n_n4205) & (n_n4204) & (!x12394x)) + ((n_n4786) & (n_n4783) & (n_n4205) & (n_n4204) & (x12394x)));
	assign x14721x = (((!n_n4782) & (!n_n4779) & (!n_n4790) & (!n_n4781) & (x14718x)) + ((!n_n4782) & (!n_n4779) & (!n_n4790) & (n_n4781) & (!x14718x)) + ((!n_n4782) & (!n_n4779) & (!n_n4790) & (n_n4781) & (x14718x)) + ((!n_n4782) & (!n_n4779) & (n_n4790) & (!n_n4781) & (!x14718x)) + ((!n_n4782) & (!n_n4779) & (n_n4790) & (!n_n4781) & (x14718x)) + ((!n_n4782) & (!n_n4779) & (n_n4790) & (n_n4781) & (!x14718x)) + ((!n_n4782) & (!n_n4779) & (n_n4790) & (n_n4781) & (x14718x)) + ((!n_n4782) & (n_n4779) & (!n_n4790) & (!n_n4781) & (!x14718x)) + ((!n_n4782) & (n_n4779) & (!n_n4790) & (!n_n4781) & (x14718x)) + ((!n_n4782) & (n_n4779) & (!n_n4790) & (n_n4781) & (!x14718x)) + ((!n_n4782) & (n_n4779) & (!n_n4790) & (n_n4781) & (x14718x)) + ((!n_n4782) & (n_n4779) & (n_n4790) & (!n_n4781) & (!x14718x)) + ((!n_n4782) & (n_n4779) & (n_n4790) & (!n_n4781) & (x14718x)) + ((!n_n4782) & (n_n4779) & (n_n4790) & (n_n4781) & (!x14718x)) + ((!n_n4782) & (n_n4779) & (n_n4790) & (n_n4781) & (x14718x)) + ((n_n4782) & (!n_n4779) & (!n_n4790) & (!n_n4781) & (!x14718x)) + ((n_n4782) & (!n_n4779) & (!n_n4790) & (!n_n4781) & (x14718x)) + ((n_n4782) & (!n_n4779) & (!n_n4790) & (n_n4781) & (!x14718x)) + ((n_n4782) & (!n_n4779) & (!n_n4790) & (n_n4781) & (x14718x)) + ((n_n4782) & (!n_n4779) & (n_n4790) & (!n_n4781) & (!x14718x)) + ((n_n4782) & (!n_n4779) & (n_n4790) & (!n_n4781) & (x14718x)) + ((n_n4782) & (!n_n4779) & (n_n4790) & (n_n4781) & (!x14718x)) + ((n_n4782) & (!n_n4779) & (n_n4790) & (n_n4781) & (x14718x)) + ((n_n4782) & (n_n4779) & (!n_n4790) & (!n_n4781) & (!x14718x)) + ((n_n4782) & (n_n4779) & (!n_n4790) & (!n_n4781) & (x14718x)) + ((n_n4782) & (n_n4779) & (!n_n4790) & (n_n4781) & (!x14718x)) + ((n_n4782) & (n_n4779) & (!n_n4790) & (n_n4781) & (x14718x)) + ((n_n4782) & (n_n4779) & (n_n4790) & (!n_n4781) & (!x14718x)) + ((n_n4782) & (n_n4779) & (n_n4790) & (!n_n4781) & (x14718x)) + ((n_n4782) & (n_n4779) & (n_n4790) & (n_n4781) & (!x14718x)) + ((n_n4782) & (n_n4779) & (n_n4790) & (n_n4781) & (x14718x)));
	assign n_n3694 = (((!n_n4885) & (!n_n4890) & (!x264x) & (!n_n3810) & (x261x)) + ((!n_n4885) & (!n_n4890) & (!x264x) & (n_n3810) & (!x261x)) + ((!n_n4885) & (!n_n4890) & (!x264x) & (n_n3810) & (x261x)) + ((!n_n4885) & (!n_n4890) & (x264x) & (!n_n3810) & (!x261x)) + ((!n_n4885) & (!n_n4890) & (x264x) & (!n_n3810) & (x261x)) + ((!n_n4885) & (!n_n4890) & (x264x) & (n_n3810) & (!x261x)) + ((!n_n4885) & (!n_n4890) & (x264x) & (n_n3810) & (x261x)) + ((!n_n4885) & (n_n4890) & (!x264x) & (!n_n3810) & (!x261x)) + ((!n_n4885) & (n_n4890) & (!x264x) & (!n_n3810) & (x261x)) + ((!n_n4885) & (n_n4890) & (!x264x) & (n_n3810) & (!x261x)) + ((!n_n4885) & (n_n4890) & (!x264x) & (n_n3810) & (x261x)) + ((!n_n4885) & (n_n4890) & (x264x) & (!n_n3810) & (!x261x)) + ((!n_n4885) & (n_n4890) & (x264x) & (!n_n3810) & (x261x)) + ((!n_n4885) & (n_n4890) & (x264x) & (n_n3810) & (!x261x)) + ((!n_n4885) & (n_n4890) & (x264x) & (n_n3810) & (x261x)) + ((n_n4885) & (!n_n4890) & (!x264x) & (!n_n3810) & (!x261x)) + ((n_n4885) & (!n_n4890) & (!x264x) & (!n_n3810) & (x261x)) + ((n_n4885) & (!n_n4890) & (!x264x) & (n_n3810) & (!x261x)) + ((n_n4885) & (!n_n4890) & (!x264x) & (n_n3810) & (x261x)) + ((n_n4885) & (!n_n4890) & (x264x) & (!n_n3810) & (!x261x)) + ((n_n4885) & (!n_n4890) & (x264x) & (!n_n3810) & (x261x)) + ((n_n4885) & (!n_n4890) & (x264x) & (n_n3810) & (!x261x)) + ((n_n4885) & (!n_n4890) & (x264x) & (n_n3810) & (x261x)) + ((n_n4885) & (n_n4890) & (!x264x) & (!n_n3810) & (!x261x)) + ((n_n4885) & (n_n4890) & (!x264x) & (!n_n3810) & (x261x)) + ((n_n4885) & (n_n4890) & (!x264x) & (n_n3810) & (!x261x)) + ((n_n4885) & (n_n4890) & (!x264x) & (n_n3810) & (x261x)) + ((n_n4885) & (n_n4890) & (x264x) & (!n_n3810) & (!x261x)) + ((n_n4885) & (n_n4890) & (x264x) & (!n_n3810) & (x261x)) + ((n_n4885) & (n_n4890) & (x264x) & (n_n3810) & (!x261x)) + ((n_n4885) & (n_n4890) & (x264x) & (n_n3810) & (x261x)));
	assign n_n3693 = (((!n_n4900) & (!n_n4903) & (!n_n4908) & (!n_n4899) & (x14739x)) + ((!n_n4900) & (!n_n4903) & (!n_n4908) & (n_n4899) & (!x14739x)) + ((!n_n4900) & (!n_n4903) & (!n_n4908) & (n_n4899) & (x14739x)) + ((!n_n4900) & (!n_n4903) & (n_n4908) & (!n_n4899) & (!x14739x)) + ((!n_n4900) & (!n_n4903) & (n_n4908) & (!n_n4899) & (x14739x)) + ((!n_n4900) & (!n_n4903) & (n_n4908) & (n_n4899) & (!x14739x)) + ((!n_n4900) & (!n_n4903) & (n_n4908) & (n_n4899) & (x14739x)) + ((!n_n4900) & (n_n4903) & (!n_n4908) & (!n_n4899) & (!x14739x)) + ((!n_n4900) & (n_n4903) & (!n_n4908) & (!n_n4899) & (x14739x)) + ((!n_n4900) & (n_n4903) & (!n_n4908) & (n_n4899) & (!x14739x)) + ((!n_n4900) & (n_n4903) & (!n_n4908) & (n_n4899) & (x14739x)) + ((!n_n4900) & (n_n4903) & (n_n4908) & (!n_n4899) & (!x14739x)) + ((!n_n4900) & (n_n4903) & (n_n4908) & (!n_n4899) & (x14739x)) + ((!n_n4900) & (n_n4903) & (n_n4908) & (n_n4899) & (!x14739x)) + ((!n_n4900) & (n_n4903) & (n_n4908) & (n_n4899) & (x14739x)) + ((n_n4900) & (!n_n4903) & (!n_n4908) & (!n_n4899) & (!x14739x)) + ((n_n4900) & (!n_n4903) & (!n_n4908) & (!n_n4899) & (x14739x)) + ((n_n4900) & (!n_n4903) & (!n_n4908) & (n_n4899) & (!x14739x)) + ((n_n4900) & (!n_n4903) & (!n_n4908) & (n_n4899) & (x14739x)) + ((n_n4900) & (!n_n4903) & (n_n4908) & (!n_n4899) & (!x14739x)) + ((n_n4900) & (!n_n4903) & (n_n4908) & (!n_n4899) & (x14739x)) + ((n_n4900) & (!n_n4903) & (n_n4908) & (n_n4899) & (!x14739x)) + ((n_n4900) & (!n_n4903) & (n_n4908) & (n_n4899) & (x14739x)) + ((n_n4900) & (n_n4903) & (!n_n4908) & (!n_n4899) & (!x14739x)) + ((n_n4900) & (n_n4903) & (!n_n4908) & (!n_n4899) & (x14739x)) + ((n_n4900) & (n_n4903) & (!n_n4908) & (n_n4899) & (!x14739x)) + ((n_n4900) & (n_n4903) & (!n_n4908) & (n_n4899) & (x14739x)) + ((n_n4900) & (n_n4903) & (n_n4908) & (!n_n4899) & (!x14739x)) + ((n_n4900) & (n_n4903) & (n_n4908) & (!n_n4899) & (x14739x)) + ((n_n4900) & (n_n4903) & (n_n4908) & (n_n4899) & (!x14739x)) + ((n_n4900) & (n_n4903) & (n_n4908) & (n_n4899) & (x14739x)));
	assign n_n3642 = (((!x142x) & (!n_n3691) & (!x14748x) & (x14749x)) + ((!x142x) & (!n_n3691) & (x14748x) & (!x14749x)) + ((!x142x) & (!n_n3691) & (x14748x) & (x14749x)) + ((!x142x) & (n_n3691) & (!x14748x) & (!x14749x)) + ((!x142x) & (n_n3691) & (!x14748x) & (x14749x)) + ((!x142x) & (n_n3691) & (x14748x) & (!x14749x)) + ((!x142x) & (n_n3691) & (x14748x) & (x14749x)) + ((x142x) & (!n_n3691) & (!x14748x) & (!x14749x)) + ((x142x) & (!n_n3691) & (!x14748x) & (x14749x)) + ((x142x) & (!n_n3691) & (x14748x) & (!x14749x)) + ((x142x) & (!n_n3691) & (x14748x) & (x14749x)) + ((x142x) & (n_n3691) & (!x14748x) & (!x14749x)) + ((x142x) & (n_n3691) & (!x14748x) & (x14749x)) + ((x142x) & (n_n3691) & (x14748x) & (!x14749x)) + ((x142x) & (n_n3691) & (x14748x) & (x14749x)));
	assign n_n3641 = (((!n_n3803) & (!n_n3802) & (!x14754x) & (!x14764x) & (x14763x)) + ((!n_n3803) & (!n_n3802) & (!x14754x) & (x14764x) & (!x14763x)) + ((!n_n3803) & (!n_n3802) & (!x14754x) & (x14764x) & (x14763x)) + ((!n_n3803) & (!n_n3802) & (x14754x) & (!x14764x) & (!x14763x)) + ((!n_n3803) & (!n_n3802) & (x14754x) & (!x14764x) & (x14763x)) + ((!n_n3803) & (!n_n3802) & (x14754x) & (x14764x) & (!x14763x)) + ((!n_n3803) & (!n_n3802) & (x14754x) & (x14764x) & (x14763x)) + ((!n_n3803) & (n_n3802) & (!x14754x) & (!x14764x) & (!x14763x)) + ((!n_n3803) & (n_n3802) & (!x14754x) & (!x14764x) & (x14763x)) + ((!n_n3803) & (n_n3802) & (!x14754x) & (x14764x) & (!x14763x)) + ((!n_n3803) & (n_n3802) & (!x14754x) & (x14764x) & (x14763x)) + ((!n_n3803) & (n_n3802) & (x14754x) & (!x14764x) & (!x14763x)) + ((!n_n3803) & (n_n3802) & (x14754x) & (!x14764x) & (x14763x)) + ((!n_n3803) & (n_n3802) & (x14754x) & (x14764x) & (!x14763x)) + ((!n_n3803) & (n_n3802) & (x14754x) & (x14764x) & (x14763x)) + ((n_n3803) & (!n_n3802) & (!x14754x) & (!x14764x) & (!x14763x)) + ((n_n3803) & (!n_n3802) & (!x14754x) & (!x14764x) & (x14763x)) + ((n_n3803) & (!n_n3802) & (!x14754x) & (x14764x) & (!x14763x)) + ((n_n3803) & (!n_n3802) & (!x14754x) & (x14764x) & (x14763x)) + ((n_n3803) & (!n_n3802) & (x14754x) & (!x14764x) & (!x14763x)) + ((n_n3803) & (!n_n3802) & (x14754x) & (!x14764x) & (x14763x)) + ((n_n3803) & (!n_n3802) & (x14754x) & (x14764x) & (!x14763x)) + ((n_n3803) & (!n_n3802) & (x14754x) & (x14764x) & (x14763x)) + ((n_n3803) & (n_n3802) & (!x14754x) & (!x14764x) & (!x14763x)) + ((n_n3803) & (n_n3802) & (!x14754x) & (!x14764x) & (x14763x)) + ((n_n3803) & (n_n3802) & (!x14754x) & (x14764x) & (!x14763x)) + ((n_n3803) & (n_n3802) & (!x14754x) & (x14764x) & (x14763x)) + ((n_n3803) & (n_n3802) & (x14754x) & (!x14764x) & (!x14763x)) + ((n_n3803) & (n_n3802) & (x14754x) & (!x14764x) & (x14763x)) + ((n_n3803) & (n_n3802) & (x14754x) & (x14764x) & (!x14763x)) + ((n_n3803) & (n_n3802) & (x14754x) & (x14764x) & (x14763x)));
	assign x14770x = (((!n_n4882) & (!n_n4881) & (!n_n4878) & (!n_n4880) & (x14769x)) + ((!n_n4882) & (!n_n4881) & (!n_n4878) & (n_n4880) & (!x14769x)) + ((!n_n4882) & (!n_n4881) & (!n_n4878) & (n_n4880) & (x14769x)) + ((!n_n4882) & (!n_n4881) & (n_n4878) & (!n_n4880) & (!x14769x)) + ((!n_n4882) & (!n_n4881) & (n_n4878) & (!n_n4880) & (x14769x)) + ((!n_n4882) & (!n_n4881) & (n_n4878) & (n_n4880) & (!x14769x)) + ((!n_n4882) & (!n_n4881) & (n_n4878) & (n_n4880) & (x14769x)) + ((!n_n4882) & (n_n4881) & (!n_n4878) & (!n_n4880) & (!x14769x)) + ((!n_n4882) & (n_n4881) & (!n_n4878) & (!n_n4880) & (x14769x)) + ((!n_n4882) & (n_n4881) & (!n_n4878) & (n_n4880) & (!x14769x)) + ((!n_n4882) & (n_n4881) & (!n_n4878) & (n_n4880) & (x14769x)) + ((!n_n4882) & (n_n4881) & (n_n4878) & (!n_n4880) & (!x14769x)) + ((!n_n4882) & (n_n4881) & (n_n4878) & (!n_n4880) & (x14769x)) + ((!n_n4882) & (n_n4881) & (n_n4878) & (n_n4880) & (!x14769x)) + ((!n_n4882) & (n_n4881) & (n_n4878) & (n_n4880) & (x14769x)) + ((n_n4882) & (!n_n4881) & (!n_n4878) & (!n_n4880) & (!x14769x)) + ((n_n4882) & (!n_n4881) & (!n_n4878) & (!n_n4880) & (x14769x)) + ((n_n4882) & (!n_n4881) & (!n_n4878) & (n_n4880) & (!x14769x)) + ((n_n4882) & (!n_n4881) & (!n_n4878) & (n_n4880) & (x14769x)) + ((n_n4882) & (!n_n4881) & (n_n4878) & (!n_n4880) & (!x14769x)) + ((n_n4882) & (!n_n4881) & (n_n4878) & (!n_n4880) & (x14769x)) + ((n_n4882) & (!n_n4881) & (n_n4878) & (n_n4880) & (!x14769x)) + ((n_n4882) & (!n_n4881) & (n_n4878) & (n_n4880) & (x14769x)) + ((n_n4882) & (n_n4881) & (!n_n4878) & (!n_n4880) & (!x14769x)) + ((n_n4882) & (n_n4881) & (!n_n4878) & (!n_n4880) & (x14769x)) + ((n_n4882) & (n_n4881) & (!n_n4878) & (n_n4880) & (!x14769x)) + ((n_n4882) & (n_n4881) & (!n_n4878) & (n_n4880) & (x14769x)) + ((n_n4882) & (n_n4881) & (n_n4878) & (!n_n4880) & (!x14769x)) + ((n_n4882) & (n_n4881) & (n_n4878) & (!n_n4880) & (x14769x)) + ((n_n4882) & (n_n4881) & (n_n4878) & (n_n4880) & (!x14769x)) + ((n_n4882) & (n_n4881) & (n_n4878) & (n_n4880) & (x14769x)));
	assign n_n3626 = (((!n_n3694) & (!n_n3693) & (!n_n3642) & (!n_n3641) & (x14770x)) + ((!n_n3694) & (!n_n3693) & (!n_n3642) & (n_n3641) & (!x14770x)) + ((!n_n3694) & (!n_n3693) & (!n_n3642) & (n_n3641) & (x14770x)) + ((!n_n3694) & (!n_n3693) & (n_n3642) & (!n_n3641) & (!x14770x)) + ((!n_n3694) & (!n_n3693) & (n_n3642) & (!n_n3641) & (x14770x)) + ((!n_n3694) & (!n_n3693) & (n_n3642) & (n_n3641) & (!x14770x)) + ((!n_n3694) & (!n_n3693) & (n_n3642) & (n_n3641) & (x14770x)) + ((!n_n3694) & (n_n3693) & (!n_n3642) & (!n_n3641) & (!x14770x)) + ((!n_n3694) & (n_n3693) & (!n_n3642) & (!n_n3641) & (x14770x)) + ((!n_n3694) & (n_n3693) & (!n_n3642) & (n_n3641) & (!x14770x)) + ((!n_n3694) & (n_n3693) & (!n_n3642) & (n_n3641) & (x14770x)) + ((!n_n3694) & (n_n3693) & (n_n3642) & (!n_n3641) & (!x14770x)) + ((!n_n3694) & (n_n3693) & (n_n3642) & (!n_n3641) & (x14770x)) + ((!n_n3694) & (n_n3693) & (n_n3642) & (n_n3641) & (!x14770x)) + ((!n_n3694) & (n_n3693) & (n_n3642) & (n_n3641) & (x14770x)) + ((n_n3694) & (!n_n3693) & (!n_n3642) & (!n_n3641) & (!x14770x)) + ((n_n3694) & (!n_n3693) & (!n_n3642) & (!n_n3641) & (x14770x)) + ((n_n3694) & (!n_n3693) & (!n_n3642) & (n_n3641) & (!x14770x)) + ((n_n3694) & (!n_n3693) & (!n_n3642) & (n_n3641) & (x14770x)) + ((n_n3694) & (!n_n3693) & (n_n3642) & (!n_n3641) & (!x14770x)) + ((n_n3694) & (!n_n3693) & (n_n3642) & (!n_n3641) & (x14770x)) + ((n_n3694) & (!n_n3693) & (n_n3642) & (n_n3641) & (!x14770x)) + ((n_n3694) & (!n_n3693) & (n_n3642) & (n_n3641) & (x14770x)) + ((n_n3694) & (n_n3693) & (!n_n3642) & (!n_n3641) & (!x14770x)) + ((n_n3694) & (n_n3693) & (!n_n3642) & (!n_n3641) & (x14770x)) + ((n_n3694) & (n_n3693) & (!n_n3642) & (n_n3641) & (!x14770x)) + ((n_n3694) & (n_n3693) & (!n_n3642) & (n_n3641) & (x14770x)) + ((n_n3694) & (n_n3693) & (n_n3642) & (!n_n3641) & (!x14770x)) + ((n_n3694) & (n_n3693) & (n_n3642) & (!n_n3641) & (x14770x)) + ((n_n3694) & (n_n3693) & (n_n3642) & (n_n3641) & (!x14770x)) + ((n_n3694) & (n_n3693) & (n_n3642) & (n_n3641) & (x14770x)));
	assign n_n5330 = (((i_7_) & (!i_8_) & (!i_6_) & (x19x) & (n_n464)));
	assign n_n524 = (((i_7_) & (!i_8_) & (!i_6_)));
	assign n_n5331 = (((!i_9_) & (n_n524) & (n_n464) & (n_n65)));
	assign x14796x = (((!n_n5059) & (!n_n5018) & (!x371x) & (!x97x) & (x14793x)) + ((!n_n5059) & (!n_n5018) & (!x371x) & (x97x) & (!x14793x)) + ((!n_n5059) & (!n_n5018) & (!x371x) & (x97x) & (x14793x)) + ((!n_n5059) & (!n_n5018) & (x371x) & (!x97x) & (!x14793x)) + ((!n_n5059) & (!n_n5018) & (x371x) & (!x97x) & (x14793x)) + ((!n_n5059) & (!n_n5018) & (x371x) & (x97x) & (!x14793x)) + ((!n_n5059) & (!n_n5018) & (x371x) & (x97x) & (x14793x)) + ((!n_n5059) & (n_n5018) & (!x371x) & (!x97x) & (!x14793x)) + ((!n_n5059) & (n_n5018) & (!x371x) & (!x97x) & (x14793x)) + ((!n_n5059) & (n_n5018) & (!x371x) & (x97x) & (!x14793x)) + ((!n_n5059) & (n_n5018) & (!x371x) & (x97x) & (x14793x)) + ((!n_n5059) & (n_n5018) & (x371x) & (!x97x) & (!x14793x)) + ((!n_n5059) & (n_n5018) & (x371x) & (!x97x) & (x14793x)) + ((!n_n5059) & (n_n5018) & (x371x) & (x97x) & (!x14793x)) + ((!n_n5059) & (n_n5018) & (x371x) & (x97x) & (x14793x)) + ((n_n5059) & (!n_n5018) & (!x371x) & (!x97x) & (!x14793x)) + ((n_n5059) & (!n_n5018) & (!x371x) & (!x97x) & (x14793x)) + ((n_n5059) & (!n_n5018) & (!x371x) & (x97x) & (!x14793x)) + ((n_n5059) & (!n_n5018) & (!x371x) & (x97x) & (x14793x)) + ((n_n5059) & (!n_n5018) & (x371x) & (!x97x) & (!x14793x)) + ((n_n5059) & (!n_n5018) & (x371x) & (!x97x) & (x14793x)) + ((n_n5059) & (!n_n5018) & (x371x) & (x97x) & (!x14793x)) + ((n_n5059) & (!n_n5018) & (x371x) & (x97x) & (x14793x)) + ((n_n5059) & (n_n5018) & (!x371x) & (!x97x) & (!x14793x)) + ((n_n5059) & (n_n5018) & (!x371x) & (!x97x) & (x14793x)) + ((n_n5059) & (n_n5018) & (!x371x) & (x97x) & (!x14793x)) + ((n_n5059) & (n_n5018) & (!x371x) & (x97x) & (x14793x)) + ((n_n5059) & (n_n5018) & (x371x) & (!x97x) & (!x14793x)) + ((n_n5059) & (n_n5018) & (x371x) & (!x97x) & (x14793x)) + ((n_n5059) & (n_n5018) & (x371x) & (x97x) & (!x14793x)) + ((n_n5059) & (n_n5018) & (x371x) & (x97x) & (x14793x)));
	assign x14797x = (((!x155x) & (!x143x) & (!x14785x) & (!x14790x) & (x14791x)) + ((!x155x) & (!x143x) & (!x14785x) & (x14790x) & (!x14791x)) + ((!x155x) & (!x143x) & (!x14785x) & (x14790x) & (x14791x)) + ((!x155x) & (!x143x) & (x14785x) & (!x14790x) & (!x14791x)) + ((!x155x) & (!x143x) & (x14785x) & (!x14790x) & (x14791x)) + ((!x155x) & (!x143x) & (x14785x) & (x14790x) & (!x14791x)) + ((!x155x) & (!x143x) & (x14785x) & (x14790x) & (x14791x)) + ((!x155x) & (x143x) & (!x14785x) & (!x14790x) & (!x14791x)) + ((!x155x) & (x143x) & (!x14785x) & (!x14790x) & (x14791x)) + ((!x155x) & (x143x) & (!x14785x) & (x14790x) & (!x14791x)) + ((!x155x) & (x143x) & (!x14785x) & (x14790x) & (x14791x)) + ((!x155x) & (x143x) & (x14785x) & (!x14790x) & (!x14791x)) + ((!x155x) & (x143x) & (x14785x) & (!x14790x) & (x14791x)) + ((!x155x) & (x143x) & (x14785x) & (x14790x) & (!x14791x)) + ((!x155x) & (x143x) & (x14785x) & (x14790x) & (x14791x)) + ((x155x) & (!x143x) & (!x14785x) & (!x14790x) & (!x14791x)) + ((x155x) & (!x143x) & (!x14785x) & (!x14790x) & (x14791x)) + ((x155x) & (!x143x) & (!x14785x) & (x14790x) & (!x14791x)) + ((x155x) & (!x143x) & (!x14785x) & (x14790x) & (x14791x)) + ((x155x) & (!x143x) & (x14785x) & (!x14790x) & (!x14791x)) + ((x155x) & (!x143x) & (x14785x) & (!x14790x) & (x14791x)) + ((x155x) & (!x143x) & (x14785x) & (x14790x) & (!x14791x)) + ((x155x) & (!x143x) & (x14785x) & (x14790x) & (x14791x)) + ((x155x) & (x143x) & (!x14785x) & (!x14790x) & (!x14791x)) + ((x155x) & (x143x) & (!x14785x) & (!x14790x) & (x14791x)) + ((x155x) & (x143x) & (!x14785x) & (x14790x) & (!x14791x)) + ((x155x) & (x143x) & (!x14785x) & (x14790x) & (x14791x)) + ((x155x) & (x143x) & (x14785x) & (!x14790x) & (!x14791x)) + ((x155x) & (x143x) & (x14785x) & (!x14790x) & (x14791x)) + ((x155x) & (x143x) & (x14785x) & (x14790x) & (!x14791x)) + ((x155x) & (x143x) & (x14785x) & (x14790x) & (x14791x)));
	assign x14829x = (((!x14807x) & (!x14803x) & (!x14804x) & (!x14825x) & (x14826x)) + ((!x14807x) & (!x14803x) & (!x14804x) & (x14825x) & (!x14826x)) + ((!x14807x) & (!x14803x) & (!x14804x) & (x14825x) & (x14826x)) + ((!x14807x) & (!x14803x) & (x14804x) & (!x14825x) & (!x14826x)) + ((!x14807x) & (!x14803x) & (x14804x) & (!x14825x) & (x14826x)) + ((!x14807x) & (!x14803x) & (x14804x) & (x14825x) & (!x14826x)) + ((!x14807x) & (!x14803x) & (x14804x) & (x14825x) & (x14826x)) + ((!x14807x) & (x14803x) & (!x14804x) & (!x14825x) & (!x14826x)) + ((!x14807x) & (x14803x) & (!x14804x) & (!x14825x) & (x14826x)) + ((!x14807x) & (x14803x) & (!x14804x) & (x14825x) & (!x14826x)) + ((!x14807x) & (x14803x) & (!x14804x) & (x14825x) & (x14826x)) + ((!x14807x) & (x14803x) & (x14804x) & (!x14825x) & (!x14826x)) + ((!x14807x) & (x14803x) & (x14804x) & (!x14825x) & (x14826x)) + ((!x14807x) & (x14803x) & (x14804x) & (x14825x) & (!x14826x)) + ((!x14807x) & (x14803x) & (x14804x) & (x14825x) & (x14826x)) + ((x14807x) & (!x14803x) & (!x14804x) & (!x14825x) & (!x14826x)) + ((x14807x) & (!x14803x) & (!x14804x) & (!x14825x) & (x14826x)) + ((x14807x) & (!x14803x) & (!x14804x) & (x14825x) & (!x14826x)) + ((x14807x) & (!x14803x) & (!x14804x) & (x14825x) & (x14826x)) + ((x14807x) & (!x14803x) & (x14804x) & (!x14825x) & (!x14826x)) + ((x14807x) & (!x14803x) & (x14804x) & (!x14825x) & (x14826x)) + ((x14807x) & (!x14803x) & (x14804x) & (x14825x) & (!x14826x)) + ((x14807x) & (!x14803x) & (x14804x) & (x14825x) & (x14826x)) + ((x14807x) & (x14803x) & (!x14804x) & (!x14825x) & (!x14826x)) + ((x14807x) & (x14803x) & (!x14804x) & (!x14825x) & (x14826x)) + ((x14807x) & (x14803x) & (!x14804x) & (x14825x) & (!x14826x)) + ((x14807x) & (x14803x) & (!x14804x) & (x14825x) & (x14826x)) + ((x14807x) & (x14803x) & (x14804x) & (!x14825x) & (!x14826x)) + ((x14807x) & (x14803x) & (x14804x) & (!x14825x) & (x14826x)) + ((x14807x) & (x14803x) & (x14804x) & (x14825x) & (!x14826x)) + ((x14807x) & (x14803x) & (x14804x) & (x14825x) & (x14826x)));
	assign x14828x = (((!x14813x) & (!x14814x) & (!x14820x) & (x14821x)) + ((!x14813x) & (!x14814x) & (x14820x) & (!x14821x)) + ((!x14813x) & (!x14814x) & (x14820x) & (x14821x)) + ((!x14813x) & (x14814x) & (!x14820x) & (!x14821x)) + ((!x14813x) & (x14814x) & (!x14820x) & (x14821x)) + ((!x14813x) & (x14814x) & (x14820x) & (!x14821x)) + ((!x14813x) & (x14814x) & (x14820x) & (x14821x)) + ((x14813x) & (!x14814x) & (!x14820x) & (!x14821x)) + ((x14813x) & (!x14814x) & (!x14820x) & (x14821x)) + ((x14813x) & (!x14814x) & (x14820x) & (!x14821x)) + ((x14813x) & (!x14814x) & (x14820x) & (x14821x)) + ((x14813x) & (x14814x) & (!x14820x) & (!x14821x)) + ((x14813x) & (x14814x) & (!x14820x) & (x14821x)) + ((x14813x) & (x14814x) & (x14820x) & (!x14821x)) + ((x14813x) & (x14814x) & (x14820x) & (x14821x)));
	assign n_n2449 = (((!x14796x) & (!x14797x) & (!x14829x) & (x14828x)) + ((!x14796x) & (!x14797x) & (x14829x) & (!x14828x)) + ((!x14796x) & (!x14797x) & (x14829x) & (x14828x)) + ((!x14796x) & (x14797x) & (!x14829x) & (!x14828x)) + ((!x14796x) & (x14797x) & (!x14829x) & (x14828x)) + ((!x14796x) & (x14797x) & (x14829x) & (!x14828x)) + ((!x14796x) & (x14797x) & (x14829x) & (x14828x)) + ((x14796x) & (!x14797x) & (!x14829x) & (!x14828x)) + ((x14796x) & (!x14797x) & (!x14829x) & (x14828x)) + ((x14796x) & (!x14797x) & (x14829x) & (!x14828x)) + ((x14796x) & (!x14797x) & (x14829x) & (x14828x)) + ((x14796x) & (x14797x) & (!x14829x) & (!x14828x)) + ((x14796x) & (x14797x) & (!x14829x) & (x14828x)) + ((x14796x) & (x14797x) & (x14829x) & (!x14828x)) + ((x14796x) & (x14797x) & (x14829x) & (x14828x)));
	assign n_n2548 = (((!n_n1217) & (!n_n4848) & (!n_n4842) & (!x14907x) & (x14904x)) + ((!n_n1217) & (!n_n4848) & (!n_n4842) & (x14907x) & (!x14904x)) + ((!n_n1217) & (!n_n4848) & (!n_n4842) & (x14907x) & (x14904x)) + ((!n_n1217) & (!n_n4848) & (n_n4842) & (!x14907x) & (!x14904x)) + ((!n_n1217) & (!n_n4848) & (n_n4842) & (!x14907x) & (x14904x)) + ((!n_n1217) & (!n_n4848) & (n_n4842) & (x14907x) & (!x14904x)) + ((!n_n1217) & (!n_n4848) & (n_n4842) & (x14907x) & (x14904x)) + ((!n_n1217) & (n_n4848) & (!n_n4842) & (!x14907x) & (!x14904x)) + ((!n_n1217) & (n_n4848) & (!n_n4842) & (!x14907x) & (x14904x)) + ((!n_n1217) & (n_n4848) & (!n_n4842) & (x14907x) & (!x14904x)) + ((!n_n1217) & (n_n4848) & (!n_n4842) & (x14907x) & (x14904x)) + ((!n_n1217) & (n_n4848) & (n_n4842) & (!x14907x) & (!x14904x)) + ((!n_n1217) & (n_n4848) & (n_n4842) & (!x14907x) & (x14904x)) + ((!n_n1217) & (n_n4848) & (n_n4842) & (x14907x) & (!x14904x)) + ((!n_n1217) & (n_n4848) & (n_n4842) & (x14907x) & (x14904x)) + ((n_n1217) & (!n_n4848) & (!n_n4842) & (!x14907x) & (!x14904x)) + ((n_n1217) & (!n_n4848) & (!n_n4842) & (!x14907x) & (x14904x)) + ((n_n1217) & (!n_n4848) & (!n_n4842) & (x14907x) & (!x14904x)) + ((n_n1217) & (!n_n4848) & (!n_n4842) & (x14907x) & (x14904x)) + ((n_n1217) & (!n_n4848) & (n_n4842) & (!x14907x) & (!x14904x)) + ((n_n1217) & (!n_n4848) & (n_n4842) & (!x14907x) & (x14904x)) + ((n_n1217) & (!n_n4848) & (n_n4842) & (x14907x) & (!x14904x)) + ((n_n1217) & (!n_n4848) & (n_n4842) & (x14907x) & (x14904x)) + ((n_n1217) & (n_n4848) & (!n_n4842) & (!x14907x) & (!x14904x)) + ((n_n1217) & (n_n4848) & (!n_n4842) & (!x14907x) & (x14904x)) + ((n_n1217) & (n_n4848) & (!n_n4842) & (x14907x) & (!x14904x)) + ((n_n1217) & (n_n4848) & (!n_n4842) & (x14907x) & (x14904x)) + ((n_n1217) & (n_n4848) & (n_n4842) & (!x14907x) & (!x14904x)) + ((n_n1217) & (n_n4848) & (n_n4842) & (!x14907x) & (x14904x)) + ((n_n1217) & (n_n4848) & (n_n4842) & (x14907x) & (!x14904x)) + ((n_n1217) & (n_n4848) & (n_n4842) & (x14907x) & (x14904x)));
	assign n_n2598 = (((!n_n3451) & (!x174x) & (!n_n4876) & (!n_n4874) & (x14908x)) + ((!n_n3451) & (!x174x) & (!n_n4876) & (n_n4874) & (!x14908x)) + ((!n_n3451) & (!x174x) & (!n_n4876) & (n_n4874) & (x14908x)) + ((!n_n3451) & (!x174x) & (n_n4876) & (!n_n4874) & (!x14908x)) + ((!n_n3451) & (!x174x) & (n_n4876) & (!n_n4874) & (x14908x)) + ((!n_n3451) & (!x174x) & (n_n4876) & (n_n4874) & (!x14908x)) + ((!n_n3451) & (!x174x) & (n_n4876) & (n_n4874) & (x14908x)) + ((!n_n3451) & (x174x) & (!n_n4876) & (!n_n4874) & (!x14908x)) + ((!n_n3451) & (x174x) & (!n_n4876) & (!n_n4874) & (x14908x)) + ((!n_n3451) & (x174x) & (!n_n4876) & (n_n4874) & (!x14908x)) + ((!n_n3451) & (x174x) & (!n_n4876) & (n_n4874) & (x14908x)) + ((!n_n3451) & (x174x) & (n_n4876) & (!n_n4874) & (!x14908x)) + ((!n_n3451) & (x174x) & (n_n4876) & (!n_n4874) & (x14908x)) + ((!n_n3451) & (x174x) & (n_n4876) & (n_n4874) & (!x14908x)) + ((!n_n3451) & (x174x) & (n_n4876) & (n_n4874) & (x14908x)) + ((n_n3451) & (!x174x) & (!n_n4876) & (!n_n4874) & (!x14908x)) + ((n_n3451) & (!x174x) & (!n_n4876) & (!n_n4874) & (x14908x)) + ((n_n3451) & (!x174x) & (!n_n4876) & (n_n4874) & (!x14908x)) + ((n_n3451) & (!x174x) & (!n_n4876) & (n_n4874) & (x14908x)) + ((n_n3451) & (!x174x) & (n_n4876) & (!n_n4874) & (!x14908x)) + ((n_n3451) & (!x174x) & (n_n4876) & (!n_n4874) & (x14908x)) + ((n_n3451) & (!x174x) & (n_n4876) & (n_n4874) & (!x14908x)) + ((n_n3451) & (!x174x) & (n_n4876) & (n_n4874) & (x14908x)) + ((n_n3451) & (x174x) & (!n_n4876) & (!n_n4874) & (!x14908x)) + ((n_n3451) & (x174x) & (!n_n4876) & (!n_n4874) & (x14908x)) + ((n_n3451) & (x174x) & (!n_n4876) & (n_n4874) & (!x14908x)) + ((n_n3451) & (x174x) & (!n_n4876) & (n_n4874) & (x14908x)) + ((n_n3451) & (x174x) & (n_n4876) & (!n_n4874) & (!x14908x)) + ((n_n3451) & (x174x) & (n_n4876) & (!n_n4874) & (x14908x)) + ((n_n3451) & (x174x) & (n_n4876) & (n_n4874) & (!x14908x)) + ((n_n3451) & (x174x) & (n_n4876) & (n_n4874) & (x14908x)));
	assign n_n2597 = (((!n_n3450) & (!n_n4894) & (!n_n4889) & (!x12179x) & (x49x)) + ((!n_n3450) & (!n_n4894) & (!n_n4889) & (x12179x) & (!x49x)) + ((!n_n3450) & (!n_n4894) & (!n_n4889) & (x12179x) & (x49x)) + ((!n_n3450) & (!n_n4894) & (n_n4889) & (!x12179x) & (!x49x)) + ((!n_n3450) & (!n_n4894) & (n_n4889) & (!x12179x) & (x49x)) + ((!n_n3450) & (!n_n4894) & (n_n4889) & (x12179x) & (!x49x)) + ((!n_n3450) & (!n_n4894) & (n_n4889) & (x12179x) & (x49x)) + ((!n_n3450) & (n_n4894) & (!n_n4889) & (!x12179x) & (!x49x)) + ((!n_n3450) & (n_n4894) & (!n_n4889) & (!x12179x) & (x49x)) + ((!n_n3450) & (n_n4894) & (!n_n4889) & (x12179x) & (!x49x)) + ((!n_n3450) & (n_n4894) & (!n_n4889) & (x12179x) & (x49x)) + ((!n_n3450) & (n_n4894) & (n_n4889) & (!x12179x) & (!x49x)) + ((!n_n3450) & (n_n4894) & (n_n4889) & (!x12179x) & (x49x)) + ((!n_n3450) & (n_n4894) & (n_n4889) & (x12179x) & (!x49x)) + ((!n_n3450) & (n_n4894) & (n_n4889) & (x12179x) & (x49x)) + ((n_n3450) & (!n_n4894) & (!n_n4889) & (!x12179x) & (!x49x)) + ((n_n3450) & (!n_n4894) & (!n_n4889) & (!x12179x) & (x49x)) + ((n_n3450) & (!n_n4894) & (!n_n4889) & (x12179x) & (!x49x)) + ((n_n3450) & (!n_n4894) & (!n_n4889) & (x12179x) & (x49x)) + ((n_n3450) & (!n_n4894) & (n_n4889) & (!x12179x) & (!x49x)) + ((n_n3450) & (!n_n4894) & (n_n4889) & (!x12179x) & (x49x)) + ((n_n3450) & (!n_n4894) & (n_n4889) & (x12179x) & (!x49x)) + ((n_n3450) & (!n_n4894) & (n_n4889) & (x12179x) & (x49x)) + ((n_n3450) & (n_n4894) & (!n_n4889) & (!x12179x) & (!x49x)) + ((n_n3450) & (n_n4894) & (!n_n4889) & (!x12179x) & (x49x)) + ((n_n3450) & (n_n4894) & (!n_n4889) & (x12179x) & (!x49x)) + ((n_n3450) & (n_n4894) & (!n_n4889) & (x12179x) & (x49x)) + ((n_n3450) & (n_n4894) & (n_n4889) & (!x12179x) & (!x49x)) + ((n_n3450) & (n_n4894) & (n_n4889) & (!x12179x) & (x49x)) + ((n_n3450) & (n_n4894) & (n_n4889) & (x12179x) & (!x49x)) + ((n_n3450) & (n_n4894) & (n_n4889) & (x12179x) & (x49x)));
	assign n_n2549 = (((!x14927x) & (!x14918x) & (!x14919x) & (x14926x)) + ((!x14927x) & (!x14918x) & (x14919x) & (!x14926x)) + ((!x14927x) & (!x14918x) & (x14919x) & (x14926x)) + ((!x14927x) & (x14918x) & (!x14919x) & (!x14926x)) + ((!x14927x) & (x14918x) & (!x14919x) & (x14926x)) + ((!x14927x) & (x14918x) & (x14919x) & (!x14926x)) + ((!x14927x) & (x14918x) & (x14919x) & (x14926x)) + ((x14927x) & (!x14918x) & (!x14919x) & (!x14926x)) + ((x14927x) & (!x14918x) & (!x14919x) & (x14926x)) + ((x14927x) & (!x14918x) & (x14919x) & (!x14926x)) + ((x14927x) & (!x14918x) & (x14919x) & (x14926x)) + ((x14927x) & (x14918x) & (!x14919x) & (!x14926x)) + ((x14927x) & (x14918x) & (!x14919x) & (x14926x)) + ((x14927x) & (x14918x) & (x14919x) & (!x14926x)) + ((x14927x) & (x14918x) & (x14919x) & (x14926x)));
	assign x14933x = (((!n_n4862) & (!n_n4870) & (!n_n4872) & (!n_n4867) & (x14932x)) + ((!n_n4862) & (!n_n4870) & (!n_n4872) & (n_n4867) & (!x14932x)) + ((!n_n4862) & (!n_n4870) & (!n_n4872) & (n_n4867) & (x14932x)) + ((!n_n4862) & (!n_n4870) & (n_n4872) & (!n_n4867) & (!x14932x)) + ((!n_n4862) & (!n_n4870) & (n_n4872) & (!n_n4867) & (x14932x)) + ((!n_n4862) & (!n_n4870) & (n_n4872) & (n_n4867) & (!x14932x)) + ((!n_n4862) & (!n_n4870) & (n_n4872) & (n_n4867) & (x14932x)) + ((!n_n4862) & (n_n4870) & (!n_n4872) & (!n_n4867) & (!x14932x)) + ((!n_n4862) & (n_n4870) & (!n_n4872) & (!n_n4867) & (x14932x)) + ((!n_n4862) & (n_n4870) & (!n_n4872) & (n_n4867) & (!x14932x)) + ((!n_n4862) & (n_n4870) & (!n_n4872) & (n_n4867) & (x14932x)) + ((!n_n4862) & (n_n4870) & (n_n4872) & (!n_n4867) & (!x14932x)) + ((!n_n4862) & (n_n4870) & (n_n4872) & (!n_n4867) & (x14932x)) + ((!n_n4862) & (n_n4870) & (n_n4872) & (n_n4867) & (!x14932x)) + ((!n_n4862) & (n_n4870) & (n_n4872) & (n_n4867) & (x14932x)) + ((n_n4862) & (!n_n4870) & (!n_n4872) & (!n_n4867) & (!x14932x)) + ((n_n4862) & (!n_n4870) & (!n_n4872) & (!n_n4867) & (x14932x)) + ((n_n4862) & (!n_n4870) & (!n_n4872) & (n_n4867) & (!x14932x)) + ((n_n4862) & (!n_n4870) & (!n_n4872) & (n_n4867) & (x14932x)) + ((n_n4862) & (!n_n4870) & (n_n4872) & (!n_n4867) & (!x14932x)) + ((n_n4862) & (!n_n4870) & (n_n4872) & (!n_n4867) & (x14932x)) + ((n_n4862) & (!n_n4870) & (n_n4872) & (n_n4867) & (!x14932x)) + ((n_n4862) & (!n_n4870) & (n_n4872) & (n_n4867) & (x14932x)) + ((n_n4862) & (n_n4870) & (!n_n4872) & (!n_n4867) & (!x14932x)) + ((n_n4862) & (n_n4870) & (!n_n4872) & (!n_n4867) & (x14932x)) + ((n_n4862) & (n_n4870) & (!n_n4872) & (n_n4867) & (!x14932x)) + ((n_n4862) & (n_n4870) & (!n_n4872) & (n_n4867) & (x14932x)) + ((n_n4862) & (n_n4870) & (n_n4872) & (!n_n4867) & (!x14932x)) + ((n_n4862) & (n_n4870) & (n_n4872) & (!n_n4867) & (x14932x)) + ((n_n4862) & (n_n4870) & (n_n4872) & (n_n4867) & (!x14932x)) + ((n_n4862) & (n_n4870) & (n_n4872) & (n_n4867) & (x14932x)));
	assign n_n2589 = (((!n_n4987) & (!n_n4993) & (!n_n1576) & (!x134x) & (x252x)) + ((!n_n4987) & (!n_n4993) & (!n_n1576) & (x134x) & (!x252x)) + ((!n_n4987) & (!n_n4993) & (!n_n1576) & (x134x) & (x252x)) + ((!n_n4987) & (!n_n4993) & (n_n1576) & (!x134x) & (!x252x)) + ((!n_n4987) & (!n_n4993) & (n_n1576) & (!x134x) & (x252x)) + ((!n_n4987) & (!n_n4993) & (n_n1576) & (x134x) & (!x252x)) + ((!n_n4987) & (!n_n4993) & (n_n1576) & (x134x) & (x252x)) + ((!n_n4987) & (n_n4993) & (!n_n1576) & (!x134x) & (!x252x)) + ((!n_n4987) & (n_n4993) & (!n_n1576) & (!x134x) & (x252x)) + ((!n_n4987) & (n_n4993) & (!n_n1576) & (x134x) & (!x252x)) + ((!n_n4987) & (n_n4993) & (!n_n1576) & (x134x) & (x252x)) + ((!n_n4987) & (n_n4993) & (n_n1576) & (!x134x) & (!x252x)) + ((!n_n4987) & (n_n4993) & (n_n1576) & (!x134x) & (x252x)) + ((!n_n4987) & (n_n4993) & (n_n1576) & (x134x) & (!x252x)) + ((!n_n4987) & (n_n4993) & (n_n1576) & (x134x) & (x252x)) + ((n_n4987) & (!n_n4993) & (!n_n1576) & (!x134x) & (!x252x)) + ((n_n4987) & (!n_n4993) & (!n_n1576) & (!x134x) & (x252x)) + ((n_n4987) & (!n_n4993) & (!n_n1576) & (x134x) & (!x252x)) + ((n_n4987) & (!n_n4993) & (!n_n1576) & (x134x) & (x252x)) + ((n_n4987) & (!n_n4993) & (n_n1576) & (!x134x) & (!x252x)) + ((n_n4987) & (!n_n4993) & (n_n1576) & (!x134x) & (x252x)) + ((n_n4987) & (!n_n4993) & (n_n1576) & (x134x) & (!x252x)) + ((n_n4987) & (!n_n4993) & (n_n1576) & (x134x) & (x252x)) + ((n_n4987) & (n_n4993) & (!n_n1576) & (!x134x) & (!x252x)) + ((n_n4987) & (n_n4993) & (!n_n1576) & (!x134x) & (x252x)) + ((n_n4987) & (n_n4993) & (!n_n1576) & (x134x) & (!x252x)) + ((n_n4987) & (n_n4993) & (!n_n1576) & (x134x) & (x252x)) + ((n_n4987) & (n_n4993) & (n_n1576) & (!x134x) & (!x252x)) + ((n_n4987) & (n_n4993) & (n_n1576) & (!x134x) & (x252x)) + ((n_n4987) & (n_n4993) & (n_n1576) & (x134x) & (!x252x)) + ((n_n4987) & (n_n4993) & (n_n1576) & (x134x) & (x252x)));
	assign n_n2588 = (((!n_n5000) & (!x136x) & (!x247x) & (!x393x) & (x14940x)) + ((!n_n5000) & (!x136x) & (!x247x) & (x393x) & (!x14940x)) + ((!n_n5000) & (!x136x) & (!x247x) & (x393x) & (x14940x)) + ((!n_n5000) & (!x136x) & (x247x) & (!x393x) & (!x14940x)) + ((!n_n5000) & (!x136x) & (x247x) & (!x393x) & (x14940x)) + ((!n_n5000) & (!x136x) & (x247x) & (x393x) & (!x14940x)) + ((!n_n5000) & (!x136x) & (x247x) & (x393x) & (x14940x)) + ((!n_n5000) & (x136x) & (!x247x) & (!x393x) & (!x14940x)) + ((!n_n5000) & (x136x) & (!x247x) & (!x393x) & (x14940x)) + ((!n_n5000) & (x136x) & (!x247x) & (x393x) & (!x14940x)) + ((!n_n5000) & (x136x) & (!x247x) & (x393x) & (x14940x)) + ((!n_n5000) & (x136x) & (x247x) & (!x393x) & (!x14940x)) + ((!n_n5000) & (x136x) & (x247x) & (!x393x) & (x14940x)) + ((!n_n5000) & (x136x) & (x247x) & (x393x) & (!x14940x)) + ((!n_n5000) & (x136x) & (x247x) & (x393x) & (x14940x)) + ((n_n5000) & (!x136x) & (!x247x) & (!x393x) & (!x14940x)) + ((n_n5000) & (!x136x) & (!x247x) & (!x393x) & (x14940x)) + ((n_n5000) & (!x136x) & (!x247x) & (x393x) & (!x14940x)) + ((n_n5000) & (!x136x) & (!x247x) & (x393x) & (x14940x)) + ((n_n5000) & (!x136x) & (x247x) & (!x393x) & (!x14940x)) + ((n_n5000) & (!x136x) & (x247x) & (!x393x) & (x14940x)) + ((n_n5000) & (!x136x) & (x247x) & (x393x) & (!x14940x)) + ((n_n5000) & (!x136x) & (x247x) & (x393x) & (x14940x)) + ((n_n5000) & (x136x) & (!x247x) & (!x393x) & (!x14940x)) + ((n_n5000) & (x136x) & (!x247x) & (!x393x) & (x14940x)) + ((n_n5000) & (x136x) & (!x247x) & (x393x) & (!x14940x)) + ((n_n5000) & (x136x) & (!x247x) & (x393x) & (x14940x)) + ((n_n5000) & (x136x) & (x247x) & (!x393x) & (!x14940x)) + ((n_n5000) & (x136x) & (x247x) & (!x393x) & (x14940x)) + ((n_n5000) & (x136x) & (x247x) & (x393x) & (!x14940x)) + ((n_n5000) & (x136x) & (x247x) & (x393x) & (x14940x)));
	assign n_n2546 = (((!x14960x) & (!x14948x) & (!x14949x) & (n_n2596)) + ((!x14960x) & (!x14948x) & (x14949x) & (!n_n2596)) + ((!x14960x) & (!x14948x) & (x14949x) & (n_n2596)) + ((!x14960x) & (x14948x) & (!x14949x) & (!n_n2596)) + ((!x14960x) & (x14948x) & (!x14949x) & (n_n2596)) + ((!x14960x) & (x14948x) & (x14949x) & (!n_n2596)) + ((!x14960x) & (x14948x) & (x14949x) & (n_n2596)) + ((x14960x) & (!x14948x) & (!x14949x) & (!n_n2596)) + ((x14960x) & (!x14948x) & (!x14949x) & (n_n2596)) + ((x14960x) & (!x14948x) & (x14949x) & (!n_n2596)) + ((x14960x) & (!x14948x) & (x14949x) & (n_n2596)) + ((x14960x) & (x14948x) & (!x14949x) & (!n_n2596)) + ((x14960x) & (x14948x) & (!x14949x) & (n_n2596)) + ((x14960x) & (x14948x) & (x14949x) & (!n_n2596)) + ((x14960x) & (x14948x) & (x14949x) & (n_n2596)));
	assign n_n2545 = (((!n_n4939) & (!x382x) & (!x14974x) & (!n_n2591) & (x14970x)) + ((!n_n4939) & (!x382x) & (!x14974x) & (n_n2591) & (!x14970x)) + ((!n_n4939) & (!x382x) & (!x14974x) & (n_n2591) & (x14970x)) + ((!n_n4939) & (!x382x) & (x14974x) & (!n_n2591) & (!x14970x)) + ((!n_n4939) & (!x382x) & (x14974x) & (!n_n2591) & (x14970x)) + ((!n_n4939) & (!x382x) & (x14974x) & (n_n2591) & (!x14970x)) + ((!n_n4939) & (!x382x) & (x14974x) & (n_n2591) & (x14970x)) + ((!n_n4939) & (x382x) & (!x14974x) & (!n_n2591) & (!x14970x)) + ((!n_n4939) & (x382x) & (!x14974x) & (!n_n2591) & (x14970x)) + ((!n_n4939) & (x382x) & (!x14974x) & (n_n2591) & (!x14970x)) + ((!n_n4939) & (x382x) & (!x14974x) & (n_n2591) & (x14970x)) + ((!n_n4939) & (x382x) & (x14974x) & (!n_n2591) & (!x14970x)) + ((!n_n4939) & (x382x) & (x14974x) & (!n_n2591) & (x14970x)) + ((!n_n4939) & (x382x) & (x14974x) & (n_n2591) & (!x14970x)) + ((!n_n4939) & (x382x) & (x14974x) & (n_n2591) & (x14970x)) + ((n_n4939) & (!x382x) & (!x14974x) & (!n_n2591) & (!x14970x)) + ((n_n4939) & (!x382x) & (!x14974x) & (!n_n2591) & (x14970x)) + ((n_n4939) & (!x382x) & (!x14974x) & (n_n2591) & (!x14970x)) + ((n_n4939) & (!x382x) & (!x14974x) & (n_n2591) & (x14970x)) + ((n_n4939) & (!x382x) & (x14974x) & (!n_n2591) & (!x14970x)) + ((n_n4939) & (!x382x) & (x14974x) & (!n_n2591) & (x14970x)) + ((n_n4939) & (!x382x) & (x14974x) & (n_n2591) & (!x14970x)) + ((n_n4939) & (!x382x) & (x14974x) & (n_n2591) & (x14970x)) + ((n_n4939) & (x382x) & (!x14974x) & (!n_n2591) & (!x14970x)) + ((n_n4939) & (x382x) & (!x14974x) & (!n_n2591) & (x14970x)) + ((n_n4939) & (x382x) & (!x14974x) & (n_n2591) & (!x14970x)) + ((n_n4939) & (x382x) & (!x14974x) & (n_n2591) & (x14970x)) + ((n_n4939) & (x382x) & (x14974x) & (!n_n2591) & (!x14970x)) + ((n_n4939) & (x382x) & (x14974x) & (!n_n2591) & (x14970x)) + ((n_n4939) & (x382x) & (x14974x) & (n_n2591) & (!x14970x)) + ((n_n4939) & (x382x) & (x14974x) & (n_n2591) & (x14970x)));
	assign x14979x = (((!n_n4978) & (!x29x) & (!n_n4965) & (!x68x) & (x228x)) + ((!n_n4978) & (!x29x) & (!n_n4965) & (x68x) & (!x228x)) + ((!n_n4978) & (!x29x) & (!n_n4965) & (x68x) & (x228x)) + ((!n_n4978) & (!x29x) & (n_n4965) & (!x68x) & (!x228x)) + ((!n_n4978) & (!x29x) & (n_n4965) & (!x68x) & (x228x)) + ((!n_n4978) & (!x29x) & (n_n4965) & (x68x) & (!x228x)) + ((!n_n4978) & (!x29x) & (n_n4965) & (x68x) & (x228x)) + ((!n_n4978) & (x29x) & (!n_n4965) & (!x68x) & (!x228x)) + ((!n_n4978) & (x29x) & (!n_n4965) & (!x68x) & (x228x)) + ((!n_n4978) & (x29x) & (!n_n4965) & (x68x) & (!x228x)) + ((!n_n4978) & (x29x) & (!n_n4965) & (x68x) & (x228x)) + ((!n_n4978) & (x29x) & (n_n4965) & (!x68x) & (!x228x)) + ((!n_n4978) & (x29x) & (n_n4965) & (!x68x) & (x228x)) + ((!n_n4978) & (x29x) & (n_n4965) & (x68x) & (!x228x)) + ((!n_n4978) & (x29x) & (n_n4965) & (x68x) & (x228x)) + ((n_n4978) & (!x29x) & (!n_n4965) & (!x68x) & (!x228x)) + ((n_n4978) & (!x29x) & (!n_n4965) & (!x68x) & (x228x)) + ((n_n4978) & (!x29x) & (!n_n4965) & (x68x) & (!x228x)) + ((n_n4978) & (!x29x) & (!n_n4965) & (x68x) & (x228x)) + ((n_n4978) & (!x29x) & (n_n4965) & (!x68x) & (!x228x)) + ((n_n4978) & (!x29x) & (n_n4965) & (!x68x) & (x228x)) + ((n_n4978) & (!x29x) & (n_n4965) & (x68x) & (!x228x)) + ((n_n4978) & (!x29x) & (n_n4965) & (x68x) & (x228x)) + ((n_n4978) & (x29x) & (!n_n4965) & (!x68x) & (!x228x)) + ((n_n4978) & (x29x) & (!n_n4965) & (!x68x) & (x228x)) + ((n_n4978) & (x29x) & (!n_n4965) & (x68x) & (!x228x)) + ((n_n4978) & (x29x) & (!n_n4965) & (x68x) & (x228x)) + ((n_n4978) & (x29x) & (n_n4965) & (!x68x) & (!x228x)) + ((n_n4978) & (x29x) & (n_n4965) & (!x68x) & (x228x)) + ((n_n4978) & (x29x) & (n_n4965) & (x68x) & (!x228x)) + ((n_n4978) & (x29x) & (n_n4965) & (x68x) & (x228x)));
	assign n_n2608 = (((!x21x) & (!x483x) & (!x20x) & (!x47x) & (x14986x)) + ((!x21x) & (!x483x) & (!x20x) & (x47x) & (!x14986x)) + ((!x21x) & (!x483x) & (!x20x) & (x47x) & (x14986x)) + ((!x21x) & (!x483x) & (x20x) & (!x47x) & (x14986x)) + ((!x21x) & (!x483x) & (x20x) & (x47x) & (!x14986x)) + ((!x21x) & (!x483x) & (x20x) & (x47x) & (x14986x)) + ((!x21x) & (x483x) & (!x20x) & (!x47x) & (x14986x)) + ((!x21x) & (x483x) & (!x20x) & (x47x) & (!x14986x)) + ((!x21x) & (x483x) & (!x20x) & (x47x) & (x14986x)) + ((!x21x) & (x483x) & (x20x) & (!x47x) & (!x14986x)) + ((!x21x) & (x483x) & (x20x) & (!x47x) & (x14986x)) + ((!x21x) & (x483x) & (x20x) & (x47x) & (!x14986x)) + ((!x21x) & (x483x) & (x20x) & (x47x) & (x14986x)) + ((x21x) & (!x483x) & (!x20x) & (!x47x) & (x14986x)) + ((x21x) & (!x483x) & (!x20x) & (x47x) & (!x14986x)) + ((x21x) & (!x483x) & (!x20x) & (x47x) & (x14986x)) + ((x21x) & (!x483x) & (x20x) & (!x47x) & (x14986x)) + ((x21x) & (!x483x) & (x20x) & (x47x) & (!x14986x)) + ((x21x) & (!x483x) & (x20x) & (x47x) & (x14986x)) + ((x21x) & (x483x) & (!x20x) & (!x47x) & (!x14986x)) + ((x21x) & (x483x) & (!x20x) & (!x47x) & (x14986x)) + ((x21x) & (x483x) & (!x20x) & (x47x) & (!x14986x)) + ((x21x) & (x483x) & (!x20x) & (x47x) & (x14986x)) + ((x21x) & (x483x) & (x20x) & (!x47x) & (!x14986x)) + ((x21x) & (x483x) & (x20x) & (!x47x) & (x14986x)) + ((x21x) & (x483x) & (x20x) & (x47x) & (!x14986x)) + ((x21x) & (x483x) & (x20x) & (x47x) & (x14986x)));
	assign n_n2607 = (((!n_n4761) & (!n_n4764) & (!n_n4763) & (!x164x) & (!x22092x)) + ((!n_n4761) & (!n_n4764) & (!n_n4763) & (x164x) & (!x22092x)) + ((!n_n4761) & (!n_n4764) & (!n_n4763) & (x164x) & (x22092x)) + ((!n_n4761) & (!n_n4764) & (n_n4763) & (!x164x) & (!x22092x)) + ((!n_n4761) & (!n_n4764) & (n_n4763) & (!x164x) & (x22092x)) + ((!n_n4761) & (!n_n4764) & (n_n4763) & (x164x) & (!x22092x)) + ((!n_n4761) & (!n_n4764) & (n_n4763) & (x164x) & (x22092x)) + ((!n_n4761) & (n_n4764) & (!n_n4763) & (!x164x) & (!x22092x)) + ((!n_n4761) & (n_n4764) & (!n_n4763) & (!x164x) & (x22092x)) + ((!n_n4761) & (n_n4764) & (!n_n4763) & (x164x) & (!x22092x)) + ((!n_n4761) & (n_n4764) & (!n_n4763) & (x164x) & (x22092x)) + ((!n_n4761) & (n_n4764) & (n_n4763) & (!x164x) & (!x22092x)) + ((!n_n4761) & (n_n4764) & (n_n4763) & (!x164x) & (x22092x)) + ((!n_n4761) & (n_n4764) & (n_n4763) & (x164x) & (!x22092x)) + ((!n_n4761) & (n_n4764) & (n_n4763) & (x164x) & (x22092x)) + ((n_n4761) & (!n_n4764) & (!n_n4763) & (!x164x) & (!x22092x)) + ((n_n4761) & (!n_n4764) & (!n_n4763) & (!x164x) & (x22092x)) + ((n_n4761) & (!n_n4764) & (!n_n4763) & (x164x) & (!x22092x)) + ((n_n4761) & (!n_n4764) & (!n_n4763) & (x164x) & (x22092x)) + ((n_n4761) & (!n_n4764) & (n_n4763) & (!x164x) & (!x22092x)) + ((n_n4761) & (!n_n4764) & (n_n4763) & (!x164x) & (x22092x)) + ((n_n4761) & (!n_n4764) & (n_n4763) & (x164x) & (!x22092x)) + ((n_n4761) & (!n_n4764) & (n_n4763) & (x164x) & (x22092x)) + ((n_n4761) & (n_n4764) & (!n_n4763) & (!x164x) & (!x22092x)) + ((n_n4761) & (n_n4764) & (!n_n4763) & (!x164x) & (x22092x)) + ((n_n4761) & (n_n4764) & (!n_n4763) & (x164x) & (!x22092x)) + ((n_n4761) & (n_n4764) & (!n_n4763) & (x164x) & (x22092x)) + ((n_n4761) & (n_n4764) & (n_n4763) & (!x164x) & (!x22092x)) + ((n_n4761) & (n_n4764) & (n_n4763) & (!x164x) & (x22092x)) + ((n_n4761) & (n_n4764) & (n_n4763) & (x164x) & (!x22092x)) + ((n_n4761) & (n_n4764) & (n_n4763) & (x164x) & (x22092x)));
	assign x15021x = (((!n_n4776) & (!n_n4774) & (!n_n4781) & (n_n4777)) + ((!n_n4776) & (!n_n4774) & (n_n4781) & (!n_n4777)) + ((!n_n4776) & (!n_n4774) & (n_n4781) & (n_n4777)) + ((!n_n4776) & (n_n4774) & (!n_n4781) & (!n_n4777)) + ((!n_n4776) & (n_n4774) & (!n_n4781) & (n_n4777)) + ((!n_n4776) & (n_n4774) & (n_n4781) & (!n_n4777)) + ((!n_n4776) & (n_n4774) & (n_n4781) & (n_n4777)) + ((n_n4776) & (!n_n4774) & (!n_n4781) & (!n_n4777)) + ((n_n4776) & (!n_n4774) & (!n_n4781) & (n_n4777)) + ((n_n4776) & (!n_n4774) & (n_n4781) & (!n_n4777)) + ((n_n4776) & (!n_n4774) & (n_n4781) & (n_n4777)) + ((n_n4776) & (n_n4774) & (!n_n4781) & (!n_n4777)) + ((n_n4776) & (n_n4774) & (!n_n4781) & (n_n4777)) + ((n_n4776) & (n_n4774) & (n_n4781) & (!n_n4777)) + ((n_n4776) & (n_n4774) & (n_n4781) & (n_n4777)));
	assign x15022x = (((!n_n4779) & (!n_n4780) & (!n_n4778) & (!n_n4773) & (n_n4775)) + ((!n_n4779) & (!n_n4780) & (!n_n4778) & (n_n4773) & (!n_n4775)) + ((!n_n4779) & (!n_n4780) & (!n_n4778) & (n_n4773) & (n_n4775)) + ((!n_n4779) & (!n_n4780) & (n_n4778) & (!n_n4773) & (!n_n4775)) + ((!n_n4779) & (!n_n4780) & (n_n4778) & (!n_n4773) & (n_n4775)) + ((!n_n4779) & (!n_n4780) & (n_n4778) & (n_n4773) & (!n_n4775)) + ((!n_n4779) & (!n_n4780) & (n_n4778) & (n_n4773) & (n_n4775)) + ((!n_n4779) & (n_n4780) & (!n_n4778) & (!n_n4773) & (!n_n4775)) + ((!n_n4779) & (n_n4780) & (!n_n4778) & (!n_n4773) & (n_n4775)) + ((!n_n4779) & (n_n4780) & (!n_n4778) & (n_n4773) & (!n_n4775)) + ((!n_n4779) & (n_n4780) & (!n_n4778) & (n_n4773) & (n_n4775)) + ((!n_n4779) & (n_n4780) & (n_n4778) & (!n_n4773) & (!n_n4775)) + ((!n_n4779) & (n_n4780) & (n_n4778) & (!n_n4773) & (n_n4775)) + ((!n_n4779) & (n_n4780) & (n_n4778) & (n_n4773) & (!n_n4775)) + ((!n_n4779) & (n_n4780) & (n_n4778) & (n_n4773) & (n_n4775)) + ((n_n4779) & (!n_n4780) & (!n_n4778) & (!n_n4773) & (!n_n4775)) + ((n_n4779) & (!n_n4780) & (!n_n4778) & (!n_n4773) & (n_n4775)) + ((n_n4779) & (!n_n4780) & (!n_n4778) & (n_n4773) & (!n_n4775)) + ((n_n4779) & (!n_n4780) & (!n_n4778) & (n_n4773) & (n_n4775)) + ((n_n4779) & (!n_n4780) & (n_n4778) & (!n_n4773) & (!n_n4775)) + ((n_n4779) & (!n_n4780) & (n_n4778) & (!n_n4773) & (n_n4775)) + ((n_n4779) & (!n_n4780) & (n_n4778) & (n_n4773) & (!n_n4775)) + ((n_n4779) & (!n_n4780) & (n_n4778) & (n_n4773) & (n_n4775)) + ((n_n4779) & (n_n4780) & (!n_n4778) & (!n_n4773) & (!n_n4775)) + ((n_n4779) & (n_n4780) & (!n_n4778) & (!n_n4773) & (n_n4775)) + ((n_n4779) & (n_n4780) & (!n_n4778) & (n_n4773) & (!n_n4775)) + ((n_n4779) & (n_n4780) & (!n_n4778) & (n_n4773) & (n_n4775)) + ((n_n4779) & (n_n4780) & (n_n4778) & (!n_n4773) & (!n_n4775)) + ((n_n4779) & (n_n4780) & (n_n4778) & (!n_n4773) & (n_n4775)) + ((n_n4779) & (n_n4780) & (n_n4778) & (n_n4773) & (!n_n4775)) + ((n_n4779) & (n_n4780) & (n_n4778) & (n_n4773) & (n_n4775)));
	assign x15025x = (((!n_n2608) & (!n_n2607) & (!x15021x) & (x15022x)) + ((!n_n2608) & (!n_n2607) & (x15021x) & (!x15022x)) + ((!n_n2608) & (!n_n2607) & (x15021x) & (x15022x)) + ((!n_n2608) & (n_n2607) & (!x15021x) & (!x15022x)) + ((!n_n2608) & (n_n2607) & (!x15021x) & (x15022x)) + ((!n_n2608) & (n_n2607) & (x15021x) & (!x15022x)) + ((!n_n2608) & (n_n2607) & (x15021x) & (x15022x)) + ((n_n2608) & (!n_n2607) & (!x15021x) & (!x15022x)) + ((n_n2608) & (!n_n2607) & (!x15021x) & (x15022x)) + ((n_n2608) & (!n_n2607) & (x15021x) & (!x15022x)) + ((n_n2608) & (!n_n2607) & (x15021x) & (x15022x)) + ((n_n2608) & (n_n2607) & (!x15021x) & (!x15022x)) + ((n_n2608) & (n_n2607) & (!x15021x) & (x15022x)) + ((n_n2608) & (n_n2607) & (x15021x) & (!x15022x)) + ((n_n2608) & (n_n2607) & (x15021x) & (x15022x)));
	assign n_n2552 = (((!n_n2614) & (!x15002x) & (!x15003x) & (x15004x)) + ((!n_n2614) & (!x15002x) & (x15003x) & (!x15004x)) + ((!n_n2614) & (!x15002x) & (x15003x) & (x15004x)) + ((!n_n2614) & (x15002x) & (!x15003x) & (!x15004x)) + ((!n_n2614) & (x15002x) & (!x15003x) & (x15004x)) + ((!n_n2614) & (x15002x) & (x15003x) & (!x15004x)) + ((!n_n2614) & (x15002x) & (x15003x) & (x15004x)) + ((n_n2614) & (!x15002x) & (!x15003x) & (!x15004x)) + ((n_n2614) & (!x15002x) & (!x15003x) & (x15004x)) + ((n_n2614) & (!x15002x) & (x15003x) & (!x15004x)) + ((n_n2614) & (!x15002x) & (x15003x) & (x15004x)) + ((n_n2614) & (x15002x) & (!x15003x) & (!x15004x)) + ((n_n2614) & (x15002x) & (!x15003x) & (x15004x)) + ((n_n2614) & (x15002x) & (x15003x) & (!x15004x)) + ((n_n2614) & (x15002x) & (x15003x) & (x15004x)));
	assign n_n2551 = (((!n_n2611) & (!x15013x) & (!x15014x) & (x15015x)) + ((!n_n2611) & (!x15013x) & (x15014x) & (!x15015x)) + ((!n_n2611) & (!x15013x) & (x15014x) & (x15015x)) + ((!n_n2611) & (x15013x) & (!x15014x) & (!x15015x)) + ((!n_n2611) & (x15013x) & (!x15014x) & (x15015x)) + ((!n_n2611) & (x15013x) & (x15014x) & (!x15015x)) + ((!n_n2611) & (x15013x) & (x15014x) & (x15015x)) + ((n_n2611) & (!x15013x) & (!x15014x) & (!x15015x)) + ((n_n2611) & (!x15013x) & (!x15014x) & (x15015x)) + ((n_n2611) & (!x15013x) & (x15014x) & (!x15015x)) + ((n_n2611) & (!x15013x) & (x15014x) & (x15015x)) + ((n_n2611) & (x15013x) & (!x15014x) & (!x15015x)) + ((n_n2611) & (x15013x) & (!x15014x) & (x15015x)) + ((n_n2611) & (x15013x) & (x15014x) & (!x15015x)) + ((n_n2611) & (x15013x) & (x15014x) & (x15015x)));
	assign n_n2531 = (((!x15025x) & (!n_n2552) & (n_n2551)) + ((!x15025x) & (n_n2552) & (!n_n2551)) + ((!x15025x) & (n_n2552) & (n_n2551)) + ((x15025x) & (!n_n2552) & (!n_n2551)) + ((x15025x) & (!n_n2552) & (n_n2551)) + ((x15025x) & (n_n2552) & (!n_n2551)) + ((x15025x) & (n_n2552) & (n_n2551)));
	assign n_n2560 = (((!n_n2637) & (!x15033x) & (!x15034x) & (x15040x)) + ((!n_n2637) & (!x15033x) & (x15034x) & (!x15040x)) + ((!n_n2637) & (!x15033x) & (x15034x) & (x15040x)) + ((!n_n2637) & (x15033x) & (!x15034x) & (!x15040x)) + ((!n_n2637) & (x15033x) & (!x15034x) & (x15040x)) + ((!n_n2637) & (x15033x) & (x15034x) & (!x15040x)) + ((!n_n2637) & (x15033x) & (x15034x) & (x15040x)) + ((n_n2637) & (!x15033x) & (!x15034x) & (!x15040x)) + ((n_n2637) & (!x15033x) & (!x15034x) & (x15040x)) + ((n_n2637) & (!x15033x) & (x15034x) & (!x15040x)) + ((n_n2637) & (!x15033x) & (x15034x) & (x15040x)) + ((n_n2637) & (x15033x) & (!x15034x) & (!x15040x)) + ((n_n2637) & (x15033x) & (!x15034x) & (x15040x)) + ((n_n2637) & (x15033x) & (x15034x) & (!x15040x)) + ((n_n2637) & (x15033x) & (x15034x) & (x15040x)));
	assign n_n2559 = (((!n_n2634) & (!x15049x) & (!x15050x) & (x15055x)) + ((!n_n2634) & (!x15049x) & (x15050x) & (!x15055x)) + ((!n_n2634) & (!x15049x) & (x15050x) & (x15055x)) + ((!n_n2634) & (x15049x) & (!x15050x) & (!x15055x)) + ((!n_n2634) & (x15049x) & (!x15050x) & (x15055x)) + ((!n_n2634) & (x15049x) & (x15050x) & (!x15055x)) + ((!n_n2634) & (x15049x) & (x15050x) & (x15055x)) + ((n_n2634) & (!x15049x) & (!x15050x) & (!x15055x)) + ((n_n2634) & (!x15049x) & (!x15050x) & (x15055x)) + ((n_n2634) & (!x15049x) & (x15050x) & (!x15055x)) + ((n_n2634) & (!x15049x) & (x15050x) & (x15055x)) + ((n_n2634) & (x15049x) & (!x15050x) & (!x15055x)) + ((n_n2634) & (x15049x) & (!x15050x) & (x15055x)) + ((n_n2634) & (x15049x) & (x15050x) & (!x15055x)) + ((n_n2634) & (x15049x) & (x15050x) & (x15055x)));
	assign x15167x = (((!x156x) & (!n_n2640) & (!n_n2641) & (!x337x) & (x15164x)) + ((!x156x) & (!n_n2640) & (!n_n2641) & (x337x) & (!x15164x)) + ((!x156x) & (!n_n2640) & (!n_n2641) & (x337x) & (x15164x)) + ((!x156x) & (!n_n2640) & (n_n2641) & (!x337x) & (!x15164x)) + ((!x156x) & (!n_n2640) & (n_n2641) & (!x337x) & (x15164x)) + ((!x156x) & (!n_n2640) & (n_n2641) & (x337x) & (!x15164x)) + ((!x156x) & (!n_n2640) & (n_n2641) & (x337x) & (x15164x)) + ((!x156x) & (n_n2640) & (!n_n2641) & (!x337x) & (!x15164x)) + ((!x156x) & (n_n2640) & (!n_n2641) & (!x337x) & (x15164x)) + ((!x156x) & (n_n2640) & (!n_n2641) & (x337x) & (!x15164x)) + ((!x156x) & (n_n2640) & (!n_n2641) & (x337x) & (x15164x)) + ((!x156x) & (n_n2640) & (n_n2641) & (!x337x) & (!x15164x)) + ((!x156x) & (n_n2640) & (n_n2641) & (!x337x) & (x15164x)) + ((!x156x) & (n_n2640) & (n_n2641) & (x337x) & (!x15164x)) + ((!x156x) & (n_n2640) & (n_n2641) & (x337x) & (x15164x)) + ((x156x) & (!n_n2640) & (!n_n2641) & (!x337x) & (!x15164x)) + ((x156x) & (!n_n2640) & (!n_n2641) & (!x337x) & (x15164x)) + ((x156x) & (!n_n2640) & (!n_n2641) & (x337x) & (!x15164x)) + ((x156x) & (!n_n2640) & (!n_n2641) & (x337x) & (x15164x)) + ((x156x) & (!n_n2640) & (n_n2641) & (!x337x) & (!x15164x)) + ((x156x) & (!n_n2640) & (n_n2641) & (!x337x) & (x15164x)) + ((x156x) & (!n_n2640) & (n_n2641) & (x337x) & (!x15164x)) + ((x156x) & (!n_n2640) & (n_n2641) & (x337x) & (x15164x)) + ((x156x) & (n_n2640) & (!n_n2641) & (!x337x) & (!x15164x)) + ((x156x) & (n_n2640) & (!n_n2641) & (!x337x) & (x15164x)) + ((x156x) & (n_n2640) & (!n_n2641) & (x337x) & (!x15164x)) + ((x156x) & (n_n2640) & (!n_n2641) & (x337x) & (x15164x)) + ((x156x) & (n_n2640) & (n_n2641) & (!x337x) & (!x15164x)) + ((x156x) & (n_n2640) & (n_n2641) & (!x337x) & (x15164x)) + ((x156x) & (n_n2640) & (n_n2641) & (x337x) & (!x15164x)) + ((x156x) & (n_n2640) & (n_n2641) & (x337x) & (x15164x)));
	assign n_n2538 = (((!n_n2570) & (!x15221x) & (x15220x)) + ((!n_n2570) & (x15221x) & (!x15220x)) + ((!n_n2570) & (x15221x) & (x15220x)) + ((n_n2570) & (!x15221x) & (!x15220x)) + ((n_n2570) & (!x15221x) & (x15220x)) + ((n_n2570) & (x15221x) & (!x15220x)) + ((n_n2570) & (x15221x) & (x15220x)));
	assign n_n2539 = (((!x15269x) & (!x15270x) & (!x15278x) & (x15277x)) + ((!x15269x) & (!x15270x) & (x15278x) & (!x15277x)) + ((!x15269x) & (!x15270x) & (x15278x) & (x15277x)) + ((!x15269x) & (x15270x) & (!x15278x) & (!x15277x)) + ((!x15269x) & (x15270x) & (!x15278x) & (x15277x)) + ((!x15269x) & (x15270x) & (x15278x) & (!x15277x)) + ((!x15269x) & (x15270x) & (x15278x) & (x15277x)) + ((x15269x) & (!x15270x) & (!x15278x) & (!x15277x)) + ((x15269x) & (!x15270x) & (!x15278x) & (x15277x)) + ((x15269x) & (!x15270x) & (x15278x) & (!x15277x)) + ((x15269x) & (!x15270x) & (x15278x) & (x15277x)) + ((x15269x) & (x15270x) & (!x15278x) & (!x15277x)) + ((x15269x) & (x15270x) & (!x15278x) & (x15277x)) + ((x15269x) & (x15270x) & (x15278x) & (!x15277x)) + ((x15269x) & (x15270x) & (x15278x) & (x15277x)));
	assign n_n2576 = (((!n_n5167) & (!n_n5164) & (!n_n5162) & (!n_n5166) & (x15284x)) + ((!n_n5167) & (!n_n5164) & (!n_n5162) & (n_n5166) & (!x15284x)) + ((!n_n5167) & (!n_n5164) & (!n_n5162) & (n_n5166) & (x15284x)) + ((!n_n5167) & (!n_n5164) & (n_n5162) & (!n_n5166) & (!x15284x)) + ((!n_n5167) & (!n_n5164) & (n_n5162) & (!n_n5166) & (x15284x)) + ((!n_n5167) & (!n_n5164) & (n_n5162) & (n_n5166) & (!x15284x)) + ((!n_n5167) & (!n_n5164) & (n_n5162) & (n_n5166) & (x15284x)) + ((!n_n5167) & (n_n5164) & (!n_n5162) & (!n_n5166) & (!x15284x)) + ((!n_n5167) & (n_n5164) & (!n_n5162) & (!n_n5166) & (x15284x)) + ((!n_n5167) & (n_n5164) & (!n_n5162) & (n_n5166) & (!x15284x)) + ((!n_n5167) & (n_n5164) & (!n_n5162) & (n_n5166) & (x15284x)) + ((!n_n5167) & (n_n5164) & (n_n5162) & (!n_n5166) & (!x15284x)) + ((!n_n5167) & (n_n5164) & (n_n5162) & (!n_n5166) & (x15284x)) + ((!n_n5167) & (n_n5164) & (n_n5162) & (n_n5166) & (!x15284x)) + ((!n_n5167) & (n_n5164) & (n_n5162) & (n_n5166) & (x15284x)) + ((n_n5167) & (!n_n5164) & (!n_n5162) & (!n_n5166) & (!x15284x)) + ((n_n5167) & (!n_n5164) & (!n_n5162) & (!n_n5166) & (x15284x)) + ((n_n5167) & (!n_n5164) & (!n_n5162) & (n_n5166) & (!x15284x)) + ((n_n5167) & (!n_n5164) & (!n_n5162) & (n_n5166) & (x15284x)) + ((n_n5167) & (!n_n5164) & (n_n5162) & (!n_n5166) & (!x15284x)) + ((n_n5167) & (!n_n5164) & (n_n5162) & (!n_n5166) & (x15284x)) + ((n_n5167) & (!n_n5164) & (n_n5162) & (n_n5166) & (!x15284x)) + ((n_n5167) & (!n_n5164) & (n_n5162) & (n_n5166) & (x15284x)) + ((n_n5167) & (n_n5164) & (!n_n5162) & (!n_n5166) & (!x15284x)) + ((n_n5167) & (n_n5164) & (!n_n5162) & (!n_n5166) & (x15284x)) + ((n_n5167) & (n_n5164) & (!n_n5162) & (n_n5166) & (!x15284x)) + ((n_n5167) & (n_n5164) & (!n_n5162) & (n_n5166) & (x15284x)) + ((n_n5167) & (n_n5164) & (n_n5162) & (!n_n5166) & (!x15284x)) + ((n_n5167) & (n_n5164) & (n_n5162) & (!n_n5166) & (x15284x)) + ((n_n5167) & (n_n5164) & (n_n5162) & (n_n5166) & (!x15284x)) + ((n_n5167) & (n_n5164) & (n_n5162) & (n_n5166) & (x15284x)));
	assign n_n2577 = (((!n_n5149) & (!n_n5152) & (!n_n5153) & (!x407x) & (!x22204x)) + ((!n_n5149) & (!n_n5152) & (!n_n5153) & (x407x) & (!x22204x)) + ((!n_n5149) & (!n_n5152) & (!n_n5153) & (x407x) & (x22204x)) + ((!n_n5149) & (!n_n5152) & (n_n5153) & (!x407x) & (!x22204x)) + ((!n_n5149) & (!n_n5152) & (n_n5153) & (!x407x) & (x22204x)) + ((!n_n5149) & (!n_n5152) & (n_n5153) & (x407x) & (!x22204x)) + ((!n_n5149) & (!n_n5152) & (n_n5153) & (x407x) & (x22204x)) + ((!n_n5149) & (n_n5152) & (!n_n5153) & (!x407x) & (!x22204x)) + ((!n_n5149) & (n_n5152) & (!n_n5153) & (!x407x) & (x22204x)) + ((!n_n5149) & (n_n5152) & (!n_n5153) & (x407x) & (!x22204x)) + ((!n_n5149) & (n_n5152) & (!n_n5153) & (x407x) & (x22204x)) + ((!n_n5149) & (n_n5152) & (n_n5153) & (!x407x) & (!x22204x)) + ((!n_n5149) & (n_n5152) & (n_n5153) & (!x407x) & (x22204x)) + ((!n_n5149) & (n_n5152) & (n_n5153) & (x407x) & (!x22204x)) + ((!n_n5149) & (n_n5152) & (n_n5153) & (x407x) & (x22204x)) + ((n_n5149) & (!n_n5152) & (!n_n5153) & (!x407x) & (!x22204x)) + ((n_n5149) & (!n_n5152) & (!n_n5153) & (!x407x) & (x22204x)) + ((n_n5149) & (!n_n5152) & (!n_n5153) & (x407x) & (!x22204x)) + ((n_n5149) & (!n_n5152) & (!n_n5153) & (x407x) & (x22204x)) + ((n_n5149) & (!n_n5152) & (n_n5153) & (!x407x) & (!x22204x)) + ((n_n5149) & (!n_n5152) & (n_n5153) & (!x407x) & (x22204x)) + ((n_n5149) & (!n_n5152) & (n_n5153) & (x407x) & (!x22204x)) + ((n_n5149) & (!n_n5152) & (n_n5153) & (x407x) & (x22204x)) + ((n_n5149) & (n_n5152) & (!n_n5153) & (!x407x) & (!x22204x)) + ((n_n5149) & (n_n5152) & (!n_n5153) & (!x407x) & (x22204x)) + ((n_n5149) & (n_n5152) & (!n_n5153) & (x407x) & (!x22204x)) + ((n_n5149) & (n_n5152) & (!n_n5153) & (x407x) & (x22204x)) + ((n_n5149) & (n_n5152) & (n_n5153) & (!x407x) & (!x22204x)) + ((n_n5149) & (n_n5152) & (n_n5153) & (!x407x) & (x22204x)) + ((n_n5149) & (n_n5152) & (n_n5153) & (x407x) & (!x22204x)) + ((n_n5149) & (n_n5152) & (n_n5153) & (x407x) & (x22204x)));
	assign x15293x = (((!n_n5138) & (!n_n2304) & (!x211x) & (!x22184x)) + ((!n_n5138) & (!n_n2304) & (x211x) & (!x22184x)) + ((!n_n5138) & (!n_n2304) & (x211x) & (x22184x)) + ((!n_n5138) & (n_n2304) & (!x211x) & (!x22184x)) + ((!n_n5138) & (n_n2304) & (!x211x) & (x22184x)) + ((!n_n5138) & (n_n2304) & (x211x) & (!x22184x)) + ((!n_n5138) & (n_n2304) & (x211x) & (x22184x)) + ((n_n5138) & (!n_n2304) & (!x211x) & (!x22184x)) + ((n_n5138) & (!n_n2304) & (!x211x) & (x22184x)) + ((n_n5138) & (!n_n2304) & (x211x) & (!x22184x)) + ((n_n5138) & (!n_n2304) & (x211x) & (x22184x)) + ((n_n5138) & (n_n2304) & (!x211x) & (!x22184x)) + ((n_n5138) & (n_n2304) & (!x211x) & (x22184x)) + ((n_n5138) & (n_n2304) & (x211x) & (!x22184x)) + ((n_n5138) & (n_n2304) & (x211x) & (x22184x)));
	assign x15297x = (((!n_n2538) & (!n_n2539) & (!n_n2576) & (!n_n2577) & (x15293x)) + ((!n_n2538) & (!n_n2539) & (!n_n2576) & (n_n2577) & (!x15293x)) + ((!n_n2538) & (!n_n2539) & (!n_n2576) & (n_n2577) & (x15293x)) + ((!n_n2538) & (!n_n2539) & (n_n2576) & (!n_n2577) & (!x15293x)) + ((!n_n2538) & (!n_n2539) & (n_n2576) & (!n_n2577) & (x15293x)) + ((!n_n2538) & (!n_n2539) & (n_n2576) & (n_n2577) & (!x15293x)) + ((!n_n2538) & (!n_n2539) & (n_n2576) & (n_n2577) & (x15293x)) + ((!n_n2538) & (n_n2539) & (!n_n2576) & (!n_n2577) & (!x15293x)) + ((!n_n2538) & (n_n2539) & (!n_n2576) & (!n_n2577) & (x15293x)) + ((!n_n2538) & (n_n2539) & (!n_n2576) & (n_n2577) & (!x15293x)) + ((!n_n2538) & (n_n2539) & (!n_n2576) & (n_n2577) & (x15293x)) + ((!n_n2538) & (n_n2539) & (n_n2576) & (!n_n2577) & (!x15293x)) + ((!n_n2538) & (n_n2539) & (n_n2576) & (!n_n2577) & (x15293x)) + ((!n_n2538) & (n_n2539) & (n_n2576) & (n_n2577) & (!x15293x)) + ((!n_n2538) & (n_n2539) & (n_n2576) & (n_n2577) & (x15293x)) + ((n_n2538) & (!n_n2539) & (!n_n2576) & (!n_n2577) & (!x15293x)) + ((n_n2538) & (!n_n2539) & (!n_n2576) & (!n_n2577) & (x15293x)) + ((n_n2538) & (!n_n2539) & (!n_n2576) & (n_n2577) & (!x15293x)) + ((n_n2538) & (!n_n2539) & (!n_n2576) & (n_n2577) & (x15293x)) + ((n_n2538) & (!n_n2539) & (n_n2576) & (!n_n2577) & (!x15293x)) + ((n_n2538) & (!n_n2539) & (n_n2576) & (!n_n2577) & (x15293x)) + ((n_n2538) & (!n_n2539) & (n_n2576) & (n_n2577) & (!x15293x)) + ((n_n2538) & (!n_n2539) & (n_n2576) & (n_n2577) & (x15293x)) + ((n_n2538) & (n_n2539) & (!n_n2576) & (!n_n2577) & (!x15293x)) + ((n_n2538) & (n_n2539) & (!n_n2576) & (!n_n2577) & (x15293x)) + ((n_n2538) & (n_n2539) & (!n_n2576) & (n_n2577) & (!x15293x)) + ((n_n2538) & (n_n2539) & (!n_n2576) & (n_n2577) & (x15293x)) + ((n_n2538) & (n_n2539) & (n_n2576) & (!n_n2577) & (!x15293x)) + ((n_n2538) & (n_n2539) & (n_n2576) & (!n_n2577) & (x15293x)) + ((n_n2538) & (n_n2539) & (n_n2576) & (n_n2577) & (!x15293x)) + ((n_n2538) & (n_n2539) & (n_n2576) & (n_n2577) & (x15293x)));
	assign n_n2526 = (((!n_n2568) & (!n_n2569) & (!x15184x) & (!x15206x) & (x15205x)) + ((!n_n2568) & (!n_n2569) & (!x15184x) & (x15206x) & (!x15205x)) + ((!n_n2568) & (!n_n2569) & (!x15184x) & (x15206x) & (x15205x)) + ((!n_n2568) & (!n_n2569) & (x15184x) & (!x15206x) & (!x15205x)) + ((!n_n2568) & (!n_n2569) & (x15184x) & (!x15206x) & (x15205x)) + ((!n_n2568) & (!n_n2569) & (x15184x) & (x15206x) & (!x15205x)) + ((!n_n2568) & (!n_n2569) & (x15184x) & (x15206x) & (x15205x)) + ((!n_n2568) & (n_n2569) & (!x15184x) & (!x15206x) & (!x15205x)) + ((!n_n2568) & (n_n2569) & (!x15184x) & (!x15206x) & (x15205x)) + ((!n_n2568) & (n_n2569) & (!x15184x) & (x15206x) & (!x15205x)) + ((!n_n2568) & (n_n2569) & (!x15184x) & (x15206x) & (x15205x)) + ((!n_n2568) & (n_n2569) & (x15184x) & (!x15206x) & (!x15205x)) + ((!n_n2568) & (n_n2569) & (x15184x) & (!x15206x) & (x15205x)) + ((!n_n2568) & (n_n2569) & (x15184x) & (x15206x) & (!x15205x)) + ((!n_n2568) & (n_n2569) & (x15184x) & (x15206x) & (x15205x)) + ((n_n2568) & (!n_n2569) & (!x15184x) & (!x15206x) & (!x15205x)) + ((n_n2568) & (!n_n2569) & (!x15184x) & (!x15206x) & (x15205x)) + ((n_n2568) & (!n_n2569) & (!x15184x) & (x15206x) & (!x15205x)) + ((n_n2568) & (!n_n2569) & (!x15184x) & (x15206x) & (x15205x)) + ((n_n2568) & (!n_n2569) & (x15184x) & (!x15206x) & (!x15205x)) + ((n_n2568) & (!n_n2569) & (x15184x) & (!x15206x) & (x15205x)) + ((n_n2568) & (!n_n2569) & (x15184x) & (x15206x) & (!x15205x)) + ((n_n2568) & (!n_n2569) & (x15184x) & (x15206x) & (x15205x)) + ((n_n2568) & (n_n2569) & (!x15184x) & (!x15206x) & (!x15205x)) + ((n_n2568) & (n_n2569) & (!x15184x) & (!x15206x) & (x15205x)) + ((n_n2568) & (n_n2569) & (!x15184x) & (x15206x) & (!x15205x)) + ((n_n2568) & (n_n2569) & (!x15184x) & (x15206x) & (x15205x)) + ((n_n2568) & (n_n2569) & (x15184x) & (!x15206x) & (!x15205x)) + ((n_n2568) & (n_n2569) & (x15184x) & (!x15206x) & (x15205x)) + ((n_n2568) & (n_n2569) & (x15184x) & (x15206x) & (!x15205x)) + ((n_n2568) & (n_n2569) & (x15184x) & (x15206x) & (x15205x)));
	assign n_n2542 = (((!x90x) & (!n_n2584) & (!x15232x) & (!x22093x)) + ((!x90x) & (!n_n2584) & (x15232x) & (!x22093x)) + ((!x90x) & (!n_n2584) & (x15232x) & (x22093x)) + ((!x90x) & (n_n2584) & (!x15232x) & (!x22093x)) + ((!x90x) & (n_n2584) & (!x15232x) & (x22093x)) + ((!x90x) & (n_n2584) & (x15232x) & (!x22093x)) + ((!x90x) & (n_n2584) & (x15232x) & (x22093x)) + ((x90x) & (!n_n2584) & (!x15232x) & (!x22093x)) + ((x90x) & (!n_n2584) & (!x15232x) & (x22093x)) + ((x90x) & (!n_n2584) & (x15232x) & (!x22093x)) + ((x90x) & (!n_n2584) & (x15232x) & (x22093x)) + ((x90x) & (n_n2584) & (!x15232x) & (!x22093x)) + ((x90x) & (n_n2584) & (!x15232x) & (x22093x)) + ((x90x) & (n_n2584) & (x15232x) & (!x22093x)) + ((x90x) & (n_n2584) & (x15232x) & (x22093x)));
	assign n_n2541 = (((!x15239x) & (!x15240x) & (!x15249x) & (x15248x)) + ((!x15239x) & (!x15240x) & (x15249x) & (!x15248x)) + ((!x15239x) & (!x15240x) & (x15249x) & (x15248x)) + ((!x15239x) & (x15240x) & (!x15249x) & (!x15248x)) + ((!x15239x) & (x15240x) & (!x15249x) & (x15248x)) + ((!x15239x) & (x15240x) & (x15249x) & (!x15248x)) + ((!x15239x) & (x15240x) & (x15249x) & (x15248x)) + ((x15239x) & (!x15240x) & (!x15249x) & (!x15248x)) + ((x15239x) & (!x15240x) & (!x15249x) & (x15248x)) + ((x15239x) & (!x15240x) & (x15249x) & (!x15248x)) + ((x15239x) & (!x15240x) & (x15249x) & (x15248x)) + ((x15239x) & (x15240x) & (!x15249x) & (!x15248x)) + ((x15239x) & (x15240x) & (!x15249x) & (x15248x)) + ((x15239x) & (x15240x) & (x15249x) & (!x15248x)) + ((x15239x) & (x15240x) & (x15249x) & (x15248x)));
	assign x15264x = (((!x15254x) & (!x15255x) & (!n_n2586) & (x15262x)) + ((!x15254x) & (!x15255x) & (n_n2586) & (!x15262x)) + ((!x15254x) & (!x15255x) & (n_n2586) & (x15262x)) + ((!x15254x) & (x15255x) & (!n_n2586) & (!x15262x)) + ((!x15254x) & (x15255x) & (!n_n2586) & (x15262x)) + ((!x15254x) & (x15255x) & (n_n2586) & (!x15262x)) + ((!x15254x) & (x15255x) & (n_n2586) & (x15262x)) + ((x15254x) & (!x15255x) & (!n_n2586) & (!x15262x)) + ((x15254x) & (!x15255x) & (!n_n2586) & (x15262x)) + ((x15254x) & (!x15255x) & (n_n2586) & (!x15262x)) + ((x15254x) & (!x15255x) & (n_n2586) & (x15262x)) + ((x15254x) & (x15255x) & (!n_n2586) & (!x15262x)) + ((x15254x) & (x15255x) & (!n_n2586) & (x15262x)) + ((x15254x) & (x15255x) & (n_n2586) & (!x15262x)) + ((x15254x) & (x15255x) & (n_n2586) & (x15262x)));
	assign n_n4359 = (((i_1_) & (i_2_) & (i_0_) & (n_n509) & (x23x)));
	assign n_n4397 = (((!i_9_) & (n_n536) & (n_n482) & (n_n530)));
	assign x15308x = (((!n_n4359) & (!n_n4391) & (!n_n4384) & (n_n4397)) + ((!n_n4359) & (!n_n4391) & (n_n4384) & (!n_n4397)) + ((!n_n4359) & (!n_n4391) & (n_n4384) & (n_n4397)) + ((!n_n4359) & (n_n4391) & (!n_n4384) & (!n_n4397)) + ((!n_n4359) & (n_n4391) & (!n_n4384) & (n_n4397)) + ((!n_n4359) & (n_n4391) & (n_n4384) & (!n_n4397)) + ((!n_n4359) & (n_n4391) & (n_n4384) & (n_n4397)) + ((n_n4359) & (!n_n4391) & (!n_n4384) & (!n_n4397)) + ((n_n4359) & (!n_n4391) & (!n_n4384) & (n_n4397)) + ((n_n4359) & (!n_n4391) & (n_n4384) & (!n_n4397)) + ((n_n4359) & (!n_n4391) & (n_n4384) & (n_n4397)) + ((n_n4359) & (n_n4391) & (!n_n4384) & (!n_n4397)) + ((n_n4359) & (n_n4391) & (!n_n4384) & (n_n4397)) + ((n_n4359) & (n_n4391) & (n_n4384) & (!n_n4397)) + ((n_n4359) & (n_n4391) & (n_n4384) & (n_n4397)));
	assign n_n4431 = (((!i_9_) & (n_n536) & (n_n528) & (n_n464)));
	assign n_n4436 = (((i_9_) & (n_n536) & (n_n522) & (n_n464)));
	assign n_n4424 = (((i_9_) & (n_n536) & (n_n534) & (n_n464)));
	assign x15309x = (((!n_n4431) & (!n_n4436) & (!n_n4371) & (!n_n4424) & (n_n4417)) + ((!n_n4431) & (!n_n4436) & (!n_n4371) & (n_n4424) & (!n_n4417)) + ((!n_n4431) & (!n_n4436) & (!n_n4371) & (n_n4424) & (n_n4417)) + ((!n_n4431) & (!n_n4436) & (n_n4371) & (!n_n4424) & (!n_n4417)) + ((!n_n4431) & (!n_n4436) & (n_n4371) & (!n_n4424) & (n_n4417)) + ((!n_n4431) & (!n_n4436) & (n_n4371) & (n_n4424) & (!n_n4417)) + ((!n_n4431) & (!n_n4436) & (n_n4371) & (n_n4424) & (n_n4417)) + ((!n_n4431) & (n_n4436) & (!n_n4371) & (!n_n4424) & (!n_n4417)) + ((!n_n4431) & (n_n4436) & (!n_n4371) & (!n_n4424) & (n_n4417)) + ((!n_n4431) & (n_n4436) & (!n_n4371) & (n_n4424) & (!n_n4417)) + ((!n_n4431) & (n_n4436) & (!n_n4371) & (n_n4424) & (n_n4417)) + ((!n_n4431) & (n_n4436) & (n_n4371) & (!n_n4424) & (!n_n4417)) + ((!n_n4431) & (n_n4436) & (n_n4371) & (!n_n4424) & (n_n4417)) + ((!n_n4431) & (n_n4436) & (n_n4371) & (n_n4424) & (!n_n4417)) + ((!n_n4431) & (n_n4436) & (n_n4371) & (n_n4424) & (n_n4417)) + ((n_n4431) & (!n_n4436) & (!n_n4371) & (!n_n4424) & (!n_n4417)) + ((n_n4431) & (!n_n4436) & (!n_n4371) & (!n_n4424) & (n_n4417)) + ((n_n4431) & (!n_n4436) & (!n_n4371) & (n_n4424) & (!n_n4417)) + ((n_n4431) & (!n_n4436) & (!n_n4371) & (n_n4424) & (n_n4417)) + ((n_n4431) & (!n_n4436) & (n_n4371) & (!n_n4424) & (!n_n4417)) + ((n_n4431) & (!n_n4436) & (n_n4371) & (!n_n4424) & (n_n4417)) + ((n_n4431) & (!n_n4436) & (n_n4371) & (n_n4424) & (!n_n4417)) + ((n_n4431) & (!n_n4436) & (n_n4371) & (n_n4424) & (n_n4417)) + ((n_n4431) & (n_n4436) & (!n_n4371) & (!n_n4424) & (!n_n4417)) + ((n_n4431) & (n_n4436) & (!n_n4371) & (!n_n4424) & (n_n4417)) + ((n_n4431) & (n_n4436) & (!n_n4371) & (n_n4424) & (!n_n4417)) + ((n_n4431) & (n_n4436) & (!n_n4371) & (n_n4424) & (n_n4417)) + ((n_n4431) & (n_n4436) & (n_n4371) & (!n_n4424) & (!n_n4417)) + ((n_n4431) & (n_n4436) & (n_n4371) & (!n_n4424) & (n_n4417)) + ((n_n4431) & (n_n4436) & (n_n4371) & (n_n4424) & (!n_n4417)) + ((n_n4431) & (n_n4436) & (n_n4371) & (n_n4424) & (n_n4417)));
	assign n_n4451 = (((!i_9_) & (n_n524) & (n_n455) & (n_n535)));
	assign n_n4476 = (((i_9_) & (n_n455) & (n_n509) & (n_n530)));
	assign x15316x = (((!n_n4453) & (!n_n4451) & (!n_n4488) & (!n_n4457) & (n_n4476)) + ((!n_n4453) & (!n_n4451) & (!n_n4488) & (n_n4457) & (!n_n4476)) + ((!n_n4453) & (!n_n4451) & (!n_n4488) & (n_n4457) & (n_n4476)) + ((!n_n4453) & (!n_n4451) & (n_n4488) & (!n_n4457) & (!n_n4476)) + ((!n_n4453) & (!n_n4451) & (n_n4488) & (!n_n4457) & (n_n4476)) + ((!n_n4453) & (!n_n4451) & (n_n4488) & (n_n4457) & (!n_n4476)) + ((!n_n4453) & (!n_n4451) & (n_n4488) & (n_n4457) & (n_n4476)) + ((!n_n4453) & (n_n4451) & (!n_n4488) & (!n_n4457) & (!n_n4476)) + ((!n_n4453) & (n_n4451) & (!n_n4488) & (!n_n4457) & (n_n4476)) + ((!n_n4453) & (n_n4451) & (!n_n4488) & (n_n4457) & (!n_n4476)) + ((!n_n4453) & (n_n4451) & (!n_n4488) & (n_n4457) & (n_n4476)) + ((!n_n4453) & (n_n4451) & (n_n4488) & (!n_n4457) & (!n_n4476)) + ((!n_n4453) & (n_n4451) & (n_n4488) & (!n_n4457) & (n_n4476)) + ((!n_n4453) & (n_n4451) & (n_n4488) & (n_n4457) & (!n_n4476)) + ((!n_n4453) & (n_n4451) & (n_n4488) & (n_n4457) & (n_n4476)) + ((n_n4453) & (!n_n4451) & (!n_n4488) & (!n_n4457) & (!n_n4476)) + ((n_n4453) & (!n_n4451) & (!n_n4488) & (!n_n4457) & (n_n4476)) + ((n_n4453) & (!n_n4451) & (!n_n4488) & (n_n4457) & (!n_n4476)) + ((n_n4453) & (!n_n4451) & (!n_n4488) & (n_n4457) & (n_n4476)) + ((n_n4453) & (!n_n4451) & (n_n4488) & (!n_n4457) & (!n_n4476)) + ((n_n4453) & (!n_n4451) & (n_n4488) & (!n_n4457) & (n_n4476)) + ((n_n4453) & (!n_n4451) & (n_n4488) & (n_n4457) & (!n_n4476)) + ((n_n4453) & (!n_n4451) & (n_n4488) & (n_n4457) & (n_n4476)) + ((n_n4453) & (n_n4451) & (!n_n4488) & (!n_n4457) & (!n_n4476)) + ((n_n4453) & (n_n4451) & (!n_n4488) & (!n_n4457) & (n_n4476)) + ((n_n4453) & (n_n4451) & (!n_n4488) & (n_n4457) & (!n_n4476)) + ((n_n4453) & (n_n4451) & (!n_n4488) & (n_n4457) & (n_n4476)) + ((n_n4453) & (n_n4451) & (n_n4488) & (!n_n4457) & (!n_n4476)) + ((n_n4453) & (n_n4451) & (n_n4488) & (!n_n4457) & (n_n4476)) + ((n_n4453) & (n_n4451) & (n_n4488) & (n_n4457) & (!n_n4476)) + ((n_n4453) & (n_n4451) & (n_n4488) & (n_n4457) & (n_n4476)));
	assign n_n4478 = (((i_9_) & (n_n455) & (n_n528) & (n_n509)));
	assign n_n2844 = (((!x15316x) & (!n_n4487) & (!n_n4478) & (!n_n4456) & (n_n4458)) + ((!x15316x) & (!n_n4487) & (!n_n4478) & (n_n4456) & (!n_n4458)) + ((!x15316x) & (!n_n4487) & (!n_n4478) & (n_n4456) & (n_n4458)) + ((!x15316x) & (!n_n4487) & (n_n4478) & (!n_n4456) & (!n_n4458)) + ((!x15316x) & (!n_n4487) & (n_n4478) & (!n_n4456) & (n_n4458)) + ((!x15316x) & (!n_n4487) & (n_n4478) & (n_n4456) & (!n_n4458)) + ((!x15316x) & (!n_n4487) & (n_n4478) & (n_n4456) & (n_n4458)) + ((!x15316x) & (n_n4487) & (!n_n4478) & (!n_n4456) & (!n_n4458)) + ((!x15316x) & (n_n4487) & (!n_n4478) & (!n_n4456) & (n_n4458)) + ((!x15316x) & (n_n4487) & (!n_n4478) & (n_n4456) & (!n_n4458)) + ((!x15316x) & (n_n4487) & (!n_n4478) & (n_n4456) & (n_n4458)) + ((!x15316x) & (n_n4487) & (n_n4478) & (!n_n4456) & (!n_n4458)) + ((!x15316x) & (n_n4487) & (n_n4478) & (!n_n4456) & (n_n4458)) + ((!x15316x) & (n_n4487) & (n_n4478) & (n_n4456) & (!n_n4458)) + ((!x15316x) & (n_n4487) & (n_n4478) & (n_n4456) & (n_n4458)) + ((x15316x) & (!n_n4487) & (!n_n4478) & (!n_n4456) & (!n_n4458)) + ((x15316x) & (!n_n4487) & (!n_n4478) & (!n_n4456) & (n_n4458)) + ((x15316x) & (!n_n4487) & (!n_n4478) & (n_n4456) & (!n_n4458)) + ((x15316x) & (!n_n4487) & (!n_n4478) & (n_n4456) & (n_n4458)) + ((x15316x) & (!n_n4487) & (n_n4478) & (!n_n4456) & (!n_n4458)) + ((x15316x) & (!n_n4487) & (n_n4478) & (!n_n4456) & (n_n4458)) + ((x15316x) & (!n_n4487) & (n_n4478) & (n_n4456) & (!n_n4458)) + ((x15316x) & (!n_n4487) & (n_n4478) & (n_n4456) & (n_n4458)) + ((x15316x) & (n_n4487) & (!n_n4478) & (!n_n4456) & (!n_n4458)) + ((x15316x) & (n_n4487) & (!n_n4478) & (!n_n4456) & (n_n4458)) + ((x15316x) & (n_n4487) & (!n_n4478) & (n_n4456) & (!n_n4458)) + ((x15316x) & (n_n4487) & (!n_n4478) & (n_n4456) & (n_n4458)) + ((x15316x) & (n_n4487) & (n_n4478) & (!n_n4456) & (!n_n4458)) + ((x15316x) & (n_n4487) & (n_n4478) & (!n_n4456) & (n_n4458)) + ((x15316x) & (n_n4487) & (n_n4478) & (n_n4456) & (!n_n4458)) + ((x15316x) & (n_n4487) & (n_n4478) & (n_n4456) & (n_n4458)));
	assign n_n4345 = (((!i_9_) & (n_n536) & (n_n534) & (n_n509)));
	assign n_n4319 = (((!i_9_) & (n_n536) & (n_n528) & (n_n535)));
	assign n_n4355 = (((!i_9_) & (n_n536) & (n_n524) & (n_n509)));
	assign n_n4335 = (((!i_9_) & (n_n536) & (n_n518) & (n_n528)));
	assign n_n4316 = (((i_9_) & (n_n536) & (n_n535) & (n_n530)));
	assign x15323x = (((!n_n4345) & (!n_n4319) & (!n_n4355) & (!n_n4335) & (n_n4316)) + ((!n_n4345) & (!n_n4319) & (!n_n4355) & (n_n4335) & (!n_n4316)) + ((!n_n4345) & (!n_n4319) & (!n_n4355) & (n_n4335) & (n_n4316)) + ((!n_n4345) & (!n_n4319) & (n_n4355) & (!n_n4335) & (!n_n4316)) + ((!n_n4345) & (!n_n4319) & (n_n4355) & (!n_n4335) & (n_n4316)) + ((!n_n4345) & (!n_n4319) & (n_n4355) & (n_n4335) & (!n_n4316)) + ((!n_n4345) & (!n_n4319) & (n_n4355) & (n_n4335) & (n_n4316)) + ((!n_n4345) & (n_n4319) & (!n_n4355) & (!n_n4335) & (!n_n4316)) + ((!n_n4345) & (n_n4319) & (!n_n4355) & (!n_n4335) & (n_n4316)) + ((!n_n4345) & (n_n4319) & (!n_n4355) & (n_n4335) & (!n_n4316)) + ((!n_n4345) & (n_n4319) & (!n_n4355) & (n_n4335) & (n_n4316)) + ((!n_n4345) & (n_n4319) & (n_n4355) & (!n_n4335) & (!n_n4316)) + ((!n_n4345) & (n_n4319) & (n_n4355) & (!n_n4335) & (n_n4316)) + ((!n_n4345) & (n_n4319) & (n_n4355) & (n_n4335) & (!n_n4316)) + ((!n_n4345) & (n_n4319) & (n_n4355) & (n_n4335) & (n_n4316)) + ((n_n4345) & (!n_n4319) & (!n_n4355) & (!n_n4335) & (!n_n4316)) + ((n_n4345) & (!n_n4319) & (!n_n4355) & (!n_n4335) & (n_n4316)) + ((n_n4345) & (!n_n4319) & (!n_n4355) & (n_n4335) & (!n_n4316)) + ((n_n4345) & (!n_n4319) & (!n_n4355) & (n_n4335) & (n_n4316)) + ((n_n4345) & (!n_n4319) & (n_n4355) & (!n_n4335) & (!n_n4316)) + ((n_n4345) & (!n_n4319) & (n_n4355) & (!n_n4335) & (n_n4316)) + ((n_n4345) & (!n_n4319) & (n_n4355) & (n_n4335) & (!n_n4316)) + ((n_n4345) & (!n_n4319) & (n_n4355) & (n_n4335) & (n_n4316)) + ((n_n4345) & (n_n4319) & (!n_n4355) & (!n_n4335) & (!n_n4316)) + ((n_n4345) & (n_n4319) & (!n_n4355) & (!n_n4335) & (n_n4316)) + ((n_n4345) & (n_n4319) & (!n_n4355) & (n_n4335) & (!n_n4316)) + ((n_n4345) & (n_n4319) & (!n_n4355) & (n_n4335) & (n_n4316)) + ((n_n4345) & (n_n4319) & (n_n4355) & (!n_n4335) & (!n_n4316)) + ((n_n4345) & (n_n4319) & (n_n4355) & (!n_n4335) & (n_n4316)) + ((n_n4345) & (n_n4319) & (n_n4355) & (n_n4335) & (!n_n4316)) + ((n_n4345) & (n_n4319) & (n_n4355) & (n_n4335) & (n_n4316)));
	assign n_n4357 = (((i_1_) & (i_2_) & (i_0_) & (n_n509) & (x20x)));
	assign n_n4348 = (((i_9_) & (n_n536) & (n_n509) & (n_n530)));
	assign n_n2846 = (((!x15323x) & (!n_n4320) & (!n_n4315) & (!n_n4357) & (n_n4348)) + ((!x15323x) & (!n_n4320) & (!n_n4315) & (n_n4357) & (!n_n4348)) + ((!x15323x) & (!n_n4320) & (!n_n4315) & (n_n4357) & (n_n4348)) + ((!x15323x) & (!n_n4320) & (n_n4315) & (!n_n4357) & (!n_n4348)) + ((!x15323x) & (!n_n4320) & (n_n4315) & (!n_n4357) & (n_n4348)) + ((!x15323x) & (!n_n4320) & (n_n4315) & (n_n4357) & (!n_n4348)) + ((!x15323x) & (!n_n4320) & (n_n4315) & (n_n4357) & (n_n4348)) + ((!x15323x) & (n_n4320) & (!n_n4315) & (!n_n4357) & (!n_n4348)) + ((!x15323x) & (n_n4320) & (!n_n4315) & (!n_n4357) & (n_n4348)) + ((!x15323x) & (n_n4320) & (!n_n4315) & (n_n4357) & (!n_n4348)) + ((!x15323x) & (n_n4320) & (!n_n4315) & (n_n4357) & (n_n4348)) + ((!x15323x) & (n_n4320) & (n_n4315) & (!n_n4357) & (!n_n4348)) + ((!x15323x) & (n_n4320) & (n_n4315) & (!n_n4357) & (n_n4348)) + ((!x15323x) & (n_n4320) & (n_n4315) & (n_n4357) & (!n_n4348)) + ((!x15323x) & (n_n4320) & (n_n4315) & (n_n4357) & (n_n4348)) + ((x15323x) & (!n_n4320) & (!n_n4315) & (!n_n4357) & (!n_n4348)) + ((x15323x) & (!n_n4320) & (!n_n4315) & (!n_n4357) & (n_n4348)) + ((x15323x) & (!n_n4320) & (!n_n4315) & (n_n4357) & (!n_n4348)) + ((x15323x) & (!n_n4320) & (!n_n4315) & (n_n4357) & (n_n4348)) + ((x15323x) & (!n_n4320) & (n_n4315) & (!n_n4357) & (!n_n4348)) + ((x15323x) & (!n_n4320) & (n_n4315) & (!n_n4357) & (n_n4348)) + ((x15323x) & (!n_n4320) & (n_n4315) & (n_n4357) & (!n_n4348)) + ((x15323x) & (!n_n4320) & (n_n4315) & (n_n4357) & (n_n4348)) + ((x15323x) & (n_n4320) & (!n_n4315) & (!n_n4357) & (!n_n4348)) + ((x15323x) & (n_n4320) & (!n_n4315) & (!n_n4357) & (n_n4348)) + ((x15323x) & (n_n4320) & (!n_n4315) & (n_n4357) & (!n_n4348)) + ((x15323x) & (n_n4320) & (!n_n4315) & (n_n4357) & (n_n4348)) + ((x15323x) & (n_n4320) & (n_n4315) & (!n_n4357) & (!n_n4348)) + ((x15323x) & (n_n4320) & (n_n4315) & (!n_n4357) & (n_n4348)) + ((x15323x) & (n_n4320) & (n_n4315) & (n_n4357) & (!n_n4348)) + ((x15323x) & (n_n4320) & (n_n4315) & (n_n4357) & (n_n4348)));
	assign n_n4514 = (((i_9_) & (n_n524) & (n_n455) & (n_n491)));
	assign n_n4511 = (((!i_9_) & (n_n455) & (n_n528) & (n_n491)));
	assign n_n4525 = (((!i_9_) & (n_n482) & (n_n455) & (n_n530)));
	assign n_n4528 = (((i_9_) & (n_n526) & (n_n482) & (n_n455)));
	assign x15341x = (((!n_n4542) & (!n_n4552) & (!n_n4543) & (!n_n4527) & (n_n4534)) + ((!n_n4542) & (!n_n4552) & (!n_n4543) & (n_n4527) & (!n_n4534)) + ((!n_n4542) & (!n_n4552) & (!n_n4543) & (n_n4527) & (n_n4534)) + ((!n_n4542) & (!n_n4552) & (n_n4543) & (!n_n4527) & (!n_n4534)) + ((!n_n4542) & (!n_n4552) & (n_n4543) & (!n_n4527) & (n_n4534)) + ((!n_n4542) & (!n_n4552) & (n_n4543) & (n_n4527) & (!n_n4534)) + ((!n_n4542) & (!n_n4552) & (n_n4543) & (n_n4527) & (n_n4534)) + ((!n_n4542) & (n_n4552) & (!n_n4543) & (!n_n4527) & (!n_n4534)) + ((!n_n4542) & (n_n4552) & (!n_n4543) & (!n_n4527) & (n_n4534)) + ((!n_n4542) & (n_n4552) & (!n_n4543) & (n_n4527) & (!n_n4534)) + ((!n_n4542) & (n_n4552) & (!n_n4543) & (n_n4527) & (n_n4534)) + ((!n_n4542) & (n_n4552) & (n_n4543) & (!n_n4527) & (!n_n4534)) + ((!n_n4542) & (n_n4552) & (n_n4543) & (!n_n4527) & (n_n4534)) + ((!n_n4542) & (n_n4552) & (n_n4543) & (n_n4527) & (!n_n4534)) + ((!n_n4542) & (n_n4552) & (n_n4543) & (n_n4527) & (n_n4534)) + ((n_n4542) & (!n_n4552) & (!n_n4543) & (!n_n4527) & (!n_n4534)) + ((n_n4542) & (!n_n4552) & (!n_n4543) & (!n_n4527) & (n_n4534)) + ((n_n4542) & (!n_n4552) & (!n_n4543) & (n_n4527) & (!n_n4534)) + ((n_n4542) & (!n_n4552) & (!n_n4543) & (n_n4527) & (n_n4534)) + ((n_n4542) & (!n_n4552) & (n_n4543) & (!n_n4527) & (!n_n4534)) + ((n_n4542) & (!n_n4552) & (n_n4543) & (!n_n4527) & (n_n4534)) + ((n_n4542) & (!n_n4552) & (n_n4543) & (n_n4527) & (!n_n4534)) + ((n_n4542) & (!n_n4552) & (n_n4543) & (n_n4527) & (n_n4534)) + ((n_n4542) & (n_n4552) & (!n_n4543) & (!n_n4527) & (!n_n4534)) + ((n_n4542) & (n_n4552) & (!n_n4543) & (!n_n4527) & (n_n4534)) + ((n_n4542) & (n_n4552) & (!n_n4543) & (n_n4527) & (!n_n4534)) + ((n_n4542) & (n_n4552) & (!n_n4543) & (n_n4527) & (n_n4534)) + ((n_n4542) & (n_n4552) & (n_n4543) & (!n_n4527) & (!n_n4534)) + ((n_n4542) & (n_n4552) & (n_n4543) & (!n_n4527) & (n_n4534)) + ((n_n4542) & (n_n4552) & (n_n4543) & (n_n4527) & (!n_n4534)) + ((n_n4542) & (n_n4552) & (n_n4543) & (n_n4527) & (n_n4534)));
	assign x15342x = (((!n_n4514) & (!n_n4511) & (!n_n4525) & (!n_n4528) & (x15341x)) + ((!n_n4514) & (!n_n4511) & (!n_n4525) & (n_n4528) & (!x15341x)) + ((!n_n4514) & (!n_n4511) & (!n_n4525) & (n_n4528) & (x15341x)) + ((!n_n4514) & (!n_n4511) & (n_n4525) & (!n_n4528) & (!x15341x)) + ((!n_n4514) & (!n_n4511) & (n_n4525) & (!n_n4528) & (x15341x)) + ((!n_n4514) & (!n_n4511) & (n_n4525) & (n_n4528) & (!x15341x)) + ((!n_n4514) & (!n_n4511) & (n_n4525) & (n_n4528) & (x15341x)) + ((!n_n4514) & (n_n4511) & (!n_n4525) & (!n_n4528) & (!x15341x)) + ((!n_n4514) & (n_n4511) & (!n_n4525) & (!n_n4528) & (x15341x)) + ((!n_n4514) & (n_n4511) & (!n_n4525) & (n_n4528) & (!x15341x)) + ((!n_n4514) & (n_n4511) & (!n_n4525) & (n_n4528) & (x15341x)) + ((!n_n4514) & (n_n4511) & (n_n4525) & (!n_n4528) & (!x15341x)) + ((!n_n4514) & (n_n4511) & (n_n4525) & (!n_n4528) & (x15341x)) + ((!n_n4514) & (n_n4511) & (n_n4525) & (n_n4528) & (!x15341x)) + ((!n_n4514) & (n_n4511) & (n_n4525) & (n_n4528) & (x15341x)) + ((n_n4514) & (!n_n4511) & (!n_n4525) & (!n_n4528) & (!x15341x)) + ((n_n4514) & (!n_n4511) & (!n_n4525) & (!n_n4528) & (x15341x)) + ((n_n4514) & (!n_n4511) & (!n_n4525) & (n_n4528) & (!x15341x)) + ((n_n4514) & (!n_n4511) & (!n_n4525) & (n_n4528) & (x15341x)) + ((n_n4514) & (!n_n4511) & (n_n4525) & (!n_n4528) & (!x15341x)) + ((n_n4514) & (!n_n4511) & (n_n4525) & (!n_n4528) & (x15341x)) + ((n_n4514) & (!n_n4511) & (n_n4525) & (n_n4528) & (!x15341x)) + ((n_n4514) & (!n_n4511) & (n_n4525) & (n_n4528) & (x15341x)) + ((n_n4514) & (n_n4511) & (!n_n4525) & (!n_n4528) & (!x15341x)) + ((n_n4514) & (n_n4511) & (!n_n4525) & (!n_n4528) & (x15341x)) + ((n_n4514) & (n_n4511) & (!n_n4525) & (n_n4528) & (!x15341x)) + ((n_n4514) & (n_n4511) & (!n_n4525) & (n_n4528) & (x15341x)) + ((n_n4514) & (n_n4511) & (n_n4525) & (!n_n4528) & (!x15341x)) + ((n_n4514) & (n_n4511) & (n_n4525) & (!n_n4528) & (x15341x)) + ((n_n4514) & (n_n4511) & (n_n4525) & (n_n4528) & (!x15341x)) + ((n_n4514) & (n_n4511) & (n_n4525) & (n_n4528) & (x15341x)));
	assign n_n2842 = (((!n_n4598) & (!n_n4612) & (!n_n4570) & (!n_n4572) & (x15329x)) + ((!n_n4598) & (!n_n4612) & (!n_n4570) & (n_n4572) & (!x15329x)) + ((!n_n4598) & (!n_n4612) & (!n_n4570) & (n_n4572) & (x15329x)) + ((!n_n4598) & (!n_n4612) & (n_n4570) & (!n_n4572) & (!x15329x)) + ((!n_n4598) & (!n_n4612) & (n_n4570) & (!n_n4572) & (x15329x)) + ((!n_n4598) & (!n_n4612) & (n_n4570) & (n_n4572) & (!x15329x)) + ((!n_n4598) & (!n_n4612) & (n_n4570) & (n_n4572) & (x15329x)) + ((!n_n4598) & (n_n4612) & (!n_n4570) & (!n_n4572) & (!x15329x)) + ((!n_n4598) & (n_n4612) & (!n_n4570) & (!n_n4572) & (x15329x)) + ((!n_n4598) & (n_n4612) & (!n_n4570) & (n_n4572) & (!x15329x)) + ((!n_n4598) & (n_n4612) & (!n_n4570) & (n_n4572) & (x15329x)) + ((!n_n4598) & (n_n4612) & (n_n4570) & (!n_n4572) & (!x15329x)) + ((!n_n4598) & (n_n4612) & (n_n4570) & (!n_n4572) & (x15329x)) + ((!n_n4598) & (n_n4612) & (n_n4570) & (n_n4572) & (!x15329x)) + ((!n_n4598) & (n_n4612) & (n_n4570) & (n_n4572) & (x15329x)) + ((n_n4598) & (!n_n4612) & (!n_n4570) & (!n_n4572) & (!x15329x)) + ((n_n4598) & (!n_n4612) & (!n_n4570) & (!n_n4572) & (x15329x)) + ((n_n4598) & (!n_n4612) & (!n_n4570) & (n_n4572) & (!x15329x)) + ((n_n4598) & (!n_n4612) & (!n_n4570) & (n_n4572) & (x15329x)) + ((n_n4598) & (!n_n4612) & (n_n4570) & (!n_n4572) & (!x15329x)) + ((n_n4598) & (!n_n4612) & (n_n4570) & (!n_n4572) & (x15329x)) + ((n_n4598) & (!n_n4612) & (n_n4570) & (n_n4572) & (!x15329x)) + ((n_n4598) & (!n_n4612) & (n_n4570) & (n_n4572) & (x15329x)) + ((n_n4598) & (n_n4612) & (!n_n4570) & (!n_n4572) & (!x15329x)) + ((n_n4598) & (n_n4612) & (!n_n4570) & (!n_n4572) & (x15329x)) + ((n_n4598) & (n_n4612) & (!n_n4570) & (n_n4572) & (!x15329x)) + ((n_n4598) & (n_n4612) & (!n_n4570) & (n_n4572) & (x15329x)) + ((n_n4598) & (n_n4612) & (n_n4570) & (!n_n4572) & (!x15329x)) + ((n_n4598) & (n_n4612) & (n_n4570) & (!n_n4572) & (x15329x)) + ((n_n4598) & (n_n4612) & (n_n4570) & (n_n4572) & (!x15329x)) + ((n_n4598) & (n_n4612) & (n_n4570) & (n_n4572) & (x15329x)));
	assign x15334x = (((!n_n4659) & (!x75x) & (!n_n4689) & (n_n4698)) + ((!n_n4659) & (!x75x) & (n_n4689) & (!n_n4698)) + ((!n_n4659) & (!x75x) & (n_n4689) & (n_n4698)) + ((!n_n4659) & (x75x) & (!n_n4689) & (!n_n4698)) + ((!n_n4659) & (x75x) & (!n_n4689) & (n_n4698)) + ((!n_n4659) & (x75x) & (n_n4689) & (!n_n4698)) + ((!n_n4659) & (x75x) & (n_n4689) & (n_n4698)) + ((n_n4659) & (!x75x) & (!n_n4689) & (!n_n4698)) + ((n_n4659) & (!x75x) & (!n_n4689) & (n_n4698)) + ((n_n4659) & (!x75x) & (n_n4689) & (!n_n4698)) + ((n_n4659) & (!x75x) & (n_n4689) & (n_n4698)) + ((n_n4659) & (x75x) & (!n_n4689) & (!n_n4698)) + ((n_n4659) & (x75x) & (!n_n4689) & (n_n4698)) + ((n_n4659) & (x75x) & (n_n4689) & (!n_n4698)) + ((n_n4659) & (x75x) & (n_n4689) & (n_n4698)));
	assign x15335x = (((!n_n4634) & (!n_n4631) & (!n_n4691) & (!n_n4686) & (n_n4687)) + ((!n_n4634) & (!n_n4631) & (!n_n4691) & (n_n4686) & (!n_n4687)) + ((!n_n4634) & (!n_n4631) & (!n_n4691) & (n_n4686) & (n_n4687)) + ((!n_n4634) & (!n_n4631) & (n_n4691) & (!n_n4686) & (!n_n4687)) + ((!n_n4634) & (!n_n4631) & (n_n4691) & (!n_n4686) & (n_n4687)) + ((!n_n4634) & (!n_n4631) & (n_n4691) & (n_n4686) & (!n_n4687)) + ((!n_n4634) & (!n_n4631) & (n_n4691) & (n_n4686) & (n_n4687)) + ((!n_n4634) & (n_n4631) & (!n_n4691) & (!n_n4686) & (!n_n4687)) + ((!n_n4634) & (n_n4631) & (!n_n4691) & (!n_n4686) & (n_n4687)) + ((!n_n4634) & (n_n4631) & (!n_n4691) & (n_n4686) & (!n_n4687)) + ((!n_n4634) & (n_n4631) & (!n_n4691) & (n_n4686) & (n_n4687)) + ((!n_n4634) & (n_n4631) & (n_n4691) & (!n_n4686) & (!n_n4687)) + ((!n_n4634) & (n_n4631) & (n_n4691) & (!n_n4686) & (n_n4687)) + ((!n_n4634) & (n_n4631) & (n_n4691) & (n_n4686) & (!n_n4687)) + ((!n_n4634) & (n_n4631) & (n_n4691) & (n_n4686) & (n_n4687)) + ((n_n4634) & (!n_n4631) & (!n_n4691) & (!n_n4686) & (!n_n4687)) + ((n_n4634) & (!n_n4631) & (!n_n4691) & (!n_n4686) & (n_n4687)) + ((n_n4634) & (!n_n4631) & (!n_n4691) & (n_n4686) & (!n_n4687)) + ((n_n4634) & (!n_n4631) & (!n_n4691) & (n_n4686) & (n_n4687)) + ((n_n4634) & (!n_n4631) & (n_n4691) & (!n_n4686) & (!n_n4687)) + ((n_n4634) & (!n_n4631) & (n_n4691) & (!n_n4686) & (n_n4687)) + ((n_n4634) & (!n_n4631) & (n_n4691) & (n_n4686) & (!n_n4687)) + ((n_n4634) & (!n_n4631) & (n_n4691) & (n_n4686) & (n_n4687)) + ((n_n4634) & (n_n4631) & (!n_n4691) & (!n_n4686) & (!n_n4687)) + ((n_n4634) & (n_n4631) & (!n_n4691) & (!n_n4686) & (n_n4687)) + ((n_n4634) & (n_n4631) & (!n_n4691) & (n_n4686) & (!n_n4687)) + ((n_n4634) & (n_n4631) & (!n_n4691) & (n_n4686) & (n_n4687)) + ((n_n4634) & (n_n4631) & (n_n4691) & (!n_n4686) & (!n_n4687)) + ((n_n4634) & (n_n4631) & (n_n4691) & (!n_n4686) & (n_n4687)) + ((n_n4634) & (n_n4631) & (n_n4691) & (n_n4686) & (!n_n4687)) + ((n_n4634) & (n_n4631) & (n_n4691) & (n_n4686) & (n_n4687)));
	assign n_n2827 = (((!x15342x) & (!n_n2842) & (!x15334x) & (x15335x)) + ((!x15342x) & (!n_n2842) & (x15334x) & (!x15335x)) + ((!x15342x) & (!n_n2842) & (x15334x) & (x15335x)) + ((!x15342x) & (n_n2842) & (!x15334x) & (!x15335x)) + ((!x15342x) & (n_n2842) & (!x15334x) & (x15335x)) + ((!x15342x) & (n_n2842) & (x15334x) & (!x15335x)) + ((!x15342x) & (n_n2842) & (x15334x) & (x15335x)) + ((x15342x) & (!n_n2842) & (!x15334x) & (!x15335x)) + ((x15342x) & (!n_n2842) & (!x15334x) & (x15335x)) + ((x15342x) & (!n_n2842) & (x15334x) & (!x15335x)) + ((x15342x) & (!n_n2842) & (x15334x) & (x15335x)) + ((x15342x) & (n_n2842) & (!x15334x) & (!x15335x)) + ((x15342x) & (n_n2842) & (!x15334x) & (x15335x)) + ((x15342x) & (n_n2842) & (x15334x) & (!x15335x)) + ((x15342x) & (n_n2842) & (x15334x) & (x15335x)));
	assign x15369x = (((!n_n5090) & (!n_n5068) & (!n_n5080) & (!x279x) & (x15367x)) + ((!n_n5090) & (!n_n5068) & (!n_n5080) & (x279x) & (!x15367x)) + ((!n_n5090) & (!n_n5068) & (!n_n5080) & (x279x) & (x15367x)) + ((!n_n5090) & (!n_n5068) & (n_n5080) & (!x279x) & (!x15367x)) + ((!n_n5090) & (!n_n5068) & (n_n5080) & (!x279x) & (x15367x)) + ((!n_n5090) & (!n_n5068) & (n_n5080) & (x279x) & (!x15367x)) + ((!n_n5090) & (!n_n5068) & (n_n5080) & (x279x) & (x15367x)) + ((!n_n5090) & (n_n5068) & (!n_n5080) & (!x279x) & (!x15367x)) + ((!n_n5090) & (n_n5068) & (!n_n5080) & (!x279x) & (x15367x)) + ((!n_n5090) & (n_n5068) & (!n_n5080) & (x279x) & (!x15367x)) + ((!n_n5090) & (n_n5068) & (!n_n5080) & (x279x) & (x15367x)) + ((!n_n5090) & (n_n5068) & (n_n5080) & (!x279x) & (!x15367x)) + ((!n_n5090) & (n_n5068) & (n_n5080) & (!x279x) & (x15367x)) + ((!n_n5090) & (n_n5068) & (n_n5080) & (x279x) & (!x15367x)) + ((!n_n5090) & (n_n5068) & (n_n5080) & (x279x) & (x15367x)) + ((n_n5090) & (!n_n5068) & (!n_n5080) & (!x279x) & (!x15367x)) + ((n_n5090) & (!n_n5068) & (!n_n5080) & (!x279x) & (x15367x)) + ((n_n5090) & (!n_n5068) & (!n_n5080) & (x279x) & (!x15367x)) + ((n_n5090) & (!n_n5068) & (!n_n5080) & (x279x) & (x15367x)) + ((n_n5090) & (!n_n5068) & (n_n5080) & (!x279x) & (!x15367x)) + ((n_n5090) & (!n_n5068) & (n_n5080) & (!x279x) & (x15367x)) + ((n_n5090) & (!n_n5068) & (n_n5080) & (x279x) & (!x15367x)) + ((n_n5090) & (!n_n5068) & (n_n5080) & (x279x) & (x15367x)) + ((n_n5090) & (n_n5068) & (!n_n5080) & (!x279x) & (!x15367x)) + ((n_n5090) & (n_n5068) & (!n_n5080) & (!x279x) & (x15367x)) + ((n_n5090) & (n_n5068) & (!n_n5080) & (x279x) & (!x15367x)) + ((n_n5090) & (n_n5068) & (!n_n5080) & (x279x) & (x15367x)) + ((n_n5090) & (n_n5068) & (n_n5080) & (!x279x) & (!x15367x)) + ((n_n5090) & (n_n5068) & (n_n5080) & (!x279x) & (x15367x)) + ((n_n5090) & (n_n5068) & (n_n5080) & (x279x) & (!x15367x)) + ((n_n5090) & (n_n5068) & (n_n5080) & (x279x) & (x15367x)));
	assign x15370x = (((!x15355x) & (!x15356x) & (!x15361x) & (x15362x)) + ((!x15355x) & (!x15356x) & (x15361x) & (!x15362x)) + ((!x15355x) & (!x15356x) & (x15361x) & (x15362x)) + ((!x15355x) & (x15356x) & (!x15361x) & (!x15362x)) + ((!x15355x) & (x15356x) & (!x15361x) & (x15362x)) + ((!x15355x) & (x15356x) & (x15361x) & (!x15362x)) + ((!x15355x) & (x15356x) & (x15361x) & (x15362x)) + ((x15355x) & (!x15356x) & (!x15361x) & (!x15362x)) + ((x15355x) & (!x15356x) & (!x15361x) & (x15362x)) + ((x15355x) & (!x15356x) & (x15361x) & (!x15362x)) + ((x15355x) & (!x15356x) & (x15361x) & (x15362x)) + ((x15355x) & (x15356x) & (!x15361x) & (!x15362x)) + ((x15355x) & (x15356x) & (!x15361x) & (x15362x)) + ((x15355x) & (x15356x) & (x15361x) & (!x15362x)) + ((x15355x) & (x15356x) & (x15361x) & (x15362x)));
	assign n_n2823 = (((!x15374x) & (!x15375x) & (!x15381x) & (!x15382x) & (x15383x)) + ((!x15374x) & (!x15375x) & (!x15381x) & (x15382x) & (!x15383x)) + ((!x15374x) & (!x15375x) & (!x15381x) & (x15382x) & (x15383x)) + ((!x15374x) & (!x15375x) & (x15381x) & (!x15382x) & (!x15383x)) + ((!x15374x) & (!x15375x) & (x15381x) & (!x15382x) & (x15383x)) + ((!x15374x) & (!x15375x) & (x15381x) & (x15382x) & (!x15383x)) + ((!x15374x) & (!x15375x) & (x15381x) & (x15382x) & (x15383x)) + ((!x15374x) & (x15375x) & (!x15381x) & (!x15382x) & (!x15383x)) + ((!x15374x) & (x15375x) & (!x15381x) & (!x15382x) & (x15383x)) + ((!x15374x) & (x15375x) & (!x15381x) & (x15382x) & (!x15383x)) + ((!x15374x) & (x15375x) & (!x15381x) & (x15382x) & (x15383x)) + ((!x15374x) & (x15375x) & (x15381x) & (!x15382x) & (!x15383x)) + ((!x15374x) & (x15375x) & (x15381x) & (!x15382x) & (x15383x)) + ((!x15374x) & (x15375x) & (x15381x) & (x15382x) & (!x15383x)) + ((!x15374x) & (x15375x) & (x15381x) & (x15382x) & (x15383x)) + ((x15374x) & (!x15375x) & (!x15381x) & (!x15382x) & (!x15383x)) + ((x15374x) & (!x15375x) & (!x15381x) & (!x15382x) & (x15383x)) + ((x15374x) & (!x15375x) & (!x15381x) & (x15382x) & (!x15383x)) + ((x15374x) & (!x15375x) & (!x15381x) & (x15382x) & (x15383x)) + ((x15374x) & (!x15375x) & (x15381x) & (!x15382x) & (!x15383x)) + ((x15374x) & (!x15375x) & (x15381x) & (!x15382x) & (x15383x)) + ((x15374x) & (!x15375x) & (x15381x) & (x15382x) & (!x15383x)) + ((x15374x) & (!x15375x) & (x15381x) & (x15382x) & (x15383x)) + ((x15374x) & (x15375x) & (!x15381x) & (!x15382x) & (!x15383x)) + ((x15374x) & (x15375x) & (!x15381x) & (!x15382x) & (x15383x)) + ((x15374x) & (x15375x) & (!x15381x) & (x15382x) & (!x15383x)) + ((x15374x) & (x15375x) & (!x15381x) & (x15382x) & (x15383x)) + ((x15374x) & (x15375x) & (x15381x) & (!x15382x) & (!x15383x)) + ((x15374x) & (x15375x) & (x15381x) & (!x15382x) & (x15383x)) + ((x15374x) & (x15375x) & (x15381x) & (x15382x) & (!x15383x)) + ((x15374x) & (x15375x) & (x15381x) & (x15382x) & (x15383x)));
	assign x15398x = (((!n_n4931) & (!n_n4948) & (!n_n4957) & (!x141x) & (x15396x)) + ((!n_n4931) & (!n_n4948) & (!n_n4957) & (x141x) & (!x15396x)) + ((!n_n4931) & (!n_n4948) & (!n_n4957) & (x141x) & (x15396x)) + ((!n_n4931) & (!n_n4948) & (n_n4957) & (!x141x) & (!x15396x)) + ((!n_n4931) & (!n_n4948) & (n_n4957) & (!x141x) & (x15396x)) + ((!n_n4931) & (!n_n4948) & (n_n4957) & (x141x) & (!x15396x)) + ((!n_n4931) & (!n_n4948) & (n_n4957) & (x141x) & (x15396x)) + ((!n_n4931) & (n_n4948) & (!n_n4957) & (!x141x) & (!x15396x)) + ((!n_n4931) & (n_n4948) & (!n_n4957) & (!x141x) & (x15396x)) + ((!n_n4931) & (n_n4948) & (!n_n4957) & (x141x) & (!x15396x)) + ((!n_n4931) & (n_n4948) & (!n_n4957) & (x141x) & (x15396x)) + ((!n_n4931) & (n_n4948) & (n_n4957) & (!x141x) & (!x15396x)) + ((!n_n4931) & (n_n4948) & (n_n4957) & (!x141x) & (x15396x)) + ((!n_n4931) & (n_n4948) & (n_n4957) & (x141x) & (!x15396x)) + ((!n_n4931) & (n_n4948) & (n_n4957) & (x141x) & (x15396x)) + ((n_n4931) & (!n_n4948) & (!n_n4957) & (!x141x) & (!x15396x)) + ((n_n4931) & (!n_n4948) & (!n_n4957) & (!x141x) & (x15396x)) + ((n_n4931) & (!n_n4948) & (!n_n4957) & (x141x) & (!x15396x)) + ((n_n4931) & (!n_n4948) & (!n_n4957) & (x141x) & (x15396x)) + ((n_n4931) & (!n_n4948) & (n_n4957) & (!x141x) & (!x15396x)) + ((n_n4931) & (!n_n4948) & (n_n4957) & (!x141x) & (x15396x)) + ((n_n4931) & (!n_n4948) & (n_n4957) & (x141x) & (!x15396x)) + ((n_n4931) & (!n_n4948) & (n_n4957) & (x141x) & (x15396x)) + ((n_n4931) & (n_n4948) & (!n_n4957) & (!x141x) & (!x15396x)) + ((n_n4931) & (n_n4948) & (!n_n4957) & (!x141x) & (x15396x)) + ((n_n4931) & (n_n4948) & (!n_n4957) & (x141x) & (!x15396x)) + ((n_n4931) & (n_n4948) & (!n_n4957) & (x141x) & (x15396x)) + ((n_n4931) & (n_n4948) & (n_n4957) & (!x141x) & (!x15396x)) + ((n_n4931) & (n_n4948) & (n_n4957) & (!x141x) & (x15396x)) + ((n_n4931) & (n_n4948) & (n_n4957) & (x141x) & (!x15396x)) + ((n_n4931) & (n_n4948) & (n_n4957) & (x141x) & (x15396x)));
	assign x15399x = (((!x15348x) & (!x15349x) & (n_n2835)) + ((!x15348x) & (x15349x) & (!n_n2835)) + ((!x15348x) & (x15349x) & (n_n2835)) + ((x15348x) & (!x15349x) & (!n_n2835)) + ((x15348x) & (!x15349x) & (n_n2835)) + ((x15348x) & (x15349x) & (!n_n2835)) + ((x15348x) & (x15349x) & (n_n2835)));
	assign n_n2821 = (((!x15369x) & (!x15370x) & (!n_n2823) & (!x15398x) & (x15399x)) + ((!x15369x) & (!x15370x) & (!n_n2823) & (x15398x) & (!x15399x)) + ((!x15369x) & (!x15370x) & (!n_n2823) & (x15398x) & (x15399x)) + ((!x15369x) & (!x15370x) & (n_n2823) & (!x15398x) & (!x15399x)) + ((!x15369x) & (!x15370x) & (n_n2823) & (!x15398x) & (x15399x)) + ((!x15369x) & (!x15370x) & (n_n2823) & (x15398x) & (!x15399x)) + ((!x15369x) & (!x15370x) & (n_n2823) & (x15398x) & (x15399x)) + ((!x15369x) & (x15370x) & (!n_n2823) & (!x15398x) & (!x15399x)) + ((!x15369x) & (x15370x) & (!n_n2823) & (!x15398x) & (x15399x)) + ((!x15369x) & (x15370x) & (!n_n2823) & (x15398x) & (!x15399x)) + ((!x15369x) & (x15370x) & (!n_n2823) & (x15398x) & (x15399x)) + ((!x15369x) & (x15370x) & (n_n2823) & (!x15398x) & (!x15399x)) + ((!x15369x) & (x15370x) & (n_n2823) & (!x15398x) & (x15399x)) + ((!x15369x) & (x15370x) & (n_n2823) & (x15398x) & (!x15399x)) + ((!x15369x) & (x15370x) & (n_n2823) & (x15398x) & (x15399x)) + ((x15369x) & (!x15370x) & (!n_n2823) & (!x15398x) & (!x15399x)) + ((x15369x) & (!x15370x) & (!n_n2823) & (!x15398x) & (x15399x)) + ((x15369x) & (!x15370x) & (!n_n2823) & (x15398x) & (!x15399x)) + ((x15369x) & (!x15370x) & (!n_n2823) & (x15398x) & (x15399x)) + ((x15369x) & (!x15370x) & (n_n2823) & (!x15398x) & (!x15399x)) + ((x15369x) & (!x15370x) & (n_n2823) & (!x15398x) & (x15399x)) + ((x15369x) & (!x15370x) & (n_n2823) & (x15398x) & (!x15399x)) + ((x15369x) & (!x15370x) & (n_n2823) & (x15398x) & (x15399x)) + ((x15369x) & (x15370x) & (!n_n2823) & (!x15398x) & (!x15399x)) + ((x15369x) & (x15370x) & (!n_n2823) & (!x15398x) & (x15399x)) + ((x15369x) & (x15370x) & (!n_n2823) & (x15398x) & (!x15399x)) + ((x15369x) & (x15370x) & (!n_n2823) & (x15398x) & (x15399x)) + ((x15369x) & (x15370x) & (n_n2823) & (!x15398x) & (!x15399x)) + ((x15369x) & (x15370x) & (n_n2823) & (!x15398x) & (x15399x)) + ((x15369x) & (x15370x) & (n_n2823) & (x15398x) & (!x15399x)) + ((x15369x) & (x15370x) & (n_n2823) & (x15398x) & (x15399x)));
	assign x73x = (((!i_9_) & (n_n532) & (n_n509) & (n_n325) & (!n_n530)) + ((!i_9_) & (n_n532) & (n_n509) & (n_n325) & (n_n530)) + ((i_9_) & (!n_n532) & (n_n509) & (n_n325) & (n_n530)) + ((i_9_) & (n_n532) & (n_n509) & (n_n325) & (n_n530)));
	assign n_n4700 = (((i_9_) & (n_n325) & (n_n535) & (n_n530)));
	assign n_n1760 = (((!n_n524) & (!n_n526) & (!n_n509) & (!x14x) & (n_n4733)) + ((!n_n524) & (!n_n526) & (!n_n509) & (x14x) & (n_n4733)) + ((!n_n524) & (!n_n526) & (n_n509) & (!x14x) & (n_n4733)) + ((!n_n524) & (!n_n526) & (n_n509) & (x14x) & (n_n4733)) + ((!n_n524) & (n_n526) & (!n_n509) & (!x14x) & (n_n4733)) + ((!n_n524) & (n_n526) & (!n_n509) & (x14x) & (n_n4733)) + ((!n_n524) & (n_n526) & (n_n509) & (!x14x) & (n_n4733)) + ((!n_n524) & (n_n526) & (n_n509) & (x14x) & (!n_n4733)) + ((!n_n524) & (n_n526) & (n_n509) & (x14x) & (n_n4733)) + ((n_n524) & (!n_n526) & (!n_n509) & (!x14x) & (n_n4733)) + ((n_n524) & (!n_n526) & (!n_n509) & (x14x) & (n_n4733)) + ((n_n524) & (!n_n526) & (n_n509) & (!x14x) & (n_n4733)) + ((n_n524) & (!n_n526) & (n_n509) & (x14x) & (!n_n4733)) + ((n_n524) & (!n_n526) & (n_n509) & (x14x) & (n_n4733)) + ((n_n524) & (n_n526) & (!n_n509) & (!x14x) & (n_n4733)) + ((n_n524) & (n_n526) & (!n_n509) & (x14x) & (n_n4733)) + ((n_n524) & (n_n526) & (n_n509) & (!x14x) & (n_n4733)) + ((n_n524) & (n_n526) & (n_n509) & (x14x) & (!n_n4733)) + ((n_n524) & (n_n526) & (n_n509) & (x14x) & (n_n4733)));
	assign x15414x = (((!i_9_) & (!n_n534) & (!n_n509) & (!n_n325) & (n_n4711)) + ((!i_9_) & (!n_n534) & (!n_n509) & (n_n325) & (n_n4711)) + ((!i_9_) & (!n_n534) & (n_n509) & (!n_n325) & (n_n4711)) + ((!i_9_) & (!n_n534) & (n_n509) & (n_n325) & (n_n4711)) + ((!i_9_) & (n_n534) & (!n_n509) & (!n_n325) & (n_n4711)) + ((!i_9_) & (n_n534) & (!n_n509) & (n_n325) & (n_n4711)) + ((!i_9_) & (n_n534) & (n_n509) & (!n_n325) & (n_n4711)) + ((!i_9_) & (n_n534) & (n_n509) & (n_n325) & (!n_n4711)) + ((!i_9_) & (n_n534) & (n_n509) & (n_n325) & (n_n4711)) + ((i_9_) & (!n_n534) & (!n_n509) & (!n_n325) & (n_n4711)) + ((i_9_) & (!n_n534) & (!n_n509) & (n_n325) & (n_n4711)) + ((i_9_) & (!n_n534) & (n_n509) & (!n_n325) & (n_n4711)) + ((i_9_) & (!n_n534) & (n_n509) & (n_n325) & (n_n4711)) + ((i_9_) & (n_n534) & (!n_n509) & (!n_n325) & (n_n4711)) + ((i_9_) & (n_n534) & (!n_n509) & (n_n325) & (n_n4711)) + ((i_9_) & (n_n534) & (n_n509) & (!n_n325) & (n_n4711)) + ((i_9_) & (n_n534) & (n_n509) & (n_n325) & (n_n4711)));
	assign x15418x = (((!n_n4718) & (!x73x) & (!n_n4700) & (!n_n1760) & (x15414x)) + ((!n_n4718) & (!x73x) & (!n_n4700) & (n_n1760) & (!x15414x)) + ((!n_n4718) & (!x73x) & (!n_n4700) & (n_n1760) & (x15414x)) + ((!n_n4718) & (!x73x) & (n_n4700) & (!n_n1760) & (!x15414x)) + ((!n_n4718) & (!x73x) & (n_n4700) & (!n_n1760) & (x15414x)) + ((!n_n4718) & (!x73x) & (n_n4700) & (n_n1760) & (!x15414x)) + ((!n_n4718) & (!x73x) & (n_n4700) & (n_n1760) & (x15414x)) + ((!n_n4718) & (x73x) & (!n_n4700) & (!n_n1760) & (!x15414x)) + ((!n_n4718) & (x73x) & (!n_n4700) & (!n_n1760) & (x15414x)) + ((!n_n4718) & (x73x) & (!n_n4700) & (n_n1760) & (!x15414x)) + ((!n_n4718) & (x73x) & (!n_n4700) & (n_n1760) & (x15414x)) + ((!n_n4718) & (x73x) & (n_n4700) & (!n_n1760) & (!x15414x)) + ((!n_n4718) & (x73x) & (n_n4700) & (!n_n1760) & (x15414x)) + ((!n_n4718) & (x73x) & (n_n4700) & (n_n1760) & (!x15414x)) + ((!n_n4718) & (x73x) & (n_n4700) & (n_n1760) & (x15414x)) + ((n_n4718) & (!x73x) & (!n_n4700) & (!n_n1760) & (!x15414x)) + ((n_n4718) & (!x73x) & (!n_n4700) & (!n_n1760) & (x15414x)) + ((n_n4718) & (!x73x) & (!n_n4700) & (n_n1760) & (!x15414x)) + ((n_n4718) & (!x73x) & (!n_n4700) & (n_n1760) & (x15414x)) + ((n_n4718) & (!x73x) & (n_n4700) & (!n_n1760) & (!x15414x)) + ((n_n4718) & (!x73x) & (n_n4700) & (!n_n1760) & (x15414x)) + ((n_n4718) & (!x73x) & (n_n4700) & (n_n1760) & (!x15414x)) + ((n_n4718) & (!x73x) & (n_n4700) & (n_n1760) & (x15414x)) + ((n_n4718) & (x73x) & (!n_n4700) & (!n_n1760) & (!x15414x)) + ((n_n4718) & (x73x) & (!n_n4700) & (!n_n1760) & (x15414x)) + ((n_n4718) & (x73x) & (!n_n4700) & (n_n1760) & (!x15414x)) + ((n_n4718) & (x73x) & (!n_n4700) & (n_n1760) & (x15414x)) + ((n_n4718) & (x73x) & (n_n4700) & (!n_n1760) & (!x15414x)) + ((n_n4718) & (x73x) & (n_n4700) & (!n_n1760) & (x15414x)) + ((n_n4718) & (x73x) & (n_n4700) & (n_n1760) & (!x15414x)) + ((n_n4718) & (x73x) & (n_n4700) & (n_n1760) & (x15414x)));
	assign x15406x = (((!n_n4788) & (!n_n4769) & (!n_n4794) & (n_n4797)) + ((!n_n4788) & (!n_n4769) & (n_n4794) & (!n_n4797)) + ((!n_n4788) & (!n_n4769) & (n_n4794) & (n_n4797)) + ((!n_n4788) & (n_n4769) & (!n_n4794) & (!n_n4797)) + ((!n_n4788) & (n_n4769) & (!n_n4794) & (n_n4797)) + ((!n_n4788) & (n_n4769) & (n_n4794) & (!n_n4797)) + ((!n_n4788) & (n_n4769) & (n_n4794) & (n_n4797)) + ((n_n4788) & (!n_n4769) & (!n_n4794) & (!n_n4797)) + ((n_n4788) & (!n_n4769) & (!n_n4794) & (n_n4797)) + ((n_n4788) & (!n_n4769) & (n_n4794) & (!n_n4797)) + ((n_n4788) & (!n_n4769) & (n_n4794) & (n_n4797)) + ((n_n4788) & (n_n4769) & (!n_n4794) & (!n_n4797)) + ((n_n4788) & (n_n4769) & (!n_n4794) & (n_n4797)) + ((n_n4788) & (n_n4769) & (n_n4794) & (!n_n4797)) + ((n_n4788) & (n_n4769) & (n_n4794) & (n_n4797)));
	assign x15407x = (((!n_n4757) & (!n_n4760) & (!n_n4778) & (!n_n4745) & (n_n4815)) + ((!n_n4757) & (!n_n4760) & (!n_n4778) & (n_n4745) & (!n_n4815)) + ((!n_n4757) & (!n_n4760) & (!n_n4778) & (n_n4745) & (n_n4815)) + ((!n_n4757) & (!n_n4760) & (n_n4778) & (!n_n4745) & (!n_n4815)) + ((!n_n4757) & (!n_n4760) & (n_n4778) & (!n_n4745) & (n_n4815)) + ((!n_n4757) & (!n_n4760) & (n_n4778) & (n_n4745) & (!n_n4815)) + ((!n_n4757) & (!n_n4760) & (n_n4778) & (n_n4745) & (n_n4815)) + ((!n_n4757) & (n_n4760) & (!n_n4778) & (!n_n4745) & (!n_n4815)) + ((!n_n4757) & (n_n4760) & (!n_n4778) & (!n_n4745) & (n_n4815)) + ((!n_n4757) & (n_n4760) & (!n_n4778) & (n_n4745) & (!n_n4815)) + ((!n_n4757) & (n_n4760) & (!n_n4778) & (n_n4745) & (n_n4815)) + ((!n_n4757) & (n_n4760) & (n_n4778) & (!n_n4745) & (!n_n4815)) + ((!n_n4757) & (n_n4760) & (n_n4778) & (!n_n4745) & (n_n4815)) + ((!n_n4757) & (n_n4760) & (n_n4778) & (n_n4745) & (!n_n4815)) + ((!n_n4757) & (n_n4760) & (n_n4778) & (n_n4745) & (n_n4815)) + ((n_n4757) & (!n_n4760) & (!n_n4778) & (!n_n4745) & (!n_n4815)) + ((n_n4757) & (!n_n4760) & (!n_n4778) & (!n_n4745) & (n_n4815)) + ((n_n4757) & (!n_n4760) & (!n_n4778) & (n_n4745) & (!n_n4815)) + ((n_n4757) & (!n_n4760) & (!n_n4778) & (n_n4745) & (n_n4815)) + ((n_n4757) & (!n_n4760) & (n_n4778) & (!n_n4745) & (!n_n4815)) + ((n_n4757) & (!n_n4760) & (n_n4778) & (!n_n4745) & (n_n4815)) + ((n_n4757) & (!n_n4760) & (n_n4778) & (n_n4745) & (!n_n4815)) + ((n_n4757) & (!n_n4760) & (n_n4778) & (n_n4745) & (n_n4815)) + ((n_n4757) & (n_n4760) & (!n_n4778) & (!n_n4745) & (!n_n4815)) + ((n_n4757) & (n_n4760) & (!n_n4778) & (!n_n4745) & (n_n4815)) + ((n_n4757) & (n_n4760) & (!n_n4778) & (n_n4745) & (!n_n4815)) + ((n_n4757) & (n_n4760) & (!n_n4778) & (n_n4745) & (n_n4815)) + ((n_n4757) & (n_n4760) & (n_n4778) & (!n_n4745) & (!n_n4815)) + ((n_n4757) & (n_n4760) & (n_n4778) & (!n_n4745) & (n_n4815)) + ((n_n4757) & (n_n4760) & (n_n4778) & (n_n4745) & (!n_n4815)) + ((n_n4757) & (n_n4760) & (n_n4778) & (n_n4745) & (n_n4815)));
	assign n_n2838 = (((!n_n4854) & (!n_n4817) & (!n_n4843) & (!n_n4823) & (x15413x)) + ((!n_n4854) & (!n_n4817) & (!n_n4843) & (n_n4823) & (!x15413x)) + ((!n_n4854) & (!n_n4817) & (!n_n4843) & (n_n4823) & (x15413x)) + ((!n_n4854) & (!n_n4817) & (n_n4843) & (!n_n4823) & (!x15413x)) + ((!n_n4854) & (!n_n4817) & (n_n4843) & (!n_n4823) & (x15413x)) + ((!n_n4854) & (!n_n4817) & (n_n4843) & (n_n4823) & (!x15413x)) + ((!n_n4854) & (!n_n4817) & (n_n4843) & (n_n4823) & (x15413x)) + ((!n_n4854) & (n_n4817) & (!n_n4843) & (!n_n4823) & (!x15413x)) + ((!n_n4854) & (n_n4817) & (!n_n4843) & (!n_n4823) & (x15413x)) + ((!n_n4854) & (n_n4817) & (!n_n4843) & (n_n4823) & (!x15413x)) + ((!n_n4854) & (n_n4817) & (!n_n4843) & (n_n4823) & (x15413x)) + ((!n_n4854) & (n_n4817) & (n_n4843) & (!n_n4823) & (!x15413x)) + ((!n_n4854) & (n_n4817) & (n_n4843) & (!n_n4823) & (x15413x)) + ((!n_n4854) & (n_n4817) & (n_n4843) & (n_n4823) & (!x15413x)) + ((!n_n4854) & (n_n4817) & (n_n4843) & (n_n4823) & (x15413x)) + ((n_n4854) & (!n_n4817) & (!n_n4843) & (!n_n4823) & (!x15413x)) + ((n_n4854) & (!n_n4817) & (!n_n4843) & (!n_n4823) & (x15413x)) + ((n_n4854) & (!n_n4817) & (!n_n4843) & (n_n4823) & (!x15413x)) + ((n_n4854) & (!n_n4817) & (!n_n4843) & (n_n4823) & (x15413x)) + ((n_n4854) & (!n_n4817) & (n_n4843) & (!n_n4823) & (!x15413x)) + ((n_n4854) & (!n_n4817) & (n_n4843) & (!n_n4823) & (x15413x)) + ((n_n4854) & (!n_n4817) & (n_n4843) & (n_n4823) & (!x15413x)) + ((n_n4854) & (!n_n4817) & (n_n4843) & (n_n4823) & (x15413x)) + ((n_n4854) & (n_n4817) & (!n_n4843) & (!n_n4823) & (!x15413x)) + ((n_n4854) & (n_n4817) & (!n_n4843) & (!n_n4823) & (x15413x)) + ((n_n4854) & (n_n4817) & (!n_n4843) & (n_n4823) & (!x15413x)) + ((n_n4854) & (n_n4817) & (!n_n4843) & (n_n4823) & (x15413x)) + ((n_n4854) & (n_n4817) & (n_n4843) & (!n_n4823) & (!x15413x)) + ((n_n4854) & (n_n4817) & (n_n4843) & (!n_n4823) & (x15413x)) + ((n_n4854) & (n_n4817) & (n_n4843) & (n_n4823) & (!x15413x)) + ((n_n4854) & (n_n4817) & (n_n4843) & (n_n4823) & (x15413x)));
	assign n_n2826 = (((!x15418x) & (!x15406x) & (!x15407x) & (n_n2838)) + ((!x15418x) & (!x15406x) & (x15407x) & (!n_n2838)) + ((!x15418x) & (!x15406x) & (x15407x) & (n_n2838)) + ((!x15418x) & (x15406x) & (!x15407x) & (!n_n2838)) + ((!x15418x) & (x15406x) & (!x15407x) & (n_n2838)) + ((!x15418x) & (x15406x) & (x15407x) & (!n_n2838)) + ((!x15418x) & (x15406x) & (x15407x) & (n_n2838)) + ((x15418x) & (!x15406x) & (!x15407x) & (!n_n2838)) + ((x15418x) & (!x15406x) & (!x15407x) & (n_n2838)) + ((x15418x) & (!x15406x) & (x15407x) & (!n_n2838)) + ((x15418x) & (!x15406x) & (x15407x) & (n_n2838)) + ((x15418x) & (x15406x) & (!x15407x) & (!n_n2838)) + ((x15418x) & (x15406x) & (!x15407x) & (n_n2838)) + ((x15418x) & (x15406x) & (x15407x) & (!n_n2838)) + ((x15418x) & (x15406x) & (x15407x) & (n_n2838)));
	assign n_n3001 = (((!n_n4466) & (!x412x) & (!n_n4472) & (!n_n4469) & (!x22082x)) + ((!n_n4466) & (!x412x) & (!n_n4472) & (n_n4469) & (!x22082x)) + ((!n_n4466) & (!x412x) & (!n_n4472) & (n_n4469) & (x22082x)) + ((!n_n4466) & (!x412x) & (n_n4472) & (!n_n4469) & (!x22082x)) + ((!n_n4466) & (!x412x) & (n_n4472) & (!n_n4469) & (x22082x)) + ((!n_n4466) & (!x412x) & (n_n4472) & (n_n4469) & (!x22082x)) + ((!n_n4466) & (!x412x) & (n_n4472) & (n_n4469) & (x22082x)) + ((!n_n4466) & (x412x) & (!n_n4472) & (!n_n4469) & (!x22082x)) + ((!n_n4466) & (x412x) & (!n_n4472) & (!n_n4469) & (x22082x)) + ((!n_n4466) & (x412x) & (!n_n4472) & (n_n4469) & (!x22082x)) + ((!n_n4466) & (x412x) & (!n_n4472) & (n_n4469) & (x22082x)) + ((!n_n4466) & (x412x) & (n_n4472) & (!n_n4469) & (!x22082x)) + ((!n_n4466) & (x412x) & (n_n4472) & (!n_n4469) & (x22082x)) + ((!n_n4466) & (x412x) & (n_n4472) & (n_n4469) & (!x22082x)) + ((!n_n4466) & (x412x) & (n_n4472) & (n_n4469) & (x22082x)) + ((n_n4466) & (!x412x) & (!n_n4472) & (!n_n4469) & (!x22082x)) + ((n_n4466) & (!x412x) & (!n_n4472) & (!n_n4469) & (x22082x)) + ((n_n4466) & (!x412x) & (!n_n4472) & (n_n4469) & (!x22082x)) + ((n_n4466) & (!x412x) & (!n_n4472) & (n_n4469) & (x22082x)) + ((n_n4466) & (!x412x) & (n_n4472) & (!n_n4469) & (!x22082x)) + ((n_n4466) & (!x412x) & (n_n4472) & (!n_n4469) & (x22082x)) + ((n_n4466) & (!x412x) & (n_n4472) & (n_n4469) & (!x22082x)) + ((n_n4466) & (!x412x) & (n_n4472) & (n_n4469) & (x22082x)) + ((n_n4466) & (x412x) & (!n_n4472) & (!n_n4469) & (!x22082x)) + ((n_n4466) & (x412x) & (!n_n4472) & (!n_n4469) & (x22082x)) + ((n_n4466) & (x412x) & (!n_n4472) & (n_n4469) & (!x22082x)) + ((n_n4466) & (x412x) & (!n_n4472) & (n_n4469) & (x22082x)) + ((n_n4466) & (x412x) & (n_n4472) & (!n_n4469) & (!x22082x)) + ((n_n4466) & (x412x) & (n_n4472) & (!n_n4469) & (x22082x)) + ((n_n4466) & (x412x) & (n_n4472) & (n_n4469) & (!x22082x)) + ((n_n4466) & (x412x) & (n_n4472) & (n_n4469) & (x22082x)));
	assign n_n3003 = (((!n_n4440) & (!x323x) & (!n_n4449) & (!x470x) & (x421x)) + ((!n_n4440) & (!x323x) & (!n_n4449) & (x470x) & (!x421x)) + ((!n_n4440) & (!x323x) & (!n_n4449) & (x470x) & (x421x)) + ((!n_n4440) & (!x323x) & (n_n4449) & (!x470x) & (!x421x)) + ((!n_n4440) & (!x323x) & (n_n4449) & (!x470x) & (x421x)) + ((!n_n4440) & (!x323x) & (n_n4449) & (x470x) & (!x421x)) + ((!n_n4440) & (!x323x) & (n_n4449) & (x470x) & (x421x)) + ((!n_n4440) & (x323x) & (!n_n4449) & (!x470x) & (!x421x)) + ((!n_n4440) & (x323x) & (!n_n4449) & (!x470x) & (x421x)) + ((!n_n4440) & (x323x) & (!n_n4449) & (x470x) & (!x421x)) + ((!n_n4440) & (x323x) & (!n_n4449) & (x470x) & (x421x)) + ((!n_n4440) & (x323x) & (n_n4449) & (!x470x) & (!x421x)) + ((!n_n4440) & (x323x) & (n_n4449) & (!x470x) & (x421x)) + ((!n_n4440) & (x323x) & (n_n4449) & (x470x) & (!x421x)) + ((!n_n4440) & (x323x) & (n_n4449) & (x470x) & (x421x)) + ((n_n4440) & (!x323x) & (!n_n4449) & (!x470x) & (!x421x)) + ((n_n4440) & (!x323x) & (!n_n4449) & (!x470x) & (x421x)) + ((n_n4440) & (!x323x) & (!n_n4449) & (x470x) & (!x421x)) + ((n_n4440) & (!x323x) & (!n_n4449) & (x470x) & (x421x)) + ((n_n4440) & (!x323x) & (n_n4449) & (!x470x) & (!x421x)) + ((n_n4440) & (!x323x) & (n_n4449) & (!x470x) & (x421x)) + ((n_n4440) & (!x323x) & (n_n4449) & (x470x) & (!x421x)) + ((n_n4440) & (!x323x) & (n_n4449) & (x470x) & (x421x)) + ((n_n4440) & (x323x) & (!n_n4449) & (!x470x) & (!x421x)) + ((n_n4440) & (x323x) & (!n_n4449) & (!x470x) & (x421x)) + ((n_n4440) & (x323x) & (!n_n4449) & (x470x) & (!x421x)) + ((n_n4440) & (x323x) & (!n_n4449) & (x470x) & (x421x)) + ((n_n4440) & (x323x) & (n_n4449) & (!x470x) & (!x421x)) + ((n_n4440) & (x323x) & (n_n4449) & (!x470x) & (x421x)) + ((n_n4440) & (x323x) & (n_n4449) & (x470x) & (!x421x)) + ((n_n4440) & (x323x) & (n_n4449) & (x470x) & (x421x)));
	assign x15459x = (((!n_n4463) & (!n_n4455) & (!n_n4450) & (n_n4452)) + ((!n_n4463) & (!n_n4455) & (n_n4450) & (!n_n4452)) + ((!n_n4463) & (!n_n4455) & (n_n4450) & (n_n4452)) + ((!n_n4463) & (n_n4455) & (!n_n4450) & (!n_n4452)) + ((!n_n4463) & (n_n4455) & (!n_n4450) & (n_n4452)) + ((!n_n4463) & (n_n4455) & (n_n4450) & (!n_n4452)) + ((!n_n4463) & (n_n4455) & (n_n4450) & (n_n4452)) + ((n_n4463) & (!n_n4455) & (!n_n4450) & (!n_n4452)) + ((n_n4463) & (!n_n4455) & (!n_n4450) & (n_n4452)) + ((n_n4463) & (!n_n4455) & (n_n4450) & (!n_n4452)) + ((n_n4463) & (!n_n4455) & (n_n4450) & (n_n4452)) + ((n_n4463) & (n_n4455) & (!n_n4450) & (!n_n4452)) + ((n_n4463) & (n_n4455) & (!n_n4450) & (n_n4452)) + ((n_n4463) & (n_n4455) & (n_n4450) & (!n_n4452)) + ((n_n4463) & (n_n4455) & (n_n4450) & (n_n4452)));
	assign x15460x = (((!n_n4459) & (!n_n4461) & (!n_n4454) & (!n_n4465) & (n_n4462)) + ((!n_n4459) & (!n_n4461) & (!n_n4454) & (n_n4465) & (!n_n4462)) + ((!n_n4459) & (!n_n4461) & (!n_n4454) & (n_n4465) & (n_n4462)) + ((!n_n4459) & (!n_n4461) & (n_n4454) & (!n_n4465) & (!n_n4462)) + ((!n_n4459) & (!n_n4461) & (n_n4454) & (!n_n4465) & (n_n4462)) + ((!n_n4459) & (!n_n4461) & (n_n4454) & (n_n4465) & (!n_n4462)) + ((!n_n4459) & (!n_n4461) & (n_n4454) & (n_n4465) & (n_n4462)) + ((!n_n4459) & (n_n4461) & (!n_n4454) & (!n_n4465) & (!n_n4462)) + ((!n_n4459) & (n_n4461) & (!n_n4454) & (!n_n4465) & (n_n4462)) + ((!n_n4459) & (n_n4461) & (!n_n4454) & (n_n4465) & (!n_n4462)) + ((!n_n4459) & (n_n4461) & (!n_n4454) & (n_n4465) & (n_n4462)) + ((!n_n4459) & (n_n4461) & (n_n4454) & (!n_n4465) & (!n_n4462)) + ((!n_n4459) & (n_n4461) & (n_n4454) & (!n_n4465) & (n_n4462)) + ((!n_n4459) & (n_n4461) & (n_n4454) & (n_n4465) & (!n_n4462)) + ((!n_n4459) & (n_n4461) & (n_n4454) & (n_n4465) & (n_n4462)) + ((n_n4459) & (!n_n4461) & (!n_n4454) & (!n_n4465) & (!n_n4462)) + ((n_n4459) & (!n_n4461) & (!n_n4454) & (!n_n4465) & (n_n4462)) + ((n_n4459) & (!n_n4461) & (!n_n4454) & (n_n4465) & (!n_n4462)) + ((n_n4459) & (!n_n4461) & (!n_n4454) & (n_n4465) & (n_n4462)) + ((n_n4459) & (!n_n4461) & (n_n4454) & (!n_n4465) & (!n_n4462)) + ((n_n4459) & (!n_n4461) & (n_n4454) & (!n_n4465) & (n_n4462)) + ((n_n4459) & (!n_n4461) & (n_n4454) & (n_n4465) & (!n_n4462)) + ((n_n4459) & (!n_n4461) & (n_n4454) & (n_n4465) & (n_n4462)) + ((n_n4459) & (n_n4461) & (!n_n4454) & (!n_n4465) & (!n_n4462)) + ((n_n4459) & (n_n4461) & (!n_n4454) & (!n_n4465) & (n_n4462)) + ((n_n4459) & (n_n4461) & (!n_n4454) & (n_n4465) & (!n_n4462)) + ((n_n4459) & (n_n4461) & (!n_n4454) & (n_n4465) & (n_n4462)) + ((n_n4459) & (n_n4461) & (n_n4454) & (!n_n4465) & (!n_n4462)) + ((n_n4459) & (n_n4461) & (n_n4454) & (!n_n4465) & (n_n4462)) + ((n_n4459) & (n_n4461) & (n_n4454) & (n_n4465) & (!n_n4462)) + ((n_n4459) & (n_n4461) & (n_n4454) & (n_n4465) & (n_n4462)));
	assign x15463x = (((!n_n3001) & (!n_n3003) & (!x15459x) & (x15460x)) + ((!n_n3001) & (!n_n3003) & (x15459x) & (!x15460x)) + ((!n_n3001) & (!n_n3003) & (x15459x) & (x15460x)) + ((!n_n3001) & (n_n3003) & (!x15459x) & (!x15460x)) + ((!n_n3001) & (n_n3003) & (!x15459x) & (x15460x)) + ((!n_n3001) & (n_n3003) & (x15459x) & (!x15460x)) + ((!n_n3001) & (n_n3003) & (x15459x) & (x15460x)) + ((n_n3001) & (!n_n3003) & (!x15459x) & (!x15460x)) + ((n_n3001) & (!n_n3003) & (!x15459x) & (x15460x)) + ((n_n3001) & (!n_n3003) & (x15459x) & (!x15460x)) + ((n_n3001) & (!n_n3003) & (x15459x) & (x15460x)) + ((n_n3001) & (n_n3003) & (!x15459x) & (!x15460x)) + ((n_n3001) & (n_n3003) & (!x15459x) & (x15460x)) + ((n_n3001) & (n_n3003) & (x15459x) & (!x15460x)) + ((n_n3001) & (n_n3003) & (x15459x) & (x15460x)));
	assign n_n2999 = (((!n_n4498) & (!n_n4499) & (!n_n4496) & (!x163x) & (!x22081x)) + ((!n_n4498) & (!n_n4499) & (!n_n4496) & (x163x) & (!x22081x)) + ((!n_n4498) & (!n_n4499) & (!n_n4496) & (x163x) & (x22081x)) + ((!n_n4498) & (!n_n4499) & (n_n4496) & (!x163x) & (!x22081x)) + ((!n_n4498) & (!n_n4499) & (n_n4496) & (!x163x) & (x22081x)) + ((!n_n4498) & (!n_n4499) & (n_n4496) & (x163x) & (!x22081x)) + ((!n_n4498) & (!n_n4499) & (n_n4496) & (x163x) & (x22081x)) + ((!n_n4498) & (n_n4499) & (!n_n4496) & (!x163x) & (!x22081x)) + ((!n_n4498) & (n_n4499) & (!n_n4496) & (!x163x) & (x22081x)) + ((!n_n4498) & (n_n4499) & (!n_n4496) & (x163x) & (!x22081x)) + ((!n_n4498) & (n_n4499) & (!n_n4496) & (x163x) & (x22081x)) + ((!n_n4498) & (n_n4499) & (n_n4496) & (!x163x) & (!x22081x)) + ((!n_n4498) & (n_n4499) & (n_n4496) & (!x163x) & (x22081x)) + ((!n_n4498) & (n_n4499) & (n_n4496) & (x163x) & (!x22081x)) + ((!n_n4498) & (n_n4499) & (n_n4496) & (x163x) & (x22081x)) + ((n_n4498) & (!n_n4499) & (!n_n4496) & (!x163x) & (!x22081x)) + ((n_n4498) & (!n_n4499) & (!n_n4496) & (!x163x) & (x22081x)) + ((n_n4498) & (!n_n4499) & (!n_n4496) & (x163x) & (!x22081x)) + ((n_n4498) & (!n_n4499) & (!n_n4496) & (x163x) & (x22081x)) + ((n_n4498) & (!n_n4499) & (n_n4496) & (!x163x) & (!x22081x)) + ((n_n4498) & (!n_n4499) & (n_n4496) & (!x163x) & (x22081x)) + ((n_n4498) & (!n_n4499) & (n_n4496) & (x163x) & (!x22081x)) + ((n_n4498) & (!n_n4499) & (n_n4496) & (x163x) & (x22081x)) + ((n_n4498) & (n_n4499) & (!n_n4496) & (!x163x) & (!x22081x)) + ((n_n4498) & (n_n4499) & (!n_n4496) & (!x163x) & (x22081x)) + ((n_n4498) & (n_n4499) & (!n_n4496) & (x163x) & (!x22081x)) + ((n_n4498) & (n_n4499) & (!n_n4496) & (x163x) & (x22081x)) + ((n_n4498) & (n_n4499) & (n_n4496) & (!x163x) & (!x22081x)) + ((n_n4498) & (n_n4499) & (n_n4496) & (!x163x) & (x22081x)) + ((n_n4498) & (n_n4499) & (n_n4496) & (x163x) & (!x22081x)) + ((n_n4498) & (n_n4499) & (n_n4496) & (x163x) & (x22081x)));
	assign x206x = (((!n_n4489) & (!x70x) & (!n_n3515) & (!n_n4486) & (n_n4484)) + ((!n_n4489) & (!x70x) & (!n_n3515) & (n_n4486) & (!n_n4484)) + ((!n_n4489) & (!x70x) & (!n_n3515) & (n_n4486) & (n_n4484)) + ((!n_n4489) & (!x70x) & (n_n3515) & (!n_n4486) & (!n_n4484)) + ((!n_n4489) & (!x70x) & (n_n3515) & (!n_n4486) & (n_n4484)) + ((!n_n4489) & (!x70x) & (n_n3515) & (n_n4486) & (!n_n4484)) + ((!n_n4489) & (!x70x) & (n_n3515) & (n_n4486) & (n_n4484)) + ((!n_n4489) & (x70x) & (!n_n3515) & (!n_n4486) & (!n_n4484)) + ((!n_n4489) & (x70x) & (!n_n3515) & (!n_n4486) & (n_n4484)) + ((!n_n4489) & (x70x) & (!n_n3515) & (n_n4486) & (!n_n4484)) + ((!n_n4489) & (x70x) & (!n_n3515) & (n_n4486) & (n_n4484)) + ((!n_n4489) & (x70x) & (n_n3515) & (!n_n4486) & (!n_n4484)) + ((!n_n4489) & (x70x) & (n_n3515) & (!n_n4486) & (n_n4484)) + ((!n_n4489) & (x70x) & (n_n3515) & (n_n4486) & (!n_n4484)) + ((!n_n4489) & (x70x) & (n_n3515) & (n_n4486) & (n_n4484)) + ((n_n4489) & (!x70x) & (!n_n3515) & (!n_n4486) & (!n_n4484)) + ((n_n4489) & (!x70x) & (!n_n3515) & (!n_n4486) & (n_n4484)) + ((n_n4489) & (!x70x) & (!n_n3515) & (n_n4486) & (!n_n4484)) + ((n_n4489) & (!x70x) & (!n_n3515) & (n_n4486) & (n_n4484)) + ((n_n4489) & (!x70x) & (n_n3515) & (!n_n4486) & (!n_n4484)) + ((n_n4489) & (!x70x) & (n_n3515) & (!n_n4486) & (n_n4484)) + ((n_n4489) & (!x70x) & (n_n3515) & (n_n4486) & (!n_n4484)) + ((n_n4489) & (!x70x) & (n_n3515) & (n_n4486) & (n_n4484)) + ((n_n4489) & (x70x) & (!n_n3515) & (!n_n4486) & (!n_n4484)) + ((n_n4489) & (x70x) & (!n_n3515) & (!n_n4486) & (n_n4484)) + ((n_n4489) & (x70x) & (!n_n3515) & (n_n4486) & (!n_n4484)) + ((n_n4489) & (x70x) & (!n_n3515) & (n_n4486) & (n_n4484)) + ((n_n4489) & (x70x) & (n_n3515) & (!n_n4486) & (!n_n4484)) + ((n_n4489) & (x70x) & (n_n3515) & (!n_n4486) & (n_n4484)) + ((n_n4489) & (x70x) & (n_n3515) & (n_n4486) & (!n_n4484)) + ((n_n4489) & (x70x) & (n_n3515) & (n_n4486) & (n_n4484)));
	assign x15437x = (((!x189x) & (!n_n4490) & (!n_n3509) & (!x162x) & (x15433x)) + ((!x189x) & (!n_n4490) & (!n_n3509) & (x162x) & (!x15433x)) + ((!x189x) & (!n_n4490) & (!n_n3509) & (x162x) & (x15433x)) + ((!x189x) & (!n_n4490) & (n_n3509) & (!x162x) & (!x15433x)) + ((!x189x) & (!n_n4490) & (n_n3509) & (!x162x) & (x15433x)) + ((!x189x) & (!n_n4490) & (n_n3509) & (x162x) & (!x15433x)) + ((!x189x) & (!n_n4490) & (n_n3509) & (x162x) & (x15433x)) + ((!x189x) & (n_n4490) & (!n_n3509) & (!x162x) & (!x15433x)) + ((!x189x) & (n_n4490) & (!n_n3509) & (!x162x) & (x15433x)) + ((!x189x) & (n_n4490) & (!n_n3509) & (x162x) & (!x15433x)) + ((!x189x) & (n_n4490) & (!n_n3509) & (x162x) & (x15433x)) + ((!x189x) & (n_n4490) & (n_n3509) & (!x162x) & (!x15433x)) + ((!x189x) & (n_n4490) & (n_n3509) & (!x162x) & (x15433x)) + ((!x189x) & (n_n4490) & (n_n3509) & (x162x) & (!x15433x)) + ((!x189x) & (n_n4490) & (n_n3509) & (x162x) & (x15433x)) + ((x189x) & (!n_n4490) & (!n_n3509) & (!x162x) & (!x15433x)) + ((x189x) & (!n_n4490) & (!n_n3509) & (!x162x) & (x15433x)) + ((x189x) & (!n_n4490) & (!n_n3509) & (x162x) & (!x15433x)) + ((x189x) & (!n_n4490) & (!n_n3509) & (x162x) & (x15433x)) + ((x189x) & (!n_n4490) & (n_n3509) & (!x162x) & (!x15433x)) + ((x189x) & (!n_n4490) & (n_n3509) & (!x162x) & (x15433x)) + ((x189x) & (!n_n4490) & (n_n3509) & (x162x) & (!x15433x)) + ((x189x) & (!n_n4490) & (n_n3509) & (x162x) & (x15433x)) + ((x189x) & (n_n4490) & (!n_n3509) & (!x162x) & (!x15433x)) + ((x189x) & (n_n4490) & (!n_n3509) & (!x162x) & (x15433x)) + ((x189x) & (n_n4490) & (!n_n3509) & (x162x) & (!x15433x)) + ((x189x) & (n_n4490) & (!n_n3509) & (x162x) & (x15433x)) + ((x189x) & (n_n4490) & (n_n3509) & (!x162x) & (!x15433x)) + ((x189x) & (n_n4490) & (n_n3509) & (!x162x) & (x15433x)) + ((x189x) & (n_n4490) & (n_n3509) & (x162x) & (!x15433x)) + ((x189x) & (n_n4490) & (n_n3509) & (x162x) & (x15433x)));
	assign n_n2929 = (((!n_n2997) & (!x15445x) & (!x15446x) & (x15453x)) + ((!n_n2997) & (!x15445x) & (x15446x) & (!x15453x)) + ((!n_n2997) & (!x15445x) & (x15446x) & (x15453x)) + ((!n_n2997) & (x15445x) & (!x15446x) & (!x15453x)) + ((!n_n2997) & (x15445x) & (!x15446x) & (x15453x)) + ((!n_n2997) & (x15445x) & (x15446x) & (!x15453x)) + ((!n_n2997) & (x15445x) & (x15446x) & (x15453x)) + ((n_n2997) & (!x15445x) & (!x15446x) & (!x15453x)) + ((n_n2997) & (!x15445x) & (!x15446x) & (x15453x)) + ((n_n2997) & (!x15445x) & (x15446x) & (!x15453x)) + ((n_n2997) & (!x15445x) & (x15446x) & (x15453x)) + ((n_n2997) & (x15445x) & (!x15446x) & (!x15453x)) + ((n_n2997) & (x15445x) & (!x15446x) & (x15453x)) + ((n_n2997) & (x15445x) & (x15446x) & (!x15453x)) + ((n_n2997) & (x15445x) & (x15446x) & (x15453x)));
	assign n_n2907 = (((!x15463x) & (!n_n2999) & (!x206x) & (!x15437x) & (n_n2929)) + ((!x15463x) & (!n_n2999) & (!x206x) & (x15437x) & (!n_n2929)) + ((!x15463x) & (!n_n2999) & (!x206x) & (x15437x) & (n_n2929)) + ((!x15463x) & (!n_n2999) & (x206x) & (!x15437x) & (!n_n2929)) + ((!x15463x) & (!n_n2999) & (x206x) & (!x15437x) & (n_n2929)) + ((!x15463x) & (!n_n2999) & (x206x) & (x15437x) & (!n_n2929)) + ((!x15463x) & (!n_n2999) & (x206x) & (x15437x) & (n_n2929)) + ((!x15463x) & (n_n2999) & (!x206x) & (!x15437x) & (!n_n2929)) + ((!x15463x) & (n_n2999) & (!x206x) & (!x15437x) & (n_n2929)) + ((!x15463x) & (n_n2999) & (!x206x) & (x15437x) & (!n_n2929)) + ((!x15463x) & (n_n2999) & (!x206x) & (x15437x) & (n_n2929)) + ((!x15463x) & (n_n2999) & (x206x) & (!x15437x) & (!n_n2929)) + ((!x15463x) & (n_n2999) & (x206x) & (!x15437x) & (n_n2929)) + ((!x15463x) & (n_n2999) & (x206x) & (x15437x) & (!n_n2929)) + ((!x15463x) & (n_n2999) & (x206x) & (x15437x) & (n_n2929)) + ((x15463x) & (!n_n2999) & (!x206x) & (!x15437x) & (!n_n2929)) + ((x15463x) & (!n_n2999) & (!x206x) & (!x15437x) & (n_n2929)) + ((x15463x) & (!n_n2999) & (!x206x) & (x15437x) & (!n_n2929)) + ((x15463x) & (!n_n2999) & (!x206x) & (x15437x) & (n_n2929)) + ((x15463x) & (!n_n2999) & (x206x) & (!x15437x) & (!n_n2929)) + ((x15463x) & (!n_n2999) & (x206x) & (!x15437x) & (n_n2929)) + ((x15463x) & (!n_n2999) & (x206x) & (x15437x) & (!n_n2929)) + ((x15463x) & (!n_n2999) & (x206x) & (x15437x) & (n_n2929)) + ((x15463x) & (n_n2999) & (!x206x) & (!x15437x) & (!n_n2929)) + ((x15463x) & (n_n2999) & (!x206x) & (!x15437x) & (n_n2929)) + ((x15463x) & (n_n2999) & (!x206x) & (x15437x) & (!n_n2929)) + ((x15463x) & (n_n2999) & (!x206x) & (x15437x) & (n_n2929)) + ((x15463x) & (n_n2999) & (x206x) & (!x15437x) & (!n_n2929)) + ((x15463x) & (n_n2999) & (x206x) & (!x15437x) & (n_n2929)) + ((x15463x) & (n_n2999) & (x206x) & (x15437x) & (!n_n2929)) + ((x15463x) & (n_n2999) & (x206x) & (x15437x) & (n_n2929)));
	assign x100x = (((!i_9_) & (!n_n518) & (!n_n390) & (!n_n534) & (n_n4583)) + ((!i_9_) & (!n_n518) & (!n_n390) & (n_n534) & (n_n4583)) + ((!i_9_) & (!n_n518) & (n_n390) & (!n_n534) & (n_n4583)) + ((!i_9_) & (!n_n518) & (n_n390) & (n_n534) & (n_n4583)) + ((!i_9_) & (n_n518) & (!n_n390) & (!n_n534) & (n_n4583)) + ((!i_9_) & (n_n518) & (!n_n390) & (n_n534) & (n_n4583)) + ((!i_9_) & (n_n518) & (n_n390) & (!n_n534) & (n_n4583)) + ((!i_9_) & (n_n518) & (n_n390) & (n_n534) & (n_n4583)) + ((i_9_) & (!n_n518) & (!n_n390) & (!n_n534) & (n_n4583)) + ((i_9_) & (!n_n518) & (!n_n390) & (n_n534) & (n_n4583)) + ((i_9_) & (!n_n518) & (n_n390) & (!n_n534) & (n_n4583)) + ((i_9_) & (!n_n518) & (n_n390) & (n_n534) & (n_n4583)) + ((i_9_) & (n_n518) & (!n_n390) & (!n_n534) & (n_n4583)) + ((i_9_) & (n_n518) & (!n_n390) & (n_n534) & (n_n4583)) + ((i_9_) & (n_n518) & (n_n390) & (!n_n534) & (n_n4583)) + ((i_9_) & (n_n518) & (n_n390) & (n_n534) & (!n_n4583)) + ((i_9_) & (n_n518) & (n_n390) & (n_n534) & (n_n4583)));
	assign x237x = (((!i_9_) & (n_n390) & (n_n535) & (!n_n520) & (x20x)) + ((!i_9_) & (n_n390) & (n_n535) & (n_n520) & (x20x)) + ((i_9_) & (n_n390) & (n_n535) & (!n_n520) & (x20x)) + ((i_9_) & (n_n390) & (n_n535) & (n_n520) & (!x20x)) + ((i_9_) & (n_n390) & (n_n535) & (n_n520) & (x20x)));
	assign n_n2993 = (((!n_n4574) & (!n_n4573) & (!n_n3870) & (!x276x) & (x222x)) + ((!n_n4574) & (!n_n4573) & (!n_n3870) & (x276x) & (!x222x)) + ((!n_n4574) & (!n_n4573) & (!n_n3870) & (x276x) & (x222x)) + ((!n_n4574) & (!n_n4573) & (n_n3870) & (!x276x) & (!x222x)) + ((!n_n4574) & (!n_n4573) & (n_n3870) & (!x276x) & (x222x)) + ((!n_n4574) & (!n_n4573) & (n_n3870) & (x276x) & (!x222x)) + ((!n_n4574) & (!n_n4573) & (n_n3870) & (x276x) & (x222x)) + ((!n_n4574) & (n_n4573) & (!n_n3870) & (!x276x) & (!x222x)) + ((!n_n4574) & (n_n4573) & (!n_n3870) & (!x276x) & (x222x)) + ((!n_n4574) & (n_n4573) & (!n_n3870) & (x276x) & (!x222x)) + ((!n_n4574) & (n_n4573) & (!n_n3870) & (x276x) & (x222x)) + ((!n_n4574) & (n_n4573) & (n_n3870) & (!x276x) & (!x222x)) + ((!n_n4574) & (n_n4573) & (n_n3870) & (!x276x) & (x222x)) + ((!n_n4574) & (n_n4573) & (n_n3870) & (x276x) & (!x222x)) + ((!n_n4574) & (n_n4573) & (n_n3870) & (x276x) & (x222x)) + ((n_n4574) & (!n_n4573) & (!n_n3870) & (!x276x) & (!x222x)) + ((n_n4574) & (!n_n4573) & (!n_n3870) & (!x276x) & (x222x)) + ((n_n4574) & (!n_n4573) & (!n_n3870) & (x276x) & (!x222x)) + ((n_n4574) & (!n_n4573) & (!n_n3870) & (x276x) & (x222x)) + ((n_n4574) & (!n_n4573) & (n_n3870) & (!x276x) & (!x222x)) + ((n_n4574) & (!n_n4573) & (n_n3870) & (!x276x) & (x222x)) + ((n_n4574) & (!n_n4573) & (n_n3870) & (x276x) & (!x222x)) + ((n_n4574) & (!n_n4573) & (n_n3870) & (x276x) & (x222x)) + ((n_n4574) & (n_n4573) & (!n_n3870) & (!x276x) & (!x222x)) + ((n_n4574) & (n_n4573) & (!n_n3870) & (!x276x) & (x222x)) + ((n_n4574) & (n_n4573) & (!n_n3870) & (x276x) & (!x222x)) + ((n_n4574) & (n_n4573) & (!n_n3870) & (x276x) & (x222x)) + ((n_n4574) & (n_n4573) & (n_n3870) & (!x276x) & (!x222x)) + ((n_n4574) & (n_n4573) & (n_n3870) & (!x276x) & (x222x)) + ((n_n4574) & (n_n4573) & (n_n3870) & (x276x) & (!x222x)) + ((n_n4574) & (n_n4573) & (n_n3870) & (x276x) & (x222x)));
	assign x15479x = (((!n_n4587) & (!x365x) & (!n_n4580) & (n_n4585)) + ((!n_n4587) & (!x365x) & (n_n4580) & (!n_n4585)) + ((!n_n4587) & (!x365x) & (n_n4580) & (n_n4585)) + ((!n_n4587) & (x365x) & (!n_n4580) & (!n_n4585)) + ((!n_n4587) & (x365x) & (!n_n4580) & (n_n4585)) + ((!n_n4587) & (x365x) & (n_n4580) & (!n_n4585)) + ((!n_n4587) & (x365x) & (n_n4580) & (n_n4585)) + ((n_n4587) & (!x365x) & (!n_n4580) & (!n_n4585)) + ((n_n4587) & (!x365x) & (!n_n4580) & (n_n4585)) + ((n_n4587) & (!x365x) & (n_n4580) & (!n_n4585)) + ((n_n4587) & (!x365x) & (n_n4580) & (n_n4585)) + ((n_n4587) & (x365x) & (!n_n4580) & (!n_n4585)) + ((n_n4587) & (x365x) & (!n_n4580) & (n_n4585)) + ((n_n4587) & (x365x) & (n_n4580) & (!n_n4585)) + ((n_n4587) & (x365x) & (n_n4580) & (n_n4585)));
	assign x15501x = (((!n_n4554) & (!n_n4555) & (!n_n4559) & (!x214x) & (!x22090x)) + ((!n_n4554) & (!n_n4555) & (!n_n4559) & (x214x) & (!x22090x)) + ((!n_n4554) & (!n_n4555) & (!n_n4559) & (x214x) & (x22090x)) + ((!n_n4554) & (!n_n4555) & (n_n4559) & (!x214x) & (!x22090x)) + ((!n_n4554) & (!n_n4555) & (n_n4559) & (!x214x) & (x22090x)) + ((!n_n4554) & (!n_n4555) & (n_n4559) & (x214x) & (!x22090x)) + ((!n_n4554) & (!n_n4555) & (n_n4559) & (x214x) & (x22090x)) + ((!n_n4554) & (n_n4555) & (!n_n4559) & (!x214x) & (!x22090x)) + ((!n_n4554) & (n_n4555) & (!n_n4559) & (!x214x) & (x22090x)) + ((!n_n4554) & (n_n4555) & (!n_n4559) & (x214x) & (!x22090x)) + ((!n_n4554) & (n_n4555) & (!n_n4559) & (x214x) & (x22090x)) + ((!n_n4554) & (n_n4555) & (n_n4559) & (!x214x) & (!x22090x)) + ((!n_n4554) & (n_n4555) & (n_n4559) & (!x214x) & (x22090x)) + ((!n_n4554) & (n_n4555) & (n_n4559) & (x214x) & (!x22090x)) + ((!n_n4554) & (n_n4555) & (n_n4559) & (x214x) & (x22090x)) + ((n_n4554) & (!n_n4555) & (!n_n4559) & (!x214x) & (!x22090x)) + ((n_n4554) & (!n_n4555) & (!n_n4559) & (!x214x) & (x22090x)) + ((n_n4554) & (!n_n4555) & (!n_n4559) & (x214x) & (!x22090x)) + ((n_n4554) & (!n_n4555) & (!n_n4559) & (x214x) & (x22090x)) + ((n_n4554) & (!n_n4555) & (n_n4559) & (!x214x) & (!x22090x)) + ((n_n4554) & (!n_n4555) & (n_n4559) & (!x214x) & (x22090x)) + ((n_n4554) & (!n_n4555) & (n_n4559) & (x214x) & (!x22090x)) + ((n_n4554) & (!n_n4555) & (n_n4559) & (x214x) & (x22090x)) + ((n_n4554) & (n_n4555) & (!n_n4559) & (!x214x) & (!x22090x)) + ((n_n4554) & (n_n4555) & (!n_n4559) & (!x214x) & (x22090x)) + ((n_n4554) & (n_n4555) & (!n_n4559) & (x214x) & (!x22090x)) + ((n_n4554) & (n_n4555) & (!n_n4559) & (x214x) & (x22090x)) + ((n_n4554) & (n_n4555) & (n_n4559) & (!x214x) & (!x22090x)) + ((n_n4554) & (n_n4555) & (n_n4559) & (!x214x) & (x22090x)) + ((n_n4554) & (n_n4555) & (n_n4559) & (x214x) & (!x22090x)) + ((n_n4554) & (n_n4555) & (n_n4559) & (x214x) & (x22090x)));
	assign x15503x = (((!x100x) & (!x237x) & (!n_n2993) & (!x15479x) & (x15501x)) + ((!x100x) & (!x237x) & (!n_n2993) & (x15479x) & (!x15501x)) + ((!x100x) & (!x237x) & (!n_n2993) & (x15479x) & (x15501x)) + ((!x100x) & (!x237x) & (n_n2993) & (!x15479x) & (!x15501x)) + ((!x100x) & (!x237x) & (n_n2993) & (!x15479x) & (x15501x)) + ((!x100x) & (!x237x) & (n_n2993) & (x15479x) & (!x15501x)) + ((!x100x) & (!x237x) & (n_n2993) & (x15479x) & (x15501x)) + ((!x100x) & (x237x) & (!n_n2993) & (!x15479x) & (!x15501x)) + ((!x100x) & (x237x) & (!n_n2993) & (!x15479x) & (x15501x)) + ((!x100x) & (x237x) & (!n_n2993) & (x15479x) & (!x15501x)) + ((!x100x) & (x237x) & (!n_n2993) & (x15479x) & (x15501x)) + ((!x100x) & (x237x) & (n_n2993) & (!x15479x) & (!x15501x)) + ((!x100x) & (x237x) & (n_n2993) & (!x15479x) & (x15501x)) + ((!x100x) & (x237x) & (n_n2993) & (x15479x) & (!x15501x)) + ((!x100x) & (x237x) & (n_n2993) & (x15479x) & (x15501x)) + ((x100x) & (!x237x) & (!n_n2993) & (!x15479x) & (!x15501x)) + ((x100x) & (!x237x) & (!n_n2993) & (!x15479x) & (x15501x)) + ((x100x) & (!x237x) & (!n_n2993) & (x15479x) & (!x15501x)) + ((x100x) & (!x237x) & (!n_n2993) & (x15479x) & (x15501x)) + ((x100x) & (!x237x) & (n_n2993) & (!x15479x) & (!x15501x)) + ((x100x) & (!x237x) & (n_n2993) & (!x15479x) & (x15501x)) + ((x100x) & (!x237x) & (n_n2993) & (x15479x) & (!x15501x)) + ((x100x) & (!x237x) & (n_n2993) & (x15479x) & (x15501x)) + ((x100x) & (x237x) & (!n_n2993) & (!x15479x) & (!x15501x)) + ((x100x) & (x237x) & (!n_n2993) & (!x15479x) & (x15501x)) + ((x100x) & (x237x) & (!n_n2993) & (x15479x) & (!x15501x)) + ((x100x) & (x237x) & (!n_n2993) & (x15479x) & (x15501x)) + ((x100x) & (x237x) & (n_n2993) & (!x15479x) & (!x15501x)) + ((x100x) & (x237x) & (n_n2993) & (!x15479x) & (x15501x)) + ((x100x) & (x237x) & (n_n2993) & (x15479x) & (!x15501x)) + ((x100x) & (x237x) & (n_n2993) & (x15479x) & (x15501x)));
	assign n_n2990 = (((!n_n4618) & (!n_n4232) & (!n_n4620) & (!x22226x)) + ((!n_n4618) & (!n_n4232) & (n_n4620) & (!x22226x)) + ((!n_n4618) & (!n_n4232) & (n_n4620) & (x22226x)) + ((!n_n4618) & (n_n4232) & (!n_n4620) & (!x22226x)) + ((!n_n4618) & (n_n4232) & (!n_n4620) & (x22226x)) + ((!n_n4618) & (n_n4232) & (n_n4620) & (!x22226x)) + ((!n_n4618) & (n_n4232) & (n_n4620) & (x22226x)) + ((n_n4618) & (!n_n4232) & (!n_n4620) & (!x22226x)) + ((n_n4618) & (!n_n4232) & (!n_n4620) & (x22226x)) + ((n_n4618) & (!n_n4232) & (n_n4620) & (!x22226x)) + ((n_n4618) & (!n_n4232) & (n_n4620) & (x22226x)) + ((n_n4618) & (n_n4232) & (!n_n4620) & (!x22226x)) + ((n_n4618) & (n_n4232) & (!n_n4620) & (x22226x)) + ((n_n4618) & (n_n4232) & (n_n4620) & (!x22226x)) + ((n_n4618) & (n_n4232) & (n_n4620) & (x22226x)));
	assign n_n2991 = (((!n_n4593) & (!n_n4601) & (!n_n4590) & (!n_n4594) & (x15489x)) + ((!n_n4593) & (!n_n4601) & (!n_n4590) & (n_n4594) & (!x15489x)) + ((!n_n4593) & (!n_n4601) & (!n_n4590) & (n_n4594) & (x15489x)) + ((!n_n4593) & (!n_n4601) & (n_n4590) & (!n_n4594) & (!x15489x)) + ((!n_n4593) & (!n_n4601) & (n_n4590) & (!n_n4594) & (x15489x)) + ((!n_n4593) & (!n_n4601) & (n_n4590) & (n_n4594) & (!x15489x)) + ((!n_n4593) & (!n_n4601) & (n_n4590) & (n_n4594) & (x15489x)) + ((!n_n4593) & (n_n4601) & (!n_n4590) & (!n_n4594) & (!x15489x)) + ((!n_n4593) & (n_n4601) & (!n_n4590) & (!n_n4594) & (x15489x)) + ((!n_n4593) & (n_n4601) & (!n_n4590) & (n_n4594) & (!x15489x)) + ((!n_n4593) & (n_n4601) & (!n_n4590) & (n_n4594) & (x15489x)) + ((!n_n4593) & (n_n4601) & (n_n4590) & (!n_n4594) & (!x15489x)) + ((!n_n4593) & (n_n4601) & (n_n4590) & (!n_n4594) & (x15489x)) + ((!n_n4593) & (n_n4601) & (n_n4590) & (n_n4594) & (!x15489x)) + ((!n_n4593) & (n_n4601) & (n_n4590) & (n_n4594) & (x15489x)) + ((n_n4593) & (!n_n4601) & (!n_n4590) & (!n_n4594) & (!x15489x)) + ((n_n4593) & (!n_n4601) & (!n_n4590) & (!n_n4594) & (x15489x)) + ((n_n4593) & (!n_n4601) & (!n_n4590) & (n_n4594) & (!x15489x)) + ((n_n4593) & (!n_n4601) & (!n_n4590) & (n_n4594) & (x15489x)) + ((n_n4593) & (!n_n4601) & (n_n4590) & (!n_n4594) & (!x15489x)) + ((n_n4593) & (!n_n4601) & (n_n4590) & (!n_n4594) & (x15489x)) + ((n_n4593) & (!n_n4601) & (n_n4590) & (n_n4594) & (!x15489x)) + ((n_n4593) & (!n_n4601) & (n_n4590) & (n_n4594) & (x15489x)) + ((n_n4593) & (n_n4601) & (!n_n4590) & (!n_n4594) & (!x15489x)) + ((n_n4593) & (n_n4601) & (!n_n4590) & (!n_n4594) & (x15489x)) + ((n_n4593) & (n_n4601) & (!n_n4590) & (n_n4594) & (!x15489x)) + ((n_n4593) & (n_n4601) & (!n_n4590) & (n_n4594) & (x15489x)) + ((n_n4593) & (n_n4601) & (n_n4590) & (!n_n4594) & (!x15489x)) + ((n_n4593) & (n_n4601) & (n_n4590) & (!n_n4594) & (x15489x)) + ((n_n4593) & (n_n4601) & (n_n4590) & (n_n4594) & (!x15489x)) + ((n_n4593) & (n_n4601) & (n_n4590) & (n_n4594) & (x15489x)));
	assign n_n2926 = (((!n_n2987) & (!x15471x) & (x15470x)) + ((!n_n2987) & (x15471x) & (!x15470x)) + ((!n_n2987) & (x15471x) & (x15470x)) + ((n_n2987) & (!x15471x) & (!x15470x)) + ((n_n2987) & (!x15471x) & (x15470x)) + ((n_n2987) & (x15471x) & (!x15470x)) + ((n_n2987) & (x15471x) & (x15470x)));
	assign x15494x = (((!n_n4628) & (!n_n4629) & (!x190x) & (x15493x)) + ((!n_n4628) & (!n_n4629) & (x190x) & (!x15493x)) + ((!n_n4628) & (!n_n4629) & (x190x) & (x15493x)) + ((!n_n4628) & (n_n4629) & (!x190x) & (!x15493x)) + ((!n_n4628) & (n_n4629) & (!x190x) & (x15493x)) + ((!n_n4628) & (n_n4629) & (x190x) & (!x15493x)) + ((!n_n4628) & (n_n4629) & (x190x) & (x15493x)) + ((n_n4628) & (!n_n4629) & (!x190x) & (!x15493x)) + ((n_n4628) & (!n_n4629) & (!x190x) & (x15493x)) + ((n_n4628) & (!n_n4629) & (x190x) & (!x15493x)) + ((n_n4628) & (!n_n4629) & (x190x) & (x15493x)) + ((n_n4628) & (n_n4629) & (!x190x) & (!x15493x)) + ((n_n4628) & (n_n4629) & (!x190x) & (x15493x)) + ((n_n4628) & (n_n4629) & (x190x) & (!x15493x)) + ((n_n4628) & (n_n4629) & (x190x) & (x15493x)));
	assign n_n3007 = (((!n_n4383) & (!n_n4389) & (!n_n4385) & (!n_n4390) & (x15508x)) + ((!n_n4383) & (!n_n4389) & (!n_n4385) & (n_n4390) & (!x15508x)) + ((!n_n4383) & (!n_n4389) & (!n_n4385) & (n_n4390) & (x15508x)) + ((!n_n4383) & (!n_n4389) & (n_n4385) & (!n_n4390) & (!x15508x)) + ((!n_n4383) & (!n_n4389) & (n_n4385) & (!n_n4390) & (x15508x)) + ((!n_n4383) & (!n_n4389) & (n_n4385) & (n_n4390) & (!x15508x)) + ((!n_n4383) & (!n_n4389) & (n_n4385) & (n_n4390) & (x15508x)) + ((!n_n4383) & (n_n4389) & (!n_n4385) & (!n_n4390) & (!x15508x)) + ((!n_n4383) & (n_n4389) & (!n_n4385) & (!n_n4390) & (x15508x)) + ((!n_n4383) & (n_n4389) & (!n_n4385) & (n_n4390) & (!x15508x)) + ((!n_n4383) & (n_n4389) & (!n_n4385) & (n_n4390) & (x15508x)) + ((!n_n4383) & (n_n4389) & (n_n4385) & (!n_n4390) & (!x15508x)) + ((!n_n4383) & (n_n4389) & (n_n4385) & (!n_n4390) & (x15508x)) + ((!n_n4383) & (n_n4389) & (n_n4385) & (n_n4390) & (!x15508x)) + ((!n_n4383) & (n_n4389) & (n_n4385) & (n_n4390) & (x15508x)) + ((n_n4383) & (!n_n4389) & (!n_n4385) & (!n_n4390) & (!x15508x)) + ((n_n4383) & (!n_n4389) & (!n_n4385) & (!n_n4390) & (x15508x)) + ((n_n4383) & (!n_n4389) & (!n_n4385) & (n_n4390) & (!x15508x)) + ((n_n4383) & (!n_n4389) & (!n_n4385) & (n_n4390) & (x15508x)) + ((n_n4383) & (!n_n4389) & (n_n4385) & (!n_n4390) & (!x15508x)) + ((n_n4383) & (!n_n4389) & (n_n4385) & (!n_n4390) & (x15508x)) + ((n_n4383) & (!n_n4389) & (n_n4385) & (n_n4390) & (!x15508x)) + ((n_n4383) & (!n_n4389) & (n_n4385) & (n_n4390) & (x15508x)) + ((n_n4383) & (n_n4389) & (!n_n4385) & (!n_n4390) & (!x15508x)) + ((n_n4383) & (n_n4389) & (!n_n4385) & (!n_n4390) & (x15508x)) + ((n_n4383) & (n_n4389) & (!n_n4385) & (n_n4390) & (!x15508x)) + ((n_n4383) & (n_n4389) & (!n_n4385) & (n_n4390) & (x15508x)) + ((n_n4383) & (n_n4389) & (n_n4385) & (!n_n4390) & (!x15508x)) + ((n_n4383) & (n_n4389) & (n_n4385) & (!n_n4390) & (x15508x)) + ((n_n4383) & (n_n4389) & (n_n4385) & (n_n4390) & (!x15508x)) + ((n_n4383) & (n_n4389) & (n_n4385) & (n_n4390) & (x15508x)));
	assign x15512x = (((!n_n4362) & (!n_n4366) & (x64x)) + ((!n_n4362) & (n_n4366) & (!x64x)) + ((!n_n4362) & (n_n4366) & (x64x)) + ((n_n4362) & (!n_n4366) & (!x64x)) + ((n_n4362) & (!n_n4366) & (x64x)) + ((n_n4362) & (n_n4366) & (!x64x)) + ((n_n4362) & (n_n4366) & (x64x)));
	assign x15513x = (((!n_n4365) & (!n_n4358) & (!n_n4356) & (!n_n4353) & (n_n4354)) + ((!n_n4365) & (!n_n4358) & (!n_n4356) & (n_n4353) & (!n_n4354)) + ((!n_n4365) & (!n_n4358) & (!n_n4356) & (n_n4353) & (n_n4354)) + ((!n_n4365) & (!n_n4358) & (n_n4356) & (!n_n4353) & (!n_n4354)) + ((!n_n4365) & (!n_n4358) & (n_n4356) & (!n_n4353) & (n_n4354)) + ((!n_n4365) & (!n_n4358) & (n_n4356) & (n_n4353) & (!n_n4354)) + ((!n_n4365) & (!n_n4358) & (n_n4356) & (n_n4353) & (n_n4354)) + ((!n_n4365) & (n_n4358) & (!n_n4356) & (!n_n4353) & (!n_n4354)) + ((!n_n4365) & (n_n4358) & (!n_n4356) & (!n_n4353) & (n_n4354)) + ((!n_n4365) & (n_n4358) & (!n_n4356) & (n_n4353) & (!n_n4354)) + ((!n_n4365) & (n_n4358) & (!n_n4356) & (n_n4353) & (n_n4354)) + ((!n_n4365) & (n_n4358) & (n_n4356) & (!n_n4353) & (!n_n4354)) + ((!n_n4365) & (n_n4358) & (n_n4356) & (!n_n4353) & (n_n4354)) + ((!n_n4365) & (n_n4358) & (n_n4356) & (n_n4353) & (!n_n4354)) + ((!n_n4365) & (n_n4358) & (n_n4356) & (n_n4353) & (n_n4354)) + ((n_n4365) & (!n_n4358) & (!n_n4356) & (!n_n4353) & (!n_n4354)) + ((n_n4365) & (!n_n4358) & (!n_n4356) & (!n_n4353) & (n_n4354)) + ((n_n4365) & (!n_n4358) & (!n_n4356) & (n_n4353) & (!n_n4354)) + ((n_n4365) & (!n_n4358) & (!n_n4356) & (n_n4353) & (n_n4354)) + ((n_n4365) & (!n_n4358) & (n_n4356) & (!n_n4353) & (!n_n4354)) + ((n_n4365) & (!n_n4358) & (n_n4356) & (!n_n4353) & (n_n4354)) + ((n_n4365) & (!n_n4358) & (n_n4356) & (n_n4353) & (!n_n4354)) + ((n_n4365) & (!n_n4358) & (n_n4356) & (n_n4353) & (n_n4354)) + ((n_n4365) & (n_n4358) & (!n_n4356) & (!n_n4353) & (!n_n4354)) + ((n_n4365) & (n_n4358) & (!n_n4356) & (!n_n4353) & (n_n4354)) + ((n_n4365) & (n_n4358) & (!n_n4356) & (n_n4353) & (!n_n4354)) + ((n_n4365) & (n_n4358) & (!n_n4356) & (n_n4353) & (n_n4354)) + ((n_n4365) & (n_n4358) & (n_n4356) & (!n_n4353) & (!n_n4354)) + ((n_n4365) & (n_n4358) & (n_n4356) & (!n_n4353) & (n_n4354)) + ((n_n4365) & (n_n4358) & (n_n4356) & (n_n4353) & (!n_n4354)) + ((n_n4365) & (n_n4358) & (n_n4356) & (n_n4353) & (n_n4354)));
	assign x15547x = (((!n_n4369) & (!n_n4373) & (!n_n4374) & (!n_n3176) & (x27x)) + ((!n_n4369) & (!n_n4373) & (!n_n4374) & (n_n3176) & (!x27x)) + ((!n_n4369) & (!n_n4373) & (!n_n4374) & (n_n3176) & (x27x)) + ((!n_n4369) & (!n_n4373) & (n_n4374) & (!n_n3176) & (!x27x)) + ((!n_n4369) & (!n_n4373) & (n_n4374) & (!n_n3176) & (x27x)) + ((!n_n4369) & (!n_n4373) & (n_n4374) & (n_n3176) & (!x27x)) + ((!n_n4369) & (!n_n4373) & (n_n4374) & (n_n3176) & (x27x)) + ((!n_n4369) & (n_n4373) & (!n_n4374) & (!n_n3176) & (!x27x)) + ((!n_n4369) & (n_n4373) & (!n_n4374) & (!n_n3176) & (x27x)) + ((!n_n4369) & (n_n4373) & (!n_n4374) & (n_n3176) & (!x27x)) + ((!n_n4369) & (n_n4373) & (!n_n4374) & (n_n3176) & (x27x)) + ((!n_n4369) & (n_n4373) & (n_n4374) & (!n_n3176) & (!x27x)) + ((!n_n4369) & (n_n4373) & (n_n4374) & (!n_n3176) & (x27x)) + ((!n_n4369) & (n_n4373) & (n_n4374) & (n_n3176) & (!x27x)) + ((!n_n4369) & (n_n4373) & (n_n4374) & (n_n3176) & (x27x)) + ((n_n4369) & (!n_n4373) & (!n_n4374) & (!n_n3176) & (!x27x)) + ((n_n4369) & (!n_n4373) & (!n_n4374) & (!n_n3176) & (x27x)) + ((n_n4369) & (!n_n4373) & (!n_n4374) & (n_n3176) & (!x27x)) + ((n_n4369) & (!n_n4373) & (!n_n4374) & (n_n3176) & (x27x)) + ((n_n4369) & (!n_n4373) & (n_n4374) & (!n_n3176) & (!x27x)) + ((n_n4369) & (!n_n4373) & (n_n4374) & (!n_n3176) & (x27x)) + ((n_n4369) & (!n_n4373) & (n_n4374) & (n_n3176) & (!x27x)) + ((n_n4369) & (!n_n4373) & (n_n4374) & (n_n3176) & (x27x)) + ((n_n4369) & (n_n4373) & (!n_n4374) & (!n_n3176) & (!x27x)) + ((n_n4369) & (n_n4373) & (!n_n4374) & (!n_n3176) & (x27x)) + ((n_n4369) & (n_n4373) & (!n_n4374) & (n_n3176) & (!x27x)) + ((n_n4369) & (n_n4373) & (!n_n4374) & (n_n3176) & (x27x)) + ((n_n4369) & (n_n4373) & (n_n4374) & (!n_n3176) & (!x27x)) + ((n_n4369) & (n_n4373) & (n_n4374) & (!n_n3176) & (x27x)) + ((n_n4369) & (n_n4373) & (n_n4374) & (n_n3176) & (!x27x)) + ((n_n4369) & (n_n4373) & (n_n4374) & (n_n3176) & (x27x)));
	assign x15549x = (((!n_n3007) & (!x15512x) & (!x15513x) & (x15547x)) + ((!n_n3007) & (!x15512x) & (x15513x) & (!x15547x)) + ((!n_n3007) & (!x15512x) & (x15513x) & (x15547x)) + ((!n_n3007) & (x15512x) & (!x15513x) & (!x15547x)) + ((!n_n3007) & (x15512x) & (!x15513x) & (x15547x)) + ((!n_n3007) & (x15512x) & (x15513x) & (!x15547x)) + ((!n_n3007) & (x15512x) & (x15513x) & (x15547x)) + ((n_n3007) & (!x15512x) & (!x15513x) & (!x15547x)) + ((n_n3007) & (!x15512x) & (!x15513x) & (x15547x)) + ((n_n3007) & (!x15512x) & (x15513x) & (!x15547x)) + ((n_n3007) & (!x15512x) & (x15513x) & (x15547x)) + ((n_n3007) & (x15512x) & (!x15513x) & (!x15547x)) + ((n_n3007) & (x15512x) & (!x15513x) & (x15547x)) + ((n_n3007) & (x15512x) & (x15513x) & (!x15547x)) + ((n_n3007) & (x15512x) & (x15513x) & (x15547x)));
	assign n_n2934 = (((!n_n3010) & (!n_n3012) & (x15527x)) + ((!n_n3010) & (n_n3012) & (!x15527x)) + ((!n_n3010) & (n_n3012) & (x15527x)) + ((n_n3010) & (!n_n3012) & (!x15527x)) + ((n_n3010) & (!n_n3012) & (x15527x)) + ((n_n3010) & (n_n3012) & (!x15527x)) + ((n_n3010) & (n_n3012) & (x15527x)));
	assign n_n3004 = (((!n_n4433) & (!n_n4438) & (!x15531x) & (!x22200x)) + ((!n_n4433) & (!n_n4438) & (x15531x) & (!x22200x)) + ((!n_n4433) & (!n_n4438) & (x15531x) & (x22200x)) + ((!n_n4433) & (n_n4438) & (!x15531x) & (!x22200x)) + ((!n_n4433) & (n_n4438) & (!x15531x) & (x22200x)) + ((!n_n4433) & (n_n4438) & (x15531x) & (!x22200x)) + ((!n_n4433) & (n_n4438) & (x15531x) & (x22200x)) + ((n_n4433) & (!n_n4438) & (!x15531x) & (!x22200x)) + ((n_n4433) & (!n_n4438) & (!x15531x) & (x22200x)) + ((n_n4433) & (!n_n4438) & (x15531x) & (!x22200x)) + ((n_n4433) & (!n_n4438) & (x15531x) & (x22200x)) + ((n_n4433) & (n_n4438) & (!x15531x) & (!x22200x)) + ((n_n4433) & (n_n4438) & (!x15531x) & (x22200x)) + ((n_n4433) & (n_n4438) & (x15531x) & (!x22200x)) + ((n_n4433) & (n_n4438) & (x15531x) & (x22200x)));
	assign n_n3005 = (((!n_n4420) & (!n_n4416) & (!n_n4414) & (!x83x) & (x15536x)) + ((!n_n4420) & (!n_n4416) & (!n_n4414) & (x83x) & (!x15536x)) + ((!n_n4420) & (!n_n4416) & (!n_n4414) & (x83x) & (x15536x)) + ((!n_n4420) & (!n_n4416) & (n_n4414) & (!x83x) & (!x15536x)) + ((!n_n4420) & (!n_n4416) & (n_n4414) & (!x83x) & (x15536x)) + ((!n_n4420) & (!n_n4416) & (n_n4414) & (x83x) & (!x15536x)) + ((!n_n4420) & (!n_n4416) & (n_n4414) & (x83x) & (x15536x)) + ((!n_n4420) & (n_n4416) & (!n_n4414) & (!x83x) & (!x15536x)) + ((!n_n4420) & (n_n4416) & (!n_n4414) & (!x83x) & (x15536x)) + ((!n_n4420) & (n_n4416) & (!n_n4414) & (x83x) & (!x15536x)) + ((!n_n4420) & (n_n4416) & (!n_n4414) & (x83x) & (x15536x)) + ((!n_n4420) & (n_n4416) & (n_n4414) & (!x83x) & (!x15536x)) + ((!n_n4420) & (n_n4416) & (n_n4414) & (!x83x) & (x15536x)) + ((!n_n4420) & (n_n4416) & (n_n4414) & (x83x) & (!x15536x)) + ((!n_n4420) & (n_n4416) & (n_n4414) & (x83x) & (x15536x)) + ((n_n4420) & (!n_n4416) & (!n_n4414) & (!x83x) & (!x15536x)) + ((n_n4420) & (!n_n4416) & (!n_n4414) & (!x83x) & (x15536x)) + ((n_n4420) & (!n_n4416) & (!n_n4414) & (x83x) & (!x15536x)) + ((n_n4420) & (!n_n4416) & (!n_n4414) & (x83x) & (x15536x)) + ((n_n4420) & (!n_n4416) & (n_n4414) & (!x83x) & (!x15536x)) + ((n_n4420) & (!n_n4416) & (n_n4414) & (!x83x) & (x15536x)) + ((n_n4420) & (!n_n4416) & (n_n4414) & (x83x) & (!x15536x)) + ((n_n4420) & (!n_n4416) & (n_n4414) & (x83x) & (x15536x)) + ((n_n4420) & (n_n4416) & (!n_n4414) & (!x83x) & (!x15536x)) + ((n_n4420) & (n_n4416) & (!n_n4414) & (!x83x) & (x15536x)) + ((n_n4420) & (n_n4416) & (!n_n4414) & (x83x) & (!x15536x)) + ((n_n4420) & (n_n4416) & (!n_n4414) & (x83x) & (x15536x)) + ((n_n4420) & (n_n4416) & (n_n4414) & (!x83x) & (!x15536x)) + ((n_n4420) & (n_n4416) & (n_n4414) & (!x83x) & (x15536x)) + ((n_n4420) & (n_n4416) & (n_n4414) & (x83x) & (!x15536x)) + ((n_n4420) & (n_n4416) & (n_n4414) & (x83x) & (x15536x)));
	assign x15543x = (((!n_n4403) & (!n_n4407) & (!n_n4409) & (!n_n4410) & (x15542x)) + ((!n_n4403) & (!n_n4407) & (!n_n4409) & (n_n4410) & (!x15542x)) + ((!n_n4403) & (!n_n4407) & (!n_n4409) & (n_n4410) & (x15542x)) + ((!n_n4403) & (!n_n4407) & (n_n4409) & (!n_n4410) & (!x15542x)) + ((!n_n4403) & (!n_n4407) & (n_n4409) & (!n_n4410) & (x15542x)) + ((!n_n4403) & (!n_n4407) & (n_n4409) & (n_n4410) & (!x15542x)) + ((!n_n4403) & (!n_n4407) & (n_n4409) & (n_n4410) & (x15542x)) + ((!n_n4403) & (n_n4407) & (!n_n4409) & (!n_n4410) & (!x15542x)) + ((!n_n4403) & (n_n4407) & (!n_n4409) & (!n_n4410) & (x15542x)) + ((!n_n4403) & (n_n4407) & (!n_n4409) & (n_n4410) & (!x15542x)) + ((!n_n4403) & (n_n4407) & (!n_n4409) & (n_n4410) & (x15542x)) + ((!n_n4403) & (n_n4407) & (n_n4409) & (!n_n4410) & (!x15542x)) + ((!n_n4403) & (n_n4407) & (n_n4409) & (!n_n4410) & (x15542x)) + ((!n_n4403) & (n_n4407) & (n_n4409) & (n_n4410) & (!x15542x)) + ((!n_n4403) & (n_n4407) & (n_n4409) & (n_n4410) & (x15542x)) + ((n_n4403) & (!n_n4407) & (!n_n4409) & (!n_n4410) & (!x15542x)) + ((n_n4403) & (!n_n4407) & (!n_n4409) & (!n_n4410) & (x15542x)) + ((n_n4403) & (!n_n4407) & (!n_n4409) & (n_n4410) & (!x15542x)) + ((n_n4403) & (!n_n4407) & (!n_n4409) & (n_n4410) & (x15542x)) + ((n_n4403) & (!n_n4407) & (n_n4409) & (!n_n4410) & (!x15542x)) + ((n_n4403) & (!n_n4407) & (n_n4409) & (!n_n4410) & (x15542x)) + ((n_n4403) & (!n_n4407) & (n_n4409) & (n_n4410) & (!x15542x)) + ((n_n4403) & (!n_n4407) & (n_n4409) & (n_n4410) & (x15542x)) + ((n_n4403) & (n_n4407) & (!n_n4409) & (!n_n4410) & (!x15542x)) + ((n_n4403) & (n_n4407) & (!n_n4409) & (!n_n4410) & (x15542x)) + ((n_n4403) & (n_n4407) & (!n_n4409) & (n_n4410) & (!x15542x)) + ((n_n4403) & (n_n4407) & (!n_n4409) & (n_n4410) & (x15542x)) + ((n_n4403) & (n_n4407) & (n_n4409) & (!n_n4410) & (!x15542x)) + ((n_n4403) & (n_n4407) & (n_n4409) & (!n_n4410) & (x15542x)) + ((n_n4403) & (n_n4407) & (n_n4409) & (n_n4410) & (!x15542x)) + ((n_n4403) & (n_n4407) & (n_n4409) & (n_n4410) & (x15542x)));
	assign n_n2915 = (((!x15607x) & (!x15611x) & (!x15618x) & (!x22087x)) + ((!x15607x) & (!x15611x) & (x15618x) & (!x22087x)) + ((!x15607x) & (!x15611x) & (x15618x) & (x22087x)) + ((!x15607x) & (x15611x) & (!x15618x) & (!x22087x)) + ((!x15607x) & (x15611x) & (!x15618x) & (x22087x)) + ((!x15607x) & (x15611x) & (x15618x) & (!x22087x)) + ((!x15607x) & (x15611x) & (x15618x) & (x22087x)) + ((x15607x) & (!x15611x) & (!x15618x) & (!x22087x)) + ((x15607x) & (!x15611x) & (!x15618x) & (x22087x)) + ((x15607x) & (!x15611x) & (x15618x) & (!x22087x)) + ((x15607x) & (!x15611x) & (x15618x) & (x22087x)) + ((x15607x) & (x15611x) & (!x15618x) & (!x22087x)) + ((x15607x) & (x15611x) & (!x15618x) & (x22087x)) + ((x15607x) & (x15611x) & (x15618x) & (!x22087x)) + ((x15607x) & (x15611x) & (x15618x) & (x22087x)));
	assign n_n2952 = (((!n_n5107) & (!n_n5108) & (!n_n5106) & (!x127x) & (!x22086x)) + ((!n_n5107) & (!n_n5108) & (!n_n5106) & (x127x) & (!x22086x)) + ((!n_n5107) & (!n_n5108) & (!n_n5106) & (x127x) & (x22086x)) + ((!n_n5107) & (!n_n5108) & (n_n5106) & (!x127x) & (!x22086x)) + ((!n_n5107) & (!n_n5108) & (n_n5106) & (!x127x) & (x22086x)) + ((!n_n5107) & (!n_n5108) & (n_n5106) & (x127x) & (!x22086x)) + ((!n_n5107) & (!n_n5108) & (n_n5106) & (x127x) & (x22086x)) + ((!n_n5107) & (n_n5108) & (!n_n5106) & (!x127x) & (!x22086x)) + ((!n_n5107) & (n_n5108) & (!n_n5106) & (!x127x) & (x22086x)) + ((!n_n5107) & (n_n5108) & (!n_n5106) & (x127x) & (!x22086x)) + ((!n_n5107) & (n_n5108) & (!n_n5106) & (x127x) & (x22086x)) + ((!n_n5107) & (n_n5108) & (n_n5106) & (!x127x) & (!x22086x)) + ((!n_n5107) & (n_n5108) & (n_n5106) & (!x127x) & (x22086x)) + ((!n_n5107) & (n_n5108) & (n_n5106) & (x127x) & (!x22086x)) + ((!n_n5107) & (n_n5108) & (n_n5106) & (x127x) & (x22086x)) + ((n_n5107) & (!n_n5108) & (!n_n5106) & (!x127x) & (!x22086x)) + ((n_n5107) & (!n_n5108) & (!n_n5106) & (!x127x) & (x22086x)) + ((n_n5107) & (!n_n5108) & (!n_n5106) & (x127x) & (!x22086x)) + ((n_n5107) & (!n_n5108) & (!n_n5106) & (x127x) & (x22086x)) + ((n_n5107) & (!n_n5108) & (n_n5106) & (!x127x) & (!x22086x)) + ((n_n5107) & (!n_n5108) & (n_n5106) & (!x127x) & (x22086x)) + ((n_n5107) & (!n_n5108) & (n_n5106) & (x127x) & (!x22086x)) + ((n_n5107) & (!n_n5108) & (n_n5106) & (x127x) & (x22086x)) + ((n_n5107) & (n_n5108) & (!n_n5106) & (!x127x) & (!x22086x)) + ((n_n5107) & (n_n5108) & (!n_n5106) & (!x127x) & (x22086x)) + ((n_n5107) & (n_n5108) & (!n_n5106) & (x127x) & (!x22086x)) + ((n_n5107) & (n_n5108) & (!n_n5106) & (x127x) & (x22086x)) + ((n_n5107) & (n_n5108) & (n_n5106) & (!x127x) & (!x22086x)) + ((n_n5107) & (n_n5108) & (n_n5106) & (!x127x) & (x22086x)) + ((n_n5107) & (n_n5108) & (n_n5106) & (x127x) & (!x22086x)) + ((n_n5107) & (n_n5108) & (n_n5106) & (x127x) & (x22086x)));
	assign x15633x = (((!n_n5138) & (!n_n5134) & (!n_n3772) & (!n_n3051) & (x15626x)) + ((!n_n5138) & (!n_n5134) & (!n_n3772) & (n_n3051) & (!x15626x)) + ((!n_n5138) & (!n_n5134) & (!n_n3772) & (n_n3051) & (x15626x)) + ((!n_n5138) & (!n_n5134) & (n_n3772) & (!n_n3051) & (!x15626x)) + ((!n_n5138) & (!n_n5134) & (n_n3772) & (!n_n3051) & (x15626x)) + ((!n_n5138) & (!n_n5134) & (n_n3772) & (n_n3051) & (!x15626x)) + ((!n_n5138) & (!n_n5134) & (n_n3772) & (n_n3051) & (x15626x)) + ((!n_n5138) & (n_n5134) & (!n_n3772) & (!n_n3051) & (!x15626x)) + ((!n_n5138) & (n_n5134) & (!n_n3772) & (!n_n3051) & (x15626x)) + ((!n_n5138) & (n_n5134) & (!n_n3772) & (n_n3051) & (!x15626x)) + ((!n_n5138) & (n_n5134) & (!n_n3772) & (n_n3051) & (x15626x)) + ((!n_n5138) & (n_n5134) & (n_n3772) & (!n_n3051) & (!x15626x)) + ((!n_n5138) & (n_n5134) & (n_n3772) & (!n_n3051) & (x15626x)) + ((!n_n5138) & (n_n5134) & (n_n3772) & (n_n3051) & (!x15626x)) + ((!n_n5138) & (n_n5134) & (n_n3772) & (n_n3051) & (x15626x)) + ((n_n5138) & (!n_n5134) & (!n_n3772) & (!n_n3051) & (!x15626x)) + ((n_n5138) & (!n_n5134) & (!n_n3772) & (!n_n3051) & (x15626x)) + ((n_n5138) & (!n_n5134) & (!n_n3772) & (n_n3051) & (!x15626x)) + ((n_n5138) & (!n_n5134) & (!n_n3772) & (n_n3051) & (x15626x)) + ((n_n5138) & (!n_n5134) & (n_n3772) & (!n_n3051) & (!x15626x)) + ((n_n5138) & (!n_n5134) & (n_n3772) & (!n_n3051) & (x15626x)) + ((n_n5138) & (!n_n5134) & (n_n3772) & (n_n3051) & (!x15626x)) + ((n_n5138) & (!n_n5134) & (n_n3772) & (n_n3051) & (x15626x)) + ((n_n5138) & (n_n5134) & (!n_n3772) & (!n_n3051) & (!x15626x)) + ((n_n5138) & (n_n5134) & (!n_n3772) & (!n_n3051) & (x15626x)) + ((n_n5138) & (n_n5134) & (!n_n3772) & (n_n3051) & (!x15626x)) + ((n_n5138) & (n_n5134) & (!n_n3772) & (n_n3051) & (x15626x)) + ((n_n5138) & (n_n5134) & (n_n3772) & (!n_n3051) & (!x15626x)) + ((n_n5138) & (n_n5134) & (n_n3772) & (!n_n3051) & (x15626x)) + ((n_n5138) & (n_n5134) & (n_n3772) & (n_n3051) & (!x15626x)) + ((n_n5138) & (n_n5134) & (n_n3772) & (n_n3051) & (x15626x)));
	assign x15642x = (((!n_n2957) & (!x15602x) & (!x15603x) & (!x15638x) & (x15639x)) + ((!n_n2957) & (!x15602x) & (!x15603x) & (x15638x) & (!x15639x)) + ((!n_n2957) & (!x15602x) & (!x15603x) & (x15638x) & (x15639x)) + ((!n_n2957) & (!x15602x) & (x15603x) & (!x15638x) & (!x15639x)) + ((!n_n2957) & (!x15602x) & (x15603x) & (!x15638x) & (x15639x)) + ((!n_n2957) & (!x15602x) & (x15603x) & (x15638x) & (!x15639x)) + ((!n_n2957) & (!x15602x) & (x15603x) & (x15638x) & (x15639x)) + ((!n_n2957) & (x15602x) & (!x15603x) & (!x15638x) & (!x15639x)) + ((!n_n2957) & (x15602x) & (!x15603x) & (!x15638x) & (x15639x)) + ((!n_n2957) & (x15602x) & (!x15603x) & (x15638x) & (!x15639x)) + ((!n_n2957) & (x15602x) & (!x15603x) & (x15638x) & (x15639x)) + ((!n_n2957) & (x15602x) & (x15603x) & (!x15638x) & (!x15639x)) + ((!n_n2957) & (x15602x) & (x15603x) & (!x15638x) & (x15639x)) + ((!n_n2957) & (x15602x) & (x15603x) & (x15638x) & (!x15639x)) + ((!n_n2957) & (x15602x) & (x15603x) & (x15638x) & (x15639x)) + ((n_n2957) & (!x15602x) & (!x15603x) & (!x15638x) & (!x15639x)) + ((n_n2957) & (!x15602x) & (!x15603x) & (!x15638x) & (x15639x)) + ((n_n2957) & (!x15602x) & (!x15603x) & (x15638x) & (!x15639x)) + ((n_n2957) & (!x15602x) & (!x15603x) & (x15638x) & (x15639x)) + ((n_n2957) & (!x15602x) & (x15603x) & (!x15638x) & (!x15639x)) + ((n_n2957) & (!x15602x) & (x15603x) & (!x15638x) & (x15639x)) + ((n_n2957) & (!x15602x) & (x15603x) & (x15638x) & (!x15639x)) + ((n_n2957) & (!x15602x) & (x15603x) & (x15638x) & (x15639x)) + ((n_n2957) & (x15602x) & (!x15603x) & (!x15638x) & (!x15639x)) + ((n_n2957) & (x15602x) & (!x15603x) & (!x15638x) & (x15639x)) + ((n_n2957) & (x15602x) & (!x15603x) & (x15638x) & (!x15639x)) + ((n_n2957) & (x15602x) & (!x15603x) & (x15638x) & (x15639x)) + ((n_n2957) & (x15602x) & (x15603x) & (!x15638x) & (!x15639x)) + ((n_n2957) & (x15602x) & (x15603x) & (!x15638x) & (x15639x)) + ((n_n2957) & (x15602x) & (x15603x) & (x15638x) & (!x15639x)) + ((n_n2957) & (x15602x) & (x15603x) & (x15638x) & (x15639x)));
	assign x15632x = (((!n_n5136) & (!n_n5124) & (!x335x) & (!x35x) & (x286x)) + ((!n_n5136) & (!n_n5124) & (!x335x) & (x35x) & (!x286x)) + ((!n_n5136) & (!n_n5124) & (!x335x) & (x35x) & (x286x)) + ((!n_n5136) & (!n_n5124) & (x335x) & (!x35x) & (!x286x)) + ((!n_n5136) & (!n_n5124) & (x335x) & (!x35x) & (x286x)) + ((!n_n5136) & (!n_n5124) & (x335x) & (x35x) & (!x286x)) + ((!n_n5136) & (!n_n5124) & (x335x) & (x35x) & (x286x)) + ((!n_n5136) & (n_n5124) & (!x335x) & (!x35x) & (!x286x)) + ((!n_n5136) & (n_n5124) & (!x335x) & (!x35x) & (x286x)) + ((!n_n5136) & (n_n5124) & (!x335x) & (x35x) & (!x286x)) + ((!n_n5136) & (n_n5124) & (!x335x) & (x35x) & (x286x)) + ((!n_n5136) & (n_n5124) & (x335x) & (!x35x) & (!x286x)) + ((!n_n5136) & (n_n5124) & (x335x) & (!x35x) & (x286x)) + ((!n_n5136) & (n_n5124) & (x335x) & (x35x) & (!x286x)) + ((!n_n5136) & (n_n5124) & (x335x) & (x35x) & (x286x)) + ((n_n5136) & (!n_n5124) & (!x335x) & (!x35x) & (!x286x)) + ((n_n5136) & (!n_n5124) & (!x335x) & (!x35x) & (x286x)) + ((n_n5136) & (!n_n5124) & (!x335x) & (x35x) & (!x286x)) + ((n_n5136) & (!n_n5124) & (!x335x) & (x35x) & (x286x)) + ((n_n5136) & (!n_n5124) & (x335x) & (!x35x) & (!x286x)) + ((n_n5136) & (!n_n5124) & (x335x) & (!x35x) & (x286x)) + ((n_n5136) & (!n_n5124) & (x335x) & (x35x) & (!x286x)) + ((n_n5136) & (!n_n5124) & (x335x) & (x35x) & (x286x)) + ((n_n5136) & (n_n5124) & (!x335x) & (!x35x) & (!x286x)) + ((n_n5136) & (n_n5124) & (!x335x) & (!x35x) & (x286x)) + ((n_n5136) & (n_n5124) & (!x335x) & (x35x) & (!x286x)) + ((n_n5136) & (n_n5124) & (!x335x) & (x35x) & (x286x)) + ((n_n5136) & (n_n5124) & (x335x) & (!x35x) & (!x286x)) + ((n_n5136) & (n_n5124) & (x335x) & (!x35x) & (x286x)) + ((n_n5136) & (n_n5124) & (x335x) & (x35x) & (!x286x)) + ((n_n5136) & (n_n5124) & (x335x) & (x35x) & (x286x)));
	assign n_n2912 = (((!x15554x) & (!x15555x) & (!x15564x) & (x15563x)) + ((!x15554x) & (!x15555x) & (x15564x) & (!x15563x)) + ((!x15554x) & (!x15555x) & (x15564x) & (x15563x)) + ((!x15554x) & (x15555x) & (!x15564x) & (!x15563x)) + ((!x15554x) & (x15555x) & (!x15564x) & (x15563x)) + ((!x15554x) & (x15555x) & (x15564x) & (!x15563x)) + ((!x15554x) & (x15555x) & (x15564x) & (x15563x)) + ((x15554x) & (!x15555x) & (!x15564x) & (!x15563x)) + ((x15554x) & (!x15555x) & (!x15564x) & (x15563x)) + ((x15554x) & (!x15555x) & (x15564x) & (!x15563x)) + ((x15554x) & (!x15555x) & (x15564x) & (x15563x)) + ((x15554x) & (x15555x) & (!x15564x) & (!x15563x)) + ((x15554x) & (x15555x) & (!x15564x) & (x15563x)) + ((x15554x) & (x15555x) & (x15564x) & (!x15563x)) + ((x15554x) & (x15555x) & (x15564x) & (x15563x)));
	assign n_n2911 = (((!n_n3031) & (!n_n2943) & (!n_n3385) & (!x15575x) & (x15577x)) + ((!n_n3031) & (!n_n2943) & (!n_n3385) & (x15575x) & (!x15577x)) + ((!n_n3031) & (!n_n2943) & (!n_n3385) & (x15575x) & (x15577x)) + ((!n_n3031) & (!n_n2943) & (n_n3385) & (!x15575x) & (!x15577x)) + ((!n_n3031) & (!n_n2943) & (n_n3385) & (!x15575x) & (x15577x)) + ((!n_n3031) & (!n_n2943) & (n_n3385) & (x15575x) & (!x15577x)) + ((!n_n3031) & (!n_n2943) & (n_n3385) & (x15575x) & (x15577x)) + ((!n_n3031) & (n_n2943) & (!n_n3385) & (!x15575x) & (!x15577x)) + ((!n_n3031) & (n_n2943) & (!n_n3385) & (!x15575x) & (x15577x)) + ((!n_n3031) & (n_n2943) & (!n_n3385) & (x15575x) & (!x15577x)) + ((!n_n3031) & (n_n2943) & (!n_n3385) & (x15575x) & (x15577x)) + ((!n_n3031) & (n_n2943) & (n_n3385) & (!x15575x) & (!x15577x)) + ((!n_n3031) & (n_n2943) & (n_n3385) & (!x15575x) & (x15577x)) + ((!n_n3031) & (n_n2943) & (n_n3385) & (x15575x) & (!x15577x)) + ((!n_n3031) & (n_n2943) & (n_n3385) & (x15575x) & (x15577x)) + ((n_n3031) & (!n_n2943) & (!n_n3385) & (!x15575x) & (!x15577x)) + ((n_n3031) & (!n_n2943) & (!n_n3385) & (!x15575x) & (x15577x)) + ((n_n3031) & (!n_n2943) & (!n_n3385) & (x15575x) & (!x15577x)) + ((n_n3031) & (!n_n2943) & (!n_n3385) & (x15575x) & (x15577x)) + ((n_n3031) & (!n_n2943) & (n_n3385) & (!x15575x) & (!x15577x)) + ((n_n3031) & (!n_n2943) & (n_n3385) & (!x15575x) & (x15577x)) + ((n_n3031) & (!n_n2943) & (n_n3385) & (x15575x) & (!x15577x)) + ((n_n3031) & (!n_n2943) & (n_n3385) & (x15575x) & (x15577x)) + ((n_n3031) & (n_n2943) & (!n_n3385) & (!x15575x) & (!x15577x)) + ((n_n3031) & (n_n2943) & (!n_n3385) & (!x15575x) & (x15577x)) + ((n_n3031) & (n_n2943) & (!n_n3385) & (x15575x) & (!x15577x)) + ((n_n3031) & (n_n2943) & (!n_n3385) & (x15575x) & (x15577x)) + ((n_n3031) & (n_n2943) & (n_n3385) & (!x15575x) & (!x15577x)) + ((n_n3031) & (n_n2943) & (n_n3385) & (!x15575x) & (x15577x)) + ((n_n3031) & (n_n2943) & (n_n3385) & (x15575x) & (!x15577x)) + ((n_n3031) & (n_n2943) & (n_n3385) & (x15575x) & (x15577x)));
	assign x15594x = (((!n_n5179) & (!n_n5173) & (!n_n2948) & (!n_n2949) & (!x22180x)) + ((!n_n5179) & (!n_n5173) & (!n_n2948) & (n_n2949) & (!x22180x)) + ((!n_n5179) & (!n_n5173) & (!n_n2948) & (n_n2949) & (x22180x)) + ((!n_n5179) & (!n_n5173) & (n_n2948) & (!n_n2949) & (!x22180x)) + ((!n_n5179) & (!n_n5173) & (n_n2948) & (!n_n2949) & (x22180x)) + ((!n_n5179) & (!n_n5173) & (n_n2948) & (n_n2949) & (!x22180x)) + ((!n_n5179) & (!n_n5173) & (n_n2948) & (n_n2949) & (x22180x)) + ((!n_n5179) & (n_n5173) & (!n_n2948) & (!n_n2949) & (!x22180x)) + ((!n_n5179) & (n_n5173) & (!n_n2948) & (!n_n2949) & (x22180x)) + ((!n_n5179) & (n_n5173) & (!n_n2948) & (n_n2949) & (!x22180x)) + ((!n_n5179) & (n_n5173) & (!n_n2948) & (n_n2949) & (x22180x)) + ((!n_n5179) & (n_n5173) & (n_n2948) & (!n_n2949) & (!x22180x)) + ((!n_n5179) & (n_n5173) & (n_n2948) & (!n_n2949) & (x22180x)) + ((!n_n5179) & (n_n5173) & (n_n2948) & (n_n2949) & (!x22180x)) + ((!n_n5179) & (n_n5173) & (n_n2948) & (n_n2949) & (x22180x)) + ((n_n5179) & (!n_n5173) & (!n_n2948) & (!n_n2949) & (!x22180x)) + ((n_n5179) & (!n_n5173) & (!n_n2948) & (!n_n2949) & (x22180x)) + ((n_n5179) & (!n_n5173) & (!n_n2948) & (n_n2949) & (!x22180x)) + ((n_n5179) & (!n_n5173) & (!n_n2948) & (n_n2949) & (x22180x)) + ((n_n5179) & (!n_n5173) & (n_n2948) & (!n_n2949) & (!x22180x)) + ((n_n5179) & (!n_n5173) & (n_n2948) & (!n_n2949) & (x22180x)) + ((n_n5179) & (!n_n5173) & (n_n2948) & (n_n2949) & (!x22180x)) + ((n_n5179) & (!n_n5173) & (n_n2948) & (n_n2949) & (x22180x)) + ((n_n5179) & (n_n5173) & (!n_n2948) & (!n_n2949) & (!x22180x)) + ((n_n5179) & (n_n5173) & (!n_n2948) & (!n_n2949) & (x22180x)) + ((n_n5179) & (n_n5173) & (!n_n2948) & (n_n2949) & (!x22180x)) + ((n_n5179) & (n_n5173) & (!n_n2948) & (n_n2949) & (x22180x)) + ((n_n5179) & (n_n5173) & (n_n2948) & (!n_n2949) & (!x22180x)) + ((n_n5179) & (n_n5173) & (n_n2948) & (!n_n2949) & (x22180x)) + ((n_n5179) & (n_n5173) & (n_n2948) & (n_n2949) & (!x22180x)) + ((n_n5179) & (n_n5173) & (n_n2948) & (n_n2949) & (x22180x)));
	assign x15674x = (((!n_n5288) & (!n_n5286) & (!x197x) & (!n_n2937) & (x15668x)) + ((!n_n5288) & (!n_n5286) & (!x197x) & (n_n2937) & (!x15668x)) + ((!n_n5288) & (!n_n5286) & (!x197x) & (n_n2937) & (x15668x)) + ((!n_n5288) & (!n_n5286) & (x197x) & (!n_n2937) & (!x15668x)) + ((!n_n5288) & (!n_n5286) & (x197x) & (!n_n2937) & (x15668x)) + ((!n_n5288) & (!n_n5286) & (x197x) & (n_n2937) & (!x15668x)) + ((!n_n5288) & (!n_n5286) & (x197x) & (n_n2937) & (x15668x)) + ((!n_n5288) & (n_n5286) & (!x197x) & (!n_n2937) & (!x15668x)) + ((!n_n5288) & (n_n5286) & (!x197x) & (!n_n2937) & (x15668x)) + ((!n_n5288) & (n_n5286) & (!x197x) & (n_n2937) & (!x15668x)) + ((!n_n5288) & (n_n5286) & (!x197x) & (n_n2937) & (x15668x)) + ((!n_n5288) & (n_n5286) & (x197x) & (!n_n2937) & (!x15668x)) + ((!n_n5288) & (n_n5286) & (x197x) & (!n_n2937) & (x15668x)) + ((!n_n5288) & (n_n5286) & (x197x) & (n_n2937) & (!x15668x)) + ((!n_n5288) & (n_n5286) & (x197x) & (n_n2937) & (x15668x)) + ((n_n5288) & (!n_n5286) & (!x197x) & (!n_n2937) & (!x15668x)) + ((n_n5288) & (!n_n5286) & (!x197x) & (!n_n2937) & (x15668x)) + ((n_n5288) & (!n_n5286) & (!x197x) & (n_n2937) & (!x15668x)) + ((n_n5288) & (!n_n5286) & (!x197x) & (n_n2937) & (x15668x)) + ((n_n5288) & (!n_n5286) & (x197x) & (!n_n2937) & (!x15668x)) + ((n_n5288) & (!n_n5286) & (x197x) & (!n_n2937) & (x15668x)) + ((n_n5288) & (!n_n5286) & (x197x) & (n_n2937) & (!x15668x)) + ((n_n5288) & (!n_n5286) & (x197x) & (n_n2937) & (x15668x)) + ((n_n5288) & (n_n5286) & (!x197x) & (!n_n2937) & (!x15668x)) + ((n_n5288) & (n_n5286) & (!x197x) & (!n_n2937) & (x15668x)) + ((n_n5288) & (n_n5286) & (!x197x) & (n_n2937) & (!x15668x)) + ((n_n5288) & (n_n5286) & (!x197x) & (n_n2937) & (x15668x)) + ((n_n5288) & (n_n5286) & (x197x) & (!n_n2937) & (!x15668x)) + ((n_n5288) & (n_n5286) & (x197x) & (!n_n2937) & (x15668x)) + ((n_n5288) & (n_n5286) & (x197x) & (n_n2937) & (!x15668x)) + ((n_n5288) & (n_n5286) & (x197x) & (n_n2937) & (x15668x)));
	assign x15675x = (((!x15649x) & (!x15650x) & (!n_n2939) & (!n_n2940) & (x15671x)) + ((!x15649x) & (!x15650x) & (!n_n2939) & (n_n2940) & (!x15671x)) + ((!x15649x) & (!x15650x) & (!n_n2939) & (n_n2940) & (x15671x)) + ((!x15649x) & (!x15650x) & (n_n2939) & (!n_n2940) & (!x15671x)) + ((!x15649x) & (!x15650x) & (n_n2939) & (!n_n2940) & (x15671x)) + ((!x15649x) & (!x15650x) & (n_n2939) & (n_n2940) & (!x15671x)) + ((!x15649x) & (!x15650x) & (n_n2939) & (n_n2940) & (x15671x)) + ((!x15649x) & (x15650x) & (!n_n2939) & (!n_n2940) & (!x15671x)) + ((!x15649x) & (x15650x) & (!n_n2939) & (!n_n2940) & (x15671x)) + ((!x15649x) & (x15650x) & (!n_n2939) & (n_n2940) & (!x15671x)) + ((!x15649x) & (x15650x) & (!n_n2939) & (n_n2940) & (x15671x)) + ((!x15649x) & (x15650x) & (n_n2939) & (!n_n2940) & (!x15671x)) + ((!x15649x) & (x15650x) & (n_n2939) & (!n_n2940) & (x15671x)) + ((!x15649x) & (x15650x) & (n_n2939) & (n_n2940) & (!x15671x)) + ((!x15649x) & (x15650x) & (n_n2939) & (n_n2940) & (x15671x)) + ((x15649x) & (!x15650x) & (!n_n2939) & (!n_n2940) & (!x15671x)) + ((x15649x) & (!x15650x) & (!n_n2939) & (!n_n2940) & (x15671x)) + ((x15649x) & (!x15650x) & (!n_n2939) & (n_n2940) & (!x15671x)) + ((x15649x) & (!x15650x) & (!n_n2939) & (n_n2940) & (x15671x)) + ((x15649x) & (!x15650x) & (n_n2939) & (!n_n2940) & (!x15671x)) + ((x15649x) & (!x15650x) & (n_n2939) & (!n_n2940) & (x15671x)) + ((x15649x) & (!x15650x) & (n_n2939) & (n_n2940) & (!x15671x)) + ((x15649x) & (!x15650x) & (n_n2939) & (n_n2940) & (x15671x)) + ((x15649x) & (x15650x) & (!n_n2939) & (!n_n2940) & (!x15671x)) + ((x15649x) & (x15650x) & (!n_n2939) & (!n_n2940) & (x15671x)) + ((x15649x) & (x15650x) & (!n_n2939) & (n_n2940) & (!x15671x)) + ((x15649x) & (x15650x) & (!n_n2939) & (n_n2940) & (x15671x)) + ((x15649x) & (x15650x) & (n_n2939) & (!n_n2940) & (!x15671x)) + ((x15649x) & (x15650x) & (n_n2939) & (!n_n2940) & (x15671x)) + ((x15649x) & (x15650x) & (n_n2939) & (n_n2940) & (!x15671x)) + ((x15649x) & (x15650x) & (n_n2939) & (n_n2940) & (x15671x)));
	assign n_n2921 = (((!n_n3460) & (!n_n3820) & (!n_n2973) & (!x15693x) & (x15695x)) + ((!n_n3460) & (!n_n3820) & (!n_n2973) & (x15693x) & (!x15695x)) + ((!n_n3460) & (!n_n3820) & (!n_n2973) & (x15693x) & (x15695x)) + ((!n_n3460) & (!n_n3820) & (n_n2973) & (!x15693x) & (!x15695x)) + ((!n_n3460) & (!n_n3820) & (n_n2973) & (!x15693x) & (x15695x)) + ((!n_n3460) & (!n_n3820) & (n_n2973) & (x15693x) & (!x15695x)) + ((!n_n3460) & (!n_n3820) & (n_n2973) & (x15693x) & (x15695x)) + ((!n_n3460) & (n_n3820) & (!n_n2973) & (!x15693x) & (!x15695x)) + ((!n_n3460) & (n_n3820) & (!n_n2973) & (!x15693x) & (x15695x)) + ((!n_n3460) & (n_n3820) & (!n_n2973) & (x15693x) & (!x15695x)) + ((!n_n3460) & (n_n3820) & (!n_n2973) & (x15693x) & (x15695x)) + ((!n_n3460) & (n_n3820) & (n_n2973) & (!x15693x) & (!x15695x)) + ((!n_n3460) & (n_n3820) & (n_n2973) & (!x15693x) & (x15695x)) + ((!n_n3460) & (n_n3820) & (n_n2973) & (x15693x) & (!x15695x)) + ((!n_n3460) & (n_n3820) & (n_n2973) & (x15693x) & (x15695x)) + ((n_n3460) & (!n_n3820) & (!n_n2973) & (!x15693x) & (!x15695x)) + ((n_n3460) & (!n_n3820) & (!n_n2973) & (!x15693x) & (x15695x)) + ((n_n3460) & (!n_n3820) & (!n_n2973) & (x15693x) & (!x15695x)) + ((n_n3460) & (!n_n3820) & (!n_n2973) & (x15693x) & (x15695x)) + ((n_n3460) & (!n_n3820) & (n_n2973) & (!x15693x) & (!x15695x)) + ((n_n3460) & (!n_n3820) & (n_n2973) & (!x15693x) & (x15695x)) + ((n_n3460) & (!n_n3820) & (n_n2973) & (x15693x) & (!x15695x)) + ((n_n3460) & (!n_n3820) & (n_n2973) & (x15693x) & (x15695x)) + ((n_n3460) & (n_n3820) & (!n_n2973) & (!x15693x) & (!x15695x)) + ((n_n3460) & (n_n3820) & (!n_n2973) & (!x15693x) & (x15695x)) + ((n_n3460) & (n_n3820) & (!n_n2973) & (x15693x) & (!x15695x)) + ((n_n3460) & (n_n3820) & (!n_n2973) & (x15693x) & (x15695x)) + ((n_n3460) & (n_n3820) & (n_n2973) & (!x15693x) & (!x15695x)) + ((n_n3460) & (n_n3820) & (n_n2973) & (!x15693x) & (x15695x)) + ((n_n3460) & (n_n3820) & (n_n2973) & (x15693x) & (!x15695x)) + ((n_n3460) & (n_n3820) & (n_n2973) & (x15693x) & (x15695x)));
	assign n_n2903 = (((!n_n2966) & (!n_n2917) & (!n_n2918) & (!n_n2965) & (x15740x)) + ((!n_n2966) & (!n_n2917) & (!n_n2918) & (n_n2965) & (!x15740x)) + ((!n_n2966) & (!n_n2917) & (!n_n2918) & (n_n2965) & (x15740x)) + ((!n_n2966) & (!n_n2917) & (n_n2918) & (!n_n2965) & (!x15740x)) + ((!n_n2966) & (!n_n2917) & (n_n2918) & (!n_n2965) & (x15740x)) + ((!n_n2966) & (!n_n2917) & (n_n2918) & (n_n2965) & (!x15740x)) + ((!n_n2966) & (!n_n2917) & (n_n2918) & (n_n2965) & (x15740x)) + ((!n_n2966) & (n_n2917) & (!n_n2918) & (!n_n2965) & (!x15740x)) + ((!n_n2966) & (n_n2917) & (!n_n2918) & (!n_n2965) & (x15740x)) + ((!n_n2966) & (n_n2917) & (!n_n2918) & (n_n2965) & (!x15740x)) + ((!n_n2966) & (n_n2917) & (!n_n2918) & (n_n2965) & (x15740x)) + ((!n_n2966) & (n_n2917) & (n_n2918) & (!n_n2965) & (!x15740x)) + ((!n_n2966) & (n_n2917) & (n_n2918) & (!n_n2965) & (x15740x)) + ((!n_n2966) & (n_n2917) & (n_n2918) & (n_n2965) & (!x15740x)) + ((!n_n2966) & (n_n2917) & (n_n2918) & (n_n2965) & (x15740x)) + ((n_n2966) & (!n_n2917) & (!n_n2918) & (!n_n2965) & (!x15740x)) + ((n_n2966) & (!n_n2917) & (!n_n2918) & (!n_n2965) & (x15740x)) + ((n_n2966) & (!n_n2917) & (!n_n2918) & (n_n2965) & (!x15740x)) + ((n_n2966) & (!n_n2917) & (!n_n2918) & (n_n2965) & (x15740x)) + ((n_n2966) & (!n_n2917) & (n_n2918) & (!n_n2965) & (!x15740x)) + ((n_n2966) & (!n_n2917) & (n_n2918) & (!n_n2965) & (x15740x)) + ((n_n2966) & (!n_n2917) & (n_n2918) & (n_n2965) & (!x15740x)) + ((n_n2966) & (!n_n2917) & (n_n2918) & (n_n2965) & (x15740x)) + ((n_n2966) & (n_n2917) & (!n_n2918) & (!n_n2965) & (!x15740x)) + ((n_n2966) & (n_n2917) & (!n_n2918) & (!n_n2965) & (x15740x)) + ((n_n2966) & (n_n2917) & (!n_n2918) & (n_n2965) & (!x15740x)) + ((n_n2966) & (n_n2917) & (!n_n2918) & (n_n2965) & (x15740x)) + ((n_n2966) & (n_n2917) & (n_n2918) & (!n_n2965) & (!x15740x)) + ((n_n2966) & (n_n2917) & (n_n2918) & (!n_n2965) & (x15740x)) + ((n_n2966) & (n_n2917) & (n_n2918) & (n_n2965) & (!x15740x)) + ((n_n2966) & (n_n2917) & (n_n2918) & (n_n2965) & (x15740x)));
	assign n_n2905 = (((!n_n2977) & (!n_n2979) & (!x15766x) & (!n_n2925) & (x15786x)) + ((!n_n2977) & (!n_n2979) & (!x15766x) & (n_n2925) & (!x15786x)) + ((!n_n2977) & (!n_n2979) & (!x15766x) & (n_n2925) & (x15786x)) + ((!n_n2977) & (!n_n2979) & (x15766x) & (!n_n2925) & (!x15786x)) + ((!n_n2977) & (!n_n2979) & (x15766x) & (!n_n2925) & (x15786x)) + ((!n_n2977) & (!n_n2979) & (x15766x) & (n_n2925) & (!x15786x)) + ((!n_n2977) & (!n_n2979) & (x15766x) & (n_n2925) & (x15786x)) + ((!n_n2977) & (n_n2979) & (!x15766x) & (!n_n2925) & (!x15786x)) + ((!n_n2977) & (n_n2979) & (!x15766x) & (!n_n2925) & (x15786x)) + ((!n_n2977) & (n_n2979) & (!x15766x) & (n_n2925) & (!x15786x)) + ((!n_n2977) & (n_n2979) & (!x15766x) & (n_n2925) & (x15786x)) + ((!n_n2977) & (n_n2979) & (x15766x) & (!n_n2925) & (!x15786x)) + ((!n_n2977) & (n_n2979) & (x15766x) & (!n_n2925) & (x15786x)) + ((!n_n2977) & (n_n2979) & (x15766x) & (n_n2925) & (!x15786x)) + ((!n_n2977) & (n_n2979) & (x15766x) & (n_n2925) & (x15786x)) + ((n_n2977) & (!n_n2979) & (!x15766x) & (!n_n2925) & (!x15786x)) + ((n_n2977) & (!n_n2979) & (!x15766x) & (!n_n2925) & (x15786x)) + ((n_n2977) & (!n_n2979) & (!x15766x) & (n_n2925) & (!x15786x)) + ((n_n2977) & (!n_n2979) & (!x15766x) & (n_n2925) & (x15786x)) + ((n_n2977) & (!n_n2979) & (x15766x) & (!n_n2925) & (!x15786x)) + ((n_n2977) & (!n_n2979) & (x15766x) & (!n_n2925) & (x15786x)) + ((n_n2977) & (!n_n2979) & (x15766x) & (n_n2925) & (!x15786x)) + ((n_n2977) & (!n_n2979) & (x15766x) & (n_n2925) & (x15786x)) + ((n_n2977) & (n_n2979) & (!x15766x) & (!n_n2925) & (!x15786x)) + ((n_n2977) & (n_n2979) & (!x15766x) & (!n_n2925) & (x15786x)) + ((n_n2977) & (n_n2979) & (!x15766x) & (n_n2925) & (!x15786x)) + ((n_n2977) & (n_n2979) & (!x15766x) & (n_n2925) & (x15786x)) + ((n_n2977) & (n_n2979) & (x15766x) & (!n_n2925) & (!x15786x)) + ((n_n2977) & (n_n2979) & (x15766x) & (!n_n2925) & (x15786x)) + ((n_n2977) & (n_n2979) & (x15766x) & (n_n2925) & (!x15786x)) + ((n_n2977) & (n_n2979) & (x15766x) & (n_n2925) & (x15786x)));
	assign n_n2922 = (((!x158x) & (!x380x) & (!x15791x) & (!x15798x) & (x15797x)) + ((!x158x) & (!x380x) & (!x15791x) & (x15798x) & (!x15797x)) + ((!x158x) & (!x380x) & (!x15791x) & (x15798x) & (x15797x)) + ((!x158x) & (!x380x) & (x15791x) & (!x15798x) & (!x15797x)) + ((!x158x) & (!x380x) & (x15791x) & (!x15798x) & (x15797x)) + ((!x158x) & (!x380x) & (x15791x) & (x15798x) & (!x15797x)) + ((!x158x) & (!x380x) & (x15791x) & (x15798x) & (x15797x)) + ((!x158x) & (x380x) & (!x15791x) & (!x15798x) & (!x15797x)) + ((!x158x) & (x380x) & (!x15791x) & (!x15798x) & (x15797x)) + ((!x158x) & (x380x) & (!x15791x) & (x15798x) & (!x15797x)) + ((!x158x) & (x380x) & (!x15791x) & (x15798x) & (x15797x)) + ((!x158x) & (x380x) & (x15791x) & (!x15798x) & (!x15797x)) + ((!x158x) & (x380x) & (x15791x) & (!x15798x) & (x15797x)) + ((!x158x) & (x380x) & (x15791x) & (x15798x) & (!x15797x)) + ((!x158x) & (x380x) & (x15791x) & (x15798x) & (x15797x)) + ((x158x) & (!x380x) & (!x15791x) & (!x15798x) & (!x15797x)) + ((x158x) & (!x380x) & (!x15791x) & (!x15798x) & (x15797x)) + ((x158x) & (!x380x) & (!x15791x) & (x15798x) & (!x15797x)) + ((x158x) & (!x380x) & (!x15791x) & (x15798x) & (x15797x)) + ((x158x) & (!x380x) & (x15791x) & (!x15798x) & (!x15797x)) + ((x158x) & (!x380x) & (x15791x) & (!x15798x) & (x15797x)) + ((x158x) & (!x380x) & (x15791x) & (x15798x) & (!x15797x)) + ((x158x) & (!x380x) & (x15791x) & (x15798x) & (x15797x)) + ((x158x) & (x380x) & (!x15791x) & (!x15798x) & (!x15797x)) + ((x158x) & (x380x) & (!x15791x) & (!x15798x) & (x15797x)) + ((x158x) & (x380x) & (!x15791x) & (x15798x) & (!x15797x)) + ((x158x) & (x380x) & (!x15791x) & (x15798x) & (x15797x)) + ((x158x) & (x380x) & (x15791x) & (!x15798x) & (!x15797x)) + ((x158x) & (x380x) & (x15791x) & (!x15798x) & (x15797x)) + ((x158x) & (x380x) & (x15791x) & (x15798x) & (!x15797x)) + ((x158x) & (x380x) & (x15791x) & (x15798x) & (x15797x)));
	assign x15806x = (((!n_n2970) & (!n_n2968) & (!x15802x) & (x15803x)) + ((!n_n2970) & (!n_n2968) & (x15802x) & (!x15803x)) + ((!n_n2970) & (!n_n2968) & (x15802x) & (x15803x)) + ((!n_n2970) & (n_n2968) & (!x15802x) & (!x15803x)) + ((!n_n2970) & (n_n2968) & (!x15802x) & (x15803x)) + ((!n_n2970) & (n_n2968) & (x15802x) & (!x15803x)) + ((!n_n2970) & (n_n2968) & (x15802x) & (x15803x)) + ((n_n2970) & (!n_n2968) & (!x15802x) & (!x15803x)) + ((n_n2970) & (!n_n2968) & (!x15802x) & (x15803x)) + ((n_n2970) & (!n_n2968) & (x15802x) & (!x15803x)) + ((n_n2970) & (!n_n2968) & (x15802x) & (x15803x)) + ((n_n2970) & (n_n2968) & (!x15802x) & (!x15803x)) + ((n_n2970) & (n_n2968) & (!x15802x) & (x15803x)) + ((n_n2970) & (n_n2968) & (x15802x) & (!x15803x)) + ((n_n2970) & (n_n2968) & (x15802x) & (x15803x)));
	assign n_n1709 = (((!x15887x) & (!x15871x) & (!x15872x) & (n_n1717)) + ((!x15887x) & (!x15871x) & (x15872x) & (!n_n1717)) + ((!x15887x) & (!x15871x) & (x15872x) & (n_n1717)) + ((!x15887x) & (x15871x) & (!x15872x) & (!n_n1717)) + ((!x15887x) & (x15871x) & (!x15872x) & (n_n1717)) + ((!x15887x) & (x15871x) & (x15872x) & (!n_n1717)) + ((!x15887x) & (x15871x) & (x15872x) & (n_n1717)) + ((x15887x) & (!x15871x) & (!x15872x) & (!n_n1717)) + ((x15887x) & (!x15871x) & (!x15872x) & (n_n1717)) + ((x15887x) & (!x15871x) & (x15872x) & (!n_n1717)) + ((x15887x) & (!x15871x) & (x15872x) & (n_n1717)) + ((x15887x) & (x15871x) & (!x15872x) & (!n_n1717)) + ((x15887x) & (x15871x) & (!x15872x) & (n_n1717)) + ((x15887x) & (x15871x) & (x15872x) & (!n_n1717)) + ((x15887x) & (x15871x) & (x15872x) & (n_n1717)));
	assign x15899x = (((!x15845x) & (!x15846x) & (x15898x)) + ((!x15845x) & (x15846x) & (!x15898x)) + ((!x15845x) & (x15846x) & (x15898x)) + ((x15845x) & (!x15846x) & (!x15898x)) + ((x15845x) & (!x15846x) & (x15898x)) + ((x15845x) & (x15846x) & (!x15898x)) + ((x15845x) & (x15846x) & (x15898x)));
	assign x15900x = (((!x15852x) & (!x15853x) & (!x15859x) & (x15860x)) + ((!x15852x) & (!x15853x) & (x15859x) & (!x15860x)) + ((!x15852x) & (!x15853x) & (x15859x) & (x15860x)) + ((!x15852x) & (x15853x) & (!x15859x) & (!x15860x)) + ((!x15852x) & (x15853x) & (!x15859x) & (x15860x)) + ((!x15852x) & (x15853x) & (x15859x) & (!x15860x)) + ((!x15852x) & (x15853x) & (x15859x) & (x15860x)) + ((x15852x) & (!x15853x) & (!x15859x) & (!x15860x)) + ((x15852x) & (!x15853x) & (!x15859x) & (x15860x)) + ((x15852x) & (!x15853x) & (x15859x) & (!x15860x)) + ((x15852x) & (!x15853x) & (x15859x) & (x15860x)) + ((x15852x) & (x15853x) & (!x15859x) & (!x15860x)) + ((x15852x) & (x15853x) & (!x15859x) & (x15860x)) + ((x15852x) & (x15853x) & (x15859x) & (!x15860x)) + ((x15852x) & (x15853x) & (x15859x) & (x15860x)));
	assign x15901x = (((!n_n1720) & (!x15894x) & (x15895x)) + ((!n_n1720) & (x15894x) & (!x15895x)) + ((!n_n1720) & (x15894x) & (x15895x)) + ((n_n1720) & (!x15894x) & (!x15895x)) + ((n_n1720) & (!x15894x) & (x15895x)) + ((n_n1720) & (x15894x) & (!x15895x)) + ((n_n1720) & (x15894x) & (x15895x)));
	assign n_n1712 = (((!x15838x) & (!x15823x) & (!x15824x) & (!x15829x) & (x15830x)) + ((!x15838x) & (!x15823x) & (!x15824x) & (x15829x) & (!x15830x)) + ((!x15838x) & (!x15823x) & (!x15824x) & (x15829x) & (x15830x)) + ((!x15838x) & (!x15823x) & (x15824x) & (!x15829x) & (!x15830x)) + ((!x15838x) & (!x15823x) & (x15824x) & (!x15829x) & (x15830x)) + ((!x15838x) & (!x15823x) & (x15824x) & (x15829x) & (!x15830x)) + ((!x15838x) & (!x15823x) & (x15824x) & (x15829x) & (x15830x)) + ((!x15838x) & (x15823x) & (!x15824x) & (!x15829x) & (!x15830x)) + ((!x15838x) & (x15823x) & (!x15824x) & (!x15829x) & (x15830x)) + ((!x15838x) & (x15823x) & (!x15824x) & (x15829x) & (!x15830x)) + ((!x15838x) & (x15823x) & (!x15824x) & (x15829x) & (x15830x)) + ((!x15838x) & (x15823x) & (x15824x) & (!x15829x) & (!x15830x)) + ((!x15838x) & (x15823x) & (x15824x) & (!x15829x) & (x15830x)) + ((!x15838x) & (x15823x) & (x15824x) & (x15829x) & (!x15830x)) + ((!x15838x) & (x15823x) & (x15824x) & (x15829x) & (x15830x)) + ((x15838x) & (!x15823x) & (!x15824x) & (!x15829x) & (!x15830x)) + ((x15838x) & (!x15823x) & (!x15824x) & (!x15829x) & (x15830x)) + ((x15838x) & (!x15823x) & (!x15824x) & (x15829x) & (!x15830x)) + ((x15838x) & (!x15823x) & (!x15824x) & (x15829x) & (x15830x)) + ((x15838x) & (!x15823x) & (x15824x) & (!x15829x) & (!x15830x)) + ((x15838x) & (!x15823x) & (x15824x) & (!x15829x) & (x15830x)) + ((x15838x) & (!x15823x) & (x15824x) & (x15829x) & (!x15830x)) + ((x15838x) & (!x15823x) & (x15824x) & (x15829x) & (x15830x)) + ((x15838x) & (x15823x) & (!x15824x) & (!x15829x) & (!x15830x)) + ((x15838x) & (x15823x) & (!x15824x) & (!x15829x) & (x15830x)) + ((x15838x) & (x15823x) & (!x15824x) & (x15829x) & (!x15830x)) + ((x15838x) & (x15823x) & (!x15824x) & (x15829x) & (x15830x)) + ((x15838x) & (x15823x) & (x15824x) & (!x15829x) & (!x15830x)) + ((x15838x) & (x15823x) & (x15824x) & (!x15829x) & (x15830x)) + ((x15838x) & (x15823x) & (x15824x) & (x15829x) & (!x15830x)) + ((x15838x) & (x15823x) & (x15824x) & (x15829x) & (x15830x)));
	assign n_n1711 = (((!x15932x) & (!x15920x) & (!x15921x) & (!x15924x) & (x15925x)) + ((!x15932x) & (!x15920x) & (!x15921x) & (x15924x) & (!x15925x)) + ((!x15932x) & (!x15920x) & (!x15921x) & (x15924x) & (x15925x)) + ((!x15932x) & (!x15920x) & (x15921x) & (!x15924x) & (!x15925x)) + ((!x15932x) & (!x15920x) & (x15921x) & (!x15924x) & (x15925x)) + ((!x15932x) & (!x15920x) & (x15921x) & (x15924x) & (!x15925x)) + ((!x15932x) & (!x15920x) & (x15921x) & (x15924x) & (x15925x)) + ((!x15932x) & (x15920x) & (!x15921x) & (!x15924x) & (!x15925x)) + ((!x15932x) & (x15920x) & (!x15921x) & (!x15924x) & (x15925x)) + ((!x15932x) & (x15920x) & (!x15921x) & (x15924x) & (!x15925x)) + ((!x15932x) & (x15920x) & (!x15921x) & (x15924x) & (x15925x)) + ((!x15932x) & (x15920x) & (x15921x) & (!x15924x) & (!x15925x)) + ((!x15932x) & (x15920x) & (x15921x) & (!x15924x) & (x15925x)) + ((!x15932x) & (x15920x) & (x15921x) & (x15924x) & (!x15925x)) + ((!x15932x) & (x15920x) & (x15921x) & (x15924x) & (x15925x)) + ((x15932x) & (!x15920x) & (!x15921x) & (!x15924x) & (!x15925x)) + ((x15932x) & (!x15920x) & (!x15921x) & (!x15924x) & (x15925x)) + ((x15932x) & (!x15920x) & (!x15921x) & (x15924x) & (!x15925x)) + ((x15932x) & (!x15920x) & (!x15921x) & (x15924x) & (x15925x)) + ((x15932x) & (!x15920x) & (x15921x) & (!x15924x) & (!x15925x)) + ((x15932x) & (!x15920x) & (x15921x) & (!x15924x) & (x15925x)) + ((x15932x) & (!x15920x) & (x15921x) & (x15924x) & (!x15925x)) + ((x15932x) & (!x15920x) & (x15921x) & (x15924x) & (x15925x)) + ((x15932x) & (x15920x) & (!x15921x) & (!x15924x) & (!x15925x)) + ((x15932x) & (x15920x) & (!x15921x) & (!x15924x) & (x15925x)) + ((x15932x) & (x15920x) & (!x15921x) & (x15924x) & (!x15925x)) + ((x15932x) & (x15920x) & (!x15921x) & (x15924x) & (x15925x)) + ((x15932x) & (x15920x) & (x15921x) & (!x15924x) & (!x15925x)) + ((x15932x) & (x15920x) & (x15921x) & (!x15924x) & (x15925x)) + ((x15932x) & (x15920x) & (x15921x) & (x15924x) & (!x15925x)) + ((x15932x) & (x15920x) & (x15921x) & (x15924x) & (x15925x)));
	assign x15939x = (((!n_n4337) & (!n_n4314) & (!x337x) & (x15938x)) + ((!n_n4337) & (!n_n4314) & (x337x) & (!x15938x)) + ((!n_n4337) & (!n_n4314) & (x337x) & (x15938x)) + ((!n_n4337) & (n_n4314) & (!x337x) & (!x15938x)) + ((!n_n4337) & (n_n4314) & (!x337x) & (x15938x)) + ((!n_n4337) & (n_n4314) & (x337x) & (!x15938x)) + ((!n_n4337) & (n_n4314) & (x337x) & (x15938x)) + ((n_n4337) & (!n_n4314) & (!x337x) & (!x15938x)) + ((n_n4337) & (!n_n4314) & (!x337x) & (x15938x)) + ((n_n4337) & (!n_n4314) & (x337x) & (!x15938x)) + ((n_n4337) & (!n_n4314) & (x337x) & (x15938x)) + ((n_n4337) & (n_n4314) & (!x337x) & (!x15938x)) + ((n_n4337) & (n_n4314) & (!x337x) & (x15938x)) + ((n_n4337) & (n_n4314) & (x337x) & (!x15938x)) + ((n_n4337) & (n_n4314) & (x337x) & (x15938x)));
	assign x15940x = (((!x15909x) & (!x15910x) & (!x15915x) & (x15916x)) + ((!x15909x) & (!x15910x) & (x15915x) & (!x15916x)) + ((!x15909x) & (!x15910x) & (x15915x) & (x15916x)) + ((!x15909x) & (x15910x) & (!x15915x) & (!x15916x)) + ((!x15909x) & (x15910x) & (!x15915x) & (x15916x)) + ((!x15909x) & (x15910x) & (x15915x) & (!x15916x)) + ((!x15909x) & (x15910x) & (x15915x) & (x15916x)) + ((x15909x) & (!x15910x) & (!x15915x) & (!x15916x)) + ((x15909x) & (!x15910x) & (!x15915x) & (x15916x)) + ((x15909x) & (!x15910x) & (x15915x) & (!x15916x)) + ((x15909x) & (!x15910x) & (x15915x) & (x15916x)) + ((x15909x) & (x15910x) & (!x15915x) & (!x15916x)) + ((x15909x) & (x15910x) & (!x15915x) & (x15916x)) + ((x15909x) & (x15910x) & (x15915x) & (!x15916x)) + ((x15909x) & (x15910x) & (x15915x) & (x15916x)));
	assign x15978x = (((!n_n524) & (!n_n482) & (!n_n528) & (!x18x) & (x97x)) + ((!n_n524) & (!n_n482) & (!n_n528) & (x18x) & (x97x)) + ((!n_n524) & (!n_n482) & (n_n528) & (!x18x) & (x97x)) + ((!n_n524) & (!n_n482) & (n_n528) & (x18x) & (x97x)) + ((!n_n524) & (n_n482) & (!n_n528) & (!x18x) & (x97x)) + ((!n_n524) & (n_n482) & (!n_n528) & (x18x) & (x97x)) + ((!n_n524) & (n_n482) & (n_n528) & (!x18x) & (x97x)) + ((!n_n524) & (n_n482) & (n_n528) & (x18x) & (!x97x)) + ((!n_n524) & (n_n482) & (n_n528) & (x18x) & (x97x)) + ((n_n524) & (!n_n482) & (!n_n528) & (!x18x) & (x97x)) + ((n_n524) & (!n_n482) & (!n_n528) & (x18x) & (x97x)) + ((n_n524) & (!n_n482) & (n_n528) & (!x18x) & (x97x)) + ((n_n524) & (!n_n482) & (n_n528) & (x18x) & (x97x)) + ((n_n524) & (n_n482) & (!n_n528) & (!x18x) & (x97x)) + ((n_n524) & (n_n482) & (!n_n528) & (x18x) & (!x97x)) + ((n_n524) & (n_n482) & (!n_n528) & (x18x) & (x97x)) + ((n_n524) & (n_n482) & (n_n528) & (!x18x) & (x97x)) + ((n_n524) & (n_n482) & (n_n528) & (x18x) & (!x97x)) + ((n_n524) & (n_n482) & (n_n528) & (x18x) & (x97x)));
	assign x15979x = (((!n_n5048) & (!n_n5044) & (!n_n5045) & (!n_n5053) & (n_n5047)) + ((!n_n5048) & (!n_n5044) & (!n_n5045) & (n_n5053) & (!n_n5047)) + ((!n_n5048) & (!n_n5044) & (!n_n5045) & (n_n5053) & (n_n5047)) + ((!n_n5048) & (!n_n5044) & (n_n5045) & (!n_n5053) & (!n_n5047)) + ((!n_n5048) & (!n_n5044) & (n_n5045) & (!n_n5053) & (n_n5047)) + ((!n_n5048) & (!n_n5044) & (n_n5045) & (n_n5053) & (!n_n5047)) + ((!n_n5048) & (!n_n5044) & (n_n5045) & (n_n5053) & (n_n5047)) + ((!n_n5048) & (n_n5044) & (!n_n5045) & (!n_n5053) & (!n_n5047)) + ((!n_n5048) & (n_n5044) & (!n_n5045) & (!n_n5053) & (n_n5047)) + ((!n_n5048) & (n_n5044) & (!n_n5045) & (n_n5053) & (!n_n5047)) + ((!n_n5048) & (n_n5044) & (!n_n5045) & (n_n5053) & (n_n5047)) + ((!n_n5048) & (n_n5044) & (n_n5045) & (!n_n5053) & (!n_n5047)) + ((!n_n5048) & (n_n5044) & (n_n5045) & (!n_n5053) & (n_n5047)) + ((!n_n5048) & (n_n5044) & (n_n5045) & (n_n5053) & (!n_n5047)) + ((!n_n5048) & (n_n5044) & (n_n5045) & (n_n5053) & (n_n5047)) + ((n_n5048) & (!n_n5044) & (!n_n5045) & (!n_n5053) & (!n_n5047)) + ((n_n5048) & (!n_n5044) & (!n_n5045) & (!n_n5053) & (n_n5047)) + ((n_n5048) & (!n_n5044) & (!n_n5045) & (n_n5053) & (!n_n5047)) + ((n_n5048) & (!n_n5044) & (!n_n5045) & (n_n5053) & (n_n5047)) + ((n_n5048) & (!n_n5044) & (n_n5045) & (!n_n5053) & (!n_n5047)) + ((n_n5048) & (!n_n5044) & (n_n5045) & (!n_n5053) & (n_n5047)) + ((n_n5048) & (!n_n5044) & (n_n5045) & (n_n5053) & (!n_n5047)) + ((n_n5048) & (!n_n5044) & (n_n5045) & (n_n5053) & (n_n5047)) + ((n_n5048) & (n_n5044) & (!n_n5045) & (!n_n5053) & (!n_n5047)) + ((n_n5048) & (n_n5044) & (!n_n5045) & (!n_n5053) & (n_n5047)) + ((n_n5048) & (n_n5044) & (!n_n5045) & (n_n5053) & (!n_n5047)) + ((n_n5048) & (n_n5044) & (!n_n5045) & (n_n5053) & (n_n5047)) + ((n_n5048) & (n_n5044) & (n_n5045) & (!n_n5053) & (!n_n5047)) + ((n_n5048) & (n_n5044) & (n_n5045) & (!n_n5053) & (n_n5047)) + ((n_n5048) & (n_n5044) & (n_n5045) & (n_n5053) & (!n_n5047)) + ((n_n5048) & (n_n5044) & (n_n5045) & (n_n5053) & (n_n5047)));
	assign n_n1844 = (((!n_n5025) & (!n_n5023) & (!n_n5021) & (!n_n5024) & (x15983x)) + ((!n_n5025) & (!n_n5023) & (!n_n5021) & (n_n5024) & (!x15983x)) + ((!n_n5025) & (!n_n5023) & (!n_n5021) & (n_n5024) & (x15983x)) + ((!n_n5025) & (!n_n5023) & (n_n5021) & (!n_n5024) & (!x15983x)) + ((!n_n5025) & (!n_n5023) & (n_n5021) & (!n_n5024) & (x15983x)) + ((!n_n5025) & (!n_n5023) & (n_n5021) & (n_n5024) & (!x15983x)) + ((!n_n5025) & (!n_n5023) & (n_n5021) & (n_n5024) & (x15983x)) + ((!n_n5025) & (n_n5023) & (!n_n5021) & (!n_n5024) & (!x15983x)) + ((!n_n5025) & (n_n5023) & (!n_n5021) & (!n_n5024) & (x15983x)) + ((!n_n5025) & (n_n5023) & (!n_n5021) & (n_n5024) & (!x15983x)) + ((!n_n5025) & (n_n5023) & (!n_n5021) & (n_n5024) & (x15983x)) + ((!n_n5025) & (n_n5023) & (n_n5021) & (!n_n5024) & (!x15983x)) + ((!n_n5025) & (n_n5023) & (n_n5021) & (!n_n5024) & (x15983x)) + ((!n_n5025) & (n_n5023) & (n_n5021) & (n_n5024) & (!x15983x)) + ((!n_n5025) & (n_n5023) & (n_n5021) & (n_n5024) & (x15983x)) + ((n_n5025) & (!n_n5023) & (!n_n5021) & (!n_n5024) & (!x15983x)) + ((n_n5025) & (!n_n5023) & (!n_n5021) & (!n_n5024) & (x15983x)) + ((n_n5025) & (!n_n5023) & (!n_n5021) & (n_n5024) & (!x15983x)) + ((n_n5025) & (!n_n5023) & (!n_n5021) & (n_n5024) & (x15983x)) + ((n_n5025) & (!n_n5023) & (n_n5021) & (!n_n5024) & (!x15983x)) + ((n_n5025) & (!n_n5023) & (n_n5021) & (!n_n5024) & (x15983x)) + ((n_n5025) & (!n_n5023) & (n_n5021) & (n_n5024) & (!x15983x)) + ((n_n5025) & (!n_n5023) & (n_n5021) & (n_n5024) & (x15983x)) + ((n_n5025) & (n_n5023) & (!n_n5021) & (!n_n5024) & (!x15983x)) + ((n_n5025) & (n_n5023) & (!n_n5021) & (!n_n5024) & (x15983x)) + ((n_n5025) & (n_n5023) & (!n_n5021) & (n_n5024) & (!x15983x)) + ((n_n5025) & (n_n5023) & (!n_n5021) & (n_n5024) & (x15983x)) + ((n_n5025) & (n_n5023) & (n_n5021) & (!n_n5024) & (!x15983x)) + ((n_n5025) & (n_n5023) & (n_n5021) & (!n_n5024) & (x15983x)) + ((n_n5025) & (n_n5023) & (n_n5021) & (n_n5024) & (!x15983x)) + ((n_n5025) & (n_n5023) & (n_n5021) & (n_n5024) & (x15983x)));
	assign x15989x = (((!n_n5027) & (!n_n5028) & (!x50x) & (!n_n5029) & (!x22069x)) + ((!n_n5027) & (!n_n5028) & (!x50x) & (n_n5029) & (!x22069x)) + ((!n_n5027) & (!n_n5028) & (!x50x) & (n_n5029) & (x22069x)) + ((!n_n5027) & (!n_n5028) & (x50x) & (!n_n5029) & (!x22069x)) + ((!n_n5027) & (!n_n5028) & (x50x) & (!n_n5029) & (x22069x)) + ((!n_n5027) & (!n_n5028) & (x50x) & (n_n5029) & (!x22069x)) + ((!n_n5027) & (!n_n5028) & (x50x) & (n_n5029) & (x22069x)) + ((!n_n5027) & (n_n5028) & (!x50x) & (!n_n5029) & (!x22069x)) + ((!n_n5027) & (n_n5028) & (!x50x) & (!n_n5029) & (x22069x)) + ((!n_n5027) & (n_n5028) & (!x50x) & (n_n5029) & (!x22069x)) + ((!n_n5027) & (n_n5028) & (!x50x) & (n_n5029) & (x22069x)) + ((!n_n5027) & (n_n5028) & (x50x) & (!n_n5029) & (!x22069x)) + ((!n_n5027) & (n_n5028) & (x50x) & (!n_n5029) & (x22069x)) + ((!n_n5027) & (n_n5028) & (x50x) & (n_n5029) & (!x22069x)) + ((!n_n5027) & (n_n5028) & (x50x) & (n_n5029) & (x22069x)) + ((n_n5027) & (!n_n5028) & (!x50x) & (!n_n5029) & (!x22069x)) + ((n_n5027) & (!n_n5028) & (!x50x) & (!n_n5029) & (x22069x)) + ((n_n5027) & (!n_n5028) & (!x50x) & (n_n5029) & (!x22069x)) + ((n_n5027) & (!n_n5028) & (!x50x) & (n_n5029) & (x22069x)) + ((n_n5027) & (!n_n5028) & (x50x) & (!n_n5029) & (!x22069x)) + ((n_n5027) & (!n_n5028) & (x50x) & (!n_n5029) & (x22069x)) + ((n_n5027) & (!n_n5028) & (x50x) & (n_n5029) & (!x22069x)) + ((n_n5027) & (!n_n5028) & (x50x) & (n_n5029) & (x22069x)) + ((n_n5027) & (n_n5028) & (!x50x) & (!n_n5029) & (!x22069x)) + ((n_n5027) & (n_n5028) & (!x50x) & (!n_n5029) & (x22069x)) + ((n_n5027) & (n_n5028) & (!x50x) & (n_n5029) & (!x22069x)) + ((n_n5027) & (n_n5028) & (!x50x) & (n_n5029) & (x22069x)) + ((n_n5027) & (n_n5028) & (x50x) & (!n_n5029) & (!x22069x)) + ((n_n5027) & (n_n5028) & (x50x) & (!n_n5029) & (x22069x)) + ((n_n5027) & (n_n5028) & (x50x) & (n_n5029) & (!x22069x)) + ((n_n5027) & (n_n5028) & (x50x) & (n_n5029) & (x22069x)));
	assign x15991x = (((!x15978x) & (!x15979x) & (!n_n1844) & (x15989x)) + ((!x15978x) & (!x15979x) & (n_n1844) & (!x15989x)) + ((!x15978x) & (!x15979x) & (n_n1844) & (x15989x)) + ((!x15978x) & (x15979x) & (!n_n1844) & (!x15989x)) + ((!x15978x) & (x15979x) & (!n_n1844) & (x15989x)) + ((!x15978x) & (x15979x) & (n_n1844) & (!x15989x)) + ((!x15978x) & (x15979x) & (n_n1844) & (x15989x)) + ((x15978x) & (!x15979x) & (!n_n1844) & (!x15989x)) + ((x15978x) & (!x15979x) & (!n_n1844) & (x15989x)) + ((x15978x) & (!x15979x) & (n_n1844) & (!x15989x)) + ((x15978x) & (!x15979x) & (n_n1844) & (x15989x)) + ((x15978x) & (x15979x) & (!n_n1844) & (!x15989x)) + ((x15978x) & (x15979x) & (!n_n1844) & (x15989x)) + ((x15978x) & (x15979x) & (n_n1844) & (!x15989x)) + ((x15978x) & (x15979x) & (n_n1844) & (x15989x)));
	assign n_n1885 = (((!n_n3883) & (!x65x) & (!n_n4492) & (!n_n4496) & (x347x)) + ((!n_n3883) & (!x65x) & (!n_n4492) & (n_n4496) & (!x347x)) + ((!n_n3883) & (!x65x) & (!n_n4492) & (n_n4496) & (x347x)) + ((!n_n3883) & (!x65x) & (n_n4492) & (!n_n4496) & (!x347x)) + ((!n_n3883) & (!x65x) & (n_n4492) & (!n_n4496) & (x347x)) + ((!n_n3883) & (!x65x) & (n_n4492) & (n_n4496) & (!x347x)) + ((!n_n3883) & (!x65x) & (n_n4492) & (n_n4496) & (x347x)) + ((!n_n3883) & (x65x) & (!n_n4492) & (!n_n4496) & (!x347x)) + ((!n_n3883) & (x65x) & (!n_n4492) & (!n_n4496) & (x347x)) + ((!n_n3883) & (x65x) & (!n_n4492) & (n_n4496) & (!x347x)) + ((!n_n3883) & (x65x) & (!n_n4492) & (n_n4496) & (x347x)) + ((!n_n3883) & (x65x) & (n_n4492) & (!n_n4496) & (!x347x)) + ((!n_n3883) & (x65x) & (n_n4492) & (!n_n4496) & (x347x)) + ((!n_n3883) & (x65x) & (n_n4492) & (n_n4496) & (!x347x)) + ((!n_n3883) & (x65x) & (n_n4492) & (n_n4496) & (x347x)) + ((n_n3883) & (!x65x) & (!n_n4492) & (!n_n4496) & (!x347x)) + ((n_n3883) & (!x65x) & (!n_n4492) & (!n_n4496) & (x347x)) + ((n_n3883) & (!x65x) & (!n_n4492) & (n_n4496) & (!x347x)) + ((n_n3883) & (!x65x) & (!n_n4492) & (n_n4496) & (x347x)) + ((n_n3883) & (!x65x) & (n_n4492) & (!n_n4496) & (!x347x)) + ((n_n3883) & (!x65x) & (n_n4492) & (!n_n4496) & (x347x)) + ((n_n3883) & (!x65x) & (n_n4492) & (n_n4496) & (!x347x)) + ((n_n3883) & (!x65x) & (n_n4492) & (n_n4496) & (x347x)) + ((n_n3883) & (x65x) & (!n_n4492) & (!n_n4496) & (!x347x)) + ((n_n3883) & (x65x) & (!n_n4492) & (!n_n4496) & (x347x)) + ((n_n3883) & (x65x) & (!n_n4492) & (n_n4496) & (!x347x)) + ((n_n3883) & (x65x) & (!n_n4492) & (n_n4496) & (x347x)) + ((n_n3883) & (x65x) & (n_n4492) & (!n_n4496) & (!x347x)) + ((n_n3883) & (x65x) & (n_n4492) & (!n_n4496) & (x347x)) + ((n_n3883) & (x65x) & (n_n4492) & (n_n4496) & (!x347x)) + ((n_n3883) & (x65x) & (n_n4492) & (n_n4496) & (x347x)));
	assign n_n1886 = (((!x78x) & (!n_n4477) & (!x184x) & (!n_n4479) & (x376x)) + ((!x78x) & (!n_n4477) & (!x184x) & (n_n4479) & (!x376x)) + ((!x78x) & (!n_n4477) & (!x184x) & (n_n4479) & (x376x)) + ((!x78x) & (!n_n4477) & (x184x) & (!n_n4479) & (!x376x)) + ((!x78x) & (!n_n4477) & (x184x) & (!n_n4479) & (x376x)) + ((!x78x) & (!n_n4477) & (x184x) & (n_n4479) & (!x376x)) + ((!x78x) & (!n_n4477) & (x184x) & (n_n4479) & (x376x)) + ((!x78x) & (n_n4477) & (!x184x) & (!n_n4479) & (!x376x)) + ((!x78x) & (n_n4477) & (!x184x) & (!n_n4479) & (x376x)) + ((!x78x) & (n_n4477) & (!x184x) & (n_n4479) & (!x376x)) + ((!x78x) & (n_n4477) & (!x184x) & (n_n4479) & (x376x)) + ((!x78x) & (n_n4477) & (x184x) & (!n_n4479) & (!x376x)) + ((!x78x) & (n_n4477) & (x184x) & (!n_n4479) & (x376x)) + ((!x78x) & (n_n4477) & (x184x) & (n_n4479) & (!x376x)) + ((!x78x) & (n_n4477) & (x184x) & (n_n4479) & (x376x)) + ((x78x) & (!n_n4477) & (!x184x) & (!n_n4479) & (!x376x)) + ((x78x) & (!n_n4477) & (!x184x) & (!n_n4479) & (x376x)) + ((x78x) & (!n_n4477) & (!x184x) & (n_n4479) & (!x376x)) + ((x78x) & (!n_n4477) & (!x184x) & (n_n4479) & (x376x)) + ((x78x) & (!n_n4477) & (x184x) & (!n_n4479) & (!x376x)) + ((x78x) & (!n_n4477) & (x184x) & (!n_n4479) & (x376x)) + ((x78x) & (!n_n4477) & (x184x) & (n_n4479) & (!x376x)) + ((x78x) & (!n_n4477) & (x184x) & (n_n4479) & (x376x)) + ((x78x) & (n_n4477) & (!x184x) & (!n_n4479) & (!x376x)) + ((x78x) & (n_n4477) & (!x184x) & (!n_n4479) & (x376x)) + ((x78x) & (n_n4477) & (!x184x) & (n_n4479) & (!x376x)) + ((x78x) & (n_n4477) & (!x184x) & (n_n4479) & (x376x)) + ((x78x) & (n_n4477) & (x184x) & (!n_n4479) & (!x376x)) + ((x78x) & (n_n4477) & (x184x) & (!n_n4479) & (x376x)) + ((x78x) & (n_n4477) & (x184x) & (n_n4479) & (!x376x)) + ((x78x) & (n_n4477) & (x184x) & (n_n4479) & (x376x)));
	assign x16023x = (((!n_n4512) & (!n_n4514) & (!n_n4504) & (n_n4503)) + ((!n_n4512) & (!n_n4514) & (n_n4504) & (!n_n4503)) + ((!n_n4512) & (!n_n4514) & (n_n4504) & (n_n4503)) + ((!n_n4512) & (n_n4514) & (!n_n4504) & (!n_n4503)) + ((!n_n4512) & (n_n4514) & (!n_n4504) & (n_n4503)) + ((!n_n4512) & (n_n4514) & (n_n4504) & (!n_n4503)) + ((!n_n4512) & (n_n4514) & (n_n4504) & (n_n4503)) + ((n_n4512) & (!n_n4514) & (!n_n4504) & (!n_n4503)) + ((n_n4512) & (!n_n4514) & (!n_n4504) & (n_n4503)) + ((n_n4512) & (!n_n4514) & (n_n4504) & (!n_n4503)) + ((n_n4512) & (!n_n4514) & (n_n4504) & (n_n4503)) + ((n_n4512) & (n_n4514) & (!n_n4504) & (!n_n4503)) + ((n_n4512) & (n_n4514) & (!n_n4504) & (n_n4503)) + ((n_n4512) & (n_n4514) & (n_n4504) & (!n_n4503)) + ((n_n4512) & (n_n4514) & (n_n4504) & (n_n4503)));
	assign x16024x = (((!x492x) & (!x13x) & (!x572x) & (!n_n4500) & (x189x)) + ((!x492x) & (!x13x) & (!x572x) & (n_n4500) & (!x189x)) + ((!x492x) & (!x13x) & (!x572x) & (n_n4500) & (x189x)) + ((!x492x) & (!x13x) & (x572x) & (!n_n4500) & (x189x)) + ((!x492x) & (!x13x) & (x572x) & (n_n4500) & (!x189x)) + ((!x492x) & (!x13x) & (x572x) & (n_n4500) & (x189x)) + ((!x492x) & (x13x) & (!x572x) & (!n_n4500) & (x189x)) + ((!x492x) & (x13x) & (!x572x) & (n_n4500) & (!x189x)) + ((!x492x) & (x13x) & (!x572x) & (n_n4500) & (x189x)) + ((!x492x) & (x13x) & (x572x) & (!n_n4500) & (!x189x)) + ((!x492x) & (x13x) & (x572x) & (!n_n4500) & (x189x)) + ((!x492x) & (x13x) & (x572x) & (n_n4500) & (!x189x)) + ((!x492x) & (x13x) & (x572x) & (n_n4500) & (x189x)) + ((x492x) & (!x13x) & (!x572x) & (!n_n4500) & (x189x)) + ((x492x) & (!x13x) & (!x572x) & (n_n4500) & (!x189x)) + ((x492x) & (!x13x) & (!x572x) & (n_n4500) & (x189x)) + ((x492x) & (!x13x) & (x572x) & (!n_n4500) & (x189x)) + ((x492x) & (!x13x) & (x572x) & (n_n4500) & (!x189x)) + ((x492x) & (!x13x) & (x572x) & (n_n4500) & (x189x)) + ((x492x) & (x13x) & (!x572x) & (!n_n4500) & (!x189x)) + ((x492x) & (x13x) & (!x572x) & (!n_n4500) & (x189x)) + ((x492x) & (x13x) & (!x572x) & (n_n4500) & (!x189x)) + ((x492x) & (x13x) & (!x572x) & (n_n4500) & (x189x)) + ((x492x) & (x13x) & (x572x) & (!n_n4500) & (!x189x)) + ((x492x) & (x13x) & (x572x) & (!n_n4500) & (x189x)) + ((x492x) & (x13x) & (x572x) & (n_n4500) & (!x189x)) + ((x492x) & (x13x) & (x572x) & (n_n4500) & (x189x)));
	assign x16027x = (((!n_n1885) & (!n_n1886) & (!x16023x) & (x16024x)) + ((!n_n1885) & (!n_n1886) & (x16023x) & (!x16024x)) + ((!n_n1885) & (!n_n1886) & (x16023x) & (x16024x)) + ((!n_n1885) & (n_n1886) & (!x16023x) & (!x16024x)) + ((!n_n1885) & (n_n1886) & (!x16023x) & (x16024x)) + ((!n_n1885) & (n_n1886) & (x16023x) & (!x16024x)) + ((!n_n1885) & (n_n1886) & (x16023x) & (x16024x)) + ((n_n1885) & (!n_n1886) & (!x16023x) & (!x16024x)) + ((n_n1885) & (!n_n1886) & (!x16023x) & (x16024x)) + ((n_n1885) & (!n_n1886) & (x16023x) & (!x16024x)) + ((n_n1885) & (!n_n1886) & (x16023x) & (x16024x)) + ((n_n1885) & (n_n1886) & (!x16023x) & (!x16024x)) + ((n_n1885) & (n_n1886) & (!x16023x) & (x16024x)) + ((n_n1885) & (n_n1886) & (x16023x) & (!x16024x)) + ((n_n1885) & (n_n1886) & (x16023x) & (x16024x)));
	assign n_n1882 = (((!n_n4532) & (!n_n4537) & (!x11532x) & (!n_n4529) & (!x22223x)) + ((!n_n4532) & (!n_n4537) & (!x11532x) & (n_n4529) & (!x22223x)) + ((!n_n4532) & (!n_n4537) & (!x11532x) & (n_n4529) & (x22223x)) + ((!n_n4532) & (!n_n4537) & (x11532x) & (!n_n4529) & (!x22223x)) + ((!n_n4532) & (!n_n4537) & (x11532x) & (!n_n4529) & (x22223x)) + ((!n_n4532) & (!n_n4537) & (x11532x) & (n_n4529) & (!x22223x)) + ((!n_n4532) & (!n_n4537) & (x11532x) & (n_n4529) & (x22223x)) + ((!n_n4532) & (n_n4537) & (!x11532x) & (!n_n4529) & (!x22223x)) + ((!n_n4532) & (n_n4537) & (!x11532x) & (!n_n4529) & (x22223x)) + ((!n_n4532) & (n_n4537) & (!x11532x) & (n_n4529) & (!x22223x)) + ((!n_n4532) & (n_n4537) & (!x11532x) & (n_n4529) & (x22223x)) + ((!n_n4532) & (n_n4537) & (x11532x) & (!n_n4529) & (!x22223x)) + ((!n_n4532) & (n_n4537) & (x11532x) & (!n_n4529) & (x22223x)) + ((!n_n4532) & (n_n4537) & (x11532x) & (n_n4529) & (!x22223x)) + ((!n_n4532) & (n_n4537) & (x11532x) & (n_n4529) & (x22223x)) + ((n_n4532) & (!n_n4537) & (!x11532x) & (!n_n4529) & (!x22223x)) + ((n_n4532) & (!n_n4537) & (!x11532x) & (!n_n4529) & (x22223x)) + ((n_n4532) & (!n_n4537) & (!x11532x) & (n_n4529) & (!x22223x)) + ((n_n4532) & (!n_n4537) & (!x11532x) & (n_n4529) & (x22223x)) + ((n_n4532) & (!n_n4537) & (x11532x) & (!n_n4529) & (!x22223x)) + ((n_n4532) & (!n_n4537) & (x11532x) & (!n_n4529) & (x22223x)) + ((n_n4532) & (!n_n4537) & (x11532x) & (n_n4529) & (!x22223x)) + ((n_n4532) & (!n_n4537) & (x11532x) & (n_n4529) & (x22223x)) + ((n_n4532) & (n_n4537) & (!x11532x) & (!n_n4529) & (!x22223x)) + ((n_n4532) & (n_n4537) & (!x11532x) & (!n_n4529) & (x22223x)) + ((n_n4532) & (n_n4537) & (!x11532x) & (n_n4529) & (!x22223x)) + ((n_n4532) & (n_n4537) & (!x11532x) & (n_n4529) & (x22223x)) + ((n_n4532) & (n_n4537) & (x11532x) & (!n_n4529) & (!x22223x)) + ((n_n4532) & (n_n4537) & (x11532x) & (!n_n4529) & (x22223x)) + ((n_n4532) & (n_n4537) & (x11532x) & (n_n4529) & (!x22223x)) + ((n_n4532) & (n_n4537) & (x11532x) & (n_n4529) & (x22223x)));
	assign n_n1817 = (((!n_n3889) & (!n_n4472) & (!x194x) & (!x16007x) & (n_n1889)) + ((!n_n3889) & (!n_n4472) & (!x194x) & (x16007x) & (!n_n1889)) + ((!n_n3889) & (!n_n4472) & (!x194x) & (x16007x) & (n_n1889)) + ((!n_n3889) & (!n_n4472) & (x194x) & (!x16007x) & (!n_n1889)) + ((!n_n3889) & (!n_n4472) & (x194x) & (!x16007x) & (n_n1889)) + ((!n_n3889) & (!n_n4472) & (x194x) & (x16007x) & (!n_n1889)) + ((!n_n3889) & (!n_n4472) & (x194x) & (x16007x) & (n_n1889)) + ((!n_n3889) & (n_n4472) & (!x194x) & (!x16007x) & (!n_n1889)) + ((!n_n3889) & (n_n4472) & (!x194x) & (!x16007x) & (n_n1889)) + ((!n_n3889) & (n_n4472) & (!x194x) & (x16007x) & (!n_n1889)) + ((!n_n3889) & (n_n4472) & (!x194x) & (x16007x) & (n_n1889)) + ((!n_n3889) & (n_n4472) & (x194x) & (!x16007x) & (!n_n1889)) + ((!n_n3889) & (n_n4472) & (x194x) & (!x16007x) & (n_n1889)) + ((!n_n3889) & (n_n4472) & (x194x) & (x16007x) & (!n_n1889)) + ((!n_n3889) & (n_n4472) & (x194x) & (x16007x) & (n_n1889)) + ((n_n3889) & (!n_n4472) & (!x194x) & (!x16007x) & (!n_n1889)) + ((n_n3889) & (!n_n4472) & (!x194x) & (!x16007x) & (n_n1889)) + ((n_n3889) & (!n_n4472) & (!x194x) & (x16007x) & (!n_n1889)) + ((n_n3889) & (!n_n4472) & (!x194x) & (x16007x) & (n_n1889)) + ((n_n3889) & (!n_n4472) & (x194x) & (!x16007x) & (!n_n1889)) + ((n_n3889) & (!n_n4472) & (x194x) & (!x16007x) & (n_n1889)) + ((n_n3889) & (!n_n4472) & (x194x) & (x16007x) & (!n_n1889)) + ((n_n3889) & (!n_n4472) & (x194x) & (x16007x) & (n_n1889)) + ((n_n3889) & (n_n4472) & (!x194x) & (!x16007x) & (!n_n1889)) + ((n_n3889) & (n_n4472) & (!x194x) & (!x16007x) & (n_n1889)) + ((n_n3889) & (n_n4472) & (!x194x) & (x16007x) & (!n_n1889)) + ((n_n3889) & (n_n4472) & (!x194x) & (x16007x) & (n_n1889)) + ((n_n3889) & (n_n4472) & (x194x) & (!x16007x) & (!n_n1889)) + ((n_n3889) & (n_n4472) & (x194x) & (!x16007x) & (n_n1889)) + ((n_n3889) & (n_n4472) & (x194x) & (x16007x) & (!n_n1889)) + ((n_n3889) & (n_n4472) & (x194x) & (x16007x) & (n_n1889)));
	assign x16018x = (((!n_n4521) & (!n_n4526) & (!n_n3504) & (!x14108x) & (x14109x)) + ((!n_n4521) & (!n_n4526) & (!n_n3504) & (x14108x) & (!x14109x)) + ((!n_n4521) & (!n_n4526) & (!n_n3504) & (x14108x) & (x14109x)) + ((!n_n4521) & (!n_n4526) & (n_n3504) & (!x14108x) & (!x14109x)) + ((!n_n4521) & (!n_n4526) & (n_n3504) & (!x14108x) & (x14109x)) + ((!n_n4521) & (!n_n4526) & (n_n3504) & (x14108x) & (!x14109x)) + ((!n_n4521) & (!n_n4526) & (n_n3504) & (x14108x) & (x14109x)) + ((!n_n4521) & (n_n4526) & (!n_n3504) & (!x14108x) & (!x14109x)) + ((!n_n4521) & (n_n4526) & (!n_n3504) & (!x14108x) & (x14109x)) + ((!n_n4521) & (n_n4526) & (!n_n3504) & (x14108x) & (!x14109x)) + ((!n_n4521) & (n_n4526) & (!n_n3504) & (x14108x) & (x14109x)) + ((!n_n4521) & (n_n4526) & (n_n3504) & (!x14108x) & (!x14109x)) + ((!n_n4521) & (n_n4526) & (n_n3504) & (!x14108x) & (x14109x)) + ((!n_n4521) & (n_n4526) & (n_n3504) & (x14108x) & (!x14109x)) + ((!n_n4521) & (n_n4526) & (n_n3504) & (x14108x) & (x14109x)) + ((n_n4521) & (!n_n4526) & (!n_n3504) & (!x14108x) & (!x14109x)) + ((n_n4521) & (!n_n4526) & (!n_n3504) & (!x14108x) & (x14109x)) + ((n_n4521) & (!n_n4526) & (!n_n3504) & (x14108x) & (!x14109x)) + ((n_n4521) & (!n_n4526) & (!n_n3504) & (x14108x) & (x14109x)) + ((n_n4521) & (!n_n4526) & (n_n3504) & (!x14108x) & (!x14109x)) + ((n_n4521) & (!n_n4526) & (n_n3504) & (!x14108x) & (x14109x)) + ((n_n4521) & (!n_n4526) & (n_n3504) & (x14108x) & (!x14109x)) + ((n_n4521) & (!n_n4526) & (n_n3504) & (x14108x) & (x14109x)) + ((n_n4521) & (n_n4526) & (!n_n3504) & (!x14108x) & (!x14109x)) + ((n_n4521) & (n_n4526) & (!n_n3504) & (!x14108x) & (x14109x)) + ((n_n4521) & (n_n4526) & (!n_n3504) & (x14108x) & (!x14109x)) + ((n_n4521) & (n_n4526) & (!n_n3504) & (x14108x) & (x14109x)) + ((n_n4521) & (n_n4526) & (n_n3504) & (!x14108x) & (!x14109x)) + ((n_n4521) & (n_n4526) & (n_n3504) & (!x14108x) & (x14109x)) + ((n_n4521) & (n_n4526) & (n_n3504) & (x14108x) & (!x14109x)) + ((n_n4521) & (n_n4526) & (n_n3504) & (x14108x) & (x14109x)));
	assign x16017x = (((!n_n4524) & (!x170x) & (!n_n4525) & (!n_n4517) & (x307x)) + ((!n_n4524) & (!x170x) & (!n_n4525) & (n_n4517) & (!x307x)) + ((!n_n4524) & (!x170x) & (!n_n4525) & (n_n4517) & (x307x)) + ((!n_n4524) & (!x170x) & (n_n4525) & (!n_n4517) & (!x307x)) + ((!n_n4524) & (!x170x) & (n_n4525) & (!n_n4517) & (x307x)) + ((!n_n4524) & (!x170x) & (n_n4525) & (n_n4517) & (!x307x)) + ((!n_n4524) & (!x170x) & (n_n4525) & (n_n4517) & (x307x)) + ((!n_n4524) & (x170x) & (!n_n4525) & (!n_n4517) & (!x307x)) + ((!n_n4524) & (x170x) & (!n_n4525) & (!n_n4517) & (x307x)) + ((!n_n4524) & (x170x) & (!n_n4525) & (n_n4517) & (!x307x)) + ((!n_n4524) & (x170x) & (!n_n4525) & (n_n4517) & (x307x)) + ((!n_n4524) & (x170x) & (n_n4525) & (!n_n4517) & (!x307x)) + ((!n_n4524) & (x170x) & (n_n4525) & (!n_n4517) & (x307x)) + ((!n_n4524) & (x170x) & (n_n4525) & (n_n4517) & (!x307x)) + ((!n_n4524) & (x170x) & (n_n4525) & (n_n4517) & (x307x)) + ((n_n4524) & (!x170x) & (!n_n4525) & (!n_n4517) & (!x307x)) + ((n_n4524) & (!x170x) & (!n_n4525) & (!n_n4517) & (x307x)) + ((n_n4524) & (!x170x) & (!n_n4525) & (n_n4517) & (!x307x)) + ((n_n4524) & (!x170x) & (!n_n4525) & (n_n4517) & (x307x)) + ((n_n4524) & (!x170x) & (n_n4525) & (!n_n4517) & (!x307x)) + ((n_n4524) & (!x170x) & (n_n4525) & (!n_n4517) & (x307x)) + ((n_n4524) & (!x170x) & (n_n4525) & (n_n4517) & (!x307x)) + ((n_n4524) & (!x170x) & (n_n4525) & (n_n4517) & (x307x)) + ((n_n4524) & (x170x) & (!n_n4525) & (!n_n4517) & (!x307x)) + ((n_n4524) & (x170x) & (!n_n4525) & (!n_n4517) & (x307x)) + ((n_n4524) & (x170x) & (!n_n4525) & (n_n4517) & (!x307x)) + ((n_n4524) & (x170x) & (!n_n4525) & (n_n4517) & (x307x)) + ((n_n4524) & (x170x) & (n_n4525) & (!n_n4517) & (!x307x)) + ((n_n4524) & (x170x) & (n_n4525) & (!n_n4517) & (x307x)) + ((n_n4524) & (x170x) & (n_n4525) & (n_n4517) & (!x307x)) + ((n_n4524) & (x170x) & (n_n4525) & (n_n4517) & (x307x)));
	assign n_n1878 = (((!n_n4584) & (!n_n4580) & (!x276x) & (!n_n2401) & (x237x)) + ((!n_n4584) & (!n_n4580) & (!x276x) & (n_n2401) & (!x237x)) + ((!n_n4584) & (!n_n4580) & (!x276x) & (n_n2401) & (x237x)) + ((!n_n4584) & (!n_n4580) & (x276x) & (!n_n2401) & (!x237x)) + ((!n_n4584) & (!n_n4580) & (x276x) & (!n_n2401) & (x237x)) + ((!n_n4584) & (!n_n4580) & (x276x) & (n_n2401) & (!x237x)) + ((!n_n4584) & (!n_n4580) & (x276x) & (n_n2401) & (x237x)) + ((!n_n4584) & (n_n4580) & (!x276x) & (!n_n2401) & (!x237x)) + ((!n_n4584) & (n_n4580) & (!x276x) & (!n_n2401) & (x237x)) + ((!n_n4584) & (n_n4580) & (!x276x) & (n_n2401) & (!x237x)) + ((!n_n4584) & (n_n4580) & (!x276x) & (n_n2401) & (x237x)) + ((!n_n4584) & (n_n4580) & (x276x) & (!n_n2401) & (!x237x)) + ((!n_n4584) & (n_n4580) & (x276x) & (!n_n2401) & (x237x)) + ((!n_n4584) & (n_n4580) & (x276x) & (n_n2401) & (!x237x)) + ((!n_n4584) & (n_n4580) & (x276x) & (n_n2401) & (x237x)) + ((n_n4584) & (!n_n4580) & (!x276x) & (!n_n2401) & (!x237x)) + ((n_n4584) & (!n_n4580) & (!x276x) & (!n_n2401) & (x237x)) + ((n_n4584) & (!n_n4580) & (!x276x) & (n_n2401) & (!x237x)) + ((n_n4584) & (!n_n4580) & (!x276x) & (n_n2401) & (x237x)) + ((n_n4584) & (!n_n4580) & (x276x) & (!n_n2401) & (!x237x)) + ((n_n4584) & (!n_n4580) & (x276x) & (!n_n2401) & (x237x)) + ((n_n4584) & (!n_n4580) & (x276x) & (n_n2401) & (!x237x)) + ((n_n4584) & (!n_n4580) & (x276x) & (n_n2401) & (x237x)) + ((n_n4584) & (n_n4580) & (!x276x) & (!n_n2401) & (!x237x)) + ((n_n4584) & (n_n4580) & (!x276x) & (!n_n2401) & (x237x)) + ((n_n4584) & (n_n4580) & (!x276x) & (n_n2401) & (!x237x)) + ((n_n4584) & (n_n4580) & (!x276x) & (n_n2401) & (x237x)) + ((n_n4584) & (n_n4580) & (x276x) & (!n_n2401) & (!x237x)) + ((n_n4584) & (n_n4580) & (x276x) & (!n_n2401) & (x237x)) + ((n_n4584) & (n_n4580) & (x276x) & (n_n2401) & (!x237x)) + ((n_n4584) & (n_n4580) & (x276x) & (n_n2401) & (x237x)));
	assign x16036x = (((!x23x) & (!x523x) & (!n_n4574) & (!n_n4573) & (x121x)) + ((!x23x) & (!x523x) & (!n_n4574) & (n_n4573) & (!x121x)) + ((!x23x) & (!x523x) & (!n_n4574) & (n_n4573) & (x121x)) + ((!x23x) & (!x523x) & (n_n4574) & (!n_n4573) & (!x121x)) + ((!x23x) & (!x523x) & (n_n4574) & (!n_n4573) & (x121x)) + ((!x23x) & (!x523x) & (n_n4574) & (n_n4573) & (!x121x)) + ((!x23x) & (!x523x) & (n_n4574) & (n_n4573) & (x121x)) + ((!x23x) & (x523x) & (!n_n4574) & (!n_n4573) & (x121x)) + ((!x23x) & (x523x) & (!n_n4574) & (n_n4573) & (!x121x)) + ((!x23x) & (x523x) & (!n_n4574) & (n_n4573) & (x121x)) + ((!x23x) & (x523x) & (n_n4574) & (!n_n4573) & (!x121x)) + ((!x23x) & (x523x) & (n_n4574) & (!n_n4573) & (x121x)) + ((!x23x) & (x523x) & (n_n4574) & (n_n4573) & (!x121x)) + ((!x23x) & (x523x) & (n_n4574) & (n_n4573) & (x121x)) + ((x23x) & (!x523x) & (!n_n4574) & (!n_n4573) & (x121x)) + ((x23x) & (!x523x) & (!n_n4574) & (n_n4573) & (!x121x)) + ((x23x) & (!x523x) & (!n_n4574) & (n_n4573) & (x121x)) + ((x23x) & (!x523x) & (n_n4574) & (!n_n4573) & (!x121x)) + ((x23x) & (!x523x) & (n_n4574) & (!n_n4573) & (x121x)) + ((x23x) & (!x523x) & (n_n4574) & (n_n4573) & (!x121x)) + ((x23x) & (!x523x) & (n_n4574) & (n_n4573) & (x121x)) + ((x23x) & (x523x) & (!n_n4574) & (!n_n4573) & (!x121x)) + ((x23x) & (x523x) & (!n_n4574) & (!n_n4573) & (x121x)) + ((x23x) & (x523x) & (!n_n4574) & (n_n4573) & (!x121x)) + ((x23x) & (x523x) & (!n_n4574) & (n_n4573) & (x121x)) + ((x23x) & (x523x) & (n_n4574) & (!n_n4573) & (!x121x)) + ((x23x) & (x523x) & (n_n4574) & (!n_n4573) & (x121x)) + ((x23x) & (x523x) & (n_n4574) & (n_n4573) & (!x121x)) + ((x23x) & (x523x) & (n_n4574) & (n_n4573) & (x121x)));
	assign x16070x = (((!n_n4560) & (!n_n4551) & (!x214x) & (!x430x) & (n_n4239)) + ((!n_n4560) & (!n_n4551) & (!x214x) & (x430x) & (!n_n4239)) + ((!n_n4560) & (!n_n4551) & (!x214x) & (x430x) & (n_n4239)) + ((!n_n4560) & (!n_n4551) & (x214x) & (!x430x) & (!n_n4239)) + ((!n_n4560) & (!n_n4551) & (x214x) & (!x430x) & (n_n4239)) + ((!n_n4560) & (!n_n4551) & (x214x) & (x430x) & (!n_n4239)) + ((!n_n4560) & (!n_n4551) & (x214x) & (x430x) & (n_n4239)) + ((!n_n4560) & (n_n4551) & (!x214x) & (!x430x) & (!n_n4239)) + ((!n_n4560) & (n_n4551) & (!x214x) & (!x430x) & (n_n4239)) + ((!n_n4560) & (n_n4551) & (!x214x) & (x430x) & (!n_n4239)) + ((!n_n4560) & (n_n4551) & (!x214x) & (x430x) & (n_n4239)) + ((!n_n4560) & (n_n4551) & (x214x) & (!x430x) & (!n_n4239)) + ((!n_n4560) & (n_n4551) & (x214x) & (!x430x) & (n_n4239)) + ((!n_n4560) & (n_n4551) & (x214x) & (x430x) & (!n_n4239)) + ((!n_n4560) & (n_n4551) & (x214x) & (x430x) & (n_n4239)) + ((n_n4560) & (!n_n4551) & (!x214x) & (!x430x) & (!n_n4239)) + ((n_n4560) & (!n_n4551) & (!x214x) & (!x430x) & (n_n4239)) + ((n_n4560) & (!n_n4551) & (!x214x) & (x430x) & (!n_n4239)) + ((n_n4560) & (!n_n4551) & (!x214x) & (x430x) & (n_n4239)) + ((n_n4560) & (!n_n4551) & (x214x) & (!x430x) & (!n_n4239)) + ((n_n4560) & (!n_n4551) & (x214x) & (!x430x) & (n_n4239)) + ((n_n4560) & (!n_n4551) & (x214x) & (x430x) & (!n_n4239)) + ((n_n4560) & (!n_n4551) & (x214x) & (x430x) & (n_n4239)) + ((n_n4560) & (n_n4551) & (!x214x) & (!x430x) & (!n_n4239)) + ((n_n4560) & (n_n4551) & (!x214x) & (!x430x) & (n_n4239)) + ((n_n4560) & (n_n4551) & (!x214x) & (x430x) & (!n_n4239)) + ((n_n4560) & (n_n4551) & (!x214x) & (x430x) & (n_n4239)) + ((n_n4560) & (n_n4551) & (x214x) & (!x430x) & (!n_n4239)) + ((n_n4560) & (n_n4551) & (x214x) & (!x430x) & (n_n4239)) + ((n_n4560) & (n_n4551) & (x214x) & (x430x) & (!n_n4239)) + ((n_n4560) & (n_n4551) & (x214x) & (x430x) & (n_n4239)));
	assign x22201x = (((!n_n4571) & (!n_n4575) & (!n_n4577) & (!n_n4576)));
	assign x16072x = (((!n_n1878) & (!x16036x) & (!x16070x) & (!x22201x)) + ((!n_n1878) & (!x16036x) & (x16070x) & (!x22201x)) + ((!n_n1878) & (!x16036x) & (x16070x) & (x22201x)) + ((!n_n1878) & (x16036x) & (!x16070x) & (!x22201x)) + ((!n_n1878) & (x16036x) & (!x16070x) & (x22201x)) + ((!n_n1878) & (x16036x) & (x16070x) & (!x22201x)) + ((!n_n1878) & (x16036x) & (x16070x) & (x22201x)) + ((n_n1878) & (!x16036x) & (!x16070x) & (!x22201x)) + ((n_n1878) & (!x16036x) & (!x16070x) & (x22201x)) + ((n_n1878) & (!x16036x) & (x16070x) & (!x22201x)) + ((n_n1878) & (!x16036x) & (x16070x) & (x22201x)) + ((n_n1878) & (x16036x) & (!x16070x) & (!x22201x)) + ((n_n1878) & (x16036x) & (!x16070x) & (x22201x)) + ((n_n1878) & (x16036x) & (x16070x) & (!x22201x)) + ((n_n1878) & (x16036x) & (x16070x) & (x22201x)));
	assign n_n1877 = (((!n_n4595) & (!x172x) & (!n_n4588) & (!x45x) & (n_n2037)) + ((!n_n4595) & (!x172x) & (!n_n4588) & (x45x) & (!n_n2037)) + ((!n_n4595) & (!x172x) & (!n_n4588) & (x45x) & (n_n2037)) + ((!n_n4595) & (!x172x) & (n_n4588) & (!x45x) & (!n_n2037)) + ((!n_n4595) & (!x172x) & (n_n4588) & (!x45x) & (n_n2037)) + ((!n_n4595) & (!x172x) & (n_n4588) & (x45x) & (!n_n2037)) + ((!n_n4595) & (!x172x) & (n_n4588) & (x45x) & (n_n2037)) + ((!n_n4595) & (x172x) & (!n_n4588) & (!x45x) & (!n_n2037)) + ((!n_n4595) & (x172x) & (!n_n4588) & (!x45x) & (n_n2037)) + ((!n_n4595) & (x172x) & (!n_n4588) & (x45x) & (!n_n2037)) + ((!n_n4595) & (x172x) & (!n_n4588) & (x45x) & (n_n2037)) + ((!n_n4595) & (x172x) & (n_n4588) & (!x45x) & (!n_n2037)) + ((!n_n4595) & (x172x) & (n_n4588) & (!x45x) & (n_n2037)) + ((!n_n4595) & (x172x) & (n_n4588) & (x45x) & (!n_n2037)) + ((!n_n4595) & (x172x) & (n_n4588) & (x45x) & (n_n2037)) + ((n_n4595) & (!x172x) & (!n_n4588) & (!x45x) & (!n_n2037)) + ((n_n4595) & (!x172x) & (!n_n4588) & (!x45x) & (n_n2037)) + ((n_n4595) & (!x172x) & (!n_n4588) & (x45x) & (!n_n2037)) + ((n_n4595) & (!x172x) & (!n_n4588) & (x45x) & (n_n2037)) + ((n_n4595) & (!x172x) & (n_n4588) & (!x45x) & (!n_n2037)) + ((n_n4595) & (!x172x) & (n_n4588) & (!x45x) & (n_n2037)) + ((n_n4595) & (!x172x) & (n_n4588) & (x45x) & (!n_n2037)) + ((n_n4595) & (!x172x) & (n_n4588) & (x45x) & (n_n2037)) + ((n_n4595) & (x172x) & (!n_n4588) & (!x45x) & (!n_n2037)) + ((n_n4595) & (x172x) & (!n_n4588) & (!x45x) & (n_n2037)) + ((n_n4595) & (x172x) & (!n_n4588) & (x45x) & (!n_n2037)) + ((n_n4595) & (x172x) & (!n_n4588) & (x45x) & (n_n2037)) + ((n_n4595) & (x172x) & (n_n4588) & (!x45x) & (!n_n2037)) + ((n_n4595) & (x172x) & (n_n4588) & (!x45x) & (n_n2037)) + ((n_n4595) & (x172x) & (n_n4588) & (x45x) & (!n_n2037)) + ((n_n4595) & (x172x) & (n_n4588) & (x45x) & (n_n2037)));
	assign x16048x = (((!n_n4617) & (!n_n4628) & (!n_n4621) & (!n_n4630) & (x16047x)) + ((!n_n4617) & (!n_n4628) & (!n_n4621) & (n_n4630) & (!x16047x)) + ((!n_n4617) & (!n_n4628) & (!n_n4621) & (n_n4630) & (x16047x)) + ((!n_n4617) & (!n_n4628) & (n_n4621) & (!n_n4630) & (!x16047x)) + ((!n_n4617) & (!n_n4628) & (n_n4621) & (!n_n4630) & (x16047x)) + ((!n_n4617) & (!n_n4628) & (n_n4621) & (n_n4630) & (!x16047x)) + ((!n_n4617) & (!n_n4628) & (n_n4621) & (n_n4630) & (x16047x)) + ((!n_n4617) & (n_n4628) & (!n_n4621) & (!n_n4630) & (!x16047x)) + ((!n_n4617) & (n_n4628) & (!n_n4621) & (!n_n4630) & (x16047x)) + ((!n_n4617) & (n_n4628) & (!n_n4621) & (n_n4630) & (!x16047x)) + ((!n_n4617) & (n_n4628) & (!n_n4621) & (n_n4630) & (x16047x)) + ((!n_n4617) & (n_n4628) & (n_n4621) & (!n_n4630) & (!x16047x)) + ((!n_n4617) & (n_n4628) & (n_n4621) & (!n_n4630) & (x16047x)) + ((!n_n4617) & (n_n4628) & (n_n4621) & (n_n4630) & (!x16047x)) + ((!n_n4617) & (n_n4628) & (n_n4621) & (n_n4630) & (x16047x)) + ((n_n4617) & (!n_n4628) & (!n_n4621) & (!n_n4630) & (!x16047x)) + ((n_n4617) & (!n_n4628) & (!n_n4621) & (!n_n4630) & (x16047x)) + ((n_n4617) & (!n_n4628) & (!n_n4621) & (n_n4630) & (!x16047x)) + ((n_n4617) & (!n_n4628) & (!n_n4621) & (n_n4630) & (x16047x)) + ((n_n4617) & (!n_n4628) & (n_n4621) & (!n_n4630) & (!x16047x)) + ((n_n4617) & (!n_n4628) & (n_n4621) & (!n_n4630) & (x16047x)) + ((n_n4617) & (!n_n4628) & (n_n4621) & (n_n4630) & (!x16047x)) + ((n_n4617) & (!n_n4628) & (n_n4621) & (n_n4630) & (x16047x)) + ((n_n4617) & (n_n4628) & (!n_n4621) & (!n_n4630) & (!x16047x)) + ((n_n4617) & (n_n4628) & (!n_n4621) & (!n_n4630) & (x16047x)) + ((n_n4617) & (n_n4628) & (!n_n4621) & (n_n4630) & (!x16047x)) + ((n_n4617) & (n_n4628) & (!n_n4621) & (n_n4630) & (x16047x)) + ((n_n4617) & (n_n4628) & (n_n4621) & (!n_n4630) & (!x16047x)) + ((n_n4617) & (n_n4628) & (n_n4621) & (!n_n4630) & (x16047x)) + ((n_n4617) & (n_n4628) & (n_n4621) & (n_n4630) & (!x16047x)) + ((n_n4617) & (n_n4628) & (n_n4621) & (n_n4630) & (x16047x)));
	assign n_n1812 = (((!x16065x) & (!x16053x) & (!x16054x) & (n_n1873)) + ((!x16065x) & (!x16053x) & (x16054x) & (!n_n1873)) + ((!x16065x) & (!x16053x) & (x16054x) & (n_n1873)) + ((!x16065x) & (x16053x) & (!x16054x) & (!n_n1873)) + ((!x16065x) & (x16053x) & (!x16054x) & (n_n1873)) + ((!x16065x) & (x16053x) & (x16054x) & (!n_n1873)) + ((!x16065x) & (x16053x) & (x16054x) & (n_n1873)) + ((x16065x) & (!x16053x) & (!x16054x) & (!n_n1873)) + ((x16065x) & (!x16053x) & (!x16054x) & (n_n1873)) + ((x16065x) & (!x16053x) & (x16054x) & (!n_n1873)) + ((x16065x) & (!x16053x) & (x16054x) & (n_n1873)) + ((x16065x) & (x16053x) & (!x16054x) & (!n_n1873)) + ((x16065x) & (x16053x) & (!x16054x) & (n_n1873)) + ((x16065x) & (x16053x) & (x16054x) & (!n_n1873)) + ((x16065x) & (x16053x) & (x16054x) & (n_n1873)));
	assign n_n1876 = (((!n_n4612) & (!n_n4609) & (!n_n4608) & (!x51x) & (n_n2036)) + ((!n_n4612) & (!n_n4609) & (!n_n4608) & (x51x) & (!n_n2036)) + ((!n_n4612) & (!n_n4609) & (!n_n4608) & (x51x) & (n_n2036)) + ((!n_n4612) & (!n_n4609) & (n_n4608) & (!x51x) & (!n_n2036)) + ((!n_n4612) & (!n_n4609) & (n_n4608) & (!x51x) & (n_n2036)) + ((!n_n4612) & (!n_n4609) & (n_n4608) & (x51x) & (!n_n2036)) + ((!n_n4612) & (!n_n4609) & (n_n4608) & (x51x) & (n_n2036)) + ((!n_n4612) & (n_n4609) & (!n_n4608) & (!x51x) & (!n_n2036)) + ((!n_n4612) & (n_n4609) & (!n_n4608) & (!x51x) & (n_n2036)) + ((!n_n4612) & (n_n4609) & (!n_n4608) & (x51x) & (!n_n2036)) + ((!n_n4612) & (n_n4609) & (!n_n4608) & (x51x) & (n_n2036)) + ((!n_n4612) & (n_n4609) & (n_n4608) & (!x51x) & (!n_n2036)) + ((!n_n4612) & (n_n4609) & (n_n4608) & (!x51x) & (n_n2036)) + ((!n_n4612) & (n_n4609) & (n_n4608) & (x51x) & (!n_n2036)) + ((!n_n4612) & (n_n4609) & (n_n4608) & (x51x) & (n_n2036)) + ((n_n4612) & (!n_n4609) & (!n_n4608) & (!x51x) & (!n_n2036)) + ((n_n4612) & (!n_n4609) & (!n_n4608) & (!x51x) & (n_n2036)) + ((n_n4612) & (!n_n4609) & (!n_n4608) & (x51x) & (!n_n2036)) + ((n_n4612) & (!n_n4609) & (!n_n4608) & (x51x) & (n_n2036)) + ((n_n4612) & (!n_n4609) & (n_n4608) & (!x51x) & (!n_n2036)) + ((n_n4612) & (!n_n4609) & (n_n4608) & (!x51x) & (n_n2036)) + ((n_n4612) & (!n_n4609) & (n_n4608) & (x51x) & (!n_n2036)) + ((n_n4612) & (!n_n4609) & (n_n4608) & (x51x) & (n_n2036)) + ((n_n4612) & (n_n4609) & (!n_n4608) & (!x51x) & (!n_n2036)) + ((n_n4612) & (n_n4609) & (!n_n4608) & (!x51x) & (n_n2036)) + ((n_n4612) & (n_n4609) & (!n_n4608) & (x51x) & (!n_n2036)) + ((n_n4612) & (n_n4609) & (!n_n4608) & (x51x) & (n_n2036)) + ((n_n4612) & (n_n4609) & (n_n4608) & (!x51x) & (!n_n2036)) + ((n_n4612) & (n_n4609) & (n_n4608) & (!x51x) & (n_n2036)) + ((n_n4612) & (n_n4609) & (n_n4608) & (x51x) & (!n_n2036)) + ((n_n4612) & (n_n4609) & (n_n4608) & (x51x) & (n_n2036)));
	assign n_n1894 = (((!n_n4369) & (!n_n4275) & (!x64x) & (x16089x)) + ((!n_n4369) & (!n_n4275) & (x64x) & (!x16089x)) + ((!n_n4369) & (!n_n4275) & (x64x) & (x16089x)) + ((!n_n4369) & (n_n4275) & (!x64x) & (!x16089x)) + ((!n_n4369) & (n_n4275) & (!x64x) & (x16089x)) + ((!n_n4369) & (n_n4275) & (x64x) & (!x16089x)) + ((!n_n4369) & (n_n4275) & (x64x) & (x16089x)) + ((n_n4369) & (!n_n4275) & (!x64x) & (!x16089x)) + ((n_n4369) & (!n_n4275) & (!x64x) & (x16089x)) + ((n_n4369) & (!n_n4275) & (x64x) & (!x16089x)) + ((n_n4369) & (!n_n4275) & (x64x) & (x16089x)) + ((n_n4369) & (n_n4275) & (!x64x) & (!x16089x)) + ((n_n4369) & (n_n4275) & (!x64x) & (x16089x)) + ((n_n4369) & (n_n4275) & (x64x) & (!x16089x)) + ((n_n4369) & (n_n4275) & (x64x) & (x16089x)));
	assign n_n1893 = (((!n_n4380) & (!x280x) & (!n_n3903) & (!x14460x) & (n_n4377)) + ((!n_n4380) & (!x280x) & (!n_n3903) & (x14460x) & (!n_n4377)) + ((!n_n4380) & (!x280x) & (!n_n3903) & (x14460x) & (n_n4377)) + ((!n_n4380) & (!x280x) & (n_n3903) & (!x14460x) & (!n_n4377)) + ((!n_n4380) & (!x280x) & (n_n3903) & (!x14460x) & (n_n4377)) + ((!n_n4380) & (!x280x) & (n_n3903) & (x14460x) & (!n_n4377)) + ((!n_n4380) & (!x280x) & (n_n3903) & (x14460x) & (n_n4377)) + ((!n_n4380) & (x280x) & (!n_n3903) & (!x14460x) & (!n_n4377)) + ((!n_n4380) & (x280x) & (!n_n3903) & (!x14460x) & (n_n4377)) + ((!n_n4380) & (x280x) & (!n_n3903) & (x14460x) & (!n_n4377)) + ((!n_n4380) & (x280x) & (!n_n3903) & (x14460x) & (n_n4377)) + ((!n_n4380) & (x280x) & (n_n3903) & (!x14460x) & (!n_n4377)) + ((!n_n4380) & (x280x) & (n_n3903) & (!x14460x) & (n_n4377)) + ((!n_n4380) & (x280x) & (n_n3903) & (x14460x) & (!n_n4377)) + ((!n_n4380) & (x280x) & (n_n3903) & (x14460x) & (n_n4377)) + ((n_n4380) & (!x280x) & (!n_n3903) & (!x14460x) & (!n_n4377)) + ((n_n4380) & (!x280x) & (!n_n3903) & (!x14460x) & (n_n4377)) + ((n_n4380) & (!x280x) & (!n_n3903) & (x14460x) & (!n_n4377)) + ((n_n4380) & (!x280x) & (!n_n3903) & (x14460x) & (n_n4377)) + ((n_n4380) & (!x280x) & (n_n3903) & (!x14460x) & (!n_n4377)) + ((n_n4380) & (!x280x) & (n_n3903) & (!x14460x) & (n_n4377)) + ((n_n4380) & (!x280x) & (n_n3903) & (x14460x) & (!n_n4377)) + ((n_n4380) & (!x280x) & (n_n3903) & (x14460x) & (n_n4377)) + ((n_n4380) & (x280x) & (!n_n3903) & (!x14460x) & (!n_n4377)) + ((n_n4380) & (x280x) & (!n_n3903) & (!x14460x) & (n_n4377)) + ((n_n4380) & (x280x) & (!n_n3903) & (x14460x) & (!n_n4377)) + ((n_n4380) & (x280x) & (!n_n3903) & (x14460x) & (n_n4377)) + ((n_n4380) & (x280x) & (n_n3903) & (!x14460x) & (!n_n4377)) + ((n_n4380) & (x280x) & (n_n3903) & (!x14460x) & (n_n4377)) + ((n_n4380) & (x280x) & (n_n3903) & (x14460x) & (!n_n4377)) + ((n_n4380) & (x280x) & (n_n3903) & (x14460x) & (n_n4377)));
	assign x16110x = (((!n_n4361) & (!n_n4363) & (!n_n4359) & (n_n4356)) + ((!n_n4361) & (!n_n4363) & (n_n4359) & (!n_n4356)) + ((!n_n4361) & (!n_n4363) & (n_n4359) & (n_n4356)) + ((!n_n4361) & (n_n4363) & (!n_n4359) & (!n_n4356)) + ((!n_n4361) & (n_n4363) & (!n_n4359) & (n_n4356)) + ((!n_n4361) & (n_n4363) & (n_n4359) & (!n_n4356)) + ((!n_n4361) & (n_n4363) & (n_n4359) & (n_n4356)) + ((n_n4361) & (!n_n4363) & (!n_n4359) & (!n_n4356)) + ((n_n4361) & (!n_n4363) & (!n_n4359) & (n_n4356)) + ((n_n4361) & (!n_n4363) & (n_n4359) & (!n_n4356)) + ((n_n4361) & (!n_n4363) & (n_n4359) & (n_n4356)) + ((n_n4361) & (n_n4363) & (!n_n4359) & (!n_n4356)) + ((n_n4361) & (n_n4363) & (!n_n4359) & (n_n4356)) + ((n_n4361) & (n_n4363) & (n_n4359) & (!n_n4356)) + ((n_n4361) & (n_n4363) & (n_n4359) & (n_n4356)));
	assign x16111x = (((!n_n4357) & (!n_n4358) & (!n_n4354) & (!n_n4350) & (n_n4355)) + ((!n_n4357) & (!n_n4358) & (!n_n4354) & (n_n4350) & (!n_n4355)) + ((!n_n4357) & (!n_n4358) & (!n_n4354) & (n_n4350) & (n_n4355)) + ((!n_n4357) & (!n_n4358) & (n_n4354) & (!n_n4350) & (!n_n4355)) + ((!n_n4357) & (!n_n4358) & (n_n4354) & (!n_n4350) & (n_n4355)) + ((!n_n4357) & (!n_n4358) & (n_n4354) & (n_n4350) & (!n_n4355)) + ((!n_n4357) & (!n_n4358) & (n_n4354) & (n_n4350) & (n_n4355)) + ((!n_n4357) & (n_n4358) & (!n_n4354) & (!n_n4350) & (!n_n4355)) + ((!n_n4357) & (n_n4358) & (!n_n4354) & (!n_n4350) & (n_n4355)) + ((!n_n4357) & (n_n4358) & (!n_n4354) & (n_n4350) & (!n_n4355)) + ((!n_n4357) & (n_n4358) & (!n_n4354) & (n_n4350) & (n_n4355)) + ((!n_n4357) & (n_n4358) & (n_n4354) & (!n_n4350) & (!n_n4355)) + ((!n_n4357) & (n_n4358) & (n_n4354) & (!n_n4350) & (n_n4355)) + ((!n_n4357) & (n_n4358) & (n_n4354) & (n_n4350) & (!n_n4355)) + ((!n_n4357) & (n_n4358) & (n_n4354) & (n_n4350) & (n_n4355)) + ((n_n4357) & (!n_n4358) & (!n_n4354) & (!n_n4350) & (!n_n4355)) + ((n_n4357) & (!n_n4358) & (!n_n4354) & (!n_n4350) & (n_n4355)) + ((n_n4357) & (!n_n4358) & (!n_n4354) & (n_n4350) & (!n_n4355)) + ((n_n4357) & (!n_n4358) & (!n_n4354) & (n_n4350) & (n_n4355)) + ((n_n4357) & (!n_n4358) & (n_n4354) & (!n_n4350) & (!n_n4355)) + ((n_n4357) & (!n_n4358) & (n_n4354) & (!n_n4350) & (n_n4355)) + ((n_n4357) & (!n_n4358) & (n_n4354) & (n_n4350) & (!n_n4355)) + ((n_n4357) & (!n_n4358) & (n_n4354) & (n_n4350) & (n_n4355)) + ((n_n4357) & (n_n4358) & (!n_n4354) & (!n_n4350) & (!n_n4355)) + ((n_n4357) & (n_n4358) & (!n_n4354) & (!n_n4350) & (n_n4355)) + ((n_n4357) & (n_n4358) & (!n_n4354) & (n_n4350) & (!n_n4355)) + ((n_n4357) & (n_n4358) & (!n_n4354) & (n_n4350) & (n_n4355)) + ((n_n4357) & (n_n4358) & (n_n4354) & (!n_n4350) & (!n_n4355)) + ((n_n4357) & (n_n4358) & (n_n4354) & (!n_n4350) & (n_n4355)) + ((n_n4357) & (n_n4358) & (n_n4354) & (n_n4350) & (!n_n4355)) + ((n_n4357) & (n_n4358) & (n_n4354) & (n_n4350) & (n_n4355)));
	assign x16114x = (((!n_n1894) & (!n_n1893) & (!x16110x) & (x16111x)) + ((!n_n1894) & (!n_n1893) & (x16110x) & (!x16111x)) + ((!n_n1894) & (!n_n1893) & (x16110x) & (x16111x)) + ((!n_n1894) & (n_n1893) & (!x16110x) & (!x16111x)) + ((!n_n1894) & (n_n1893) & (!x16110x) & (x16111x)) + ((!n_n1894) & (n_n1893) & (x16110x) & (!x16111x)) + ((!n_n1894) & (n_n1893) & (x16110x) & (x16111x)) + ((n_n1894) & (!n_n1893) & (!x16110x) & (!x16111x)) + ((n_n1894) & (!n_n1893) & (!x16110x) & (x16111x)) + ((n_n1894) & (!n_n1893) & (x16110x) & (!x16111x)) + ((n_n1894) & (!n_n1893) & (x16110x) & (x16111x)) + ((n_n1894) & (n_n1893) & (!x16110x) & (!x16111x)) + ((n_n1894) & (n_n1893) & (!x16110x) & (x16111x)) + ((n_n1894) & (n_n1893) & (x16110x) & (!x16111x)) + ((n_n1894) & (n_n1893) & (x16110x) & (x16111x)));
	assign n_n1896 = (((!n_n4338) & (!n_n4339) & (!n_n4335) & (!x124x) & (!x22078x)) + ((!n_n4338) & (!n_n4339) & (!n_n4335) & (x124x) & (!x22078x)) + ((!n_n4338) & (!n_n4339) & (!n_n4335) & (x124x) & (x22078x)) + ((!n_n4338) & (!n_n4339) & (n_n4335) & (!x124x) & (!x22078x)) + ((!n_n4338) & (!n_n4339) & (n_n4335) & (!x124x) & (x22078x)) + ((!n_n4338) & (!n_n4339) & (n_n4335) & (x124x) & (!x22078x)) + ((!n_n4338) & (!n_n4339) & (n_n4335) & (x124x) & (x22078x)) + ((!n_n4338) & (n_n4339) & (!n_n4335) & (!x124x) & (!x22078x)) + ((!n_n4338) & (n_n4339) & (!n_n4335) & (!x124x) & (x22078x)) + ((!n_n4338) & (n_n4339) & (!n_n4335) & (x124x) & (!x22078x)) + ((!n_n4338) & (n_n4339) & (!n_n4335) & (x124x) & (x22078x)) + ((!n_n4338) & (n_n4339) & (n_n4335) & (!x124x) & (!x22078x)) + ((!n_n4338) & (n_n4339) & (n_n4335) & (!x124x) & (x22078x)) + ((!n_n4338) & (n_n4339) & (n_n4335) & (x124x) & (!x22078x)) + ((!n_n4338) & (n_n4339) & (n_n4335) & (x124x) & (x22078x)) + ((n_n4338) & (!n_n4339) & (!n_n4335) & (!x124x) & (!x22078x)) + ((n_n4338) & (!n_n4339) & (!n_n4335) & (!x124x) & (x22078x)) + ((n_n4338) & (!n_n4339) & (!n_n4335) & (x124x) & (!x22078x)) + ((n_n4338) & (!n_n4339) & (!n_n4335) & (x124x) & (x22078x)) + ((n_n4338) & (!n_n4339) & (n_n4335) & (!x124x) & (!x22078x)) + ((n_n4338) & (!n_n4339) & (n_n4335) & (!x124x) & (x22078x)) + ((n_n4338) & (!n_n4339) & (n_n4335) & (x124x) & (!x22078x)) + ((n_n4338) & (!n_n4339) & (n_n4335) & (x124x) & (x22078x)) + ((n_n4338) & (n_n4339) & (!n_n4335) & (!x124x) & (!x22078x)) + ((n_n4338) & (n_n4339) & (!n_n4335) & (!x124x) & (x22078x)) + ((n_n4338) & (n_n4339) & (!n_n4335) & (x124x) & (!x22078x)) + ((n_n4338) & (n_n4339) & (!n_n4335) & (x124x) & (x22078x)) + ((n_n4338) & (n_n4339) & (n_n4335) & (!x124x) & (!x22078x)) + ((n_n4338) & (n_n4339) & (n_n4335) & (!x124x) & (x22078x)) + ((n_n4338) & (n_n4339) & (n_n4335) & (x124x) & (!x22078x)) + ((n_n4338) & (n_n4339) & (n_n4335) & (x124x) & (x22078x)));
	assign x16086x = (((!n_n4318) & (!n_n4331) & (!n_n4279) & (!n_n1703) & (x16080x)) + ((!n_n4318) & (!n_n4331) & (!n_n4279) & (n_n1703) & (!x16080x)) + ((!n_n4318) & (!n_n4331) & (!n_n4279) & (n_n1703) & (x16080x)) + ((!n_n4318) & (!n_n4331) & (n_n4279) & (!n_n1703) & (!x16080x)) + ((!n_n4318) & (!n_n4331) & (n_n4279) & (!n_n1703) & (x16080x)) + ((!n_n4318) & (!n_n4331) & (n_n4279) & (n_n1703) & (!x16080x)) + ((!n_n4318) & (!n_n4331) & (n_n4279) & (n_n1703) & (x16080x)) + ((!n_n4318) & (n_n4331) & (!n_n4279) & (!n_n1703) & (!x16080x)) + ((!n_n4318) & (n_n4331) & (!n_n4279) & (!n_n1703) & (x16080x)) + ((!n_n4318) & (n_n4331) & (!n_n4279) & (n_n1703) & (!x16080x)) + ((!n_n4318) & (n_n4331) & (!n_n4279) & (n_n1703) & (x16080x)) + ((!n_n4318) & (n_n4331) & (n_n4279) & (!n_n1703) & (!x16080x)) + ((!n_n4318) & (n_n4331) & (n_n4279) & (!n_n1703) & (x16080x)) + ((!n_n4318) & (n_n4331) & (n_n4279) & (n_n1703) & (!x16080x)) + ((!n_n4318) & (n_n4331) & (n_n4279) & (n_n1703) & (x16080x)) + ((n_n4318) & (!n_n4331) & (!n_n4279) & (!n_n1703) & (!x16080x)) + ((n_n4318) & (!n_n4331) & (!n_n4279) & (!n_n1703) & (x16080x)) + ((n_n4318) & (!n_n4331) & (!n_n4279) & (n_n1703) & (!x16080x)) + ((n_n4318) & (!n_n4331) & (!n_n4279) & (n_n1703) & (x16080x)) + ((n_n4318) & (!n_n4331) & (n_n4279) & (!n_n1703) & (!x16080x)) + ((n_n4318) & (!n_n4331) & (n_n4279) & (!n_n1703) & (x16080x)) + ((n_n4318) & (!n_n4331) & (n_n4279) & (n_n1703) & (!x16080x)) + ((n_n4318) & (!n_n4331) & (n_n4279) & (n_n1703) & (x16080x)) + ((n_n4318) & (n_n4331) & (!n_n4279) & (!n_n1703) & (!x16080x)) + ((n_n4318) & (n_n4331) & (!n_n4279) & (!n_n1703) & (x16080x)) + ((n_n4318) & (n_n4331) & (!n_n4279) & (n_n1703) & (!x16080x)) + ((n_n4318) & (n_n4331) & (!n_n4279) & (n_n1703) & (x16080x)) + ((n_n4318) & (n_n4331) & (n_n4279) & (!n_n1703) & (!x16080x)) + ((n_n4318) & (n_n4331) & (n_n4279) & (!n_n1703) & (x16080x)) + ((n_n4318) & (n_n4331) & (n_n4279) & (n_n1703) & (!x16080x)) + ((n_n4318) & (n_n4331) & (n_n4279) & (n_n1703) & (x16080x)));
	assign n_n1818 = (((!n_n1890) & (!x16099x) & (!x16100x) & (x16105x)) + ((!n_n1890) & (!x16099x) & (x16100x) & (!x16105x)) + ((!n_n1890) & (!x16099x) & (x16100x) & (x16105x)) + ((!n_n1890) & (x16099x) & (!x16100x) & (!x16105x)) + ((!n_n1890) & (x16099x) & (!x16100x) & (x16105x)) + ((!n_n1890) & (x16099x) & (x16100x) & (!x16105x)) + ((!n_n1890) & (x16099x) & (x16100x) & (x16105x)) + ((n_n1890) & (!x16099x) & (!x16100x) & (!x16105x)) + ((n_n1890) & (!x16099x) & (!x16100x) & (x16105x)) + ((n_n1890) & (!x16099x) & (x16100x) & (!x16105x)) + ((n_n1890) & (!x16099x) & (x16100x) & (x16105x)) + ((n_n1890) & (x16099x) & (!x16100x) & (!x16105x)) + ((n_n1890) & (x16099x) & (!x16100x) & (x16105x)) + ((n_n1890) & (x16099x) & (x16100x) & (!x16105x)) + ((n_n1890) & (x16099x) & (x16100x) & (x16105x)));
	assign x16085x = (((!n_n4319) & (!n_n4321) & (!x364x) & (!x443x) & (x106x)) + ((!n_n4319) & (!n_n4321) & (!x364x) & (x443x) & (!x106x)) + ((!n_n4319) & (!n_n4321) & (!x364x) & (x443x) & (x106x)) + ((!n_n4319) & (!n_n4321) & (x364x) & (!x443x) & (!x106x)) + ((!n_n4319) & (!n_n4321) & (x364x) & (!x443x) & (x106x)) + ((!n_n4319) & (!n_n4321) & (x364x) & (x443x) & (!x106x)) + ((!n_n4319) & (!n_n4321) & (x364x) & (x443x) & (x106x)) + ((!n_n4319) & (n_n4321) & (!x364x) & (!x443x) & (!x106x)) + ((!n_n4319) & (n_n4321) & (!x364x) & (!x443x) & (x106x)) + ((!n_n4319) & (n_n4321) & (!x364x) & (x443x) & (!x106x)) + ((!n_n4319) & (n_n4321) & (!x364x) & (x443x) & (x106x)) + ((!n_n4319) & (n_n4321) & (x364x) & (!x443x) & (!x106x)) + ((!n_n4319) & (n_n4321) & (x364x) & (!x443x) & (x106x)) + ((!n_n4319) & (n_n4321) & (x364x) & (x443x) & (!x106x)) + ((!n_n4319) & (n_n4321) & (x364x) & (x443x) & (x106x)) + ((n_n4319) & (!n_n4321) & (!x364x) & (!x443x) & (!x106x)) + ((n_n4319) & (!n_n4321) & (!x364x) & (!x443x) & (x106x)) + ((n_n4319) & (!n_n4321) & (!x364x) & (x443x) & (!x106x)) + ((n_n4319) & (!n_n4321) & (!x364x) & (x443x) & (x106x)) + ((n_n4319) & (!n_n4321) & (x364x) & (!x443x) & (!x106x)) + ((n_n4319) & (!n_n4321) & (x364x) & (!x443x) & (x106x)) + ((n_n4319) & (!n_n4321) & (x364x) & (x443x) & (!x106x)) + ((n_n4319) & (!n_n4321) & (x364x) & (x443x) & (x106x)) + ((n_n4319) & (n_n4321) & (!x364x) & (!x443x) & (!x106x)) + ((n_n4319) & (n_n4321) & (!x364x) & (!x443x) & (x106x)) + ((n_n4319) & (n_n4321) & (!x364x) & (x443x) & (!x106x)) + ((n_n4319) & (n_n4321) & (!x364x) & (x443x) & (x106x)) + ((n_n4319) & (n_n4321) & (x364x) & (!x443x) & (!x106x)) + ((n_n4319) & (n_n4321) & (x364x) & (!x443x) & (x106x)) + ((n_n4319) & (n_n4321) & (x364x) & (x443x) & (!x106x)) + ((n_n4319) & (n_n4321) & (x364x) & (x443x) & (x106x)));
	assign n_n1867 = (((!n_n4735) & (!n_n4744) & (!x374x) & (!x22073x)) + ((!n_n4735) & (!n_n4744) & (x374x) & (!x22073x)) + ((!n_n4735) & (!n_n4744) & (x374x) & (x22073x)) + ((!n_n4735) & (n_n4744) & (!x374x) & (!x22073x)) + ((!n_n4735) & (n_n4744) & (!x374x) & (x22073x)) + ((!n_n4735) & (n_n4744) & (x374x) & (!x22073x)) + ((!n_n4735) & (n_n4744) & (x374x) & (x22073x)) + ((n_n4735) & (!n_n4744) & (!x374x) & (!x22073x)) + ((n_n4735) & (!n_n4744) & (!x374x) & (x22073x)) + ((n_n4735) & (!n_n4744) & (x374x) & (!x22073x)) + ((n_n4735) & (!n_n4744) & (x374x) & (x22073x)) + ((n_n4735) & (n_n4744) & (!x374x) & (!x22073x)) + ((n_n4735) & (n_n4744) & (!x374x) & (x22073x)) + ((n_n4735) & (n_n4744) & (x374x) & (!x22073x)) + ((n_n4735) & (n_n4744) & (x374x) & (x22073x)));
	assign n_n1866 = (((!n_n4751) & (!n_n4750) & (!n_n4745) & (!x258x) & (!x22072x)) + ((!n_n4751) & (!n_n4750) & (!n_n4745) & (x258x) & (!x22072x)) + ((!n_n4751) & (!n_n4750) & (!n_n4745) & (x258x) & (x22072x)) + ((!n_n4751) & (!n_n4750) & (n_n4745) & (!x258x) & (!x22072x)) + ((!n_n4751) & (!n_n4750) & (n_n4745) & (!x258x) & (x22072x)) + ((!n_n4751) & (!n_n4750) & (n_n4745) & (x258x) & (!x22072x)) + ((!n_n4751) & (!n_n4750) & (n_n4745) & (x258x) & (x22072x)) + ((!n_n4751) & (n_n4750) & (!n_n4745) & (!x258x) & (!x22072x)) + ((!n_n4751) & (n_n4750) & (!n_n4745) & (!x258x) & (x22072x)) + ((!n_n4751) & (n_n4750) & (!n_n4745) & (x258x) & (!x22072x)) + ((!n_n4751) & (n_n4750) & (!n_n4745) & (x258x) & (x22072x)) + ((!n_n4751) & (n_n4750) & (n_n4745) & (!x258x) & (!x22072x)) + ((!n_n4751) & (n_n4750) & (n_n4745) & (!x258x) & (x22072x)) + ((!n_n4751) & (n_n4750) & (n_n4745) & (x258x) & (!x22072x)) + ((!n_n4751) & (n_n4750) & (n_n4745) & (x258x) & (x22072x)) + ((n_n4751) & (!n_n4750) & (!n_n4745) & (!x258x) & (!x22072x)) + ((n_n4751) & (!n_n4750) & (!n_n4745) & (!x258x) & (x22072x)) + ((n_n4751) & (!n_n4750) & (!n_n4745) & (x258x) & (!x22072x)) + ((n_n4751) & (!n_n4750) & (!n_n4745) & (x258x) & (x22072x)) + ((n_n4751) & (!n_n4750) & (n_n4745) & (!x258x) & (!x22072x)) + ((n_n4751) & (!n_n4750) & (n_n4745) & (!x258x) & (x22072x)) + ((n_n4751) & (!n_n4750) & (n_n4745) & (x258x) & (!x22072x)) + ((n_n4751) & (!n_n4750) & (n_n4745) & (x258x) & (x22072x)) + ((n_n4751) & (n_n4750) & (!n_n4745) & (!x258x) & (!x22072x)) + ((n_n4751) & (n_n4750) & (!n_n4745) & (!x258x) & (x22072x)) + ((n_n4751) & (n_n4750) & (!n_n4745) & (x258x) & (!x22072x)) + ((n_n4751) & (n_n4750) & (!n_n4745) & (x258x) & (x22072x)) + ((n_n4751) & (n_n4750) & (n_n4745) & (!x258x) & (!x22072x)) + ((n_n4751) & (n_n4750) & (n_n4745) & (!x258x) & (x22072x)) + ((n_n4751) & (n_n4750) & (n_n4745) & (x258x) & (!x22072x)) + ((n_n4751) & (n_n4750) & (n_n4745) & (x258x) & (x22072x)));
	assign x16130x = (((!n_n4724) & (!n_n4723) & (!n_n4722) & (!x242x) & (!x22177x)) + ((!n_n4724) & (!n_n4723) & (!n_n4722) & (x242x) & (!x22177x)) + ((!n_n4724) & (!n_n4723) & (!n_n4722) & (x242x) & (x22177x)) + ((!n_n4724) & (!n_n4723) & (n_n4722) & (!x242x) & (!x22177x)) + ((!n_n4724) & (!n_n4723) & (n_n4722) & (!x242x) & (x22177x)) + ((!n_n4724) & (!n_n4723) & (n_n4722) & (x242x) & (!x22177x)) + ((!n_n4724) & (!n_n4723) & (n_n4722) & (x242x) & (x22177x)) + ((!n_n4724) & (n_n4723) & (!n_n4722) & (!x242x) & (!x22177x)) + ((!n_n4724) & (n_n4723) & (!n_n4722) & (!x242x) & (x22177x)) + ((!n_n4724) & (n_n4723) & (!n_n4722) & (x242x) & (!x22177x)) + ((!n_n4724) & (n_n4723) & (!n_n4722) & (x242x) & (x22177x)) + ((!n_n4724) & (n_n4723) & (n_n4722) & (!x242x) & (!x22177x)) + ((!n_n4724) & (n_n4723) & (n_n4722) & (!x242x) & (x22177x)) + ((!n_n4724) & (n_n4723) & (n_n4722) & (x242x) & (!x22177x)) + ((!n_n4724) & (n_n4723) & (n_n4722) & (x242x) & (x22177x)) + ((n_n4724) & (!n_n4723) & (!n_n4722) & (!x242x) & (!x22177x)) + ((n_n4724) & (!n_n4723) & (!n_n4722) & (!x242x) & (x22177x)) + ((n_n4724) & (!n_n4723) & (!n_n4722) & (x242x) & (!x22177x)) + ((n_n4724) & (!n_n4723) & (!n_n4722) & (x242x) & (x22177x)) + ((n_n4724) & (!n_n4723) & (n_n4722) & (!x242x) & (!x22177x)) + ((n_n4724) & (!n_n4723) & (n_n4722) & (!x242x) & (x22177x)) + ((n_n4724) & (!n_n4723) & (n_n4722) & (x242x) & (!x22177x)) + ((n_n4724) & (!n_n4723) & (n_n4722) & (x242x) & (x22177x)) + ((n_n4724) & (n_n4723) & (!n_n4722) & (!x242x) & (!x22177x)) + ((n_n4724) & (n_n4723) & (!n_n4722) & (!x242x) & (x22177x)) + ((n_n4724) & (n_n4723) & (!n_n4722) & (x242x) & (!x22177x)) + ((n_n4724) & (n_n4723) & (!n_n4722) & (x242x) & (x22177x)) + ((n_n4724) & (n_n4723) & (n_n4722) & (!x242x) & (!x22177x)) + ((n_n4724) & (n_n4723) & (n_n4722) & (!x242x) & (x22177x)) + ((n_n4724) & (n_n4723) & (n_n4722) & (x242x) & (!x22177x)) + ((n_n4724) & (n_n4723) & (n_n4722) & (x242x) & (x22177x)));
	assign n_n1811 = (((!x16135x) & (!x16144x) & (!x16141x) & (!x22071x)) + ((!x16135x) & (!x16144x) & (x16141x) & (!x22071x)) + ((!x16135x) & (!x16144x) & (x16141x) & (x22071x)) + ((!x16135x) & (x16144x) & (!x16141x) & (!x22071x)) + ((!x16135x) & (x16144x) & (!x16141x) & (x22071x)) + ((!x16135x) & (x16144x) & (x16141x) & (!x22071x)) + ((!x16135x) & (x16144x) & (x16141x) & (x22071x)) + ((x16135x) & (!x16144x) & (!x16141x) & (!x22071x)) + ((x16135x) & (!x16144x) & (!x16141x) & (x22071x)) + ((x16135x) & (!x16144x) & (x16141x) & (!x22071x)) + ((x16135x) & (!x16144x) & (x16141x) & (x22071x)) + ((x16135x) & (x16144x) & (!x16141x) & (!x22071x)) + ((x16135x) & (x16144x) & (!x16141x) & (x22071x)) + ((x16135x) & (x16144x) & (x16141x) & (!x22071x)) + ((x16135x) & (x16144x) & (x16141x) & (x22071x)));
	assign x16240x = (((!n_n1863) & (!x16233x) & (!x16234x) & (x16238x)) + ((!n_n1863) & (!x16233x) & (x16234x) & (!x16238x)) + ((!n_n1863) & (!x16233x) & (x16234x) & (x16238x)) + ((!n_n1863) & (x16233x) & (!x16234x) & (!x16238x)) + ((!n_n1863) & (x16233x) & (!x16234x) & (x16238x)) + ((!n_n1863) & (x16233x) & (x16234x) & (!x16238x)) + ((!n_n1863) & (x16233x) & (x16234x) & (x16238x)) + ((n_n1863) & (!x16233x) & (!x16234x) & (!x16238x)) + ((n_n1863) & (!x16233x) & (!x16234x) & (x16238x)) + ((n_n1863) & (!x16233x) & (x16234x) & (!x16238x)) + ((n_n1863) & (!x16233x) & (x16234x) & (x16238x)) + ((n_n1863) & (x16233x) & (!x16234x) & (!x16238x)) + ((n_n1863) & (x16233x) & (!x16234x) & (x16238x)) + ((n_n1863) & (x16233x) & (x16234x) & (!x16238x)) + ((n_n1863) & (x16233x) & (x16234x) & (x16238x)));
	assign x16242x = (((!n_n1867) & (!n_n1866) & (!x16130x) & (!n_n1811) & (x16240x)) + ((!n_n1867) & (!n_n1866) & (!x16130x) & (n_n1811) & (!x16240x)) + ((!n_n1867) & (!n_n1866) & (!x16130x) & (n_n1811) & (x16240x)) + ((!n_n1867) & (!n_n1866) & (x16130x) & (!n_n1811) & (!x16240x)) + ((!n_n1867) & (!n_n1866) & (x16130x) & (!n_n1811) & (x16240x)) + ((!n_n1867) & (!n_n1866) & (x16130x) & (n_n1811) & (!x16240x)) + ((!n_n1867) & (!n_n1866) & (x16130x) & (n_n1811) & (x16240x)) + ((!n_n1867) & (n_n1866) & (!x16130x) & (!n_n1811) & (!x16240x)) + ((!n_n1867) & (n_n1866) & (!x16130x) & (!n_n1811) & (x16240x)) + ((!n_n1867) & (n_n1866) & (!x16130x) & (n_n1811) & (!x16240x)) + ((!n_n1867) & (n_n1866) & (!x16130x) & (n_n1811) & (x16240x)) + ((!n_n1867) & (n_n1866) & (x16130x) & (!n_n1811) & (!x16240x)) + ((!n_n1867) & (n_n1866) & (x16130x) & (!n_n1811) & (x16240x)) + ((!n_n1867) & (n_n1866) & (x16130x) & (n_n1811) & (!x16240x)) + ((!n_n1867) & (n_n1866) & (x16130x) & (n_n1811) & (x16240x)) + ((n_n1867) & (!n_n1866) & (!x16130x) & (!n_n1811) & (!x16240x)) + ((n_n1867) & (!n_n1866) & (!x16130x) & (!n_n1811) & (x16240x)) + ((n_n1867) & (!n_n1866) & (!x16130x) & (n_n1811) & (!x16240x)) + ((n_n1867) & (!n_n1866) & (!x16130x) & (n_n1811) & (x16240x)) + ((n_n1867) & (!n_n1866) & (x16130x) & (!n_n1811) & (!x16240x)) + ((n_n1867) & (!n_n1866) & (x16130x) & (!n_n1811) & (x16240x)) + ((n_n1867) & (!n_n1866) & (x16130x) & (n_n1811) & (!x16240x)) + ((n_n1867) & (!n_n1866) & (x16130x) & (n_n1811) & (x16240x)) + ((n_n1867) & (n_n1866) & (!x16130x) & (!n_n1811) & (!x16240x)) + ((n_n1867) & (n_n1866) & (!x16130x) & (!n_n1811) & (x16240x)) + ((n_n1867) & (n_n1866) & (!x16130x) & (n_n1811) & (!x16240x)) + ((n_n1867) & (n_n1866) & (!x16130x) & (n_n1811) & (x16240x)) + ((n_n1867) & (n_n1866) & (x16130x) & (!n_n1811) & (!x16240x)) + ((n_n1867) & (n_n1866) & (x16130x) & (!n_n1811) & (x16240x)) + ((n_n1867) & (n_n1866) & (x16130x) & (n_n1811) & (!x16240x)) + ((n_n1867) & (n_n1866) & (x16130x) & (n_n1811) & (x16240x)));
	assign n_n1789 = (((!n_n1846) & (!x16157x) & (!n_n1805) & (!x16180x) & (x16156x)) + ((!n_n1846) & (!x16157x) & (!n_n1805) & (x16180x) & (!x16156x)) + ((!n_n1846) & (!x16157x) & (!n_n1805) & (x16180x) & (x16156x)) + ((!n_n1846) & (!x16157x) & (n_n1805) & (!x16180x) & (!x16156x)) + ((!n_n1846) & (!x16157x) & (n_n1805) & (!x16180x) & (x16156x)) + ((!n_n1846) & (!x16157x) & (n_n1805) & (x16180x) & (!x16156x)) + ((!n_n1846) & (!x16157x) & (n_n1805) & (x16180x) & (x16156x)) + ((!n_n1846) & (x16157x) & (!n_n1805) & (!x16180x) & (!x16156x)) + ((!n_n1846) & (x16157x) & (!n_n1805) & (!x16180x) & (x16156x)) + ((!n_n1846) & (x16157x) & (!n_n1805) & (x16180x) & (!x16156x)) + ((!n_n1846) & (x16157x) & (!n_n1805) & (x16180x) & (x16156x)) + ((!n_n1846) & (x16157x) & (n_n1805) & (!x16180x) & (!x16156x)) + ((!n_n1846) & (x16157x) & (n_n1805) & (!x16180x) & (x16156x)) + ((!n_n1846) & (x16157x) & (n_n1805) & (x16180x) & (!x16156x)) + ((!n_n1846) & (x16157x) & (n_n1805) & (x16180x) & (x16156x)) + ((n_n1846) & (!x16157x) & (!n_n1805) & (!x16180x) & (!x16156x)) + ((n_n1846) & (!x16157x) & (!n_n1805) & (!x16180x) & (x16156x)) + ((n_n1846) & (!x16157x) & (!n_n1805) & (x16180x) & (!x16156x)) + ((n_n1846) & (!x16157x) & (!n_n1805) & (x16180x) & (x16156x)) + ((n_n1846) & (!x16157x) & (n_n1805) & (!x16180x) & (!x16156x)) + ((n_n1846) & (!x16157x) & (n_n1805) & (!x16180x) & (x16156x)) + ((n_n1846) & (!x16157x) & (n_n1805) & (x16180x) & (!x16156x)) + ((n_n1846) & (!x16157x) & (n_n1805) & (x16180x) & (x16156x)) + ((n_n1846) & (x16157x) & (!n_n1805) & (!x16180x) & (!x16156x)) + ((n_n1846) & (x16157x) & (!n_n1805) & (!x16180x) & (x16156x)) + ((n_n1846) & (x16157x) & (!n_n1805) & (x16180x) & (!x16156x)) + ((n_n1846) & (x16157x) & (!n_n1805) & (x16180x) & (x16156x)) + ((n_n1846) & (x16157x) & (n_n1805) & (!x16180x) & (!x16156x)) + ((n_n1846) & (x16157x) & (n_n1805) & (!x16180x) & (x16156x)) + ((n_n1846) & (x16157x) & (n_n1805) & (x16180x) & (!x16156x)) + ((n_n1846) & (x16157x) & (n_n1805) & (x16180x) & (x16156x)));
	assign n_n1790 = (((!n_n1854) & (!n_n1808) & (!n_n1807) & (!n_n1856) & (x16222x)) + ((!n_n1854) & (!n_n1808) & (!n_n1807) & (n_n1856) & (!x16222x)) + ((!n_n1854) & (!n_n1808) & (!n_n1807) & (n_n1856) & (x16222x)) + ((!n_n1854) & (!n_n1808) & (n_n1807) & (!n_n1856) & (!x16222x)) + ((!n_n1854) & (!n_n1808) & (n_n1807) & (!n_n1856) & (x16222x)) + ((!n_n1854) & (!n_n1808) & (n_n1807) & (n_n1856) & (!x16222x)) + ((!n_n1854) & (!n_n1808) & (n_n1807) & (n_n1856) & (x16222x)) + ((!n_n1854) & (n_n1808) & (!n_n1807) & (!n_n1856) & (!x16222x)) + ((!n_n1854) & (n_n1808) & (!n_n1807) & (!n_n1856) & (x16222x)) + ((!n_n1854) & (n_n1808) & (!n_n1807) & (n_n1856) & (!x16222x)) + ((!n_n1854) & (n_n1808) & (!n_n1807) & (n_n1856) & (x16222x)) + ((!n_n1854) & (n_n1808) & (n_n1807) & (!n_n1856) & (!x16222x)) + ((!n_n1854) & (n_n1808) & (n_n1807) & (!n_n1856) & (x16222x)) + ((!n_n1854) & (n_n1808) & (n_n1807) & (n_n1856) & (!x16222x)) + ((!n_n1854) & (n_n1808) & (n_n1807) & (n_n1856) & (x16222x)) + ((n_n1854) & (!n_n1808) & (!n_n1807) & (!n_n1856) & (!x16222x)) + ((n_n1854) & (!n_n1808) & (!n_n1807) & (!n_n1856) & (x16222x)) + ((n_n1854) & (!n_n1808) & (!n_n1807) & (n_n1856) & (!x16222x)) + ((n_n1854) & (!n_n1808) & (!n_n1807) & (n_n1856) & (x16222x)) + ((n_n1854) & (!n_n1808) & (n_n1807) & (!n_n1856) & (!x16222x)) + ((n_n1854) & (!n_n1808) & (n_n1807) & (!n_n1856) & (x16222x)) + ((n_n1854) & (!n_n1808) & (n_n1807) & (n_n1856) & (!x16222x)) + ((n_n1854) & (!n_n1808) & (n_n1807) & (n_n1856) & (x16222x)) + ((n_n1854) & (n_n1808) & (!n_n1807) & (!n_n1856) & (!x16222x)) + ((n_n1854) & (n_n1808) & (!n_n1807) & (!n_n1856) & (x16222x)) + ((n_n1854) & (n_n1808) & (!n_n1807) & (n_n1856) & (!x16222x)) + ((n_n1854) & (n_n1808) & (!n_n1807) & (n_n1856) & (x16222x)) + ((n_n1854) & (n_n1808) & (n_n1807) & (!n_n1856) & (!x16222x)) + ((n_n1854) & (n_n1808) & (n_n1807) & (!n_n1856) & (x16222x)) + ((n_n1854) & (n_n1808) & (n_n1807) & (n_n1856) & (!x16222x)) + ((n_n1854) & (n_n1808) & (n_n1807) & (n_n1856) & (x16222x)));
	assign x466x = (((!n_n5156) & (!n_n5155) & (!n_n5157) & (!x195x) & (n_n5160)) + ((!n_n5156) & (!n_n5155) & (!n_n5157) & (x195x) & (!n_n5160)) + ((!n_n5156) & (!n_n5155) & (!n_n5157) & (x195x) & (n_n5160)) + ((!n_n5156) & (!n_n5155) & (n_n5157) & (!x195x) & (!n_n5160)) + ((!n_n5156) & (!n_n5155) & (n_n5157) & (!x195x) & (n_n5160)) + ((!n_n5156) & (!n_n5155) & (n_n5157) & (x195x) & (!n_n5160)) + ((!n_n5156) & (!n_n5155) & (n_n5157) & (x195x) & (n_n5160)) + ((!n_n5156) & (n_n5155) & (!n_n5157) & (!x195x) & (!n_n5160)) + ((!n_n5156) & (n_n5155) & (!n_n5157) & (!x195x) & (n_n5160)) + ((!n_n5156) & (n_n5155) & (!n_n5157) & (x195x) & (!n_n5160)) + ((!n_n5156) & (n_n5155) & (!n_n5157) & (x195x) & (n_n5160)) + ((!n_n5156) & (n_n5155) & (n_n5157) & (!x195x) & (!n_n5160)) + ((!n_n5156) & (n_n5155) & (n_n5157) & (!x195x) & (n_n5160)) + ((!n_n5156) & (n_n5155) & (n_n5157) & (x195x) & (!n_n5160)) + ((!n_n5156) & (n_n5155) & (n_n5157) & (x195x) & (n_n5160)) + ((n_n5156) & (!n_n5155) & (!n_n5157) & (!x195x) & (!n_n5160)) + ((n_n5156) & (!n_n5155) & (!n_n5157) & (!x195x) & (n_n5160)) + ((n_n5156) & (!n_n5155) & (!n_n5157) & (x195x) & (!n_n5160)) + ((n_n5156) & (!n_n5155) & (!n_n5157) & (x195x) & (n_n5160)) + ((n_n5156) & (!n_n5155) & (n_n5157) & (!x195x) & (!n_n5160)) + ((n_n5156) & (!n_n5155) & (n_n5157) & (!x195x) & (n_n5160)) + ((n_n5156) & (!n_n5155) & (n_n5157) & (x195x) & (!n_n5160)) + ((n_n5156) & (!n_n5155) & (n_n5157) & (x195x) & (n_n5160)) + ((n_n5156) & (n_n5155) & (!n_n5157) & (!x195x) & (!n_n5160)) + ((n_n5156) & (n_n5155) & (!n_n5157) & (!x195x) & (n_n5160)) + ((n_n5156) & (n_n5155) & (!n_n5157) & (x195x) & (!n_n5160)) + ((n_n5156) & (n_n5155) & (!n_n5157) & (x195x) & (n_n5160)) + ((n_n5156) & (n_n5155) & (n_n5157) & (!x195x) & (!n_n5160)) + ((n_n5156) & (n_n5155) & (n_n5157) & (!x195x) & (n_n5160)) + ((n_n5156) & (n_n5155) & (n_n5157) & (x195x) & (!n_n5160)) + ((n_n5156) & (n_n5155) & (n_n5157) & (x195x) & (n_n5160)));
	assign x16245x = (((!i_9_) & (n_n482) & (!n_n532) & (n_n534) & (n_n130)) + ((!i_9_) & (n_n482) & (n_n532) & (!n_n534) & (n_n130)) + ((!i_9_) & (n_n482) & (n_n532) & (n_n534) & (n_n130)) + ((i_9_) & (n_n482) & (n_n532) & (!n_n534) & (n_n130)) + ((i_9_) & (n_n482) & (n_n532) & (n_n534) & (n_n130)));
	assign n_n1833 = (((!n_n5174) & (!n_n5164) & (!n_n5170) & (!x254x) & (x16248x)) + ((!n_n5174) & (!n_n5164) & (!n_n5170) & (x254x) & (!x16248x)) + ((!n_n5174) & (!n_n5164) & (!n_n5170) & (x254x) & (x16248x)) + ((!n_n5174) & (!n_n5164) & (n_n5170) & (!x254x) & (!x16248x)) + ((!n_n5174) & (!n_n5164) & (n_n5170) & (!x254x) & (x16248x)) + ((!n_n5174) & (!n_n5164) & (n_n5170) & (x254x) & (!x16248x)) + ((!n_n5174) & (!n_n5164) & (n_n5170) & (x254x) & (x16248x)) + ((!n_n5174) & (n_n5164) & (!n_n5170) & (!x254x) & (!x16248x)) + ((!n_n5174) & (n_n5164) & (!n_n5170) & (!x254x) & (x16248x)) + ((!n_n5174) & (n_n5164) & (!n_n5170) & (x254x) & (!x16248x)) + ((!n_n5174) & (n_n5164) & (!n_n5170) & (x254x) & (x16248x)) + ((!n_n5174) & (n_n5164) & (n_n5170) & (!x254x) & (!x16248x)) + ((!n_n5174) & (n_n5164) & (n_n5170) & (!x254x) & (x16248x)) + ((!n_n5174) & (n_n5164) & (n_n5170) & (x254x) & (!x16248x)) + ((!n_n5174) & (n_n5164) & (n_n5170) & (x254x) & (x16248x)) + ((n_n5174) & (!n_n5164) & (!n_n5170) & (!x254x) & (!x16248x)) + ((n_n5174) & (!n_n5164) & (!n_n5170) & (!x254x) & (x16248x)) + ((n_n5174) & (!n_n5164) & (!n_n5170) & (x254x) & (!x16248x)) + ((n_n5174) & (!n_n5164) & (!n_n5170) & (x254x) & (x16248x)) + ((n_n5174) & (!n_n5164) & (n_n5170) & (!x254x) & (!x16248x)) + ((n_n5174) & (!n_n5164) & (n_n5170) & (!x254x) & (x16248x)) + ((n_n5174) & (!n_n5164) & (n_n5170) & (x254x) & (!x16248x)) + ((n_n5174) & (!n_n5164) & (n_n5170) & (x254x) & (x16248x)) + ((n_n5174) & (n_n5164) & (!n_n5170) & (!x254x) & (!x16248x)) + ((n_n5174) & (n_n5164) & (!n_n5170) & (!x254x) & (x16248x)) + ((n_n5174) & (n_n5164) & (!n_n5170) & (x254x) & (!x16248x)) + ((n_n5174) & (n_n5164) & (!n_n5170) & (x254x) & (x16248x)) + ((n_n5174) & (n_n5164) & (n_n5170) & (!x254x) & (!x16248x)) + ((n_n5174) & (n_n5164) & (n_n5170) & (!x254x) & (x16248x)) + ((n_n5174) & (n_n5164) & (n_n5170) & (x254x) & (!x16248x)) + ((n_n5174) & (n_n5164) & (n_n5170) & (x254x) & (x16248x)));
	assign x16287x = (((!n_n5142) & (!n_n5148) & (!x196x) & (!n_n5143) & (!x22077x)) + ((!n_n5142) & (!n_n5148) & (!x196x) & (n_n5143) & (!x22077x)) + ((!n_n5142) & (!n_n5148) & (!x196x) & (n_n5143) & (x22077x)) + ((!n_n5142) & (!n_n5148) & (x196x) & (!n_n5143) & (!x22077x)) + ((!n_n5142) & (!n_n5148) & (x196x) & (!n_n5143) & (x22077x)) + ((!n_n5142) & (!n_n5148) & (x196x) & (n_n5143) & (!x22077x)) + ((!n_n5142) & (!n_n5148) & (x196x) & (n_n5143) & (x22077x)) + ((!n_n5142) & (n_n5148) & (!x196x) & (!n_n5143) & (!x22077x)) + ((!n_n5142) & (n_n5148) & (!x196x) & (!n_n5143) & (x22077x)) + ((!n_n5142) & (n_n5148) & (!x196x) & (n_n5143) & (!x22077x)) + ((!n_n5142) & (n_n5148) & (!x196x) & (n_n5143) & (x22077x)) + ((!n_n5142) & (n_n5148) & (x196x) & (!n_n5143) & (!x22077x)) + ((!n_n5142) & (n_n5148) & (x196x) & (!n_n5143) & (x22077x)) + ((!n_n5142) & (n_n5148) & (x196x) & (n_n5143) & (!x22077x)) + ((!n_n5142) & (n_n5148) & (x196x) & (n_n5143) & (x22077x)) + ((n_n5142) & (!n_n5148) & (!x196x) & (!n_n5143) & (!x22077x)) + ((n_n5142) & (!n_n5148) & (!x196x) & (!n_n5143) & (x22077x)) + ((n_n5142) & (!n_n5148) & (!x196x) & (n_n5143) & (!x22077x)) + ((n_n5142) & (!n_n5148) & (!x196x) & (n_n5143) & (x22077x)) + ((n_n5142) & (!n_n5148) & (x196x) & (!n_n5143) & (!x22077x)) + ((n_n5142) & (!n_n5148) & (x196x) & (!n_n5143) & (x22077x)) + ((n_n5142) & (!n_n5148) & (x196x) & (n_n5143) & (!x22077x)) + ((n_n5142) & (!n_n5148) & (x196x) & (n_n5143) & (x22077x)) + ((n_n5142) & (n_n5148) & (!x196x) & (!n_n5143) & (!x22077x)) + ((n_n5142) & (n_n5148) & (!x196x) & (!n_n5143) & (x22077x)) + ((n_n5142) & (n_n5148) & (!x196x) & (n_n5143) & (!x22077x)) + ((n_n5142) & (n_n5148) & (!x196x) & (n_n5143) & (x22077x)) + ((n_n5142) & (n_n5148) & (x196x) & (!n_n5143) & (!x22077x)) + ((n_n5142) & (n_n5148) & (x196x) & (!n_n5143) & (x22077x)) + ((n_n5142) & (n_n5148) & (x196x) & (n_n5143) & (!x22077x)) + ((n_n5142) & (n_n5148) & (x196x) & (n_n5143) & (x22077x)));
	assign x16289x = (((!x466x) & (!x16245x) & (!n_n1833) & (x16287x)) + ((!x466x) & (!x16245x) & (n_n1833) & (!x16287x)) + ((!x466x) & (!x16245x) & (n_n1833) & (x16287x)) + ((!x466x) & (x16245x) & (!n_n1833) & (!x16287x)) + ((!x466x) & (x16245x) & (!n_n1833) & (x16287x)) + ((!x466x) & (x16245x) & (n_n1833) & (!x16287x)) + ((!x466x) & (x16245x) & (n_n1833) & (x16287x)) + ((x466x) & (!x16245x) & (!n_n1833) & (!x16287x)) + ((x466x) & (!x16245x) & (!n_n1833) & (x16287x)) + ((x466x) & (!x16245x) & (n_n1833) & (!x16287x)) + ((x466x) & (!x16245x) & (n_n1833) & (x16287x)) + ((x466x) & (x16245x) & (!n_n1833) & (!x16287x)) + ((x466x) & (x16245x) & (!n_n1833) & (x16287x)) + ((x466x) & (x16245x) & (n_n1833) & (!x16287x)) + ((x466x) & (x16245x) & (n_n1833) & (x16287x)));
	assign n_n1832 = (((!n_n5186) & (!n_n5187) & (!n_n5182) & (!x152x) & (!x22076x)) + ((!n_n5186) & (!n_n5187) & (!n_n5182) & (x152x) & (!x22076x)) + ((!n_n5186) & (!n_n5187) & (!n_n5182) & (x152x) & (x22076x)) + ((!n_n5186) & (!n_n5187) & (n_n5182) & (!x152x) & (!x22076x)) + ((!n_n5186) & (!n_n5187) & (n_n5182) & (!x152x) & (x22076x)) + ((!n_n5186) & (!n_n5187) & (n_n5182) & (x152x) & (!x22076x)) + ((!n_n5186) & (!n_n5187) & (n_n5182) & (x152x) & (x22076x)) + ((!n_n5186) & (n_n5187) & (!n_n5182) & (!x152x) & (!x22076x)) + ((!n_n5186) & (n_n5187) & (!n_n5182) & (!x152x) & (x22076x)) + ((!n_n5186) & (n_n5187) & (!n_n5182) & (x152x) & (!x22076x)) + ((!n_n5186) & (n_n5187) & (!n_n5182) & (x152x) & (x22076x)) + ((!n_n5186) & (n_n5187) & (n_n5182) & (!x152x) & (!x22076x)) + ((!n_n5186) & (n_n5187) & (n_n5182) & (!x152x) & (x22076x)) + ((!n_n5186) & (n_n5187) & (n_n5182) & (x152x) & (!x22076x)) + ((!n_n5186) & (n_n5187) & (n_n5182) & (x152x) & (x22076x)) + ((n_n5186) & (!n_n5187) & (!n_n5182) & (!x152x) & (!x22076x)) + ((n_n5186) & (!n_n5187) & (!n_n5182) & (!x152x) & (x22076x)) + ((n_n5186) & (!n_n5187) & (!n_n5182) & (x152x) & (!x22076x)) + ((n_n5186) & (!n_n5187) & (!n_n5182) & (x152x) & (x22076x)) + ((n_n5186) & (!n_n5187) & (n_n5182) & (!x152x) & (!x22076x)) + ((n_n5186) & (!n_n5187) & (n_n5182) & (!x152x) & (x22076x)) + ((n_n5186) & (!n_n5187) & (n_n5182) & (x152x) & (!x22076x)) + ((n_n5186) & (!n_n5187) & (n_n5182) & (x152x) & (x22076x)) + ((n_n5186) & (n_n5187) & (!n_n5182) & (!x152x) & (!x22076x)) + ((n_n5186) & (n_n5187) & (!n_n5182) & (!x152x) & (x22076x)) + ((n_n5186) & (n_n5187) & (!n_n5182) & (x152x) & (!x22076x)) + ((n_n5186) & (n_n5187) & (!n_n5182) & (x152x) & (x22076x)) + ((n_n5186) & (n_n5187) & (n_n5182) & (!x152x) & (!x22076x)) + ((n_n5186) & (n_n5187) & (n_n5182) & (!x152x) & (x22076x)) + ((n_n5186) & (n_n5187) & (n_n5182) & (x152x) & (!x22076x)) + ((n_n5186) & (n_n5187) & (n_n5182) & (x152x) & (x22076x)));
	assign x16262x = (((!n_n5212) & (!n_n5189) & (!n_n5194) & (!x453x) & (!x22218x)) + ((!n_n5212) & (!n_n5189) & (!n_n5194) & (x453x) & (!x22218x)) + ((!n_n5212) & (!n_n5189) & (!n_n5194) & (x453x) & (x22218x)) + ((!n_n5212) & (!n_n5189) & (n_n5194) & (!x453x) & (!x22218x)) + ((!n_n5212) & (!n_n5189) & (n_n5194) & (!x453x) & (x22218x)) + ((!n_n5212) & (!n_n5189) & (n_n5194) & (x453x) & (!x22218x)) + ((!n_n5212) & (!n_n5189) & (n_n5194) & (x453x) & (x22218x)) + ((!n_n5212) & (n_n5189) & (!n_n5194) & (!x453x) & (!x22218x)) + ((!n_n5212) & (n_n5189) & (!n_n5194) & (!x453x) & (x22218x)) + ((!n_n5212) & (n_n5189) & (!n_n5194) & (x453x) & (!x22218x)) + ((!n_n5212) & (n_n5189) & (!n_n5194) & (x453x) & (x22218x)) + ((!n_n5212) & (n_n5189) & (n_n5194) & (!x453x) & (!x22218x)) + ((!n_n5212) & (n_n5189) & (n_n5194) & (!x453x) & (x22218x)) + ((!n_n5212) & (n_n5189) & (n_n5194) & (x453x) & (!x22218x)) + ((!n_n5212) & (n_n5189) & (n_n5194) & (x453x) & (x22218x)) + ((n_n5212) & (!n_n5189) & (!n_n5194) & (!x453x) & (!x22218x)) + ((n_n5212) & (!n_n5189) & (!n_n5194) & (!x453x) & (x22218x)) + ((n_n5212) & (!n_n5189) & (!n_n5194) & (x453x) & (!x22218x)) + ((n_n5212) & (!n_n5189) & (!n_n5194) & (x453x) & (x22218x)) + ((n_n5212) & (!n_n5189) & (n_n5194) & (!x453x) & (!x22218x)) + ((n_n5212) & (!n_n5189) & (n_n5194) & (!x453x) & (x22218x)) + ((n_n5212) & (!n_n5189) & (n_n5194) & (x453x) & (!x22218x)) + ((n_n5212) & (!n_n5189) & (n_n5194) & (x453x) & (x22218x)) + ((n_n5212) & (n_n5189) & (!n_n5194) & (!x453x) & (!x22218x)) + ((n_n5212) & (n_n5189) & (!n_n5194) & (!x453x) & (x22218x)) + ((n_n5212) & (n_n5189) & (!n_n5194) & (x453x) & (!x22218x)) + ((n_n5212) & (n_n5189) & (!n_n5194) & (x453x) & (x22218x)) + ((n_n5212) & (n_n5189) & (n_n5194) & (!x453x) & (!x22218x)) + ((n_n5212) & (n_n5189) & (n_n5194) & (!x453x) & (x22218x)) + ((n_n5212) & (n_n5189) & (n_n5194) & (x453x) & (!x22218x)) + ((n_n5212) & (n_n5189) & (n_n5194) & (x453x) & (x22218x)));
	assign n_n1797 = (((!x16267x) & (!x16268x) & (!n_n1829) & (!x16278x) & (x16279x)) + ((!x16267x) & (!x16268x) & (!n_n1829) & (x16278x) & (!x16279x)) + ((!x16267x) & (!x16268x) & (!n_n1829) & (x16278x) & (x16279x)) + ((!x16267x) & (!x16268x) & (n_n1829) & (!x16278x) & (!x16279x)) + ((!x16267x) & (!x16268x) & (n_n1829) & (!x16278x) & (x16279x)) + ((!x16267x) & (!x16268x) & (n_n1829) & (x16278x) & (!x16279x)) + ((!x16267x) & (!x16268x) & (n_n1829) & (x16278x) & (x16279x)) + ((!x16267x) & (x16268x) & (!n_n1829) & (!x16278x) & (!x16279x)) + ((!x16267x) & (x16268x) & (!n_n1829) & (!x16278x) & (x16279x)) + ((!x16267x) & (x16268x) & (!n_n1829) & (x16278x) & (!x16279x)) + ((!x16267x) & (x16268x) & (!n_n1829) & (x16278x) & (x16279x)) + ((!x16267x) & (x16268x) & (n_n1829) & (!x16278x) & (!x16279x)) + ((!x16267x) & (x16268x) & (n_n1829) & (!x16278x) & (x16279x)) + ((!x16267x) & (x16268x) & (n_n1829) & (x16278x) & (!x16279x)) + ((!x16267x) & (x16268x) & (n_n1829) & (x16278x) & (x16279x)) + ((x16267x) & (!x16268x) & (!n_n1829) & (!x16278x) & (!x16279x)) + ((x16267x) & (!x16268x) & (!n_n1829) & (!x16278x) & (x16279x)) + ((x16267x) & (!x16268x) & (!n_n1829) & (x16278x) & (!x16279x)) + ((x16267x) & (!x16268x) & (!n_n1829) & (x16278x) & (x16279x)) + ((x16267x) & (!x16268x) & (n_n1829) & (!x16278x) & (!x16279x)) + ((x16267x) & (!x16268x) & (n_n1829) & (!x16278x) & (x16279x)) + ((x16267x) & (!x16268x) & (n_n1829) & (x16278x) & (!x16279x)) + ((x16267x) & (!x16268x) & (n_n1829) & (x16278x) & (x16279x)) + ((x16267x) & (x16268x) & (!n_n1829) & (!x16278x) & (!x16279x)) + ((x16267x) & (x16268x) & (!n_n1829) & (!x16278x) & (x16279x)) + ((x16267x) & (x16268x) & (!n_n1829) & (x16278x) & (!x16279x)) + ((x16267x) & (x16268x) & (!n_n1829) & (x16278x) & (x16279x)) + ((x16267x) & (x16268x) & (n_n1829) & (!x16278x) & (!x16279x)) + ((x16267x) & (x16268x) & (n_n1829) & (!x16278x) & (x16279x)) + ((x16267x) & (x16268x) & (n_n1829) & (x16278x) & (!x16279x)) + ((x16267x) & (x16268x) & (n_n1829) & (x16278x) & (x16279x)));
	assign x16261x = (((!n_n5191) & (!x220x) & (!x454x) & (!n_n5192) & (x452x)) + ((!n_n5191) & (!x220x) & (!x454x) & (n_n5192) & (!x452x)) + ((!n_n5191) & (!x220x) & (!x454x) & (n_n5192) & (x452x)) + ((!n_n5191) & (!x220x) & (x454x) & (!n_n5192) & (!x452x)) + ((!n_n5191) & (!x220x) & (x454x) & (!n_n5192) & (x452x)) + ((!n_n5191) & (!x220x) & (x454x) & (n_n5192) & (!x452x)) + ((!n_n5191) & (!x220x) & (x454x) & (n_n5192) & (x452x)) + ((!n_n5191) & (x220x) & (!x454x) & (!n_n5192) & (!x452x)) + ((!n_n5191) & (x220x) & (!x454x) & (!n_n5192) & (x452x)) + ((!n_n5191) & (x220x) & (!x454x) & (n_n5192) & (!x452x)) + ((!n_n5191) & (x220x) & (!x454x) & (n_n5192) & (x452x)) + ((!n_n5191) & (x220x) & (x454x) & (!n_n5192) & (!x452x)) + ((!n_n5191) & (x220x) & (x454x) & (!n_n5192) & (x452x)) + ((!n_n5191) & (x220x) & (x454x) & (n_n5192) & (!x452x)) + ((!n_n5191) & (x220x) & (x454x) & (n_n5192) & (x452x)) + ((n_n5191) & (!x220x) & (!x454x) & (!n_n5192) & (!x452x)) + ((n_n5191) & (!x220x) & (!x454x) & (!n_n5192) & (x452x)) + ((n_n5191) & (!x220x) & (!x454x) & (n_n5192) & (!x452x)) + ((n_n5191) & (!x220x) & (!x454x) & (n_n5192) & (x452x)) + ((n_n5191) & (!x220x) & (x454x) & (!n_n5192) & (!x452x)) + ((n_n5191) & (!x220x) & (x454x) & (!n_n5192) & (x452x)) + ((n_n5191) & (!x220x) & (x454x) & (n_n5192) & (!x452x)) + ((n_n5191) & (!x220x) & (x454x) & (n_n5192) & (x452x)) + ((n_n5191) & (x220x) & (!x454x) & (!n_n5192) & (!x452x)) + ((n_n5191) & (x220x) & (!x454x) & (!n_n5192) & (x452x)) + ((n_n5191) & (x220x) & (!x454x) & (n_n5192) & (!x452x)) + ((n_n5191) & (x220x) & (!x454x) & (n_n5192) & (x452x)) + ((n_n5191) & (x220x) & (x454x) & (!n_n5192) & (!x452x)) + ((n_n5191) & (x220x) & (x454x) & (!n_n5192) & (x452x)) + ((n_n5191) & (x220x) & (x454x) & (n_n5192) & (!x452x)) + ((n_n5191) & (x220x) & (x454x) & (n_n5192) & (x452x)));
	assign n_n5307 = (((!i_9_) & (n_n473) & (n_n532) & (n_n65)));
	assign n_n5308 = (((i_5_) & (!i_3_) & (!i_4_) & (x19x) & (n_n530)));
	assign x63x = (((!x19x) & (n_n482) & (!n_n522) & (x20x) & (n_n65)) + ((!x19x) & (n_n482) & (n_n522) & (x20x) & (n_n65)) + ((x19x) & (n_n482) & (!n_n522) & (x20x) & (n_n65)) + ((x19x) & (n_n482) & (n_n522) & (!x20x) & (!n_n65)) + ((x19x) & (n_n482) & (n_n522) & (!x20x) & (n_n65)) + ((x19x) & (n_n482) & (n_n522) & (x20x) & (!n_n65)) + ((x19x) & (n_n482) & (n_n522) & (x20x) & (n_n65)));
	assign x16315x = (((!n_n5319) & (!n_n5326) & (!n_n5332) & (!n_n5329) & (x117x)) + ((!n_n5319) & (!n_n5326) & (!n_n5332) & (n_n5329) & (!x117x)) + ((!n_n5319) & (!n_n5326) & (!n_n5332) & (n_n5329) & (x117x)) + ((!n_n5319) & (!n_n5326) & (n_n5332) & (!n_n5329) & (!x117x)) + ((!n_n5319) & (!n_n5326) & (n_n5332) & (!n_n5329) & (x117x)) + ((!n_n5319) & (!n_n5326) & (n_n5332) & (n_n5329) & (!x117x)) + ((!n_n5319) & (!n_n5326) & (n_n5332) & (n_n5329) & (x117x)) + ((!n_n5319) & (n_n5326) & (!n_n5332) & (!n_n5329) & (!x117x)) + ((!n_n5319) & (n_n5326) & (!n_n5332) & (!n_n5329) & (x117x)) + ((!n_n5319) & (n_n5326) & (!n_n5332) & (n_n5329) & (!x117x)) + ((!n_n5319) & (n_n5326) & (!n_n5332) & (n_n5329) & (x117x)) + ((!n_n5319) & (n_n5326) & (n_n5332) & (!n_n5329) & (!x117x)) + ((!n_n5319) & (n_n5326) & (n_n5332) & (!n_n5329) & (x117x)) + ((!n_n5319) & (n_n5326) & (n_n5332) & (n_n5329) & (!x117x)) + ((!n_n5319) & (n_n5326) & (n_n5332) & (n_n5329) & (x117x)) + ((n_n5319) & (!n_n5326) & (!n_n5332) & (!n_n5329) & (!x117x)) + ((n_n5319) & (!n_n5326) & (!n_n5332) & (!n_n5329) & (x117x)) + ((n_n5319) & (!n_n5326) & (!n_n5332) & (n_n5329) & (!x117x)) + ((n_n5319) & (!n_n5326) & (!n_n5332) & (n_n5329) & (x117x)) + ((n_n5319) & (!n_n5326) & (n_n5332) & (!n_n5329) & (!x117x)) + ((n_n5319) & (!n_n5326) & (n_n5332) & (!n_n5329) & (x117x)) + ((n_n5319) & (!n_n5326) & (n_n5332) & (n_n5329) & (!x117x)) + ((n_n5319) & (!n_n5326) & (n_n5332) & (n_n5329) & (x117x)) + ((n_n5319) & (n_n5326) & (!n_n5332) & (!n_n5329) & (!x117x)) + ((n_n5319) & (n_n5326) & (!n_n5332) & (!n_n5329) & (x117x)) + ((n_n5319) & (n_n5326) & (!n_n5332) & (n_n5329) & (!x117x)) + ((n_n5319) & (n_n5326) & (!n_n5332) & (n_n5329) & (x117x)) + ((n_n5319) & (n_n5326) & (n_n5332) & (!n_n5329) & (!x117x)) + ((n_n5319) & (n_n5326) & (n_n5332) & (!n_n5329) & (x117x)) + ((n_n5319) & (n_n5326) & (n_n5332) & (n_n5329) & (!x117x)) + ((n_n5319) & (n_n5326) & (n_n5332) & (n_n5329) & (x117x)));
	assign x22068x = (((!n_n5305) & (!n_n5310) & (!n_n5311) & (!n_n5309) & (!n_n5304)));
	assign x16318x = (((!n_n5307) & (!n_n5308) & (!x63x) & (!x16315x) & (!x22068x)) + ((!n_n5307) & (!n_n5308) & (!x63x) & (x16315x) & (!x22068x)) + ((!n_n5307) & (!n_n5308) & (!x63x) & (x16315x) & (x22068x)) + ((!n_n5307) & (!n_n5308) & (x63x) & (!x16315x) & (!x22068x)) + ((!n_n5307) & (!n_n5308) & (x63x) & (!x16315x) & (x22068x)) + ((!n_n5307) & (!n_n5308) & (x63x) & (x16315x) & (!x22068x)) + ((!n_n5307) & (!n_n5308) & (x63x) & (x16315x) & (x22068x)) + ((!n_n5307) & (n_n5308) & (!x63x) & (!x16315x) & (!x22068x)) + ((!n_n5307) & (n_n5308) & (!x63x) & (!x16315x) & (x22068x)) + ((!n_n5307) & (n_n5308) & (!x63x) & (x16315x) & (!x22068x)) + ((!n_n5307) & (n_n5308) & (!x63x) & (x16315x) & (x22068x)) + ((!n_n5307) & (n_n5308) & (x63x) & (!x16315x) & (!x22068x)) + ((!n_n5307) & (n_n5308) & (x63x) & (!x16315x) & (x22068x)) + ((!n_n5307) & (n_n5308) & (x63x) & (x16315x) & (!x22068x)) + ((!n_n5307) & (n_n5308) & (x63x) & (x16315x) & (x22068x)) + ((n_n5307) & (!n_n5308) & (!x63x) & (!x16315x) & (!x22068x)) + ((n_n5307) & (!n_n5308) & (!x63x) & (!x16315x) & (x22068x)) + ((n_n5307) & (!n_n5308) & (!x63x) & (x16315x) & (!x22068x)) + ((n_n5307) & (!n_n5308) & (!x63x) & (x16315x) & (x22068x)) + ((n_n5307) & (!n_n5308) & (x63x) & (!x16315x) & (!x22068x)) + ((n_n5307) & (!n_n5308) & (x63x) & (!x16315x) & (x22068x)) + ((n_n5307) & (!n_n5308) & (x63x) & (x16315x) & (!x22068x)) + ((n_n5307) & (!n_n5308) & (x63x) & (x16315x) & (x22068x)) + ((n_n5307) & (n_n5308) & (!x63x) & (!x16315x) & (!x22068x)) + ((n_n5307) & (n_n5308) & (!x63x) & (!x16315x) & (x22068x)) + ((n_n5307) & (n_n5308) & (!x63x) & (x16315x) & (!x22068x)) + ((n_n5307) & (n_n5308) & (!x63x) & (x16315x) & (x22068x)) + ((n_n5307) & (n_n5308) & (x63x) & (!x16315x) & (!x22068x)) + ((n_n5307) & (n_n5308) & (x63x) & (!x16315x) & (x22068x)) + ((n_n5307) & (n_n5308) & (x63x) & (x16315x) & (!x22068x)) + ((n_n5307) & (n_n5308) & (x63x) & (x16315x) & (x22068x)));
	assign n_n1825 = (((!n_n5284) & (!n_n5285) & (!n_n5279) & (!x218x) & (!x22067x)) + ((!n_n5284) & (!n_n5285) & (!n_n5279) & (x218x) & (!x22067x)) + ((!n_n5284) & (!n_n5285) & (!n_n5279) & (x218x) & (x22067x)) + ((!n_n5284) & (!n_n5285) & (n_n5279) & (!x218x) & (!x22067x)) + ((!n_n5284) & (!n_n5285) & (n_n5279) & (!x218x) & (x22067x)) + ((!n_n5284) & (!n_n5285) & (n_n5279) & (x218x) & (!x22067x)) + ((!n_n5284) & (!n_n5285) & (n_n5279) & (x218x) & (x22067x)) + ((!n_n5284) & (n_n5285) & (!n_n5279) & (!x218x) & (!x22067x)) + ((!n_n5284) & (n_n5285) & (!n_n5279) & (!x218x) & (x22067x)) + ((!n_n5284) & (n_n5285) & (!n_n5279) & (x218x) & (!x22067x)) + ((!n_n5284) & (n_n5285) & (!n_n5279) & (x218x) & (x22067x)) + ((!n_n5284) & (n_n5285) & (n_n5279) & (!x218x) & (!x22067x)) + ((!n_n5284) & (n_n5285) & (n_n5279) & (!x218x) & (x22067x)) + ((!n_n5284) & (n_n5285) & (n_n5279) & (x218x) & (!x22067x)) + ((!n_n5284) & (n_n5285) & (n_n5279) & (x218x) & (x22067x)) + ((n_n5284) & (!n_n5285) & (!n_n5279) & (!x218x) & (!x22067x)) + ((n_n5284) & (!n_n5285) & (!n_n5279) & (!x218x) & (x22067x)) + ((n_n5284) & (!n_n5285) & (!n_n5279) & (x218x) & (!x22067x)) + ((n_n5284) & (!n_n5285) & (!n_n5279) & (x218x) & (x22067x)) + ((n_n5284) & (!n_n5285) & (n_n5279) & (!x218x) & (!x22067x)) + ((n_n5284) & (!n_n5285) & (n_n5279) & (!x218x) & (x22067x)) + ((n_n5284) & (!n_n5285) & (n_n5279) & (x218x) & (!x22067x)) + ((n_n5284) & (!n_n5285) & (n_n5279) & (x218x) & (x22067x)) + ((n_n5284) & (n_n5285) & (!n_n5279) & (!x218x) & (!x22067x)) + ((n_n5284) & (n_n5285) & (!n_n5279) & (!x218x) & (x22067x)) + ((n_n5284) & (n_n5285) & (!n_n5279) & (x218x) & (!x22067x)) + ((n_n5284) & (n_n5285) & (!n_n5279) & (x218x) & (x22067x)) + ((n_n5284) & (n_n5285) & (n_n5279) & (!x218x) & (!x22067x)) + ((n_n5284) & (n_n5285) & (n_n5279) & (!x218x) & (x22067x)) + ((n_n5284) & (n_n5285) & (n_n5279) & (x218x) & (!x22067x)) + ((n_n5284) & (n_n5285) & (n_n5279) & (x218x) & (x22067x)));
	assign n_n1824 = (((!n_n5297) & (!n_n5298) & (!x197x) & (x16301x)) + ((!n_n5297) & (!n_n5298) & (x197x) & (!x16301x)) + ((!n_n5297) & (!n_n5298) & (x197x) & (x16301x)) + ((!n_n5297) & (n_n5298) & (!x197x) & (!x16301x)) + ((!n_n5297) & (n_n5298) & (!x197x) & (x16301x)) + ((!n_n5297) & (n_n5298) & (x197x) & (!x16301x)) + ((!n_n5297) & (n_n5298) & (x197x) & (x16301x)) + ((n_n5297) & (!n_n5298) & (!x197x) & (!x16301x)) + ((n_n5297) & (!n_n5298) & (!x197x) & (x16301x)) + ((n_n5297) & (!n_n5298) & (x197x) & (!x16301x)) + ((n_n5297) & (!n_n5298) & (x197x) & (x16301x)) + ((n_n5297) & (n_n5298) & (!x197x) & (!x16301x)) + ((n_n5297) & (n_n5298) & (!x197x) & (x16301x)) + ((n_n5297) & (n_n5298) & (x197x) & (!x16301x)) + ((n_n5297) & (n_n5298) & (x197x) & (x16301x)));
	assign n_n1826 = (((!n_n5264) & (!x77x) & (!x334x) & (!x203x) & (x16302x)) + ((!n_n5264) & (!x77x) & (!x334x) & (x203x) & (!x16302x)) + ((!n_n5264) & (!x77x) & (!x334x) & (x203x) & (x16302x)) + ((!n_n5264) & (!x77x) & (x334x) & (!x203x) & (!x16302x)) + ((!n_n5264) & (!x77x) & (x334x) & (!x203x) & (x16302x)) + ((!n_n5264) & (!x77x) & (x334x) & (x203x) & (!x16302x)) + ((!n_n5264) & (!x77x) & (x334x) & (x203x) & (x16302x)) + ((!n_n5264) & (x77x) & (!x334x) & (!x203x) & (!x16302x)) + ((!n_n5264) & (x77x) & (!x334x) & (!x203x) & (x16302x)) + ((!n_n5264) & (x77x) & (!x334x) & (x203x) & (!x16302x)) + ((!n_n5264) & (x77x) & (!x334x) & (x203x) & (x16302x)) + ((!n_n5264) & (x77x) & (x334x) & (!x203x) & (!x16302x)) + ((!n_n5264) & (x77x) & (x334x) & (!x203x) & (x16302x)) + ((!n_n5264) & (x77x) & (x334x) & (x203x) & (!x16302x)) + ((!n_n5264) & (x77x) & (x334x) & (x203x) & (x16302x)) + ((n_n5264) & (!x77x) & (!x334x) & (!x203x) & (!x16302x)) + ((n_n5264) & (!x77x) & (!x334x) & (!x203x) & (x16302x)) + ((n_n5264) & (!x77x) & (!x334x) & (x203x) & (!x16302x)) + ((n_n5264) & (!x77x) & (!x334x) & (x203x) & (x16302x)) + ((n_n5264) & (!x77x) & (x334x) & (!x203x) & (!x16302x)) + ((n_n5264) & (!x77x) & (x334x) & (!x203x) & (x16302x)) + ((n_n5264) & (!x77x) & (x334x) & (x203x) & (!x16302x)) + ((n_n5264) & (!x77x) & (x334x) & (x203x) & (x16302x)) + ((n_n5264) & (x77x) & (!x334x) & (!x203x) & (!x16302x)) + ((n_n5264) & (x77x) & (!x334x) & (!x203x) & (x16302x)) + ((n_n5264) & (x77x) & (!x334x) & (x203x) & (!x16302x)) + ((n_n5264) & (x77x) & (!x334x) & (x203x) & (x16302x)) + ((n_n5264) & (x77x) & (x334x) & (!x203x) & (!x16302x)) + ((n_n5264) & (x77x) & (x334x) & (!x203x) & (x16302x)) + ((n_n5264) & (x77x) & (x334x) & (x203x) & (!x16302x)) + ((n_n5264) & (x77x) & (x334x) & (x203x) & (x16302x)));
	assign x16314x = (((!x19x) & (!x516x) & (!x506x) & (!n_n5320) & (n_n1900)) + ((!x19x) & (!x516x) & (!x506x) & (n_n5320) & (!n_n1900)) + ((!x19x) & (!x516x) & (!x506x) & (n_n5320) & (n_n1900)) + ((!x19x) & (!x516x) & (x506x) & (!n_n5320) & (n_n1900)) + ((!x19x) & (!x516x) & (x506x) & (n_n5320) & (!n_n1900)) + ((!x19x) & (!x516x) & (x506x) & (n_n5320) & (n_n1900)) + ((!x19x) & (x516x) & (!x506x) & (!n_n5320) & (n_n1900)) + ((!x19x) & (x516x) & (!x506x) & (n_n5320) & (!n_n1900)) + ((!x19x) & (x516x) & (!x506x) & (n_n5320) & (n_n1900)) + ((!x19x) & (x516x) & (x506x) & (!n_n5320) & (n_n1900)) + ((!x19x) & (x516x) & (x506x) & (n_n5320) & (!n_n1900)) + ((!x19x) & (x516x) & (x506x) & (n_n5320) & (n_n1900)) + ((x19x) & (!x516x) & (!x506x) & (!n_n5320) & (n_n1900)) + ((x19x) & (!x516x) & (!x506x) & (n_n5320) & (!n_n1900)) + ((x19x) & (!x516x) & (!x506x) & (n_n5320) & (n_n1900)) + ((x19x) & (!x516x) & (x506x) & (!n_n5320) & (!n_n1900)) + ((x19x) & (!x516x) & (x506x) & (!n_n5320) & (n_n1900)) + ((x19x) & (!x516x) & (x506x) & (n_n5320) & (!n_n1900)) + ((x19x) & (!x516x) & (x506x) & (n_n5320) & (n_n1900)) + ((x19x) & (x516x) & (!x506x) & (!n_n5320) & (!n_n1900)) + ((x19x) & (x516x) & (!x506x) & (!n_n5320) & (n_n1900)) + ((x19x) & (x516x) & (!x506x) & (n_n5320) & (!n_n1900)) + ((x19x) & (x516x) & (!x506x) & (n_n5320) & (n_n1900)) + ((x19x) & (x516x) & (x506x) & (!n_n5320) & (!n_n1900)) + ((x19x) & (x516x) & (x506x) & (!n_n5320) & (n_n1900)) + ((x19x) & (x516x) & (x506x) & (n_n5320) & (!n_n1900)) + ((x19x) & (x516x) & (x506x) & (n_n5320) & (n_n1900)));
	assign x16319x = (((!n_n1825) & (!n_n1824) & (!n_n1826) & (x16314x)) + ((!n_n1825) & (!n_n1824) & (n_n1826) & (!x16314x)) + ((!n_n1825) & (!n_n1824) & (n_n1826) & (x16314x)) + ((!n_n1825) & (n_n1824) & (!n_n1826) & (!x16314x)) + ((!n_n1825) & (n_n1824) & (!n_n1826) & (x16314x)) + ((!n_n1825) & (n_n1824) & (n_n1826) & (!x16314x)) + ((!n_n1825) & (n_n1824) & (n_n1826) & (x16314x)) + ((n_n1825) & (!n_n1824) & (!n_n1826) & (!x16314x)) + ((n_n1825) & (!n_n1824) & (!n_n1826) & (x16314x)) + ((n_n1825) & (!n_n1824) & (n_n1826) & (!x16314x)) + ((n_n1825) & (!n_n1824) & (n_n1826) & (x16314x)) + ((n_n1825) & (n_n1824) & (!n_n1826) & (!x16314x)) + ((n_n1825) & (n_n1824) & (!n_n1826) & (x16314x)) + ((n_n1825) & (n_n1824) & (n_n1826) & (!x16314x)) + ((n_n1825) & (n_n1824) & (n_n1826) & (x16314x)));
	assign n_n2175 = (((!n_n2218) & (!x16435x) & (!x16436x) & (!x16440x) & (x16441x)) + ((!n_n2218) & (!x16435x) & (!x16436x) & (x16440x) & (!x16441x)) + ((!n_n2218) & (!x16435x) & (!x16436x) & (x16440x) & (x16441x)) + ((!n_n2218) & (!x16435x) & (x16436x) & (!x16440x) & (!x16441x)) + ((!n_n2218) & (!x16435x) & (x16436x) & (!x16440x) & (x16441x)) + ((!n_n2218) & (!x16435x) & (x16436x) & (x16440x) & (!x16441x)) + ((!n_n2218) & (!x16435x) & (x16436x) & (x16440x) & (x16441x)) + ((!n_n2218) & (x16435x) & (!x16436x) & (!x16440x) & (!x16441x)) + ((!n_n2218) & (x16435x) & (!x16436x) & (!x16440x) & (x16441x)) + ((!n_n2218) & (x16435x) & (!x16436x) & (x16440x) & (!x16441x)) + ((!n_n2218) & (x16435x) & (!x16436x) & (x16440x) & (x16441x)) + ((!n_n2218) & (x16435x) & (x16436x) & (!x16440x) & (!x16441x)) + ((!n_n2218) & (x16435x) & (x16436x) & (!x16440x) & (x16441x)) + ((!n_n2218) & (x16435x) & (x16436x) & (x16440x) & (!x16441x)) + ((!n_n2218) & (x16435x) & (x16436x) & (x16440x) & (x16441x)) + ((n_n2218) & (!x16435x) & (!x16436x) & (!x16440x) & (!x16441x)) + ((n_n2218) & (!x16435x) & (!x16436x) & (!x16440x) & (x16441x)) + ((n_n2218) & (!x16435x) & (!x16436x) & (x16440x) & (!x16441x)) + ((n_n2218) & (!x16435x) & (!x16436x) & (x16440x) & (x16441x)) + ((n_n2218) & (!x16435x) & (x16436x) & (!x16440x) & (!x16441x)) + ((n_n2218) & (!x16435x) & (x16436x) & (!x16440x) & (x16441x)) + ((n_n2218) & (!x16435x) & (x16436x) & (x16440x) & (!x16441x)) + ((n_n2218) & (!x16435x) & (x16436x) & (x16440x) & (x16441x)) + ((n_n2218) & (x16435x) & (!x16436x) & (!x16440x) & (!x16441x)) + ((n_n2218) & (x16435x) & (!x16436x) & (!x16440x) & (x16441x)) + ((n_n2218) & (x16435x) & (!x16436x) & (x16440x) & (!x16441x)) + ((n_n2218) & (x16435x) & (!x16436x) & (x16440x) & (x16441x)) + ((n_n2218) & (x16435x) & (x16436x) & (!x16440x) & (!x16441x)) + ((n_n2218) & (x16435x) & (x16436x) & (!x16440x) & (x16441x)) + ((n_n2218) & (x16435x) & (x16436x) & (x16440x) & (!x16441x)) + ((n_n2218) & (x16435x) & (x16436x) & (x16440x) & (x16441x)));
	assign x16456x = (((!x351x) & (!n_n4918) & (!n_n4917) & (!n_n4915) & (!x22064x)) + ((!x351x) & (!n_n4918) & (!n_n4917) & (n_n4915) & (!x22064x)) + ((!x351x) & (!n_n4918) & (!n_n4917) & (n_n4915) & (x22064x)) + ((!x351x) & (!n_n4918) & (n_n4917) & (!n_n4915) & (!x22064x)) + ((!x351x) & (!n_n4918) & (n_n4917) & (!n_n4915) & (x22064x)) + ((!x351x) & (!n_n4918) & (n_n4917) & (n_n4915) & (!x22064x)) + ((!x351x) & (!n_n4918) & (n_n4917) & (n_n4915) & (x22064x)) + ((!x351x) & (n_n4918) & (!n_n4917) & (!n_n4915) & (!x22064x)) + ((!x351x) & (n_n4918) & (!n_n4917) & (!n_n4915) & (x22064x)) + ((!x351x) & (n_n4918) & (!n_n4917) & (n_n4915) & (!x22064x)) + ((!x351x) & (n_n4918) & (!n_n4917) & (n_n4915) & (x22064x)) + ((!x351x) & (n_n4918) & (n_n4917) & (!n_n4915) & (!x22064x)) + ((!x351x) & (n_n4918) & (n_n4917) & (!n_n4915) & (x22064x)) + ((!x351x) & (n_n4918) & (n_n4917) & (n_n4915) & (!x22064x)) + ((!x351x) & (n_n4918) & (n_n4917) & (n_n4915) & (x22064x)) + ((x351x) & (!n_n4918) & (!n_n4917) & (!n_n4915) & (!x22064x)) + ((x351x) & (!n_n4918) & (!n_n4917) & (!n_n4915) & (x22064x)) + ((x351x) & (!n_n4918) & (!n_n4917) & (n_n4915) & (!x22064x)) + ((x351x) & (!n_n4918) & (!n_n4917) & (n_n4915) & (x22064x)) + ((x351x) & (!n_n4918) & (n_n4917) & (!n_n4915) & (!x22064x)) + ((x351x) & (!n_n4918) & (n_n4917) & (!n_n4915) & (x22064x)) + ((x351x) & (!n_n4918) & (n_n4917) & (n_n4915) & (!x22064x)) + ((x351x) & (!n_n4918) & (n_n4917) & (n_n4915) & (x22064x)) + ((x351x) & (n_n4918) & (!n_n4917) & (!n_n4915) & (!x22064x)) + ((x351x) & (n_n4918) & (!n_n4917) & (!n_n4915) & (x22064x)) + ((x351x) & (n_n4918) & (!n_n4917) & (n_n4915) & (!x22064x)) + ((x351x) & (n_n4918) & (!n_n4917) & (n_n4915) & (x22064x)) + ((x351x) & (n_n4918) & (n_n4917) & (!n_n4915) & (!x22064x)) + ((x351x) & (n_n4918) & (n_n4917) & (!n_n4915) & (x22064x)) + ((x351x) & (n_n4918) & (n_n4917) & (n_n4915) & (!x22064x)) + ((x351x) & (n_n4918) & (n_n4917) & (n_n4915) & (x22064x)));
	assign n_n2223 = (((!x31x) & (!n_n4937) & (!n_n4933) & (!n_n4935) & (x249x)) + ((!x31x) & (!n_n4937) & (!n_n4933) & (n_n4935) & (!x249x)) + ((!x31x) & (!n_n4937) & (!n_n4933) & (n_n4935) & (x249x)) + ((!x31x) & (!n_n4937) & (n_n4933) & (!n_n4935) & (!x249x)) + ((!x31x) & (!n_n4937) & (n_n4933) & (!n_n4935) & (x249x)) + ((!x31x) & (!n_n4937) & (n_n4933) & (n_n4935) & (!x249x)) + ((!x31x) & (!n_n4937) & (n_n4933) & (n_n4935) & (x249x)) + ((!x31x) & (n_n4937) & (!n_n4933) & (!n_n4935) & (!x249x)) + ((!x31x) & (n_n4937) & (!n_n4933) & (!n_n4935) & (x249x)) + ((!x31x) & (n_n4937) & (!n_n4933) & (n_n4935) & (!x249x)) + ((!x31x) & (n_n4937) & (!n_n4933) & (n_n4935) & (x249x)) + ((!x31x) & (n_n4937) & (n_n4933) & (!n_n4935) & (!x249x)) + ((!x31x) & (n_n4937) & (n_n4933) & (!n_n4935) & (x249x)) + ((!x31x) & (n_n4937) & (n_n4933) & (n_n4935) & (!x249x)) + ((!x31x) & (n_n4937) & (n_n4933) & (n_n4935) & (x249x)) + ((x31x) & (!n_n4937) & (!n_n4933) & (!n_n4935) & (!x249x)) + ((x31x) & (!n_n4937) & (!n_n4933) & (!n_n4935) & (x249x)) + ((x31x) & (!n_n4937) & (!n_n4933) & (n_n4935) & (!x249x)) + ((x31x) & (!n_n4937) & (!n_n4933) & (n_n4935) & (x249x)) + ((x31x) & (!n_n4937) & (n_n4933) & (!n_n4935) & (!x249x)) + ((x31x) & (!n_n4937) & (n_n4933) & (!n_n4935) & (x249x)) + ((x31x) & (!n_n4937) & (n_n4933) & (n_n4935) & (!x249x)) + ((x31x) & (!n_n4937) & (n_n4933) & (n_n4935) & (x249x)) + ((x31x) & (n_n4937) & (!n_n4933) & (!n_n4935) & (!x249x)) + ((x31x) & (n_n4937) & (!n_n4933) & (!n_n4935) & (x249x)) + ((x31x) & (n_n4937) & (!n_n4933) & (n_n4935) & (!x249x)) + ((x31x) & (n_n4937) & (!n_n4933) & (n_n4935) & (x249x)) + ((x31x) & (n_n4937) & (n_n4933) & (!n_n4935) & (!x249x)) + ((x31x) & (n_n4937) & (n_n4933) & (!n_n4935) & (x249x)) + ((x31x) & (n_n4937) & (n_n4933) & (n_n4935) & (!x249x)) + ((x31x) & (n_n4937) & (n_n4933) & (n_n4935) & (x249x)));
	assign n_n2225 = (((!n_n4901) & (!n_n4903) & (!x226x) & (!n_n3810) & (x16447x)) + ((!n_n4901) & (!n_n4903) & (!x226x) & (n_n3810) & (!x16447x)) + ((!n_n4901) & (!n_n4903) & (!x226x) & (n_n3810) & (x16447x)) + ((!n_n4901) & (!n_n4903) & (x226x) & (!n_n3810) & (!x16447x)) + ((!n_n4901) & (!n_n4903) & (x226x) & (!n_n3810) & (x16447x)) + ((!n_n4901) & (!n_n4903) & (x226x) & (n_n3810) & (!x16447x)) + ((!n_n4901) & (!n_n4903) & (x226x) & (n_n3810) & (x16447x)) + ((!n_n4901) & (n_n4903) & (!x226x) & (!n_n3810) & (!x16447x)) + ((!n_n4901) & (n_n4903) & (!x226x) & (!n_n3810) & (x16447x)) + ((!n_n4901) & (n_n4903) & (!x226x) & (n_n3810) & (!x16447x)) + ((!n_n4901) & (n_n4903) & (!x226x) & (n_n3810) & (x16447x)) + ((!n_n4901) & (n_n4903) & (x226x) & (!n_n3810) & (!x16447x)) + ((!n_n4901) & (n_n4903) & (x226x) & (!n_n3810) & (x16447x)) + ((!n_n4901) & (n_n4903) & (x226x) & (n_n3810) & (!x16447x)) + ((!n_n4901) & (n_n4903) & (x226x) & (n_n3810) & (x16447x)) + ((n_n4901) & (!n_n4903) & (!x226x) & (!n_n3810) & (!x16447x)) + ((n_n4901) & (!n_n4903) & (!x226x) & (!n_n3810) & (x16447x)) + ((n_n4901) & (!n_n4903) & (!x226x) & (n_n3810) & (!x16447x)) + ((n_n4901) & (!n_n4903) & (!x226x) & (n_n3810) & (x16447x)) + ((n_n4901) & (!n_n4903) & (x226x) & (!n_n3810) & (!x16447x)) + ((n_n4901) & (!n_n4903) & (x226x) & (!n_n3810) & (x16447x)) + ((n_n4901) & (!n_n4903) & (x226x) & (n_n3810) & (!x16447x)) + ((n_n4901) & (!n_n4903) & (x226x) & (n_n3810) & (x16447x)) + ((n_n4901) & (n_n4903) & (!x226x) & (!n_n3810) & (!x16447x)) + ((n_n4901) & (n_n4903) & (!x226x) & (!n_n3810) & (x16447x)) + ((n_n4901) & (n_n4903) & (!x226x) & (n_n3810) & (!x16447x)) + ((n_n4901) & (n_n4903) & (!x226x) & (n_n3810) & (x16447x)) + ((n_n4901) & (n_n4903) & (x226x) & (!n_n3810) & (!x16447x)) + ((n_n4901) & (n_n4903) & (x226x) & (!n_n3810) & (x16447x)) + ((n_n4901) & (n_n4903) & (x226x) & (n_n3810) & (!x16447x)) + ((n_n4901) & (n_n4903) & (x226x) & (n_n3810) & (x16447x)));
	assign x16468x = (((!n_n3803) & (!n_n3805) & (!x16327x) & (!n_n2220) & (x16466x)) + ((!n_n3803) & (!n_n3805) & (!x16327x) & (n_n2220) & (!x16466x)) + ((!n_n3803) & (!n_n3805) & (!x16327x) & (n_n2220) & (x16466x)) + ((!n_n3803) & (!n_n3805) & (x16327x) & (!n_n2220) & (!x16466x)) + ((!n_n3803) & (!n_n3805) & (x16327x) & (!n_n2220) & (x16466x)) + ((!n_n3803) & (!n_n3805) & (x16327x) & (n_n2220) & (!x16466x)) + ((!n_n3803) & (!n_n3805) & (x16327x) & (n_n2220) & (x16466x)) + ((!n_n3803) & (n_n3805) & (!x16327x) & (!n_n2220) & (!x16466x)) + ((!n_n3803) & (n_n3805) & (!x16327x) & (!n_n2220) & (x16466x)) + ((!n_n3803) & (n_n3805) & (!x16327x) & (n_n2220) & (!x16466x)) + ((!n_n3803) & (n_n3805) & (!x16327x) & (n_n2220) & (x16466x)) + ((!n_n3803) & (n_n3805) & (x16327x) & (!n_n2220) & (!x16466x)) + ((!n_n3803) & (n_n3805) & (x16327x) & (!n_n2220) & (x16466x)) + ((!n_n3803) & (n_n3805) & (x16327x) & (n_n2220) & (!x16466x)) + ((!n_n3803) & (n_n3805) & (x16327x) & (n_n2220) & (x16466x)) + ((n_n3803) & (!n_n3805) & (!x16327x) & (!n_n2220) & (!x16466x)) + ((n_n3803) & (!n_n3805) & (!x16327x) & (!n_n2220) & (x16466x)) + ((n_n3803) & (!n_n3805) & (!x16327x) & (n_n2220) & (!x16466x)) + ((n_n3803) & (!n_n3805) & (!x16327x) & (n_n2220) & (x16466x)) + ((n_n3803) & (!n_n3805) & (x16327x) & (!n_n2220) & (!x16466x)) + ((n_n3803) & (!n_n3805) & (x16327x) & (!n_n2220) & (x16466x)) + ((n_n3803) & (!n_n3805) & (x16327x) & (n_n2220) & (!x16466x)) + ((n_n3803) & (!n_n3805) & (x16327x) & (n_n2220) & (x16466x)) + ((n_n3803) & (n_n3805) & (!x16327x) & (!n_n2220) & (!x16466x)) + ((n_n3803) & (n_n3805) & (!x16327x) & (!n_n2220) & (x16466x)) + ((n_n3803) & (n_n3805) & (!x16327x) & (n_n2220) & (!x16466x)) + ((n_n3803) & (n_n3805) & (!x16327x) & (n_n2220) & (x16466x)) + ((n_n3803) & (n_n3805) & (x16327x) & (!n_n2220) & (!x16466x)) + ((n_n3803) & (n_n3805) & (x16327x) & (!n_n2220) & (x16466x)) + ((n_n3803) & (n_n3805) & (x16327x) & (n_n2220) & (!x16466x)) + ((n_n3803) & (n_n3805) & (x16327x) & (n_n2220) & (x16466x)));
	assign n_n4400 = (((i_9_) & (n_n536) & (n_n526) & (n_n482)));
	assign x16476x = (((!n_n4400) & (!n_n4389) & (!n_n4420) & (n_n4407)) + ((!n_n4400) & (!n_n4389) & (n_n4420) & (!n_n4407)) + ((!n_n4400) & (!n_n4389) & (n_n4420) & (n_n4407)) + ((!n_n4400) & (n_n4389) & (!n_n4420) & (!n_n4407)) + ((!n_n4400) & (n_n4389) & (!n_n4420) & (n_n4407)) + ((!n_n4400) & (n_n4389) & (n_n4420) & (!n_n4407)) + ((!n_n4400) & (n_n4389) & (n_n4420) & (n_n4407)) + ((n_n4400) & (!n_n4389) & (!n_n4420) & (!n_n4407)) + ((n_n4400) & (!n_n4389) & (!n_n4420) & (n_n4407)) + ((n_n4400) & (!n_n4389) & (n_n4420) & (!n_n4407)) + ((n_n4400) & (!n_n4389) & (n_n4420) & (n_n4407)) + ((n_n4400) & (n_n4389) & (!n_n4420) & (!n_n4407)) + ((n_n4400) & (n_n4389) & (!n_n4420) & (n_n4407)) + ((n_n4400) & (n_n4389) & (n_n4420) & (!n_n4407)) + ((n_n4400) & (n_n4389) & (n_n4420) & (n_n4407)));
	assign n_n4416 = (((i_9_) & (n_n536) & (n_n526) & (n_n473)));
	assign n_n4405 = (((i_1_) & (i_2_) & (i_0_) & (n_n482) & (x20x)));
	assign n_n4406 = (((i_9_) & (n_n536) & (n_n482) & (n_n520)));
	assign x16477x = (((!n_n4416) & (!n_n4404) & (!n_n4413) & (!n_n4405) & (n_n4406)) + ((!n_n4416) & (!n_n4404) & (!n_n4413) & (n_n4405) & (!n_n4406)) + ((!n_n4416) & (!n_n4404) & (!n_n4413) & (n_n4405) & (n_n4406)) + ((!n_n4416) & (!n_n4404) & (n_n4413) & (!n_n4405) & (!n_n4406)) + ((!n_n4416) & (!n_n4404) & (n_n4413) & (!n_n4405) & (n_n4406)) + ((!n_n4416) & (!n_n4404) & (n_n4413) & (n_n4405) & (!n_n4406)) + ((!n_n4416) & (!n_n4404) & (n_n4413) & (n_n4405) & (n_n4406)) + ((!n_n4416) & (n_n4404) & (!n_n4413) & (!n_n4405) & (!n_n4406)) + ((!n_n4416) & (n_n4404) & (!n_n4413) & (!n_n4405) & (n_n4406)) + ((!n_n4416) & (n_n4404) & (!n_n4413) & (n_n4405) & (!n_n4406)) + ((!n_n4416) & (n_n4404) & (!n_n4413) & (n_n4405) & (n_n4406)) + ((!n_n4416) & (n_n4404) & (n_n4413) & (!n_n4405) & (!n_n4406)) + ((!n_n4416) & (n_n4404) & (n_n4413) & (!n_n4405) & (n_n4406)) + ((!n_n4416) & (n_n4404) & (n_n4413) & (n_n4405) & (!n_n4406)) + ((!n_n4416) & (n_n4404) & (n_n4413) & (n_n4405) & (n_n4406)) + ((n_n4416) & (!n_n4404) & (!n_n4413) & (!n_n4405) & (!n_n4406)) + ((n_n4416) & (!n_n4404) & (!n_n4413) & (!n_n4405) & (n_n4406)) + ((n_n4416) & (!n_n4404) & (!n_n4413) & (n_n4405) & (!n_n4406)) + ((n_n4416) & (!n_n4404) & (!n_n4413) & (n_n4405) & (n_n4406)) + ((n_n4416) & (!n_n4404) & (n_n4413) & (!n_n4405) & (!n_n4406)) + ((n_n4416) & (!n_n4404) & (n_n4413) & (!n_n4405) & (n_n4406)) + ((n_n4416) & (!n_n4404) & (n_n4413) & (n_n4405) & (!n_n4406)) + ((n_n4416) & (!n_n4404) & (n_n4413) & (n_n4405) & (n_n4406)) + ((n_n4416) & (n_n4404) & (!n_n4413) & (!n_n4405) & (!n_n4406)) + ((n_n4416) & (n_n4404) & (!n_n4413) & (!n_n4405) & (n_n4406)) + ((n_n4416) & (n_n4404) & (!n_n4413) & (n_n4405) & (!n_n4406)) + ((n_n4416) & (n_n4404) & (!n_n4413) & (n_n4405) & (n_n4406)) + ((n_n4416) & (n_n4404) & (n_n4413) & (!n_n4405) & (!n_n4406)) + ((n_n4416) & (n_n4404) & (n_n4413) & (!n_n4405) & (n_n4406)) + ((n_n4416) & (n_n4404) & (n_n4413) & (n_n4405) & (!n_n4406)) + ((n_n4416) & (n_n4404) & (n_n4413) & (n_n4405) & (n_n4406)));
	assign n_n2102 = (((!n_n4513) & (!x16483x) & (!n_n4518) & (!n_n4492) & (n_n4496)) + ((!n_n4513) & (!x16483x) & (!n_n4518) & (n_n4492) & (!n_n4496)) + ((!n_n4513) & (!x16483x) & (!n_n4518) & (n_n4492) & (n_n4496)) + ((!n_n4513) & (!x16483x) & (n_n4518) & (!n_n4492) & (!n_n4496)) + ((!n_n4513) & (!x16483x) & (n_n4518) & (!n_n4492) & (n_n4496)) + ((!n_n4513) & (!x16483x) & (n_n4518) & (n_n4492) & (!n_n4496)) + ((!n_n4513) & (!x16483x) & (n_n4518) & (n_n4492) & (n_n4496)) + ((!n_n4513) & (x16483x) & (!n_n4518) & (!n_n4492) & (!n_n4496)) + ((!n_n4513) & (x16483x) & (!n_n4518) & (!n_n4492) & (n_n4496)) + ((!n_n4513) & (x16483x) & (!n_n4518) & (n_n4492) & (!n_n4496)) + ((!n_n4513) & (x16483x) & (!n_n4518) & (n_n4492) & (n_n4496)) + ((!n_n4513) & (x16483x) & (n_n4518) & (!n_n4492) & (!n_n4496)) + ((!n_n4513) & (x16483x) & (n_n4518) & (!n_n4492) & (n_n4496)) + ((!n_n4513) & (x16483x) & (n_n4518) & (n_n4492) & (!n_n4496)) + ((!n_n4513) & (x16483x) & (n_n4518) & (n_n4492) & (n_n4496)) + ((n_n4513) & (!x16483x) & (!n_n4518) & (!n_n4492) & (!n_n4496)) + ((n_n4513) & (!x16483x) & (!n_n4518) & (!n_n4492) & (n_n4496)) + ((n_n4513) & (!x16483x) & (!n_n4518) & (n_n4492) & (!n_n4496)) + ((n_n4513) & (!x16483x) & (!n_n4518) & (n_n4492) & (n_n4496)) + ((n_n4513) & (!x16483x) & (n_n4518) & (!n_n4492) & (!n_n4496)) + ((n_n4513) & (!x16483x) & (n_n4518) & (!n_n4492) & (n_n4496)) + ((n_n4513) & (!x16483x) & (n_n4518) & (n_n4492) & (!n_n4496)) + ((n_n4513) & (!x16483x) & (n_n4518) & (n_n4492) & (n_n4496)) + ((n_n4513) & (x16483x) & (!n_n4518) & (!n_n4492) & (!n_n4496)) + ((n_n4513) & (x16483x) & (!n_n4518) & (!n_n4492) & (n_n4496)) + ((n_n4513) & (x16483x) & (!n_n4518) & (n_n4492) & (!n_n4496)) + ((n_n4513) & (x16483x) & (!n_n4518) & (n_n4492) & (n_n4496)) + ((n_n4513) & (x16483x) & (n_n4518) & (!n_n4492) & (!n_n4496)) + ((n_n4513) & (x16483x) & (n_n4518) & (!n_n4492) & (n_n4496)) + ((n_n4513) & (x16483x) & (n_n4518) & (n_n4492) & (!n_n4496)) + ((n_n4513) & (x16483x) & (n_n4518) & (n_n4492) & (n_n4496)));
	assign x16487x = (((!n_n4617) & (!n_n4612) & (!n_n4574) & (n_n4572)) + ((!n_n4617) & (!n_n4612) & (n_n4574) & (!n_n4572)) + ((!n_n4617) & (!n_n4612) & (n_n4574) & (n_n4572)) + ((!n_n4617) & (n_n4612) & (!n_n4574) & (!n_n4572)) + ((!n_n4617) & (n_n4612) & (!n_n4574) & (n_n4572)) + ((!n_n4617) & (n_n4612) & (n_n4574) & (!n_n4572)) + ((!n_n4617) & (n_n4612) & (n_n4574) & (n_n4572)) + ((n_n4617) & (!n_n4612) & (!n_n4574) & (!n_n4572)) + ((n_n4617) & (!n_n4612) & (!n_n4574) & (n_n4572)) + ((n_n4617) & (!n_n4612) & (n_n4574) & (!n_n4572)) + ((n_n4617) & (!n_n4612) & (n_n4574) & (n_n4572)) + ((n_n4617) & (n_n4612) & (!n_n4574) & (!n_n4572)) + ((n_n4617) & (n_n4612) & (!n_n4574) & (n_n4572)) + ((n_n4617) & (n_n4612) & (n_n4574) & (!n_n4572)) + ((n_n4617) & (n_n4612) & (n_n4574) & (n_n4572)));
	assign x16488x = (((!n_n4640) & (!n_n4581) & (!x256x) & (n_n4623)) + ((!n_n4640) & (!n_n4581) & (x256x) & (!n_n4623)) + ((!n_n4640) & (!n_n4581) & (x256x) & (n_n4623)) + ((!n_n4640) & (n_n4581) & (!x256x) & (!n_n4623)) + ((!n_n4640) & (n_n4581) & (!x256x) & (n_n4623)) + ((!n_n4640) & (n_n4581) & (x256x) & (!n_n4623)) + ((!n_n4640) & (n_n4581) & (x256x) & (n_n4623)) + ((n_n4640) & (!n_n4581) & (!x256x) & (!n_n4623)) + ((n_n4640) & (!n_n4581) & (!x256x) & (n_n4623)) + ((n_n4640) & (!n_n4581) & (x256x) & (!n_n4623)) + ((n_n4640) & (!n_n4581) & (x256x) & (n_n4623)) + ((n_n4640) & (n_n4581) & (!x256x) & (!n_n4623)) + ((n_n4640) & (n_n4581) & (!x256x) & (n_n4623)) + ((n_n4640) & (n_n4581) & (x256x) & (!n_n4623)) + ((n_n4640) & (n_n4581) & (x256x) & (n_n4623)));
	assign x16494x = (((!n_n4547) & (!n_n4539) & (!n_n4521) & (n_n4544)) + ((!n_n4547) & (!n_n4539) & (n_n4521) & (!n_n4544)) + ((!n_n4547) & (!n_n4539) & (n_n4521) & (n_n4544)) + ((!n_n4547) & (n_n4539) & (!n_n4521) & (!n_n4544)) + ((!n_n4547) & (n_n4539) & (!n_n4521) & (n_n4544)) + ((!n_n4547) & (n_n4539) & (n_n4521) & (!n_n4544)) + ((!n_n4547) & (n_n4539) & (n_n4521) & (n_n4544)) + ((n_n4547) & (!n_n4539) & (!n_n4521) & (!n_n4544)) + ((n_n4547) & (!n_n4539) & (!n_n4521) & (n_n4544)) + ((n_n4547) & (!n_n4539) & (n_n4521) & (!n_n4544)) + ((n_n4547) & (!n_n4539) & (n_n4521) & (n_n4544)) + ((n_n4547) & (n_n4539) & (!n_n4521) & (!n_n4544)) + ((n_n4547) & (n_n4539) & (!n_n4521) & (n_n4544)) + ((n_n4547) & (n_n4539) & (n_n4521) & (!n_n4544)) + ((n_n4547) & (n_n4539) & (n_n4521) & (n_n4544)));
	assign x16495x = (((!n_n4571) & (!n_n4523) & (!n_n4557) & (!n_n4560) & (n_n4553)) + ((!n_n4571) & (!n_n4523) & (!n_n4557) & (n_n4560) & (!n_n4553)) + ((!n_n4571) & (!n_n4523) & (!n_n4557) & (n_n4560) & (n_n4553)) + ((!n_n4571) & (!n_n4523) & (n_n4557) & (!n_n4560) & (!n_n4553)) + ((!n_n4571) & (!n_n4523) & (n_n4557) & (!n_n4560) & (n_n4553)) + ((!n_n4571) & (!n_n4523) & (n_n4557) & (n_n4560) & (!n_n4553)) + ((!n_n4571) & (!n_n4523) & (n_n4557) & (n_n4560) & (n_n4553)) + ((!n_n4571) & (n_n4523) & (!n_n4557) & (!n_n4560) & (!n_n4553)) + ((!n_n4571) & (n_n4523) & (!n_n4557) & (!n_n4560) & (n_n4553)) + ((!n_n4571) & (n_n4523) & (!n_n4557) & (n_n4560) & (!n_n4553)) + ((!n_n4571) & (n_n4523) & (!n_n4557) & (n_n4560) & (n_n4553)) + ((!n_n4571) & (n_n4523) & (n_n4557) & (!n_n4560) & (!n_n4553)) + ((!n_n4571) & (n_n4523) & (n_n4557) & (!n_n4560) & (n_n4553)) + ((!n_n4571) & (n_n4523) & (n_n4557) & (n_n4560) & (!n_n4553)) + ((!n_n4571) & (n_n4523) & (n_n4557) & (n_n4560) & (n_n4553)) + ((n_n4571) & (!n_n4523) & (!n_n4557) & (!n_n4560) & (!n_n4553)) + ((n_n4571) & (!n_n4523) & (!n_n4557) & (!n_n4560) & (n_n4553)) + ((n_n4571) & (!n_n4523) & (!n_n4557) & (n_n4560) & (!n_n4553)) + ((n_n4571) & (!n_n4523) & (!n_n4557) & (n_n4560) & (n_n4553)) + ((n_n4571) & (!n_n4523) & (n_n4557) & (!n_n4560) & (!n_n4553)) + ((n_n4571) & (!n_n4523) & (n_n4557) & (!n_n4560) & (n_n4553)) + ((n_n4571) & (!n_n4523) & (n_n4557) & (n_n4560) & (!n_n4553)) + ((n_n4571) & (!n_n4523) & (n_n4557) & (n_n4560) & (n_n4553)) + ((n_n4571) & (n_n4523) & (!n_n4557) & (!n_n4560) & (!n_n4553)) + ((n_n4571) & (n_n4523) & (!n_n4557) & (!n_n4560) & (n_n4553)) + ((n_n4571) & (n_n4523) & (!n_n4557) & (n_n4560) & (!n_n4553)) + ((n_n4571) & (n_n4523) & (!n_n4557) & (n_n4560) & (n_n4553)) + ((n_n4571) & (n_n4523) & (n_n4557) & (!n_n4560) & (!n_n4553)) + ((n_n4571) & (n_n4523) & (n_n4557) & (!n_n4560) & (n_n4553)) + ((n_n4571) & (n_n4523) & (n_n4557) & (n_n4560) & (!n_n4553)) + ((n_n4571) & (n_n4523) & (n_n4557) & (n_n4560) & (n_n4553)));
	assign n_n2087 = (((!n_n2102) & (!x16487x) & (!x16488x) & (!x16494x) & (x16495x)) + ((!n_n2102) & (!x16487x) & (!x16488x) & (x16494x) & (!x16495x)) + ((!n_n2102) & (!x16487x) & (!x16488x) & (x16494x) & (x16495x)) + ((!n_n2102) & (!x16487x) & (x16488x) & (!x16494x) & (!x16495x)) + ((!n_n2102) & (!x16487x) & (x16488x) & (!x16494x) & (x16495x)) + ((!n_n2102) & (!x16487x) & (x16488x) & (x16494x) & (!x16495x)) + ((!n_n2102) & (!x16487x) & (x16488x) & (x16494x) & (x16495x)) + ((!n_n2102) & (x16487x) & (!x16488x) & (!x16494x) & (!x16495x)) + ((!n_n2102) & (x16487x) & (!x16488x) & (!x16494x) & (x16495x)) + ((!n_n2102) & (x16487x) & (!x16488x) & (x16494x) & (!x16495x)) + ((!n_n2102) & (x16487x) & (!x16488x) & (x16494x) & (x16495x)) + ((!n_n2102) & (x16487x) & (x16488x) & (!x16494x) & (!x16495x)) + ((!n_n2102) & (x16487x) & (x16488x) & (!x16494x) & (x16495x)) + ((!n_n2102) & (x16487x) & (x16488x) & (x16494x) & (!x16495x)) + ((!n_n2102) & (x16487x) & (x16488x) & (x16494x) & (x16495x)) + ((n_n2102) & (!x16487x) & (!x16488x) & (!x16494x) & (!x16495x)) + ((n_n2102) & (!x16487x) & (!x16488x) & (!x16494x) & (x16495x)) + ((n_n2102) & (!x16487x) & (!x16488x) & (x16494x) & (!x16495x)) + ((n_n2102) & (!x16487x) & (!x16488x) & (x16494x) & (x16495x)) + ((n_n2102) & (!x16487x) & (x16488x) & (!x16494x) & (!x16495x)) + ((n_n2102) & (!x16487x) & (x16488x) & (!x16494x) & (x16495x)) + ((n_n2102) & (!x16487x) & (x16488x) & (x16494x) & (!x16495x)) + ((n_n2102) & (!x16487x) & (x16488x) & (x16494x) & (x16495x)) + ((n_n2102) & (x16487x) & (!x16488x) & (!x16494x) & (!x16495x)) + ((n_n2102) & (x16487x) & (!x16488x) & (!x16494x) & (x16495x)) + ((n_n2102) & (x16487x) & (!x16488x) & (x16494x) & (!x16495x)) + ((n_n2102) & (x16487x) & (!x16488x) & (x16494x) & (x16495x)) + ((n_n2102) & (x16487x) & (x16488x) & (!x16494x) & (!x16495x)) + ((n_n2102) & (x16487x) & (x16488x) & (!x16494x) & (x16495x)) + ((n_n2102) & (x16487x) & (x16488x) & (x16494x) & (!x16495x)) + ((n_n2102) & (x16487x) & (x16488x) & (x16494x) & (x16495x)));
	assign x24x = (((!i_9_) & (i_7_) & (!i_8_) & (i_6_)));
	assign x530x = (((!i_1_) & (!i_2_) & (i_0_) & (n_n464)));
	assign n_n2130 = (((!n_n482) & (!n_n532) & (!x14x) & (!n_n530) & (n_n4777)) + ((!n_n482) & (!n_n532) & (!x14x) & (n_n530) & (n_n4777)) + ((!n_n482) & (!n_n532) & (x14x) & (!n_n530) & (n_n4777)) + ((!n_n482) & (!n_n532) & (x14x) & (n_n530) & (n_n4777)) + ((!n_n482) & (n_n532) & (!x14x) & (!n_n530) & (n_n4777)) + ((!n_n482) & (n_n532) & (!x14x) & (n_n530) & (n_n4777)) + ((!n_n482) & (n_n532) & (x14x) & (!n_n530) & (n_n4777)) + ((!n_n482) & (n_n532) & (x14x) & (n_n530) & (n_n4777)) + ((n_n482) & (!n_n532) & (!x14x) & (!n_n530) & (n_n4777)) + ((n_n482) & (!n_n532) & (!x14x) & (n_n530) & (n_n4777)) + ((n_n482) & (!n_n532) & (x14x) & (!n_n530) & (n_n4777)) + ((n_n482) & (!n_n532) & (x14x) & (n_n530) & (!n_n4777)) + ((n_n482) & (!n_n532) & (x14x) & (n_n530) & (n_n4777)) + ((n_n482) & (n_n532) & (!x14x) & (!n_n530) & (n_n4777)) + ((n_n482) & (n_n532) & (!x14x) & (n_n530) & (n_n4777)) + ((n_n482) & (n_n532) & (x14x) & (!n_n530) & (!n_n4777)) + ((n_n482) & (n_n532) & (x14x) & (!n_n530) & (n_n4777)) + ((n_n482) & (n_n532) & (x14x) & (n_n530) & (!n_n4777)) + ((n_n482) & (n_n532) & (x14x) & (n_n530) & (n_n4777)));
	assign n_n4781 = (((!i_9_) & (n_n482) & (n_n325) & (n_n530)));
	assign x16514x = (((!n_n4800) & (!n_n4803) & (!n_n4783) & (n_n4812)) + ((!n_n4800) & (!n_n4803) & (n_n4783) & (!n_n4812)) + ((!n_n4800) & (!n_n4803) & (n_n4783) & (n_n4812)) + ((!n_n4800) & (n_n4803) & (!n_n4783) & (!n_n4812)) + ((!n_n4800) & (n_n4803) & (!n_n4783) & (n_n4812)) + ((!n_n4800) & (n_n4803) & (n_n4783) & (!n_n4812)) + ((!n_n4800) & (n_n4803) & (n_n4783) & (n_n4812)) + ((n_n4800) & (!n_n4803) & (!n_n4783) & (!n_n4812)) + ((n_n4800) & (!n_n4803) & (!n_n4783) & (n_n4812)) + ((n_n4800) & (!n_n4803) & (n_n4783) & (!n_n4812)) + ((n_n4800) & (!n_n4803) & (n_n4783) & (n_n4812)) + ((n_n4800) & (n_n4803) & (!n_n4783) & (!n_n4812)) + ((n_n4800) & (n_n4803) & (!n_n4783) & (n_n4812)) + ((n_n4800) & (n_n4803) & (n_n4783) & (!n_n4812)) + ((n_n4800) & (n_n4803) & (n_n4783) & (n_n4812)));
	assign x16516x = (((!x24x) & (!x530x) & (!n_n2130) & (!n_n4781) & (x16514x)) + ((!x24x) & (!x530x) & (!n_n2130) & (n_n4781) & (!x16514x)) + ((!x24x) & (!x530x) & (!n_n2130) & (n_n4781) & (x16514x)) + ((!x24x) & (!x530x) & (n_n2130) & (!n_n4781) & (!x16514x)) + ((!x24x) & (!x530x) & (n_n2130) & (!n_n4781) & (x16514x)) + ((!x24x) & (!x530x) & (n_n2130) & (n_n4781) & (!x16514x)) + ((!x24x) & (!x530x) & (n_n2130) & (n_n4781) & (x16514x)) + ((!x24x) & (x530x) & (!n_n2130) & (!n_n4781) & (x16514x)) + ((!x24x) & (x530x) & (!n_n2130) & (n_n4781) & (!x16514x)) + ((!x24x) & (x530x) & (!n_n2130) & (n_n4781) & (x16514x)) + ((!x24x) & (x530x) & (n_n2130) & (!n_n4781) & (!x16514x)) + ((!x24x) & (x530x) & (n_n2130) & (!n_n4781) & (x16514x)) + ((!x24x) & (x530x) & (n_n2130) & (n_n4781) & (!x16514x)) + ((!x24x) & (x530x) & (n_n2130) & (n_n4781) & (x16514x)) + ((x24x) & (!x530x) & (!n_n2130) & (!n_n4781) & (x16514x)) + ((x24x) & (!x530x) & (!n_n2130) & (n_n4781) & (!x16514x)) + ((x24x) & (!x530x) & (!n_n2130) & (n_n4781) & (x16514x)) + ((x24x) & (!x530x) & (n_n2130) & (!n_n4781) & (!x16514x)) + ((x24x) & (!x530x) & (n_n2130) & (!n_n4781) & (x16514x)) + ((x24x) & (!x530x) & (n_n2130) & (n_n4781) & (!x16514x)) + ((x24x) & (!x530x) & (n_n2130) & (n_n4781) & (x16514x)) + ((x24x) & (x530x) & (!n_n2130) & (!n_n4781) & (!x16514x)) + ((x24x) & (x530x) & (!n_n2130) & (!n_n4781) & (x16514x)) + ((x24x) & (x530x) & (!n_n2130) & (n_n4781) & (!x16514x)) + ((x24x) & (x530x) & (!n_n2130) & (n_n4781) & (x16514x)) + ((x24x) & (x530x) & (n_n2130) & (!n_n4781) & (!x16514x)) + ((x24x) & (x530x) & (n_n2130) & (!n_n4781) & (x16514x)) + ((x24x) & (x530x) & (n_n2130) & (n_n4781) & (!x16514x)) + ((x24x) & (x530x) & (n_n2130) & (n_n4781) & (x16514x)));
	assign x16503x = (((!n_n4740) & (!n_n4710) & (!n_n4719) & (n_n4708)) + ((!n_n4740) & (!n_n4710) & (n_n4719) & (!n_n4708)) + ((!n_n4740) & (!n_n4710) & (n_n4719) & (n_n4708)) + ((!n_n4740) & (n_n4710) & (!n_n4719) & (!n_n4708)) + ((!n_n4740) & (n_n4710) & (!n_n4719) & (n_n4708)) + ((!n_n4740) & (n_n4710) & (n_n4719) & (!n_n4708)) + ((!n_n4740) & (n_n4710) & (n_n4719) & (n_n4708)) + ((n_n4740) & (!n_n4710) & (!n_n4719) & (!n_n4708)) + ((n_n4740) & (!n_n4710) & (!n_n4719) & (n_n4708)) + ((n_n4740) & (!n_n4710) & (n_n4719) & (!n_n4708)) + ((n_n4740) & (!n_n4710) & (n_n4719) & (n_n4708)) + ((n_n4740) & (n_n4710) & (!n_n4719) & (!n_n4708)) + ((n_n4740) & (n_n4710) & (!n_n4719) & (n_n4708)) + ((n_n4740) & (n_n4710) & (n_n4719) & (!n_n4708)) + ((n_n4740) & (n_n4710) & (n_n4719) & (n_n4708)));
	assign x16504x = (((!n_n4764) & (!n_n4772) & (!n_n4706) & (!n_n4699) & (n_n4687)) + ((!n_n4764) & (!n_n4772) & (!n_n4706) & (n_n4699) & (!n_n4687)) + ((!n_n4764) & (!n_n4772) & (!n_n4706) & (n_n4699) & (n_n4687)) + ((!n_n4764) & (!n_n4772) & (n_n4706) & (!n_n4699) & (!n_n4687)) + ((!n_n4764) & (!n_n4772) & (n_n4706) & (!n_n4699) & (n_n4687)) + ((!n_n4764) & (!n_n4772) & (n_n4706) & (n_n4699) & (!n_n4687)) + ((!n_n4764) & (!n_n4772) & (n_n4706) & (n_n4699) & (n_n4687)) + ((!n_n4764) & (n_n4772) & (!n_n4706) & (!n_n4699) & (!n_n4687)) + ((!n_n4764) & (n_n4772) & (!n_n4706) & (!n_n4699) & (n_n4687)) + ((!n_n4764) & (n_n4772) & (!n_n4706) & (n_n4699) & (!n_n4687)) + ((!n_n4764) & (n_n4772) & (!n_n4706) & (n_n4699) & (n_n4687)) + ((!n_n4764) & (n_n4772) & (n_n4706) & (!n_n4699) & (!n_n4687)) + ((!n_n4764) & (n_n4772) & (n_n4706) & (!n_n4699) & (n_n4687)) + ((!n_n4764) & (n_n4772) & (n_n4706) & (n_n4699) & (!n_n4687)) + ((!n_n4764) & (n_n4772) & (n_n4706) & (n_n4699) & (n_n4687)) + ((n_n4764) & (!n_n4772) & (!n_n4706) & (!n_n4699) & (!n_n4687)) + ((n_n4764) & (!n_n4772) & (!n_n4706) & (!n_n4699) & (n_n4687)) + ((n_n4764) & (!n_n4772) & (!n_n4706) & (n_n4699) & (!n_n4687)) + ((n_n4764) & (!n_n4772) & (!n_n4706) & (n_n4699) & (n_n4687)) + ((n_n4764) & (!n_n4772) & (n_n4706) & (!n_n4699) & (!n_n4687)) + ((n_n4764) & (!n_n4772) & (n_n4706) & (!n_n4699) & (n_n4687)) + ((n_n4764) & (!n_n4772) & (n_n4706) & (n_n4699) & (!n_n4687)) + ((n_n4764) & (!n_n4772) & (n_n4706) & (n_n4699) & (n_n4687)) + ((n_n4764) & (n_n4772) & (!n_n4706) & (!n_n4699) & (!n_n4687)) + ((n_n4764) & (n_n4772) & (!n_n4706) & (!n_n4699) & (n_n4687)) + ((n_n4764) & (n_n4772) & (!n_n4706) & (n_n4699) & (!n_n4687)) + ((n_n4764) & (n_n4772) & (!n_n4706) & (n_n4699) & (n_n4687)) + ((n_n4764) & (n_n4772) & (n_n4706) & (!n_n4699) & (!n_n4687)) + ((n_n4764) & (n_n4772) & (n_n4706) & (!n_n4699) & (n_n4687)) + ((n_n4764) & (n_n4772) & (n_n4706) & (n_n4699) & (!n_n4687)) + ((n_n4764) & (n_n4772) & (n_n4706) & (n_n4699) & (n_n4687)));
	assign x16509x = (((!n_n4647) & (!n_n4656) & (!n_n4659) & (n_n4675)) + ((!n_n4647) & (!n_n4656) & (n_n4659) & (!n_n4675)) + ((!n_n4647) & (!n_n4656) & (n_n4659) & (n_n4675)) + ((!n_n4647) & (n_n4656) & (!n_n4659) & (!n_n4675)) + ((!n_n4647) & (n_n4656) & (!n_n4659) & (n_n4675)) + ((!n_n4647) & (n_n4656) & (n_n4659) & (!n_n4675)) + ((!n_n4647) & (n_n4656) & (n_n4659) & (n_n4675)) + ((n_n4647) & (!n_n4656) & (!n_n4659) & (!n_n4675)) + ((n_n4647) & (!n_n4656) & (!n_n4659) & (n_n4675)) + ((n_n4647) & (!n_n4656) & (n_n4659) & (!n_n4675)) + ((n_n4647) & (!n_n4656) & (n_n4659) & (n_n4675)) + ((n_n4647) & (n_n4656) & (!n_n4659) & (!n_n4675)) + ((n_n4647) & (n_n4656) & (!n_n4659) & (n_n4675)) + ((n_n4647) & (n_n4656) & (n_n4659) & (!n_n4675)) + ((n_n4647) & (n_n4656) & (n_n4659) & (n_n4675)));
	assign x16510x = (((!n_n4674) & (!n_n4661) & (!n_n4671) & (!n_n4672) & (n_n4685)) + ((!n_n4674) & (!n_n4661) & (!n_n4671) & (n_n4672) & (!n_n4685)) + ((!n_n4674) & (!n_n4661) & (!n_n4671) & (n_n4672) & (n_n4685)) + ((!n_n4674) & (!n_n4661) & (n_n4671) & (!n_n4672) & (!n_n4685)) + ((!n_n4674) & (!n_n4661) & (n_n4671) & (!n_n4672) & (n_n4685)) + ((!n_n4674) & (!n_n4661) & (n_n4671) & (n_n4672) & (!n_n4685)) + ((!n_n4674) & (!n_n4661) & (n_n4671) & (n_n4672) & (n_n4685)) + ((!n_n4674) & (n_n4661) & (!n_n4671) & (!n_n4672) & (!n_n4685)) + ((!n_n4674) & (n_n4661) & (!n_n4671) & (!n_n4672) & (n_n4685)) + ((!n_n4674) & (n_n4661) & (!n_n4671) & (n_n4672) & (!n_n4685)) + ((!n_n4674) & (n_n4661) & (!n_n4671) & (n_n4672) & (n_n4685)) + ((!n_n4674) & (n_n4661) & (n_n4671) & (!n_n4672) & (!n_n4685)) + ((!n_n4674) & (n_n4661) & (n_n4671) & (!n_n4672) & (n_n4685)) + ((!n_n4674) & (n_n4661) & (n_n4671) & (n_n4672) & (!n_n4685)) + ((!n_n4674) & (n_n4661) & (n_n4671) & (n_n4672) & (n_n4685)) + ((n_n4674) & (!n_n4661) & (!n_n4671) & (!n_n4672) & (!n_n4685)) + ((n_n4674) & (!n_n4661) & (!n_n4671) & (!n_n4672) & (n_n4685)) + ((n_n4674) & (!n_n4661) & (!n_n4671) & (n_n4672) & (!n_n4685)) + ((n_n4674) & (!n_n4661) & (!n_n4671) & (n_n4672) & (n_n4685)) + ((n_n4674) & (!n_n4661) & (n_n4671) & (!n_n4672) & (!n_n4685)) + ((n_n4674) & (!n_n4661) & (n_n4671) & (!n_n4672) & (n_n4685)) + ((n_n4674) & (!n_n4661) & (n_n4671) & (n_n4672) & (!n_n4685)) + ((n_n4674) & (!n_n4661) & (n_n4671) & (n_n4672) & (n_n4685)) + ((n_n4674) & (n_n4661) & (!n_n4671) & (!n_n4672) & (!n_n4685)) + ((n_n4674) & (n_n4661) & (!n_n4671) & (!n_n4672) & (n_n4685)) + ((n_n4674) & (n_n4661) & (!n_n4671) & (n_n4672) & (!n_n4685)) + ((n_n4674) & (n_n4661) & (!n_n4671) & (n_n4672) & (n_n4685)) + ((n_n4674) & (n_n4661) & (n_n4671) & (!n_n4672) & (!n_n4685)) + ((n_n4674) & (n_n4661) & (n_n4671) & (!n_n4672) & (n_n4685)) + ((n_n4674) & (n_n4661) & (n_n4671) & (n_n4672) & (!n_n4685)) + ((n_n4674) & (n_n4661) & (n_n4671) & (n_n4672) & (n_n4685)));
	assign x16517x = (((!x16503x) & (!x16504x) & (!x16509x) & (x16510x)) + ((!x16503x) & (!x16504x) & (x16509x) & (!x16510x)) + ((!x16503x) & (!x16504x) & (x16509x) & (x16510x)) + ((!x16503x) & (x16504x) & (!x16509x) & (!x16510x)) + ((!x16503x) & (x16504x) & (!x16509x) & (x16510x)) + ((!x16503x) & (x16504x) & (x16509x) & (!x16510x)) + ((!x16503x) & (x16504x) & (x16509x) & (x16510x)) + ((x16503x) & (!x16504x) & (!x16509x) & (!x16510x)) + ((x16503x) & (!x16504x) & (!x16509x) & (x16510x)) + ((x16503x) & (!x16504x) & (x16509x) & (!x16510x)) + ((x16503x) & (!x16504x) & (x16509x) & (x16510x)) + ((x16503x) & (x16504x) & (!x16509x) & (!x16510x)) + ((x16503x) & (x16504x) & (!x16509x) & (x16510x)) + ((x16503x) & (x16504x) & (x16509x) & (!x16510x)) + ((x16503x) & (x16504x) & (x16509x) & (x16510x)));
	assign n_n2267 = (((!n_n4363) & (!n_n4359) & (!n_n4275) & (!x74x) & (x345x)) + ((!n_n4363) & (!n_n4359) & (!n_n4275) & (x74x) & (!x345x)) + ((!n_n4363) & (!n_n4359) & (!n_n4275) & (x74x) & (x345x)) + ((!n_n4363) & (!n_n4359) & (n_n4275) & (!x74x) & (!x345x)) + ((!n_n4363) & (!n_n4359) & (n_n4275) & (!x74x) & (x345x)) + ((!n_n4363) & (!n_n4359) & (n_n4275) & (x74x) & (!x345x)) + ((!n_n4363) & (!n_n4359) & (n_n4275) & (x74x) & (x345x)) + ((!n_n4363) & (n_n4359) & (!n_n4275) & (!x74x) & (!x345x)) + ((!n_n4363) & (n_n4359) & (!n_n4275) & (!x74x) & (x345x)) + ((!n_n4363) & (n_n4359) & (!n_n4275) & (x74x) & (!x345x)) + ((!n_n4363) & (n_n4359) & (!n_n4275) & (x74x) & (x345x)) + ((!n_n4363) & (n_n4359) & (n_n4275) & (!x74x) & (!x345x)) + ((!n_n4363) & (n_n4359) & (n_n4275) & (!x74x) & (x345x)) + ((!n_n4363) & (n_n4359) & (n_n4275) & (x74x) & (!x345x)) + ((!n_n4363) & (n_n4359) & (n_n4275) & (x74x) & (x345x)) + ((n_n4363) & (!n_n4359) & (!n_n4275) & (!x74x) & (!x345x)) + ((n_n4363) & (!n_n4359) & (!n_n4275) & (!x74x) & (x345x)) + ((n_n4363) & (!n_n4359) & (!n_n4275) & (x74x) & (!x345x)) + ((n_n4363) & (!n_n4359) & (!n_n4275) & (x74x) & (x345x)) + ((n_n4363) & (!n_n4359) & (n_n4275) & (!x74x) & (!x345x)) + ((n_n4363) & (!n_n4359) & (n_n4275) & (!x74x) & (x345x)) + ((n_n4363) & (!n_n4359) & (n_n4275) & (x74x) & (!x345x)) + ((n_n4363) & (!n_n4359) & (n_n4275) & (x74x) & (x345x)) + ((n_n4363) & (n_n4359) & (!n_n4275) & (!x74x) & (!x345x)) + ((n_n4363) & (n_n4359) & (!n_n4275) & (!x74x) & (x345x)) + ((n_n4363) & (n_n4359) & (!n_n4275) & (x74x) & (!x345x)) + ((n_n4363) & (n_n4359) & (!n_n4275) & (x74x) & (x345x)) + ((n_n4363) & (n_n4359) & (n_n4275) & (!x74x) & (!x345x)) + ((n_n4363) & (n_n4359) & (n_n4275) & (!x74x) & (x345x)) + ((n_n4363) & (n_n4359) & (n_n4275) & (x74x) & (!x345x)) + ((n_n4363) & (n_n4359) & (n_n4275) & (x74x) & (x345x)));
	assign x16554x = (((!n_n4382) & (!n_n4379) & (!n_n4373) & (!x300x) & (x423x)) + ((!n_n4382) & (!n_n4379) & (!n_n4373) & (x300x) & (!x423x)) + ((!n_n4382) & (!n_n4379) & (!n_n4373) & (x300x) & (x423x)) + ((!n_n4382) & (!n_n4379) & (n_n4373) & (!x300x) & (!x423x)) + ((!n_n4382) & (!n_n4379) & (n_n4373) & (!x300x) & (x423x)) + ((!n_n4382) & (!n_n4379) & (n_n4373) & (x300x) & (!x423x)) + ((!n_n4382) & (!n_n4379) & (n_n4373) & (x300x) & (x423x)) + ((!n_n4382) & (n_n4379) & (!n_n4373) & (!x300x) & (!x423x)) + ((!n_n4382) & (n_n4379) & (!n_n4373) & (!x300x) & (x423x)) + ((!n_n4382) & (n_n4379) & (!n_n4373) & (x300x) & (!x423x)) + ((!n_n4382) & (n_n4379) & (!n_n4373) & (x300x) & (x423x)) + ((!n_n4382) & (n_n4379) & (n_n4373) & (!x300x) & (!x423x)) + ((!n_n4382) & (n_n4379) & (n_n4373) & (!x300x) & (x423x)) + ((!n_n4382) & (n_n4379) & (n_n4373) & (x300x) & (!x423x)) + ((!n_n4382) & (n_n4379) & (n_n4373) & (x300x) & (x423x)) + ((n_n4382) & (!n_n4379) & (!n_n4373) & (!x300x) & (!x423x)) + ((n_n4382) & (!n_n4379) & (!n_n4373) & (!x300x) & (x423x)) + ((n_n4382) & (!n_n4379) & (!n_n4373) & (x300x) & (!x423x)) + ((n_n4382) & (!n_n4379) & (!n_n4373) & (x300x) & (x423x)) + ((n_n4382) & (!n_n4379) & (n_n4373) & (!x300x) & (!x423x)) + ((n_n4382) & (!n_n4379) & (n_n4373) & (!x300x) & (x423x)) + ((n_n4382) & (!n_n4379) & (n_n4373) & (x300x) & (!x423x)) + ((n_n4382) & (!n_n4379) & (n_n4373) & (x300x) & (x423x)) + ((n_n4382) & (n_n4379) & (!n_n4373) & (!x300x) & (!x423x)) + ((n_n4382) & (n_n4379) & (!n_n4373) & (!x300x) & (x423x)) + ((n_n4382) & (n_n4379) & (!n_n4373) & (x300x) & (!x423x)) + ((n_n4382) & (n_n4379) & (!n_n4373) & (x300x) & (x423x)) + ((n_n4382) & (n_n4379) & (n_n4373) & (!x300x) & (!x423x)) + ((n_n4382) & (n_n4379) & (n_n4373) & (!x300x) & (x423x)) + ((n_n4382) & (n_n4379) & (n_n4373) & (x300x) & (!x423x)) + ((n_n4382) & (n_n4379) & (n_n4373) & (x300x) & (x423x)));
	assign x16555x = (((!n_n4386) & (!n_n2435) & (!x14460x) & (!x282x) & (x12447x)) + ((!n_n4386) & (!n_n2435) & (!x14460x) & (x282x) & (!x12447x)) + ((!n_n4386) & (!n_n2435) & (!x14460x) & (x282x) & (x12447x)) + ((!n_n4386) & (!n_n2435) & (x14460x) & (!x282x) & (!x12447x)) + ((!n_n4386) & (!n_n2435) & (x14460x) & (!x282x) & (x12447x)) + ((!n_n4386) & (!n_n2435) & (x14460x) & (x282x) & (!x12447x)) + ((!n_n4386) & (!n_n2435) & (x14460x) & (x282x) & (x12447x)) + ((!n_n4386) & (n_n2435) & (!x14460x) & (!x282x) & (!x12447x)) + ((!n_n4386) & (n_n2435) & (!x14460x) & (!x282x) & (x12447x)) + ((!n_n4386) & (n_n2435) & (!x14460x) & (x282x) & (!x12447x)) + ((!n_n4386) & (n_n2435) & (!x14460x) & (x282x) & (x12447x)) + ((!n_n4386) & (n_n2435) & (x14460x) & (!x282x) & (!x12447x)) + ((!n_n4386) & (n_n2435) & (x14460x) & (!x282x) & (x12447x)) + ((!n_n4386) & (n_n2435) & (x14460x) & (x282x) & (!x12447x)) + ((!n_n4386) & (n_n2435) & (x14460x) & (x282x) & (x12447x)) + ((n_n4386) & (!n_n2435) & (!x14460x) & (!x282x) & (!x12447x)) + ((n_n4386) & (!n_n2435) & (!x14460x) & (!x282x) & (x12447x)) + ((n_n4386) & (!n_n2435) & (!x14460x) & (x282x) & (!x12447x)) + ((n_n4386) & (!n_n2435) & (!x14460x) & (x282x) & (x12447x)) + ((n_n4386) & (!n_n2435) & (x14460x) & (!x282x) & (!x12447x)) + ((n_n4386) & (!n_n2435) & (x14460x) & (!x282x) & (x12447x)) + ((n_n4386) & (!n_n2435) & (x14460x) & (x282x) & (!x12447x)) + ((n_n4386) & (!n_n2435) & (x14460x) & (x282x) & (x12447x)) + ((n_n4386) & (n_n2435) & (!x14460x) & (!x282x) & (!x12447x)) + ((n_n4386) & (n_n2435) & (!x14460x) & (!x282x) & (x12447x)) + ((n_n4386) & (n_n2435) & (!x14460x) & (x282x) & (!x12447x)) + ((n_n4386) & (n_n2435) & (!x14460x) & (x282x) & (x12447x)) + ((n_n4386) & (n_n2435) & (x14460x) & (!x282x) & (!x12447x)) + ((n_n4386) & (n_n2435) & (x14460x) & (!x282x) & (x12447x)) + ((n_n4386) & (n_n2435) & (x14460x) & (x282x) & (!x12447x)) + ((n_n4386) & (n_n2435) & (x14460x) & (x282x) & (x12447x)));
	assign x16557x = (((!n_n2267) & (!x16554x) & (x16555x)) + ((!n_n2267) & (x16554x) & (!x16555x)) + ((!n_n2267) & (x16554x) & (x16555x)) + ((n_n2267) & (!x16554x) & (!x16555x)) + ((n_n2267) & (!x16554x) & (x16555x)) + ((n_n2267) & (x16554x) & (!x16555x)) + ((n_n2267) & (x16554x) & (x16555x)));
	assign n_n2190 = (((!n_n2263) & (!x16526x) & (!x16527x) & (x16533x)) + ((!n_n2263) & (!x16526x) & (x16527x) & (!x16533x)) + ((!n_n2263) & (!x16526x) & (x16527x) & (x16533x)) + ((!n_n2263) & (x16526x) & (!x16527x) & (!x16533x)) + ((!n_n2263) & (x16526x) & (!x16527x) & (x16533x)) + ((!n_n2263) & (x16526x) & (x16527x) & (!x16533x)) + ((!n_n2263) & (x16526x) & (x16527x) & (x16533x)) + ((n_n2263) & (!x16526x) & (!x16527x) & (!x16533x)) + ((n_n2263) & (!x16526x) & (!x16527x) & (x16533x)) + ((n_n2263) & (!x16526x) & (x16527x) & (!x16533x)) + ((n_n2263) & (!x16526x) & (x16527x) & (x16533x)) + ((n_n2263) & (x16526x) & (!x16527x) & (!x16533x)) + ((n_n2263) & (x16526x) & (!x16527x) & (x16533x)) + ((n_n2263) & (x16526x) & (x16527x) & (!x16533x)) + ((n_n2263) & (x16526x) & (x16527x) & (x16533x)));
	assign n_n2268 = (((!n_n4343) & (!n_n4352) & (!x399x) & (!x22197x)) + ((!n_n4343) & (!n_n4352) & (x399x) & (!x22197x)) + ((!n_n4343) & (!n_n4352) & (x399x) & (x22197x)) + ((!n_n4343) & (n_n4352) & (!x399x) & (!x22197x)) + ((!n_n4343) & (n_n4352) & (!x399x) & (x22197x)) + ((!n_n4343) & (n_n4352) & (x399x) & (!x22197x)) + ((!n_n4343) & (n_n4352) & (x399x) & (x22197x)) + ((n_n4343) & (!n_n4352) & (!x399x) & (!x22197x)) + ((n_n4343) & (!n_n4352) & (!x399x) & (x22197x)) + ((n_n4343) & (!n_n4352) & (x399x) & (!x22197x)) + ((n_n4343) & (!n_n4352) & (x399x) & (x22197x)) + ((n_n4343) & (n_n4352) & (!x399x) & (!x22197x)) + ((n_n4343) & (n_n4352) & (!x399x) & (x22197x)) + ((n_n4343) & (n_n4352) & (x399x) & (!x22197x)) + ((n_n4343) & (n_n4352) & (x399x) & (x22197x)));
	assign x16545x = (((!n_n4317) & (!n_n4312) & (!n_n2446) & (!n_n2443) & (n_n2445)) + ((!n_n4317) & (!n_n4312) & (!n_n2446) & (n_n2443) & (!n_n2445)) + ((!n_n4317) & (!n_n4312) & (!n_n2446) & (n_n2443) & (n_n2445)) + ((!n_n4317) & (!n_n4312) & (n_n2446) & (!n_n2443) & (!n_n2445)) + ((!n_n4317) & (!n_n4312) & (n_n2446) & (!n_n2443) & (n_n2445)) + ((!n_n4317) & (!n_n4312) & (n_n2446) & (n_n2443) & (!n_n2445)) + ((!n_n4317) & (!n_n4312) & (n_n2446) & (n_n2443) & (n_n2445)) + ((!n_n4317) & (n_n4312) & (!n_n2446) & (!n_n2443) & (!n_n2445)) + ((!n_n4317) & (n_n4312) & (!n_n2446) & (!n_n2443) & (n_n2445)) + ((!n_n4317) & (n_n4312) & (!n_n2446) & (n_n2443) & (!n_n2445)) + ((!n_n4317) & (n_n4312) & (!n_n2446) & (n_n2443) & (n_n2445)) + ((!n_n4317) & (n_n4312) & (n_n2446) & (!n_n2443) & (!n_n2445)) + ((!n_n4317) & (n_n4312) & (n_n2446) & (!n_n2443) & (n_n2445)) + ((!n_n4317) & (n_n4312) & (n_n2446) & (n_n2443) & (!n_n2445)) + ((!n_n4317) & (n_n4312) & (n_n2446) & (n_n2443) & (n_n2445)) + ((n_n4317) & (!n_n4312) & (!n_n2446) & (!n_n2443) & (!n_n2445)) + ((n_n4317) & (!n_n4312) & (!n_n2446) & (!n_n2443) & (n_n2445)) + ((n_n4317) & (!n_n4312) & (!n_n2446) & (n_n2443) & (!n_n2445)) + ((n_n4317) & (!n_n4312) & (!n_n2446) & (n_n2443) & (n_n2445)) + ((n_n4317) & (!n_n4312) & (n_n2446) & (!n_n2443) & (!n_n2445)) + ((n_n4317) & (!n_n4312) & (n_n2446) & (!n_n2443) & (n_n2445)) + ((n_n4317) & (!n_n4312) & (n_n2446) & (n_n2443) & (!n_n2445)) + ((n_n4317) & (!n_n4312) & (n_n2446) & (n_n2443) & (n_n2445)) + ((n_n4317) & (n_n4312) & (!n_n2446) & (!n_n2443) & (!n_n2445)) + ((n_n4317) & (n_n4312) & (!n_n2446) & (!n_n2443) & (n_n2445)) + ((n_n4317) & (n_n4312) & (!n_n2446) & (n_n2443) & (!n_n2445)) + ((n_n4317) & (n_n4312) & (!n_n2446) & (n_n2443) & (n_n2445)) + ((n_n4317) & (n_n4312) & (n_n2446) & (!n_n2443) & (!n_n2445)) + ((n_n4317) & (n_n4312) & (n_n2446) & (!n_n2443) & (n_n2445)) + ((n_n4317) & (n_n4312) & (n_n2446) & (n_n2443) & (!n_n2445)) + ((n_n4317) & (n_n4312) & (n_n2446) & (n_n2443) & (n_n2445)));
	assign x16544x = (((!n_n4319) & (!n_n4336) & (!n_n4321) & (!x198x) & (x283x)) + ((!n_n4319) & (!n_n4336) & (!n_n4321) & (x198x) & (!x283x)) + ((!n_n4319) & (!n_n4336) & (!n_n4321) & (x198x) & (x283x)) + ((!n_n4319) & (!n_n4336) & (n_n4321) & (!x198x) & (!x283x)) + ((!n_n4319) & (!n_n4336) & (n_n4321) & (!x198x) & (x283x)) + ((!n_n4319) & (!n_n4336) & (n_n4321) & (x198x) & (!x283x)) + ((!n_n4319) & (!n_n4336) & (n_n4321) & (x198x) & (x283x)) + ((!n_n4319) & (n_n4336) & (!n_n4321) & (!x198x) & (!x283x)) + ((!n_n4319) & (n_n4336) & (!n_n4321) & (!x198x) & (x283x)) + ((!n_n4319) & (n_n4336) & (!n_n4321) & (x198x) & (!x283x)) + ((!n_n4319) & (n_n4336) & (!n_n4321) & (x198x) & (x283x)) + ((!n_n4319) & (n_n4336) & (n_n4321) & (!x198x) & (!x283x)) + ((!n_n4319) & (n_n4336) & (n_n4321) & (!x198x) & (x283x)) + ((!n_n4319) & (n_n4336) & (n_n4321) & (x198x) & (!x283x)) + ((!n_n4319) & (n_n4336) & (n_n4321) & (x198x) & (x283x)) + ((n_n4319) & (!n_n4336) & (!n_n4321) & (!x198x) & (!x283x)) + ((n_n4319) & (!n_n4336) & (!n_n4321) & (!x198x) & (x283x)) + ((n_n4319) & (!n_n4336) & (!n_n4321) & (x198x) & (!x283x)) + ((n_n4319) & (!n_n4336) & (!n_n4321) & (x198x) & (x283x)) + ((n_n4319) & (!n_n4336) & (n_n4321) & (!x198x) & (!x283x)) + ((n_n4319) & (!n_n4336) & (n_n4321) & (!x198x) & (x283x)) + ((n_n4319) & (!n_n4336) & (n_n4321) & (x198x) & (!x283x)) + ((n_n4319) & (!n_n4336) & (n_n4321) & (x198x) & (x283x)) + ((n_n4319) & (n_n4336) & (!n_n4321) & (!x198x) & (!x283x)) + ((n_n4319) & (n_n4336) & (!n_n4321) & (!x198x) & (x283x)) + ((n_n4319) & (n_n4336) & (!n_n4321) & (x198x) & (!x283x)) + ((n_n4319) & (n_n4336) & (!n_n4321) & (x198x) & (x283x)) + ((n_n4319) & (n_n4336) & (n_n4321) & (!x198x) & (!x283x)) + ((n_n4319) & (n_n4336) & (n_n4321) & (!x198x) & (x283x)) + ((n_n4319) & (n_n4336) & (n_n4321) & (x198x) & (!x283x)) + ((n_n4319) & (n_n4336) & (n_n4321) & (x198x) & (x283x)));
	assign n_n2257 = (((!n_n4491) & (!n_n4497) & (!n_n3883) & (!x65x) & (x66x)) + ((!n_n4491) & (!n_n4497) & (!n_n3883) & (x65x) & (!x66x)) + ((!n_n4491) & (!n_n4497) & (!n_n3883) & (x65x) & (x66x)) + ((!n_n4491) & (!n_n4497) & (n_n3883) & (!x65x) & (!x66x)) + ((!n_n4491) & (!n_n4497) & (n_n3883) & (!x65x) & (x66x)) + ((!n_n4491) & (!n_n4497) & (n_n3883) & (x65x) & (!x66x)) + ((!n_n4491) & (!n_n4497) & (n_n3883) & (x65x) & (x66x)) + ((!n_n4491) & (n_n4497) & (!n_n3883) & (!x65x) & (!x66x)) + ((!n_n4491) & (n_n4497) & (!n_n3883) & (!x65x) & (x66x)) + ((!n_n4491) & (n_n4497) & (!n_n3883) & (x65x) & (!x66x)) + ((!n_n4491) & (n_n4497) & (!n_n3883) & (x65x) & (x66x)) + ((!n_n4491) & (n_n4497) & (n_n3883) & (!x65x) & (!x66x)) + ((!n_n4491) & (n_n4497) & (n_n3883) & (!x65x) & (x66x)) + ((!n_n4491) & (n_n4497) & (n_n3883) & (x65x) & (!x66x)) + ((!n_n4491) & (n_n4497) & (n_n3883) & (x65x) & (x66x)) + ((n_n4491) & (!n_n4497) & (!n_n3883) & (!x65x) & (!x66x)) + ((n_n4491) & (!n_n4497) & (!n_n3883) & (!x65x) & (x66x)) + ((n_n4491) & (!n_n4497) & (!n_n3883) & (x65x) & (!x66x)) + ((n_n4491) & (!n_n4497) & (!n_n3883) & (x65x) & (x66x)) + ((n_n4491) & (!n_n4497) & (n_n3883) & (!x65x) & (!x66x)) + ((n_n4491) & (!n_n4497) & (n_n3883) & (!x65x) & (x66x)) + ((n_n4491) & (!n_n4497) & (n_n3883) & (x65x) & (!x66x)) + ((n_n4491) & (!n_n4497) & (n_n3883) & (x65x) & (x66x)) + ((n_n4491) & (n_n4497) & (!n_n3883) & (!x65x) & (!x66x)) + ((n_n4491) & (n_n4497) & (!n_n3883) & (!x65x) & (x66x)) + ((n_n4491) & (n_n4497) & (!n_n3883) & (x65x) & (!x66x)) + ((n_n4491) & (n_n4497) & (!n_n3883) & (x65x) & (x66x)) + ((n_n4491) & (n_n4497) & (n_n3883) & (!x65x) & (!x66x)) + ((n_n4491) & (n_n4497) & (n_n3883) & (!x65x) & (x66x)) + ((n_n4491) & (n_n4497) & (n_n3883) & (x65x) & (!x66x)) + ((n_n4491) & (n_n4497) & (n_n3883) & (x65x) & (x66x)));
	assign n_n2258 = (((!n_n4487) & (!n_n4478) & (!n_n4254) & (!x70x) & (x184x)) + ((!n_n4487) & (!n_n4478) & (!n_n4254) & (x70x) & (!x184x)) + ((!n_n4487) & (!n_n4478) & (!n_n4254) & (x70x) & (x184x)) + ((!n_n4487) & (!n_n4478) & (n_n4254) & (!x70x) & (!x184x)) + ((!n_n4487) & (!n_n4478) & (n_n4254) & (!x70x) & (x184x)) + ((!n_n4487) & (!n_n4478) & (n_n4254) & (x70x) & (!x184x)) + ((!n_n4487) & (!n_n4478) & (n_n4254) & (x70x) & (x184x)) + ((!n_n4487) & (n_n4478) & (!n_n4254) & (!x70x) & (!x184x)) + ((!n_n4487) & (n_n4478) & (!n_n4254) & (!x70x) & (x184x)) + ((!n_n4487) & (n_n4478) & (!n_n4254) & (x70x) & (!x184x)) + ((!n_n4487) & (n_n4478) & (!n_n4254) & (x70x) & (x184x)) + ((!n_n4487) & (n_n4478) & (n_n4254) & (!x70x) & (!x184x)) + ((!n_n4487) & (n_n4478) & (n_n4254) & (!x70x) & (x184x)) + ((!n_n4487) & (n_n4478) & (n_n4254) & (x70x) & (!x184x)) + ((!n_n4487) & (n_n4478) & (n_n4254) & (x70x) & (x184x)) + ((n_n4487) & (!n_n4478) & (!n_n4254) & (!x70x) & (!x184x)) + ((n_n4487) & (!n_n4478) & (!n_n4254) & (!x70x) & (x184x)) + ((n_n4487) & (!n_n4478) & (!n_n4254) & (x70x) & (!x184x)) + ((n_n4487) & (!n_n4478) & (!n_n4254) & (x70x) & (x184x)) + ((n_n4487) & (!n_n4478) & (n_n4254) & (!x70x) & (!x184x)) + ((n_n4487) & (!n_n4478) & (n_n4254) & (!x70x) & (x184x)) + ((n_n4487) & (!n_n4478) & (n_n4254) & (x70x) & (!x184x)) + ((n_n4487) & (!n_n4478) & (n_n4254) & (x70x) & (x184x)) + ((n_n4487) & (n_n4478) & (!n_n4254) & (!x70x) & (!x184x)) + ((n_n4487) & (n_n4478) & (!n_n4254) & (!x70x) & (x184x)) + ((n_n4487) & (n_n4478) & (!n_n4254) & (x70x) & (!x184x)) + ((n_n4487) & (n_n4478) & (!n_n4254) & (x70x) & (x184x)) + ((n_n4487) & (n_n4478) & (n_n4254) & (!x70x) & (!x184x)) + ((n_n4487) & (n_n4478) & (n_n4254) & (!x70x) & (x184x)) + ((n_n4487) & (n_n4478) & (n_n4254) & (x70x) & (!x184x)) + ((n_n4487) & (n_n4478) & (n_n4254) & (x70x) & (x184x)));
	assign x16596x = (((!n_n4504) & (!n_n4503) & (!n_n4506) & (!n_n4505) & (x16595x)) + ((!n_n4504) & (!n_n4503) & (!n_n4506) & (n_n4505) & (!x16595x)) + ((!n_n4504) & (!n_n4503) & (!n_n4506) & (n_n4505) & (x16595x)) + ((!n_n4504) & (!n_n4503) & (n_n4506) & (!n_n4505) & (!x16595x)) + ((!n_n4504) & (!n_n4503) & (n_n4506) & (!n_n4505) & (x16595x)) + ((!n_n4504) & (!n_n4503) & (n_n4506) & (n_n4505) & (!x16595x)) + ((!n_n4504) & (!n_n4503) & (n_n4506) & (n_n4505) & (x16595x)) + ((!n_n4504) & (n_n4503) & (!n_n4506) & (!n_n4505) & (!x16595x)) + ((!n_n4504) & (n_n4503) & (!n_n4506) & (!n_n4505) & (x16595x)) + ((!n_n4504) & (n_n4503) & (!n_n4506) & (n_n4505) & (!x16595x)) + ((!n_n4504) & (n_n4503) & (!n_n4506) & (n_n4505) & (x16595x)) + ((!n_n4504) & (n_n4503) & (n_n4506) & (!n_n4505) & (!x16595x)) + ((!n_n4504) & (n_n4503) & (n_n4506) & (!n_n4505) & (x16595x)) + ((!n_n4504) & (n_n4503) & (n_n4506) & (n_n4505) & (!x16595x)) + ((!n_n4504) & (n_n4503) & (n_n4506) & (n_n4505) & (x16595x)) + ((n_n4504) & (!n_n4503) & (!n_n4506) & (!n_n4505) & (!x16595x)) + ((n_n4504) & (!n_n4503) & (!n_n4506) & (!n_n4505) & (x16595x)) + ((n_n4504) & (!n_n4503) & (!n_n4506) & (n_n4505) & (!x16595x)) + ((n_n4504) & (!n_n4503) & (!n_n4506) & (n_n4505) & (x16595x)) + ((n_n4504) & (!n_n4503) & (n_n4506) & (!n_n4505) & (!x16595x)) + ((n_n4504) & (!n_n4503) & (n_n4506) & (!n_n4505) & (x16595x)) + ((n_n4504) & (!n_n4503) & (n_n4506) & (n_n4505) & (!x16595x)) + ((n_n4504) & (!n_n4503) & (n_n4506) & (n_n4505) & (x16595x)) + ((n_n4504) & (n_n4503) & (!n_n4506) & (!n_n4505) & (!x16595x)) + ((n_n4504) & (n_n4503) & (!n_n4506) & (!n_n4505) & (x16595x)) + ((n_n4504) & (n_n4503) & (!n_n4506) & (n_n4505) & (!x16595x)) + ((n_n4504) & (n_n4503) & (!n_n4506) & (n_n4505) & (x16595x)) + ((n_n4504) & (n_n4503) & (n_n4506) & (!n_n4505) & (!x16595x)) + ((n_n4504) & (n_n4503) & (n_n4506) & (!n_n4505) & (x16595x)) + ((n_n4504) & (n_n4503) & (n_n4506) & (n_n4505) & (!x16595x)) + ((n_n4504) & (n_n4503) & (n_n4506) & (n_n4505) & (x16595x)));
	assign x16598x = (((!n_n2257) & (!n_n2258) & (x16596x)) + ((!n_n2257) & (n_n2258) & (!x16596x)) + ((!n_n2257) & (n_n2258) & (x16596x)) + ((n_n2257) & (!n_n2258) & (!x16596x)) + ((n_n2257) & (!n_n2258) & (x16596x)) + ((n_n2257) & (n_n2258) & (!x16596x)) + ((n_n2257) & (n_n2258) & (x16596x)));
	assign n_n2189 = (((!n_n2261) & (!x321x) & (!x16568x) & (x16569x)) + ((!n_n2261) & (!x321x) & (x16568x) & (!x16569x)) + ((!n_n2261) & (!x321x) & (x16568x) & (x16569x)) + ((!n_n2261) & (x321x) & (!x16568x) & (!x16569x)) + ((!n_n2261) & (x321x) & (!x16568x) & (x16569x)) + ((!n_n2261) & (x321x) & (x16568x) & (!x16569x)) + ((!n_n2261) & (x321x) & (x16568x) & (x16569x)) + ((n_n2261) & (!x321x) & (!x16568x) & (!x16569x)) + ((n_n2261) & (!x321x) & (!x16568x) & (x16569x)) + ((n_n2261) & (!x321x) & (x16568x) & (!x16569x)) + ((n_n2261) & (!x321x) & (x16568x) & (x16569x)) + ((n_n2261) & (x321x) & (!x16568x) & (!x16569x)) + ((n_n2261) & (x321x) & (!x16568x) & (x16569x)) + ((n_n2261) & (x321x) & (x16568x) & (!x16569x)) + ((n_n2261) & (x321x) & (x16568x) & (x16569x)));
	assign x16590x = (((!n_n4247) & (!n_n4511) & (!n_n4510) & (!n_n4528) & (!x22063x)) + ((!n_n4247) & (!n_n4511) & (!n_n4510) & (n_n4528) & (!x22063x)) + ((!n_n4247) & (!n_n4511) & (!n_n4510) & (n_n4528) & (x22063x)) + ((!n_n4247) & (!n_n4511) & (n_n4510) & (!n_n4528) & (!x22063x)) + ((!n_n4247) & (!n_n4511) & (n_n4510) & (!n_n4528) & (x22063x)) + ((!n_n4247) & (!n_n4511) & (n_n4510) & (n_n4528) & (!x22063x)) + ((!n_n4247) & (!n_n4511) & (n_n4510) & (n_n4528) & (x22063x)) + ((!n_n4247) & (n_n4511) & (!n_n4510) & (!n_n4528) & (!x22063x)) + ((!n_n4247) & (n_n4511) & (!n_n4510) & (!n_n4528) & (x22063x)) + ((!n_n4247) & (n_n4511) & (!n_n4510) & (n_n4528) & (!x22063x)) + ((!n_n4247) & (n_n4511) & (!n_n4510) & (n_n4528) & (x22063x)) + ((!n_n4247) & (n_n4511) & (n_n4510) & (!n_n4528) & (!x22063x)) + ((!n_n4247) & (n_n4511) & (n_n4510) & (!n_n4528) & (x22063x)) + ((!n_n4247) & (n_n4511) & (n_n4510) & (n_n4528) & (!x22063x)) + ((!n_n4247) & (n_n4511) & (n_n4510) & (n_n4528) & (x22063x)) + ((n_n4247) & (!n_n4511) & (!n_n4510) & (!n_n4528) & (!x22063x)) + ((n_n4247) & (!n_n4511) & (!n_n4510) & (!n_n4528) & (x22063x)) + ((n_n4247) & (!n_n4511) & (!n_n4510) & (n_n4528) & (!x22063x)) + ((n_n4247) & (!n_n4511) & (!n_n4510) & (n_n4528) & (x22063x)) + ((n_n4247) & (!n_n4511) & (n_n4510) & (!n_n4528) & (!x22063x)) + ((n_n4247) & (!n_n4511) & (n_n4510) & (!n_n4528) & (x22063x)) + ((n_n4247) & (!n_n4511) & (n_n4510) & (n_n4528) & (!x22063x)) + ((n_n4247) & (!n_n4511) & (n_n4510) & (n_n4528) & (x22063x)) + ((n_n4247) & (n_n4511) & (!n_n4510) & (!n_n4528) & (!x22063x)) + ((n_n4247) & (n_n4511) & (!n_n4510) & (!n_n4528) & (x22063x)) + ((n_n4247) & (n_n4511) & (!n_n4510) & (n_n4528) & (!x22063x)) + ((n_n4247) & (n_n4511) & (!n_n4510) & (n_n4528) & (x22063x)) + ((n_n4247) & (n_n4511) & (n_n4510) & (!n_n4528) & (!x22063x)) + ((n_n4247) & (n_n4511) & (n_n4510) & (!n_n4528) & (x22063x)) + ((n_n4247) & (n_n4511) & (n_n4510) & (n_n4528) & (!x22063x)) + ((n_n4247) & (n_n4511) & (n_n4510) & (n_n4528) & (x22063x)));
	assign n_n2253 = (((!n_n482) & (!n_n455) & (!x20x) & (!x23x) & (!x22208x)) + ((!n_n482) & (!n_n455) & (!x20x) & (x23x) & (!x22208x)) + ((!n_n482) & (!n_n455) & (x20x) & (!x23x) & (!x22208x)) + ((!n_n482) & (!n_n455) & (x20x) & (x23x) & (!x22208x)) + ((!n_n482) & (n_n455) & (!x20x) & (!x23x) & (!x22208x)) + ((!n_n482) & (n_n455) & (!x20x) & (x23x) & (!x22208x)) + ((!n_n482) & (n_n455) & (x20x) & (!x23x) & (!x22208x)) + ((!n_n482) & (n_n455) & (x20x) & (x23x) & (!x22208x)) + ((n_n482) & (!n_n455) & (!x20x) & (!x23x) & (!x22208x)) + ((n_n482) & (!n_n455) & (!x20x) & (x23x) & (!x22208x)) + ((n_n482) & (!n_n455) & (x20x) & (!x23x) & (!x22208x)) + ((n_n482) & (!n_n455) & (x20x) & (x23x) & (!x22208x)) + ((n_n482) & (n_n455) & (!x20x) & (!x23x) & (!x22208x)) + ((n_n482) & (n_n455) & (!x20x) & (x23x) & (!x22208x)) + ((n_n482) & (n_n455) & (!x20x) & (x23x) & (x22208x)) + ((n_n482) & (n_n455) & (x20x) & (!x23x) & (!x22208x)) + ((n_n482) & (n_n455) & (x20x) & (!x23x) & (x22208x)) + ((n_n482) & (n_n455) & (x20x) & (x23x) & (!x22208x)) + ((n_n482) & (n_n455) & (x20x) & (x23x) & (x22208x)));
	assign x16589x = (((!n_n4524) & (!n_n4525) & (!x178x) & (!x307x) & (x378x)) + ((!n_n4524) & (!n_n4525) & (!x178x) & (x307x) & (!x378x)) + ((!n_n4524) & (!n_n4525) & (!x178x) & (x307x) & (x378x)) + ((!n_n4524) & (!n_n4525) & (x178x) & (!x307x) & (!x378x)) + ((!n_n4524) & (!n_n4525) & (x178x) & (!x307x) & (x378x)) + ((!n_n4524) & (!n_n4525) & (x178x) & (x307x) & (!x378x)) + ((!n_n4524) & (!n_n4525) & (x178x) & (x307x) & (x378x)) + ((!n_n4524) & (n_n4525) & (!x178x) & (!x307x) & (!x378x)) + ((!n_n4524) & (n_n4525) & (!x178x) & (!x307x) & (x378x)) + ((!n_n4524) & (n_n4525) & (!x178x) & (x307x) & (!x378x)) + ((!n_n4524) & (n_n4525) & (!x178x) & (x307x) & (x378x)) + ((!n_n4524) & (n_n4525) & (x178x) & (!x307x) & (!x378x)) + ((!n_n4524) & (n_n4525) & (x178x) & (!x307x) & (x378x)) + ((!n_n4524) & (n_n4525) & (x178x) & (x307x) & (!x378x)) + ((!n_n4524) & (n_n4525) & (x178x) & (x307x) & (x378x)) + ((n_n4524) & (!n_n4525) & (!x178x) & (!x307x) & (!x378x)) + ((n_n4524) & (!n_n4525) & (!x178x) & (!x307x) & (x378x)) + ((n_n4524) & (!n_n4525) & (!x178x) & (x307x) & (!x378x)) + ((n_n4524) & (!n_n4525) & (!x178x) & (x307x) & (x378x)) + ((n_n4524) & (!n_n4525) & (x178x) & (!x307x) & (!x378x)) + ((n_n4524) & (!n_n4525) & (x178x) & (!x307x) & (x378x)) + ((n_n4524) & (!n_n4525) & (x178x) & (x307x) & (!x378x)) + ((n_n4524) & (!n_n4525) & (x178x) & (x307x) & (x378x)) + ((n_n4524) & (n_n4525) & (!x178x) & (!x307x) & (!x378x)) + ((n_n4524) & (n_n4525) & (!x178x) & (!x307x) & (x378x)) + ((n_n4524) & (n_n4525) & (!x178x) & (x307x) & (!x378x)) + ((n_n4524) & (n_n4525) & (!x178x) & (x307x) & (x378x)) + ((n_n4524) & (n_n4525) & (x178x) & (!x307x) & (!x378x)) + ((n_n4524) & (n_n4525) & (x178x) & (!x307x) & (x378x)) + ((n_n4524) & (n_n4525) & (x178x) & (x307x) & (!x378x)) + ((n_n4524) & (n_n4525) & (x178x) & (x307x) & (x378x)));
	assign n_n2251 = (((!n_n4561) & (!n_n4568) & (!x455x) & (!x121x) & (n_n4239)) + ((!n_n4561) & (!n_n4568) & (!x455x) & (x121x) & (!n_n4239)) + ((!n_n4561) & (!n_n4568) & (!x455x) & (x121x) & (n_n4239)) + ((!n_n4561) & (!n_n4568) & (x455x) & (!x121x) & (!n_n4239)) + ((!n_n4561) & (!n_n4568) & (x455x) & (!x121x) & (n_n4239)) + ((!n_n4561) & (!n_n4568) & (x455x) & (x121x) & (!n_n4239)) + ((!n_n4561) & (!n_n4568) & (x455x) & (x121x) & (n_n4239)) + ((!n_n4561) & (n_n4568) & (!x455x) & (!x121x) & (!n_n4239)) + ((!n_n4561) & (n_n4568) & (!x455x) & (!x121x) & (n_n4239)) + ((!n_n4561) & (n_n4568) & (!x455x) & (x121x) & (!n_n4239)) + ((!n_n4561) & (n_n4568) & (!x455x) & (x121x) & (n_n4239)) + ((!n_n4561) & (n_n4568) & (x455x) & (!x121x) & (!n_n4239)) + ((!n_n4561) & (n_n4568) & (x455x) & (!x121x) & (n_n4239)) + ((!n_n4561) & (n_n4568) & (x455x) & (x121x) & (!n_n4239)) + ((!n_n4561) & (n_n4568) & (x455x) & (x121x) & (n_n4239)) + ((n_n4561) & (!n_n4568) & (!x455x) & (!x121x) & (!n_n4239)) + ((n_n4561) & (!n_n4568) & (!x455x) & (!x121x) & (n_n4239)) + ((n_n4561) & (!n_n4568) & (!x455x) & (x121x) & (!n_n4239)) + ((n_n4561) & (!n_n4568) & (!x455x) & (x121x) & (n_n4239)) + ((n_n4561) & (!n_n4568) & (x455x) & (!x121x) & (!n_n4239)) + ((n_n4561) & (!n_n4568) & (x455x) & (!x121x) & (n_n4239)) + ((n_n4561) & (!n_n4568) & (x455x) & (x121x) & (!n_n4239)) + ((n_n4561) & (!n_n4568) & (x455x) & (x121x) & (n_n4239)) + ((n_n4561) & (n_n4568) & (!x455x) & (!x121x) & (!n_n4239)) + ((n_n4561) & (n_n4568) & (!x455x) & (!x121x) & (n_n4239)) + ((n_n4561) & (n_n4568) & (!x455x) & (x121x) & (!n_n4239)) + ((n_n4561) & (n_n4568) & (!x455x) & (x121x) & (n_n4239)) + ((n_n4561) & (n_n4568) & (x455x) & (!x121x) & (!n_n4239)) + ((n_n4561) & (n_n4568) & (x455x) & (!x121x) & (n_n4239)) + ((n_n4561) & (n_n4568) & (x455x) & (x121x) & (!n_n4239)) + ((n_n4561) & (n_n4568) & (x455x) & (x121x) & (n_n4239)));
	assign x16606x = (((!n_n4584) & (!n_n4577) & (!n_n4576) & (!n_n4583) & (n_n4580)) + ((!n_n4584) & (!n_n4577) & (!n_n4576) & (n_n4583) & (!n_n4580)) + ((!n_n4584) & (!n_n4577) & (!n_n4576) & (n_n4583) & (n_n4580)) + ((!n_n4584) & (!n_n4577) & (n_n4576) & (!n_n4583) & (!n_n4580)) + ((!n_n4584) & (!n_n4577) & (n_n4576) & (!n_n4583) & (n_n4580)) + ((!n_n4584) & (!n_n4577) & (n_n4576) & (n_n4583) & (!n_n4580)) + ((!n_n4584) & (!n_n4577) & (n_n4576) & (n_n4583) & (n_n4580)) + ((!n_n4584) & (n_n4577) & (!n_n4576) & (!n_n4583) & (!n_n4580)) + ((!n_n4584) & (n_n4577) & (!n_n4576) & (!n_n4583) & (n_n4580)) + ((!n_n4584) & (n_n4577) & (!n_n4576) & (n_n4583) & (!n_n4580)) + ((!n_n4584) & (n_n4577) & (!n_n4576) & (n_n4583) & (n_n4580)) + ((!n_n4584) & (n_n4577) & (n_n4576) & (!n_n4583) & (!n_n4580)) + ((!n_n4584) & (n_n4577) & (n_n4576) & (!n_n4583) & (n_n4580)) + ((!n_n4584) & (n_n4577) & (n_n4576) & (n_n4583) & (!n_n4580)) + ((!n_n4584) & (n_n4577) & (n_n4576) & (n_n4583) & (n_n4580)) + ((n_n4584) & (!n_n4577) & (!n_n4576) & (!n_n4583) & (!n_n4580)) + ((n_n4584) & (!n_n4577) & (!n_n4576) & (!n_n4583) & (n_n4580)) + ((n_n4584) & (!n_n4577) & (!n_n4576) & (n_n4583) & (!n_n4580)) + ((n_n4584) & (!n_n4577) & (!n_n4576) & (n_n4583) & (n_n4580)) + ((n_n4584) & (!n_n4577) & (n_n4576) & (!n_n4583) & (!n_n4580)) + ((n_n4584) & (!n_n4577) & (n_n4576) & (!n_n4583) & (n_n4580)) + ((n_n4584) & (!n_n4577) & (n_n4576) & (n_n4583) & (!n_n4580)) + ((n_n4584) & (!n_n4577) & (n_n4576) & (n_n4583) & (n_n4580)) + ((n_n4584) & (n_n4577) & (!n_n4576) & (!n_n4583) & (!n_n4580)) + ((n_n4584) & (n_n4577) & (!n_n4576) & (!n_n4583) & (n_n4580)) + ((n_n4584) & (n_n4577) & (!n_n4576) & (n_n4583) & (!n_n4580)) + ((n_n4584) & (n_n4577) & (!n_n4576) & (n_n4583) & (n_n4580)) + ((n_n4584) & (n_n4577) & (n_n4576) & (!n_n4583) & (!n_n4580)) + ((n_n4584) & (n_n4577) & (n_n4576) & (!n_n4583) & (n_n4580)) + ((n_n4584) & (n_n4577) & (n_n4576) & (n_n4583) & (!n_n4580)) + ((n_n4584) & (n_n4577) & (n_n4576) & (n_n4583) & (n_n4580)));
	assign x16642x = (((!n_n4554) & (!n_n4546) & (!n_n4555) & (!n_n4549) & (n_n4548)) + ((!n_n4554) & (!n_n4546) & (!n_n4555) & (n_n4549) & (!n_n4548)) + ((!n_n4554) & (!n_n4546) & (!n_n4555) & (n_n4549) & (n_n4548)) + ((!n_n4554) & (!n_n4546) & (n_n4555) & (!n_n4549) & (!n_n4548)) + ((!n_n4554) & (!n_n4546) & (n_n4555) & (!n_n4549) & (n_n4548)) + ((!n_n4554) & (!n_n4546) & (n_n4555) & (n_n4549) & (!n_n4548)) + ((!n_n4554) & (!n_n4546) & (n_n4555) & (n_n4549) & (n_n4548)) + ((!n_n4554) & (n_n4546) & (!n_n4555) & (!n_n4549) & (!n_n4548)) + ((!n_n4554) & (n_n4546) & (!n_n4555) & (!n_n4549) & (n_n4548)) + ((!n_n4554) & (n_n4546) & (!n_n4555) & (n_n4549) & (!n_n4548)) + ((!n_n4554) & (n_n4546) & (!n_n4555) & (n_n4549) & (n_n4548)) + ((!n_n4554) & (n_n4546) & (n_n4555) & (!n_n4549) & (!n_n4548)) + ((!n_n4554) & (n_n4546) & (n_n4555) & (!n_n4549) & (n_n4548)) + ((!n_n4554) & (n_n4546) & (n_n4555) & (n_n4549) & (!n_n4548)) + ((!n_n4554) & (n_n4546) & (n_n4555) & (n_n4549) & (n_n4548)) + ((n_n4554) & (!n_n4546) & (!n_n4555) & (!n_n4549) & (!n_n4548)) + ((n_n4554) & (!n_n4546) & (!n_n4555) & (!n_n4549) & (n_n4548)) + ((n_n4554) & (!n_n4546) & (!n_n4555) & (n_n4549) & (!n_n4548)) + ((n_n4554) & (!n_n4546) & (!n_n4555) & (n_n4549) & (n_n4548)) + ((n_n4554) & (!n_n4546) & (n_n4555) & (!n_n4549) & (!n_n4548)) + ((n_n4554) & (!n_n4546) & (n_n4555) & (!n_n4549) & (n_n4548)) + ((n_n4554) & (!n_n4546) & (n_n4555) & (n_n4549) & (!n_n4548)) + ((n_n4554) & (!n_n4546) & (n_n4555) & (n_n4549) & (n_n4548)) + ((n_n4554) & (n_n4546) & (!n_n4555) & (!n_n4549) & (!n_n4548)) + ((n_n4554) & (n_n4546) & (!n_n4555) & (!n_n4549) & (n_n4548)) + ((n_n4554) & (n_n4546) & (!n_n4555) & (n_n4549) & (!n_n4548)) + ((n_n4554) & (n_n4546) & (!n_n4555) & (n_n4549) & (n_n4548)) + ((n_n4554) & (n_n4546) & (n_n4555) & (!n_n4549) & (!n_n4548)) + ((n_n4554) & (n_n4546) & (n_n4555) & (!n_n4549) & (n_n4548)) + ((n_n4554) & (n_n4546) & (n_n4555) & (n_n4549) & (!n_n4548)) + ((n_n4554) & (n_n4546) & (n_n4555) & (n_n4549) & (n_n4548)));
	assign x22062x = (((!x213x) & (!n_n4551) & (!n_n4552) & (!x238x) & (!x276x)));
	assign x16645x = (((!n_n2251) & (!x16606x) & (!x16642x) & (!x22062x)) + ((!n_n2251) & (!x16606x) & (x16642x) & (!x22062x)) + ((!n_n2251) & (!x16606x) & (x16642x) & (x22062x)) + ((!n_n2251) & (x16606x) & (!x16642x) & (!x22062x)) + ((!n_n2251) & (x16606x) & (!x16642x) & (x22062x)) + ((!n_n2251) & (x16606x) & (x16642x) & (!x22062x)) + ((!n_n2251) & (x16606x) & (x16642x) & (x22062x)) + ((n_n2251) & (!x16606x) & (!x16642x) & (!x22062x)) + ((n_n2251) & (!x16606x) & (!x16642x) & (x22062x)) + ((n_n2251) & (!x16606x) & (x16642x) & (!x22062x)) + ((n_n2251) & (!x16606x) & (x16642x) & (x22062x)) + ((n_n2251) & (x16606x) & (!x16642x) & (!x22062x)) + ((n_n2251) & (x16606x) & (!x16642x) & (x22062x)) + ((n_n2251) & (x16606x) & (x16642x) & (!x22062x)) + ((n_n2251) & (x16606x) & (x16642x) & (x22062x)));
	assign n_n2185 = (((!x16622x) & (!x16611x) & (!x16612x) & (!x16617x) & (x16618x)) + ((!x16622x) & (!x16611x) & (!x16612x) & (x16617x) & (!x16618x)) + ((!x16622x) & (!x16611x) & (!x16612x) & (x16617x) & (x16618x)) + ((!x16622x) & (!x16611x) & (x16612x) & (!x16617x) & (!x16618x)) + ((!x16622x) & (!x16611x) & (x16612x) & (!x16617x) & (x16618x)) + ((!x16622x) & (!x16611x) & (x16612x) & (x16617x) & (!x16618x)) + ((!x16622x) & (!x16611x) & (x16612x) & (x16617x) & (x16618x)) + ((!x16622x) & (x16611x) & (!x16612x) & (!x16617x) & (!x16618x)) + ((!x16622x) & (x16611x) & (!x16612x) & (!x16617x) & (x16618x)) + ((!x16622x) & (x16611x) & (!x16612x) & (x16617x) & (!x16618x)) + ((!x16622x) & (x16611x) & (!x16612x) & (x16617x) & (x16618x)) + ((!x16622x) & (x16611x) & (x16612x) & (!x16617x) & (!x16618x)) + ((!x16622x) & (x16611x) & (x16612x) & (!x16617x) & (x16618x)) + ((!x16622x) & (x16611x) & (x16612x) & (x16617x) & (!x16618x)) + ((!x16622x) & (x16611x) & (x16612x) & (x16617x) & (x16618x)) + ((x16622x) & (!x16611x) & (!x16612x) & (!x16617x) & (!x16618x)) + ((x16622x) & (!x16611x) & (!x16612x) & (!x16617x) & (x16618x)) + ((x16622x) & (!x16611x) & (!x16612x) & (x16617x) & (!x16618x)) + ((x16622x) & (!x16611x) & (!x16612x) & (x16617x) & (x16618x)) + ((x16622x) & (!x16611x) & (x16612x) & (!x16617x) & (!x16618x)) + ((x16622x) & (!x16611x) & (x16612x) & (!x16617x) & (x16618x)) + ((x16622x) & (!x16611x) & (x16612x) & (x16617x) & (!x16618x)) + ((x16622x) & (!x16611x) & (x16612x) & (x16617x) & (x16618x)) + ((x16622x) & (x16611x) & (!x16612x) & (!x16617x) & (!x16618x)) + ((x16622x) & (x16611x) & (!x16612x) & (!x16617x) & (x16618x)) + ((x16622x) & (x16611x) & (!x16612x) & (x16617x) & (!x16618x)) + ((x16622x) & (x16611x) & (!x16612x) & (x16617x) & (x16618x)) + ((x16622x) & (x16611x) & (x16612x) & (!x16617x) & (!x16618x)) + ((x16622x) & (x16611x) & (x16612x) & (!x16617x) & (x16618x)) + ((x16622x) & (x16611x) & (x16612x) & (x16617x) & (!x16618x)) + ((x16622x) & (x16611x) & (x16612x) & (x16617x) & (x16618x)));
	assign n_n2184 = (((!x16628x) & (!n_n2246) & (!x16636x) & (!x22061x)) + ((!x16628x) & (!n_n2246) & (x16636x) & (!x22061x)) + ((!x16628x) & (!n_n2246) & (x16636x) & (x22061x)) + ((!x16628x) & (n_n2246) & (!x16636x) & (!x22061x)) + ((!x16628x) & (n_n2246) & (!x16636x) & (x22061x)) + ((!x16628x) & (n_n2246) & (x16636x) & (!x22061x)) + ((!x16628x) & (n_n2246) & (x16636x) & (x22061x)) + ((x16628x) & (!n_n2246) & (!x16636x) & (!x22061x)) + ((x16628x) & (!n_n2246) & (!x16636x) & (x22061x)) + ((x16628x) & (!n_n2246) & (x16636x) & (!x22061x)) + ((x16628x) & (!n_n2246) & (x16636x) & (x22061x)) + ((x16628x) & (n_n2246) & (!x16636x) & (!x22061x)) + ((x16628x) & (n_n2246) & (!x16636x) & (x22061x)) + ((x16628x) & (n_n2246) & (x16636x) & (!x22061x)) + ((x16628x) & (n_n2246) & (x16636x) & (x22061x)));
	assign n_n4380 = (((i_9_) & (n_n536) & (n_n491) & (n_n530)));
	assign x16651x = (((!n_n4338) & (!n_n4325) & (!n_n4380) & (n_n4345)) + ((!n_n4338) & (!n_n4325) & (n_n4380) & (!n_n4345)) + ((!n_n4338) & (!n_n4325) & (n_n4380) & (n_n4345)) + ((!n_n4338) & (n_n4325) & (!n_n4380) & (!n_n4345)) + ((!n_n4338) & (n_n4325) & (!n_n4380) & (n_n4345)) + ((!n_n4338) & (n_n4325) & (n_n4380) & (!n_n4345)) + ((!n_n4338) & (n_n4325) & (n_n4380) & (n_n4345)) + ((n_n4338) & (!n_n4325) & (!n_n4380) & (!n_n4345)) + ((n_n4338) & (!n_n4325) & (!n_n4380) & (n_n4345)) + ((n_n4338) & (!n_n4325) & (n_n4380) & (!n_n4345)) + ((n_n4338) & (!n_n4325) & (n_n4380) & (n_n4345)) + ((n_n4338) & (n_n4325) & (!n_n4380) & (!n_n4345)) + ((n_n4338) & (n_n4325) & (!n_n4380) & (n_n4345)) + ((n_n4338) & (n_n4325) & (n_n4380) & (!n_n4345)) + ((n_n4338) & (n_n4325) & (n_n4380) & (n_n4345)));
	assign n_n4367 = (((!i_9_) & (n_n536) & (n_n528) & (n_n500)));
	assign n_n4374 = (((i_9_) & (n_n536) & (n_n520) & (n_n500)));
	assign x16652x = (((!n_n4367) & (!n_n4374) & (!n_n4341) & (!n_n4357) & (n_n4358)) + ((!n_n4367) & (!n_n4374) & (!n_n4341) & (n_n4357) & (!n_n4358)) + ((!n_n4367) & (!n_n4374) & (!n_n4341) & (n_n4357) & (n_n4358)) + ((!n_n4367) & (!n_n4374) & (n_n4341) & (!n_n4357) & (!n_n4358)) + ((!n_n4367) & (!n_n4374) & (n_n4341) & (!n_n4357) & (n_n4358)) + ((!n_n4367) & (!n_n4374) & (n_n4341) & (n_n4357) & (!n_n4358)) + ((!n_n4367) & (!n_n4374) & (n_n4341) & (n_n4357) & (n_n4358)) + ((!n_n4367) & (n_n4374) & (!n_n4341) & (!n_n4357) & (!n_n4358)) + ((!n_n4367) & (n_n4374) & (!n_n4341) & (!n_n4357) & (n_n4358)) + ((!n_n4367) & (n_n4374) & (!n_n4341) & (n_n4357) & (!n_n4358)) + ((!n_n4367) & (n_n4374) & (!n_n4341) & (n_n4357) & (n_n4358)) + ((!n_n4367) & (n_n4374) & (n_n4341) & (!n_n4357) & (!n_n4358)) + ((!n_n4367) & (n_n4374) & (n_n4341) & (!n_n4357) & (n_n4358)) + ((!n_n4367) & (n_n4374) & (n_n4341) & (n_n4357) & (!n_n4358)) + ((!n_n4367) & (n_n4374) & (n_n4341) & (n_n4357) & (n_n4358)) + ((n_n4367) & (!n_n4374) & (!n_n4341) & (!n_n4357) & (!n_n4358)) + ((n_n4367) & (!n_n4374) & (!n_n4341) & (!n_n4357) & (n_n4358)) + ((n_n4367) & (!n_n4374) & (!n_n4341) & (n_n4357) & (!n_n4358)) + ((n_n4367) & (!n_n4374) & (!n_n4341) & (n_n4357) & (n_n4358)) + ((n_n4367) & (!n_n4374) & (n_n4341) & (!n_n4357) & (!n_n4358)) + ((n_n4367) & (!n_n4374) & (n_n4341) & (!n_n4357) & (n_n4358)) + ((n_n4367) & (!n_n4374) & (n_n4341) & (n_n4357) & (!n_n4358)) + ((n_n4367) & (!n_n4374) & (n_n4341) & (n_n4357) & (n_n4358)) + ((n_n4367) & (n_n4374) & (!n_n4341) & (!n_n4357) & (!n_n4358)) + ((n_n4367) & (n_n4374) & (!n_n4341) & (!n_n4357) & (n_n4358)) + ((n_n4367) & (n_n4374) & (!n_n4341) & (n_n4357) & (!n_n4358)) + ((n_n4367) & (n_n4374) & (!n_n4341) & (n_n4357) & (n_n4358)) + ((n_n4367) & (n_n4374) & (n_n4341) & (!n_n4357) & (!n_n4358)) + ((n_n4367) & (n_n4374) & (n_n4341) & (!n_n4357) & (n_n4358)) + ((n_n4367) & (n_n4374) & (n_n4341) & (n_n4357) & (!n_n4358)) + ((n_n4367) & (n_n4374) & (n_n4341) & (n_n4357) & (n_n4358)));
	assign x467x = (((!n_n5031) & (!n_n5024) & (!x13400x) & (!x111x) & (x253x)) + ((!n_n5031) & (!n_n5024) & (!x13400x) & (x111x) & (!x253x)) + ((!n_n5031) & (!n_n5024) & (!x13400x) & (x111x) & (x253x)) + ((!n_n5031) & (!n_n5024) & (x13400x) & (!x111x) & (!x253x)) + ((!n_n5031) & (!n_n5024) & (x13400x) & (!x111x) & (x253x)) + ((!n_n5031) & (!n_n5024) & (x13400x) & (x111x) & (!x253x)) + ((!n_n5031) & (!n_n5024) & (x13400x) & (x111x) & (x253x)) + ((!n_n5031) & (n_n5024) & (!x13400x) & (!x111x) & (!x253x)) + ((!n_n5031) & (n_n5024) & (!x13400x) & (!x111x) & (x253x)) + ((!n_n5031) & (n_n5024) & (!x13400x) & (x111x) & (!x253x)) + ((!n_n5031) & (n_n5024) & (!x13400x) & (x111x) & (x253x)) + ((!n_n5031) & (n_n5024) & (x13400x) & (!x111x) & (!x253x)) + ((!n_n5031) & (n_n5024) & (x13400x) & (!x111x) & (x253x)) + ((!n_n5031) & (n_n5024) & (x13400x) & (x111x) & (!x253x)) + ((!n_n5031) & (n_n5024) & (x13400x) & (x111x) & (x253x)) + ((n_n5031) & (!n_n5024) & (!x13400x) & (!x111x) & (!x253x)) + ((n_n5031) & (!n_n5024) & (!x13400x) & (!x111x) & (x253x)) + ((n_n5031) & (!n_n5024) & (!x13400x) & (x111x) & (!x253x)) + ((n_n5031) & (!n_n5024) & (!x13400x) & (x111x) & (x253x)) + ((n_n5031) & (!n_n5024) & (x13400x) & (!x111x) & (!x253x)) + ((n_n5031) & (!n_n5024) & (x13400x) & (!x111x) & (x253x)) + ((n_n5031) & (!n_n5024) & (x13400x) & (x111x) & (!x253x)) + ((n_n5031) & (!n_n5024) & (x13400x) & (x111x) & (x253x)) + ((n_n5031) & (n_n5024) & (!x13400x) & (!x111x) & (!x253x)) + ((n_n5031) & (n_n5024) & (!x13400x) & (!x111x) & (x253x)) + ((n_n5031) & (n_n5024) & (!x13400x) & (x111x) & (!x253x)) + ((n_n5031) & (n_n5024) & (!x13400x) & (x111x) & (x253x)) + ((n_n5031) & (n_n5024) & (x13400x) & (!x111x) & (!x253x)) + ((n_n5031) & (n_n5024) & (x13400x) & (!x111x) & (x253x)) + ((n_n5031) & (n_n5024) & (x13400x) & (x111x) & (!x253x)) + ((n_n5031) & (n_n5024) & (x13400x) & (x111x) & (x253x)));
	assign n_n2173 = (((!x16715x) & (!x90x) & (!x16711x) & (x16713x)) + ((!x16715x) & (!x90x) & (x16711x) & (!x16713x)) + ((!x16715x) & (!x90x) & (x16711x) & (x16713x)) + ((!x16715x) & (x90x) & (!x16711x) & (!x16713x)) + ((!x16715x) & (x90x) & (!x16711x) & (x16713x)) + ((!x16715x) & (x90x) & (x16711x) & (!x16713x)) + ((!x16715x) & (x90x) & (x16711x) & (x16713x)) + ((x16715x) & (!x90x) & (!x16711x) & (!x16713x)) + ((x16715x) & (!x90x) & (!x16711x) & (x16713x)) + ((x16715x) & (!x90x) & (x16711x) & (!x16713x)) + ((x16715x) & (!x90x) & (x16711x) & (x16713x)) + ((x16715x) & (x90x) & (!x16711x) & (!x16713x)) + ((x16715x) & (x90x) & (!x16711x) & (x16713x)) + ((x16715x) & (x90x) & (x16711x) & (!x16713x)) + ((x16715x) & (x90x) & (x16711x) & (x16713x)));
	assign n_n2172 = (((!n_n2210) & (!n_n2209) & (!x16728x) & (x16729x)) + ((!n_n2210) & (!n_n2209) & (x16728x) & (!x16729x)) + ((!n_n2210) & (!n_n2209) & (x16728x) & (x16729x)) + ((!n_n2210) & (n_n2209) & (!x16728x) & (!x16729x)) + ((!n_n2210) & (n_n2209) & (!x16728x) & (x16729x)) + ((!n_n2210) & (n_n2209) & (x16728x) & (!x16729x)) + ((!n_n2210) & (n_n2209) & (x16728x) & (x16729x)) + ((n_n2210) & (!n_n2209) & (!x16728x) & (!x16729x)) + ((n_n2210) & (!n_n2209) & (!x16728x) & (x16729x)) + ((n_n2210) & (!n_n2209) & (x16728x) & (!x16729x)) + ((n_n2210) & (!n_n2209) & (x16728x) & (x16729x)) + ((n_n2210) & (n_n2209) & (!x16728x) & (!x16729x)) + ((n_n2210) & (n_n2209) & (!x16728x) & (x16729x)) + ((n_n2210) & (n_n2209) & (x16728x) & (!x16729x)) + ((n_n2210) & (n_n2209) & (x16728x) & (x16729x)));
	assign n_n2214 = (((!n_n5059) & (!n_n5053) & (!n_n5052) & (!x275x) & (!x22221x)) + ((!n_n5059) & (!n_n5053) & (!n_n5052) & (x275x) & (!x22221x)) + ((!n_n5059) & (!n_n5053) & (!n_n5052) & (x275x) & (x22221x)) + ((!n_n5059) & (!n_n5053) & (n_n5052) & (!x275x) & (!x22221x)) + ((!n_n5059) & (!n_n5053) & (n_n5052) & (!x275x) & (x22221x)) + ((!n_n5059) & (!n_n5053) & (n_n5052) & (x275x) & (!x22221x)) + ((!n_n5059) & (!n_n5053) & (n_n5052) & (x275x) & (x22221x)) + ((!n_n5059) & (n_n5053) & (!n_n5052) & (!x275x) & (!x22221x)) + ((!n_n5059) & (n_n5053) & (!n_n5052) & (!x275x) & (x22221x)) + ((!n_n5059) & (n_n5053) & (!n_n5052) & (x275x) & (!x22221x)) + ((!n_n5059) & (n_n5053) & (!n_n5052) & (x275x) & (x22221x)) + ((!n_n5059) & (n_n5053) & (n_n5052) & (!x275x) & (!x22221x)) + ((!n_n5059) & (n_n5053) & (n_n5052) & (!x275x) & (x22221x)) + ((!n_n5059) & (n_n5053) & (n_n5052) & (x275x) & (!x22221x)) + ((!n_n5059) & (n_n5053) & (n_n5052) & (x275x) & (x22221x)) + ((n_n5059) & (!n_n5053) & (!n_n5052) & (!x275x) & (!x22221x)) + ((n_n5059) & (!n_n5053) & (!n_n5052) & (!x275x) & (x22221x)) + ((n_n5059) & (!n_n5053) & (!n_n5052) & (x275x) & (!x22221x)) + ((n_n5059) & (!n_n5053) & (!n_n5052) & (x275x) & (x22221x)) + ((n_n5059) & (!n_n5053) & (n_n5052) & (!x275x) & (!x22221x)) + ((n_n5059) & (!n_n5053) & (n_n5052) & (!x275x) & (x22221x)) + ((n_n5059) & (!n_n5053) & (n_n5052) & (x275x) & (!x22221x)) + ((n_n5059) & (!n_n5053) & (n_n5052) & (x275x) & (x22221x)) + ((n_n5059) & (n_n5053) & (!n_n5052) & (!x275x) & (!x22221x)) + ((n_n5059) & (n_n5053) & (!n_n5052) & (!x275x) & (x22221x)) + ((n_n5059) & (n_n5053) & (!n_n5052) & (x275x) & (!x22221x)) + ((n_n5059) & (n_n5053) & (!n_n5052) & (x275x) & (x22221x)) + ((n_n5059) & (n_n5053) & (n_n5052) & (!x275x) & (!x22221x)) + ((n_n5059) & (n_n5053) & (n_n5052) & (!x275x) & (x22221x)) + ((n_n5059) & (n_n5053) & (n_n5052) & (x275x) & (!x22221x)) + ((n_n5059) & (n_n5053) & (n_n5052) & (x275x) & (x22221x)));
	assign x16742x = (((!n_n5040) & (!n_n5048) & (!n_n5036) & (!n_n5047) & (x16741x)) + ((!n_n5040) & (!n_n5048) & (!n_n5036) & (n_n5047) & (!x16741x)) + ((!n_n5040) & (!n_n5048) & (!n_n5036) & (n_n5047) & (x16741x)) + ((!n_n5040) & (!n_n5048) & (n_n5036) & (!n_n5047) & (!x16741x)) + ((!n_n5040) & (!n_n5048) & (n_n5036) & (!n_n5047) & (x16741x)) + ((!n_n5040) & (!n_n5048) & (n_n5036) & (n_n5047) & (!x16741x)) + ((!n_n5040) & (!n_n5048) & (n_n5036) & (n_n5047) & (x16741x)) + ((!n_n5040) & (n_n5048) & (!n_n5036) & (!n_n5047) & (!x16741x)) + ((!n_n5040) & (n_n5048) & (!n_n5036) & (!n_n5047) & (x16741x)) + ((!n_n5040) & (n_n5048) & (!n_n5036) & (n_n5047) & (!x16741x)) + ((!n_n5040) & (n_n5048) & (!n_n5036) & (n_n5047) & (x16741x)) + ((!n_n5040) & (n_n5048) & (n_n5036) & (!n_n5047) & (!x16741x)) + ((!n_n5040) & (n_n5048) & (n_n5036) & (!n_n5047) & (x16741x)) + ((!n_n5040) & (n_n5048) & (n_n5036) & (n_n5047) & (!x16741x)) + ((!n_n5040) & (n_n5048) & (n_n5036) & (n_n5047) & (x16741x)) + ((n_n5040) & (!n_n5048) & (!n_n5036) & (!n_n5047) & (!x16741x)) + ((n_n5040) & (!n_n5048) & (!n_n5036) & (!n_n5047) & (x16741x)) + ((n_n5040) & (!n_n5048) & (!n_n5036) & (n_n5047) & (!x16741x)) + ((n_n5040) & (!n_n5048) & (!n_n5036) & (n_n5047) & (x16741x)) + ((n_n5040) & (!n_n5048) & (n_n5036) & (!n_n5047) & (!x16741x)) + ((n_n5040) & (!n_n5048) & (n_n5036) & (!n_n5047) & (x16741x)) + ((n_n5040) & (!n_n5048) & (n_n5036) & (n_n5047) & (!x16741x)) + ((n_n5040) & (!n_n5048) & (n_n5036) & (n_n5047) & (x16741x)) + ((n_n5040) & (n_n5048) & (!n_n5036) & (!n_n5047) & (!x16741x)) + ((n_n5040) & (n_n5048) & (!n_n5036) & (!n_n5047) & (x16741x)) + ((n_n5040) & (n_n5048) & (!n_n5036) & (n_n5047) & (!x16741x)) + ((n_n5040) & (n_n5048) & (!n_n5036) & (n_n5047) & (x16741x)) + ((n_n5040) & (n_n5048) & (n_n5036) & (!n_n5047) & (!x16741x)) + ((n_n5040) & (n_n5048) & (n_n5036) & (!n_n5047) & (x16741x)) + ((n_n5040) & (n_n5048) & (n_n5036) & (n_n5047) & (!x16741x)) + ((n_n5040) & (n_n5048) & (n_n5036) & (n_n5047) & (x16741x)));
	assign n_n2170 = (((!x16682x) & (!n_n2204) & (x16681x)) + ((!x16682x) & (n_n2204) & (!x16681x)) + ((!x16682x) & (n_n2204) & (x16681x)) + ((x16682x) & (!n_n2204) & (!x16681x)) + ((x16682x) & (!n_n2204) & (x16681x)) + ((x16682x) & (n_n2204) & (!x16681x)) + ((x16682x) & (n_n2204) & (x16681x)));
	assign n_n2169 = (((!n_n5251) & (!x435x) & (!n_n1139) & (!x16697x) & (x16693x)) + ((!n_n5251) & (!x435x) & (!n_n1139) & (x16697x) & (!x16693x)) + ((!n_n5251) & (!x435x) & (!n_n1139) & (x16697x) & (x16693x)) + ((!n_n5251) & (!x435x) & (n_n1139) & (!x16697x) & (!x16693x)) + ((!n_n5251) & (!x435x) & (n_n1139) & (!x16697x) & (x16693x)) + ((!n_n5251) & (!x435x) & (n_n1139) & (x16697x) & (!x16693x)) + ((!n_n5251) & (!x435x) & (n_n1139) & (x16697x) & (x16693x)) + ((!n_n5251) & (x435x) & (!n_n1139) & (!x16697x) & (!x16693x)) + ((!n_n5251) & (x435x) & (!n_n1139) & (!x16697x) & (x16693x)) + ((!n_n5251) & (x435x) & (!n_n1139) & (x16697x) & (!x16693x)) + ((!n_n5251) & (x435x) & (!n_n1139) & (x16697x) & (x16693x)) + ((!n_n5251) & (x435x) & (n_n1139) & (!x16697x) & (!x16693x)) + ((!n_n5251) & (x435x) & (n_n1139) & (!x16697x) & (x16693x)) + ((!n_n5251) & (x435x) & (n_n1139) & (x16697x) & (!x16693x)) + ((!n_n5251) & (x435x) & (n_n1139) & (x16697x) & (x16693x)) + ((n_n5251) & (!x435x) & (!n_n1139) & (!x16697x) & (!x16693x)) + ((n_n5251) & (!x435x) & (!n_n1139) & (!x16697x) & (x16693x)) + ((n_n5251) & (!x435x) & (!n_n1139) & (x16697x) & (!x16693x)) + ((n_n5251) & (!x435x) & (!n_n1139) & (x16697x) & (x16693x)) + ((n_n5251) & (!x435x) & (n_n1139) & (!x16697x) & (!x16693x)) + ((n_n5251) & (!x435x) & (n_n1139) & (!x16697x) & (x16693x)) + ((n_n5251) & (!x435x) & (n_n1139) & (x16697x) & (!x16693x)) + ((n_n5251) & (!x435x) & (n_n1139) & (x16697x) & (x16693x)) + ((n_n5251) & (x435x) & (!n_n1139) & (!x16697x) & (!x16693x)) + ((n_n5251) & (x435x) & (!n_n1139) & (!x16697x) & (x16693x)) + ((n_n5251) & (x435x) & (!n_n1139) & (x16697x) & (!x16693x)) + ((n_n5251) & (x435x) & (!n_n1139) & (x16697x) & (x16693x)) + ((n_n5251) & (x435x) & (n_n1139) & (!x16697x) & (!x16693x)) + ((n_n5251) & (x435x) & (n_n1139) & (!x16697x) & (x16693x)) + ((n_n5251) & (x435x) & (n_n1139) & (x16697x) & (!x16693x)) + ((n_n5251) & (x435x) & (n_n1139) & (x16697x) & (x16693x)));
	assign x16705x = (((!x358x) & (!x16666x) & (!n_n2205) & (!x125x) & (x16703x)) + ((!x358x) & (!x16666x) & (!n_n2205) & (x125x) & (!x16703x)) + ((!x358x) & (!x16666x) & (!n_n2205) & (x125x) & (x16703x)) + ((!x358x) & (!x16666x) & (n_n2205) & (!x125x) & (!x16703x)) + ((!x358x) & (!x16666x) & (n_n2205) & (!x125x) & (x16703x)) + ((!x358x) & (!x16666x) & (n_n2205) & (x125x) & (!x16703x)) + ((!x358x) & (!x16666x) & (n_n2205) & (x125x) & (x16703x)) + ((!x358x) & (x16666x) & (!n_n2205) & (!x125x) & (!x16703x)) + ((!x358x) & (x16666x) & (!n_n2205) & (!x125x) & (x16703x)) + ((!x358x) & (x16666x) & (!n_n2205) & (x125x) & (!x16703x)) + ((!x358x) & (x16666x) & (!n_n2205) & (x125x) & (x16703x)) + ((!x358x) & (x16666x) & (n_n2205) & (!x125x) & (!x16703x)) + ((!x358x) & (x16666x) & (n_n2205) & (!x125x) & (x16703x)) + ((!x358x) & (x16666x) & (n_n2205) & (x125x) & (!x16703x)) + ((!x358x) & (x16666x) & (n_n2205) & (x125x) & (x16703x)) + ((x358x) & (!x16666x) & (!n_n2205) & (!x125x) & (!x16703x)) + ((x358x) & (!x16666x) & (!n_n2205) & (!x125x) & (x16703x)) + ((x358x) & (!x16666x) & (!n_n2205) & (x125x) & (!x16703x)) + ((x358x) & (!x16666x) & (!n_n2205) & (x125x) & (x16703x)) + ((x358x) & (!x16666x) & (n_n2205) & (!x125x) & (!x16703x)) + ((x358x) & (!x16666x) & (n_n2205) & (!x125x) & (x16703x)) + ((x358x) & (!x16666x) & (n_n2205) & (x125x) & (!x16703x)) + ((x358x) & (!x16666x) & (n_n2205) & (x125x) & (x16703x)) + ((x358x) & (x16666x) & (!n_n2205) & (!x125x) & (!x16703x)) + ((x358x) & (x16666x) & (!n_n2205) & (!x125x) & (x16703x)) + ((x358x) & (x16666x) & (!n_n2205) & (x125x) & (!x16703x)) + ((x358x) & (x16666x) & (!n_n2205) & (x125x) & (x16703x)) + ((x358x) & (x16666x) & (n_n2205) & (!x125x) & (!x16703x)) + ((x358x) & (x16666x) & (n_n2205) & (!x125x) & (x16703x)) + ((x358x) & (x16666x) & (n_n2205) & (x125x) & (!x16703x)) + ((x358x) & (x16666x) & (n_n2205) & (x125x) & (x16703x)));
	assign n_n2168 = (((!x16758x) & (!n_n2196) & (x16757x)) + ((!x16758x) & (n_n2196) & (!x16757x)) + ((!x16758x) & (n_n2196) & (x16757x)) + ((x16758x) & (!n_n2196) & (!x16757x)) + ((x16758x) & (!n_n2196) & (x16757x)) + ((x16758x) & (n_n2196) & (!x16757x)) + ((x16758x) & (n_n2196) & (x16757x)));
	assign x16762x = (((!x117x) & (!x462x) & (!x16659x) & (!x16660x) & (x16761x)) + ((!x117x) & (!x462x) & (!x16659x) & (x16660x) & (!x16761x)) + ((!x117x) & (!x462x) & (!x16659x) & (x16660x) & (x16761x)) + ((!x117x) & (!x462x) & (x16659x) & (!x16660x) & (!x16761x)) + ((!x117x) & (!x462x) & (x16659x) & (!x16660x) & (x16761x)) + ((!x117x) & (!x462x) & (x16659x) & (x16660x) & (!x16761x)) + ((!x117x) & (!x462x) & (x16659x) & (x16660x) & (x16761x)) + ((!x117x) & (x462x) & (!x16659x) & (!x16660x) & (!x16761x)) + ((!x117x) & (x462x) & (!x16659x) & (!x16660x) & (x16761x)) + ((!x117x) & (x462x) & (!x16659x) & (x16660x) & (!x16761x)) + ((!x117x) & (x462x) & (!x16659x) & (x16660x) & (x16761x)) + ((!x117x) & (x462x) & (x16659x) & (!x16660x) & (!x16761x)) + ((!x117x) & (x462x) & (x16659x) & (!x16660x) & (x16761x)) + ((!x117x) & (x462x) & (x16659x) & (x16660x) & (!x16761x)) + ((!x117x) & (x462x) & (x16659x) & (x16660x) & (x16761x)) + ((x117x) & (!x462x) & (!x16659x) & (!x16660x) & (!x16761x)) + ((x117x) & (!x462x) & (!x16659x) & (!x16660x) & (x16761x)) + ((x117x) & (!x462x) & (!x16659x) & (x16660x) & (!x16761x)) + ((x117x) & (!x462x) & (!x16659x) & (x16660x) & (x16761x)) + ((x117x) & (!x462x) & (x16659x) & (!x16660x) & (!x16761x)) + ((x117x) & (!x462x) & (x16659x) & (!x16660x) & (x16761x)) + ((x117x) & (!x462x) & (x16659x) & (x16660x) & (!x16761x)) + ((x117x) & (!x462x) & (x16659x) & (x16660x) & (x16761x)) + ((x117x) & (x462x) & (!x16659x) & (!x16660x) & (!x16761x)) + ((x117x) & (x462x) & (!x16659x) & (!x16660x) & (x16761x)) + ((x117x) & (x462x) & (!x16659x) & (x16660x) & (!x16761x)) + ((x117x) & (x462x) & (!x16659x) & (x16660x) & (x16761x)) + ((x117x) & (x462x) & (x16659x) & (!x16660x) & (!x16761x)) + ((x117x) & (x462x) & (x16659x) & (!x16660x) & (x16761x)) + ((x117x) & (x462x) & (x16659x) & (x16660x) & (!x16761x)) + ((x117x) & (x462x) & (x16659x) & (x16660x) & (x16761x)));
	assign n_n4432 = (((i_9_) & (n_n536) & (n_n526) & (n_n464)));
	assign n_n4438 = (((i_9_) & (n_n536) & (n_n520) & (n_n464)));
	assign n_n4461 = (((!i_9_) & (n_n518) & (n_n455) & (n_n530)));
	assign n_n4421 = (((i_1_) & (i_2_) & (i_0_) & (n_n473) & (x20x)));
	assign x16769x = (((!n_n4432) & (!n_n4438) & (!n_n4461) & (n_n4421)) + ((!n_n4432) & (!n_n4438) & (n_n4461) & (!n_n4421)) + ((!n_n4432) & (!n_n4438) & (n_n4461) & (n_n4421)) + ((!n_n4432) & (n_n4438) & (!n_n4461) & (!n_n4421)) + ((!n_n4432) & (n_n4438) & (!n_n4461) & (n_n4421)) + ((!n_n4432) & (n_n4438) & (n_n4461) & (!n_n4421)) + ((!n_n4432) & (n_n4438) & (n_n4461) & (n_n4421)) + ((n_n4432) & (!n_n4438) & (!n_n4461) & (!n_n4421)) + ((n_n4432) & (!n_n4438) & (!n_n4461) & (n_n4421)) + ((n_n4432) & (!n_n4438) & (n_n4461) & (!n_n4421)) + ((n_n4432) & (!n_n4438) & (n_n4461) & (n_n4421)) + ((n_n4432) & (n_n4438) & (!n_n4461) & (!n_n4421)) + ((n_n4432) & (n_n4438) & (!n_n4461) & (n_n4421)) + ((n_n4432) & (n_n4438) & (n_n4461) & (!n_n4421)) + ((n_n4432) & (n_n4438) & (n_n4461) & (n_n4421)));
	assign x84x = (((!i_9_) & (n_n536) & (n_n532) & (n_n464)) + ((i_9_) & (n_n536) & (n_n532) & (n_n464)));
	assign n_n4465 = (((!i_9_) & (n_n518) & (n_n526) & (n_n455)));
	assign n_n4443 = (((!i_9_) & (n_n455) & (n_n532) & (n_n535)));
	assign n_n4429 = (((!i_9_) & (n_n536) & (n_n530) & (n_n464)));
	assign n_n2103 = (((!x16769x) & (!x84x) & (!n_n4465) & (!n_n4443) & (n_n4429)) + ((!x16769x) & (!x84x) & (!n_n4465) & (n_n4443) & (!n_n4429)) + ((!x16769x) & (!x84x) & (!n_n4465) & (n_n4443) & (n_n4429)) + ((!x16769x) & (!x84x) & (n_n4465) & (!n_n4443) & (!n_n4429)) + ((!x16769x) & (!x84x) & (n_n4465) & (!n_n4443) & (n_n4429)) + ((!x16769x) & (!x84x) & (n_n4465) & (n_n4443) & (!n_n4429)) + ((!x16769x) & (!x84x) & (n_n4465) & (n_n4443) & (n_n4429)) + ((!x16769x) & (x84x) & (!n_n4465) & (!n_n4443) & (!n_n4429)) + ((!x16769x) & (x84x) & (!n_n4465) & (!n_n4443) & (n_n4429)) + ((!x16769x) & (x84x) & (!n_n4465) & (n_n4443) & (!n_n4429)) + ((!x16769x) & (x84x) & (!n_n4465) & (n_n4443) & (n_n4429)) + ((!x16769x) & (x84x) & (n_n4465) & (!n_n4443) & (!n_n4429)) + ((!x16769x) & (x84x) & (n_n4465) & (!n_n4443) & (n_n4429)) + ((!x16769x) & (x84x) & (n_n4465) & (n_n4443) & (!n_n4429)) + ((!x16769x) & (x84x) & (n_n4465) & (n_n4443) & (n_n4429)) + ((x16769x) & (!x84x) & (!n_n4465) & (!n_n4443) & (!n_n4429)) + ((x16769x) & (!x84x) & (!n_n4465) & (!n_n4443) & (n_n4429)) + ((x16769x) & (!x84x) & (!n_n4465) & (n_n4443) & (!n_n4429)) + ((x16769x) & (!x84x) & (!n_n4465) & (n_n4443) & (n_n4429)) + ((x16769x) & (!x84x) & (n_n4465) & (!n_n4443) & (!n_n4429)) + ((x16769x) & (!x84x) & (n_n4465) & (!n_n4443) & (n_n4429)) + ((x16769x) & (!x84x) & (n_n4465) & (n_n4443) & (!n_n4429)) + ((x16769x) & (!x84x) & (n_n4465) & (n_n4443) & (n_n4429)) + ((x16769x) & (x84x) & (!n_n4465) & (!n_n4443) & (!n_n4429)) + ((x16769x) & (x84x) & (!n_n4465) & (!n_n4443) & (n_n4429)) + ((x16769x) & (x84x) & (!n_n4465) & (n_n4443) & (!n_n4429)) + ((x16769x) & (x84x) & (!n_n4465) & (n_n4443) & (n_n4429)) + ((x16769x) & (x84x) & (n_n4465) & (!n_n4443) & (!n_n4429)) + ((x16769x) & (x84x) & (n_n4465) & (!n_n4443) & (n_n4429)) + ((x16769x) & (x84x) & (n_n4465) & (n_n4443) & (!n_n4429)) + ((x16769x) & (x84x) & (n_n4465) & (n_n4443) & (n_n4429)));
	assign x16790x = (((!n_n5034) & (!n_n5099) & (!n_n5019) & (n_n5097)) + ((!n_n5034) & (!n_n5099) & (n_n5019) & (!n_n5097)) + ((!n_n5034) & (!n_n5099) & (n_n5019) & (n_n5097)) + ((!n_n5034) & (n_n5099) & (!n_n5019) & (!n_n5097)) + ((!n_n5034) & (n_n5099) & (!n_n5019) & (n_n5097)) + ((!n_n5034) & (n_n5099) & (n_n5019) & (!n_n5097)) + ((!n_n5034) & (n_n5099) & (n_n5019) & (n_n5097)) + ((n_n5034) & (!n_n5099) & (!n_n5019) & (!n_n5097)) + ((n_n5034) & (!n_n5099) & (!n_n5019) & (n_n5097)) + ((n_n5034) & (!n_n5099) & (n_n5019) & (!n_n5097)) + ((n_n5034) & (!n_n5099) & (n_n5019) & (n_n5097)) + ((n_n5034) & (n_n5099) & (!n_n5019) & (!n_n5097)) + ((n_n5034) & (n_n5099) & (!n_n5019) & (n_n5097)) + ((n_n5034) & (n_n5099) & (n_n5019) & (!n_n5097)) + ((n_n5034) & (n_n5099) & (n_n5019) & (n_n5097)));
	assign x16791x = (((!n_n5104) & (!n_n5106) & (!n_n5117) & (!n_n5121) & (n_n5122)) + ((!n_n5104) & (!n_n5106) & (!n_n5117) & (n_n5121) & (!n_n5122)) + ((!n_n5104) & (!n_n5106) & (!n_n5117) & (n_n5121) & (n_n5122)) + ((!n_n5104) & (!n_n5106) & (n_n5117) & (!n_n5121) & (!n_n5122)) + ((!n_n5104) & (!n_n5106) & (n_n5117) & (!n_n5121) & (n_n5122)) + ((!n_n5104) & (!n_n5106) & (n_n5117) & (n_n5121) & (!n_n5122)) + ((!n_n5104) & (!n_n5106) & (n_n5117) & (n_n5121) & (n_n5122)) + ((!n_n5104) & (n_n5106) & (!n_n5117) & (!n_n5121) & (!n_n5122)) + ((!n_n5104) & (n_n5106) & (!n_n5117) & (!n_n5121) & (n_n5122)) + ((!n_n5104) & (n_n5106) & (!n_n5117) & (n_n5121) & (!n_n5122)) + ((!n_n5104) & (n_n5106) & (!n_n5117) & (n_n5121) & (n_n5122)) + ((!n_n5104) & (n_n5106) & (n_n5117) & (!n_n5121) & (!n_n5122)) + ((!n_n5104) & (n_n5106) & (n_n5117) & (!n_n5121) & (n_n5122)) + ((!n_n5104) & (n_n5106) & (n_n5117) & (n_n5121) & (!n_n5122)) + ((!n_n5104) & (n_n5106) & (n_n5117) & (n_n5121) & (n_n5122)) + ((n_n5104) & (!n_n5106) & (!n_n5117) & (!n_n5121) & (!n_n5122)) + ((n_n5104) & (!n_n5106) & (!n_n5117) & (!n_n5121) & (n_n5122)) + ((n_n5104) & (!n_n5106) & (!n_n5117) & (n_n5121) & (!n_n5122)) + ((n_n5104) & (!n_n5106) & (!n_n5117) & (n_n5121) & (n_n5122)) + ((n_n5104) & (!n_n5106) & (n_n5117) & (!n_n5121) & (!n_n5122)) + ((n_n5104) & (!n_n5106) & (n_n5117) & (!n_n5121) & (n_n5122)) + ((n_n5104) & (!n_n5106) & (n_n5117) & (n_n5121) & (!n_n5122)) + ((n_n5104) & (!n_n5106) & (n_n5117) & (n_n5121) & (n_n5122)) + ((n_n5104) & (n_n5106) & (!n_n5117) & (!n_n5121) & (!n_n5122)) + ((n_n5104) & (n_n5106) & (!n_n5117) & (!n_n5121) & (n_n5122)) + ((n_n5104) & (n_n5106) & (!n_n5117) & (n_n5121) & (!n_n5122)) + ((n_n5104) & (n_n5106) & (!n_n5117) & (n_n5121) & (n_n5122)) + ((n_n5104) & (n_n5106) & (n_n5117) & (!n_n5121) & (!n_n5122)) + ((n_n5104) & (n_n5106) & (n_n5117) & (!n_n5121) & (n_n5122)) + ((n_n5104) & (n_n5106) & (n_n5117) & (n_n5121) & (!n_n5122)) + ((n_n5104) & (n_n5106) & (n_n5117) & (n_n5121) & (n_n5122)));
	assign x16796x = (((!n_n5123) & (!n_n5131) & (!n_n5137) & (n_n5146)) + ((!n_n5123) & (!n_n5131) & (n_n5137) & (!n_n5146)) + ((!n_n5123) & (!n_n5131) & (n_n5137) & (n_n5146)) + ((!n_n5123) & (n_n5131) & (!n_n5137) & (!n_n5146)) + ((!n_n5123) & (n_n5131) & (!n_n5137) & (n_n5146)) + ((!n_n5123) & (n_n5131) & (n_n5137) & (!n_n5146)) + ((!n_n5123) & (n_n5131) & (n_n5137) & (n_n5146)) + ((n_n5123) & (!n_n5131) & (!n_n5137) & (!n_n5146)) + ((n_n5123) & (!n_n5131) & (!n_n5137) & (n_n5146)) + ((n_n5123) & (!n_n5131) & (n_n5137) & (!n_n5146)) + ((n_n5123) & (!n_n5131) & (n_n5137) & (n_n5146)) + ((n_n5123) & (n_n5131) & (!n_n5137) & (!n_n5146)) + ((n_n5123) & (n_n5131) & (!n_n5137) & (n_n5146)) + ((n_n5123) & (n_n5131) & (n_n5137) & (!n_n5146)) + ((n_n5123) & (n_n5131) & (n_n5137) & (n_n5146)));
	assign x16797x = (((!n_n5193) & (!n_n5182) & (!n_n5168) & (x126x)) + ((!n_n5193) & (!n_n5182) & (n_n5168) & (!x126x)) + ((!n_n5193) & (!n_n5182) & (n_n5168) & (x126x)) + ((!n_n5193) & (n_n5182) & (!n_n5168) & (!x126x)) + ((!n_n5193) & (n_n5182) & (!n_n5168) & (x126x)) + ((!n_n5193) & (n_n5182) & (n_n5168) & (!x126x)) + ((!n_n5193) & (n_n5182) & (n_n5168) & (x126x)) + ((n_n5193) & (!n_n5182) & (!n_n5168) & (!x126x)) + ((n_n5193) & (!n_n5182) & (!n_n5168) & (x126x)) + ((n_n5193) & (!n_n5182) & (n_n5168) & (!x126x)) + ((n_n5193) & (!n_n5182) & (n_n5168) & (x126x)) + ((n_n5193) & (n_n5182) & (!n_n5168) & (!x126x)) + ((n_n5193) & (n_n5182) & (!n_n5168) & (x126x)) + ((n_n5193) & (n_n5182) & (n_n5168) & (!x126x)) + ((n_n5193) & (n_n5182) & (n_n5168) & (x126x)));
	assign x16805x = (((!n_n4996) & (!n_n4992) & (!n_n4981) & (!n_n5005) & (x16804x)) + ((!n_n4996) & (!n_n4992) & (!n_n4981) & (n_n5005) & (!x16804x)) + ((!n_n4996) & (!n_n4992) & (!n_n4981) & (n_n5005) & (x16804x)) + ((!n_n4996) & (!n_n4992) & (n_n4981) & (!n_n5005) & (!x16804x)) + ((!n_n4996) & (!n_n4992) & (n_n4981) & (!n_n5005) & (x16804x)) + ((!n_n4996) & (!n_n4992) & (n_n4981) & (n_n5005) & (!x16804x)) + ((!n_n4996) & (!n_n4992) & (n_n4981) & (n_n5005) & (x16804x)) + ((!n_n4996) & (n_n4992) & (!n_n4981) & (!n_n5005) & (!x16804x)) + ((!n_n4996) & (n_n4992) & (!n_n4981) & (!n_n5005) & (x16804x)) + ((!n_n4996) & (n_n4992) & (!n_n4981) & (n_n5005) & (!x16804x)) + ((!n_n4996) & (n_n4992) & (!n_n4981) & (n_n5005) & (x16804x)) + ((!n_n4996) & (n_n4992) & (n_n4981) & (!n_n5005) & (!x16804x)) + ((!n_n4996) & (n_n4992) & (n_n4981) & (!n_n5005) & (x16804x)) + ((!n_n4996) & (n_n4992) & (n_n4981) & (n_n5005) & (!x16804x)) + ((!n_n4996) & (n_n4992) & (n_n4981) & (n_n5005) & (x16804x)) + ((n_n4996) & (!n_n4992) & (!n_n4981) & (!n_n5005) & (!x16804x)) + ((n_n4996) & (!n_n4992) & (!n_n4981) & (!n_n5005) & (x16804x)) + ((n_n4996) & (!n_n4992) & (!n_n4981) & (n_n5005) & (!x16804x)) + ((n_n4996) & (!n_n4992) & (!n_n4981) & (n_n5005) & (x16804x)) + ((n_n4996) & (!n_n4992) & (n_n4981) & (!n_n5005) & (!x16804x)) + ((n_n4996) & (!n_n4992) & (n_n4981) & (!n_n5005) & (x16804x)) + ((n_n4996) & (!n_n4992) & (n_n4981) & (n_n5005) & (!x16804x)) + ((n_n4996) & (!n_n4992) & (n_n4981) & (n_n5005) & (x16804x)) + ((n_n4996) & (n_n4992) & (!n_n4981) & (!n_n5005) & (!x16804x)) + ((n_n4996) & (n_n4992) & (!n_n4981) & (!n_n5005) & (x16804x)) + ((n_n4996) & (n_n4992) & (!n_n4981) & (n_n5005) & (!x16804x)) + ((n_n4996) & (n_n4992) & (!n_n4981) & (n_n5005) & (x16804x)) + ((n_n4996) & (n_n4992) & (n_n4981) & (!n_n5005) & (!x16804x)) + ((n_n4996) & (n_n4992) & (n_n4981) & (!n_n5005) & (x16804x)) + ((n_n4996) & (n_n4992) & (n_n4981) & (n_n5005) & (!x16804x)) + ((n_n4996) & (n_n4992) & (n_n4981) & (n_n5005) & (x16804x)));
	assign n_n2084 = (((!x16790x) & (!x16791x) & (!x16796x) & (!x16797x) & (x16805x)) + ((!x16790x) & (!x16791x) & (!x16796x) & (x16797x) & (!x16805x)) + ((!x16790x) & (!x16791x) & (!x16796x) & (x16797x) & (x16805x)) + ((!x16790x) & (!x16791x) & (x16796x) & (!x16797x) & (!x16805x)) + ((!x16790x) & (!x16791x) & (x16796x) & (!x16797x) & (x16805x)) + ((!x16790x) & (!x16791x) & (x16796x) & (x16797x) & (!x16805x)) + ((!x16790x) & (!x16791x) & (x16796x) & (x16797x) & (x16805x)) + ((!x16790x) & (x16791x) & (!x16796x) & (!x16797x) & (!x16805x)) + ((!x16790x) & (x16791x) & (!x16796x) & (!x16797x) & (x16805x)) + ((!x16790x) & (x16791x) & (!x16796x) & (x16797x) & (!x16805x)) + ((!x16790x) & (x16791x) & (!x16796x) & (x16797x) & (x16805x)) + ((!x16790x) & (x16791x) & (x16796x) & (!x16797x) & (!x16805x)) + ((!x16790x) & (x16791x) & (x16796x) & (!x16797x) & (x16805x)) + ((!x16790x) & (x16791x) & (x16796x) & (x16797x) & (!x16805x)) + ((!x16790x) & (x16791x) & (x16796x) & (x16797x) & (x16805x)) + ((x16790x) & (!x16791x) & (!x16796x) & (!x16797x) & (!x16805x)) + ((x16790x) & (!x16791x) & (!x16796x) & (!x16797x) & (x16805x)) + ((x16790x) & (!x16791x) & (!x16796x) & (x16797x) & (!x16805x)) + ((x16790x) & (!x16791x) & (!x16796x) & (x16797x) & (x16805x)) + ((x16790x) & (!x16791x) & (x16796x) & (!x16797x) & (!x16805x)) + ((x16790x) & (!x16791x) & (x16796x) & (!x16797x) & (x16805x)) + ((x16790x) & (!x16791x) & (x16796x) & (x16797x) & (!x16805x)) + ((x16790x) & (!x16791x) & (x16796x) & (x16797x) & (x16805x)) + ((x16790x) & (x16791x) & (!x16796x) & (!x16797x) & (!x16805x)) + ((x16790x) & (x16791x) & (!x16796x) & (!x16797x) & (x16805x)) + ((x16790x) & (x16791x) & (!x16796x) & (x16797x) & (!x16805x)) + ((x16790x) & (x16791x) & (!x16796x) & (x16797x) & (x16805x)) + ((x16790x) & (x16791x) & (x16796x) & (!x16797x) & (!x16805x)) + ((x16790x) & (x16791x) & (x16796x) & (!x16797x) & (x16805x)) + ((x16790x) & (x16791x) & (x16796x) & (x16797x) & (!x16805x)) + ((x16790x) & (x16791x) & (x16796x) & (x16797x) & (x16805x)));
	assign n_n536 = (((i_1_) & (i_2_) & (i_0_)));
	assign n_n518 = (((!i_5_) & (i_3_) & (i_4_)));
	assign x21x = (((!i_9_) & (i_7_) & (!i_8_) & (!i_6_)));
	assign n_n4337 = (((!i_9_) & (n_n536) & (n_n518) & (n_n526)));
	assign n_n4403 = (((!i_9_) & (n_n536) & (n_n524) & (n_n482)));
	assign n_n455 = (((i_1_) & (!i_2_) & (i_0_)));
	assign x13x = (((i_9_) & (i_1_) & (!i_2_) & (i_0_)));
	assign n_n4464 = (((i_9_) & (n_n518) & (n_n526) & (n_n455)));
	assign n_n4467 = (((!i_9_) & (n_n524) & (n_n518) & (n_n455)));
	assign n_n528 = (((!i_7_) & (!i_8_) & (i_6_)));
	assign x11x = (((!i_9_) & (!i_7_) & (!i_8_) & (i_6_)));
	assign n_n4463 = (((!i_9_) & (n_n518) & (n_n455) & (n_n528)));
	assign n_n390 = (((!i_1_) & (i_2_) & (i_0_)));
	assign x10x = (((i_9_) & (!i_1_) & (i_2_) & (i_0_)));
	assign n_n532 = (((i_7_) & (!i_8_) & (i_6_)));
	assign n_n4666 = (((i_9_) & (n_n390) & (n_n473) & (n_n532)));
	assign n_n4667 = (((!i_9_) & (n_n390) & (n_n473) & (n_n532)));
	assign n_n4664 = (((i_9_) & (n_n390) & (n_n473) & (n_n534)));
	assign n_n509 = (((i_5_) & (i_3_) & (!i_4_)));
	assign n_n325 = (((!i_1_) & (!i_2_) & (i_0_)));
	assign x483x = (((i_5_) & (i_3_) & (!i_4_) & (n_n325)));
	assign n_n4737 = (((!i_9_) & (n_n526) & (n_n509) & (n_n325)));
	assign x14x = (((i_9_) & (!i_1_) & (!i_2_) & (i_0_)));
	assign n_n4738 = (((i_9_) & (n_n524) & (n_n509) & (n_n325)));
	assign n_n4735 = (((!i_9_) & (n_n528) & (n_n509) & (n_n325)));
	assign n_n4782 = (((i_9_) & (n_n482) & (n_n528) & (n_n325)));
	assign n_n4784 = (((i_9_) & (n_n526) & (n_n482) & (n_n325)));
	assign n_n4779 = (((!i_9_) & (n_n482) & (n_n532) & (n_n325)));
	assign n_n260 = (((i_1_) & (i_2_) & (!i_0_)));
	assign x17x = (((i_9_) & (i_1_) & (i_2_) & (!i_0_)));
	assign n_n535 = (((i_5_) & (i_3_) & (i_4_)));
	assign n_n4830 = (((i_9_) & (n_n528) & (n_n260) & (n_n535)));
	assign x552x = (((i_1_) & (i_2_) & (!i_0_) & (n_n535)));
	assign n_n4831 = (((!i_9_) & (n_n528) & (n_n260) & (n_n535)));
	assign n_n4900 = (((i_9_) & (n_n260) & (n_n522) & (n_n491)));
	assign n_n4902 = (((i_9_) & (n_n260) & (n_n491) & (n_n520)));
	assign n_n4898 = (((i_9_) & (n_n524) & (n_n260) & (n_n491)));
	assign n_n195 = (((i_1_) & (!i_2_) & (!i_0_)));
	assign x18x = (((i_9_) & (i_1_) & (!i_2_) & (!i_0_)));
	assign n_n4976 = (((i_9_) & (n_n518) & (n_n526) & (n_n195)));
	assign n_n4977 = (((!i_9_) & (n_n518) & (n_n526) & (n_n195)));
	assign n_n4975 = (((!i_9_) & (n_n518) & (n_n528) & (n_n195)));
	assign n_n5038 = (((i_9_) & (n_n482) & (n_n528) & (n_n195)));
	assign n_n5040 = (((i_9_) & (n_n526) & (n_n482) & (n_n195)));
	assign n_n5034 = (((i_9_) & (n_n482) & (n_n532) & (n_n195)));
	assign n_n130 = (((!i_1_) & (i_2_) & (!i_0_)));
	assign x12x = (((i_9_) & (!i_1_) & (i_2_) & (!i_0_)));
	assign n_n5092 = (((i_5_) & (i_3_) & (i_4_) & (n_n522) & (x12x)));
	assign n_n5093 = (((i_5_) & (i_3_) & (i_4_) & (n_n130) & (x20x)));
	assign n_n5091 = (((!i_9_) & (n_n524) & (n_n535) & (n_n130)));
	assign n_n4148 = (((!i_9_) & (!n_n524) & (n_n535) & (n_n522) & (n_n130)) + ((!i_9_) & (n_n524) & (n_n535) & (!n_n522) & (n_n130)) + ((!i_9_) & (n_n524) & (n_n535) & (n_n522) & (n_n130)) + ((i_9_) & (!n_n524) & (n_n535) & (n_n522) & (n_n130)) + ((i_9_) & (n_n524) & (n_n535) & (n_n522) & (n_n130)));
	assign n_n4440 = (((i_9_) & (n_n455) & (n_n534) & (n_n535)));
	assign x516x = (((i_7_) & (!i_8_) & (!i_6_) & (n_n464)));
	assign n_n4434 = (((i_9_) & (n_n536) & (n_n524) & (n_n464)));
	assign n_n4433 = (((!i_9_) & (n_n536) & (n_n526) & (n_n464)));
	assign x98x = (((!i_9_) & (n_n536) & (!n_n526) & (n_n528) & (n_n464)) + ((!i_9_) & (n_n536) & (n_n526) & (!n_n528) & (n_n464)) + ((!i_9_) & (n_n536) & (n_n526) & (n_n528) & (n_n464)));
	assign x23x = (((!i_9_) & (!i_7_) & (!i_8_) & (!i_6_)));
	assign x233x = (((!i_9_) & (n_n536) & (!n_n520) & (x23x) & (n_n464)) + ((!i_9_) & (n_n536) & (n_n520) & (x23x) & (n_n464)) + ((i_9_) & (n_n536) & (!n_n520) & (x23x) & (n_n464)) + ((i_9_) & (n_n536) & (n_n520) & (!x23x) & (n_n464)) + ((i_9_) & (n_n536) & (n_n520) & (x23x) & (n_n464)));
	assign x236x = (((!i_9_) & (n_n536) & (!n_n522) & (x20x) & (n_n464)) + ((!i_9_) & (n_n536) & (n_n522) & (x20x) & (n_n464)) + ((i_9_) & (n_n536) & (!n_n522) & (x20x) & (n_n464)) + ((i_9_) & (n_n536) & (n_n522) & (!x20x) & (n_n464)) + ((i_9_) & (n_n536) & (n_n522) & (x20x) & (n_n464)));
	assign x13428x = (((!n_n536) & (!n_n4438) & (x236x) & (!x23x) & (!n_n464)) + ((!n_n536) & (!n_n4438) & (x236x) & (!x23x) & (n_n464)) + ((!n_n536) & (!n_n4438) & (x236x) & (x23x) & (!n_n464)) + ((!n_n536) & (!n_n4438) & (x236x) & (x23x) & (n_n464)) + ((!n_n536) & (n_n4438) & (!x236x) & (!x23x) & (!n_n464)) + ((!n_n536) & (n_n4438) & (!x236x) & (!x23x) & (n_n464)) + ((!n_n536) & (n_n4438) & (!x236x) & (x23x) & (!n_n464)) + ((!n_n536) & (n_n4438) & (!x236x) & (x23x) & (n_n464)) + ((!n_n536) & (n_n4438) & (x236x) & (!x23x) & (!n_n464)) + ((!n_n536) & (n_n4438) & (x236x) & (!x23x) & (n_n464)) + ((!n_n536) & (n_n4438) & (x236x) & (x23x) & (!n_n464)) + ((!n_n536) & (n_n4438) & (x236x) & (x23x) & (n_n464)) + ((n_n536) & (!n_n4438) & (!x236x) & (x23x) & (n_n464)) + ((n_n536) & (!n_n4438) & (x236x) & (!x23x) & (!n_n464)) + ((n_n536) & (!n_n4438) & (x236x) & (!x23x) & (n_n464)) + ((n_n536) & (!n_n4438) & (x236x) & (x23x) & (!n_n464)) + ((n_n536) & (!n_n4438) & (x236x) & (x23x) & (n_n464)) + ((n_n536) & (n_n4438) & (!x236x) & (!x23x) & (!n_n464)) + ((n_n536) & (n_n4438) & (!x236x) & (!x23x) & (n_n464)) + ((n_n536) & (n_n4438) & (!x236x) & (x23x) & (!n_n464)) + ((n_n536) & (n_n4438) & (!x236x) & (x23x) & (n_n464)) + ((n_n536) & (n_n4438) & (x236x) & (!x23x) & (!n_n464)) + ((n_n536) & (n_n4438) & (x236x) & (!x23x) & (n_n464)) + ((n_n536) & (n_n4438) & (x236x) & (x23x) & (!n_n464)) + ((n_n536) & (n_n4438) & (x236x) & (x23x) & (n_n464)));
	assign n_n4095 = (((!n_n4440) & (!n_n4434) & (!n_n4432) & (!x98x) & (x13428x)) + ((!n_n4440) & (!n_n4434) & (!n_n4432) & (x98x) & (!x13428x)) + ((!n_n4440) & (!n_n4434) & (!n_n4432) & (x98x) & (x13428x)) + ((!n_n4440) & (!n_n4434) & (n_n4432) & (!x98x) & (!x13428x)) + ((!n_n4440) & (!n_n4434) & (n_n4432) & (!x98x) & (x13428x)) + ((!n_n4440) & (!n_n4434) & (n_n4432) & (x98x) & (!x13428x)) + ((!n_n4440) & (!n_n4434) & (n_n4432) & (x98x) & (x13428x)) + ((!n_n4440) & (n_n4434) & (!n_n4432) & (!x98x) & (!x13428x)) + ((!n_n4440) & (n_n4434) & (!n_n4432) & (!x98x) & (x13428x)) + ((!n_n4440) & (n_n4434) & (!n_n4432) & (x98x) & (!x13428x)) + ((!n_n4440) & (n_n4434) & (!n_n4432) & (x98x) & (x13428x)) + ((!n_n4440) & (n_n4434) & (n_n4432) & (!x98x) & (!x13428x)) + ((!n_n4440) & (n_n4434) & (n_n4432) & (!x98x) & (x13428x)) + ((!n_n4440) & (n_n4434) & (n_n4432) & (x98x) & (!x13428x)) + ((!n_n4440) & (n_n4434) & (n_n4432) & (x98x) & (x13428x)) + ((n_n4440) & (!n_n4434) & (!n_n4432) & (!x98x) & (!x13428x)) + ((n_n4440) & (!n_n4434) & (!n_n4432) & (!x98x) & (x13428x)) + ((n_n4440) & (!n_n4434) & (!n_n4432) & (x98x) & (!x13428x)) + ((n_n4440) & (!n_n4434) & (!n_n4432) & (x98x) & (x13428x)) + ((n_n4440) & (!n_n4434) & (n_n4432) & (!x98x) & (!x13428x)) + ((n_n4440) & (!n_n4434) & (n_n4432) & (!x98x) & (x13428x)) + ((n_n4440) & (!n_n4434) & (n_n4432) & (x98x) & (!x13428x)) + ((n_n4440) & (!n_n4434) & (n_n4432) & (x98x) & (x13428x)) + ((n_n4440) & (n_n4434) & (!n_n4432) & (!x98x) & (!x13428x)) + ((n_n4440) & (n_n4434) & (!n_n4432) & (!x98x) & (x13428x)) + ((n_n4440) & (n_n4434) & (!n_n4432) & (x98x) & (!x13428x)) + ((n_n4440) & (n_n4434) & (!n_n4432) & (x98x) & (x13428x)) + ((n_n4440) & (n_n4434) & (n_n4432) & (!x98x) & (!x13428x)) + ((n_n4440) & (n_n4434) & (n_n4432) & (!x98x) & (x13428x)) + ((n_n4440) & (n_n4434) & (n_n4432) & (x98x) & (!x13428x)) + ((n_n4440) & (n_n4434) & (n_n4432) & (x98x) & (x13428x)));
	assign n_n4720 = (((i_9_) & (n_n518) & (n_n526) & (n_n325)));
	assign n_n4717 = (((!i_9_) & (n_n518) & (n_n325) & (n_n530)));
	assign x241x = (((!i_9_) & (n_n518) & (!n_n528) & (n_n325) & (n_n530)) + ((!i_9_) & (n_n518) & (n_n528) & (n_n325) & (n_n530)) + ((i_9_) & (n_n518) & (n_n528) & (n_n325) & (!n_n530)) + ((i_9_) & (n_n518) & (n_n528) & (n_n325) & (n_n530)));
	assign n_n4857 = (((!i_9_) & (n_n534) & (n_n509) & (n_n260)));
	assign n_n4862 = (((i_9_) & (n_n528) & (n_n509) & (n_n260)));
	assign n_n4856 = (((i_9_) & (n_n534) & (n_n509) & (n_n260)));
	assign n_n4863 = (((!i_9_) & (n_n528) & (n_n509) & (n_n260)));
	assign n_n4865 = (((!i_9_) & (n_n526) & (n_n509) & (n_n260)));
	assign x40x = (((!i_9_) & (!n_n526) & (n_n528) & (n_n509) & (n_n260)) + ((!i_9_) & (n_n526) & (!n_n528) & (n_n509) & (n_n260)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n509) & (n_n260)));
	assign n_n4854 = (((i_9_) & (n_n518) & (n_n260) & (n_n520)));
	assign n_n4855 = (((!i_5_) & (i_3_) & (i_4_) & (n_n260) & (x23x)));
	assign x102x = (((!i_9_) & (n_n518) & (n_n260) & (!n_n520) & (x23x)) + ((!i_9_) & (n_n518) & (n_n260) & (n_n520) & (x23x)) + ((i_9_) & (n_n518) & (n_n260) & (!n_n520) & (x23x)) + ((i_9_) & (n_n518) & (n_n260) & (n_n520) & (!x23x)) + ((i_9_) & (n_n518) & (n_n260) & (n_n520) & (x23x)));
	assign n_n4859 = (((!i_9_) & (n_n532) & (n_n509) & (n_n260)));
	assign n_n4858 = (((i_9_) & (n_n532) & (n_n509) & (n_n260)));
	assign x245x = (((!i_9_) & (n_n532) & (n_n509) & (n_n260)) + ((i_9_) & (n_n532) & (n_n509) & (n_n260)));
	assign x13171x = (((!n_n4857) & (!n_n4862) & (!n_n4856) & (!n_n4863) & (n_n4865)) + ((!n_n4857) & (!n_n4862) & (!n_n4856) & (n_n4863) & (!n_n4865)) + ((!n_n4857) & (!n_n4862) & (!n_n4856) & (n_n4863) & (n_n4865)) + ((!n_n4857) & (!n_n4862) & (n_n4856) & (!n_n4863) & (!n_n4865)) + ((!n_n4857) & (!n_n4862) & (n_n4856) & (!n_n4863) & (n_n4865)) + ((!n_n4857) & (!n_n4862) & (n_n4856) & (n_n4863) & (!n_n4865)) + ((!n_n4857) & (!n_n4862) & (n_n4856) & (n_n4863) & (n_n4865)) + ((!n_n4857) & (n_n4862) & (!n_n4856) & (!n_n4863) & (!n_n4865)) + ((!n_n4857) & (n_n4862) & (!n_n4856) & (!n_n4863) & (n_n4865)) + ((!n_n4857) & (n_n4862) & (!n_n4856) & (n_n4863) & (!n_n4865)) + ((!n_n4857) & (n_n4862) & (!n_n4856) & (n_n4863) & (n_n4865)) + ((!n_n4857) & (n_n4862) & (n_n4856) & (!n_n4863) & (!n_n4865)) + ((!n_n4857) & (n_n4862) & (n_n4856) & (!n_n4863) & (n_n4865)) + ((!n_n4857) & (n_n4862) & (n_n4856) & (n_n4863) & (!n_n4865)) + ((!n_n4857) & (n_n4862) & (n_n4856) & (n_n4863) & (n_n4865)) + ((n_n4857) & (!n_n4862) & (!n_n4856) & (!n_n4863) & (!n_n4865)) + ((n_n4857) & (!n_n4862) & (!n_n4856) & (!n_n4863) & (n_n4865)) + ((n_n4857) & (!n_n4862) & (!n_n4856) & (n_n4863) & (!n_n4865)) + ((n_n4857) & (!n_n4862) & (!n_n4856) & (n_n4863) & (n_n4865)) + ((n_n4857) & (!n_n4862) & (n_n4856) & (!n_n4863) & (!n_n4865)) + ((n_n4857) & (!n_n4862) & (n_n4856) & (!n_n4863) & (n_n4865)) + ((n_n4857) & (!n_n4862) & (n_n4856) & (n_n4863) & (!n_n4865)) + ((n_n4857) & (!n_n4862) & (n_n4856) & (n_n4863) & (n_n4865)) + ((n_n4857) & (n_n4862) & (!n_n4856) & (!n_n4863) & (!n_n4865)) + ((n_n4857) & (n_n4862) & (!n_n4856) & (!n_n4863) & (n_n4865)) + ((n_n4857) & (n_n4862) & (!n_n4856) & (n_n4863) & (!n_n4865)) + ((n_n4857) & (n_n4862) & (!n_n4856) & (n_n4863) & (n_n4865)) + ((n_n4857) & (n_n4862) & (n_n4856) & (!n_n4863) & (!n_n4865)) + ((n_n4857) & (n_n4862) & (n_n4856) & (!n_n4863) & (n_n4865)) + ((n_n4857) & (n_n4862) & (n_n4856) & (n_n4863) & (!n_n4865)) + ((n_n4857) & (n_n4862) & (n_n4856) & (n_n4863) & (n_n4865)));
	assign n_n4991 = (((!i_9_) & (n_n528) & (n_n509) & (n_n195)));
	assign n_n4996 = (((i_9_) & (n_n509) & (n_n522) & (n_n195)));
	assign n_n4992 = (((i_9_) & (n_n526) & (n_n509) & (n_n195)));
	assign n_n4995 = (((!i_9_) & (n_n524) & (n_n509) & (n_n195)));
	assign n_n4990 = (((i_9_) & (n_n528) & (n_n509) & (n_n195)));
	assign n_n4998 = (((i_9_) & (n_n509) & (n_n520) & (n_n195)));
	assign n_n4999 = (((i_5_) & (i_3_) & (!i_4_) & (n_n195) & (x23x)));
	assign n_n500 = (((!i_5_) & (i_3_) & (!i_4_)));
	assign n_n5000 = (((i_9_) & (n_n534) & (n_n195) & (n_n500)));
	assign n_n5001 = (((!i_9_) & (n_n534) & (n_n195) & (n_n500)));
	assign x103x = (((!i_9_) & (n_n534) & (n_n195) & (n_n500)) + ((i_9_) & (n_n534) & (n_n195) & (n_n500)));
	assign x13381x = (((!n_n4990) & (!n_n4998) & (!n_n4999) & (!n_n5000) & (n_n5001)) + ((!n_n4990) & (!n_n4998) & (!n_n4999) & (n_n5000) & (!n_n5001)) + ((!n_n4990) & (!n_n4998) & (!n_n4999) & (n_n5000) & (n_n5001)) + ((!n_n4990) & (!n_n4998) & (n_n4999) & (!n_n5000) & (!n_n5001)) + ((!n_n4990) & (!n_n4998) & (n_n4999) & (!n_n5000) & (n_n5001)) + ((!n_n4990) & (!n_n4998) & (n_n4999) & (n_n5000) & (!n_n5001)) + ((!n_n4990) & (!n_n4998) & (n_n4999) & (n_n5000) & (n_n5001)) + ((!n_n4990) & (n_n4998) & (!n_n4999) & (!n_n5000) & (!n_n5001)) + ((!n_n4990) & (n_n4998) & (!n_n4999) & (!n_n5000) & (n_n5001)) + ((!n_n4990) & (n_n4998) & (!n_n4999) & (n_n5000) & (!n_n5001)) + ((!n_n4990) & (n_n4998) & (!n_n4999) & (n_n5000) & (n_n5001)) + ((!n_n4990) & (n_n4998) & (n_n4999) & (!n_n5000) & (!n_n5001)) + ((!n_n4990) & (n_n4998) & (n_n4999) & (!n_n5000) & (n_n5001)) + ((!n_n4990) & (n_n4998) & (n_n4999) & (n_n5000) & (!n_n5001)) + ((!n_n4990) & (n_n4998) & (n_n4999) & (n_n5000) & (n_n5001)) + ((n_n4990) & (!n_n4998) & (!n_n4999) & (!n_n5000) & (!n_n5001)) + ((n_n4990) & (!n_n4998) & (!n_n4999) & (!n_n5000) & (n_n5001)) + ((n_n4990) & (!n_n4998) & (!n_n4999) & (n_n5000) & (!n_n5001)) + ((n_n4990) & (!n_n4998) & (!n_n4999) & (n_n5000) & (n_n5001)) + ((n_n4990) & (!n_n4998) & (n_n4999) & (!n_n5000) & (!n_n5001)) + ((n_n4990) & (!n_n4998) & (n_n4999) & (!n_n5000) & (n_n5001)) + ((n_n4990) & (!n_n4998) & (n_n4999) & (n_n5000) & (!n_n5001)) + ((n_n4990) & (!n_n4998) & (n_n4999) & (n_n5000) & (n_n5001)) + ((n_n4990) & (n_n4998) & (!n_n4999) & (!n_n5000) & (!n_n5001)) + ((n_n4990) & (n_n4998) & (!n_n4999) & (!n_n5000) & (n_n5001)) + ((n_n4990) & (n_n4998) & (!n_n4999) & (n_n5000) & (!n_n5001)) + ((n_n4990) & (n_n4998) & (!n_n4999) & (n_n5000) & (n_n5001)) + ((n_n4990) & (n_n4998) & (n_n4999) & (!n_n5000) & (!n_n5001)) + ((n_n4990) & (n_n4998) & (n_n4999) & (!n_n5000) & (n_n5001)) + ((n_n4990) & (n_n4998) & (n_n4999) & (n_n5000) & (!n_n5001)) + ((n_n4990) & (n_n4998) & (n_n4999) & (n_n5000) & (n_n5001)));
	assign n_n4051 = (((!n_n4991) & (!n_n4996) & (!n_n4992) & (!n_n4995) & (x13381x)) + ((!n_n4991) & (!n_n4996) & (!n_n4992) & (n_n4995) & (!x13381x)) + ((!n_n4991) & (!n_n4996) & (!n_n4992) & (n_n4995) & (x13381x)) + ((!n_n4991) & (!n_n4996) & (n_n4992) & (!n_n4995) & (!x13381x)) + ((!n_n4991) & (!n_n4996) & (n_n4992) & (!n_n4995) & (x13381x)) + ((!n_n4991) & (!n_n4996) & (n_n4992) & (n_n4995) & (!x13381x)) + ((!n_n4991) & (!n_n4996) & (n_n4992) & (n_n4995) & (x13381x)) + ((!n_n4991) & (n_n4996) & (!n_n4992) & (!n_n4995) & (!x13381x)) + ((!n_n4991) & (n_n4996) & (!n_n4992) & (!n_n4995) & (x13381x)) + ((!n_n4991) & (n_n4996) & (!n_n4992) & (n_n4995) & (!x13381x)) + ((!n_n4991) & (n_n4996) & (!n_n4992) & (n_n4995) & (x13381x)) + ((!n_n4991) & (n_n4996) & (n_n4992) & (!n_n4995) & (!x13381x)) + ((!n_n4991) & (n_n4996) & (n_n4992) & (!n_n4995) & (x13381x)) + ((!n_n4991) & (n_n4996) & (n_n4992) & (n_n4995) & (!x13381x)) + ((!n_n4991) & (n_n4996) & (n_n4992) & (n_n4995) & (x13381x)) + ((n_n4991) & (!n_n4996) & (!n_n4992) & (!n_n4995) & (!x13381x)) + ((n_n4991) & (!n_n4996) & (!n_n4992) & (!n_n4995) & (x13381x)) + ((n_n4991) & (!n_n4996) & (!n_n4992) & (n_n4995) & (!x13381x)) + ((n_n4991) & (!n_n4996) & (!n_n4992) & (n_n4995) & (x13381x)) + ((n_n4991) & (!n_n4996) & (n_n4992) & (!n_n4995) & (!x13381x)) + ((n_n4991) & (!n_n4996) & (n_n4992) & (!n_n4995) & (x13381x)) + ((n_n4991) & (!n_n4996) & (n_n4992) & (n_n4995) & (!x13381x)) + ((n_n4991) & (!n_n4996) & (n_n4992) & (n_n4995) & (x13381x)) + ((n_n4991) & (n_n4996) & (!n_n4992) & (!n_n4995) & (!x13381x)) + ((n_n4991) & (n_n4996) & (!n_n4992) & (!n_n4995) & (x13381x)) + ((n_n4991) & (n_n4996) & (!n_n4992) & (n_n4995) & (!x13381x)) + ((n_n4991) & (n_n4996) & (!n_n4992) & (n_n4995) & (x13381x)) + ((n_n4991) & (n_n4996) & (n_n4992) & (!n_n4995) & (!x13381x)) + ((n_n4991) & (n_n4996) & (n_n4992) & (!n_n4995) & (x13381x)) + ((n_n4991) & (n_n4996) & (n_n4992) & (n_n4995) & (!x13381x)) + ((n_n4991) & (n_n4996) & (n_n4992) & (n_n4995) & (x13381x)));
	assign n_n4617 = (((!i_9_) & (n_n390) & (n_n534) & (n_n500)));
	assign n_n4637 = (((!i_9_) & (n_n390) & (n_n491) & (n_n530)));
	assign n_n4613 = (((!i_1_) & (i_2_) & (i_0_) & (n_n509) & (x20x)));
	assign n_n4927 = (((!i_9_) & (n_n528) & (n_n473) & (n_n260)));
	assign n_n4958 = (((i_9_) & (n_n528) & (n_n535) & (n_n195)));
	assign n_n4920 = (((i_9_) & (n_n473) & (n_n534) & (n_n260)));
	assign n_n4324 = (((i_9_) & (n_n536) & (n_n535) & (n_n522)));
	assign n_n4382 = (((i_9_) & (n_n536) & (n_n528) & (n_n491)));
	assign n_n4383 = (((!i_9_) & (n_n536) & (n_n528) & (n_n491)));
	assign x572x = (((i_5_) & (!i_3_) & (i_4_) & (n_n530)));
	assign n_n4923 = (((!i_9_) & (n_n473) & (n_n532) & (n_n260)));
	assign n_n4924 = (((i_9_) & (n_n473) & (n_n260) & (n_n530)));
	assign n_n4921 = (((!i_9_) & (n_n473) & (n_n534) & (n_n260)));
	assign n_n4982 = (((i_9_) & (n_n518) & (n_n520) & (n_n195)));
	assign n_n4983 = (((!i_5_) & (i_3_) & (i_4_) & (n_n195) & (x23x)));
	assign n_n4981 = (((!i_5_) & (i_3_) & (i_4_) & (n_n195) & (x20x)));
	assign n_n5035 = (((!i_9_) & (n_n482) & (n_n532) & (n_n195)));
	assign n_n5032 = (((i_9_) & (n_n482) & (n_n534) & (n_n195)));
	assign n_n5111 = (((!i_5_) & (i_3_) & (i_4_) & (n_n130) & (x23x)));
	assign n_n5112 = (((i_7_) & (i_8_) & (i_6_) & (n_n509) & (x12x)));
	assign n_n5109 = (((!i_5_) & (i_3_) & (i_4_) & (n_n130) & (x20x)));
	assign n_n5171 = (((!i_9_) & (n_n524) & (n_n482) & (n_n130)));
	assign n_n5174 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n520) & (x12x)));
	assign n_n5167 = (((!i_9_) & (n_n482) & (n_n528) & (n_n130)));
	assign x583x = (((!i_5_) & (i_3_) & (i_4_) & (n_n390)));
	assign n_n4597 = (((!i_5_) & (i_3_) & (i_4_) & (n_n390) & (x20x)));
	assign n_n4598 = (((i_9_) & (n_n518) & (n_n390) & (n_n520)));
	assign n_n4602 = (((i_9_) & (n_n390) & (n_n532) & (n_n509)));
	assign n_n4593 = (((!i_9_) & (n_n518) & (n_n526) & (n_n390)));
	assign n_n4601 = (((!i_9_) & (n_n390) & (n_n534) & (n_n509)));
	assign n_n4605 = (((!i_9_) & (n_n390) & (n_n509) & (n_n530)));
	assign x108x = (((!i_9_) & (n_n390) & (n_n509) & (n_n530)) + ((i_9_) & (n_n390) & (n_n509) & (n_n530)));
	assign n_n4595 = (((!i_9_) & (n_n524) & (n_n518) & (n_n390)));
	assign n_n4596 = (((i_9_) & (n_n518) & (n_n390) & (n_n522)));
	assign x257x = (((!i_9_) & (n_n524) & (n_n518) & (n_n390) & (!n_n522)) + ((!i_9_) & (n_n524) & (n_n518) & (n_n390) & (n_n522)) + ((i_9_) & (!n_n524) & (n_n518) & (n_n390) & (n_n522)) + ((i_9_) & (n_n524) & (n_n518) & (n_n390) & (n_n522)));
	assign x22114x = (((!x20x) & (!x583x) & (!n_n4598) & (!n_n4601) & (!x108x)) + ((!x20x) & (x583x) & (!n_n4598) & (!n_n4601) & (!x108x)) + ((x20x) & (!x583x) & (!n_n4598) & (!n_n4601) & (!x108x)));
	assign n_n3347 = (((!n_n4602) & (!n_n4593) & (!n_n4595) & (!n_n4596) & (!x22114x)) + ((!n_n4602) & (!n_n4593) & (!n_n4595) & (n_n4596) & (!x22114x)) + ((!n_n4602) & (!n_n4593) & (!n_n4595) & (n_n4596) & (x22114x)) + ((!n_n4602) & (!n_n4593) & (n_n4595) & (!n_n4596) & (!x22114x)) + ((!n_n4602) & (!n_n4593) & (n_n4595) & (!n_n4596) & (x22114x)) + ((!n_n4602) & (!n_n4593) & (n_n4595) & (n_n4596) & (!x22114x)) + ((!n_n4602) & (!n_n4593) & (n_n4595) & (n_n4596) & (x22114x)) + ((!n_n4602) & (n_n4593) & (!n_n4595) & (!n_n4596) & (!x22114x)) + ((!n_n4602) & (n_n4593) & (!n_n4595) & (!n_n4596) & (x22114x)) + ((!n_n4602) & (n_n4593) & (!n_n4595) & (n_n4596) & (!x22114x)) + ((!n_n4602) & (n_n4593) & (!n_n4595) & (n_n4596) & (x22114x)) + ((!n_n4602) & (n_n4593) & (n_n4595) & (!n_n4596) & (!x22114x)) + ((!n_n4602) & (n_n4593) & (n_n4595) & (!n_n4596) & (x22114x)) + ((!n_n4602) & (n_n4593) & (n_n4595) & (n_n4596) & (!x22114x)) + ((!n_n4602) & (n_n4593) & (n_n4595) & (n_n4596) & (x22114x)) + ((n_n4602) & (!n_n4593) & (!n_n4595) & (!n_n4596) & (!x22114x)) + ((n_n4602) & (!n_n4593) & (!n_n4595) & (!n_n4596) & (x22114x)) + ((n_n4602) & (!n_n4593) & (!n_n4595) & (n_n4596) & (!x22114x)) + ((n_n4602) & (!n_n4593) & (!n_n4595) & (n_n4596) & (x22114x)) + ((n_n4602) & (!n_n4593) & (n_n4595) & (!n_n4596) & (!x22114x)) + ((n_n4602) & (!n_n4593) & (n_n4595) & (!n_n4596) & (x22114x)) + ((n_n4602) & (!n_n4593) & (n_n4595) & (n_n4596) & (!x22114x)) + ((n_n4602) & (!n_n4593) & (n_n4595) & (n_n4596) & (x22114x)) + ((n_n4602) & (n_n4593) & (!n_n4595) & (!n_n4596) & (!x22114x)) + ((n_n4602) & (n_n4593) & (!n_n4595) & (!n_n4596) & (x22114x)) + ((n_n4602) & (n_n4593) & (!n_n4595) & (n_n4596) & (!x22114x)) + ((n_n4602) & (n_n4593) & (!n_n4595) & (n_n4596) & (x22114x)) + ((n_n4602) & (n_n4593) & (n_n4595) & (!n_n4596) & (!x22114x)) + ((n_n4602) & (n_n4593) & (n_n4595) & (!n_n4596) & (x22114x)) + ((n_n4602) & (n_n4593) & (n_n4595) & (n_n4596) & (!x22114x)) + ((n_n4602) & (n_n4593) & (n_n4595) & (n_n4596) & (x22114x)));
	assign n_n4744 = (((i_9_) & (n_n534) & (n_n325) & (n_n500)));
	assign n_n4754 = (((i_9_) & (n_n524) & (n_n325) & (n_n500)));
	assign n_n4757 = (((!i_1_) & (!i_2_) & (i_0_) & (x20x) & (n_n500)));
	assign n_n4749 = (((!i_9_) & (n_n325) & (n_n500) & (n_n530)));
	assign n_n4756 = (((i_9_) & (n_n325) & (n_n522) & (n_n500)));
	assign n_n4751 = (((!i_9_) & (n_n528) & (n_n325) & (n_n500)));
	assign n_n4750 = (((i_9_) & (n_n528) & (n_n325) & (n_n500)));
	assign x109x = (((!i_9_) & (n_n528) & (n_n325) & (n_n500)) + ((i_9_) & (n_n528) & (n_n325) & (n_n500)));
	assign n_n4747 = (((!i_9_) & (n_n532) & (n_n325) & (n_n500)));
	assign x22117x = (((!n_n4744) & (!n_n4754) & (!n_n4757) & (!n_n4749)));
	assign n_n3336 = (((!n_n4756) & (!x109x) & (!n_n4748) & (!n_n4747) & (!x22117x)) + ((!n_n4756) & (!x109x) & (!n_n4748) & (n_n4747) & (!x22117x)) + ((!n_n4756) & (!x109x) & (!n_n4748) & (n_n4747) & (x22117x)) + ((!n_n4756) & (!x109x) & (n_n4748) & (!n_n4747) & (!x22117x)) + ((!n_n4756) & (!x109x) & (n_n4748) & (!n_n4747) & (x22117x)) + ((!n_n4756) & (!x109x) & (n_n4748) & (n_n4747) & (!x22117x)) + ((!n_n4756) & (!x109x) & (n_n4748) & (n_n4747) & (x22117x)) + ((!n_n4756) & (x109x) & (!n_n4748) & (!n_n4747) & (!x22117x)) + ((!n_n4756) & (x109x) & (!n_n4748) & (!n_n4747) & (x22117x)) + ((!n_n4756) & (x109x) & (!n_n4748) & (n_n4747) & (!x22117x)) + ((!n_n4756) & (x109x) & (!n_n4748) & (n_n4747) & (x22117x)) + ((!n_n4756) & (x109x) & (n_n4748) & (!n_n4747) & (!x22117x)) + ((!n_n4756) & (x109x) & (n_n4748) & (!n_n4747) & (x22117x)) + ((!n_n4756) & (x109x) & (n_n4748) & (n_n4747) & (!x22117x)) + ((!n_n4756) & (x109x) & (n_n4748) & (n_n4747) & (x22117x)) + ((n_n4756) & (!x109x) & (!n_n4748) & (!n_n4747) & (!x22117x)) + ((n_n4756) & (!x109x) & (!n_n4748) & (!n_n4747) & (x22117x)) + ((n_n4756) & (!x109x) & (!n_n4748) & (n_n4747) & (!x22117x)) + ((n_n4756) & (!x109x) & (!n_n4748) & (n_n4747) & (x22117x)) + ((n_n4756) & (!x109x) & (n_n4748) & (!n_n4747) & (!x22117x)) + ((n_n4756) & (!x109x) & (n_n4748) & (!n_n4747) & (x22117x)) + ((n_n4756) & (!x109x) & (n_n4748) & (n_n4747) & (!x22117x)) + ((n_n4756) & (!x109x) & (n_n4748) & (n_n4747) & (x22117x)) + ((n_n4756) & (x109x) & (!n_n4748) & (!n_n4747) & (!x22117x)) + ((n_n4756) & (x109x) & (!n_n4748) & (!n_n4747) & (x22117x)) + ((n_n4756) & (x109x) & (!n_n4748) & (n_n4747) & (!x22117x)) + ((n_n4756) & (x109x) & (!n_n4748) & (n_n4747) & (x22117x)) + ((n_n4756) & (x109x) & (n_n4748) & (!n_n4747) & (!x22117x)) + ((n_n4756) & (x109x) & (n_n4748) & (!n_n4747) & (x22117x)) + ((n_n4756) & (x109x) & (n_n4748) & (n_n4747) & (!x22117x)) + ((n_n4756) & (x109x) & (n_n4748) & (n_n4747) & (x22117x)));
	assign n_n4887 = (((i_1_) & (i_2_) & (!i_0_) & (x23x) & (n_n500)));
	assign n_n4888 = (((i_9_) & (n_n534) & (n_n260) & (n_n491)));
	assign n_n4885 = (((i_1_) & (i_2_) & (!i_0_) & (x20x) & (n_n500)));
	assign n_n3450 = (((!n_n260) & (!x20x) & (!x23x) & (!n_n500) & (n_n4888)) + ((!n_n260) & (!x20x) & (!x23x) & (n_n500) & (n_n4888)) + ((!n_n260) & (!x20x) & (x23x) & (!n_n500) & (n_n4888)) + ((!n_n260) & (!x20x) & (x23x) & (n_n500) & (n_n4888)) + ((!n_n260) & (x20x) & (!x23x) & (!n_n500) & (n_n4888)) + ((!n_n260) & (x20x) & (!x23x) & (n_n500) & (n_n4888)) + ((!n_n260) & (x20x) & (x23x) & (!n_n500) & (n_n4888)) + ((!n_n260) & (x20x) & (x23x) & (n_n500) & (n_n4888)) + ((n_n260) & (!x20x) & (!x23x) & (!n_n500) & (n_n4888)) + ((n_n260) & (!x20x) & (!x23x) & (n_n500) & (n_n4888)) + ((n_n260) & (!x20x) & (x23x) & (!n_n500) & (n_n4888)) + ((n_n260) & (!x20x) & (x23x) & (n_n500) & (!n_n4888)) + ((n_n260) & (!x20x) & (x23x) & (n_n500) & (n_n4888)) + ((n_n260) & (x20x) & (!x23x) & (!n_n500) & (n_n4888)) + ((n_n260) & (x20x) & (!x23x) & (n_n500) & (!n_n4888)) + ((n_n260) & (x20x) & (!x23x) & (n_n500) & (n_n4888)) + ((n_n260) & (x20x) & (x23x) & (!n_n500) & (n_n4888)) + ((n_n260) & (x20x) & (x23x) & (n_n500) & (!n_n4888)) + ((n_n260) & (x20x) & (x23x) & (n_n500) & (n_n4888)));
	assign n_n4882 = (((i_9_) & (n_n524) & (n_n260) & (n_n500)));
	assign n_n4883 = (((!i_9_) & (n_n524) & (n_n260) & (n_n500)));
	assign x262x = (((!i_9_) & (n_n524) & (n_n260) & (!n_n522) & (n_n500)) + ((!i_9_) & (n_n524) & (n_n260) & (n_n522) & (n_n500)) + ((i_9_) & (!n_n524) & (n_n260) & (n_n522) & (n_n500)) + ((i_9_) & (n_n524) & (n_n260) & (n_n522) & (n_n500)));
	assign n_n3451 = (((!i_9_) & (n_n524) & (n_n260) & (!n_n522) & (n_n500)) + ((!i_9_) & (n_n524) & (n_n260) & (n_n522) & (n_n500)) + ((i_9_) & (!n_n524) & (n_n260) & (n_n522) & (n_n500)) + ((i_9_) & (n_n524) & (n_n260) & (!n_n522) & (n_n500)) + ((i_9_) & (n_n524) & (n_n260) & (n_n522) & (n_n500)));
	assign n_n5026 = (((i_9_) & (n_n524) & (n_n491) & (n_n195)));
	assign n_n5027 = (((!i_9_) & (n_n524) & (n_n491) & (n_n195)));
	assign n_n5025 = (((!i_9_) & (n_n526) & (n_n491) & (n_n195)));
	assign n_n3424 = (((!i_9_) & (!n_n524) & (n_n526) & (n_n491) & (n_n195)) + ((!i_9_) & (n_n524) & (!n_n526) & (n_n491) & (n_n195)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n491) & (n_n195)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n491) & (n_n195)) + ((i_9_) & (n_n524) & (n_n526) & (n_n491) & (n_n195)));
	assign n_n5179 = (((!i_9_) & (n_n473) & (n_n532) & (n_n130)));
	assign n_n5178 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n532) & (x12x)));
	assign n_n3399 = (((!n_n473) & (!n_n532) & (!x12x) & (!n_n530) & (n_n5179)) + ((!n_n473) & (!n_n532) & (!x12x) & (n_n530) & (n_n5179)) + ((!n_n473) & (!n_n532) & (x12x) & (!n_n530) & (n_n5179)) + ((!n_n473) & (!n_n532) & (x12x) & (n_n530) & (n_n5179)) + ((!n_n473) & (n_n532) & (!x12x) & (!n_n530) & (n_n5179)) + ((!n_n473) & (n_n532) & (!x12x) & (n_n530) & (n_n5179)) + ((!n_n473) & (n_n532) & (x12x) & (!n_n530) & (n_n5179)) + ((!n_n473) & (n_n532) & (x12x) & (n_n530) & (n_n5179)) + ((n_n473) & (!n_n532) & (!x12x) & (!n_n530) & (n_n5179)) + ((n_n473) & (!n_n532) & (!x12x) & (n_n530) & (n_n5179)) + ((n_n473) & (!n_n532) & (x12x) & (!n_n530) & (n_n5179)) + ((n_n473) & (!n_n532) & (x12x) & (n_n530) & (!n_n5179)) + ((n_n473) & (!n_n532) & (x12x) & (n_n530) & (n_n5179)) + ((n_n473) & (n_n532) & (!x12x) & (!n_n530) & (n_n5179)) + ((n_n473) & (n_n532) & (!x12x) & (n_n530) & (n_n5179)) + ((n_n473) & (n_n532) & (x12x) & (!n_n530) & (!n_n5179)) + ((n_n473) & (n_n532) & (x12x) & (!n_n530) & (n_n5179)) + ((n_n473) & (n_n532) & (x12x) & (n_n530) & (!n_n5179)) + ((n_n473) & (n_n532) & (x12x) & (n_n530) & (n_n5179)));
	assign n_n5181 = (((!i_9_) & (n_n473) & (n_n130) & (n_n530)));
	assign n_n5184 = (((i_7_) & (i_8_) & (!i_6_) & (n_n473) & (x12x)));
	assign n_n5185 = (((!i_9_) & (n_n526) & (n_n473) & (n_n130)));
	assign n_n5183 = (((!i_9_) & (n_n528) & (n_n473) & (n_n130)));
	assign n_n5186 = (((i_7_) & (!i_8_) & (!i_6_) & (n_n473) & (x12x)));
	assign n_n5187 = (((!i_9_) & (n_n524) & (n_n473) & (n_n130)));
	assign x112x = (((!i_9_) & (n_n524) & (n_n473) & (!n_n130) & (x12x)) + ((!i_9_) & (n_n524) & (n_n473) & (n_n130) & (!x12x)) + ((!i_9_) & (n_n524) & (n_n473) & (n_n130) & (x12x)) + ((i_9_) & (n_n524) & (n_n473) & (!n_n130) & (x12x)) + ((i_9_) & (n_n524) & (n_n473) & (n_n130) & (x12x)));
	assign x14026x = (((!i_9_) & (!n_n473) & (!n_n130) & (!n_n530) & (n_n5184)) + ((!i_9_) & (!n_n473) & (!n_n130) & (n_n530) & (n_n5184)) + ((!i_9_) & (!n_n473) & (n_n130) & (!n_n530) & (n_n5184)) + ((!i_9_) & (!n_n473) & (n_n130) & (n_n530) & (n_n5184)) + ((!i_9_) & (n_n473) & (!n_n130) & (!n_n530) & (n_n5184)) + ((!i_9_) & (n_n473) & (!n_n130) & (n_n530) & (n_n5184)) + ((!i_9_) & (n_n473) & (n_n130) & (!n_n530) & (n_n5184)) + ((!i_9_) & (n_n473) & (n_n130) & (n_n530) & (!n_n5184)) + ((!i_9_) & (n_n473) & (n_n130) & (n_n530) & (n_n5184)) + ((i_9_) & (!n_n473) & (!n_n130) & (!n_n530) & (n_n5184)) + ((i_9_) & (!n_n473) & (!n_n130) & (n_n530) & (n_n5184)) + ((i_9_) & (!n_n473) & (n_n130) & (!n_n530) & (n_n5184)) + ((i_9_) & (!n_n473) & (n_n130) & (n_n530) & (n_n5184)) + ((i_9_) & (n_n473) & (!n_n130) & (!n_n530) & (n_n5184)) + ((i_9_) & (n_n473) & (!n_n130) & (n_n530) & (n_n5184)) + ((i_9_) & (n_n473) & (n_n130) & (!n_n530) & (n_n5184)) + ((i_9_) & (n_n473) & (n_n130) & (n_n530) & (n_n5184)));
	assign n_n3303 = (((!n_n3399) & (!n_n5185) & (!n_n5183) & (!x112x) & (x14026x)) + ((!n_n3399) & (!n_n5185) & (!n_n5183) & (x112x) & (!x14026x)) + ((!n_n3399) & (!n_n5185) & (!n_n5183) & (x112x) & (x14026x)) + ((!n_n3399) & (!n_n5185) & (n_n5183) & (!x112x) & (!x14026x)) + ((!n_n3399) & (!n_n5185) & (n_n5183) & (!x112x) & (x14026x)) + ((!n_n3399) & (!n_n5185) & (n_n5183) & (x112x) & (!x14026x)) + ((!n_n3399) & (!n_n5185) & (n_n5183) & (x112x) & (x14026x)) + ((!n_n3399) & (n_n5185) & (!n_n5183) & (!x112x) & (!x14026x)) + ((!n_n3399) & (n_n5185) & (!n_n5183) & (!x112x) & (x14026x)) + ((!n_n3399) & (n_n5185) & (!n_n5183) & (x112x) & (!x14026x)) + ((!n_n3399) & (n_n5185) & (!n_n5183) & (x112x) & (x14026x)) + ((!n_n3399) & (n_n5185) & (n_n5183) & (!x112x) & (!x14026x)) + ((!n_n3399) & (n_n5185) & (n_n5183) & (!x112x) & (x14026x)) + ((!n_n3399) & (n_n5185) & (n_n5183) & (x112x) & (!x14026x)) + ((!n_n3399) & (n_n5185) & (n_n5183) & (x112x) & (x14026x)) + ((n_n3399) & (!n_n5185) & (!n_n5183) & (!x112x) & (!x14026x)) + ((n_n3399) & (!n_n5185) & (!n_n5183) & (!x112x) & (x14026x)) + ((n_n3399) & (!n_n5185) & (!n_n5183) & (x112x) & (!x14026x)) + ((n_n3399) & (!n_n5185) & (!n_n5183) & (x112x) & (x14026x)) + ((n_n3399) & (!n_n5185) & (n_n5183) & (!x112x) & (!x14026x)) + ((n_n3399) & (!n_n5185) & (n_n5183) & (!x112x) & (x14026x)) + ((n_n3399) & (!n_n5185) & (n_n5183) & (x112x) & (!x14026x)) + ((n_n3399) & (!n_n5185) & (n_n5183) & (x112x) & (x14026x)) + ((n_n3399) & (n_n5185) & (!n_n5183) & (!x112x) & (!x14026x)) + ((n_n3399) & (n_n5185) & (!n_n5183) & (!x112x) & (x14026x)) + ((n_n3399) & (n_n5185) & (!n_n5183) & (x112x) & (!x14026x)) + ((n_n3399) & (n_n5185) & (!n_n5183) & (x112x) & (x14026x)) + ((n_n3399) & (n_n5185) & (n_n5183) & (!x112x) & (!x14026x)) + ((n_n3399) & (n_n5185) & (n_n5183) & (!x112x) & (x14026x)) + ((n_n3399) & (n_n5185) & (n_n5183) & (x112x) & (!x14026x)) + ((n_n3399) & (n_n5185) & (n_n5183) & (x112x) & (x14026x)));
	assign n_n5310 = (((!i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n473)));
	assign x506x = (((i_5_) & (!i_3_) & (!i_4_) & (n_n520)));
	assign n_n5318 = (((i_5_) & (!i_3_) & (!i_4_) & (x19x) & (n_n520)));
	assign n_n5316 = (((i_5_) & (!i_3_) & (!i_4_) & (x19x) & (n_n522)));
	assign x502x = (((i_7_) & (!i_8_) & (!i_6_) & (n_n473)));
	assign n_n5320 = (((i_7_) & (i_8_) & (i_6_) & (x19x) & (n_n464)));
	assign n_n5321 = (((!i_9_) & (n_n534) & (n_n464) & (n_n65)));
	assign n_n5319 = (((i_5_) & (!i_3_) & (!i_4_) & (x23x) & (n_n65)));
	assign x268x = (((!i_9_) & (!n_n534) & (n_n5319) & (!n_n464) & (!n_n65)) + ((!i_9_) & (!n_n534) & (n_n5319) & (!n_n464) & (n_n65)) + ((!i_9_) & (!n_n534) & (n_n5319) & (n_n464) & (!n_n65)) + ((!i_9_) & (!n_n534) & (n_n5319) & (n_n464) & (n_n65)) + ((!i_9_) & (n_n534) & (!n_n5319) & (n_n464) & (n_n65)) + ((!i_9_) & (n_n534) & (n_n5319) & (!n_n464) & (!n_n65)) + ((!i_9_) & (n_n534) & (n_n5319) & (!n_n464) & (n_n65)) + ((!i_9_) & (n_n534) & (n_n5319) & (n_n464) & (!n_n65)) + ((!i_9_) & (n_n534) & (n_n5319) & (n_n464) & (n_n65)) + ((i_9_) & (!n_n534) & (n_n5319) & (!n_n464) & (!n_n65)) + ((i_9_) & (!n_n534) & (n_n5319) & (!n_n464) & (n_n65)) + ((i_9_) & (!n_n534) & (n_n5319) & (n_n464) & (!n_n65)) + ((i_9_) & (!n_n534) & (n_n5319) & (n_n464) & (n_n65)) + ((i_9_) & (n_n534) & (n_n5319) & (!n_n464) & (!n_n65)) + ((i_9_) & (n_n534) & (n_n5319) & (!n_n464) & (n_n65)) + ((i_9_) & (n_n534) & (n_n5319) & (n_n464) & (!n_n65)) + ((i_9_) & (n_n534) & (n_n5319) & (n_n464) & (n_n65)));
	assign n_n5312 = (((i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n473)));
	assign n_n5313 = (((!i_9_) & (n_n526) & (n_n473) & (n_n65)));
	assign x459x = (((!i_9_) & (!x19x) & (n_n526) & (n_n473) & (n_n65)) + ((!i_9_) & (x19x) & (n_n526) & (n_n473) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n526) & (n_n473) & (n_n65)) + ((i_9_) & (x19x) & (n_n526) & (n_n473) & (!n_n65)) + ((i_9_) & (x19x) & (n_n526) & (n_n473) & (n_n65)));
	assign x13935x = (((!x19x) & (!n_n5316) & (!x502x) & (!n_n5320) & (x268x)) + ((!x19x) & (!n_n5316) & (!x502x) & (n_n5320) & (!x268x)) + ((!x19x) & (!n_n5316) & (!x502x) & (n_n5320) & (x268x)) + ((!x19x) & (!n_n5316) & (x502x) & (!n_n5320) & (x268x)) + ((!x19x) & (!n_n5316) & (x502x) & (n_n5320) & (!x268x)) + ((!x19x) & (!n_n5316) & (x502x) & (n_n5320) & (x268x)) + ((!x19x) & (n_n5316) & (!x502x) & (!n_n5320) & (!x268x)) + ((!x19x) & (n_n5316) & (!x502x) & (!n_n5320) & (x268x)) + ((!x19x) & (n_n5316) & (!x502x) & (n_n5320) & (!x268x)) + ((!x19x) & (n_n5316) & (!x502x) & (n_n5320) & (x268x)) + ((!x19x) & (n_n5316) & (x502x) & (!n_n5320) & (!x268x)) + ((!x19x) & (n_n5316) & (x502x) & (!n_n5320) & (x268x)) + ((!x19x) & (n_n5316) & (x502x) & (n_n5320) & (!x268x)) + ((!x19x) & (n_n5316) & (x502x) & (n_n5320) & (x268x)) + ((x19x) & (!n_n5316) & (!x502x) & (!n_n5320) & (x268x)) + ((x19x) & (!n_n5316) & (!x502x) & (n_n5320) & (!x268x)) + ((x19x) & (!n_n5316) & (!x502x) & (n_n5320) & (x268x)) + ((x19x) & (!n_n5316) & (x502x) & (!n_n5320) & (!x268x)) + ((x19x) & (!n_n5316) & (x502x) & (!n_n5320) & (x268x)) + ((x19x) & (!n_n5316) & (x502x) & (n_n5320) & (!x268x)) + ((x19x) & (!n_n5316) & (x502x) & (n_n5320) & (x268x)) + ((x19x) & (n_n5316) & (!x502x) & (!n_n5320) & (!x268x)) + ((x19x) & (n_n5316) & (!x502x) & (!n_n5320) & (x268x)) + ((x19x) & (n_n5316) & (!x502x) & (n_n5320) & (!x268x)) + ((x19x) & (n_n5316) & (!x502x) & (n_n5320) & (x268x)) + ((x19x) & (n_n5316) & (x502x) & (!n_n5320) & (!x268x)) + ((x19x) & (n_n5316) & (x502x) & (!n_n5320) & (x268x)) + ((x19x) & (n_n5316) & (x502x) & (n_n5320) & (!x268x)) + ((x19x) & (n_n5316) & (x502x) & (n_n5320) & (x268x)));
	assign n_n3292 = (((!x19x) & (!n_n5310) & (!x506x) & (!x459x) & (x13935x)) + ((!x19x) & (!n_n5310) & (!x506x) & (x459x) & (!x13935x)) + ((!x19x) & (!n_n5310) & (!x506x) & (x459x) & (x13935x)) + ((!x19x) & (!n_n5310) & (x506x) & (!x459x) & (x13935x)) + ((!x19x) & (!n_n5310) & (x506x) & (x459x) & (!x13935x)) + ((!x19x) & (!n_n5310) & (x506x) & (x459x) & (x13935x)) + ((!x19x) & (n_n5310) & (!x506x) & (!x459x) & (!x13935x)) + ((!x19x) & (n_n5310) & (!x506x) & (!x459x) & (x13935x)) + ((!x19x) & (n_n5310) & (!x506x) & (x459x) & (!x13935x)) + ((!x19x) & (n_n5310) & (!x506x) & (x459x) & (x13935x)) + ((!x19x) & (n_n5310) & (x506x) & (!x459x) & (!x13935x)) + ((!x19x) & (n_n5310) & (x506x) & (!x459x) & (x13935x)) + ((!x19x) & (n_n5310) & (x506x) & (x459x) & (!x13935x)) + ((!x19x) & (n_n5310) & (x506x) & (x459x) & (x13935x)) + ((x19x) & (!n_n5310) & (!x506x) & (!x459x) & (x13935x)) + ((x19x) & (!n_n5310) & (!x506x) & (x459x) & (!x13935x)) + ((x19x) & (!n_n5310) & (!x506x) & (x459x) & (x13935x)) + ((x19x) & (!n_n5310) & (x506x) & (!x459x) & (!x13935x)) + ((x19x) & (!n_n5310) & (x506x) & (!x459x) & (x13935x)) + ((x19x) & (!n_n5310) & (x506x) & (x459x) & (!x13935x)) + ((x19x) & (!n_n5310) & (x506x) & (x459x) & (x13935x)) + ((x19x) & (n_n5310) & (!x506x) & (!x459x) & (!x13935x)) + ((x19x) & (n_n5310) & (!x506x) & (!x459x) & (x13935x)) + ((x19x) & (n_n5310) & (!x506x) & (x459x) & (!x13935x)) + ((x19x) & (n_n5310) & (!x506x) & (x459x) & (x13935x)) + ((x19x) & (n_n5310) & (x506x) & (!x459x) & (!x13935x)) + ((x19x) & (n_n5310) & (x506x) & (!x459x) & (x13935x)) + ((x19x) & (n_n5310) & (x506x) & (x459x) & (!x13935x)) + ((x19x) & (n_n5310) & (x506x) & (x459x) & (x13935x)));
	assign n_n4615 = (((!i_1_) & (i_2_) & (i_0_) & (n_n509) & (x23x)));
	assign n_n4616 = (((i_9_) & (n_n390) & (n_n534) & (n_n500)));
	assign n_n4607 = (((!i_9_) & (n_n528) & (n_n390) & (n_n509)));
	assign n_n4612 = (((i_9_) & (n_n390) & (n_n509) & (n_n522)));
	assign n_n4609 = (((!i_9_) & (n_n526) & (n_n390) & (n_n509)));
	assign n_n4608 = (((i_9_) & (n_n526) & (n_n390) & (n_n509)));
	assign n_n4606 = (((i_9_) & (n_n528) & (n_n390) & (n_n509)));
	assign x14072x = (((!n_n4617) & (!n_n4613) & (!n_n4608) & (n_n4606)) + ((!n_n4617) & (!n_n4613) & (n_n4608) & (!n_n4606)) + ((!n_n4617) & (!n_n4613) & (n_n4608) & (n_n4606)) + ((!n_n4617) & (n_n4613) & (!n_n4608) & (!n_n4606)) + ((!n_n4617) & (n_n4613) & (!n_n4608) & (n_n4606)) + ((!n_n4617) & (n_n4613) & (n_n4608) & (!n_n4606)) + ((!n_n4617) & (n_n4613) & (n_n4608) & (n_n4606)) + ((n_n4617) & (!n_n4613) & (!n_n4608) & (!n_n4606)) + ((n_n4617) & (!n_n4613) & (!n_n4608) & (n_n4606)) + ((n_n4617) & (!n_n4613) & (n_n4608) & (!n_n4606)) + ((n_n4617) & (!n_n4613) & (n_n4608) & (n_n4606)) + ((n_n4617) & (n_n4613) & (!n_n4608) & (!n_n4606)) + ((n_n4617) & (n_n4613) & (!n_n4608) & (n_n4606)) + ((n_n4617) & (n_n4613) & (n_n4608) & (!n_n4606)) + ((n_n4617) & (n_n4613) & (n_n4608) & (n_n4606)));
	assign x14073x = (((!n_n4615) & (!n_n4616) & (!n_n4607) & (!n_n4612) & (n_n4609)) + ((!n_n4615) & (!n_n4616) & (!n_n4607) & (n_n4612) & (!n_n4609)) + ((!n_n4615) & (!n_n4616) & (!n_n4607) & (n_n4612) & (n_n4609)) + ((!n_n4615) & (!n_n4616) & (n_n4607) & (!n_n4612) & (!n_n4609)) + ((!n_n4615) & (!n_n4616) & (n_n4607) & (!n_n4612) & (n_n4609)) + ((!n_n4615) & (!n_n4616) & (n_n4607) & (n_n4612) & (!n_n4609)) + ((!n_n4615) & (!n_n4616) & (n_n4607) & (n_n4612) & (n_n4609)) + ((!n_n4615) & (n_n4616) & (!n_n4607) & (!n_n4612) & (!n_n4609)) + ((!n_n4615) & (n_n4616) & (!n_n4607) & (!n_n4612) & (n_n4609)) + ((!n_n4615) & (n_n4616) & (!n_n4607) & (n_n4612) & (!n_n4609)) + ((!n_n4615) & (n_n4616) & (!n_n4607) & (n_n4612) & (n_n4609)) + ((!n_n4615) & (n_n4616) & (n_n4607) & (!n_n4612) & (!n_n4609)) + ((!n_n4615) & (n_n4616) & (n_n4607) & (!n_n4612) & (n_n4609)) + ((!n_n4615) & (n_n4616) & (n_n4607) & (n_n4612) & (!n_n4609)) + ((!n_n4615) & (n_n4616) & (n_n4607) & (n_n4612) & (n_n4609)) + ((n_n4615) & (!n_n4616) & (!n_n4607) & (!n_n4612) & (!n_n4609)) + ((n_n4615) & (!n_n4616) & (!n_n4607) & (!n_n4612) & (n_n4609)) + ((n_n4615) & (!n_n4616) & (!n_n4607) & (n_n4612) & (!n_n4609)) + ((n_n4615) & (!n_n4616) & (!n_n4607) & (n_n4612) & (n_n4609)) + ((n_n4615) & (!n_n4616) & (n_n4607) & (!n_n4612) & (!n_n4609)) + ((n_n4615) & (!n_n4616) & (n_n4607) & (!n_n4612) & (n_n4609)) + ((n_n4615) & (!n_n4616) & (n_n4607) & (n_n4612) & (!n_n4609)) + ((n_n4615) & (!n_n4616) & (n_n4607) & (n_n4612) & (n_n4609)) + ((n_n4615) & (n_n4616) & (!n_n4607) & (!n_n4612) & (!n_n4609)) + ((n_n4615) & (n_n4616) & (!n_n4607) & (!n_n4612) & (n_n4609)) + ((n_n4615) & (n_n4616) & (!n_n4607) & (n_n4612) & (!n_n4609)) + ((n_n4615) & (n_n4616) & (!n_n4607) & (n_n4612) & (n_n4609)) + ((n_n4615) & (n_n4616) & (n_n4607) & (!n_n4612) & (!n_n4609)) + ((n_n4615) & (n_n4616) & (n_n4607) & (!n_n4612) & (n_n4609)) + ((n_n4615) & (n_n4616) & (n_n4607) & (n_n4612) & (!n_n4609)) + ((n_n4615) & (n_n4616) & (n_n4607) & (n_n4612) & (n_n4609)));
	assign n_n4641 = (((!i_9_) & (n_n526) & (n_n390) & (n_n491)));
	assign n_n4634 = (((i_9_) & (n_n390) & (n_n532) & (n_n491)));
	assign n_n4648 = (((i_9_) & (n_n482) & (n_n390) & (n_n534)));
	assign n_n4618 = (((i_9_) & (n_n390) & (n_n532) & (n_n500)));
	assign n_n4628 = (((i_9_) & (n_n390) & (n_n522) & (n_n500)));
	assign n_n4625 = (((!i_9_) & (n_n526) & (n_n390) & (n_n500)));
	assign n_n1649 = (((!i_9_) & (!n_n524) & (n_n526) & (n_n390) & (n_n500)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n390) & (n_n500)) + ((i_9_) & (!n_n524) & (n_n526) & (n_n390) & (n_n500)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n390) & (n_n500)) + ((i_9_) & (n_n524) & (n_n526) & (n_n390) & (n_n500)));
	assign x26x = (((!i_9_) & (n_n390) & (n_n491) & (n_n530)) + ((i_9_) & (n_n390) & (n_n491) & (n_n530)));
	assign n_n4621 = (((!i_9_) & (n_n390) & (n_n500) & (n_n530)));
	assign n_n4619 = (((!i_9_) & (n_n390) & (n_n532) & (n_n500)));
	assign x118x = (((!i_9_) & (n_n390) & (!n_n532) & (n_n500) & (n_n530)) + ((!i_9_) & (n_n390) & (n_n532) & (n_n500) & (!n_n530)) + ((!i_9_) & (n_n390) & (n_n532) & (n_n500) & (n_n530)));
	assign n_n4643 = (((!i_9_) & (n_n524) & (n_n390) & (n_n491)));
	assign n_n4645 = (((!i_1_) & (i_2_) & (i_0_) & (n_n491) & (x20x)));
	assign x309x = (((!i_9_) & (!n_n524) & (n_n390) & (n_n491) & (x20x)) + ((!i_9_) & (n_n524) & (n_n390) & (n_n491) & (!x20x)) + ((!i_9_) & (n_n524) & (n_n390) & (n_n491) & (x20x)) + ((i_9_) & (!n_n524) & (n_n390) & (n_n491) & (x20x)) + ((i_9_) & (n_n524) & (n_n390) & (n_n491) & (x20x)));
	assign n_n4639 = (((!i_9_) & (n_n528) & (n_n390) & (n_n491)));
	assign n_n4642 = (((i_9_) & (n_n524) & (n_n390) & (n_n491)));
	assign x348x = (((!i_9_) & (!n_n524) & (n_n528) & (n_n390) & (n_n491)) + ((!i_9_) & (n_n524) & (n_n528) & (n_n390) & (n_n491)) + ((i_9_) & (n_n524) & (!n_n528) & (n_n390) & (n_n491)) + ((i_9_) & (n_n524) & (n_n528) & (n_n390) & (n_n491)));
	assign n_n4631 = (((!i_1_) & (i_2_) & (i_0_) & (x23x) & (n_n500)));
	assign n_n4632 = (((i_9_) & (n_n390) & (n_n534) & (n_n491)));
	assign x349x = (((!n_n390) & (!x23x) & (!n_n500) & (n_n4632)) + ((!n_n390) & (!x23x) & (n_n500) & (n_n4632)) + ((!n_n390) & (x23x) & (!n_n500) & (n_n4632)) + ((!n_n390) & (x23x) & (n_n500) & (n_n4632)) + ((n_n390) & (!x23x) & (!n_n500) & (n_n4632)) + ((n_n390) & (!x23x) & (n_n500) & (n_n4632)) + ((n_n390) & (x23x) & (!n_n500) & (n_n4632)) + ((n_n390) & (x23x) & (n_n500) & (!n_n4632)) + ((n_n390) & (x23x) & (n_n500) & (n_n4632)));
	assign x14080x = (((!x10x) & (!n_n522) & (!n_n500) & (!n_n1649) & (x26x)) + ((!x10x) & (!n_n522) & (!n_n500) & (n_n1649) & (!x26x)) + ((!x10x) & (!n_n522) & (!n_n500) & (n_n1649) & (x26x)) + ((!x10x) & (!n_n522) & (n_n500) & (!n_n1649) & (x26x)) + ((!x10x) & (!n_n522) & (n_n500) & (n_n1649) & (!x26x)) + ((!x10x) & (!n_n522) & (n_n500) & (n_n1649) & (x26x)) + ((!x10x) & (n_n522) & (!n_n500) & (!n_n1649) & (x26x)) + ((!x10x) & (n_n522) & (!n_n500) & (n_n1649) & (!x26x)) + ((!x10x) & (n_n522) & (!n_n500) & (n_n1649) & (x26x)) + ((!x10x) & (n_n522) & (n_n500) & (!n_n1649) & (x26x)) + ((!x10x) & (n_n522) & (n_n500) & (n_n1649) & (!x26x)) + ((!x10x) & (n_n522) & (n_n500) & (n_n1649) & (x26x)) + ((x10x) & (!n_n522) & (!n_n500) & (!n_n1649) & (x26x)) + ((x10x) & (!n_n522) & (!n_n500) & (n_n1649) & (!x26x)) + ((x10x) & (!n_n522) & (!n_n500) & (n_n1649) & (x26x)) + ((x10x) & (!n_n522) & (n_n500) & (!n_n1649) & (x26x)) + ((x10x) & (!n_n522) & (n_n500) & (n_n1649) & (!x26x)) + ((x10x) & (!n_n522) & (n_n500) & (n_n1649) & (x26x)) + ((x10x) & (n_n522) & (!n_n500) & (!n_n1649) & (x26x)) + ((x10x) & (n_n522) & (!n_n500) & (n_n1649) & (!x26x)) + ((x10x) & (n_n522) & (!n_n500) & (n_n1649) & (x26x)) + ((x10x) & (n_n522) & (n_n500) & (!n_n1649) & (!x26x)) + ((x10x) & (n_n522) & (n_n500) & (!n_n1649) & (x26x)) + ((x10x) & (n_n522) & (n_n500) & (n_n1649) & (!x26x)) + ((x10x) & (n_n522) & (n_n500) & (n_n1649) & (x26x)));
	assign x14082x = (((!n_n4641) & (!n_n4634) & (!n_n4648) & (!n_n4618) & (x14080x)) + ((!n_n4641) & (!n_n4634) & (!n_n4648) & (n_n4618) & (!x14080x)) + ((!n_n4641) & (!n_n4634) & (!n_n4648) & (n_n4618) & (x14080x)) + ((!n_n4641) & (!n_n4634) & (n_n4648) & (!n_n4618) & (!x14080x)) + ((!n_n4641) & (!n_n4634) & (n_n4648) & (!n_n4618) & (x14080x)) + ((!n_n4641) & (!n_n4634) & (n_n4648) & (n_n4618) & (!x14080x)) + ((!n_n4641) & (!n_n4634) & (n_n4648) & (n_n4618) & (x14080x)) + ((!n_n4641) & (n_n4634) & (!n_n4648) & (!n_n4618) & (!x14080x)) + ((!n_n4641) & (n_n4634) & (!n_n4648) & (!n_n4618) & (x14080x)) + ((!n_n4641) & (n_n4634) & (!n_n4648) & (n_n4618) & (!x14080x)) + ((!n_n4641) & (n_n4634) & (!n_n4648) & (n_n4618) & (x14080x)) + ((!n_n4641) & (n_n4634) & (n_n4648) & (!n_n4618) & (!x14080x)) + ((!n_n4641) & (n_n4634) & (n_n4648) & (!n_n4618) & (x14080x)) + ((!n_n4641) & (n_n4634) & (n_n4648) & (n_n4618) & (!x14080x)) + ((!n_n4641) & (n_n4634) & (n_n4648) & (n_n4618) & (x14080x)) + ((n_n4641) & (!n_n4634) & (!n_n4648) & (!n_n4618) & (!x14080x)) + ((n_n4641) & (!n_n4634) & (!n_n4648) & (!n_n4618) & (x14080x)) + ((n_n4641) & (!n_n4634) & (!n_n4648) & (n_n4618) & (!x14080x)) + ((n_n4641) & (!n_n4634) & (!n_n4648) & (n_n4618) & (x14080x)) + ((n_n4641) & (!n_n4634) & (n_n4648) & (!n_n4618) & (!x14080x)) + ((n_n4641) & (!n_n4634) & (n_n4648) & (!n_n4618) & (x14080x)) + ((n_n4641) & (!n_n4634) & (n_n4648) & (n_n4618) & (!x14080x)) + ((n_n4641) & (!n_n4634) & (n_n4648) & (n_n4618) & (x14080x)) + ((n_n4641) & (n_n4634) & (!n_n4648) & (!n_n4618) & (!x14080x)) + ((n_n4641) & (n_n4634) & (!n_n4648) & (!n_n4618) & (x14080x)) + ((n_n4641) & (n_n4634) & (!n_n4648) & (n_n4618) & (!x14080x)) + ((n_n4641) & (n_n4634) & (!n_n4648) & (n_n4618) & (x14080x)) + ((n_n4641) & (n_n4634) & (n_n4648) & (!n_n4618) & (!x14080x)) + ((n_n4641) & (n_n4634) & (n_n4648) & (!n_n4618) & (x14080x)) + ((n_n4641) & (n_n4634) & (n_n4648) & (n_n4618) & (!x14080x)) + ((n_n4641) & (n_n4634) & (n_n4648) & (n_n4618) & (x14080x)));
	assign x14081x = (((!n_n4621) & (!n_n4619) & (!x309x) & (!x348x) & (x349x)) + ((!n_n4621) & (!n_n4619) & (!x309x) & (x348x) & (!x349x)) + ((!n_n4621) & (!n_n4619) & (!x309x) & (x348x) & (x349x)) + ((!n_n4621) & (!n_n4619) & (x309x) & (!x348x) & (!x349x)) + ((!n_n4621) & (!n_n4619) & (x309x) & (!x348x) & (x349x)) + ((!n_n4621) & (!n_n4619) & (x309x) & (x348x) & (!x349x)) + ((!n_n4621) & (!n_n4619) & (x309x) & (x348x) & (x349x)) + ((!n_n4621) & (n_n4619) & (!x309x) & (!x348x) & (!x349x)) + ((!n_n4621) & (n_n4619) & (!x309x) & (!x348x) & (x349x)) + ((!n_n4621) & (n_n4619) & (!x309x) & (x348x) & (!x349x)) + ((!n_n4621) & (n_n4619) & (!x309x) & (x348x) & (x349x)) + ((!n_n4621) & (n_n4619) & (x309x) & (!x348x) & (!x349x)) + ((!n_n4621) & (n_n4619) & (x309x) & (!x348x) & (x349x)) + ((!n_n4621) & (n_n4619) & (x309x) & (x348x) & (!x349x)) + ((!n_n4621) & (n_n4619) & (x309x) & (x348x) & (x349x)) + ((n_n4621) & (!n_n4619) & (!x309x) & (!x348x) & (!x349x)) + ((n_n4621) & (!n_n4619) & (!x309x) & (!x348x) & (x349x)) + ((n_n4621) & (!n_n4619) & (!x309x) & (x348x) & (!x349x)) + ((n_n4621) & (!n_n4619) & (!x309x) & (x348x) & (x349x)) + ((n_n4621) & (!n_n4619) & (x309x) & (!x348x) & (!x349x)) + ((n_n4621) & (!n_n4619) & (x309x) & (!x348x) & (x349x)) + ((n_n4621) & (!n_n4619) & (x309x) & (x348x) & (!x349x)) + ((n_n4621) & (!n_n4619) & (x309x) & (x348x) & (x349x)) + ((n_n4621) & (n_n4619) & (!x309x) & (!x348x) & (!x349x)) + ((n_n4621) & (n_n4619) & (!x309x) & (!x348x) & (x349x)) + ((n_n4621) & (n_n4619) & (!x309x) & (x348x) & (!x349x)) + ((n_n4621) & (n_n4619) & (!x309x) & (x348x) & (x349x)) + ((n_n4621) & (n_n4619) & (x309x) & (!x348x) & (!x349x)) + ((n_n4621) & (n_n4619) & (x309x) & (!x348x) & (x349x)) + ((n_n4621) & (n_n4619) & (x309x) & (x348x) & (!x349x)) + ((n_n4621) & (n_n4619) & (x309x) & (x348x) & (x349x)));
	assign n_n3281 = (((!x14072x) & (!x14073x) & (!x14082x) & (x14081x)) + ((!x14072x) & (!x14073x) & (x14082x) & (!x14081x)) + ((!x14072x) & (!x14073x) & (x14082x) & (x14081x)) + ((!x14072x) & (x14073x) & (!x14082x) & (!x14081x)) + ((!x14072x) & (x14073x) & (!x14082x) & (x14081x)) + ((!x14072x) & (x14073x) & (x14082x) & (!x14081x)) + ((!x14072x) & (x14073x) & (x14082x) & (x14081x)) + ((x14072x) & (!x14073x) & (!x14082x) & (!x14081x)) + ((x14072x) & (!x14073x) & (!x14082x) & (x14081x)) + ((x14072x) & (!x14073x) & (x14082x) & (!x14081x)) + ((x14072x) & (!x14073x) & (x14082x) & (x14081x)) + ((x14072x) & (x14073x) & (!x14082x) & (!x14081x)) + ((x14072x) & (x14073x) & (!x14082x) & (x14081x)) + ((x14072x) & (x14073x) & (x14082x) & (!x14081x)) + ((x14072x) & (x14073x) & (x14082x) & (x14081x)));
	assign n_n5050 = (((i_9_) & (n_n473) & (n_n532) & (n_n195)));
	assign n_n5060 = (((i_9_) & (n_n473) & (n_n522) & (n_n195)));
	assign n_n5055 = (((!i_9_) & (n_n528) & (n_n473) & (n_n195)));
	assign n_n5054 = (((i_9_) & (n_n528) & (n_n473) & (n_n195)));
	assign n_n5059 = (((!i_9_) & (n_n524) & (n_n473) & (n_n195)));
	assign n_n5064 = (((i_9_) & (n_n534) & (n_n195) & (n_n464)));
	assign x120x = (((!i_9_) & (!n_n473) & (!n_n520) & (!n_n195) & (n_n5064)) + ((!i_9_) & (!n_n473) & (!n_n520) & (n_n195) & (n_n5064)) + ((!i_9_) & (!n_n473) & (n_n520) & (!n_n195) & (n_n5064)) + ((!i_9_) & (!n_n473) & (n_n520) & (n_n195) & (n_n5064)) + ((!i_9_) & (n_n473) & (!n_n520) & (!n_n195) & (n_n5064)) + ((!i_9_) & (n_n473) & (!n_n520) & (n_n195) & (n_n5064)) + ((!i_9_) & (n_n473) & (n_n520) & (!n_n195) & (n_n5064)) + ((!i_9_) & (n_n473) & (n_n520) & (n_n195) & (n_n5064)) + ((i_9_) & (!n_n473) & (!n_n520) & (!n_n195) & (n_n5064)) + ((i_9_) & (!n_n473) & (!n_n520) & (n_n195) & (n_n5064)) + ((i_9_) & (!n_n473) & (n_n520) & (!n_n195) & (n_n5064)) + ((i_9_) & (!n_n473) & (n_n520) & (n_n195) & (n_n5064)) + ((i_9_) & (n_n473) & (!n_n520) & (!n_n195) & (n_n5064)) + ((i_9_) & (n_n473) & (!n_n520) & (n_n195) & (n_n5064)) + ((i_9_) & (n_n473) & (n_n520) & (!n_n195) & (n_n5064)) + ((i_9_) & (n_n473) & (n_n520) & (n_n195) & (!n_n5064)) + ((i_9_) & (n_n473) & (n_n520) & (n_n195) & (n_n5064)));
	assign n_n5057 = (((!i_9_) & (n_n526) & (n_n473) & (n_n195)));
	assign n_n5058 = (((i_9_) & (n_n524) & (n_n473) & (n_n195)));
	assign x13982x = (((!n_n5055) & (!n_n5054) & (!n_n5059) & (x120x)) + ((!n_n5055) & (!n_n5054) & (n_n5059) & (!x120x)) + ((!n_n5055) & (!n_n5054) & (n_n5059) & (x120x)) + ((!n_n5055) & (n_n5054) & (!n_n5059) & (!x120x)) + ((!n_n5055) & (n_n5054) & (!n_n5059) & (x120x)) + ((!n_n5055) & (n_n5054) & (n_n5059) & (!x120x)) + ((!n_n5055) & (n_n5054) & (n_n5059) & (x120x)) + ((n_n5055) & (!n_n5054) & (!n_n5059) & (!x120x)) + ((n_n5055) & (!n_n5054) & (!n_n5059) & (x120x)) + ((n_n5055) & (!n_n5054) & (n_n5059) & (!x120x)) + ((n_n5055) & (!n_n5054) & (n_n5059) & (x120x)) + ((n_n5055) & (n_n5054) & (!n_n5059) & (!x120x)) + ((n_n5055) & (n_n5054) & (!n_n5059) & (x120x)) + ((n_n5055) & (n_n5054) & (n_n5059) & (!x120x)) + ((n_n5055) & (n_n5054) & (n_n5059) & (x120x)));
	assign n_n5048 = (((i_9_) & (n_n473) & (n_n534) & (n_n195)));
	assign n_n5028 = (((i_9_) & (n_n522) & (n_n491) & (n_n195)));
	assign n_n5036 = (((i_9_) & (n_n482) & (n_n195) & (n_n530)));
	assign n_n5031 = (((i_5_) & (!i_3_) & (i_4_) & (n_n195) & (x23x)));
	assign x50x = (((!i_9_) & (n_n491) & (!n_n520) & (n_n195) & (x23x)) + ((!i_9_) & (n_n491) & (n_n520) & (n_n195) & (x23x)) + ((i_9_) & (n_n491) & (!n_n520) & (n_n195) & (x23x)) + ((i_9_) & (n_n491) & (n_n520) & (n_n195) & (!x23x)) + ((i_9_) & (n_n491) & (n_n520) & (n_n195) & (x23x)));
	assign x13983x = (((!i_7_) & (!i_8_) & (i_6_) & (n_n482) & (x18x)) + ((i_7_) & (!i_8_) & (!i_6_) & (n_n482) & (x18x)));
	assign x13984x = (((!i_9_) & (!n_n526) & (n_n482) & (n_n528) & (n_n195)) + ((!i_9_) & (n_n526) & (n_n482) & (!n_n528) & (n_n195)) + ((!i_9_) & (n_n526) & (n_n482) & (n_n528) & (n_n195)) + ((i_9_) & (n_n526) & (n_n482) & (!n_n528) & (n_n195)) + ((i_9_) & (n_n526) & (n_n482) & (n_n528) & (n_n195)));
	assign x231x = (((!i_9_) & (n_n482) & (n_n532) & (n_n195)) + ((i_9_) & (n_n482) & (n_n532) & (n_n195)));
	assign n_n5046 = (((i_9_) & (n_n482) & (n_n520) & (n_n195)));
	assign n_n5044 = (((i_9_) & (n_n482) & (n_n522) & (n_n195)));
	assign x356x = (((!i_7_) & (!i_8_) & (!i_6_) & (n_n482) & (x18x)) + ((!i_7_) & (i_8_) & (!i_6_) & (n_n482) & (x18x)));
	assign x13991x = (((!n_n3424) & (!n_n5028) & (!n_n5036) & (!x13983x) & (x13984x)) + ((!n_n3424) & (!n_n5028) & (!n_n5036) & (x13983x) & (!x13984x)) + ((!n_n3424) & (!n_n5028) & (!n_n5036) & (x13983x) & (x13984x)) + ((!n_n3424) & (!n_n5028) & (n_n5036) & (!x13983x) & (!x13984x)) + ((!n_n3424) & (!n_n5028) & (n_n5036) & (!x13983x) & (x13984x)) + ((!n_n3424) & (!n_n5028) & (n_n5036) & (x13983x) & (!x13984x)) + ((!n_n3424) & (!n_n5028) & (n_n5036) & (x13983x) & (x13984x)) + ((!n_n3424) & (n_n5028) & (!n_n5036) & (!x13983x) & (!x13984x)) + ((!n_n3424) & (n_n5028) & (!n_n5036) & (!x13983x) & (x13984x)) + ((!n_n3424) & (n_n5028) & (!n_n5036) & (x13983x) & (!x13984x)) + ((!n_n3424) & (n_n5028) & (!n_n5036) & (x13983x) & (x13984x)) + ((!n_n3424) & (n_n5028) & (n_n5036) & (!x13983x) & (!x13984x)) + ((!n_n3424) & (n_n5028) & (n_n5036) & (!x13983x) & (x13984x)) + ((!n_n3424) & (n_n5028) & (n_n5036) & (x13983x) & (!x13984x)) + ((!n_n3424) & (n_n5028) & (n_n5036) & (x13983x) & (x13984x)) + ((n_n3424) & (!n_n5028) & (!n_n5036) & (!x13983x) & (!x13984x)) + ((n_n3424) & (!n_n5028) & (!n_n5036) & (!x13983x) & (x13984x)) + ((n_n3424) & (!n_n5028) & (!n_n5036) & (x13983x) & (!x13984x)) + ((n_n3424) & (!n_n5028) & (!n_n5036) & (x13983x) & (x13984x)) + ((n_n3424) & (!n_n5028) & (n_n5036) & (!x13983x) & (!x13984x)) + ((n_n3424) & (!n_n5028) & (n_n5036) & (!x13983x) & (x13984x)) + ((n_n3424) & (!n_n5028) & (n_n5036) & (x13983x) & (!x13984x)) + ((n_n3424) & (!n_n5028) & (n_n5036) & (x13983x) & (x13984x)) + ((n_n3424) & (n_n5028) & (!n_n5036) & (!x13983x) & (!x13984x)) + ((n_n3424) & (n_n5028) & (!n_n5036) & (!x13983x) & (x13984x)) + ((n_n3424) & (n_n5028) & (!n_n5036) & (x13983x) & (!x13984x)) + ((n_n3424) & (n_n5028) & (!n_n5036) & (x13983x) & (x13984x)) + ((n_n3424) & (n_n5028) & (n_n5036) & (!x13983x) & (!x13984x)) + ((n_n3424) & (n_n5028) & (n_n5036) & (!x13983x) & (x13984x)) + ((n_n3424) & (n_n5028) & (n_n5036) & (x13983x) & (!x13984x)) + ((n_n3424) & (n_n5028) & (n_n5036) & (x13983x) & (x13984x)));
	assign x13990x = (((!n_n5032) & (!n_n5048) & (!x50x) & (!x231x) & (x356x)) + ((!n_n5032) & (!n_n5048) & (!x50x) & (x231x) & (!x356x)) + ((!n_n5032) & (!n_n5048) & (!x50x) & (x231x) & (x356x)) + ((!n_n5032) & (!n_n5048) & (x50x) & (!x231x) & (!x356x)) + ((!n_n5032) & (!n_n5048) & (x50x) & (!x231x) & (x356x)) + ((!n_n5032) & (!n_n5048) & (x50x) & (x231x) & (!x356x)) + ((!n_n5032) & (!n_n5048) & (x50x) & (x231x) & (x356x)) + ((!n_n5032) & (n_n5048) & (!x50x) & (!x231x) & (!x356x)) + ((!n_n5032) & (n_n5048) & (!x50x) & (!x231x) & (x356x)) + ((!n_n5032) & (n_n5048) & (!x50x) & (x231x) & (!x356x)) + ((!n_n5032) & (n_n5048) & (!x50x) & (x231x) & (x356x)) + ((!n_n5032) & (n_n5048) & (x50x) & (!x231x) & (!x356x)) + ((!n_n5032) & (n_n5048) & (x50x) & (!x231x) & (x356x)) + ((!n_n5032) & (n_n5048) & (x50x) & (x231x) & (!x356x)) + ((!n_n5032) & (n_n5048) & (x50x) & (x231x) & (x356x)) + ((n_n5032) & (!n_n5048) & (!x50x) & (!x231x) & (!x356x)) + ((n_n5032) & (!n_n5048) & (!x50x) & (!x231x) & (x356x)) + ((n_n5032) & (!n_n5048) & (!x50x) & (x231x) & (!x356x)) + ((n_n5032) & (!n_n5048) & (!x50x) & (x231x) & (x356x)) + ((n_n5032) & (!n_n5048) & (x50x) & (!x231x) & (!x356x)) + ((n_n5032) & (!n_n5048) & (x50x) & (!x231x) & (x356x)) + ((n_n5032) & (!n_n5048) & (x50x) & (x231x) & (!x356x)) + ((n_n5032) & (!n_n5048) & (x50x) & (x231x) & (x356x)) + ((n_n5032) & (n_n5048) & (!x50x) & (!x231x) & (!x356x)) + ((n_n5032) & (n_n5048) & (!x50x) & (!x231x) & (x356x)) + ((n_n5032) & (n_n5048) & (!x50x) & (x231x) & (!x356x)) + ((n_n5032) & (n_n5048) & (!x50x) & (x231x) & (x356x)) + ((n_n5032) & (n_n5048) & (x50x) & (!x231x) & (!x356x)) + ((n_n5032) & (n_n5048) & (x50x) & (!x231x) & (x356x)) + ((n_n5032) & (n_n5048) & (x50x) & (x231x) & (!x356x)) + ((n_n5032) & (n_n5048) & (x50x) & (x231x) & (x356x)));
	assign x22222x = (((!n_n5050) & (!n_n5060) & (!n_n5057) & (!n_n5058)));
	assign n_n3270 = (((!x13982x) & (!x13991x) & (!x13990x) & (!x22222x)) + ((!x13982x) & (!x13991x) & (x13990x) & (!x22222x)) + ((!x13982x) & (!x13991x) & (x13990x) & (x22222x)) + ((!x13982x) & (x13991x) & (!x13990x) & (!x22222x)) + ((!x13982x) & (x13991x) & (!x13990x) & (x22222x)) + ((!x13982x) & (x13991x) & (x13990x) & (!x22222x)) + ((!x13982x) & (x13991x) & (x13990x) & (x22222x)) + ((x13982x) & (!x13991x) & (!x13990x) & (!x22222x)) + ((x13982x) & (!x13991x) & (!x13990x) & (x22222x)) + ((x13982x) & (!x13991x) & (x13990x) & (!x22222x)) + ((x13982x) & (!x13991x) & (x13990x) & (x22222x)) + ((x13982x) & (x13991x) & (!x13990x) & (!x22222x)) + ((x13982x) & (x13991x) & (!x13990x) & (x22222x)) + ((x13982x) & (x13991x) & (x13990x) & (!x22222x)) + ((x13982x) & (x13991x) & (x13990x) & (x22222x)));
	assign n_n4571 = (((!i_9_) & (n_n390) & (n_n532) & (n_n535)));
	assign n_n4578 = (((i_9_) & (n_n524) & (n_n390) & (n_n535)));
	assign n_n4570 = (((i_9_) & (n_n390) & (n_n532) & (n_n535)));
	assign n_n4849 = (((!i_9_) & (n_n518) & (n_n526) & (n_n260)));
	assign n_n5096 = (((!i_5_) & (i_3_) & (i_4_) & (n_n534) & (x12x)));
	assign n_n5099 = (((!i_9_) & (n_n518) & (n_n532) & (n_n130)));
	assign n_n5085 = (((!i_9_) & (n_n535) & (n_n130) & (n_n530)));
	assign x280x = (((!i_9_) & (n_n536) & (n_n532) & (n_n491)) + ((i_9_) & (n_n536) & (n_n532) & (n_n491)));
	assign n_n5101 = (((!i_9_) & (n_n518) & (n_n130) & (n_n530)));
	assign n_n5110 = (((!i_5_) & (i_3_) & (i_4_) & (n_n520) & (x12x)));
	assign n_n5142 = (((!i_7_) & (!i_8_) & (!i_6_) & (x12x) & (n_n500)));
	assign n_n5107 = (((!i_9_) & (n_n524) & (n_n518) & (n_n130)));
	assign n_n5130 = (((i_7_) & (!i_8_) & (i_6_) & (x12x) & (n_n500)));
	assign n_n5123 = (((!i_9_) & (n_n524) & (n_n509) & (n_n130)));
	assign n_n5129 = (((!i_9_) & (n_n534) & (n_n130) & (n_n500)));
	assign n_n5145 = (((!i_9_) & (n_n534) & (n_n491) & (n_n130)));
	assign n_n5156 = (((!i_7_) & (i_8_) & (!i_6_) & (n_n491) & (x12x)));
	assign x13696x = (((!n_n5142) & (!n_n5107) & (!n_n5130) & (n_n5123)) + ((!n_n5142) & (!n_n5107) & (n_n5130) & (!n_n5123)) + ((!n_n5142) & (!n_n5107) & (n_n5130) & (n_n5123)) + ((!n_n5142) & (n_n5107) & (!n_n5130) & (!n_n5123)) + ((!n_n5142) & (n_n5107) & (!n_n5130) & (n_n5123)) + ((!n_n5142) & (n_n5107) & (n_n5130) & (!n_n5123)) + ((!n_n5142) & (n_n5107) & (n_n5130) & (n_n5123)) + ((n_n5142) & (!n_n5107) & (!n_n5130) & (!n_n5123)) + ((n_n5142) & (!n_n5107) & (!n_n5130) & (n_n5123)) + ((n_n5142) & (!n_n5107) & (n_n5130) & (!n_n5123)) + ((n_n5142) & (!n_n5107) & (n_n5130) & (n_n5123)) + ((n_n5142) & (n_n5107) & (!n_n5130) & (!n_n5123)) + ((n_n5142) & (n_n5107) & (!n_n5130) & (n_n5123)) + ((n_n5142) & (n_n5107) & (n_n5130) & (!n_n5123)) + ((n_n5142) & (n_n5107) & (n_n5130) & (n_n5123)));
	assign x13697x = (((!n_n5101) & (!n_n5110) & (!n_n5129) & (!n_n5145) & (n_n5156)) + ((!n_n5101) & (!n_n5110) & (!n_n5129) & (n_n5145) & (!n_n5156)) + ((!n_n5101) & (!n_n5110) & (!n_n5129) & (n_n5145) & (n_n5156)) + ((!n_n5101) & (!n_n5110) & (n_n5129) & (!n_n5145) & (!n_n5156)) + ((!n_n5101) & (!n_n5110) & (n_n5129) & (!n_n5145) & (n_n5156)) + ((!n_n5101) & (!n_n5110) & (n_n5129) & (n_n5145) & (!n_n5156)) + ((!n_n5101) & (!n_n5110) & (n_n5129) & (n_n5145) & (n_n5156)) + ((!n_n5101) & (n_n5110) & (!n_n5129) & (!n_n5145) & (!n_n5156)) + ((!n_n5101) & (n_n5110) & (!n_n5129) & (!n_n5145) & (n_n5156)) + ((!n_n5101) & (n_n5110) & (!n_n5129) & (n_n5145) & (!n_n5156)) + ((!n_n5101) & (n_n5110) & (!n_n5129) & (n_n5145) & (n_n5156)) + ((!n_n5101) & (n_n5110) & (n_n5129) & (!n_n5145) & (!n_n5156)) + ((!n_n5101) & (n_n5110) & (n_n5129) & (!n_n5145) & (n_n5156)) + ((!n_n5101) & (n_n5110) & (n_n5129) & (n_n5145) & (!n_n5156)) + ((!n_n5101) & (n_n5110) & (n_n5129) & (n_n5145) & (n_n5156)) + ((n_n5101) & (!n_n5110) & (!n_n5129) & (!n_n5145) & (!n_n5156)) + ((n_n5101) & (!n_n5110) & (!n_n5129) & (!n_n5145) & (n_n5156)) + ((n_n5101) & (!n_n5110) & (!n_n5129) & (n_n5145) & (!n_n5156)) + ((n_n5101) & (!n_n5110) & (!n_n5129) & (n_n5145) & (n_n5156)) + ((n_n5101) & (!n_n5110) & (n_n5129) & (!n_n5145) & (!n_n5156)) + ((n_n5101) & (!n_n5110) & (n_n5129) & (!n_n5145) & (n_n5156)) + ((n_n5101) & (!n_n5110) & (n_n5129) & (n_n5145) & (!n_n5156)) + ((n_n5101) & (!n_n5110) & (n_n5129) & (n_n5145) & (n_n5156)) + ((n_n5101) & (n_n5110) & (!n_n5129) & (!n_n5145) & (!n_n5156)) + ((n_n5101) & (n_n5110) & (!n_n5129) & (!n_n5145) & (n_n5156)) + ((n_n5101) & (n_n5110) & (!n_n5129) & (n_n5145) & (!n_n5156)) + ((n_n5101) & (n_n5110) & (!n_n5129) & (n_n5145) & (n_n5156)) + ((n_n5101) & (n_n5110) & (n_n5129) & (!n_n5145) & (!n_n5156)) + ((n_n5101) & (n_n5110) & (n_n5129) & (!n_n5145) & (n_n5156)) + ((n_n5101) & (n_n5110) & (n_n5129) & (n_n5145) & (!n_n5156)) + ((n_n5101) & (n_n5110) & (n_n5129) & (n_n5145) & (n_n5156)));
	assign n_n4318 = (((i_9_) & (n_n536) & (n_n528) & (n_n535)));
	assign n_n4385 = (((!i_9_) & (n_n536) & (n_n526) & (n_n491)));
	assign n_n4455 = (((i_1_) & (!i_2_) & (i_0_) & (n_n535) & (x23x)));
	assign n_n4513 = (((!i_9_) & (n_n526) & (n_n455) & (n_n491)));
	assign n_n4515 = (((!i_9_) & (n_n524) & (n_n455) & (n_n491)));
	assign n_n4790 = (((i_9_) & (n_n482) & (n_n325) & (n_n520)));
	assign n_n4791 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n325) & (x23x)));
	assign n_n4787 = (((!i_9_) & (n_n524) & (n_n482) & (n_n325)));
	assign n_n4860 = (((i_9_) & (n_n509) & (n_n260) & (n_n530)));
	assign n_n4926 = (((i_9_) & (n_n528) & (n_n473) & (n_n260)));
	assign n_n4928 = (((i_9_) & (n_n526) & (n_n473) & (n_n260)));
	assign n_n4925 = (((!i_9_) & (n_n473) & (n_n260) & (n_n530)));
	assign n_n4988 = (((i_9_) & (n_n509) & (n_n195) & (n_n530)));
	assign n_n4987 = (((!i_9_) & (n_n532) & (n_n509) & (n_n195)));
	assign n_n5041 = (((!i_9_) & (n_n526) & (n_n482) & (n_n195)));
	assign n_n5042 = (((i_9_) & (n_n524) & (n_n482) & (n_n195)));
	assign n_n5100 = (((!i_5_) & (i_3_) & (i_4_) & (x12x) & (n_n530)));
	assign n_n4724 = (((i_9_) & (n_n518) & (n_n325) & (n_n522)));
	assign n_n4734 = (((i_9_) & (n_n528) & (n_n509) & (n_n325)));
	assign x95x = (((!i_9_) & (n_n528) & (n_n509) & (n_n325)) + ((i_9_) & (n_n528) & (n_n509) & (n_n325)));
	assign n_n4726 = (((i_9_) & (n_n518) & (n_n325) & (n_n520)));
	assign x101x = (((!i_9_) & (n_n518) & (n_n325) & (!n_n520) & (x20x)) + ((!i_9_) & (n_n518) & (n_n325) & (n_n520) & (x20x)) + ((i_9_) & (n_n518) & (n_n325) & (!n_n520) & (x20x)) + ((i_9_) & (n_n518) & (n_n325) & (n_n520) & (!x20x)) + ((i_9_) & (n_n518) & (n_n325) & (n_n520) & (x20x)));
	assign n_n4728 = (((i_9_) & (n_n534) & (n_n509) & (n_n325)));
	assign x244x = (((i_7_) & (!i_8_) & (i_6_) & (n_n509) & (x14x)) + ((i_7_) & (i_8_) & (i_6_) & (n_n509) & (x14x)));
	assign x15745x = (((!i_9_) & (!n_n524) & (n_n528) & (n_n509) & (n_n325)) + ((!i_9_) & (n_n524) & (!n_n528) & (n_n509) & (n_n325)) + ((!i_9_) & (n_n524) & (n_n528) & (n_n509) & (n_n325)) + ((i_9_) & (!n_n524) & (n_n528) & (n_n509) & (n_n325)) + ((i_9_) & (n_n524) & (n_n528) & (n_n509) & (n_n325)));
	assign n_n2981 = (((!n_n4724) & (!n_n4727) & (!x101x) & (!x244x) & (x15745x)) + ((!n_n4724) & (!n_n4727) & (!x101x) & (x244x) & (!x15745x)) + ((!n_n4724) & (!n_n4727) & (!x101x) & (x244x) & (x15745x)) + ((!n_n4724) & (!n_n4727) & (x101x) & (!x244x) & (!x15745x)) + ((!n_n4724) & (!n_n4727) & (x101x) & (!x244x) & (x15745x)) + ((!n_n4724) & (!n_n4727) & (x101x) & (x244x) & (!x15745x)) + ((!n_n4724) & (!n_n4727) & (x101x) & (x244x) & (x15745x)) + ((!n_n4724) & (n_n4727) & (!x101x) & (!x244x) & (!x15745x)) + ((!n_n4724) & (n_n4727) & (!x101x) & (!x244x) & (x15745x)) + ((!n_n4724) & (n_n4727) & (!x101x) & (x244x) & (!x15745x)) + ((!n_n4724) & (n_n4727) & (!x101x) & (x244x) & (x15745x)) + ((!n_n4724) & (n_n4727) & (x101x) & (!x244x) & (!x15745x)) + ((!n_n4724) & (n_n4727) & (x101x) & (!x244x) & (x15745x)) + ((!n_n4724) & (n_n4727) & (x101x) & (x244x) & (!x15745x)) + ((!n_n4724) & (n_n4727) & (x101x) & (x244x) & (x15745x)) + ((n_n4724) & (!n_n4727) & (!x101x) & (!x244x) & (!x15745x)) + ((n_n4724) & (!n_n4727) & (!x101x) & (!x244x) & (x15745x)) + ((n_n4724) & (!n_n4727) & (!x101x) & (x244x) & (!x15745x)) + ((n_n4724) & (!n_n4727) & (!x101x) & (x244x) & (x15745x)) + ((n_n4724) & (!n_n4727) & (x101x) & (!x244x) & (!x15745x)) + ((n_n4724) & (!n_n4727) & (x101x) & (!x244x) & (x15745x)) + ((n_n4724) & (!n_n4727) & (x101x) & (x244x) & (!x15745x)) + ((n_n4724) & (!n_n4727) & (x101x) & (x244x) & (x15745x)) + ((n_n4724) & (n_n4727) & (!x101x) & (!x244x) & (!x15745x)) + ((n_n4724) & (n_n4727) & (!x101x) & (!x244x) & (x15745x)) + ((n_n4724) & (n_n4727) & (!x101x) & (x244x) & (!x15745x)) + ((n_n4724) & (n_n4727) & (!x101x) & (x244x) & (x15745x)) + ((n_n4724) & (n_n4727) & (x101x) & (!x244x) & (!x15745x)) + ((n_n4724) & (n_n4727) & (x101x) & (!x244x) & (x15745x)) + ((n_n4724) & (n_n4727) & (x101x) & (x244x) & (!x15745x)) + ((n_n4724) & (n_n4727) & (x101x) & (x244x) & (x15745x)));
	assign n_n4868 = (((i_9_) & (n_n509) & (n_n260) & (n_n522)));
	assign n_n4861 = (((!i_9_) & (n_n509) & (n_n260) & (n_n530)));
	assign x246x = (((!i_9_) & (!n_n528) & (n_n509) & (n_n260) & (n_n530)) + ((!i_9_) & (n_n528) & (n_n509) & (n_n260) & (n_n530)) + ((i_9_) & (n_n528) & (n_n509) & (n_n260) & (!n_n530)) + ((i_9_) & (n_n528) & (n_n509) & (n_n260) & (n_n530)));
	assign n_n4869 = (((i_5_) & (i_3_) & (!i_4_) & (n_n260) & (x20x)));
	assign n_n4870 = (((i_9_) & (n_n509) & (n_n260) & (n_n520)));
	assign x294x = (((!i_9_) & (n_n509) & (n_n260) & (!n_n520) & (x20x)) + ((!i_9_) & (n_n509) & (n_n260) & (n_n520) & (x20x)) + ((i_9_) & (n_n509) & (n_n260) & (!n_n520) & (x20x)) + ((i_9_) & (n_n509) & (n_n260) & (n_n520) & (!x20x)) + ((i_9_) & (n_n509) & (n_n260) & (n_n520) & (x20x)));
	assign x15678x = (((!i_7_) & (i_8_) & (i_6_) & (n_n509) & (x17x)) + ((i_7_) & (i_8_) & (!i_6_) & (n_n509) & (x17x)));
	assign n_n2970 = (((!x245x) & (!n_n4868) & (!x246x) & (!x294x) & (x15678x)) + ((!x245x) & (!n_n4868) & (!x246x) & (x294x) & (!x15678x)) + ((!x245x) & (!n_n4868) & (!x246x) & (x294x) & (x15678x)) + ((!x245x) & (!n_n4868) & (x246x) & (!x294x) & (!x15678x)) + ((!x245x) & (!n_n4868) & (x246x) & (!x294x) & (x15678x)) + ((!x245x) & (!n_n4868) & (x246x) & (x294x) & (!x15678x)) + ((!x245x) & (!n_n4868) & (x246x) & (x294x) & (x15678x)) + ((!x245x) & (n_n4868) & (!x246x) & (!x294x) & (!x15678x)) + ((!x245x) & (n_n4868) & (!x246x) & (!x294x) & (x15678x)) + ((!x245x) & (n_n4868) & (!x246x) & (x294x) & (!x15678x)) + ((!x245x) & (n_n4868) & (!x246x) & (x294x) & (x15678x)) + ((!x245x) & (n_n4868) & (x246x) & (!x294x) & (!x15678x)) + ((!x245x) & (n_n4868) & (x246x) & (!x294x) & (x15678x)) + ((!x245x) & (n_n4868) & (x246x) & (x294x) & (!x15678x)) + ((!x245x) & (n_n4868) & (x246x) & (x294x) & (x15678x)) + ((x245x) & (!n_n4868) & (!x246x) & (!x294x) & (!x15678x)) + ((x245x) & (!n_n4868) & (!x246x) & (!x294x) & (x15678x)) + ((x245x) & (!n_n4868) & (!x246x) & (x294x) & (!x15678x)) + ((x245x) & (!n_n4868) & (!x246x) & (x294x) & (x15678x)) + ((x245x) & (!n_n4868) & (x246x) & (!x294x) & (!x15678x)) + ((x245x) & (!n_n4868) & (x246x) & (!x294x) & (x15678x)) + ((x245x) & (!n_n4868) & (x246x) & (x294x) & (!x15678x)) + ((x245x) & (!n_n4868) & (x246x) & (x294x) & (x15678x)) + ((x245x) & (n_n4868) & (!x246x) & (!x294x) & (!x15678x)) + ((x245x) & (n_n4868) & (!x246x) & (!x294x) & (x15678x)) + ((x245x) & (n_n4868) & (!x246x) & (x294x) & (!x15678x)) + ((x245x) & (n_n4868) & (!x246x) & (x294x) & (x15678x)) + ((x245x) & (n_n4868) & (x246x) & (!x294x) & (!x15678x)) + ((x245x) & (n_n4868) & (x246x) & (!x294x) & (x15678x)) + ((x245x) & (n_n4868) & (x246x) & (x294x) & (!x15678x)) + ((x245x) & (n_n4868) & (x246x) & (x294x) & (x15678x)));
	assign n_n5018 = (((i_9_) & (n_n532) & (n_n491) & (n_n195)));
	assign n_n5022 = (((i_9_) & (n_n528) & (n_n491) & (n_n195)));
	assign n_n5017 = (((!i_9_) & (n_n534) & (n_n491) & (n_n195)));
	assign n_n5014 = (((i_9_) & (n_n520) & (n_n195) & (n_n500)));
	assign n_n5015 = (((i_1_) & (!i_2_) & (!i_0_) & (x23x) & (n_n500)));
	assign n_n5023 = (((!i_9_) & (n_n528) & (n_n491) & (n_n195)));
	assign n_n5021 = (((!i_9_) & (n_n491) & (n_n195) & (n_n530)));
	assign x296x = (((!i_9_) & (!n_n528) & (n_n491) & (n_n195) & (n_n530)) + ((!i_9_) & (n_n528) & (n_n491) & (n_n195) & (!n_n530)) + ((!i_9_) & (n_n528) & (n_n491) & (n_n195) & (n_n530)));
	assign n_n5019 = (((!i_9_) & (n_n532) & (n_n491) & (n_n195)));
	assign n_n5020 = (((i_9_) & (n_n491) & (n_n195) & (n_n530)));
	assign x298x = (((!i_9_) & (n_n532) & (n_n491) & (n_n195) & (!n_n530)) + ((!i_9_) & (n_n532) & (n_n491) & (n_n195) & (n_n530)) + ((i_9_) & (!n_n532) & (n_n491) & (n_n195) & (n_n530)) + ((i_9_) & (n_n532) & (n_n491) & (n_n195) & (n_n530)));
	assign x15705x = (((!n_n5018) & (!n_n5022) & (!n_n5017) & (!n_n5014) & (n_n5015)) + ((!n_n5018) & (!n_n5022) & (!n_n5017) & (n_n5014) & (!n_n5015)) + ((!n_n5018) & (!n_n5022) & (!n_n5017) & (n_n5014) & (n_n5015)) + ((!n_n5018) & (!n_n5022) & (n_n5017) & (!n_n5014) & (!n_n5015)) + ((!n_n5018) & (!n_n5022) & (n_n5017) & (!n_n5014) & (n_n5015)) + ((!n_n5018) & (!n_n5022) & (n_n5017) & (n_n5014) & (!n_n5015)) + ((!n_n5018) & (!n_n5022) & (n_n5017) & (n_n5014) & (n_n5015)) + ((!n_n5018) & (n_n5022) & (!n_n5017) & (!n_n5014) & (!n_n5015)) + ((!n_n5018) & (n_n5022) & (!n_n5017) & (!n_n5014) & (n_n5015)) + ((!n_n5018) & (n_n5022) & (!n_n5017) & (n_n5014) & (!n_n5015)) + ((!n_n5018) & (n_n5022) & (!n_n5017) & (n_n5014) & (n_n5015)) + ((!n_n5018) & (n_n5022) & (n_n5017) & (!n_n5014) & (!n_n5015)) + ((!n_n5018) & (n_n5022) & (n_n5017) & (!n_n5014) & (n_n5015)) + ((!n_n5018) & (n_n5022) & (n_n5017) & (n_n5014) & (!n_n5015)) + ((!n_n5018) & (n_n5022) & (n_n5017) & (n_n5014) & (n_n5015)) + ((n_n5018) & (!n_n5022) & (!n_n5017) & (!n_n5014) & (!n_n5015)) + ((n_n5018) & (!n_n5022) & (!n_n5017) & (!n_n5014) & (n_n5015)) + ((n_n5018) & (!n_n5022) & (!n_n5017) & (n_n5014) & (!n_n5015)) + ((n_n5018) & (!n_n5022) & (!n_n5017) & (n_n5014) & (n_n5015)) + ((n_n5018) & (!n_n5022) & (n_n5017) & (!n_n5014) & (!n_n5015)) + ((n_n5018) & (!n_n5022) & (n_n5017) & (!n_n5014) & (n_n5015)) + ((n_n5018) & (!n_n5022) & (n_n5017) & (n_n5014) & (!n_n5015)) + ((n_n5018) & (!n_n5022) & (n_n5017) & (n_n5014) & (n_n5015)) + ((n_n5018) & (n_n5022) & (!n_n5017) & (!n_n5014) & (!n_n5015)) + ((n_n5018) & (n_n5022) & (!n_n5017) & (!n_n5014) & (n_n5015)) + ((n_n5018) & (n_n5022) & (!n_n5017) & (n_n5014) & (!n_n5015)) + ((n_n5018) & (n_n5022) & (!n_n5017) & (n_n5014) & (n_n5015)) + ((n_n5018) & (n_n5022) & (n_n5017) & (!n_n5014) & (!n_n5015)) + ((n_n5018) & (n_n5022) & (n_n5017) & (!n_n5014) & (n_n5015)) + ((n_n5018) & (n_n5022) & (n_n5017) & (n_n5014) & (!n_n5015)) + ((n_n5018) & (n_n5022) & (n_n5017) & (n_n5014) & (n_n5015)));
	assign n_n4993 = (((!i_9_) & (n_n526) & (n_n509) & (n_n195)));
	assign n_n4994 = (((i_9_) & (n_n524) & (n_n509) & (n_n195)));
	assign n_n1576 = (((!i_9_) & (n_n524) & (n_n509) & (!n_n522) & (n_n195)) + ((!i_9_) & (n_n524) & (n_n509) & (n_n522) & (n_n195)) + ((i_9_) & (!n_n524) & (n_n509) & (n_n522) & (n_n195)) + ((i_9_) & (n_n524) & (n_n509) & (!n_n522) & (n_n195)) + ((i_9_) & (n_n524) & (n_n509) & (n_n522) & (n_n195)));
	assign n_n4989 = (((!i_9_) & (n_n509) & (n_n195) & (n_n530)));
	assign x134x = (((!i_9_) & (n_n509) & (n_n195) & (n_n530)) + ((i_9_) & (n_n509) & (n_n195) & (n_n530)));
	assign n_n4980 = (((i_9_) & (n_n518) & (n_n522) & (n_n195)));
	assign x252x = (((!i_7_) & (!i_8_) & (!i_6_) & (n_n518) & (x18x)) + ((!i_7_) & (i_8_) & (!i_6_) & (n_n518) & (x18x)));
	assign n_n5005 = (((!i_9_) & (n_n195) & (n_n500) & (n_n530)));
	assign n_n5004 = (((i_9_) & (n_n195) & (n_n500) & (n_n530)));
	assign n_n5006 = (((i_9_) & (n_n528) & (n_n195) & (n_n500)));
	assign n_n5007 = (((!i_9_) & (n_n528) & (n_n195) & (n_n500)));
	assign x136x = (((!i_9_) & (n_n528) & (n_n195) & (n_n500)) + ((i_9_) & (n_n528) & (n_n195) & (n_n500)));
	assign x247x = (((!i_9_) & (n_n509) & (!n_n520) & (n_n195) & (x20x)) + ((!i_9_) & (n_n509) & (n_n520) & (n_n195) & (x20x)) + ((i_9_) & (n_n509) & (!n_n520) & (n_n195) & (x20x)) + ((i_9_) & (n_n509) & (n_n520) & (n_n195) & (!x20x)) + ((i_9_) & (n_n509) & (n_n520) & (n_n195) & (x20x)));
	assign n_n5003 = (((!i_9_) & (n_n532) & (n_n195) & (n_n500)));
	assign n_n5002 = (((i_9_) & (n_n532) & (n_n195) & (n_n500)));
	assign x393x = (((!i_9_) & (n_n532) & (n_n195) & (n_n500)) + ((i_9_) & (n_n532) & (n_n195) & (n_n500)));
	assign x14940x = (((!i_9_) & (n_n195) & (n_n500) & (n_n530)) + ((i_9_) & (n_n195) & (n_n500) & (n_n530)));
	assign n_n4907 = (((!i_9_) & (n_n482) & (n_n532) & (n_n260)));
	assign n_n4913 = (((!i_9_) & (n_n526) & (n_n482) & (n_n260)));
	assign n_n4922 = (((i_9_) & (n_n473) & (n_n532) & (n_n260)));
	assign x371x = (((!i_9_) & (!n_n473) & (!n_n534) & (!n_n195) & (n_n5047)) + ((!i_9_) & (!n_n473) & (!n_n534) & (n_n195) & (n_n5047)) + ((!i_9_) & (!n_n473) & (n_n534) & (!n_n195) & (n_n5047)) + ((!i_9_) & (!n_n473) & (n_n534) & (n_n195) & (n_n5047)) + ((!i_9_) & (n_n473) & (!n_n534) & (!n_n195) & (n_n5047)) + ((!i_9_) & (n_n473) & (!n_n534) & (n_n195) & (n_n5047)) + ((!i_9_) & (n_n473) & (n_n534) & (!n_n195) & (n_n5047)) + ((!i_9_) & (n_n473) & (n_n534) & (n_n195) & (n_n5047)) + ((i_9_) & (!n_n473) & (!n_n534) & (!n_n195) & (n_n5047)) + ((i_9_) & (!n_n473) & (!n_n534) & (n_n195) & (n_n5047)) + ((i_9_) & (!n_n473) & (n_n534) & (!n_n195) & (n_n5047)) + ((i_9_) & (!n_n473) & (n_n534) & (n_n195) & (n_n5047)) + ((i_9_) & (n_n473) & (!n_n534) & (!n_n195) & (n_n5047)) + ((i_9_) & (n_n473) & (!n_n534) & (n_n195) & (n_n5047)) + ((i_9_) & (n_n473) & (n_n534) & (!n_n195) & (n_n5047)) + ((i_9_) & (n_n473) & (n_n534) & (n_n195) & (!n_n5047)) + ((i_9_) & (n_n473) & (n_n534) & (n_n195) & (n_n5047)));
	assign x97x = (((!i_9_) & (n_n526) & (n_n482) & (n_n195)) + ((i_9_) & (n_n526) & (n_n482) & (n_n195)));
	assign x14793x = (((!i_9_) & (n_n482) & (!n_n532) & (n_n195) & (x20x)) + ((!i_9_) & (n_n482) & (n_n532) & (n_n195) & (!x20x)) + ((!i_9_) & (n_n482) & (n_n532) & (n_n195) & (x20x)) + ((i_9_) & (n_n482) & (!n_n532) & (n_n195) & (x20x)) + ((i_9_) & (n_n482) & (n_n532) & (n_n195) & (!x20x)) + ((i_9_) & (n_n482) & (n_n532) & (n_n195) & (x20x)));
	assign x155x = (((!i_9_) & (!n_n532) & (!n_n130) & (!n_n500) & (n_n5132)) + ((!i_9_) & (!n_n532) & (!n_n130) & (n_n500) & (n_n5132)) + ((!i_9_) & (!n_n532) & (n_n130) & (!n_n500) & (n_n5132)) + ((!i_9_) & (!n_n532) & (n_n130) & (n_n500) & (n_n5132)) + ((!i_9_) & (n_n532) & (!n_n130) & (!n_n500) & (n_n5132)) + ((!i_9_) & (n_n532) & (!n_n130) & (n_n500) & (n_n5132)) + ((!i_9_) & (n_n532) & (n_n130) & (!n_n500) & (n_n5132)) + ((!i_9_) & (n_n532) & (n_n130) & (n_n500) & (!n_n5132)) + ((!i_9_) & (n_n532) & (n_n130) & (n_n500) & (n_n5132)) + ((i_9_) & (!n_n532) & (!n_n130) & (!n_n500) & (n_n5132)) + ((i_9_) & (!n_n532) & (!n_n130) & (n_n500) & (n_n5132)) + ((i_9_) & (!n_n532) & (n_n130) & (!n_n500) & (n_n5132)) + ((i_9_) & (!n_n532) & (n_n130) & (n_n500) & (n_n5132)) + ((i_9_) & (n_n532) & (!n_n130) & (!n_n500) & (n_n5132)) + ((i_9_) & (n_n532) & (!n_n130) & (n_n500) & (n_n5132)) + ((i_9_) & (n_n532) & (n_n130) & (!n_n500) & (n_n5132)) + ((i_9_) & (n_n532) & (n_n130) & (n_n500) & (n_n5132)));
	assign x143x = (((!i_9_) & (!n_n528) & (!n_n535) & (!n_n130) & (n_n5088)) + ((!i_9_) & (!n_n528) & (!n_n535) & (n_n130) & (n_n5088)) + ((!i_9_) & (!n_n528) & (n_n535) & (!n_n130) & (n_n5088)) + ((!i_9_) & (!n_n528) & (n_n535) & (n_n130) & (n_n5088)) + ((!i_9_) & (n_n528) & (!n_n535) & (!n_n130) & (n_n5088)) + ((!i_9_) & (n_n528) & (!n_n535) & (n_n130) & (n_n5088)) + ((!i_9_) & (n_n528) & (n_n535) & (!n_n130) & (n_n5088)) + ((!i_9_) & (n_n528) & (n_n535) & (n_n130) & (!n_n5088)) + ((!i_9_) & (n_n528) & (n_n535) & (n_n130) & (n_n5088)) + ((i_9_) & (!n_n528) & (!n_n535) & (!n_n130) & (n_n5088)) + ((i_9_) & (!n_n528) & (!n_n535) & (n_n130) & (n_n5088)) + ((i_9_) & (!n_n528) & (n_n535) & (!n_n130) & (n_n5088)) + ((i_9_) & (!n_n528) & (n_n535) & (n_n130) & (n_n5088)) + ((i_9_) & (n_n528) & (!n_n535) & (!n_n130) & (n_n5088)) + ((i_9_) & (n_n528) & (!n_n535) & (n_n130) & (n_n5088)) + ((i_9_) & (n_n528) & (n_n535) & (!n_n130) & (n_n5088)) + ((i_9_) & (n_n528) & (n_n535) & (n_n130) & (n_n5088)));
	assign x14785x = (((!n_n5113) & (!n_n5081) & (!n_n5098) & (!n_n5104) & (n_n5095)) + ((!n_n5113) & (!n_n5081) & (!n_n5098) & (n_n5104) & (!n_n5095)) + ((!n_n5113) & (!n_n5081) & (!n_n5098) & (n_n5104) & (n_n5095)) + ((!n_n5113) & (!n_n5081) & (n_n5098) & (!n_n5104) & (!n_n5095)) + ((!n_n5113) & (!n_n5081) & (n_n5098) & (!n_n5104) & (n_n5095)) + ((!n_n5113) & (!n_n5081) & (n_n5098) & (n_n5104) & (!n_n5095)) + ((!n_n5113) & (!n_n5081) & (n_n5098) & (n_n5104) & (n_n5095)) + ((!n_n5113) & (n_n5081) & (!n_n5098) & (!n_n5104) & (!n_n5095)) + ((!n_n5113) & (n_n5081) & (!n_n5098) & (!n_n5104) & (n_n5095)) + ((!n_n5113) & (n_n5081) & (!n_n5098) & (n_n5104) & (!n_n5095)) + ((!n_n5113) & (n_n5081) & (!n_n5098) & (n_n5104) & (n_n5095)) + ((!n_n5113) & (n_n5081) & (n_n5098) & (!n_n5104) & (!n_n5095)) + ((!n_n5113) & (n_n5081) & (n_n5098) & (!n_n5104) & (n_n5095)) + ((!n_n5113) & (n_n5081) & (n_n5098) & (n_n5104) & (!n_n5095)) + ((!n_n5113) & (n_n5081) & (n_n5098) & (n_n5104) & (n_n5095)) + ((n_n5113) & (!n_n5081) & (!n_n5098) & (!n_n5104) & (!n_n5095)) + ((n_n5113) & (!n_n5081) & (!n_n5098) & (!n_n5104) & (n_n5095)) + ((n_n5113) & (!n_n5081) & (!n_n5098) & (n_n5104) & (!n_n5095)) + ((n_n5113) & (!n_n5081) & (!n_n5098) & (n_n5104) & (n_n5095)) + ((n_n5113) & (!n_n5081) & (n_n5098) & (!n_n5104) & (!n_n5095)) + ((n_n5113) & (!n_n5081) & (n_n5098) & (!n_n5104) & (n_n5095)) + ((n_n5113) & (!n_n5081) & (n_n5098) & (n_n5104) & (!n_n5095)) + ((n_n5113) & (!n_n5081) & (n_n5098) & (n_n5104) & (n_n5095)) + ((n_n5113) & (n_n5081) & (!n_n5098) & (!n_n5104) & (!n_n5095)) + ((n_n5113) & (n_n5081) & (!n_n5098) & (!n_n5104) & (n_n5095)) + ((n_n5113) & (n_n5081) & (!n_n5098) & (n_n5104) & (!n_n5095)) + ((n_n5113) & (n_n5081) & (!n_n5098) & (n_n5104) & (n_n5095)) + ((n_n5113) & (n_n5081) & (n_n5098) & (!n_n5104) & (!n_n5095)) + ((n_n5113) & (n_n5081) & (n_n5098) & (!n_n5104) & (n_n5095)) + ((n_n5113) & (n_n5081) & (n_n5098) & (n_n5104) & (!n_n5095)) + ((n_n5113) & (n_n5081) & (n_n5098) & (n_n5104) & (n_n5095)));
	assign x14790x = (((!n_n5174) & (!n_n5184) & (!n_n5212) & (n_n5172)) + ((!n_n5174) & (!n_n5184) & (n_n5212) & (!n_n5172)) + ((!n_n5174) & (!n_n5184) & (n_n5212) & (n_n5172)) + ((!n_n5174) & (n_n5184) & (!n_n5212) & (!n_n5172)) + ((!n_n5174) & (n_n5184) & (!n_n5212) & (n_n5172)) + ((!n_n5174) & (n_n5184) & (n_n5212) & (!n_n5172)) + ((!n_n5174) & (n_n5184) & (n_n5212) & (n_n5172)) + ((n_n5174) & (!n_n5184) & (!n_n5212) & (!n_n5172)) + ((n_n5174) & (!n_n5184) & (!n_n5212) & (n_n5172)) + ((n_n5174) & (!n_n5184) & (n_n5212) & (!n_n5172)) + ((n_n5174) & (!n_n5184) & (n_n5212) & (n_n5172)) + ((n_n5174) & (n_n5184) & (!n_n5212) & (!n_n5172)) + ((n_n5174) & (n_n5184) & (!n_n5212) & (n_n5172)) + ((n_n5174) & (n_n5184) & (n_n5212) & (!n_n5172)) + ((n_n5174) & (n_n5184) & (n_n5212) & (n_n5172)));
	assign x14791x = (((!x12x) & (!x572x) & (!n_n5170) & (!n_n5234) & (x385x)) + ((!x12x) & (!x572x) & (!n_n5170) & (n_n5234) & (!x385x)) + ((!x12x) & (!x572x) & (!n_n5170) & (n_n5234) & (x385x)) + ((!x12x) & (!x572x) & (n_n5170) & (!n_n5234) & (!x385x)) + ((!x12x) & (!x572x) & (n_n5170) & (!n_n5234) & (x385x)) + ((!x12x) & (!x572x) & (n_n5170) & (n_n5234) & (!x385x)) + ((!x12x) & (!x572x) & (n_n5170) & (n_n5234) & (x385x)) + ((!x12x) & (x572x) & (!n_n5170) & (!n_n5234) & (x385x)) + ((!x12x) & (x572x) & (!n_n5170) & (n_n5234) & (!x385x)) + ((!x12x) & (x572x) & (!n_n5170) & (n_n5234) & (x385x)) + ((!x12x) & (x572x) & (n_n5170) & (!n_n5234) & (!x385x)) + ((!x12x) & (x572x) & (n_n5170) & (!n_n5234) & (x385x)) + ((!x12x) & (x572x) & (n_n5170) & (n_n5234) & (!x385x)) + ((!x12x) & (x572x) & (n_n5170) & (n_n5234) & (x385x)) + ((x12x) & (!x572x) & (!n_n5170) & (!n_n5234) & (x385x)) + ((x12x) & (!x572x) & (!n_n5170) & (n_n5234) & (!x385x)) + ((x12x) & (!x572x) & (!n_n5170) & (n_n5234) & (x385x)) + ((x12x) & (!x572x) & (n_n5170) & (!n_n5234) & (!x385x)) + ((x12x) & (!x572x) & (n_n5170) & (!n_n5234) & (x385x)) + ((x12x) & (!x572x) & (n_n5170) & (n_n5234) & (!x385x)) + ((x12x) & (!x572x) & (n_n5170) & (n_n5234) & (x385x)) + ((x12x) & (x572x) & (!n_n5170) & (!n_n5234) & (!x385x)) + ((x12x) & (x572x) & (!n_n5170) & (!n_n5234) & (x385x)) + ((x12x) & (x572x) & (!n_n5170) & (n_n5234) & (!x385x)) + ((x12x) & (x572x) & (!n_n5170) & (n_n5234) & (x385x)) + ((x12x) & (x572x) & (n_n5170) & (!n_n5234) & (!x385x)) + ((x12x) & (x572x) & (n_n5170) & (!n_n5234) & (x385x)) + ((x12x) & (x572x) & (n_n5170) & (n_n5234) & (!x385x)) + ((x12x) & (x572x) & (n_n5170) & (n_n5234) & (x385x)));
	assign n_n4934 = (((i_9_) & (n_n473) & (n_n260) & (n_n520)));
	assign n_n5324 = (((!i_7_) & (i_8_) & (i_6_) & (x19x) & (n_n464)));
	assign n_n5335 = (((!i_5_) & (!i_3_) & (!i_4_) & (x23x) & (n_n65)));
	assign x14807x = (((!n_n5296) & (!n_n5320) & (!n_n5324) & (n_n5335)) + ((!n_n5296) & (!n_n5320) & (n_n5324) & (!n_n5335)) + ((!n_n5296) & (!n_n5320) & (n_n5324) & (n_n5335)) + ((!n_n5296) & (n_n5320) & (!n_n5324) & (!n_n5335)) + ((!n_n5296) & (n_n5320) & (!n_n5324) & (n_n5335)) + ((!n_n5296) & (n_n5320) & (n_n5324) & (!n_n5335)) + ((!n_n5296) & (n_n5320) & (n_n5324) & (n_n5335)) + ((n_n5296) & (!n_n5320) & (!n_n5324) & (!n_n5335)) + ((n_n5296) & (!n_n5320) & (!n_n5324) & (n_n5335)) + ((n_n5296) & (!n_n5320) & (n_n5324) & (!n_n5335)) + ((n_n5296) & (!n_n5320) & (n_n5324) & (n_n5335)) + ((n_n5296) & (n_n5320) & (!n_n5324) & (!n_n5335)) + ((n_n5296) & (n_n5320) & (!n_n5324) & (n_n5335)) + ((n_n5296) & (n_n5320) & (n_n5324) & (!n_n5335)) + ((n_n5296) & (n_n5320) & (n_n5324) & (n_n5335)));
	assign x531x = (((i_1_) & (i_2_) & (!i_0_) & (n_n464)));
	assign n_n5010 = (((i_9_) & (n_n524) & (n_n195) & (n_n500)));
	assign n_n4967 = (((i_5_) & (i_3_) & (i_4_) & (n_n195) & (x23x)));
	assign x14813x = (((!x23x) & (!n_n5015) & (!x531x) & (!n_n5010) & (n_n4967)) + ((!x23x) & (!n_n5015) & (!x531x) & (n_n5010) & (!n_n4967)) + ((!x23x) & (!n_n5015) & (!x531x) & (n_n5010) & (n_n4967)) + ((!x23x) & (!n_n5015) & (x531x) & (!n_n5010) & (n_n4967)) + ((!x23x) & (!n_n5015) & (x531x) & (n_n5010) & (!n_n4967)) + ((!x23x) & (!n_n5015) & (x531x) & (n_n5010) & (n_n4967)) + ((!x23x) & (n_n5015) & (!x531x) & (!n_n5010) & (!n_n4967)) + ((!x23x) & (n_n5015) & (!x531x) & (!n_n5010) & (n_n4967)) + ((!x23x) & (n_n5015) & (!x531x) & (n_n5010) & (!n_n4967)) + ((!x23x) & (n_n5015) & (!x531x) & (n_n5010) & (n_n4967)) + ((!x23x) & (n_n5015) & (x531x) & (!n_n5010) & (!n_n4967)) + ((!x23x) & (n_n5015) & (x531x) & (!n_n5010) & (n_n4967)) + ((!x23x) & (n_n5015) & (x531x) & (n_n5010) & (!n_n4967)) + ((!x23x) & (n_n5015) & (x531x) & (n_n5010) & (n_n4967)) + ((x23x) & (!n_n5015) & (!x531x) & (!n_n5010) & (n_n4967)) + ((x23x) & (!n_n5015) & (!x531x) & (n_n5010) & (!n_n4967)) + ((x23x) & (!n_n5015) & (!x531x) & (n_n5010) & (n_n4967)) + ((x23x) & (!n_n5015) & (x531x) & (!n_n5010) & (!n_n4967)) + ((x23x) & (!n_n5015) & (x531x) & (!n_n5010) & (n_n4967)) + ((x23x) & (!n_n5015) & (x531x) & (n_n5010) & (!n_n4967)) + ((x23x) & (!n_n5015) & (x531x) & (n_n5010) & (n_n4967)) + ((x23x) & (n_n5015) & (!x531x) & (!n_n5010) & (!n_n4967)) + ((x23x) & (n_n5015) & (!x531x) & (!n_n5010) & (n_n4967)) + ((x23x) & (n_n5015) & (!x531x) & (n_n5010) & (!n_n4967)) + ((x23x) & (n_n5015) & (!x531x) & (n_n5010) & (n_n4967)) + ((x23x) & (n_n5015) & (x531x) & (!n_n5010) & (!n_n4967)) + ((x23x) & (n_n5015) & (x531x) & (!n_n5010) & (n_n4967)) + ((x23x) & (n_n5015) & (x531x) & (n_n5010) & (!n_n4967)) + ((x23x) & (n_n5015) & (x531x) & (n_n5010) & (n_n4967)));
	assign n_n4985 = (((!i_9_) & (n_n534) & (n_n509) & (n_n195)));
	assign n_n4986 = (((i_9_) & (n_n532) & (n_n509) & (n_n195)));
	assign n_n4962 = (((i_9_) & (n_n524) & (n_n535) & (n_n195)));
	assign x14814x = (((!n_n4975) & (!n_n4983) & (!n_n4985) & (!n_n4986) & (n_n4962)) + ((!n_n4975) & (!n_n4983) & (!n_n4985) & (n_n4986) & (!n_n4962)) + ((!n_n4975) & (!n_n4983) & (!n_n4985) & (n_n4986) & (n_n4962)) + ((!n_n4975) & (!n_n4983) & (n_n4985) & (!n_n4986) & (!n_n4962)) + ((!n_n4975) & (!n_n4983) & (n_n4985) & (!n_n4986) & (n_n4962)) + ((!n_n4975) & (!n_n4983) & (n_n4985) & (n_n4986) & (!n_n4962)) + ((!n_n4975) & (!n_n4983) & (n_n4985) & (n_n4986) & (n_n4962)) + ((!n_n4975) & (n_n4983) & (!n_n4985) & (!n_n4986) & (!n_n4962)) + ((!n_n4975) & (n_n4983) & (!n_n4985) & (!n_n4986) & (n_n4962)) + ((!n_n4975) & (n_n4983) & (!n_n4985) & (n_n4986) & (!n_n4962)) + ((!n_n4975) & (n_n4983) & (!n_n4985) & (n_n4986) & (n_n4962)) + ((!n_n4975) & (n_n4983) & (n_n4985) & (!n_n4986) & (!n_n4962)) + ((!n_n4975) & (n_n4983) & (n_n4985) & (!n_n4986) & (n_n4962)) + ((!n_n4975) & (n_n4983) & (n_n4985) & (n_n4986) & (!n_n4962)) + ((!n_n4975) & (n_n4983) & (n_n4985) & (n_n4986) & (n_n4962)) + ((n_n4975) & (!n_n4983) & (!n_n4985) & (!n_n4986) & (!n_n4962)) + ((n_n4975) & (!n_n4983) & (!n_n4985) & (!n_n4986) & (n_n4962)) + ((n_n4975) & (!n_n4983) & (!n_n4985) & (n_n4986) & (!n_n4962)) + ((n_n4975) & (!n_n4983) & (!n_n4985) & (n_n4986) & (n_n4962)) + ((n_n4975) & (!n_n4983) & (n_n4985) & (!n_n4986) & (!n_n4962)) + ((n_n4975) & (!n_n4983) & (n_n4985) & (!n_n4986) & (n_n4962)) + ((n_n4975) & (!n_n4983) & (n_n4985) & (n_n4986) & (!n_n4962)) + ((n_n4975) & (!n_n4983) & (n_n4985) & (n_n4986) & (n_n4962)) + ((n_n4975) & (n_n4983) & (!n_n4985) & (!n_n4986) & (!n_n4962)) + ((n_n4975) & (n_n4983) & (!n_n4985) & (!n_n4986) & (n_n4962)) + ((n_n4975) & (n_n4983) & (!n_n4985) & (n_n4986) & (!n_n4962)) + ((n_n4975) & (n_n4983) & (!n_n4985) & (n_n4986) & (n_n4962)) + ((n_n4975) & (n_n4983) & (n_n4985) & (!n_n4986) & (!n_n4962)) + ((n_n4975) & (n_n4983) & (n_n4985) & (!n_n4986) & (n_n4962)) + ((n_n4975) & (n_n4983) & (n_n4985) & (n_n4986) & (!n_n4962)) + ((n_n4975) & (n_n4983) & (n_n4985) & (n_n4986) & (n_n4962)));
	assign n_n4828 = (((i_9_) & (n_n260) & (n_n535) & (n_n530)));
	assign n_n4844 = (((i_9_) & (n_n518) & (n_n260) & (n_n530)));
	assign n_n4899 = (((!i_9_) & (n_n524) & (n_n260) & (n_n491)));
	assign n_n4897 = (((!i_9_) & (n_n526) & (n_n260) & (n_n491)));
	assign x14820x = (((!n_n4828) & (!n_n4844) & (!n_n4899) & (n_n4897)) + ((!n_n4828) & (!n_n4844) & (n_n4899) & (!n_n4897)) + ((!n_n4828) & (!n_n4844) & (n_n4899) & (n_n4897)) + ((!n_n4828) & (n_n4844) & (!n_n4899) & (!n_n4897)) + ((!n_n4828) & (n_n4844) & (!n_n4899) & (n_n4897)) + ((!n_n4828) & (n_n4844) & (n_n4899) & (!n_n4897)) + ((!n_n4828) & (n_n4844) & (n_n4899) & (n_n4897)) + ((n_n4828) & (!n_n4844) & (!n_n4899) & (!n_n4897)) + ((n_n4828) & (!n_n4844) & (!n_n4899) & (n_n4897)) + ((n_n4828) & (!n_n4844) & (n_n4899) & (!n_n4897)) + ((n_n4828) & (!n_n4844) & (n_n4899) & (n_n4897)) + ((n_n4828) & (n_n4844) & (!n_n4899) & (!n_n4897)) + ((n_n4828) & (n_n4844) & (!n_n4899) & (n_n4897)) + ((n_n4828) & (n_n4844) & (n_n4899) & (!n_n4897)) + ((n_n4828) & (n_n4844) & (n_n4899) & (n_n4897)));
	assign n_n4886 = (((i_9_) & (n_n260) & (n_n520) & (n_n500)));
	assign n_n4871 = (((i_5_) & (i_3_) & (!i_4_) & (n_n260) & (x23x)));
	assign x14821x = (((!n_n4865) & (!n_n4847) & (!n_n4868) & (!n_n4886) & (n_n4871)) + ((!n_n4865) & (!n_n4847) & (!n_n4868) & (n_n4886) & (!n_n4871)) + ((!n_n4865) & (!n_n4847) & (!n_n4868) & (n_n4886) & (n_n4871)) + ((!n_n4865) & (!n_n4847) & (n_n4868) & (!n_n4886) & (!n_n4871)) + ((!n_n4865) & (!n_n4847) & (n_n4868) & (!n_n4886) & (n_n4871)) + ((!n_n4865) & (!n_n4847) & (n_n4868) & (n_n4886) & (!n_n4871)) + ((!n_n4865) & (!n_n4847) & (n_n4868) & (n_n4886) & (n_n4871)) + ((!n_n4865) & (n_n4847) & (!n_n4868) & (!n_n4886) & (!n_n4871)) + ((!n_n4865) & (n_n4847) & (!n_n4868) & (!n_n4886) & (n_n4871)) + ((!n_n4865) & (n_n4847) & (!n_n4868) & (n_n4886) & (!n_n4871)) + ((!n_n4865) & (n_n4847) & (!n_n4868) & (n_n4886) & (n_n4871)) + ((!n_n4865) & (n_n4847) & (n_n4868) & (!n_n4886) & (!n_n4871)) + ((!n_n4865) & (n_n4847) & (n_n4868) & (!n_n4886) & (n_n4871)) + ((!n_n4865) & (n_n4847) & (n_n4868) & (n_n4886) & (!n_n4871)) + ((!n_n4865) & (n_n4847) & (n_n4868) & (n_n4886) & (n_n4871)) + ((n_n4865) & (!n_n4847) & (!n_n4868) & (!n_n4886) & (!n_n4871)) + ((n_n4865) & (!n_n4847) & (!n_n4868) & (!n_n4886) & (n_n4871)) + ((n_n4865) & (!n_n4847) & (!n_n4868) & (n_n4886) & (!n_n4871)) + ((n_n4865) & (!n_n4847) & (!n_n4868) & (n_n4886) & (n_n4871)) + ((n_n4865) & (!n_n4847) & (n_n4868) & (!n_n4886) & (!n_n4871)) + ((n_n4865) & (!n_n4847) & (n_n4868) & (!n_n4886) & (n_n4871)) + ((n_n4865) & (!n_n4847) & (n_n4868) & (n_n4886) & (!n_n4871)) + ((n_n4865) & (!n_n4847) & (n_n4868) & (n_n4886) & (n_n4871)) + ((n_n4865) & (n_n4847) & (!n_n4868) & (!n_n4886) & (!n_n4871)) + ((n_n4865) & (n_n4847) & (!n_n4868) & (!n_n4886) & (n_n4871)) + ((n_n4865) & (n_n4847) & (!n_n4868) & (n_n4886) & (!n_n4871)) + ((n_n4865) & (n_n4847) & (!n_n4868) & (n_n4886) & (n_n4871)) + ((n_n4865) & (n_n4847) & (n_n4868) & (!n_n4886) & (!n_n4871)) + ((n_n4865) & (n_n4847) & (n_n4868) & (!n_n4886) & (n_n4871)) + ((n_n4865) & (n_n4847) & (n_n4868) & (n_n4886) & (!n_n4871)) + ((n_n4865) & (n_n4847) & (n_n4868) & (n_n4886) & (n_n4871)));
	assign n_n4929 = (((!i_9_) & (n_n526) & (n_n473) & (n_n260)));
	assign x31x = (((!i_9_) & (n_n526) & (n_n473) & (n_n260)) + ((i_9_) & (n_n526) & (n_n473) & (n_n260)));
	assign n_n4901 = (((i_1_) & (i_2_) & (!i_0_) & (n_n491) & (x20x)));
	assign n_n4904 = (((i_9_) & (n_n482) & (n_n534) & (n_n260)));
	assign x353x = (((!n_n260) & (!n_n491) & (!x20x) & (n_n4904)) + ((!n_n260) & (!n_n491) & (x20x) & (n_n4904)) + ((!n_n260) & (n_n491) & (!x20x) & (n_n4904)) + ((!n_n260) & (n_n491) & (x20x) & (n_n4904)) + ((n_n260) & (!n_n491) & (!x20x) & (n_n4904)) + ((n_n260) & (!n_n491) & (x20x) & (n_n4904)) + ((n_n260) & (n_n491) & (!x20x) & (n_n4904)) + ((n_n260) & (n_n491) & (x20x) & (!n_n4904)) + ((n_n260) & (n_n491) & (x20x) & (n_n4904)));
	assign x14803x = (((!n_n5245) & (!n_n5278) & (!n_n5287) & (n_n5261)) + ((!n_n5245) & (!n_n5278) & (n_n5287) & (!n_n5261)) + ((!n_n5245) & (!n_n5278) & (n_n5287) & (n_n5261)) + ((!n_n5245) & (n_n5278) & (!n_n5287) & (!n_n5261)) + ((!n_n5245) & (n_n5278) & (!n_n5287) & (n_n5261)) + ((!n_n5245) & (n_n5278) & (n_n5287) & (!n_n5261)) + ((!n_n5245) & (n_n5278) & (n_n5287) & (n_n5261)) + ((n_n5245) & (!n_n5278) & (!n_n5287) & (!n_n5261)) + ((n_n5245) & (!n_n5278) & (!n_n5287) & (n_n5261)) + ((n_n5245) & (!n_n5278) & (n_n5287) & (!n_n5261)) + ((n_n5245) & (!n_n5278) & (n_n5287) & (n_n5261)) + ((n_n5245) & (n_n5278) & (!n_n5287) & (!n_n5261)) + ((n_n5245) & (n_n5278) & (!n_n5287) & (n_n5261)) + ((n_n5245) & (n_n5278) & (n_n5287) & (!n_n5261)) + ((n_n5245) & (n_n5278) & (n_n5287) & (n_n5261)));
	assign x14804x = (((!n_n5284) & (!n_n5240) & (!n_n5292) & (!n_n5235) & (n_n5248)) + ((!n_n5284) & (!n_n5240) & (!n_n5292) & (n_n5235) & (!n_n5248)) + ((!n_n5284) & (!n_n5240) & (!n_n5292) & (n_n5235) & (n_n5248)) + ((!n_n5284) & (!n_n5240) & (n_n5292) & (!n_n5235) & (!n_n5248)) + ((!n_n5284) & (!n_n5240) & (n_n5292) & (!n_n5235) & (n_n5248)) + ((!n_n5284) & (!n_n5240) & (n_n5292) & (n_n5235) & (!n_n5248)) + ((!n_n5284) & (!n_n5240) & (n_n5292) & (n_n5235) & (n_n5248)) + ((!n_n5284) & (n_n5240) & (!n_n5292) & (!n_n5235) & (!n_n5248)) + ((!n_n5284) & (n_n5240) & (!n_n5292) & (!n_n5235) & (n_n5248)) + ((!n_n5284) & (n_n5240) & (!n_n5292) & (n_n5235) & (!n_n5248)) + ((!n_n5284) & (n_n5240) & (!n_n5292) & (n_n5235) & (n_n5248)) + ((!n_n5284) & (n_n5240) & (n_n5292) & (!n_n5235) & (!n_n5248)) + ((!n_n5284) & (n_n5240) & (n_n5292) & (!n_n5235) & (n_n5248)) + ((!n_n5284) & (n_n5240) & (n_n5292) & (n_n5235) & (!n_n5248)) + ((!n_n5284) & (n_n5240) & (n_n5292) & (n_n5235) & (n_n5248)) + ((n_n5284) & (!n_n5240) & (!n_n5292) & (!n_n5235) & (!n_n5248)) + ((n_n5284) & (!n_n5240) & (!n_n5292) & (!n_n5235) & (n_n5248)) + ((n_n5284) & (!n_n5240) & (!n_n5292) & (n_n5235) & (!n_n5248)) + ((n_n5284) & (!n_n5240) & (!n_n5292) & (n_n5235) & (n_n5248)) + ((n_n5284) & (!n_n5240) & (n_n5292) & (!n_n5235) & (!n_n5248)) + ((n_n5284) & (!n_n5240) & (n_n5292) & (!n_n5235) & (n_n5248)) + ((n_n5284) & (!n_n5240) & (n_n5292) & (n_n5235) & (!n_n5248)) + ((n_n5284) & (!n_n5240) & (n_n5292) & (n_n5235) & (n_n5248)) + ((n_n5284) & (n_n5240) & (!n_n5292) & (!n_n5235) & (!n_n5248)) + ((n_n5284) & (n_n5240) & (!n_n5292) & (!n_n5235) & (n_n5248)) + ((n_n5284) & (n_n5240) & (!n_n5292) & (n_n5235) & (!n_n5248)) + ((n_n5284) & (n_n5240) & (!n_n5292) & (n_n5235) & (n_n5248)) + ((n_n5284) & (n_n5240) & (n_n5292) & (!n_n5235) & (!n_n5248)) + ((n_n5284) & (n_n5240) & (n_n5292) & (!n_n5235) & (n_n5248)) + ((n_n5284) & (n_n5240) & (n_n5292) & (n_n5235) & (!n_n5248)) + ((n_n5284) & (n_n5240) & (n_n5292) & (n_n5235) & (n_n5248)));
	assign x14825x = (((!n_n4925) & (!n_n4907) & (!n_n4901) & (n_n4904)) + ((!n_n4925) & (!n_n4907) & (n_n4901) & (!n_n4904)) + ((!n_n4925) & (!n_n4907) & (n_n4901) & (n_n4904)) + ((!n_n4925) & (n_n4907) & (!n_n4901) & (!n_n4904)) + ((!n_n4925) & (n_n4907) & (!n_n4901) & (n_n4904)) + ((!n_n4925) & (n_n4907) & (n_n4901) & (!n_n4904)) + ((!n_n4925) & (n_n4907) & (n_n4901) & (n_n4904)) + ((n_n4925) & (!n_n4907) & (!n_n4901) & (!n_n4904)) + ((n_n4925) & (!n_n4907) & (!n_n4901) & (n_n4904)) + ((n_n4925) & (!n_n4907) & (n_n4901) & (!n_n4904)) + ((n_n4925) & (!n_n4907) & (n_n4901) & (n_n4904)) + ((n_n4925) & (n_n4907) & (!n_n4901) & (!n_n4904)) + ((n_n4925) & (n_n4907) & (!n_n4901) & (n_n4904)) + ((n_n4925) & (n_n4907) & (n_n4901) & (!n_n4904)) + ((n_n4925) & (n_n4907) & (n_n4901) & (n_n4904)));
	assign x14826x = (((!n_n4913) & (!n_n4922) & (!n_n4934) & (x31x)) + ((!n_n4913) & (!n_n4922) & (n_n4934) & (!x31x)) + ((!n_n4913) & (!n_n4922) & (n_n4934) & (x31x)) + ((!n_n4913) & (n_n4922) & (!n_n4934) & (!x31x)) + ((!n_n4913) & (n_n4922) & (!n_n4934) & (x31x)) + ((!n_n4913) & (n_n4922) & (n_n4934) & (!x31x)) + ((!n_n4913) & (n_n4922) & (n_n4934) & (x31x)) + ((n_n4913) & (!n_n4922) & (!n_n4934) & (!x31x)) + ((n_n4913) & (!n_n4922) & (!n_n4934) & (x31x)) + ((n_n4913) & (!n_n4922) & (n_n4934) & (!x31x)) + ((n_n4913) & (!n_n4922) & (n_n4934) & (x31x)) + ((n_n4913) & (n_n4922) & (!n_n4934) & (!x31x)) + ((n_n4913) & (n_n4922) & (!n_n4934) & (x31x)) + ((n_n4913) & (n_n4922) & (n_n4934) & (!x31x)) + ((n_n4913) & (n_n4922) & (n_n4934) & (x31x)));
	assign x14834x = (((!n_n4616) & (!n_n4608) & (!n_n4606) & (!n_n4628) & (n_n4629)) + ((!n_n4616) & (!n_n4608) & (!n_n4606) & (n_n4628) & (!n_n4629)) + ((!n_n4616) & (!n_n4608) & (!n_n4606) & (n_n4628) & (n_n4629)) + ((!n_n4616) & (!n_n4608) & (n_n4606) & (!n_n4628) & (!n_n4629)) + ((!n_n4616) & (!n_n4608) & (n_n4606) & (!n_n4628) & (n_n4629)) + ((!n_n4616) & (!n_n4608) & (n_n4606) & (n_n4628) & (!n_n4629)) + ((!n_n4616) & (!n_n4608) & (n_n4606) & (n_n4628) & (n_n4629)) + ((!n_n4616) & (n_n4608) & (!n_n4606) & (!n_n4628) & (!n_n4629)) + ((!n_n4616) & (n_n4608) & (!n_n4606) & (!n_n4628) & (n_n4629)) + ((!n_n4616) & (n_n4608) & (!n_n4606) & (n_n4628) & (!n_n4629)) + ((!n_n4616) & (n_n4608) & (!n_n4606) & (n_n4628) & (n_n4629)) + ((!n_n4616) & (n_n4608) & (n_n4606) & (!n_n4628) & (!n_n4629)) + ((!n_n4616) & (n_n4608) & (n_n4606) & (!n_n4628) & (n_n4629)) + ((!n_n4616) & (n_n4608) & (n_n4606) & (n_n4628) & (!n_n4629)) + ((!n_n4616) & (n_n4608) & (n_n4606) & (n_n4628) & (n_n4629)) + ((n_n4616) & (!n_n4608) & (!n_n4606) & (!n_n4628) & (!n_n4629)) + ((n_n4616) & (!n_n4608) & (!n_n4606) & (!n_n4628) & (n_n4629)) + ((n_n4616) & (!n_n4608) & (!n_n4606) & (n_n4628) & (!n_n4629)) + ((n_n4616) & (!n_n4608) & (!n_n4606) & (n_n4628) & (n_n4629)) + ((n_n4616) & (!n_n4608) & (n_n4606) & (!n_n4628) & (!n_n4629)) + ((n_n4616) & (!n_n4608) & (n_n4606) & (!n_n4628) & (n_n4629)) + ((n_n4616) & (!n_n4608) & (n_n4606) & (n_n4628) & (!n_n4629)) + ((n_n4616) & (!n_n4608) & (n_n4606) & (n_n4628) & (n_n4629)) + ((n_n4616) & (n_n4608) & (!n_n4606) & (!n_n4628) & (!n_n4629)) + ((n_n4616) & (n_n4608) & (!n_n4606) & (!n_n4628) & (n_n4629)) + ((n_n4616) & (n_n4608) & (!n_n4606) & (n_n4628) & (!n_n4629)) + ((n_n4616) & (n_n4608) & (!n_n4606) & (n_n4628) & (n_n4629)) + ((n_n4616) & (n_n4608) & (n_n4606) & (!n_n4628) & (!n_n4629)) + ((n_n4616) & (n_n4608) & (n_n4606) & (!n_n4628) & (n_n4629)) + ((n_n4616) & (n_n4608) & (n_n4606) & (n_n4628) & (!n_n4629)) + ((n_n4616) & (n_n4608) & (n_n4606) & (n_n4628) & (n_n4629)));
	assign x14839x = (((!n_n4463) & (!n_n4494) & (!n_n4470) & (n_n4460)) + ((!n_n4463) & (!n_n4494) & (n_n4470) & (!n_n4460)) + ((!n_n4463) & (!n_n4494) & (n_n4470) & (n_n4460)) + ((!n_n4463) & (n_n4494) & (!n_n4470) & (!n_n4460)) + ((!n_n4463) & (n_n4494) & (!n_n4470) & (n_n4460)) + ((!n_n4463) & (n_n4494) & (n_n4470) & (!n_n4460)) + ((!n_n4463) & (n_n4494) & (n_n4470) & (n_n4460)) + ((n_n4463) & (!n_n4494) & (!n_n4470) & (!n_n4460)) + ((n_n4463) & (!n_n4494) & (!n_n4470) & (n_n4460)) + ((n_n4463) & (!n_n4494) & (n_n4470) & (!n_n4460)) + ((n_n4463) & (!n_n4494) & (n_n4470) & (n_n4460)) + ((n_n4463) & (n_n4494) & (!n_n4470) & (!n_n4460)) + ((n_n4463) & (n_n4494) & (!n_n4470) & (n_n4460)) + ((n_n4463) & (n_n4494) & (n_n4470) & (!n_n4460)) + ((n_n4463) & (n_n4494) & (n_n4470) & (n_n4460)));
	assign x14840x = (((!n_n4504) & (!n_n4525) & (!n_n4457) & (!n_n4475) & (n_n4476)) + ((!n_n4504) & (!n_n4525) & (!n_n4457) & (n_n4475) & (!n_n4476)) + ((!n_n4504) & (!n_n4525) & (!n_n4457) & (n_n4475) & (n_n4476)) + ((!n_n4504) & (!n_n4525) & (n_n4457) & (!n_n4475) & (!n_n4476)) + ((!n_n4504) & (!n_n4525) & (n_n4457) & (!n_n4475) & (n_n4476)) + ((!n_n4504) & (!n_n4525) & (n_n4457) & (n_n4475) & (!n_n4476)) + ((!n_n4504) & (!n_n4525) & (n_n4457) & (n_n4475) & (n_n4476)) + ((!n_n4504) & (n_n4525) & (!n_n4457) & (!n_n4475) & (!n_n4476)) + ((!n_n4504) & (n_n4525) & (!n_n4457) & (!n_n4475) & (n_n4476)) + ((!n_n4504) & (n_n4525) & (!n_n4457) & (n_n4475) & (!n_n4476)) + ((!n_n4504) & (n_n4525) & (!n_n4457) & (n_n4475) & (n_n4476)) + ((!n_n4504) & (n_n4525) & (n_n4457) & (!n_n4475) & (!n_n4476)) + ((!n_n4504) & (n_n4525) & (n_n4457) & (!n_n4475) & (n_n4476)) + ((!n_n4504) & (n_n4525) & (n_n4457) & (n_n4475) & (!n_n4476)) + ((!n_n4504) & (n_n4525) & (n_n4457) & (n_n4475) & (n_n4476)) + ((n_n4504) & (!n_n4525) & (!n_n4457) & (!n_n4475) & (!n_n4476)) + ((n_n4504) & (!n_n4525) & (!n_n4457) & (!n_n4475) & (n_n4476)) + ((n_n4504) & (!n_n4525) & (!n_n4457) & (n_n4475) & (!n_n4476)) + ((n_n4504) & (!n_n4525) & (!n_n4457) & (n_n4475) & (n_n4476)) + ((n_n4504) & (!n_n4525) & (n_n4457) & (!n_n4475) & (!n_n4476)) + ((n_n4504) & (!n_n4525) & (n_n4457) & (!n_n4475) & (n_n4476)) + ((n_n4504) & (!n_n4525) & (n_n4457) & (n_n4475) & (!n_n4476)) + ((n_n4504) & (!n_n4525) & (n_n4457) & (n_n4475) & (n_n4476)) + ((n_n4504) & (n_n4525) & (!n_n4457) & (!n_n4475) & (!n_n4476)) + ((n_n4504) & (n_n4525) & (!n_n4457) & (!n_n4475) & (n_n4476)) + ((n_n4504) & (n_n4525) & (!n_n4457) & (n_n4475) & (!n_n4476)) + ((n_n4504) & (n_n4525) & (!n_n4457) & (n_n4475) & (n_n4476)) + ((n_n4504) & (n_n4525) & (n_n4457) & (!n_n4475) & (!n_n4476)) + ((n_n4504) & (n_n4525) & (n_n4457) & (!n_n4475) & (n_n4476)) + ((n_n4504) & (n_n4525) & (n_n4457) & (n_n4475) & (!n_n4476)) + ((n_n4504) & (n_n4525) & (n_n4457) & (n_n4475) & (n_n4476)));
	assign x14849x = (((!x118x) & (!x349x) & (!x14834x) & (!x14839x) & (x14840x)) + ((!x118x) & (!x349x) & (!x14834x) & (x14839x) & (!x14840x)) + ((!x118x) & (!x349x) & (!x14834x) & (x14839x) & (x14840x)) + ((!x118x) & (!x349x) & (x14834x) & (!x14839x) & (!x14840x)) + ((!x118x) & (!x349x) & (x14834x) & (!x14839x) & (x14840x)) + ((!x118x) & (!x349x) & (x14834x) & (x14839x) & (!x14840x)) + ((!x118x) & (!x349x) & (x14834x) & (x14839x) & (x14840x)) + ((!x118x) & (x349x) & (!x14834x) & (!x14839x) & (!x14840x)) + ((!x118x) & (x349x) & (!x14834x) & (!x14839x) & (x14840x)) + ((!x118x) & (x349x) & (!x14834x) & (x14839x) & (!x14840x)) + ((!x118x) & (x349x) & (!x14834x) & (x14839x) & (x14840x)) + ((!x118x) & (x349x) & (x14834x) & (!x14839x) & (!x14840x)) + ((!x118x) & (x349x) & (x14834x) & (!x14839x) & (x14840x)) + ((!x118x) & (x349x) & (x14834x) & (x14839x) & (!x14840x)) + ((!x118x) & (x349x) & (x14834x) & (x14839x) & (x14840x)) + ((x118x) & (!x349x) & (!x14834x) & (!x14839x) & (!x14840x)) + ((x118x) & (!x349x) & (!x14834x) & (!x14839x) & (x14840x)) + ((x118x) & (!x349x) & (!x14834x) & (x14839x) & (!x14840x)) + ((x118x) & (!x349x) & (!x14834x) & (x14839x) & (x14840x)) + ((x118x) & (!x349x) & (x14834x) & (!x14839x) & (!x14840x)) + ((x118x) & (!x349x) & (x14834x) & (!x14839x) & (x14840x)) + ((x118x) & (!x349x) & (x14834x) & (x14839x) & (!x14840x)) + ((x118x) & (!x349x) & (x14834x) & (x14839x) & (x14840x)) + ((x118x) & (x349x) & (!x14834x) & (!x14839x) & (!x14840x)) + ((x118x) & (x349x) & (!x14834x) & (!x14839x) & (x14840x)) + ((x118x) & (x349x) & (!x14834x) & (x14839x) & (!x14840x)) + ((x118x) & (x349x) & (!x14834x) & (x14839x) & (x14840x)) + ((x118x) & (x349x) & (x14834x) & (!x14839x) & (!x14840x)) + ((x118x) & (x349x) & (x14834x) & (!x14839x) & (x14840x)) + ((x118x) & (x349x) & (x14834x) & (x14839x) & (!x14840x)) + ((x118x) & (x349x) & (x14834x) & (x14839x) & (x14840x)));
	assign n_n4803 = (((!i_9_) & (n_n524) & (n_n473) & (n_n325)));
	assign n_n4770 = (((i_9_) & (n_n524) & (n_n325) & (n_n491)));
	assign n_n4771 = (((!i_9_) & (n_n524) & (n_n325) & (n_n491)));
	assign n_n4772 = (((i_9_) & (n_n325) & (n_n522) & (n_n491)));
	assign x14869x = (((!n_n4790) & (!n_n4800) & (!n_n4766) & (!n_n4826) & (n_n4805)) + ((!n_n4790) & (!n_n4800) & (!n_n4766) & (n_n4826) & (!n_n4805)) + ((!n_n4790) & (!n_n4800) & (!n_n4766) & (n_n4826) & (n_n4805)) + ((!n_n4790) & (!n_n4800) & (n_n4766) & (!n_n4826) & (!n_n4805)) + ((!n_n4790) & (!n_n4800) & (n_n4766) & (!n_n4826) & (n_n4805)) + ((!n_n4790) & (!n_n4800) & (n_n4766) & (n_n4826) & (!n_n4805)) + ((!n_n4790) & (!n_n4800) & (n_n4766) & (n_n4826) & (n_n4805)) + ((!n_n4790) & (n_n4800) & (!n_n4766) & (!n_n4826) & (!n_n4805)) + ((!n_n4790) & (n_n4800) & (!n_n4766) & (!n_n4826) & (n_n4805)) + ((!n_n4790) & (n_n4800) & (!n_n4766) & (n_n4826) & (!n_n4805)) + ((!n_n4790) & (n_n4800) & (!n_n4766) & (n_n4826) & (n_n4805)) + ((!n_n4790) & (n_n4800) & (n_n4766) & (!n_n4826) & (!n_n4805)) + ((!n_n4790) & (n_n4800) & (n_n4766) & (!n_n4826) & (n_n4805)) + ((!n_n4790) & (n_n4800) & (n_n4766) & (n_n4826) & (!n_n4805)) + ((!n_n4790) & (n_n4800) & (n_n4766) & (n_n4826) & (n_n4805)) + ((n_n4790) & (!n_n4800) & (!n_n4766) & (!n_n4826) & (!n_n4805)) + ((n_n4790) & (!n_n4800) & (!n_n4766) & (!n_n4826) & (n_n4805)) + ((n_n4790) & (!n_n4800) & (!n_n4766) & (n_n4826) & (!n_n4805)) + ((n_n4790) & (!n_n4800) & (!n_n4766) & (n_n4826) & (n_n4805)) + ((n_n4790) & (!n_n4800) & (n_n4766) & (!n_n4826) & (!n_n4805)) + ((n_n4790) & (!n_n4800) & (n_n4766) & (!n_n4826) & (n_n4805)) + ((n_n4790) & (!n_n4800) & (n_n4766) & (n_n4826) & (!n_n4805)) + ((n_n4790) & (!n_n4800) & (n_n4766) & (n_n4826) & (n_n4805)) + ((n_n4790) & (n_n4800) & (!n_n4766) & (!n_n4826) & (!n_n4805)) + ((n_n4790) & (n_n4800) & (!n_n4766) & (!n_n4826) & (n_n4805)) + ((n_n4790) & (n_n4800) & (!n_n4766) & (n_n4826) & (!n_n4805)) + ((n_n4790) & (n_n4800) & (!n_n4766) & (n_n4826) & (n_n4805)) + ((n_n4790) & (n_n4800) & (n_n4766) & (!n_n4826) & (!n_n4805)) + ((n_n4790) & (n_n4800) & (n_n4766) & (!n_n4826) & (n_n4805)) + ((n_n4790) & (n_n4800) & (n_n4766) & (n_n4826) & (!n_n4805)) + ((n_n4790) & (n_n4800) & (n_n4766) & (n_n4826) & (n_n4805)));
	assign x14870x = (((!n_n4803) & (!n_n4770) & (!n_n4771) & (!n_n4772) & (x14869x)) + ((!n_n4803) & (!n_n4770) & (!n_n4771) & (n_n4772) & (!x14869x)) + ((!n_n4803) & (!n_n4770) & (!n_n4771) & (n_n4772) & (x14869x)) + ((!n_n4803) & (!n_n4770) & (n_n4771) & (!n_n4772) & (!x14869x)) + ((!n_n4803) & (!n_n4770) & (n_n4771) & (!n_n4772) & (x14869x)) + ((!n_n4803) & (!n_n4770) & (n_n4771) & (n_n4772) & (!x14869x)) + ((!n_n4803) & (!n_n4770) & (n_n4771) & (n_n4772) & (x14869x)) + ((!n_n4803) & (n_n4770) & (!n_n4771) & (!n_n4772) & (!x14869x)) + ((!n_n4803) & (n_n4770) & (!n_n4771) & (!n_n4772) & (x14869x)) + ((!n_n4803) & (n_n4770) & (!n_n4771) & (n_n4772) & (!x14869x)) + ((!n_n4803) & (n_n4770) & (!n_n4771) & (n_n4772) & (x14869x)) + ((!n_n4803) & (n_n4770) & (n_n4771) & (!n_n4772) & (!x14869x)) + ((!n_n4803) & (n_n4770) & (n_n4771) & (!n_n4772) & (x14869x)) + ((!n_n4803) & (n_n4770) & (n_n4771) & (n_n4772) & (!x14869x)) + ((!n_n4803) & (n_n4770) & (n_n4771) & (n_n4772) & (x14869x)) + ((n_n4803) & (!n_n4770) & (!n_n4771) & (!n_n4772) & (!x14869x)) + ((n_n4803) & (!n_n4770) & (!n_n4771) & (!n_n4772) & (x14869x)) + ((n_n4803) & (!n_n4770) & (!n_n4771) & (n_n4772) & (!x14869x)) + ((n_n4803) & (!n_n4770) & (!n_n4771) & (n_n4772) & (x14869x)) + ((n_n4803) & (!n_n4770) & (n_n4771) & (!n_n4772) & (!x14869x)) + ((n_n4803) & (!n_n4770) & (n_n4771) & (!n_n4772) & (x14869x)) + ((n_n4803) & (!n_n4770) & (n_n4771) & (n_n4772) & (!x14869x)) + ((n_n4803) & (!n_n4770) & (n_n4771) & (n_n4772) & (x14869x)) + ((n_n4803) & (n_n4770) & (!n_n4771) & (!n_n4772) & (!x14869x)) + ((n_n4803) & (n_n4770) & (!n_n4771) & (!n_n4772) & (x14869x)) + ((n_n4803) & (n_n4770) & (!n_n4771) & (n_n4772) & (!x14869x)) + ((n_n4803) & (n_n4770) & (!n_n4771) & (n_n4772) & (x14869x)) + ((n_n4803) & (n_n4770) & (n_n4771) & (!n_n4772) & (!x14869x)) + ((n_n4803) & (n_n4770) & (n_n4771) & (!n_n4772) & (x14869x)) + ((n_n4803) & (n_n4770) & (n_n4771) & (n_n4772) & (!x14869x)) + ((n_n4803) & (n_n4770) & (n_n4771) & (n_n4772) & (x14869x)));
	assign x14855x = (((!n_n4656) & (!n_n4697) & (!n_n4681) & (n_n4660)) + ((!n_n4656) & (!n_n4697) & (n_n4681) & (!n_n4660)) + ((!n_n4656) & (!n_n4697) & (n_n4681) & (n_n4660)) + ((!n_n4656) & (n_n4697) & (!n_n4681) & (!n_n4660)) + ((!n_n4656) & (n_n4697) & (!n_n4681) & (n_n4660)) + ((!n_n4656) & (n_n4697) & (n_n4681) & (!n_n4660)) + ((!n_n4656) & (n_n4697) & (n_n4681) & (n_n4660)) + ((n_n4656) & (!n_n4697) & (!n_n4681) & (!n_n4660)) + ((n_n4656) & (!n_n4697) & (!n_n4681) & (n_n4660)) + ((n_n4656) & (!n_n4697) & (n_n4681) & (!n_n4660)) + ((n_n4656) & (!n_n4697) & (n_n4681) & (n_n4660)) + ((n_n4656) & (n_n4697) & (!n_n4681) & (!n_n4660)) + ((n_n4656) & (n_n4697) & (!n_n4681) & (n_n4660)) + ((n_n4656) & (n_n4697) & (n_n4681) & (!n_n4660)) + ((n_n4656) & (n_n4697) & (n_n4681) & (n_n4660)));
	assign x14856x = (((!n_n4673) & (!n_n4690) & (!n_n4665) & (!n_n4708) & (n_n4692)) + ((!n_n4673) & (!n_n4690) & (!n_n4665) & (n_n4708) & (!n_n4692)) + ((!n_n4673) & (!n_n4690) & (!n_n4665) & (n_n4708) & (n_n4692)) + ((!n_n4673) & (!n_n4690) & (n_n4665) & (!n_n4708) & (!n_n4692)) + ((!n_n4673) & (!n_n4690) & (n_n4665) & (!n_n4708) & (n_n4692)) + ((!n_n4673) & (!n_n4690) & (n_n4665) & (n_n4708) & (!n_n4692)) + ((!n_n4673) & (!n_n4690) & (n_n4665) & (n_n4708) & (n_n4692)) + ((!n_n4673) & (n_n4690) & (!n_n4665) & (!n_n4708) & (!n_n4692)) + ((!n_n4673) & (n_n4690) & (!n_n4665) & (!n_n4708) & (n_n4692)) + ((!n_n4673) & (n_n4690) & (!n_n4665) & (n_n4708) & (!n_n4692)) + ((!n_n4673) & (n_n4690) & (!n_n4665) & (n_n4708) & (n_n4692)) + ((!n_n4673) & (n_n4690) & (n_n4665) & (!n_n4708) & (!n_n4692)) + ((!n_n4673) & (n_n4690) & (n_n4665) & (!n_n4708) & (n_n4692)) + ((!n_n4673) & (n_n4690) & (n_n4665) & (n_n4708) & (!n_n4692)) + ((!n_n4673) & (n_n4690) & (n_n4665) & (n_n4708) & (n_n4692)) + ((n_n4673) & (!n_n4690) & (!n_n4665) & (!n_n4708) & (!n_n4692)) + ((n_n4673) & (!n_n4690) & (!n_n4665) & (!n_n4708) & (n_n4692)) + ((n_n4673) & (!n_n4690) & (!n_n4665) & (n_n4708) & (!n_n4692)) + ((n_n4673) & (!n_n4690) & (!n_n4665) & (n_n4708) & (n_n4692)) + ((n_n4673) & (!n_n4690) & (n_n4665) & (!n_n4708) & (!n_n4692)) + ((n_n4673) & (!n_n4690) & (n_n4665) & (!n_n4708) & (n_n4692)) + ((n_n4673) & (!n_n4690) & (n_n4665) & (n_n4708) & (!n_n4692)) + ((n_n4673) & (!n_n4690) & (n_n4665) & (n_n4708) & (n_n4692)) + ((n_n4673) & (n_n4690) & (!n_n4665) & (!n_n4708) & (!n_n4692)) + ((n_n4673) & (n_n4690) & (!n_n4665) & (!n_n4708) & (n_n4692)) + ((n_n4673) & (n_n4690) & (!n_n4665) & (n_n4708) & (!n_n4692)) + ((n_n4673) & (n_n4690) & (!n_n4665) & (n_n4708) & (n_n4692)) + ((n_n4673) & (n_n4690) & (n_n4665) & (!n_n4708) & (!n_n4692)) + ((n_n4673) & (n_n4690) & (n_n4665) & (!n_n4708) & (n_n4692)) + ((n_n4673) & (n_n4690) & (n_n4665) & (n_n4708) & (!n_n4692)) + ((n_n4673) & (n_n4690) & (n_n4665) & (n_n4708) & (n_n4692)));
	assign x14861x = (((!n_n4735) & (!n_n4724) & (!n_n4725) & (n_n4733)) + ((!n_n4735) & (!n_n4724) & (n_n4725) & (!n_n4733)) + ((!n_n4735) & (!n_n4724) & (n_n4725) & (n_n4733)) + ((!n_n4735) & (n_n4724) & (!n_n4725) & (!n_n4733)) + ((!n_n4735) & (n_n4724) & (!n_n4725) & (n_n4733)) + ((!n_n4735) & (n_n4724) & (n_n4725) & (!n_n4733)) + ((!n_n4735) & (n_n4724) & (n_n4725) & (n_n4733)) + ((n_n4735) & (!n_n4724) & (!n_n4725) & (!n_n4733)) + ((n_n4735) & (!n_n4724) & (!n_n4725) & (n_n4733)) + ((n_n4735) & (!n_n4724) & (n_n4725) & (!n_n4733)) + ((n_n4735) & (!n_n4724) & (n_n4725) & (n_n4733)) + ((n_n4735) & (n_n4724) & (!n_n4725) & (!n_n4733)) + ((n_n4735) & (n_n4724) & (!n_n4725) & (n_n4733)) + ((n_n4735) & (n_n4724) & (n_n4725) & (!n_n4733)) + ((n_n4735) & (n_n4724) & (n_n4725) & (n_n4733)));
	assign x14862x = (((!n_n4747) & (!n_n4760) & (!n_n4758) & (!n_n4745) & (n_n4714)) + ((!n_n4747) & (!n_n4760) & (!n_n4758) & (n_n4745) & (!n_n4714)) + ((!n_n4747) & (!n_n4760) & (!n_n4758) & (n_n4745) & (n_n4714)) + ((!n_n4747) & (!n_n4760) & (n_n4758) & (!n_n4745) & (!n_n4714)) + ((!n_n4747) & (!n_n4760) & (n_n4758) & (!n_n4745) & (n_n4714)) + ((!n_n4747) & (!n_n4760) & (n_n4758) & (n_n4745) & (!n_n4714)) + ((!n_n4747) & (!n_n4760) & (n_n4758) & (n_n4745) & (n_n4714)) + ((!n_n4747) & (n_n4760) & (!n_n4758) & (!n_n4745) & (!n_n4714)) + ((!n_n4747) & (n_n4760) & (!n_n4758) & (!n_n4745) & (n_n4714)) + ((!n_n4747) & (n_n4760) & (!n_n4758) & (n_n4745) & (!n_n4714)) + ((!n_n4747) & (n_n4760) & (!n_n4758) & (n_n4745) & (n_n4714)) + ((!n_n4747) & (n_n4760) & (n_n4758) & (!n_n4745) & (!n_n4714)) + ((!n_n4747) & (n_n4760) & (n_n4758) & (!n_n4745) & (n_n4714)) + ((!n_n4747) & (n_n4760) & (n_n4758) & (n_n4745) & (!n_n4714)) + ((!n_n4747) & (n_n4760) & (n_n4758) & (n_n4745) & (n_n4714)) + ((n_n4747) & (!n_n4760) & (!n_n4758) & (!n_n4745) & (!n_n4714)) + ((n_n4747) & (!n_n4760) & (!n_n4758) & (!n_n4745) & (n_n4714)) + ((n_n4747) & (!n_n4760) & (!n_n4758) & (n_n4745) & (!n_n4714)) + ((n_n4747) & (!n_n4760) & (!n_n4758) & (n_n4745) & (n_n4714)) + ((n_n4747) & (!n_n4760) & (n_n4758) & (!n_n4745) & (!n_n4714)) + ((n_n4747) & (!n_n4760) & (n_n4758) & (!n_n4745) & (n_n4714)) + ((n_n4747) & (!n_n4760) & (n_n4758) & (n_n4745) & (!n_n4714)) + ((n_n4747) & (!n_n4760) & (n_n4758) & (n_n4745) & (n_n4714)) + ((n_n4747) & (n_n4760) & (!n_n4758) & (!n_n4745) & (!n_n4714)) + ((n_n4747) & (n_n4760) & (!n_n4758) & (!n_n4745) & (n_n4714)) + ((n_n4747) & (n_n4760) & (!n_n4758) & (n_n4745) & (!n_n4714)) + ((n_n4747) & (n_n4760) & (!n_n4758) & (n_n4745) & (n_n4714)) + ((n_n4747) & (n_n4760) & (n_n4758) & (!n_n4745) & (!n_n4714)) + ((n_n4747) & (n_n4760) & (n_n4758) & (!n_n4745) & (n_n4714)) + ((n_n4747) & (n_n4760) & (n_n4758) & (n_n4745) & (!n_n4714)) + ((n_n4747) & (n_n4760) & (n_n4758) & (n_n4745) & (n_n4714)));
	assign x14871x = (((!x14855x) & (!x14856x) & (!x14861x) & (x14862x)) + ((!x14855x) & (!x14856x) & (x14861x) & (!x14862x)) + ((!x14855x) & (!x14856x) & (x14861x) & (x14862x)) + ((!x14855x) & (x14856x) & (!x14861x) & (!x14862x)) + ((!x14855x) & (x14856x) & (!x14861x) & (x14862x)) + ((!x14855x) & (x14856x) & (x14861x) & (!x14862x)) + ((!x14855x) & (x14856x) & (x14861x) & (x14862x)) + ((x14855x) & (!x14856x) & (!x14861x) & (!x14862x)) + ((x14855x) & (!x14856x) & (!x14861x) & (x14862x)) + ((x14855x) & (!x14856x) & (x14861x) & (!x14862x)) + ((x14855x) & (!x14856x) & (x14861x) & (x14862x)) + ((x14855x) & (x14856x) & (!x14861x) & (!x14862x)) + ((x14855x) & (x14856x) & (!x14861x) & (x14862x)) + ((x14855x) & (x14856x) & (x14861x) & (!x14862x)) + ((x14855x) & (x14856x) & (x14861x) & (x14862x)));
	assign n_n4373 = (((i_1_) & (i_2_) & (i_0_) & (x20x) & (n_n500)));
	assign x14876x = (((!n_n4403) & (!n_n4382) & (!n_n4373) & (n_n4371)) + ((!n_n4403) & (!n_n4382) & (n_n4373) & (!n_n4371)) + ((!n_n4403) & (!n_n4382) & (n_n4373) & (n_n4371)) + ((!n_n4403) & (n_n4382) & (!n_n4373) & (!n_n4371)) + ((!n_n4403) & (n_n4382) & (!n_n4373) & (n_n4371)) + ((!n_n4403) & (n_n4382) & (n_n4373) & (!n_n4371)) + ((!n_n4403) & (n_n4382) & (n_n4373) & (n_n4371)) + ((n_n4403) & (!n_n4382) & (!n_n4373) & (!n_n4371)) + ((n_n4403) & (!n_n4382) & (!n_n4373) & (n_n4371)) + ((n_n4403) & (!n_n4382) & (n_n4373) & (!n_n4371)) + ((n_n4403) & (!n_n4382) & (n_n4373) & (n_n4371)) + ((n_n4403) & (n_n4382) & (!n_n4373) & (!n_n4371)) + ((n_n4403) & (n_n4382) & (!n_n4373) & (n_n4371)) + ((n_n4403) & (n_n4382) & (n_n4373) & (!n_n4371)) + ((n_n4403) & (n_n4382) & (n_n4373) & (n_n4371)));
	assign n_n4396 = (((i_9_) & (n_n536) & (n_n482) & (n_n530)));
	assign n_n4375 = (((i_1_) & (i_2_) & (i_0_) & (x23x) & (n_n500)));
	assign x14877x = (((!n_n4391) & (!n_n4362) & (!n_n4396) & (!n_n4399) & (n_n4375)) + ((!n_n4391) & (!n_n4362) & (!n_n4396) & (n_n4399) & (!n_n4375)) + ((!n_n4391) & (!n_n4362) & (!n_n4396) & (n_n4399) & (n_n4375)) + ((!n_n4391) & (!n_n4362) & (n_n4396) & (!n_n4399) & (!n_n4375)) + ((!n_n4391) & (!n_n4362) & (n_n4396) & (!n_n4399) & (n_n4375)) + ((!n_n4391) & (!n_n4362) & (n_n4396) & (n_n4399) & (!n_n4375)) + ((!n_n4391) & (!n_n4362) & (n_n4396) & (n_n4399) & (n_n4375)) + ((!n_n4391) & (n_n4362) & (!n_n4396) & (!n_n4399) & (!n_n4375)) + ((!n_n4391) & (n_n4362) & (!n_n4396) & (!n_n4399) & (n_n4375)) + ((!n_n4391) & (n_n4362) & (!n_n4396) & (n_n4399) & (!n_n4375)) + ((!n_n4391) & (n_n4362) & (!n_n4396) & (n_n4399) & (n_n4375)) + ((!n_n4391) & (n_n4362) & (n_n4396) & (!n_n4399) & (!n_n4375)) + ((!n_n4391) & (n_n4362) & (n_n4396) & (!n_n4399) & (n_n4375)) + ((!n_n4391) & (n_n4362) & (n_n4396) & (n_n4399) & (!n_n4375)) + ((!n_n4391) & (n_n4362) & (n_n4396) & (n_n4399) & (n_n4375)) + ((n_n4391) & (!n_n4362) & (!n_n4396) & (!n_n4399) & (!n_n4375)) + ((n_n4391) & (!n_n4362) & (!n_n4396) & (!n_n4399) & (n_n4375)) + ((n_n4391) & (!n_n4362) & (!n_n4396) & (n_n4399) & (!n_n4375)) + ((n_n4391) & (!n_n4362) & (!n_n4396) & (n_n4399) & (n_n4375)) + ((n_n4391) & (!n_n4362) & (n_n4396) & (!n_n4399) & (!n_n4375)) + ((n_n4391) & (!n_n4362) & (n_n4396) & (!n_n4399) & (n_n4375)) + ((n_n4391) & (!n_n4362) & (n_n4396) & (n_n4399) & (!n_n4375)) + ((n_n4391) & (!n_n4362) & (n_n4396) & (n_n4399) & (n_n4375)) + ((n_n4391) & (n_n4362) & (!n_n4396) & (!n_n4399) & (!n_n4375)) + ((n_n4391) & (n_n4362) & (!n_n4396) & (!n_n4399) & (n_n4375)) + ((n_n4391) & (n_n4362) & (!n_n4396) & (n_n4399) & (!n_n4375)) + ((n_n4391) & (n_n4362) & (!n_n4396) & (n_n4399) & (n_n4375)) + ((n_n4391) & (n_n4362) & (n_n4396) & (!n_n4399) & (!n_n4375)) + ((n_n4391) & (n_n4362) & (n_n4396) & (!n_n4399) & (n_n4375)) + ((n_n4391) & (n_n4362) & (n_n4396) & (n_n4399) & (!n_n4375)) + ((n_n4391) & (n_n4362) & (n_n4396) & (n_n4399) & (n_n4375)));
	assign n_n4344 = (((i_9_) & (n_n536) & (n_n534) & (n_n509)));
	assign x14882x = (((!n_n4318) & (!n_n4344) & (!n_n4320) & (n_n4341)) + ((!n_n4318) & (!n_n4344) & (n_n4320) & (!n_n4341)) + ((!n_n4318) & (!n_n4344) & (n_n4320) & (n_n4341)) + ((!n_n4318) & (n_n4344) & (!n_n4320) & (!n_n4341)) + ((!n_n4318) & (n_n4344) & (!n_n4320) & (n_n4341)) + ((!n_n4318) & (n_n4344) & (n_n4320) & (!n_n4341)) + ((!n_n4318) & (n_n4344) & (n_n4320) & (n_n4341)) + ((n_n4318) & (!n_n4344) & (!n_n4320) & (!n_n4341)) + ((n_n4318) & (!n_n4344) & (!n_n4320) & (n_n4341)) + ((n_n4318) & (!n_n4344) & (n_n4320) & (!n_n4341)) + ((n_n4318) & (!n_n4344) & (n_n4320) & (n_n4341)) + ((n_n4318) & (n_n4344) & (!n_n4320) & (!n_n4341)) + ((n_n4318) & (n_n4344) & (!n_n4320) & (n_n4341)) + ((n_n4318) & (n_n4344) & (n_n4320) & (!n_n4341)) + ((n_n4318) & (n_n4344) & (n_n4320) & (n_n4341)));
	assign n_n4330 = (((i_9_) & (n_n536) & (n_n518) & (n_n532)));
	assign n_n4352 = (((i_9_) & (n_n536) & (n_n526) & (n_n509)));
	assign n_n4351 = (((!i_9_) & (n_n536) & (n_n528) & (n_n509)));
	assign n_n4313 = (((!i_9_) & (n_n536) & (n_n534) & (n_n535)));
	assign x14883x = (((!n_n4330) & (!n_n4352) & (!n_n4351) & (!n_n4316) & (n_n4313)) + ((!n_n4330) & (!n_n4352) & (!n_n4351) & (n_n4316) & (!n_n4313)) + ((!n_n4330) & (!n_n4352) & (!n_n4351) & (n_n4316) & (n_n4313)) + ((!n_n4330) & (!n_n4352) & (n_n4351) & (!n_n4316) & (!n_n4313)) + ((!n_n4330) & (!n_n4352) & (n_n4351) & (!n_n4316) & (n_n4313)) + ((!n_n4330) & (!n_n4352) & (n_n4351) & (n_n4316) & (!n_n4313)) + ((!n_n4330) & (!n_n4352) & (n_n4351) & (n_n4316) & (n_n4313)) + ((!n_n4330) & (n_n4352) & (!n_n4351) & (!n_n4316) & (!n_n4313)) + ((!n_n4330) & (n_n4352) & (!n_n4351) & (!n_n4316) & (n_n4313)) + ((!n_n4330) & (n_n4352) & (!n_n4351) & (n_n4316) & (!n_n4313)) + ((!n_n4330) & (n_n4352) & (!n_n4351) & (n_n4316) & (n_n4313)) + ((!n_n4330) & (n_n4352) & (n_n4351) & (!n_n4316) & (!n_n4313)) + ((!n_n4330) & (n_n4352) & (n_n4351) & (!n_n4316) & (n_n4313)) + ((!n_n4330) & (n_n4352) & (n_n4351) & (n_n4316) & (!n_n4313)) + ((!n_n4330) & (n_n4352) & (n_n4351) & (n_n4316) & (n_n4313)) + ((n_n4330) & (!n_n4352) & (!n_n4351) & (!n_n4316) & (!n_n4313)) + ((n_n4330) & (!n_n4352) & (!n_n4351) & (!n_n4316) & (n_n4313)) + ((n_n4330) & (!n_n4352) & (!n_n4351) & (n_n4316) & (!n_n4313)) + ((n_n4330) & (!n_n4352) & (!n_n4351) & (n_n4316) & (n_n4313)) + ((n_n4330) & (!n_n4352) & (n_n4351) & (!n_n4316) & (!n_n4313)) + ((n_n4330) & (!n_n4352) & (n_n4351) & (!n_n4316) & (n_n4313)) + ((n_n4330) & (!n_n4352) & (n_n4351) & (n_n4316) & (!n_n4313)) + ((n_n4330) & (!n_n4352) & (n_n4351) & (n_n4316) & (n_n4313)) + ((n_n4330) & (n_n4352) & (!n_n4351) & (!n_n4316) & (!n_n4313)) + ((n_n4330) & (n_n4352) & (!n_n4351) & (!n_n4316) & (n_n4313)) + ((n_n4330) & (n_n4352) & (!n_n4351) & (n_n4316) & (!n_n4313)) + ((n_n4330) & (n_n4352) & (!n_n4351) & (n_n4316) & (n_n4313)) + ((n_n4330) & (n_n4352) & (n_n4351) & (!n_n4316) & (!n_n4313)) + ((n_n4330) & (n_n4352) & (n_n4351) & (!n_n4316) & (n_n4313)) + ((n_n4330) & (n_n4352) & (n_n4351) & (n_n4316) & (!n_n4313)) + ((n_n4330) & (n_n4352) & (n_n4351) & (n_n4316) & (n_n4313)));
	assign n_n4444 = (((i_9_) & (n_n455) & (n_n535) & (n_n530)));
	assign x234x = (((!i_7_) & (i_8_) & (i_6_) & (x13x) & (n_n535)) + ((i_7_) & (i_8_) & (i_6_) & (x13x) & (n_n535)));
	assign n_n4448 = (((i_9_) & (n_n526) & (n_n455) & (n_n535)));
	assign n_n4447 = (((!i_9_) & (n_n455) & (n_n528) & (n_n535)));
	assign x323x = (((!i_9_) & (!n_n526) & (n_n455) & (n_n528) & (n_n535)) + ((!i_9_) & (n_n526) & (n_n455) & (n_n528) & (n_n535)) + ((i_9_) & (n_n526) & (n_n455) & (!n_n528) & (n_n535)) + ((i_9_) & (n_n526) & (n_n455) & (n_n528) & (n_n535)));
	assign n_n4415 = (((!i_9_) & (n_n536) & (n_n528) & (n_n473)));
	assign n_n4372 = (((i_9_) & (n_n536) & (n_n522) & (n_n500)));
	assign n_n4430 = (((i_9_) & (n_n536) & (n_n528) & (n_n464)));
	assign n_n4494 = (((i_9_) & (n_n455) & (n_n528) & (n_n500)));
	assign n_n4495 = (((!i_9_) & (n_n455) & (n_n528) & (n_n500)));
	assign n_n4491 = (((!i_9_) & (n_n455) & (n_n532) & (n_n500)));
	assign n_n4834 = (((i_9_) & (n_n524) & (n_n260) & (n_n535)));
	assign n_n4835 = (((!i_9_) & (n_n524) & (n_n260) & (n_n535)));
	assign n_n4832 = (((i_9_) & (n_n526) & (n_n260) & (n_n535)));
	assign n_n4909 = (((!i_9_) & (n_n482) & (n_n260) & (n_n530)));
	assign n_n4911 = (((!i_9_) & (n_n482) & (n_n528) & (n_n260)));
	assign n_n4903 = (((i_1_) & (i_2_) & (!i_0_) & (n_n491) & (x23x)));
	assign n_n5049 = (((!i_9_) & (n_n473) & (n_n534) & (n_n195)));
	assign n_n5239 = (((!i_5_) & (i_3_) & (i_4_) & (x23x) & (n_n65)));
	assign n_n5240 = (((i_7_) & (i_8_) & (i_6_) & (x19x) & (n_n509)));
	assign n_n5238 = (((!i_5_) & (i_3_) & (i_4_) & (x19x) & (n_n520)));
	assign x130x = (((!i_9_) & (n_n524) & (n_n455) & (!n_n522) & (n_n491)) + ((!i_9_) & (n_n524) & (n_n455) & (n_n522) & (n_n491)) + ((i_9_) & (!n_n524) & (n_n455) & (n_n522) & (n_n491)) + ((i_9_) & (n_n524) & (n_n455) & (n_n522) & (n_n491)));
	assign n_n4247 = (((!i_9_) & (n_n524) & (n_n455) & (!n_n522) & (n_n491)) + ((!i_9_) & (n_n524) & (n_n455) & (n_n522) & (n_n491)) + ((i_9_) & (!n_n524) & (n_n455) & (n_n522) & (n_n491)) + ((i_9_) & (n_n524) & (n_n455) & (!n_n522) & (n_n491)) + ((i_9_) & (n_n524) & (n_n455) & (n_n522) & (n_n491)));
	assign n_n4646 = (((i_9_) & (n_n390) & (n_n491) & (n_n520)));
	assign n_n4644 = (((i_9_) & (n_n390) & (n_n522) & (n_n491)));
	assign n_n4651 = (((!i_9_) & (n_n482) & (n_n390) & (n_n532)));
	assign n_n4649 = (((!i_9_) & (n_n482) & (n_n390) & (n_n534)));
	assign n_n4652 = (((i_9_) & (n_n482) & (n_n390) & (n_n530)));
	assign x311x = (((!i_9_) & (n_n482) & (n_n390) & (n_n530)) + ((i_9_) & (n_n482) & (n_n390) & (n_n530)));
	assign x16628x = (((!n_n4643) & (!n_n4645) & (!n_n4644) & (!n_n4651) & (n_n4649)) + ((!n_n4643) & (!n_n4645) & (!n_n4644) & (n_n4651) & (!n_n4649)) + ((!n_n4643) & (!n_n4645) & (!n_n4644) & (n_n4651) & (n_n4649)) + ((!n_n4643) & (!n_n4645) & (n_n4644) & (!n_n4651) & (!n_n4649)) + ((!n_n4643) & (!n_n4645) & (n_n4644) & (!n_n4651) & (n_n4649)) + ((!n_n4643) & (!n_n4645) & (n_n4644) & (n_n4651) & (!n_n4649)) + ((!n_n4643) & (!n_n4645) & (n_n4644) & (n_n4651) & (n_n4649)) + ((!n_n4643) & (n_n4645) & (!n_n4644) & (!n_n4651) & (!n_n4649)) + ((!n_n4643) & (n_n4645) & (!n_n4644) & (!n_n4651) & (n_n4649)) + ((!n_n4643) & (n_n4645) & (!n_n4644) & (n_n4651) & (!n_n4649)) + ((!n_n4643) & (n_n4645) & (!n_n4644) & (n_n4651) & (n_n4649)) + ((!n_n4643) & (n_n4645) & (n_n4644) & (!n_n4651) & (!n_n4649)) + ((!n_n4643) & (n_n4645) & (n_n4644) & (!n_n4651) & (n_n4649)) + ((!n_n4643) & (n_n4645) & (n_n4644) & (n_n4651) & (!n_n4649)) + ((!n_n4643) & (n_n4645) & (n_n4644) & (n_n4651) & (n_n4649)) + ((n_n4643) & (!n_n4645) & (!n_n4644) & (!n_n4651) & (!n_n4649)) + ((n_n4643) & (!n_n4645) & (!n_n4644) & (!n_n4651) & (n_n4649)) + ((n_n4643) & (!n_n4645) & (!n_n4644) & (n_n4651) & (!n_n4649)) + ((n_n4643) & (!n_n4645) & (!n_n4644) & (n_n4651) & (n_n4649)) + ((n_n4643) & (!n_n4645) & (n_n4644) & (!n_n4651) & (!n_n4649)) + ((n_n4643) & (!n_n4645) & (n_n4644) & (!n_n4651) & (n_n4649)) + ((n_n4643) & (!n_n4645) & (n_n4644) & (n_n4651) & (!n_n4649)) + ((n_n4643) & (!n_n4645) & (n_n4644) & (n_n4651) & (n_n4649)) + ((n_n4643) & (n_n4645) & (!n_n4644) & (!n_n4651) & (!n_n4649)) + ((n_n4643) & (n_n4645) & (!n_n4644) & (!n_n4651) & (n_n4649)) + ((n_n4643) & (n_n4645) & (!n_n4644) & (n_n4651) & (!n_n4649)) + ((n_n4643) & (n_n4645) & (!n_n4644) & (n_n4651) & (n_n4649)) + ((n_n4643) & (n_n4645) & (n_n4644) & (!n_n4651) & (!n_n4649)) + ((n_n4643) & (n_n4645) & (n_n4644) & (!n_n4651) & (n_n4649)) + ((n_n4643) & (n_n4645) & (n_n4644) & (n_n4651) & (!n_n4649)) + ((n_n4643) & (n_n4645) & (n_n4644) & (n_n4651) & (n_n4649)));
	assign n_n4952 = (((i_9_) & (n_n534) & (n_n535) & (n_n195)));
	assign n_n4950 = (((i_9_) & (n_n260) & (n_n520) & (n_n464)));
	assign n_n3803 = (((!n_n260) & (!x23x) & (!n_n464) & (!n_n4952) & (n_n4950)) + ((!n_n260) & (!x23x) & (!n_n464) & (n_n4952) & (!n_n4950)) + ((!n_n260) & (!x23x) & (!n_n464) & (n_n4952) & (n_n4950)) + ((!n_n260) & (!x23x) & (n_n464) & (!n_n4952) & (n_n4950)) + ((!n_n260) & (!x23x) & (n_n464) & (n_n4952) & (!n_n4950)) + ((!n_n260) & (!x23x) & (n_n464) & (n_n4952) & (n_n4950)) + ((!n_n260) & (x23x) & (!n_n464) & (!n_n4952) & (n_n4950)) + ((!n_n260) & (x23x) & (!n_n464) & (n_n4952) & (!n_n4950)) + ((!n_n260) & (x23x) & (!n_n464) & (n_n4952) & (n_n4950)) + ((!n_n260) & (x23x) & (n_n464) & (!n_n4952) & (n_n4950)) + ((!n_n260) & (x23x) & (n_n464) & (n_n4952) & (!n_n4950)) + ((!n_n260) & (x23x) & (n_n464) & (n_n4952) & (n_n4950)) + ((n_n260) & (!x23x) & (!n_n464) & (!n_n4952) & (n_n4950)) + ((n_n260) & (!x23x) & (!n_n464) & (n_n4952) & (!n_n4950)) + ((n_n260) & (!x23x) & (!n_n464) & (n_n4952) & (n_n4950)) + ((n_n260) & (!x23x) & (n_n464) & (!n_n4952) & (n_n4950)) + ((n_n260) & (!x23x) & (n_n464) & (n_n4952) & (!n_n4950)) + ((n_n260) & (!x23x) & (n_n464) & (n_n4952) & (n_n4950)) + ((n_n260) & (x23x) & (!n_n464) & (!n_n4952) & (n_n4950)) + ((n_n260) & (x23x) & (!n_n464) & (n_n4952) & (!n_n4950)) + ((n_n260) & (x23x) & (!n_n464) & (n_n4952) & (n_n4950)) + ((n_n260) & (x23x) & (n_n464) & (!n_n4952) & (!n_n4950)) + ((n_n260) & (x23x) & (n_n464) & (!n_n4952) & (n_n4950)) + ((n_n260) & (x23x) & (n_n464) & (n_n4952) & (!n_n4950)) + ((n_n260) & (x23x) & (n_n464) & (n_n4952) & (n_n4950)));
	assign n_n4942 = (((i_9_) & (n_n528) & (n_n260) & (n_n464)));
	assign n_n3805 = (((!i_9_) & (!n_n528) & (n_n260) & (n_n530) & (n_n464)) + ((!i_9_) & (n_n528) & (n_n260) & (!n_n530) & (n_n464)) + ((!i_9_) & (n_n528) & (n_n260) & (n_n530) & (n_n464)) + ((i_9_) & (n_n528) & (n_n260) & (!n_n530) & (n_n464)) + ((i_9_) & (n_n528) & (n_n260) & (n_n530) & (n_n464)));
	assign n_n4945 = (((!i_9_) & (n_n526) & (n_n260) & (n_n464)));
	assign n_n4946 = (((i_9_) & (n_n524) & (n_n260) & (n_n464)));
	assign n_n4949 = (((i_1_) & (i_2_) & (!i_0_) & (x20x) & (n_n464)));
	assign x16327x = (((!i_9_) & (!n_n260) & (!x516x) & (!n_n4945) & (n_n4949)) + ((!i_9_) & (!n_n260) & (!x516x) & (n_n4945) & (!n_n4949)) + ((!i_9_) & (!n_n260) & (!x516x) & (n_n4945) & (n_n4949)) + ((!i_9_) & (!n_n260) & (x516x) & (!n_n4945) & (n_n4949)) + ((!i_9_) & (!n_n260) & (x516x) & (n_n4945) & (!n_n4949)) + ((!i_9_) & (!n_n260) & (x516x) & (n_n4945) & (n_n4949)) + ((!i_9_) & (n_n260) & (!x516x) & (!n_n4945) & (n_n4949)) + ((!i_9_) & (n_n260) & (!x516x) & (n_n4945) & (!n_n4949)) + ((!i_9_) & (n_n260) & (!x516x) & (n_n4945) & (n_n4949)) + ((!i_9_) & (n_n260) & (x516x) & (!n_n4945) & (n_n4949)) + ((!i_9_) & (n_n260) & (x516x) & (n_n4945) & (!n_n4949)) + ((!i_9_) & (n_n260) & (x516x) & (n_n4945) & (n_n4949)) + ((i_9_) & (!n_n260) & (!x516x) & (!n_n4945) & (n_n4949)) + ((i_9_) & (!n_n260) & (!x516x) & (n_n4945) & (!n_n4949)) + ((i_9_) & (!n_n260) & (!x516x) & (n_n4945) & (n_n4949)) + ((i_9_) & (!n_n260) & (x516x) & (!n_n4945) & (n_n4949)) + ((i_9_) & (!n_n260) & (x516x) & (n_n4945) & (!n_n4949)) + ((i_9_) & (!n_n260) & (x516x) & (n_n4945) & (n_n4949)) + ((i_9_) & (n_n260) & (!x516x) & (!n_n4945) & (n_n4949)) + ((i_9_) & (n_n260) & (!x516x) & (n_n4945) & (!n_n4949)) + ((i_9_) & (n_n260) & (!x516x) & (n_n4945) & (n_n4949)) + ((i_9_) & (n_n260) & (x516x) & (!n_n4945) & (!n_n4949)) + ((i_9_) & (n_n260) & (x516x) & (!n_n4945) & (n_n4949)) + ((i_9_) & (n_n260) & (x516x) & (n_n4945) & (!n_n4949)) + ((i_9_) & (n_n260) & (x516x) & (n_n4945) & (n_n4949)));
	assign n_n5244 = (((i_5_) & (i_3_) & (!i_4_) & (x19x) & (n_n530)));
	assign n_n5245 = (((!i_9_) & (n_n509) & (n_n530) & (n_n65)));
	assign n_n5241 = (((!i_9_) & (n_n534) & (n_n509) & (n_n65)));
	assign n_n5242 = (((i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n509)));
	assign n_n5247 = (((!i_9_) & (n_n528) & (n_n509) & (n_n65)));
	assign n_n5246 = (((!i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n509)));
	assign x319x = (((!n_n518) & (!x23x) & (!n_n65) & (n_n5240)) + ((!n_n518) & (!x23x) & (n_n65) & (n_n5240)) + ((!n_n518) & (x23x) & (!n_n65) & (n_n5240)) + ((!n_n518) & (x23x) & (n_n65) & (n_n5240)) + ((n_n518) & (!x23x) & (!n_n65) & (n_n5240)) + ((n_n518) & (!x23x) & (n_n65) & (n_n5240)) + ((n_n518) & (x23x) & (!n_n65) & (n_n5240)) + ((n_n518) & (x23x) & (n_n65) & (!n_n5240)) + ((n_n518) & (x23x) & (n_n65) & (n_n5240)));
	assign x16687x = (((!n_n5238) & (!n_n5244) & (!n_n5245) & (!n_n5241) & (n_n5242)) + ((!n_n5238) & (!n_n5244) & (!n_n5245) & (n_n5241) & (!n_n5242)) + ((!n_n5238) & (!n_n5244) & (!n_n5245) & (n_n5241) & (n_n5242)) + ((!n_n5238) & (!n_n5244) & (n_n5245) & (!n_n5241) & (!n_n5242)) + ((!n_n5238) & (!n_n5244) & (n_n5245) & (!n_n5241) & (n_n5242)) + ((!n_n5238) & (!n_n5244) & (n_n5245) & (n_n5241) & (!n_n5242)) + ((!n_n5238) & (!n_n5244) & (n_n5245) & (n_n5241) & (n_n5242)) + ((!n_n5238) & (n_n5244) & (!n_n5245) & (!n_n5241) & (!n_n5242)) + ((!n_n5238) & (n_n5244) & (!n_n5245) & (!n_n5241) & (n_n5242)) + ((!n_n5238) & (n_n5244) & (!n_n5245) & (n_n5241) & (!n_n5242)) + ((!n_n5238) & (n_n5244) & (!n_n5245) & (n_n5241) & (n_n5242)) + ((!n_n5238) & (n_n5244) & (n_n5245) & (!n_n5241) & (!n_n5242)) + ((!n_n5238) & (n_n5244) & (n_n5245) & (!n_n5241) & (n_n5242)) + ((!n_n5238) & (n_n5244) & (n_n5245) & (n_n5241) & (!n_n5242)) + ((!n_n5238) & (n_n5244) & (n_n5245) & (n_n5241) & (n_n5242)) + ((n_n5238) & (!n_n5244) & (!n_n5245) & (!n_n5241) & (!n_n5242)) + ((n_n5238) & (!n_n5244) & (!n_n5245) & (!n_n5241) & (n_n5242)) + ((n_n5238) & (!n_n5244) & (!n_n5245) & (n_n5241) & (!n_n5242)) + ((n_n5238) & (!n_n5244) & (!n_n5245) & (n_n5241) & (n_n5242)) + ((n_n5238) & (!n_n5244) & (n_n5245) & (!n_n5241) & (!n_n5242)) + ((n_n5238) & (!n_n5244) & (n_n5245) & (!n_n5241) & (n_n5242)) + ((n_n5238) & (!n_n5244) & (n_n5245) & (n_n5241) & (!n_n5242)) + ((n_n5238) & (!n_n5244) & (n_n5245) & (n_n5241) & (n_n5242)) + ((n_n5238) & (n_n5244) & (!n_n5245) & (!n_n5241) & (!n_n5242)) + ((n_n5238) & (n_n5244) & (!n_n5245) & (!n_n5241) & (n_n5242)) + ((n_n5238) & (n_n5244) & (!n_n5245) & (n_n5241) & (!n_n5242)) + ((n_n5238) & (n_n5244) & (!n_n5245) & (n_n5241) & (n_n5242)) + ((n_n5238) & (n_n5244) & (n_n5245) & (!n_n5241) & (!n_n5242)) + ((n_n5238) & (n_n5244) & (n_n5245) & (!n_n5241) & (n_n5242)) + ((n_n5238) & (n_n5244) & (n_n5245) & (n_n5241) & (!n_n5242)) + ((n_n5238) & (n_n5244) & (n_n5245) & (n_n5241) & (n_n5242)));
	assign n_n4445 = (((!i_9_) & (n_n455) & (n_n535) & (n_n530)));
	assign n_n4449 = (((!i_9_) & (n_n526) & (n_n455) & (n_n535)));
	assign x368x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n455) & (n_n535)) + ((!i_9_) & (n_n524) & (!n_n526) & (n_n455) & (n_n535)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n455) & (n_n535)));
	assign x16563x = (((!n_n4444) & (!n_n4448) & (!n_n4447) & (!n_n4442) & (n_n4441)) + ((!n_n4444) & (!n_n4448) & (!n_n4447) & (n_n4442) & (!n_n4441)) + ((!n_n4444) & (!n_n4448) & (!n_n4447) & (n_n4442) & (n_n4441)) + ((!n_n4444) & (!n_n4448) & (n_n4447) & (!n_n4442) & (!n_n4441)) + ((!n_n4444) & (!n_n4448) & (n_n4447) & (!n_n4442) & (n_n4441)) + ((!n_n4444) & (!n_n4448) & (n_n4447) & (n_n4442) & (!n_n4441)) + ((!n_n4444) & (!n_n4448) & (n_n4447) & (n_n4442) & (n_n4441)) + ((!n_n4444) & (n_n4448) & (!n_n4447) & (!n_n4442) & (!n_n4441)) + ((!n_n4444) & (n_n4448) & (!n_n4447) & (!n_n4442) & (n_n4441)) + ((!n_n4444) & (n_n4448) & (!n_n4447) & (n_n4442) & (!n_n4441)) + ((!n_n4444) & (n_n4448) & (!n_n4447) & (n_n4442) & (n_n4441)) + ((!n_n4444) & (n_n4448) & (n_n4447) & (!n_n4442) & (!n_n4441)) + ((!n_n4444) & (n_n4448) & (n_n4447) & (!n_n4442) & (n_n4441)) + ((!n_n4444) & (n_n4448) & (n_n4447) & (n_n4442) & (!n_n4441)) + ((!n_n4444) & (n_n4448) & (n_n4447) & (n_n4442) & (n_n4441)) + ((n_n4444) & (!n_n4448) & (!n_n4447) & (!n_n4442) & (!n_n4441)) + ((n_n4444) & (!n_n4448) & (!n_n4447) & (!n_n4442) & (n_n4441)) + ((n_n4444) & (!n_n4448) & (!n_n4447) & (n_n4442) & (!n_n4441)) + ((n_n4444) & (!n_n4448) & (!n_n4447) & (n_n4442) & (n_n4441)) + ((n_n4444) & (!n_n4448) & (n_n4447) & (!n_n4442) & (!n_n4441)) + ((n_n4444) & (!n_n4448) & (n_n4447) & (!n_n4442) & (n_n4441)) + ((n_n4444) & (!n_n4448) & (n_n4447) & (n_n4442) & (!n_n4441)) + ((n_n4444) & (!n_n4448) & (n_n4447) & (n_n4442) & (n_n4441)) + ((n_n4444) & (n_n4448) & (!n_n4447) & (!n_n4442) & (!n_n4441)) + ((n_n4444) & (n_n4448) & (!n_n4447) & (!n_n4442) & (n_n4441)) + ((n_n4444) & (n_n4448) & (!n_n4447) & (n_n4442) & (!n_n4441)) + ((n_n4444) & (n_n4448) & (!n_n4447) & (n_n4442) & (n_n4441)) + ((n_n4444) & (n_n4448) & (n_n4447) & (!n_n4442) & (!n_n4441)) + ((n_n4444) & (n_n4448) & (n_n4447) & (!n_n4442) & (n_n4441)) + ((n_n4444) & (n_n4448) & (n_n4447) & (n_n4442) & (!n_n4441)) + ((n_n4444) & (n_n4448) & (n_n4447) & (n_n4442) & (n_n4441)));
	assign n_n2261 = (((!n_n4450) & (!n_n4445) & (!x368x) & (x16563x)) + ((!n_n4450) & (!n_n4445) & (x368x) & (!x16563x)) + ((!n_n4450) & (!n_n4445) & (x368x) & (x16563x)) + ((!n_n4450) & (n_n4445) & (!x368x) & (!x16563x)) + ((!n_n4450) & (n_n4445) & (!x368x) & (x16563x)) + ((!n_n4450) & (n_n4445) & (x368x) & (!x16563x)) + ((!n_n4450) & (n_n4445) & (x368x) & (x16563x)) + ((n_n4450) & (!n_n4445) & (!x368x) & (!x16563x)) + ((n_n4450) & (!n_n4445) & (!x368x) & (x16563x)) + ((n_n4450) & (!n_n4445) & (x368x) & (!x16563x)) + ((n_n4450) & (!n_n4445) & (x368x) & (x16563x)) + ((n_n4450) & (n_n4445) & (!x368x) & (!x16563x)) + ((n_n4450) & (n_n4445) & (!x368x) & (x16563x)) + ((n_n4450) & (n_n4445) & (x368x) & (!x16563x)) + ((n_n4450) & (n_n4445) & (x368x) & (x16563x)));
	assign n_n4466 = (((i_9_) & (n_n524) & (n_n518) & (n_n455)));
	assign x147x = (((!i_9_) & (n_n518) & (!n_n526) & (n_n455) & (n_n528)) + ((!i_9_) & (n_n518) & (n_n526) & (n_n455) & (n_n528)) + ((i_9_) & (n_n518) & (n_n526) & (n_n455) & (!n_n528)) + ((i_9_) & (n_n518) & (n_n526) & (n_n455) & (n_n528)));
	assign n_n3889 = (((!i_9_) & (n_n455) & (n_n535) & (n_n522) & (!n_n520)) + ((!i_9_) & (n_n455) & (n_n535) & (n_n522) & (n_n520)) + ((i_9_) & (n_n455) & (n_n535) & (!n_n522) & (n_n520)) + ((i_9_) & (n_n455) & (n_n535) & (n_n522) & (!n_n520)) + ((i_9_) & (n_n455) & (n_n535) & (n_n522) & (n_n520)));
	assign x321x = (((!n_n4455) & (!n_n3889) & (!n_n4456) & (!n_n4457) & (n_n4462)) + ((!n_n4455) & (!n_n3889) & (!n_n4456) & (n_n4457) & (!n_n4462)) + ((!n_n4455) & (!n_n3889) & (!n_n4456) & (n_n4457) & (n_n4462)) + ((!n_n4455) & (!n_n3889) & (n_n4456) & (!n_n4457) & (!n_n4462)) + ((!n_n4455) & (!n_n3889) & (n_n4456) & (!n_n4457) & (n_n4462)) + ((!n_n4455) & (!n_n3889) & (n_n4456) & (n_n4457) & (!n_n4462)) + ((!n_n4455) & (!n_n3889) & (n_n4456) & (n_n4457) & (n_n4462)) + ((!n_n4455) & (n_n3889) & (!n_n4456) & (!n_n4457) & (!n_n4462)) + ((!n_n4455) & (n_n3889) & (!n_n4456) & (!n_n4457) & (n_n4462)) + ((!n_n4455) & (n_n3889) & (!n_n4456) & (n_n4457) & (!n_n4462)) + ((!n_n4455) & (n_n3889) & (!n_n4456) & (n_n4457) & (n_n4462)) + ((!n_n4455) & (n_n3889) & (n_n4456) & (!n_n4457) & (!n_n4462)) + ((!n_n4455) & (n_n3889) & (n_n4456) & (!n_n4457) & (n_n4462)) + ((!n_n4455) & (n_n3889) & (n_n4456) & (n_n4457) & (!n_n4462)) + ((!n_n4455) & (n_n3889) & (n_n4456) & (n_n4457) & (n_n4462)) + ((n_n4455) & (!n_n3889) & (!n_n4456) & (!n_n4457) & (!n_n4462)) + ((n_n4455) & (!n_n3889) & (!n_n4456) & (!n_n4457) & (n_n4462)) + ((n_n4455) & (!n_n3889) & (!n_n4456) & (n_n4457) & (!n_n4462)) + ((n_n4455) & (!n_n3889) & (!n_n4456) & (n_n4457) & (n_n4462)) + ((n_n4455) & (!n_n3889) & (n_n4456) & (!n_n4457) & (!n_n4462)) + ((n_n4455) & (!n_n3889) & (n_n4456) & (!n_n4457) & (n_n4462)) + ((n_n4455) & (!n_n3889) & (n_n4456) & (n_n4457) & (!n_n4462)) + ((n_n4455) & (!n_n3889) & (n_n4456) & (n_n4457) & (n_n4462)) + ((n_n4455) & (n_n3889) & (!n_n4456) & (!n_n4457) & (!n_n4462)) + ((n_n4455) & (n_n3889) & (!n_n4456) & (!n_n4457) & (n_n4462)) + ((n_n4455) & (n_n3889) & (!n_n4456) & (n_n4457) & (!n_n4462)) + ((n_n4455) & (n_n3889) & (!n_n4456) & (n_n4457) & (n_n4462)) + ((n_n4455) & (n_n3889) & (n_n4456) & (!n_n4457) & (!n_n4462)) + ((n_n4455) & (n_n3889) & (n_n4456) & (!n_n4457) & (n_n4462)) + ((n_n4455) & (n_n3889) & (n_n4456) & (n_n4457) & (!n_n4462)) + ((n_n4455) & (n_n3889) & (n_n4456) & (n_n4457) & (n_n4462)));
	assign n_n4468 = (((i_9_) & (n_n518) & (n_n455) & (n_n522)));
	assign x412x = (((!i_9_) & (n_n524) & (n_n518) & (n_n455) & (!n_n522)) + ((!i_9_) & (n_n524) & (n_n518) & (n_n455) & (n_n522)) + ((i_9_) & (!n_n524) & (n_n518) & (n_n455) & (n_n522)) + ((i_9_) & (n_n524) & (n_n518) & (n_n455) & (n_n522)));
	assign x16568x = (((!n_n4459) & (!n_n4470) & (!n_n4460) & (n_n4473)) + ((!n_n4459) & (!n_n4470) & (n_n4460) & (!n_n4473)) + ((!n_n4459) & (!n_n4470) & (n_n4460) & (n_n4473)) + ((!n_n4459) & (n_n4470) & (!n_n4460) & (!n_n4473)) + ((!n_n4459) & (n_n4470) & (!n_n4460) & (n_n4473)) + ((!n_n4459) & (n_n4470) & (n_n4460) & (!n_n4473)) + ((!n_n4459) & (n_n4470) & (n_n4460) & (n_n4473)) + ((n_n4459) & (!n_n4470) & (!n_n4460) & (!n_n4473)) + ((n_n4459) & (!n_n4470) & (!n_n4460) & (n_n4473)) + ((n_n4459) & (!n_n4470) & (n_n4460) & (!n_n4473)) + ((n_n4459) & (!n_n4470) & (n_n4460) & (n_n4473)) + ((n_n4459) & (n_n4470) & (!n_n4460) & (!n_n4473)) + ((n_n4459) & (n_n4470) & (!n_n4460) & (n_n4473)) + ((n_n4459) & (n_n4470) & (n_n4460) & (!n_n4473)) + ((n_n4459) & (n_n4470) & (n_n4460) & (n_n4473)));
	assign x16569x = (((!n_n4466) & (!x147x) & (!x412x) & (!n_n4471) & (n_n4472)) + ((!n_n4466) & (!x147x) & (!x412x) & (n_n4471) & (!n_n4472)) + ((!n_n4466) & (!x147x) & (!x412x) & (n_n4471) & (n_n4472)) + ((!n_n4466) & (!x147x) & (x412x) & (!n_n4471) & (!n_n4472)) + ((!n_n4466) & (!x147x) & (x412x) & (!n_n4471) & (n_n4472)) + ((!n_n4466) & (!x147x) & (x412x) & (n_n4471) & (!n_n4472)) + ((!n_n4466) & (!x147x) & (x412x) & (n_n4471) & (n_n4472)) + ((!n_n4466) & (x147x) & (!x412x) & (!n_n4471) & (!n_n4472)) + ((!n_n4466) & (x147x) & (!x412x) & (!n_n4471) & (n_n4472)) + ((!n_n4466) & (x147x) & (!x412x) & (n_n4471) & (!n_n4472)) + ((!n_n4466) & (x147x) & (!x412x) & (n_n4471) & (n_n4472)) + ((!n_n4466) & (x147x) & (x412x) & (!n_n4471) & (!n_n4472)) + ((!n_n4466) & (x147x) & (x412x) & (!n_n4471) & (n_n4472)) + ((!n_n4466) & (x147x) & (x412x) & (n_n4471) & (!n_n4472)) + ((!n_n4466) & (x147x) & (x412x) & (n_n4471) & (n_n4472)) + ((n_n4466) & (!x147x) & (!x412x) & (!n_n4471) & (!n_n4472)) + ((n_n4466) & (!x147x) & (!x412x) & (!n_n4471) & (n_n4472)) + ((n_n4466) & (!x147x) & (!x412x) & (n_n4471) & (!n_n4472)) + ((n_n4466) & (!x147x) & (!x412x) & (n_n4471) & (n_n4472)) + ((n_n4466) & (!x147x) & (x412x) & (!n_n4471) & (!n_n4472)) + ((n_n4466) & (!x147x) & (x412x) & (!n_n4471) & (n_n4472)) + ((n_n4466) & (!x147x) & (x412x) & (n_n4471) & (!n_n4472)) + ((n_n4466) & (!x147x) & (x412x) & (n_n4471) & (n_n4472)) + ((n_n4466) & (x147x) & (!x412x) & (!n_n4471) & (!n_n4472)) + ((n_n4466) & (x147x) & (!x412x) & (!n_n4471) & (n_n4472)) + ((n_n4466) & (x147x) & (!x412x) & (n_n4471) & (!n_n4472)) + ((n_n4466) & (x147x) & (!x412x) & (n_n4471) & (n_n4472)) + ((n_n4466) & (x147x) & (x412x) & (!n_n4471) & (!n_n4472)) + ((n_n4466) & (x147x) & (x412x) & (!n_n4471) & (n_n4472)) + ((n_n4466) & (x147x) & (x412x) & (n_n4471) & (!n_n4472)) + ((n_n4466) & (x147x) & (x412x) & (n_n4471) & (n_n4472)));
	assign n_n4895 = (((!i_9_) & (n_n528) & (n_n260) & (n_n491)));
	assign n_n4890 = (((i_9_) & (n_n532) & (n_n260) & (n_n491)));
	assign x260x = (((!i_9_) & (n_n260) & (!n_n520) & (x23x) & (n_n500)) + ((!i_9_) & (n_n260) & (n_n520) & (x23x) & (n_n500)) + ((i_9_) & (n_n260) & (!n_n520) & (x23x) & (n_n500)) + ((i_9_) & (n_n260) & (n_n520) & (!x23x) & (n_n500)) + ((i_9_) & (n_n260) & (n_n520) & (x23x) & (n_n500)));
	assign x16330x = (((!i_9_) & (n_n528) & (!n_n532) & (n_n260) & (n_n491)) + ((!i_9_) & (n_n528) & (n_n532) & (n_n260) & (n_n491)) + ((i_9_) & (!n_n528) & (n_n532) & (n_n260) & (n_n491)) + ((i_9_) & (n_n528) & (n_n532) & (n_n260) & (n_n491)));
	assign n_n2226 = (((!n_n4888) & (!n_n4885) & (!n_n3451) & (!x260x) & (x16330x)) + ((!n_n4888) & (!n_n4885) & (!n_n3451) & (x260x) & (!x16330x)) + ((!n_n4888) & (!n_n4885) & (!n_n3451) & (x260x) & (x16330x)) + ((!n_n4888) & (!n_n4885) & (n_n3451) & (!x260x) & (!x16330x)) + ((!n_n4888) & (!n_n4885) & (n_n3451) & (!x260x) & (x16330x)) + ((!n_n4888) & (!n_n4885) & (n_n3451) & (x260x) & (!x16330x)) + ((!n_n4888) & (!n_n4885) & (n_n3451) & (x260x) & (x16330x)) + ((!n_n4888) & (n_n4885) & (!n_n3451) & (!x260x) & (!x16330x)) + ((!n_n4888) & (n_n4885) & (!n_n3451) & (!x260x) & (x16330x)) + ((!n_n4888) & (n_n4885) & (!n_n3451) & (x260x) & (!x16330x)) + ((!n_n4888) & (n_n4885) & (!n_n3451) & (x260x) & (x16330x)) + ((!n_n4888) & (n_n4885) & (n_n3451) & (!x260x) & (!x16330x)) + ((!n_n4888) & (n_n4885) & (n_n3451) & (!x260x) & (x16330x)) + ((!n_n4888) & (n_n4885) & (n_n3451) & (x260x) & (!x16330x)) + ((!n_n4888) & (n_n4885) & (n_n3451) & (x260x) & (x16330x)) + ((n_n4888) & (!n_n4885) & (!n_n3451) & (!x260x) & (!x16330x)) + ((n_n4888) & (!n_n4885) & (!n_n3451) & (!x260x) & (x16330x)) + ((n_n4888) & (!n_n4885) & (!n_n3451) & (x260x) & (!x16330x)) + ((n_n4888) & (!n_n4885) & (!n_n3451) & (x260x) & (x16330x)) + ((n_n4888) & (!n_n4885) & (n_n3451) & (!x260x) & (!x16330x)) + ((n_n4888) & (!n_n4885) & (n_n3451) & (!x260x) & (x16330x)) + ((n_n4888) & (!n_n4885) & (n_n3451) & (x260x) & (!x16330x)) + ((n_n4888) & (!n_n4885) & (n_n3451) & (x260x) & (x16330x)) + ((n_n4888) & (n_n4885) & (!n_n3451) & (!x260x) & (!x16330x)) + ((n_n4888) & (n_n4885) & (!n_n3451) & (!x260x) & (x16330x)) + ((n_n4888) & (n_n4885) & (!n_n3451) & (x260x) & (!x16330x)) + ((n_n4888) & (n_n4885) & (!n_n3451) & (x260x) & (x16330x)) + ((n_n4888) & (n_n4885) & (n_n3451) & (!x260x) & (!x16330x)) + ((n_n4888) & (n_n4885) & (n_n3451) & (!x260x) & (x16330x)) + ((n_n4888) & (n_n4885) & (n_n3451) & (x260x) & (!x16330x)) + ((n_n4888) & (n_n4885) & (n_n3451) & (x260x) & (x16330x)));
	assign n_n4850 = (((i_9_) & (n_n524) & (n_n518) & (n_n260)));
	assign n_n4852 = (((i_9_) & (n_n518) & (n_n260) & (n_n522)));
	assign x277x = (((!i_9_) & (n_n518) & (n_n260) & (!n_n522) & (x20x)) + ((!i_9_) & (n_n518) & (n_n260) & (n_n522) & (x20x)) + ((i_9_) & (n_n518) & (n_n260) & (!n_n522) & (x20x)) + ((i_9_) & (n_n518) & (n_n260) & (n_n522) & (!x20x)) + ((i_9_) & (n_n518) & (n_n260) & (n_n522) & (x20x)));
	assign x295x = (((!i_7_) & (i_8_) & (!i_6_) & (n_n509) & (x17x)) + ((i_7_) & (!i_8_) & (!i_6_) & (n_n509) & (x17x)));
	assign x16336x = (((!n_n4862) & (!n_n4859) & (!n_n4864) & (!n_n4861) & (n_n4850)) + ((!n_n4862) & (!n_n4859) & (!n_n4864) & (n_n4861) & (!n_n4850)) + ((!n_n4862) & (!n_n4859) & (!n_n4864) & (n_n4861) & (n_n4850)) + ((!n_n4862) & (!n_n4859) & (n_n4864) & (!n_n4861) & (!n_n4850)) + ((!n_n4862) & (!n_n4859) & (n_n4864) & (!n_n4861) & (n_n4850)) + ((!n_n4862) & (!n_n4859) & (n_n4864) & (n_n4861) & (!n_n4850)) + ((!n_n4862) & (!n_n4859) & (n_n4864) & (n_n4861) & (n_n4850)) + ((!n_n4862) & (n_n4859) & (!n_n4864) & (!n_n4861) & (!n_n4850)) + ((!n_n4862) & (n_n4859) & (!n_n4864) & (!n_n4861) & (n_n4850)) + ((!n_n4862) & (n_n4859) & (!n_n4864) & (n_n4861) & (!n_n4850)) + ((!n_n4862) & (n_n4859) & (!n_n4864) & (n_n4861) & (n_n4850)) + ((!n_n4862) & (n_n4859) & (n_n4864) & (!n_n4861) & (!n_n4850)) + ((!n_n4862) & (n_n4859) & (n_n4864) & (!n_n4861) & (n_n4850)) + ((!n_n4862) & (n_n4859) & (n_n4864) & (n_n4861) & (!n_n4850)) + ((!n_n4862) & (n_n4859) & (n_n4864) & (n_n4861) & (n_n4850)) + ((n_n4862) & (!n_n4859) & (!n_n4864) & (!n_n4861) & (!n_n4850)) + ((n_n4862) & (!n_n4859) & (!n_n4864) & (!n_n4861) & (n_n4850)) + ((n_n4862) & (!n_n4859) & (!n_n4864) & (n_n4861) & (!n_n4850)) + ((n_n4862) & (!n_n4859) & (!n_n4864) & (n_n4861) & (n_n4850)) + ((n_n4862) & (!n_n4859) & (n_n4864) & (!n_n4861) & (!n_n4850)) + ((n_n4862) & (!n_n4859) & (n_n4864) & (!n_n4861) & (n_n4850)) + ((n_n4862) & (!n_n4859) & (n_n4864) & (n_n4861) & (!n_n4850)) + ((n_n4862) & (!n_n4859) & (n_n4864) & (n_n4861) & (n_n4850)) + ((n_n4862) & (n_n4859) & (!n_n4864) & (!n_n4861) & (!n_n4850)) + ((n_n4862) & (n_n4859) & (!n_n4864) & (!n_n4861) & (n_n4850)) + ((n_n4862) & (n_n4859) & (!n_n4864) & (n_n4861) & (!n_n4850)) + ((n_n4862) & (n_n4859) & (!n_n4864) & (n_n4861) & (n_n4850)) + ((n_n4862) & (n_n4859) & (n_n4864) & (!n_n4861) & (!n_n4850)) + ((n_n4862) & (n_n4859) & (n_n4864) & (!n_n4861) & (n_n4850)) + ((n_n4862) & (n_n4859) & (n_n4864) & (n_n4861) & (!n_n4850)) + ((n_n4862) & (n_n4859) & (n_n4864) & (n_n4861) & (n_n4850)));
	assign n_n2228 = (((!n_n4853) & (!n_n4852) & (!x295x) & (x16336x)) + ((!n_n4853) & (!n_n4852) & (x295x) & (!x16336x)) + ((!n_n4853) & (!n_n4852) & (x295x) & (x16336x)) + ((!n_n4853) & (n_n4852) & (!x295x) & (!x16336x)) + ((!n_n4853) & (n_n4852) & (!x295x) & (x16336x)) + ((!n_n4853) & (n_n4852) & (x295x) & (!x16336x)) + ((!n_n4853) & (n_n4852) & (x295x) & (x16336x)) + ((n_n4853) & (!n_n4852) & (!x295x) & (!x16336x)) + ((n_n4853) & (!n_n4852) & (!x295x) & (x16336x)) + ((n_n4853) & (!n_n4852) & (x295x) & (!x16336x)) + ((n_n4853) & (!n_n4852) & (x295x) & (x16336x)) + ((n_n4853) & (n_n4852) & (!x295x) & (!x16336x)) + ((n_n4853) & (n_n4852) & (!x295x) & (x16336x)) + ((n_n4853) & (n_n4852) & (x295x) & (!x16336x)) + ((n_n4853) & (n_n4852) & (x295x) & (x16336x)));
	assign n_n4881 = (((!i_9_) & (n_n526) & (n_n260) & (n_n500)));
	assign n_n4878 = (((i_9_) & (n_n528) & (n_n260) & (n_n500)));
	assign n_n4880 = (((i_9_) & (n_n526) & (n_n260) & (n_n500)));
	assign n_n4877 = (((!i_9_) & (n_n260) & (n_n500) & (n_n530)));
	assign n_n4872 = (((i_9_) & (n_n534) & (n_n260) & (n_n500)));
	assign n_n4875 = (((!i_9_) & (n_n532) & (n_n260) & (n_n500)));
	assign n_n4873 = (((!i_9_) & (n_n534) & (n_n260) & (n_n500)));
	assign x174x = (((!i_9_) & (!n_n532) & (n_n534) & (n_n260) & (n_n500)) + ((!i_9_) & (n_n532) & (!n_n534) & (n_n260) & (n_n500)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n260) & (n_n500)));
	assign x16340x = (((!n_n4881) & (!n_n4878) & (!n_n4875) & (n_n4873)) + ((!n_n4881) & (!n_n4878) & (n_n4875) & (!n_n4873)) + ((!n_n4881) & (!n_n4878) & (n_n4875) & (n_n4873)) + ((!n_n4881) & (n_n4878) & (!n_n4875) & (!n_n4873)) + ((!n_n4881) & (n_n4878) & (!n_n4875) & (n_n4873)) + ((!n_n4881) & (n_n4878) & (n_n4875) & (!n_n4873)) + ((!n_n4881) & (n_n4878) & (n_n4875) & (n_n4873)) + ((n_n4881) & (!n_n4878) & (!n_n4875) & (!n_n4873)) + ((n_n4881) & (!n_n4878) & (!n_n4875) & (n_n4873)) + ((n_n4881) & (!n_n4878) & (n_n4875) & (!n_n4873)) + ((n_n4881) & (!n_n4878) & (n_n4875) & (n_n4873)) + ((n_n4881) & (n_n4878) & (!n_n4875) & (!n_n4873)) + ((n_n4881) & (n_n4878) & (!n_n4875) & (n_n4873)) + ((n_n4881) & (n_n4878) & (n_n4875) & (!n_n4873)) + ((n_n4881) & (n_n4878) & (n_n4875) & (n_n4873)));
	assign x16341x = (((!n_n4869) & (!n_n4870) & (!n_n4880) & (!n_n4877) & (n_n4872)) + ((!n_n4869) & (!n_n4870) & (!n_n4880) & (n_n4877) & (!n_n4872)) + ((!n_n4869) & (!n_n4870) & (!n_n4880) & (n_n4877) & (n_n4872)) + ((!n_n4869) & (!n_n4870) & (n_n4880) & (!n_n4877) & (!n_n4872)) + ((!n_n4869) & (!n_n4870) & (n_n4880) & (!n_n4877) & (n_n4872)) + ((!n_n4869) & (!n_n4870) & (n_n4880) & (n_n4877) & (!n_n4872)) + ((!n_n4869) & (!n_n4870) & (n_n4880) & (n_n4877) & (n_n4872)) + ((!n_n4869) & (n_n4870) & (!n_n4880) & (!n_n4877) & (!n_n4872)) + ((!n_n4869) & (n_n4870) & (!n_n4880) & (!n_n4877) & (n_n4872)) + ((!n_n4869) & (n_n4870) & (!n_n4880) & (n_n4877) & (!n_n4872)) + ((!n_n4869) & (n_n4870) & (!n_n4880) & (n_n4877) & (n_n4872)) + ((!n_n4869) & (n_n4870) & (n_n4880) & (!n_n4877) & (!n_n4872)) + ((!n_n4869) & (n_n4870) & (n_n4880) & (!n_n4877) & (n_n4872)) + ((!n_n4869) & (n_n4870) & (n_n4880) & (n_n4877) & (!n_n4872)) + ((!n_n4869) & (n_n4870) & (n_n4880) & (n_n4877) & (n_n4872)) + ((n_n4869) & (!n_n4870) & (!n_n4880) & (!n_n4877) & (!n_n4872)) + ((n_n4869) & (!n_n4870) & (!n_n4880) & (!n_n4877) & (n_n4872)) + ((n_n4869) & (!n_n4870) & (!n_n4880) & (n_n4877) & (!n_n4872)) + ((n_n4869) & (!n_n4870) & (!n_n4880) & (n_n4877) & (n_n4872)) + ((n_n4869) & (!n_n4870) & (n_n4880) & (!n_n4877) & (!n_n4872)) + ((n_n4869) & (!n_n4870) & (n_n4880) & (!n_n4877) & (n_n4872)) + ((n_n4869) & (!n_n4870) & (n_n4880) & (n_n4877) & (!n_n4872)) + ((n_n4869) & (!n_n4870) & (n_n4880) & (n_n4877) & (n_n4872)) + ((n_n4869) & (n_n4870) & (!n_n4880) & (!n_n4877) & (!n_n4872)) + ((n_n4869) & (n_n4870) & (!n_n4880) & (!n_n4877) & (n_n4872)) + ((n_n4869) & (n_n4870) & (!n_n4880) & (n_n4877) & (!n_n4872)) + ((n_n4869) & (n_n4870) & (!n_n4880) & (n_n4877) & (n_n4872)) + ((n_n4869) & (n_n4870) & (n_n4880) & (!n_n4877) & (!n_n4872)) + ((n_n4869) & (n_n4870) & (n_n4880) & (!n_n4877) & (n_n4872)) + ((n_n4869) & (n_n4870) & (n_n4880) & (n_n4877) & (!n_n4872)) + ((n_n4869) & (n_n4870) & (n_n4880) & (n_n4877) & (n_n4872)));
	assign n_n2178 = (((!n_n2226) & (!n_n2228) & (!x16340x) & (x16341x)) + ((!n_n2226) & (!n_n2228) & (x16340x) & (!x16341x)) + ((!n_n2226) & (!n_n2228) & (x16340x) & (x16341x)) + ((!n_n2226) & (n_n2228) & (!x16340x) & (!x16341x)) + ((!n_n2226) & (n_n2228) & (!x16340x) & (x16341x)) + ((!n_n2226) & (n_n2228) & (x16340x) & (!x16341x)) + ((!n_n2226) & (n_n2228) & (x16340x) & (x16341x)) + ((n_n2226) & (!n_n2228) & (!x16340x) & (!x16341x)) + ((n_n2226) & (!n_n2228) & (!x16340x) & (x16341x)) + ((n_n2226) & (!n_n2228) & (x16340x) & (!x16341x)) + ((n_n2226) & (!n_n2228) & (x16340x) & (x16341x)) + ((n_n2226) & (n_n2228) & (!x16340x) & (!x16341x)) + ((n_n2226) & (n_n2228) & (!x16340x) & (x16341x)) + ((n_n2226) & (n_n2228) & (x16340x) & (!x16341x)) + ((n_n2226) & (n_n2228) & (x16340x) & (x16341x)));
	assign n_n5322 = (((i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n464)));
	assign n_n2274 = (((!i_9_) & (!n_n532) & (!n_n464) & (!n_n65) & (n_n5324)) + ((!i_9_) & (!n_n532) & (!n_n464) & (n_n65) & (n_n5324)) + ((!i_9_) & (!n_n532) & (n_n464) & (!n_n65) & (n_n5324)) + ((!i_9_) & (!n_n532) & (n_n464) & (n_n65) & (n_n5324)) + ((!i_9_) & (n_n532) & (!n_n464) & (!n_n65) & (n_n5324)) + ((!i_9_) & (n_n532) & (!n_n464) & (n_n65) & (n_n5324)) + ((!i_9_) & (n_n532) & (n_n464) & (!n_n65) & (n_n5324)) + ((!i_9_) & (n_n532) & (n_n464) & (n_n65) & (!n_n5324)) + ((!i_9_) & (n_n532) & (n_n464) & (n_n65) & (n_n5324)) + ((i_9_) & (!n_n532) & (!n_n464) & (!n_n65) & (n_n5324)) + ((i_9_) & (!n_n532) & (!n_n464) & (n_n65) & (n_n5324)) + ((i_9_) & (!n_n532) & (n_n464) & (!n_n65) & (n_n5324)) + ((i_9_) & (!n_n532) & (n_n464) & (n_n65) & (n_n5324)) + ((i_9_) & (n_n532) & (!n_n464) & (!n_n65) & (n_n5324)) + ((i_9_) & (n_n532) & (!n_n464) & (n_n65) & (n_n5324)) + ((i_9_) & (n_n532) & (n_n464) & (!n_n65) & (n_n5324)) + ((i_9_) & (n_n532) & (n_n464) & (n_n65) & (!n_n5324)) + ((i_9_) & (n_n532) & (n_n464) & (n_n65) & (n_n5324)));
	assign n_n5326 = (((!i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n464)));
	assign n_n5325 = (((!i_9_) & (n_n530) & (n_n464) & (n_n65)));
	assign n_n5332 = (((!i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n464)));
	assign n_n5329 = (((!i_9_) & (n_n526) & (n_n464) & (n_n65)));
	assign x115x = (((!x19x) & (n_n473) & (!n_n522) & (x20x) & (n_n65)) + ((!x19x) & (n_n473) & (n_n522) & (x20x) & (n_n65)) + ((x19x) & (n_n473) & (!n_n522) & (x20x) & (n_n65)) + ((x19x) & (n_n473) & (n_n522) & (!x20x) & (!n_n65)) + ((x19x) & (n_n473) & (n_n522) & (!x20x) & (n_n65)) + ((x19x) & (n_n473) & (n_n522) & (x20x) & (!n_n65)) + ((x19x) & (n_n473) & (n_n522) & (x20x) & (n_n65)));
	assign x16292x = (((!i_9_) & (!n_n526) & (!n_n473) & (!n_n65) & (x115x)) + ((!i_9_) & (!n_n526) & (!n_n473) & (n_n65) & (x115x)) + ((!i_9_) & (!n_n526) & (n_n473) & (!n_n65) & (x115x)) + ((!i_9_) & (!n_n526) & (n_n473) & (n_n65) & (x115x)) + ((!i_9_) & (n_n526) & (!n_n473) & (!n_n65) & (x115x)) + ((!i_9_) & (n_n526) & (!n_n473) & (n_n65) & (x115x)) + ((!i_9_) & (n_n526) & (n_n473) & (!n_n65) & (x115x)) + ((!i_9_) & (n_n526) & (n_n473) & (n_n65) & (!x115x)) + ((!i_9_) & (n_n526) & (n_n473) & (n_n65) & (x115x)) + ((i_9_) & (!n_n526) & (!n_n473) & (!n_n65) & (x115x)) + ((i_9_) & (!n_n526) & (!n_n473) & (n_n65) & (x115x)) + ((i_9_) & (!n_n526) & (n_n473) & (!n_n65) & (x115x)) + ((i_9_) & (!n_n526) & (n_n473) & (n_n65) & (x115x)) + ((i_9_) & (n_n526) & (!n_n473) & (!n_n65) & (x115x)) + ((i_9_) & (n_n526) & (!n_n473) & (n_n65) & (x115x)) + ((i_9_) & (n_n526) & (n_n473) & (!n_n65) & (x115x)) + ((i_9_) & (n_n526) & (n_n473) & (n_n65) & (!x115x)) + ((i_9_) & (n_n526) & (n_n473) & (n_n65) & (x115x)));
	assign n_n5315 = (((!i_9_) & (n_n524) & (n_n473) & (n_n65)));
	assign x117x = (((!x19x) & (!n_n524) & (!n_n473) & (!x16292x) & (n_n5315)) + ((!x19x) & (!n_n524) & (!n_n473) & (x16292x) & (!n_n5315)) + ((!x19x) & (!n_n524) & (!n_n473) & (x16292x) & (n_n5315)) + ((!x19x) & (!n_n524) & (n_n473) & (!x16292x) & (n_n5315)) + ((!x19x) & (!n_n524) & (n_n473) & (x16292x) & (!n_n5315)) + ((!x19x) & (!n_n524) & (n_n473) & (x16292x) & (n_n5315)) + ((!x19x) & (n_n524) & (!n_n473) & (!x16292x) & (n_n5315)) + ((!x19x) & (n_n524) & (!n_n473) & (x16292x) & (!n_n5315)) + ((!x19x) & (n_n524) & (!n_n473) & (x16292x) & (n_n5315)) + ((!x19x) & (n_n524) & (n_n473) & (!x16292x) & (n_n5315)) + ((!x19x) & (n_n524) & (n_n473) & (x16292x) & (!n_n5315)) + ((!x19x) & (n_n524) & (n_n473) & (x16292x) & (n_n5315)) + ((x19x) & (!n_n524) & (!n_n473) & (!x16292x) & (n_n5315)) + ((x19x) & (!n_n524) & (!n_n473) & (x16292x) & (!n_n5315)) + ((x19x) & (!n_n524) & (!n_n473) & (x16292x) & (n_n5315)) + ((x19x) & (!n_n524) & (n_n473) & (!x16292x) & (n_n5315)) + ((x19x) & (!n_n524) & (n_n473) & (x16292x) & (!n_n5315)) + ((x19x) & (!n_n524) & (n_n473) & (x16292x) & (n_n5315)) + ((x19x) & (n_n524) & (!n_n473) & (!x16292x) & (n_n5315)) + ((x19x) & (n_n524) & (!n_n473) & (x16292x) & (!n_n5315)) + ((x19x) & (n_n524) & (!n_n473) & (x16292x) & (n_n5315)) + ((x19x) & (n_n524) & (n_n473) & (!x16292x) & (!n_n5315)) + ((x19x) & (n_n524) & (n_n473) & (!x16292x) & (n_n5315)) + ((x19x) & (n_n524) & (n_n473) & (x16292x) & (!n_n5315)) + ((x19x) & (n_n524) & (n_n473) & (x16292x) & (n_n5315)));
	assign n_n5311 = (((!i_9_) & (n_n528) & (n_n473) & (n_n65)));
	assign n_n5302 = (((!i_5_) & (!i_3_) & (i_4_) & (x19x) & (n_n520)));
	assign n_n5303 = (((!i_5_) & (!i_3_) & (i_4_) & (x23x) & (n_n65)));
	assign n_n5306 = (((i_5_) & (!i_3_) & (!i_4_) & (x19x) & (n_n532)));
	assign n_n5304 = (((i_5_) & (!i_3_) & (!i_4_) & (x19x) & (n_n534)));
	assign x462x = (((!n_n5302) & (!n_n5303) & (!n_n5306) & (!x63x) & (n_n5304)) + ((!n_n5302) & (!n_n5303) & (!n_n5306) & (x63x) & (!n_n5304)) + ((!n_n5302) & (!n_n5303) & (!n_n5306) & (x63x) & (n_n5304)) + ((!n_n5302) & (!n_n5303) & (n_n5306) & (!x63x) & (!n_n5304)) + ((!n_n5302) & (!n_n5303) & (n_n5306) & (!x63x) & (n_n5304)) + ((!n_n5302) & (!n_n5303) & (n_n5306) & (x63x) & (!n_n5304)) + ((!n_n5302) & (!n_n5303) & (n_n5306) & (x63x) & (n_n5304)) + ((!n_n5302) & (n_n5303) & (!n_n5306) & (!x63x) & (!n_n5304)) + ((!n_n5302) & (n_n5303) & (!n_n5306) & (!x63x) & (n_n5304)) + ((!n_n5302) & (n_n5303) & (!n_n5306) & (x63x) & (!n_n5304)) + ((!n_n5302) & (n_n5303) & (!n_n5306) & (x63x) & (n_n5304)) + ((!n_n5302) & (n_n5303) & (n_n5306) & (!x63x) & (!n_n5304)) + ((!n_n5302) & (n_n5303) & (n_n5306) & (!x63x) & (n_n5304)) + ((!n_n5302) & (n_n5303) & (n_n5306) & (x63x) & (!n_n5304)) + ((!n_n5302) & (n_n5303) & (n_n5306) & (x63x) & (n_n5304)) + ((n_n5302) & (!n_n5303) & (!n_n5306) & (!x63x) & (!n_n5304)) + ((n_n5302) & (!n_n5303) & (!n_n5306) & (!x63x) & (n_n5304)) + ((n_n5302) & (!n_n5303) & (!n_n5306) & (x63x) & (!n_n5304)) + ((n_n5302) & (!n_n5303) & (!n_n5306) & (x63x) & (n_n5304)) + ((n_n5302) & (!n_n5303) & (n_n5306) & (!x63x) & (!n_n5304)) + ((n_n5302) & (!n_n5303) & (n_n5306) & (!x63x) & (n_n5304)) + ((n_n5302) & (!n_n5303) & (n_n5306) & (x63x) & (!n_n5304)) + ((n_n5302) & (!n_n5303) & (n_n5306) & (x63x) & (n_n5304)) + ((n_n5302) & (n_n5303) & (!n_n5306) & (!x63x) & (!n_n5304)) + ((n_n5302) & (n_n5303) & (!n_n5306) & (!x63x) & (n_n5304)) + ((n_n5302) & (n_n5303) & (!n_n5306) & (x63x) & (!n_n5304)) + ((n_n5302) & (n_n5303) & (!n_n5306) & (x63x) & (n_n5304)) + ((n_n5302) & (n_n5303) & (n_n5306) & (!x63x) & (!n_n5304)) + ((n_n5302) & (n_n5303) & (n_n5306) & (!x63x) & (n_n5304)) + ((n_n5302) & (n_n5303) & (n_n5306) & (x63x) & (!n_n5304)) + ((n_n5302) & (n_n5303) & (n_n5306) & (x63x) & (n_n5304)));
	assign n_n4793 = (((!i_9_) & (n_n473) & (n_n534) & (n_n325)));
	assign n_n4804 = (((i_9_) & (n_n473) & (n_n325) & (n_n522)));
	assign n_n4794 = (((i_9_) & (n_n473) & (n_n532) & (n_n325)));
	assign n_n4795 = (((!i_9_) & (n_n473) & (n_n532) & (n_n325)));
	assign x16349x = (((!n_n4793) & (!n_n4804) & (!n_n4794) & (n_n4795)) + ((!n_n4793) & (!n_n4804) & (n_n4794) & (!n_n4795)) + ((!n_n4793) & (!n_n4804) & (n_n4794) & (n_n4795)) + ((!n_n4793) & (n_n4804) & (!n_n4794) & (!n_n4795)) + ((!n_n4793) & (n_n4804) & (!n_n4794) & (n_n4795)) + ((!n_n4793) & (n_n4804) & (n_n4794) & (!n_n4795)) + ((!n_n4793) & (n_n4804) & (n_n4794) & (n_n4795)) + ((n_n4793) & (!n_n4804) & (!n_n4794) & (!n_n4795)) + ((n_n4793) & (!n_n4804) & (!n_n4794) & (n_n4795)) + ((n_n4793) & (!n_n4804) & (n_n4794) & (!n_n4795)) + ((n_n4793) & (!n_n4804) & (n_n4794) & (n_n4795)) + ((n_n4793) & (n_n4804) & (!n_n4794) & (!n_n4795)) + ((n_n4793) & (n_n4804) & (!n_n4794) & (n_n4795)) + ((n_n4793) & (n_n4804) & (n_n4794) & (!n_n4795)) + ((n_n4793) & (n_n4804) & (n_n4794) & (n_n4795)));
	assign n_n4798 = (((i_9_) & (n_n528) & (n_n473) & (n_n325)));
	assign n_n4796 = (((i_9_) & (n_n473) & (n_n325) & (n_n530)));
	assign n_n4797 = (((!i_9_) & (n_n473) & (n_n325) & (n_n530)));
	assign n_n4801 = (((!i_9_) & (n_n526) & (n_n473) & (n_n325)));
	assign x16350x = (((!n_n4791) & (!n_n4798) & (!n_n4796) & (!n_n4797) & (n_n4801)) + ((!n_n4791) & (!n_n4798) & (!n_n4796) & (n_n4797) & (!n_n4801)) + ((!n_n4791) & (!n_n4798) & (!n_n4796) & (n_n4797) & (n_n4801)) + ((!n_n4791) & (!n_n4798) & (n_n4796) & (!n_n4797) & (!n_n4801)) + ((!n_n4791) & (!n_n4798) & (n_n4796) & (!n_n4797) & (n_n4801)) + ((!n_n4791) & (!n_n4798) & (n_n4796) & (n_n4797) & (!n_n4801)) + ((!n_n4791) & (!n_n4798) & (n_n4796) & (n_n4797) & (n_n4801)) + ((!n_n4791) & (n_n4798) & (!n_n4796) & (!n_n4797) & (!n_n4801)) + ((!n_n4791) & (n_n4798) & (!n_n4796) & (!n_n4797) & (n_n4801)) + ((!n_n4791) & (n_n4798) & (!n_n4796) & (n_n4797) & (!n_n4801)) + ((!n_n4791) & (n_n4798) & (!n_n4796) & (n_n4797) & (n_n4801)) + ((!n_n4791) & (n_n4798) & (n_n4796) & (!n_n4797) & (!n_n4801)) + ((!n_n4791) & (n_n4798) & (n_n4796) & (!n_n4797) & (n_n4801)) + ((!n_n4791) & (n_n4798) & (n_n4796) & (n_n4797) & (!n_n4801)) + ((!n_n4791) & (n_n4798) & (n_n4796) & (n_n4797) & (n_n4801)) + ((n_n4791) & (!n_n4798) & (!n_n4796) & (!n_n4797) & (!n_n4801)) + ((n_n4791) & (!n_n4798) & (!n_n4796) & (!n_n4797) & (n_n4801)) + ((n_n4791) & (!n_n4798) & (!n_n4796) & (n_n4797) & (!n_n4801)) + ((n_n4791) & (!n_n4798) & (!n_n4796) & (n_n4797) & (n_n4801)) + ((n_n4791) & (!n_n4798) & (n_n4796) & (!n_n4797) & (!n_n4801)) + ((n_n4791) & (!n_n4798) & (n_n4796) & (!n_n4797) & (n_n4801)) + ((n_n4791) & (!n_n4798) & (n_n4796) & (n_n4797) & (!n_n4801)) + ((n_n4791) & (!n_n4798) & (n_n4796) & (n_n4797) & (n_n4801)) + ((n_n4791) & (n_n4798) & (!n_n4796) & (!n_n4797) & (!n_n4801)) + ((n_n4791) & (n_n4798) & (!n_n4796) & (!n_n4797) & (n_n4801)) + ((n_n4791) & (n_n4798) & (!n_n4796) & (n_n4797) & (!n_n4801)) + ((n_n4791) & (n_n4798) & (!n_n4796) & (n_n4797) & (n_n4801)) + ((n_n4791) & (n_n4798) & (n_n4796) & (!n_n4797) & (!n_n4801)) + ((n_n4791) & (n_n4798) & (n_n4796) & (!n_n4797) & (n_n4801)) + ((n_n4791) & (n_n4798) & (n_n4796) & (n_n4797) & (!n_n4801)) + ((n_n4791) & (n_n4798) & (n_n4796) & (n_n4797) & (n_n4801)));
	assign n_n4845 = (((!i_9_) & (n_n518) & (n_n260) & (n_n530)));
	assign x177x = (((!n_n260) & (!n_n535) & (!x23x) & (n_n4840)) + ((!n_n260) & (!n_n535) & (x23x) & (n_n4840)) + ((!n_n260) & (n_n535) & (!x23x) & (n_n4840)) + ((!n_n260) & (n_n535) & (x23x) & (n_n4840)) + ((n_n260) & (!n_n535) & (!x23x) & (n_n4840)) + ((n_n260) & (!n_n535) & (x23x) & (n_n4840)) + ((n_n260) & (n_n535) & (!x23x) & (n_n4840)) + ((n_n260) & (n_n535) & (x23x) & (!n_n4840)) + ((n_n260) & (n_n535) & (x23x) & (n_n4840)));
	assign n_n2230 = (((!n_n4834) & (!n_n4835) & (!n_n4832) & (!x185x) & (x388x)) + ((!n_n4834) & (!n_n4835) & (!n_n4832) & (x185x) & (!x388x)) + ((!n_n4834) & (!n_n4835) & (!n_n4832) & (x185x) & (x388x)) + ((!n_n4834) & (!n_n4835) & (n_n4832) & (!x185x) & (!x388x)) + ((!n_n4834) & (!n_n4835) & (n_n4832) & (!x185x) & (x388x)) + ((!n_n4834) & (!n_n4835) & (n_n4832) & (x185x) & (!x388x)) + ((!n_n4834) & (!n_n4835) & (n_n4832) & (x185x) & (x388x)) + ((!n_n4834) & (n_n4835) & (!n_n4832) & (!x185x) & (!x388x)) + ((!n_n4834) & (n_n4835) & (!n_n4832) & (!x185x) & (x388x)) + ((!n_n4834) & (n_n4835) & (!n_n4832) & (x185x) & (!x388x)) + ((!n_n4834) & (n_n4835) & (!n_n4832) & (x185x) & (x388x)) + ((!n_n4834) & (n_n4835) & (n_n4832) & (!x185x) & (!x388x)) + ((!n_n4834) & (n_n4835) & (n_n4832) & (!x185x) & (x388x)) + ((!n_n4834) & (n_n4835) & (n_n4832) & (x185x) & (!x388x)) + ((!n_n4834) & (n_n4835) & (n_n4832) & (x185x) & (x388x)) + ((n_n4834) & (!n_n4835) & (!n_n4832) & (!x185x) & (!x388x)) + ((n_n4834) & (!n_n4835) & (!n_n4832) & (!x185x) & (x388x)) + ((n_n4834) & (!n_n4835) & (!n_n4832) & (x185x) & (!x388x)) + ((n_n4834) & (!n_n4835) & (!n_n4832) & (x185x) & (x388x)) + ((n_n4834) & (!n_n4835) & (n_n4832) & (!x185x) & (!x388x)) + ((n_n4834) & (!n_n4835) & (n_n4832) & (!x185x) & (x388x)) + ((n_n4834) & (!n_n4835) & (n_n4832) & (x185x) & (!x388x)) + ((n_n4834) & (!n_n4835) & (n_n4832) & (x185x) & (x388x)) + ((n_n4834) & (n_n4835) & (!n_n4832) & (!x185x) & (!x388x)) + ((n_n4834) & (n_n4835) & (!n_n4832) & (!x185x) & (x388x)) + ((n_n4834) & (n_n4835) & (!n_n4832) & (x185x) & (!x388x)) + ((n_n4834) & (n_n4835) & (!n_n4832) & (x185x) & (x388x)) + ((n_n4834) & (n_n4835) & (n_n4832) & (!x185x) & (!x388x)) + ((n_n4834) & (n_n4835) & (n_n4832) & (!x185x) & (x388x)) + ((n_n4834) & (n_n4835) & (n_n4832) & (x185x) & (!x388x)) + ((n_n4834) & (n_n4835) & (n_n4832) & (x185x) & (x388x)));
	assign x16357x = (((!n_n4843) & (!n_n4846) & (!n_n4842) & (!n_n4841) & (n_n4837)) + ((!n_n4843) & (!n_n4846) & (!n_n4842) & (n_n4841) & (!n_n4837)) + ((!n_n4843) & (!n_n4846) & (!n_n4842) & (n_n4841) & (n_n4837)) + ((!n_n4843) & (!n_n4846) & (n_n4842) & (!n_n4841) & (!n_n4837)) + ((!n_n4843) & (!n_n4846) & (n_n4842) & (!n_n4841) & (n_n4837)) + ((!n_n4843) & (!n_n4846) & (n_n4842) & (n_n4841) & (!n_n4837)) + ((!n_n4843) & (!n_n4846) & (n_n4842) & (n_n4841) & (n_n4837)) + ((!n_n4843) & (n_n4846) & (!n_n4842) & (!n_n4841) & (!n_n4837)) + ((!n_n4843) & (n_n4846) & (!n_n4842) & (!n_n4841) & (n_n4837)) + ((!n_n4843) & (n_n4846) & (!n_n4842) & (n_n4841) & (!n_n4837)) + ((!n_n4843) & (n_n4846) & (!n_n4842) & (n_n4841) & (n_n4837)) + ((!n_n4843) & (n_n4846) & (n_n4842) & (!n_n4841) & (!n_n4837)) + ((!n_n4843) & (n_n4846) & (n_n4842) & (!n_n4841) & (n_n4837)) + ((!n_n4843) & (n_n4846) & (n_n4842) & (n_n4841) & (!n_n4837)) + ((!n_n4843) & (n_n4846) & (n_n4842) & (n_n4841) & (n_n4837)) + ((n_n4843) & (!n_n4846) & (!n_n4842) & (!n_n4841) & (!n_n4837)) + ((n_n4843) & (!n_n4846) & (!n_n4842) & (!n_n4841) & (n_n4837)) + ((n_n4843) & (!n_n4846) & (!n_n4842) & (n_n4841) & (!n_n4837)) + ((n_n4843) & (!n_n4846) & (!n_n4842) & (n_n4841) & (n_n4837)) + ((n_n4843) & (!n_n4846) & (n_n4842) & (!n_n4841) & (!n_n4837)) + ((n_n4843) & (!n_n4846) & (n_n4842) & (!n_n4841) & (n_n4837)) + ((n_n4843) & (!n_n4846) & (n_n4842) & (n_n4841) & (!n_n4837)) + ((n_n4843) & (!n_n4846) & (n_n4842) & (n_n4841) & (n_n4837)) + ((n_n4843) & (n_n4846) & (!n_n4842) & (!n_n4841) & (!n_n4837)) + ((n_n4843) & (n_n4846) & (!n_n4842) & (!n_n4841) & (n_n4837)) + ((n_n4843) & (n_n4846) & (!n_n4842) & (n_n4841) & (!n_n4837)) + ((n_n4843) & (n_n4846) & (!n_n4842) & (n_n4841) & (n_n4837)) + ((n_n4843) & (n_n4846) & (n_n4842) & (!n_n4841) & (!n_n4837)) + ((n_n4843) & (n_n4846) & (n_n4842) & (!n_n4841) & (n_n4837)) + ((n_n4843) & (n_n4846) & (n_n4842) & (n_n4841) & (!n_n4837)) + ((n_n4843) & (n_n4846) & (n_n4842) & (n_n4841) & (n_n4837)));
	assign x16365x = (((!n_n4845) & (!x177x) & (!n_n4844) & (!n_n2230) & (x16357x)) + ((!n_n4845) & (!x177x) & (!n_n4844) & (n_n2230) & (!x16357x)) + ((!n_n4845) & (!x177x) & (!n_n4844) & (n_n2230) & (x16357x)) + ((!n_n4845) & (!x177x) & (n_n4844) & (!n_n2230) & (!x16357x)) + ((!n_n4845) & (!x177x) & (n_n4844) & (!n_n2230) & (x16357x)) + ((!n_n4845) & (!x177x) & (n_n4844) & (n_n2230) & (!x16357x)) + ((!n_n4845) & (!x177x) & (n_n4844) & (n_n2230) & (x16357x)) + ((!n_n4845) & (x177x) & (!n_n4844) & (!n_n2230) & (!x16357x)) + ((!n_n4845) & (x177x) & (!n_n4844) & (!n_n2230) & (x16357x)) + ((!n_n4845) & (x177x) & (!n_n4844) & (n_n2230) & (!x16357x)) + ((!n_n4845) & (x177x) & (!n_n4844) & (n_n2230) & (x16357x)) + ((!n_n4845) & (x177x) & (n_n4844) & (!n_n2230) & (!x16357x)) + ((!n_n4845) & (x177x) & (n_n4844) & (!n_n2230) & (x16357x)) + ((!n_n4845) & (x177x) & (n_n4844) & (n_n2230) & (!x16357x)) + ((!n_n4845) & (x177x) & (n_n4844) & (n_n2230) & (x16357x)) + ((n_n4845) & (!x177x) & (!n_n4844) & (!n_n2230) & (!x16357x)) + ((n_n4845) & (!x177x) & (!n_n4844) & (!n_n2230) & (x16357x)) + ((n_n4845) & (!x177x) & (!n_n4844) & (n_n2230) & (!x16357x)) + ((n_n4845) & (!x177x) & (!n_n4844) & (n_n2230) & (x16357x)) + ((n_n4845) & (!x177x) & (n_n4844) & (!n_n2230) & (!x16357x)) + ((n_n4845) & (!x177x) & (n_n4844) & (!n_n2230) & (x16357x)) + ((n_n4845) & (!x177x) & (n_n4844) & (n_n2230) & (!x16357x)) + ((n_n4845) & (!x177x) & (n_n4844) & (n_n2230) & (x16357x)) + ((n_n4845) & (x177x) & (!n_n4844) & (!n_n2230) & (!x16357x)) + ((n_n4845) & (x177x) & (!n_n4844) & (!n_n2230) & (x16357x)) + ((n_n4845) & (x177x) & (!n_n4844) & (n_n2230) & (!x16357x)) + ((n_n4845) & (x177x) & (!n_n4844) & (n_n2230) & (x16357x)) + ((n_n4845) & (x177x) & (n_n4844) & (!n_n2230) & (!x16357x)) + ((n_n4845) & (x177x) & (n_n4844) & (!n_n2230) & (x16357x)) + ((n_n4845) & (x177x) & (n_n4844) & (n_n2230) & (!x16357x)) + ((n_n4845) & (x177x) & (n_n4844) & (n_n2230) & (x16357x)));
	assign n_n4767 = (((!i_9_) & (n_n528) & (n_n325) & (n_n491)));
	assign n_n4763 = (((!i_9_) & (n_n532) & (n_n325) & (n_n491)));
	assign n_n3469 = (((!i_9_) & (!n_n524) & (n_n325) & (n_n491) & (x20x)) + ((!i_9_) & (n_n524) & (n_n325) & (n_n491) & (!x20x)) + ((!i_9_) & (n_n524) & (n_n325) & (n_n491) & (x20x)) + ((i_9_) & (!n_n524) & (n_n325) & (n_n491) & (x20x)) + ((i_9_) & (n_n524) & (n_n325) & (n_n491) & (!x20x)) + ((i_9_) & (n_n524) & (n_n325) & (n_n491) & (x20x)));
	assign x164x = (((!i_9_) & (n_n526) & (n_n325) & (n_n491)) + ((i_9_) & (n_n526) & (n_n325) & (n_n491)));
	assign n_n2234 = (((!n_n4767) & (!x165x) & (!n_n4763) & (!n_n3469) & (x164x)) + ((!n_n4767) & (!x165x) & (!n_n4763) & (n_n3469) & (!x164x)) + ((!n_n4767) & (!x165x) & (!n_n4763) & (n_n3469) & (x164x)) + ((!n_n4767) & (!x165x) & (n_n4763) & (!n_n3469) & (!x164x)) + ((!n_n4767) & (!x165x) & (n_n4763) & (!n_n3469) & (x164x)) + ((!n_n4767) & (!x165x) & (n_n4763) & (n_n3469) & (!x164x)) + ((!n_n4767) & (!x165x) & (n_n4763) & (n_n3469) & (x164x)) + ((!n_n4767) & (x165x) & (!n_n4763) & (!n_n3469) & (!x164x)) + ((!n_n4767) & (x165x) & (!n_n4763) & (!n_n3469) & (x164x)) + ((!n_n4767) & (x165x) & (!n_n4763) & (n_n3469) & (!x164x)) + ((!n_n4767) & (x165x) & (!n_n4763) & (n_n3469) & (x164x)) + ((!n_n4767) & (x165x) & (n_n4763) & (!n_n3469) & (!x164x)) + ((!n_n4767) & (x165x) & (n_n4763) & (!n_n3469) & (x164x)) + ((!n_n4767) & (x165x) & (n_n4763) & (n_n3469) & (!x164x)) + ((!n_n4767) & (x165x) & (n_n4763) & (n_n3469) & (x164x)) + ((n_n4767) & (!x165x) & (!n_n4763) & (!n_n3469) & (!x164x)) + ((n_n4767) & (!x165x) & (!n_n4763) & (!n_n3469) & (x164x)) + ((n_n4767) & (!x165x) & (!n_n4763) & (n_n3469) & (!x164x)) + ((n_n4767) & (!x165x) & (!n_n4763) & (n_n3469) & (x164x)) + ((n_n4767) & (!x165x) & (n_n4763) & (!n_n3469) & (!x164x)) + ((n_n4767) & (!x165x) & (n_n4763) & (!n_n3469) & (x164x)) + ((n_n4767) & (!x165x) & (n_n4763) & (n_n3469) & (!x164x)) + ((n_n4767) & (!x165x) & (n_n4763) & (n_n3469) & (x164x)) + ((n_n4767) & (x165x) & (!n_n4763) & (!n_n3469) & (!x164x)) + ((n_n4767) & (x165x) & (!n_n4763) & (!n_n3469) & (x164x)) + ((n_n4767) & (x165x) & (!n_n4763) & (n_n3469) & (!x164x)) + ((n_n4767) & (x165x) & (!n_n4763) & (n_n3469) & (x164x)) + ((n_n4767) & (x165x) & (n_n4763) & (!n_n3469) & (!x164x)) + ((n_n4767) & (x165x) & (n_n4763) & (!n_n3469) & (x164x)) + ((n_n4767) & (x165x) & (n_n4763) & (n_n3469) & (!x164x)) + ((n_n4767) & (x165x) & (n_n4763) & (n_n3469) & (x164x)));
	assign n_n4776 = (((i_9_) & (n_n482) & (n_n534) & (n_n325)));
	assign n_n4774 = (((i_9_) & (n_n325) & (n_n491) & (n_n520)));
	assign n_n4786 = (((i_9_) & (n_n524) & (n_n482) & (n_n325)));
	assign x131x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n482) & (n_n325)) + ((!i_9_) & (n_n524) & (!n_n526) & (n_n482) & (n_n325)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n482) & (n_n325)));
	assign n_n4789 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n325) & (x20x)));
	assign x313x = (((!i_9_) & (n_n482) & (n_n325) & (!n_n522) & (x20x)) + ((!i_9_) & (n_n482) & (n_n325) & (n_n522) & (x20x)) + ((i_9_) & (n_n482) & (n_n325) & (!n_n522) & (x20x)) + ((i_9_) & (n_n482) & (n_n325) & (n_n522) & (!x20x)) + ((i_9_) & (n_n482) & (n_n325) & (n_n522) & (x20x)));
	assign x16374x = (((!n_n4786) & (!x131x) & (!n_n4789) & (!n_n4788) & (!x22060x)) + ((!n_n4786) & (!x131x) & (!n_n4789) & (n_n4788) & (!x22060x)) + ((!n_n4786) & (!x131x) & (!n_n4789) & (n_n4788) & (x22060x)) + ((!n_n4786) & (!x131x) & (n_n4789) & (!n_n4788) & (!x22060x)) + ((!n_n4786) & (!x131x) & (n_n4789) & (!n_n4788) & (x22060x)) + ((!n_n4786) & (!x131x) & (n_n4789) & (n_n4788) & (!x22060x)) + ((!n_n4786) & (!x131x) & (n_n4789) & (n_n4788) & (x22060x)) + ((!n_n4786) & (x131x) & (!n_n4789) & (!n_n4788) & (!x22060x)) + ((!n_n4786) & (x131x) & (!n_n4789) & (!n_n4788) & (x22060x)) + ((!n_n4786) & (x131x) & (!n_n4789) & (n_n4788) & (!x22060x)) + ((!n_n4786) & (x131x) & (!n_n4789) & (n_n4788) & (x22060x)) + ((!n_n4786) & (x131x) & (n_n4789) & (!n_n4788) & (!x22060x)) + ((!n_n4786) & (x131x) & (n_n4789) & (!n_n4788) & (x22060x)) + ((!n_n4786) & (x131x) & (n_n4789) & (n_n4788) & (!x22060x)) + ((!n_n4786) & (x131x) & (n_n4789) & (n_n4788) & (x22060x)) + ((n_n4786) & (!x131x) & (!n_n4789) & (!n_n4788) & (!x22060x)) + ((n_n4786) & (!x131x) & (!n_n4789) & (!n_n4788) & (x22060x)) + ((n_n4786) & (!x131x) & (!n_n4789) & (n_n4788) & (!x22060x)) + ((n_n4786) & (!x131x) & (!n_n4789) & (n_n4788) & (x22060x)) + ((n_n4786) & (!x131x) & (n_n4789) & (!n_n4788) & (!x22060x)) + ((n_n4786) & (!x131x) & (n_n4789) & (!n_n4788) & (x22060x)) + ((n_n4786) & (!x131x) & (n_n4789) & (n_n4788) & (!x22060x)) + ((n_n4786) & (!x131x) & (n_n4789) & (n_n4788) & (x22060x)) + ((n_n4786) & (x131x) & (!n_n4789) & (!n_n4788) & (!x22060x)) + ((n_n4786) & (x131x) & (!n_n4789) & (!n_n4788) & (x22060x)) + ((n_n4786) & (x131x) & (!n_n4789) & (n_n4788) & (!x22060x)) + ((n_n4786) & (x131x) & (!n_n4789) & (n_n4788) & (x22060x)) + ((n_n4786) & (x131x) & (n_n4789) & (!n_n4788) & (!x22060x)) + ((n_n4786) & (x131x) & (n_n4789) & (!n_n4788) & (x22060x)) + ((n_n4786) & (x131x) & (n_n4789) & (n_n4788) & (!x22060x)) + ((n_n4786) & (x131x) & (n_n4789) & (n_n4788) & (x22060x)));
	assign x16376x = (((!x16349x) & (!x16350x) & (!n_n2234) & (x16374x)) + ((!x16349x) & (!x16350x) & (n_n2234) & (!x16374x)) + ((!x16349x) & (!x16350x) & (n_n2234) & (x16374x)) + ((!x16349x) & (x16350x) & (!n_n2234) & (!x16374x)) + ((!x16349x) & (x16350x) & (!n_n2234) & (x16374x)) + ((!x16349x) & (x16350x) & (n_n2234) & (!x16374x)) + ((!x16349x) & (x16350x) & (n_n2234) & (x16374x)) + ((x16349x) & (!x16350x) & (!n_n2234) & (!x16374x)) + ((x16349x) & (!x16350x) & (!n_n2234) & (x16374x)) + ((x16349x) & (!x16350x) & (n_n2234) & (!x16374x)) + ((x16349x) & (!x16350x) & (n_n2234) & (x16374x)) + ((x16349x) & (x16350x) & (!n_n2234) & (!x16374x)) + ((x16349x) & (x16350x) & (!n_n2234) & (x16374x)) + ((x16349x) & (x16350x) & (n_n2234) & (!x16374x)) + ((x16349x) & (x16350x) & (n_n2234) & (x16374x)));
	assign x16362x = (((!x23x) & (!x530x) & (!n_n4824) & (!n_n4822) & (n_n4806)) + ((!x23x) & (!x530x) & (!n_n4824) & (n_n4822) & (!n_n4806)) + ((!x23x) & (!x530x) & (!n_n4824) & (n_n4822) & (n_n4806)) + ((!x23x) & (!x530x) & (n_n4824) & (!n_n4822) & (!n_n4806)) + ((!x23x) & (!x530x) & (n_n4824) & (!n_n4822) & (n_n4806)) + ((!x23x) & (!x530x) & (n_n4824) & (n_n4822) & (!n_n4806)) + ((!x23x) & (!x530x) & (n_n4824) & (n_n4822) & (n_n4806)) + ((!x23x) & (x530x) & (!n_n4824) & (!n_n4822) & (n_n4806)) + ((!x23x) & (x530x) & (!n_n4824) & (n_n4822) & (!n_n4806)) + ((!x23x) & (x530x) & (!n_n4824) & (n_n4822) & (n_n4806)) + ((!x23x) & (x530x) & (n_n4824) & (!n_n4822) & (!n_n4806)) + ((!x23x) & (x530x) & (n_n4824) & (!n_n4822) & (n_n4806)) + ((!x23x) & (x530x) & (n_n4824) & (n_n4822) & (!n_n4806)) + ((!x23x) & (x530x) & (n_n4824) & (n_n4822) & (n_n4806)) + ((x23x) & (!x530x) & (!n_n4824) & (!n_n4822) & (n_n4806)) + ((x23x) & (!x530x) & (!n_n4824) & (n_n4822) & (!n_n4806)) + ((x23x) & (!x530x) & (!n_n4824) & (n_n4822) & (n_n4806)) + ((x23x) & (!x530x) & (n_n4824) & (!n_n4822) & (!n_n4806)) + ((x23x) & (!x530x) & (n_n4824) & (!n_n4822) & (n_n4806)) + ((x23x) & (!x530x) & (n_n4824) & (n_n4822) & (!n_n4806)) + ((x23x) & (!x530x) & (n_n4824) & (n_n4822) & (n_n4806)) + ((x23x) & (x530x) & (!n_n4824) & (!n_n4822) & (!n_n4806)) + ((x23x) & (x530x) & (!n_n4824) & (!n_n4822) & (n_n4806)) + ((x23x) & (x530x) & (!n_n4824) & (n_n4822) & (!n_n4806)) + ((x23x) & (x530x) & (!n_n4824) & (n_n4822) & (n_n4806)) + ((x23x) & (x530x) & (n_n4824) & (!n_n4822) & (!n_n4806)) + ((x23x) & (x530x) & (n_n4824) & (!n_n4822) & (n_n4806)) + ((x23x) & (x530x) & (n_n4824) & (n_n4822) & (!n_n4806)) + ((x23x) & (x530x) & (n_n4824) & (n_n4822) & (n_n4806)));
	assign x16363x = (((!n_n4821) & (!n_n4820) & (!n_n4818) & (!n_n4810) & (n_n4819)) + ((!n_n4821) & (!n_n4820) & (!n_n4818) & (n_n4810) & (!n_n4819)) + ((!n_n4821) & (!n_n4820) & (!n_n4818) & (n_n4810) & (n_n4819)) + ((!n_n4821) & (!n_n4820) & (n_n4818) & (!n_n4810) & (!n_n4819)) + ((!n_n4821) & (!n_n4820) & (n_n4818) & (!n_n4810) & (n_n4819)) + ((!n_n4821) & (!n_n4820) & (n_n4818) & (n_n4810) & (!n_n4819)) + ((!n_n4821) & (!n_n4820) & (n_n4818) & (n_n4810) & (n_n4819)) + ((!n_n4821) & (n_n4820) & (!n_n4818) & (!n_n4810) & (!n_n4819)) + ((!n_n4821) & (n_n4820) & (!n_n4818) & (!n_n4810) & (n_n4819)) + ((!n_n4821) & (n_n4820) & (!n_n4818) & (n_n4810) & (!n_n4819)) + ((!n_n4821) & (n_n4820) & (!n_n4818) & (n_n4810) & (n_n4819)) + ((!n_n4821) & (n_n4820) & (n_n4818) & (!n_n4810) & (!n_n4819)) + ((!n_n4821) & (n_n4820) & (n_n4818) & (!n_n4810) & (n_n4819)) + ((!n_n4821) & (n_n4820) & (n_n4818) & (n_n4810) & (!n_n4819)) + ((!n_n4821) & (n_n4820) & (n_n4818) & (n_n4810) & (n_n4819)) + ((n_n4821) & (!n_n4820) & (!n_n4818) & (!n_n4810) & (!n_n4819)) + ((n_n4821) & (!n_n4820) & (!n_n4818) & (!n_n4810) & (n_n4819)) + ((n_n4821) & (!n_n4820) & (!n_n4818) & (n_n4810) & (!n_n4819)) + ((n_n4821) & (!n_n4820) & (!n_n4818) & (n_n4810) & (n_n4819)) + ((n_n4821) & (!n_n4820) & (n_n4818) & (!n_n4810) & (!n_n4819)) + ((n_n4821) & (!n_n4820) & (n_n4818) & (!n_n4810) & (n_n4819)) + ((n_n4821) & (!n_n4820) & (n_n4818) & (n_n4810) & (!n_n4819)) + ((n_n4821) & (!n_n4820) & (n_n4818) & (n_n4810) & (n_n4819)) + ((n_n4821) & (n_n4820) & (!n_n4818) & (!n_n4810) & (!n_n4819)) + ((n_n4821) & (n_n4820) & (!n_n4818) & (!n_n4810) & (n_n4819)) + ((n_n4821) & (n_n4820) & (!n_n4818) & (n_n4810) & (!n_n4819)) + ((n_n4821) & (n_n4820) & (!n_n4818) & (n_n4810) & (n_n4819)) + ((n_n4821) & (n_n4820) & (n_n4818) & (!n_n4810) & (!n_n4819)) + ((n_n4821) & (n_n4820) & (n_n4818) & (!n_n4810) & (n_n4819)) + ((n_n4821) & (n_n4820) & (n_n4818) & (n_n4810) & (!n_n4819)) + ((n_n4821) & (n_n4820) & (n_n4818) & (n_n4810) & (n_n4819)));
	assign n_n4755 = (((!i_9_) & (n_n524) & (n_n325) & (n_n500)));
	assign n_n4743 = (((i_5_) & (i_3_) & (!i_4_) & (n_n325) & (x23x)));
	assign n_n4742 = (((i_9_) & (n_n509) & (n_n325) & (n_n520)));
	assign n_n4752 = (((i_9_) & (n_n526) & (n_n325) & (n_n500)));
	assign x16383x = (((!n_n4751) & (!n_n4750) & (!n_n4743) & (!n_n4742) & (n_n4752)) + ((!n_n4751) & (!n_n4750) & (!n_n4743) & (n_n4742) & (!n_n4752)) + ((!n_n4751) & (!n_n4750) & (!n_n4743) & (n_n4742) & (n_n4752)) + ((!n_n4751) & (!n_n4750) & (n_n4743) & (!n_n4742) & (!n_n4752)) + ((!n_n4751) & (!n_n4750) & (n_n4743) & (!n_n4742) & (n_n4752)) + ((!n_n4751) & (!n_n4750) & (n_n4743) & (n_n4742) & (!n_n4752)) + ((!n_n4751) & (!n_n4750) & (n_n4743) & (n_n4742) & (n_n4752)) + ((!n_n4751) & (n_n4750) & (!n_n4743) & (!n_n4742) & (!n_n4752)) + ((!n_n4751) & (n_n4750) & (!n_n4743) & (!n_n4742) & (n_n4752)) + ((!n_n4751) & (n_n4750) & (!n_n4743) & (n_n4742) & (!n_n4752)) + ((!n_n4751) & (n_n4750) & (!n_n4743) & (n_n4742) & (n_n4752)) + ((!n_n4751) & (n_n4750) & (n_n4743) & (!n_n4742) & (!n_n4752)) + ((!n_n4751) & (n_n4750) & (n_n4743) & (!n_n4742) & (n_n4752)) + ((!n_n4751) & (n_n4750) & (n_n4743) & (n_n4742) & (!n_n4752)) + ((!n_n4751) & (n_n4750) & (n_n4743) & (n_n4742) & (n_n4752)) + ((n_n4751) & (!n_n4750) & (!n_n4743) & (!n_n4742) & (!n_n4752)) + ((n_n4751) & (!n_n4750) & (!n_n4743) & (!n_n4742) & (n_n4752)) + ((n_n4751) & (!n_n4750) & (!n_n4743) & (n_n4742) & (!n_n4752)) + ((n_n4751) & (!n_n4750) & (!n_n4743) & (n_n4742) & (n_n4752)) + ((n_n4751) & (!n_n4750) & (n_n4743) & (!n_n4742) & (!n_n4752)) + ((n_n4751) & (!n_n4750) & (n_n4743) & (!n_n4742) & (n_n4752)) + ((n_n4751) & (!n_n4750) & (n_n4743) & (n_n4742) & (!n_n4752)) + ((n_n4751) & (!n_n4750) & (n_n4743) & (n_n4742) & (n_n4752)) + ((n_n4751) & (n_n4750) & (!n_n4743) & (!n_n4742) & (!n_n4752)) + ((n_n4751) & (n_n4750) & (!n_n4743) & (!n_n4742) & (n_n4752)) + ((n_n4751) & (n_n4750) & (!n_n4743) & (n_n4742) & (!n_n4752)) + ((n_n4751) & (n_n4750) & (!n_n4743) & (n_n4742) & (n_n4752)) + ((n_n4751) & (n_n4750) & (n_n4743) & (!n_n4742) & (!n_n4752)) + ((n_n4751) & (n_n4750) & (n_n4743) & (!n_n4742) & (n_n4752)) + ((n_n4751) & (n_n4750) & (n_n4743) & (n_n4742) & (!n_n4752)) + ((n_n4751) & (n_n4750) & (n_n4743) & (n_n4742) & (n_n4752)));
	assign n_n4753 = (((!i_9_) & (n_n526) & (n_n325) & (n_n500)));
	assign n_n2236 = (((!n_n4749) & (!n_n4748) & (!n_n4747) & (!x16383x) & (n_n4753)) + ((!n_n4749) & (!n_n4748) & (!n_n4747) & (x16383x) & (!n_n4753)) + ((!n_n4749) & (!n_n4748) & (!n_n4747) & (x16383x) & (n_n4753)) + ((!n_n4749) & (!n_n4748) & (n_n4747) & (!x16383x) & (!n_n4753)) + ((!n_n4749) & (!n_n4748) & (n_n4747) & (!x16383x) & (n_n4753)) + ((!n_n4749) & (!n_n4748) & (n_n4747) & (x16383x) & (!n_n4753)) + ((!n_n4749) & (!n_n4748) & (n_n4747) & (x16383x) & (n_n4753)) + ((!n_n4749) & (n_n4748) & (!n_n4747) & (!x16383x) & (!n_n4753)) + ((!n_n4749) & (n_n4748) & (!n_n4747) & (!x16383x) & (n_n4753)) + ((!n_n4749) & (n_n4748) & (!n_n4747) & (x16383x) & (!n_n4753)) + ((!n_n4749) & (n_n4748) & (!n_n4747) & (x16383x) & (n_n4753)) + ((!n_n4749) & (n_n4748) & (n_n4747) & (!x16383x) & (!n_n4753)) + ((!n_n4749) & (n_n4748) & (n_n4747) & (!x16383x) & (n_n4753)) + ((!n_n4749) & (n_n4748) & (n_n4747) & (x16383x) & (!n_n4753)) + ((!n_n4749) & (n_n4748) & (n_n4747) & (x16383x) & (n_n4753)) + ((n_n4749) & (!n_n4748) & (!n_n4747) & (!x16383x) & (!n_n4753)) + ((n_n4749) & (!n_n4748) & (!n_n4747) & (!x16383x) & (n_n4753)) + ((n_n4749) & (!n_n4748) & (!n_n4747) & (x16383x) & (!n_n4753)) + ((n_n4749) & (!n_n4748) & (!n_n4747) & (x16383x) & (n_n4753)) + ((n_n4749) & (!n_n4748) & (n_n4747) & (!x16383x) & (!n_n4753)) + ((n_n4749) & (!n_n4748) & (n_n4747) & (!x16383x) & (n_n4753)) + ((n_n4749) & (!n_n4748) & (n_n4747) & (x16383x) & (!n_n4753)) + ((n_n4749) & (!n_n4748) & (n_n4747) & (x16383x) & (n_n4753)) + ((n_n4749) & (n_n4748) & (!n_n4747) & (!x16383x) & (!n_n4753)) + ((n_n4749) & (n_n4748) & (!n_n4747) & (!x16383x) & (n_n4753)) + ((n_n4749) & (n_n4748) & (!n_n4747) & (x16383x) & (!n_n4753)) + ((n_n4749) & (n_n4748) & (!n_n4747) & (x16383x) & (n_n4753)) + ((n_n4749) & (n_n4748) & (n_n4747) & (!x16383x) & (!n_n4753)) + ((n_n4749) & (n_n4748) & (n_n4747) & (!x16383x) & (n_n4753)) + ((n_n4749) & (n_n4748) & (n_n4747) & (x16383x) & (!n_n4753)) + ((n_n4749) & (n_n4748) & (n_n4747) & (x16383x) & (n_n4753)));
	assign x293x = (((!i_9_) & (!i_7_) & (i_8_) & (!i_6_) & (x483x)) + ((!i_9_) & (i_7_) & (!i_8_) & (!i_6_) & (x483x)));
	assign n_n3475 = (((!i_9_) & (!n_n526) & (n_n528) & (n_n509) & (n_n325)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n509) & (n_n325)) + ((i_9_) & (!n_n526) & (n_n528) & (n_n509) & (n_n325)) + ((i_9_) & (n_n526) & (!n_n528) & (n_n509) & (n_n325)) + ((i_9_) & (n_n526) & (n_n528) & (n_n509) & (n_n325)));
	assign n_n2237 = (((!n_n4738) & (!n_n4733) & (!x73x) & (!x293x) & (n_n3475)) + ((!n_n4738) & (!n_n4733) & (!x73x) & (x293x) & (!n_n3475)) + ((!n_n4738) & (!n_n4733) & (!x73x) & (x293x) & (n_n3475)) + ((!n_n4738) & (!n_n4733) & (x73x) & (!x293x) & (!n_n3475)) + ((!n_n4738) & (!n_n4733) & (x73x) & (!x293x) & (n_n3475)) + ((!n_n4738) & (!n_n4733) & (x73x) & (x293x) & (!n_n3475)) + ((!n_n4738) & (!n_n4733) & (x73x) & (x293x) & (n_n3475)) + ((!n_n4738) & (n_n4733) & (!x73x) & (!x293x) & (!n_n3475)) + ((!n_n4738) & (n_n4733) & (!x73x) & (!x293x) & (n_n3475)) + ((!n_n4738) & (n_n4733) & (!x73x) & (x293x) & (!n_n3475)) + ((!n_n4738) & (n_n4733) & (!x73x) & (x293x) & (n_n3475)) + ((!n_n4738) & (n_n4733) & (x73x) & (!x293x) & (!n_n3475)) + ((!n_n4738) & (n_n4733) & (x73x) & (!x293x) & (n_n3475)) + ((!n_n4738) & (n_n4733) & (x73x) & (x293x) & (!n_n3475)) + ((!n_n4738) & (n_n4733) & (x73x) & (x293x) & (n_n3475)) + ((n_n4738) & (!n_n4733) & (!x73x) & (!x293x) & (!n_n3475)) + ((n_n4738) & (!n_n4733) & (!x73x) & (!x293x) & (n_n3475)) + ((n_n4738) & (!n_n4733) & (!x73x) & (x293x) & (!n_n3475)) + ((n_n4738) & (!n_n4733) & (!x73x) & (x293x) & (n_n3475)) + ((n_n4738) & (!n_n4733) & (x73x) & (!x293x) & (!n_n3475)) + ((n_n4738) & (!n_n4733) & (x73x) & (!x293x) & (n_n3475)) + ((n_n4738) & (!n_n4733) & (x73x) & (x293x) & (!n_n3475)) + ((n_n4738) & (!n_n4733) & (x73x) & (x293x) & (n_n3475)) + ((n_n4738) & (n_n4733) & (!x73x) & (!x293x) & (!n_n3475)) + ((n_n4738) & (n_n4733) & (!x73x) & (!x293x) & (n_n3475)) + ((n_n4738) & (n_n4733) & (!x73x) & (x293x) & (!n_n3475)) + ((n_n4738) & (n_n4733) & (!x73x) & (x293x) & (n_n3475)) + ((n_n4738) & (n_n4733) & (x73x) & (!x293x) & (!n_n3475)) + ((n_n4738) & (n_n4733) & (x73x) & (!x293x) & (n_n3475)) + ((n_n4738) & (n_n4733) & (x73x) & (x293x) & (!n_n3475)) + ((n_n4738) & (n_n4733) & (x73x) & (x293x) & (n_n3475)));
	assign n_n4759 = (((!i_1_) & (!i_2_) & (i_0_) & (x23x) & (n_n500)));
	assign n_n4760 = (((i_9_) & (n_n534) & (n_n325) & (n_n491)));
	assign n_n4758 = (((i_9_) & (n_n325) & (n_n520) & (n_n500)));
	assign n_n4707 = (((!i_9_) & (n_n524) & (n_n325) & (n_n535)));
	assign n_n4702 = (((i_9_) & (n_n528) & (n_n325) & (n_n535)));
	assign n_n2378 = (((!i_9_) & (!n_n526) & (n_n528) & (n_n325) & (n_n535)) + ((!i_9_) & (n_n526) & (!n_n528) & (n_n325) & (n_n535)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n325) & (n_n535)) + ((i_9_) & (n_n526) & (!n_n528) & (n_n325) & (n_n535)) + ((i_9_) & (n_n526) & (n_n528) & (n_n325) & (n_n535)));
	assign x22219x = (((!n_n4720) & (!x241x) & (!n_n4709) & (!n_n4698)));
	assign x16399x = (((!n_n4707) & (!n_n4702) & (!n_n2378) & (!x22219x)) + ((!n_n4707) & (!n_n4702) & (n_n2378) & (!x22219x)) + ((!n_n4707) & (!n_n4702) & (n_n2378) & (x22219x)) + ((!n_n4707) & (n_n4702) & (!n_n2378) & (!x22219x)) + ((!n_n4707) & (n_n4702) & (!n_n2378) & (x22219x)) + ((!n_n4707) & (n_n4702) & (n_n2378) & (!x22219x)) + ((!n_n4707) & (n_n4702) & (n_n2378) & (x22219x)) + ((n_n4707) & (!n_n4702) & (!n_n2378) & (!x22219x)) + ((n_n4707) & (!n_n4702) & (!n_n2378) & (x22219x)) + ((n_n4707) & (!n_n4702) & (n_n2378) & (!x22219x)) + ((n_n4707) & (!n_n4702) & (n_n2378) & (x22219x)) + ((n_n4707) & (n_n4702) & (!n_n2378) & (!x22219x)) + ((n_n4707) & (n_n4702) & (!n_n2378) & (x22219x)) + ((n_n4707) & (n_n4702) & (n_n2378) & (!x22219x)) + ((n_n4707) & (n_n4702) & (n_n2378) & (x22219x)));
	assign n_n4696 = (((i_9_) & (n_n534) & (n_n325) & (n_n535)));
	assign n_n4695 = (((!i_1_) & (i_2_) & (i_0_) & (x23x) & (n_n464)));
	assign x16395x = (((!n_n4711) & (!n_n4712) & (!n_n4701) & (n_n4700)) + ((!n_n4711) & (!n_n4712) & (n_n4701) & (!n_n4700)) + ((!n_n4711) & (!n_n4712) & (n_n4701) & (n_n4700)) + ((!n_n4711) & (n_n4712) & (!n_n4701) & (!n_n4700)) + ((!n_n4711) & (n_n4712) & (!n_n4701) & (n_n4700)) + ((!n_n4711) & (n_n4712) & (n_n4701) & (!n_n4700)) + ((!n_n4711) & (n_n4712) & (n_n4701) & (n_n4700)) + ((n_n4711) & (!n_n4712) & (!n_n4701) & (!n_n4700)) + ((n_n4711) & (!n_n4712) & (!n_n4701) & (n_n4700)) + ((n_n4711) & (!n_n4712) & (n_n4701) & (!n_n4700)) + ((n_n4711) & (!n_n4712) & (n_n4701) & (n_n4700)) + ((n_n4711) & (n_n4712) & (!n_n4701) & (!n_n4700)) + ((n_n4711) & (n_n4712) & (!n_n4701) & (n_n4700)) + ((n_n4711) & (n_n4712) & (n_n4701) & (!n_n4700)) + ((n_n4711) & (n_n4712) & (n_n4701) & (n_n4700)));
	assign x22176x = (((!x244x) & (!x39x) & (!n_n4715) & (!n_n4714) & (!x16390x)));
	assign n_n2182 = (((!x16399x) & (!n_n4696) & (!n_n4695) & (!x16395x) & (!x22176x)) + ((!x16399x) & (!n_n4696) & (!n_n4695) & (x16395x) & (!x22176x)) + ((!x16399x) & (!n_n4696) & (!n_n4695) & (x16395x) & (x22176x)) + ((!x16399x) & (!n_n4696) & (n_n4695) & (!x16395x) & (!x22176x)) + ((!x16399x) & (!n_n4696) & (n_n4695) & (!x16395x) & (x22176x)) + ((!x16399x) & (!n_n4696) & (n_n4695) & (x16395x) & (!x22176x)) + ((!x16399x) & (!n_n4696) & (n_n4695) & (x16395x) & (x22176x)) + ((!x16399x) & (n_n4696) & (!n_n4695) & (!x16395x) & (!x22176x)) + ((!x16399x) & (n_n4696) & (!n_n4695) & (!x16395x) & (x22176x)) + ((!x16399x) & (n_n4696) & (!n_n4695) & (x16395x) & (!x22176x)) + ((!x16399x) & (n_n4696) & (!n_n4695) & (x16395x) & (x22176x)) + ((!x16399x) & (n_n4696) & (n_n4695) & (!x16395x) & (!x22176x)) + ((!x16399x) & (n_n4696) & (n_n4695) & (!x16395x) & (x22176x)) + ((!x16399x) & (n_n4696) & (n_n4695) & (x16395x) & (!x22176x)) + ((!x16399x) & (n_n4696) & (n_n4695) & (x16395x) & (x22176x)) + ((x16399x) & (!n_n4696) & (!n_n4695) & (!x16395x) & (!x22176x)) + ((x16399x) & (!n_n4696) & (!n_n4695) & (!x16395x) & (x22176x)) + ((x16399x) & (!n_n4696) & (!n_n4695) & (x16395x) & (!x22176x)) + ((x16399x) & (!n_n4696) & (!n_n4695) & (x16395x) & (x22176x)) + ((x16399x) & (!n_n4696) & (n_n4695) & (!x16395x) & (!x22176x)) + ((x16399x) & (!n_n4696) & (n_n4695) & (!x16395x) & (x22176x)) + ((x16399x) & (!n_n4696) & (n_n4695) & (x16395x) & (!x22176x)) + ((x16399x) & (!n_n4696) & (n_n4695) & (x16395x) & (x22176x)) + ((x16399x) & (n_n4696) & (!n_n4695) & (!x16395x) & (!x22176x)) + ((x16399x) & (n_n4696) & (!n_n4695) & (!x16395x) & (x22176x)) + ((x16399x) & (n_n4696) & (!n_n4695) & (x16395x) & (!x22176x)) + ((x16399x) & (n_n4696) & (!n_n4695) & (x16395x) & (x22176x)) + ((x16399x) & (n_n4696) & (n_n4695) & (!x16395x) & (!x22176x)) + ((x16399x) & (n_n4696) & (n_n4695) & (!x16395x) & (x22176x)) + ((x16399x) & (n_n4696) & (n_n4695) & (x16395x) & (!x22176x)) + ((x16399x) & (n_n4696) & (n_n4695) & (x16395x) & (x22176x)));
	assign n_n1764 = (((!x10x) & (!n_n473) & (!n_n4667) & (!n_n534) & (n_n4663)) + ((!x10x) & (!n_n473) & (!n_n4667) & (n_n534) & (n_n4663)) + ((!x10x) & (!n_n473) & (n_n4667) & (!n_n534) & (!n_n4663)) + ((!x10x) & (!n_n473) & (n_n4667) & (!n_n534) & (n_n4663)) + ((!x10x) & (!n_n473) & (n_n4667) & (n_n534) & (!n_n4663)) + ((!x10x) & (!n_n473) & (n_n4667) & (n_n534) & (n_n4663)) + ((!x10x) & (n_n473) & (!n_n4667) & (!n_n534) & (n_n4663)) + ((!x10x) & (n_n473) & (!n_n4667) & (n_n534) & (n_n4663)) + ((!x10x) & (n_n473) & (n_n4667) & (!n_n534) & (!n_n4663)) + ((!x10x) & (n_n473) & (n_n4667) & (!n_n534) & (n_n4663)) + ((!x10x) & (n_n473) & (n_n4667) & (n_n534) & (!n_n4663)) + ((!x10x) & (n_n473) & (n_n4667) & (n_n534) & (n_n4663)) + ((x10x) & (!n_n473) & (!n_n4667) & (!n_n534) & (n_n4663)) + ((x10x) & (!n_n473) & (!n_n4667) & (n_n534) & (n_n4663)) + ((x10x) & (!n_n473) & (n_n4667) & (!n_n534) & (!n_n4663)) + ((x10x) & (!n_n473) & (n_n4667) & (!n_n534) & (n_n4663)) + ((x10x) & (!n_n473) & (n_n4667) & (n_n534) & (!n_n4663)) + ((x10x) & (!n_n473) & (n_n4667) & (n_n534) & (n_n4663)) + ((x10x) & (n_n473) & (!n_n4667) & (!n_n534) & (n_n4663)) + ((x10x) & (n_n473) & (!n_n4667) & (n_n534) & (!n_n4663)) + ((x10x) & (n_n473) & (!n_n4667) & (n_n534) & (n_n4663)) + ((x10x) & (n_n473) & (n_n4667) & (!n_n534) & (!n_n4663)) + ((x10x) & (n_n473) & (n_n4667) & (!n_n534) & (n_n4663)) + ((x10x) & (n_n473) & (n_n4667) & (n_n534) & (!n_n4663)) + ((x10x) & (n_n473) & (n_n4667) & (n_n534) & (n_n4663)));
	assign n_n4688 = (((i_9_) & (n_n526) & (n_n390) & (n_n464)));
	assign n_n3849 = (((!i_9_) & (!n_n524) & (n_n526) & (n_n390) & (n_n464)) + ((!i_9_) & (n_n524) & (!n_n526) & (n_n390) & (n_n464)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n390) & (n_n464)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n390) & (n_n464)) + ((i_9_) & (n_n524) & (n_n526) & (n_n390) & (n_n464)));
	assign n_n4686 = (((i_9_) & (n_n528) & (n_n390) & (n_n464)));
	assign n_n3848 = (((!i_9_) & (n_n390) & (n_n522) & (!n_n520) & (n_n464)) + ((!i_9_) & (n_n390) & (n_n522) & (n_n520) & (n_n464)) + ((i_9_) & (n_n390) & (!n_n522) & (n_n520) & (n_n464)) + ((i_9_) & (n_n390) & (n_n522) & (!n_n520) & (n_n464)) + ((i_9_) & (n_n390) & (n_n522) & (n_n520) & (n_n464)));
	assign x16415x = (((!n_n1764) & (!n_n4688) & (!n_n3849) & (!n_n4686) & (n_n3848)) + ((!n_n1764) & (!n_n4688) & (!n_n3849) & (n_n4686) & (!n_n3848)) + ((!n_n1764) & (!n_n4688) & (!n_n3849) & (n_n4686) & (n_n3848)) + ((!n_n1764) & (!n_n4688) & (n_n3849) & (!n_n4686) & (!n_n3848)) + ((!n_n1764) & (!n_n4688) & (n_n3849) & (!n_n4686) & (n_n3848)) + ((!n_n1764) & (!n_n4688) & (n_n3849) & (n_n4686) & (!n_n3848)) + ((!n_n1764) & (!n_n4688) & (n_n3849) & (n_n4686) & (n_n3848)) + ((!n_n1764) & (n_n4688) & (!n_n3849) & (!n_n4686) & (!n_n3848)) + ((!n_n1764) & (n_n4688) & (!n_n3849) & (!n_n4686) & (n_n3848)) + ((!n_n1764) & (n_n4688) & (!n_n3849) & (n_n4686) & (!n_n3848)) + ((!n_n1764) & (n_n4688) & (!n_n3849) & (n_n4686) & (n_n3848)) + ((!n_n1764) & (n_n4688) & (n_n3849) & (!n_n4686) & (!n_n3848)) + ((!n_n1764) & (n_n4688) & (n_n3849) & (!n_n4686) & (n_n3848)) + ((!n_n1764) & (n_n4688) & (n_n3849) & (n_n4686) & (!n_n3848)) + ((!n_n1764) & (n_n4688) & (n_n3849) & (n_n4686) & (n_n3848)) + ((n_n1764) & (!n_n4688) & (!n_n3849) & (!n_n4686) & (!n_n3848)) + ((n_n1764) & (!n_n4688) & (!n_n3849) & (!n_n4686) & (n_n3848)) + ((n_n1764) & (!n_n4688) & (!n_n3849) & (n_n4686) & (!n_n3848)) + ((n_n1764) & (!n_n4688) & (!n_n3849) & (n_n4686) & (n_n3848)) + ((n_n1764) & (!n_n4688) & (n_n3849) & (!n_n4686) & (!n_n3848)) + ((n_n1764) & (!n_n4688) & (n_n3849) & (!n_n4686) & (n_n3848)) + ((n_n1764) & (!n_n4688) & (n_n3849) & (n_n4686) & (!n_n3848)) + ((n_n1764) & (!n_n4688) & (n_n3849) & (n_n4686) & (n_n3848)) + ((n_n1764) & (n_n4688) & (!n_n3849) & (!n_n4686) & (!n_n3848)) + ((n_n1764) & (n_n4688) & (!n_n3849) & (!n_n4686) & (n_n3848)) + ((n_n1764) & (n_n4688) & (!n_n3849) & (n_n4686) & (!n_n3848)) + ((n_n1764) & (n_n4688) & (!n_n3849) & (n_n4686) & (n_n3848)) + ((n_n1764) & (n_n4688) & (n_n3849) & (!n_n4686) & (!n_n3848)) + ((n_n1764) & (n_n4688) & (n_n3849) & (!n_n4686) & (n_n3848)) + ((n_n1764) & (n_n4688) & (n_n3849) & (n_n4686) & (!n_n3848)) + ((n_n1764) & (n_n4688) & (n_n3849) & (n_n4686) & (n_n3848)));
	assign n_n2242 = (((!n_n4673) & (!n_n4676) & (!n_n4681) & (!n_n4679) & (x16406x)) + ((!n_n4673) & (!n_n4676) & (!n_n4681) & (n_n4679) & (!x16406x)) + ((!n_n4673) & (!n_n4676) & (!n_n4681) & (n_n4679) & (x16406x)) + ((!n_n4673) & (!n_n4676) & (n_n4681) & (!n_n4679) & (!x16406x)) + ((!n_n4673) & (!n_n4676) & (n_n4681) & (!n_n4679) & (x16406x)) + ((!n_n4673) & (!n_n4676) & (n_n4681) & (n_n4679) & (!x16406x)) + ((!n_n4673) & (!n_n4676) & (n_n4681) & (n_n4679) & (x16406x)) + ((!n_n4673) & (n_n4676) & (!n_n4681) & (!n_n4679) & (!x16406x)) + ((!n_n4673) & (n_n4676) & (!n_n4681) & (!n_n4679) & (x16406x)) + ((!n_n4673) & (n_n4676) & (!n_n4681) & (n_n4679) & (!x16406x)) + ((!n_n4673) & (n_n4676) & (!n_n4681) & (n_n4679) & (x16406x)) + ((!n_n4673) & (n_n4676) & (n_n4681) & (!n_n4679) & (!x16406x)) + ((!n_n4673) & (n_n4676) & (n_n4681) & (!n_n4679) & (x16406x)) + ((!n_n4673) & (n_n4676) & (n_n4681) & (n_n4679) & (!x16406x)) + ((!n_n4673) & (n_n4676) & (n_n4681) & (n_n4679) & (x16406x)) + ((n_n4673) & (!n_n4676) & (!n_n4681) & (!n_n4679) & (!x16406x)) + ((n_n4673) & (!n_n4676) & (!n_n4681) & (!n_n4679) & (x16406x)) + ((n_n4673) & (!n_n4676) & (!n_n4681) & (n_n4679) & (!x16406x)) + ((n_n4673) & (!n_n4676) & (!n_n4681) & (n_n4679) & (x16406x)) + ((n_n4673) & (!n_n4676) & (n_n4681) & (!n_n4679) & (!x16406x)) + ((n_n4673) & (!n_n4676) & (n_n4681) & (!n_n4679) & (x16406x)) + ((n_n4673) & (!n_n4676) & (n_n4681) & (n_n4679) & (!x16406x)) + ((n_n4673) & (!n_n4676) & (n_n4681) & (n_n4679) & (x16406x)) + ((n_n4673) & (n_n4676) & (!n_n4681) & (!n_n4679) & (!x16406x)) + ((n_n4673) & (n_n4676) & (!n_n4681) & (!n_n4679) & (x16406x)) + ((n_n4673) & (n_n4676) & (!n_n4681) & (n_n4679) & (!x16406x)) + ((n_n4673) & (n_n4676) & (!n_n4681) & (n_n4679) & (x16406x)) + ((n_n4673) & (n_n4676) & (n_n4681) & (!n_n4679) & (!x16406x)) + ((n_n4673) & (n_n4676) & (n_n4681) & (!n_n4679) & (x16406x)) + ((n_n4673) & (n_n4676) & (n_n4681) & (n_n4679) & (!x16406x)) + ((n_n4673) & (n_n4676) & (n_n4681) & (n_n4679) & (x16406x)));
	assign x16414x = (((!n_n4662) & (!n_n4683) & (!n_n4657) & (!x431x) & (x16408x)) + ((!n_n4662) & (!n_n4683) & (!n_n4657) & (x431x) & (!x16408x)) + ((!n_n4662) & (!n_n4683) & (!n_n4657) & (x431x) & (x16408x)) + ((!n_n4662) & (!n_n4683) & (n_n4657) & (!x431x) & (!x16408x)) + ((!n_n4662) & (!n_n4683) & (n_n4657) & (!x431x) & (x16408x)) + ((!n_n4662) & (!n_n4683) & (n_n4657) & (x431x) & (!x16408x)) + ((!n_n4662) & (!n_n4683) & (n_n4657) & (x431x) & (x16408x)) + ((!n_n4662) & (n_n4683) & (!n_n4657) & (!x431x) & (!x16408x)) + ((!n_n4662) & (n_n4683) & (!n_n4657) & (!x431x) & (x16408x)) + ((!n_n4662) & (n_n4683) & (!n_n4657) & (x431x) & (!x16408x)) + ((!n_n4662) & (n_n4683) & (!n_n4657) & (x431x) & (x16408x)) + ((!n_n4662) & (n_n4683) & (n_n4657) & (!x431x) & (!x16408x)) + ((!n_n4662) & (n_n4683) & (n_n4657) & (!x431x) & (x16408x)) + ((!n_n4662) & (n_n4683) & (n_n4657) & (x431x) & (!x16408x)) + ((!n_n4662) & (n_n4683) & (n_n4657) & (x431x) & (x16408x)) + ((n_n4662) & (!n_n4683) & (!n_n4657) & (!x431x) & (!x16408x)) + ((n_n4662) & (!n_n4683) & (!n_n4657) & (!x431x) & (x16408x)) + ((n_n4662) & (!n_n4683) & (!n_n4657) & (x431x) & (!x16408x)) + ((n_n4662) & (!n_n4683) & (!n_n4657) & (x431x) & (x16408x)) + ((n_n4662) & (!n_n4683) & (n_n4657) & (!x431x) & (!x16408x)) + ((n_n4662) & (!n_n4683) & (n_n4657) & (!x431x) & (x16408x)) + ((n_n4662) & (!n_n4683) & (n_n4657) & (x431x) & (!x16408x)) + ((n_n4662) & (!n_n4683) & (n_n4657) & (x431x) & (x16408x)) + ((n_n4662) & (n_n4683) & (!n_n4657) & (!x431x) & (!x16408x)) + ((n_n4662) & (n_n4683) & (!n_n4657) & (!x431x) & (x16408x)) + ((n_n4662) & (n_n4683) & (!n_n4657) & (x431x) & (!x16408x)) + ((n_n4662) & (n_n4683) & (!n_n4657) & (x431x) & (x16408x)) + ((n_n4662) & (n_n4683) & (n_n4657) & (!x431x) & (!x16408x)) + ((n_n4662) & (n_n4683) & (n_n4657) & (!x431x) & (x16408x)) + ((n_n4662) & (n_n4683) & (n_n4657) & (x431x) & (!x16408x)) + ((n_n4662) & (n_n4683) & (n_n4657) & (x431x) & (x16408x)));
	assign n_n2183 = (((!x16415x) & (!n_n2242) & (x16414x)) + ((!x16415x) & (n_n2242) & (!x16414x)) + ((!x16415x) & (n_n2242) & (x16414x)) + ((x16415x) & (!n_n2242) & (!x16414x)) + ((x16415x) & (!n_n2242) & (x16414x)) + ((x16415x) & (n_n2242) & (!x16414x)) + ((x16415x) & (n_n2242) & (x16414x)));
	assign n_n4761 = (((!i_9_) & (n_n534) & (n_n325) & (n_n491)));
	assign n_n4762 = (((i_9_) & (n_n532) & (n_n325) & (n_n491)));
	assign x69x = (((!i_9_) & (!n_n532) & (n_n534) & (n_n325) & (n_n491)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n325) & (n_n491)) + ((i_9_) & (n_n532) & (!n_n534) & (n_n325) & (n_n491)) + ((i_9_) & (n_n532) & (n_n534) & (n_n325) & (n_n491)));
	assign x16423x = (((!n_n4759) & (!n_n4760) & (!n_n4758) & (!x69x) & (x16421x)) + ((!n_n4759) & (!n_n4760) & (!n_n4758) & (x69x) & (!x16421x)) + ((!n_n4759) & (!n_n4760) & (!n_n4758) & (x69x) & (x16421x)) + ((!n_n4759) & (!n_n4760) & (n_n4758) & (!x69x) & (!x16421x)) + ((!n_n4759) & (!n_n4760) & (n_n4758) & (!x69x) & (x16421x)) + ((!n_n4759) & (!n_n4760) & (n_n4758) & (x69x) & (!x16421x)) + ((!n_n4759) & (!n_n4760) & (n_n4758) & (x69x) & (x16421x)) + ((!n_n4759) & (n_n4760) & (!n_n4758) & (!x69x) & (!x16421x)) + ((!n_n4759) & (n_n4760) & (!n_n4758) & (!x69x) & (x16421x)) + ((!n_n4759) & (n_n4760) & (!n_n4758) & (x69x) & (!x16421x)) + ((!n_n4759) & (n_n4760) & (!n_n4758) & (x69x) & (x16421x)) + ((!n_n4759) & (n_n4760) & (n_n4758) & (!x69x) & (!x16421x)) + ((!n_n4759) & (n_n4760) & (n_n4758) & (!x69x) & (x16421x)) + ((!n_n4759) & (n_n4760) & (n_n4758) & (x69x) & (!x16421x)) + ((!n_n4759) & (n_n4760) & (n_n4758) & (x69x) & (x16421x)) + ((n_n4759) & (!n_n4760) & (!n_n4758) & (!x69x) & (!x16421x)) + ((n_n4759) & (!n_n4760) & (!n_n4758) & (!x69x) & (x16421x)) + ((n_n4759) & (!n_n4760) & (!n_n4758) & (x69x) & (!x16421x)) + ((n_n4759) & (!n_n4760) & (!n_n4758) & (x69x) & (x16421x)) + ((n_n4759) & (!n_n4760) & (n_n4758) & (!x69x) & (!x16421x)) + ((n_n4759) & (!n_n4760) & (n_n4758) & (!x69x) & (x16421x)) + ((n_n4759) & (!n_n4760) & (n_n4758) & (x69x) & (!x16421x)) + ((n_n4759) & (!n_n4760) & (n_n4758) & (x69x) & (x16421x)) + ((n_n4759) & (n_n4760) & (!n_n4758) & (!x69x) & (!x16421x)) + ((n_n4759) & (n_n4760) & (!n_n4758) & (!x69x) & (x16421x)) + ((n_n4759) & (n_n4760) & (!n_n4758) & (x69x) & (!x16421x)) + ((n_n4759) & (n_n4760) & (!n_n4758) & (x69x) & (x16421x)) + ((n_n4759) & (n_n4760) & (n_n4758) & (!x69x) & (!x16421x)) + ((n_n4759) & (n_n4760) & (n_n4758) & (!x69x) & (x16421x)) + ((n_n4759) & (n_n4760) & (n_n4758) & (x69x) & (!x16421x)) + ((n_n4759) & (n_n4760) & (n_n4758) & (x69x) & (x16421x)));
	assign n_n4963 = (((!i_9_) & (n_n524) & (n_n535) & (n_n195)));
	assign n_n4959 = (((!i_9_) & (n_n528) & (n_n535) & (n_n195)));
	assign n_n4960 = (((i_9_) & (n_n526) & (n_n535) & (n_n195)));
	assign n_n4964 = (((i_9_) & (n_n535) & (n_n522) & (n_n195)));
	assign n_n2218 = (((!n_n5001) & (!n_n5006) & (!n_n5007) & (!x393x) & (!x22065x)) + ((!n_n5001) & (!n_n5006) & (!n_n5007) & (x393x) & (!x22065x)) + ((!n_n5001) & (!n_n5006) & (!n_n5007) & (x393x) & (x22065x)) + ((!n_n5001) & (!n_n5006) & (n_n5007) & (!x393x) & (!x22065x)) + ((!n_n5001) & (!n_n5006) & (n_n5007) & (!x393x) & (x22065x)) + ((!n_n5001) & (!n_n5006) & (n_n5007) & (x393x) & (!x22065x)) + ((!n_n5001) & (!n_n5006) & (n_n5007) & (x393x) & (x22065x)) + ((!n_n5001) & (n_n5006) & (!n_n5007) & (!x393x) & (!x22065x)) + ((!n_n5001) & (n_n5006) & (!n_n5007) & (!x393x) & (x22065x)) + ((!n_n5001) & (n_n5006) & (!n_n5007) & (x393x) & (!x22065x)) + ((!n_n5001) & (n_n5006) & (!n_n5007) & (x393x) & (x22065x)) + ((!n_n5001) & (n_n5006) & (n_n5007) & (!x393x) & (!x22065x)) + ((!n_n5001) & (n_n5006) & (n_n5007) & (!x393x) & (x22065x)) + ((!n_n5001) & (n_n5006) & (n_n5007) & (x393x) & (!x22065x)) + ((!n_n5001) & (n_n5006) & (n_n5007) & (x393x) & (x22065x)) + ((n_n5001) & (!n_n5006) & (!n_n5007) & (!x393x) & (!x22065x)) + ((n_n5001) & (!n_n5006) & (!n_n5007) & (!x393x) & (x22065x)) + ((n_n5001) & (!n_n5006) & (!n_n5007) & (x393x) & (!x22065x)) + ((n_n5001) & (!n_n5006) & (!n_n5007) & (x393x) & (x22065x)) + ((n_n5001) & (!n_n5006) & (n_n5007) & (!x393x) & (!x22065x)) + ((n_n5001) & (!n_n5006) & (n_n5007) & (!x393x) & (x22065x)) + ((n_n5001) & (!n_n5006) & (n_n5007) & (x393x) & (!x22065x)) + ((n_n5001) & (!n_n5006) & (n_n5007) & (x393x) & (x22065x)) + ((n_n5001) & (n_n5006) & (!n_n5007) & (!x393x) & (!x22065x)) + ((n_n5001) & (n_n5006) & (!n_n5007) & (!x393x) & (x22065x)) + ((n_n5001) & (n_n5006) & (!n_n5007) & (x393x) & (!x22065x)) + ((n_n5001) & (n_n5006) & (!n_n5007) & (x393x) & (x22065x)) + ((n_n5001) & (n_n5006) & (n_n5007) & (!x393x) & (!x22065x)) + ((n_n5001) & (n_n5006) & (n_n5007) & (!x393x) & (x22065x)) + ((n_n5001) & (n_n5006) & (n_n5007) & (x393x) & (!x22065x)) + ((n_n5001) & (n_n5006) & (n_n5007) & (x393x) & (x22065x)));
	assign x16435x = (((!n_n5018) & (!n_n5015) & (!n_n5010) & (n_n5012)) + ((!n_n5018) & (!n_n5015) & (n_n5010) & (!n_n5012)) + ((!n_n5018) & (!n_n5015) & (n_n5010) & (n_n5012)) + ((!n_n5018) & (n_n5015) & (!n_n5010) & (!n_n5012)) + ((!n_n5018) & (n_n5015) & (!n_n5010) & (n_n5012)) + ((!n_n5018) & (n_n5015) & (n_n5010) & (!n_n5012)) + ((!n_n5018) & (n_n5015) & (n_n5010) & (n_n5012)) + ((n_n5018) & (!n_n5015) & (!n_n5010) & (!n_n5012)) + ((n_n5018) & (!n_n5015) & (!n_n5010) & (n_n5012)) + ((n_n5018) & (!n_n5015) & (n_n5010) & (!n_n5012)) + ((n_n5018) & (!n_n5015) & (n_n5010) & (n_n5012)) + ((n_n5018) & (n_n5015) & (!n_n5010) & (!n_n5012)) + ((n_n5018) & (n_n5015) & (!n_n5010) & (n_n5012)) + ((n_n5018) & (n_n5015) & (n_n5010) & (!n_n5012)) + ((n_n5018) & (n_n5015) & (n_n5010) & (n_n5012)));
	assign x16436x = (((!n_n5017) & (!n_n5021) & (!n_n5016) & (!n_n5009) & (n_n5013)) + ((!n_n5017) & (!n_n5021) & (!n_n5016) & (n_n5009) & (!n_n5013)) + ((!n_n5017) & (!n_n5021) & (!n_n5016) & (n_n5009) & (n_n5013)) + ((!n_n5017) & (!n_n5021) & (n_n5016) & (!n_n5009) & (!n_n5013)) + ((!n_n5017) & (!n_n5021) & (n_n5016) & (!n_n5009) & (n_n5013)) + ((!n_n5017) & (!n_n5021) & (n_n5016) & (n_n5009) & (!n_n5013)) + ((!n_n5017) & (!n_n5021) & (n_n5016) & (n_n5009) & (n_n5013)) + ((!n_n5017) & (n_n5021) & (!n_n5016) & (!n_n5009) & (!n_n5013)) + ((!n_n5017) & (n_n5021) & (!n_n5016) & (!n_n5009) & (n_n5013)) + ((!n_n5017) & (n_n5021) & (!n_n5016) & (n_n5009) & (!n_n5013)) + ((!n_n5017) & (n_n5021) & (!n_n5016) & (n_n5009) & (n_n5013)) + ((!n_n5017) & (n_n5021) & (n_n5016) & (!n_n5009) & (!n_n5013)) + ((!n_n5017) & (n_n5021) & (n_n5016) & (!n_n5009) & (n_n5013)) + ((!n_n5017) & (n_n5021) & (n_n5016) & (n_n5009) & (!n_n5013)) + ((!n_n5017) & (n_n5021) & (n_n5016) & (n_n5009) & (n_n5013)) + ((n_n5017) & (!n_n5021) & (!n_n5016) & (!n_n5009) & (!n_n5013)) + ((n_n5017) & (!n_n5021) & (!n_n5016) & (!n_n5009) & (n_n5013)) + ((n_n5017) & (!n_n5021) & (!n_n5016) & (n_n5009) & (!n_n5013)) + ((n_n5017) & (!n_n5021) & (!n_n5016) & (n_n5009) & (n_n5013)) + ((n_n5017) & (!n_n5021) & (n_n5016) & (!n_n5009) & (!n_n5013)) + ((n_n5017) & (!n_n5021) & (n_n5016) & (!n_n5009) & (n_n5013)) + ((n_n5017) & (!n_n5021) & (n_n5016) & (n_n5009) & (!n_n5013)) + ((n_n5017) & (!n_n5021) & (n_n5016) & (n_n5009) & (n_n5013)) + ((n_n5017) & (n_n5021) & (!n_n5016) & (!n_n5009) & (!n_n5013)) + ((n_n5017) & (n_n5021) & (!n_n5016) & (!n_n5009) & (n_n5013)) + ((n_n5017) & (n_n5021) & (!n_n5016) & (n_n5009) & (!n_n5013)) + ((n_n5017) & (n_n5021) & (!n_n5016) & (n_n5009) & (n_n5013)) + ((n_n5017) & (n_n5021) & (n_n5016) & (!n_n5009) & (!n_n5013)) + ((n_n5017) & (n_n5021) & (n_n5016) & (!n_n5009) & (n_n5013)) + ((n_n5017) & (n_n5021) & (n_n5016) & (n_n5009) & (!n_n5013)) + ((n_n5017) & (n_n5021) & (n_n5016) & (n_n5009) & (n_n5013)));
	assign x16440x = (((!n_n4990) & (!n_n4988) & (!n_n4987) & (n_n4979)) + ((!n_n4990) & (!n_n4988) & (n_n4987) & (!n_n4979)) + ((!n_n4990) & (!n_n4988) & (n_n4987) & (n_n4979)) + ((!n_n4990) & (n_n4988) & (!n_n4987) & (!n_n4979)) + ((!n_n4990) & (n_n4988) & (!n_n4987) & (n_n4979)) + ((!n_n4990) & (n_n4988) & (n_n4987) & (!n_n4979)) + ((!n_n4990) & (n_n4988) & (n_n4987) & (n_n4979)) + ((n_n4990) & (!n_n4988) & (!n_n4987) & (!n_n4979)) + ((n_n4990) & (!n_n4988) & (!n_n4987) & (n_n4979)) + ((n_n4990) & (!n_n4988) & (n_n4987) & (!n_n4979)) + ((n_n4990) & (!n_n4988) & (n_n4987) & (n_n4979)) + ((n_n4990) & (n_n4988) & (!n_n4987) & (!n_n4979)) + ((n_n4990) & (n_n4988) & (!n_n4987) & (n_n4979)) + ((n_n4990) & (n_n4988) & (n_n4987) & (!n_n4979)) + ((n_n4990) & (n_n4988) & (n_n4987) & (n_n4979)));
	assign x16441x = (((!n_n4982) & (!n_n4983) & (!n_n4985) & (!n_n4984) & (n_n4986)) + ((!n_n4982) & (!n_n4983) & (!n_n4985) & (n_n4984) & (!n_n4986)) + ((!n_n4982) & (!n_n4983) & (!n_n4985) & (n_n4984) & (n_n4986)) + ((!n_n4982) & (!n_n4983) & (n_n4985) & (!n_n4984) & (!n_n4986)) + ((!n_n4982) & (!n_n4983) & (n_n4985) & (!n_n4984) & (n_n4986)) + ((!n_n4982) & (!n_n4983) & (n_n4985) & (n_n4984) & (!n_n4986)) + ((!n_n4982) & (!n_n4983) & (n_n4985) & (n_n4984) & (n_n4986)) + ((!n_n4982) & (n_n4983) & (!n_n4985) & (!n_n4984) & (!n_n4986)) + ((!n_n4982) & (n_n4983) & (!n_n4985) & (!n_n4984) & (n_n4986)) + ((!n_n4982) & (n_n4983) & (!n_n4985) & (n_n4984) & (!n_n4986)) + ((!n_n4982) & (n_n4983) & (!n_n4985) & (n_n4984) & (n_n4986)) + ((!n_n4982) & (n_n4983) & (n_n4985) & (!n_n4984) & (!n_n4986)) + ((!n_n4982) & (n_n4983) & (n_n4985) & (!n_n4984) & (n_n4986)) + ((!n_n4982) & (n_n4983) & (n_n4985) & (n_n4984) & (!n_n4986)) + ((!n_n4982) & (n_n4983) & (n_n4985) & (n_n4984) & (n_n4986)) + ((n_n4982) & (!n_n4983) & (!n_n4985) & (!n_n4984) & (!n_n4986)) + ((n_n4982) & (!n_n4983) & (!n_n4985) & (!n_n4984) & (n_n4986)) + ((n_n4982) & (!n_n4983) & (!n_n4985) & (n_n4984) & (!n_n4986)) + ((n_n4982) & (!n_n4983) & (!n_n4985) & (n_n4984) & (n_n4986)) + ((n_n4982) & (!n_n4983) & (n_n4985) & (!n_n4984) & (!n_n4986)) + ((n_n4982) & (!n_n4983) & (n_n4985) & (!n_n4984) & (n_n4986)) + ((n_n4982) & (!n_n4983) & (n_n4985) & (n_n4984) & (!n_n4986)) + ((n_n4982) & (!n_n4983) & (n_n4985) & (n_n4984) & (n_n4986)) + ((n_n4982) & (n_n4983) & (!n_n4985) & (!n_n4984) & (!n_n4986)) + ((n_n4982) & (n_n4983) & (!n_n4985) & (!n_n4984) & (n_n4986)) + ((n_n4982) & (n_n4983) & (!n_n4985) & (n_n4984) & (!n_n4986)) + ((n_n4982) & (n_n4983) & (!n_n4985) & (n_n4984) & (n_n4986)) + ((n_n4982) & (n_n4983) & (n_n4985) & (!n_n4984) & (!n_n4986)) + ((n_n4982) & (n_n4983) & (n_n4985) & (!n_n4984) & (n_n4986)) + ((n_n4982) & (n_n4983) & (n_n4985) & (n_n4984) & (!n_n4986)) + ((n_n4982) & (n_n4983) & (n_n4985) & (n_n4984) & (n_n4986)));
	assign x351x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n482) & (n_n260)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n482) & (n_n260)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n482) & (n_n260)) + ((i_9_) & (n_n524) & (n_n526) & (n_n482) & (n_n260)));
	assign n_n4918 = (((i_9_) & (n_n482) & (n_n260) & (n_n520)));
	assign n_n4917 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n260) & (x20x)));
	assign n_n4915 = (((!i_9_) & (n_n524) & (n_n482) & (n_n260)));
	assign x22064x = (((!n_n4920) & (!n_n4923) & (!n_n4921) & (!n_n4919)));
	assign x228x = (((!i_9_) & (n_n518) & (n_n526) & (n_n195)) + ((i_9_) & (n_n518) & (n_n526) & (n_n195)));
	assign n_n4972 = (((i_9_) & (n_n518) & (n_n195) & (n_n530)));
	assign x341x = (((!i_9_) & (n_n518) & (n_n534) & (n_n195)) + ((i_9_) & (n_n518) & (n_n534) & (n_n195)));
	assign x362x = (((n_n535) & (n_n195) & (!x20x) & (x23x)) + ((n_n535) & (n_n195) & (x20x) & (!x23x)) + ((n_n535) & (n_n195) & (x20x) & (x23x)));
	assign x16458x = (((!i_9_) & (!n_n535) & (!n_n520) & (!n_n195) & (n_n4978)) + ((!i_9_) & (!n_n535) & (!n_n520) & (n_n195) & (n_n4978)) + ((!i_9_) & (!n_n535) & (n_n520) & (!n_n195) & (n_n4978)) + ((!i_9_) & (!n_n535) & (n_n520) & (n_n195) & (n_n4978)) + ((!i_9_) & (n_n535) & (!n_n520) & (!n_n195) & (n_n4978)) + ((!i_9_) & (n_n535) & (!n_n520) & (n_n195) & (n_n4978)) + ((!i_9_) & (n_n535) & (n_n520) & (!n_n195) & (n_n4978)) + ((!i_9_) & (n_n535) & (n_n520) & (n_n195) & (n_n4978)) + ((i_9_) & (!n_n535) & (!n_n520) & (!n_n195) & (n_n4978)) + ((i_9_) & (!n_n535) & (!n_n520) & (n_n195) & (n_n4978)) + ((i_9_) & (!n_n535) & (n_n520) & (!n_n195) & (n_n4978)) + ((i_9_) & (!n_n535) & (n_n520) & (n_n195) & (n_n4978)) + ((i_9_) & (n_n535) & (!n_n520) & (!n_n195) & (n_n4978)) + ((i_9_) & (n_n535) & (!n_n520) & (n_n195) & (n_n4978)) + ((i_9_) & (n_n535) & (n_n520) & (!n_n195) & (n_n4978)) + ((i_9_) & (n_n535) & (n_n520) & (n_n195) & (!n_n4978)) + ((i_9_) & (n_n535) & (n_n520) & (n_n195) & (n_n4978)));
	assign n_n2220 = (((!x228x) & (!n_n4972) & (!x341x) & (!x362x) & (x16458x)) + ((!x228x) & (!n_n4972) & (!x341x) & (x362x) & (!x16458x)) + ((!x228x) & (!n_n4972) & (!x341x) & (x362x) & (x16458x)) + ((!x228x) & (!n_n4972) & (x341x) & (!x362x) & (!x16458x)) + ((!x228x) & (!n_n4972) & (x341x) & (!x362x) & (x16458x)) + ((!x228x) & (!n_n4972) & (x341x) & (x362x) & (!x16458x)) + ((!x228x) & (!n_n4972) & (x341x) & (x362x) & (x16458x)) + ((!x228x) & (n_n4972) & (!x341x) & (!x362x) & (!x16458x)) + ((!x228x) & (n_n4972) & (!x341x) & (!x362x) & (x16458x)) + ((!x228x) & (n_n4972) & (!x341x) & (x362x) & (!x16458x)) + ((!x228x) & (n_n4972) & (!x341x) & (x362x) & (x16458x)) + ((!x228x) & (n_n4972) & (x341x) & (!x362x) & (!x16458x)) + ((!x228x) & (n_n4972) & (x341x) & (!x362x) & (x16458x)) + ((!x228x) & (n_n4972) & (x341x) & (x362x) & (!x16458x)) + ((!x228x) & (n_n4972) & (x341x) & (x362x) & (x16458x)) + ((x228x) & (!n_n4972) & (!x341x) & (!x362x) & (!x16458x)) + ((x228x) & (!n_n4972) & (!x341x) & (!x362x) & (x16458x)) + ((x228x) & (!n_n4972) & (!x341x) & (x362x) & (!x16458x)) + ((x228x) & (!n_n4972) & (!x341x) & (x362x) & (x16458x)) + ((x228x) & (!n_n4972) & (x341x) & (!x362x) & (!x16458x)) + ((x228x) & (!n_n4972) & (x341x) & (!x362x) & (x16458x)) + ((x228x) & (!n_n4972) & (x341x) & (x362x) & (!x16458x)) + ((x228x) & (!n_n4972) & (x341x) & (x362x) & (x16458x)) + ((x228x) & (n_n4972) & (!x341x) & (!x362x) & (!x16458x)) + ((x228x) & (n_n4972) & (!x341x) & (!x362x) & (x16458x)) + ((x228x) & (n_n4972) & (!x341x) & (x362x) & (!x16458x)) + ((x228x) & (n_n4972) & (!x341x) & (x362x) & (x16458x)) + ((x228x) & (n_n4972) & (x341x) & (!x362x) & (!x16458x)) + ((x228x) & (n_n4972) & (x341x) & (!x362x) & (x16458x)) + ((x228x) & (n_n4972) & (x341x) & (x362x) & (!x16458x)) + ((x228x) & (n_n4972) & (x341x) & (x362x) & (x16458x)));
	assign n_n4953 = (((!i_9_) & (n_n534) & (n_n535) & (n_n195)));
	assign n_n3802 = (((!i_9_) & (!n_n532) & (n_n534) & (n_n535) & (n_n195)) + ((!i_9_) & (n_n532) & (!n_n534) & (n_n535) & (n_n195)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n535) & (n_n195)) + ((i_9_) & (n_n532) & (!n_n534) & (n_n535) & (n_n195)) + ((i_9_) & (n_n532) & (n_n534) & (n_n535) & (n_n195)));
	assign n_n4956 = (((i_9_) & (n_n535) & (n_n195) & (n_n530)));
	assign x250x = (((!i_7_) & (!i_8_) & (i_6_) & (n_n535) & (x18x)) + ((!i_7_) & (i_8_) & (i_6_) & (n_n535) & (x18x)));
	assign n_n4817 = (((!i_9_) & (n_n526) & (n_n325) & (n_n464)));
	assign n_n4827 = (((!i_9_) & (n_n532) & (n_n260) & (n_n535)));
	assign n_n4816 = (((i_9_) & (n_n526) & (n_n325) & (n_n464)));
	assign n_n5097 = (((!i_9_) & (n_n518) & (n_n534) & (n_n130)));
	assign n_n4523 = (((!i_9_) & (n_n482) & (n_n455) & (n_n532)));
	assign n_n4547 = (((!i_9_) & (n_n524) & (n_n455) & (n_n473)));
	assign n_n4474 = (((i_9_) & (n_n455) & (n_n532) & (n_n509)));
	assign n_n4486 = (((i_9_) & (n_n455) & (n_n509) & (n_n520)));
	assign x199x = (((!i_9_) & (!n_n526) & (n_n455) & (n_n528) & (n_n509)) + ((!i_9_) & (n_n526) & (n_n455) & (!n_n528) & (n_n509)) + ((!i_9_) & (n_n526) & (n_n455) & (n_n528) & (n_n509)));
	assign x16483x = (((!n_n4474) & (!n_n4486) & (!n_n4484) & (x199x)) + ((!n_n4474) & (!n_n4486) & (n_n4484) & (!x199x)) + ((!n_n4474) & (!n_n4486) & (n_n4484) & (x199x)) + ((!n_n4474) & (n_n4486) & (!n_n4484) & (!x199x)) + ((!n_n4474) & (n_n4486) & (!n_n4484) & (x199x)) + ((!n_n4474) & (n_n4486) & (n_n4484) & (!x199x)) + ((!n_n4474) & (n_n4486) & (n_n4484) & (x199x)) + ((n_n4474) & (!n_n4486) & (!n_n4484) & (!x199x)) + ((n_n4474) & (!n_n4486) & (!n_n4484) & (x199x)) + ((n_n4474) & (!n_n4486) & (n_n4484) & (!x199x)) + ((n_n4474) & (!n_n4486) & (n_n4484) & (x199x)) + ((n_n4474) & (n_n4486) & (!n_n4484) & (!x199x)) + ((n_n4474) & (n_n4486) & (!n_n4484) & (x199x)) + ((n_n4474) & (n_n4486) & (n_n4484) & (!x199x)) + ((n_n4474) & (n_n4486) & (n_n4484) & (x199x)));
	assign n_n4518 = (((i_9_) & (n_n455) & (n_n491) & (n_n520)));
	assign n_n4492 = (((i_9_) & (n_n455) & (n_n500) & (n_n530)));
	assign n_n4496 = (((i_9_) & (n_n526) & (n_n455) & (n_n500)));
	assign n_n4574 = (((i_9_) & (n_n528) & (n_n390) & (n_n535)));
	assign n_n4572 = (((i_9_) & (n_n390) & (n_n535) & (n_n530)));
	assign n_n4581 = (((!i_1_) & (i_2_) & (i_0_) & (n_n535) & (x20x)));
	assign x256x = (((!i_7_) & (i_8_) & (i_6_) & (x10x) & (n_n509)) + ((i_7_) & (!i_8_) & (i_6_) & (x10x) & (n_n509)));
	assign n_n4623 = (((!i_9_) & (n_n528) & (n_n390) & (n_n500)));
	assign n_n4521 = (((!i_9_) & (n_n482) & (n_n455) & (n_n534)));
	assign x523x = (((i_1_) & (!i_2_) & (i_0_) & (n_n464)));
	assign n_n4557 = (((!i_9_) & (n_n455) & (n_n530) & (n_n464)));
	assign n_n4560 = (((i_9_) & (n_n526) & (n_n455) & (n_n464)));
	assign n_n4553 = (((!i_9_) & (n_n455) & (n_n534) & (n_n464)));
	assign n_n4800 = (((i_9_) & (n_n526) & (n_n473) & (n_n325)));
	assign n_n4780 = (((i_9_) & (n_n482) & (n_n325) & (n_n530)));
	assign n_n4777 = (((!i_9_) & (n_n482) & (n_n534) & (n_n325)));
	assign n_n4783 = (((!i_9_) & (n_n482) & (n_n528) & (n_n325)));
	assign n_n4812 = (((i_9_) & (n_n325) & (n_n530) & (n_n464)));
	assign n_n4811 = (((!i_9_) & (n_n532) & (n_n325) & (n_n464)));
	assign n_n4740 = (((i_9_) & (n_n509) & (n_n325) & (n_n522)));
	assign n_n4710 = (((i_9_) & (n_n325) & (n_n535) & (n_n520)));
	assign n_n4719 = (((!i_9_) & (n_n518) & (n_n528) & (n_n325)));
	assign n_n4708 = (((i_9_) & (n_n325) & (n_n535) & (n_n522)));
	assign n_n4764 = (((i_9_) & (n_n325) & (n_n491) & (n_n530)));
	assign n_n4706 = (((i_9_) & (n_n524) & (n_n325) & (n_n535)));
	assign n_n4699 = (((!i_9_) & (n_n532) & (n_n325) & (n_n535)));
	assign n_n4687 = (((!i_9_) & (n_n528) & (n_n390) & (n_n464)));
	assign n_n4647 = (((!i_1_) & (i_2_) & (i_0_) & (n_n491) & (x23x)));
	assign n_n4656 = (((i_9_) & (n_n526) & (n_n482) & (n_n390)));
	assign n_n4659 = (((!i_9_) & (n_n524) & (n_n482) & (n_n390)));
	assign n_n4675 = (((!i_9_) & (n_n524) & (n_n390) & (n_n473)));
	assign n_n4674 = (((i_9_) & (n_n524) & (n_n390) & (n_n473)));
	assign n_n4661 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n390) & (x20x)));
	assign n_n4671 = (((!i_9_) & (n_n528) & (n_n390) & (n_n473)));
	assign n_n4672 = (((i_9_) & (n_n526) & (n_n390) & (n_n473)));
	assign n_n4685 = (((!i_9_) & (n_n390) & (n_n530) & (n_n464)));
	assign n_n4361 = (((!i_9_) & (n_n536) & (n_n534) & (n_n500)));
	assign n_n4825 = (((!i_9_) & (n_n534) & (n_n260) & (n_n535)));
	assign n_n4824 = (((i_9_) & (n_n534) & (n_n260) & (n_n535)));
	assign n_n4879 = (((!i_9_) & (n_n528) & (n_n260) & (n_n500)));
	assign n_n4937 = (((!i_9_) & (n_n534) & (n_n260) & (n_n464)));
	assign n_n4938 = (((i_9_) & (n_n532) & (n_n260) & (n_n464)));
	assign n_n4936 = (((i_9_) & (n_n534) & (n_n260) & (n_n464)));
	assign n_n5037 = (((!i_9_) & (n_n482) & (n_n195) & (n_n530)));
	assign n_n5043 = (((!i_9_) & (n_n524) & (n_n482) & (n_n195)));
	assign n_n5045 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n195) & (x20x)));
	assign n_n5294 = (((!i_5_) & (!i_3_) & (i_4_) & (x19x) & (n_n528)));
	assign n_n4894 = (((i_9_) & (n_n528) & (n_n260) & (n_n491)));
	assign n_n4916 = (((i_9_) & (n_n482) & (n_n260) & (n_n522)));
	assign n_n4930 = (((i_9_) & (n_n524) & (n_n473) & (n_n260)));
	assign n_n4947 = (((!i_9_) & (n_n524) & (n_n260) & (n_n464)));
	assign x96x = (((!i_7_) & (!i_8_) & (!i_6_) & (x17x) & (n_n491)) + ((!i_7_) & (i_8_) & (!i_6_) & (x17x) & (n_n491)));
	assign x12089x = (((!n_n4920) & (!n_n4907) & (!n_n4950) & (n_n4894)) + ((!n_n4920) & (!n_n4907) & (n_n4950) & (!n_n4894)) + ((!n_n4920) & (!n_n4907) & (n_n4950) & (n_n4894)) + ((!n_n4920) & (n_n4907) & (!n_n4950) & (!n_n4894)) + ((!n_n4920) & (n_n4907) & (!n_n4950) & (n_n4894)) + ((!n_n4920) & (n_n4907) & (n_n4950) & (!n_n4894)) + ((!n_n4920) & (n_n4907) & (n_n4950) & (n_n4894)) + ((n_n4920) & (!n_n4907) & (!n_n4950) & (!n_n4894)) + ((n_n4920) & (!n_n4907) & (!n_n4950) & (n_n4894)) + ((n_n4920) & (!n_n4907) & (n_n4950) & (!n_n4894)) + ((n_n4920) & (!n_n4907) & (n_n4950) & (n_n4894)) + ((n_n4920) & (n_n4907) & (!n_n4950) & (!n_n4894)) + ((n_n4920) & (n_n4907) & (!n_n4950) & (n_n4894)) + ((n_n4920) & (n_n4907) & (n_n4950) & (!n_n4894)) + ((n_n4920) & (n_n4907) & (n_n4950) & (n_n4894)));
	assign x12090x = (((!x17x) & (!x502x) & (!n_n4916) & (!n_n4947) & (x96x)) + ((!x17x) & (!x502x) & (!n_n4916) & (n_n4947) & (!x96x)) + ((!x17x) & (!x502x) & (!n_n4916) & (n_n4947) & (x96x)) + ((!x17x) & (!x502x) & (n_n4916) & (!n_n4947) & (!x96x)) + ((!x17x) & (!x502x) & (n_n4916) & (!n_n4947) & (x96x)) + ((!x17x) & (!x502x) & (n_n4916) & (n_n4947) & (!x96x)) + ((!x17x) & (!x502x) & (n_n4916) & (n_n4947) & (x96x)) + ((!x17x) & (x502x) & (!n_n4916) & (!n_n4947) & (x96x)) + ((!x17x) & (x502x) & (!n_n4916) & (n_n4947) & (!x96x)) + ((!x17x) & (x502x) & (!n_n4916) & (n_n4947) & (x96x)) + ((!x17x) & (x502x) & (n_n4916) & (!n_n4947) & (!x96x)) + ((!x17x) & (x502x) & (n_n4916) & (!n_n4947) & (x96x)) + ((!x17x) & (x502x) & (n_n4916) & (n_n4947) & (!x96x)) + ((!x17x) & (x502x) & (n_n4916) & (n_n4947) & (x96x)) + ((x17x) & (!x502x) & (!n_n4916) & (!n_n4947) & (x96x)) + ((x17x) & (!x502x) & (!n_n4916) & (n_n4947) & (!x96x)) + ((x17x) & (!x502x) & (!n_n4916) & (n_n4947) & (x96x)) + ((x17x) & (!x502x) & (n_n4916) & (!n_n4947) & (!x96x)) + ((x17x) & (!x502x) & (n_n4916) & (!n_n4947) & (x96x)) + ((x17x) & (!x502x) & (n_n4916) & (n_n4947) & (!x96x)) + ((x17x) & (!x502x) & (n_n4916) & (n_n4947) & (x96x)) + ((x17x) & (x502x) & (!n_n4916) & (!n_n4947) & (!x96x)) + ((x17x) & (x502x) & (!n_n4916) & (!n_n4947) & (x96x)) + ((x17x) & (x502x) & (!n_n4916) & (n_n4947) & (!x96x)) + ((x17x) & (x502x) & (!n_n4916) & (n_n4947) & (x96x)) + ((x17x) & (x502x) & (n_n4916) & (!n_n4947) & (!x96x)) + ((x17x) & (x502x) & (n_n4916) & (!n_n4947) & (x96x)) + ((x17x) & (x502x) & (n_n4916) & (n_n4947) & (!x96x)) + ((x17x) & (x502x) & (n_n4916) & (n_n4947) & (x96x)));
	assign n_n5131 = (((!i_9_) & (n_n532) & (n_n130) & (n_n500)));
	assign n_n5137 = (((!i_9_) & (n_n526) & (n_n130) & (n_n500)));
	assign n_n5136 = (((i_7_) & (i_8_) & (!i_6_) & (x12x) & (n_n500)));
	assign n_n5200 = (((i_7_) & (i_8_) & (!i_6_) & (x12x) & (n_n464)));
	assign n_n5206 = (((!i_7_) & (!i_8_) & (!i_6_) & (x12x) & (n_n464)));
	assign n_n5146 = (((i_7_) & (!i_8_) & (i_6_) & (n_n491) & (x12x)));
	assign n_n5204 = (((!i_7_) & (i_8_) & (!i_6_) & (x12x) & (n_n464)));
	assign n_n5191 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n130) & (x23x)));
	assign x12091x = (((!i_9_) & (!n_n532) & (n_n534) & (n_n130) & (n_n500)) + ((!i_9_) & (n_n532) & (!n_n534) & (n_n130) & (n_n500)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n130) & (n_n500)));
	assign x12097x = (((!n_n5146) & (!n_n5204) & (!n_n5191) & (x12091x)) + ((!n_n5146) & (!n_n5204) & (n_n5191) & (!x12091x)) + ((!n_n5146) & (!n_n5204) & (n_n5191) & (x12091x)) + ((!n_n5146) & (n_n5204) & (!n_n5191) & (!x12091x)) + ((!n_n5146) & (n_n5204) & (!n_n5191) & (x12091x)) + ((!n_n5146) & (n_n5204) & (n_n5191) & (!x12091x)) + ((!n_n5146) & (n_n5204) & (n_n5191) & (x12091x)) + ((n_n5146) & (!n_n5204) & (!n_n5191) & (!x12091x)) + ((n_n5146) & (!n_n5204) & (!n_n5191) & (x12091x)) + ((n_n5146) & (!n_n5204) & (n_n5191) & (!x12091x)) + ((n_n5146) & (!n_n5204) & (n_n5191) & (x12091x)) + ((n_n5146) & (n_n5204) & (!n_n5191) & (!x12091x)) + ((n_n5146) & (n_n5204) & (!n_n5191) & (x12091x)) + ((n_n5146) & (n_n5204) & (n_n5191) & (!x12091x)) + ((n_n5146) & (n_n5204) & (n_n5191) & (x12091x)));
	assign n_n1330 = (((!n_n5137) & (!n_n5136) & (!n_n5200) & (!n_n5206) & (x12097x)) + ((!n_n5137) & (!n_n5136) & (!n_n5200) & (n_n5206) & (!x12097x)) + ((!n_n5137) & (!n_n5136) & (!n_n5200) & (n_n5206) & (x12097x)) + ((!n_n5137) & (!n_n5136) & (n_n5200) & (!n_n5206) & (!x12097x)) + ((!n_n5137) & (!n_n5136) & (n_n5200) & (!n_n5206) & (x12097x)) + ((!n_n5137) & (!n_n5136) & (n_n5200) & (n_n5206) & (!x12097x)) + ((!n_n5137) & (!n_n5136) & (n_n5200) & (n_n5206) & (x12097x)) + ((!n_n5137) & (n_n5136) & (!n_n5200) & (!n_n5206) & (!x12097x)) + ((!n_n5137) & (n_n5136) & (!n_n5200) & (!n_n5206) & (x12097x)) + ((!n_n5137) & (n_n5136) & (!n_n5200) & (n_n5206) & (!x12097x)) + ((!n_n5137) & (n_n5136) & (!n_n5200) & (n_n5206) & (x12097x)) + ((!n_n5137) & (n_n5136) & (n_n5200) & (!n_n5206) & (!x12097x)) + ((!n_n5137) & (n_n5136) & (n_n5200) & (!n_n5206) & (x12097x)) + ((!n_n5137) & (n_n5136) & (n_n5200) & (n_n5206) & (!x12097x)) + ((!n_n5137) & (n_n5136) & (n_n5200) & (n_n5206) & (x12097x)) + ((n_n5137) & (!n_n5136) & (!n_n5200) & (!n_n5206) & (!x12097x)) + ((n_n5137) & (!n_n5136) & (!n_n5200) & (!n_n5206) & (x12097x)) + ((n_n5137) & (!n_n5136) & (!n_n5200) & (n_n5206) & (!x12097x)) + ((n_n5137) & (!n_n5136) & (!n_n5200) & (n_n5206) & (x12097x)) + ((n_n5137) & (!n_n5136) & (n_n5200) & (!n_n5206) & (!x12097x)) + ((n_n5137) & (!n_n5136) & (n_n5200) & (!n_n5206) & (x12097x)) + ((n_n5137) & (!n_n5136) & (n_n5200) & (n_n5206) & (!x12097x)) + ((n_n5137) & (!n_n5136) & (n_n5200) & (n_n5206) & (x12097x)) + ((n_n5137) & (n_n5136) & (!n_n5200) & (!n_n5206) & (!x12097x)) + ((n_n5137) & (n_n5136) & (!n_n5200) & (!n_n5206) & (x12097x)) + ((n_n5137) & (n_n5136) & (!n_n5200) & (n_n5206) & (!x12097x)) + ((n_n5137) & (n_n5136) & (!n_n5200) & (n_n5206) & (x12097x)) + ((n_n5137) & (n_n5136) & (n_n5200) & (!n_n5206) & (!x12097x)) + ((n_n5137) & (n_n5136) & (n_n5200) & (!n_n5206) & (x12097x)) + ((n_n5137) & (n_n5136) & (n_n5200) & (n_n5206) & (!x12097x)) + ((n_n5137) & (n_n5136) & (n_n5200) & (n_n5206) & (x12097x)));
	assign n_n5113 = (((!i_9_) & (n_n534) & (n_n509) & (n_n130)));
	assign n_n5081 = (((!i_9_) & (n_n534) & (n_n535) & (n_n130)));
	assign n_n5089 = (((!i_9_) & (n_n526) & (n_n535) & (n_n130)));
	assign n_n5124 = (((i_5_) & (i_3_) & (!i_4_) & (n_n522) & (x12x)));
	assign n_n5114 = (((i_7_) & (!i_8_) & (i_6_) & (n_n509) & (x12x)));
	assign n_n5116 = (((i_5_) & (i_3_) & (!i_4_) & (x12x) & (n_n530)));
	assign x335x = (((!i_7_) & (i_8_) & (i_6_) & (n_n509) & (x12x)) + ((i_7_) & (!i_8_) & (i_6_) & (n_n509) & (x12x)));
	assign n_n5063 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n195) & (x23x)));
	assign x344x = (((!i_9_) & (!n_n532) & (!n_n195) & (!n_n464) & (n_n5063)) + ((!i_9_) & (!n_n532) & (!n_n195) & (n_n464) & (n_n5063)) + ((!i_9_) & (!n_n532) & (n_n195) & (!n_n464) & (n_n5063)) + ((!i_9_) & (!n_n532) & (n_n195) & (n_n464) & (n_n5063)) + ((!i_9_) & (n_n532) & (!n_n195) & (!n_n464) & (n_n5063)) + ((!i_9_) & (n_n532) & (!n_n195) & (n_n464) & (n_n5063)) + ((!i_9_) & (n_n532) & (n_n195) & (!n_n464) & (n_n5063)) + ((!i_9_) & (n_n532) & (n_n195) & (n_n464) & (n_n5063)) + ((i_9_) & (!n_n532) & (!n_n195) & (!n_n464) & (n_n5063)) + ((i_9_) & (!n_n532) & (!n_n195) & (n_n464) & (n_n5063)) + ((i_9_) & (!n_n532) & (n_n195) & (!n_n464) & (n_n5063)) + ((i_9_) & (!n_n532) & (n_n195) & (n_n464) & (n_n5063)) + ((i_9_) & (n_n532) & (!n_n195) & (!n_n464) & (n_n5063)) + ((i_9_) & (n_n532) & (!n_n195) & (n_n464) & (n_n5063)) + ((i_9_) & (n_n532) & (n_n195) & (!n_n464) & (n_n5063)) + ((i_9_) & (n_n532) & (n_n195) & (n_n464) & (!n_n5063)) + ((i_9_) & (n_n532) & (n_n195) & (n_n464) & (n_n5063)));
	assign x12099x = (((!i_9_) & (!n_n526) & (n_n534) & (n_n535) & (n_n130)) + ((!i_9_) & (n_n526) & (!n_n534) & (n_n535) & (n_n130)) + ((!i_9_) & (n_n526) & (n_n534) & (n_n535) & (n_n130)));
	assign x12100x = (((!i_7_) & (i_8_) & (!i_6_) & (n_n509) & (x12x)) + ((!i_7_) & (i_8_) & (i_6_) & (n_n509) & (x12x)) + ((i_7_) & (!i_8_) & (i_6_) & (n_n509) & (x12x)));
	assign n_n1331 = (((!n_n5096) & (!n_n5113) & (!x344x) & (!x12099x) & (x12100x)) + ((!n_n5096) & (!n_n5113) & (!x344x) & (x12099x) & (!x12100x)) + ((!n_n5096) & (!n_n5113) & (!x344x) & (x12099x) & (x12100x)) + ((!n_n5096) & (!n_n5113) & (x344x) & (!x12099x) & (!x12100x)) + ((!n_n5096) & (!n_n5113) & (x344x) & (!x12099x) & (x12100x)) + ((!n_n5096) & (!n_n5113) & (x344x) & (x12099x) & (!x12100x)) + ((!n_n5096) & (!n_n5113) & (x344x) & (x12099x) & (x12100x)) + ((!n_n5096) & (n_n5113) & (!x344x) & (!x12099x) & (!x12100x)) + ((!n_n5096) & (n_n5113) & (!x344x) & (!x12099x) & (x12100x)) + ((!n_n5096) & (n_n5113) & (!x344x) & (x12099x) & (!x12100x)) + ((!n_n5096) & (n_n5113) & (!x344x) & (x12099x) & (x12100x)) + ((!n_n5096) & (n_n5113) & (x344x) & (!x12099x) & (!x12100x)) + ((!n_n5096) & (n_n5113) & (x344x) & (!x12099x) & (x12100x)) + ((!n_n5096) & (n_n5113) & (x344x) & (x12099x) & (!x12100x)) + ((!n_n5096) & (n_n5113) & (x344x) & (x12099x) & (x12100x)) + ((n_n5096) & (!n_n5113) & (!x344x) & (!x12099x) & (!x12100x)) + ((n_n5096) & (!n_n5113) & (!x344x) & (!x12099x) & (x12100x)) + ((n_n5096) & (!n_n5113) & (!x344x) & (x12099x) & (!x12100x)) + ((n_n5096) & (!n_n5113) & (!x344x) & (x12099x) & (x12100x)) + ((n_n5096) & (!n_n5113) & (x344x) & (!x12099x) & (!x12100x)) + ((n_n5096) & (!n_n5113) & (x344x) & (!x12099x) & (x12100x)) + ((n_n5096) & (!n_n5113) & (x344x) & (x12099x) & (!x12100x)) + ((n_n5096) & (!n_n5113) & (x344x) & (x12099x) & (x12100x)) + ((n_n5096) & (n_n5113) & (!x344x) & (!x12099x) & (!x12100x)) + ((n_n5096) & (n_n5113) & (!x344x) & (!x12099x) & (x12100x)) + ((n_n5096) & (n_n5113) & (!x344x) & (x12099x) & (!x12100x)) + ((n_n5096) & (n_n5113) & (!x344x) & (x12099x) & (x12100x)) + ((n_n5096) & (n_n5113) & (x344x) & (!x12099x) & (!x12100x)) + ((n_n5096) & (n_n5113) & (x344x) & (!x12099x) & (x12100x)) + ((n_n5096) & (n_n5113) & (x344x) & (x12099x) & (!x12100x)) + ((n_n5096) & (n_n5113) & (x344x) & (x12099x) & (x12100x)));
	assign n_n5258 = (((i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n500)));
	assign n_n5274 = (((i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n491)));
	assign n_n5232 = (((!i_5_) & (i_3_) & (i_4_) & (x19x) & (n_n526)));
	assign n_n5255 = (((i_5_) & (i_3_) & (!i_4_) & (x23x) & (n_n65)));
	assign n_n5267 = (((!i_9_) & (n_n524) & (n_n500) & (n_n65)));
	assign n_n5216 = (((i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n535)));
	assign n_n5222 = (((i_5_) & (i_3_) & (i_4_) & (x19x) & (n_n520)));
	assign n_n5212 = (((i_5_) & (i_3_) & (i_4_) & (x19x) & (n_n530)));
	assign x12109x = (((!n_n5244) & (!n_n5258) & (!n_n5216) & (!n_n5222) & (n_n5212)) + ((!n_n5244) & (!n_n5258) & (!n_n5216) & (n_n5222) & (!n_n5212)) + ((!n_n5244) & (!n_n5258) & (!n_n5216) & (n_n5222) & (n_n5212)) + ((!n_n5244) & (!n_n5258) & (n_n5216) & (!n_n5222) & (!n_n5212)) + ((!n_n5244) & (!n_n5258) & (n_n5216) & (!n_n5222) & (n_n5212)) + ((!n_n5244) & (!n_n5258) & (n_n5216) & (n_n5222) & (!n_n5212)) + ((!n_n5244) & (!n_n5258) & (n_n5216) & (n_n5222) & (n_n5212)) + ((!n_n5244) & (n_n5258) & (!n_n5216) & (!n_n5222) & (!n_n5212)) + ((!n_n5244) & (n_n5258) & (!n_n5216) & (!n_n5222) & (n_n5212)) + ((!n_n5244) & (n_n5258) & (!n_n5216) & (n_n5222) & (!n_n5212)) + ((!n_n5244) & (n_n5258) & (!n_n5216) & (n_n5222) & (n_n5212)) + ((!n_n5244) & (n_n5258) & (n_n5216) & (!n_n5222) & (!n_n5212)) + ((!n_n5244) & (n_n5258) & (n_n5216) & (!n_n5222) & (n_n5212)) + ((!n_n5244) & (n_n5258) & (n_n5216) & (n_n5222) & (!n_n5212)) + ((!n_n5244) & (n_n5258) & (n_n5216) & (n_n5222) & (n_n5212)) + ((n_n5244) & (!n_n5258) & (!n_n5216) & (!n_n5222) & (!n_n5212)) + ((n_n5244) & (!n_n5258) & (!n_n5216) & (!n_n5222) & (n_n5212)) + ((n_n5244) & (!n_n5258) & (!n_n5216) & (n_n5222) & (!n_n5212)) + ((n_n5244) & (!n_n5258) & (!n_n5216) & (n_n5222) & (n_n5212)) + ((n_n5244) & (!n_n5258) & (n_n5216) & (!n_n5222) & (!n_n5212)) + ((n_n5244) & (!n_n5258) & (n_n5216) & (!n_n5222) & (n_n5212)) + ((n_n5244) & (!n_n5258) & (n_n5216) & (n_n5222) & (!n_n5212)) + ((n_n5244) & (!n_n5258) & (n_n5216) & (n_n5222) & (n_n5212)) + ((n_n5244) & (n_n5258) & (!n_n5216) & (!n_n5222) & (!n_n5212)) + ((n_n5244) & (n_n5258) & (!n_n5216) & (!n_n5222) & (n_n5212)) + ((n_n5244) & (n_n5258) & (!n_n5216) & (n_n5222) & (!n_n5212)) + ((n_n5244) & (n_n5258) & (!n_n5216) & (n_n5222) & (n_n5212)) + ((n_n5244) & (n_n5258) & (n_n5216) & (!n_n5222) & (!n_n5212)) + ((n_n5244) & (n_n5258) & (n_n5216) & (!n_n5222) & (n_n5212)) + ((n_n5244) & (n_n5258) & (n_n5216) & (n_n5222) & (!n_n5212)) + ((n_n5244) & (n_n5258) & (n_n5216) & (n_n5222) & (n_n5212)));
	assign x12110x = (((!n_n5274) & (!n_n5232) & (!n_n5255) & (!n_n5267) & (x12109x)) + ((!n_n5274) & (!n_n5232) & (!n_n5255) & (n_n5267) & (!x12109x)) + ((!n_n5274) & (!n_n5232) & (!n_n5255) & (n_n5267) & (x12109x)) + ((!n_n5274) & (!n_n5232) & (n_n5255) & (!n_n5267) & (!x12109x)) + ((!n_n5274) & (!n_n5232) & (n_n5255) & (!n_n5267) & (x12109x)) + ((!n_n5274) & (!n_n5232) & (n_n5255) & (n_n5267) & (!x12109x)) + ((!n_n5274) & (!n_n5232) & (n_n5255) & (n_n5267) & (x12109x)) + ((!n_n5274) & (n_n5232) & (!n_n5255) & (!n_n5267) & (!x12109x)) + ((!n_n5274) & (n_n5232) & (!n_n5255) & (!n_n5267) & (x12109x)) + ((!n_n5274) & (n_n5232) & (!n_n5255) & (n_n5267) & (!x12109x)) + ((!n_n5274) & (n_n5232) & (!n_n5255) & (n_n5267) & (x12109x)) + ((!n_n5274) & (n_n5232) & (n_n5255) & (!n_n5267) & (!x12109x)) + ((!n_n5274) & (n_n5232) & (n_n5255) & (!n_n5267) & (x12109x)) + ((!n_n5274) & (n_n5232) & (n_n5255) & (n_n5267) & (!x12109x)) + ((!n_n5274) & (n_n5232) & (n_n5255) & (n_n5267) & (x12109x)) + ((n_n5274) & (!n_n5232) & (!n_n5255) & (!n_n5267) & (!x12109x)) + ((n_n5274) & (!n_n5232) & (!n_n5255) & (!n_n5267) & (x12109x)) + ((n_n5274) & (!n_n5232) & (!n_n5255) & (n_n5267) & (!x12109x)) + ((n_n5274) & (!n_n5232) & (!n_n5255) & (n_n5267) & (x12109x)) + ((n_n5274) & (!n_n5232) & (n_n5255) & (!n_n5267) & (!x12109x)) + ((n_n5274) & (!n_n5232) & (n_n5255) & (!n_n5267) & (x12109x)) + ((n_n5274) & (!n_n5232) & (n_n5255) & (n_n5267) & (!x12109x)) + ((n_n5274) & (!n_n5232) & (n_n5255) & (n_n5267) & (x12109x)) + ((n_n5274) & (n_n5232) & (!n_n5255) & (!n_n5267) & (!x12109x)) + ((n_n5274) & (n_n5232) & (!n_n5255) & (!n_n5267) & (x12109x)) + ((n_n5274) & (n_n5232) & (!n_n5255) & (n_n5267) & (!x12109x)) + ((n_n5274) & (n_n5232) & (!n_n5255) & (n_n5267) & (x12109x)) + ((n_n5274) & (n_n5232) & (n_n5255) & (!n_n5267) & (!x12109x)) + ((n_n5274) & (n_n5232) & (n_n5255) & (!n_n5267) & (x12109x)) + ((n_n5274) & (n_n5232) & (n_n5255) & (n_n5267) & (!x12109x)) + ((n_n5274) & (n_n5232) & (n_n5255) & (n_n5267) & (x12109x)));
	assign n_n4343 = (((i_1_) & (i_2_) & (i_0_) & (n_n518) & (x23x)));
	assign n_n4393 = (((!i_9_) & (n_n536) & (n_n482) & (n_n534)));
	assign n_n4611 = (((!i_9_) & (n_n524) & (n_n390) & (n_n509)));
	assign n_n4669 = (((!i_9_) & (n_n390) & (n_n473) & (n_n530)));
	assign n_n4673 = (((!i_9_) & (n_n526) & (n_n390) & (n_n473)));
	assign n_n4668 = (((i_9_) & (n_n390) & (n_n473) & (n_n530)));
	assign n_n4792 = (((i_9_) & (n_n473) & (n_n534) & (n_n325)));
	assign n_n4908 = (((i_9_) & (n_n482) & (n_n260) & (n_n530)));
	assign n_n4966 = (((i_9_) & (n_n535) & (n_n520) & (n_n195)));
	assign n_n4968 = (((i_9_) & (n_n518) & (n_n534) & (n_n195)));
	assign n_n5012 = (((i_9_) & (n_n522) & (n_n195) & (n_n500)));
	assign n_n5067 = (((!i_9_) & (n_n532) & (n_n195) & (n_n464)));
	assign n_n5069 = (((!i_9_) & (n_n195) & (n_n530) & (n_n464)));
	assign n_n5243 = (((!i_9_) & (n_n532) & (n_n509) & (n_n65)));
	assign n_n5300 = (((!i_5_) & (!i_3_) & (i_4_) & (x19x) & (n_n522)));
	assign n_n5299 = (((!i_9_) & (n_n524) & (n_n482) & (n_n65)));
	assign n_n4364 = (((i_9_) & (n_n536) & (n_n500) & (n_n530)));
	assign n_n3533 = (((!i_9_) & (n_n536) & (n_n532) & (n_n500) & (!n_n530)) + ((!i_9_) & (n_n536) & (n_n532) & (n_n500) & (n_n530)) + ((i_9_) & (n_n536) & (!n_n532) & (n_n500) & (n_n530)) + ((i_9_) & (n_n536) & (n_n532) & (n_n500) & (!n_n530)) + ((i_9_) & (n_n536) & (n_n532) & (n_n500) & (n_n530)));
	assign n_n4366 = (((i_9_) & (n_n536) & (n_n528) & (n_n500)));
	assign n_n4365 = (((!i_9_) & (n_n536) & (n_n500) & (n_n530)));
	assign n_n1308 = (((!i_9_) & (n_n536) & (!n_n528) & (n_n500) & (n_n530)) + ((!i_9_) & (n_n536) & (n_n528) & (n_n500) & (!n_n530)) + ((!i_9_) & (n_n536) & (n_n528) & (n_n500) & (n_n530)) + ((i_9_) & (n_n536) & (n_n528) & (n_n500) & (!n_n530)) + ((i_9_) & (n_n536) & (n_n528) & (n_n500) & (n_n530)));
	assign n_n4769 = (((!i_9_) & (n_n526) & (n_n325) & (n_n491)));
	assign n_n4765 = (((!i_9_) & (n_n325) & (n_n491) & (n_n530)));
	assign n_n4766 = (((i_9_) & (n_n528) & (n_n325) & (n_n491)));
	assign x316x = (((!x14x) & (!n_n522) & (!n_n491) & (!n_n520) & (n_n4771)) + ((!x14x) & (!n_n522) & (!n_n491) & (n_n520) & (n_n4771)) + ((!x14x) & (!n_n522) & (n_n491) & (!n_n520) & (n_n4771)) + ((!x14x) & (!n_n522) & (n_n491) & (n_n520) & (n_n4771)) + ((!x14x) & (n_n522) & (!n_n491) & (!n_n520) & (n_n4771)) + ((!x14x) & (n_n522) & (!n_n491) & (n_n520) & (n_n4771)) + ((!x14x) & (n_n522) & (n_n491) & (!n_n520) & (n_n4771)) + ((!x14x) & (n_n522) & (n_n491) & (n_n520) & (n_n4771)) + ((x14x) & (!n_n522) & (!n_n491) & (!n_n520) & (n_n4771)) + ((x14x) & (!n_n522) & (!n_n491) & (n_n520) & (n_n4771)) + ((x14x) & (!n_n522) & (n_n491) & (!n_n520) & (n_n4771)) + ((x14x) & (!n_n522) & (n_n491) & (n_n520) & (!n_n4771)) + ((x14x) & (!n_n522) & (n_n491) & (n_n520) & (n_n4771)) + ((x14x) & (n_n522) & (!n_n491) & (!n_n520) & (n_n4771)) + ((x14x) & (n_n522) & (!n_n491) & (n_n520) & (n_n4771)) + ((x14x) & (n_n522) & (n_n491) & (!n_n520) & (!n_n4771)) + ((x14x) & (n_n522) & (n_n491) & (!n_n520) & (n_n4771)) + ((x14x) & (n_n522) & (n_n491) & (n_n520) & (!n_n4771)) + ((x14x) & (n_n522) & (n_n491) & (n_n520) & (n_n4771)));
	assign x11749x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n325) & (n_n491)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n325) & (n_n491)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n325) & (n_n491)) + ((i_9_) & (n_n524) & (n_n526) & (n_n325) & (n_n491)));
	assign n_n1086 = (((!n_n4767) & (!n_n4764) & (!x165x) & (!x316x) & (x11749x)) + ((!n_n4767) & (!n_n4764) & (!x165x) & (x316x) & (!x11749x)) + ((!n_n4767) & (!n_n4764) & (!x165x) & (x316x) & (x11749x)) + ((!n_n4767) & (!n_n4764) & (x165x) & (!x316x) & (!x11749x)) + ((!n_n4767) & (!n_n4764) & (x165x) & (!x316x) & (x11749x)) + ((!n_n4767) & (!n_n4764) & (x165x) & (x316x) & (!x11749x)) + ((!n_n4767) & (!n_n4764) & (x165x) & (x316x) & (x11749x)) + ((!n_n4767) & (n_n4764) & (!x165x) & (!x316x) & (!x11749x)) + ((!n_n4767) & (n_n4764) & (!x165x) & (!x316x) & (x11749x)) + ((!n_n4767) & (n_n4764) & (!x165x) & (x316x) & (!x11749x)) + ((!n_n4767) & (n_n4764) & (!x165x) & (x316x) & (x11749x)) + ((!n_n4767) & (n_n4764) & (x165x) & (!x316x) & (!x11749x)) + ((!n_n4767) & (n_n4764) & (x165x) & (!x316x) & (x11749x)) + ((!n_n4767) & (n_n4764) & (x165x) & (x316x) & (!x11749x)) + ((!n_n4767) & (n_n4764) & (x165x) & (x316x) & (x11749x)) + ((n_n4767) & (!n_n4764) & (!x165x) & (!x316x) & (!x11749x)) + ((n_n4767) & (!n_n4764) & (!x165x) & (!x316x) & (x11749x)) + ((n_n4767) & (!n_n4764) & (!x165x) & (x316x) & (!x11749x)) + ((n_n4767) & (!n_n4764) & (!x165x) & (x316x) & (x11749x)) + ((n_n4767) & (!n_n4764) & (x165x) & (!x316x) & (!x11749x)) + ((n_n4767) & (!n_n4764) & (x165x) & (!x316x) & (x11749x)) + ((n_n4767) & (!n_n4764) & (x165x) & (x316x) & (!x11749x)) + ((n_n4767) & (!n_n4764) & (x165x) & (x316x) & (x11749x)) + ((n_n4767) & (n_n4764) & (!x165x) & (!x316x) & (!x11749x)) + ((n_n4767) & (n_n4764) & (!x165x) & (!x316x) & (x11749x)) + ((n_n4767) & (n_n4764) & (!x165x) & (x316x) & (!x11749x)) + ((n_n4767) & (n_n4764) & (!x165x) & (x316x) & (x11749x)) + ((n_n4767) & (n_n4764) & (x165x) & (!x316x) & (!x11749x)) + ((n_n4767) & (n_n4764) & (x165x) & (!x316x) & (x11749x)) + ((n_n4767) & (n_n4764) & (x165x) & (x316x) & (!x11749x)) + ((n_n4767) & (n_n4764) & (x165x) & (x316x) & (x11749x)));
	assign n_n4905 = (((!i_9_) & (n_n482) & (n_n534) & (n_n260)));
	assign x306x = (((!i_9_) & (!n_n526) & (n_n482) & (n_n528) & (n_n260)) + ((!i_9_) & (n_n526) & (n_n482) & (n_n528) & (n_n260)) + ((i_9_) & (n_n526) & (n_n482) & (!n_n528) & (n_n260)) + ((i_9_) & (n_n526) & (n_n482) & (n_n528) & (n_n260)));
	assign n_n4914 = (((i_9_) & (n_n524) & (n_n482) & (n_n260)));
	assign x352x = (((i_7_) & (!i_8_) & (i_6_) & (n_n482) & (x17x)) + ((i_7_) & (i_8_) & (i_6_) & (n_n482) & (x17x)));
	assign x11786x = (((!n_n4911) & (!n_n4916) & (!n_n4912) & (!n_n4908) & (n_n4905)) + ((!n_n4911) & (!n_n4916) & (!n_n4912) & (n_n4908) & (!n_n4905)) + ((!n_n4911) & (!n_n4916) & (!n_n4912) & (n_n4908) & (n_n4905)) + ((!n_n4911) & (!n_n4916) & (n_n4912) & (!n_n4908) & (!n_n4905)) + ((!n_n4911) & (!n_n4916) & (n_n4912) & (!n_n4908) & (n_n4905)) + ((!n_n4911) & (!n_n4916) & (n_n4912) & (n_n4908) & (!n_n4905)) + ((!n_n4911) & (!n_n4916) & (n_n4912) & (n_n4908) & (n_n4905)) + ((!n_n4911) & (n_n4916) & (!n_n4912) & (!n_n4908) & (!n_n4905)) + ((!n_n4911) & (n_n4916) & (!n_n4912) & (!n_n4908) & (n_n4905)) + ((!n_n4911) & (n_n4916) & (!n_n4912) & (n_n4908) & (!n_n4905)) + ((!n_n4911) & (n_n4916) & (!n_n4912) & (n_n4908) & (n_n4905)) + ((!n_n4911) & (n_n4916) & (n_n4912) & (!n_n4908) & (!n_n4905)) + ((!n_n4911) & (n_n4916) & (n_n4912) & (!n_n4908) & (n_n4905)) + ((!n_n4911) & (n_n4916) & (n_n4912) & (n_n4908) & (!n_n4905)) + ((!n_n4911) & (n_n4916) & (n_n4912) & (n_n4908) & (n_n4905)) + ((n_n4911) & (!n_n4916) & (!n_n4912) & (!n_n4908) & (!n_n4905)) + ((n_n4911) & (!n_n4916) & (!n_n4912) & (!n_n4908) & (n_n4905)) + ((n_n4911) & (!n_n4916) & (!n_n4912) & (n_n4908) & (!n_n4905)) + ((n_n4911) & (!n_n4916) & (!n_n4912) & (n_n4908) & (n_n4905)) + ((n_n4911) & (!n_n4916) & (n_n4912) & (!n_n4908) & (!n_n4905)) + ((n_n4911) & (!n_n4916) & (n_n4912) & (!n_n4908) & (n_n4905)) + ((n_n4911) & (!n_n4916) & (n_n4912) & (n_n4908) & (!n_n4905)) + ((n_n4911) & (!n_n4916) & (n_n4912) & (n_n4908) & (n_n4905)) + ((n_n4911) & (n_n4916) & (!n_n4912) & (!n_n4908) & (!n_n4905)) + ((n_n4911) & (n_n4916) & (!n_n4912) & (!n_n4908) & (n_n4905)) + ((n_n4911) & (n_n4916) & (!n_n4912) & (n_n4908) & (!n_n4905)) + ((n_n4911) & (n_n4916) & (!n_n4912) & (n_n4908) & (n_n4905)) + ((n_n4911) & (n_n4916) & (n_n4912) & (!n_n4908) & (!n_n4905)) + ((n_n4911) & (n_n4916) & (n_n4912) & (!n_n4908) & (n_n4905)) + ((n_n4911) & (n_n4916) & (n_n4912) & (n_n4908) & (!n_n4905)) + ((n_n4911) & (n_n4916) & (n_n4912) & (n_n4908) & (n_n4905)));
	assign n_n1075 = (((!x351x) & (!x352x) & (x11786x)) + ((!x351x) & (x352x) & (!x11786x)) + ((!x351x) & (x352x) & (x11786x)) + ((x351x) & (!x352x) & (!x11786x)) + ((x351x) & (!x352x) & (x11786x)) + ((x351x) & (x352x) & (!x11786x)) + ((x351x) & (x352x) & (x11786x)));
	assign n_n5056 = (((i_9_) & (n_n526) & (n_n473) & (n_n195)));
	assign n_n5053 = (((!i_9_) & (n_n473) & (n_n195) & (n_n530)));
	assign n_n5052 = (((i_9_) & (n_n473) & (n_n195) & (n_n530)));
	assign x166x = (((!i_9_) & (n_n473) & (n_n195) & (n_n530)) + ((i_9_) & (n_n473) & (n_n195) & (n_n530)));
	assign x22155x = (((!n_n5050) & (!n_n5055) & (!n_n5059) & (!n_n5045)));
	assign n_n1064 = (((!n_n5057) & (!n_n5046) & (!n_n5056) & (!x166x) & (!x22155x)) + ((!n_n5057) & (!n_n5046) & (!n_n5056) & (x166x) & (!x22155x)) + ((!n_n5057) & (!n_n5046) & (!n_n5056) & (x166x) & (x22155x)) + ((!n_n5057) & (!n_n5046) & (n_n5056) & (!x166x) & (!x22155x)) + ((!n_n5057) & (!n_n5046) & (n_n5056) & (!x166x) & (x22155x)) + ((!n_n5057) & (!n_n5046) & (n_n5056) & (x166x) & (!x22155x)) + ((!n_n5057) & (!n_n5046) & (n_n5056) & (x166x) & (x22155x)) + ((!n_n5057) & (n_n5046) & (!n_n5056) & (!x166x) & (!x22155x)) + ((!n_n5057) & (n_n5046) & (!n_n5056) & (!x166x) & (x22155x)) + ((!n_n5057) & (n_n5046) & (!n_n5056) & (x166x) & (!x22155x)) + ((!n_n5057) & (n_n5046) & (!n_n5056) & (x166x) & (x22155x)) + ((!n_n5057) & (n_n5046) & (n_n5056) & (!x166x) & (!x22155x)) + ((!n_n5057) & (n_n5046) & (n_n5056) & (!x166x) & (x22155x)) + ((!n_n5057) & (n_n5046) & (n_n5056) & (x166x) & (!x22155x)) + ((!n_n5057) & (n_n5046) & (n_n5056) & (x166x) & (x22155x)) + ((n_n5057) & (!n_n5046) & (!n_n5056) & (!x166x) & (!x22155x)) + ((n_n5057) & (!n_n5046) & (!n_n5056) & (!x166x) & (x22155x)) + ((n_n5057) & (!n_n5046) & (!n_n5056) & (x166x) & (!x22155x)) + ((n_n5057) & (!n_n5046) & (!n_n5056) & (x166x) & (x22155x)) + ((n_n5057) & (!n_n5046) & (n_n5056) & (!x166x) & (!x22155x)) + ((n_n5057) & (!n_n5046) & (n_n5056) & (!x166x) & (x22155x)) + ((n_n5057) & (!n_n5046) & (n_n5056) & (x166x) & (!x22155x)) + ((n_n5057) & (!n_n5046) & (n_n5056) & (x166x) & (x22155x)) + ((n_n5057) & (n_n5046) & (!n_n5056) & (!x166x) & (!x22155x)) + ((n_n5057) & (n_n5046) & (!n_n5056) & (!x166x) & (x22155x)) + ((n_n5057) & (n_n5046) & (!n_n5056) & (x166x) & (!x22155x)) + ((n_n5057) & (n_n5046) & (!n_n5056) & (x166x) & (x22155x)) + ((n_n5057) & (n_n5046) & (n_n5056) & (!x166x) & (!x22155x)) + ((n_n5057) & (n_n5046) & (n_n5056) & (!x166x) & (x22155x)) + ((n_n5057) & (n_n5046) & (n_n5056) & (x166x) & (!x22155x)) + ((n_n5057) & (n_n5046) & (n_n5056) & (x166x) & (x22155x)));
	assign x179x = (((!i_9_) & (n_n473) & (n_n532) & (n_n325)) + ((i_9_) & (n_n473) & (n_n532) & (n_n325)));
	assign n_n2003 = (((!i_9_) & (n_n473) & (!n_n532) & (n_n534) & (n_n325)) + ((!i_9_) & (n_n473) & (n_n532) & (!n_n534) & (n_n325)) + ((!i_9_) & (n_n473) & (n_n532) & (n_n534) & (n_n325)) + ((i_9_) & (n_n473) & (n_n532) & (!n_n534) & (n_n325)) + ((i_9_) & (n_n473) & (n_n532) & (n_n534) & (n_n325)));
	assign n_n4806 = (((i_9_) & (n_n473) & (n_n325) & (n_n520)));
	assign n_n4807 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n325) & (x23x)));
	assign x11757x = (((!n_n4803) & (!n_n4804) & (!n_n4806) & (!n_n4802) & (n_n4807)) + ((!n_n4803) & (!n_n4804) & (!n_n4806) & (n_n4802) & (!n_n4807)) + ((!n_n4803) & (!n_n4804) & (!n_n4806) & (n_n4802) & (n_n4807)) + ((!n_n4803) & (!n_n4804) & (n_n4806) & (!n_n4802) & (!n_n4807)) + ((!n_n4803) & (!n_n4804) & (n_n4806) & (!n_n4802) & (n_n4807)) + ((!n_n4803) & (!n_n4804) & (n_n4806) & (n_n4802) & (!n_n4807)) + ((!n_n4803) & (!n_n4804) & (n_n4806) & (n_n4802) & (n_n4807)) + ((!n_n4803) & (n_n4804) & (!n_n4806) & (!n_n4802) & (!n_n4807)) + ((!n_n4803) & (n_n4804) & (!n_n4806) & (!n_n4802) & (n_n4807)) + ((!n_n4803) & (n_n4804) & (!n_n4806) & (n_n4802) & (!n_n4807)) + ((!n_n4803) & (n_n4804) & (!n_n4806) & (n_n4802) & (n_n4807)) + ((!n_n4803) & (n_n4804) & (n_n4806) & (!n_n4802) & (!n_n4807)) + ((!n_n4803) & (n_n4804) & (n_n4806) & (!n_n4802) & (n_n4807)) + ((!n_n4803) & (n_n4804) & (n_n4806) & (n_n4802) & (!n_n4807)) + ((!n_n4803) & (n_n4804) & (n_n4806) & (n_n4802) & (n_n4807)) + ((n_n4803) & (!n_n4804) & (!n_n4806) & (!n_n4802) & (!n_n4807)) + ((n_n4803) & (!n_n4804) & (!n_n4806) & (!n_n4802) & (n_n4807)) + ((n_n4803) & (!n_n4804) & (!n_n4806) & (n_n4802) & (!n_n4807)) + ((n_n4803) & (!n_n4804) & (!n_n4806) & (n_n4802) & (n_n4807)) + ((n_n4803) & (!n_n4804) & (n_n4806) & (!n_n4802) & (!n_n4807)) + ((n_n4803) & (!n_n4804) & (n_n4806) & (!n_n4802) & (n_n4807)) + ((n_n4803) & (!n_n4804) & (n_n4806) & (n_n4802) & (!n_n4807)) + ((n_n4803) & (!n_n4804) & (n_n4806) & (n_n4802) & (n_n4807)) + ((n_n4803) & (n_n4804) & (!n_n4806) & (!n_n4802) & (!n_n4807)) + ((n_n4803) & (n_n4804) & (!n_n4806) & (!n_n4802) & (n_n4807)) + ((n_n4803) & (n_n4804) & (!n_n4806) & (n_n4802) & (!n_n4807)) + ((n_n4803) & (n_n4804) & (!n_n4806) & (n_n4802) & (n_n4807)) + ((n_n4803) & (n_n4804) & (n_n4806) & (!n_n4802) & (!n_n4807)) + ((n_n4803) & (n_n4804) & (n_n4806) & (!n_n4802) & (n_n4807)) + ((n_n4803) & (n_n4804) & (n_n4806) & (n_n4802) & (!n_n4807)) + ((n_n4803) & (n_n4804) & (n_n4806) & (n_n4802) & (n_n4807)));
	assign x439x = (((!i_9_) & (!n_n532) & (n_n534) & (n_n325) & (n_n464)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n325) & (n_n464)) + ((i_9_) & (n_n532) & (!n_n534) & (n_n325) & (n_n464)) + ((i_9_) & (n_n532) & (n_n534) & (n_n325) & (n_n464)));
	assign n_n4821 = (((!i_1_) & (!i_2_) & (i_0_) & (x20x) & (n_n464)));
	assign n_n4822 = (((i_9_) & (n_n325) & (n_n520) & (n_n464)));
	assign n_n4818 = (((i_9_) & (n_n524) & (n_n325) & (n_n464)));
	assign n_n4819 = (((!i_9_) & (n_n524) & (n_n325) & (n_n464)));
	assign x85x = (((i_9_) & (n_n528) & (n_n325) & (n_n464)));
	assign x11762x = (((!n_n4821) & (!n_n4822) & (!n_n4818) & (!n_n4819) & (x85x)) + ((!n_n4821) & (!n_n4822) & (!n_n4818) & (n_n4819) & (!x85x)) + ((!n_n4821) & (!n_n4822) & (!n_n4818) & (n_n4819) & (x85x)) + ((!n_n4821) & (!n_n4822) & (n_n4818) & (!n_n4819) & (!x85x)) + ((!n_n4821) & (!n_n4822) & (n_n4818) & (!n_n4819) & (x85x)) + ((!n_n4821) & (!n_n4822) & (n_n4818) & (n_n4819) & (!x85x)) + ((!n_n4821) & (!n_n4822) & (n_n4818) & (n_n4819) & (x85x)) + ((!n_n4821) & (n_n4822) & (!n_n4818) & (!n_n4819) & (!x85x)) + ((!n_n4821) & (n_n4822) & (!n_n4818) & (!n_n4819) & (x85x)) + ((!n_n4821) & (n_n4822) & (!n_n4818) & (n_n4819) & (!x85x)) + ((!n_n4821) & (n_n4822) & (!n_n4818) & (n_n4819) & (x85x)) + ((!n_n4821) & (n_n4822) & (n_n4818) & (!n_n4819) & (!x85x)) + ((!n_n4821) & (n_n4822) & (n_n4818) & (!n_n4819) & (x85x)) + ((!n_n4821) & (n_n4822) & (n_n4818) & (n_n4819) & (!x85x)) + ((!n_n4821) & (n_n4822) & (n_n4818) & (n_n4819) & (x85x)) + ((n_n4821) & (!n_n4822) & (!n_n4818) & (!n_n4819) & (!x85x)) + ((n_n4821) & (!n_n4822) & (!n_n4818) & (!n_n4819) & (x85x)) + ((n_n4821) & (!n_n4822) & (!n_n4818) & (n_n4819) & (!x85x)) + ((n_n4821) & (!n_n4822) & (!n_n4818) & (n_n4819) & (x85x)) + ((n_n4821) & (!n_n4822) & (n_n4818) & (!n_n4819) & (!x85x)) + ((n_n4821) & (!n_n4822) & (n_n4818) & (!n_n4819) & (x85x)) + ((n_n4821) & (!n_n4822) & (n_n4818) & (n_n4819) & (!x85x)) + ((n_n4821) & (!n_n4822) & (n_n4818) & (n_n4819) & (x85x)) + ((n_n4821) & (n_n4822) & (!n_n4818) & (!n_n4819) & (!x85x)) + ((n_n4821) & (n_n4822) & (!n_n4818) & (!n_n4819) & (x85x)) + ((n_n4821) & (n_n4822) & (!n_n4818) & (n_n4819) & (!x85x)) + ((n_n4821) & (n_n4822) & (!n_n4818) & (n_n4819) & (x85x)) + ((n_n4821) & (n_n4822) & (n_n4818) & (!n_n4819) & (!x85x)) + ((n_n4821) & (n_n4822) & (n_n4818) & (!n_n4819) & (x85x)) + ((n_n4821) & (n_n4822) & (n_n4818) & (n_n4819) & (!x85x)) + ((n_n4821) & (n_n4822) & (n_n4818) & (n_n4819) & (x85x)));
	assign x151x = (((!i_9_) & (!n_n526) & (n_n528) & (n_n325) & (n_n464)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n325) & (n_n464)) + ((i_9_) & (n_n526) & (!n_n528) & (n_n325) & (n_n464)) + ((i_9_) & (n_n526) & (n_n528) & (n_n325) & (n_n464)));
	assign x292x = (((!i_9_) & (n_n482) & (n_n325) & (!n_n520) & (x23x)) + ((!i_9_) & (n_n482) & (n_n325) & (n_n520) & (x23x)) + ((i_9_) & (n_n482) & (n_n325) & (!n_n520) & (x23x)) + ((i_9_) & (n_n482) & (n_n325) & (n_n520) & (!x23x)) + ((i_9_) & (n_n482) & (n_n325) & (n_n520) & (x23x)));
	assign n_n4851 = (((!i_9_) & (n_n524) & (n_n518) & (n_n260)));
	assign n_n1217 = (((!n_n518) & (!x17x) & (!n_n522) & (!n_n4849) & (n_n4851)) + ((!n_n518) & (!x17x) & (!n_n522) & (n_n4849) & (!n_n4851)) + ((!n_n518) & (!x17x) & (!n_n522) & (n_n4849) & (n_n4851)) + ((!n_n518) & (!x17x) & (n_n522) & (!n_n4849) & (n_n4851)) + ((!n_n518) & (!x17x) & (n_n522) & (n_n4849) & (!n_n4851)) + ((!n_n518) & (!x17x) & (n_n522) & (n_n4849) & (n_n4851)) + ((!n_n518) & (x17x) & (!n_n522) & (!n_n4849) & (n_n4851)) + ((!n_n518) & (x17x) & (!n_n522) & (n_n4849) & (!n_n4851)) + ((!n_n518) & (x17x) & (!n_n522) & (n_n4849) & (n_n4851)) + ((!n_n518) & (x17x) & (n_n522) & (!n_n4849) & (n_n4851)) + ((!n_n518) & (x17x) & (n_n522) & (n_n4849) & (!n_n4851)) + ((!n_n518) & (x17x) & (n_n522) & (n_n4849) & (n_n4851)) + ((n_n518) & (!x17x) & (!n_n522) & (!n_n4849) & (n_n4851)) + ((n_n518) & (!x17x) & (!n_n522) & (n_n4849) & (!n_n4851)) + ((n_n518) & (!x17x) & (!n_n522) & (n_n4849) & (n_n4851)) + ((n_n518) & (!x17x) & (n_n522) & (!n_n4849) & (n_n4851)) + ((n_n518) & (!x17x) & (n_n522) & (n_n4849) & (!n_n4851)) + ((n_n518) & (!x17x) & (n_n522) & (n_n4849) & (n_n4851)) + ((n_n518) & (x17x) & (!n_n522) & (!n_n4849) & (n_n4851)) + ((n_n518) & (x17x) & (!n_n522) & (n_n4849) & (!n_n4851)) + ((n_n518) & (x17x) & (!n_n522) & (n_n4849) & (n_n4851)) + ((n_n518) & (x17x) & (n_n522) & (!n_n4849) & (!n_n4851)) + ((n_n518) & (x17x) & (n_n522) & (!n_n4849) & (n_n4851)) + ((n_n518) & (x17x) & (n_n522) & (n_n4849) & (!n_n4851)) + ((n_n518) & (x17x) & (n_n522) & (n_n4849) & (n_n4851)));
	assign n_n4843 = (((!i_9_) & (n_n518) & (n_n532) & (n_n260)));
	assign n_n4846 = (((i_9_) & (n_n518) & (n_n528) & (n_n260)));
	assign n_n4848 = (((i_9_) & (n_n518) & (n_n526) & (n_n260)));
	assign n_n4836 = (((i_9_) & (n_n260) & (n_n535) & (n_n522)));
	assign n_n3460 = (((!i_9_) & (!n_n524) & (n_n260) & (n_n535) & (n_n522)) + ((!i_9_) & (n_n524) & (n_n260) & (n_n535) & (!n_n522)) + ((!i_9_) & (n_n524) & (n_n260) & (n_n535) & (n_n522)) + ((i_9_) & (!n_n524) & (n_n260) & (n_n535) & (n_n522)) + ((i_9_) & (n_n524) & (n_n260) & (n_n535) & (n_n522)));
	assign x11773x = (((!n_n4856) & (!n_n4854) & (!n_n4855) & (!n_n4853) & (n_n4860)) + ((!n_n4856) & (!n_n4854) & (!n_n4855) & (n_n4853) & (!n_n4860)) + ((!n_n4856) & (!n_n4854) & (!n_n4855) & (n_n4853) & (n_n4860)) + ((!n_n4856) & (!n_n4854) & (n_n4855) & (!n_n4853) & (!n_n4860)) + ((!n_n4856) & (!n_n4854) & (n_n4855) & (!n_n4853) & (n_n4860)) + ((!n_n4856) & (!n_n4854) & (n_n4855) & (n_n4853) & (!n_n4860)) + ((!n_n4856) & (!n_n4854) & (n_n4855) & (n_n4853) & (n_n4860)) + ((!n_n4856) & (n_n4854) & (!n_n4855) & (!n_n4853) & (!n_n4860)) + ((!n_n4856) & (n_n4854) & (!n_n4855) & (!n_n4853) & (n_n4860)) + ((!n_n4856) & (n_n4854) & (!n_n4855) & (n_n4853) & (!n_n4860)) + ((!n_n4856) & (n_n4854) & (!n_n4855) & (n_n4853) & (n_n4860)) + ((!n_n4856) & (n_n4854) & (n_n4855) & (!n_n4853) & (!n_n4860)) + ((!n_n4856) & (n_n4854) & (n_n4855) & (!n_n4853) & (n_n4860)) + ((!n_n4856) & (n_n4854) & (n_n4855) & (n_n4853) & (!n_n4860)) + ((!n_n4856) & (n_n4854) & (n_n4855) & (n_n4853) & (n_n4860)) + ((n_n4856) & (!n_n4854) & (!n_n4855) & (!n_n4853) & (!n_n4860)) + ((n_n4856) & (!n_n4854) & (!n_n4855) & (!n_n4853) & (n_n4860)) + ((n_n4856) & (!n_n4854) & (!n_n4855) & (n_n4853) & (!n_n4860)) + ((n_n4856) & (!n_n4854) & (!n_n4855) & (n_n4853) & (n_n4860)) + ((n_n4856) & (!n_n4854) & (n_n4855) & (!n_n4853) & (!n_n4860)) + ((n_n4856) & (!n_n4854) & (n_n4855) & (!n_n4853) & (n_n4860)) + ((n_n4856) & (!n_n4854) & (n_n4855) & (n_n4853) & (!n_n4860)) + ((n_n4856) & (!n_n4854) & (n_n4855) & (n_n4853) & (n_n4860)) + ((n_n4856) & (n_n4854) & (!n_n4855) & (!n_n4853) & (!n_n4860)) + ((n_n4856) & (n_n4854) & (!n_n4855) & (!n_n4853) & (n_n4860)) + ((n_n4856) & (n_n4854) & (!n_n4855) & (n_n4853) & (!n_n4860)) + ((n_n4856) & (n_n4854) & (!n_n4855) & (n_n4853) & (n_n4860)) + ((n_n4856) & (n_n4854) & (n_n4855) & (!n_n4853) & (!n_n4860)) + ((n_n4856) & (n_n4854) & (n_n4855) & (!n_n4853) & (n_n4860)) + ((n_n4856) & (n_n4854) & (n_n4855) & (n_n4853) & (!n_n4860)) + ((n_n4856) & (n_n4854) & (n_n4855) & (n_n4853) & (n_n4860)));
	assign n_n4840 = (((i_9_) & (n_n518) & (n_n534) & (n_n260)));
	assign n_n4838 = (((i_9_) & (n_n260) & (n_n535) & (n_n520)));
	assign n_n3820 = (((!n_n260) & (!n_n535) & (!x23x) & (!n_n4838) & (n_n4840)) + ((!n_n260) & (!n_n535) & (!x23x) & (n_n4838) & (!n_n4840)) + ((!n_n260) & (!n_n535) & (!x23x) & (n_n4838) & (n_n4840)) + ((!n_n260) & (!n_n535) & (x23x) & (!n_n4838) & (n_n4840)) + ((!n_n260) & (!n_n535) & (x23x) & (n_n4838) & (!n_n4840)) + ((!n_n260) & (!n_n535) & (x23x) & (n_n4838) & (n_n4840)) + ((!n_n260) & (n_n535) & (!x23x) & (!n_n4838) & (n_n4840)) + ((!n_n260) & (n_n535) & (!x23x) & (n_n4838) & (!n_n4840)) + ((!n_n260) & (n_n535) & (!x23x) & (n_n4838) & (n_n4840)) + ((!n_n260) & (n_n535) & (x23x) & (!n_n4838) & (n_n4840)) + ((!n_n260) & (n_n535) & (x23x) & (n_n4838) & (!n_n4840)) + ((!n_n260) & (n_n535) & (x23x) & (n_n4838) & (n_n4840)) + ((n_n260) & (!n_n535) & (!x23x) & (!n_n4838) & (n_n4840)) + ((n_n260) & (!n_n535) & (!x23x) & (n_n4838) & (!n_n4840)) + ((n_n260) & (!n_n535) & (!x23x) & (n_n4838) & (n_n4840)) + ((n_n260) & (!n_n535) & (x23x) & (!n_n4838) & (n_n4840)) + ((n_n260) & (!n_n535) & (x23x) & (n_n4838) & (!n_n4840)) + ((n_n260) & (!n_n535) & (x23x) & (n_n4838) & (n_n4840)) + ((n_n260) & (n_n535) & (!x23x) & (!n_n4838) & (n_n4840)) + ((n_n260) & (n_n535) & (!x23x) & (n_n4838) & (!n_n4840)) + ((n_n260) & (n_n535) & (!x23x) & (n_n4838) & (n_n4840)) + ((n_n260) & (n_n535) & (x23x) & (!n_n4838) & (!n_n4840)) + ((n_n260) & (n_n535) & (x23x) & (!n_n4838) & (n_n4840)) + ((n_n260) & (n_n535) & (x23x) & (n_n4838) & (!n_n4840)) + ((n_n260) & (n_n535) & (x23x) & (n_n4838) & (n_n4840)));
	assign n_n4826 = (((i_9_) & (n_n532) & (n_n260) & (n_n535)));
	assign x185x = (((!i_9_) & (!n_n532) & (n_n534) & (n_n260) & (n_n535)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n260) & (n_n535)) + ((i_9_) & (n_n532) & (!n_n534) & (n_n260) & (n_n535)) + ((i_9_) & (n_n532) & (n_n534) & (n_n260) & (n_n535)));
	assign n_n4842 = (((i_9_) & (n_n518) & (n_n532) & (n_n260)));
	assign n_n4841 = (((!i_9_) & (n_n518) & (n_n534) & (n_n260)));
	assign x372x = (((!i_9_) & (n_n518) & (!n_n532) & (n_n534) & (n_n260)) + ((!i_9_) & (n_n518) & (n_n532) & (n_n534) & (n_n260)) + ((i_9_) & (n_n518) & (n_n532) & (!n_n534) & (n_n260)) + ((i_9_) & (n_n518) & (n_n532) & (n_n534) & (n_n260)));
	assign x11780x = (((!n_n4827) & (!n_n4843) & (!n_n4848) & (!x185x) & (x372x)) + ((!n_n4827) & (!n_n4843) & (!n_n4848) & (x185x) & (!x372x)) + ((!n_n4827) & (!n_n4843) & (!n_n4848) & (x185x) & (x372x)) + ((!n_n4827) & (!n_n4843) & (n_n4848) & (!x185x) & (!x372x)) + ((!n_n4827) & (!n_n4843) & (n_n4848) & (!x185x) & (x372x)) + ((!n_n4827) & (!n_n4843) & (n_n4848) & (x185x) & (!x372x)) + ((!n_n4827) & (!n_n4843) & (n_n4848) & (x185x) & (x372x)) + ((!n_n4827) & (n_n4843) & (!n_n4848) & (!x185x) & (!x372x)) + ((!n_n4827) & (n_n4843) & (!n_n4848) & (!x185x) & (x372x)) + ((!n_n4827) & (n_n4843) & (!n_n4848) & (x185x) & (!x372x)) + ((!n_n4827) & (n_n4843) & (!n_n4848) & (x185x) & (x372x)) + ((!n_n4827) & (n_n4843) & (n_n4848) & (!x185x) & (!x372x)) + ((!n_n4827) & (n_n4843) & (n_n4848) & (!x185x) & (x372x)) + ((!n_n4827) & (n_n4843) & (n_n4848) & (x185x) & (!x372x)) + ((!n_n4827) & (n_n4843) & (n_n4848) & (x185x) & (x372x)) + ((n_n4827) & (!n_n4843) & (!n_n4848) & (!x185x) & (!x372x)) + ((n_n4827) & (!n_n4843) & (!n_n4848) & (!x185x) & (x372x)) + ((n_n4827) & (!n_n4843) & (!n_n4848) & (x185x) & (!x372x)) + ((n_n4827) & (!n_n4843) & (!n_n4848) & (x185x) & (x372x)) + ((n_n4827) & (!n_n4843) & (n_n4848) & (!x185x) & (!x372x)) + ((n_n4827) & (!n_n4843) & (n_n4848) & (!x185x) & (x372x)) + ((n_n4827) & (!n_n4843) & (n_n4848) & (x185x) & (!x372x)) + ((n_n4827) & (!n_n4843) & (n_n4848) & (x185x) & (x372x)) + ((n_n4827) & (n_n4843) & (!n_n4848) & (!x185x) & (!x372x)) + ((n_n4827) & (n_n4843) & (!n_n4848) & (!x185x) & (x372x)) + ((n_n4827) & (n_n4843) & (!n_n4848) & (x185x) & (!x372x)) + ((n_n4827) & (n_n4843) & (!n_n4848) & (x185x) & (x372x)) + ((n_n4827) & (n_n4843) & (n_n4848) & (!x185x) & (!x372x)) + ((n_n4827) & (n_n4843) & (n_n4848) & (!x185x) & (x372x)) + ((n_n4827) & (n_n4843) & (n_n4848) & (x185x) & (!x372x)) + ((n_n4827) & (n_n4843) & (n_n4848) & (x185x) & (x372x)));
	assign x11782x = (((!n_n4862) & (!x245x) & (!n_n4861) & (!x11773x) & (x11780x)) + ((!n_n4862) & (!x245x) & (!n_n4861) & (x11773x) & (!x11780x)) + ((!n_n4862) & (!x245x) & (!n_n4861) & (x11773x) & (x11780x)) + ((!n_n4862) & (!x245x) & (n_n4861) & (!x11773x) & (!x11780x)) + ((!n_n4862) & (!x245x) & (n_n4861) & (!x11773x) & (x11780x)) + ((!n_n4862) & (!x245x) & (n_n4861) & (x11773x) & (!x11780x)) + ((!n_n4862) & (!x245x) & (n_n4861) & (x11773x) & (x11780x)) + ((!n_n4862) & (x245x) & (!n_n4861) & (!x11773x) & (!x11780x)) + ((!n_n4862) & (x245x) & (!n_n4861) & (!x11773x) & (x11780x)) + ((!n_n4862) & (x245x) & (!n_n4861) & (x11773x) & (!x11780x)) + ((!n_n4862) & (x245x) & (!n_n4861) & (x11773x) & (x11780x)) + ((!n_n4862) & (x245x) & (n_n4861) & (!x11773x) & (!x11780x)) + ((!n_n4862) & (x245x) & (n_n4861) & (!x11773x) & (x11780x)) + ((!n_n4862) & (x245x) & (n_n4861) & (x11773x) & (!x11780x)) + ((!n_n4862) & (x245x) & (n_n4861) & (x11773x) & (x11780x)) + ((n_n4862) & (!x245x) & (!n_n4861) & (!x11773x) & (!x11780x)) + ((n_n4862) & (!x245x) & (!n_n4861) & (!x11773x) & (x11780x)) + ((n_n4862) & (!x245x) & (!n_n4861) & (x11773x) & (!x11780x)) + ((n_n4862) & (!x245x) & (!n_n4861) & (x11773x) & (x11780x)) + ((n_n4862) & (!x245x) & (n_n4861) & (!x11773x) & (!x11780x)) + ((n_n4862) & (!x245x) & (n_n4861) & (!x11773x) & (x11780x)) + ((n_n4862) & (!x245x) & (n_n4861) & (x11773x) & (!x11780x)) + ((n_n4862) & (!x245x) & (n_n4861) & (x11773x) & (x11780x)) + ((n_n4862) & (x245x) & (!n_n4861) & (!x11773x) & (!x11780x)) + ((n_n4862) & (x245x) & (!n_n4861) & (!x11773x) & (x11780x)) + ((n_n4862) & (x245x) & (!n_n4861) & (x11773x) & (!x11780x)) + ((n_n4862) & (x245x) & (!n_n4861) & (x11773x) & (x11780x)) + ((n_n4862) & (x245x) & (n_n4861) & (!x11773x) & (!x11780x)) + ((n_n4862) & (x245x) & (n_n4861) & (!x11773x) & (x11780x)) + ((n_n4862) & (x245x) & (n_n4861) & (x11773x) & (!x11780x)) + ((n_n4862) & (x245x) & (n_n4861) & (x11773x) & (x11780x)));
	assign x11778x = (((!n_n4849) & (!n_n4852) & (!n_n4845) & (!n_n4846) & (n_n4851)) + ((!n_n4849) & (!n_n4852) & (!n_n4845) & (n_n4846) & (!n_n4851)) + ((!n_n4849) & (!n_n4852) & (!n_n4845) & (n_n4846) & (n_n4851)) + ((!n_n4849) & (!n_n4852) & (n_n4845) & (!n_n4846) & (!n_n4851)) + ((!n_n4849) & (!n_n4852) & (n_n4845) & (!n_n4846) & (n_n4851)) + ((!n_n4849) & (!n_n4852) & (n_n4845) & (n_n4846) & (!n_n4851)) + ((!n_n4849) & (!n_n4852) & (n_n4845) & (n_n4846) & (n_n4851)) + ((!n_n4849) & (n_n4852) & (!n_n4845) & (!n_n4846) & (!n_n4851)) + ((!n_n4849) & (n_n4852) & (!n_n4845) & (!n_n4846) & (n_n4851)) + ((!n_n4849) & (n_n4852) & (!n_n4845) & (n_n4846) & (!n_n4851)) + ((!n_n4849) & (n_n4852) & (!n_n4845) & (n_n4846) & (n_n4851)) + ((!n_n4849) & (n_n4852) & (n_n4845) & (!n_n4846) & (!n_n4851)) + ((!n_n4849) & (n_n4852) & (n_n4845) & (!n_n4846) & (n_n4851)) + ((!n_n4849) & (n_n4852) & (n_n4845) & (n_n4846) & (!n_n4851)) + ((!n_n4849) & (n_n4852) & (n_n4845) & (n_n4846) & (n_n4851)) + ((n_n4849) & (!n_n4852) & (!n_n4845) & (!n_n4846) & (!n_n4851)) + ((n_n4849) & (!n_n4852) & (!n_n4845) & (!n_n4846) & (n_n4851)) + ((n_n4849) & (!n_n4852) & (!n_n4845) & (n_n4846) & (!n_n4851)) + ((n_n4849) & (!n_n4852) & (!n_n4845) & (n_n4846) & (n_n4851)) + ((n_n4849) & (!n_n4852) & (n_n4845) & (!n_n4846) & (!n_n4851)) + ((n_n4849) & (!n_n4852) & (n_n4845) & (!n_n4846) & (n_n4851)) + ((n_n4849) & (!n_n4852) & (n_n4845) & (n_n4846) & (!n_n4851)) + ((n_n4849) & (!n_n4852) & (n_n4845) & (n_n4846) & (n_n4851)) + ((n_n4849) & (n_n4852) & (!n_n4845) & (!n_n4846) & (!n_n4851)) + ((n_n4849) & (n_n4852) & (!n_n4845) & (!n_n4846) & (n_n4851)) + ((n_n4849) & (n_n4852) & (!n_n4845) & (n_n4846) & (!n_n4851)) + ((n_n4849) & (n_n4852) & (!n_n4845) & (n_n4846) & (n_n4851)) + ((n_n4849) & (n_n4852) & (n_n4845) & (!n_n4846) & (!n_n4851)) + ((n_n4849) & (n_n4852) & (n_n4845) & (!n_n4846) & (n_n4851)) + ((n_n4849) & (n_n4852) & (n_n4845) & (n_n4846) & (!n_n4851)) + ((n_n4849) & (n_n4852) & (n_n4845) & (n_n4846) & (n_n4851)));
	assign n_n4390 = (((i_9_) & (n_n536) & (n_n491) & (n_n520)));
	assign n_n4633 = (((!i_9_) & (n_n390) & (n_n534) & (n_n491)));
	assign n_n5155 = (((!i_9_) & (n_n524) & (n_n491) & (n_n130)));
	assign n_n5161 = (((!i_9_) & (n_n482) & (n_n534) & (n_n130)));
	assign n_n4482 = (((i_9_) & (n_n524) & (n_n455) & (n_n509)));
	assign n_n4489 = (((!i_9_) & (n_n455) & (n_n534) & (n_n500)));
	assign n_n4504 = (((i_9_) & (n_n455) & (n_n534) & (n_n491)));
	assign n_n4526 = (((i_9_) & (n_n482) & (n_n455) & (n_n528)));
	assign n_n4554 = (((i_9_) & (n_n455) & (n_n532) & (n_n464)));
	assign n_n4561 = (((!i_9_) & (n_n526) & (n_n455) & (n_n464)));
	assign n_n4568 = (((i_9_) & (n_n390) & (n_n534) & (n_n535)));
	assign n_n4575 = (((!i_9_) & (n_n528) & (n_n390) & (n_n535)));
	assign n_n4590 = (((i_9_) & (n_n518) & (n_n528) & (n_n390)));
	assign n_n4690 = (((i_9_) & (n_n524) & (n_n390) & (n_n464)));
	assign n_n4704 = (((i_9_) & (n_n526) & (n_n325) & (n_n535)));
	assign n_n4711 = (((!i_1_) & (!i_2_) & (i_0_) & (n_n535) & (x23x)));
	assign n_n4974 = (((i_9_) & (n_n518) & (n_n528) & (n_n195)));
	assign n_n5047 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n195) & (x23x)));
	assign n_n5098 = (((!i_5_) & (i_3_) & (i_4_) & (n_n532) & (x12x)));
	assign n_n5105 = (((!i_9_) & (n_n518) & (n_n526) & (n_n130)));
	assign n_n5120 = (((i_7_) & (i_8_) & (!i_6_) & (n_n509) & (x12x)));
	assign n_n5127 = (((i_5_) & (i_3_) & (!i_4_) & (n_n130) & (x23x)));
	assign n_n5164 = (((!i_5_) & (!i_3_) & (i_4_) & (x12x) & (n_n530)));
	assign n_n5193 = (((!i_9_) & (n_n534) & (n_n130) & (n_n464)));
	assign n_n5251 = (((!i_9_) & (n_n524) & (n_n509) & (n_n65)));
	assign n_n5266 = (((i_7_) & (!i_8_) & (!i_6_) & (x19x) & (n_n500)));
	assign n_n5273 = (((!i_9_) & (n_n534) & (n_n491) & (n_n65)));
	assign n_n4398 = (((i_9_) & (n_n536) & (n_n482) & (n_n528)));
	assign n_n4524 = (((i_9_) & (n_n482) & (n_n455) & (n_n530)));
	assign n_n4522 = (((i_9_) & (n_n482) & (n_n455) & (n_n532)));
	assign x170x = (((!i_9_) & (n_n482) & (n_n455) & (n_n532)) + ((i_9_) & (n_n482) & (n_n455) & (n_n532)));
	assign n_n4246 = (((!i_9_) & (n_n482) & (n_n455) & (n_n532) & (!n_n530)) + ((!i_9_) & (n_n482) & (n_n455) & (n_n532) & (n_n530)) + ((i_9_) & (n_n482) & (n_n455) & (!n_n532) & (n_n530)) + ((i_9_) & (n_n482) & (n_n455) & (n_n532) & (!n_n530)) + ((i_9_) & (n_n482) & (n_n455) & (n_n532) & (n_n530)));
	assign n_n4670 = (((i_9_) & (n_n528) & (n_n390) & (n_n473)));
	assign n_n4732 = (((i_9_) & (n_n509) & (n_n325) & (n_n530)));
	assign n_n5086 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n535) & (x12x)));
	assign n_n5087 = (((!i_9_) & (n_n528) & (n_n535) & (n_n130)));
	assign n_n4587 = (((!i_9_) & (n_n518) & (n_n390) & (n_n532)));
	assign n_n881 = (((!x15x) & (!n_n518) & (!n_n390) & (!x24x) & (n_n4590)) + ((!x15x) & (!n_n518) & (!n_n390) & (x24x) & (n_n4590)) + ((!x15x) & (!n_n518) & (n_n390) & (!x24x) & (n_n4590)) + ((!x15x) & (!n_n518) & (n_n390) & (x24x) & (n_n4590)) + ((!x15x) & (n_n518) & (!n_n390) & (!x24x) & (n_n4590)) + ((!x15x) & (n_n518) & (!n_n390) & (x24x) & (n_n4590)) + ((!x15x) & (n_n518) & (n_n390) & (!x24x) & (n_n4590)) + ((!x15x) & (n_n518) & (n_n390) & (x24x) & (!n_n4590)) + ((!x15x) & (n_n518) & (n_n390) & (x24x) & (n_n4590)) + ((x15x) & (!n_n518) & (!n_n390) & (!x24x) & (n_n4590)) + ((x15x) & (!n_n518) & (!n_n390) & (x24x) & (n_n4590)) + ((x15x) & (!n_n518) & (n_n390) & (!x24x) & (n_n4590)) + ((x15x) & (!n_n518) & (n_n390) & (x24x) & (n_n4590)) + ((x15x) & (n_n518) & (!n_n390) & (!x24x) & (n_n4590)) + ((x15x) & (n_n518) & (!n_n390) & (x24x) & (n_n4590)) + ((x15x) & (n_n518) & (n_n390) & (!x24x) & (!n_n4590)) + ((x15x) & (n_n518) & (n_n390) & (!x24x) & (n_n4590)) + ((x15x) & (n_n518) & (n_n390) & (x24x) & (!n_n4590)) + ((x15x) & (n_n518) & (n_n390) & (x24x) & (n_n4590)));
	assign n_n4594 = (((i_9_) & (n_n524) & (n_n518) & (n_n390)));
	assign n_n4591 = (((!i_9_) & (n_n518) & (n_n528) & (n_n390)));
	assign n_n4592 = (((i_9_) & (n_n518) & (n_n526) & (n_n390)));
	assign x172x = (((!i_9_) & (n_n518) & (!n_n526) & (n_n528) & (n_n390)) + ((!i_9_) & (n_n518) & (n_n526) & (n_n528) & (n_n390)) + ((i_9_) & (n_n518) & (n_n526) & (!n_n528) & (n_n390)) + ((i_9_) & (n_n518) & (n_n526) & (n_n528) & (n_n390)));
	assign n_n4083 = (((!n_n4593) & (!x257x) & (!n_n881) & (!n_n4594) & (x172x)) + ((!n_n4593) & (!x257x) & (!n_n881) & (n_n4594) & (!x172x)) + ((!n_n4593) & (!x257x) & (!n_n881) & (n_n4594) & (x172x)) + ((!n_n4593) & (!x257x) & (n_n881) & (!n_n4594) & (!x172x)) + ((!n_n4593) & (!x257x) & (n_n881) & (!n_n4594) & (x172x)) + ((!n_n4593) & (!x257x) & (n_n881) & (n_n4594) & (!x172x)) + ((!n_n4593) & (!x257x) & (n_n881) & (n_n4594) & (x172x)) + ((!n_n4593) & (x257x) & (!n_n881) & (!n_n4594) & (!x172x)) + ((!n_n4593) & (x257x) & (!n_n881) & (!n_n4594) & (x172x)) + ((!n_n4593) & (x257x) & (!n_n881) & (n_n4594) & (!x172x)) + ((!n_n4593) & (x257x) & (!n_n881) & (n_n4594) & (x172x)) + ((!n_n4593) & (x257x) & (n_n881) & (!n_n4594) & (!x172x)) + ((!n_n4593) & (x257x) & (n_n881) & (!n_n4594) & (x172x)) + ((!n_n4593) & (x257x) & (n_n881) & (n_n4594) & (!x172x)) + ((!n_n4593) & (x257x) & (n_n881) & (n_n4594) & (x172x)) + ((n_n4593) & (!x257x) & (!n_n881) & (!n_n4594) & (!x172x)) + ((n_n4593) & (!x257x) & (!n_n881) & (!n_n4594) & (x172x)) + ((n_n4593) & (!x257x) & (!n_n881) & (n_n4594) & (!x172x)) + ((n_n4593) & (!x257x) & (!n_n881) & (n_n4594) & (x172x)) + ((n_n4593) & (!x257x) & (n_n881) & (!n_n4594) & (!x172x)) + ((n_n4593) & (!x257x) & (n_n881) & (!n_n4594) & (x172x)) + ((n_n4593) & (!x257x) & (n_n881) & (n_n4594) & (!x172x)) + ((n_n4593) & (!x257x) & (n_n881) & (n_n4594) & (x172x)) + ((n_n4593) & (x257x) & (!n_n881) & (!n_n4594) & (!x172x)) + ((n_n4593) & (x257x) & (!n_n881) & (!n_n4594) & (x172x)) + ((n_n4593) & (x257x) & (!n_n881) & (n_n4594) & (!x172x)) + ((n_n4593) & (x257x) & (!n_n881) & (n_n4594) & (x172x)) + ((n_n4593) & (x257x) & (n_n881) & (!n_n4594) & (!x172x)) + ((n_n4593) & (x257x) & (n_n881) & (!n_n4594) & (x172x)) + ((n_n4593) & (x257x) & (n_n881) & (n_n4594) & (!x172x)) + ((n_n4593) & (x257x) & (n_n881) & (n_n4594) & (x172x)));
	assign n_n4452 = (((i_9_) & (n_n455) & (n_n535) & (n_n522)));
	assign n_n3520 = (((!i_9_) & (!n_n524) & (n_n455) & (n_n535) & (n_n522)) + ((!i_9_) & (n_n524) & (n_n455) & (n_n535) & (!n_n522)) + ((!i_9_) & (n_n524) & (n_n455) & (n_n535) & (n_n522)) + ((i_9_) & (!n_n524) & (n_n455) & (n_n535) & (n_n522)) + ((i_9_) & (n_n524) & (n_n455) & (n_n535) & (n_n522)));
	assign n_n4919 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n260) & (x23x)));
	assign n_n4984 = (((i_9_) & (n_n534) & (n_n509) & (n_n195)));
	assign n_n5162 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n532) & (x12x)));
	assign n_n4582 = (((i_9_) & (n_n390) & (n_n535) & (n_n520)));
	assign n_n4584 = (((i_9_) & (n_n518) & (n_n390) & (n_n534)));
	assign n_n4586 = (((i_9_) & (n_n518) & (n_n390) & (n_n532)));
	assign n_n4588 = (((i_9_) & (n_n518) & (n_n390) & (n_n530)));
	assign x365x = (((!i_9_) & (n_n518) & (n_n390) & (n_n530)) + ((i_9_) & (n_n518) & (n_n390) & (n_n530)));
	assign x14093x = (((!n_n4591) & (!n_n4592) & (!n_n4582) & (!n_n4584) & (n_n4586)) + ((!n_n4591) & (!n_n4592) & (!n_n4582) & (n_n4584) & (!n_n4586)) + ((!n_n4591) & (!n_n4592) & (!n_n4582) & (n_n4584) & (n_n4586)) + ((!n_n4591) & (!n_n4592) & (n_n4582) & (!n_n4584) & (!n_n4586)) + ((!n_n4591) & (!n_n4592) & (n_n4582) & (!n_n4584) & (n_n4586)) + ((!n_n4591) & (!n_n4592) & (n_n4582) & (n_n4584) & (!n_n4586)) + ((!n_n4591) & (!n_n4592) & (n_n4582) & (n_n4584) & (n_n4586)) + ((!n_n4591) & (n_n4592) & (!n_n4582) & (!n_n4584) & (!n_n4586)) + ((!n_n4591) & (n_n4592) & (!n_n4582) & (!n_n4584) & (n_n4586)) + ((!n_n4591) & (n_n4592) & (!n_n4582) & (n_n4584) & (!n_n4586)) + ((!n_n4591) & (n_n4592) & (!n_n4582) & (n_n4584) & (n_n4586)) + ((!n_n4591) & (n_n4592) & (n_n4582) & (!n_n4584) & (!n_n4586)) + ((!n_n4591) & (n_n4592) & (n_n4582) & (!n_n4584) & (n_n4586)) + ((!n_n4591) & (n_n4592) & (n_n4582) & (n_n4584) & (!n_n4586)) + ((!n_n4591) & (n_n4592) & (n_n4582) & (n_n4584) & (n_n4586)) + ((n_n4591) & (!n_n4592) & (!n_n4582) & (!n_n4584) & (!n_n4586)) + ((n_n4591) & (!n_n4592) & (!n_n4582) & (!n_n4584) & (n_n4586)) + ((n_n4591) & (!n_n4592) & (!n_n4582) & (n_n4584) & (!n_n4586)) + ((n_n4591) & (!n_n4592) & (!n_n4582) & (n_n4584) & (n_n4586)) + ((n_n4591) & (!n_n4592) & (n_n4582) & (!n_n4584) & (!n_n4586)) + ((n_n4591) & (!n_n4592) & (n_n4582) & (!n_n4584) & (n_n4586)) + ((n_n4591) & (!n_n4592) & (n_n4582) & (n_n4584) & (!n_n4586)) + ((n_n4591) & (!n_n4592) & (n_n4582) & (n_n4584) & (n_n4586)) + ((n_n4591) & (n_n4592) & (!n_n4582) & (!n_n4584) & (!n_n4586)) + ((n_n4591) & (n_n4592) & (!n_n4582) & (!n_n4584) & (n_n4586)) + ((n_n4591) & (n_n4592) & (!n_n4582) & (n_n4584) & (!n_n4586)) + ((n_n4591) & (n_n4592) & (!n_n4582) & (n_n4584) & (n_n4586)) + ((n_n4591) & (n_n4592) & (n_n4582) & (!n_n4584) & (!n_n4586)) + ((n_n4591) & (n_n4592) & (n_n4582) & (!n_n4584) & (n_n4586)) + ((n_n4591) & (n_n4592) & (n_n4582) & (n_n4584) & (!n_n4586)) + ((n_n4591) & (n_n4592) & (n_n4582) & (n_n4584) & (n_n4586)));
	assign n_n3348 = (((!n_n4590) & (!n_n4587) & (!x365x) & (x14093x)) + ((!n_n4590) & (!n_n4587) & (x365x) & (!x14093x)) + ((!n_n4590) & (!n_n4587) & (x365x) & (x14093x)) + ((!n_n4590) & (n_n4587) & (!x365x) & (!x14093x)) + ((!n_n4590) & (n_n4587) & (!x365x) & (x14093x)) + ((!n_n4590) & (n_n4587) & (x365x) & (!x14093x)) + ((!n_n4590) & (n_n4587) & (x365x) & (x14093x)) + ((n_n4590) & (!n_n4587) & (!x365x) & (!x14093x)) + ((n_n4590) & (!n_n4587) & (!x365x) & (x14093x)) + ((n_n4590) & (!n_n4587) & (x365x) & (!x14093x)) + ((n_n4590) & (!n_n4587) & (x365x) & (x14093x)) + ((n_n4590) & (n_n4587) & (!x365x) & (!x14093x)) + ((n_n4590) & (n_n4587) & (!x365x) & (x14093x)) + ((n_n4590) & (n_n4587) & (x365x) & (!x14093x)) + ((n_n4590) & (n_n4587) & (x365x) & (x14093x)));
	assign n_n4876 = (((i_9_) & (n_n260) & (n_n500) & (n_n530)));
	assign x461x = (((!n_n509) & (!x17x) & (!n_n520) & (!n_n4872) & (n_n4871)) + ((!n_n509) & (!x17x) & (!n_n520) & (n_n4872) & (!n_n4871)) + ((!n_n509) & (!x17x) & (!n_n520) & (n_n4872) & (n_n4871)) + ((!n_n509) & (!x17x) & (n_n520) & (!n_n4872) & (n_n4871)) + ((!n_n509) & (!x17x) & (n_n520) & (n_n4872) & (!n_n4871)) + ((!n_n509) & (!x17x) & (n_n520) & (n_n4872) & (n_n4871)) + ((!n_n509) & (x17x) & (!n_n520) & (!n_n4872) & (n_n4871)) + ((!n_n509) & (x17x) & (!n_n520) & (n_n4872) & (!n_n4871)) + ((!n_n509) & (x17x) & (!n_n520) & (n_n4872) & (n_n4871)) + ((!n_n509) & (x17x) & (n_n520) & (!n_n4872) & (n_n4871)) + ((!n_n509) & (x17x) & (n_n520) & (n_n4872) & (!n_n4871)) + ((!n_n509) & (x17x) & (n_n520) & (n_n4872) & (n_n4871)) + ((n_n509) & (!x17x) & (!n_n520) & (!n_n4872) & (n_n4871)) + ((n_n509) & (!x17x) & (!n_n520) & (n_n4872) & (!n_n4871)) + ((n_n509) & (!x17x) & (!n_n520) & (n_n4872) & (n_n4871)) + ((n_n509) & (!x17x) & (n_n520) & (!n_n4872) & (n_n4871)) + ((n_n509) & (!x17x) & (n_n520) & (n_n4872) & (!n_n4871)) + ((n_n509) & (!x17x) & (n_n520) & (n_n4872) & (n_n4871)) + ((n_n509) & (x17x) & (!n_n520) & (!n_n4872) & (n_n4871)) + ((n_n509) & (x17x) & (!n_n520) & (n_n4872) & (!n_n4871)) + ((n_n509) & (x17x) & (!n_n520) & (n_n4872) & (n_n4871)) + ((n_n509) & (x17x) & (n_n520) & (!n_n4872) & (!n_n4871)) + ((n_n509) & (x17x) & (n_n520) & (!n_n4872) & (n_n4871)) + ((n_n509) & (x17x) & (n_n520) & (n_n4872) & (!n_n4871)) + ((n_n509) & (x17x) & (n_n520) & (n_n4872) & (n_n4871)));
	assign x22120x = (((!n_n4881) & (!n_n4878) & (!n_n4880) & (!n_n4877)));
	assign n_n3326 = (((!n_n4879) & (!n_n4876) & (!x461x) & (!x22120x)) + ((!n_n4879) & (!n_n4876) & (x461x) & (!x22120x)) + ((!n_n4879) & (!n_n4876) & (x461x) & (x22120x)) + ((!n_n4879) & (n_n4876) & (!x461x) & (!x22120x)) + ((!n_n4879) & (n_n4876) & (!x461x) & (x22120x)) + ((!n_n4879) & (n_n4876) & (x461x) & (!x22120x)) + ((!n_n4879) & (n_n4876) & (x461x) & (x22120x)) + ((n_n4879) & (!n_n4876) & (!x461x) & (!x22120x)) + ((n_n4879) & (!n_n4876) & (!x461x) & (x22120x)) + ((n_n4879) & (!n_n4876) & (x461x) & (!x22120x)) + ((n_n4879) & (!n_n4876) & (x461x) & (x22120x)) + ((n_n4879) & (n_n4876) & (!x461x) & (!x22120x)) + ((n_n4879) & (n_n4876) & (!x461x) & (x22120x)) + ((n_n4879) & (n_n4876) & (x461x) & (!x22120x)) + ((n_n4879) & (n_n4876) & (x461x) & (x22120x)));
	assign n_n5327 = (((!i_9_) & (n_n528) & (n_n464) & (n_n65)));
	assign n_n2643 = (((!i_9_) & (!n_n528) & (n_n530) & (n_n464) & (n_n65)) + ((!i_9_) & (n_n528) & (!n_n530) & (n_n464) & (n_n65)) + ((!i_9_) & (n_n528) & (n_n530) & (n_n464) & (n_n65)) + ((i_9_) & (n_n528) & (!n_n530) & (n_n464) & (n_n65)) + ((i_9_) & (n_n528) & (n_n530) & (n_n464) & (n_n65)));
	assign n_n5323 = (((!i_9_) & (n_n532) & (n_n464) & (n_n65)));
	assign n_n4577 = (((!i_9_) & (n_n526) & (n_n390) & (n_n535)));
	assign n_n4576 = (((i_9_) & (n_n526) & (n_n390) & (n_n535)));
	assign n_n4569 = (((!i_9_) & (n_n390) & (n_n534) & (n_n535)));
	assign n_n4573 = (((!i_9_) & (n_n390) & (n_n535) & (n_n530)));
	assign n_n4579 = (((!i_9_) & (n_n524) & (n_n390) & (n_n535)));
	assign x14100x = (((!n_n4575) & (!n_n4577) & (!n_n4572) & (!n_n4573) & (n_n4579)) + ((!n_n4575) & (!n_n4577) & (!n_n4572) & (n_n4573) & (!n_n4579)) + ((!n_n4575) & (!n_n4577) & (!n_n4572) & (n_n4573) & (n_n4579)) + ((!n_n4575) & (!n_n4577) & (n_n4572) & (!n_n4573) & (!n_n4579)) + ((!n_n4575) & (!n_n4577) & (n_n4572) & (!n_n4573) & (n_n4579)) + ((!n_n4575) & (!n_n4577) & (n_n4572) & (n_n4573) & (!n_n4579)) + ((!n_n4575) & (!n_n4577) & (n_n4572) & (n_n4573) & (n_n4579)) + ((!n_n4575) & (n_n4577) & (!n_n4572) & (!n_n4573) & (!n_n4579)) + ((!n_n4575) & (n_n4577) & (!n_n4572) & (!n_n4573) & (n_n4579)) + ((!n_n4575) & (n_n4577) & (!n_n4572) & (n_n4573) & (!n_n4579)) + ((!n_n4575) & (n_n4577) & (!n_n4572) & (n_n4573) & (n_n4579)) + ((!n_n4575) & (n_n4577) & (n_n4572) & (!n_n4573) & (!n_n4579)) + ((!n_n4575) & (n_n4577) & (n_n4572) & (!n_n4573) & (n_n4579)) + ((!n_n4575) & (n_n4577) & (n_n4572) & (n_n4573) & (!n_n4579)) + ((!n_n4575) & (n_n4577) & (n_n4572) & (n_n4573) & (n_n4579)) + ((n_n4575) & (!n_n4577) & (!n_n4572) & (!n_n4573) & (!n_n4579)) + ((n_n4575) & (!n_n4577) & (!n_n4572) & (!n_n4573) & (n_n4579)) + ((n_n4575) & (!n_n4577) & (!n_n4572) & (n_n4573) & (!n_n4579)) + ((n_n4575) & (!n_n4577) & (!n_n4572) & (n_n4573) & (n_n4579)) + ((n_n4575) & (!n_n4577) & (n_n4572) & (!n_n4573) & (!n_n4579)) + ((n_n4575) & (!n_n4577) & (n_n4572) & (!n_n4573) & (n_n4579)) + ((n_n4575) & (!n_n4577) & (n_n4572) & (n_n4573) & (!n_n4579)) + ((n_n4575) & (!n_n4577) & (n_n4572) & (n_n4573) & (n_n4579)) + ((n_n4575) & (n_n4577) & (!n_n4572) & (!n_n4573) & (!n_n4579)) + ((n_n4575) & (n_n4577) & (!n_n4572) & (!n_n4573) & (n_n4579)) + ((n_n4575) & (n_n4577) & (!n_n4572) & (n_n4573) & (!n_n4579)) + ((n_n4575) & (n_n4577) & (!n_n4572) & (n_n4573) & (n_n4579)) + ((n_n4575) & (n_n4577) & (n_n4572) & (!n_n4573) & (!n_n4579)) + ((n_n4575) & (n_n4577) & (n_n4572) & (!n_n4573) & (n_n4579)) + ((n_n4575) & (n_n4577) & (n_n4572) & (n_n4573) & (!n_n4579)) + ((n_n4575) & (n_n4577) & (n_n4572) & (n_n4573) & (n_n4579)));
	assign x14101x = (((!n_n4576) & (!n_n4569) & (!n_n4574) & (!n_n4581) & (x14100x)) + ((!n_n4576) & (!n_n4569) & (!n_n4574) & (n_n4581) & (!x14100x)) + ((!n_n4576) & (!n_n4569) & (!n_n4574) & (n_n4581) & (x14100x)) + ((!n_n4576) & (!n_n4569) & (n_n4574) & (!n_n4581) & (!x14100x)) + ((!n_n4576) & (!n_n4569) & (n_n4574) & (!n_n4581) & (x14100x)) + ((!n_n4576) & (!n_n4569) & (n_n4574) & (n_n4581) & (!x14100x)) + ((!n_n4576) & (!n_n4569) & (n_n4574) & (n_n4581) & (x14100x)) + ((!n_n4576) & (n_n4569) & (!n_n4574) & (!n_n4581) & (!x14100x)) + ((!n_n4576) & (n_n4569) & (!n_n4574) & (!n_n4581) & (x14100x)) + ((!n_n4576) & (n_n4569) & (!n_n4574) & (n_n4581) & (!x14100x)) + ((!n_n4576) & (n_n4569) & (!n_n4574) & (n_n4581) & (x14100x)) + ((!n_n4576) & (n_n4569) & (n_n4574) & (!n_n4581) & (!x14100x)) + ((!n_n4576) & (n_n4569) & (n_n4574) & (!n_n4581) & (x14100x)) + ((!n_n4576) & (n_n4569) & (n_n4574) & (n_n4581) & (!x14100x)) + ((!n_n4576) & (n_n4569) & (n_n4574) & (n_n4581) & (x14100x)) + ((n_n4576) & (!n_n4569) & (!n_n4574) & (!n_n4581) & (!x14100x)) + ((n_n4576) & (!n_n4569) & (!n_n4574) & (!n_n4581) & (x14100x)) + ((n_n4576) & (!n_n4569) & (!n_n4574) & (n_n4581) & (!x14100x)) + ((n_n4576) & (!n_n4569) & (!n_n4574) & (n_n4581) & (x14100x)) + ((n_n4576) & (!n_n4569) & (n_n4574) & (!n_n4581) & (!x14100x)) + ((n_n4576) & (!n_n4569) & (n_n4574) & (!n_n4581) & (x14100x)) + ((n_n4576) & (!n_n4569) & (n_n4574) & (n_n4581) & (!x14100x)) + ((n_n4576) & (!n_n4569) & (n_n4574) & (n_n4581) & (x14100x)) + ((n_n4576) & (n_n4569) & (!n_n4574) & (!n_n4581) & (!x14100x)) + ((n_n4576) & (n_n4569) & (!n_n4574) & (!n_n4581) & (x14100x)) + ((n_n4576) & (n_n4569) & (!n_n4574) & (n_n4581) & (!x14100x)) + ((n_n4576) & (n_n4569) & (!n_n4574) & (n_n4581) & (x14100x)) + ((n_n4576) & (n_n4569) & (n_n4574) & (!n_n4581) & (!x14100x)) + ((n_n4576) & (n_n4569) & (n_n4574) & (!n_n4581) & (x14100x)) + ((n_n4576) & (n_n4569) & (n_n4574) & (n_n4581) & (!x14100x)) + ((n_n4576) & (n_n4569) & (n_n4574) & (n_n4581) & (x14100x)));
	assign n_n4538 = (((i_9_) & (n_n455) & (n_n473) & (n_n532)));
	assign n_n4542 = (((i_9_) & (n_n455) & (n_n528) & (n_n473)));
	assign x201x = (((!i_9_) & (n_n455) & (n_n473) & (n_n530)) + ((i_9_) & (n_n455) & (n_n473) & (n_n530)));
	assign n_n3504 = (((!i_9_) & (n_n455) & (!n_n528) & (n_n473) & (n_n530)) + ((!i_9_) & (n_n455) & (n_n528) & (n_n473) & (n_n530)) + ((i_9_) & (n_n455) & (!n_n528) & (n_n473) & (n_n530)) + ((i_9_) & (n_n455) & (n_n528) & (n_n473) & (!n_n530)) + ((i_9_) & (n_n455) & (n_n528) & (n_n473) & (n_n530)));
	assign n_n4531 = (((!i_9_) & (n_n524) & (n_n482) & (n_n455)));
	assign n_n4551 = (((i_1_) & (!i_2_) & (i_0_) & (n_n473) & (x23x)));
	assign n_n3871 = (((!i_9_) & (!n_n455) & (!n_n534) & (!n_n464) & (n_n4551)) + ((!i_9_) & (!n_n455) & (!n_n534) & (n_n464) & (n_n4551)) + ((!i_9_) & (!n_n455) & (n_n534) & (!n_n464) & (n_n4551)) + ((!i_9_) & (!n_n455) & (n_n534) & (n_n464) & (n_n4551)) + ((!i_9_) & (n_n455) & (!n_n534) & (!n_n464) & (n_n4551)) + ((!i_9_) & (n_n455) & (!n_n534) & (n_n464) & (n_n4551)) + ((!i_9_) & (n_n455) & (n_n534) & (!n_n464) & (n_n4551)) + ((!i_9_) & (n_n455) & (n_n534) & (n_n464) & (!n_n4551)) + ((!i_9_) & (n_n455) & (n_n534) & (n_n464) & (n_n4551)) + ((i_9_) & (!n_n455) & (!n_n534) & (!n_n464) & (n_n4551)) + ((i_9_) & (!n_n455) & (!n_n534) & (n_n464) & (n_n4551)) + ((i_9_) & (!n_n455) & (n_n534) & (!n_n464) & (n_n4551)) + ((i_9_) & (!n_n455) & (n_n534) & (n_n464) & (n_n4551)) + ((i_9_) & (n_n455) & (!n_n534) & (!n_n464) & (n_n4551)) + ((i_9_) & (n_n455) & (!n_n534) & (n_n464) & (n_n4551)) + ((i_9_) & (n_n455) & (n_n534) & (!n_n464) & (n_n4551)) + ((i_9_) & (n_n455) & (n_n534) & (n_n464) & (!n_n4551)) + ((i_9_) & (n_n455) & (n_n534) & (n_n464) & (n_n4551)));
	assign x213x = (((!i_9_) & (n_n455) & (n_n528) & (n_n464)) + ((i_9_) & (n_n455) & (n_n528) & (n_n464)));
	assign n_n4556 = (((i_9_) & (n_n455) & (n_n530) & (n_n464)));
	assign x430x = (((!i_9_) & (n_n455) & (n_n532) & (n_n464)) + ((i_9_) & (n_n455) & (n_n532) & (n_n464)));
	assign x222x = (((!n_n455) & (!x23x) & (!n_n464) & (n_n4568)) + ((!n_n455) & (!x23x) & (n_n464) & (n_n4568)) + ((!n_n455) & (x23x) & (!n_n464) & (n_n4568)) + ((!n_n455) & (x23x) & (n_n464) & (n_n4568)) + ((n_n455) & (!x23x) & (!n_n464) & (n_n4568)) + ((n_n455) & (!x23x) & (n_n464) & (n_n4568)) + ((n_n455) & (x23x) & (!n_n464) & (n_n4568)) + ((n_n455) & (x23x) & (n_n464) & (!n_n4568)) + ((n_n455) & (x23x) & (n_n464) & (n_n4568)));
	assign x14103x = (((!i_9_) & (n_n526) & (n_n455) & (n_n464)) + ((i_9_) & (n_n526) & (n_n455) & (n_n464)));
	assign n_n3350 = (((!x213x) & (!n_n4556) & (!x430x) & (!x222x) & (x14103x)) + ((!x213x) & (!n_n4556) & (!x430x) & (x222x) & (!x14103x)) + ((!x213x) & (!n_n4556) & (!x430x) & (x222x) & (x14103x)) + ((!x213x) & (!n_n4556) & (x430x) & (!x222x) & (!x14103x)) + ((!x213x) & (!n_n4556) & (x430x) & (!x222x) & (x14103x)) + ((!x213x) & (!n_n4556) & (x430x) & (x222x) & (!x14103x)) + ((!x213x) & (!n_n4556) & (x430x) & (x222x) & (x14103x)) + ((!x213x) & (n_n4556) & (!x430x) & (!x222x) & (!x14103x)) + ((!x213x) & (n_n4556) & (!x430x) & (!x222x) & (x14103x)) + ((!x213x) & (n_n4556) & (!x430x) & (x222x) & (!x14103x)) + ((!x213x) & (n_n4556) & (!x430x) & (x222x) & (x14103x)) + ((!x213x) & (n_n4556) & (x430x) & (!x222x) & (!x14103x)) + ((!x213x) & (n_n4556) & (x430x) & (!x222x) & (x14103x)) + ((!x213x) & (n_n4556) & (x430x) & (x222x) & (!x14103x)) + ((!x213x) & (n_n4556) & (x430x) & (x222x) & (x14103x)) + ((x213x) & (!n_n4556) & (!x430x) & (!x222x) & (!x14103x)) + ((x213x) & (!n_n4556) & (!x430x) & (!x222x) & (x14103x)) + ((x213x) & (!n_n4556) & (!x430x) & (x222x) & (!x14103x)) + ((x213x) & (!n_n4556) & (!x430x) & (x222x) & (x14103x)) + ((x213x) & (!n_n4556) & (x430x) & (!x222x) & (!x14103x)) + ((x213x) & (!n_n4556) & (x430x) & (!x222x) & (x14103x)) + ((x213x) & (!n_n4556) & (x430x) & (x222x) & (!x14103x)) + ((x213x) & (!n_n4556) & (x430x) & (x222x) & (x14103x)) + ((x213x) & (n_n4556) & (!x430x) & (!x222x) & (!x14103x)) + ((x213x) & (n_n4556) & (!x430x) & (!x222x) & (x14103x)) + ((x213x) & (n_n4556) & (!x430x) & (x222x) & (!x14103x)) + ((x213x) & (n_n4556) & (!x430x) & (x222x) & (x14103x)) + ((x213x) & (n_n4556) & (x430x) & (!x222x) & (!x14103x)) + ((x213x) & (n_n4556) & (x430x) & (!x222x) & (x14103x)) + ((x213x) & (n_n4556) & (x430x) & (x222x) & (!x14103x)) + ((x213x) & (n_n4556) & (x430x) & (x222x) & (x14103x)));
	assign x14108x = (((!i_9_) & (n_n455) & (n_n528) & (n_n473) & (!n_n520)) + ((!i_9_) & (n_n455) & (n_n528) & (n_n473) & (n_n520)) + ((i_9_) & (n_n455) & (!n_n528) & (n_n473) & (n_n520)) + ((i_9_) & (n_n455) & (n_n528) & (n_n473) & (n_n520)));
	assign x212x = (((!i_9_) & (n_n455) & (n_n473) & (!n_n522) & (x20x)) + ((!i_9_) & (n_n455) & (n_n473) & (n_n522) & (x20x)) + ((i_9_) & (n_n455) & (n_n473) & (!n_n522) & (x20x)) + ((i_9_) & (n_n455) & (n_n473) & (n_n522) & (!x20x)) + ((i_9_) & (n_n455) & (n_n473) & (n_n522) & (x20x)));
	assign x14109x = (((!i_9_) & (!n_n524) & (!n_n455) & (!n_n473) & (x212x)) + ((!i_9_) & (!n_n524) & (!n_n455) & (n_n473) & (x212x)) + ((!i_9_) & (!n_n524) & (n_n455) & (!n_n473) & (x212x)) + ((!i_9_) & (!n_n524) & (n_n455) & (n_n473) & (x212x)) + ((!i_9_) & (n_n524) & (!n_n455) & (!n_n473) & (x212x)) + ((!i_9_) & (n_n524) & (!n_n455) & (n_n473) & (x212x)) + ((!i_9_) & (n_n524) & (n_n455) & (!n_n473) & (x212x)) + ((!i_9_) & (n_n524) & (n_n455) & (n_n473) & (!x212x)) + ((!i_9_) & (n_n524) & (n_n455) & (n_n473) & (x212x)) + ((i_9_) & (!n_n524) & (!n_n455) & (!n_n473) & (x212x)) + ((i_9_) & (!n_n524) & (!n_n455) & (n_n473) & (x212x)) + ((i_9_) & (!n_n524) & (n_n455) & (!n_n473) & (x212x)) + ((i_9_) & (!n_n524) & (n_n455) & (n_n473) & (x212x)) + ((i_9_) & (n_n524) & (!n_n455) & (!n_n473) & (x212x)) + ((i_9_) & (n_n524) & (!n_n455) & (n_n473) & (x212x)) + ((i_9_) & (n_n524) & (n_n455) & (!n_n473) & (x212x)) + ((i_9_) & (n_n524) & (n_n455) & (n_n473) & (!x212x)) + ((i_9_) & (n_n524) & (n_n455) & (n_n473) & (x212x)));
	assign n_n4535 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n455) & (x23x)));
	assign n_n4536 = (((i_9_) & (n_n455) & (n_n473) & (n_n534)));
	assign x14112x = (((!n_n4526) & (!n_n4538) & (!n_n4535) & (n_n4536)) + ((!n_n4526) & (!n_n4538) & (n_n4535) & (!n_n4536)) + ((!n_n4526) & (!n_n4538) & (n_n4535) & (n_n4536)) + ((!n_n4526) & (n_n4538) & (!n_n4535) & (!n_n4536)) + ((!n_n4526) & (n_n4538) & (!n_n4535) & (n_n4536)) + ((!n_n4526) & (n_n4538) & (n_n4535) & (!n_n4536)) + ((!n_n4526) & (n_n4538) & (n_n4535) & (n_n4536)) + ((n_n4526) & (!n_n4538) & (!n_n4535) & (!n_n4536)) + ((n_n4526) & (!n_n4538) & (!n_n4535) & (n_n4536)) + ((n_n4526) & (!n_n4538) & (n_n4535) & (!n_n4536)) + ((n_n4526) & (!n_n4538) & (n_n4535) & (n_n4536)) + ((n_n4526) & (n_n4538) & (!n_n4535) & (!n_n4536)) + ((n_n4526) & (n_n4538) & (!n_n4535) & (n_n4536)) + ((n_n4526) & (n_n4538) & (n_n4535) & (!n_n4536)) + ((n_n4526) & (n_n4538) & (n_n4535) & (n_n4536)));
	assign x14115x = (((!n_n4525) & (!n_n3504) & (!n_n4531) & (!x14108x) & (x14109x)) + ((!n_n4525) & (!n_n3504) & (!n_n4531) & (x14108x) & (!x14109x)) + ((!n_n4525) & (!n_n3504) & (!n_n4531) & (x14108x) & (x14109x)) + ((!n_n4525) & (!n_n3504) & (n_n4531) & (!x14108x) & (!x14109x)) + ((!n_n4525) & (!n_n3504) & (n_n4531) & (!x14108x) & (x14109x)) + ((!n_n4525) & (!n_n3504) & (n_n4531) & (x14108x) & (!x14109x)) + ((!n_n4525) & (!n_n3504) & (n_n4531) & (x14108x) & (x14109x)) + ((!n_n4525) & (n_n3504) & (!n_n4531) & (!x14108x) & (!x14109x)) + ((!n_n4525) & (n_n3504) & (!n_n4531) & (!x14108x) & (x14109x)) + ((!n_n4525) & (n_n3504) & (!n_n4531) & (x14108x) & (!x14109x)) + ((!n_n4525) & (n_n3504) & (!n_n4531) & (x14108x) & (x14109x)) + ((!n_n4525) & (n_n3504) & (n_n4531) & (!x14108x) & (!x14109x)) + ((!n_n4525) & (n_n3504) & (n_n4531) & (!x14108x) & (x14109x)) + ((!n_n4525) & (n_n3504) & (n_n4531) & (x14108x) & (!x14109x)) + ((!n_n4525) & (n_n3504) & (n_n4531) & (x14108x) & (x14109x)) + ((n_n4525) & (!n_n3504) & (!n_n4531) & (!x14108x) & (!x14109x)) + ((n_n4525) & (!n_n3504) & (!n_n4531) & (!x14108x) & (x14109x)) + ((n_n4525) & (!n_n3504) & (!n_n4531) & (x14108x) & (!x14109x)) + ((n_n4525) & (!n_n3504) & (!n_n4531) & (x14108x) & (x14109x)) + ((n_n4525) & (!n_n3504) & (n_n4531) & (!x14108x) & (!x14109x)) + ((n_n4525) & (!n_n3504) & (n_n4531) & (!x14108x) & (x14109x)) + ((n_n4525) & (!n_n3504) & (n_n4531) & (x14108x) & (!x14109x)) + ((n_n4525) & (!n_n3504) & (n_n4531) & (x14108x) & (x14109x)) + ((n_n4525) & (n_n3504) & (!n_n4531) & (!x14108x) & (!x14109x)) + ((n_n4525) & (n_n3504) & (!n_n4531) & (!x14108x) & (x14109x)) + ((n_n4525) & (n_n3504) & (!n_n4531) & (x14108x) & (!x14109x)) + ((n_n4525) & (n_n3504) & (!n_n4531) & (x14108x) & (x14109x)) + ((n_n4525) & (n_n3504) & (n_n4531) & (!x14108x) & (!x14109x)) + ((n_n4525) & (n_n3504) & (n_n4531) & (!x14108x) & (x14109x)) + ((n_n4525) & (n_n3504) & (n_n4531) & (x14108x) & (!x14109x)) + ((n_n4525) & (n_n3504) & (n_n4531) & (x14108x) & (x14109x)));
	assign x14117x = (((!n_n3871) & (!n_n3350) & (!x14112x) & (x14115x)) + ((!n_n3871) & (!n_n3350) & (x14112x) & (!x14115x)) + ((!n_n3871) & (!n_n3350) & (x14112x) & (x14115x)) + ((!n_n3871) & (n_n3350) & (!x14112x) & (!x14115x)) + ((!n_n3871) & (n_n3350) & (!x14112x) & (x14115x)) + ((!n_n3871) & (n_n3350) & (x14112x) & (!x14115x)) + ((!n_n3871) & (n_n3350) & (x14112x) & (x14115x)) + ((n_n3871) & (!n_n3350) & (!x14112x) & (!x14115x)) + ((n_n3871) & (!n_n3350) & (!x14112x) & (x14115x)) + ((n_n3871) & (!n_n3350) & (x14112x) & (!x14115x)) + ((n_n3871) & (!n_n3350) & (x14112x) & (x14115x)) + ((n_n3871) & (n_n3350) & (!x14112x) & (!x14115x)) + ((n_n3871) & (n_n3350) & (!x14112x) & (x14115x)) + ((n_n3871) & (n_n3350) & (x14112x) & (!x14115x)) + ((n_n3871) & (n_n3350) & (x14112x) & (x14115x)));
	assign n_n3260 = (((!n_n3347) & (!n_n3281) & (!n_n3348) & (!x14101x) & (x14117x)) + ((!n_n3347) & (!n_n3281) & (!n_n3348) & (x14101x) & (!x14117x)) + ((!n_n3347) & (!n_n3281) & (!n_n3348) & (x14101x) & (x14117x)) + ((!n_n3347) & (!n_n3281) & (n_n3348) & (!x14101x) & (!x14117x)) + ((!n_n3347) & (!n_n3281) & (n_n3348) & (!x14101x) & (x14117x)) + ((!n_n3347) & (!n_n3281) & (n_n3348) & (x14101x) & (!x14117x)) + ((!n_n3347) & (!n_n3281) & (n_n3348) & (x14101x) & (x14117x)) + ((!n_n3347) & (n_n3281) & (!n_n3348) & (!x14101x) & (!x14117x)) + ((!n_n3347) & (n_n3281) & (!n_n3348) & (!x14101x) & (x14117x)) + ((!n_n3347) & (n_n3281) & (!n_n3348) & (x14101x) & (!x14117x)) + ((!n_n3347) & (n_n3281) & (!n_n3348) & (x14101x) & (x14117x)) + ((!n_n3347) & (n_n3281) & (n_n3348) & (!x14101x) & (!x14117x)) + ((!n_n3347) & (n_n3281) & (n_n3348) & (!x14101x) & (x14117x)) + ((!n_n3347) & (n_n3281) & (n_n3348) & (x14101x) & (!x14117x)) + ((!n_n3347) & (n_n3281) & (n_n3348) & (x14101x) & (x14117x)) + ((n_n3347) & (!n_n3281) & (!n_n3348) & (!x14101x) & (!x14117x)) + ((n_n3347) & (!n_n3281) & (!n_n3348) & (!x14101x) & (x14117x)) + ((n_n3347) & (!n_n3281) & (!n_n3348) & (x14101x) & (!x14117x)) + ((n_n3347) & (!n_n3281) & (!n_n3348) & (x14101x) & (x14117x)) + ((n_n3347) & (!n_n3281) & (n_n3348) & (!x14101x) & (!x14117x)) + ((n_n3347) & (!n_n3281) & (n_n3348) & (!x14101x) & (x14117x)) + ((n_n3347) & (!n_n3281) & (n_n3348) & (x14101x) & (!x14117x)) + ((n_n3347) & (!n_n3281) & (n_n3348) & (x14101x) & (x14117x)) + ((n_n3347) & (n_n3281) & (!n_n3348) & (!x14101x) & (!x14117x)) + ((n_n3347) & (n_n3281) & (!n_n3348) & (!x14101x) & (x14117x)) + ((n_n3347) & (n_n3281) & (!n_n3348) & (x14101x) & (!x14117x)) + ((n_n3347) & (n_n3281) & (!n_n3348) & (x14101x) & (x14117x)) + ((n_n3347) & (n_n3281) & (n_n3348) & (!x14101x) & (!x14117x)) + ((n_n3347) & (n_n3281) & (n_n3348) & (!x14101x) & (x14117x)) + ((n_n3347) & (n_n3281) & (n_n3348) & (x14101x) & (!x14117x)) + ((n_n3347) & (n_n3281) & (n_n3348) & (x14101x) & (x14117x)));
	assign n_n4629 = (((!i_1_) & (i_2_) & (i_0_) & (x20x) & (n_n500)));
	assign n_n4583 = (((!i_1_) & (i_2_) & (i_0_) & (n_n535) & (x23x)));
	assign n_n5182 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n473) & (x12x)));
	assign n_n5173 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n130) & (x20x)));
	assign n_n5165 = (((!i_9_) & (n_n482) & (n_n130) & (n_n530)));
	assign n_n5230 = (((!i_5_) & (i_3_) & (i_4_) & (x19x) & (n_n528)));
	assign n_n5166 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n528) & (x12x)));
	assign n_n5163 = (((!i_9_) & (n_n482) & (n_n532) & (n_n130)));
	assign n_n5214 = (((!i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n535)));
	assign n_n5033 = (((!i_9_) & (n_n482) & (n_n534) & (n_n195)));
	assign n_n5051 = (((!i_9_) & (n_n473) & (n_n532) & (n_n195)));
	assign n_n5072 = (((i_9_) & (n_n526) & (n_n195) & (n_n464)));
	assign n_n5082 = (((i_7_) & (!i_8_) & (i_6_) & (n_n535) & (x12x)));
	assign n_n5075 = (((!i_9_) & (n_n524) & (n_n195) & (n_n464)));
	assign x13719x = (((!n_n5085) & (!n_n5072) & (!n_n5082) & (n_n5075)) + ((!n_n5085) & (!n_n5072) & (n_n5082) & (!n_n5075)) + ((!n_n5085) & (!n_n5072) & (n_n5082) & (n_n5075)) + ((!n_n5085) & (n_n5072) & (!n_n5082) & (!n_n5075)) + ((!n_n5085) & (n_n5072) & (!n_n5082) & (n_n5075)) + ((!n_n5085) & (n_n5072) & (n_n5082) & (!n_n5075)) + ((!n_n5085) & (n_n5072) & (n_n5082) & (n_n5075)) + ((n_n5085) & (!n_n5072) & (!n_n5082) & (!n_n5075)) + ((n_n5085) & (!n_n5072) & (!n_n5082) & (n_n5075)) + ((n_n5085) & (!n_n5072) & (n_n5082) & (!n_n5075)) + ((n_n5085) & (!n_n5072) & (n_n5082) & (n_n5075)) + ((n_n5085) & (n_n5072) & (!n_n5082) & (!n_n5075)) + ((n_n5085) & (n_n5072) & (!n_n5082) & (n_n5075)) + ((n_n5085) & (n_n5072) & (n_n5082) & (!n_n5075)) + ((n_n5085) & (n_n5072) & (n_n5082) & (n_n5075)));
	assign n_n5079 = (((i_1_) & (!i_2_) & (!i_0_) & (x23x) & (n_n464)));
	assign n_n5065 = (((!i_9_) & (n_n534) & (n_n195) & (n_n464)));
	assign x13720x = (((!n_n5096) & (!n_n5099) & (!n_n5063) & (!n_n5079) & (n_n5065)) + ((!n_n5096) & (!n_n5099) & (!n_n5063) & (n_n5079) & (!n_n5065)) + ((!n_n5096) & (!n_n5099) & (!n_n5063) & (n_n5079) & (n_n5065)) + ((!n_n5096) & (!n_n5099) & (n_n5063) & (!n_n5079) & (!n_n5065)) + ((!n_n5096) & (!n_n5099) & (n_n5063) & (!n_n5079) & (n_n5065)) + ((!n_n5096) & (!n_n5099) & (n_n5063) & (n_n5079) & (!n_n5065)) + ((!n_n5096) & (!n_n5099) & (n_n5063) & (n_n5079) & (n_n5065)) + ((!n_n5096) & (n_n5099) & (!n_n5063) & (!n_n5079) & (!n_n5065)) + ((!n_n5096) & (n_n5099) & (!n_n5063) & (!n_n5079) & (n_n5065)) + ((!n_n5096) & (n_n5099) & (!n_n5063) & (n_n5079) & (!n_n5065)) + ((!n_n5096) & (n_n5099) & (!n_n5063) & (n_n5079) & (n_n5065)) + ((!n_n5096) & (n_n5099) & (n_n5063) & (!n_n5079) & (!n_n5065)) + ((!n_n5096) & (n_n5099) & (n_n5063) & (!n_n5079) & (n_n5065)) + ((!n_n5096) & (n_n5099) & (n_n5063) & (n_n5079) & (!n_n5065)) + ((!n_n5096) & (n_n5099) & (n_n5063) & (n_n5079) & (n_n5065)) + ((n_n5096) & (!n_n5099) & (!n_n5063) & (!n_n5079) & (!n_n5065)) + ((n_n5096) & (!n_n5099) & (!n_n5063) & (!n_n5079) & (n_n5065)) + ((n_n5096) & (!n_n5099) & (!n_n5063) & (n_n5079) & (!n_n5065)) + ((n_n5096) & (!n_n5099) & (!n_n5063) & (n_n5079) & (n_n5065)) + ((n_n5096) & (!n_n5099) & (n_n5063) & (!n_n5079) & (!n_n5065)) + ((n_n5096) & (!n_n5099) & (n_n5063) & (!n_n5079) & (n_n5065)) + ((n_n5096) & (!n_n5099) & (n_n5063) & (n_n5079) & (!n_n5065)) + ((n_n5096) & (!n_n5099) & (n_n5063) & (n_n5079) & (n_n5065)) + ((n_n5096) & (n_n5099) & (!n_n5063) & (!n_n5079) & (!n_n5065)) + ((n_n5096) & (n_n5099) & (!n_n5063) & (!n_n5079) & (n_n5065)) + ((n_n5096) & (n_n5099) & (!n_n5063) & (n_n5079) & (!n_n5065)) + ((n_n5096) & (n_n5099) & (!n_n5063) & (n_n5079) & (n_n5065)) + ((n_n5096) & (n_n5099) & (n_n5063) & (!n_n5079) & (!n_n5065)) + ((n_n5096) & (n_n5099) & (n_n5063) & (!n_n5079) & (n_n5065)) + ((n_n5096) & (n_n5099) & (n_n5063) & (n_n5079) & (!n_n5065)) + ((n_n5096) & (n_n5099) & (n_n5063) & (n_n5079) & (n_n5065)));
	assign n_n4454 = (((i_9_) & (n_n455) & (n_n535) & (n_n520)));
	assign n_n4517 = (((i_1_) & (!i_2_) & (i_0_) & (n_n491) & (x20x)));
	assign n_n3152 = (((!i_9_) & (n_n455) & (n_n491) & (!n_n520) & (x20x)) + ((!i_9_) & (n_n455) & (n_n491) & (n_n520) & (!x20x)) + ((!i_9_) & (n_n455) & (n_n491) & (n_n520) & (x20x)) + ((i_9_) & (n_n455) & (n_n491) & (!n_n520) & (x20x)) + ((i_9_) & (n_n455) & (n_n491) & (n_n520) & (!x20x)) + ((i_9_) & (n_n455) & (n_n491) & (n_n520) & (x20x)));
	assign n_n5039 = (((!i_9_) & (n_n482) & (n_n528) & (n_n195)));
	assign n_n5103 = (((!i_9_) & (n_n518) & (n_n528) & (n_n130)));
	assign n_n5104 = (((!i_5_) & (i_3_) & (i_4_) & (n_n526) & (x12x)));
	assign n_n5102 = (((!i_5_) & (i_3_) & (i_4_) & (n_n528) & (x12x)));
	assign n_n4395 = (((!i_9_) & (n_n536) & (n_n482) & (n_n532)));
	assign x281x = (((!i_9_) & (n_n536) & (n_n532) & (n_n491) & (!n_n530)) + ((!i_9_) & (n_n536) & (n_n532) & (n_n491) & (n_n530)) + ((i_9_) & (n_n536) & (!n_n532) & (n_n491) & (n_n530)) + ((i_9_) & (n_n536) & (n_n532) & (n_n491) & (n_n530)));
	assign n_n3176 = (((!i_9_) & (n_n536) & (!n_n532) & (n_n534) & (n_n491)) + ((!i_9_) & (n_n536) & (n_n532) & (n_n534) & (n_n491)) + ((i_9_) & (n_n536) & (!n_n532) & (n_n534) & (n_n491)) + ((i_9_) & (n_n536) & (n_n532) & (!n_n534) & (n_n491)) + ((i_9_) & (n_n536) & (n_n532) & (n_n534) & (n_n491)));
	assign x64x = (((!i_9_) & (n_n536) & (!n_n526) & (n_n528) & (n_n500)) + ((!i_9_) & (n_n536) & (n_n526) & (n_n528) & (n_n500)) + ((i_9_) & (n_n536) & (n_n526) & (!n_n528) & (n_n500)) + ((i_9_) & (n_n536) & (n_n526) & (n_n528) & (n_n500)));
	assign n_n2637 = (((!n_n4384) & (!n_n4374) & (!x281x) & (!n_n3176) & (x64x)) + ((!n_n4384) & (!n_n4374) & (!x281x) & (n_n3176) & (!x64x)) + ((!n_n4384) & (!n_n4374) & (!x281x) & (n_n3176) & (x64x)) + ((!n_n4384) & (!n_n4374) & (x281x) & (!n_n3176) & (!x64x)) + ((!n_n4384) & (!n_n4374) & (x281x) & (!n_n3176) & (x64x)) + ((!n_n4384) & (!n_n4374) & (x281x) & (n_n3176) & (!x64x)) + ((!n_n4384) & (!n_n4374) & (x281x) & (n_n3176) & (x64x)) + ((!n_n4384) & (n_n4374) & (!x281x) & (!n_n3176) & (!x64x)) + ((!n_n4384) & (n_n4374) & (!x281x) & (!n_n3176) & (x64x)) + ((!n_n4384) & (n_n4374) & (!x281x) & (n_n3176) & (!x64x)) + ((!n_n4384) & (n_n4374) & (!x281x) & (n_n3176) & (x64x)) + ((!n_n4384) & (n_n4374) & (x281x) & (!n_n3176) & (!x64x)) + ((!n_n4384) & (n_n4374) & (x281x) & (!n_n3176) & (x64x)) + ((!n_n4384) & (n_n4374) & (x281x) & (n_n3176) & (!x64x)) + ((!n_n4384) & (n_n4374) & (x281x) & (n_n3176) & (x64x)) + ((n_n4384) & (!n_n4374) & (!x281x) & (!n_n3176) & (!x64x)) + ((n_n4384) & (!n_n4374) & (!x281x) & (!n_n3176) & (x64x)) + ((n_n4384) & (!n_n4374) & (!x281x) & (n_n3176) & (!x64x)) + ((n_n4384) & (!n_n4374) & (!x281x) & (n_n3176) & (x64x)) + ((n_n4384) & (!n_n4374) & (x281x) & (!n_n3176) & (!x64x)) + ((n_n4384) & (!n_n4374) & (x281x) & (!n_n3176) & (x64x)) + ((n_n4384) & (!n_n4374) & (x281x) & (n_n3176) & (!x64x)) + ((n_n4384) & (!n_n4374) & (x281x) & (n_n3176) & (x64x)) + ((n_n4384) & (n_n4374) & (!x281x) & (!n_n3176) & (!x64x)) + ((n_n4384) & (n_n4374) & (!x281x) & (!n_n3176) & (x64x)) + ((n_n4384) & (n_n4374) & (!x281x) & (n_n3176) & (!x64x)) + ((n_n4384) & (n_n4374) & (!x281x) & (n_n3176) & (x64x)) + ((n_n4384) & (n_n4374) & (x281x) & (!n_n3176) & (!x64x)) + ((n_n4384) & (n_n4374) & (x281x) & (!n_n3176) & (x64x)) + ((n_n4384) & (n_n4374) & (x281x) & (n_n3176) & (!x64x)) + ((n_n4384) & (n_n4374) & (x281x) & (n_n3176) & (x64x)));
	assign x15033x = (((!n_n4361) & (!n_n4363) & (!n_n4359) & (n_n4364)) + ((!n_n4361) & (!n_n4363) & (n_n4359) & (!n_n4364)) + ((!n_n4361) & (!n_n4363) & (n_n4359) & (n_n4364)) + ((!n_n4361) & (n_n4363) & (!n_n4359) & (!n_n4364)) + ((!n_n4361) & (n_n4363) & (!n_n4359) & (n_n4364)) + ((!n_n4361) & (n_n4363) & (n_n4359) & (!n_n4364)) + ((!n_n4361) & (n_n4363) & (n_n4359) & (n_n4364)) + ((n_n4361) & (!n_n4363) & (!n_n4359) & (!n_n4364)) + ((n_n4361) & (!n_n4363) & (!n_n4359) & (n_n4364)) + ((n_n4361) & (!n_n4363) & (n_n4359) & (!n_n4364)) + ((n_n4361) & (!n_n4363) & (n_n4359) & (n_n4364)) + ((n_n4361) & (n_n4363) & (!n_n4359) & (!n_n4364)) + ((n_n4361) & (n_n4363) & (!n_n4359) & (n_n4364)) + ((n_n4361) & (n_n4363) & (n_n4359) & (!n_n4364)) + ((n_n4361) & (n_n4363) & (n_n4359) & (n_n4364)));
	assign n_n4356 = (((i_9_) & (n_n536) & (n_n509) & (n_n522)));
	assign x15034x = (((!n_n4366) & (!n_n4357) & (!n_n4358) & (!n_n4356) & (n_n4355)) + ((!n_n4366) & (!n_n4357) & (!n_n4358) & (n_n4356) & (!n_n4355)) + ((!n_n4366) & (!n_n4357) & (!n_n4358) & (n_n4356) & (n_n4355)) + ((!n_n4366) & (!n_n4357) & (n_n4358) & (!n_n4356) & (!n_n4355)) + ((!n_n4366) & (!n_n4357) & (n_n4358) & (!n_n4356) & (n_n4355)) + ((!n_n4366) & (!n_n4357) & (n_n4358) & (n_n4356) & (!n_n4355)) + ((!n_n4366) & (!n_n4357) & (n_n4358) & (n_n4356) & (n_n4355)) + ((!n_n4366) & (n_n4357) & (!n_n4358) & (!n_n4356) & (!n_n4355)) + ((!n_n4366) & (n_n4357) & (!n_n4358) & (!n_n4356) & (n_n4355)) + ((!n_n4366) & (n_n4357) & (!n_n4358) & (n_n4356) & (!n_n4355)) + ((!n_n4366) & (n_n4357) & (!n_n4358) & (n_n4356) & (n_n4355)) + ((!n_n4366) & (n_n4357) & (n_n4358) & (!n_n4356) & (!n_n4355)) + ((!n_n4366) & (n_n4357) & (n_n4358) & (!n_n4356) & (n_n4355)) + ((!n_n4366) & (n_n4357) & (n_n4358) & (n_n4356) & (!n_n4355)) + ((!n_n4366) & (n_n4357) & (n_n4358) & (n_n4356) & (n_n4355)) + ((n_n4366) & (!n_n4357) & (!n_n4358) & (!n_n4356) & (!n_n4355)) + ((n_n4366) & (!n_n4357) & (!n_n4358) & (!n_n4356) & (n_n4355)) + ((n_n4366) & (!n_n4357) & (!n_n4358) & (n_n4356) & (!n_n4355)) + ((n_n4366) & (!n_n4357) & (!n_n4358) & (n_n4356) & (n_n4355)) + ((n_n4366) & (!n_n4357) & (n_n4358) & (!n_n4356) & (!n_n4355)) + ((n_n4366) & (!n_n4357) & (n_n4358) & (!n_n4356) & (n_n4355)) + ((n_n4366) & (!n_n4357) & (n_n4358) & (n_n4356) & (!n_n4355)) + ((n_n4366) & (!n_n4357) & (n_n4358) & (n_n4356) & (n_n4355)) + ((n_n4366) & (n_n4357) & (!n_n4358) & (!n_n4356) & (!n_n4355)) + ((n_n4366) & (n_n4357) & (!n_n4358) & (!n_n4356) & (n_n4355)) + ((n_n4366) & (n_n4357) & (!n_n4358) & (n_n4356) & (!n_n4355)) + ((n_n4366) & (n_n4357) & (!n_n4358) & (n_n4356) & (n_n4355)) + ((n_n4366) & (n_n4357) & (n_n4358) & (!n_n4356) & (!n_n4355)) + ((n_n4366) & (n_n4357) & (n_n4358) & (!n_n4356) & (n_n4355)) + ((n_n4366) & (n_n4357) & (n_n4358) & (n_n4356) & (!n_n4355)) + ((n_n4366) & (n_n4357) & (n_n4358) & (n_n4356) & (n_n4355)));
	assign n_n4394 = (((i_9_) & (n_n536) & (n_n482) & (n_n532)));
	assign x216x = (((!i_9_) & (n_n536) & (n_n482) & (!n_n532) & (n_n534)) + ((!i_9_) & (n_n536) & (n_n482) & (n_n532) & (n_n534)) + ((i_9_) & (n_n536) & (n_n482) & (n_n532) & (!n_n534)) + ((i_9_) & (n_n536) & (n_n482) & (n_n532) & (n_n534)));
	assign n_n4386 = (((i_9_) & (n_n536) & (n_n524) & (n_n491)));
	assign n_n4387 = (((!i_9_) & (n_n536) & (n_n524) & (n_n491)));
	assign x425x = (((!i_9_) & (n_n536) & (n_n524) & (n_n491)) + ((i_9_) & (n_n536) & (n_n524) & (n_n491)));
	assign x22099x = (((!n_n4389) & (!n_n4385) & (!n_n4388) & (!n_n4392)));
	assign x15040x = (((!n_n4393) & (!n_n4395) & (!n_n4394) & (!x425x) & (!x22099x)) + ((!n_n4393) & (!n_n4395) & (!n_n4394) & (x425x) & (!x22099x)) + ((!n_n4393) & (!n_n4395) & (!n_n4394) & (x425x) & (x22099x)) + ((!n_n4393) & (!n_n4395) & (n_n4394) & (!x425x) & (!x22099x)) + ((!n_n4393) & (!n_n4395) & (n_n4394) & (!x425x) & (x22099x)) + ((!n_n4393) & (!n_n4395) & (n_n4394) & (x425x) & (!x22099x)) + ((!n_n4393) & (!n_n4395) & (n_n4394) & (x425x) & (x22099x)) + ((!n_n4393) & (n_n4395) & (!n_n4394) & (!x425x) & (!x22099x)) + ((!n_n4393) & (n_n4395) & (!n_n4394) & (!x425x) & (x22099x)) + ((!n_n4393) & (n_n4395) & (!n_n4394) & (x425x) & (!x22099x)) + ((!n_n4393) & (n_n4395) & (!n_n4394) & (x425x) & (x22099x)) + ((!n_n4393) & (n_n4395) & (n_n4394) & (!x425x) & (!x22099x)) + ((!n_n4393) & (n_n4395) & (n_n4394) & (!x425x) & (x22099x)) + ((!n_n4393) & (n_n4395) & (n_n4394) & (x425x) & (!x22099x)) + ((!n_n4393) & (n_n4395) & (n_n4394) & (x425x) & (x22099x)) + ((n_n4393) & (!n_n4395) & (!n_n4394) & (!x425x) & (!x22099x)) + ((n_n4393) & (!n_n4395) & (!n_n4394) & (!x425x) & (x22099x)) + ((n_n4393) & (!n_n4395) & (!n_n4394) & (x425x) & (!x22099x)) + ((n_n4393) & (!n_n4395) & (!n_n4394) & (x425x) & (x22099x)) + ((n_n4393) & (!n_n4395) & (n_n4394) & (!x425x) & (!x22099x)) + ((n_n4393) & (!n_n4395) & (n_n4394) & (!x425x) & (x22099x)) + ((n_n4393) & (!n_n4395) & (n_n4394) & (x425x) & (!x22099x)) + ((n_n4393) & (!n_n4395) & (n_n4394) & (x425x) & (x22099x)) + ((n_n4393) & (n_n4395) & (!n_n4394) & (!x425x) & (!x22099x)) + ((n_n4393) & (n_n4395) & (!n_n4394) & (!x425x) & (x22099x)) + ((n_n4393) & (n_n4395) & (!n_n4394) & (x425x) & (!x22099x)) + ((n_n4393) & (n_n4395) & (!n_n4394) & (x425x) & (x22099x)) + ((n_n4393) & (n_n4395) & (n_n4394) & (!x425x) & (!x22099x)) + ((n_n4393) & (n_n4395) & (n_n4394) & (!x425x) & (x22099x)) + ((n_n4393) & (n_n4395) & (n_n4394) & (x425x) & (!x22099x)) + ((n_n4393) & (n_n4395) & (n_n4394) & (x425x) & (x22099x)));
	assign n_n4426 = (((i_9_) & (n_n536) & (n_n532) & (n_n464)));
	assign n_n4414 = (((i_9_) & (n_n536) & (n_n528) & (n_n473)));
	assign x215x = (((!i_9_) & (n_n536) & (n_n473) & (!n_n520) & (x23x)) + ((!i_9_) & (n_n536) & (n_n473) & (n_n520) & (x23x)) + ((i_9_) & (n_n536) & (n_n473) & (!n_n520) & (x23x)) + ((i_9_) & (n_n536) & (n_n473) & (n_n520) & (!x23x)) + ((i_9_) & (n_n536) & (n_n473) & (n_n520) & (x23x)));
	assign x15045x = (((!n_n4421) & (!n_n4410) & (!n_n4414) & (x215x)) + ((!n_n4421) & (!n_n4410) & (n_n4414) & (!x215x)) + ((!n_n4421) & (!n_n4410) & (n_n4414) & (x215x)) + ((!n_n4421) & (n_n4410) & (!n_n4414) & (!x215x)) + ((!n_n4421) & (n_n4410) & (!n_n4414) & (x215x)) + ((!n_n4421) & (n_n4410) & (n_n4414) & (!x215x)) + ((!n_n4421) & (n_n4410) & (n_n4414) & (x215x)) + ((n_n4421) & (!n_n4410) & (!n_n4414) & (!x215x)) + ((n_n4421) & (!n_n4410) & (!n_n4414) & (x215x)) + ((n_n4421) & (!n_n4410) & (n_n4414) & (!x215x)) + ((n_n4421) & (!n_n4410) & (n_n4414) & (x215x)) + ((n_n4421) & (n_n4410) & (!n_n4414) & (!x215x)) + ((n_n4421) & (n_n4410) & (!n_n4414) & (x215x)) + ((n_n4421) & (n_n4410) & (n_n4414) & (!x215x)) + ((n_n4421) & (n_n4410) & (n_n4414) & (x215x)));
	assign n_n4419 = (((!i_9_) & (n_n536) & (n_n524) & (n_n473)));
	assign n_n4411 = (((!i_9_) & (n_n536) & (n_n473) & (n_n532)));
	assign n_n4412 = (((i_9_) & (n_n536) & (n_n473) & (n_n530)));
	assign n_n2634 = (((!x15045x) & (!n_n4419) & (!n_n4417) & (!n_n4411) & (n_n4412)) + ((!x15045x) & (!n_n4419) & (!n_n4417) & (n_n4411) & (!n_n4412)) + ((!x15045x) & (!n_n4419) & (!n_n4417) & (n_n4411) & (n_n4412)) + ((!x15045x) & (!n_n4419) & (n_n4417) & (!n_n4411) & (!n_n4412)) + ((!x15045x) & (!n_n4419) & (n_n4417) & (!n_n4411) & (n_n4412)) + ((!x15045x) & (!n_n4419) & (n_n4417) & (n_n4411) & (!n_n4412)) + ((!x15045x) & (!n_n4419) & (n_n4417) & (n_n4411) & (n_n4412)) + ((!x15045x) & (n_n4419) & (!n_n4417) & (!n_n4411) & (!n_n4412)) + ((!x15045x) & (n_n4419) & (!n_n4417) & (!n_n4411) & (n_n4412)) + ((!x15045x) & (n_n4419) & (!n_n4417) & (n_n4411) & (!n_n4412)) + ((!x15045x) & (n_n4419) & (!n_n4417) & (n_n4411) & (n_n4412)) + ((!x15045x) & (n_n4419) & (n_n4417) & (!n_n4411) & (!n_n4412)) + ((!x15045x) & (n_n4419) & (n_n4417) & (!n_n4411) & (n_n4412)) + ((!x15045x) & (n_n4419) & (n_n4417) & (n_n4411) & (!n_n4412)) + ((!x15045x) & (n_n4419) & (n_n4417) & (n_n4411) & (n_n4412)) + ((x15045x) & (!n_n4419) & (!n_n4417) & (!n_n4411) & (!n_n4412)) + ((x15045x) & (!n_n4419) & (!n_n4417) & (!n_n4411) & (n_n4412)) + ((x15045x) & (!n_n4419) & (!n_n4417) & (n_n4411) & (!n_n4412)) + ((x15045x) & (!n_n4419) & (!n_n4417) & (n_n4411) & (n_n4412)) + ((x15045x) & (!n_n4419) & (n_n4417) & (!n_n4411) & (!n_n4412)) + ((x15045x) & (!n_n4419) & (n_n4417) & (!n_n4411) & (n_n4412)) + ((x15045x) & (!n_n4419) & (n_n4417) & (n_n4411) & (!n_n4412)) + ((x15045x) & (!n_n4419) & (n_n4417) & (n_n4411) & (n_n4412)) + ((x15045x) & (n_n4419) & (!n_n4417) & (!n_n4411) & (!n_n4412)) + ((x15045x) & (n_n4419) & (!n_n4417) & (!n_n4411) & (n_n4412)) + ((x15045x) & (n_n4419) & (!n_n4417) & (n_n4411) & (!n_n4412)) + ((x15045x) & (n_n4419) & (!n_n4417) & (n_n4411) & (n_n4412)) + ((x15045x) & (n_n4419) & (n_n4417) & (!n_n4411) & (!n_n4412)) + ((x15045x) & (n_n4419) & (n_n4417) & (!n_n4411) & (n_n4412)) + ((x15045x) & (n_n4419) & (n_n4417) & (n_n4411) & (!n_n4412)) + ((x15045x) & (n_n4419) & (n_n4417) & (n_n4411) & (n_n4412)));
	assign x15049x = (((!n_n4401) & (!n_n4400) & (!n_n4397) & (n_n4398)) + ((!n_n4401) & (!n_n4400) & (n_n4397) & (!n_n4398)) + ((!n_n4401) & (!n_n4400) & (n_n4397) & (n_n4398)) + ((!n_n4401) & (n_n4400) & (!n_n4397) & (!n_n4398)) + ((!n_n4401) & (n_n4400) & (!n_n4397) & (n_n4398)) + ((!n_n4401) & (n_n4400) & (n_n4397) & (!n_n4398)) + ((!n_n4401) & (n_n4400) & (n_n4397) & (n_n4398)) + ((n_n4401) & (!n_n4400) & (!n_n4397) & (!n_n4398)) + ((n_n4401) & (!n_n4400) & (!n_n4397) & (n_n4398)) + ((n_n4401) & (!n_n4400) & (n_n4397) & (!n_n4398)) + ((n_n4401) & (!n_n4400) & (n_n4397) & (n_n4398)) + ((n_n4401) & (n_n4400) & (!n_n4397) & (!n_n4398)) + ((n_n4401) & (n_n4400) & (!n_n4397) & (n_n4398)) + ((n_n4401) & (n_n4400) & (n_n4397) & (!n_n4398)) + ((n_n4401) & (n_n4400) & (n_n4397) & (n_n4398)));
	assign x15050x = (((!n_n4404) & (!n_n4405) & (!n_n4406) & (!n_n4409) & (n_n4408)) + ((!n_n4404) & (!n_n4405) & (!n_n4406) & (n_n4409) & (!n_n4408)) + ((!n_n4404) & (!n_n4405) & (!n_n4406) & (n_n4409) & (n_n4408)) + ((!n_n4404) & (!n_n4405) & (n_n4406) & (!n_n4409) & (!n_n4408)) + ((!n_n4404) & (!n_n4405) & (n_n4406) & (!n_n4409) & (n_n4408)) + ((!n_n4404) & (!n_n4405) & (n_n4406) & (n_n4409) & (!n_n4408)) + ((!n_n4404) & (!n_n4405) & (n_n4406) & (n_n4409) & (n_n4408)) + ((!n_n4404) & (n_n4405) & (!n_n4406) & (!n_n4409) & (!n_n4408)) + ((!n_n4404) & (n_n4405) & (!n_n4406) & (!n_n4409) & (n_n4408)) + ((!n_n4404) & (n_n4405) & (!n_n4406) & (n_n4409) & (!n_n4408)) + ((!n_n4404) & (n_n4405) & (!n_n4406) & (n_n4409) & (n_n4408)) + ((!n_n4404) & (n_n4405) & (n_n4406) & (!n_n4409) & (!n_n4408)) + ((!n_n4404) & (n_n4405) & (n_n4406) & (!n_n4409) & (n_n4408)) + ((!n_n4404) & (n_n4405) & (n_n4406) & (n_n4409) & (!n_n4408)) + ((!n_n4404) & (n_n4405) & (n_n4406) & (n_n4409) & (n_n4408)) + ((n_n4404) & (!n_n4405) & (!n_n4406) & (!n_n4409) & (!n_n4408)) + ((n_n4404) & (!n_n4405) & (!n_n4406) & (!n_n4409) & (n_n4408)) + ((n_n4404) & (!n_n4405) & (!n_n4406) & (n_n4409) & (!n_n4408)) + ((n_n4404) & (!n_n4405) & (!n_n4406) & (n_n4409) & (n_n4408)) + ((n_n4404) & (!n_n4405) & (n_n4406) & (!n_n4409) & (!n_n4408)) + ((n_n4404) & (!n_n4405) & (n_n4406) & (!n_n4409) & (n_n4408)) + ((n_n4404) & (!n_n4405) & (n_n4406) & (n_n4409) & (!n_n4408)) + ((n_n4404) & (!n_n4405) & (n_n4406) & (n_n4409) & (n_n4408)) + ((n_n4404) & (n_n4405) & (!n_n4406) & (!n_n4409) & (!n_n4408)) + ((n_n4404) & (n_n4405) & (!n_n4406) & (!n_n4409) & (n_n4408)) + ((n_n4404) & (n_n4405) & (!n_n4406) & (n_n4409) & (!n_n4408)) + ((n_n4404) & (n_n4405) & (!n_n4406) & (n_n4409) & (n_n4408)) + ((n_n4404) & (n_n4405) & (n_n4406) & (!n_n4409) & (!n_n4408)) + ((n_n4404) & (n_n4405) & (n_n4406) & (!n_n4409) & (n_n4408)) + ((n_n4404) & (n_n4405) & (n_n4406) & (n_n4409) & (!n_n4408)) + ((n_n4404) & (n_n4405) & (n_n4406) & (n_n4409) & (n_n4408)));
	assign n_n2802 = (((!i_9_) & (n_n536) & (!n_n532) & (n_n530) & (n_n464)) + ((!i_9_) & (n_n536) & (n_n532) & (!n_n530) & (n_n464)) + ((!i_9_) & (n_n536) & (n_n532) & (n_n530) & (n_n464)) + ((i_9_) & (n_n536) & (!n_n532) & (n_n530) & (n_n464)) + ((i_9_) & (n_n536) & (n_n532) & (n_n530) & (n_n464)));
	assign x37x = (((!i_9_) & (n_n536) & (n_n534) & (n_n464)) + ((i_9_) & (n_n536) & (n_n534) & (n_n464)));
	assign x15051x = (((!i_9_) & (n_n536) & (!n_n526) & (n_n528) & (n_n464)) + ((!i_9_) & (n_n536) & (n_n526) & (n_n528) & (n_n464)) + ((i_9_) & (n_n536) & (n_n526) & (!n_n528) & (n_n464)) + ((i_9_) & (n_n536) & (n_n526) & (n_n528) & (n_n464)));
	assign x15055x = (((!n_n4430) & (!n_n4426) & (!n_n2802) & (!x37x) & (x15051x)) + ((!n_n4430) & (!n_n4426) & (!n_n2802) & (x37x) & (!x15051x)) + ((!n_n4430) & (!n_n4426) & (!n_n2802) & (x37x) & (x15051x)) + ((!n_n4430) & (!n_n4426) & (n_n2802) & (!x37x) & (!x15051x)) + ((!n_n4430) & (!n_n4426) & (n_n2802) & (!x37x) & (x15051x)) + ((!n_n4430) & (!n_n4426) & (n_n2802) & (x37x) & (!x15051x)) + ((!n_n4430) & (!n_n4426) & (n_n2802) & (x37x) & (x15051x)) + ((!n_n4430) & (n_n4426) & (!n_n2802) & (!x37x) & (!x15051x)) + ((!n_n4430) & (n_n4426) & (!n_n2802) & (!x37x) & (x15051x)) + ((!n_n4430) & (n_n4426) & (!n_n2802) & (x37x) & (!x15051x)) + ((!n_n4430) & (n_n4426) & (!n_n2802) & (x37x) & (x15051x)) + ((!n_n4430) & (n_n4426) & (n_n2802) & (!x37x) & (!x15051x)) + ((!n_n4430) & (n_n4426) & (n_n2802) & (!x37x) & (x15051x)) + ((!n_n4430) & (n_n4426) & (n_n2802) & (x37x) & (!x15051x)) + ((!n_n4430) & (n_n4426) & (n_n2802) & (x37x) & (x15051x)) + ((n_n4430) & (!n_n4426) & (!n_n2802) & (!x37x) & (!x15051x)) + ((n_n4430) & (!n_n4426) & (!n_n2802) & (!x37x) & (x15051x)) + ((n_n4430) & (!n_n4426) & (!n_n2802) & (x37x) & (!x15051x)) + ((n_n4430) & (!n_n4426) & (!n_n2802) & (x37x) & (x15051x)) + ((n_n4430) & (!n_n4426) & (n_n2802) & (!x37x) & (!x15051x)) + ((n_n4430) & (!n_n4426) & (n_n2802) & (!x37x) & (x15051x)) + ((n_n4430) & (!n_n4426) & (n_n2802) & (x37x) & (!x15051x)) + ((n_n4430) & (!n_n4426) & (n_n2802) & (x37x) & (x15051x)) + ((n_n4430) & (n_n4426) & (!n_n2802) & (!x37x) & (!x15051x)) + ((n_n4430) & (n_n4426) & (!n_n2802) & (!x37x) & (x15051x)) + ((n_n4430) & (n_n4426) & (!n_n2802) & (x37x) & (!x15051x)) + ((n_n4430) & (n_n4426) & (!n_n2802) & (x37x) & (x15051x)) + ((n_n4430) & (n_n4426) & (n_n2802) & (!x37x) & (!x15051x)) + ((n_n4430) & (n_n4426) & (n_n2802) & (!x37x) & (x15051x)) + ((n_n4430) & (n_n4426) & (n_n2802) & (x37x) & (!x15051x)) + ((n_n4430) & (n_n4426) & (n_n2802) & (x37x) & (x15051x)));
	assign n_n4360 = (((i_9_) & (n_n536) & (n_n534) & (n_n500)));
	assign n_n4483 = (((!i_9_) & (n_n524) & (n_n455) & (n_n509)));
	assign n_n4837 = (((i_1_) & (i_2_) & (!i_0_) & (n_n535) & (x20x)));
	assign n_n5115 = (((!i_9_) & (n_n532) & (n_n509) & (n_n130)));
	assign n_n5175 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n130) & (x23x)));
	assign n_n5177 = (((!i_9_) & (n_n473) & (n_n534) & (n_n130)));
	assign n_n4933 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n260) & (x20x)));
	assign n_n4935 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n260) & (x23x)));
	assign x249x = (((!i_9_) & (!n_n528) & (n_n473) & (n_n260) & (n_n530)) + ((!i_9_) & (n_n528) & (n_n473) & (n_n260) & (!n_n530)) + ((!i_9_) & (n_n528) & (n_n473) & (n_n260) & (n_n530)) + ((i_9_) & (!n_n528) & (n_n473) & (n_n260) & (n_n530)) + ((i_9_) & (n_n528) & (n_n473) & (n_n260) & (!n_n530)) + ((i_9_) & (n_n528) & (n_n473) & (n_n260) & (n_n530)));
	assign n_n5108 = (((!i_5_) & (i_3_) & (i_4_) & (n_n522) & (x12x)));
	assign x290x = (((!i_9_) & (!n_n524) & (!n_n518) & (!n_n130) & (n_n5108)) + ((!i_9_) & (!n_n524) & (!n_n518) & (n_n130) & (n_n5108)) + ((!i_9_) & (!n_n524) & (n_n518) & (!n_n130) & (n_n5108)) + ((!i_9_) & (!n_n524) & (n_n518) & (n_n130) & (n_n5108)) + ((!i_9_) & (n_n524) & (!n_n518) & (!n_n130) & (n_n5108)) + ((!i_9_) & (n_n524) & (!n_n518) & (n_n130) & (n_n5108)) + ((!i_9_) & (n_n524) & (n_n518) & (!n_n130) & (n_n5108)) + ((!i_9_) & (n_n524) & (n_n518) & (n_n130) & (!n_n5108)) + ((!i_9_) & (n_n524) & (n_n518) & (n_n130) & (n_n5108)) + ((i_9_) & (!n_n524) & (!n_n518) & (!n_n130) & (n_n5108)) + ((i_9_) & (!n_n524) & (!n_n518) & (n_n130) & (n_n5108)) + ((i_9_) & (!n_n524) & (n_n518) & (!n_n130) & (n_n5108)) + ((i_9_) & (!n_n524) & (n_n518) & (n_n130) & (n_n5108)) + ((i_9_) & (n_n524) & (!n_n518) & (!n_n130) & (n_n5108)) + ((i_9_) & (n_n524) & (!n_n518) & (n_n130) & (n_n5108)) + ((i_9_) & (n_n524) & (n_n518) & (!n_n130) & (n_n5108)) + ((i_9_) & (n_n524) & (n_n518) & (n_n130) & (n_n5108)));
	assign n_n4144 = (((!n_n518) & (!x21x) & (!n_n130) & (!x20x) & (n_n5108)) + ((!n_n518) & (!x21x) & (!n_n130) & (x20x) & (n_n5108)) + ((!n_n518) & (!x21x) & (n_n130) & (!x20x) & (n_n5108)) + ((!n_n518) & (!x21x) & (n_n130) & (x20x) & (n_n5108)) + ((!n_n518) & (x21x) & (!n_n130) & (!x20x) & (n_n5108)) + ((!n_n518) & (x21x) & (!n_n130) & (x20x) & (n_n5108)) + ((!n_n518) & (x21x) & (n_n130) & (!x20x) & (n_n5108)) + ((!n_n518) & (x21x) & (n_n130) & (x20x) & (n_n5108)) + ((n_n518) & (!x21x) & (!n_n130) & (!x20x) & (n_n5108)) + ((n_n518) & (!x21x) & (!n_n130) & (x20x) & (n_n5108)) + ((n_n518) & (!x21x) & (n_n130) & (!x20x) & (n_n5108)) + ((n_n518) & (!x21x) & (n_n130) & (x20x) & (!n_n5108)) + ((n_n518) & (!x21x) & (n_n130) & (x20x) & (n_n5108)) + ((n_n518) & (x21x) & (!n_n130) & (!x20x) & (n_n5108)) + ((n_n518) & (x21x) & (!n_n130) & (x20x) & (n_n5108)) + ((n_n518) & (x21x) & (n_n130) & (!x20x) & (!n_n5108)) + ((n_n518) & (x21x) & (n_n130) & (!x20x) & (n_n5108)) + ((n_n518) & (x21x) & (n_n130) & (x20x) & (!n_n5108)) + ((n_n518) & (x21x) & (n_n130) & (x20x) & (n_n5108)));
	assign n_n5095 = (((i_5_) & (i_3_) & (i_4_) & (n_n130) & (x23x)));
	assign x34x = (((!n_n518) & (!n_n532) & (!x12x) & (n_n5095)) + ((!n_n518) & (!n_n532) & (x12x) & (n_n5095)) + ((!n_n518) & (n_n532) & (!x12x) & (n_n5095)) + ((!n_n518) & (n_n532) & (x12x) & (n_n5095)) + ((n_n518) & (!n_n532) & (!x12x) & (n_n5095)) + ((n_n518) & (!n_n532) & (x12x) & (n_n5095)) + ((n_n518) & (n_n532) & (!x12x) & (n_n5095)) + ((n_n518) & (n_n532) & (x12x) & (!n_n5095)) + ((n_n518) & (n_n532) & (x12x) & (n_n5095)));
	assign x289x = (((!i_9_) & (n_n518) & (!n_n526) & (n_n130) & (n_n530)) + ((!i_9_) & (n_n518) & (n_n526) & (n_n130) & (!n_n530)) + ((!i_9_) & (n_n518) & (n_n526) & (n_n130) & (n_n530)));
	assign n_n2210 = (((!n_n5096) & (!n_n5100) & (!n_n4144) & (!x34x) & (x289x)) + ((!n_n5096) & (!n_n5100) & (!n_n4144) & (x34x) & (!x289x)) + ((!n_n5096) & (!n_n5100) & (!n_n4144) & (x34x) & (x289x)) + ((!n_n5096) & (!n_n5100) & (n_n4144) & (!x34x) & (!x289x)) + ((!n_n5096) & (!n_n5100) & (n_n4144) & (!x34x) & (x289x)) + ((!n_n5096) & (!n_n5100) & (n_n4144) & (x34x) & (!x289x)) + ((!n_n5096) & (!n_n5100) & (n_n4144) & (x34x) & (x289x)) + ((!n_n5096) & (n_n5100) & (!n_n4144) & (!x34x) & (!x289x)) + ((!n_n5096) & (n_n5100) & (!n_n4144) & (!x34x) & (x289x)) + ((!n_n5096) & (n_n5100) & (!n_n4144) & (x34x) & (!x289x)) + ((!n_n5096) & (n_n5100) & (!n_n4144) & (x34x) & (x289x)) + ((!n_n5096) & (n_n5100) & (n_n4144) & (!x34x) & (!x289x)) + ((!n_n5096) & (n_n5100) & (n_n4144) & (!x34x) & (x289x)) + ((!n_n5096) & (n_n5100) & (n_n4144) & (x34x) & (!x289x)) + ((!n_n5096) & (n_n5100) & (n_n4144) & (x34x) & (x289x)) + ((n_n5096) & (!n_n5100) & (!n_n4144) & (!x34x) & (!x289x)) + ((n_n5096) & (!n_n5100) & (!n_n4144) & (!x34x) & (x289x)) + ((n_n5096) & (!n_n5100) & (!n_n4144) & (x34x) & (!x289x)) + ((n_n5096) & (!n_n5100) & (!n_n4144) & (x34x) & (x289x)) + ((n_n5096) & (!n_n5100) & (n_n4144) & (!x34x) & (!x289x)) + ((n_n5096) & (!n_n5100) & (n_n4144) & (!x34x) & (x289x)) + ((n_n5096) & (!n_n5100) & (n_n4144) & (x34x) & (!x289x)) + ((n_n5096) & (!n_n5100) & (n_n4144) & (x34x) & (x289x)) + ((n_n5096) & (n_n5100) & (!n_n4144) & (!x34x) & (!x289x)) + ((n_n5096) & (n_n5100) & (!n_n4144) & (!x34x) & (x289x)) + ((n_n5096) & (n_n5100) & (!n_n4144) & (x34x) & (!x289x)) + ((n_n5096) & (n_n5100) & (!n_n4144) & (x34x) & (x289x)) + ((n_n5096) & (n_n5100) & (n_n4144) & (!x34x) & (!x289x)) + ((n_n5096) & (n_n5100) & (n_n4144) & (!x34x) & (x289x)) + ((n_n5096) & (n_n5100) & (n_n4144) & (x34x) & (!x289x)) + ((n_n5096) & (n_n5100) & (n_n4144) & (x34x) & (x289x)));
	assign n_n4497 = (((!i_9_) & (n_n526) & (n_n455) & (n_n500)));
	assign x428x = (((!i_9_) & (n_n455) & (!n_n532) & (n_n534) & (n_n500)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n534) & (n_n500)) + ((i_9_) & (n_n455) & (n_n532) & (!n_n534) & (n_n500)) + ((i_9_) & (n_n455) & (n_n532) & (n_n534) & (n_n500)));
	assign n_n3883 = (((!i_9_) & (n_n455) & (!n_n532) & (n_n534) & (n_n500)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n534) & (n_n500)) + ((i_9_) & (n_n455) & (!n_n532) & (n_n534) & (n_n500)) + ((i_9_) & (n_n455) & (n_n532) & (!n_n534) & (n_n500)) + ((i_9_) & (n_n455) & (n_n532) & (n_n534) & (n_n500)));
	assign n_n4498 = (((i_9_) & (n_n524) & (n_n455) & (n_n500)));
	assign x65x = (((!i_9_) & (n_n524) & (n_n455) & (n_n500)) + ((i_9_) & (n_n524) & (n_n455) & (n_n500)));
	assign x66x = (((!i_9_) & (n_n455) & (n_n528) & (n_n500)) + ((i_9_) & (n_n455) & (n_n528) & (n_n500)));
	assign x78x = (((!i_9_) & (n_n455) & (n_n532) & (n_n509) & (!n_n530)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n509) & (n_n530)) + ((i_9_) & (n_n455) & (!n_n532) & (n_n509) & (n_n530)) + ((i_9_) & (n_n455) & (n_n532) & (n_n509) & (n_n530)));
	assign n_n4477 = (((!i_9_) & (n_n455) & (n_n509) & (n_n530)));
	assign n_n4254 = (((!i_9_) & (n_n455) & (!n_n532) & (n_n509) & (n_n530)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n509) & (!n_n530)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n509) & (n_n530)) + ((i_9_) & (n_n455) & (!n_n532) & (n_n509) & (n_n530)) + ((i_9_) & (n_n455) & (n_n532) & (n_n509) & (n_n530)));
	assign x70x = (((!i_9_) & (!n_n524) & (n_n455) & (n_n509) & (x20x)) + ((!i_9_) & (n_n524) & (n_n455) & (n_n509) & (!x20x)) + ((!i_9_) & (n_n524) & (n_n455) & (n_n509) & (x20x)) + ((i_9_) & (!n_n524) & (n_n455) & (n_n509) & (x20x)) + ((i_9_) & (n_n524) & (n_n455) & (n_n509) & (x20x)));
	assign x184x = (((i_7_) & (!i_8_) & (!i_6_) & (x13x) & (n_n509)) + ((i_7_) & (i_8_) & (!i_6_) & (x13x) & (n_n509)));
	assign x38x = (((!i_9_) & (!n_n528) & (n_n260) & (n_n535) & (n_n530)) + ((!i_9_) & (n_n528) & (n_n260) & (n_n535) & (n_n530)) + ((i_9_) & (n_n528) & (n_n260) & (n_n535) & (!n_n530)) + ((i_9_) & (n_n528) & (n_n260) & (n_n535) & (n_n530)));
	assign x388x = (((!i_9_) & (!n_n528) & (n_n260) & (n_n535) & (n_n530)) + ((!i_9_) & (n_n528) & (n_n260) & (n_n535) & (!n_n530)) + ((!i_9_) & (n_n528) & (n_n260) & (n_n535) & (n_n530)) + ((i_9_) & (!n_n528) & (n_n260) & (n_n535) & (n_n530)) + ((i_9_) & (n_n528) & (n_n260) & (n_n535) & (!n_n530)) + ((i_9_) & (n_n528) & (n_n260) & (n_n535) & (n_n530)));
	assign x176x = (((!i_9_) & (n_n518) & (n_n260) & (n_n530)) + ((i_9_) & (n_n518) & (n_n260) & (n_n530)));
	assign n_n4823 = (((!i_1_) & (!i_2_) & (i_0_) & (x23x) & (n_n464)));
	assign n_n4820 = (((i_9_) & (n_n325) & (n_n522) & (n_n464)));
	assign n_n4810 = (((i_9_) & (n_n532) & (n_n325) & (n_n464)));
	assign x186x = (((!i_9_) & (!n_n524) & (n_n325) & (x20x) & (n_n464)) + ((!i_9_) & (n_n524) & (n_n325) & (!x20x) & (n_n464)) + ((!i_9_) & (n_n524) & (n_n325) & (x20x) & (n_n464)) + ((i_9_) & (!n_n524) & (n_n325) & (x20x) & (n_n464)) + ((i_9_) & (n_n524) & (n_n325) & (x20x) & (n_n464)));
	assign x16522x = (((!n_n4415) & (!n_n4408) & (!n_n4414) & (!n_n4411) & (n_n4412)) + ((!n_n4415) & (!n_n4408) & (!n_n4414) & (n_n4411) & (!n_n4412)) + ((!n_n4415) & (!n_n4408) & (!n_n4414) & (n_n4411) & (n_n4412)) + ((!n_n4415) & (!n_n4408) & (n_n4414) & (!n_n4411) & (!n_n4412)) + ((!n_n4415) & (!n_n4408) & (n_n4414) & (!n_n4411) & (n_n4412)) + ((!n_n4415) & (!n_n4408) & (n_n4414) & (n_n4411) & (!n_n4412)) + ((!n_n4415) & (!n_n4408) & (n_n4414) & (n_n4411) & (n_n4412)) + ((!n_n4415) & (n_n4408) & (!n_n4414) & (!n_n4411) & (!n_n4412)) + ((!n_n4415) & (n_n4408) & (!n_n4414) & (!n_n4411) & (n_n4412)) + ((!n_n4415) & (n_n4408) & (!n_n4414) & (n_n4411) & (!n_n4412)) + ((!n_n4415) & (n_n4408) & (!n_n4414) & (n_n4411) & (n_n4412)) + ((!n_n4415) & (n_n4408) & (n_n4414) & (!n_n4411) & (!n_n4412)) + ((!n_n4415) & (n_n4408) & (n_n4414) & (!n_n4411) & (n_n4412)) + ((!n_n4415) & (n_n4408) & (n_n4414) & (n_n4411) & (!n_n4412)) + ((!n_n4415) & (n_n4408) & (n_n4414) & (n_n4411) & (n_n4412)) + ((n_n4415) & (!n_n4408) & (!n_n4414) & (!n_n4411) & (!n_n4412)) + ((n_n4415) & (!n_n4408) & (!n_n4414) & (!n_n4411) & (n_n4412)) + ((n_n4415) & (!n_n4408) & (!n_n4414) & (n_n4411) & (!n_n4412)) + ((n_n4415) & (!n_n4408) & (!n_n4414) & (n_n4411) & (n_n4412)) + ((n_n4415) & (!n_n4408) & (n_n4414) & (!n_n4411) & (!n_n4412)) + ((n_n4415) & (!n_n4408) & (n_n4414) & (!n_n4411) & (n_n4412)) + ((n_n4415) & (!n_n4408) & (n_n4414) & (n_n4411) & (!n_n4412)) + ((n_n4415) & (!n_n4408) & (n_n4414) & (n_n4411) & (n_n4412)) + ((n_n4415) & (n_n4408) & (!n_n4414) & (!n_n4411) & (!n_n4412)) + ((n_n4415) & (n_n4408) & (!n_n4414) & (!n_n4411) & (n_n4412)) + ((n_n4415) & (n_n4408) & (!n_n4414) & (n_n4411) & (!n_n4412)) + ((n_n4415) & (n_n4408) & (!n_n4414) & (n_n4411) & (n_n4412)) + ((n_n4415) & (n_n4408) & (n_n4414) & (!n_n4411) & (!n_n4412)) + ((n_n4415) & (n_n4408) & (n_n4414) & (!n_n4411) & (n_n4412)) + ((n_n4415) & (n_n4408) & (n_n4414) & (n_n4411) & (!n_n4412)) + ((n_n4415) & (n_n4408) & (n_n4414) & (n_n4411) & (n_n4412)));
	assign n_n2263 = (((!x16522x) & (!n_n4419) & (!n_n4409) & (!n_n4417) & (n_n4410)) + ((!x16522x) & (!n_n4419) & (!n_n4409) & (n_n4417) & (!n_n4410)) + ((!x16522x) & (!n_n4419) & (!n_n4409) & (n_n4417) & (n_n4410)) + ((!x16522x) & (!n_n4419) & (n_n4409) & (!n_n4417) & (!n_n4410)) + ((!x16522x) & (!n_n4419) & (n_n4409) & (!n_n4417) & (n_n4410)) + ((!x16522x) & (!n_n4419) & (n_n4409) & (n_n4417) & (!n_n4410)) + ((!x16522x) & (!n_n4419) & (n_n4409) & (n_n4417) & (n_n4410)) + ((!x16522x) & (n_n4419) & (!n_n4409) & (!n_n4417) & (!n_n4410)) + ((!x16522x) & (n_n4419) & (!n_n4409) & (!n_n4417) & (n_n4410)) + ((!x16522x) & (n_n4419) & (!n_n4409) & (n_n4417) & (!n_n4410)) + ((!x16522x) & (n_n4419) & (!n_n4409) & (n_n4417) & (n_n4410)) + ((!x16522x) & (n_n4419) & (n_n4409) & (!n_n4417) & (!n_n4410)) + ((!x16522x) & (n_n4419) & (n_n4409) & (!n_n4417) & (n_n4410)) + ((!x16522x) & (n_n4419) & (n_n4409) & (n_n4417) & (!n_n4410)) + ((!x16522x) & (n_n4419) & (n_n4409) & (n_n4417) & (n_n4410)) + ((x16522x) & (!n_n4419) & (!n_n4409) & (!n_n4417) & (!n_n4410)) + ((x16522x) & (!n_n4419) & (!n_n4409) & (!n_n4417) & (n_n4410)) + ((x16522x) & (!n_n4419) & (!n_n4409) & (n_n4417) & (!n_n4410)) + ((x16522x) & (!n_n4419) & (!n_n4409) & (n_n4417) & (n_n4410)) + ((x16522x) & (!n_n4419) & (n_n4409) & (!n_n4417) & (!n_n4410)) + ((x16522x) & (!n_n4419) & (n_n4409) & (!n_n4417) & (n_n4410)) + ((x16522x) & (!n_n4419) & (n_n4409) & (n_n4417) & (!n_n4410)) + ((x16522x) & (!n_n4419) & (n_n4409) & (n_n4417) & (n_n4410)) + ((x16522x) & (n_n4419) & (!n_n4409) & (!n_n4417) & (!n_n4410)) + ((x16522x) & (n_n4419) & (!n_n4409) & (!n_n4417) & (n_n4410)) + ((x16522x) & (n_n4419) & (!n_n4409) & (n_n4417) & (!n_n4410)) + ((x16522x) & (n_n4419) & (!n_n4409) & (n_n4417) & (n_n4410)) + ((x16522x) & (n_n4419) & (n_n4409) & (!n_n4417) & (!n_n4410)) + ((x16522x) & (n_n4419) & (n_n4409) & (!n_n4417) & (n_n4410)) + ((x16522x) & (n_n4419) & (n_n4409) & (n_n4417) & (!n_n4410)) + ((x16522x) & (n_n4419) & (n_n4409) & (n_n4417) & (n_n4410)));
	assign x16526x = (((!i_9_) & (!n_n536) & (!n_n4440) & (!x516x) & (x215x)) + ((!i_9_) & (!n_n536) & (!n_n4440) & (x516x) & (x215x)) + ((!i_9_) & (!n_n536) & (n_n4440) & (!x516x) & (!x215x)) + ((!i_9_) & (!n_n536) & (n_n4440) & (!x516x) & (x215x)) + ((!i_9_) & (!n_n536) & (n_n4440) & (x516x) & (!x215x)) + ((!i_9_) & (!n_n536) & (n_n4440) & (x516x) & (x215x)) + ((!i_9_) & (n_n536) & (!n_n4440) & (!x516x) & (x215x)) + ((!i_9_) & (n_n536) & (!n_n4440) & (x516x) & (x215x)) + ((!i_9_) & (n_n536) & (n_n4440) & (!x516x) & (!x215x)) + ((!i_9_) & (n_n536) & (n_n4440) & (!x516x) & (x215x)) + ((!i_9_) & (n_n536) & (n_n4440) & (x516x) & (!x215x)) + ((!i_9_) & (n_n536) & (n_n4440) & (x516x) & (x215x)) + ((i_9_) & (!n_n536) & (!n_n4440) & (!x516x) & (x215x)) + ((i_9_) & (!n_n536) & (!n_n4440) & (x516x) & (x215x)) + ((i_9_) & (!n_n536) & (n_n4440) & (!x516x) & (!x215x)) + ((i_9_) & (!n_n536) & (n_n4440) & (!x516x) & (x215x)) + ((i_9_) & (!n_n536) & (n_n4440) & (x516x) & (!x215x)) + ((i_9_) & (!n_n536) & (n_n4440) & (x516x) & (x215x)) + ((i_9_) & (n_n536) & (!n_n4440) & (!x516x) & (x215x)) + ((i_9_) & (n_n536) & (!n_n4440) & (x516x) & (!x215x)) + ((i_9_) & (n_n536) & (!n_n4440) & (x516x) & (x215x)) + ((i_9_) & (n_n536) & (n_n4440) & (!x516x) & (!x215x)) + ((i_9_) & (n_n536) & (n_n4440) & (!x516x) & (x215x)) + ((i_9_) & (n_n536) & (n_n4440) & (x516x) & (!x215x)) + ((i_9_) & (n_n536) & (n_n4440) & (x516x) & (x215x)));
	assign x16527x = (((!x98x) & (!x23x) & (!x496x) & (!n_n4430) & (n_n4428)) + ((!x98x) & (!x23x) & (!x496x) & (n_n4430) & (!n_n4428)) + ((!x98x) & (!x23x) & (!x496x) & (n_n4430) & (n_n4428)) + ((!x98x) & (!x23x) & (x496x) & (!n_n4430) & (n_n4428)) + ((!x98x) & (!x23x) & (x496x) & (n_n4430) & (!n_n4428)) + ((!x98x) & (!x23x) & (x496x) & (n_n4430) & (n_n4428)) + ((!x98x) & (x23x) & (!x496x) & (!n_n4430) & (n_n4428)) + ((!x98x) & (x23x) & (!x496x) & (n_n4430) & (!n_n4428)) + ((!x98x) & (x23x) & (!x496x) & (n_n4430) & (n_n4428)) + ((!x98x) & (x23x) & (x496x) & (!n_n4430) & (!n_n4428)) + ((!x98x) & (x23x) & (x496x) & (!n_n4430) & (n_n4428)) + ((!x98x) & (x23x) & (x496x) & (n_n4430) & (!n_n4428)) + ((!x98x) & (x23x) & (x496x) & (n_n4430) & (n_n4428)) + ((x98x) & (!x23x) & (!x496x) & (!n_n4430) & (!n_n4428)) + ((x98x) & (!x23x) & (!x496x) & (!n_n4430) & (n_n4428)) + ((x98x) & (!x23x) & (!x496x) & (n_n4430) & (!n_n4428)) + ((x98x) & (!x23x) & (!x496x) & (n_n4430) & (n_n4428)) + ((x98x) & (!x23x) & (x496x) & (!n_n4430) & (!n_n4428)) + ((x98x) & (!x23x) & (x496x) & (!n_n4430) & (n_n4428)) + ((x98x) & (!x23x) & (x496x) & (n_n4430) & (!n_n4428)) + ((x98x) & (!x23x) & (x496x) & (n_n4430) & (n_n4428)) + ((x98x) & (x23x) & (!x496x) & (!n_n4430) & (!n_n4428)) + ((x98x) & (x23x) & (!x496x) & (!n_n4430) & (n_n4428)) + ((x98x) & (x23x) & (!x496x) & (n_n4430) & (!n_n4428)) + ((x98x) & (x23x) & (!x496x) & (n_n4430) & (n_n4428)) + ((x98x) & (x23x) & (x496x) & (!n_n4430) & (!n_n4428)) + ((x98x) & (x23x) & (x496x) & (!n_n4430) & (n_n4428)) + ((x98x) & (x23x) & (x496x) & (n_n4430) & (!n_n4428)) + ((x98x) & (x23x) & (x496x) & (n_n4430) & (n_n4428)));
	assign x16532x = (((!n_n4401) & (!n_n4393) & (!n_n4398) & (!n_n4395) & (n_n4402)) + ((!n_n4401) & (!n_n4393) & (!n_n4398) & (n_n4395) & (!n_n4402)) + ((!n_n4401) & (!n_n4393) & (!n_n4398) & (n_n4395) & (n_n4402)) + ((!n_n4401) & (!n_n4393) & (n_n4398) & (!n_n4395) & (!n_n4402)) + ((!n_n4401) & (!n_n4393) & (n_n4398) & (!n_n4395) & (n_n4402)) + ((!n_n4401) & (!n_n4393) & (n_n4398) & (n_n4395) & (!n_n4402)) + ((!n_n4401) & (!n_n4393) & (n_n4398) & (n_n4395) & (n_n4402)) + ((!n_n4401) & (n_n4393) & (!n_n4398) & (!n_n4395) & (!n_n4402)) + ((!n_n4401) & (n_n4393) & (!n_n4398) & (!n_n4395) & (n_n4402)) + ((!n_n4401) & (n_n4393) & (!n_n4398) & (n_n4395) & (!n_n4402)) + ((!n_n4401) & (n_n4393) & (!n_n4398) & (n_n4395) & (n_n4402)) + ((!n_n4401) & (n_n4393) & (n_n4398) & (!n_n4395) & (!n_n4402)) + ((!n_n4401) & (n_n4393) & (n_n4398) & (!n_n4395) & (n_n4402)) + ((!n_n4401) & (n_n4393) & (n_n4398) & (n_n4395) & (!n_n4402)) + ((!n_n4401) & (n_n4393) & (n_n4398) & (n_n4395) & (n_n4402)) + ((n_n4401) & (!n_n4393) & (!n_n4398) & (!n_n4395) & (!n_n4402)) + ((n_n4401) & (!n_n4393) & (!n_n4398) & (!n_n4395) & (n_n4402)) + ((n_n4401) & (!n_n4393) & (!n_n4398) & (n_n4395) & (!n_n4402)) + ((n_n4401) & (!n_n4393) & (!n_n4398) & (n_n4395) & (n_n4402)) + ((n_n4401) & (!n_n4393) & (n_n4398) & (!n_n4395) & (!n_n4402)) + ((n_n4401) & (!n_n4393) & (n_n4398) & (!n_n4395) & (n_n4402)) + ((n_n4401) & (!n_n4393) & (n_n4398) & (n_n4395) & (!n_n4402)) + ((n_n4401) & (!n_n4393) & (n_n4398) & (n_n4395) & (n_n4402)) + ((n_n4401) & (n_n4393) & (!n_n4398) & (!n_n4395) & (!n_n4402)) + ((n_n4401) & (n_n4393) & (!n_n4398) & (!n_n4395) & (n_n4402)) + ((n_n4401) & (n_n4393) & (!n_n4398) & (n_n4395) & (!n_n4402)) + ((n_n4401) & (n_n4393) & (!n_n4398) & (n_n4395) & (n_n4402)) + ((n_n4401) & (n_n4393) & (n_n4398) & (!n_n4395) & (!n_n4402)) + ((n_n4401) & (n_n4393) & (n_n4398) & (!n_n4395) & (n_n4402)) + ((n_n4401) & (n_n4393) & (n_n4398) & (n_n4395) & (!n_n4402)) + ((n_n4401) & (n_n4393) & (n_n4398) & (n_n4395) & (n_n4402)));
	assign x16533x = (((!n_n4403) & (!n_n4392) & (!n_n4396) & (!n_n4399) & (x16532x)) + ((!n_n4403) & (!n_n4392) & (!n_n4396) & (n_n4399) & (!x16532x)) + ((!n_n4403) & (!n_n4392) & (!n_n4396) & (n_n4399) & (x16532x)) + ((!n_n4403) & (!n_n4392) & (n_n4396) & (!n_n4399) & (!x16532x)) + ((!n_n4403) & (!n_n4392) & (n_n4396) & (!n_n4399) & (x16532x)) + ((!n_n4403) & (!n_n4392) & (n_n4396) & (n_n4399) & (!x16532x)) + ((!n_n4403) & (!n_n4392) & (n_n4396) & (n_n4399) & (x16532x)) + ((!n_n4403) & (n_n4392) & (!n_n4396) & (!n_n4399) & (!x16532x)) + ((!n_n4403) & (n_n4392) & (!n_n4396) & (!n_n4399) & (x16532x)) + ((!n_n4403) & (n_n4392) & (!n_n4396) & (n_n4399) & (!x16532x)) + ((!n_n4403) & (n_n4392) & (!n_n4396) & (n_n4399) & (x16532x)) + ((!n_n4403) & (n_n4392) & (n_n4396) & (!n_n4399) & (!x16532x)) + ((!n_n4403) & (n_n4392) & (n_n4396) & (!n_n4399) & (x16532x)) + ((!n_n4403) & (n_n4392) & (n_n4396) & (n_n4399) & (!x16532x)) + ((!n_n4403) & (n_n4392) & (n_n4396) & (n_n4399) & (x16532x)) + ((n_n4403) & (!n_n4392) & (!n_n4396) & (!n_n4399) & (!x16532x)) + ((n_n4403) & (!n_n4392) & (!n_n4396) & (!n_n4399) & (x16532x)) + ((n_n4403) & (!n_n4392) & (!n_n4396) & (n_n4399) & (!x16532x)) + ((n_n4403) & (!n_n4392) & (!n_n4396) & (n_n4399) & (x16532x)) + ((n_n4403) & (!n_n4392) & (n_n4396) & (!n_n4399) & (!x16532x)) + ((n_n4403) & (!n_n4392) & (n_n4396) & (!n_n4399) & (x16532x)) + ((n_n4403) & (!n_n4392) & (n_n4396) & (n_n4399) & (!x16532x)) + ((n_n4403) & (!n_n4392) & (n_n4396) & (n_n4399) & (x16532x)) + ((n_n4403) & (n_n4392) & (!n_n4396) & (!n_n4399) & (!x16532x)) + ((n_n4403) & (n_n4392) & (!n_n4396) & (!n_n4399) & (x16532x)) + ((n_n4403) & (n_n4392) & (!n_n4396) & (n_n4399) & (!x16532x)) + ((n_n4403) & (n_n4392) & (!n_n4396) & (n_n4399) & (x16532x)) + ((n_n4403) & (n_n4392) & (n_n4396) & (!n_n4399) & (!x16532x)) + ((n_n4403) & (n_n4392) & (n_n4396) & (!n_n4399) & (x16532x)) + ((n_n4403) & (n_n4392) & (n_n4396) & (n_n4399) & (!x16532x)) + ((n_n4403) & (n_n4392) & (n_n4396) & (n_n4399) & (x16532x)));
	assign n_n2446 = (((!i_9_) & (n_n536) & (n_n535) & (!n_n522) & (n_n520)) + ((!i_9_) & (n_n536) & (n_n535) & (n_n522) & (n_n520)) + ((i_9_) & (n_n536) & (n_n535) & (!n_n522) & (n_n520)) + ((i_9_) & (n_n536) & (n_n535) & (n_n522) & (!n_n520)) + ((i_9_) & (n_n536) & (n_n535) & (n_n522) & (n_n520)));
	assign x399x = (((!i_9_) & (n_n536) & (n_n528) & (n_n509)) + ((i_9_) & (n_n536) & (n_n528) & (n_n509)));
	assign x22197x = (((!x67x) & (!n_n4353) & (!n_n4354) & (!n_n4349)));
	assign n_n4336 = (((i_9_) & (n_n536) & (n_n518) & (n_n526)));
	assign n_n2443 = (((!n_n536) & (!n_n518) & (!x21x) & (!n_n4337) & (n_n4340)) + ((!n_n536) & (!n_n518) & (!x21x) & (n_n4337) & (!n_n4340)) + ((!n_n536) & (!n_n518) & (!x21x) & (n_n4337) & (n_n4340)) + ((!n_n536) & (!n_n518) & (x21x) & (!n_n4337) & (n_n4340)) + ((!n_n536) & (!n_n518) & (x21x) & (n_n4337) & (!n_n4340)) + ((!n_n536) & (!n_n518) & (x21x) & (n_n4337) & (n_n4340)) + ((!n_n536) & (n_n518) & (!x21x) & (!n_n4337) & (n_n4340)) + ((!n_n536) & (n_n518) & (!x21x) & (n_n4337) & (!n_n4340)) + ((!n_n536) & (n_n518) & (!x21x) & (n_n4337) & (n_n4340)) + ((!n_n536) & (n_n518) & (x21x) & (!n_n4337) & (n_n4340)) + ((!n_n536) & (n_n518) & (x21x) & (n_n4337) & (!n_n4340)) + ((!n_n536) & (n_n518) & (x21x) & (n_n4337) & (n_n4340)) + ((n_n536) & (!n_n518) & (!x21x) & (!n_n4337) & (n_n4340)) + ((n_n536) & (!n_n518) & (!x21x) & (n_n4337) & (!n_n4340)) + ((n_n536) & (!n_n518) & (!x21x) & (n_n4337) & (n_n4340)) + ((n_n536) & (!n_n518) & (x21x) & (!n_n4337) & (n_n4340)) + ((n_n536) & (!n_n518) & (x21x) & (n_n4337) & (!n_n4340)) + ((n_n536) & (!n_n518) & (x21x) & (n_n4337) & (n_n4340)) + ((n_n536) & (n_n518) & (!x21x) & (!n_n4337) & (n_n4340)) + ((n_n536) & (n_n518) & (!x21x) & (n_n4337) & (!n_n4340)) + ((n_n536) & (n_n518) & (!x21x) & (n_n4337) & (n_n4340)) + ((n_n536) & (n_n518) & (x21x) & (!n_n4337) & (!n_n4340)) + ((n_n536) & (n_n518) & (x21x) & (!n_n4337) & (n_n4340)) + ((n_n536) & (n_n518) & (x21x) & (n_n4337) & (!n_n4340)) + ((n_n536) & (n_n518) & (x21x) & (n_n4337) & (n_n4340)));
	assign n_n2445 = (((!i_9_) & (n_n536) & (n_n518) & (n_n532) & (!n_n534)) + ((!i_9_) & (n_n536) & (n_n518) & (n_n532) & (n_n534)) + ((i_9_) & (n_n536) & (n_n518) & (!n_n532) & (n_n534)) + ((i_9_) & (n_n536) & (n_n518) & (n_n532) & (!n_n534)) + ((i_9_) & (n_n536) & (n_n518) & (n_n532) & (n_n534)));
	assign n_n4321 = (((!i_9_) & (n_n536) & (n_n526) & (n_n535)));
	assign x171x = (((!i_9_) & (n_n536) & (!n_n526) & (n_n528) & (n_n535)) + ((!i_9_) & (n_n536) & (n_n526) & (!n_n528) & (n_n535)) + ((!i_9_) & (n_n536) & (n_n526) & (n_n528) & (n_n535)));
	assign n_n4332 = (((i_9_) & (n_n536) & (n_n518) & (n_n530)));
	assign x198x = (((!i_9_) & (n_n536) & (n_n518) & (n_n530)) + ((i_9_) & (n_n536) & (n_n518) & (n_n530)));
	assign x283x = (((!i_9_) & (n_n536) & (n_n532) & (n_n535)) + ((i_9_) & (n_n536) & (n_n532) & (n_n535)));
	assign n_n4275 = (((!i_9_) & (n_n536) & (!n_n528) & (n_n500) & (n_n530)) + ((!i_9_) & (n_n536) & (n_n528) & (n_n500) & (n_n530)) + ((i_9_) & (n_n536) & (!n_n528) & (n_n500) & (n_n530)) + ((i_9_) & (n_n536) & (n_n528) & (n_n500) & (!n_n530)) + ((i_9_) & (n_n536) & (n_n528) & (n_n500) & (n_n530)));
	assign x74x = (((!i_9_) & (n_n536) & (n_n524) & (n_n509) & (!n_n522)) + ((!i_9_) & (n_n536) & (n_n524) & (n_n509) & (n_n522)) + ((i_9_) & (n_n536) & (!n_n524) & (n_n509) & (n_n522)) + ((i_9_) & (n_n536) & (n_n524) & (n_n509) & (n_n522)));
	assign x345x = (((i_9_) & (n_n536) & (!n_n532) & (n_n534) & (n_n500)) + ((i_9_) & (n_n536) & (n_n532) & (!n_n534) & (n_n500)) + ((i_9_) & (n_n536) & (n_n532) & (n_n534) & (n_n500)));
	assign n_n2435 = (((!i_9_) & (n_n536) & (!n_n522) & (n_n491) & (n_n520)) + ((!i_9_) & (n_n536) & (n_n522) & (n_n491) & (n_n520)) + ((i_9_) & (n_n536) & (!n_n522) & (n_n491) & (n_n520)) + ((i_9_) & (n_n536) & (n_n522) & (n_n491) & (!n_n520)) + ((i_9_) & (n_n536) & (n_n522) & (n_n491) & (n_n520)));
	assign n_n3903 = (((!i_9_) & (n_n536) & (!n_n524) & (n_n526) & (n_n491)) + ((!i_9_) & (n_n536) & (n_n524) & (n_n526) & (n_n491)) + ((i_9_) & (n_n536) & (!n_n524) & (n_n526) & (n_n491)) + ((i_9_) & (n_n536) & (n_n524) & (!n_n526) & (n_n491)) + ((i_9_) & (n_n536) & (n_n524) & (n_n526) & (n_n491)));
	assign x14460x = (((!i_9_) & (n_n536) & (!n_n528) & (n_n491) & (n_n530)) + ((!i_9_) & (n_n536) & (n_n528) & (n_n491) & (!n_n530)) + ((!i_9_) & (n_n536) & (n_n528) & (n_n491) & (n_n530)));
	assign x282x = (((!i_9_) & (n_n536) & (!n_n524) & (n_n526) & (n_n500)) + ((!i_9_) & (n_n536) & (n_n524) & (n_n526) & (n_n500)) + ((i_9_) & (n_n536) & (!n_n524) & (n_n526) & (n_n500)) + ((i_9_) & (n_n536) & (n_n524) & (!n_n526) & (n_n500)) + ((i_9_) & (n_n536) & (n_n524) & (n_n526) & (n_n500)));
	assign x300x = (((!i_9_) & (n_n536) & (n_n524) & (!n_n522) & (n_n500)) + ((!i_9_) & (n_n536) & (n_n524) & (n_n522) & (n_n500)) + ((i_9_) & (n_n536) & (!n_n524) & (n_n522) & (n_n500)) + ((i_9_) & (n_n536) & (n_n524) & (n_n522) & (n_n500)));
	assign n_n4377 = (((!i_9_) & (n_n536) & (n_n534) & (n_n491)));
	assign n_n4376 = (((i_9_) & (n_n536) & (n_n534) & (n_n491)));
	assign x423x = (((!i_9_) & (n_n536) & (n_n534) & (n_n491)) + ((i_9_) & (n_n536) & (n_n534) & (n_n491)));
	assign n_n4503 = (((i_1_) & (!i_2_) & (i_0_) & (x23x) & (n_n500)));
	assign n_n4502 = (((i_9_) & (n_n455) & (n_n520) & (n_n500)));
	assign n_n4500 = (((i_9_) & (n_n455) & (n_n522) & (n_n500)));
	assign n_n4510 = (((i_9_) & (n_n455) & (n_n528) & (n_n491)));
	assign x22063x = (((!n_n4512) & (!n_n4522) & (!n_n4531) & (!n_n4517)));
	assign n_n4505 = (((!i_9_) & (n_n455) & (n_n534) & (n_n491)));
	assign x189x = (((!i_9_) & (n_n455) & (!n_n532) & (n_n534) & (n_n491)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n534) & (n_n491)) + ((i_9_) & (n_n455) & (n_n532) & (!n_n534) & (n_n491)) + ((i_9_) & (n_n455) & (n_n532) & (n_n534) & (n_n491)));
	assign x387x = (((!i_9_) & (n_n455) & (!n_n532) & (n_n491) & (n_n530)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n491) & (!n_n530)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n491) & (n_n530)) + ((i_9_) & (n_n455) & (!n_n532) & (n_n491) & (n_n530)) + ((i_9_) & (n_n455) & (n_n532) & (n_n491) & (n_n530)));
	assign n_n4546 = (((i_9_) & (n_n524) & (n_n455) & (n_n473)));
	assign n_n4555 = (((!i_9_) & (n_n455) & (n_n532) & (n_n464)));
	assign x455x = (((!i_9_) & (n_n524) & (n_n455) & (n_n464)) + ((i_9_) & (n_n524) & (n_n455) & (n_n464)));
	assign x121x = (((!i_9_) & (n_n390) & (!n_n532) & (n_n534) & (n_n535)) + ((!i_9_) & (n_n390) & (n_n532) & (n_n534) & (n_n535)) + ((i_9_) & (n_n390) & (n_n532) & (!n_n534) & (n_n535)) + ((i_9_) & (n_n390) & (n_n532) & (n_n534) & (n_n535)));
	assign n_n4239 = (((!i_9_) & (!n_n455) & (!n_n520) & (!n_n464) & (x471x)) + ((!i_9_) & (!n_n455) & (!n_n520) & (n_n464) & (x471x)) + ((!i_9_) & (!n_n455) & (n_n520) & (!n_n464) & (x471x)) + ((!i_9_) & (!n_n455) & (n_n520) & (n_n464) & (x471x)) + ((!i_9_) & (n_n455) & (!n_n520) & (!n_n464) & (x471x)) + ((!i_9_) & (n_n455) & (!n_n520) & (n_n464) & (x471x)) + ((!i_9_) & (n_n455) & (n_n520) & (!n_n464) & (x471x)) + ((!i_9_) & (n_n455) & (n_n520) & (n_n464) & (x471x)) + ((i_9_) & (!n_n455) & (!n_n520) & (!n_n464) & (x471x)) + ((i_9_) & (!n_n455) & (!n_n520) & (n_n464) & (x471x)) + ((i_9_) & (!n_n455) & (n_n520) & (!n_n464) & (x471x)) + ((i_9_) & (!n_n455) & (n_n520) & (n_n464) & (x471x)) + ((i_9_) & (n_n455) & (!n_n520) & (!n_n464) & (x471x)) + ((i_9_) & (n_n455) & (!n_n520) & (n_n464) & (x471x)) + ((i_9_) & (n_n455) & (n_n520) & (!n_n464) & (x471x)) + ((i_9_) & (n_n455) & (n_n520) & (n_n464) & (!x471x)) + ((i_9_) & (n_n455) & (n_n520) & (n_n464) & (x471x)));
	assign n_n4580 = (((i_9_) & (n_n390) & (n_n535) & (n_n522)));
	assign n_n2401 = (((!i_9_) & (n_n518) & (n_n390) & (!n_n532) & (n_n534)) + ((!i_9_) & (n_n518) & (n_n390) & (n_n532) & (!n_n534)) + ((!i_9_) & (n_n518) & (n_n390) & (n_n532) & (n_n534)) + ((i_9_) & (n_n518) & (n_n390) & (n_n532) & (!n_n534)) + ((i_9_) & (n_n518) & (n_n390) & (n_n532) & (n_n534)));
	assign x16622x = (((!n_n4593) & (!n_n4590) & (!x172x) & (!x365x) & (n_n2401)) + ((!n_n4593) & (!n_n4590) & (!x172x) & (x365x) & (!n_n2401)) + ((!n_n4593) & (!n_n4590) & (!x172x) & (x365x) & (n_n2401)) + ((!n_n4593) & (!n_n4590) & (x172x) & (!x365x) & (!n_n2401)) + ((!n_n4593) & (!n_n4590) & (x172x) & (!x365x) & (n_n2401)) + ((!n_n4593) & (!n_n4590) & (x172x) & (x365x) & (!n_n2401)) + ((!n_n4593) & (!n_n4590) & (x172x) & (x365x) & (n_n2401)) + ((!n_n4593) & (n_n4590) & (!x172x) & (!x365x) & (!n_n2401)) + ((!n_n4593) & (n_n4590) & (!x172x) & (!x365x) & (n_n2401)) + ((!n_n4593) & (n_n4590) & (!x172x) & (x365x) & (!n_n2401)) + ((!n_n4593) & (n_n4590) & (!x172x) & (x365x) & (n_n2401)) + ((!n_n4593) & (n_n4590) & (x172x) & (!x365x) & (!n_n2401)) + ((!n_n4593) & (n_n4590) & (x172x) & (!x365x) & (n_n2401)) + ((!n_n4593) & (n_n4590) & (x172x) & (x365x) & (!n_n2401)) + ((!n_n4593) & (n_n4590) & (x172x) & (x365x) & (n_n2401)) + ((n_n4593) & (!n_n4590) & (!x172x) & (!x365x) & (!n_n2401)) + ((n_n4593) & (!n_n4590) & (!x172x) & (!x365x) & (n_n2401)) + ((n_n4593) & (!n_n4590) & (!x172x) & (x365x) & (!n_n2401)) + ((n_n4593) & (!n_n4590) & (!x172x) & (x365x) & (n_n2401)) + ((n_n4593) & (!n_n4590) & (x172x) & (!x365x) & (!n_n2401)) + ((n_n4593) & (!n_n4590) & (x172x) & (!x365x) & (n_n2401)) + ((n_n4593) & (!n_n4590) & (x172x) & (x365x) & (!n_n2401)) + ((n_n4593) & (!n_n4590) & (x172x) & (x365x) & (n_n2401)) + ((n_n4593) & (n_n4590) & (!x172x) & (!x365x) & (!n_n2401)) + ((n_n4593) & (n_n4590) & (!x172x) & (!x365x) & (n_n2401)) + ((n_n4593) & (n_n4590) & (!x172x) & (x365x) & (!n_n2401)) + ((n_n4593) & (n_n4590) & (!x172x) & (x365x) & (n_n2401)) + ((n_n4593) & (n_n4590) & (x172x) & (!x365x) & (!n_n2401)) + ((n_n4593) & (n_n4590) & (x172x) & (!x365x) & (n_n2401)) + ((n_n4593) & (n_n4590) & (x172x) & (x365x) & (!n_n2401)) + ((n_n4593) & (n_n4590) & (x172x) & (x365x) & (n_n2401)));
	assign x16611x = (((!n_n4616) & (!n_n4607) & (!n_n4618) & (n_n4611)) + ((!n_n4616) & (!n_n4607) & (n_n4618) & (!n_n4611)) + ((!n_n4616) & (!n_n4607) & (n_n4618) & (n_n4611)) + ((!n_n4616) & (n_n4607) & (!n_n4618) & (!n_n4611)) + ((!n_n4616) & (n_n4607) & (!n_n4618) & (n_n4611)) + ((!n_n4616) & (n_n4607) & (n_n4618) & (!n_n4611)) + ((!n_n4616) & (n_n4607) & (n_n4618) & (n_n4611)) + ((n_n4616) & (!n_n4607) & (!n_n4618) & (!n_n4611)) + ((n_n4616) & (!n_n4607) & (!n_n4618) & (n_n4611)) + ((n_n4616) & (!n_n4607) & (n_n4618) & (!n_n4611)) + ((n_n4616) & (!n_n4607) & (n_n4618) & (n_n4611)) + ((n_n4616) & (n_n4607) & (!n_n4618) & (!n_n4611)) + ((n_n4616) & (n_n4607) & (!n_n4618) & (n_n4611)) + ((n_n4616) & (n_n4607) & (n_n4618) & (!n_n4611)) + ((n_n4616) & (n_n4607) & (n_n4618) & (n_n4611)));
	assign x16612x = (((!n_n4613) & (!n_n4609) & (!n_n4608) & (!n_n4610) & (n_n4614)) + ((!n_n4613) & (!n_n4609) & (!n_n4608) & (n_n4610) & (!n_n4614)) + ((!n_n4613) & (!n_n4609) & (!n_n4608) & (n_n4610) & (n_n4614)) + ((!n_n4613) & (!n_n4609) & (n_n4608) & (!n_n4610) & (!n_n4614)) + ((!n_n4613) & (!n_n4609) & (n_n4608) & (!n_n4610) & (n_n4614)) + ((!n_n4613) & (!n_n4609) & (n_n4608) & (n_n4610) & (!n_n4614)) + ((!n_n4613) & (!n_n4609) & (n_n4608) & (n_n4610) & (n_n4614)) + ((!n_n4613) & (n_n4609) & (!n_n4608) & (!n_n4610) & (!n_n4614)) + ((!n_n4613) & (n_n4609) & (!n_n4608) & (!n_n4610) & (n_n4614)) + ((!n_n4613) & (n_n4609) & (!n_n4608) & (n_n4610) & (!n_n4614)) + ((!n_n4613) & (n_n4609) & (!n_n4608) & (n_n4610) & (n_n4614)) + ((!n_n4613) & (n_n4609) & (n_n4608) & (!n_n4610) & (!n_n4614)) + ((!n_n4613) & (n_n4609) & (n_n4608) & (!n_n4610) & (n_n4614)) + ((!n_n4613) & (n_n4609) & (n_n4608) & (n_n4610) & (!n_n4614)) + ((!n_n4613) & (n_n4609) & (n_n4608) & (n_n4610) & (n_n4614)) + ((n_n4613) & (!n_n4609) & (!n_n4608) & (!n_n4610) & (!n_n4614)) + ((n_n4613) & (!n_n4609) & (!n_n4608) & (!n_n4610) & (n_n4614)) + ((n_n4613) & (!n_n4609) & (!n_n4608) & (n_n4610) & (!n_n4614)) + ((n_n4613) & (!n_n4609) & (!n_n4608) & (n_n4610) & (n_n4614)) + ((n_n4613) & (!n_n4609) & (n_n4608) & (!n_n4610) & (!n_n4614)) + ((n_n4613) & (!n_n4609) & (n_n4608) & (!n_n4610) & (n_n4614)) + ((n_n4613) & (!n_n4609) & (n_n4608) & (n_n4610) & (!n_n4614)) + ((n_n4613) & (!n_n4609) & (n_n4608) & (n_n4610) & (n_n4614)) + ((n_n4613) & (n_n4609) & (!n_n4608) & (!n_n4610) & (!n_n4614)) + ((n_n4613) & (n_n4609) & (!n_n4608) & (!n_n4610) & (n_n4614)) + ((n_n4613) & (n_n4609) & (!n_n4608) & (n_n4610) & (!n_n4614)) + ((n_n4613) & (n_n4609) & (!n_n4608) & (n_n4610) & (n_n4614)) + ((n_n4613) & (n_n4609) & (n_n4608) & (!n_n4610) & (!n_n4614)) + ((n_n4613) & (n_n4609) & (n_n4608) & (!n_n4610) & (n_n4614)) + ((n_n4613) & (n_n4609) & (n_n4608) & (n_n4610) & (!n_n4614)) + ((n_n4613) & (n_n4609) & (n_n4608) & (n_n4610) & (n_n4614)));
	assign x16617x = (((!n_n4598) & (!n_n4601) & (!n_n4606) & (n_n4594)) + ((!n_n4598) & (!n_n4601) & (n_n4606) & (!n_n4594)) + ((!n_n4598) & (!n_n4601) & (n_n4606) & (n_n4594)) + ((!n_n4598) & (n_n4601) & (!n_n4606) & (!n_n4594)) + ((!n_n4598) & (n_n4601) & (!n_n4606) & (n_n4594)) + ((!n_n4598) & (n_n4601) & (n_n4606) & (!n_n4594)) + ((!n_n4598) & (n_n4601) & (n_n4606) & (n_n4594)) + ((n_n4598) & (!n_n4601) & (!n_n4606) & (!n_n4594)) + ((n_n4598) & (!n_n4601) & (!n_n4606) & (n_n4594)) + ((n_n4598) & (!n_n4601) & (n_n4606) & (!n_n4594)) + ((n_n4598) & (!n_n4601) & (n_n4606) & (n_n4594)) + ((n_n4598) & (n_n4601) & (!n_n4606) & (!n_n4594)) + ((n_n4598) & (n_n4601) & (!n_n4606) & (n_n4594)) + ((n_n4598) & (n_n4601) & (n_n4606) & (!n_n4594)) + ((n_n4598) & (n_n4601) & (n_n4606) & (n_n4594)));
	assign x16618x = (((!n_n4597) & (!n_n4605) & (!n_n4596) & (!n_n4600) & (n_n4603)) + ((!n_n4597) & (!n_n4605) & (!n_n4596) & (n_n4600) & (!n_n4603)) + ((!n_n4597) & (!n_n4605) & (!n_n4596) & (n_n4600) & (n_n4603)) + ((!n_n4597) & (!n_n4605) & (n_n4596) & (!n_n4600) & (!n_n4603)) + ((!n_n4597) & (!n_n4605) & (n_n4596) & (!n_n4600) & (n_n4603)) + ((!n_n4597) & (!n_n4605) & (n_n4596) & (n_n4600) & (!n_n4603)) + ((!n_n4597) & (!n_n4605) & (n_n4596) & (n_n4600) & (n_n4603)) + ((!n_n4597) & (n_n4605) & (!n_n4596) & (!n_n4600) & (!n_n4603)) + ((!n_n4597) & (n_n4605) & (!n_n4596) & (!n_n4600) & (n_n4603)) + ((!n_n4597) & (n_n4605) & (!n_n4596) & (n_n4600) & (!n_n4603)) + ((!n_n4597) & (n_n4605) & (!n_n4596) & (n_n4600) & (n_n4603)) + ((!n_n4597) & (n_n4605) & (n_n4596) & (!n_n4600) & (!n_n4603)) + ((!n_n4597) & (n_n4605) & (n_n4596) & (!n_n4600) & (n_n4603)) + ((!n_n4597) & (n_n4605) & (n_n4596) & (n_n4600) & (!n_n4603)) + ((!n_n4597) & (n_n4605) & (n_n4596) & (n_n4600) & (n_n4603)) + ((n_n4597) & (!n_n4605) & (!n_n4596) & (!n_n4600) & (!n_n4603)) + ((n_n4597) & (!n_n4605) & (!n_n4596) & (!n_n4600) & (n_n4603)) + ((n_n4597) & (!n_n4605) & (!n_n4596) & (n_n4600) & (!n_n4603)) + ((n_n4597) & (!n_n4605) & (!n_n4596) & (n_n4600) & (n_n4603)) + ((n_n4597) & (!n_n4605) & (n_n4596) & (!n_n4600) & (!n_n4603)) + ((n_n4597) & (!n_n4605) & (n_n4596) & (!n_n4600) & (n_n4603)) + ((n_n4597) & (!n_n4605) & (n_n4596) & (n_n4600) & (!n_n4603)) + ((n_n4597) & (!n_n4605) & (n_n4596) & (n_n4600) & (n_n4603)) + ((n_n4597) & (n_n4605) & (!n_n4596) & (!n_n4600) & (!n_n4603)) + ((n_n4597) & (n_n4605) & (!n_n4596) & (!n_n4600) & (n_n4603)) + ((n_n4597) & (n_n4605) & (!n_n4596) & (n_n4600) & (!n_n4603)) + ((n_n4597) & (n_n4605) & (!n_n4596) & (n_n4600) & (n_n4603)) + ((n_n4597) & (n_n4605) & (n_n4596) & (!n_n4600) & (!n_n4603)) + ((n_n4597) & (n_n4605) & (n_n4596) & (!n_n4600) & (n_n4603)) + ((n_n4597) & (n_n4605) & (n_n4596) & (n_n4600) & (!n_n4603)) + ((n_n4597) & (n_n4605) & (n_n4596) & (n_n4600) & (n_n4603)));
	assign n_n2246 = (((!n_n4629) & (!n_n4630) & (!x16632x) & (x190x)) + ((!n_n4629) & (!n_n4630) & (x16632x) & (!x190x)) + ((!n_n4629) & (!n_n4630) & (x16632x) & (x190x)) + ((!n_n4629) & (n_n4630) & (!x16632x) & (!x190x)) + ((!n_n4629) & (n_n4630) & (!x16632x) & (x190x)) + ((!n_n4629) & (n_n4630) & (x16632x) & (!x190x)) + ((!n_n4629) & (n_n4630) & (x16632x) & (x190x)) + ((n_n4629) & (!n_n4630) & (!x16632x) & (!x190x)) + ((n_n4629) & (!n_n4630) & (!x16632x) & (x190x)) + ((n_n4629) & (!n_n4630) & (x16632x) & (!x190x)) + ((n_n4629) & (!n_n4630) & (x16632x) & (x190x)) + ((n_n4629) & (n_n4630) & (!x16632x) & (!x190x)) + ((n_n4629) & (n_n4630) & (!x16632x) & (x190x)) + ((n_n4629) & (n_n4630) & (x16632x) & (!x190x)) + ((n_n4629) & (n_n4630) & (x16632x) & (x190x)));
	assign x16636x = (((!n_n4641) & (!n_n4639) & (!n_n4642) & (!n_n4633) & (n_n4635)) + ((!n_n4641) & (!n_n4639) & (!n_n4642) & (n_n4633) & (!n_n4635)) + ((!n_n4641) & (!n_n4639) & (!n_n4642) & (n_n4633) & (n_n4635)) + ((!n_n4641) & (!n_n4639) & (n_n4642) & (!n_n4633) & (!n_n4635)) + ((!n_n4641) & (!n_n4639) & (n_n4642) & (!n_n4633) & (n_n4635)) + ((!n_n4641) & (!n_n4639) & (n_n4642) & (n_n4633) & (!n_n4635)) + ((!n_n4641) & (!n_n4639) & (n_n4642) & (n_n4633) & (n_n4635)) + ((!n_n4641) & (n_n4639) & (!n_n4642) & (!n_n4633) & (!n_n4635)) + ((!n_n4641) & (n_n4639) & (!n_n4642) & (!n_n4633) & (n_n4635)) + ((!n_n4641) & (n_n4639) & (!n_n4642) & (n_n4633) & (!n_n4635)) + ((!n_n4641) & (n_n4639) & (!n_n4642) & (n_n4633) & (n_n4635)) + ((!n_n4641) & (n_n4639) & (n_n4642) & (!n_n4633) & (!n_n4635)) + ((!n_n4641) & (n_n4639) & (n_n4642) & (!n_n4633) & (n_n4635)) + ((!n_n4641) & (n_n4639) & (n_n4642) & (n_n4633) & (!n_n4635)) + ((!n_n4641) & (n_n4639) & (n_n4642) & (n_n4633) & (n_n4635)) + ((n_n4641) & (!n_n4639) & (!n_n4642) & (!n_n4633) & (!n_n4635)) + ((n_n4641) & (!n_n4639) & (!n_n4642) & (!n_n4633) & (n_n4635)) + ((n_n4641) & (!n_n4639) & (!n_n4642) & (n_n4633) & (!n_n4635)) + ((n_n4641) & (!n_n4639) & (!n_n4642) & (n_n4633) & (n_n4635)) + ((n_n4641) & (!n_n4639) & (n_n4642) & (!n_n4633) & (!n_n4635)) + ((n_n4641) & (!n_n4639) & (n_n4642) & (!n_n4633) & (n_n4635)) + ((n_n4641) & (!n_n4639) & (n_n4642) & (n_n4633) & (!n_n4635)) + ((n_n4641) & (!n_n4639) & (n_n4642) & (n_n4633) & (n_n4635)) + ((n_n4641) & (n_n4639) & (!n_n4642) & (!n_n4633) & (!n_n4635)) + ((n_n4641) & (n_n4639) & (!n_n4642) & (!n_n4633) & (n_n4635)) + ((n_n4641) & (n_n4639) & (!n_n4642) & (n_n4633) & (!n_n4635)) + ((n_n4641) & (n_n4639) & (!n_n4642) & (n_n4633) & (n_n4635)) + ((n_n4641) & (n_n4639) & (n_n4642) & (!n_n4633) & (!n_n4635)) + ((n_n4641) & (n_n4639) & (n_n4642) & (!n_n4633) & (n_n4635)) + ((n_n4641) & (n_n4639) & (n_n4642) & (n_n4633) & (!n_n4635)) + ((n_n4641) & (n_n4639) & (n_n4642) & (n_n4633) & (n_n4635)));
	assign x22061x = (((!n_n4648) & (!n_n4646) & (!x311x) & (!x119x) & (!x271x)));
	assign n_n4549 = (((i_1_) & (!i_2_) & (i_0_) & (n_n473) & (x20x)));
	assign n_n4548 = (((i_9_) & (n_n455) & (n_n473) & (n_n522)));
	assign n_n4559 = (((!i_9_) & (n_n455) & (n_n528) & (n_n464)));
	assign n_n4552 = (((i_9_) & (n_n455) & (n_n534) & (n_n464)));
	assign n_n5106 = (((i_7_) & (!i_8_) & (!i_6_) & (n_n518) & (x12x)));
	assign n_n5117 = (((!i_9_) & (n_n509) & (n_n130) & (n_n530)));
	assign n_n5121 = (((!i_9_) & (n_n526) & (n_n509) & (n_n130)));
	assign n_n5122 = (((i_7_) & (!i_8_) & (!i_6_) & (n_n509) & (x12x)));
	assign x35x = (((!n_n524) & (!n_n509) & (!x12x) & (n_n5121)) + ((!n_n524) & (!n_n509) & (x12x) & (n_n5121)) + ((!n_n524) & (n_n509) & (!x12x) & (n_n5121)) + ((!n_n524) & (n_n509) & (x12x) & (n_n5121)) + ((n_n524) & (!n_n509) & (!x12x) & (n_n5121)) + ((n_n524) & (!n_n509) & (x12x) & (n_n5121)) + ((n_n524) & (n_n509) & (!x12x) & (n_n5121)) + ((n_n524) & (n_n509) & (x12x) & (!n_n5121)) + ((n_n524) & (n_n509) & (x12x) & (n_n5121)));
	assign n_n5223 = (((i_5_) & (i_3_) & (i_4_) & (x23x) & (n_n65)));
	assign n_n5328 = (((i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n464)));
	assign n_n5254 = (((i_5_) & (i_3_) & (!i_4_) & (x19x) & (n_n520)));
	assign n_n5249 = (((!i_9_) & (n_n526) & (n_n509) & (n_n65)));
	assign n_n5233 = (((!i_9_) & (n_n518) & (n_n526) & (n_n65)));
	assign n_n5236 = (((!i_5_) & (i_3_) & (i_4_) & (x19x) & (n_n522)));
	assign n_n5262 = (((!i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n500)));
	assign n_n5278 = (((!i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n491)));
	assign n_n5290 = (((!i_5_) & (!i_3_) & (i_4_) & (x19x) & (n_n532)));
	assign n_n5289 = (((!i_9_) & (n_n482) & (n_n534) & (n_n65)));
	assign x392x = (((!x25x) & (x19x) & (n_n482) & (n_n532) & (!n_n65)) + ((!x25x) & (x19x) & (n_n482) & (n_n532) & (n_n65)) + ((x25x) & (!x19x) & (n_n482) & (!n_n532) & (n_n65)) + ((x25x) & (!x19x) & (n_n482) & (n_n532) & (n_n65)) + ((x25x) & (x19x) & (n_n482) & (!n_n532) & (n_n65)) + ((x25x) & (x19x) & (n_n482) & (n_n532) & (!n_n65)) + ((x25x) & (x19x) & (n_n482) & (n_n532) & (n_n65)));
	assign n_n5217 = (((!i_9_) & (n_n526) & (n_n535) & (n_n65)));
	assign x449x = (((!i_9_) & (!x19x) & (n_n526) & (n_n535) & (n_n65)) + ((!i_9_) & (x19x) & (n_n526) & (n_n535) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n526) & (n_n535) & (n_n65)) + ((i_9_) & (x19x) & (n_n526) & (n_n535) & (!n_n65)) + ((i_9_) & (x19x) & (n_n526) & (n_n535) & (n_n65)));
	assign x16778x = (((!n_n5236) & (!n_n5262) & (!n_n5278) & (!n_n5290) & (n_n5289)) + ((!n_n5236) & (!n_n5262) & (!n_n5278) & (n_n5290) & (!n_n5289)) + ((!n_n5236) & (!n_n5262) & (!n_n5278) & (n_n5290) & (n_n5289)) + ((!n_n5236) & (!n_n5262) & (n_n5278) & (!n_n5290) & (!n_n5289)) + ((!n_n5236) & (!n_n5262) & (n_n5278) & (!n_n5290) & (n_n5289)) + ((!n_n5236) & (!n_n5262) & (n_n5278) & (n_n5290) & (!n_n5289)) + ((!n_n5236) & (!n_n5262) & (n_n5278) & (n_n5290) & (n_n5289)) + ((!n_n5236) & (n_n5262) & (!n_n5278) & (!n_n5290) & (!n_n5289)) + ((!n_n5236) & (n_n5262) & (!n_n5278) & (!n_n5290) & (n_n5289)) + ((!n_n5236) & (n_n5262) & (!n_n5278) & (n_n5290) & (!n_n5289)) + ((!n_n5236) & (n_n5262) & (!n_n5278) & (n_n5290) & (n_n5289)) + ((!n_n5236) & (n_n5262) & (n_n5278) & (!n_n5290) & (!n_n5289)) + ((!n_n5236) & (n_n5262) & (n_n5278) & (!n_n5290) & (n_n5289)) + ((!n_n5236) & (n_n5262) & (n_n5278) & (n_n5290) & (!n_n5289)) + ((!n_n5236) & (n_n5262) & (n_n5278) & (n_n5290) & (n_n5289)) + ((n_n5236) & (!n_n5262) & (!n_n5278) & (!n_n5290) & (!n_n5289)) + ((n_n5236) & (!n_n5262) & (!n_n5278) & (!n_n5290) & (n_n5289)) + ((n_n5236) & (!n_n5262) & (!n_n5278) & (n_n5290) & (!n_n5289)) + ((n_n5236) & (!n_n5262) & (!n_n5278) & (n_n5290) & (n_n5289)) + ((n_n5236) & (!n_n5262) & (n_n5278) & (!n_n5290) & (!n_n5289)) + ((n_n5236) & (!n_n5262) & (n_n5278) & (!n_n5290) & (n_n5289)) + ((n_n5236) & (!n_n5262) & (n_n5278) & (n_n5290) & (!n_n5289)) + ((n_n5236) & (!n_n5262) & (n_n5278) & (n_n5290) & (n_n5289)) + ((n_n5236) & (n_n5262) & (!n_n5278) & (!n_n5290) & (!n_n5289)) + ((n_n5236) & (n_n5262) & (!n_n5278) & (!n_n5290) & (n_n5289)) + ((n_n5236) & (n_n5262) & (!n_n5278) & (n_n5290) & (!n_n5289)) + ((n_n5236) & (n_n5262) & (!n_n5278) & (n_n5290) & (n_n5289)) + ((n_n5236) & (n_n5262) & (n_n5278) & (!n_n5290) & (!n_n5289)) + ((n_n5236) & (n_n5262) & (n_n5278) & (!n_n5290) & (n_n5289)) + ((n_n5236) & (n_n5262) & (n_n5278) & (n_n5290) & (!n_n5289)) + ((n_n5236) & (n_n5262) & (n_n5278) & (n_n5290) & (n_n5289)));
	assign x16777x = (((!n_n5328) & (!n_n5254) & (!n_n5249) & (n_n5233)) + ((!n_n5328) & (!n_n5254) & (n_n5249) & (!n_n5233)) + ((!n_n5328) & (!n_n5254) & (n_n5249) & (n_n5233)) + ((!n_n5328) & (n_n5254) & (!n_n5249) & (!n_n5233)) + ((!n_n5328) & (n_n5254) & (!n_n5249) & (n_n5233)) + ((!n_n5328) & (n_n5254) & (n_n5249) & (!n_n5233)) + ((!n_n5328) & (n_n5254) & (n_n5249) & (n_n5233)) + ((n_n5328) & (!n_n5254) & (!n_n5249) & (!n_n5233)) + ((n_n5328) & (!n_n5254) & (!n_n5249) & (n_n5233)) + ((n_n5328) & (!n_n5254) & (n_n5249) & (!n_n5233)) + ((n_n5328) & (!n_n5254) & (n_n5249) & (n_n5233)) + ((n_n5328) & (n_n5254) & (!n_n5249) & (!n_n5233)) + ((n_n5328) & (n_n5254) & (!n_n5249) & (n_n5233)) + ((n_n5328) & (n_n5254) & (n_n5249) & (!n_n5233)) + ((n_n5328) & (n_n5254) & (n_n5249) & (n_n5233)));
	assign x16779x = (((!n_n5206) & (!n_n5216) & (!n_n5223) & (!n_n5217) & (x16777x)) + ((!n_n5206) & (!n_n5216) & (!n_n5223) & (n_n5217) & (!x16777x)) + ((!n_n5206) & (!n_n5216) & (!n_n5223) & (n_n5217) & (x16777x)) + ((!n_n5206) & (!n_n5216) & (n_n5223) & (!n_n5217) & (!x16777x)) + ((!n_n5206) & (!n_n5216) & (n_n5223) & (!n_n5217) & (x16777x)) + ((!n_n5206) & (!n_n5216) & (n_n5223) & (n_n5217) & (!x16777x)) + ((!n_n5206) & (!n_n5216) & (n_n5223) & (n_n5217) & (x16777x)) + ((!n_n5206) & (n_n5216) & (!n_n5223) & (!n_n5217) & (!x16777x)) + ((!n_n5206) & (n_n5216) & (!n_n5223) & (!n_n5217) & (x16777x)) + ((!n_n5206) & (n_n5216) & (!n_n5223) & (n_n5217) & (!x16777x)) + ((!n_n5206) & (n_n5216) & (!n_n5223) & (n_n5217) & (x16777x)) + ((!n_n5206) & (n_n5216) & (n_n5223) & (!n_n5217) & (!x16777x)) + ((!n_n5206) & (n_n5216) & (n_n5223) & (!n_n5217) & (x16777x)) + ((!n_n5206) & (n_n5216) & (n_n5223) & (n_n5217) & (!x16777x)) + ((!n_n5206) & (n_n5216) & (n_n5223) & (n_n5217) & (x16777x)) + ((n_n5206) & (!n_n5216) & (!n_n5223) & (!n_n5217) & (!x16777x)) + ((n_n5206) & (!n_n5216) & (!n_n5223) & (!n_n5217) & (x16777x)) + ((n_n5206) & (!n_n5216) & (!n_n5223) & (n_n5217) & (!x16777x)) + ((n_n5206) & (!n_n5216) & (!n_n5223) & (n_n5217) & (x16777x)) + ((n_n5206) & (!n_n5216) & (n_n5223) & (!n_n5217) & (!x16777x)) + ((n_n5206) & (!n_n5216) & (n_n5223) & (!n_n5217) & (x16777x)) + ((n_n5206) & (!n_n5216) & (n_n5223) & (n_n5217) & (!x16777x)) + ((n_n5206) & (!n_n5216) & (n_n5223) & (n_n5217) & (x16777x)) + ((n_n5206) & (n_n5216) & (!n_n5223) & (!n_n5217) & (!x16777x)) + ((n_n5206) & (n_n5216) & (!n_n5223) & (!n_n5217) & (x16777x)) + ((n_n5206) & (n_n5216) & (!n_n5223) & (n_n5217) & (!x16777x)) + ((n_n5206) & (n_n5216) & (!n_n5223) & (n_n5217) & (x16777x)) + ((n_n5206) & (n_n5216) & (n_n5223) & (!n_n5217) & (!x16777x)) + ((n_n5206) & (n_n5216) & (n_n5223) & (!n_n5217) & (x16777x)) + ((n_n5206) & (n_n5216) & (n_n5223) & (n_n5217) & (!x16777x)) + ((n_n5206) & (n_n5216) & (n_n5223) & (n_n5217) & (x16777x)));
	assign n_n4833 = (((!i_9_) & (n_n526) & (n_n260) & (n_n535)));
	assign n_n4940 = (((i_9_) & (n_n260) & (n_n530) & (n_n464)));
	assign n_n4939 = (((!i_9_) & (n_n532) & (n_n260) & (n_n464)));
	assign x373x = (((!i_9_) & (n_n509) & (n_n325) & (!n_n520) & (x23x)) + ((!i_9_) & (n_n509) & (n_n325) & (n_n520) & (x23x)) + ((i_9_) & (n_n509) & (n_n325) & (!n_n520) & (x23x)) + ((i_9_) & (n_n509) & (n_n325) & (n_n520) & (!x23x)) + ((i_9_) & (n_n509) & (n_n325) & (n_n520) & (x23x)));
	assign x374x = (((!i_9_) & (n_n509) & (n_n325) & (!n_n522) & (x20x)) + ((!i_9_) & (n_n509) & (n_n325) & (n_n522) & (x20x)) + ((i_9_) & (n_n509) & (n_n325) & (!n_n522) & (x20x)) + ((i_9_) & (n_n509) & (n_n325) & (n_n522) & (!x20x)) + ((i_9_) & (n_n509) & (n_n325) & (n_n522) & (x20x)));
	assign x22073x = (((!x25x) & (!x483x) & (!n_n4734) & (!n_n4728) & (!x373x)) + ((!x25x) & (x483x) & (!n_n4734) & (!n_n4728) & (!x373x)) + ((x25x) & (!x483x) & (!n_n4734) & (!n_n4728) & (!x373x)));
	assign n_n5132 = (((!i_5_) & (i_3_) & (!i_4_) & (x12x) & (n_n530)));
	assign n_n5128 = (((i_7_) & (i_8_) & (i_6_) & (x12x) & (n_n500)));
	assign n_n5016 = (((i_9_) & (n_n534) & (n_n491) & (n_n195)));
	assign x12253x = (((!n_n5026) & (!n_n5017) & (!n_n5014) & (!n_n5015) & (n_n5016)) + ((!n_n5026) & (!n_n5017) & (!n_n5014) & (n_n5015) & (!n_n5016)) + ((!n_n5026) & (!n_n5017) & (!n_n5014) & (n_n5015) & (n_n5016)) + ((!n_n5026) & (!n_n5017) & (n_n5014) & (!n_n5015) & (!n_n5016)) + ((!n_n5026) & (!n_n5017) & (n_n5014) & (!n_n5015) & (n_n5016)) + ((!n_n5026) & (!n_n5017) & (n_n5014) & (n_n5015) & (!n_n5016)) + ((!n_n5026) & (!n_n5017) & (n_n5014) & (n_n5015) & (n_n5016)) + ((!n_n5026) & (n_n5017) & (!n_n5014) & (!n_n5015) & (!n_n5016)) + ((!n_n5026) & (n_n5017) & (!n_n5014) & (!n_n5015) & (n_n5016)) + ((!n_n5026) & (n_n5017) & (!n_n5014) & (n_n5015) & (!n_n5016)) + ((!n_n5026) & (n_n5017) & (!n_n5014) & (n_n5015) & (n_n5016)) + ((!n_n5026) & (n_n5017) & (n_n5014) & (!n_n5015) & (!n_n5016)) + ((!n_n5026) & (n_n5017) & (n_n5014) & (!n_n5015) & (n_n5016)) + ((!n_n5026) & (n_n5017) & (n_n5014) & (n_n5015) & (!n_n5016)) + ((!n_n5026) & (n_n5017) & (n_n5014) & (n_n5015) & (n_n5016)) + ((n_n5026) & (!n_n5017) & (!n_n5014) & (!n_n5015) & (!n_n5016)) + ((n_n5026) & (!n_n5017) & (!n_n5014) & (!n_n5015) & (n_n5016)) + ((n_n5026) & (!n_n5017) & (!n_n5014) & (n_n5015) & (!n_n5016)) + ((n_n5026) & (!n_n5017) & (!n_n5014) & (n_n5015) & (n_n5016)) + ((n_n5026) & (!n_n5017) & (n_n5014) & (!n_n5015) & (!n_n5016)) + ((n_n5026) & (!n_n5017) & (n_n5014) & (!n_n5015) & (n_n5016)) + ((n_n5026) & (!n_n5017) & (n_n5014) & (n_n5015) & (!n_n5016)) + ((n_n5026) & (!n_n5017) & (n_n5014) & (n_n5015) & (n_n5016)) + ((n_n5026) & (n_n5017) & (!n_n5014) & (!n_n5015) & (!n_n5016)) + ((n_n5026) & (n_n5017) & (!n_n5014) & (!n_n5015) & (n_n5016)) + ((n_n5026) & (n_n5017) & (!n_n5014) & (n_n5015) & (!n_n5016)) + ((n_n5026) & (n_n5017) & (!n_n5014) & (n_n5015) & (n_n5016)) + ((n_n5026) & (n_n5017) & (n_n5014) & (!n_n5015) & (!n_n5016)) + ((n_n5026) & (n_n5017) & (n_n5014) & (!n_n5015) & (n_n5016)) + ((n_n5026) & (n_n5017) & (n_n5014) & (n_n5015) & (!n_n5016)) + ((n_n5026) & (n_n5017) & (n_n5014) & (n_n5015) & (n_n5016)));
	assign n_n1453 = (((!n_n5023) & (!n_n5021) & (!n_n5019) & (!n_n5020) & (x12253x)) + ((!n_n5023) & (!n_n5021) & (!n_n5019) & (n_n5020) & (!x12253x)) + ((!n_n5023) & (!n_n5021) & (!n_n5019) & (n_n5020) & (x12253x)) + ((!n_n5023) & (!n_n5021) & (n_n5019) & (!n_n5020) & (!x12253x)) + ((!n_n5023) & (!n_n5021) & (n_n5019) & (!n_n5020) & (x12253x)) + ((!n_n5023) & (!n_n5021) & (n_n5019) & (n_n5020) & (!x12253x)) + ((!n_n5023) & (!n_n5021) & (n_n5019) & (n_n5020) & (x12253x)) + ((!n_n5023) & (n_n5021) & (!n_n5019) & (!n_n5020) & (!x12253x)) + ((!n_n5023) & (n_n5021) & (!n_n5019) & (!n_n5020) & (x12253x)) + ((!n_n5023) & (n_n5021) & (!n_n5019) & (n_n5020) & (!x12253x)) + ((!n_n5023) & (n_n5021) & (!n_n5019) & (n_n5020) & (x12253x)) + ((!n_n5023) & (n_n5021) & (n_n5019) & (!n_n5020) & (!x12253x)) + ((!n_n5023) & (n_n5021) & (n_n5019) & (!n_n5020) & (x12253x)) + ((!n_n5023) & (n_n5021) & (n_n5019) & (n_n5020) & (!x12253x)) + ((!n_n5023) & (n_n5021) & (n_n5019) & (n_n5020) & (x12253x)) + ((n_n5023) & (!n_n5021) & (!n_n5019) & (!n_n5020) & (!x12253x)) + ((n_n5023) & (!n_n5021) & (!n_n5019) & (!n_n5020) & (x12253x)) + ((n_n5023) & (!n_n5021) & (!n_n5019) & (n_n5020) & (!x12253x)) + ((n_n5023) & (!n_n5021) & (!n_n5019) & (n_n5020) & (x12253x)) + ((n_n5023) & (!n_n5021) & (n_n5019) & (!n_n5020) & (!x12253x)) + ((n_n5023) & (!n_n5021) & (n_n5019) & (!n_n5020) & (x12253x)) + ((n_n5023) & (!n_n5021) & (n_n5019) & (n_n5020) & (!x12253x)) + ((n_n5023) & (!n_n5021) & (n_n5019) & (n_n5020) & (x12253x)) + ((n_n5023) & (n_n5021) & (!n_n5019) & (!n_n5020) & (!x12253x)) + ((n_n5023) & (n_n5021) & (!n_n5019) & (!n_n5020) & (x12253x)) + ((n_n5023) & (n_n5021) & (!n_n5019) & (n_n5020) & (!x12253x)) + ((n_n5023) & (n_n5021) & (!n_n5019) & (n_n5020) & (x12253x)) + ((n_n5023) & (n_n5021) & (n_n5019) & (!n_n5020) & (!x12253x)) + ((n_n5023) & (n_n5021) & (n_n5019) & (!n_n5020) & (x12253x)) + ((n_n5023) & (n_n5021) & (n_n5019) & (n_n5020) & (!x12253x)) + ((n_n5023) & (n_n5021) & (n_n5019) & (n_n5020) & (x12253x)));
	assign n_n4129 = (((!i_9_) & (!n_n473) & (!n_n130) & (!n_n530) & (n_n5182)) + ((!i_9_) & (!n_n473) & (!n_n130) & (n_n530) & (n_n5182)) + ((!i_9_) & (!n_n473) & (n_n130) & (!n_n530) & (n_n5182)) + ((!i_9_) & (!n_n473) & (n_n130) & (n_n530) & (n_n5182)) + ((!i_9_) & (n_n473) & (!n_n130) & (!n_n530) & (n_n5182)) + ((!i_9_) & (n_n473) & (!n_n130) & (n_n530) & (n_n5182)) + ((!i_9_) & (n_n473) & (n_n130) & (!n_n530) & (n_n5182)) + ((!i_9_) & (n_n473) & (n_n130) & (n_n530) & (!n_n5182)) + ((!i_9_) & (n_n473) & (n_n130) & (n_n530) & (n_n5182)) + ((i_9_) & (!n_n473) & (!n_n130) & (!n_n530) & (n_n5182)) + ((i_9_) & (!n_n473) & (!n_n130) & (n_n530) & (n_n5182)) + ((i_9_) & (!n_n473) & (n_n130) & (!n_n530) & (n_n5182)) + ((i_9_) & (!n_n473) & (n_n130) & (n_n530) & (n_n5182)) + ((i_9_) & (n_n473) & (!n_n130) & (!n_n530) & (n_n5182)) + ((i_9_) & (n_n473) & (!n_n130) & (n_n530) & (n_n5182)) + ((i_9_) & (n_n473) & (n_n130) & (!n_n530) & (n_n5182)) + ((i_9_) & (n_n473) & (n_n130) & (n_n530) & (!n_n5182)) + ((i_9_) & (n_n473) & (n_n130) & (n_n530) & (n_n5182)));
	assign n_n3019 = (((!x19x) & (!n_n473) & (!n_n532) & (!n_n530) & (n_n5307)) + ((!x19x) & (!n_n473) & (!n_n532) & (n_n530) & (n_n5307)) + ((!x19x) & (!n_n473) & (n_n532) & (!n_n530) & (n_n5307)) + ((!x19x) & (!n_n473) & (n_n532) & (n_n530) & (n_n5307)) + ((!x19x) & (n_n473) & (!n_n532) & (!n_n530) & (n_n5307)) + ((!x19x) & (n_n473) & (!n_n532) & (n_n530) & (n_n5307)) + ((!x19x) & (n_n473) & (n_n532) & (!n_n530) & (n_n5307)) + ((!x19x) & (n_n473) & (n_n532) & (n_n530) & (n_n5307)) + ((x19x) & (!n_n473) & (!n_n532) & (!n_n530) & (n_n5307)) + ((x19x) & (!n_n473) & (!n_n532) & (n_n530) & (n_n5307)) + ((x19x) & (!n_n473) & (n_n532) & (!n_n530) & (n_n5307)) + ((x19x) & (!n_n473) & (n_n532) & (n_n530) & (n_n5307)) + ((x19x) & (n_n473) & (!n_n532) & (!n_n530) & (n_n5307)) + ((x19x) & (n_n473) & (!n_n532) & (n_n530) & (!n_n5307)) + ((x19x) & (n_n473) & (!n_n532) & (n_n530) & (n_n5307)) + ((x19x) & (n_n473) & (n_n532) & (!n_n530) & (!n_n5307)) + ((x19x) & (n_n473) & (n_n532) & (!n_n530) & (n_n5307)) + ((x19x) & (n_n473) & (n_n532) & (n_n530) & (!n_n5307)) + ((x19x) & (n_n473) & (n_n532) & (n_n530) & (n_n5307)));
	assign n_n5009 = (((!i_9_) & (n_n526) & (n_n195) & (n_n500)));
	assign n_n4562 = (((i_9_) & (n_n524) & (n_n455) & (n_n464)));
	assign x12048x = (((!n_n4617) & (!n_n4618) & (!n_n4576) & (n_n4569)) + ((!n_n4617) & (!n_n4618) & (n_n4576) & (!n_n4569)) + ((!n_n4617) & (!n_n4618) & (n_n4576) & (n_n4569)) + ((!n_n4617) & (n_n4618) & (!n_n4576) & (!n_n4569)) + ((!n_n4617) & (n_n4618) & (!n_n4576) & (n_n4569)) + ((!n_n4617) & (n_n4618) & (n_n4576) & (!n_n4569)) + ((!n_n4617) & (n_n4618) & (n_n4576) & (n_n4569)) + ((n_n4617) & (!n_n4618) & (!n_n4576) & (!n_n4569)) + ((n_n4617) & (!n_n4618) & (!n_n4576) & (n_n4569)) + ((n_n4617) & (!n_n4618) & (n_n4576) & (!n_n4569)) + ((n_n4617) & (!n_n4618) & (n_n4576) & (n_n4569)) + ((n_n4617) & (n_n4618) & (!n_n4576) & (!n_n4569)) + ((n_n4617) & (n_n4618) & (!n_n4576) & (n_n4569)) + ((n_n4617) & (n_n4618) & (n_n4576) & (!n_n4569)) + ((n_n4617) & (n_n4618) & (n_n4576) & (n_n4569)));
	assign n_n4635 = (((!i_9_) & (n_n390) & (n_n532) & (n_n491)));
	assign x12049x = (((!x10x) & (!x572x) & (!x172x) & (!n_n4580) & (n_n4635)) + ((!x10x) & (!x572x) & (!x172x) & (n_n4580) & (!n_n4635)) + ((!x10x) & (!x572x) & (!x172x) & (n_n4580) & (n_n4635)) + ((!x10x) & (!x572x) & (x172x) & (!n_n4580) & (!n_n4635)) + ((!x10x) & (!x572x) & (x172x) & (!n_n4580) & (n_n4635)) + ((!x10x) & (!x572x) & (x172x) & (n_n4580) & (!n_n4635)) + ((!x10x) & (!x572x) & (x172x) & (n_n4580) & (n_n4635)) + ((!x10x) & (x572x) & (!x172x) & (!n_n4580) & (n_n4635)) + ((!x10x) & (x572x) & (!x172x) & (n_n4580) & (!n_n4635)) + ((!x10x) & (x572x) & (!x172x) & (n_n4580) & (n_n4635)) + ((!x10x) & (x572x) & (x172x) & (!n_n4580) & (!n_n4635)) + ((!x10x) & (x572x) & (x172x) & (!n_n4580) & (n_n4635)) + ((!x10x) & (x572x) & (x172x) & (n_n4580) & (!n_n4635)) + ((!x10x) & (x572x) & (x172x) & (n_n4580) & (n_n4635)) + ((x10x) & (!x572x) & (!x172x) & (!n_n4580) & (n_n4635)) + ((x10x) & (!x572x) & (!x172x) & (n_n4580) & (!n_n4635)) + ((x10x) & (!x572x) & (!x172x) & (n_n4580) & (n_n4635)) + ((x10x) & (!x572x) & (x172x) & (!n_n4580) & (!n_n4635)) + ((x10x) & (!x572x) & (x172x) & (!n_n4580) & (n_n4635)) + ((x10x) & (!x572x) & (x172x) & (n_n4580) & (!n_n4635)) + ((x10x) & (!x572x) & (x172x) & (n_n4580) & (n_n4635)) + ((x10x) & (x572x) & (!x172x) & (!n_n4580) & (!n_n4635)) + ((x10x) & (x572x) & (!x172x) & (!n_n4580) & (n_n4635)) + ((x10x) & (x572x) & (!x172x) & (n_n4580) & (!n_n4635)) + ((x10x) & (x572x) & (!x172x) & (n_n4580) & (n_n4635)) + ((x10x) & (x572x) & (x172x) & (!n_n4580) & (!n_n4635)) + ((x10x) & (x572x) & (x172x) & (!n_n4580) & (n_n4635)) + ((x10x) & (x572x) & (x172x) & (n_n4580) & (!n_n4635)) + ((x10x) & (x572x) & (x172x) & (n_n4580) & (n_n4635)));
	assign x12053x = (((!n_n455) & (!x24x) & (!n_n4438) & (!n_n500) & (x184x)) + ((!n_n455) & (!x24x) & (!n_n4438) & (n_n500) & (x184x)) + ((!n_n455) & (!x24x) & (n_n4438) & (!n_n500) & (!x184x)) + ((!n_n455) & (!x24x) & (n_n4438) & (!n_n500) & (x184x)) + ((!n_n455) & (!x24x) & (n_n4438) & (n_n500) & (!x184x)) + ((!n_n455) & (!x24x) & (n_n4438) & (n_n500) & (x184x)) + ((!n_n455) & (x24x) & (!n_n4438) & (!n_n500) & (x184x)) + ((!n_n455) & (x24x) & (!n_n4438) & (n_n500) & (x184x)) + ((!n_n455) & (x24x) & (n_n4438) & (!n_n500) & (!x184x)) + ((!n_n455) & (x24x) & (n_n4438) & (!n_n500) & (x184x)) + ((!n_n455) & (x24x) & (n_n4438) & (n_n500) & (!x184x)) + ((!n_n455) & (x24x) & (n_n4438) & (n_n500) & (x184x)) + ((n_n455) & (!x24x) & (!n_n4438) & (!n_n500) & (x184x)) + ((n_n455) & (!x24x) & (!n_n4438) & (n_n500) & (x184x)) + ((n_n455) & (!x24x) & (n_n4438) & (!n_n500) & (!x184x)) + ((n_n455) & (!x24x) & (n_n4438) & (!n_n500) & (x184x)) + ((n_n455) & (!x24x) & (n_n4438) & (n_n500) & (!x184x)) + ((n_n455) & (!x24x) & (n_n4438) & (n_n500) & (x184x)) + ((n_n455) & (x24x) & (!n_n4438) & (!n_n500) & (x184x)) + ((n_n455) & (x24x) & (!n_n4438) & (n_n500) & (!x184x)) + ((n_n455) & (x24x) & (!n_n4438) & (n_n500) & (x184x)) + ((n_n455) & (x24x) & (n_n4438) & (!n_n500) & (!x184x)) + ((n_n455) & (x24x) & (n_n4438) & (!n_n500) & (x184x)) + ((n_n455) & (x24x) & (n_n4438) & (n_n500) & (!x184x)) + ((n_n455) & (x24x) & (n_n4438) & (n_n500) & (x184x)));
	assign x12054x = (((!n_n4436) & (!x70x) & (!n_n4458) & (n_n4474)) + ((!n_n4436) & (!x70x) & (n_n4458) & (!n_n4474)) + ((!n_n4436) & (!x70x) & (n_n4458) & (n_n4474)) + ((!n_n4436) & (x70x) & (!n_n4458) & (!n_n4474)) + ((!n_n4436) & (x70x) & (!n_n4458) & (n_n4474)) + ((!n_n4436) & (x70x) & (n_n4458) & (!n_n4474)) + ((!n_n4436) & (x70x) & (n_n4458) & (n_n4474)) + ((n_n4436) & (!x70x) & (!n_n4458) & (!n_n4474)) + ((n_n4436) & (!x70x) & (!n_n4458) & (n_n4474)) + ((n_n4436) & (!x70x) & (n_n4458) & (!n_n4474)) + ((n_n4436) & (!x70x) & (n_n4458) & (n_n4474)) + ((n_n4436) & (x70x) & (!n_n4458) & (!n_n4474)) + ((n_n4436) & (x70x) & (!n_n4458) & (n_n4474)) + ((n_n4436) & (x70x) & (n_n4458) & (!n_n4474)) + ((n_n4436) & (x70x) & (n_n4458) & (n_n4474)));
	assign x12061x = (((!n_n4512) & (!n_n4526) & (!n_n4535) & (!n_n4492) & (n_n4496)) + ((!n_n4512) & (!n_n4526) & (!n_n4535) & (n_n4492) & (!n_n4496)) + ((!n_n4512) & (!n_n4526) & (!n_n4535) & (n_n4492) & (n_n4496)) + ((!n_n4512) & (!n_n4526) & (n_n4535) & (!n_n4492) & (!n_n4496)) + ((!n_n4512) & (!n_n4526) & (n_n4535) & (!n_n4492) & (n_n4496)) + ((!n_n4512) & (!n_n4526) & (n_n4535) & (n_n4492) & (!n_n4496)) + ((!n_n4512) & (!n_n4526) & (n_n4535) & (n_n4492) & (n_n4496)) + ((!n_n4512) & (n_n4526) & (!n_n4535) & (!n_n4492) & (!n_n4496)) + ((!n_n4512) & (n_n4526) & (!n_n4535) & (!n_n4492) & (n_n4496)) + ((!n_n4512) & (n_n4526) & (!n_n4535) & (n_n4492) & (!n_n4496)) + ((!n_n4512) & (n_n4526) & (!n_n4535) & (n_n4492) & (n_n4496)) + ((!n_n4512) & (n_n4526) & (n_n4535) & (!n_n4492) & (!n_n4496)) + ((!n_n4512) & (n_n4526) & (n_n4535) & (!n_n4492) & (n_n4496)) + ((!n_n4512) & (n_n4526) & (n_n4535) & (n_n4492) & (!n_n4496)) + ((!n_n4512) & (n_n4526) & (n_n4535) & (n_n4492) & (n_n4496)) + ((n_n4512) & (!n_n4526) & (!n_n4535) & (!n_n4492) & (!n_n4496)) + ((n_n4512) & (!n_n4526) & (!n_n4535) & (!n_n4492) & (n_n4496)) + ((n_n4512) & (!n_n4526) & (!n_n4535) & (n_n4492) & (!n_n4496)) + ((n_n4512) & (!n_n4526) & (!n_n4535) & (n_n4492) & (n_n4496)) + ((n_n4512) & (!n_n4526) & (n_n4535) & (!n_n4492) & (!n_n4496)) + ((n_n4512) & (!n_n4526) & (n_n4535) & (!n_n4492) & (n_n4496)) + ((n_n4512) & (!n_n4526) & (n_n4535) & (n_n4492) & (!n_n4496)) + ((n_n4512) & (!n_n4526) & (n_n4535) & (n_n4492) & (n_n4496)) + ((n_n4512) & (n_n4526) & (!n_n4535) & (!n_n4492) & (!n_n4496)) + ((n_n4512) & (n_n4526) & (!n_n4535) & (!n_n4492) & (n_n4496)) + ((n_n4512) & (n_n4526) & (!n_n4535) & (n_n4492) & (!n_n4496)) + ((n_n4512) & (n_n4526) & (!n_n4535) & (n_n4492) & (n_n4496)) + ((n_n4512) & (n_n4526) & (n_n4535) & (!n_n4492) & (!n_n4496)) + ((n_n4512) & (n_n4526) & (n_n4535) & (!n_n4492) & (n_n4496)) + ((n_n4512) & (n_n4526) & (n_n4535) & (n_n4492) & (!n_n4496)) + ((n_n4512) & (n_n4526) & (n_n4535) & (n_n4492) & (n_n4496)));
	assign x12068x = (((!n_n4737) & (!n_n4756) & (!n_n4724) & (n_n4759)) + ((!n_n4737) & (!n_n4756) & (n_n4724) & (!n_n4759)) + ((!n_n4737) & (!n_n4756) & (n_n4724) & (n_n4759)) + ((!n_n4737) & (n_n4756) & (!n_n4724) & (!n_n4759)) + ((!n_n4737) & (n_n4756) & (!n_n4724) & (n_n4759)) + ((!n_n4737) & (n_n4756) & (n_n4724) & (!n_n4759)) + ((!n_n4737) & (n_n4756) & (n_n4724) & (n_n4759)) + ((n_n4737) & (!n_n4756) & (!n_n4724) & (!n_n4759)) + ((n_n4737) & (!n_n4756) & (!n_n4724) & (n_n4759)) + ((n_n4737) & (!n_n4756) & (n_n4724) & (!n_n4759)) + ((n_n4737) & (!n_n4756) & (n_n4724) & (n_n4759)) + ((n_n4737) & (n_n4756) & (!n_n4724) & (!n_n4759)) + ((n_n4737) & (n_n4756) & (!n_n4724) & (n_n4759)) + ((n_n4737) & (n_n4756) & (n_n4724) & (!n_n4759)) + ((n_n4737) & (n_n4756) & (n_n4724) & (n_n4759)));
	assign x12069x = (((!x483x) & (!x23x) & (!n_n4751) & (!n_n4732) & (x350x)) + ((!x483x) & (!x23x) & (!n_n4751) & (n_n4732) & (!x350x)) + ((!x483x) & (!x23x) & (!n_n4751) & (n_n4732) & (x350x)) + ((!x483x) & (!x23x) & (n_n4751) & (!n_n4732) & (!x350x)) + ((!x483x) & (!x23x) & (n_n4751) & (!n_n4732) & (x350x)) + ((!x483x) & (!x23x) & (n_n4751) & (n_n4732) & (!x350x)) + ((!x483x) & (!x23x) & (n_n4751) & (n_n4732) & (x350x)) + ((!x483x) & (x23x) & (!n_n4751) & (!n_n4732) & (x350x)) + ((!x483x) & (x23x) & (!n_n4751) & (n_n4732) & (!x350x)) + ((!x483x) & (x23x) & (!n_n4751) & (n_n4732) & (x350x)) + ((!x483x) & (x23x) & (n_n4751) & (!n_n4732) & (!x350x)) + ((!x483x) & (x23x) & (n_n4751) & (!n_n4732) & (x350x)) + ((!x483x) & (x23x) & (n_n4751) & (n_n4732) & (!x350x)) + ((!x483x) & (x23x) & (n_n4751) & (n_n4732) & (x350x)) + ((x483x) & (!x23x) & (!n_n4751) & (!n_n4732) & (x350x)) + ((x483x) & (!x23x) & (!n_n4751) & (n_n4732) & (!x350x)) + ((x483x) & (!x23x) & (!n_n4751) & (n_n4732) & (x350x)) + ((x483x) & (!x23x) & (n_n4751) & (!n_n4732) & (!x350x)) + ((x483x) & (!x23x) & (n_n4751) & (!n_n4732) & (x350x)) + ((x483x) & (!x23x) & (n_n4751) & (n_n4732) & (!x350x)) + ((x483x) & (!x23x) & (n_n4751) & (n_n4732) & (x350x)) + ((x483x) & (x23x) & (!n_n4751) & (!n_n4732) & (!x350x)) + ((x483x) & (x23x) & (!n_n4751) & (!n_n4732) & (x350x)) + ((x483x) & (x23x) & (!n_n4751) & (n_n4732) & (!x350x)) + ((x483x) & (x23x) & (!n_n4751) & (n_n4732) & (x350x)) + ((x483x) & (x23x) & (n_n4751) & (!n_n4732) & (!x350x)) + ((x483x) & (x23x) & (n_n4751) & (!n_n4732) & (x350x)) + ((x483x) & (x23x) & (n_n4751) & (n_n4732) & (!x350x)) + ((x483x) & (x23x) & (n_n4751) & (n_n4732) & (x350x)));
	assign n_n4655 = (((!i_9_) & (n_n482) & (n_n528) & (n_n390)));
	assign x12074x = (((!n_n4666) & (!n_n4649) & (!n_n4638) & (n_n4655)) + ((!n_n4666) & (!n_n4649) & (n_n4638) & (!n_n4655)) + ((!n_n4666) & (!n_n4649) & (n_n4638) & (n_n4655)) + ((!n_n4666) & (n_n4649) & (!n_n4638) & (!n_n4655)) + ((!n_n4666) & (n_n4649) & (!n_n4638) & (n_n4655)) + ((!n_n4666) & (n_n4649) & (n_n4638) & (!n_n4655)) + ((!n_n4666) & (n_n4649) & (n_n4638) & (n_n4655)) + ((n_n4666) & (!n_n4649) & (!n_n4638) & (!n_n4655)) + ((n_n4666) & (!n_n4649) & (!n_n4638) & (n_n4655)) + ((n_n4666) & (!n_n4649) & (n_n4638) & (!n_n4655)) + ((n_n4666) & (!n_n4649) & (n_n4638) & (n_n4655)) + ((n_n4666) & (n_n4649) & (!n_n4638) & (!n_n4655)) + ((n_n4666) & (n_n4649) & (!n_n4638) & (n_n4655)) + ((n_n4666) & (n_n4649) & (n_n4638) & (!n_n4655)) + ((n_n4666) & (n_n4649) & (n_n4638) & (n_n4655)));
	assign n_n4712 = (((i_9_) & (n_n518) & (n_n534) & (n_n325)));
	assign n_n4658 = (((i_9_) & (n_n524) & (n_n482) & (n_n390)));
	assign n_n4714 = (((i_9_) & (n_n518) & (n_n532) & (n_n325)));
	assign x12075x = (((!n_n4712) & (!n_n4658) & (!n_n4714) & (!n_n4708) & (n_n4706)) + ((!n_n4712) & (!n_n4658) & (!n_n4714) & (n_n4708) & (!n_n4706)) + ((!n_n4712) & (!n_n4658) & (!n_n4714) & (n_n4708) & (n_n4706)) + ((!n_n4712) & (!n_n4658) & (n_n4714) & (!n_n4708) & (!n_n4706)) + ((!n_n4712) & (!n_n4658) & (n_n4714) & (!n_n4708) & (n_n4706)) + ((!n_n4712) & (!n_n4658) & (n_n4714) & (n_n4708) & (!n_n4706)) + ((!n_n4712) & (!n_n4658) & (n_n4714) & (n_n4708) & (n_n4706)) + ((!n_n4712) & (n_n4658) & (!n_n4714) & (!n_n4708) & (!n_n4706)) + ((!n_n4712) & (n_n4658) & (!n_n4714) & (!n_n4708) & (n_n4706)) + ((!n_n4712) & (n_n4658) & (!n_n4714) & (n_n4708) & (!n_n4706)) + ((!n_n4712) & (n_n4658) & (!n_n4714) & (n_n4708) & (n_n4706)) + ((!n_n4712) & (n_n4658) & (n_n4714) & (!n_n4708) & (!n_n4706)) + ((!n_n4712) & (n_n4658) & (n_n4714) & (!n_n4708) & (n_n4706)) + ((!n_n4712) & (n_n4658) & (n_n4714) & (n_n4708) & (!n_n4706)) + ((!n_n4712) & (n_n4658) & (n_n4714) & (n_n4708) & (n_n4706)) + ((n_n4712) & (!n_n4658) & (!n_n4714) & (!n_n4708) & (!n_n4706)) + ((n_n4712) & (!n_n4658) & (!n_n4714) & (!n_n4708) & (n_n4706)) + ((n_n4712) & (!n_n4658) & (!n_n4714) & (n_n4708) & (!n_n4706)) + ((n_n4712) & (!n_n4658) & (!n_n4714) & (n_n4708) & (n_n4706)) + ((n_n4712) & (!n_n4658) & (n_n4714) & (!n_n4708) & (!n_n4706)) + ((n_n4712) & (!n_n4658) & (n_n4714) & (!n_n4708) & (n_n4706)) + ((n_n4712) & (!n_n4658) & (n_n4714) & (n_n4708) & (!n_n4706)) + ((n_n4712) & (!n_n4658) & (n_n4714) & (n_n4708) & (n_n4706)) + ((n_n4712) & (n_n4658) & (!n_n4714) & (!n_n4708) & (!n_n4706)) + ((n_n4712) & (n_n4658) & (!n_n4714) & (!n_n4708) & (n_n4706)) + ((n_n4712) & (n_n4658) & (!n_n4714) & (n_n4708) & (!n_n4706)) + ((n_n4712) & (n_n4658) & (!n_n4714) & (n_n4708) & (n_n4706)) + ((n_n4712) & (n_n4658) & (n_n4714) & (!n_n4708) & (!n_n4706)) + ((n_n4712) & (n_n4658) & (n_n4714) & (!n_n4708) & (n_n4706)) + ((n_n4712) & (n_n4658) & (n_n4714) & (n_n4708) & (!n_n4706)) + ((n_n4712) & (n_n4658) & (n_n4714) & (n_n4708) & (n_n4706)));
	assign x12082x = (((!n_n4790) & (!n_n4835) & (!n_n4788) & (!n_n4823) & (n_n4806)) + ((!n_n4790) & (!n_n4835) & (!n_n4788) & (n_n4823) & (!n_n4806)) + ((!n_n4790) & (!n_n4835) & (!n_n4788) & (n_n4823) & (n_n4806)) + ((!n_n4790) & (!n_n4835) & (n_n4788) & (!n_n4823) & (!n_n4806)) + ((!n_n4790) & (!n_n4835) & (n_n4788) & (!n_n4823) & (n_n4806)) + ((!n_n4790) & (!n_n4835) & (n_n4788) & (n_n4823) & (!n_n4806)) + ((!n_n4790) & (!n_n4835) & (n_n4788) & (n_n4823) & (n_n4806)) + ((!n_n4790) & (n_n4835) & (!n_n4788) & (!n_n4823) & (!n_n4806)) + ((!n_n4790) & (n_n4835) & (!n_n4788) & (!n_n4823) & (n_n4806)) + ((!n_n4790) & (n_n4835) & (!n_n4788) & (n_n4823) & (!n_n4806)) + ((!n_n4790) & (n_n4835) & (!n_n4788) & (n_n4823) & (n_n4806)) + ((!n_n4790) & (n_n4835) & (n_n4788) & (!n_n4823) & (!n_n4806)) + ((!n_n4790) & (n_n4835) & (n_n4788) & (!n_n4823) & (n_n4806)) + ((!n_n4790) & (n_n4835) & (n_n4788) & (n_n4823) & (!n_n4806)) + ((!n_n4790) & (n_n4835) & (n_n4788) & (n_n4823) & (n_n4806)) + ((n_n4790) & (!n_n4835) & (!n_n4788) & (!n_n4823) & (!n_n4806)) + ((n_n4790) & (!n_n4835) & (!n_n4788) & (!n_n4823) & (n_n4806)) + ((n_n4790) & (!n_n4835) & (!n_n4788) & (n_n4823) & (!n_n4806)) + ((n_n4790) & (!n_n4835) & (!n_n4788) & (n_n4823) & (n_n4806)) + ((n_n4790) & (!n_n4835) & (n_n4788) & (!n_n4823) & (!n_n4806)) + ((n_n4790) & (!n_n4835) & (n_n4788) & (!n_n4823) & (n_n4806)) + ((n_n4790) & (!n_n4835) & (n_n4788) & (n_n4823) & (!n_n4806)) + ((n_n4790) & (!n_n4835) & (n_n4788) & (n_n4823) & (n_n4806)) + ((n_n4790) & (n_n4835) & (!n_n4788) & (!n_n4823) & (!n_n4806)) + ((n_n4790) & (n_n4835) & (!n_n4788) & (!n_n4823) & (n_n4806)) + ((n_n4790) & (n_n4835) & (!n_n4788) & (n_n4823) & (!n_n4806)) + ((n_n4790) & (n_n4835) & (!n_n4788) & (n_n4823) & (n_n4806)) + ((n_n4790) & (n_n4835) & (n_n4788) & (!n_n4823) & (!n_n4806)) + ((n_n4790) & (n_n4835) & (n_n4788) & (!n_n4823) & (n_n4806)) + ((n_n4790) & (n_n4835) & (n_n4788) & (n_n4823) & (!n_n4806)) + ((n_n4790) & (n_n4835) & (n_n4788) & (n_n4823) & (n_n4806)));
	assign n_n4342 = (((i_9_) & (n_n536) & (n_n518) & (n_n520)));
	assign n_n4610 = (((i_9_) & (n_n524) & (n_n390) & (n_n509)));
	assign n_n4676 = (((i_9_) & (n_n390) & (n_n473) & (n_n522)));
	assign n_n5189 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n130) & (x20x)));
	assign n_n5190 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n520) & (x12x)));
	assign n_n5188 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n522) & (x12x)));
	assign x67x = (((!i_9_) & (n_n536) & (n_n532) & (n_n509)) + ((i_9_) & (n_n536) & (n_n532) & (n_n509)));
	assign n_n4353 = (((!i_9_) & (n_n536) & (n_n526) & (n_n509)));
	assign x22196x = (((!n_n4357) & (!n_n4358) & (!n_n4352) & (!n_n4351)));
	assign n_n1120 = (((!n_n4356) & (!x67x) & (!n_n4353) & (!n_n4354) & (!x22196x)) + ((!n_n4356) & (!x67x) & (!n_n4353) & (n_n4354) & (!x22196x)) + ((!n_n4356) & (!x67x) & (!n_n4353) & (n_n4354) & (x22196x)) + ((!n_n4356) & (!x67x) & (n_n4353) & (!n_n4354) & (!x22196x)) + ((!n_n4356) & (!x67x) & (n_n4353) & (!n_n4354) & (x22196x)) + ((!n_n4356) & (!x67x) & (n_n4353) & (n_n4354) & (!x22196x)) + ((!n_n4356) & (!x67x) & (n_n4353) & (n_n4354) & (x22196x)) + ((!n_n4356) & (x67x) & (!n_n4353) & (!n_n4354) & (!x22196x)) + ((!n_n4356) & (x67x) & (!n_n4353) & (!n_n4354) & (x22196x)) + ((!n_n4356) & (x67x) & (!n_n4353) & (n_n4354) & (!x22196x)) + ((!n_n4356) & (x67x) & (!n_n4353) & (n_n4354) & (x22196x)) + ((!n_n4356) & (x67x) & (n_n4353) & (!n_n4354) & (!x22196x)) + ((!n_n4356) & (x67x) & (n_n4353) & (!n_n4354) & (x22196x)) + ((!n_n4356) & (x67x) & (n_n4353) & (n_n4354) & (!x22196x)) + ((!n_n4356) & (x67x) & (n_n4353) & (n_n4354) & (x22196x)) + ((n_n4356) & (!x67x) & (!n_n4353) & (!n_n4354) & (!x22196x)) + ((n_n4356) & (!x67x) & (!n_n4353) & (!n_n4354) & (x22196x)) + ((n_n4356) & (!x67x) & (!n_n4353) & (n_n4354) & (!x22196x)) + ((n_n4356) & (!x67x) & (!n_n4353) & (n_n4354) & (x22196x)) + ((n_n4356) & (!x67x) & (n_n4353) & (!n_n4354) & (!x22196x)) + ((n_n4356) & (!x67x) & (n_n4353) & (!n_n4354) & (x22196x)) + ((n_n4356) & (!x67x) & (n_n4353) & (n_n4354) & (!x22196x)) + ((n_n4356) & (!x67x) & (n_n4353) & (n_n4354) & (x22196x)) + ((n_n4356) & (x67x) & (!n_n4353) & (!n_n4354) & (!x22196x)) + ((n_n4356) & (x67x) & (!n_n4353) & (!n_n4354) & (x22196x)) + ((n_n4356) & (x67x) & (!n_n4353) & (n_n4354) & (!x22196x)) + ((n_n4356) & (x67x) & (!n_n4353) & (n_n4354) & (x22196x)) + ((n_n4356) & (x67x) & (n_n4353) & (!n_n4354) & (!x22196x)) + ((n_n4356) & (x67x) & (n_n4353) & (!n_n4354) & (x22196x)) + ((n_n4356) & (x67x) & (n_n4353) & (n_n4354) & (!x22196x)) + ((n_n4356) & (x67x) & (n_n4353) & (n_n4354) & (x22196x)));
	assign n_n4509 = (((!i_9_) & (n_n455) & (n_n491) & (n_n530)));
	assign x129x = (((!i_9_) & (n_n526) & (n_n455) & (n_n491)) + ((i_9_) & (n_n526) & (n_n455) & (n_n491)));
	assign x308x = (((!i_9_) & (n_n455) & (n_n528) & (n_n491)) + ((i_9_) & (n_n455) & (n_n528) & (n_n491)));
	assign x22163x = (((!n_n4514) & (!n_n4506) & (!n_n4507) & (!n_n4509)));
	assign n_n4622 = (((i_9_) & (n_n528) & (n_n390) & (n_n500)));
	assign x75x = (((i_9_) & (n_n526) & (n_n390) & (n_n500)));
	assign n_n5073 = (((!i_9_) & (n_n526) & (n_n195) & (n_n464)));
	assign n_n4152 = (((!i_9_) & (!n_n524) & (n_n526) & (n_n195) & (n_n464)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n195) & (n_n464)) + ((i_9_) & (!n_n524) & (n_n526) & (n_n195) & (n_n464)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n195) & (n_n464)) + ((i_9_) & (n_n524) & (n_n526) & (n_n195) & (n_n464)));
	assign x11790x = (((!n_n4924) & (!n_n4921) & (!n_n4926) & (n_n4925)) + ((!n_n4924) & (!n_n4921) & (n_n4926) & (!n_n4925)) + ((!n_n4924) & (!n_n4921) & (n_n4926) & (n_n4925)) + ((!n_n4924) & (n_n4921) & (!n_n4926) & (!n_n4925)) + ((!n_n4924) & (n_n4921) & (!n_n4926) & (n_n4925)) + ((!n_n4924) & (n_n4921) & (n_n4926) & (!n_n4925)) + ((!n_n4924) & (n_n4921) & (n_n4926) & (n_n4925)) + ((n_n4924) & (!n_n4921) & (!n_n4926) & (!n_n4925)) + ((n_n4924) & (!n_n4921) & (!n_n4926) & (n_n4925)) + ((n_n4924) & (!n_n4921) & (n_n4926) & (!n_n4925)) + ((n_n4924) & (!n_n4921) & (n_n4926) & (n_n4925)) + ((n_n4924) & (n_n4921) & (!n_n4926) & (!n_n4925)) + ((n_n4924) & (n_n4921) & (!n_n4926) & (n_n4925)) + ((n_n4924) & (n_n4921) & (n_n4926) & (!n_n4925)) + ((n_n4924) & (n_n4921) & (n_n4926) & (n_n4925)));
	assign x11791x = (((!n_n4920) & (!n_n4922) & (!n_n4930) & (!n_n4918) & (n_n4919)) + ((!n_n4920) & (!n_n4922) & (!n_n4930) & (n_n4918) & (!n_n4919)) + ((!n_n4920) & (!n_n4922) & (!n_n4930) & (n_n4918) & (n_n4919)) + ((!n_n4920) & (!n_n4922) & (n_n4930) & (!n_n4918) & (!n_n4919)) + ((!n_n4920) & (!n_n4922) & (n_n4930) & (!n_n4918) & (n_n4919)) + ((!n_n4920) & (!n_n4922) & (n_n4930) & (n_n4918) & (!n_n4919)) + ((!n_n4920) & (!n_n4922) & (n_n4930) & (n_n4918) & (n_n4919)) + ((!n_n4920) & (n_n4922) & (!n_n4930) & (!n_n4918) & (!n_n4919)) + ((!n_n4920) & (n_n4922) & (!n_n4930) & (!n_n4918) & (n_n4919)) + ((!n_n4920) & (n_n4922) & (!n_n4930) & (n_n4918) & (!n_n4919)) + ((!n_n4920) & (n_n4922) & (!n_n4930) & (n_n4918) & (n_n4919)) + ((!n_n4920) & (n_n4922) & (n_n4930) & (!n_n4918) & (!n_n4919)) + ((!n_n4920) & (n_n4922) & (n_n4930) & (!n_n4918) & (n_n4919)) + ((!n_n4920) & (n_n4922) & (n_n4930) & (n_n4918) & (!n_n4919)) + ((!n_n4920) & (n_n4922) & (n_n4930) & (n_n4918) & (n_n4919)) + ((n_n4920) & (!n_n4922) & (!n_n4930) & (!n_n4918) & (!n_n4919)) + ((n_n4920) & (!n_n4922) & (!n_n4930) & (!n_n4918) & (n_n4919)) + ((n_n4920) & (!n_n4922) & (!n_n4930) & (n_n4918) & (!n_n4919)) + ((n_n4920) & (!n_n4922) & (!n_n4930) & (n_n4918) & (n_n4919)) + ((n_n4920) & (!n_n4922) & (n_n4930) & (!n_n4918) & (!n_n4919)) + ((n_n4920) & (!n_n4922) & (n_n4930) & (!n_n4918) & (n_n4919)) + ((n_n4920) & (!n_n4922) & (n_n4930) & (n_n4918) & (!n_n4919)) + ((n_n4920) & (!n_n4922) & (n_n4930) & (n_n4918) & (n_n4919)) + ((n_n4920) & (n_n4922) & (!n_n4930) & (!n_n4918) & (!n_n4919)) + ((n_n4920) & (n_n4922) & (!n_n4930) & (!n_n4918) & (n_n4919)) + ((n_n4920) & (n_n4922) & (!n_n4930) & (n_n4918) & (!n_n4919)) + ((n_n4920) & (n_n4922) & (!n_n4930) & (n_n4918) & (n_n4919)) + ((n_n4920) & (n_n4922) & (n_n4930) & (!n_n4918) & (!n_n4919)) + ((n_n4920) & (n_n4922) & (n_n4930) & (!n_n4918) & (n_n4919)) + ((n_n4920) & (n_n4922) & (n_n4930) & (n_n4918) & (!n_n4919)) + ((n_n4920) & (n_n4922) & (n_n4930) & (n_n4918) & (n_n4919)));
	assign n_n4931 = (((!i_9_) & (n_n524) & (n_n473) & (n_n260)));
	assign n_n4932 = (((i_9_) & (n_n473) & (n_n260) & (n_n522)));
	assign x382x = (((!i_9_) & (n_n473) & (n_n260) & (!n_n522) & (x20x)) + ((!i_9_) & (n_n473) & (n_n260) & (n_n522) & (x20x)) + ((i_9_) & (n_n473) & (n_n260) & (!n_n522) & (x20x)) + ((i_9_) & (n_n473) & (n_n260) & (n_n522) & (!x20x)) + ((i_9_) & (n_n473) & (n_n260) & (n_n522) & (x20x)));
	assign x411x = (((!i_9_) & (n_n532) & (n_n260) & (!n_n530) & (n_n464)) + ((!i_9_) & (n_n532) & (n_n260) & (n_n530) & (n_n464)) + ((i_9_) & (!n_n532) & (n_n260) & (n_n530) & (n_n464)) + ((i_9_) & (n_n532) & (n_n260) & (n_n530) & (n_n464)));
	assign x22175x = (((!n_n4934) & (!n_n4937) & (!n_n4938) & (!n_n4935)));
	assign x11796x = (((!n_n4933) & (!n_n4931) & (!n_n4932) & (!x411x) & (!x22175x)) + ((!n_n4933) & (!n_n4931) & (!n_n4932) & (x411x) & (!x22175x)) + ((!n_n4933) & (!n_n4931) & (!n_n4932) & (x411x) & (x22175x)) + ((!n_n4933) & (!n_n4931) & (n_n4932) & (!x411x) & (!x22175x)) + ((!n_n4933) & (!n_n4931) & (n_n4932) & (!x411x) & (x22175x)) + ((!n_n4933) & (!n_n4931) & (n_n4932) & (x411x) & (!x22175x)) + ((!n_n4933) & (!n_n4931) & (n_n4932) & (x411x) & (x22175x)) + ((!n_n4933) & (n_n4931) & (!n_n4932) & (!x411x) & (!x22175x)) + ((!n_n4933) & (n_n4931) & (!n_n4932) & (!x411x) & (x22175x)) + ((!n_n4933) & (n_n4931) & (!n_n4932) & (x411x) & (!x22175x)) + ((!n_n4933) & (n_n4931) & (!n_n4932) & (x411x) & (x22175x)) + ((!n_n4933) & (n_n4931) & (n_n4932) & (!x411x) & (!x22175x)) + ((!n_n4933) & (n_n4931) & (n_n4932) & (!x411x) & (x22175x)) + ((!n_n4933) & (n_n4931) & (n_n4932) & (x411x) & (!x22175x)) + ((!n_n4933) & (n_n4931) & (n_n4932) & (x411x) & (x22175x)) + ((n_n4933) & (!n_n4931) & (!n_n4932) & (!x411x) & (!x22175x)) + ((n_n4933) & (!n_n4931) & (!n_n4932) & (!x411x) & (x22175x)) + ((n_n4933) & (!n_n4931) & (!n_n4932) & (x411x) & (!x22175x)) + ((n_n4933) & (!n_n4931) & (!n_n4932) & (x411x) & (x22175x)) + ((n_n4933) & (!n_n4931) & (n_n4932) & (!x411x) & (!x22175x)) + ((n_n4933) & (!n_n4931) & (n_n4932) & (!x411x) & (x22175x)) + ((n_n4933) & (!n_n4931) & (n_n4932) & (x411x) & (!x22175x)) + ((n_n4933) & (!n_n4931) & (n_n4932) & (x411x) & (x22175x)) + ((n_n4933) & (n_n4931) & (!n_n4932) & (!x411x) & (!x22175x)) + ((n_n4933) & (n_n4931) & (!n_n4932) & (!x411x) & (x22175x)) + ((n_n4933) & (n_n4931) & (!n_n4932) & (x411x) & (!x22175x)) + ((n_n4933) & (n_n4931) & (!n_n4932) & (x411x) & (x22175x)) + ((n_n4933) & (n_n4931) & (n_n4932) & (!x411x) & (!x22175x)) + ((n_n4933) & (n_n4931) & (n_n4932) & (!x411x) & (x22175x)) + ((n_n4933) & (n_n4931) & (n_n4932) & (x411x) & (!x22175x)) + ((n_n4933) & (n_n4931) & (n_n4932) & (x411x) & (x22175x)));
	assign n_n1026 = (((!n_n1075) & (!x11790x) & (!x11791x) & (x11796x)) + ((!n_n1075) & (!x11790x) & (x11791x) & (!x11796x)) + ((!n_n1075) & (!x11790x) & (x11791x) & (x11796x)) + ((!n_n1075) & (x11790x) & (!x11791x) & (!x11796x)) + ((!n_n1075) & (x11790x) & (!x11791x) & (x11796x)) + ((!n_n1075) & (x11790x) & (x11791x) & (!x11796x)) + ((!n_n1075) & (x11790x) & (x11791x) & (x11796x)) + ((n_n1075) & (!x11790x) & (!x11791x) & (!x11796x)) + ((n_n1075) & (!x11790x) & (!x11791x) & (x11796x)) + ((n_n1075) & (!x11790x) & (x11791x) & (!x11796x)) + ((n_n1075) & (!x11790x) & (x11791x) & (x11796x)) + ((n_n1075) & (x11790x) & (!x11791x) & (!x11796x)) + ((n_n1075) & (x11790x) & (!x11791x) & (x11796x)) + ((n_n1075) & (x11790x) & (x11791x) & (!x11796x)) + ((n_n1075) & (x11790x) & (x11791x) & (x11796x)));
	assign n_n4971 = (((!i_9_) & (n_n518) & (n_n532) & (n_n195)));
	assign x11802x = (((!n_n4958) & (!n_n4956) & (!n_n4968) & (!n_n4962) & (n_n4971)) + ((!n_n4958) & (!n_n4956) & (!n_n4968) & (n_n4962) & (!n_n4971)) + ((!n_n4958) & (!n_n4956) & (!n_n4968) & (n_n4962) & (n_n4971)) + ((!n_n4958) & (!n_n4956) & (n_n4968) & (!n_n4962) & (!n_n4971)) + ((!n_n4958) & (!n_n4956) & (n_n4968) & (!n_n4962) & (n_n4971)) + ((!n_n4958) & (!n_n4956) & (n_n4968) & (n_n4962) & (!n_n4971)) + ((!n_n4958) & (!n_n4956) & (n_n4968) & (n_n4962) & (n_n4971)) + ((!n_n4958) & (n_n4956) & (!n_n4968) & (!n_n4962) & (!n_n4971)) + ((!n_n4958) & (n_n4956) & (!n_n4968) & (!n_n4962) & (n_n4971)) + ((!n_n4958) & (n_n4956) & (!n_n4968) & (n_n4962) & (!n_n4971)) + ((!n_n4958) & (n_n4956) & (!n_n4968) & (n_n4962) & (n_n4971)) + ((!n_n4958) & (n_n4956) & (n_n4968) & (!n_n4962) & (!n_n4971)) + ((!n_n4958) & (n_n4956) & (n_n4968) & (!n_n4962) & (n_n4971)) + ((!n_n4958) & (n_n4956) & (n_n4968) & (n_n4962) & (!n_n4971)) + ((!n_n4958) & (n_n4956) & (n_n4968) & (n_n4962) & (n_n4971)) + ((n_n4958) & (!n_n4956) & (!n_n4968) & (!n_n4962) & (!n_n4971)) + ((n_n4958) & (!n_n4956) & (!n_n4968) & (!n_n4962) & (n_n4971)) + ((n_n4958) & (!n_n4956) & (!n_n4968) & (n_n4962) & (!n_n4971)) + ((n_n4958) & (!n_n4956) & (!n_n4968) & (n_n4962) & (n_n4971)) + ((n_n4958) & (!n_n4956) & (n_n4968) & (!n_n4962) & (!n_n4971)) + ((n_n4958) & (!n_n4956) & (n_n4968) & (!n_n4962) & (n_n4971)) + ((n_n4958) & (!n_n4956) & (n_n4968) & (n_n4962) & (!n_n4971)) + ((n_n4958) & (!n_n4956) & (n_n4968) & (n_n4962) & (n_n4971)) + ((n_n4958) & (n_n4956) & (!n_n4968) & (!n_n4962) & (!n_n4971)) + ((n_n4958) & (n_n4956) & (!n_n4968) & (!n_n4962) & (n_n4971)) + ((n_n4958) & (n_n4956) & (!n_n4968) & (n_n4962) & (!n_n4971)) + ((n_n4958) & (n_n4956) & (!n_n4968) & (n_n4962) & (n_n4971)) + ((n_n4958) & (n_n4956) & (n_n4968) & (!n_n4962) & (!n_n4971)) + ((n_n4958) & (n_n4956) & (n_n4968) & (!n_n4962) & (n_n4971)) + ((n_n4958) & (n_n4956) & (n_n4968) & (n_n4962) & (!n_n4971)) + ((n_n4958) & (n_n4956) & (n_n4968) & (n_n4962) & (n_n4971)));
	assign x68x = (((!i_9_) & (n_n518) & (!n_n532) & (n_n534) & (n_n195)) + ((!i_9_) & (n_n518) & (n_n532) & (n_n534) & (n_n195)) + ((i_9_) & (n_n518) & (n_n532) & (!n_n534) & (n_n195)) + ((i_9_) & (n_n518) & (n_n532) & (n_n534) & (n_n195)));
	assign n_n1071 = (((!n_n4963) & (!n_n4966) & (!x11802x) & (x68x)) + ((!n_n4963) & (!n_n4966) & (x11802x) & (!x68x)) + ((!n_n4963) & (!n_n4966) & (x11802x) & (x68x)) + ((!n_n4963) & (n_n4966) & (!x11802x) & (!x68x)) + ((!n_n4963) & (n_n4966) & (!x11802x) & (x68x)) + ((!n_n4963) & (n_n4966) & (x11802x) & (!x68x)) + ((!n_n4963) & (n_n4966) & (x11802x) & (x68x)) + ((n_n4963) & (!n_n4966) & (!x11802x) & (!x68x)) + ((n_n4963) & (!n_n4966) & (!x11802x) & (x68x)) + ((n_n4963) & (!n_n4966) & (x11802x) & (!x68x)) + ((n_n4963) & (!n_n4966) & (x11802x) & (x68x)) + ((n_n4963) & (n_n4966) & (!x11802x) & (!x68x)) + ((n_n4963) & (n_n4966) & (!x11802x) & (x68x)) + ((n_n4963) & (n_n4966) & (x11802x) & (!x68x)) + ((n_n4963) & (n_n4966) & (x11802x) & (x68x)));
	assign n_n4948 = (((i_9_) & (n_n260) & (n_n522) & (n_n464)));
	assign x11806x = (((!i_9_) & (n_n532) & (!n_n534) & (n_n535) & (n_n195)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n535) & (n_n195)) + ((i_9_) & (!n_n532) & (n_n534) & (n_n535) & (n_n195)) + ((i_9_) & (n_n532) & (!n_n534) & (n_n535) & (n_n195)) + ((i_9_) & (n_n532) & (n_n534) & (n_n535) & (n_n195)));
	assign x22160x = (((!x11x) & (!x531x) & (!n_n4950) & (!n_n4942) & (!n_n4945)) + ((!x11x) & (x531x) & (!n_n4950) & (!n_n4942) & (!n_n4945)) + ((x11x) & (!x531x) & (!n_n4950) & (!n_n4942) & (!n_n4945)));
	assign n_n1072 = (((!x17x) & (!x516x) & (!n_n4948) & (!x11806x) & (!x22160x)) + ((!x17x) & (!x516x) & (!n_n4948) & (x11806x) & (!x22160x)) + ((!x17x) & (!x516x) & (!n_n4948) & (x11806x) & (x22160x)) + ((!x17x) & (!x516x) & (n_n4948) & (!x11806x) & (!x22160x)) + ((!x17x) & (!x516x) & (n_n4948) & (!x11806x) & (x22160x)) + ((!x17x) & (!x516x) & (n_n4948) & (x11806x) & (!x22160x)) + ((!x17x) & (!x516x) & (n_n4948) & (x11806x) & (x22160x)) + ((!x17x) & (x516x) & (!n_n4948) & (!x11806x) & (!x22160x)) + ((!x17x) & (x516x) & (!n_n4948) & (x11806x) & (!x22160x)) + ((!x17x) & (x516x) & (!n_n4948) & (x11806x) & (x22160x)) + ((!x17x) & (x516x) & (n_n4948) & (!x11806x) & (!x22160x)) + ((!x17x) & (x516x) & (n_n4948) & (!x11806x) & (x22160x)) + ((!x17x) & (x516x) & (n_n4948) & (x11806x) & (!x22160x)) + ((!x17x) & (x516x) & (n_n4948) & (x11806x) & (x22160x)) + ((x17x) & (!x516x) & (!n_n4948) & (!x11806x) & (!x22160x)) + ((x17x) & (!x516x) & (!n_n4948) & (x11806x) & (!x22160x)) + ((x17x) & (!x516x) & (!n_n4948) & (x11806x) & (x22160x)) + ((x17x) & (!x516x) & (n_n4948) & (!x11806x) & (!x22160x)) + ((x17x) & (!x516x) & (n_n4948) & (!x11806x) & (x22160x)) + ((x17x) & (!x516x) & (n_n4948) & (x11806x) & (!x22160x)) + ((x17x) & (!x516x) & (n_n4948) & (x11806x) & (x22160x)) + ((x17x) & (x516x) & (!n_n4948) & (!x11806x) & (!x22160x)) + ((x17x) & (x516x) & (!n_n4948) & (!x11806x) & (x22160x)) + ((x17x) & (x516x) & (!n_n4948) & (x11806x) & (!x22160x)) + ((x17x) & (x516x) & (!n_n4948) & (x11806x) & (x22160x)) + ((x17x) & (x516x) & (n_n4948) & (!x11806x) & (!x22160x)) + ((x17x) & (x516x) & (n_n4948) & (!x11806x) & (x22160x)) + ((x17x) & (x516x) & (n_n4948) & (x11806x) & (!x22160x)) + ((x17x) & (x516x) & (n_n4948) & (x11806x) & (x22160x)));
	assign n_n4973 = (((!i_9_) & (n_n518) & (n_n195) & (n_n530)));
	assign x29x = (((!i_9_) & (n_n518) & (!n_n528) & (n_n195) & (n_n530)) + ((!i_9_) & (n_n518) & (n_n528) & (n_n195) & (n_n530)) + ((i_9_) & (n_n518) & (!n_n528) & (n_n195) & (n_n530)) + ((i_9_) & (n_n518) & (n_n528) & (n_n195) & (!n_n530)) + ((i_9_) & (n_n518) & (n_n528) & (n_n195) & (n_n530)));
	assign x11814x = (((!n_n524) & (!n_n518) & (!n_n522) & (!x18x) & (x29x)) + ((!n_n524) & (!n_n518) & (!n_n522) & (x18x) & (x29x)) + ((!n_n524) & (!n_n518) & (n_n522) & (!x18x) & (x29x)) + ((!n_n524) & (!n_n518) & (n_n522) & (x18x) & (x29x)) + ((!n_n524) & (n_n518) & (!n_n522) & (!x18x) & (x29x)) + ((!n_n524) & (n_n518) & (!n_n522) & (x18x) & (x29x)) + ((!n_n524) & (n_n518) & (n_n522) & (!x18x) & (x29x)) + ((!n_n524) & (n_n518) & (n_n522) & (x18x) & (!x29x)) + ((!n_n524) & (n_n518) & (n_n522) & (x18x) & (x29x)) + ((n_n524) & (!n_n518) & (!n_n522) & (!x18x) & (x29x)) + ((n_n524) & (!n_n518) & (!n_n522) & (x18x) & (x29x)) + ((n_n524) & (!n_n518) & (n_n522) & (!x18x) & (x29x)) + ((n_n524) & (!n_n518) & (n_n522) & (x18x) & (x29x)) + ((n_n524) & (n_n518) & (!n_n522) & (!x18x) & (x29x)) + ((n_n524) & (n_n518) & (!n_n522) & (x18x) & (!x29x)) + ((n_n524) & (n_n518) & (!n_n522) & (x18x) & (x29x)) + ((n_n524) & (n_n518) & (n_n522) & (!x18x) & (x29x)) + ((n_n524) & (n_n518) & (n_n522) & (x18x) & (!x29x)) + ((n_n524) & (n_n518) & (n_n522) & (x18x) & (x29x)));
	assign x11815x = (((!n_n4977) & (!n_n4975) & (!n_n4981) & (!n_n4979) & (x11814x)) + ((!n_n4977) & (!n_n4975) & (!n_n4981) & (n_n4979) & (!x11814x)) + ((!n_n4977) & (!n_n4975) & (!n_n4981) & (n_n4979) & (x11814x)) + ((!n_n4977) & (!n_n4975) & (n_n4981) & (!n_n4979) & (!x11814x)) + ((!n_n4977) & (!n_n4975) & (n_n4981) & (!n_n4979) & (x11814x)) + ((!n_n4977) & (!n_n4975) & (n_n4981) & (n_n4979) & (!x11814x)) + ((!n_n4977) & (!n_n4975) & (n_n4981) & (n_n4979) & (x11814x)) + ((!n_n4977) & (n_n4975) & (!n_n4981) & (!n_n4979) & (!x11814x)) + ((!n_n4977) & (n_n4975) & (!n_n4981) & (!n_n4979) & (x11814x)) + ((!n_n4977) & (n_n4975) & (!n_n4981) & (n_n4979) & (!x11814x)) + ((!n_n4977) & (n_n4975) & (!n_n4981) & (n_n4979) & (x11814x)) + ((!n_n4977) & (n_n4975) & (n_n4981) & (!n_n4979) & (!x11814x)) + ((!n_n4977) & (n_n4975) & (n_n4981) & (!n_n4979) & (x11814x)) + ((!n_n4977) & (n_n4975) & (n_n4981) & (n_n4979) & (!x11814x)) + ((!n_n4977) & (n_n4975) & (n_n4981) & (n_n4979) & (x11814x)) + ((n_n4977) & (!n_n4975) & (!n_n4981) & (!n_n4979) & (!x11814x)) + ((n_n4977) & (!n_n4975) & (!n_n4981) & (!n_n4979) & (x11814x)) + ((n_n4977) & (!n_n4975) & (!n_n4981) & (n_n4979) & (!x11814x)) + ((n_n4977) & (!n_n4975) & (!n_n4981) & (n_n4979) & (x11814x)) + ((n_n4977) & (!n_n4975) & (n_n4981) & (!n_n4979) & (!x11814x)) + ((n_n4977) & (!n_n4975) & (n_n4981) & (!n_n4979) & (x11814x)) + ((n_n4977) & (!n_n4975) & (n_n4981) & (n_n4979) & (!x11814x)) + ((n_n4977) & (!n_n4975) & (n_n4981) & (n_n4979) & (x11814x)) + ((n_n4977) & (n_n4975) & (!n_n4981) & (!n_n4979) & (!x11814x)) + ((n_n4977) & (n_n4975) & (!n_n4981) & (!n_n4979) & (x11814x)) + ((n_n4977) & (n_n4975) & (!n_n4981) & (n_n4979) & (!x11814x)) + ((n_n4977) & (n_n4975) & (!n_n4981) & (n_n4979) & (x11814x)) + ((n_n4977) & (n_n4975) & (n_n4981) & (!n_n4979) & (!x11814x)) + ((n_n4977) & (n_n4975) & (n_n4981) & (!n_n4979) & (x11814x)) + ((n_n4977) & (n_n4975) & (n_n4981) & (n_n4979) & (!x11814x)) + ((n_n4977) & (n_n4975) & (n_n4981) & (n_n4979) & (x11814x)));
	assign n_n1985 = (((!n_n260) & (!x20x) & (!n_n500) & (x262x)) + ((!n_n260) & (!x20x) & (n_n500) & (x262x)) + ((!n_n260) & (x20x) & (!n_n500) & (x262x)) + ((!n_n260) & (x20x) & (n_n500) & (x262x)) + ((n_n260) & (!x20x) & (!n_n500) & (x262x)) + ((n_n260) & (!x20x) & (n_n500) & (x262x)) + ((n_n260) & (x20x) & (!n_n500) & (x262x)) + ((n_n260) & (x20x) & (n_n500) & (!x262x)) + ((n_n260) & (x20x) & (n_n500) & (x262x)));
	assign n_n3815 = (((!i_9_) & (n_n532) & (n_n260) & (n_n500) & (!n_n530)) + ((!i_9_) & (n_n532) & (n_n260) & (n_n500) & (n_n530)) + ((i_9_) & (!n_n532) & (n_n260) & (n_n500) & (n_n530)) + ((i_9_) & (n_n532) & (n_n260) & (n_n500) & (!n_n530)) + ((i_9_) & (n_n532) & (n_n260) & (n_n500) & (n_n530)));
	assign n_n1077 = (((!n_n4882) & (!n_n4880) & (!n_n4877) & (!n_n1985) & (n_n3815)) + ((!n_n4882) & (!n_n4880) & (!n_n4877) & (n_n1985) & (!n_n3815)) + ((!n_n4882) & (!n_n4880) & (!n_n4877) & (n_n1985) & (n_n3815)) + ((!n_n4882) & (!n_n4880) & (n_n4877) & (!n_n1985) & (!n_n3815)) + ((!n_n4882) & (!n_n4880) & (n_n4877) & (!n_n1985) & (n_n3815)) + ((!n_n4882) & (!n_n4880) & (n_n4877) & (n_n1985) & (!n_n3815)) + ((!n_n4882) & (!n_n4880) & (n_n4877) & (n_n1985) & (n_n3815)) + ((!n_n4882) & (n_n4880) & (!n_n4877) & (!n_n1985) & (!n_n3815)) + ((!n_n4882) & (n_n4880) & (!n_n4877) & (!n_n1985) & (n_n3815)) + ((!n_n4882) & (n_n4880) & (!n_n4877) & (n_n1985) & (!n_n3815)) + ((!n_n4882) & (n_n4880) & (!n_n4877) & (n_n1985) & (n_n3815)) + ((!n_n4882) & (n_n4880) & (n_n4877) & (!n_n1985) & (!n_n3815)) + ((!n_n4882) & (n_n4880) & (n_n4877) & (!n_n1985) & (n_n3815)) + ((!n_n4882) & (n_n4880) & (n_n4877) & (n_n1985) & (!n_n3815)) + ((!n_n4882) & (n_n4880) & (n_n4877) & (n_n1985) & (n_n3815)) + ((n_n4882) & (!n_n4880) & (!n_n4877) & (!n_n1985) & (!n_n3815)) + ((n_n4882) & (!n_n4880) & (!n_n4877) & (!n_n1985) & (n_n3815)) + ((n_n4882) & (!n_n4880) & (!n_n4877) & (n_n1985) & (!n_n3815)) + ((n_n4882) & (!n_n4880) & (!n_n4877) & (n_n1985) & (n_n3815)) + ((n_n4882) & (!n_n4880) & (n_n4877) & (!n_n1985) & (!n_n3815)) + ((n_n4882) & (!n_n4880) & (n_n4877) & (!n_n1985) & (n_n3815)) + ((n_n4882) & (!n_n4880) & (n_n4877) & (n_n1985) & (!n_n3815)) + ((n_n4882) & (!n_n4880) & (n_n4877) & (n_n1985) & (n_n3815)) + ((n_n4882) & (n_n4880) & (!n_n4877) & (!n_n1985) & (!n_n3815)) + ((n_n4882) & (n_n4880) & (!n_n4877) & (!n_n1985) & (n_n3815)) + ((n_n4882) & (n_n4880) & (!n_n4877) & (n_n1985) & (!n_n3815)) + ((n_n4882) & (n_n4880) & (!n_n4877) & (n_n1985) & (n_n3815)) + ((n_n4882) & (n_n4880) & (n_n4877) & (!n_n1985) & (!n_n3815)) + ((n_n4882) & (n_n4880) & (n_n4877) & (!n_n1985) & (n_n3815)) + ((n_n4882) & (n_n4880) & (n_n4877) & (n_n1985) & (!n_n3815)) + ((n_n4882) & (n_n4880) & (n_n4877) & (n_n1985) & (n_n3815)));
	assign n_n4867 = (((!i_9_) & (n_n524) & (n_n509) & (n_n260)));
	assign x11824x = (((!n_n4863) & (!n_n4865) & (!n_n4864) & (!n_n4873) & (n_n4867)) + ((!n_n4863) & (!n_n4865) & (!n_n4864) & (n_n4873) & (!n_n4867)) + ((!n_n4863) & (!n_n4865) & (!n_n4864) & (n_n4873) & (n_n4867)) + ((!n_n4863) & (!n_n4865) & (n_n4864) & (!n_n4873) & (!n_n4867)) + ((!n_n4863) & (!n_n4865) & (n_n4864) & (!n_n4873) & (n_n4867)) + ((!n_n4863) & (!n_n4865) & (n_n4864) & (n_n4873) & (!n_n4867)) + ((!n_n4863) & (!n_n4865) & (n_n4864) & (n_n4873) & (n_n4867)) + ((!n_n4863) & (n_n4865) & (!n_n4864) & (!n_n4873) & (!n_n4867)) + ((!n_n4863) & (n_n4865) & (!n_n4864) & (!n_n4873) & (n_n4867)) + ((!n_n4863) & (n_n4865) & (!n_n4864) & (n_n4873) & (!n_n4867)) + ((!n_n4863) & (n_n4865) & (!n_n4864) & (n_n4873) & (n_n4867)) + ((!n_n4863) & (n_n4865) & (n_n4864) & (!n_n4873) & (!n_n4867)) + ((!n_n4863) & (n_n4865) & (n_n4864) & (!n_n4873) & (n_n4867)) + ((!n_n4863) & (n_n4865) & (n_n4864) & (n_n4873) & (!n_n4867)) + ((!n_n4863) & (n_n4865) & (n_n4864) & (n_n4873) & (n_n4867)) + ((n_n4863) & (!n_n4865) & (!n_n4864) & (!n_n4873) & (!n_n4867)) + ((n_n4863) & (!n_n4865) & (!n_n4864) & (!n_n4873) & (n_n4867)) + ((n_n4863) & (!n_n4865) & (!n_n4864) & (n_n4873) & (!n_n4867)) + ((n_n4863) & (!n_n4865) & (!n_n4864) & (n_n4873) & (n_n4867)) + ((n_n4863) & (!n_n4865) & (n_n4864) & (!n_n4873) & (!n_n4867)) + ((n_n4863) & (!n_n4865) & (n_n4864) & (!n_n4873) & (n_n4867)) + ((n_n4863) & (!n_n4865) & (n_n4864) & (n_n4873) & (!n_n4867)) + ((n_n4863) & (!n_n4865) & (n_n4864) & (n_n4873) & (n_n4867)) + ((n_n4863) & (n_n4865) & (!n_n4864) & (!n_n4873) & (!n_n4867)) + ((n_n4863) & (n_n4865) & (!n_n4864) & (!n_n4873) & (n_n4867)) + ((n_n4863) & (n_n4865) & (!n_n4864) & (n_n4873) & (!n_n4867)) + ((n_n4863) & (n_n4865) & (!n_n4864) & (n_n4873) & (n_n4867)) + ((n_n4863) & (n_n4865) & (n_n4864) & (!n_n4873) & (!n_n4867)) + ((n_n4863) & (n_n4865) & (n_n4864) & (!n_n4873) & (n_n4867)) + ((n_n4863) & (n_n4865) & (n_n4864) & (n_n4873) & (!n_n4867)) + ((n_n4863) & (n_n4865) & (n_n4864) & (n_n4873) & (n_n4867)));
	assign x226x = (((!i_9_) & (n_n524) & (n_n260) & (!n_n522) & (n_n491)) + ((!i_9_) & (n_n524) & (n_n260) & (n_n522) & (n_n491)) + ((i_9_) & (!n_n524) & (n_n260) & (n_n522) & (n_n491)) + ((i_9_) & (n_n524) & (n_n260) & (n_n522) & (n_n491)));
	assign n_n4892 = (((i_9_) & (n_n260) & (n_n491) & (n_n530)));
	assign x264x = (((!i_7_) & (!i_8_) & (i_6_) & (x17x) & (n_n491)) + ((!i_7_) & (i_8_) & (i_6_) & (x17x) & (n_n491)));
	assign x11830x = (((!n_n4901) & (!n_n4903) & (!n_n4897) & (!x226x) & (x11828x)) + ((!n_n4901) & (!n_n4903) & (!n_n4897) & (x226x) & (!x11828x)) + ((!n_n4901) & (!n_n4903) & (!n_n4897) & (x226x) & (x11828x)) + ((!n_n4901) & (!n_n4903) & (n_n4897) & (!x226x) & (!x11828x)) + ((!n_n4901) & (!n_n4903) & (n_n4897) & (!x226x) & (x11828x)) + ((!n_n4901) & (!n_n4903) & (n_n4897) & (x226x) & (!x11828x)) + ((!n_n4901) & (!n_n4903) & (n_n4897) & (x226x) & (x11828x)) + ((!n_n4901) & (n_n4903) & (!n_n4897) & (!x226x) & (!x11828x)) + ((!n_n4901) & (n_n4903) & (!n_n4897) & (!x226x) & (x11828x)) + ((!n_n4901) & (n_n4903) & (!n_n4897) & (x226x) & (!x11828x)) + ((!n_n4901) & (n_n4903) & (!n_n4897) & (x226x) & (x11828x)) + ((!n_n4901) & (n_n4903) & (n_n4897) & (!x226x) & (!x11828x)) + ((!n_n4901) & (n_n4903) & (n_n4897) & (!x226x) & (x11828x)) + ((!n_n4901) & (n_n4903) & (n_n4897) & (x226x) & (!x11828x)) + ((!n_n4901) & (n_n4903) & (n_n4897) & (x226x) & (x11828x)) + ((n_n4901) & (!n_n4903) & (!n_n4897) & (!x226x) & (!x11828x)) + ((n_n4901) & (!n_n4903) & (!n_n4897) & (!x226x) & (x11828x)) + ((n_n4901) & (!n_n4903) & (!n_n4897) & (x226x) & (!x11828x)) + ((n_n4901) & (!n_n4903) & (!n_n4897) & (x226x) & (x11828x)) + ((n_n4901) & (!n_n4903) & (n_n4897) & (!x226x) & (!x11828x)) + ((n_n4901) & (!n_n4903) & (n_n4897) & (!x226x) & (x11828x)) + ((n_n4901) & (!n_n4903) & (n_n4897) & (x226x) & (!x11828x)) + ((n_n4901) & (!n_n4903) & (n_n4897) & (x226x) & (x11828x)) + ((n_n4901) & (n_n4903) & (!n_n4897) & (!x226x) & (!x11828x)) + ((n_n4901) & (n_n4903) & (!n_n4897) & (!x226x) & (x11828x)) + ((n_n4901) & (n_n4903) & (!n_n4897) & (x226x) & (!x11828x)) + ((n_n4901) & (n_n4903) & (!n_n4897) & (x226x) & (x11828x)) + ((n_n4901) & (n_n4903) & (n_n4897) & (!x226x) & (!x11828x)) + ((n_n4901) & (n_n4903) & (n_n4897) & (!x226x) & (x11828x)) + ((n_n4901) & (n_n4903) & (n_n4897) & (x226x) & (!x11828x)) + ((n_n4901) & (n_n4903) & (n_n4897) & (x226x) & (x11828x)));
	assign x11832x = (((!x294x) & (!x295x) & (!n_n1077) & (!x11824x) & (x11830x)) + ((!x294x) & (!x295x) & (!n_n1077) & (x11824x) & (!x11830x)) + ((!x294x) & (!x295x) & (!n_n1077) & (x11824x) & (x11830x)) + ((!x294x) & (!x295x) & (n_n1077) & (!x11824x) & (!x11830x)) + ((!x294x) & (!x295x) & (n_n1077) & (!x11824x) & (x11830x)) + ((!x294x) & (!x295x) & (n_n1077) & (x11824x) & (!x11830x)) + ((!x294x) & (!x295x) & (n_n1077) & (x11824x) & (x11830x)) + ((!x294x) & (x295x) & (!n_n1077) & (!x11824x) & (!x11830x)) + ((!x294x) & (x295x) & (!n_n1077) & (!x11824x) & (x11830x)) + ((!x294x) & (x295x) & (!n_n1077) & (x11824x) & (!x11830x)) + ((!x294x) & (x295x) & (!n_n1077) & (x11824x) & (x11830x)) + ((!x294x) & (x295x) & (n_n1077) & (!x11824x) & (!x11830x)) + ((!x294x) & (x295x) & (n_n1077) & (!x11824x) & (x11830x)) + ((!x294x) & (x295x) & (n_n1077) & (x11824x) & (!x11830x)) + ((!x294x) & (x295x) & (n_n1077) & (x11824x) & (x11830x)) + ((x294x) & (!x295x) & (!n_n1077) & (!x11824x) & (!x11830x)) + ((x294x) & (!x295x) & (!n_n1077) & (!x11824x) & (x11830x)) + ((x294x) & (!x295x) & (!n_n1077) & (x11824x) & (!x11830x)) + ((x294x) & (!x295x) & (!n_n1077) & (x11824x) & (x11830x)) + ((x294x) & (!x295x) & (n_n1077) & (!x11824x) & (!x11830x)) + ((x294x) & (!x295x) & (n_n1077) & (!x11824x) & (x11830x)) + ((x294x) & (!x295x) & (n_n1077) & (x11824x) & (!x11830x)) + ((x294x) & (!x295x) & (n_n1077) & (x11824x) & (x11830x)) + ((x294x) & (x295x) & (!n_n1077) & (!x11824x) & (!x11830x)) + ((x294x) & (x295x) & (!n_n1077) & (!x11824x) & (x11830x)) + ((x294x) & (x295x) & (!n_n1077) & (x11824x) & (!x11830x)) + ((x294x) & (x295x) & (!n_n1077) & (x11824x) & (x11830x)) + ((x294x) & (x295x) & (n_n1077) & (!x11824x) & (!x11830x)) + ((x294x) & (x295x) & (n_n1077) & (!x11824x) & (x11830x)) + ((x294x) & (x295x) & (n_n1077) & (x11824x) & (!x11830x)) + ((x294x) & (x295x) & (n_n1077) & (x11824x) & (x11830x)));
	assign n_n4349 = (((!i_9_) & (n_n536) & (n_n509) & (n_n530)));
	assign n_n1002 = (((!i_9_) & (n_n536) & (!n_n528) & (n_n509) & (n_n530)) + ((!i_9_) & (n_n536) & (n_n528) & (n_n509) & (n_n530)) + ((i_9_) & (n_n536) & (!n_n528) & (n_n509) & (n_n530)) + ((i_9_) & (n_n536) & (n_n528) & (n_n509) & (!n_n530)) + ((i_9_) & (n_n536) & (n_n528) & (n_n509) & (n_n530)));
	assign n_n5172 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n522) & (x12x)));
	assign n_n4689 = (((!i_9_) & (n_n526) & (n_n390) & (n_n464)));
	assign n_n4697 = (((!i_9_) & (n_n534) & (n_n325) & (n_n535)));
	assign n_n4703 = (((!i_9_) & (n_n528) & (n_n325) & (n_n535)));
	assign n_n4778 = (((i_9_) & (n_n482) & (n_n532) & (n_n325)));
	assign n_n5011 = (((!i_9_) & (n_n524) & (n_n195) & (n_n500)));
	assign n_n5061 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n195) & (x20x)));
	assign n_n5070 = (((i_9_) & (n_n528) & (n_n195) & (n_n464)));
	assign n_n5076 = (((i_9_) & (n_n522) & (n_n195) & (n_n464)));
	assign n_n5135 = (((!i_9_) & (n_n528) & (n_n130) & (n_n500)));
	assign n_n5157 = (((i_5_) & (!i_3_) & (i_4_) & (n_n130) & (x20x)));
	assign n_n5201 = (((!i_9_) & (n_n526) & (n_n130) & (n_n464)));
	assign n_n5207 = (((!i_1_) & (i_2_) & (!i_0_) & (x23x) & (n_n464)));
	assign n_n5237 = (((!i_5_) & (i_3_) & (i_4_) & (x20x) & (n_n65)));
	assign n_n5252 = (((i_5_) & (i_3_) & (!i_4_) & (x19x) & (n_n522)));
	assign n_n4773 = (((!i_1_) & (!i_2_) & (i_0_) & (n_n491) & (x20x)));
	assign n_n4205 = (((!x21x) & (!n_n325) & (!n_n491) & (!x20x) & (n_n4772)) + ((!x21x) & (!n_n325) & (!n_n491) & (x20x) & (n_n4772)) + ((!x21x) & (!n_n325) & (n_n491) & (!x20x) & (n_n4772)) + ((!x21x) & (!n_n325) & (n_n491) & (x20x) & (n_n4772)) + ((!x21x) & (n_n325) & (!n_n491) & (!x20x) & (n_n4772)) + ((!x21x) & (n_n325) & (!n_n491) & (x20x) & (n_n4772)) + ((!x21x) & (n_n325) & (n_n491) & (!x20x) & (n_n4772)) + ((!x21x) & (n_n325) & (n_n491) & (x20x) & (!n_n4772)) + ((!x21x) & (n_n325) & (n_n491) & (x20x) & (n_n4772)) + ((x21x) & (!n_n325) & (!n_n491) & (!x20x) & (n_n4772)) + ((x21x) & (!n_n325) & (!n_n491) & (x20x) & (n_n4772)) + ((x21x) & (!n_n325) & (n_n491) & (!x20x) & (n_n4772)) + ((x21x) & (!n_n325) & (n_n491) & (x20x) & (n_n4772)) + ((x21x) & (n_n325) & (!n_n491) & (!x20x) & (n_n4772)) + ((x21x) & (n_n325) & (!n_n491) & (x20x) & (n_n4772)) + ((x21x) & (n_n325) & (n_n491) & (!x20x) & (!n_n4772)) + ((x21x) & (n_n325) & (n_n491) & (!x20x) & (n_n4772)) + ((x21x) & (n_n325) & (n_n491) & (x20x) & (!n_n4772)) + ((x21x) & (n_n325) & (n_n491) & (x20x) & (n_n4772)));
	assign n_n5024 = (((i_9_) & (n_n526) & (n_n491) & (n_n195)));
	assign x13400x = (((!i_9_) & (n_n528) & (n_n491) & (n_n195)) + ((i_9_) & (n_n528) & (n_n491) & (n_n195)));
	assign n_n4161 = (((!i_9_) & (!n_n526) & (n_n528) & (n_n491) & (n_n195)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n491) & (n_n195)) + ((i_9_) & (!n_n526) & (n_n528) & (n_n491) & (n_n195)) + ((i_9_) & (n_n526) & (!n_n528) & (n_n491) & (n_n195)) + ((i_9_) & (n_n526) & (n_n528) & (n_n491) & (n_n195)));
	assign n_n5084 = (((i_5_) & (i_3_) & (i_4_) & (x12x) & (n_n530)));
	assign n_n5275 = (((!i_9_) & (n_n532) & (n_n491) & (n_n65)));
	assign n_n5276 = (((i_5_) & (!i_3_) & (i_4_) & (x19x) & (n_n530)));
	assign n_n4600 = (((i_9_) & (n_n390) & (n_n534) & (n_n509)));
	assign x45x = (((!i_9_) & (n_n518) & (n_n390) & (!n_n520) & (x23x)) + ((!i_9_) & (n_n518) & (n_n390) & (n_n520) & (x23x)) + ((i_9_) & (n_n518) & (n_n390) & (!n_n520) & (x23x)) + ((i_9_) & (n_n518) & (n_n390) & (n_n520) & (!x23x)) + ((i_9_) & (n_n518) & (n_n390) & (n_n520) & (x23x)));
	assign x22215x = (((!n_n4612) & (!n_n4609) & (!n_n4606) & (!n_n4610)));
	assign n_n4082 = (((!x108x) & (!n_n4600) & (!x45x) & (!x22215x)) + ((!x108x) & (!n_n4600) & (x45x) & (!x22215x)) + ((!x108x) & (!n_n4600) & (x45x) & (x22215x)) + ((!x108x) & (n_n4600) & (!x45x) & (!x22215x)) + ((!x108x) & (n_n4600) & (!x45x) & (x22215x)) + ((!x108x) & (n_n4600) & (x45x) & (!x22215x)) + ((!x108x) & (n_n4600) & (x45x) & (x22215x)) + ((x108x) & (!n_n4600) & (!x45x) & (!x22215x)) + ((x108x) & (!n_n4600) & (!x45x) & (x22215x)) + ((x108x) & (!n_n4600) & (x45x) & (!x22215x)) + ((x108x) & (!n_n4600) & (x45x) & (x22215x)) + ((x108x) & (n_n4600) & (!x45x) & (!x22215x)) + ((x108x) & (n_n4600) & (!x45x) & (x22215x)) + ((x108x) & (n_n4600) & (x45x) & (!x22215x)) + ((x108x) & (n_n4600) & (x45x) & (x22215x)));
	assign n_n4775 = (((!i_1_) & (!i_2_) & (i_0_) & (n_n491) & (x23x)));
	assign n_n4204 = (((!n_n482) & (!n_n534) & (!x14x) & (!n_n4774) & (n_n4775)) + ((!n_n482) & (!n_n534) & (!x14x) & (n_n4774) & (!n_n4775)) + ((!n_n482) & (!n_n534) & (!x14x) & (n_n4774) & (n_n4775)) + ((!n_n482) & (!n_n534) & (x14x) & (!n_n4774) & (n_n4775)) + ((!n_n482) & (!n_n534) & (x14x) & (n_n4774) & (!n_n4775)) + ((!n_n482) & (!n_n534) & (x14x) & (n_n4774) & (n_n4775)) + ((!n_n482) & (n_n534) & (!x14x) & (!n_n4774) & (n_n4775)) + ((!n_n482) & (n_n534) & (!x14x) & (n_n4774) & (!n_n4775)) + ((!n_n482) & (n_n534) & (!x14x) & (n_n4774) & (n_n4775)) + ((!n_n482) & (n_n534) & (x14x) & (!n_n4774) & (n_n4775)) + ((!n_n482) & (n_n534) & (x14x) & (n_n4774) & (!n_n4775)) + ((!n_n482) & (n_n534) & (x14x) & (n_n4774) & (n_n4775)) + ((n_n482) & (!n_n534) & (!x14x) & (!n_n4774) & (n_n4775)) + ((n_n482) & (!n_n534) & (!x14x) & (n_n4774) & (!n_n4775)) + ((n_n482) & (!n_n534) & (!x14x) & (n_n4774) & (n_n4775)) + ((n_n482) & (!n_n534) & (x14x) & (!n_n4774) & (n_n4775)) + ((n_n482) & (!n_n534) & (x14x) & (n_n4774) & (!n_n4775)) + ((n_n482) & (!n_n534) & (x14x) & (n_n4774) & (n_n4775)) + ((n_n482) & (n_n534) & (!x14x) & (!n_n4774) & (n_n4775)) + ((n_n482) & (n_n534) & (!x14x) & (n_n4774) & (!n_n4775)) + ((n_n482) & (n_n534) & (!x14x) & (n_n4774) & (n_n4775)) + ((n_n482) & (n_n534) & (x14x) & (!n_n4774) & (!n_n4775)) + ((n_n482) & (n_n534) & (x14x) & (!n_n4774) & (n_n4775)) + ((n_n482) & (n_n534) & (x14x) & (n_n4774) & (!n_n4775)) + ((n_n482) & (n_n534) & (x14x) & (n_n4774) & (n_n4775)));
	assign x13149x = (((!i_9_) & (n_n528) & (n_n325) & (n_n491) & (!n_n530)) + ((!i_9_) & (n_n528) & (n_n325) & (n_n491) & (n_n530)) + ((i_9_) & (!n_n528) & (n_n325) & (n_n491) & (n_n530)) + ((i_9_) & (n_n528) & (n_n325) & (n_n491) & (!n_n530)) + ((i_9_) & (n_n528) & (n_n325) & (n_n491) & (n_n530)));
	assign n_n4799 = (((!i_9_) & (n_n528) & (n_n473) & (n_n325)));
	assign x22121x = (((!n_n4790) & (!n_n4798) & (!n_n4796) & (!n_n4797)));
	assign n_n4068 = (((!n_n4792) & (!n_n4793) & (!x179x) & (!n_n4799) & (!x22121x)) + ((!n_n4792) & (!n_n4793) & (!x179x) & (n_n4799) & (!x22121x)) + ((!n_n4792) & (!n_n4793) & (!x179x) & (n_n4799) & (x22121x)) + ((!n_n4792) & (!n_n4793) & (x179x) & (!n_n4799) & (!x22121x)) + ((!n_n4792) & (!n_n4793) & (x179x) & (!n_n4799) & (x22121x)) + ((!n_n4792) & (!n_n4793) & (x179x) & (n_n4799) & (!x22121x)) + ((!n_n4792) & (!n_n4793) & (x179x) & (n_n4799) & (x22121x)) + ((!n_n4792) & (n_n4793) & (!x179x) & (!n_n4799) & (!x22121x)) + ((!n_n4792) & (n_n4793) & (!x179x) & (!n_n4799) & (x22121x)) + ((!n_n4792) & (n_n4793) & (!x179x) & (n_n4799) & (!x22121x)) + ((!n_n4792) & (n_n4793) & (!x179x) & (n_n4799) & (x22121x)) + ((!n_n4792) & (n_n4793) & (x179x) & (!n_n4799) & (!x22121x)) + ((!n_n4792) & (n_n4793) & (x179x) & (!n_n4799) & (x22121x)) + ((!n_n4792) & (n_n4793) & (x179x) & (n_n4799) & (!x22121x)) + ((!n_n4792) & (n_n4793) & (x179x) & (n_n4799) & (x22121x)) + ((n_n4792) & (!n_n4793) & (!x179x) & (!n_n4799) & (!x22121x)) + ((n_n4792) & (!n_n4793) & (!x179x) & (!n_n4799) & (x22121x)) + ((n_n4792) & (!n_n4793) & (!x179x) & (n_n4799) & (!x22121x)) + ((n_n4792) & (!n_n4793) & (!x179x) & (n_n4799) & (x22121x)) + ((n_n4792) & (!n_n4793) & (x179x) & (!n_n4799) & (!x22121x)) + ((n_n4792) & (!n_n4793) & (x179x) & (!n_n4799) & (x22121x)) + ((n_n4792) & (!n_n4793) & (x179x) & (n_n4799) & (!x22121x)) + ((n_n4792) & (!n_n4793) & (x179x) & (n_n4799) & (x22121x)) + ((n_n4792) & (n_n4793) & (!x179x) & (!n_n4799) & (!x22121x)) + ((n_n4792) & (n_n4793) & (!x179x) & (!n_n4799) & (x22121x)) + ((n_n4792) & (n_n4793) & (!x179x) & (n_n4799) & (!x22121x)) + ((n_n4792) & (n_n4793) & (!x179x) & (n_n4799) & (x22121x)) + ((n_n4792) & (n_n4793) & (x179x) & (!n_n4799) & (!x22121x)) + ((n_n4792) & (n_n4793) & (x179x) & (!n_n4799) & (x22121x)) + ((n_n4792) & (n_n4793) & (x179x) & (n_n4799) & (!x22121x)) + ((n_n4792) & (n_n4793) & (x179x) & (n_n4799) & (x22121x)));
	assign n_n4197 = (((!i_9_) & (!n_n532) & (n_n534) & (n_n325) & (n_n464)) + ((!i_9_) & (n_n532) & (!n_n534) & (n_n325) & (n_n464)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n325) & (n_n464)) + ((i_9_) & (n_n532) & (!n_n534) & (n_n325) & (n_n464)) + ((i_9_) & (n_n532) & (n_n534) & (n_n325) & (n_n464)));
	assign x390x = (((!x14x) & (!n_n522) & (!n_n464) & (!n_n4819) & (n_n4196)) + ((!x14x) & (!n_n522) & (!n_n464) & (n_n4819) & (!n_n4196)) + ((!x14x) & (!n_n522) & (!n_n464) & (n_n4819) & (n_n4196)) + ((!x14x) & (!n_n522) & (n_n464) & (!n_n4819) & (n_n4196)) + ((!x14x) & (!n_n522) & (n_n464) & (n_n4819) & (!n_n4196)) + ((!x14x) & (!n_n522) & (n_n464) & (n_n4819) & (n_n4196)) + ((!x14x) & (n_n522) & (!n_n464) & (!n_n4819) & (n_n4196)) + ((!x14x) & (n_n522) & (!n_n464) & (n_n4819) & (!n_n4196)) + ((!x14x) & (n_n522) & (!n_n464) & (n_n4819) & (n_n4196)) + ((!x14x) & (n_n522) & (n_n464) & (!n_n4819) & (n_n4196)) + ((!x14x) & (n_n522) & (n_n464) & (n_n4819) & (!n_n4196)) + ((!x14x) & (n_n522) & (n_n464) & (n_n4819) & (n_n4196)) + ((x14x) & (!n_n522) & (!n_n464) & (!n_n4819) & (n_n4196)) + ((x14x) & (!n_n522) & (!n_n464) & (n_n4819) & (!n_n4196)) + ((x14x) & (!n_n522) & (!n_n464) & (n_n4819) & (n_n4196)) + ((x14x) & (!n_n522) & (n_n464) & (!n_n4819) & (n_n4196)) + ((x14x) & (!n_n522) & (n_n464) & (n_n4819) & (!n_n4196)) + ((x14x) & (!n_n522) & (n_n464) & (n_n4819) & (n_n4196)) + ((x14x) & (n_n522) & (!n_n464) & (!n_n4819) & (n_n4196)) + ((x14x) & (n_n522) & (!n_n464) & (n_n4819) & (!n_n4196)) + ((x14x) & (n_n522) & (!n_n464) & (n_n4819) & (n_n4196)) + ((x14x) & (n_n522) & (n_n464) & (!n_n4819) & (!n_n4196)) + ((x14x) & (n_n522) & (n_n464) & (!n_n4819) & (n_n4196)) + ((x14x) & (n_n522) & (n_n464) & (n_n4819) & (!n_n4196)) + ((x14x) & (n_n522) & (n_n464) & (n_n4819) & (n_n4196)));
	assign x13166x = (((!n_n4801) & (!n_n4818) & (!n_n4197) & (x390x)) + ((!n_n4801) & (!n_n4818) & (n_n4197) & (!x390x)) + ((!n_n4801) & (!n_n4818) & (n_n4197) & (x390x)) + ((!n_n4801) & (n_n4818) & (!n_n4197) & (!x390x)) + ((!n_n4801) & (n_n4818) & (!n_n4197) & (x390x)) + ((!n_n4801) & (n_n4818) & (n_n4197) & (!x390x)) + ((!n_n4801) & (n_n4818) & (n_n4197) & (x390x)) + ((n_n4801) & (!n_n4818) & (!n_n4197) & (!x390x)) + ((n_n4801) & (!n_n4818) & (!n_n4197) & (x390x)) + ((n_n4801) & (!n_n4818) & (n_n4197) & (!x390x)) + ((n_n4801) & (!n_n4818) & (n_n4197) & (x390x)) + ((n_n4801) & (n_n4818) & (!n_n4197) & (!x390x)) + ((n_n4801) & (n_n4818) & (!n_n4197) & (x390x)) + ((n_n4801) & (n_n4818) & (n_n4197) & (!x390x)) + ((n_n4801) & (n_n4818) & (n_n4197) & (x390x)));
	assign x395x = (((!i_9_) & (n_n473) & (n_n325) & (!n_n520) & (x20x)) + ((!i_9_) & (n_n473) & (n_n325) & (n_n520) & (x20x)) + ((i_9_) & (n_n473) & (n_n325) & (!n_n520) & (x20x)) + ((i_9_) & (n_n473) & (n_n325) & (n_n520) & (!x20x)) + ((i_9_) & (n_n473) & (n_n325) & (n_n520) & (x20x)));
	assign n_n4065 = (((!x23x) & (!x530x) & (!x388x) & (!x389x) & (x326x)) + ((!x23x) & (!x530x) & (!x388x) & (x389x) & (!x326x)) + ((!x23x) & (!x530x) & (!x388x) & (x389x) & (x326x)) + ((!x23x) & (!x530x) & (x388x) & (!x389x) & (!x326x)) + ((!x23x) & (!x530x) & (x388x) & (!x389x) & (x326x)) + ((!x23x) & (!x530x) & (x388x) & (x389x) & (!x326x)) + ((!x23x) & (!x530x) & (x388x) & (x389x) & (x326x)) + ((!x23x) & (x530x) & (!x388x) & (!x389x) & (x326x)) + ((!x23x) & (x530x) & (!x388x) & (x389x) & (!x326x)) + ((!x23x) & (x530x) & (!x388x) & (x389x) & (x326x)) + ((!x23x) & (x530x) & (x388x) & (!x389x) & (!x326x)) + ((!x23x) & (x530x) & (x388x) & (!x389x) & (x326x)) + ((!x23x) & (x530x) & (x388x) & (x389x) & (!x326x)) + ((!x23x) & (x530x) & (x388x) & (x389x) & (x326x)) + ((x23x) & (!x530x) & (!x388x) & (!x389x) & (x326x)) + ((x23x) & (!x530x) & (!x388x) & (x389x) & (!x326x)) + ((x23x) & (!x530x) & (!x388x) & (x389x) & (x326x)) + ((x23x) & (!x530x) & (x388x) & (!x389x) & (!x326x)) + ((x23x) & (!x530x) & (x388x) & (!x389x) & (x326x)) + ((x23x) & (!x530x) & (x388x) & (x389x) & (!x326x)) + ((x23x) & (!x530x) & (x388x) & (x389x) & (x326x)) + ((x23x) & (x530x) & (!x388x) & (!x389x) & (!x326x)) + ((x23x) & (x530x) & (!x388x) & (!x389x) & (x326x)) + ((x23x) & (x530x) & (!x388x) & (x389x) & (!x326x)) + ((x23x) & (x530x) & (!x388x) & (x389x) & (x326x)) + ((x23x) & (x530x) & (x388x) & (!x389x) & (!x326x)) + ((x23x) & (x530x) & (x388x) & (!x389x) & (x326x)) + ((x23x) & (x530x) & (x388x) & (x389x) & (!x326x)) + ((x23x) & (x530x) & (x388x) & (x389x) & (x326x)));
	assign x13163x = (((!n_n4817) & (!n_n4800) & (!n_n4803) & (n_n4804)) + ((!n_n4817) & (!n_n4800) & (n_n4803) & (!n_n4804)) + ((!n_n4817) & (!n_n4800) & (n_n4803) & (n_n4804)) + ((!n_n4817) & (n_n4800) & (!n_n4803) & (!n_n4804)) + ((!n_n4817) & (n_n4800) & (!n_n4803) & (n_n4804)) + ((!n_n4817) & (n_n4800) & (n_n4803) & (!n_n4804)) + ((!n_n4817) & (n_n4800) & (n_n4803) & (n_n4804)) + ((n_n4817) & (!n_n4800) & (!n_n4803) & (!n_n4804)) + ((n_n4817) & (!n_n4800) & (!n_n4803) & (n_n4804)) + ((n_n4817) & (!n_n4800) & (n_n4803) & (!n_n4804)) + ((n_n4817) & (!n_n4800) & (n_n4803) & (n_n4804)) + ((n_n4817) & (n_n4800) & (!n_n4803) & (!n_n4804)) + ((n_n4817) & (n_n4800) & (!n_n4803) & (n_n4804)) + ((n_n4817) & (n_n4800) & (n_n4803) & (!n_n4804)) + ((n_n4817) & (n_n4800) & (n_n4803) & (n_n4804)));
	assign n_n4010 = (((!x13166x) & (!x395x) & (!x151x) & (!n_n4065) & (x13163x)) + ((!x13166x) & (!x395x) & (!x151x) & (n_n4065) & (!x13163x)) + ((!x13166x) & (!x395x) & (!x151x) & (n_n4065) & (x13163x)) + ((!x13166x) & (!x395x) & (x151x) & (!n_n4065) & (!x13163x)) + ((!x13166x) & (!x395x) & (x151x) & (!n_n4065) & (x13163x)) + ((!x13166x) & (!x395x) & (x151x) & (n_n4065) & (!x13163x)) + ((!x13166x) & (!x395x) & (x151x) & (n_n4065) & (x13163x)) + ((!x13166x) & (x395x) & (!x151x) & (!n_n4065) & (!x13163x)) + ((!x13166x) & (x395x) & (!x151x) & (!n_n4065) & (x13163x)) + ((!x13166x) & (x395x) & (!x151x) & (n_n4065) & (!x13163x)) + ((!x13166x) & (x395x) & (!x151x) & (n_n4065) & (x13163x)) + ((!x13166x) & (x395x) & (x151x) & (!n_n4065) & (!x13163x)) + ((!x13166x) & (x395x) & (x151x) & (!n_n4065) & (x13163x)) + ((!x13166x) & (x395x) & (x151x) & (n_n4065) & (!x13163x)) + ((!x13166x) & (x395x) & (x151x) & (n_n4065) & (x13163x)) + ((x13166x) & (!x395x) & (!x151x) & (!n_n4065) & (!x13163x)) + ((x13166x) & (!x395x) & (!x151x) & (!n_n4065) & (x13163x)) + ((x13166x) & (!x395x) & (!x151x) & (n_n4065) & (!x13163x)) + ((x13166x) & (!x395x) & (!x151x) & (n_n4065) & (x13163x)) + ((x13166x) & (!x395x) & (x151x) & (!n_n4065) & (!x13163x)) + ((x13166x) & (!x395x) & (x151x) & (!n_n4065) & (x13163x)) + ((x13166x) & (!x395x) & (x151x) & (n_n4065) & (!x13163x)) + ((x13166x) & (!x395x) & (x151x) & (n_n4065) & (x13163x)) + ((x13166x) & (x395x) & (!x151x) & (!n_n4065) & (!x13163x)) + ((x13166x) & (x395x) & (!x151x) & (!n_n4065) & (x13163x)) + ((x13166x) & (x395x) & (!x151x) & (n_n4065) & (!x13163x)) + ((x13166x) & (x395x) & (!x151x) & (n_n4065) & (x13163x)) + ((x13166x) & (x395x) & (x151x) & (!n_n4065) & (!x13163x)) + ((x13166x) & (x395x) & (x151x) & (!n_n4065) & (x13163x)) + ((x13166x) & (x395x) & (x151x) & (n_n4065) & (!x13163x)) + ((x13166x) & (x395x) & (x151x) & (n_n4065) & (x13163x)));
	assign x13178x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n260) & (n_n535)) + ((!i_9_) & (n_n524) & (!n_n526) & (n_n260) & (n_n535)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n260) & (n_n535)) + ((i_9_) & (!n_n524) & (n_n526) & (n_n260) & (n_n535)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n260) & (n_n535)) + ((i_9_) & (n_n524) & (n_n526) & (n_n260) & (n_n535)));
	assign x13180x = (((!n_n4843) & (!x177x) & (!n_n4838) & (!n_n4837) & (x13178x)) + ((!n_n4843) & (!x177x) & (!n_n4838) & (n_n4837) & (!x13178x)) + ((!n_n4843) & (!x177x) & (!n_n4838) & (n_n4837) & (x13178x)) + ((!n_n4843) & (!x177x) & (n_n4838) & (!n_n4837) & (!x13178x)) + ((!n_n4843) & (!x177x) & (n_n4838) & (!n_n4837) & (x13178x)) + ((!n_n4843) & (!x177x) & (n_n4838) & (n_n4837) & (!x13178x)) + ((!n_n4843) & (!x177x) & (n_n4838) & (n_n4837) & (x13178x)) + ((!n_n4843) & (x177x) & (!n_n4838) & (!n_n4837) & (!x13178x)) + ((!n_n4843) & (x177x) & (!n_n4838) & (!n_n4837) & (x13178x)) + ((!n_n4843) & (x177x) & (!n_n4838) & (n_n4837) & (!x13178x)) + ((!n_n4843) & (x177x) & (!n_n4838) & (n_n4837) & (x13178x)) + ((!n_n4843) & (x177x) & (n_n4838) & (!n_n4837) & (!x13178x)) + ((!n_n4843) & (x177x) & (n_n4838) & (!n_n4837) & (x13178x)) + ((!n_n4843) & (x177x) & (n_n4838) & (n_n4837) & (!x13178x)) + ((!n_n4843) & (x177x) & (n_n4838) & (n_n4837) & (x13178x)) + ((n_n4843) & (!x177x) & (!n_n4838) & (!n_n4837) & (!x13178x)) + ((n_n4843) & (!x177x) & (!n_n4838) & (!n_n4837) & (x13178x)) + ((n_n4843) & (!x177x) & (!n_n4838) & (n_n4837) & (!x13178x)) + ((n_n4843) & (!x177x) & (!n_n4838) & (n_n4837) & (x13178x)) + ((n_n4843) & (!x177x) & (n_n4838) & (!n_n4837) & (!x13178x)) + ((n_n4843) & (!x177x) & (n_n4838) & (!n_n4837) & (x13178x)) + ((n_n4843) & (!x177x) & (n_n4838) & (n_n4837) & (!x13178x)) + ((n_n4843) & (!x177x) & (n_n4838) & (n_n4837) & (x13178x)) + ((n_n4843) & (x177x) & (!n_n4838) & (!n_n4837) & (!x13178x)) + ((n_n4843) & (x177x) & (!n_n4838) & (!n_n4837) & (x13178x)) + ((n_n4843) & (x177x) & (!n_n4838) & (n_n4837) & (!x13178x)) + ((n_n4843) & (x177x) & (!n_n4838) & (n_n4837) & (x13178x)) + ((n_n4843) & (x177x) & (n_n4838) & (!n_n4837) & (!x13178x)) + ((n_n4843) & (x177x) & (n_n4838) & (!n_n4837) & (x13178x)) + ((n_n4843) & (x177x) & (n_n4838) & (n_n4837) & (!x13178x)) + ((n_n4843) & (x177x) & (n_n4838) & (n_n4837) & (x13178x)));
	assign n_n4063 = (((!n_n4847) & (!x277x) & (!x176x) & (!n_n4851) & (n_n834)) + ((!n_n4847) & (!x277x) & (!x176x) & (n_n4851) & (!n_n834)) + ((!n_n4847) & (!x277x) & (!x176x) & (n_n4851) & (n_n834)) + ((!n_n4847) & (!x277x) & (x176x) & (!n_n4851) & (!n_n834)) + ((!n_n4847) & (!x277x) & (x176x) & (!n_n4851) & (n_n834)) + ((!n_n4847) & (!x277x) & (x176x) & (n_n4851) & (!n_n834)) + ((!n_n4847) & (!x277x) & (x176x) & (n_n4851) & (n_n834)) + ((!n_n4847) & (x277x) & (!x176x) & (!n_n4851) & (!n_n834)) + ((!n_n4847) & (x277x) & (!x176x) & (!n_n4851) & (n_n834)) + ((!n_n4847) & (x277x) & (!x176x) & (n_n4851) & (!n_n834)) + ((!n_n4847) & (x277x) & (!x176x) & (n_n4851) & (n_n834)) + ((!n_n4847) & (x277x) & (x176x) & (!n_n4851) & (!n_n834)) + ((!n_n4847) & (x277x) & (x176x) & (!n_n4851) & (n_n834)) + ((!n_n4847) & (x277x) & (x176x) & (n_n4851) & (!n_n834)) + ((!n_n4847) & (x277x) & (x176x) & (n_n4851) & (n_n834)) + ((n_n4847) & (!x277x) & (!x176x) & (!n_n4851) & (!n_n834)) + ((n_n4847) & (!x277x) & (!x176x) & (!n_n4851) & (n_n834)) + ((n_n4847) & (!x277x) & (!x176x) & (n_n4851) & (!n_n834)) + ((n_n4847) & (!x277x) & (!x176x) & (n_n4851) & (n_n834)) + ((n_n4847) & (!x277x) & (x176x) & (!n_n4851) & (!n_n834)) + ((n_n4847) & (!x277x) & (x176x) & (!n_n4851) & (n_n834)) + ((n_n4847) & (!x277x) & (x176x) & (n_n4851) & (!n_n834)) + ((n_n4847) & (!x277x) & (x176x) & (n_n4851) & (n_n834)) + ((n_n4847) & (x277x) & (!x176x) & (!n_n4851) & (!n_n834)) + ((n_n4847) & (x277x) & (!x176x) & (!n_n4851) & (n_n834)) + ((n_n4847) & (x277x) & (!x176x) & (n_n4851) & (!n_n834)) + ((n_n4847) & (x277x) & (!x176x) & (n_n4851) & (n_n834)) + ((n_n4847) & (x277x) & (x176x) & (!n_n4851) & (!n_n834)) + ((n_n4847) & (x277x) & (x176x) & (!n_n4851) & (n_n834)) + ((n_n4847) & (x277x) & (x176x) & (n_n4851) & (!n_n834)) + ((n_n4847) & (x277x) & (x176x) & (n_n4851) & (n_n834)));
	assign n_n4009 = (((!x102x) & (!x245x) & (!x13171x) & (!x13180x) & (n_n4063)) + ((!x102x) & (!x245x) & (!x13171x) & (x13180x) & (!n_n4063)) + ((!x102x) & (!x245x) & (!x13171x) & (x13180x) & (n_n4063)) + ((!x102x) & (!x245x) & (x13171x) & (!x13180x) & (!n_n4063)) + ((!x102x) & (!x245x) & (x13171x) & (!x13180x) & (n_n4063)) + ((!x102x) & (!x245x) & (x13171x) & (x13180x) & (!n_n4063)) + ((!x102x) & (!x245x) & (x13171x) & (x13180x) & (n_n4063)) + ((!x102x) & (x245x) & (!x13171x) & (!x13180x) & (!n_n4063)) + ((!x102x) & (x245x) & (!x13171x) & (!x13180x) & (n_n4063)) + ((!x102x) & (x245x) & (!x13171x) & (x13180x) & (!n_n4063)) + ((!x102x) & (x245x) & (!x13171x) & (x13180x) & (n_n4063)) + ((!x102x) & (x245x) & (x13171x) & (!x13180x) & (!n_n4063)) + ((!x102x) & (x245x) & (x13171x) & (!x13180x) & (n_n4063)) + ((!x102x) & (x245x) & (x13171x) & (x13180x) & (!n_n4063)) + ((!x102x) & (x245x) & (x13171x) & (x13180x) & (n_n4063)) + ((x102x) & (!x245x) & (!x13171x) & (!x13180x) & (!n_n4063)) + ((x102x) & (!x245x) & (!x13171x) & (!x13180x) & (n_n4063)) + ((x102x) & (!x245x) & (!x13171x) & (x13180x) & (!n_n4063)) + ((x102x) & (!x245x) & (!x13171x) & (x13180x) & (n_n4063)) + ((x102x) & (!x245x) & (x13171x) & (!x13180x) & (!n_n4063)) + ((x102x) & (!x245x) & (x13171x) & (!x13180x) & (n_n4063)) + ((x102x) & (!x245x) & (x13171x) & (x13180x) & (!n_n4063)) + ((x102x) & (!x245x) & (x13171x) & (x13180x) & (n_n4063)) + ((x102x) & (x245x) & (!x13171x) & (!x13180x) & (!n_n4063)) + ((x102x) & (x245x) & (!x13171x) & (!x13180x) & (n_n4063)) + ((x102x) & (x245x) & (!x13171x) & (x13180x) & (!n_n4063)) + ((x102x) & (x245x) & (!x13171x) & (x13180x) & (n_n4063)) + ((x102x) & (x245x) & (x13171x) & (!x13180x) & (!n_n4063)) + ((x102x) & (x245x) & (x13171x) & (!x13180x) & (n_n4063)) + ((x102x) & (x245x) & (x13171x) & (x13180x) & (!n_n4063)) + ((x102x) & (x245x) & (x13171x) & (x13180x) & (n_n4063)));
	assign x12394x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n325) & (n_n491)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n325) & (n_n491)) + ((i_9_) & (!n_n524) & (n_n526) & (n_n325) & (n_n491)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n325) & (n_n491)) + ((i_9_) & (n_n524) & (n_n526) & (n_n325) & (n_n491)));
	assign x13186x = (((!n_n4779) & (!x131x) & (!n_n4789) & (!n_n4204) & (x13182x)) + ((!n_n4779) & (!x131x) & (!n_n4789) & (n_n4204) & (!x13182x)) + ((!n_n4779) & (!x131x) & (!n_n4789) & (n_n4204) & (x13182x)) + ((!n_n4779) & (!x131x) & (n_n4789) & (!n_n4204) & (!x13182x)) + ((!n_n4779) & (!x131x) & (n_n4789) & (!n_n4204) & (x13182x)) + ((!n_n4779) & (!x131x) & (n_n4789) & (n_n4204) & (!x13182x)) + ((!n_n4779) & (!x131x) & (n_n4789) & (n_n4204) & (x13182x)) + ((!n_n4779) & (x131x) & (!n_n4789) & (!n_n4204) & (!x13182x)) + ((!n_n4779) & (x131x) & (!n_n4789) & (!n_n4204) & (x13182x)) + ((!n_n4779) & (x131x) & (!n_n4789) & (n_n4204) & (!x13182x)) + ((!n_n4779) & (x131x) & (!n_n4789) & (n_n4204) & (x13182x)) + ((!n_n4779) & (x131x) & (n_n4789) & (!n_n4204) & (!x13182x)) + ((!n_n4779) & (x131x) & (n_n4789) & (!n_n4204) & (x13182x)) + ((!n_n4779) & (x131x) & (n_n4789) & (n_n4204) & (!x13182x)) + ((!n_n4779) & (x131x) & (n_n4789) & (n_n4204) & (x13182x)) + ((n_n4779) & (!x131x) & (!n_n4789) & (!n_n4204) & (!x13182x)) + ((n_n4779) & (!x131x) & (!n_n4789) & (!n_n4204) & (x13182x)) + ((n_n4779) & (!x131x) & (!n_n4789) & (n_n4204) & (!x13182x)) + ((n_n4779) & (!x131x) & (!n_n4789) & (n_n4204) & (x13182x)) + ((n_n4779) & (!x131x) & (n_n4789) & (!n_n4204) & (!x13182x)) + ((n_n4779) & (!x131x) & (n_n4789) & (!n_n4204) & (x13182x)) + ((n_n4779) & (!x131x) & (n_n4789) & (n_n4204) & (!x13182x)) + ((n_n4779) & (!x131x) & (n_n4789) & (n_n4204) & (x13182x)) + ((n_n4779) & (x131x) & (!n_n4789) & (!n_n4204) & (!x13182x)) + ((n_n4779) & (x131x) & (!n_n4789) & (!n_n4204) & (x13182x)) + ((n_n4779) & (x131x) & (!n_n4789) & (n_n4204) & (!x13182x)) + ((n_n4779) & (x131x) & (!n_n4789) & (n_n4204) & (x13182x)) + ((n_n4779) & (x131x) & (n_n4789) & (!n_n4204) & (!x13182x)) + ((n_n4779) & (x131x) & (n_n4789) & (!n_n4204) & (x13182x)) + ((n_n4779) & (x131x) & (n_n4789) & (n_n4204) & (!x13182x)) + ((n_n4779) & (x131x) & (n_n4789) & (n_n4204) & (x13182x)));
	assign x13188x = (((!n_n4205) & (!x13149x) & (!n_n4068) & (!x12394x) & (x13186x)) + ((!n_n4205) & (!x13149x) & (!n_n4068) & (x12394x) & (!x13186x)) + ((!n_n4205) & (!x13149x) & (!n_n4068) & (x12394x) & (x13186x)) + ((!n_n4205) & (!x13149x) & (n_n4068) & (!x12394x) & (!x13186x)) + ((!n_n4205) & (!x13149x) & (n_n4068) & (!x12394x) & (x13186x)) + ((!n_n4205) & (!x13149x) & (n_n4068) & (x12394x) & (!x13186x)) + ((!n_n4205) & (!x13149x) & (n_n4068) & (x12394x) & (x13186x)) + ((!n_n4205) & (x13149x) & (!n_n4068) & (!x12394x) & (!x13186x)) + ((!n_n4205) & (x13149x) & (!n_n4068) & (!x12394x) & (x13186x)) + ((!n_n4205) & (x13149x) & (!n_n4068) & (x12394x) & (!x13186x)) + ((!n_n4205) & (x13149x) & (!n_n4068) & (x12394x) & (x13186x)) + ((!n_n4205) & (x13149x) & (n_n4068) & (!x12394x) & (!x13186x)) + ((!n_n4205) & (x13149x) & (n_n4068) & (!x12394x) & (x13186x)) + ((!n_n4205) & (x13149x) & (n_n4068) & (x12394x) & (!x13186x)) + ((!n_n4205) & (x13149x) & (n_n4068) & (x12394x) & (x13186x)) + ((n_n4205) & (!x13149x) & (!n_n4068) & (!x12394x) & (!x13186x)) + ((n_n4205) & (!x13149x) & (!n_n4068) & (!x12394x) & (x13186x)) + ((n_n4205) & (!x13149x) & (!n_n4068) & (x12394x) & (!x13186x)) + ((n_n4205) & (!x13149x) & (!n_n4068) & (x12394x) & (x13186x)) + ((n_n4205) & (!x13149x) & (n_n4068) & (!x12394x) & (!x13186x)) + ((n_n4205) & (!x13149x) & (n_n4068) & (!x12394x) & (x13186x)) + ((n_n4205) & (!x13149x) & (n_n4068) & (x12394x) & (!x13186x)) + ((n_n4205) & (!x13149x) & (n_n4068) & (x12394x) & (x13186x)) + ((n_n4205) & (x13149x) & (!n_n4068) & (!x12394x) & (!x13186x)) + ((n_n4205) & (x13149x) & (!n_n4068) & (!x12394x) & (x13186x)) + ((n_n4205) & (x13149x) & (!n_n4068) & (x12394x) & (!x13186x)) + ((n_n4205) & (x13149x) & (!n_n4068) & (x12394x) & (x13186x)) + ((n_n4205) & (x13149x) & (n_n4068) & (!x12394x) & (!x13186x)) + ((n_n4205) & (x13149x) & (n_n4068) & (!x12394x) & (x13186x)) + ((n_n4205) & (x13149x) & (n_n4068) & (x12394x) & (!x13186x)) + ((n_n4205) & (x13149x) & (n_n4068) & (x12394x) & (x13186x)));
	assign n_n4889 = (((!i_9_) & (n_n534) & (n_n260) & (n_n491)));
	assign x22127x = (((!n_n4887) & (!n_n4885) & (!n_n4882) & (!n_n4883) & (!n_n4886)));
	assign n_n4060 = (((!n_n4878) & (!n_n4880) & (!n_n4879) & (!n_n4889) & (!x22127x)) + ((!n_n4878) & (!n_n4880) & (!n_n4879) & (n_n4889) & (!x22127x)) + ((!n_n4878) & (!n_n4880) & (!n_n4879) & (n_n4889) & (x22127x)) + ((!n_n4878) & (!n_n4880) & (n_n4879) & (!n_n4889) & (!x22127x)) + ((!n_n4878) & (!n_n4880) & (n_n4879) & (!n_n4889) & (x22127x)) + ((!n_n4878) & (!n_n4880) & (n_n4879) & (n_n4889) & (!x22127x)) + ((!n_n4878) & (!n_n4880) & (n_n4879) & (n_n4889) & (x22127x)) + ((!n_n4878) & (n_n4880) & (!n_n4879) & (!n_n4889) & (!x22127x)) + ((!n_n4878) & (n_n4880) & (!n_n4879) & (!n_n4889) & (x22127x)) + ((!n_n4878) & (n_n4880) & (!n_n4879) & (n_n4889) & (!x22127x)) + ((!n_n4878) & (n_n4880) & (!n_n4879) & (n_n4889) & (x22127x)) + ((!n_n4878) & (n_n4880) & (n_n4879) & (!n_n4889) & (!x22127x)) + ((!n_n4878) & (n_n4880) & (n_n4879) & (!n_n4889) & (x22127x)) + ((!n_n4878) & (n_n4880) & (n_n4879) & (n_n4889) & (!x22127x)) + ((!n_n4878) & (n_n4880) & (n_n4879) & (n_n4889) & (x22127x)) + ((n_n4878) & (!n_n4880) & (!n_n4879) & (!n_n4889) & (!x22127x)) + ((n_n4878) & (!n_n4880) & (!n_n4879) & (!n_n4889) & (x22127x)) + ((n_n4878) & (!n_n4880) & (!n_n4879) & (n_n4889) & (!x22127x)) + ((n_n4878) & (!n_n4880) & (!n_n4879) & (n_n4889) & (x22127x)) + ((n_n4878) & (!n_n4880) & (n_n4879) & (!n_n4889) & (!x22127x)) + ((n_n4878) & (!n_n4880) & (n_n4879) & (!n_n4889) & (x22127x)) + ((n_n4878) & (!n_n4880) & (n_n4879) & (n_n4889) & (!x22127x)) + ((n_n4878) & (!n_n4880) & (n_n4879) & (n_n4889) & (x22127x)) + ((n_n4878) & (n_n4880) & (!n_n4879) & (!n_n4889) & (!x22127x)) + ((n_n4878) & (n_n4880) & (!n_n4879) & (!n_n4889) & (x22127x)) + ((n_n4878) & (n_n4880) & (!n_n4879) & (n_n4889) & (!x22127x)) + ((n_n4878) & (n_n4880) & (!n_n4879) & (n_n4889) & (x22127x)) + ((n_n4878) & (n_n4880) & (n_n4879) & (!n_n4889) & (!x22127x)) + ((n_n4878) & (n_n4880) & (n_n4879) & (!n_n4889) & (x22127x)) + ((n_n4878) & (n_n4880) & (n_n4879) & (n_n4889) & (!x22127x)) + ((n_n4878) & (n_n4880) & (n_n4879) & (n_n4889) & (x22127x)));
	assign n_n4891 = (((!i_9_) & (n_n532) & (n_n260) & (n_n491)));
	assign x13199x = (((!n_n4900) & (!n_n4902) & (!n_n4894) & (!n_n4897) & (n_n4891)) + ((!n_n4900) & (!n_n4902) & (!n_n4894) & (n_n4897) & (!n_n4891)) + ((!n_n4900) & (!n_n4902) & (!n_n4894) & (n_n4897) & (n_n4891)) + ((!n_n4900) & (!n_n4902) & (n_n4894) & (!n_n4897) & (!n_n4891)) + ((!n_n4900) & (!n_n4902) & (n_n4894) & (!n_n4897) & (n_n4891)) + ((!n_n4900) & (!n_n4902) & (n_n4894) & (n_n4897) & (!n_n4891)) + ((!n_n4900) & (!n_n4902) & (n_n4894) & (n_n4897) & (n_n4891)) + ((!n_n4900) & (n_n4902) & (!n_n4894) & (!n_n4897) & (!n_n4891)) + ((!n_n4900) & (n_n4902) & (!n_n4894) & (!n_n4897) & (n_n4891)) + ((!n_n4900) & (n_n4902) & (!n_n4894) & (n_n4897) & (!n_n4891)) + ((!n_n4900) & (n_n4902) & (!n_n4894) & (n_n4897) & (n_n4891)) + ((!n_n4900) & (n_n4902) & (n_n4894) & (!n_n4897) & (!n_n4891)) + ((!n_n4900) & (n_n4902) & (n_n4894) & (!n_n4897) & (n_n4891)) + ((!n_n4900) & (n_n4902) & (n_n4894) & (n_n4897) & (!n_n4891)) + ((!n_n4900) & (n_n4902) & (n_n4894) & (n_n4897) & (n_n4891)) + ((n_n4900) & (!n_n4902) & (!n_n4894) & (!n_n4897) & (!n_n4891)) + ((n_n4900) & (!n_n4902) & (!n_n4894) & (!n_n4897) & (n_n4891)) + ((n_n4900) & (!n_n4902) & (!n_n4894) & (n_n4897) & (!n_n4891)) + ((n_n4900) & (!n_n4902) & (!n_n4894) & (n_n4897) & (n_n4891)) + ((n_n4900) & (!n_n4902) & (n_n4894) & (!n_n4897) & (!n_n4891)) + ((n_n4900) & (!n_n4902) & (n_n4894) & (!n_n4897) & (n_n4891)) + ((n_n4900) & (!n_n4902) & (n_n4894) & (n_n4897) & (!n_n4891)) + ((n_n4900) & (!n_n4902) & (n_n4894) & (n_n4897) & (n_n4891)) + ((n_n4900) & (n_n4902) & (!n_n4894) & (!n_n4897) & (!n_n4891)) + ((n_n4900) & (n_n4902) & (!n_n4894) & (!n_n4897) & (n_n4891)) + ((n_n4900) & (n_n4902) & (!n_n4894) & (n_n4897) & (!n_n4891)) + ((n_n4900) & (n_n4902) & (!n_n4894) & (n_n4897) & (n_n4891)) + ((n_n4900) & (n_n4902) & (n_n4894) & (!n_n4897) & (!n_n4891)) + ((n_n4900) & (n_n4902) & (n_n4894) & (!n_n4897) & (n_n4891)) + ((n_n4900) & (n_n4902) & (n_n4894) & (n_n4897) & (!n_n4891)) + ((n_n4900) & (n_n4902) & (n_n4894) & (n_n4897) & (n_n4891)));
	assign n_n1592 = (((!x25x) & (!n_n473) & (!n_n260) & (!n_n4918) & (n_n4919)) + ((!x25x) & (!n_n473) & (!n_n260) & (n_n4918) & (!n_n4919)) + ((!x25x) & (!n_n473) & (!n_n260) & (n_n4918) & (n_n4919)) + ((!x25x) & (!n_n473) & (n_n260) & (!n_n4918) & (n_n4919)) + ((!x25x) & (!n_n473) & (n_n260) & (n_n4918) & (!n_n4919)) + ((!x25x) & (!n_n473) & (n_n260) & (n_n4918) & (n_n4919)) + ((!x25x) & (n_n473) & (!n_n260) & (!n_n4918) & (n_n4919)) + ((!x25x) & (n_n473) & (!n_n260) & (n_n4918) & (!n_n4919)) + ((!x25x) & (n_n473) & (!n_n260) & (n_n4918) & (n_n4919)) + ((!x25x) & (n_n473) & (n_n260) & (!n_n4918) & (n_n4919)) + ((!x25x) & (n_n473) & (n_n260) & (n_n4918) & (!n_n4919)) + ((!x25x) & (n_n473) & (n_n260) & (n_n4918) & (n_n4919)) + ((x25x) & (!n_n473) & (!n_n260) & (!n_n4918) & (n_n4919)) + ((x25x) & (!n_n473) & (!n_n260) & (n_n4918) & (!n_n4919)) + ((x25x) & (!n_n473) & (!n_n260) & (n_n4918) & (n_n4919)) + ((x25x) & (!n_n473) & (n_n260) & (!n_n4918) & (n_n4919)) + ((x25x) & (!n_n473) & (n_n260) & (n_n4918) & (!n_n4919)) + ((x25x) & (!n_n473) & (n_n260) & (n_n4918) & (n_n4919)) + ((x25x) & (n_n473) & (!n_n260) & (!n_n4918) & (n_n4919)) + ((x25x) & (n_n473) & (!n_n260) & (n_n4918) & (!n_n4919)) + ((x25x) & (n_n473) & (!n_n260) & (n_n4918) & (n_n4919)) + ((x25x) & (n_n473) & (n_n260) & (!n_n4918) & (!n_n4919)) + ((x25x) & (n_n473) & (n_n260) & (!n_n4918) & (n_n4919)) + ((x25x) & (n_n473) & (n_n260) & (n_n4918) & (!n_n4919)) + ((x25x) & (n_n473) & (n_n260) & (n_n4918) & (n_n4919)));
	assign x42x = (((!i_9_) & (n_n473) & (n_n532) & (n_n260)) + ((i_9_) & (n_n473) & (n_n532) & (n_n260)));
	assign x13213x = (((!n_n4926) & (!n_n4925) & (!x31x) & (!n_n1592) & (x42x)) + ((!n_n4926) & (!n_n4925) & (!x31x) & (n_n1592) & (!x42x)) + ((!n_n4926) & (!n_n4925) & (!x31x) & (n_n1592) & (x42x)) + ((!n_n4926) & (!n_n4925) & (x31x) & (!n_n1592) & (!x42x)) + ((!n_n4926) & (!n_n4925) & (x31x) & (!n_n1592) & (x42x)) + ((!n_n4926) & (!n_n4925) & (x31x) & (n_n1592) & (!x42x)) + ((!n_n4926) & (!n_n4925) & (x31x) & (n_n1592) & (x42x)) + ((!n_n4926) & (n_n4925) & (!x31x) & (!n_n1592) & (!x42x)) + ((!n_n4926) & (n_n4925) & (!x31x) & (!n_n1592) & (x42x)) + ((!n_n4926) & (n_n4925) & (!x31x) & (n_n1592) & (!x42x)) + ((!n_n4926) & (n_n4925) & (!x31x) & (n_n1592) & (x42x)) + ((!n_n4926) & (n_n4925) & (x31x) & (!n_n1592) & (!x42x)) + ((!n_n4926) & (n_n4925) & (x31x) & (!n_n1592) & (x42x)) + ((!n_n4926) & (n_n4925) & (x31x) & (n_n1592) & (!x42x)) + ((!n_n4926) & (n_n4925) & (x31x) & (n_n1592) & (x42x)) + ((n_n4926) & (!n_n4925) & (!x31x) & (!n_n1592) & (!x42x)) + ((n_n4926) & (!n_n4925) & (!x31x) & (!n_n1592) & (x42x)) + ((n_n4926) & (!n_n4925) & (!x31x) & (n_n1592) & (!x42x)) + ((n_n4926) & (!n_n4925) & (!x31x) & (n_n1592) & (x42x)) + ((n_n4926) & (!n_n4925) & (x31x) & (!n_n1592) & (!x42x)) + ((n_n4926) & (!n_n4925) & (x31x) & (!n_n1592) & (x42x)) + ((n_n4926) & (!n_n4925) & (x31x) & (n_n1592) & (!x42x)) + ((n_n4926) & (!n_n4925) & (x31x) & (n_n1592) & (x42x)) + ((n_n4926) & (n_n4925) & (!x31x) & (!n_n1592) & (!x42x)) + ((n_n4926) & (n_n4925) & (!x31x) & (!n_n1592) & (x42x)) + ((n_n4926) & (n_n4925) & (!x31x) & (n_n1592) & (!x42x)) + ((n_n4926) & (n_n4925) & (!x31x) & (n_n1592) & (x42x)) + ((n_n4926) & (n_n4925) & (x31x) & (!n_n1592) & (!x42x)) + ((n_n4926) & (n_n4925) & (x31x) & (!n_n1592) & (x42x)) + ((n_n4926) & (n_n4925) & (x31x) & (n_n1592) & (!x42x)) + ((n_n4926) & (n_n4925) & (x31x) & (n_n1592) & (x42x)));
	assign n_n4058 = (((!n_n4909) & (!n_n4916) & (!x154x) & (x13204x)) + ((!n_n4909) & (!n_n4916) & (x154x) & (!x13204x)) + ((!n_n4909) & (!n_n4916) & (x154x) & (x13204x)) + ((!n_n4909) & (n_n4916) & (!x154x) & (!x13204x)) + ((!n_n4909) & (n_n4916) & (!x154x) & (x13204x)) + ((!n_n4909) & (n_n4916) & (x154x) & (!x13204x)) + ((!n_n4909) & (n_n4916) & (x154x) & (x13204x)) + ((n_n4909) & (!n_n4916) & (!x154x) & (!x13204x)) + ((n_n4909) & (!n_n4916) & (!x154x) & (x13204x)) + ((n_n4909) & (!n_n4916) & (x154x) & (!x13204x)) + ((n_n4909) & (!n_n4916) & (x154x) & (x13204x)) + ((n_n4909) & (n_n4916) & (!x154x) & (!x13204x)) + ((n_n4909) & (n_n4916) & (!x154x) & (x13204x)) + ((n_n4909) & (n_n4916) & (x154x) & (!x13204x)) + ((n_n4909) & (n_n4916) & (x154x) & (x13204x)));
	assign x13208x = (((!i_9_) & (!n_n528) & (!x531x) & (!n_n4936) & (x331x)) + ((!i_9_) & (!n_n528) & (!x531x) & (n_n4936) & (!x331x)) + ((!i_9_) & (!n_n528) & (!x531x) & (n_n4936) & (x331x)) + ((!i_9_) & (!n_n528) & (x531x) & (!n_n4936) & (x331x)) + ((!i_9_) & (!n_n528) & (x531x) & (n_n4936) & (!x331x)) + ((!i_9_) & (!n_n528) & (x531x) & (n_n4936) & (x331x)) + ((!i_9_) & (n_n528) & (!x531x) & (!n_n4936) & (x331x)) + ((!i_9_) & (n_n528) & (!x531x) & (n_n4936) & (!x331x)) + ((!i_9_) & (n_n528) & (!x531x) & (n_n4936) & (x331x)) + ((!i_9_) & (n_n528) & (x531x) & (!n_n4936) & (!x331x)) + ((!i_9_) & (n_n528) & (x531x) & (!n_n4936) & (x331x)) + ((!i_9_) & (n_n528) & (x531x) & (n_n4936) & (!x331x)) + ((!i_9_) & (n_n528) & (x531x) & (n_n4936) & (x331x)) + ((i_9_) & (!n_n528) & (!x531x) & (!n_n4936) & (x331x)) + ((i_9_) & (!n_n528) & (!x531x) & (n_n4936) & (!x331x)) + ((i_9_) & (!n_n528) & (!x531x) & (n_n4936) & (x331x)) + ((i_9_) & (!n_n528) & (x531x) & (!n_n4936) & (x331x)) + ((i_9_) & (!n_n528) & (x531x) & (n_n4936) & (!x331x)) + ((i_9_) & (!n_n528) & (x531x) & (n_n4936) & (x331x)) + ((i_9_) & (n_n528) & (!x531x) & (!n_n4936) & (x331x)) + ((i_9_) & (n_n528) & (!x531x) & (n_n4936) & (!x331x)) + ((i_9_) & (n_n528) & (!x531x) & (n_n4936) & (x331x)) + ((i_9_) & (n_n528) & (x531x) & (!n_n4936) & (x331x)) + ((i_9_) & (n_n528) & (x531x) & (n_n4936) & (!x331x)) + ((i_9_) & (n_n528) & (x531x) & (n_n4936) & (x331x)));
	assign x13209x = (((!n_n4934) & (!n_n4930) & (!n_n4935) & (!n_n4939) & (n_n4944)) + ((!n_n4934) & (!n_n4930) & (!n_n4935) & (n_n4939) & (!n_n4944)) + ((!n_n4934) & (!n_n4930) & (!n_n4935) & (n_n4939) & (n_n4944)) + ((!n_n4934) & (!n_n4930) & (n_n4935) & (!n_n4939) & (!n_n4944)) + ((!n_n4934) & (!n_n4930) & (n_n4935) & (!n_n4939) & (n_n4944)) + ((!n_n4934) & (!n_n4930) & (n_n4935) & (n_n4939) & (!n_n4944)) + ((!n_n4934) & (!n_n4930) & (n_n4935) & (n_n4939) & (n_n4944)) + ((!n_n4934) & (n_n4930) & (!n_n4935) & (!n_n4939) & (!n_n4944)) + ((!n_n4934) & (n_n4930) & (!n_n4935) & (!n_n4939) & (n_n4944)) + ((!n_n4934) & (n_n4930) & (!n_n4935) & (n_n4939) & (!n_n4944)) + ((!n_n4934) & (n_n4930) & (!n_n4935) & (n_n4939) & (n_n4944)) + ((!n_n4934) & (n_n4930) & (n_n4935) & (!n_n4939) & (!n_n4944)) + ((!n_n4934) & (n_n4930) & (n_n4935) & (!n_n4939) & (n_n4944)) + ((!n_n4934) & (n_n4930) & (n_n4935) & (n_n4939) & (!n_n4944)) + ((!n_n4934) & (n_n4930) & (n_n4935) & (n_n4939) & (n_n4944)) + ((n_n4934) & (!n_n4930) & (!n_n4935) & (!n_n4939) & (!n_n4944)) + ((n_n4934) & (!n_n4930) & (!n_n4935) & (!n_n4939) & (n_n4944)) + ((n_n4934) & (!n_n4930) & (!n_n4935) & (n_n4939) & (!n_n4944)) + ((n_n4934) & (!n_n4930) & (!n_n4935) & (n_n4939) & (n_n4944)) + ((n_n4934) & (!n_n4930) & (n_n4935) & (!n_n4939) & (!n_n4944)) + ((n_n4934) & (!n_n4930) & (n_n4935) & (!n_n4939) & (n_n4944)) + ((n_n4934) & (!n_n4930) & (n_n4935) & (n_n4939) & (!n_n4944)) + ((n_n4934) & (!n_n4930) & (n_n4935) & (n_n4939) & (n_n4944)) + ((n_n4934) & (n_n4930) & (!n_n4935) & (!n_n4939) & (!n_n4944)) + ((n_n4934) & (n_n4930) & (!n_n4935) & (!n_n4939) & (n_n4944)) + ((n_n4934) & (n_n4930) & (!n_n4935) & (n_n4939) & (!n_n4944)) + ((n_n4934) & (n_n4930) & (!n_n4935) & (n_n4939) & (n_n4944)) + ((n_n4934) & (n_n4930) & (n_n4935) & (!n_n4939) & (!n_n4944)) + ((n_n4934) & (n_n4930) & (n_n4935) & (!n_n4939) & (n_n4944)) + ((n_n4934) & (n_n4930) & (n_n4935) & (n_n4939) & (!n_n4944)) + ((n_n4934) & (n_n4930) & (n_n4935) & (n_n4939) & (n_n4944)));
	assign n_n4007 = (((!x13213x) & (!n_n4058) & (!x13208x) & (x13209x)) + ((!x13213x) & (!n_n4058) & (x13208x) & (!x13209x)) + ((!x13213x) & (!n_n4058) & (x13208x) & (x13209x)) + ((!x13213x) & (n_n4058) & (!x13208x) & (!x13209x)) + ((!x13213x) & (n_n4058) & (!x13208x) & (x13209x)) + ((!x13213x) & (n_n4058) & (x13208x) & (!x13209x)) + ((!x13213x) & (n_n4058) & (x13208x) & (x13209x)) + ((x13213x) & (!n_n4058) & (!x13208x) & (!x13209x)) + ((x13213x) & (!n_n4058) & (!x13208x) & (x13209x)) + ((x13213x) & (!n_n4058) & (x13208x) & (!x13209x)) + ((x13213x) & (!n_n4058) & (x13208x) & (x13209x)) + ((x13213x) & (n_n4058) & (!x13208x) & (!x13209x)) + ((x13213x) & (n_n4058) & (!x13208x) & (x13209x)) + ((x13213x) & (n_n4058) & (x13208x) & (!x13209x)) + ((x13213x) & (n_n4058) & (x13208x) & (x13209x)));
	assign x13226x = (((!x68x) & (!x210x) & (n_n814)) + ((!x68x) & (x210x) & (!n_n814)) + ((!x68x) & (x210x) & (n_n814)) + ((x68x) & (!x210x) & (!n_n814)) + ((x68x) & (!x210x) & (n_n814)) + ((x68x) & (x210x) & (!n_n814)) + ((x68x) & (x210x) & (n_n814)));
	assign x13227x = (((!n_n4952) & (!n_n4954) & (!x317x) & (x13224x)) + ((!n_n4952) & (!n_n4954) & (x317x) & (!x13224x)) + ((!n_n4952) & (!n_n4954) & (x317x) & (x13224x)) + ((!n_n4952) & (n_n4954) & (!x317x) & (!x13224x)) + ((!n_n4952) & (n_n4954) & (!x317x) & (x13224x)) + ((!n_n4952) & (n_n4954) & (x317x) & (!x13224x)) + ((!n_n4952) & (n_n4954) & (x317x) & (x13224x)) + ((n_n4952) & (!n_n4954) & (!x317x) & (!x13224x)) + ((n_n4952) & (!n_n4954) & (!x317x) & (x13224x)) + ((n_n4952) & (!n_n4954) & (x317x) & (!x13224x)) + ((n_n4952) & (!n_n4954) & (x317x) & (x13224x)) + ((n_n4952) & (n_n4954) & (!x317x) & (!x13224x)) + ((n_n4952) & (n_n4954) & (!x317x) & (x13224x)) + ((n_n4952) & (n_n4954) & (x317x) & (!x13224x)) + ((n_n4952) & (n_n4954) & (x317x) & (x13224x)));
	assign x13232x = (((!n_n509) & (!n_n260) & (!x20x) & (!n_n4876) & (x461x)) + ((!n_n509) & (!n_n260) & (!x20x) & (n_n4876) & (!x461x)) + ((!n_n509) & (!n_n260) & (!x20x) & (n_n4876) & (x461x)) + ((!n_n509) & (!n_n260) & (x20x) & (!n_n4876) & (x461x)) + ((!n_n509) & (!n_n260) & (x20x) & (n_n4876) & (!x461x)) + ((!n_n509) & (!n_n260) & (x20x) & (n_n4876) & (x461x)) + ((!n_n509) & (n_n260) & (!x20x) & (!n_n4876) & (x461x)) + ((!n_n509) & (n_n260) & (!x20x) & (n_n4876) & (!x461x)) + ((!n_n509) & (n_n260) & (!x20x) & (n_n4876) & (x461x)) + ((!n_n509) & (n_n260) & (x20x) & (!n_n4876) & (x461x)) + ((!n_n509) & (n_n260) & (x20x) & (n_n4876) & (!x461x)) + ((!n_n509) & (n_n260) & (x20x) & (n_n4876) & (x461x)) + ((n_n509) & (!n_n260) & (!x20x) & (!n_n4876) & (x461x)) + ((n_n509) & (!n_n260) & (!x20x) & (n_n4876) & (!x461x)) + ((n_n509) & (!n_n260) & (!x20x) & (n_n4876) & (x461x)) + ((n_n509) & (!n_n260) & (x20x) & (!n_n4876) & (x461x)) + ((n_n509) & (!n_n260) & (x20x) & (n_n4876) & (!x461x)) + ((n_n509) & (!n_n260) & (x20x) & (n_n4876) & (x461x)) + ((n_n509) & (n_n260) & (!x20x) & (!n_n4876) & (x461x)) + ((n_n509) & (n_n260) & (!x20x) & (n_n4876) & (!x461x)) + ((n_n509) & (n_n260) & (!x20x) & (n_n4876) & (x461x)) + ((n_n509) & (n_n260) & (x20x) & (!n_n4876) & (!x461x)) + ((n_n509) & (n_n260) & (x20x) & (!n_n4876) & (x461x)) + ((n_n509) & (n_n260) & (x20x) & (n_n4876) & (!x461x)) + ((n_n509) & (n_n260) & (x20x) & (n_n4876) & (x461x)));
	assign x22128x = (((!x295x) & (!x174x) & (!n_n4172) & (!n_n1970) & (!x137x)));
	assign x13235x = (((!x13226x) & (!x13227x) & (!x13232x) & (!x22128x)) + ((!x13226x) & (!x13227x) & (x13232x) & (!x22128x)) + ((!x13226x) & (!x13227x) & (x13232x) & (x22128x)) + ((!x13226x) & (x13227x) & (!x13232x) & (!x22128x)) + ((!x13226x) & (x13227x) & (!x13232x) & (x22128x)) + ((!x13226x) & (x13227x) & (x13232x) & (!x22128x)) + ((!x13226x) & (x13227x) & (x13232x) & (x22128x)) + ((x13226x) & (!x13227x) & (!x13232x) & (!x22128x)) + ((x13226x) & (!x13227x) & (!x13232x) & (x22128x)) + ((x13226x) & (!x13227x) & (x13232x) & (!x22128x)) + ((x13226x) & (!x13227x) & (x13232x) & (x22128x)) + ((x13226x) & (x13227x) & (!x13232x) & (!x22128x)) + ((x13226x) & (x13227x) & (!x13232x) & (x22128x)) + ((x13226x) & (x13227x) & (x13232x) & (!x22128x)) + ((x13226x) & (x13227x) & (x13232x) & (x22128x)));
	assign x13234x = (((!n_n4898) & (!n_n4895) & (!n_n4060) & (!x13199x) & (x49x)) + ((!n_n4898) & (!n_n4895) & (!n_n4060) & (x13199x) & (!x49x)) + ((!n_n4898) & (!n_n4895) & (!n_n4060) & (x13199x) & (x49x)) + ((!n_n4898) & (!n_n4895) & (n_n4060) & (!x13199x) & (!x49x)) + ((!n_n4898) & (!n_n4895) & (n_n4060) & (!x13199x) & (x49x)) + ((!n_n4898) & (!n_n4895) & (n_n4060) & (x13199x) & (!x49x)) + ((!n_n4898) & (!n_n4895) & (n_n4060) & (x13199x) & (x49x)) + ((!n_n4898) & (n_n4895) & (!n_n4060) & (!x13199x) & (!x49x)) + ((!n_n4898) & (n_n4895) & (!n_n4060) & (!x13199x) & (x49x)) + ((!n_n4898) & (n_n4895) & (!n_n4060) & (x13199x) & (!x49x)) + ((!n_n4898) & (n_n4895) & (!n_n4060) & (x13199x) & (x49x)) + ((!n_n4898) & (n_n4895) & (n_n4060) & (!x13199x) & (!x49x)) + ((!n_n4898) & (n_n4895) & (n_n4060) & (!x13199x) & (x49x)) + ((!n_n4898) & (n_n4895) & (n_n4060) & (x13199x) & (!x49x)) + ((!n_n4898) & (n_n4895) & (n_n4060) & (x13199x) & (x49x)) + ((n_n4898) & (!n_n4895) & (!n_n4060) & (!x13199x) & (!x49x)) + ((n_n4898) & (!n_n4895) & (!n_n4060) & (!x13199x) & (x49x)) + ((n_n4898) & (!n_n4895) & (!n_n4060) & (x13199x) & (!x49x)) + ((n_n4898) & (!n_n4895) & (!n_n4060) & (x13199x) & (x49x)) + ((n_n4898) & (!n_n4895) & (n_n4060) & (!x13199x) & (!x49x)) + ((n_n4898) & (!n_n4895) & (n_n4060) & (!x13199x) & (x49x)) + ((n_n4898) & (!n_n4895) & (n_n4060) & (x13199x) & (!x49x)) + ((n_n4898) & (!n_n4895) & (n_n4060) & (x13199x) & (x49x)) + ((n_n4898) & (n_n4895) & (!n_n4060) & (!x13199x) & (!x49x)) + ((n_n4898) & (n_n4895) & (!n_n4060) & (!x13199x) & (x49x)) + ((n_n4898) & (n_n4895) & (!n_n4060) & (x13199x) & (!x49x)) + ((n_n4898) & (n_n4895) & (!n_n4060) & (x13199x) & (x49x)) + ((n_n4898) & (n_n4895) & (n_n4060) & (!x13199x) & (!x49x)) + ((n_n4898) & (n_n4895) & (n_n4060) & (!x13199x) & (x49x)) + ((n_n4898) & (n_n4895) & (n_n4060) & (x13199x) & (!x49x)) + ((n_n4898) & (n_n4895) & (n_n4060) & (x13199x) & (x49x)));
	assign x94x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n509) & (n_n325)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n509) & (n_n325)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n509) & (n_n325)) + ((i_9_) & (n_n524) & (n_n526) & (n_n509) & (n_n325)));
	assign x13237x = (((!i_9_) & (n_n528) & (n_n509) & (n_n325)) + ((i_9_) & (n_n528) & (n_n509) & (n_n325)));
	assign n_n4072 = (((!n_n4743) & (!x374x) & (!x73x) & (!x94x) & (x13237x)) + ((!n_n4743) & (!x374x) & (!x73x) & (x94x) & (!x13237x)) + ((!n_n4743) & (!x374x) & (!x73x) & (x94x) & (x13237x)) + ((!n_n4743) & (!x374x) & (x73x) & (!x94x) & (!x13237x)) + ((!n_n4743) & (!x374x) & (x73x) & (!x94x) & (x13237x)) + ((!n_n4743) & (!x374x) & (x73x) & (x94x) & (!x13237x)) + ((!n_n4743) & (!x374x) & (x73x) & (x94x) & (x13237x)) + ((!n_n4743) & (x374x) & (!x73x) & (!x94x) & (!x13237x)) + ((!n_n4743) & (x374x) & (!x73x) & (!x94x) & (x13237x)) + ((!n_n4743) & (x374x) & (!x73x) & (x94x) & (!x13237x)) + ((!n_n4743) & (x374x) & (!x73x) & (x94x) & (x13237x)) + ((!n_n4743) & (x374x) & (x73x) & (!x94x) & (!x13237x)) + ((!n_n4743) & (x374x) & (x73x) & (!x94x) & (x13237x)) + ((!n_n4743) & (x374x) & (x73x) & (x94x) & (!x13237x)) + ((!n_n4743) & (x374x) & (x73x) & (x94x) & (x13237x)) + ((n_n4743) & (!x374x) & (!x73x) & (!x94x) & (!x13237x)) + ((n_n4743) & (!x374x) & (!x73x) & (!x94x) & (x13237x)) + ((n_n4743) & (!x374x) & (!x73x) & (x94x) & (!x13237x)) + ((n_n4743) & (!x374x) & (!x73x) & (x94x) & (x13237x)) + ((n_n4743) & (!x374x) & (x73x) & (!x94x) & (!x13237x)) + ((n_n4743) & (!x374x) & (x73x) & (!x94x) & (x13237x)) + ((n_n4743) & (!x374x) & (x73x) & (x94x) & (!x13237x)) + ((n_n4743) & (!x374x) & (x73x) & (x94x) & (x13237x)) + ((n_n4743) & (x374x) & (!x73x) & (!x94x) & (!x13237x)) + ((n_n4743) & (x374x) & (!x73x) & (!x94x) & (x13237x)) + ((n_n4743) & (x374x) & (!x73x) & (x94x) & (!x13237x)) + ((n_n4743) & (x374x) & (!x73x) & (x94x) & (x13237x)) + ((n_n4743) & (x374x) & (x73x) & (!x94x) & (!x13237x)) + ((n_n4743) & (x374x) & (x73x) & (!x94x) & (x13237x)) + ((n_n4743) & (x374x) & (x73x) & (x94x) & (!x13237x)) + ((n_n4743) & (x374x) & (x73x) & (x94x) & (x13237x)));
	assign n_n4210 = (((!x21x) & (!n_n325) & (!x20x) & (!n_n500) & (n_n4756)) + ((!x21x) & (!n_n325) & (!x20x) & (n_n500) & (n_n4756)) + ((!x21x) & (!n_n325) & (x20x) & (!n_n500) & (n_n4756)) + ((!x21x) & (!n_n325) & (x20x) & (n_n500) & (n_n4756)) + ((!x21x) & (n_n325) & (!x20x) & (!n_n500) & (n_n4756)) + ((!x21x) & (n_n325) & (!x20x) & (n_n500) & (n_n4756)) + ((!x21x) & (n_n325) & (x20x) & (!n_n500) & (n_n4756)) + ((!x21x) & (n_n325) & (x20x) & (n_n500) & (!n_n4756)) + ((!x21x) & (n_n325) & (x20x) & (n_n500) & (n_n4756)) + ((x21x) & (!n_n325) & (!x20x) & (!n_n500) & (n_n4756)) + ((x21x) & (!n_n325) & (!x20x) & (n_n500) & (n_n4756)) + ((x21x) & (!n_n325) & (x20x) & (!n_n500) & (n_n4756)) + ((x21x) & (!n_n325) & (x20x) & (n_n500) & (n_n4756)) + ((x21x) & (n_n325) & (!x20x) & (!n_n500) & (n_n4756)) + ((x21x) & (n_n325) & (!x20x) & (n_n500) & (!n_n4756)) + ((x21x) & (n_n325) & (!x20x) & (n_n500) & (n_n4756)) + ((x21x) & (n_n325) & (x20x) & (!n_n500) & (n_n4756)) + ((x21x) & (n_n325) & (x20x) & (n_n500) & (!n_n4756)) + ((x21x) & (n_n325) & (x20x) & (n_n500) & (n_n4756)));
	assign n_n1087 = (((!n_n4759) & (!x69x) & (!n_n4763) & (!n_n4210) & (x370x)) + ((!n_n4759) & (!x69x) & (!n_n4763) & (n_n4210) & (!x370x)) + ((!n_n4759) & (!x69x) & (!n_n4763) & (n_n4210) & (x370x)) + ((!n_n4759) & (!x69x) & (n_n4763) & (!n_n4210) & (!x370x)) + ((!n_n4759) & (!x69x) & (n_n4763) & (!n_n4210) & (x370x)) + ((!n_n4759) & (!x69x) & (n_n4763) & (n_n4210) & (!x370x)) + ((!n_n4759) & (!x69x) & (n_n4763) & (n_n4210) & (x370x)) + ((!n_n4759) & (x69x) & (!n_n4763) & (!n_n4210) & (!x370x)) + ((!n_n4759) & (x69x) & (!n_n4763) & (!n_n4210) & (x370x)) + ((!n_n4759) & (x69x) & (!n_n4763) & (n_n4210) & (!x370x)) + ((!n_n4759) & (x69x) & (!n_n4763) & (n_n4210) & (x370x)) + ((!n_n4759) & (x69x) & (n_n4763) & (!n_n4210) & (!x370x)) + ((!n_n4759) & (x69x) & (n_n4763) & (!n_n4210) & (x370x)) + ((!n_n4759) & (x69x) & (n_n4763) & (n_n4210) & (!x370x)) + ((!n_n4759) & (x69x) & (n_n4763) & (n_n4210) & (x370x)) + ((n_n4759) & (!x69x) & (!n_n4763) & (!n_n4210) & (!x370x)) + ((n_n4759) & (!x69x) & (!n_n4763) & (!n_n4210) & (x370x)) + ((n_n4759) & (!x69x) & (!n_n4763) & (n_n4210) & (!x370x)) + ((n_n4759) & (!x69x) & (!n_n4763) & (n_n4210) & (x370x)) + ((n_n4759) & (!x69x) & (n_n4763) & (!n_n4210) & (!x370x)) + ((n_n4759) & (!x69x) & (n_n4763) & (!n_n4210) & (x370x)) + ((n_n4759) & (!x69x) & (n_n4763) & (n_n4210) & (!x370x)) + ((n_n4759) & (!x69x) & (n_n4763) & (n_n4210) & (x370x)) + ((n_n4759) & (x69x) & (!n_n4763) & (!n_n4210) & (!x370x)) + ((n_n4759) & (x69x) & (!n_n4763) & (!n_n4210) & (x370x)) + ((n_n4759) & (x69x) & (!n_n4763) & (n_n4210) & (!x370x)) + ((n_n4759) & (x69x) & (!n_n4763) & (n_n4210) & (x370x)) + ((n_n4759) & (x69x) & (n_n4763) & (!n_n4210) & (!x370x)) + ((n_n4759) & (x69x) & (n_n4763) & (!n_n4210) & (x370x)) + ((n_n4759) & (x69x) & (n_n4763) & (n_n4210) & (!x370x)) + ((n_n4759) & (x69x) & (n_n4763) & (n_n4210) & (x370x)));
	assign x13244x = (((!x25x) & (!n_n325) & (!n_n535) & (!n_n4695) & (x221x)) + ((!x25x) & (!n_n325) & (!n_n535) & (n_n4695) & (!x221x)) + ((!x25x) & (!n_n325) & (!n_n535) & (n_n4695) & (x221x)) + ((!x25x) & (!n_n325) & (n_n535) & (!n_n4695) & (x221x)) + ((!x25x) & (!n_n325) & (n_n535) & (n_n4695) & (!x221x)) + ((!x25x) & (!n_n325) & (n_n535) & (n_n4695) & (x221x)) + ((!x25x) & (n_n325) & (!n_n535) & (!n_n4695) & (x221x)) + ((!x25x) & (n_n325) & (!n_n535) & (n_n4695) & (!x221x)) + ((!x25x) & (n_n325) & (!n_n535) & (n_n4695) & (x221x)) + ((!x25x) & (n_n325) & (n_n535) & (!n_n4695) & (x221x)) + ((!x25x) & (n_n325) & (n_n535) & (n_n4695) & (!x221x)) + ((!x25x) & (n_n325) & (n_n535) & (n_n4695) & (x221x)) + ((x25x) & (!n_n325) & (!n_n535) & (!n_n4695) & (x221x)) + ((x25x) & (!n_n325) & (!n_n535) & (n_n4695) & (!x221x)) + ((x25x) & (!n_n325) & (!n_n535) & (n_n4695) & (x221x)) + ((x25x) & (!n_n325) & (n_n535) & (!n_n4695) & (x221x)) + ((x25x) & (!n_n325) & (n_n535) & (n_n4695) & (!x221x)) + ((x25x) & (!n_n325) & (n_n535) & (n_n4695) & (x221x)) + ((x25x) & (n_n325) & (!n_n535) & (!n_n4695) & (x221x)) + ((x25x) & (n_n325) & (!n_n535) & (n_n4695) & (!x221x)) + ((x25x) & (n_n325) & (!n_n535) & (n_n4695) & (x221x)) + ((x25x) & (n_n325) & (n_n535) & (!n_n4695) & (!x221x)) + ((x25x) & (n_n325) & (n_n535) & (!n_n4695) & (x221x)) + ((x25x) & (n_n325) & (n_n535) & (n_n4695) & (!x221x)) + ((x25x) & (n_n325) & (n_n535) & (n_n4695) & (x221x)));
	assign x13245x = (((!x10x) & (!n_n520) & (!n_n464) & (!n_n4700) & (n_n4219)) + ((!x10x) & (!n_n520) & (!n_n464) & (n_n4700) & (!n_n4219)) + ((!x10x) & (!n_n520) & (!n_n464) & (n_n4700) & (n_n4219)) + ((!x10x) & (!n_n520) & (n_n464) & (!n_n4700) & (n_n4219)) + ((!x10x) & (!n_n520) & (n_n464) & (n_n4700) & (!n_n4219)) + ((!x10x) & (!n_n520) & (n_n464) & (n_n4700) & (n_n4219)) + ((!x10x) & (n_n520) & (!n_n464) & (!n_n4700) & (n_n4219)) + ((!x10x) & (n_n520) & (!n_n464) & (n_n4700) & (!n_n4219)) + ((!x10x) & (n_n520) & (!n_n464) & (n_n4700) & (n_n4219)) + ((!x10x) & (n_n520) & (n_n464) & (!n_n4700) & (n_n4219)) + ((!x10x) & (n_n520) & (n_n464) & (n_n4700) & (!n_n4219)) + ((!x10x) & (n_n520) & (n_n464) & (n_n4700) & (n_n4219)) + ((x10x) & (!n_n520) & (!n_n464) & (!n_n4700) & (n_n4219)) + ((x10x) & (!n_n520) & (!n_n464) & (n_n4700) & (!n_n4219)) + ((x10x) & (!n_n520) & (!n_n464) & (n_n4700) & (n_n4219)) + ((x10x) & (!n_n520) & (n_n464) & (!n_n4700) & (n_n4219)) + ((x10x) & (!n_n520) & (n_n464) & (n_n4700) & (!n_n4219)) + ((x10x) & (!n_n520) & (n_n464) & (n_n4700) & (n_n4219)) + ((x10x) & (n_n520) & (!n_n464) & (!n_n4700) & (n_n4219)) + ((x10x) & (n_n520) & (!n_n464) & (n_n4700) & (!n_n4219)) + ((x10x) & (n_n520) & (!n_n464) & (n_n4700) & (n_n4219)) + ((x10x) & (n_n520) & (n_n464) & (!n_n4700) & (!n_n4219)) + ((x10x) & (n_n520) & (n_n464) & (!n_n4700) & (n_n4219)) + ((x10x) & (n_n520) & (n_n464) & (n_n4700) & (!n_n4219)) + ((x10x) & (n_n520) & (n_n464) & (n_n4700) & (n_n4219)));
	assign x13251x = (((!n_n4708) & (!n_n4716) & (!n_n4723) & (n_n4713)) + ((!n_n4708) & (!n_n4716) & (n_n4723) & (!n_n4713)) + ((!n_n4708) & (!n_n4716) & (n_n4723) & (n_n4713)) + ((!n_n4708) & (n_n4716) & (!n_n4723) & (!n_n4713)) + ((!n_n4708) & (n_n4716) & (!n_n4723) & (n_n4713)) + ((!n_n4708) & (n_n4716) & (n_n4723) & (!n_n4713)) + ((!n_n4708) & (n_n4716) & (n_n4723) & (n_n4713)) + ((n_n4708) & (!n_n4716) & (!n_n4723) & (!n_n4713)) + ((n_n4708) & (!n_n4716) & (!n_n4723) & (n_n4713)) + ((n_n4708) & (!n_n4716) & (n_n4723) & (!n_n4713)) + ((n_n4708) & (!n_n4716) & (n_n4723) & (n_n4713)) + ((n_n4708) & (n_n4716) & (!n_n4723) & (!n_n4713)) + ((n_n4708) & (n_n4716) & (!n_n4723) & (n_n4713)) + ((n_n4708) & (n_n4716) & (n_n4723) & (!n_n4713)) + ((n_n4708) & (n_n4716) & (n_n4723) & (n_n4713)));
	assign x13252x = (((!n_n4720) & (!x241x) & (!n_n4727) & (!n_n4726) & (n_n4728)) + ((!n_n4720) & (!x241x) & (!n_n4727) & (n_n4726) & (!n_n4728)) + ((!n_n4720) & (!x241x) & (!n_n4727) & (n_n4726) & (n_n4728)) + ((!n_n4720) & (!x241x) & (n_n4727) & (!n_n4726) & (!n_n4728)) + ((!n_n4720) & (!x241x) & (n_n4727) & (!n_n4726) & (n_n4728)) + ((!n_n4720) & (!x241x) & (n_n4727) & (n_n4726) & (!n_n4728)) + ((!n_n4720) & (!x241x) & (n_n4727) & (n_n4726) & (n_n4728)) + ((!n_n4720) & (x241x) & (!n_n4727) & (!n_n4726) & (!n_n4728)) + ((!n_n4720) & (x241x) & (!n_n4727) & (!n_n4726) & (n_n4728)) + ((!n_n4720) & (x241x) & (!n_n4727) & (n_n4726) & (!n_n4728)) + ((!n_n4720) & (x241x) & (!n_n4727) & (n_n4726) & (n_n4728)) + ((!n_n4720) & (x241x) & (n_n4727) & (!n_n4726) & (!n_n4728)) + ((!n_n4720) & (x241x) & (n_n4727) & (!n_n4726) & (n_n4728)) + ((!n_n4720) & (x241x) & (n_n4727) & (n_n4726) & (!n_n4728)) + ((!n_n4720) & (x241x) & (n_n4727) & (n_n4726) & (n_n4728)) + ((n_n4720) & (!x241x) & (!n_n4727) & (!n_n4726) & (!n_n4728)) + ((n_n4720) & (!x241x) & (!n_n4727) & (!n_n4726) & (n_n4728)) + ((n_n4720) & (!x241x) & (!n_n4727) & (n_n4726) & (!n_n4728)) + ((n_n4720) & (!x241x) & (!n_n4727) & (n_n4726) & (n_n4728)) + ((n_n4720) & (!x241x) & (n_n4727) & (!n_n4726) & (!n_n4728)) + ((n_n4720) & (!x241x) & (n_n4727) & (!n_n4726) & (n_n4728)) + ((n_n4720) & (!x241x) & (n_n4727) & (n_n4726) & (!n_n4728)) + ((n_n4720) & (!x241x) & (n_n4727) & (n_n4726) & (n_n4728)) + ((n_n4720) & (x241x) & (!n_n4727) & (!n_n4726) & (!n_n4728)) + ((n_n4720) & (x241x) & (!n_n4727) & (!n_n4726) & (n_n4728)) + ((n_n4720) & (x241x) & (!n_n4727) & (n_n4726) & (!n_n4728)) + ((n_n4720) & (x241x) & (!n_n4727) & (n_n4726) & (n_n4728)) + ((n_n4720) & (x241x) & (n_n4727) & (!n_n4726) & (!n_n4728)) + ((n_n4720) & (x241x) & (n_n4727) & (!n_n4726) & (n_n4728)) + ((n_n4720) & (x241x) & (n_n4727) & (n_n4726) & (!n_n4728)) + ((n_n4720) & (x241x) & (n_n4727) & (n_n4726) & (n_n4728)));
	assign x13253x = (((!x39x) & (!n_n4715) & (!n_n4714) & (!x367x) & (x30x)) + ((!x39x) & (!n_n4715) & (!n_n4714) & (x367x) & (!x30x)) + ((!x39x) & (!n_n4715) & (!n_n4714) & (x367x) & (x30x)) + ((!x39x) & (!n_n4715) & (n_n4714) & (!x367x) & (!x30x)) + ((!x39x) & (!n_n4715) & (n_n4714) & (!x367x) & (x30x)) + ((!x39x) & (!n_n4715) & (n_n4714) & (x367x) & (!x30x)) + ((!x39x) & (!n_n4715) & (n_n4714) & (x367x) & (x30x)) + ((!x39x) & (n_n4715) & (!n_n4714) & (!x367x) & (!x30x)) + ((!x39x) & (n_n4715) & (!n_n4714) & (!x367x) & (x30x)) + ((!x39x) & (n_n4715) & (!n_n4714) & (x367x) & (!x30x)) + ((!x39x) & (n_n4715) & (!n_n4714) & (x367x) & (x30x)) + ((!x39x) & (n_n4715) & (n_n4714) & (!x367x) & (!x30x)) + ((!x39x) & (n_n4715) & (n_n4714) & (!x367x) & (x30x)) + ((!x39x) & (n_n4715) & (n_n4714) & (x367x) & (!x30x)) + ((!x39x) & (n_n4715) & (n_n4714) & (x367x) & (x30x)) + ((x39x) & (!n_n4715) & (!n_n4714) & (!x367x) & (!x30x)) + ((x39x) & (!n_n4715) & (!n_n4714) & (!x367x) & (x30x)) + ((x39x) & (!n_n4715) & (!n_n4714) & (x367x) & (!x30x)) + ((x39x) & (!n_n4715) & (!n_n4714) & (x367x) & (x30x)) + ((x39x) & (!n_n4715) & (n_n4714) & (!x367x) & (!x30x)) + ((x39x) & (!n_n4715) & (n_n4714) & (!x367x) & (x30x)) + ((x39x) & (!n_n4715) & (n_n4714) & (x367x) & (!x30x)) + ((x39x) & (!n_n4715) & (n_n4714) & (x367x) & (x30x)) + ((x39x) & (n_n4715) & (!n_n4714) & (!x367x) & (!x30x)) + ((x39x) & (n_n4715) & (!n_n4714) & (!x367x) & (x30x)) + ((x39x) & (n_n4715) & (!n_n4714) & (x367x) & (!x30x)) + ((x39x) & (n_n4715) & (!n_n4714) & (x367x) & (x30x)) + ((x39x) & (n_n4715) & (n_n4714) & (!x367x) & (!x30x)) + ((x39x) & (n_n4715) & (n_n4714) & (!x367x) & (x30x)) + ((x39x) & (n_n4715) & (n_n4714) & (x367x) & (!x30x)) + ((x39x) & (n_n4715) & (n_n4714) & (x367x) & (x30x)));
	assign n_n4013 = (((!x13244x) & (!x13245x) & (!x13251x) & (!x13252x) & (x13253x)) + ((!x13244x) & (!x13245x) & (!x13251x) & (x13252x) & (!x13253x)) + ((!x13244x) & (!x13245x) & (!x13251x) & (x13252x) & (x13253x)) + ((!x13244x) & (!x13245x) & (x13251x) & (!x13252x) & (!x13253x)) + ((!x13244x) & (!x13245x) & (x13251x) & (!x13252x) & (x13253x)) + ((!x13244x) & (!x13245x) & (x13251x) & (x13252x) & (!x13253x)) + ((!x13244x) & (!x13245x) & (x13251x) & (x13252x) & (x13253x)) + ((!x13244x) & (x13245x) & (!x13251x) & (!x13252x) & (!x13253x)) + ((!x13244x) & (x13245x) & (!x13251x) & (!x13252x) & (x13253x)) + ((!x13244x) & (x13245x) & (!x13251x) & (x13252x) & (!x13253x)) + ((!x13244x) & (x13245x) & (!x13251x) & (x13252x) & (x13253x)) + ((!x13244x) & (x13245x) & (x13251x) & (!x13252x) & (!x13253x)) + ((!x13244x) & (x13245x) & (x13251x) & (!x13252x) & (x13253x)) + ((!x13244x) & (x13245x) & (x13251x) & (x13252x) & (!x13253x)) + ((!x13244x) & (x13245x) & (x13251x) & (x13252x) & (x13253x)) + ((x13244x) & (!x13245x) & (!x13251x) & (!x13252x) & (!x13253x)) + ((x13244x) & (!x13245x) & (!x13251x) & (!x13252x) & (x13253x)) + ((x13244x) & (!x13245x) & (!x13251x) & (x13252x) & (!x13253x)) + ((x13244x) & (!x13245x) & (!x13251x) & (x13252x) & (x13253x)) + ((x13244x) & (!x13245x) & (x13251x) & (!x13252x) & (!x13253x)) + ((x13244x) & (!x13245x) & (x13251x) & (!x13252x) & (x13253x)) + ((x13244x) & (!x13245x) & (x13251x) & (x13252x) & (!x13253x)) + ((x13244x) & (!x13245x) & (x13251x) & (x13252x) & (x13253x)) + ((x13244x) & (x13245x) & (!x13251x) & (!x13252x) & (!x13253x)) + ((x13244x) & (x13245x) & (!x13251x) & (!x13252x) & (x13253x)) + ((x13244x) & (x13245x) & (!x13251x) & (x13252x) & (!x13253x)) + ((x13244x) & (x13245x) & (!x13251x) & (x13252x) & (x13253x)) + ((x13244x) & (x13245x) & (x13251x) & (!x13252x) & (!x13253x)) + ((x13244x) & (x13245x) & (x13251x) & (!x13252x) & (x13253x)) + ((x13244x) & (x13245x) & (x13251x) & (x13252x) & (!x13253x)) + ((x13244x) & (x13245x) & (x13251x) & (x13252x) & (x13253x)));
	assign n_n4691 = (((!i_9_) & (n_n524) & (n_n390) & (n_n464)));
	assign n_n4693 = (((!i_1_) & (i_2_) & (i_0_) & (x20x) & (n_n464)));
	assign x22220x = (((!x10x) & (!x516x) & (!x81x) & (!x426x) & (!n_n4688)) + ((!x10x) & (x516x) & (!x81x) & (!x426x) & (!n_n4688)) + ((x10x) & (!x516x) & (!x81x) & (!x426x) & (!n_n4688)));
	assign x13269x = (((!n_n4685) & (!n_n4691) & (!n_n4687) & (!n_n4693) & (!x22220x)) + ((!n_n4685) & (!n_n4691) & (!n_n4687) & (n_n4693) & (!x22220x)) + ((!n_n4685) & (!n_n4691) & (!n_n4687) & (n_n4693) & (x22220x)) + ((!n_n4685) & (!n_n4691) & (n_n4687) & (!n_n4693) & (!x22220x)) + ((!n_n4685) & (!n_n4691) & (n_n4687) & (!n_n4693) & (x22220x)) + ((!n_n4685) & (!n_n4691) & (n_n4687) & (n_n4693) & (!x22220x)) + ((!n_n4685) & (!n_n4691) & (n_n4687) & (n_n4693) & (x22220x)) + ((!n_n4685) & (n_n4691) & (!n_n4687) & (!n_n4693) & (!x22220x)) + ((!n_n4685) & (n_n4691) & (!n_n4687) & (!n_n4693) & (x22220x)) + ((!n_n4685) & (n_n4691) & (!n_n4687) & (n_n4693) & (!x22220x)) + ((!n_n4685) & (n_n4691) & (!n_n4687) & (n_n4693) & (x22220x)) + ((!n_n4685) & (n_n4691) & (n_n4687) & (!n_n4693) & (!x22220x)) + ((!n_n4685) & (n_n4691) & (n_n4687) & (!n_n4693) & (x22220x)) + ((!n_n4685) & (n_n4691) & (n_n4687) & (n_n4693) & (!x22220x)) + ((!n_n4685) & (n_n4691) & (n_n4687) & (n_n4693) & (x22220x)) + ((n_n4685) & (!n_n4691) & (!n_n4687) & (!n_n4693) & (!x22220x)) + ((n_n4685) & (!n_n4691) & (!n_n4687) & (!n_n4693) & (x22220x)) + ((n_n4685) & (!n_n4691) & (!n_n4687) & (n_n4693) & (!x22220x)) + ((n_n4685) & (!n_n4691) & (!n_n4687) & (n_n4693) & (x22220x)) + ((n_n4685) & (!n_n4691) & (n_n4687) & (!n_n4693) & (!x22220x)) + ((n_n4685) & (!n_n4691) & (n_n4687) & (!n_n4693) & (x22220x)) + ((n_n4685) & (!n_n4691) & (n_n4687) & (n_n4693) & (!x22220x)) + ((n_n4685) & (!n_n4691) & (n_n4687) & (n_n4693) & (x22220x)) + ((n_n4685) & (n_n4691) & (!n_n4687) & (!n_n4693) & (!x22220x)) + ((n_n4685) & (n_n4691) & (!n_n4687) & (!n_n4693) & (x22220x)) + ((n_n4685) & (n_n4691) & (!n_n4687) & (n_n4693) & (!x22220x)) + ((n_n4685) & (n_n4691) & (!n_n4687) & (n_n4693) & (x22220x)) + ((n_n4685) & (n_n4691) & (n_n4687) & (!n_n4693) & (!x22220x)) + ((n_n4685) & (n_n4691) & (n_n4687) & (!n_n4693) & (x22220x)) + ((n_n4685) & (n_n4691) & (n_n4687) & (n_n4693) & (!x22220x)) + ((n_n4685) & (n_n4691) & (n_n4687) & (n_n4693) & (x22220x)));
	assign n_n4078 = (((!n_n4659) & (!n_n4661) & (!n_n4657) & (!x312x) & (!x22126x)) + ((!n_n4659) & (!n_n4661) & (!n_n4657) & (x312x) & (!x22126x)) + ((!n_n4659) & (!n_n4661) & (!n_n4657) & (x312x) & (x22126x)) + ((!n_n4659) & (!n_n4661) & (n_n4657) & (!x312x) & (!x22126x)) + ((!n_n4659) & (!n_n4661) & (n_n4657) & (!x312x) & (x22126x)) + ((!n_n4659) & (!n_n4661) & (n_n4657) & (x312x) & (!x22126x)) + ((!n_n4659) & (!n_n4661) & (n_n4657) & (x312x) & (x22126x)) + ((!n_n4659) & (n_n4661) & (!n_n4657) & (!x312x) & (!x22126x)) + ((!n_n4659) & (n_n4661) & (!n_n4657) & (!x312x) & (x22126x)) + ((!n_n4659) & (n_n4661) & (!n_n4657) & (x312x) & (!x22126x)) + ((!n_n4659) & (n_n4661) & (!n_n4657) & (x312x) & (x22126x)) + ((!n_n4659) & (n_n4661) & (n_n4657) & (!x312x) & (!x22126x)) + ((!n_n4659) & (n_n4661) & (n_n4657) & (!x312x) & (x22126x)) + ((!n_n4659) & (n_n4661) & (n_n4657) & (x312x) & (!x22126x)) + ((!n_n4659) & (n_n4661) & (n_n4657) & (x312x) & (x22126x)) + ((n_n4659) & (!n_n4661) & (!n_n4657) & (!x312x) & (!x22126x)) + ((n_n4659) & (!n_n4661) & (!n_n4657) & (!x312x) & (x22126x)) + ((n_n4659) & (!n_n4661) & (!n_n4657) & (x312x) & (!x22126x)) + ((n_n4659) & (!n_n4661) & (!n_n4657) & (x312x) & (x22126x)) + ((n_n4659) & (!n_n4661) & (n_n4657) & (!x312x) & (!x22126x)) + ((n_n4659) & (!n_n4661) & (n_n4657) & (!x312x) & (x22126x)) + ((n_n4659) & (!n_n4661) & (n_n4657) & (x312x) & (!x22126x)) + ((n_n4659) & (!n_n4661) & (n_n4657) & (x312x) & (x22126x)) + ((n_n4659) & (n_n4661) & (!n_n4657) & (!x312x) & (!x22126x)) + ((n_n4659) & (n_n4661) & (!n_n4657) & (!x312x) & (x22126x)) + ((n_n4659) & (n_n4661) & (!n_n4657) & (x312x) & (!x22126x)) + ((n_n4659) & (n_n4661) & (!n_n4657) & (x312x) & (x22126x)) + ((n_n4659) & (n_n4661) & (n_n4657) & (!x312x) & (!x22126x)) + ((n_n4659) & (n_n4661) & (n_n4657) & (!x312x) & (x22126x)) + ((n_n4659) & (n_n4661) & (n_n4657) & (x312x) & (!x22126x)) + ((n_n4659) & (n_n4661) & (n_n4657) & (x312x) & (x22126x)));
	assign x157x = (((!i_9_) & (n_n390) & (n_n473) & (n_n530)) + ((i_9_) & (n_n390) & (n_n473) & (n_n530)));
	assign x339x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n390) & (n_n473)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n390) & (n_n473)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n390) & (n_n473)) + ((i_9_) & (n_n524) & (n_n526) & (n_n390) & (n_n473)));
	assign x13264x = (((!n_n4670) & (!n_n4671) & (!n_n4680) & (x80x)) + ((!n_n4670) & (!n_n4671) & (n_n4680) & (!x80x)) + ((!n_n4670) & (!n_n4671) & (n_n4680) & (x80x)) + ((!n_n4670) & (n_n4671) & (!n_n4680) & (!x80x)) + ((!n_n4670) & (n_n4671) & (!n_n4680) & (x80x)) + ((!n_n4670) & (n_n4671) & (n_n4680) & (!x80x)) + ((!n_n4670) & (n_n4671) & (n_n4680) & (x80x)) + ((n_n4670) & (!n_n4671) & (!n_n4680) & (!x80x)) + ((n_n4670) & (!n_n4671) & (!n_n4680) & (x80x)) + ((n_n4670) & (!n_n4671) & (n_n4680) & (!x80x)) + ((n_n4670) & (!n_n4671) & (n_n4680) & (x80x)) + ((n_n4670) & (n_n4671) & (!n_n4680) & (!x80x)) + ((n_n4670) & (n_n4671) & (!n_n4680) & (x80x)) + ((n_n4670) & (n_n4671) & (n_n4680) & (!x80x)) + ((n_n4670) & (n_n4671) & (n_n4680) & (x80x)));
	assign n_n4014 = (((!x13269x) & (!n_n4078) & (!x157x) & (!x339x) & (x13264x)) + ((!x13269x) & (!n_n4078) & (!x157x) & (x339x) & (!x13264x)) + ((!x13269x) & (!n_n4078) & (!x157x) & (x339x) & (x13264x)) + ((!x13269x) & (!n_n4078) & (x157x) & (!x339x) & (!x13264x)) + ((!x13269x) & (!n_n4078) & (x157x) & (!x339x) & (x13264x)) + ((!x13269x) & (!n_n4078) & (x157x) & (x339x) & (!x13264x)) + ((!x13269x) & (!n_n4078) & (x157x) & (x339x) & (x13264x)) + ((!x13269x) & (n_n4078) & (!x157x) & (!x339x) & (!x13264x)) + ((!x13269x) & (n_n4078) & (!x157x) & (!x339x) & (x13264x)) + ((!x13269x) & (n_n4078) & (!x157x) & (x339x) & (!x13264x)) + ((!x13269x) & (n_n4078) & (!x157x) & (x339x) & (x13264x)) + ((!x13269x) & (n_n4078) & (x157x) & (!x339x) & (!x13264x)) + ((!x13269x) & (n_n4078) & (x157x) & (!x339x) & (x13264x)) + ((!x13269x) & (n_n4078) & (x157x) & (x339x) & (!x13264x)) + ((!x13269x) & (n_n4078) & (x157x) & (x339x) & (x13264x)) + ((x13269x) & (!n_n4078) & (!x157x) & (!x339x) & (!x13264x)) + ((x13269x) & (!n_n4078) & (!x157x) & (!x339x) & (x13264x)) + ((x13269x) & (!n_n4078) & (!x157x) & (x339x) & (!x13264x)) + ((x13269x) & (!n_n4078) & (!x157x) & (x339x) & (x13264x)) + ((x13269x) & (!n_n4078) & (x157x) & (!x339x) & (!x13264x)) + ((x13269x) & (!n_n4078) & (x157x) & (!x339x) & (x13264x)) + ((x13269x) & (!n_n4078) & (x157x) & (x339x) & (!x13264x)) + ((x13269x) & (!n_n4078) & (x157x) & (x339x) & (x13264x)) + ((x13269x) & (n_n4078) & (!x157x) & (!x339x) & (!x13264x)) + ((x13269x) & (n_n4078) & (!x157x) & (!x339x) & (x13264x)) + ((x13269x) & (n_n4078) & (!x157x) & (x339x) & (!x13264x)) + ((x13269x) & (n_n4078) & (!x157x) & (x339x) & (x13264x)) + ((x13269x) & (n_n4078) & (x157x) & (!x339x) & (!x13264x)) + ((x13269x) & (n_n4078) & (x157x) & (!x339x) & (x13264x)) + ((x13269x) & (n_n4078) & (x157x) & (x339x) & (!x13264x)) + ((x13269x) & (n_n4078) & (x157x) & (x339x) & (x13264x)));
	assign x47x = (((i_7_) & (!i_8_) & (i_6_) & (x14x) & (n_n500)) + ((i_7_) & (i_8_) & (i_6_) & (x14x) & (n_n500)));
	assign x13276x = (((!n_n4751) & (!n_n4750) & (!n_n4752) & (!x47x) & (!x22125x)) + ((!n_n4751) & (!n_n4750) & (!n_n4752) & (x47x) & (!x22125x)) + ((!n_n4751) & (!n_n4750) & (!n_n4752) & (x47x) & (x22125x)) + ((!n_n4751) & (!n_n4750) & (n_n4752) & (!x47x) & (!x22125x)) + ((!n_n4751) & (!n_n4750) & (n_n4752) & (!x47x) & (x22125x)) + ((!n_n4751) & (!n_n4750) & (n_n4752) & (x47x) & (!x22125x)) + ((!n_n4751) & (!n_n4750) & (n_n4752) & (x47x) & (x22125x)) + ((!n_n4751) & (n_n4750) & (!n_n4752) & (!x47x) & (!x22125x)) + ((!n_n4751) & (n_n4750) & (!n_n4752) & (!x47x) & (x22125x)) + ((!n_n4751) & (n_n4750) & (!n_n4752) & (x47x) & (!x22125x)) + ((!n_n4751) & (n_n4750) & (!n_n4752) & (x47x) & (x22125x)) + ((!n_n4751) & (n_n4750) & (n_n4752) & (!x47x) & (!x22125x)) + ((!n_n4751) & (n_n4750) & (n_n4752) & (!x47x) & (x22125x)) + ((!n_n4751) & (n_n4750) & (n_n4752) & (x47x) & (!x22125x)) + ((!n_n4751) & (n_n4750) & (n_n4752) & (x47x) & (x22125x)) + ((n_n4751) & (!n_n4750) & (!n_n4752) & (!x47x) & (!x22125x)) + ((n_n4751) & (!n_n4750) & (!n_n4752) & (!x47x) & (x22125x)) + ((n_n4751) & (!n_n4750) & (!n_n4752) & (x47x) & (!x22125x)) + ((n_n4751) & (!n_n4750) & (!n_n4752) & (x47x) & (x22125x)) + ((n_n4751) & (!n_n4750) & (n_n4752) & (!x47x) & (!x22125x)) + ((n_n4751) & (!n_n4750) & (n_n4752) & (!x47x) & (x22125x)) + ((n_n4751) & (!n_n4750) & (n_n4752) & (x47x) & (!x22125x)) + ((n_n4751) & (!n_n4750) & (n_n4752) & (x47x) & (x22125x)) + ((n_n4751) & (n_n4750) & (!n_n4752) & (!x47x) & (!x22125x)) + ((n_n4751) & (n_n4750) & (!n_n4752) & (!x47x) & (x22125x)) + ((n_n4751) & (n_n4750) & (!n_n4752) & (x47x) & (!x22125x)) + ((n_n4751) & (n_n4750) & (!n_n4752) & (x47x) & (x22125x)) + ((n_n4751) & (n_n4750) & (n_n4752) & (!x47x) & (!x22125x)) + ((n_n4751) & (n_n4750) & (n_n4752) & (!x47x) & (x22125x)) + ((n_n4751) & (n_n4750) & (n_n4752) & (x47x) & (!x22125x)) + ((n_n4751) & (n_n4750) & (n_n4752) & (x47x) & (x22125x)));
	assign n_n5088 = (((i_7_) & (i_8_) & (!i_6_) & (n_n535) & (x12x)));
	assign n_n5078 = (((i_9_) & (n_n520) & (n_n195) & (n_n464)));
	assign n_n5083 = (((!i_9_) & (n_n532) & (n_n535) & (n_n130)));
	assign x123x = (((!i_9_) & (n_n535) & (!n_n130) & (x12x) & (n_n530)) + ((!i_9_) & (n_n535) & (n_n130) & (!x12x) & (n_n530)) + ((!i_9_) & (n_n535) & (n_n130) & (x12x) & (n_n530)) + ((i_9_) & (n_n535) & (!n_n130) & (x12x) & (n_n530)) + ((i_9_) & (n_n535) & (n_n130) & (x12x) & (n_n530)));
	assign x14644x = (((!n_n5081) & (!n_n5076) & (!n_n5075) & (n_n5079)) + ((!n_n5081) & (!n_n5076) & (n_n5075) & (!n_n5079)) + ((!n_n5081) & (!n_n5076) & (n_n5075) & (n_n5079)) + ((!n_n5081) & (n_n5076) & (!n_n5075) & (!n_n5079)) + ((!n_n5081) & (n_n5076) & (!n_n5075) & (n_n5079)) + ((!n_n5081) & (n_n5076) & (n_n5075) & (!n_n5079)) + ((!n_n5081) & (n_n5076) & (n_n5075) & (n_n5079)) + ((n_n5081) & (!n_n5076) & (!n_n5075) & (!n_n5079)) + ((n_n5081) & (!n_n5076) & (!n_n5075) & (n_n5079)) + ((n_n5081) & (!n_n5076) & (n_n5075) & (!n_n5079)) + ((n_n5081) & (!n_n5076) & (n_n5075) & (n_n5079)) + ((n_n5081) & (n_n5076) & (!n_n5075) & (!n_n5079)) + ((n_n5081) & (n_n5076) & (!n_n5075) & (n_n5079)) + ((n_n5081) & (n_n5076) & (n_n5075) & (!n_n5079)) + ((n_n5081) & (n_n5076) & (n_n5075) & (n_n5079)));
	assign x14645x = (((!n_n5085) & (!n_n5084) & (!n_n5088) & (!n_n5078) & (n_n5083)) + ((!n_n5085) & (!n_n5084) & (!n_n5088) & (n_n5078) & (!n_n5083)) + ((!n_n5085) & (!n_n5084) & (!n_n5088) & (n_n5078) & (n_n5083)) + ((!n_n5085) & (!n_n5084) & (n_n5088) & (!n_n5078) & (!n_n5083)) + ((!n_n5085) & (!n_n5084) & (n_n5088) & (!n_n5078) & (n_n5083)) + ((!n_n5085) & (!n_n5084) & (n_n5088) & (n_n5078) & (!n_n5083)) + ((!n_n5085) & (!n_n5084) & (n_n5088) & (n_n5078) & (n_n5083)) + ((!n_n5085) & (n_n5084) & (!n_n5088) & (!n_n5078) & (!n_n5083)) + ((!n_n5085) & (n_n5084) & (!n_n5088) & (!n_n5078) & (n_n5083)) + ((!n_n5085) & (n_n5084) & (!n_n5088) & (n_n5078) & (!n_n5083)) + ((!n_n5085) & (n_n5084) & (!n_n5088) & (n_n5078) & (n_n5083)) + ((!n_n5085) & (n_n5084) & (n_n5088) & (!n_n5078) & (!n_n5083)) + ((!n_n5085) & (n_n5084) & (n_n5088) & (!n_n5078) & (n_n5083)) + ((!n_n5085) & (n_n5084) & (n_n5088) & (n_n5078) & (!n_n5083)) + ((!n_n5085) & (n_n5084) & (n_n5088) & (n_n5078) & (n_n5083)) + ((n_n5085) & (!n_n5084) & (!n_n5088) & (!n_n5078) & (!n_n5083)) + ((n_n5085) & (!n_n5084) & (!n_n5088) & (!n_n5078) & (n_n5083)) + ((n_n5085) & (!n_n5084) & (!n_n5088) & (n_n5078) & (!n_n5083)) + ((n_n5085) & (!n_n5084) & (!n_n5088) & (n_n5078) & (n_n5083)) + ((n_n5085) & (!n_n5084) & (n_n5088) & (!n_n5078) & (!n_n5083)) + ((n_n5085) & (!n_n5084) & (n_n5088) & (!n_n5078) & (n_n5083)) + ((n_n5085) & (!n_n5084) & (n_n5088) & (n_n5078) & (!n_n5083)) + ((n_n5085) & (!n_n5084) & (n_n5088) & (n_n5078) & (n_n5083)) + ((n_n5085) & (n_n5084) & (!n_n5088) & (!n_n5078) & (!n_n5083)) + ((n_n5085) & (n_n5084) & (!n_n5088) & (!n_n5078) & (n_n5083)) + ((n_n5085) & (n_n5084) & (!n_n5088) & (n_n5078) & (!n_n5083)) + ((n_n5085) & (n_n5084) & (!n_n5088) & (n_n5078) & (n_n5083)) + ((n_n5085) & (n_n5084) & (n_n5088) & (!n_n5078) & (!n_n5083)) + ((n_n5085) & (n_n5084) & (n_n5088) & (!n_n5078) & (n_n5083)) + ((n_n5085) & (n_n5084) & (n_n5088) & (n_n5078) & (!n_n5083)) + ((n_n5085) & (n_n5084) & (n_n5088) & (n_n5078) & (n_n5083)));
	assign x122x = (((!i_9_) & (n_n518) & (!n_n532) & (n_n130) & (n_n530)) + ((!i_9_) & (n_n518) & (n_n532) & (n_n130) & (!n_n530)) + ((!i_9_) & (n_n518) & (n_n532) & (n_n130) & (n_n530)));
	assign n_n5090 = (((i_7_) & (!i_8_) & (!i_6_) & (n_n535) & (x12x)));
	assign x232x = (((!i_9_) & (n_n524) & (n_n535) & (!n_n130) & (x12x)) + ((!i_9_) & (n_n524) & (n_n535) & (n_n130) & (!x12x)) + ((!i_9_) & (n_n524) & (n_n535) & (n_n130) & (x12x)) + ((i_9_) & (n_n524) & (n_n535) & (!n_n130) & (x12x)) + ((i_9_) & (n_n524) & (n_n535) & (n_n130) & (x12x)));
	assign x14648x = (((!n_n5091) & (!n_n5099) & (!n_n5101) & (n_n5090)) + ((!n_n5091) & (!n_n5099) & (n_n5101) & (!n_n5090)) + ((!n_n5091) & (!n_n5099) & (n_n5101) & (n_n5090)) + ((!n_n5091) & (n_n5099) & (!n_n5101) & (!n_n5090)) + ((!n_n5091) & (n_n5099) & (!n_n5101) & (n_n5090)) + ((!n_n5091) & (n_n5099) & (n_n5101) & (!n_n5090)) + ((!n_n5091) & (n_n5099) & (n_n5101) & (n_n5090)) + ((n_n5091) & (!n_n5099) & (!n_n5101) & (!n_n5090)) + ((n_n5091) & (!n_n5099) & (!n_n5101) & (n_n5090)) + ((n_n5091) & (!n_n5099) & (n_n5101) & (!n_n5090)) + ((n_n5091) & (!n_n5099) & (n_n5101) & (n_n5090)) + ((n_n5091) & (n_n5099) & (!n_n5101) & (!n_n5090)) + ((n_n5091) & (n_n5099) & (!n_n5101) & (n_n5090)) + ((n_n5091) & (n_n5099) & (n_n5101) & (!n_n5090)) + ((n_n5091) & (n_n5099) & (n_n5101) & (n_n5090)));
	assign x14649x = (((!n_n5093) & (!n_n5089) & (!n_n5098) & (!n_n5103) & (n_n5095)) + ((!n_n5093) & (!n_n5089) & (!n_n5098) & (n_n5103) & (!n_n5095)) + ((!n_n5093) & (!n_n5089) & (!n_n5098) & (n_n5103) & (n_n5095)) + ((!n_n5093) & (!n_n5089) & (n_n5098) & (!n_n5103) & (!n_n5095)) + ((!n_n5093) & (!n_n5089) & (n_n5098) & (!n_n5103) & (n_n5095)) + ((!n_n5093) & (!n_n5089) & (n_n5098) & (n_n5103) & (!n_n5095)) + ((!n_n5093) & (!n_n5089) & (n_n5098) & (n_n5103) & (n_n5095)) + ((!n_n5093) & (n_n5089) & (!n_n5098) & (!n_n5103) & (!n_n5095)) + ((!n_n5093) & (n_n5089) & (!n_n5098) & (!n_n5103) & (n_n5095)) + ((!n_n5093) & (n_n5089) & (!n_n5098) & (n_n5103) & (!n_n5095)) + ((!n_n5093) & (n_n5089) & (!n_n5098) & (n_n5103) & (n_n5095)) + ((!n_n5093) & (n_n5089) & (n_n5098) & (!n_n5103) & (!n_n5095)) + ((!n_n5093) & (n_n5089) & (n_n5098) & (!n_n5103) & (n_n5095)) + ((!n_n5093) & (n_n5089) & (n_n5098) & (n_n5103) & (!n_n5095)) + ((!n_n5093) & (n_n5089) & (n_n5098) & (n_n5103) & (n_n5095)) + ((n_n5093) & (!n_n5089) & (!n_n5098) & (!n_n5103) & (!n_n5095)) + ((n_n5093) & (!n_n5089) & (!n_n5098) & (!n_n5103) & (n_n5095)) + ((n_n5093) & (!n_n5089) & (!n_n5098) & (n_n5103) & (!n_n5095)) + ((n_n5093) & (!n_n5089) & (!n_n5098) & (n_n5103) & (n_n5095)) + ((n_n5093) & (!n_n5089) & (n_n5098) & (!n_n5103) & (!n_n5095)) + ((n_n5093) & (!n_n5089) & (n_n5098) & (!n_n5103) & (n_n5095)) + ((n_n5093) & (!n_n5089) & (n_n5098) & (n_n5103) & (!n_n5095)) + ((n_n5093) & (!n_n5089) & (n_n5098) & (n_n5103) & (n_n5095)) + ((n_n5093) & (n_n5089) & (!n_n5098) & (!n_n5103) & (!n_n5095)) + ((n_n5093) & (n_n5089) & (!n_n5098) & (!n_n5103) & (n_n5095)) + ((n_n5093) & (n_n5089) & (!n_n5098) & (n_n5103) & (!n_n5095)) + ((n_n5093) & (n_n5089) & (!n_n5098) & (n_n5103) & (n_n5095)) + ((n_n5093) & (n_n5089) & (n_n5098) & (!n_n5103) & (!n_n5095)) + ((n_n5093) & (n_n5089) & (n_n5098) & (!n_n5103) & (n_n5095)) + ((n_n5093) & (n_n5089) & (n_n5098) & (n_n5103) & (!n_n5095)) + ((n_n5093) & (n_n5089) & (n_n5098) & (n_n5103) & (n_n5095)));
	assign n_n5068 = (((i_9_) & (n_n195) & (n_n530) & (n_n464)));
	assign x160x = (((!i_7_) & (i_8_) & (i_6_) & (x18x) & (n_n464)) + ((i_7_) & (!i_8_) & (i_6_) & (x18x) & (n_n464)));
	assign x14653x = (((!n_n524) & (!n_n473) & (!x18x) & (!n_n5063) & (n_n4152)) + ((!n_n524) & (!n_n473) & (!x18x) & (n_n5063) & (!n_n4152)) + ((!n_n524) & (!n_n473) & (!x18x) & (n_n5063) & (n_n4152)) + ((!n_n524) & (!n_n473) & (x18x) & (!n_n5063) & (n_n4152)) + ((!n_n524) & (!n_n473) & (x18x) & (n_n5063) & (!n_n4152)) + ((!n_n524) & (!n_n473) & (x18x) & (n_n5063) & (n_n4152)) + ((!n_n524) & (n_n473) & (!x18x) & (!n_n5063) & (n_n4152)) + ((!n_n524) & (n_n473) & (!x18x) & (n_n5063) & (!n_n4152)) + ((!n_n524) & (n_n473) & (!x18x) & (n_n5063) & (n_n4152)) + ((!n_n524) & (n_n473) & (x18x) & (!n_n5063) & (n_n4152)) + ((!n_n524) & (n_n473) & (x18x) & (n_n5063) & (!n_n4152)) + ((!n_n524) & (n_n473) & (x18x) & (n_n5063) & (n_n4152)) + ((n_n524) & (!n_n473) & (!x18x) & (!n_n5063) & (n_n4152)) + ((n_n524) & (!n_n473) & (!x18x) & (n_n5063) & (!n_n4152)) + ((n_n524) & (!n_n473) & (!x18x) & (n_n5063) & (n_n4152)) + ((n_n524) & (!n_n473) & (x18x) & (!n_n5063) & (n_n4152)) + ((n_n524) & (!n_n473) & (x18x) & (n_n5063) & (!n_n4152)) + ((n_n524) & (!n_n473) & (x18x) & (n_n5063) & (n_n4152)) + ((n_n524) & (n_n473) & (!x18x) & (!n_n5063) & (n_n4152)) + ((n_n524) & (n_n473) & (!x18x) & (n_n5063) & (!n_n4152)) + ((n_n524) & (n_n473) & (!x18x) & (n_n5063) & (n_n4152)) + ((n_n524) & (n_n473) & (x18x) & (!n_n5063) & (!n_n4152)) + ((n_n524) & (n_n473) & (x18x) & (!n_n5063) & (n_n4152)) + ((n_n524) & (n_n473) & (x18x) & (n_n5063) & (!n_n4152)) + ((n_n524) & (n_n473) & (x18x) & (n_n5063) & (n_n4152)));
	assign x14654x = (((!n_n5060) & (!n_n5070) & (!x160x) & (x14653x)) + ((!n_n5060) & (!n_n5070) & (x160x) & (!x14653x)) + ((!n_n5060) & (!n_n5070) & (x160x) & (x14653x)) + ((!n_n5060) & (n_n5070) & (!x160x) & (!x14653x)) + ((!n_n5060) & (n_n5070) & (!x160x) & (x14653x)) + ((!n_n5060) & (n_n5070) & (x160x) & (!x14653x)) + ((!n_n5060) & (n_n5070) & (x160x) & (x14653x)) + ((n_n5060) & (!n_n5070) & (!x160x) & (!x14653x)) + ((n_n5060) & (!n_n5070) & (!x160x) & (x14653x)) + ((n_n5060) & (!n_n5070) & (x160x) & (!x14653x)) + ((n_n5060) & (!n_n5070) & (x160x) & (x14653x)) + ((n_n5060) & (n_n5070) & (!x160x) & (!x14653x)) + ((n_n5060) & (n_n5070) & (!x160x) & (x14653x)) + ((n_n5060) & (n_n5070) & (x160x) & (!x14653x)) + ((n_n5060) & (n_n5070) & (x160x) & (x14653x)));
	assign n_n5077 = (((i_1_) & (!i_2_) & (!i_0_) & (x20x) & (n_n464)));
	assign x159x = (((!i_9_) & (!n_n528) & (n_n532) & (n_n195) & (n_n464)) + ((!i_9_) & (n_n528) & (!n_n532) & (n_n195) & (n_n464)) + ((!i_9_) & (n_n528) & (n_n532) & (n_n195) & (n_n464)));
	assign x22100x = (((!n_n5092) & (!n_n5110) & (!n_n5100) & (!n_n5097)));
	assign x14240x = (((!n_n5087) & (!n_n5065) & (!n_n5077) & (!x159x) & (!x22100x)) + ((!n_n5087) & (!n_n5065) & (!n_n5077) & (x159x) & (!x22100x)) + ((!n_n5087) & (!n_n5065) & (!n_n5077) & (x159x) & (x22100x)) + ((!n_n5087) & (!n_n5065) & (n_n5077) & (!x159x) & (!x22100x)) + ((!n_n5087) & (!n_n5065) & (n_n5077) & (!x159x) & (x22100x)) + ((!n_n5087) & (!n_n5065) & (n_n5077) & (x159x) & (!x22100x)) + ((!n_n5087) & (!n_n5065) & (n_n5077) & (x159x) & (x22100x)) + ((!n_n5087) & (n_n5065) & (!n_n5077) & (!x159x) & (!x22100x)) + ((!n_n5087) & (n_n5065) & (!n_n5077) & (!x159x) & (x22100x)) + ((!n_n5087) & (n_n5065) & (!n_n5077) & (x159x) & (!x22100x)) + ((!n_n5087) & (n_n5065) & (!n_n5077) & (x159x) & (x22100x)) + ((!n_n5087) & (n_n5065) & (n_n5077) & (!x159x) & (!x22100x)) + ((!n_n5087) & (n_n5065) & (n_n5077) & (!x159x) & (x22100x)) + ((!n_n5087) & (n_n5065) & (n_n5077) & (x159x) & (!x22100x)) + ((!n_n5087) & (n_n5065) & (n_n5077) & (x159x) & (x22100x)) + ((n_n5087) & (!n_n5065) & (!n_n5077) & (!x159x) & (!x22100x)) + ((n_n5087) & (!n_n5065) & (!n_n5077) & (!x159x) & (x22100x)) + ((n_n5087) & (!n_n5065) & (!n_n5077) & (x159x) & (!x22100x)) + ((n_n5087) & (!n_n5065) & (!n_n5077) & (x159x) & (x22100x)) + ((n_n5087) & (!n_n5065) & (n_n5077) & (!x159x) & (!x22100x)) + ((n_n5087) & (!n_n5065) & (n_n5077) & (!x159x) & (x22100x)) + ((n_n5087) & (!n_n5065) & (n_n5077) & (x159x) & (!x22100x)) + ((n_n5087) & (!n_n5065) & (n_n5077) & (x159x) & (x22100x)) + ((n_n5087) & (n_n5065) & (!n_n5077) & (!x159x) & (!x22100x)) + ((n_n5087) & (n_n5065) & (!n_n5077) & (!x159x) & (x22100x)) + ((n_n5087) & (n_n5065) & (!n_n5077) & (x159x) & (!x22100x)) + ((n_n5087) & (n_n5065) & (!n_n5077) & (x159x) & (x22100x)) + ((n_n5087) & (n_n5065) & (n_n5077) & (!x159x) & (!x22100x)) + ((n_n5087) & (n_n5065) & (n_n5077) & (!x159x) & (x22100x)) + ((n_n5087) & (n_n5065) & (n_n5077) & (x159x) & (!x22100x)) + ((n_n5087) & (n_n5065) & (n_n5077) & (x159x) & (x22100x)));
	assign x14226x = (((!n_n509) & (!n_n522) & (!x12x) & (!n_n5117) & (x125x)) + ((!n_n509) & (!n_n522) & (!x12x) & (n_n5117) & (!x125x)) + ((!n_n509) & (!n_n522) & (!x12x) & (n_n5117) & (x125x)) + ((!n_n509) & (!n_n522) & (x12x) & (!n_n5117) & (x125x)) + ((!n_n509) & (!n_n522) & (x12x) & (n_n5117) & (!x125x)) + ((!n_n509) & (!n_n522) & (x12x) & (n_n5117) & (x125x)) + ((!n_n509) & (n_n522) & (!x12x) & (!n_n5117) & (x125x)) + ((!n_n509) & (n_n522) & (!x12x) & (n_n5117) & (!x125x)) + ((!n_n509) & (n_n522) & (!x12x) & (n_n5117) & (x125x)) + ((!n_n509) & (n_n522) & (x12x) & (!n_n5117) & (x125x)) + ((!n_n509) & (n_n522) & (x12x) & (n_n5117) & (!x125x)) + ((!n_n509) & (n_n522) & (x12x) & (n_n5117) & (x125x)) + ((n_n509) & (!n_n522) & (!x12x) & (!n_n5117) & (x125x)) + ((n_n509) & (!n_n522) & (!x12x) & (n_n5117) & (!x125x)) + ((n_n509) & (!n_n522) & (!x12x) & (n_n5117) & (x125x)) + ((n_n509) & (!n_n522) & (x12x) & (!n_n5117) & (x125x)) + ((n_n509) & (!n_n522) & (x12x) & (n_n5117) & (!x125x)) + ((n_n509) & (!n_n522) & (x12x) & (n_n5117) & (x125x)) + ((n_n509) & (n_n522) & (!x12x) & (!n_n5117) & (x125x)) + ((n_n509) & (n_n522) & (!x12x) & (n_n5117) & (!x125x)) + ((n_n509) & (n_n522) & (!x12x) & (n_n5117) & (x125x)) + ((n_n509) & (n_n522) & (x12x) & (!n_n5117) & (!x125x)) + ((n_n509) & (n_n522) & (x12x) & (!n_n5117) & (x125x)) + ((n_n509) & (n_n522) & (x12x) & (n_n5117) & (!x125x)) + ((n_n509) & (n_n522) & (x12x) & (n_n5117) & (x125x)));
	assign x14227x = (((!n_n5161) & (!n_n5135) & (!n_n5152) & (!n_n5153) & (n_n5160)) + ((!n_n5161) & (!n_n5135) & (!n_n5152) & (n_n5153) & (!n_n5160)) + ((!n_n5161) & (!n_n5135) & (!n_n5152) & (n_n5153) & (n_n5160)) + ((!n_n5161) & (!n_n5135) & (n_n5152) & (!n_n5153) & (!n_n5160)) + ((!n_n5161) & (!n_n5135) & (n_n5152) & (!n_n5153) & (n_n5160)) + ((!n_n5161) & (!n_n5135) & (n_n5152) & (n_n5153) & (!n_n5160)) + ((!n_n5161) & (!n_n5135) & (n_n5152) & (n_n5153) & (n_n5160)) + ((!n_n5161) & (n_n5135) & (!n_n5152) & (!n_n5153) & (!n_n5160)) + ((!n_n5161) & (n_n5135) & (!n_n5152) & (!n_n5153) & (n_n5160)) + ((!n_n5161) & (n_n5135) & (!n_n5152) & (n_n5153) & (!n_n5160)) + ((!n_n5161) & (n_n5135) & (!n_n5152) & (n_n5153) & (n_n5160)) + ((!n_n5161) & (n_n5135) & (n_n5152) & (!n_n5153) & (!n_n5160)) + ((!n_n5161) & (n_n5135) & (n_n5152) & (!n_n5153) & (n_n5160)) + ((!n_n5161) & (n_n5135) & (n_n5152) & (n_n5153) & (!n_n5160)) + ((!n_n5161) & (n_n5135) & (n_n5152) & (n_n5153) & (n_n5160)) + ((n_n5161) & (!n_n5135) & (!n_n5152) & (!n_n5153) & (!n_n5160)) + ((n_n5161) & (!n_n5135) & (!n_n5152) & (!n_n5153) & (n_n5160)) + ((n_n5161) & (!n_n5135) & (!n_n5152) & (n_n5153) & (!n_n5160)) + ((n_n5161) & (!n_n5135) & (!n_n5152) & (n_n5153) & (n_n5160)) + ((n_n5161) & (!n_n5135) & (n_n5152) & (!n_n5153) & (!n_n5160)) + ((n_n5161) & (!n_n5135) & (n_n5152) & (!n_n5153) & (n_n5160)) + ((n_n5161) & (!n_n5135) & (n_n5152) & (n_n5153) & (!n_n5160)) + ((n_n5161) & (!n_n5135) & (n_n5152) & (n_n5153) & (n_n5160)) + ((n_n5161) & (n_n5135) & (!n_n5152) & (!n_n5153) & (!n_n5160)) + ((n_n5161) & (n_n5135) & (!n_n5152) & (!n_n5153) & (n_n5160)) + ((n_n5161) & (n_n5135) & (!n_n5152) & (n_n5153) & (!n_n5160)) + ((n_n5161) & (n_n5135) & (!n_n5152) & (n_n5153) & (n_n5160)) + ((n_n5161) & (n_n5135) & (n_n5152) & (!n_n5153) & (!n_n5160)) + ((n_n5161) & (n_n5135) & (n_n5152) & (!n_n5153) & (n_n5160)) + ((n_n5161) & (n_n5135) & (n_n5152) & (n_n5153) & (!n_n5160)) + ((n_n5161) & (n_n5135) & (n_n5152) & (n_n5153) & (n_n5160)));
	assign x14232x = (((!n_n5172) & (!n_n5207) & (!n_n5169) & (n_n5197)) + ((!n_n5172) & (!n_n5207) & (n_n5169) & (!n_n5197)) + ((!n_n5172) & (!n_n5207) & (n_n5169) & (n_n5197)) + ((!n_n5172) & (n_n5207) & (!n_n5169) & (!n_n5197)) + ((!n_n5172) & (n_n5207) & (!n_n5169) & (n_n5197)) + ((!n_n5172) & (n_n5207) & (n_n5169) & (!n_n5197)) + ((!n_n5172) & (n_n5207) & (n_n5169) & (n_n5197)) + ((n_n5172) & (!n_n5207) & (!n_n5169) & (!n_n5197)) + ((n_n5172) & (!n_n5207) & (!n_n5169) & (n_n5197)) + ((n_n5172) & (!n_n5207) & (n_n5169) & (!n_n5197)) + ((n_n5172) & (!n_n5207) & (n_n5169) & (n_n5197)) + ((n_n5172) & (n_n5207) & (!n_n5169) & (!n_n5197)) + ((n_n5172) & (n_n5207) & (!n_n5169) & (n_n5197)) + ((n_n5172) & (n_n5207) & (n_n5169) & (!n_n5197)) + ((n_n5172) & (n_n5207) & (n_n5169) & (n_n5197)));
	assign x14233x = (((!n_n5167) & (!n_n5166) & (!n_n5176) & (!n_n5205) & (n_n5211)) + ((!n_n5167) & (!n_n5166) & (!n_n5176) & (n_n5205) & (!n_n5211)) + ((!n_n5167) & (!n_n5166) & (!n_n5176) & (n_n5205) & (n_n5211)) + ((!n_n5167) & (!n_n5166) & (n_n5176) & (!n_n5205) & (!n_n5211)) + ((!n_n5167) & (!n_n5166) & (n_n5176) & (!n_n5205) & (n_n5211)) + ((!n_n5167) & (!n_n5166) & (n_n5176) & (n_n5205) & (!n_n5211)) + ((!n_n5167) & (!n_n5166) & (n_n5176) & (n_n5205) & (n_n5211)) + ((!n_n5167) & (n_n5166) & (!n_n5176) & (!n_n5205) & (!n_n5211)) + ((!n_n5167) & (n_n5166) & (!n_n5176) & (!n_n5205) & (n_n5211)) + ((!n_n5167) & (n_n5166) & (!n_n5176) & (n_n5205) & (!n_n5211)) + ((!n_n5167) & (n_n5166) & (!n_n5176) & (n_n5205) & (n_n5211)) + ((!n_n5167) & (n_n5166) & (n_n5176) & (!n_n5205) & (!n_n5211)) + ((!n_n5167) & (n_n5166) & (n_n5176) & (!n_n5205) & (n_n5211)) + ((!n_n5167) & (n_n5166) & (n_n5176) & (n_n5205) & (!n_n5211)) + ((!n_n5167) & (n_n5166) & (n_n5176) & (n_n5205) & (n_n5211)) + ((n_n5167) & (!n_n5166) & (!n_n5176) & (!n_n5205) & (!n_n5211)) + ((n_n5167) & (!n_n5166) & (!n_n5176) & (!n_n5205) & (n_n5211)) + ((n_n5167) & (!n_n5166) & (!n_n5176) & (n_n5205) & (!n_n5211)) + ((n_n5167) & (!n_n5166) & (!n_n5176) & (n_n5205) & (n_n5211)) + ((n_n5167) & (!n_n5166) & (n_n5176) & (!n_n5205) & (!n_n5211)) + ((n_n5167) & (!n_n5166) & (n_n5176) & (!n_n5205) & (n_n5211)) + ((n_n5167) & (!n_n5166) & (n_n5176) & (n_n5205) & (!n_n5211)) + ((n_n5167) & (!n_n5166) & (n_n5176) & (n_n5205) & (n_n5211)) + ((n_n5167) & (n_n5166) & (!n_n5176) & (!n_n5205) & (!n_n5211)) + ((n_n5167) & (n_n5166) & (!n_n5176) & (!n_n5205) & (n_n5211)) + ((n_n5167) & (n_n5166) & (!n_n5176) & (n_n5205) & (!n_n5211)) + ((n_n5167) & (n_n5166) & (!n_n5176) & (n_n5205) & (n_n5211)) + ((n_n5167) & (n_n5166) & (n_n5176) & (!n_n5205) & (!n_n5211)) + ((n_n5167) & (n_n5166) & (n_n5176) & (!n_n5205) & (n_n5211)) + ((n_n5167) & (n_n5166) & (n_n5176) & (n_n5205) & (!n_n5211)) + ((n_n5167) & (n_n5166) & (n_n5176) & (n_n5205) & (n_n5211)));
	assign x435x = (((!i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n509)) + ((i_7_) & (!i_8_) & (!i_6_) & (x19x) & (n_n509)));
	assign x14253x = (((!n_n5232) & (!n_n5255) & (!n_n5212) & (n_n5249)) + ((!n_n5232) & (!n_n5255) & (n_n5212) & (!n_n5249)) + ((!n_n5232) & (!n_n5255) & (n_n5212) & (n_n5249)) + ((!n_n5232) & (n_n5255) & (!n_n5212) & (!n_n5249)) + ((!n_n5232) & (n_n5255) & (!n_n5212) & (n_n5249)) + ((!n_n5232) & (n_n5255) & (n_n5212) & (!n_n5249)) + ((!n_n5232) & (n_n5255) & (n_n5212) & (n_n5249)) + ((n_n5232) & (!n_n5255) & (!n_n5212) & (!n_n5249)) + ((n_n5232) & (!n_n5255) & (!n_n5212) & (n_n5249)) + ((n_n5232) & (!n_n5255) & (n_n5212) & (!n_n5249)) + ((n_n5232) & (!n_n5255) & (n_n5212) & (n_n5249)) + ((n_n5232) & (n_n5255) & (!n_n5212) & (!n_n5249)) + ((n_n5232) & (n_n5255) & (!n_n5212) & (n_n5249)) + ((n_n5232) & (n_n5255) & (n_n5212) & (!n_n5249)) + ((n_n5232) & (n_n5255) & (n_n5212) & (n_n5249)));
	assign x14254x = (((!n_n5308) & (!n_n5237) & (!n_n5226) & (n_n5218)) + ((!n_n5308) & (!n_n5237) & (n_n5226) & (!n_n5218)) + ((!n_n5308) & (!n_n5237) & (n_n5226) & (n_n5218)) + ((!n_n5308) & (n_n5237) & (!n_n5226) & (!n_n5218)) + ((!n_n5308) & (n_n5237) & (!n_n5226) & (n_n5218)) + ((!n_n5308) & (n_n5237) & (n_n5226) & (!n_n5218)) + ((!n_n5308) & (n_n5237) & (n_n5226) & (n_n5218)) + ((n_n5308) & (!n_n5237) & (!n_n5226) & (!n_n5218)) + ((n_n5308) & (!n_n5237) & (!n_n5226) & (n_n5218)) + ((n_n5308) & (!n_n5237) & (n_n5226) & (!n_n5218)) + ((n_n5308) & (!n_n5237) & (n_n5226) & (n_n5218)) + ((n_n5308) & (n_n5237) & (!n_n5226) & (!n_n5218)) + ((n_n5308) & (n_n5237) & (!n_n5226) & (n_n5218)) + ((n_n5308) & (n_n5237) & (n_n5226) & (!n_n5218)) + ((n_n5308) & (n_n5237) & (n_n5226) & (n_n5218)));
	assign x14256x = (((!n_n5320) & (!n_n5325) & (!x435x) & (!x14253x) & (x14254x)) + ((!n_n5320) & (!n_n5325) & (!x435x) & (x14253x) & (!x14254x)) + ((!n_n5320) & (!n_n5325) & (!x435x) & (x14253x) & (x14254x)) + ((!n_n5320) & (!n_n5325) & (x435x) & (!x14253x) & (!x14254x)) + ((!n_n5320) & (!n_n5325) & (x435x) & (!x14253x) & (x14254x)) + ((!n_n5320) & (!n_n5325) & (x435x) & (x14253x) & (!x14254x)) + ((!n_n5320) & (!n_n5325) & (x435x) & (x14253x) & (x14254x)) + ((!n_n5320) & (n_n5325) & (!x435x) & (!x14253x) & (!x14254x)) + ((!n_n5320) & (n_n5325) & (!x435x) & (!x14253x) & (x14254x)) + ((!n_n5320) & (n_n5325) & (!x435x) & (x14253x) & (!x14254x)) + ((!n_n5320) & (n_n5325) & (!x435x) & (x14253x) & (x14254x)) + ((!n_n5320) & (n_n5325) & (x435x) & (!x14253x) & (!x14254x)) + ((!n_n5320) & (n_n5325) & (x435x) & (!x14253x) & (x14254x)) + ((!n_n5320) & (n_n5325) & (x435x) & (x14253x) & (!x14254x)) + ((!n_n5320) & (n_n5325) & (x435x) & (x14253x) & (x14254x)) + ((n_n5320) & (!n_n5325) & (!x435x) & (!x14253x) & (!x14254x)) + ((n_n5320) & (!n_n5325) & (!x435x) & (!x14253x) & (x14254x)) + ((n_n5320) & (!n_n5325) & (!x435x) & (x14253x) & (!x14254x)) + ((n_n5320) & (!n_n5325) & (!x435x) & (x14253x) & (x14254x)) + ((n_n5320) & (!n_n5325) & (x435x) & (!x14253x) & (!x14254x)) + ((n_n5320) & (!n_n5325) & (x435x) & (!x14253x) & (x14254x)) + ((n_n5320) & (!n_n5325) & (x435x) & (x14253x) & (!x14254x)) + ((n_n5320) & (!n_n5325) & (x435x) & (x14253x) & (x14254x)) + ((n_n5320) & (n_n5325) & (!x435x) & (!x14253x) & (!x14254x)) + ((n_n5320) & (n_n5325) & (!x435x) & (!x14253x) & (x14254x)) + ((n_n5320) & (n_n5325) & (!x435x) & (x14253x) & (!x14254x)) + ((n_n5320) & (n_n5325) & (!x435x) & (x14253x) & (x14254x)) + ((n_n5320) & (n_n5325) & (x435x) & (!x14253x) & (!x14254x)) + ((n_n5320) & (n_n5325) & (x435x) & (!x14253x) & (x14254x)) + ((n_n5320) & (n_n5325) & (x435x) & (x14253x) & (!x14254x)) + ((n_n5320) & (n_n5325) & (x435x) & (x14253x) & (x14254x)));
	assign x14246x = (((!n_n5290) & (!n_n5295) & (!n_n5256) & (!n_n5257) & (n_n5283)) + ((!n_n5290) & (!n_n5295) & (!n_n5256) & (n_n5257) & (!n_n5283)) + ((!n_n5290) & (!n_n5295) & (!n_n5256) & (n_n5257) & (n_n5283)) + ((!n_n5290) & (!n_n5295) & (n_n5256) & (!n_n5257) & (!n_n5283)) + ((!n_n5290) & (!n_n5295) & (n_n5256) & (!n_n5257) & (n_n5283)) + ((!n_n5290) & (!n_n5295) & (n_n5256) & (n_n5257) & (!n_n5283)) + ((!n_n5290) & (!n_n5295) & (n_n5256) & (n_n5257) & (n_n5283)) + ((!n_n5290) & (n_n5295) & (!n_n5256) & (!n_n5257) & (!n_n5283)) + ((!n_n5290) & (n_n5295) & (!n_n5256) & (!n_n5257) & (n_n5283)) + ((!n_n5290) & (n_n5295) & (!n_n5256) & (n_n5257) & (!n_n5283)) + ((!n_n5290) & (n_n5295) & (!n_n5256) & (n_n5257) & (n_n5283)) + ((!n_n5290) & (n_n5295) & (n_n5256) & (!n_n5257) & (!n_n5283)) + ((!n_n5290) & (n_n5295) & (n_n5256) & (!n_n5257) & (n_n5283)) + ((!n_n5290) & (n_n5295) & (n_n5256) & (n_n5257) & (!n_n5283)) + ((!n_n5290) & (n_n5295) & (n_n5256) & (n_n5257) & (n_n5283)) + ((n_n5290) & (!n_n5295) & (!n_n5256) & (!n_n5257) & (!n_n5283)) + ((n_n5290) & (!n_n5295) & (!n_n5256) & (!n_n5257) & (n_n5283)) + ((n_n5290) & (!n_n5295) & (!n_n5256) & (n_n5257) & (!n_n5283)) + ((n_n5290) & (!n_n5295) & (!n_n5256) & (n_n5257) & (n_n5283)) + ((n_n5290) & (!n_n5295) & (n_n5256) & (!n_n5257) & (!n_n5283)) + ((n_n5290) & (!n_n5295) & (n_n5256) & (!n_n5257) & (n_n5283)) + ((n_n5290) & (!n_n5295) & (n_n5256) & (n_n5257) & (!n_n5283)) + ((n_n5290) & (!n_n5295) & (n_n5256) & (n_n5257) & (n_n5283)) + ((n_n5290) & (n_n5295) & (!n_n5256) & (!n_n5257) & (!n_n5283)) + ((n_n5290) & (n_n5295) & (!n_n5256) & (!n_n5257) & (n_n5283)) + ((n_n5290) & (n_n5295) & (!n_n5256) & (n_n5257) & (!n_n5283)) + ((n_n5290) & (n_n5295) & (!n_n5256) & (n_n5257) & (n_n5283)) + ((n_n5290) & (n_n5295) & (n_n5256) & (!n_n5257) & (!n_n5283)) + ((n_n5290) & (n_n5295) & (n_n5256) & (!n_n5257) & (n_n5283)) + ((n_n5290) & (n_n5295) & (n_n5256) & (n_n5257) & (!n_n5283)) + ((n_n5290) & (n_n5295) & (n_n5256) & (n_n5257) & (n_n5283)));
	assign x14261x = (((!n_n4895) & (!n_n4825) & (!n_n4879) & (n_n4841)) + ((!n_n4895) & (!n_n4825) & (n_n4879) & (!n_n4841)) + ((!n_n4895) & (!n_n4825) & (n_n4879) & (n_n4841)) + ((!n_n4895) & (n_n4825) & (!n_n4879) & (!n_n4841)) + ((!n_n4895) & (n_n4825) & (!n_n4879) & (n_n4841)) + ((!n_n4895) & (n_n4825) & (n_n4879) & (!n_n4841)) + ((!n_n4895) & (n_n4825) & (n_n4879) & (n_n4841)) + ((n_n4895) & (!n_n4825) & (!n_n4879) & (!n_n4841)) + ((n_n4895) & (!n_n4825) & (!n_n4879) & (n_n4841)) + ((n_n4895) & (!n_n4825) & (n_n4879) & (!n_n4841)) + ((n_n4895) & (!n_n4825) & (n_n4879) & (n_n4841)) + ((n_n4895) & (n_n4825) & (!n_n4879) & (!n_n4841)) + ((n_n4895) & (n_n4825) & (!n_n4879) & (n_n4841)) + ((n_n4895) & (n_n4825) & (n_n4879) & (!n_n4841)) + ((n_n4895) & (n_n4825) & (n_n4879) & (n_n4841)));
	assign x14262x = (((!n_n4883) & (!n_n4869) & (!n_n4870) & (!n_n4836) & (n_n4891)) + ((!n_n4883) & (!n_n4869) & (!n_n4870) & (n_n4836) & (!n_n4891)) + ((!n_n4883) & (!n_n4869) & (!n_n4870) & (n_n4836) & (n_n4891)) + ((!n_n4883) & (!n_n4869) & (n_n4870) & (!n_n4836) & (!n_n4891)) + ((!n_n4883) & (!n_n4869) & (n_n4870) & (!n_n4836) & (n_n4891)) + ((!n_n4883) & (!n_n4869) & (n_n4870) & (n_n4836) & (!n_n4891)) + ((!n_n4883) & (!n_n4869) & (n_n4870) & (n_n4836) & (n_n4891)) + ((!n_n4883) & (n_n4869) & (!n_n4870) & (!n_n4836) & (!n_n4891)) + ((!n_n4883) & (n_n4869) & (!n_n4870) & (!n_n4836) & (n_n4891)) + ((!n_n4883) & (n_n4869) & (!n_n4870) & (n_n4836) & (!n_n4891)) + ((!n_n4883) & (n_n4869) & (!n_n4870) & (n_n4836) & (n_n4891)) + ((!n_n4883) & (n_n4869) & (n_n4870) & (!n_n4836) & (!n_n4891)) + ((!n_n4883) & (n_n4869) & (n_n4870) & (!n_n4836) & (n_n4891)) + ((!n_n4883) & (n_n4869) & (n_n4870) & (n_n4836) & (!n_n4891)) + ((!n_n4883) & (n_n4869) & (n_n4870) & (n_n4836) & (n_n4891)) + ((n_n4883) & (!n_n4869) & (!n_n4870) & (!n_n4836) & (!n_n4891)) + ((n_n4883) & (!n_n4869) & (!n_n4870) & (!n_n4836) & (n_n4891)) + ((n_n4883) & (!n_n4869) & (!n_n4870) & (n_n4836) & (!n_n4891)) + ((n_n4883) & (!n_n4869) & (!n_n4870) & (n_n4836) & (n_n4891)) + ((n_n4883) & (!n_n4869) & (n_n4870) & (!n_n4836) & (!n_n4891)) + ((n_n4883) & (!n_n4869) & (n_n4870) & (!n_n4836) & (n_n4891)) + ((n_n4883) & (!n_n4869) & (n_n4870) & (n_n4836) & (!n_n4891)) + ((n_n4883) & (!n_n4869) & (n_n4870) & (n_n4836) & (n_n4891)) + ((n_n4883) & (n_n4869) & (!n_n4870) & (!n_n4836) & (!n_n4891)) + ((n_n4883) & (n_n4869) & (!n_n4870) & (!n_n4836) & (n_n4891)) + ((n_n4883) & (n_n4869) & (!n_n4870) & (n_n4836) & (!n_n4891)) + ((n_n4883) & (n_n4869) & (!n_n4870) & (n_n4836) & (n_n4891)) + ((n_n4883) & (n_n4869) & (n_n4870) & (!n_n4836) & (!n_n4891)) + ((n_n4883) & (n_n4869) & (n_n4870) & (!n_n4836) & (n_n4891)) + ((n_n4883) & (n_n4869) & (n_n4870) & (n_n4836) & (!n_n4891)) + ((n_n4883) & (n_n4869) & (n_n4870) & (n_n4836) & (n_n4891)));
	assign x14267x = (((!n_n4958) & (!n_n4921) & (!n_n4963) & (n_n4916)) + ((!n_n4958) & (!n_n4921) & (n_n4963) & (!n_n4916)) + ((!n_n4958) & (!n_n4921) & (n_n4963) & (n_n4916)) + ((!n_n4958) & (n_n4921) & (!n_n4963) & (!n_n4916)) + ((!n_n4958) & (n_n4921) & (!n_n4963) & (n_n4916)) + ((!n_n4958) & (n_n4921) & (n_n4963) & (!n_n4916)) + ((!n_n4958) & (n_n4921) & (n_n4963) & (n_n4916)) + ((n_n4958) & (!n_n4921) & (!n_n4963) & (!n_n4916)) + ((n_n4958) & (!n_n4921) & (!n_n4963) & (n_n4916)) + ((n_n4958) & (!n_n4921) & (n_n4963) & (!n_n4916)) + ((n_n4958) & (!n_n4921) & (n_n4963) & (n_n4916)) + ((n_n4958) & (n_n4921) & (!n_n4963) & (!n_n4916)) + ((n_n4958) & (n_n4921) & (!n_n4963) & (n_n4916)) + ((n_n4958) & (n_n4921) & (n_n4963) & (!n_n4916)) + ((n_n4958) & (n_n4921) & (n_n4963) & (n_n4916)));
	assign x14268x = (((!x352x) & (!n_n4933) & (!n_n4973) & (n_n4948)) + ((!x352x) & (!n_n4933) & (n_n4973) & (!n_n4948)) + ((!x352x) & (!n_n4933) & (n_n4973) & (n_n4948)) + ((!x352x) & (n_n4933) & (!n_n4973) & (!n_n4948)) + ((!x352x) & (n_n4933) & (!n_n4973) & (n_n4948)) + ((!x352x) & (n_n4933) & (n_n4973) & (!n_n4948)) + ((!x352x) & (n_n4933) & (n_n4973) & (n_n4948)) + ((x352x) & (!n_n4933) & (!n_n4973) & (!n_n4948)) + ((x352x) & (!n_n4933) & (!n_n4973) & (n_n4948)) + ((x352x) & (!n_n4933) & (n_n4973) & (!n_n4948)) + ((x352x) & (!n_n4933) & (n_n4973) & (n_n4948)) + ((x352x) & (n_n4933) & (!n_n4973) & (!n_n4948)) + ((x352x) & (n_n4933) & (!n_n4973) & (n_n4948)) + ((x352x) & (n_n4933) & (n_n4973) & (!n_n4948)) + ((x352x) & (n_n4933) & (n_n4973) & (n_n4948)));
	assign x275x = (((!i_9_) & (n_n473) & (!n_n520) & (n_n195) & (x20x)) + ((!i_9_) & (n_n473) & (n_n520) & (n_n195) & (x20x)) + ((i_9_) & (n_n473) & (!n_n520) & (n_n195) & (x20x)) + ((i_9_) & (n_n473) & (n_n520) & (n_n195) & (!x20x)) + ((i_9_) & (n_n473) & (n_n520) & (n_n195) & (x20x)));
	assign n_n4370 = (((i_9_) & (n_n536) & (n_n524) & (n_n500)));
	assign n_n4435 = (((!i_9_) & (n_n536) & (n_n524) & (n_n464)));
	assign n_n4493 = (((!i_9_) & (n_n455) & (n_n500) & (n_n530)));
	assign x14284x = (((!n_n4432) & (!n_n4480) & (!n_n4486) & (!n_n4435) & (n_n4493)) + ((!n_n4432) & (!n_n4480) & (!n_n4486) & (n_n4435) & (!n_n4493)) + ((!n_n4432) & (!n_n4480) & (!n_n4486) & (n_n4435) & (n_n4493)) + ((!n_n4432) & (!n_n4480) & (n_n4486) & (!n_n4435) & (!n_n4493)) + ((!n_n4432) & (!n_n4480) & (n_n4486) & (!n_n4435) & (n_n4493)) + ((!n_n4432) & (!n_n4480) & (n_n4486) & (n_n4435) & (!n_n4493)) + ((!n_n4432) & (!n_n4480) & (n_n4486) & (n_n4435) & (n_n4493)) + ((!n_n4432) & (n_n4480) & (!n_n4486) & (!n_n4435) & (!n_n4493)) + ((!n_n4432) & (n_n4480) & (!n_n4486) & (!n_n4435) & (n_n4493)) + ((!n_n4432) & (n_n4480) & (!n_n4486) & (n_n4435) & (!n_n4493)) + ((!n_n4432) & (n_n4480) & (!n_n4486) & (n_n4435) & (n_n4493)) + ((!n_n4432) & (n_n4480) & (n_n4486) & (!n_n4435) & (!n_n4493)) + ((!n_n4432) & (n_n4480) & (n_n4486) & (!n_n4435) & (n_n4493)) + ((!n_n4432) & (n_n4480) & (n_n4486) & (n_n4435) & (!n_n4493)) + ((!n_n4432) & (n_n4480) & (n_n4486) & (n_n4435) & (n_n4493)) + ((n_n4432) & (!n_n4480) & (!n_n4486) & (!n_n4435) & (!n_n4493)) + ((n_n4432) & (!n_n4480) & (!n_n4486) & (!n_n4435) & (n_n4493)) + ((n_n4432) & (!n_n4480) & (!n_n4486) & (n_n4435) & (!n_n4493)) + ((n_n4432) & (!n_n4480) & (!n_n4486) & (n_n4435) & (n_n4493)) + ((n_n4432) & (!n_n4480) & (n_n4486) & (!n_n4435) & (!n_n4493)) + ((n_n4432) & (!n_n4480) & (n_n4486) & (!n_n4435) & (n_n4493)) + ((n_n4432) & (!n_n4480) & (n_n4486) & (n_n4435) & (!n_n4493)) + ((n_n4432) & (!n_n4480) & (n_n4486) & (n_n4435) & (n_n4493)) + ((n_n4432) & (n_n4480) & (!n_n4486) & (!n_n4435) & (!n_n4493)) + ((n_n4432) & (n_n4480) & (!n_n4486) & (!n_n4435) & (n_n4493)) + ((n_n4432) & (n_n4480) & (!n_n4486) & (n_n4435) & (!n_n4493)) + ((n_n4432) & (n_n4480) & (!n_n4486) & (n_n4435) & (n_n4493)) + ((n_n4432) & (n_n4480) & (n_n4486) & (!n_n4435) & (!n_n4493)) + ((n_n4432) & (n_n4480) & (n_n4486) & (!n_n4435) & (n_n4493)) + ((n_n4432) & (n_n4480) & (n_n4486) & (n_n4435) & (!n_n4493)) + ((n_n4432) & (n_n4480) & (n_n4486) & (n_n4435) & (n_n4493)));
	assign n_n3565 = (((!n_n4464) & (!n_n4467) & (!n_n4451) & (!n_n4449) & (x14284x)) + ((!n_n4464) & (!n_n4467) & (!n_n4451) & (n_n4449) & (!x14284x)) + ((!n_n4464) & (!n_n4467) & (!n_n4451) & (n_n4449) & (x14284x)) + ((!n_n4464) & (!n_n4467) & (n_n4451) & (!n_n4449) & (!x14284x)) + ((!n_n4464) & (!n_n4467) & (n_n4451) & (!n_n4449) & (x14284x)) + ((!n_n4464) & (!n_n4467) & (n_n4451) & (n_n4449) & (!x14284x)) + ((!n_n4464) & (!n_n4467) & (n_n4451) & (n_n4449) & (x14284x)) + ((!n_n4464) & (n_n4467) & (!n_n4451) & (!n_n4449) & (!x14284x)) + ((!n_n4464) & (n_n4467) & (!n_n4451) & (!n_n4449) & (x14284x)) + ((!n_n4464) & (n_n4467) & (!n_n4451) & (n_n4449) & (!x14284x)) + ((!n_n4464) & (n_n4467) & (!n_n4451) & (n_n4449) & (x14284x)) + ((!n_n4464) & (n_n4467) & (n_n4451) & (!n_n4449) & (!x14284x)) + ((!n_n4464) & (n_n4467) & (n_n4451) & (!n_n4449) & (x14284x)) + ((!n_n4464) & (n_n4467) & (n_n4451) & (n_n4449) & (!x14284x)) + ((!n_n4464) & (n_n4467) & (n_n4451) & (n_n4449) & (x14284x)) + ((n_n4464) & (!n_n4467) & (!n_n4451) & (!n_n4449) & (!x14284x)) + ((n_n4464) & (!n_n4467) & (!n_n4451) & (!n_n4449) & (x14284x)) + ((n_n4464) & (!n_n4467) & (!n_n4451) & (n_n4449) & (!x14284x)) + ((n_n4464) & (!n_n4467) & (!n_n4451) & (n_n4449) & (x14284x)) + ((n_n4464) & (!n_n4467) & (n_n4451) & (!n_n4449) & (!x14284x)) + ((n_n4464) & (!n_n4467) & (n_n4451) & (!n_n4449) & (x14284x)) + ((n_n4464) & (!n_n4467) & (n_n4451) & (n_n4449) & (!x14284x)) + ((n_n4464) & (!n_n4467) & (n_n4451) & (n_n4449) & (x14284x)) + ((n_n4464) & (n_n4467) & (!n_n4451) & (!n_n4449) & (!x14284x)) + ((n_n4464) & (n_n4467) & (!n_n4451) & (!n_n4449) & (x14284x)) + ((n_n4464) & (n_n4467) & (!n_n4451) & (n_n4449) & (!x14284x)) + ((n_n4464) & (n_n4467) & (!n_n4451) & (n_n4449) & (x14284x)) + ((n_n4464) & (n_n4467) & (n_n4451) & (!n_n4449) & (!x14284x)) + ((n_n4464) & (n_n4467) & (n_n4451) & (!n_n4449) & (x14284x)) + ((n_n4464) & (n_n4467) & (n_n4451) & (n_n4449) & (!x14284x)) + ((n_n4464) & (n_n4467) & (n_n4451) & (n_n4449) & (x14284x)));
	assign x14290x = (((!n_n4317) & (!n_n4362) & (!n_n4319) & (n_n4336)) + ((!n_n4317) & (!n_n4362) & (n_n4319) & (!n_n4336)) + ((!n_n4317) & (!n_n4362) & (n_n4319) & (n_n4336)) + ((!n_n4317) & (n_n4362) & (!n_n4319) & (!n_n4336)) + ((!n_n4317) & (n_n4362) & (!n_n4319) & (n_n4336)) + ((!n_n4317) & (n_n4362) & (n_n4319) & (!n_n4336)) + ((!n_n4317) & (n_n4362) & (n_n4319) & (n_n4336)) + ((n_n4317) & (!n_n4362) & (!n_n4319) & (!n_n4336)) + ((n_n4317) & (!n_n4362) & (!n_n4319) & (n_n4336)) + ((n_n4317) & (!n_n4362) & (n_n4319) & (!n_n4336)) + ((n_n4317) & (!n_n4362) & (n_n4319) & (n_n4336)) + ((n_n4317) & (n_n4362) & (!n_n4319) & (!n_n4336)) + ((n_n4317) & (n_n4362) & (!n_n4319) & (n_n4336)) + ((n_n4317) & (n_n4362) & (n_n4319) & (!n_n4336)) + ((n_n4317) & (n_n4362) & (n_n4319) & (n_n4336)));
	assign x14291x = (((!n_n4324) & (!n_n4314) & (!n_n4321) & (!n_n4348) & (n_n4355)) + ((!n_n4324) & (!n_n4314) & (!n_n4321) & (n_n4348) & (!n_n4355)) + ((!n_n4324) & (!n_n4314) & (!n_n4321) & (n_n4348) & (n_n4355)) + ((!n_n4324) & (!n_n4314) & (n_n4321) & (!n_n4348) & (!n_n4355)) + ((!n_n4324) & (!n_n4314) & (n_n4321) & (!n_n4348) & (n_n4355)) + ((!n_n4324) & (!n_n4314) & (n_n4321) & (n_n4348) & (!n_n4355)) + ((!n_n4324) & (!n_n4314) & (n_n4321) & (n_n4348) & (n_n4355)) + ((!n_n4324) & (n_n4314) & (!n_n4321) & (!n_n4348) & (!n_n4355)) + ((!n_n4324) & (n_n4314) & (!n_n4321) & (!n_n4348) & (n_n4355)) + ((!n_n4324) & (n_n4314) & (!n_n4321) & (n_n4348) & (!n_n4355)) + ((!n_n4324) & (n_n4314) & (!n_n4321) & (n_n4348) & (n_n4355)) + ((!n_n4324) & (n_n4314) & (n_n4321) & (!n_n4348) & (!n_n4355)) + ((!n_n4324) & (n_n4314) & (n_n4321) & (!n_n4348) & (n_n4355)) + ((!n_n4324) & (n_n4314) & (n_n4321) & (n_n4348) & (!n_n4355)) + ((!n_n4324) & (n_n4314) & (n_n4321) & (n_n4348) & (n_n4355)) + ((n_n4324) & (!n_n4314) & (!n_n4321) & (!n_n4348) & (!n_n4355)) + ((n_n4324) & (!n_n4314) & (!n_n4321) & (!n_n4348) & (n_n4355)) + ((n_n4324) & (!n_n4314) & (!n_n4321) & (n_n4348) & (!n_n4355)) + ((n_n4324) & (!n_n4314) & (!n_n4321) & (n_n4348) & (n_n4355)) + ((n_n4324) & (!n_n4314) & (n_n4321) & (!n_n4348) & (!n_n4355)) + ((n_n4324) & (!n_n4314) & (n_n4321) & (!n_n4348) & (n_n4355)) + ((n_n4324) & (!n_n4314) & (n_n4321) & (n_n4348) & (!n_n4355)) + ((n_n4324) & (!n_n4314) & (n_n4321) & (n_n4348) & (n_n4355)) + ((n_n4324) & (n_n4314) & (!n_n4321) & (!n_n4348) & (!n_n4355)) + ((n_n4324) & (n_n4314) & (!n_n4321) & (!n_n4348) & (n_n4355)) + ((n_n4324) & (n_n4314) & (!n_n4321) & (n_n4348) & (!n_n4355)) + ((n_n4324) & (n_n4314) & (!n_n4321) & (n_n4348) & (n_n4355)) + ((n_n4324) & (n_n4314) & (n_n4321) & (!n_n4348) & (!n_n4355)) + ((n_n4324) & (n_n4314) & (n_n4321) & (!n_n4348) & (n_n4355)) + ((n_n4324) & (n_n4314) & (n_n4321) & (n_n4348) & (!n_n4355)) + ((n_n4324) & (n_n4314) & (n_n4321) & (n_n4348) & (n_n4355)));
	assign n_n3562 = (((!n_n4617) & (!n_n4637) & (!n_n4638) & (!n_n4626) & (x14296x)) + ((!n_n4617) & (!n_n4637) & (!n_n4638) & (n_n4626) & (!x14296x)) + ((!n_n4617) & (!n_n4637) & (!n_n4638) & (n_n4626) & (x14296x)) + ((!n_n4617) & (!n_n4637) & (n_n4638) & (!n_n4626) & (!x14296x)) + ((!n_n4617) & (!n_n4637) & (n_n4638) & (!n_n4626) & (x14296x)) + ((!n_n4617) & (!n_n4637) & (n_n4638) & (n_n4626) & (!x14296x)) + ((!n_n4617) & (!n_n4637) & (n_n4638) & (n_n4626) & (x14296x)) + ((!n_n4617) & (n_n4637) & (!n_n4638) & (!n_n4626) & (!x14296x)) + ((!n_n4617) & (n_n4637) & (!n_n4638) & (!n_n4626) & (x14296x)) + ((!n_n4617) & (n_n4637) & (!n_n4638) & (n_n4626) & (!x14296x)) + ((!n_n4617) & (n_n4637) & (!n_n4638) & (n_n4626) & (x14296x)) + ((!n_n4617) & (n_n4637) & (n_n4638) & (!n_n4626) & (!x14296x)) + ((!n_n4617) & (n_n4637) & (n_n4638) & (!n_n4626) & (x14296x)) + ((!n_n4617) & (n_n4637) & (n_n4638) & (n_n4626) & (!x14296x)) + ((!n_n4617) & (n_n4637) & (n_n4638) & (n_n4626) & (x14296x)) + ((n_n4617) & (!n_n4637) & (!n_n4638) & (!n_n4626) & (!x14296x)) + ((n_n4617) & (!n_n4637) & (!n_n4638) & (!n_n4626) & (x14296x)) + ((n_n4617) & (!n_n4637) & (!n_n4638) & (n_n4626) & (!x14296x)) + ((n_n4617) & (!n_n4637) & (!n_n4638) & (n_n4626) & (x14296x)) + ((n_n4617) & (!n_n4637) & (n_n4638) & (!n_n4626) & (!x14296x)) + ((n_n4617) & (!n_n4637) & (n_n4638) & (!n_n4626) & (x14296x)) + ((n_n4617) & (!n_n4637) & (n_n4638) & (n_n4626) & (!x14296x)) + ((n_n4617) & (!n_n4637) & (n_n4638) & (n_n4626) & (x14296x)) + ((n_n4617) & (n_n4637) & (!n_n4638) & (!n_n4626) & (!x14296x)) + ((n_n4617) & (n_n4637) & (!n_n4638) & (!n_n4626) & (x14296x)) + ((n_n4617) & (n_n4637) & (!n_n4638) & (n_n4626) & (!x14296x)) + ((n_n4617) & (n_n4637) & (!n_n4638) & (n_n4626) & (x14296x)) + ((n_n4617) & (n_n4637) & (n_n4638) & (!n_n4626) & (!x14296x)) + ((n_n4617) & (n_n4637) & (n_n4638) & (!n_n4626) & (x14296x)) + ((n_n4617) & (n_n4637) & (n_n4638) & (n_n4626) & (!x14296x)) + ((n_n4617) & (n_n4637) & (n_n4638) & (n_n4626) & (x14296x)));
	assign x14301x = (((!n_n4514) & (!n_n4544) & (!n_n4561) & (n_n4522)) + ((!n_n4514) & (!n_n4544) & (n_n4561) & (!n_n4522)) + ((!n_n4514) & (!n_n4544) & (n_n4561) & (n_n4522)) + ((!n_n4514) & (n_n4544) & (!n_n4561) & (!n_n4522)) + ((!n_n4514) & (n_n4544) & (!n_n4561) & (n_n4522)) + ((!n_n4514) & (n_n4544) & (n_n4561) & (!n_n4522)) + ((!n_n4514) & (n_n4544) & (n_n4561) & (n_n4522)) + ((n_n4514) & (!n_n4544) & (!n_n4561) & (!n_n4522)) + ((n_n4514) & (!n_n4544) & (!n_n4561) & (n_n4522)) + ((n_n4514) & (!n_n4544) & (n_n4561) & (!n_n4522)) + ((n_n4514) & (!n_n4544) & (n_n4561) & (n_n4522)) + ((n_n4514) & (n_n4544) & (!n_n4561) & (!n_n4522)) + ((n_n4514) & (n_n4544) & (!n_n4561) & (n_n4522)) + ((n_n4514) & (n_n4544) & (n_n4561) & (!n_n4522)) + ((n_n4514) & (n_n4544) & (n_n4561) & (n_n4522)));
	assign x14302x = (((!n_n4525) & (!n_n4542) & (!n_n4498) & (!n_n4499) & (n_n4559)) + ((!n_n4525) & (!n_n4542) & (!n_n4498) & (n_n4499) & (!n_n4559)) + ((!n_n4525) & (!n_n4542) & (!n_n4498) & (n_n4499) & (n_n4559)) + ((!n_n4525) & (!n_n4542) & (n_n4498) & (!n_n4499) & (!n_n4559)) + ((!n_n4525) & (!n_n4542) & (n_n4498) & (!n_n4499) & (n_n4559)) + ((!n_n4525) & (!n_n4542) & (n_n4498) & (n_n4499) & (!n_n4559)) + ((!n_n4525) & (!n_n4542) & (n_n4498) & (n_n4499) & (n_n4559)) + ((!n_n4525) & (n_n4542) & (!n_n4498) & (!n_n4499) & (!n_n4559)) + ((!n_n4525) & (n_n4542) & (!n_n4498) & (!n_n4499) & (n_n4559)) + ((!n_n4525) & (n_n4542) & (!n_n4498) & (n_n4499) & (!n_n4559)) + ((!n_n4525) & (n_n4542) & (!n_n4498) & (n_n4499) & (n_n4559)) + ((!n_n4525) & (n_n4542) & (n_n4498) & (!n_n4499) & (!n_n4559)) + ((!n_n4525) & (n_n4542) & (n_n4498) & (!n_n4499) & (n_n4559)) + ((!n_n4525) & (n_n4542) & (n_n4498) & (n_n4499) & (!n_n4559)) + ((!n_n4525) & (n_n4542) & (n_n4498) & (n_n4499) & (n_n4559)) + ((n_n4525) & (!n_n4542) & (!n_n4498) & (!n_n4499) & (!n_n4559)) + ((n_n4525) & (!n_n4542) & (!n_n4498) & (!n_n4499) & (n_n4559)) + ((n_n4525) & (!n_n4542) & (!n_n4498) & (n_n4499) & (!n_n4559)) + ((n_n4525) & (!n_n4542) & (!n_n4498) & (n_n4499) & (n_n4559)) + ((n_n4525) & (!n_n4542) & (n_n4498) & (!n_n4499) & (!n_n4559)) + ((n_n4525) & (!n_n4542) & (n_n4498) & (!n_n4499) & (n_n4559)) + ((n_n4525) & (!n_n4542) & (n_n4498) & (n_n4499) & (!n_n4559)) + ((n_n4525) & (!n_n4542) & (n_n4498) & (n_n4499) & (n_n4559)) + ((n_n4525) & (n_n4542) & (!n_n4498) & (!n_n4499) & (!n_n4559)) + ((n_n4525) & (n_n4542) & (!n_n4498) & (!n_n4499) & (n_n4559)) + ((n_n4525) & (n_n4542) & (!n_n4498) & (n_n4499) & (!n_n4559)) + ((n_n4525) & (n_n4542) & (!n_n4498) & (n_n4499) & (n_n4559)) + ((n_n4525) & (n_n4542) & (n_n4498) & (!n_n4499) & (!n_n4559)) + ((n_n4525) & (n_n4542) & (n_n4498) & (!n_n4499) & (n_n4559)) + ((n_n4525) & (n_n4542) & (n_n4498) & (n_n4499) & (!n_n4559)) + ((n_n4525) & (n_n4542) & (n_n4498) & (n_n4499) & (n_n4559)));
	assign x14308x = (((!n_n4568) & (!n_n4590) & (!n_n4582) & (n_n4581)) + ((!n_n4568) & (!n_n4590) & (n_n4582) & (!n_n4581)) + ((!n_n4568) & (!n_n4590) & (n_n4582) & (n_n4581)) + ((!n_n4568) & (n_n4590) & (!n_n4582) & (!n_n4581)) + ((!n_n4568) & (n_n4590) & (!n_n4582) & (n_n4581)) + ((!n_n4568) & (n_n4590) & (n_n4582) & (!n_n4581)) + ((!n_n4568) & (n_n4590) & (n_n4582) & (n_n4581)) + ((n_n4568) & (!n_n4590) & (!n_n4582) & (!n_n4581)) + ((n_n4568) & (!n_n4590) & (!n_n4582) & (n_n4581)) + ((n_n4568) & (!n_n4590) & (n_n4582) & (!n_n4581)) + ((n_n4568) & (!n_n4590) & (n_n4582) & (n_n4581)) + ((n_n4568) & (n_n4590) & (!n_n4582) & (!n_n4581)) + ((n_n4568) & (n_n4590) & (!n_n4582) & (n_n4581)) + ((n_n4568) & (n_n4590) & (n_n4582) & (!n_n4581)) + ((n_n4568) & (n_n4590) & (n_n4582) & (n_n4581)));
	assign x14309x = (((!n_n4602) & (!n_n4601) & (!n_n4595) & (!n_n4608) & (n_n4579)) + ((!n_n4602) & (!n_n4601) & (!n_n4595) & (n_n4608) & (!n_n4579)) + ((!n_n4602) & (!n_n4601) & (!n_n4595) & (n_n4608) & (n_n4579)) + ((!n_n4602) & (!n_n4601) & (n_n4595) & (!n_n4608) & (!n_n4579)) + ((!n_n4602) & (!n_n4601) & (n_n4595) & (!n_n4608) & (n_n4579)) + ((!n_n4602) & (!n_n4601) & (n_n4595) & (n_n4608) & (!n_n4579)) + ((!n_n4602) & (!n_n4601) & (n_n4595) & (n_n4608) & (n_n4579)) + ((!n_n4602) & (n_n4601) & (!n_n4595) & (!n_n4608) & (!n_n4579)) + ((!n_n4602) & (n_n4601) & (!n_n4595) & (!n_n4608) & (n_n4579)) + ((!n_n4602) & (n_n4601) & (!n_n4595) & (n_n4608) & (!n_n4579)) + ((!n_n4602) & (n_n4601) & (!n_n4595) & (n_n4608) & (n_n4579)) + ((!n_n4602) & (n_n4601) & (n_n4595) & (!n_n4608) & (!n_n4579)) + ((!n_n4602) & (n_n4601) & (n_n4595) & (!n_n4608) & (n_n4579)) + ((!n_n4602) & (n_n4601) & (n_n4595) & (n_n4608) & (!n_n4579)) + ((!n_n4602) & (n_n4601) & (n_n4595) & (n_n4608) & (n_n4579)) + ((n_n4602) & (!n_n4601) & (!n_n4595) & (!n_n4608) & (!n_n4579)) + ((n_n4602) & (!n_n4601) & (!n_n4595) & (!n_n4608) & (n_n4579)) + ((n_n4602) & (!n_n4601) & (!n_n4595) & (n_n4608) & (!n_n4579)) + ((n_n4602) & (!n_n4601) & (!n_n4595) & (n_n4608) & (n_n4579)) + ((n_n4602) & (!n_n4601) & (n_n4595) & (!n_n4608) & (!n_n4579)) + ((n_n4602) & (!n_n4601) & (n_n4595) & (!n_n4608) & (n_n4579)) + ((n_n4602) & (!n_n4601) & (n_n4595) & (n_n4608) & (!n_n4579)) + ((n_n4602) & (!n_n4601) & (n_n4595) & (n_n4608) & (n_n4579)) + ((n_n4602) & (n_n4601) & (!n_n4595) & (!n_n4608) & (!n_n4579)) + ((n_n4602) & (n_n4601) & (!n_n4595) & (!n_n4608) & (n_n4579)) + ((n_n4602) & (n_n4601) & (!n_n4595) & (n_n4608) & (!n_n4579)) + ((n_n4602) & (n_n4601) & (!n_n4595) & (n_n4608) & (n_n4579)) + ((n_n4602) & (n_n4601) & (n_n4595) & (!n_n4608) & (!n_n4579)) + ((n_n4602) & (n_n4601) & (n_n4595) & (!n_n4608) & (n_n4579)) + ((n_n4602) & (n_n4601) & (n_n4595) & (n_n4608) & (!n_n4579)) + ((n_n4602) & (n_n4601) & (n_n4595) & (n_n4608) & (n_n4579)));
	assign x14331x = (((!n_n4784) & (!n_n4747) & (!n_n4787) & (!n_n4780) & (n_n4752)) + ((!n_n4784) & (!n_n4747) & (!n_n4787) & (n_n4780) & (!n_n4752)) + ((!n_n4784) & (!n_n4747) & (!n_n4787) & (n_n4780) & (n_n4752)) + ((!n_n4784) & (!n_n4747) & (n_n4787) & (!n_n4780) & (!n_n4752)) + ((!n_n4784) & (!n_n4747) & (n_n4787) & (!n_n4780) & (n_n4752)) + ((!n_n4784) & (!n_n4747) & (n_n4787) & (n_n4780) & (!n_n4752)) + ((!n_n4784) & (!n_n4747) & (n_n4787) & (n_n4780) & (n_n4752)) + ((!n_n4784) & (n_n4747) & (!n_n4787) & (!n_n4780) & (!n_n4752)) + ((!n_n4784) & (n_n4747) & (!n_n4787) & (!n_n4780) & (n_n4752)) + ((!n_n4784) & (n_n4747) & (!n_n4787) & (n_n4780) & (!n_n4752)) + ((!n_n4784) & (n_n4747) & (!n_n4787) & (n_n4780) & (n_n4752)) + ((!n_n4784) & (n_n4747) & (n_n4787) & (!n_n4780) & (!n_n4752)) + ((!n_n4784) & (n_n4747) & (n_n4787) & (!n_n4780) & (n_n4752)) + ((!n_n4784) & (n_n4747) & (n_n4787) & (n_n4780) & (!n_n4752)) + ((!n_n4784) & (n_n4747) & (n_n4787) & (n_n4780) & (n_n4752)) + ((n_n4784) & (!n_n4747) & (!n_n4787) & (!n_n4780) & (!n_n4752)) + ((n_n4784) & (!n_n4747) & (!n_n4787) & (!n_n4780) & (n_n4752)) + ((n_n4784) & (!n_n4747) & (!n_n4787) & (n_n4780) & (!n_n4752)) + ((n_n4784) & (!n_n4747) & (!n_n4787) & (n_n4780) & (n_n4752)) + ((n_n4784) & (!n_n4747) & (n_n4787) & (!n_n4780) & (!n_n4752)) + ((n_n4784) & (!n_n4747) & (n_n4787) & (!n_n4780) & (n_n4752)) + ((n_n4784) & (!n_n4747) & (n_n4787) & (n_n4780) & (!n_n4752)) + ((n_n4784) & (!n_n4747) & (n_n4787) & (n_n4780) & (n_n4752)) + ((n_n4784) & (n_n4747) & (!n_n4787) & (!n_n4780) & (!n_n4752)) + ((n_n4784) & (n_n4747) & (!n_n4787) & (!n_n4780) & (n_n4752)) + ((n_n4784) & (n_n4747) & (!n_n4787) & (n_n4780) & (!n_n4752)) + ((n_n4784) & (n_n4747) & (!n_n4787) & (n_n4780) & (n_n4752)) + ((n_n4784) & (n_n4747) & (n_n4787) & (!n_n4780) & (!n_n4752)) + ((n_n4784) & (n_n4747) & (n_n4787) & (!n_n4780) & (n_n4752)) + ((n_n4784) & (n_n4747) & (n_n4787) & (n_n4780) & (!n_n4752)) + ((n_n4784) & (n_n4747) & (n_n4787) & (n_n4780) & (n_n4752)));
	assign x14317x = (((!x483x) & (!x20x) & (!n_n4717) & (!n_n4703) & (n_n4736)) + ((!x483x) & (!x20x) & (!n_n4717) & (n_n4703) & (!n_n4736)) + ((!x483x) & (!x20x) & (!n_n4717) & (n_n4703) & (n_n4736)) + ((!x483x) & (!x20x) & (n_n4717) & (!n_n4703) & (!n_n4736)) + ((!x483x) & (!x20x) & (n_n4717) & (!n_n4703) & (n_n4736)) + ((!x483x) & (!x20x) & (n_n4717) & (n_n4703) & (!n_n4736)) + ((!x483x) & (!x20x) & (n_n4717) & (n_n4703) & (n_n4736)) + ((!x483x) & (x20x) & (!n_n4717) & (!n_n4703) & (n_n4736)) + ((!x483x) & (x20x) & (!n_n4717) & (n_n4703) & (!n_n4736)) + ((!x483x) & (x20x) & (!n_n4717) & (n_n4703) & (n_n4736)) + ((!x483x) & (x20x) & (n_n4717) & (!n_n4703) & (!n_n4736)) + ((!x483x) & (x20x) & (n_n4717) & (!n_n4703) & (n_n4736)) + ((!x483x) & (x20x) & (n_n4717) & (n_n4703) & (!n_n4736)) + ((!x483x) & (x20x) & (n_n4717) & (n_n4703) & (n_n4736)) + ((x483x) & (!x20x) & (!n_n4717) & (!n_n4703) & (n_n4736)) + ((x483x) & (!x20x) & (!n_n4717) & (n_n4703) & (!n_n4736)) + ((x483x) & (!x20x) & (!n_n4717) & (n_n4703) & (n_n4736)) + ((x483x) & (!x20x) & (n_n4717) & (!n_n4703) & (!n_n4736)) + ((x483x) & (!x20x) & (n_n4717) & (!n_n4703) & (n_n4736)) + ((x483x) & (!x20x) & (n_n4717) & (n_n4703) & (!n_n4736)) + ((x483x) & (!x20x) & (n_n4717) & (n_n4703) & (n_n4736)) + ((x483x) & (x20x) & (!n_n4717) & (!n_n4703) & (!n_n4736)) + ((x483x) & (x20x) & (!n_n4717) & (!n_n4703) & (n_n4736)) + ((x483x) & (x20x) & (!n_n4717) & (n_n4703) & (!n_n4736)) + ((x483x) & (x20x) & (!n_n4717) & (n_n4703) & (n_n4736)) + ((x483x) & (x20x) & (n_n4717) & (!n_n4703) & (!n_n4736)) + ((x483x) & (x20x) & (n_n4717) & (!n_n4703) & (n_n4736)) + ((x483x) & (x20x) & (n_n4717) & (n_n4703) & (!n_n4736)) + ((x483x) & (x20x) & (n_n4717) & (n_n4703) & (n_n4736)));
	assign x14318x = (((!n_n4744) & (!n_n4697) & (!n_n4708) & (!n_n4695) & (n_n4721)) + ((!n_n4744) & (!n_n4697) & (!n_n4708) & (n_n4695) & (!n_n4721)) + ((!n_n4744) & (!n_n4697) & (!n_n4708) & (n_n4695) & (n_n4721)) + ((!n_n4744) & (!n_n4697) & (n_n4708) & (!n_n4695) & (!n_n4721)) + ((!n_n4744) & (!n_n4697) & (n_n4708) & (!n_n4695) & (n_n4721)) + ((!n_n4744) & (!n_n4697) & (n_n4708) & (n_n4695) & (!n_n4721)) + ((!n_n4744) & (!n_n4697) & (n_n4708) & (n_n4695) & (n_n4721)) + ((!n_n4744) & (n_n4697) & (!n_n4708) & (!n_n4695) & (!n_n4721)) + ((!n_n4744) & (n_n4697) & (!n_n4708) & (!n_n4695) & (n_n4721)) + ((!n_n4744) & (n_n4697) & (!n_n4708) & (n_n4695) & (!n_n4721)) + ((!n_n4744) & (n_n4697) & (!n_n4708) & (n_n4695) & (n_n4721)) + ((!n_n4744) & (n_n4697) & (n_n4708) & (!n_n4695) & (!n_n4721)) + ((!n_n4744) & (n_n4697) & (n_n4708) & (!n_n4695) & (n_n4721)) + ((!n_n4744) & (n_n4697) & (n_n4708) & (n_n4695) & (!n_n4721)) + ((!n_n4744) & (n_n4697) & (n_n4708) & (n_n4695) & (n_n4721)) + ((n_n4744) & (!n_n4697) & (!n_n4708) & (!n_n4695) & (!n_n4721)) + ((n_n4744) & (!n_n4697) & (!n_n4708) & (!n_n4695) & (n_n4721)) + ((n_n4744) & (!n_n4697) & (!n_n4708) & (n_n4695) & (!n_n4721)) + ((n_n4744) & (!n_n4697) & (!n_n4708) & (n_n4695) & (n_n4721)) + ((n_n4744) & (!n_n4697) & (n_n4708) & (!n_n4695) & (!n_n4721)) + ((n_n4744) & (!n_n4697) & (n_n4708) & (!n_n4695) & (n_n4721)) + ((n_n4744) & (!n_n4697) & (n_n4708) & (n_n4695) & (!n_n4721)) + ((n_n4744) & (!n_n4697) & (n_n4708) & (n_n4695) & (n_n4721)) + ((n_n4744) & (n_n4697) & (!n_n4708) & (!n_n4695) & (!n_n4721)) + ((n_n4744) & (n_n4697) & (!n_n4708) & (!n_n4695) & (n_n4721)) + ((n_n4744) & (n_n4697) & (!n_n4708) & (n_n4695) & (!n_n4721)) + ((n_n4744) & (n_n4697) & (!n_n4708) & (n_n4695) & (n_n4721)) + ((n_n4744) & (n_n4697) & (n_n4708) & (!n_n4695) & (!n_n4721)) + ((n_n4744) & (n_n4697) & (n_n4708) & (!n_n4695) & (n_n4721)) + ((n_n4744) & (n_n4697) & (n_n4708) & (n_n4695) & (!n_n4721)) + ((n_n4744) & (n_n4697) & (n_n4708) & (n_n4695) & (n_n4721)));
	assign x14323x = (((!n_n4646) & (!n_n4668) & (!n_n4670) & (n_n4678)) + ((!n_n4646) & (!n_n4668) & (n_n4670) & (!n_n4678)) + ((!n_n4646) & (!n_n4668) & (n_n4670) & (n_n4678)) + ((!n_n4646) & (n_n4668) & (!n_n4670) & (!n_n4678)) + ((!n_n4646) & (n_n4668) & (!n_n4670) & (n_n4678)) + ((!n_n4646) & (n_n4668) & (n_n4670) & (!n_n4678)) + ((!n_n4646) & (n_n4668) & (n_n4670) & (n_n4678)) + ((n_n4646) & (!n_n4668) & (!n_n4670) & (!n_n4678)) + ((n_n4646) & (!n_n4668) & (!n_n4670) & (n_n4678)) + ((n_n4646) & (!n_n4668) & (n_n4670) & (!n_n4678)) + ((n_n4646) & (!n_n4668) & (n_n4670) & (n_n4678)) + ((n_n4646) & (n_n4668) & (!n_n4670) & (!n_n4678)) + ((n_n4646) & (n_n4668) & (!n_n4670) & (n_n4678)) + ((n_n4646) & (n_n4668) & (n_n4670) & (!n_n4678)) + ((n_n4646) & (n_n4668) & (n_n4670) & (n_n4678)));
	assign x14324x = (((!n_n4660) & (!n_n4665) & (!x312x) & (n_n4687)) + ((!n_n4660) & (!n_n4665) & (x312x) & (!n_n4687)) + ((!n_n4660) & (!n_n4665) & (x312x) & (n_n4687)) + ((!n_n4660) & (n_n4665) & (!x312x) & (!n_n4687)) + ((!n_n4660) & (n_n4665) & (!x312x) & (n_n4687)) + ((!n_n4660) & (n_n4665) & (x312x) & (!n_n4687)) + ((!n_n4660) & (n_n4665) & (x312x) & (n_n4687)) + ((n_n4660) & (!n_n4665) & (!x312x) & (!n_n4687)) + ((n_n4660) & (!n_n4665) & (!x312x) & (n_n4687)) + ((n_n4660) & (!n_n4665) & (x312x) & (!n_n4687)) + ((n_n4660) & (!n_n4665) & (x312x) & (n_n4687)) + ((n_n4660) & (n_n4665) & (!x312x) & (!n_n4687)) + ((n_n4660) & (n_n4665) & (!x312x) & (n_n4687)) + ((n_n4660) & (n_n4665) & (x312x) & (!n_n4687)) + ((n_n4660) & (n_n4665) & (x312x) & (n_n4687)));
	assign n_n5158 = (((i_5_) & (!i_3_) & (i_4_) & (n_n520) & (x12x)));
	assign n_n5154 = (((i_7_) & (!i_8_) & (!i_6_) & (n_n491) & (x12x)));
	assign n_n5013 = (((i_1_) & (!i_2_) & (!i_0_) & (x20x) & (n_n500)));
	assign n_n3427 = (((!i_9_) & (n_n522) & (!n_n520) & (n_n195) & (n_n500)) + ((!i_9_) & (n_n522) & (n_n520) & (n_n195) & (n_n500)) + ((i_9_) & (!n_n522) & (n_n520) & (n_n195) & (n_n500)) + ((i_9_) & (n_n522) & (!n_n520) & (n_n195) & (n_n500)) + ((i_9_) & (n_n522) & (n_n520) & (n_n195) & (n_n500)));
	assign n_n5150 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n491) & (x12x)));
	assign n_n5147 = (((!i_9_) & (n_n532) & (n_n491) & (n_n130)));
	assign n_n5149 = (((!i_9_) & (n_n491) & (n_n130) & (n_n530)));
	assign n_n5148 = (((i_5_) & (!i_3_) & (i_4_) & (x12x) & (n_n530)));
	assign x76x = (((!i_9_) & (n_n491) & (!n_n130) & (x12x) & (n_n530)) + ((!i_9_) & (n_n491) & (n_n130) & (!x12x) & (n_n530)) + ((!i_9_) & (n_n491) & (n_n130) & (x12x) & (n_n530)) + ((i_9_) & (n_n491) & (!n_n130) & (x12x) & (n_n530)) + ((i_9_) & (n_n491) & (n_n130) & (x12x) & (n_n530)));
	assign n_n5152 = (((i_7_) & (i_8_) & (!i_6_) & (n_n491) & (x12x)));
	assign n_n5153 = (((!i_9_) & (n_n526) & (n_n491) & (n_n130)));
	assign x196x = (((!i_9_) & (n_n526) & (n_n491) & (!n_n130) & (x12x)) + ((!i_9_) & (n_n526) & (n_n491) & (n_n130) & (!x12x)) + ((!i_9_) & (n_n526) & (n_n491) & (n_n130) & (x12x)) + ((i_9_) & (n_n526) & (n_n491) & (!n_n130) & (x12x)) + ((i_9_) & (n_n526) & (n_n491) & (n_n130) & (x12x)));
	assign x22115x = (((!n_n5157) & (!n_n5158) & (!n_n5154) & (!n_n5150)));
	assign n_n3305 = (((!n_n5147) & (!n_n5149) & (!n_n5148) & (!x196x) & (!x22115x)) + ((!n_n5147) & (!n_n5149) & (!n_n5148) & (x196x) & (!x22115x)) + ((!n_n5147) & (!n_n5149) & (!n_n5148) & (x196x) & (x22115x)) + ((!n_n5147) & (!n_n5149) & (n_n5148) & (!x196x) & (!x22115x)) + ((!n_n5147) & (!n_n5149) & (n_n5148) & (!x196x) & (x22115x)) + ((!n_n5147) & (!n_n5149) & (n_n5148) & (x196x) & (!x22115x)) + ((!n_n5147) & (!n_n5149) & (n_n5148) & (x196x) & (x22115x)) + ((!n_n5147) & (n_n5149) & (!n_n5148) & (!x196x) & (!x22115x)) + ((!n_n5147) & (n_n5149) & (!n_n5148) & (!x196x) & (x22115x)) + ((!n_n5147) & (n_n5149) & (!n_n5148) & (x196x) & (!x22115x)) + ((!n_n5147) & (n_n5149) & (!n_n5148) & (x196x) & (x22115x)) + ((!n_n5147) & (n_n5149) & (n_n5148) & (!x196x) & (!x22115x)) + ((!n_n5147) & (n_n5149) & (n_n5148) & (!x196x) & (x22115x)) + ((!n_n5147) & (n_n5149) & (n_n5148) & (x196x) & (!x22115x)) + ((!n_n5147) & (n_n5149) & (n_n5148) & (x196x) & (x22115x)) + ((n_n5147) & (!n_n5149) & (!n_n5148) & (!x196x) & (!x22115x)) + ((n_n5147) & (!n_n5149) & (!n_n5148) & (!x196x) & (x22115x)) + ((n_n5147) & (!n_n5149) & (!n_n5148) & (x196x) & (!x22115x)) + ((n_n5147) & (!n_n5149) & (!n_n5148) & (x196x) & (x22115x)) + ((n_n5147) & (!n_n5149) & (n_n5148) & (!x196x) & (!x22115x)) + ((n_n5147) & (!n_n5149) & (n_n5148) & (!x196x) & (x22115x)) + ((n_n5147) & (!n_n5149) & (n_n5148) & (x196x) & (!x22115x)) + ((n_n5147) & (!n_n5149) & (n_n5148) & (x196x) & (x22115x)) + ((n_n5147) & (n_n5149) & (!n_n5148) & (!x196x) & (!x22115x)) + ((n_n5147) & (n_n5149) & (!n_n5148) & (!x196x) & (x22115x)) + ((n_n5147) & (n_n5149) & (!n_n5148) & (x196x) & (!x22115x)) + ((n_n5147) & (n_n5149) & (!n_n5148) & (x196x) & (x22115x)) + ((n_n5147) & (n_n5149) & (n_n5148) & (!x196x) & (!x22115x)) + ((n_n5147) & (n_n5149) & (n_n5148) & (!x196x) & (x22115x)) + ((n_n5147) & (n_n5149) & (n_n5148) & (x196x) & (!x22115x)) + ((n_n5147) & (n_n5149) & (n_n5148) & (x196x) & (x22115x)));
	assign x13834x = (((!n_n4988) & (!n_n4979) & (!n_n4985) & (!n_n4984) & (n_n4978)) + ((!n_n4988) & (!n_n4979) & (!n_n4985) & (n_n4984) & (!n_n4978)) + ((!n_n4988) & (!n_n4979) & (!n_n4985) & (n_n4984) & (n_n4978)) + ((!n_n4988) & (!n_n4979) & (n_n4985) & (!n_n4984) & (!n_n4978)) + ((!n_n4988) & (!n_n4979) & (n_n4985) & (!n_n4984) & (n_n4978)) + ((!n_n4988) & (!n_n4979) & (n_n4985) & (n_n4984) & (!n_n4978)) + ((!n_n4988) & (!n_n4979) & (n_n4985) & (n_n4984) & (n_n4978)) + ((!n_n4988) & (n_n4979) & (!n_n4985) & (!n_n4984) & (!n_n4978)) + ((!n_n4988) & (n_n4979) & (!n_n4985) & (!n_n4984) & (n_n4978)) + ((!n_n4988) & (n_n4979) & (!n_n4985) & (n_n4984) & (!n_n4978)) + ((!n_n4988) & (n_n4979) & (!n_n4985) & (n_n4984) & (n_n4978)) + ((!n_n4988) & (n_n4979) & (n_n4985) & (!n_n4984) & (!n_n4978)) + ((!n_n4988) & (n_n4979) & (n_n4985) & (!n_n4984) & (n_n4978)) + ((!n_n4988) & (n_n4979) & (n_n4985) & (n_n4984) & (!n_n4978)) + ((!n_n4988) & (n_n4979) & (n_n4985) & (n_n4984) & (n_n4978)) + ((n_n4988) & (!n_n4979) & (!n_n4985) & (!n_n4984) & (!n_n4978)) + ((n_n4988) & (!n_n4979) & (!n_n4985) & (!n_n4984) & (n_n4978)) + ((n_n4988) & (!n_n4979) & (!n_n4985) & (n_n4984) & (!n_n4978)) + ((n_n4988) & (!n_n4979) & (!n_n4985) & (n_n4984) & (n_n4978)) + ((n_n4988) & (!n_n4979) & (n_n4985) & (!n_n4984) & (!n_n4978)) + ((n_n4988) & (!n_n4979) & (n_n4985) & (!n_n4984) & (n_n4978)) + ((n_n4988) & (!n_n4979) & (n_n4985) & (n_n4984) & (!n_n4978)) + ((n_n4988) & (!n_n4979) & (n_n4985) & (n_n4984) & (n_n4978)) + ((n_n4988) & (n_n4979) & (!n_n4985) & (!n_n4984) & (!n_n4978)) + ((n_n4988) & (n_n4979) & (!n_n4985) & (!n_n4984) & (n_n4978)) + ((n_n4988) & (n_n4979) & (!n_n4985) & (n_n4984) & (!n_n4978)) + ((n_n4988) & (n_n4979) & (!n_n4985) & (n_n4984) & (n_n4978)) + ((n_n4988) & (n_n4979) & (n_n4985) & (!n_n4984) & (!n_n4978)) + ((n_n4988) & (n_n4979) & (n_n4985) & (!n_n4984) & (n_n4978)) + ((n_n4988) & (n_n4979) & (n_n4985) & (n_n4984) & (!n_n4978)) + ((n_n4988) & (n_n4979) & (n_n4985) & (n_n4984) & (n_n4978)));
	assign n_n3318 = (((!n_n4976) & (!n_n4982) & (!n_n4983) & (!n_n4981) & (x13834x)) + ((!n_n4976) & (!n_n4982) & (!n_n4983) & (n_n4981) & (!x13834x)) + ((!n_n4976) & (!n_n4982) & (!n_n4983) & (n_n4981) & (x13834x)) + ((!n_n4976) & (!n_n4982) & (n_n4983) & (!n_n4981) & (!x13834x)) + ((!n_n4976) & (!n_n4982) & (n_n4983) & (!n_n4981) & (x13834x)) + ((!n_n4976) & (!n_n4982) & (n_n4983) & (n_n4981) & (!x13834x)) + ((!n_n4976) & (!n_n4982) & (n_n4983) & (n_n4981) & (x13834x)) + ((!n_n4976) & (n_n4982) & (!n_n4983) & (!n_n4981) & (!x13834x)) + ((!n_n4976) & (n_n4982) & (!n_n4983) & (!n_n4981) & (x13834x)) + ((!n_n4976) & (n_n4982) & (!n_n4983) & (n_n4981) & (!x13834x)) + ((!n_n4976) & (n_n4982) & (!n_n4983) & (n_n4981) & (x13834x)) + ((!n_n4976) & (n_n4982) & (n_n4983) & (!n_n4981) & (!x13834x)) + ((!n_n4976) & (n_n4982) & (n_n4983) & (!n_n4981) & (x13834x)) + ((!n_n4976) & (n_n4982) & (n_n4983) & (n_n4981) & (!x13834x)) + ((!n_n4976) & (n_n4982) & (n_n4983) & (n_n4981) & (x13834x)) + ((n_n4976) & (!n_n4982) & (!n_n4983) & (!n_n4981) & (!x13834x)) + ((n_n4976) & (!n_n4982) & (!n_n4983) & (!n_n4981) & (x13834x)) + ((n_n4976) & (!n_n4982) & (!n_n4983) & (n_n4981) & (!x13834x)) + ((n_n4976) & (!n_n4982) & (!n_n4983) & (n_n4981) & (x13834x)) + ((n_n4976) & (!n_n4982) & (n_n4983) & (!n_n4981) & (!x13834x)) + ((n_n4976) & (!n_n4982) & (n_n4983) & (!n_n4981) & (x13834x)) + ((n_n4976) & (!n_n4982) & (n_n4983) & (n_n4981) & (!x13834x)) + ((n_n4976) & (!n_n4982) & (n_n4983) & (n_n4981) & (x13834x)) + ((n_n4976) & (n_n4982) & (!n_n4983) & (!n_n4981) & (!x13834x)) + ((n_n4976) & (n_n4982) & (!n_n4983) & (!n_n4981) & (x13834x)) + ((n_n4976) & (n_n4982) & (!n_n4983) & (n_n4981) & (!x13834x)) + ((n_n4976) & (n_n4982) & (!n_n4983) & (n_n4981) & (x13834x)) + ((n_n4976) & (n_n4982) & (n_n4983) & (!n_n4981) & (!x13834x)) + ((n_n4976) & (n_n4982) & (n_n4983) & (!n_n4981) & (x13834x)) + ((n_n4976) & (n_n4982) & (n_n4983) & (n_n4981) & (!x13834x)) + ((n_n4976) & (n_n4982) & (n_n4983) & (n_n4981) & (x13834x)));
	assign n_n4957 = (((!i_9_) & (n_n535) & (n_n195) & (n_n530)));
	assign n_n4172 = (((!i_9_) & (n_n535) & (n_n522) & (!n_n520) & (n_n195)) + ((!i_9_) & (n_n535) & (n_n522) & (n_n520) & (n_n195)) + ((i_9_) & (n_n535) & (!n_n522) & (n_n520) & (n_n195)) + ((i_9_) & (n_n535) & (n_n522) & (!n_n520) & (n_n195)) + ((i_9_) & (n_n535) & (n_n522) & (n_n520) & (n_n195)));
	assign x229x = (((!n_n4975) & (!n_n4968) & (!n_n4172) & (x68x)) + ((!n_n4975) & (!n_n4968) & (n_n4172) & (!x68x)) + ((!n_n4975) & (!n_n4968) & (n_n4172) & (x68x)) + ((!n_n4975) & (n_n4968) & (!n_n4172) & (!x68x)) + ((!n_n4975) & (n_n4968) & (!n_n4172) & (x68x)) + ((!n_n4975) & (n_n4968) & (n_n4172) & (!x68x)) + ((!n_n4975) & (n_n4968) & (n_n4172) & (x68x)) + ((n_n4975) & (!n_n4968) & (!n_n4172) & (!x68x)) + ((n_n4975) & (!n_n4968) & (!n_n4172) & (x68x)) + ((n_n4975) & (!n_n4968) & (n_n4172) & (!x68x)) + ((n_n4975) & (!n_n4968) & (n_n4172) & (x68x)) + ((n_n4975) & (n_n4968) & (!n_n4172) & (!x68x)) + ((n_n4975) & (n_n4968) & (!n_n4172) & (x68x)) + ((n_n4975) & (n_n4968) & (n_n4172) & (!x68x)) + ((n_n4975) & (n_n4968) & (n_n4172) & (x68x)));
	assign x13841x = (((!n_n4974) & (!n_n4948) & (!n_n4957) & (n_n4971)) + ((!n_n4974) & (!n_n4948) & (n_n4957) & (!n_n4971)) + ((!n_n4974) & (!n_n4948) & (n_n4957) & (n_n4971)) + ((!n_n4974) & (n_n4948) & (!n_n4957) & (!n_n4971)) + ((!n_n4974) & (n_n4948) & (!n_n4957) & (n_n4971)) + ((!n_n4974) & (n_n4948) & (n_n4957) & (!n_n4971)) + ((!n_n4974) & (n_n4948) & (n_n4957) & (n_n4971)) + ((n_n4974) & (!n_n4948) & (!n_n4957) & (!n_n4971)) + ((n_n4974) & (!n_n4948) & (!n_n4957) & (n_n4971)) + ((n_n4974) & (!n_n4948) & (n_n4957) & (!n_n4971)) + ((n_n4974) & (!n_n4948) & (n_n4957) & (n_n4971)) + ((n_n4974) & (n_n4948) & (!n_n4957) & (!n_n4971)) + ((n_n4974) & (n_n4948) & (!n_n4957) & (n_n4971)) + ((n_n4974) & (n_n4948) & (n_n4957) & (!n_n4971)) + ((n_n4974) & (n_n4948) & (n_n4957) & (n_n4971)));
	assign x13842x = (((!n_n3803) & (!n_n4949) & (!n_n4963) & (!n_n4947) & (n_n4962)) + ((!n_n3803) & (!n_n4949) & (!n_n4963) & (n_n4947) & (!n_n4962)) + ((!n_n3803) & (!n_n4949) & (!n_n4963) & (n_n4947) & (n_n4962)) + ((!n_n3803) & (!n_n4949) & (n_n4963) & (!n_n4947) & (!n_n4962)) + ((!n_n3803) & (!n_n4949) & (n_n4963) & (!n_n4947) & (n_n4962)) + ((!n_n3803) & (!n_n4949) & (n_n4963) & (n_n4947) & (!n_n4962)) + ((!n_n3803) & (!n_n4949) & (n_n4963) & (n_n4947) & (n_n4962)) + ((!n_n3803) & (n_n4949) & (!n_n4963) & (!n_n4947) & (!n_n4962)) + ((!n_n3803) & (n_n4949) & (!n_n4963) & (!n_n4947) & (n_n4962)) + ((!n_n3803) & (n_n4949) & (!n_n4963) & (n_n4947) & (!n_n4962)) + ((!n_n3803) & (n_n4949) & (!n_n4963) & (n_n4947) & (n_n4962)) + ((!n_n3803) & (n_n4949) & (n_n4963) & (!n_n4947) & (!n_n4962)) + ((!n_n3803) & (n_n4949) & (n_n4963) & (!n_n4947) & (n_n4962)) + ((!n_n3803) & (n_n4949) & (n_n4963) & (n_n4947) & (!n_n4962)) + ((!n_n3803) & (n_n4949) & (n_n4963) & (n_n4947) & (n_n4962)) + ((n_n3803) & (!n_n4949) & (!n_n4963) & (!n_n4947) & (!n_n4962)) + ((n_n3803) & (!n_n4949) & (!n_n4963) & (!n_n4947) & (n_n4962)) + ((n_n3803) & (!n_n4949) & (!n_n4963) & (n_n4947) & (!n_n4962)) + ((n_n3803) & (!n_n4949) & (!n_n4963) & (n_n4947) & (n_n4962)) + ((n_n3803) & (!n_n4949) & (n_n4963) & (!n_n4947) & (!n_n4962)) + ((n_n3803) & (!n_n4949) & (n_n4963) & (!n_n4947) & (n_n4962)) + ((n_n3803) & (!n_n4949) & (n_n4963) & (n_n4947) & (!n_n4962)) + ((n_n3803) & (!n_n4949) & (n_n4963) & (n_n4947) & (n_n4962)) + ((n_n3803) & (n_n4949) & (!n_n4963) & (!n_n4947) & (!n_n4962)) + ((n_n3803) & (n_n4949) & (!n_n4963) & (!n_n4947) & (n_n4962)) + ((n_n3803) & (n_n4949) & (!n_n4963) & (n_n4947) & (!n_n4962)) + ((n_n3803) & (n_n4949) & (!n_n4963) & (n_n4947) & (n_n4962)) + ((n_n3803) & (n_n4949) & (n_n4963) & (!n_n4947) & (!n_n4962)) + ((n_n3803) & (n_n4949) & (n_n4963) & (!n_n4947) & (n_n4962)) + ((n_n3803) & (n_n4949) & (n_n4963) & (n_n4947) & (!n_n4962)) + ((n_n3803) & (n_n4949) & (n_n4963) & (n_n4947) & (n_n4962)));
	assign n_n3272 = (((!n_n3318) & (!x229x) & (!x13841x) & (x13842x)) + ((!n_n3318) & (!x229x) & (x13841x) & (!x13842x)) + ((!n_n3318) & (!x229x) & (x13841x) & (x13842x)) + ((!n_n3318) & (x229x) & (!x13841x) & (!x13842x)) + ((!n_n3318) & (x229x) & (!x13841x) & (x13842x)) + ((!n_n3318) & (x229x) & (x13841x) & (!x13842x)) + ((!n_n3318) & (x229x) & (x13841x) & (x13842x)) + ((n_n3318) & (!x229x) & (!x13841x) & (!x13842x)) + ((n_n3318) & (!x229x) & (!x13841x) & (x13842x)) + ((n_n3318) & (!x229x) & (x13841x) & (!x13842x)) + ((n_n3318) & (!x229x) & (x13841x) & (x13842x)) + ((n_n3318) & (x229x) & (!x13841x) & (!x13842x)) + ((n_n3318) & (x229x) & (!x13841x) & (x13842x)) + ((n_n3318) & (x229x) & (x13841x) & (!x13842x)) + ((n_n3318) & (x229x) & (x13841x) & (x13842x)));
	assign n_n3515 = (((!i_9_) & (!n_n524) & (n_n526) & (n_n455) & (n_n509)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n455) & (n_n509)) + ((i_9_) & (!n_n524) & (n_n526) & (n_n455) & (n_n509)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n455) & (n_n509)) + ((i_9_) & (n_n524) & (n_n526) & (n_n455) & (n_n509)));
	assign n_n4490 = (((i_9_) & (n_n455) & (n_n532) & (n_n500)));
	assign n_n4479 = (((!i_9_) & (n_n455) & (n_n528) & (n_n509)));
	assign n_n901 = (((!i_9_) & (n_n455) & (!n_n528) & (n_n509) & (n_n530)) + ((!i_9_) & (n_n455) & (n_n528) & (n_n509) & (!n_n530)) + ((!i_9_) & (n_n455) & (n_n528) & (n_n509) & (n_n530)) + ((i_9_) & (n_n455) & (n_n528) & (n_n509) & (!n_n530)) + ((i_9_) & (n_n455) & (n_n528) & (n_n509) & (n_n530)));
	assign x14122x = (((!n_n4463) & (!n_n4460) & (!n_n4466) & (!n_n4457) & (n_n4465)) + ((!n_n4463) & (!n_n4460) & (!n_n4466) & (n_n4457) & (!n_n4465)) + ((!n_n4463) & (!n_n4460) & (!n_n4466) & (n_n4457) & (n_n4465)) + ((!n_n4463) & (!n_n4460) & (n_n4466) & (!n_n4457) & (!n_n4465)) + ((!n_n4463) & (!n_n4460) & (n_n4466) & (!n_n4457) & (n_n4465)) + ((!n_n4463) & (!n_n4460) & (n_n4466) & (n_n4457) & (!n_n4465)) + ((!n_n4463) & (!n_n4460) & (n_n4466) & (n_n4457) & (n_n4465)) + ((!n_n4463) & (n_n4460) & (!n_n4466) & (!n_n4457) & (!n_n4465)) + ((!n_n4463) & (n_n4460) & (!n_n4466) & (!n_n4457) & (n_n4465)) + ((!n_n4463) & (n_n4460) & (!n_n4466) & (n_n4457) & (!n_n4465)) + ((!n_n4463) & (n_n4460) & (!n_n4466) & (n_n4457) & (n_n4465)) + ((!n_n4463) & (n_n4460) & (n_n4466) & (!n_n4457) & (!n_n4465)) + ((!n_n4463) & (n_n4460) & (n_n4466) & (!n_n4457) & (n_n4465)) + ((!n_n4463) & (n_n4460) & (n_n4466) & (n_n4457) & (!n_n4465)) + ((!n_n4463) & (n_n4460) & (n_n4466) & (n_n4457) & (n_n4465)) + ((n_n4463) & (!n_n4460) & (!n_n4466) & (!n_n4457) & (!n_n4465)) + ((n_n4463) & (!n_n4460) & (!n_n4466) & (!n_n4457) & (n_n4465)) + ((n_n4463) & (!n_n4460) & (!n_n4466) & (n_n4457) & (!n_n4465)) + ((n_n4463) & (!n_n4460) & (!n_n4466) & (n_n4457) & (n_n4465)) + ((n_n4463) & (!n_n4460) & (n_n4466) & (!n_n4457) & (!n_n4465)) + ((n_n4463) & (!n_n4460) & (n_n4466) & (!n_n4457) & (n_n4465)) + ((n_n4463) & (!n_n4460) & (n_n4466) & (n_n4457) & (!n_n4465)) + ((n_n4463) & (!n_n4460) & (n_n4466) & (n_n4457) & (n_n4465)) + ((n_n4463) & (n_n4460) & (!n_n4466) & (!n_n4457) & (!n_n4465)) + ((n_n4463) & (n_n4460) & (!n_n4466) & (!n_n4457) & (n_n4465)) + ((n_n4463) & (n_n4460) & (!n_n4466) & (n_n4457) & (!n_n4465)) + ((n_n4463) & (n_n4460) & (!n_n4466) & (n_n4457) & (n_n4465)) + ((n_n4463) & (n_n4460) & (n_n4466) & (!n_n4457) & (!n_n4465)) + ((n_n4463) & (n_n4460) & (n_n4466) & (!n_n4457) & (n_n4465)) + ((n_n4463) & (n_n4460) & (n_n4466) & (n_n4457) & (!n_n4465)) + ((n_n4463) & (n_n4460) & (n_n4466) & (n_n4457) & (n_n4465)));
	assign n_n3358 = (((!n_n4459) & (!n_n4461) & (!n_n4455) & (!n_n4454) & (x14122x)) + ((!n_n4459) & (!n_n4461) & (!n_n4455) & (n_n4454) & (!x14122x)) + ((!n_n4459) & (!n_n4461) & (!n_n4455) & (n_n4454) & (x14122x)) + ((!n_n4459) & (!n_n4461) & (n_n4455) & (!n_n4454) & (!x14122x)) + ((!n_n4459) & (!n_n4461) & (n_n4455) & (!n_n4454) & (x14122x)) + ((!n_n4459) & (!n_n4461) & (n_n4455) & (n_n4454) & (!x14122x)) + ((!n_n4459) & (!n_n4461) & (n_n4455) & (n_n4454) & (x14122x)) + ((!n_n4459) & (n_n4461) & (!n_n4455) & (!n_n4454) & (!x14122x)) + ((!n_n4459) & (n_n4461) & (!n_n4455) & (!n_n4454) & (x14122x)) + ((!n_n4459) & (n_n4461) & (!n_n4455) & (n_n4454) & (!x14122x)) + ((!n_n4459) & (n_n4461) & (!n_n4455) & (n_n4454) & (x14122x)) + ((!n_n4459) & (n_n4461) & (n_n4455) & (!n_n4454) & (!x14122x)) + ((!n_n4459) & (n_n4461) & (n_n4455) & (!n_n4454) & (x14122x)) + ((!n_n4459) & (n_n4461) & (n_n4455) & (n_n4454) & (!x14122x)) + ((!n_n4459) & (n_n4461) & (n_n4455) & (n_n4454) & (x14122x)) + ((n_n4459) & (!n_n4461) & (!n_n4455) & (!n_n4454) & (!x14122x)) + ((n_n4459) & (!n_n4461) & (!n_n4455) & (!n_n4454) & (x14122x)) + ((n_n4459) & (!n_n4461) & (!n_n4455) & (n_n4454) & (!x14122x)) + ((n_n4459) & (!n_n4461) & (!n_n4455) & (n_n4454) & (x14122x)) + ((n_n4459) & (!n_n4461) & (n_n4455) & (!n_n4454) & (!x14122x)) + ((n_n4459) & (!n_n4461) & (n_n4455) & (!n_n4454) & (x14122x)) + ((n_n4459) & (!n_n4461) & (n_n4455) & (n_n4454) & (!x14122x)) + ((n_n4459) & (!n_n4461) & (n_n4455) & (n_n4454) & (x14122x)) + ((n_n4459) & (n_n4461) & (!n_n4455) & (!n_n4454) & (!x14122x)) + ((n_n4459) & (n_n4461) & (!n_n4455) & (!n_n4454) & (x14122x)) + ((n_n4459) & (n_n4461) & (!n_n4455) & (n_n4454) & (!x14122x)) + ((n_n4459) & (n_n4461) & (!n_n4455) & (n_n4454) & (x14122x)) + ((n_n4459) & (n_n4461) & (n_n4455) & (!n_n4454) & (!x14122x)) + ((n_n4459) & (n_n4461) & (n_n4455) & (!n_n4454) & (x14122x)) + ((n_n4459) & (n_n4461) & (n_n4455) & (n_n4454) & (!x14122x)) + ((n_n4459) & (n_n4461) & (n_n4455) & (n_n4454) & (x14122x)));
	assign n_n4475 = (((!i_9_) & (n_n455) & (n_n532) & (n_n509)));
	assign x163x = (((!i_9_) & (n_n455) & (n_n532) & (n_n500) & (!n_n530)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n500) & (n_n530)) + ((i_9_) & (n_n455) & (!n_n532) & (n_n500) & (n_n530)) + ((i_9_) & (n_n455) & (n_n532) & (n_n500) & (n_n530)));
	assign n_n4469 = (((!i_5_) & (i_3_) & (i_4_) & (n_n455) & (x20x)));
	assign x194x = (((!i_9_) & (n_n518) & (n_n455) & (!n_n520) & (x20x)) + ((!i_9_) & (n_n518) & (n_n455) & (n_n520) & (x20x)) + ((i_9_) & (n_n518) & (n_n455) & (!n_n520) & (x20x)) + ((i_9_) & (n_n518) & (n_n455) & (n_n520) & (!x20x)) + ((i_9_) & (n_n518) & (n_n455) & (n_n520) & (x20x)));
	assign x14128x = (((!n_n4471) & (!n_n4483) & (!n_n4488) & (n_n4490)) + ((!n_n4471) & (!n_n4483) & (n_n4488) & (!n_n4490)) + ((!n_n4471) & (!n_n4483) & (n_n4488) & (n_n4490)) + ((!n_n4471) & (n_n4483) & (!n_n4488) & (!n_n4490)) + ((!n_n4471) & (n_n4483) & (!n_n4488) & (n_n4490)) + ((!n_n4471) & (n_n4483) & (n_n4488) & (!n_n4490)) + ((!n_n4471) & (n_n4483) & (n_n4488) & (n_n4490)) + ((n_n4471) & (!n_n4483) & (!n_n4488) & (!n_n4490)) + ((n_n4471) & (!n_n4483) & (!n_n4488) & (n_n4490)) + ((n_n4471) & (!n_n4483) & (n_n4488) & (!n_n4490)) + ((n_n4471) & (!n_n4483) & (n_n4488) & (n_n4490)) + ((n_n4471) & (n_n4483) & (!n_n4488) & (!n_n4490)) + ((n_n4471) & (n_n4483) & (!n_n4488) & (n_n4490)) + ((n_n4471) & (n_n4483) & (n_n4488) & (!n_n4490)) + ((n_n4471) & (n_n4483) & (n_n4488) & (n_n4490)));
	assign x14130x = (((!n_n4467) & (!n_n4489) & (!x78x) & (!x163x) & (x194x)) + ((!n_n4467) & (!n_n4489) & (!x78x) & (x163x) & (!x194x)) + ((!n_n4467) & (!n_n4489) & (!x78x) & (x163x) & (x194x)) + ((!n_n4467) & (!n_n4489) & (x78x) & (!x163x) & (!x194x)) + ((!n_n4467) & (!n_n4489) & (x78x) & (!x163x) & (x194x)) + ((!n_n4467) & (!n_n4489) & (x78x) & (x163x) & (!x194x)) + ((!n_n4467) & (!n_n4489) & (x78x) & (x163x) & (x194x)) + ((!n_n4467) & (n_n4489) & (!x78x) & (!x163x) & (!x194x)) + ((!n_n4467) & (n_n4489) & (!x78x) & (!x163x) & (x194x)) + ((!n_n4467) & (n_n4489) & (!x78x) & (x163x) & (!x194x)) + ((!n_n4467) & (n_n4489) & (!x78x) & (x163x) & (x194x)) + ((!n_n4467) & (n_n4489) & (x78x) & (!x163x) & (!x194x)) + ((!n_n4467) & (n_n4489) & (x78x) & (!x163x) & (x194x)) + ((!n_n4467) & (n_n4489) & (x78x) & (x163x) & (!x194x)) + ((!n_n4467) & (n_n4489) & (x78x) & (x163x) & (x194x)) + ((n_n4467) & (!n_n4489) & (!x78x) & (!x163x) & (!x194x)) + ((n_n4467) & (!n_n4489) & (!x78x) & (!x163x) & (x194x)) + ((n_n4467) & (!n_n4489) & (!x78x) & (x163x) & (!x194x)) + ((n_n4467) & (!n_n4489) & (!x78x) & (x163x) & (x194x)) + ((n_n4467) & (!n_n4489) & (x78x) & (!x163x) & (!x194x)) + ((n_n4467) & (!n_n4489) & (x78x) & (!x163x) & (x194x)) + ((n_n4467) & (!n_n4489) & (x78x) & (x163x) & (!x194x)) + ((n_n4467) & (!n_n4489) & (x78x) & (x163x) & (x194x)) + ((n_n4467) & (n_n4489) & (!x78x) & (!x163x) & (!x194x)) + ((n_n4467) & (n_n4489) & (!x78x) & (!x163x) & (x194x)) + ((n_n4467) & (n_n4489) & (!x78x) & (x163x) & (!x194x)) + ((n_n4467) & (n_n4489) & (!x78x) & (x163x) & (x194x)) + ((n_n4467) & (n_n4489) & (x78x) & (!x163x) & (!x194x)) + ((n_n4467) & (n_n4489) & (x78x) & (!x163x) & (x194x)) + ((n_n4467) & (n_n4489) & (x78x) & (x163x) & (!x194x)) + ((n_n4467) & (n_n4489) & (x78x) & (x163x) & (x194x)));
	assign n_n3285 = (((!n_n3515) & (!n_n901) & (!n_n3358) & (!x14128x) & (x14130x)) + ((!n_n3515) & (!n_n901) & (!n_n3358) & (x14128x) & (!x14130x)) + ((!n_n3515) & (!n_n901) & (!n_n3358) & (x14128x) & (x14130x)) + ((!n_n3515) & (!n_n901) & (n_n3358) & (!x14128x) & (!x14130x)) + ((!n_n3515) & (!n_n901) & (n_n3358) & (!x14128x) & (x14130x)) + ((!n_n3515) & (!n_n901) & (n_n3358) & (x14128x) & (!x14130x)) + ((!n_n3515) & (!n_n901) & (n_n3358) & (x14128x) & (x14130x)) + ((!n_n3515) & (n_n901) & (!n_n3358) & (!x14128x) & (!x14130x)) + ((!n_n3515) & (n_n901) & (!n_n3358) & (!x14128x) & (x14130x)) + ((!n_n3515) & (n_n901) & (!n_n3358) & (x14128x) & (!x14130x)) + ((!n_n3515) & (n_n901) & (!n_n3358) & (x14128x) & (x14130x)) + ((!n_n3515) & (n_n901) & (n_n3358) & (!x14128x) & (!x14130x)) + ((!n_n3515) & (n_n901) & (n_n3358) & (!x14128x) & (x14130x)) + ((!n_n3515) & (n_n901) & (n_n3358) & (x14128x) & (!x14130x)) + ((!n_n3515) & (n_n901) & (n_n3358) & (x14128x) & (x14130x)) + ((n_n3515) & (!n_n901) & (!n_n3358) & (!x14128x) & (!x14130x)) + ((n_n3515) & (!n_n901) & (!n_n3358) & (!x14128x) & (x14130x)) + ((n_n3515) & (!n_n901) & (!n_n3358) & (x14128x) & (!x14130x)) + ((n_n3515) & (!n_n901) & (!n_n3358) & (x14128x) & (x14130x)) + ((n_n3515) & (!n_n901) & (n_n3358) & (!x14128x) & (!x14130x)) + ((n_n3515) & (!n_n901) & (n_n3358) & (!x14128x) & (x14130x)) + ((n_n3515) & (!n_n901) & (n_n3358) & (x14128x) & (!x14130x)) + ((n_n3515) & (!n_n901) & (n_n3358) & (x14128x) & (x14130x)) + ((n_n3515) & (n_n901) & (!n_n3358) & (!x14128x) & (!x14130x)) + ((n_n3515) & (n_n901) & (!n_n3358) & (!x14128x) & (x14130x)) + ((n_n3515) & (n_n901) & (!n_n3358) & (x14128x) & (!x14130x)) + ((n_n3515) & (n_n901) & (!n_n3358) & (x14128x) & (x14130x)) + ((n_n3515) & (n_n901) & (n_n3358) & (!x14128x) & (!x14130x)) + ((n_n3515) & (n_n901) & (n_n3358) & (!x14128x) & (x14130x)) + ((n_n3515) & (n_n901) & (n_n3358) & (x14128x) & (!x14130x)) + ((n_n3515) & (n_n901) & (n_n3358) & (x14128x) & (x14130x)));
	assign n_n2059 = (((!i_9_) & (!n_n524) & (n_n526) & (n_n455) & (n_n535)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n455) & (n_n535)) + ((i_9_) & (!n_n524) & (n_n526) & (n_n455) & (n_n535)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n455) & (n_n535)) + ((i_9_) & (n_n524) & (n_n526) & (n_n455) & (n_n535)));
	assign n_n4423 = (((i_1_) & (i_2_) & (i_0_) & (n_n473) & (x23x)));
	assign x14138x = (((!n_n4434) & (!n_n4432) & (!n_n4431) & (n_n4441)) + ((!n_n4434) & (!n_n4432) & (n_n4431) & (!n_n4441)) + ((!n_n4434) & (!n_n4432) & (n_n4431) & (n_n4441)) + ((!n_n4434) & (n_n4432) & (!n_n4431) & (!n_n4441)) + ((!n_n4434) & (n_n4432) & (!n_n4431) & (n_n4441)) + ((!n_n4434) & (n_n4432) & (n_n4431) & (!n_n4441)) + ((!n_n4434) & (n_n4432) & (n_n4431) & (n_n4441)) + ((n_n4434) & (!n_n4432) & (!n_n4431) & (!n_n4441)) + ((n_n4434) & (!n_n4432) & (!n_n4431) & (n_n4441)) + ((n_n4434) & (!n_n4432) & (n_n4431) & (!n_n4441)) + ((n_n4434) & (!n_n4432) & (n_n4431) & (n_n4441)) + ((n_n4434) & (n_n4432) & (!n_n4431) & (!n_n4441)) + ((n_n4434) & (n_n4432) & (!n_n4431) & (n_n4441)) + ((n_n4434) & (n_n4432) & (n_n4431) & (!n_n4441)) + ((n_n4434) & (n_n4432) & (n_n4431) & (n_n4441)));
	assign x421x = (((!i_9_) & (n_n455) & (n_n532) & (n_n535)) + ((i_9_) & (n_n455) & (n_n532) & (n_n535)));
	assign x14139x = (((!n_n4436) & (!x23x) & (!x496x) & (!n_n4435) & (x421x)) + ((!n_n4436) & (!x23x) & (!x496x) & (n_n4435) & (!x421x)) + ((!n_n4436) & (!x23x) & (!x496x) & (n_n4435) & (x421x)) + ((!n_n4436) & (!x23x) & (x496x) & (!n_n4435) & (x421x)) + ((!n_n4436) & (!x23x) & (x496x) & (n_n4435) & (!x421x)) + ((!n_n4436) & (!x23x) & (x496x) & (n_n4435) & (x421x)) + ((!n_n4436) & (x23x) & (!x496x) & (!n_n4435) & (x421x)) + ((!n_n4436) & (x23x) & (!x496x) & (n_n4435) & (!x421x)) + ((!n_n4436) & (x23x) & (!x496x) & (n_n4435) & (x421x)) + ((!n_n4436) & (x23x) & (x496x) & (!n_n4435) & (!x421x)) + ((!n_n4436) & (x23x) & (x496x) & (!n_n4435) & (x421x)) + ((!n_n4436) & (x23x) & (x496x) & (n_n4435) & (!x421x)) + ((!n_n4436) & (x23x) & (x496x) & (n_n4435) & (x421x)) + ((n_n4436) & (!x23x) & (!x496x) & (!n_n4435) & (!x421x)) + ((n_n4436) & (!x23x) & (!x496x) & (!n_n4435) & (x421x)) + ((n_n4436) & (!x23x) & (!x496x) & (n_n4435) & (!x421x)) + ((n_n4436) & (!x23x) & (!x496x) & (n_n4435) & (x421x)) + ((n_n4436) & (!x23x) & (x496x) & (!n_n4435) & (!x421x)) + ((n_n4436) & (!x23x) & (x496x) & (!n_n4435) & (x421x)) + ((n_n4436) & (!x23x) & (x496x) & (n_n4435) & (!x421x)) + ((n_n4436) & (!x23x) & (x496x) & (n_n4435) & (x421x)) + ((n_n4436) & (x23x) & (!x496x) & (!n_n4435) & (!x421x)) + ((n_n4436) & (x23x) & (!x496x) & (!n_n4435) & (x421x)) + ((n_n4436) & (x23x) & (!x496x) & (n_n4435) & (!x421x)) + ((n_n4436) & (x23x) & (!x496x) & (n_n4435) & (x421x)) + ((n_n4436) & (x23x) & (x496x) & (!n_n4435) & (!x421x)) + ((n_n4436) & (x23x) & (x496x) & (!n_n4435) & (x421x)) + ((n_n4436) & (x23x) & (x496x) & (n_n4435) & (!x421x)) + ((n_n4436) & (x23x) & (x496x) & (n_n4435) & (x421x)));
	assign x32x = (((!i_9_) & (n_n455) & (!n_n528) & (n_n535) & (n_n530)) + ((!i_9_) & (n_n455) & (n_n528) & (n_n535) & (n_n530)) + ((i_9_) & (n_n455) & (n_n528) & (n_n535) & (!n_n530)) + ((i_9_) & (n_n455) & (n_n528) & (n_n535) & (n_n530)));
	assign x470x = (((!i_9_) & (n_n455) & (!n_n528) & (n_n535) & (n_n530)) + ((!i_9_) & (n_n455) & (n_n528) & (n_n535) & (n_n530)) + ((i_9_) & (n_n455) & (!n_n528) & (n_n535) & (n_n530)) + ((i_9_) & (n_n455) & (n_n528) & (n_n535) & (!n_n530)) + ((i_9_) & (n_n455) & (n_n528) & (n_n535) & (n_n530)));
	assign x14147x = (((!n_n3520) & (!n_n2059) & (!n_n4423) & (!n_n4421) & (x470x)) + ((!n_n3520) & (!n_n2059) & (!n_n4423) & (n_n4421) & (!x470x)) + ((!n_n3520) & (!n_n2059) & (!n_n4423) & (n_n4421) & (x470x)) + ((!n_n3520) & (!n_n2059) & (n_n4423) & (!n_n4421) & (!x470x)) + ((!n_n3520) & (!n_n2059) & (n_n4423) & (!n_n4421) & (x470x)) + ((!n_n3520) & (!n_n2059) & (n_n4423) & (n_n4421) & (!x470x)) + ((!n_n3520) & (!n_n2059) & (n_n4423) & (n_n4421) & (x470x)) + ((!n_n3520) & (n_n2059) & (!n_n4423) & (!n_n4421) & (!x470x)) + ((!n_n3520) & (n_n2059) & (!n_n4423) & (!n_n4421) & (x470x)) + ((!n_n3520) & (n_n2059) & (!n_n4423) & (n_n4421) & (!x470x)) + ((!n_n3520) & (n_n2059) & (!n_n4423) & (n_n4421) & (x470x)) + ((!n_n3520) & (n_n2059) & (n_n4423) & (!n_n4421) & (!x470x)) + ((!n_n3520) & (n_n2059) & (n_n4423) & (!n_n4421) & (x470x)) + ((!n_n3520) & (n_n2059) & (n_n4423) & (n_n4421) & (!x470x)) + ((!n_n3520) & (n_n2059) & (n_n4423) & (n_n4421) & (x470x)) + ((n_n3520) & (!n_n2059) & (!n_n4423) & (!n_n4421) & (!x470x)) + ((n_n3520) & (!n_n2059) & (!n_n4423) & (!n_n4421) & (x470x)) + ((n_n3520) & (!n_n2059) & (!n_n4423) & (n_n4421) & (!x470x)) + ((n_n3520) & (!n_n2059) & (!n_n4423) & (n_n4421) & (x470x)) + ((n_n3520) & (!n_n2059) & (n_n4423) & (!n_n4421) & (!x470x)) + ((n_n3520) & (!n_n2059) & (n_n4423) & (!n_n4421) & (x470x)) + ((n_n3520) & (!n_n2059) & (n_n4423) & (n_n4421) & (!x470x)) + ((n_n3520) & (!n_n2059) & (n_n4423) & (n_n4421) & (x470x)) + ((n_n3520) & (n_n2059) & (!n_n4423) & (!n_n4421) & (!x470x)) + ((n_n3520) & (n_n2059) & (!n_n4423) & (!n_n4421) & (x470x)) + ((n_n3520) & (n_n2059) & (!n_n4423) & (n_n4421) & (!x470x)) + ((n_n3520) & (n_n2059) & (!n_n4423) & (n_n4421) & (x470x)) + ((n_n3520) & (n_n2059) & (n_n4423) & (!n_n4421) & (!x470x)) + ((n_n3520) & (n_n2059) & (n_n4423) & (!n_n4421) & (x470x)) + ((n_n3520) & (n_n2059) & (n_n4423) & (n_n4421) & (!x470x)) + ((n_n3520) & (n_n2059) & (n_n4423) & (n_n4421) & (x470x)));
	assign x14146x = (((!i_9_) & (!n_n536) & (!x506x) & (!x37x) & (x14143x)) + ((!i_9_) & (!n_n536) & (!x506x) & (x37x) & (!x14143x)) + ((!i_9_) & (!n_n536) & (!x506x) & (x37x) & (x14143x)) + ((!i_9_) & (!n_n536) & (x506x) & (!x37x) & (x14143x)) + ((!i_9_) & (!n_n536) & (x506x) & (x37x) & (!x14143x)) + ((!i_9_) & (!n_n536) & (x506x) & (x37x) & (x14143x)) + ((!i_9_) & (n_n536) & (!x506x) & (!x37x) & (x14143x)) + ((!i_9_) & (n_n536) & (!x506x) & (x37x) & (!x14143x)) + ((!i_9_) & (n_n536) & (!x506x) & (x37x) & (x14143x)) + ((!i_9_) & (n_n536) & (x506x) & (!x37x) & (x14143x)) + ((!i_9_) & (n_n536) & (x506x) & (x37x) & (!x14143x)) + ((!i_9_) & (n_n536) & (x506x) & (x37x) & (x14143x)) + ((i_9_) & (!n_n536) & (!x506x) & (!x37x) & (x14143x)) + ((i_9_) & (!n_n536) & (!x506x) & (x37x) & (!x14143x)) + ((i_9_) & (!n_n536) & (!x506x) & (x37x) & (x14143x)) + ((i_9_) & (!n_n536) & (x506x) & (!x37x) & (x14143x)) + ((i_9_) & (!n_n536) & (x506x) & (x37x) & (!x14143x)) + ((i_9_) & (!n_n536) & (x506x) & (x37x) & (x14143x)) + ((i_9_) & (n_n536) & (!x506x) & (!x37x) & (x14143x)) + ((i_9_) & (n_n536) & (!x506x) & (x37x) & (!x14143x)) + ((i_9_) & (n_n536) & (!x506x) & (x37x) & (x14143x)) + ((i_9_) & (n_n536) & (x506x) & (!x37x) & (!x14143x)) + ((i_9_) & (n_n536) & (x506x) & (!x37x) & (x14143x)) + ((i_9_) & (n_n536) & (x506x) & (x37x) & (!x14143x)) + ((i_9_) & (n_n536) & (x506x) & (x37x) & (x14143x)));
	assign n_n3286 = (((!x14138x) & (!x14139x) & (!x14147x) & (x14146x)) + ((!x14138x) & (!x14139x) & (x14147x) & (!x14146x)) + ((!x14138x) & (!x14139x) & (x14147x) & (x14146x)) + ((!x14138x) & (x14139x) & (!x14147x) & (!x14146x)) + ((!x14138x) & (x14139x) & (!x14147x) & (x14146x)) + ((!x14138x) & (x14139x) & (x14147x) & (!x14146x)) + ((!x14138x) & (x14139x) & (x14147x) & (x14146x)) + ((x14138x) & (!x14139x) & (!x14147x) & (!x14146x)) + ((x14138x) & (!x14139x) & (!x14147x) & (x14146x)) + ((x14138x) & (!x14139x) & (x14147x) & (!x14146x)) + ((x14138x) & (!x14139x) & (x14147x) & (x14146x)) + ((x14138x) & (x14139x) & (!x14147x) & (!x14146x)) + ((x14138x) & (x14139x) & (!x14147x) & (x14146x)) + ((x14138x) & (x14139x) & (x14147x) & (!x14146x)) + ((x14138x) & (x14139x) & (x14147x) & (x14146x)));
	assign n_n4630 = (((i_9_) & (n_n390) & (n_n520) & (n_n500)));
	assign n_n5287 = (((i_5_) & (!i_3_) & (i_4_) & (x23x) & (n_n65)));
	assign n_n5281 = (((!i_9_) & (n_n526) & (n_n491) & (n_n65)));
	assign n_n5268 = (((!i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n500)));
	assign n_n5261 = (((!i_9_) & (n_n500) & (n_n530) & (n_n65)));
	assign n_n5029 = (((i_5_) & (!i_3_) & (i_4_) & (n_n195) & (x20x)));
	assign n_n3162 = (((!i_9_) & (n_n524) & (n_n518) & (n_n455) & (!n_n522)) + ((!i_9_) & (n_n524) & (n_n518) & (n_n455) & (n_n522)) + ((i_9_) & (!n_n524) & (n_n518) & (n_n455) & (n_n522)) + ((i_9_) & (n_n524) & (n_n518) & (n_n455) & (!n_n522)) + ((i_9_) & (n_n524) & (n_n518) & (n_n455) & (n_n522)));
	assign x22082x = (((!n_n4477) & (!n_n4479) & (!n_n4475) & (!n_n4474)));
	assign n_n4614 = (((i_9_) & (n_n390) & (n_n509) & (n_n520)));
	assign n_n4232 = (((!n_n390) & (!n_n509) & (!x23x) & (!n_n4616) & (n_n4614)) + ((!n_n390) & (!n_n509) & (!x23x) & (n_n4616) & (!n_n4614)) + ((!n_n390) & (!n_n509) & (!x23x) & (n_n4616) & (n_n4614)) + ((!n_n390) & (!n_n509) & (x23x) & (!n_n4616) & (n_n4614)) + ((!n_n390) & (!n_n509) & (x23x) & (n_n4616) & (!n_n4614)) + ((!n_n390) & (!n_n509) & (x23x) & (n_n4616) & (n_n4614)) + ((!n_n390) & (n_n509) & (!x23x) & (!n_n4616) & (n_n4614)) + ((!n_n390) & (n_n509) & (!x23x) & (n_n4616) & (!n_n4614)) + ((!n_n390) & (n_n509) & (!x23x) & (n_n4616) & (n_n4614)) + ((!n_n390) & (n_n509) & (x23x) & (!n_n4616) & (n_n4614)) + ((!n_n390) & (n_n509) & (x23x) & (n_n4616) & (!n_n4614)) + ((!n_n390) & (n_n509) & (x23x) & (n_n4616) & (n_n4614)) + ((n_n390) & (!n_n509) & (!x23x) & (!n_n4616) & (n_n4614)) + ((n_n390) & (!n_n509) & (!x23x) & (n_n4616) & (!n_n4614)) + ((n_n390) & (!n_n509) & (!x23x) & (n_n4616) & (n_n4614)) + ((n_n390) & (!n_n509) & (x23x) & (!n_n4616) & (n_n4614)) + ((n_n390) & (!n_n509) & (x23x) & (n_n4616) & (!n_n4614)) + ((n_n390) & (!n_n509) & (x23x) & (n_n4616) & (n_n4614)) + ((n_n390) & (n_n509) & (!x23x) & (!n_n4616) & (n_n4614)) + ((n_n390) & (n_n509) & (!x23x) & (n_n4616) & (!n_n4614)) + ((n_n390) & (n_n509) & (!x23x) & (n_n4616) & (n_n4614)) + ((n_n390) & (n_n509) & (x23x) & (!n_n4616) & (!n_n4614)) + ((n_n390) & (n_n509) & (x23x) & (!n_n4616) & (n_n4614)) + ((n_n390) & (n_n509) & (x23x) & (n_n4616) & (!n_n4614)) + ((n_n390) & (n_n509) & (x23x) & (n_n4616) & (n_n4614)));
	assign n_n4620 = (((i_9_) & (n_n390) & (n_n500) & (n_n530)));
	assign x22226x = (((!n_n4617) & (!n_n4613) & (!n_n4607) & (!n_n4610)));
	assign x153x = (((!i_9_) & (n_n524) & (n_n482) & (!n_n522) & (n_n195)) + ((!i_9_) & (n_n524) & (n_n482) & (n_n522) & (n_n195)) + ((i_9_) & (!n_n524) & (n_n482) & (n_n522) & (n_n195)) + ((i_9_) & (n_n524) & (n_n482) & (n_n522) & (n_n195)));
	assign n_n2957 = (((!x13983x) & (!x13984x) & (!n_n5037) & (!n_n5045) & (x153x)) + ((!x13983x) & (!x13984x) & (!n_n5037) & (n_n5045) & (!x153x)) + ((!x13983x) & (!x13984x) & (!n_n5037) & (n_n5045) & (x153x)) + ((!x13983x) & (!x13984x) & (n_n5037) & (!n_n5045) & (!x153x)) + ((!x13983x) & (!x13984x) & (n_n5037) & (!n_n5045) & (x153x)) + ((!x13983x) & (!x13984x) & (n_n5037) & (n_n5045) & (!x153x)) + ((!x13983x) & (!x13984x) & (n_n5037) & (n_n5045) & (x153x)) + ((!x13983x) & (x13984x) & (!n_n5037) & (!n_n5045) & (!x153x)) + ((!x13983x) & (x13984x) & (!n_n5037) & (!n_n5045) & (x153x)) + ((!x13983x) & (x13984x) & (!n_n5037) & (n_n5045) & (!x153x)) + ((!x13983x) & (x13984x) & (!n_n5037) & (n_n5045) & (x153x)) + ((!x13983x) & (x13984x) & (n_n5037) & (!n_n5045) & (!x153x)) + ((!x13983x) & (x13984x) & (n_n5037) & (!n_n5045) & (x153x)) + ((!x13983x) & (x13984x) & (n_n5037) & (n_n5045) & (!x153x)) + ((!x13983x) & (x13984x) & (n_n5037) & (n_n5045) & (x153x)) + ((x13983x) & (!x13984x) & (!n_n5037) & (!n_n5045) & (!x153x)) + ((x13983x) & (!x13984x) & (!n_n5037) & (!n_n5045) & (x153x)) + ((x13983x) & (!x13984x) & (!n_n5037) & (n_n5045) & (!x153x)) + ((x13983x) & (!x13984x) & (!n_n5037) & (n_n5045) & (x153x)) + ((x13983x) & (!x13984x) & (n_n5037) & (!n_n5045) & (!x153x)) + ((x13983x) & (!x13984x) & (n_n5037) & (!n_n5045) & (x153x)) + ((x13983x) & (!x13984x) & (n_n5037) & (n_n5045) & (!x153x)) + ((x13983x) & (!x13984x) & (n_n5037) & (n_n5045) & (x153x)) + ((x13983x) & (x13984x) & (!n_n5037) & (!n_n5045) & (!x153x)) + ((x13983x) & (x13984x) & (!n_n5037) & (!n_n5045) & (x153x)) + ((x13983x) & (x13984x) & (!n_n5037) & (n_n5045) & (!x153x)) + ((x13983x) & (x13984x) & (!n_n5037) & (n_n5045) & (x153x)) + ((x13983x) & (x13984x) & (n_n5037) & (!n_n5045) & (!x153x)) + ((x13983x) & (x13984x) & (n_n5037) & (!n_n5045) & (x153x)) + ((x13983x) & (x13984x) & (n_n5037) & (n_n5045) & (!x153x)) + ((x13983x) & (x13984x) & (n_n5037) & (n_n5045) & (x153x)));
	assign n_n2601 = (((!x177x) & (!n_n4841) & (!n_n4837) & (!n_n3461) & (x304x)) + ((!x177x) & (!n_n4841) & (!n_n4837) & (n_n3461) & (!x304x)) + ((!x177x) & (!n_n4841) & (!n_n4837) & (n_n3461) & (x304x)) + ((!x177x) & (!n_n4841) & (n_n4837) & (!n_n3461) & (!x304x)) + ((!x177x) & (!n_n4841) & (n_n4837) & (!n_n3461) & (x304x)) + ((!x177x) & (!n_n4841) & (n_n4837) & (n_n3461) & (!x304x)) + ((!x177x) & (!n_n4841) & (n_n4837) & (n_n3461) & (x304x)) + ((!x177x) & (n_n4841) & (!n_n4837) & (!n_n3461) & (!x304x)) + ((!x177x) & (n_n4841) & (!n_n4837) & (!n_n3461) & (x304x)) + ((!x177x) & (n_n4841) & (!n_n4837) & (n_n3461) & (!x304x)) + ((!x177x) & (n_n4841) & (!n_n4837) & (n_n3461) & (x304x)) + ((!x177x) & (n_n4841) & (n_n4837) & (!n_n3461) & (!x304x)) + ((!x177x) & (n_n4841) & (n_n4837) & (!n_n3461) & (x304x)) + ((!x177x) & (n_n4841) & (n_n4837) & (n_n3461) & (!x304x)) + ((!x177x) & (n_n4841) & (n_n4837) & (n_n3461) & (x304x)) + ((x177x) & (!n_n4841) & (!n_n4837) & (!n_n3461) & (!x304x)) + ((x177x) & (!n_n4841) & (!n_n4837) & (!n_n3461) & (x304x)) + ((x177x) & (!n_n4841) & (!n_n4837) & (n_n3461) & (!x304x)) + ((x177x) & (!n_n4841) & (!n_n4837) & (n_n3461) & (x304x)) + ((x177x) & (!n_n4841) & (n_n4837) & (!n_n3461) & (!x304x)) + ((x177x) & (!n_n4841) & (n_n4837) & (!n_n3461) & (x304x)) + ((x177x) & (!n_n4841) & (n_n4837) & (n_n3461) & (!x304x)) + ((x177x) & (!n_n4841) & (n_n4837) & (n_n3461) & (x304x)) + ((x177x) & (n_n4841) & (!n_n4837) & (!n_n3461) & (!x304x)) + ((x177x) & (n_n4841) & (!n_n4837) & (!n_n3461) & (x304x)) + ((x177x) & (n_n4841) & (!n_n4837) & (n_n3461) & (!x304x)) + ((x177x) & (n_n4841) & (!n_n4837) & (n_n3461) & (x304x)) + ((x177x) & (n_n4841) & (n_n4837) & (!n_n3461) & (!x304x)) + ((x177x) & (n_n4841) & (n_n4837) & (!n_n3461) & (x304x)) + ((x177x) & (n_n4841) & (n_n4837) & (n_n3461) & (!x304x)) + ((x177x) & (n_n4841) & (n_n4837) & (n_n3461) & (x304x)));
	assign x389x = (((!i_9_) & (n_n325) & (!n_n520) & (x20x) & (n_n464)) + ((!i_9_) & (n_n325) & (n_n520) & (x20x) & (n_n464)) + ((i_9_) & (n_n325) & (!n_n520) & (x20x) & (n_n464)) + ((i_9_) & (n_n325) & (n_n520) & (!x20x) & (n_n464)) + ((i_9_) & (n_n325) & (n_n520) & (x20x) & (n_n464)));
	assign x14900x = (((!x23x) & (!x530x) & (!n_n4824) & (!x38x) & (n_n4818)) + ((!x23x) & (!x530x) & (!n_n4824) & (x38x) & (!n_n4818)) + ((!x23x) & (!x530x) & (!n_n4824) & (x38x) & (n_n4818)) + ((!x23x) & (!x530x) & (n_n4824) & (!x38x) & (!n_n4818)) + ((!x23x) & (!x530x) & (n_n4824) & (!x38x) & (n_n4818)) + ((!x23x) & (!x530x) & (n_n4824) & (x38x) & (!n_n4818)) + ((!x23x) & (!x530x) & (n_n4824) & (x38x) & (n_n4818)) + ((!x23x) & (x530x) & (!n_n4824) & (!x38x) & (n_n4818)) + ((!x23x) & (x530x) & (!n_n4824) & (x38x) & (!n_n4818)) + ((!x23x) & (x530x) & (!n_n4824) & (x38x) & (n_n4818)) + ((!x23x) & (x530x) & (n_n4824) & (!x38x) & (!n_n4818)) + ((!x23x) & (x530x) & (n_n4824) & (!x38x) & (n_n4818)) + ((!x23x) & (x530x) & (n_n4824) & (x38x) & (!n_n4818)) + ((!x23x) & (x530x) & (n_n4824) & (x38x) & (n_n4818)) + ((x23x) & (!x530x) & (!n_n4824) & (!x38x) & (n_n4818)) + ((x23x) & (!x530x) & (!n_n4824) & (x38x) & (!n_n4818)) + ((x23x) & (!x530x) & (!n_n4824) & (x38x) & (n_n4818)) + ((x23x) & (!x530x) & (n_n4824) & (!x38x) & (!n_n4818)) + ((x23x) & (!x530x) & (n_n4824) & (!x38x) & (n_n4818)) + ((x23x) & (!x530x) & (n_n4824) & (x38x) & (!n_n4818)) + ((x23x) & (!x530x) & (n_n4824) & (x38x) & (n_n4818)) + ((x23x) & (x530x) & (!n_n4824) & (!x38x) & (!n_n4818)) + ((x23x) & (x530x) & (!n_n4824) & (!x38x) & (n_n4818)) + ((x23x) & (x530x) & (!n_n4824) & (x38x) & (!n_n4818)) + ((x23x) & (x530x) & (!n_n4824) & (x38x) & (n_n4818)) + ((x23x) & (x530x) & (n_n4824) & (!x38x) & (!n_n4818)) + ((x23x) & (x530x) & (n_n4824) & (!x38x) & (n_n4818)) + ((x23x) & (x530x) & (n_n4824) & (x38x) & (!n_n4818)) + ((x23x) & (x530x) & (n_n4824) & (x38x) & (n_n4818)));
	assign x14907x = (((!n_n4827) & (!n_n4825) & (!n_n2601) & (!x389x) & (x14900x)) + ((!n_n4827) & (!n_n4825) & (!n_n2601) & (x389x) & (!x14900x)) + ((!n_n4827) & (!n_n4825) & (!n_n2601) & (x389x) & (x14900x)) + ((!n_n4827) & (!n_n4825) & (n_n2601) & (!x389x) & (!x14900x)) + ((!n_n4827) & (!n_n4825) & (n_n2601) & (!x389x) & (x14900x)) + ((!n_n4827) & (!n_n4825) & (n_n2601) & (x389x) & (!x14900x)) + ((!n_n4827) & (!n_n4825) & (n_n2601) & (x389x) & (x14900x)) + ((!n_n4827) & (n_n4825) & (!n_n2601) & (!x389x) & (!x14900x)) + ((!n_n4827) & (n_n4825) & (!n_n2601) & (!x389x) & (x14900x)) + ((!n_n4827) & (n_n4825) & (!n_n2601) & (x389x) & (!x14900x)) + ((!n_n4827) & (n_n4825) & (!n_n2601) & (x389x) & (x14900x)) + ((!n_n4827) & (n_n4825) & (n_n2601) & (!x389x) & (!x14900x)) + ((!n_n4827) & (n_n4825) & (n_n2601) & (!x389x) & (x14900x)) + ((!n_n4827) & (n_n4825) & (n_n2601) & (x389x) & (!x14900x)) + ((!n_n4827) & (n_n4825) & (n_n2601) & (x389x) & (x14900x)) + ((n_n4827) & (!n_n4825) & (!n_n2601) & (!x389x) & (!x14900x)) + ((n_n4827) & (!n_n4825) & (!n_n2601) & (!x389x) & (x14900x)) + ((n_n4827) & (!n_n4825) & (!n_n2601) & (x389x) & (!x14900x)) + ((n_n4827) & (!n_n4825) & (!n_n2601) & (x389x) & (x14900x)) + ((n_n4827) & (!n_n4825) & (n_n2601) & (!x389x) & (!x14900x)) + ((n_n4827) & (!n_n4825) & (n_n2601) & (!x389x) & (x14900x)) + ((n_n4827) & (!n_n4825) & (n_n2601) & (x389x) & (!x14900x)) + ((n_n4827) & (!n_n4825) & (n_n2601) & (x389x) & (x14900x)) + ((n_n4827) & (n_n4825) & (!n_n2601) & (!x389x) & (!x14900x)) + ((n_n4827) & (n_n4825) & (!n_n2601) & (!x389x) & (x14900x)) + ((n_n4827) & (n_n4825) & (!n_n2601) & (x389x) & (!x14900x)) + ((n_n4827) & (n_n4825) & (!n_n2601) & (x389x) & (x14900x)) + ((n_n4827) & (n_n4825) & (n_n2601) & (!x389x) & (!x14900x)) + ((n_n4827) & (n_n4825) & (n_n2601) & (!x389x) & (x14900x)) + ((n_n4827) & (n_n4825) & (n_n2601) & (x389x) & (!x14900x)) + ((n_n4827) & (n_n4825) & (n_n2601) & (x389x) & (x14900x)));
	assign x14904x = (((!n_n4856) & (!n_n4858) & (!n_n4853) & (n_n4845)) + ((!n_n4856) & (!n_n4858) & (n_n4853) & (!n_n4845)) + ((!n_n4856) & (!n_n4858) & (n_n4853) & (n_n4845)) + ((!n_n4856) & (n_n4858) & (!n_n4853) & (!n_n4845)) + ((!n_n4856) & (n_n4858) & (!n_n4853) & (n_n4845)) + ((!n_n4856) & (n_n4858) & (n_n4853) & (!n_n4845)) + ((!n_n4856) & (n_n4858) & (n_n4853) & (n_n4845)) + ((n_n4856) & (!n_n4858) & (!n_n4853) & (!n_n4845)) + ((n_n4856) & (!n_n4858) & (!n_n4853) & (n_n4845)) + ((n_n4856) & (!n_n4858) & (n_n4853) & (!n_n4845)) + ((n_n4856) & (!n_n4858) & (n_n4853) & (n_n4845)) + ((n_n4856) & (n_n4858) & (!n_n4853) & (!n_n4845)) + ((n_n4856) & (n_n4858) & (!n_n4853) & (n_n4845)) + ((n_n4856) & (n_n4858) & (n_n4853) & (!n_n4845)) + ((n_n4856) & (n_n4858) & (n_n4853) & (n_n4845)));
	assign n_n4874 = (((i_9_) & (n_n532) & (n_n260) & (n_n500)));
	assign x14908x = (((!i_9_) & (!n_n526) & (n_n528) & (n_n260) & (n_n500)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n260) & (n_n500)) + ((i_9_) & (n_n526) & (!n_n528) & (n_n260) & (n_n500)) + ((i_9_) & (n_n526) & (n_n528) & (n_n260) & (n_n500)));
	assign x12179x = (((!i_9_) & (n_n532) & (n_n260) & (n_n491)) + ((i_9_) & (n_n532) & (n_n260) & (n_n491)));
	assign x49x = (((!i_9_) & (n_n260) & (n_n491) & (n_n530)) + ((i_9_) & (n_n260) & (n_n491) & (n_n530)));
	assign n_n2727 = (((!i_9_) & (!n_n532) & (n_n509) & (n_n260) & (n_n530)) + ((!i_9_) & (n_n532) & (n_n509) & (n_n260) & (!n_n530)) + ((!i_9_) & (n_n532) & (n_n509) & (n_n260) & (n_n530)) + ((i_9_) & (!n_n532) & (n_n509) & (n_n260) & (n_n530)) + ((i_9_) & (n_n532) & (n_n509) & (n_n260) & (n_n530)));
	assign n_n4196 = (((!i_9_) & (!n_n528) & (n_n325) & (n_n530) & (n_n464)) + ((!i_9_) & (n_n528) & (n_n325) & (n_n530) & (n_n464)) + ((i_9_) & (!n_n528) & (n_n325) & (n_n530) & (n_n464)) + ((i_9_) & (n_n528) & (n_n325) & (!n_n530) & (n_n464)) + ((i_9_) & (n_n528) & (n_n325) & (n_n530) & (n_n464)));
	assign x14920x = (((!i_7_) & (!i_8_) & (i_6_) & (n_n482) & (x14x)) + ((i_7_) & (!i_8_) & (!i_6_) & (n_n482) & (x14x)));
	assign x14927x = (((!n_n4817) & (!n_n4792) & (!n_n4196) & (!n_n4197) & (x14920x)) + ((!n_n4817) & (!n_n4792) & (!n_n4196) & (n_n4197) & (!x14920x)) + ((!n_n4817) & (!n_n4792) & (!n_n4196) & (n_n4197) & (x14920x)) + ((!n_n4817) & (!n_n4792) & (n_n4196) & (!n_n4197) & (!x14920x)) + ((!n_n4817) & (!n_n4792) & (n_n4196) & (!n_n4197) & (x14920x)) + ((!n_n4817) & (!n_n4792) & (n_n4196) & (n_n4197) & (!x14920x)) + ((!n_n4817) & (!n_n4792) & (n_n4196) & (n_n4197) & (x14920x)) + ((!n_n4817) & (n_n4792) & (!n_n4196) & (!n_n4197) & (!x14920x)) + ((!n_n4817) & (n_n4792) & (!n_n4196) & (!n_n4197) & (x14920x)) + ((!n_n4817) & (n_n4792) & (!n_n4196) & (n_n4197) & (!x14920x)) + ((!n_n4817) & (n_n4792) & (!n_n4196) & (n_n4197) & (x14920x)) + ((!n_n4817) & (n_n4792) & (n_n4196) & (!n_n4197) & (!x14920x)) + ((!n_n4817) & (n_n4792) & (n_n4196) & (!n_n4197) & (x14920x)) + ((!n_n4817) & (n_n4792) & (n_n4196) & (n_n4197) & (!x14920x)) + ((!n_n4817) & (n_n4792) & (n_n4196) & (n_n4197) & (x14920x)) + ((n_n4817) & (!n_n4792) & (!n_n4196) & (!n_n4197) & (!x14920x)) + ((n_n4817) & (!n_n4792) & (!n_n4196) & (!n_n4197) & (x14920x)) + ((n_n4817) & (!n_n4792) & (!n_n4196) & (n_n4197) & (!x14920x)) + ((n_n4817) & (!n_n4792) & (!n_n4196) & (n_n4197) & (x14920x)) + ((n_n4817) & (!n_n4792) & (n_n4196) & (!n_n4197) & (!x14920x)) + ((n_n4817) & (!n_n4792) & (n_n4196) & (!n_n4197) & (x14920x)) + ((n_n4817) & (!n_n4792) & (n_n4196) & (n_n4197) & (!x14920x)) + ((n_n4817) & (!n_n4792) & (n_n4196) & (n_n4197) & (x14920x)) + ((n_n4817) & (n_n4792) & (!n_n4196) & (!n_n4197) & (!x14920x)) + ((n_n4817) & (n_n4792) & (!n_n4196) & (!n_n4197) & (x14920x)) + ((n_n4817) & (n_n4792) & (!n_n4196) & (n_n4197) & (!x14920x)) + ((n_n4817) & (n_n4792) & (!n_n4196) & (n_n4197) & (x14920x)) + ((n_n4817) & (n_n4792) & (n_n4196) & (!n_n4197) & (!x14920x)) + ((n_n4817) & (n_n4792) & (n_n4196) & (!n_n4197) & (x14920x)) + ((n_n4817) & (n_n4792) & (n_n4196) & (n_n4197) & (!x14920x)) + ((n_n4817) & (n_n4792) & (n_n4196) & (n_n4197) & (x14920x)));
	assign x14918x = (((!n_n4793) & (!n_n4798) & (!n_n4804) & (n_n4795)) + ((!n_n4793) & (!n_n4798) & (n_n4804) & (!n_n4795)) + ((!n_n4793) & (!n_n4798) & (n_n4804) & (n_n4795)) + ((!n_n4793) & (n_n4798) & (!n_n4804) & (!n_n4795)) + ((!n_n4793) & (n_n4798) & (!n_n4804) & (n_n4795)) + ((!n_n4793) & (n_n4798) & (n_n4804) & (!n_n4795)) + ((!n_n4793) & (n_n4798) & (n_n4804) & (n_n4795)) + ((n_n4793) & (!n_n4798) & (!n_n4804) & (!n_n4795)) + ((n_n4793) & (!n_n4798) & (!n_n4804) & (n_n4795)) + ((n_n4793) & (!n_n4798) & (n_n4804) & (!n_n4795)) + ((n_n4793) & (!n_n4798) & (n_n4804) & (n_n4795)) + ((n_n4793) & (n_n4798) & (!n_n4804) & (!n_n4795)) + ((n_n4793) & (n_n4798) & (!n_n4804) & (n_n4795)) + ((n_n4793) & (n_n4798) & (n_n4804) & (!n_n4795)) + ((n_n4793) & (n_n4798) & (n_n4804) & (n_n4795)));
	assign x14919x = (((!n_n4797) & (!n_n4802) & (!n_n4807) & (!n_n4808) & (n_n4799)) + ((!n_n4797) & (!n_n4802) & (!n_n4807) & (n_n4808) & (!n_n4799)) + ((!n_n4797) & (!n_n4802) & (!n_n4807) & (n_n4808) & (n_n4799)) + ((!n_n4797) & (!n_n4802) & (n_n4807) & (!n_n4808) & (!n_n4799)) + ((!n_n4797) & (!n_n4802) & (n_n4807) & (!n_n4808) & (n_n4799)) + ((!n_n4797) & (!n_n4802) & (n_n4807) & (n_n4808) & (!n_n4799)) + ((!n_n4797) & (!n_n4802) & (n_n4807) & (n_n4808) & (n_n4799)) + ((!n_n4797) & (n_n4802) & (!n_n4807) & (!n_n4808) & (!n_n4799)) + ((!n_n4797) & (n_n4802) & (!n_n4807) & (!n_n4808) & (n_n4799)) + ((!n_n4797) & (n_n4802) & (!n_n4807) & (n_n4808) & (!n_n4799)) + ((!n_n4797) & (n_n4802) & (!n_n4807) & (n_n4808) & (n_n4799)) + ((!n_n4797) & (n_n4802) & (n_n4807) & (!n_n4808) & (!n_n4799)) + ((!n_n4797) & (n_n4802) & (n_n4807) & (!n_n4808) & (n_n4799)) + ((!n_n4797) & (n_n4802) & (n_n4807) & (n_n4808) & (!n_n4799)) + ((!n_n4797) & (n_n4802) & (n_n4807) & (n_n4808) & (n_n4799)) + ((n_n4797) & (!n_n4802) & (!n_n4807) & (!n_n4808) & (!n_n4799)) + ((n_n4797) & (!n_n4802) & (!n_n4807) & (!n_n4808) & (n_n4799)) + ((n_n4797) & (!n_n4802) & (!n_n4807) & (n_n4808) & (!n_n4799)) + ((n_n4797) & (!n_n4802) & (!n_n4807) & (n_n4808) & (n_n4799)) + ((n_n4797) & (!n_n4802) & (n_n4807) & (!n_n4808) & (!n_n4799)) + ((n_n4797) & (!n_n4802) & (n_n4807) & (!n_n4808) & (n_n4799)) + ((n_n4797) & (!n_n4802) & (n_n4807) & (n_n4808) & (!n_n4799)) + ((n_n4797) & (!n_n4802) & (n_n4807) & (n_n4808) & (n_n4799)) + ((n_n4797) & (n_n4802) & (!n_n4807) & (!n_n4808) & (!n_n4799)) + ((n_n4797) & (n_n4802) & (!n_n4807) & (!n_n4808) & (n_n4799)) + ((n_n4797) & (n_n4802) & (!n_n4807) & (n_n4808) & (!n_n4799)) + ((n_n4797) & (n_n4802) & (!n_n4807) & (n_n4808) & (n_n4799)) + ((n_n4797) & (n_n4802) & (n_n4807) & (!n_n4808) & (!n_n4799)) + ((n_n4797) & (n_n4802) & (n_n4807) & (!n_n4808) & (n_n4799)) + ((n_n4797) & (n_n4802) & (n_n4807) & (n_n4808) & (!n_n4799)) + ((n_n4797) & (n_n4802) & (n_n4807) & (n_n4808) & (n_n4799)));
	assign x14926x = (((!x131x) & (!n_n4789) & (!n_n4788) & (!x191x) & (x151x)) + ((!x131x) & (!n_n4789) & (!n_n4788) & (x191x) & (!x151x)) + ((!x131x) & (!n_n4789) & (!n_n4788) & (x191x) & (x151x)) + ((!x131x) & (!n_n4789) & (n_n4788) & (!x191x) & (!x151x)) + ((!x131x) & (!n_n4789) & (n_n4788) & (!x191x) & (x151x)) + ((!x131x) & (!n_n4789) & (n_n4788) & (x191x) & (!x151x)) + ((!x131x) & (!n_n4789) & (n_n4788) & (x191x) & (x151x)) + ((!x131x) & (n_n4789) & (!n_n4788) & (!x191x) & (!x151x)) + ((!x131x) & (n_n4789) & (!n_n4788) & (!x191x) & (x151x)) + ((!x131x) & (n_n4789) & (!n_n4788) & (x191x) & (!x151x)) + ((!x131x) & (n_n4789) & (!n_n4788) & (x191x) & (x151x)) + ((!x131x) & (n_n4789) & (n_n4788) & (!x191x) & (!x151x)) + ((!x131x) & (n_n4789) & (n_n4788) & (!x191x) & (x151x)) + ((!x131x) & (n_n4789) & (n_n4788) & (x191x) & (!x151x)) + ((!x131x) & (n_n4789) & (n_n4788) & (x191x) & (x151x)) + ((x131x) & (!n_n4789) & (!n_n4788) & (!x191x) & (!x151x)) + ((x131x) & (!n_n4789) & (!n_n4788) & (!x191x) & (x151x)) + ((x131x) & (!n_n4789) & (!n_n4788) & (x191x) & (!x151x)) + ((x131x) & (!n_n4789) & (!n_n4788) & (x191x) & (x151x)) + ((x131x) & (!n_n4789) & (n_n4788) & (!x191x) & (!x151x)) + ((x131x) & (!n_n4789) & (n_n4788) & (!x191x) & (x151x)) + ((x131x) & (!n_n4789) & (n_n4788) & (x191x) & (!x151x)) + ((x131x) & (!n_n4789) & (n_n4788) & (x191x) & (x151x)) + ((x131x) & (n_n4789) & (!n_n4788) & (!x191x) & (!x151x)) + ((x131x) & (n_n4789) & (!n_n4788) & (!x191x) & (x151x)) + ((x131x) & (n_n4789) & (!n_n4788) & (x191x) & (!x151x)) + ((x131x) & (n_n4789) & (!n_n4788) & (x191x) & (x151x)) + ((x131x) & (n_n4789) & (n_n4788) & (!x191x) & (!x151x)) + ((x131x) & (n_n4789) & (n_n4788) & (!x191x) & (x151x)) + ((x131x) & (n_n4789) & (n_n4788) & (x191x) & (!x151x)) + ((x131x) & (n_n4789) & (n_n4788) & (x191x) & (x151x)));
	assign n_n4965 = (((i_5_) & (i_3_) & (i_4_) & (n_n195) & (x20x)));
	assign x22210x = (((!n_n4914) & (!n_n4918) & (!n_n4917) & (!n_n4915) & (!n_n2718)));
	assign x14960x = (((!n_n526) & (!n_n482) & (!x17x) & (!n_n522) & (!x22210x)) + ((!n_n526) & (!n_n482) & (!x17x) & (n_n522) & (!x22210x)) + ((!n_n526) & (!n_n482) & (x17x) & (!n_n522) & (!x22210x)) + ((!n_n526) & (!n_n482) & (x17x) & (n_n522) & (!x22210x)) + ((!n_n526) & (n_n482) & (!x17x) & (!n_n522) & (!x22210x)) + ((!n_n526) & (n_n482) & (!x17x) & (n_n522) & (!x22210x)) + ((!n_n526) & (n_n482) & (x17x) & (!n_n522) & (!x22210x)) + ((!n_n526) & (n_n482) & (x17x) & (n_n522) & (!x22210x)) + ((!n_n526) & (n_n482) & (x17x) & (n_n522) & (x22210x)) + ((n_n526) & (!n_n482) & (!x17x) & (!n_n522) & (!x22210x)) + ((n_n526) & (!n_n482) & (!x17x) & (n_n522) & (!x22210x)) + ((n_n526) & (!n_n482) & (x17x) & (!n_n522) & (!x22210x)) + ((n_n526) & (!n_n482) & (x17x) & (n_n522) & (!x22210x)) + ((n_n526) & (n_n482) & (!x17x) & (!n_n522) & (!x22210x)) + ((n_n526) & (n_n482) & (!x17x) & (n_n522) & (!x22210x)) + ((n_n526) & (n_n482) & (x17x) & (!n_n522) & (!x22210x)) + ((n_n526) & (n_n482) & (x17x) & (!n_n522) & (x22210x)) + ((n_n526) & (n_n482) & (x17x) & (n_n522) & (!x22210x)) + ((n_n526) & (n_n482) & (x17x) & (n_n522) & (x22210x)));
	assign x14948x = (((!n_n4927) & (!n_n4923) & (!n_n4924) & (n_n4921)) + ((!n_n4927) & (!n_n4923) & (n_n4924) & (!n_n4921)) + ((!n_n4927) & (!n_n4923) & (n_n4924) & (n_n4921)) + ((!n_n4927) & (n_n4923) & (!n_n4924) & (!n_n4921)) + ((!n_n4927) & (n_n4923) & (!n_n4924) & (n_n4921)) + ((!n_n4927) & (n_n4923) & (n_n4924) & (!n_n4921)) + ((!n_n4927) & (n_n4923) & (n_n4924) & (n_n4921)) + ((n_n4927) & (!n_n4923) & (!n_n4924) & (!n_n4921)) + ((n_n4927) & (!n_n4923) & (!n_n4924) & (n_n4921)) + ((n_n4927) & (!n_n4923) & (n_n4924) & (!n_n4921)) + ((n_n4927) & (!n_n4923) & (n_n4924) & (n_n4921)) + ((n_n4927) & (n_n4923) & (!n_n4924) & (!n_n4921)) + ((n_n4927) & (n_n4923) & (!n_n4924) & (n_n4921)) + ((n_n4927) & (n_n4923) & (n_n4924) & (!n_n4921)) + ((n_n4927) & (n_n4923) & (n_n4924) & (n_n4921)));
	assign x14949x = (((!n_n4920) & (!n_n4926) & (!n_n4930) & (!n_n4919) & (n_n4931)) + ((!n_n4920) & (!n_n4926) & (!n_n4930) & (n_n4919) & (!n_n4931)) + ((!n_n4920) & (!n_n4926) & (!n_n4930) & (n_n4919) & (n_n4931)) + ((!n_n4920) & (!n_n4926) & (n_n4930) & (!n_n4919) & (!n_n4931)) + ((!n_n4920) & (!n_n4926) & (n_n4930) & (!n_n4919) & (n_n4931)) + ((!n_n4920) & (!n_n4926) & (n_n4930) & (n_n4919) & (!n_n4931)) + ((!n_n4920) & (!n_n4926) & (n_n4930) & (n_n4919) & (n_n4931)) + ((!n_n4920) & (n_n4926) & (!n_n4930) & (!n_n4919) & (!n_n4931)) + ((!n_n4920) & (n_n4926) & (!n_n4930) & (!n_n4919) & (n_n4931)) + ((!n_n4920) & (n_n4926) & (!n_n4930) & (n_n4919) & (!n_n4931)) + ((!n_n4920) & (n_n4926) & (!n_n4930) & (n_n4919) & (n_n4931)) + ((!n_n4920) & (n_n4926) & (n_n4930) & (!n_n4919) & (!n_n4931)) + ((!n_n4920) & (n_n4926) & (n_n4930) & (!n_n4919) & (n_n4931)) + ((!n_n4920) & (n_n4926) & (n_n4930) & (n_n4919) & (!n_n4931)) + ((!n_n4920) & (n_n4926) & (n_n4930) & (n_n4919) & (n_n4931)) + ((n_n4920) & (!n_n4926) & (!n_n4930) & (!n_n4919) & (!n_n4931)) + ((n_n4920) & (!n_n4926) & (!n_n4930) & (!n_n4919) & (n_n4931)) + ((n_n4920) & (!n_n4926) & (!n_n4930) & (n_n4919) & (!n_n4931)) + ((n_n4920) & (!n_n4926) & (!n_n4930) & (n_n4919) & (n_n4931)) + ((n_n4920) & (!n_n4926) & (n_n4930) & (!n_n4919) & (!n_n4931)) + ((n_n4920) & (!n_n4926) & (n_n4930) & (!n_n4919) & (n_n4931)) + ((n_n4920) & (!n_n4926) & (n_n4930) & (n_n4919) & (!n_n4931)) + ((n_n4920) & (!n_n4926) & (n_n4930) & (n_n4919) & (n_n4931)) + ((n_n4920) & (n_n4926) & (!n_n4930) & (!n_n4919) & (!n_n4931)) + ((n_n4920) & (n_n4926) & (!n_n4930) & (!n_n4919) & (n_n4931)) + ((n_n4920) & (n_n4926) & (!n_n4930) & (n_n4919) & (!n_n4931)) + ((n_n4920) & (n_n4926) & (!n_n4930) & (n_n4919) & (n_n4931)) + ((n_n4920) & (n_n4926) & (n_n4930) & (!n_n4919) & (!n_n4931)) + ((n_n4920) & (n_n4926) & (n_n4930) & (!n_n4919) & (n_n4931)) + ((n_n4920) & (n_n4926) & (n_n4930) & (n_n4919) & (!n_n4931)) + ((n_n4920) & (n_n4926) & (n_n4930) & (n_n4919) & (n_n4931)));
	assign n_n2596 = (((!n_n4898) & (!n_n4903) & (!n_n4895) & (!n_n4908) & (x14955x)) + ((!n_n4898) & (!n_n4903) & (!n_n4895) & (n_n4908) & (!x14955x)) + ((!n_n4898) & (!n_n4903) & (!n_n4895) & (n_n4908) & (x14955x)) + ((!n_n4898) & (!n_n4903) & (n_n4895) & (!n_n4908) & (!x14955x)) + ((!n_n4898) & (!n_n4903) & (n_n4895) & (!n_n4908) & (x14955x)) + ((!n_n4898) & (!n_n4903) & (n_n4895) & (n_n4908) & (!x14955x)) + ((!n_n4898) & (!n_n4903) & (n_n4895) & (n_n4908) & (x14955x)) + ((!n_n4898) & (n_n4903) & (!n_n4895) & (!n_n4908) & (!x14955x)) + ((!n_n4898) & (n_n4903) & (!n_n4895) & (!n_n4908) & (x14955x)) + ((!n_n4898) & (n_n4903) & (!n_n4895) & (n_n4908) & (!x14955x)) + ((!n_n4898) & (n_n4903) & (!n_n4895) & (n_n4908) & (x14955x)) + ((!n_n4898) & (n_n4903) & (n_n4895) & (!n_n4908) & (!x14955x)) + ((!n_n4898) & (n_n4903) & (n_n4895) & (!n_n4908) & (x14955x)) + ((!n_n4898) & (n_n4903) & (n_n4895) & (n_n4908) & (!x14955x)) + ((!n_n4898) & (n_n4903) & (n_n4895) & (n_n4908) & (x14955x)) + ((n_n4898) & (!n_n4903) & (!n_n4895) & (!n_n4908) & (!x14955x)) + ((n_n4898) & (!n_n4903) & (!n_n4895) & (!n_n4908) & (x14955x)) + ((n_n4898) & (!n_n4903) & (!n_n4895) & (n_n4908) & (!x14955x)) + ((n_n4898) & (!n_n4903) & (!n_n4895) & (n_n4908) & (x14955x)) + ((n_n4898) & (!n_n4903) & (n_n4895) & (!n_n4908) & (!x14955x)) + ((n_n4898) & (!n_n4903) & (n_n4895) & (!n_n4908) & (x14955x)) + ((n_n4898) & (!n_n4903) & (n_n4895) & (n_n4908) & (!x14955x)) + ((n_n4898) & (!n_n4903) & (n_n4895) & (n_n4908) & (x14955x)) + ((n_n4898) & (n_n4903) & (!n_n4895) & (!n_n4908) & (!x14955x)) + ((n_n4898) & (n_n4903) & (!n_n4895) & (!n_n4908) & (x14955x)) + ((n_n4898) & (n_n4903) & (!n_n4895) & (n_n4908) & (!x14955x)) + ((n_n4898) & (n_n4903) & (!n_n4895) & (n_n4908) & (x14955x)) + ((n_n4898) & (n_n4903) & (n_n4895) & (!n_n4908) & (!x14955x)) + ((n_n4898) & (n_n4903) & (n_n4895) & (!n_n4908) & (x14955x)) + ((n_n4898) & (n_n4903) & (n_n4895) & (n_n4908) & (!x14955x)) + ((n_n4898) & (n_n4903) & (n_n4895) & (n_n4908) & (x14955x)));
	assign n_n1973 = (((!i_9_) & (n_n524) & (n_n260) & (!n_n522) & (n_n464)) + ((!i_9_) & (n_n524) & (n_n260) & (n_n522) & (n_n464)) + ((i_9_) & (!n_n524) & (n_n260) & (n_n522) & (n_n464)) + ((i_9_) & (n_n524) & (n_n260) & (!n_n522) & (n_n464)) + ((i_9_) & (n_n524) & (n_n260) & (n_n522) & (n_n464)));
	assign n_n2710 = (((!i_9_) & (!n_n528) & (n_n260) & (n_n530) & (n_n464)) + ((!i_9_) & (n_n528) & (n_n260) & (n_n530) & (n_n464)) + ((i_9_) & (!n_n528) & (n_n260) & (n_n530) & (n_n464)) + ((i_9_) & (n_n528) & (n_n260) & (!n_n530) & (n_n464)) + ((i_9_) & (n_n528) & (n_n260) & (n_n530) & (n_n464)));
	assign x58x = (((!i_9_) & (!n_n526) & (n_n528) & (n_n260) & (n_n464)) + ((!i_9_) & (n_n526) & (!n_n528) & (n_n260) & (n_n464)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n260) & (n_n464)) + ((i_9_) & (n_n526) & (!n_n528) & (n_n260) & (n_n464)) + ((i_9_) & (n_n526) & (n_n528) & (n_n260) & (n_n464)));
	assign x14974x = (((!n_n4936) & (!n_n4935) & (!n_n1973) & (!n_n2710) & (x58x)) + ((!n_n4936) & (!n_n4935) & (!n_n1973) & (n_n2710) & (!x58x)) + ((!n_n4936) & (!n_n4935) & (!n_n1973) & (n_n2710) & (x58x)) + ((!n_n4936) & (!n_n4935) & (n_n1973) & (!n_n2710) & (!x58x)) + ((!n_n4936) & (!n_n4935) & (n_n1973) & (!n_n2710) & (x58x)) + ((!n_n4936) & (!n_n4935) & (n_n1973) & (n_n2710) & (!x58x)) + ((!n_n4936) & (!n_n4935) & (n_n1973) & (n_n2710) & (x58x)) + ((!n_n4936) & (n_n4935) & (!n_n1973) & (!n_n2710) & (!x58x)) + ((!n_n4936) & (n_n4935) & (!n_n1973) & (!n_n2710) & (x58x)) + ((!n_n4936) & (n_n4935) & (!n_n1973) & (n_n2710) & (!x58x)) + ((!n_n4936) & (n_n4935) & (!n_n1973) & (n_n2710) & (x58x)) + ((!n_n4936) & (n_n4935) & (n_n1973) & (!n_n2710) & (!x58x)) + ((!n_n4936) & (n_n4935) & (n_n1973) & (!n_n2710) & (x58x)) + ((!n_n4936) & (n_n4935) & (n_n1973) & (n_n2710) & (!x58x)) + ((!n_n4936) & (n_n4935) & (n_n1973) & (n_n2710) & (x58x)) + ((n_n4936) & (!n_n4935) & (!n_n1973) & (!n_n2710) & (!x58x)) + ((n_n4936) & (!n_n4935) & (!n_n1973) & (!n_n2710) & (x58x)) + ((n_n4936) & (!n_n4935) & (!n_n1973) & (n_n2710) & (!x58x)) + ((n_n4936) & (!n_n4935) & (!n_n1973) & (n_n2710) & (x58x)) + ((n_n4936) & (!n_n4935) & (n_n1973) & (!n_n2710) & (!x58x)) + ((n_n4936) & (!n_n4935) & (n_n1973) & (!n_n2710) & (x58x)) + ((n_n4936) & (!n_n4935) & (n_n1973) & (n_n2710) & (!x58x)) + ((n_n4936) & (!n_n4935) & (n_n1973) & (n_n2710) & (x58x)) + ((n_n4936) & (n_n4935) & (!n_n1973) & (!n_n2710) & (!x58x)) + ((n_n4936) & (n_n4935) & (!n_n1973) & (!n_n2710) & (x58x)) + ((n_n4936) & (n_n4935) & (!n_n1973) & (n_n2710) & (!x58x)) + ((n_n4936) & (n_n4935) & (!n_n1973) & (n_n2710) & (x58x)) + ((n_n4936) & (n_n4935) & (n_n1973) & (!n_n2710) & (!x58x)) + ((n_n4936) & (n_n4935) & (n_n1973) & (!n_n2710) & (x58x)) + ((n_n4936) & (n_n4935) & (n_n1973) & (n_n2710) & (!x58x)) + ((n_n4936) & (n_n4935) & (n_n1973) & (n_n2710) & (x58x)));
	assign n_n2591 = (((!n_n4964) & (!n_n3802) & (!x250x) & (!n_n4957) & (x210x)) + ((!n_n4964) & (!n_n3802) & (!x250x) & (n_n4957) & (!x210x)) + ((!n_n4964) & (!n_n3802) & (!x250x) & (n_n4957) & (x210x)) + ((!n_n4964) & (!n_n3802) & (x250x) & (!n_n4957) & (!x210x)) + ((!n_n4964) & (!n_n3802) & (x250x) & (!n_n4957) & (x210x)) + ((!n_n4964) & (!n_n3802) & (x250x) & (n_n4957) & (!x210x)) + ((!n_n4964) & (!n_n3802) & (x250x) & (n_n4957) & (x210x)) + ((!n_n4964) & (n_n3802) & (!x250x) & (!n_n4957) & (!x210x)) + ((!n_n4964) & (n_n3802) & (!x250x) & (!n_n4957) & (x210x)) + ((!n_n4964) & (n_n3802) & (!x250x) & (n_n4957) & (!x210x)) + ((!n_n4964) & (n_n3802) & (!x250x) & (n_n4957) & (x210x)) + ((!n_n4964) & (n_n3802) & (x250x) & (!n_n4957) & (!x210x)) + ((!n_n4964) & (n_n3802) & (x250x) & (!n_n4957) & (x210x)) + ((!n_n4964) & (n_n3802) & (x250x) & (n_n4957) & (!x210x)) + ((!n_n4964) & (n_n3802) & (x250x) & (n_n4957) & (x210x)) + ((n_n4964) & (!n_n3802) & (!x250x) & (!n_n4957) & (!x210x)) + ((n_n4964) & (!n_n3802) & (!x250x) & (!n_n4957) & (x210x)) + ((n_n4964) & (!n_n3802) & (!x250x) & (n_n4957) & (!x210x)) + ((n_n4964) & (!n_n3802) & (!x250x) & (n_n4957) & (x210x)) + ((n_n4964) & (!n_n3802) & (x250x) & (!n_n4957) & (!x210x)) + ((n_n4964) & (!n_n3802) & (x250x) & (!n_n4957) & (x210x)) + ((n_n4964) & (!n_n3802) & (x250x) & (n_n4957) & (!x210x)) + ((n_n4964) & (!n_n3802) & (x250x) & (n_n4957) & (x210x)) + ((n_n4964) & (n_n3802) & (!x250x) & (!n_n4957) & (!x210x)) + ((n_n4964) & (n_n3802) & (!x250x) & (!n_n4957) & (x210x)) + ((n_n4964) & (n_n3802) & (!x250x) & (n_n4957) & (!x210x)) + ((n_n4964) & (n_n3802) & (!x250x) & (n_n4957) & (x210x)) + ((n_n4964) & (n_n3802) & (x250x) & (!n_n4957) & (!x210x)) + ((n_n4964) & (n_n3802) & (x250x) & (!n_n4957) & (x210x)) + ((n_n4964) & (n_n3802) & (x250x) & (n_n4957) & (!x210x)) + ((n_n4964) & (n_n3802) & (x250x) & (n_n4957) & (x210x)));
	assign x14970x = (((!x20x) & (!x531x) & (!n_n4952) & (!n_n4950) & (n_n4937)) + ((!x20x) & (!x531x) & (!n_n4952) & (n_n4950) & (!n_n4937)) + ((!x20x) & (!x531x) & (!n_n4952) & (n_n4950) & (n_n4937)) + ((!x20x) & (!x531x) & (n_n4952) & (!n_n4950) & (!n_n4937)) + ((!x20x) & (!x531x) & (n_n4952) & (!n_n4950) & (n_n4937)) + ((!x20x) & (!x531x) & (n_n4952) & (n_n4950) & (!n_n4937)) + ((!x20x) & (!x531x) & (n_n4952) & (n_n4950) & (n_n4937)) + ((!x20x) & (x531x) & (!n_n4952) & (!n_n4950) & (n_n4937)) + ((!x20x) & (x531x) & (!n_n4952) & (n_n4950) & (!n_n4937)) + ((!x20x) & (x531x) & (!n_n4952) & (n_n4950) & (n_n4937)) + ((!x20x) & (x531x) & (n_n4952) & (!n_n4950) & (!n_n4937)) + ((!x20x) & (x531x) & (n_n4952) & (!n_n4950) & (n_n4937)) + ((!x20x) & (x531x) & (n_n4952) & (n_n4950) & (!n_n4937)) + ((!x20x) & (x531x) & (n_n4952) & (n_n4950) & (n_n4937)) + ((x20x) & (!x531x) & (!n_n4952) & (!n_n4950) & (n_n4937)) + ((x20x) & (!x531x) & (!n_n4952) & (n_n4950) & (!n_n4937)) + ((x20x) & (!x531x) & (!n_n4952) & (n_n4950) & (n_n4937)) + ((x20x) & (!x531x) & (n_n4952) & (!n_n4950) & (!n_n4937)) + ((x20x) & (!x531x) & (n_n4952) & (!n_n4950) & (n_n4937)) + ((x20x) & (!x531x) & (n_n4952) & (n_n4950) & (!n_n4937)) + ((x20x) & (!x531x) & (n_n4952) & (n_n4950) & (n_n4937)) + ((x20x) & (x531x) & (!n_n4952) & (!n_n4950) & (!n_n4937)) + ((x20x) & (x531x) & (!n_n4952) & (!n_n4950) & (n_n4937)) + ((x20x) & (x531x) & (!n_n4952) & (n_n4950) & (!n_n4937)) + ((x20x) & (x531x) & (!n_n4952) & (n_n4950) & (n_n4937)) + ((x20x) & (x531x) & (n_n4952) & (!n_n4950) & (!n_n4937)) + ((x20x) & (x531x) & (n_n4952) & (!n_n4950) & (n_n4937)) + ((x20x) & (x531x) & (n_n4952) & (n_n4950) & (!n_n4937)) + ((x20x) & (x531x) & (n_n4952) & (n_n4950) & (n_n4937)));
	assign x14986x = (((!n_n4749) & (!n_n4751) & (!n_n4750) & (!n_n4742) & (n_n4753)) + ((!n_n4749) & (!n_n4751) & (!n_n4750) & (n_n4742) & (!n_n4753)) + ((!n_n4749) & (!n_n4751) & (!n_n4750) & (n_n4742) & (n_n4753)) + ((!n_n4749) & (!n_n4751) & (n_n4750) & (!n_n4742) & (!n_n4753)) + ((!n_n4749) & (!n_n4751) & (n_n4750) & (!n_n4742) & (n_n4753)) + ((!n_n4749) & (!n_n4751) & (n_n4750) & (n_n4742) & (!n_n4753)) + ((!n_n4749) & (!n_n4751) & (n_n4750) & (n_n4742) & (n_n4753)) + ((!n_n4749) & (n_n4751) & (!n_n4750) & (!n_n4742) & (!n_n4753)) + ((!n_n4749) & (n_n4751) & (!n_n4750) & (!n_n4742) & (n_n4753)) + ((!n_n4749) & (n_n4751) & (!n_n4750) & (n_n4742) & (!n_n4753)) + ((!n_n4749) & (n_n4751) & (!n_n4750) & (n_n4742) & (n_n4753)) + ((!n_n4749) & (n_n4751) & (n_n4750) & (!n_n4742) & (!n_n4753)) + ((!n_n4749) & (n_n4751) & (n_n4750) & (!n_n4742) & (n_n4753)) + ((!n_n4749) & (n_n4751) & (n_n4750) & (n_n4742) & (!n_n4753)) + ((!n_n4749) & (n_n4751) & (n_n4750) & (n_n4742) & (n_n4753)) + ((n_n4749) & (!n_n4751) & (!n_n4750) & (!n_n4742) & (!n_n4753)) + ((n_n4749) & (!n_n4751) & (!n_n4750) & (!n_n4742) & (n_n4753)) + ((n_n4749) & (!n_n4751) & (!n_n4750) & (n_n4742) & (!n_n4753)) + ((n_n4749) & (!n_n4751) & (!n_n4750) & (n_n4742) & (n_n4753)) + ((n_n4749) & (!n_n4751) & (n_n4750) & (!n_n4742) & (!n_n4753)) + ((n_n4749) & (!n_n4751) & (n_n4750) & (!n_n4742) & (n_n4753)) + ((n_n4749) & (!n_n4751) & (n_n4750) & (n_n4742) & (!n_n4753)) + ((n_n4749) & (!n_n4751) & (n_n4750) & (n_n4742) & (n_n4753)) + ((n_n4749) & (n_n4751) & (!n_n4750) & (!n_n4742) & (!n_n4753)) + ((n_n4749) & (n_n4751) & (!n_n4750) & (!n_n4742) & (n_n4753)) + ((n_n4749) & (n_n4751) & (!n_n4750) & (n_n4742) & (!n_n4753)) + ((n_n4749) & (n_n4751) & (!n_n4750) & (n_n4742) & (n_n4753)) + ((n_n4749) & (n_n4751) & (n_n4750) & (!n_n4742) & (!n_n4753)) + ((n_n4749) & (n_n4751) & (n_n4750) & (!n_n4742) & (n_n4753)) + ((n_n4749) & (n_n4751) & (n_n4750) & (n_n4742) & (!n_n4753)) + ((n_n4749) & (n_n4751) & (n_n4750) & (n_n4742) & (n_n4753)));
	assign x22092x = (((!n_n4755) & (!n_n4759) & (!n_n4767) & (!n_n4765)));
	assign n_n2614 = (((!n_n4669) & (!n_n4668) & (!n_n4671) & (!x80x) & (!x22091x)) + ((!n_n4669) & (!n_n4668) & (!n_n4671) & (x80x) & (!x22091x)) + ((!n_n4669) & (!n_n4668) & (!n_n4671) & (x80x) & (x22091x)) + ((!n_n4669) & (!n_n4668) & (n_n4671) & (!x80x) & (!x22091x)) + ((!n_n4669) & (!n_n4668) & (n_n4671) & (!x80x) & (x22091x)) + ((!n_n4669) & (!n_n4668) & (n_n4671) & (x80x) & (!x22091x)) + ((!n_n4669) & (!n_n4668) & (n_n4671) & (x80x) & (x22091x)) + ((!n_n4669) & (n_n4668) & (!n_n4671) & (!x80x) & (!x22091x)) + ((!n_n4669) & (n_n4668) & (!n_n4671) & (!x80x) & (x22091x)) + ((!n_n4669) & (n_n4668) & (!n_n4671) & (x80x) & (!x22091x)) + ((!n_n4669) & (n_n4668) & (!n_n4671) & (x80x) & (x22091x)) + ((!n_n4669) & (n_n4668) & (n_n4671) & (!x80x) & (!x22091x)) + ((!n_n4669) & (n_n4668) & (n_n4671) & (!x80x) & (x22091x)) + ((!n_n4669) & (n_n4668) & (n_n4671) & (x80x) & (!x22091x)) + ((!n_n4669) & (n_n4668) & (n_n4671) & (x80x) & (x22091x)) + ((n_n4669) & (!n_n4668) & (!n_n4671) & (!x80x) & (!x22091x)) + ((n_n4669) & (!n_n4668) & (!n_n4671) & (!x80x) & (x22091x)) + ((n_n4669) & (!n_n4668) & (!n_n4671) & (x80x) & (!x22091x)) + ((n_n4669) & (!n_n4668) & (!n_n4671) & (x80x) & (x22091x)) + ((n_n4669) & (!n_n4668) & (n_n4671) & (!x80x) & (!x22091x)) + ((n_n4669) & (!n_n4668) & (n_n4671) & (!x80x) & (x22091x)) + ((n_n4669) & (!n_n4668) & (n_n4671) & (x80x) & (!x22091x)) + ((n_n4669) & (!n_n4668) & (n_n4671) & (x80x) & (x22091x)) + ((n_n4669) & (n_n4668) & (!n_n4671) & (!x80x) & (!x22091x)) + ((n_n4669) & (n_n4668) & (!n_n4671) & (!x80x) & (x22091x)) + ((n_n4669) & (n_n4668) & (!n_n4671) & (x80x) & (!x22091x)) + ((n_n4669) & (n_n4668) & (!n_n4671) & (x80x) & (x22091x)) + ((n_n4669) & (n_n4668) & (n_n4671) & (!x80x) & (!x22091x)) + ((n_n4669) & (n_n4668) & (n_n4671) & (!x80x) & (x22091x)) + ((n_n4669) & (n_n4668) & (n_n4671) & (x80x) & (!x22091x)) + ((n_n4669) & (n_n4668) & (n_n4671) & (x80x) & (x22091x)));
	assign x15002x = (((!n_n4698) & (!n_n4680) & (!n_n4688) & (n_n4687)) + ((!n_n4698) & (!n_n4680) & (n_n4688) & (!n_n4687)) + ((!n_n4698) & (!n_n4680) & (n_n4688) & (n_n4687)) + ((!n_n4698) & (n_n4680) & (!n_n4688) & (!n_n4687)) + ((!n_n4698) & (n_n4680) & (!n_n4688) & (n_n4687)) + ((!n_n4698) & (n_n4680) & (n_n4688) & (!n_n4687)) + ((!n_n4698) & (n_n4680) & (n_n4688) & (n_n4687)) + ((n_n4698) & (!n_n4680) & (!n_n4688) & (!n_n4687)) + ((n_n4698) & (!n_n4680) & (!n_n4688) & (n_n4687)) + ((n_n4698) & (!n_n4680) & (n_n4688) & (!n_n4687)) + ((n_n4698) & (!n_n4680) & (n_n4688) & (n_n4687)) + ((n_n4698) & (n_n4680) & (!n_n4688) & (!n_n4687)) + ((n_n4698) & (n_n4680) & (!n_n4688) & (n_n4687)) + ((n_n4698) & (n_n4680) & (n_n4688) & (!n_n4687)) + ((n_n4698) & (n_n4680) & (n_n4688) & (n_n4687)));
	assign x15003x = (((!n_n4683) & (!x81x) & (!n_n4684) & (!x86x) & (n_n4694)) + ((!n_n4683) & (!x81x) & (!n_n4684) & (x86x) & (!n_n4694)) + ((!n_n4683) & (!x81x) & (!n_n4684) & (x86x) & (n_n4694)) + ((!n_n4683) & (!x81x) & (n_n4684) & (!x86x) & (!n_n4694)) + ((!n_n4683) & (!x81x) & (n_n4684) & (!x86x) & (n_n4694)) + ((!n_n4683) & (!x81x) & (n_n4684) & (x86x) & (!n_n4694)) + ((!n_n4683) & (!x81x) & (n_n4684) & (x86x) & (n_n4694)) + ((!n_n4683) & (x81x) & (!n_n4684) & (!x86x) & (!n_n4694)) + ((!n_n4683) & (x81x) & (!n_n4684) & (!x86x) & (n_n4694)) + ((!n_n4683) & (x81x) & (!n_n4684) & (x86x) & (!n_n4694)) + ((!n_n4683) & (x81x) & (!n_n4684) & (x86x) & (n_n4694)) + ((!n_n4683) & (x81x) & (n_n4684) & (!x86x) & (!n_n4694)) + ((!n_n4683) & (x81x) & (n_n4684) & (!x86x) & (n_n4694)) + ((!n_n4683) & (x81x) & (n_n4684) & (x86x) & (!n_n4694)) + ((!n_n4683) & (x81x) & (n_n4684) & (x86x) & (n_n4694)) + ((n_n4683) & (!x81x) & (!n_n4684) & (!x86x) & (!n_n4694)) + ((n_n4683) & (!x81x) & (!n_n4684) & (!x86x) & (n_n4694)) + ((n_n4683) & (!x81x) & (!n_n4684) & (x86x) & (!n_n4694)) + ((n_n4683) & (!x81x) & (!n_n4684) & (x86x) & (n_n4694)) + ((n_n4683) & (!x81x) & (n_n4684) & (!x86x) & (!n_n4694)) + ((n_n4683) & (!x81x) & (n_n4684) & (!x86x) & (n_n4694)) + ((n_n4683) & (!x81x) & (n_n4684) & (x86x) & (!n_n4694)) + ((n_n4683) & (!x81x) & (n_n4684) & (x86x) & (n_n4694)) + ((n_n4683) & (x81x) & (!n_n4684) & (!x86x) & (!n_n4694)) + ((n_n4683) & (x81x) & (!n_n4684) & (!x86x) & (n_n4694)) + ((n_n4683) & (x81x) & (!n_n4684) & (x86x) & (!n_n4694)) + ((n_n4683) & (x81x) & (!n_n4684) & (x86x) & (n_n4694)) + ((n_n4683) & (x81x) & (n_n4684) & (!x86x) & (!n_n4694)) + ((n_n4683) & (x81x) & (n_n4684) & (!x86x) & (n_n4694)) + ((n_n4683) & (x81x) & (n_n4684) & (x86x) & (!n_n4694)) + ((n_n4683) & (x81x) & (n_n4684) & (x86x) & (n_n4694)));
	assign x15004x = (((!n_n4691) & (!x219x) & (!x417x) & (!n_n4693) & (x442x)) + ((!n_n4691) & (!x219x) & (!x417x) & (n_n4693) & (!x442x)) + ((!n_n4691) & (!x219x) & (!x417x) & (n_n4693) & (x442x)) + ((!n_n4691) & (!x219x) & (x417x) & (!n_n4693) & (!x442x)) + ((!n_n4691) & (!x219x) & (x417x) & (!n_n4693) & (x442x)) + ((!n_n4691) & (!x219x) & (x417x) & (n_n4693) & (!x442x)) + ((!n_n4691) & (!x219x) & (x417x) & (n_n4693) & (x442x)) + ((!n_n4691) & (x219x) & (!x417x) & (!n_n4693) & (!x442x)) + ((!n_n4691) & (x219x) & (!x417x) & (!n_n4693) & (x442x)) + ((!n_n4691) & (x219x) & (!x417x) & (n_n4693) & (!x442x)) + ((!n_n4691) & (x219x) & (!x417x) & (n_n4693) & (x442x)) + ((!n_n4691) & (x219x) & (x417x) & (!n_n4693) & (!x442x)) + ((!n_n4691) & (x219x) & (x417x) & (!n_n4693) & (x442x)) + ((!n_n4691) & (x219x) & (x417x) & (n_n4693) & (!x442x)) + ((!n_n4691) & (x219x) & (x417x) & (n_n4693) & (x442x)) + ((n_n4691) & (!x219x) & (!x417x) & (!n_n4693) & (!x442x)) + ((n_n4691) & (!x219x) & (!x417x) & (!n_n4693) & (x442x)) + ((n_n4691) & (!x219x) & (!x417x) & (n_n4693) & (!x442x)) + ((n_n4691) & (!x219x) & (!x417x) & (n_n4693) & (x442x)) + ((n_n4691) & (!x219x) & (x417x) & (!n_n4693) & (!x442x)) + ((n_n4691) & (!x219x) & (x417x) & (!n_n4693) & (x442x)) + ((n_n4691) & (!x219x) & (x417x) & (n_n4693) & (!x442x)) + ((n_n4691) & (!x219x) & (x417x) & (n_n4693) & (x442x)) + ((n_n4691) & (x219x) & (!x417x) & (!n_n4693) & (!x442x)) + ((n_n4691) & (x219x) & (!x417x) & (!n_n4693) & (x442x)) + ((n_n4691) & (x219x) & (!x417x) & (n_n4693) & (!x442x)) + ((n_n4691) & (x219x) & (!x417x) & (n_n4693) & (x442x)) + ((n_n4691) & (x219x) & (x417x) & (!n_n4693) & (!x442x)) + ((n_n4691) & (x219x) & (x417x) & (!n_n4693) & (x442x)) + ((n_n4691) & (x219x) & (x417x) & (n_n4693) & (!x442x)) + ((n_n4691) & (x219x) & (x417x) & (n_n4693) & (x442x)));
	assign n_n2611 = (((!n_n4711) & (!n_n4705) & (!n_n4706) & (!n_n4707) & (x464x)) + ((!n_n4711) & (!n_n4705) & (!n_n4706) & (n_n4707) & (!x464x)) + ((!n_n4711) & (!n_n4705) & (!n_n4706) & (n_n4707) & (x464x)) + ((!n_n4711) & (!n_n4705) & (n_n4706) & (!n_n4707) & (!x464x)) + ((!n_n4711) & (!n_n4705) & (n_n4706) & (!n_n4707) & (x464x)) + ((!n_n4711) & (!n_n4705) & (n_n4706) & (n_n4707) & (!x464x)) + ((!n_n4711) & (!n_n4705) & (n_n4706) & (n_n4707) & (x464x)) + ((!n_n4711) & (n_n4705) & (!n_n4706) & (!n_n4707) & (!x464x)) + ((!n_n4711) & (n_n4705) & (!n_n4706) & (!n_n4707) & (x464x)) + ((!n_n4711) & (n_n4705) & (!n_n4706) & (n_n4707) & (!x464x)) + ((!n_n4711) & (n_n4705) & (!n_n4706) & (n_n4707) & (x464x)) + ((!n_n4711) & (n_n4705) & (n_n4706) & (!n_n4707) & (!x464x)) + ((!n_n4711) & (n_n4705) & (n_n4706) & (!n_n4707) & (x464x)) + ((!n_n4711) & (n_n4705) & (n_n4706) & (n_n4707) & (!x464x)) + ((!n_n4711) & (n_n4705) & (n_n4706) & (n_n4707) & (x464x)) + ((n_n4711) & (!n_n4705) & (!n_n4706) & (!n_n4707) & (!x464x)) + ((n_n4711) & (!n_n4705) & (!n_n4706) & (!n_n4707) & (x464x)) + ((n_n4711) & (!n_n4705) & (!n_n4706) & (n_n4707) & (!x464x)) + ((n_n4711) & (!n_n4705) & (!n_n4706) & (n_n4707) & (x464x)) + ((n_n4711) & (!n_n4705) & (n_n4706) & (!n_n4707) & (!x464x)) + ((n_n4711) & (!n_n4705) & (n_n4706) & (!n_n4707) & (x464x)) + ((n_n4711) & (!n_n4705) & (n_n4706) & (n_n4707) & (!x464x)) + ((n_n4711) & (!n_n4705) & (n_n4706) & (n_n4707) & (x464x)) + ((n_n4711) & (n_n4705) & (!n_n4706) & (!n_n4707) & (!x464x)) + ((n_n4711) & (n_n4705) & (!n_n4706) & (!n_n4707) & (x464x)) + ((n_n4711) & (n_n4705) & (!n_n4706) & (n_n4707) & (!x464x)) + ((n_n4711) & (n_n4705) & (!n_n4706) & (n_n4707) & (x464x)) + ((n_n4711) & (n_n4705) & (n_n4706) & (!n_n4707) & (!x464x)) + ((n_n4711) & (n_n4705) & (n_n4706) & (!n_n4707) & (x464x)) + ((n_n4711) & (n_n4705) & (n_n4706) & (n_n4707) & (!x464x)) + ((n_n4711) & (n_n4705) & (n_n4706) & (n_n4707) & (x464x)));
	assign x15013x = (((!n_n4720) & (!x241x) & (!n_n4716) & (n_n4713)) + ((!n_n4720) & (!x241x) & (n_n4716) & (!n_n4713)) + ((!n_n4720) & (!x241x) & (n_n4716) & (n_n4713)) + ((!n_n4720) & (x241x) & (!n_n4716) & (!n_n4713)) + ((!n_n4720) & (x241x) & (!n_n4716) & (n_n4713)) + ((!n_n4720) & (x241x) & (n_n4716) & (!n_n4713)) + ((!n_n4720) & (x241x) & (n_n4716) & (n_n4713)) + ((n_n4720) & (!x241x) & (!n_n4716) & (!n_n4713)) + ((n_n4720) & (!x241x) & (!n_n4716) & (n_n4713)) + ((n_n4720) & (!x241x) & (n_n4716) & (!n_n4713)) + ((n_n4720) & (!x241x) & (n_n4716) & (n_n4713)) + ((n_n4720) & (x241x) & (!n_n4716) & (!n_n4713)) + ((n_n4720) & (x241x) & (!n_n4716) & (n_n4713)) + ((n_n4720) & (x241x) & (n_n4716) & (!n_n4713)) + ((n_n4720) & (x241x) & (n_n4716) & (n_n4713)));
	assign x15014x = (((!n_n4727) & (!n_n4726) & (!n_n4728) & (n_n856)) + ((!n_n4727) & (!n_n4726) & (n_n4728) & (!n_n856)) + ((!n_n4727) & (!n_n4726) & (n_n4728) & (n_n856)) + ((!n_n4727) & (n_n4726) & (!n_n4728) & (!n_n856)) + ((!n_n4727) & (n_n4726) & (!n_n4728) & (n_n856)) + ((!n_n4727) & (n_n4726) & (n_n4728) & (!n_n856)) + ((!n_n4727) & (n_n4726) & (n_n4728) & (n_n856)) + ((n_n4727) & (!n_n4726) & (!n_n4728) & (!n_n856)) + ((n_n4727) & (!n_n4726) & (!n_n4728) & (n_n856)) + ((n_n4727) & (!n_n4726) & (n_n4728) & (!n_n856)) + ((n_n4727) & (!n_n4726) & (n_n4728) & (n_n856)) + ((n_n4727) & (n_n4726) & (!n_n4728) & (!n_n856)) + ((n_n4727) & (n_n4726) & (!n_n4728) & (n_n856)) + ((n_n4727) & (n_n4726) & (n_n4728) & (!n_n856)) + ((n_n4727) & (n_n4726) & (n_n4728) & (n_n856)));
	assign x15015x = (((!n_n4712) & (!n_n4736) & (!x94x) & (!x39x) & (n_n4723)) + ((!n_n4712) & (!n_n4736) & (!x94x) & (x39x) & (!n_n4723)) + ((!n_n4712) & (!n_n4736) & (!x94x) & (x39x) & (n_n4723)) + ((!n_n4712) & (!n_n4736) & (x94x) & (!x39x) & (!n_n4723)) + ((!n_n4712) & (!n_n4736) & (x94x) & (!x39x) & (n_n4723)) + ((!n_n4712) & (!n_n4736) & (x94x) & (x39x) & (!n_n4723)) + ((!n_n4712) & (!n_n4736) & (x94x) & (x39x) & (n_n4723)) + ((!n_n4712) & (n_n4736) & (!x94x) & (!x39x) & (!n_n4723)) + ((!n_n4712) & (n_n4736) & (!x94x) & (!x39x) & (n_n4723)) + ((!n_n4712) & (n_n4736) & (!x94x) & (x39x) & (!n_n4723)) + ((!n_n4712) & (n_n4736) & (!x94x) & (x39x) & (n_n4723)) + ((!n_n4712) & (n_n4736) & (x94x) & (!x39x) & (!n_n4723)) + ((!n_n4712) & (n_n4736) & (x94x) & (!x39x) & (n_n4723)) + ((!n_n4712) & (n_n4736) & (x94x) & (x39x) & (!n_n4723)) + ((!n_n4712) & (n_n4736) & (x94x) & (x39x) & (n_n4723)) + ((n_n4712) & (!n_n4736) & (!x94x) & (!x39x) & (!n_n4723)) + ((n_n4712) & (!n_n4736) & (!x94x) & (!x39x) & (n_n4723)) + ((n_n4712) & (!n_n4736) & (!x94x) & (x39x) & (!n_n4723)) + ((n_n4712) & (!n_n4736) & (!x94x) & (x39x) & (n_n4723)) + ((n_n4712) & (!n_n4736) & (x94x) & (!x39x) & (!n_n4723)) + ((n_n4712) & (!n_n4736) & (x94x) & (!x39x) & (n_n4723)) + ((n_n4712) & (!n_n4736) & (x94x) & (x39x) & (!n_n4723)) + ((n_n4712) & (!n_n4736) & (x94x) & (x39x) & (n_n4723)) + ((n_n4712) & (n_n4736) & (!x94x) & (!x39x) & (!n_n4723)) + ((n_n4712) & (n_n4736) & (!x94x) & (!x39x) & (n_n4723)) + ((n_n4712) & (n_n4736) & (!x94x) & (x39x) & (!n_n4723)) + ((n_n4712) & (n_n4736) & (!x94x) & (x39x) & (n_n4723)) + ((n_n4712) & (n_n4736) & (x94x) & (!x39x) & (!n_n4723)) + ((n_n4712) & (n_n4736) & (x94x) & (!x39x) & (n_n4723)) + ((n_n4712) & (n_n4736) & (x94x) & (x39x) & (!n_n4723)) + ((n_n4712) & (n_n4736) & (x94x) & (x39x) & (n_n4723)));
	assign n_n5118 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n509) & (x12x)));
	assign n_n5119 = (((!i_9_) & (n_n528) & (n_n509) & (n_n130)));
	assign n_n5229 = (((!i_9_) & (n_n518) & (n_n530) & (n_n65)));
	assign n_n5228 = (((!i_5_) & (i_3_) & (i_4_) & (x19x) & (n_n530)));
	assign n_n5295 = (((!i_9_) & (n_n482) & (n_n528) & (n_n65)));
	assign n_n4540 = (((i_9_) & (n_n455) & (n_n473) & (n_n530)));
	assign n_n889 = (((!i_7_) & (i_8_) & (i_6_) & (x13x) & (n_n473)) + ((i_7_) & (!i_8_) & (i_6_) & (x13x) & (n_n473)) + ((i_7_) & (i_8_) & (i_6_) & (x13x) & (n_n473)));
	assign n_n4541 = (((!i_9_) & (n_n455) & (n_n473) & (n_n530)));
	assign n_n4543 = (((!i_9_) & (n_n455) & (n_n528) & (n_n473)));
	assign x22208x = (((!n_n4542) & (!n_n889) & (!n_n4532) & (!n_n4541) & (!n_n4543)));
	assign n_n4681 = (((!i_9_) & (n_n390) & (n_n534) & (n_n464)));
	assign n_n4679 = (((!i_1_) & (i_2_) & (i_0_) & (n_n473) & (x23x)));
	assign n_n4677 = (((!i_1_) & (i_2_) & (i_0_) & (n_n473) & (x20x)));
	assign n_n4678 = (((i_9_) & (n_n390) & (n_n473) & (n_n520)));
	assign x81x = (((i_9_) & (n_n390) & (n_n532) & (n_n464)));
	assign x338x = (((!i_9_) & (!n_n528) & (n_n390) & (n_n473) & (n_n530)) + ((!i_9_) & (n_n528) & (n_n390) & (n_n473) & (n_n530)) + ((i_9_) & (n_n528) & (n_n390) & (n_n473) & (!n_n530)) + ((i_9_) & (n_n528) & (n_n390) & (n_n473) & (n_n530)));
	assign x16406x = (((!n_n4669) & (!n_n4670) & (!n_n4677) & (!n_n4678) & (x81x)) + ((!n_n4669) & (!n_n4670) & (!n_n4677) & (n_n4678) & (!x81x)) + ((!n_n4669) & (!n_n4670) & (!n_n4677) & (n_n4678) & (x81x)) + ((!n_n4669) & (!n_n4670) & (n_n4677) & (!n_n4678) & (!x81x)) + ((!n_n4669) & (!n_n4670) & (n_n4677) & (!n_n4678) & (x81x)) + ((!n_n4669) & (!n_n4670) & (n_n4677) & (n_n4678) & (!x81x)) + ((!n_n4669) & (!n_n4670) & (n_n4677) & (n_n4678) & (x81x)) + ((!n_n4669) & (n_n4670) & (!n_n4677) & (!n_n4678) & (!x81x)) + ((!n_n4669) & (n_n4670) & (!n_n4677) & (!n_n4678) & (x81x)) + ((!n_n4669) & (n_n4670) & (!n_n4677) & (n_n4678) & (!x81x)) + ((!n_n4669) & (n_n4670) & (!n_n4677) & (n_n4678) & (x81x)) + ((!n_n4669) & (n_n4670) & (n_n4677) & (!n_n4678) & (!x81x)) + ((!n_n4669) & (n_n4670) & (n_n4677) & (!n_n4678) & (x81x)) + ((!n_n4669) & (n_n4670) & (n_n4677) & (n_n4678) & (!x81x)) + ((!n_n4669) & (n_n4670) & (n_n4677) & (n_n4678) & (x81x)) + ((n_n4669) & (!n_n4670) & (!n_n4677) & (!n_n4678) & (!x81x)) + ((n_n4669) & (!n_n4670) & (!n_n4677) & (!n_n4678) & (x81x)) + ((n_n4669) & (!n_n4670) & (!n_n4677) & (n_n4678) & (!x81x)) + ((n_n4669) & (!n_n4670) & (!n_n4677) & (n_n4678) & (x81x)) + ((n_n4669) & (!n_n4670) & (n_n4677) & (!n_n4678) & (!x81x)) + ((n_n4669) & (!n_n4670) & (n_n4677) & (!n_n4678) & (x81x)) + ((n_n4669) & (!n_n4670) & (n_n4677) & (n_n4678) & (!x81x)) + ((n_n4669) & (!n_n4670) & (n_n4677) & (n_n4678) & (x81x)) + ((n_n4669) & (n_n4670) & (!n_n4677) & (!n_n4678) & (!x81x)) + ((n_n4669) & (n_n4670) & (!n_n4677) & (!n_n4678) & (x81x)) + ((n_n4669) & (n_n4670) & (!n_n4677) & (n_n4678) & (!x81x)) + ((n_n4669) & (n_n4670) & (!n_n4677) & (n_n4678) & (x81x)) + ((n_n4669) & (n_n4670) & (n_n4677) & (!n_n4678) & (!x81x)) + ((n_n4669) & (n_n4670) & (n_n4677) & (!n_n4678) & (x81x)) + ((n_n4669) & (n_n4670) & (n_n4677) & (n_n4678) & (!x81x)) + ((n_n4669) & (n_n4670) & (n_n4677) & (n_n4678) & (x81x)));
	assign x127x = (((!n_n518) & (n_n534) & (n_n509) & (!n_n520) & (x12x)) + ((!n_n518) & (n_n534) & (n_n509) & (n_n520) & (x12x)) + ((n_n518) & (!n_n534) & (!n_n509) & (n_n520) & (x12x)) + ((n_n518) & (!n_n534) & (n_n509) & (n_n520) & (x12x)) + ((n_n518) & (n_n534) & (!n_n509) & (n_n520) & (x12x)) + ((n_n518) & (n_n534) & (n_n509) & (!n_n520) & (x12x)) + ((n_n518) & (n_n534) & (n_n509) & (n_n520) & (x12x)));
	assign x414x = (((!i_9_) & (n_n528) & (n_n509) & (!n_n130) & (x12x)) + ((!i_9_) & (n_n528) & (n_n509) & (n_n130) & (!x12x)) + ((!i_9_) & (n_n528) & (n_n509) & (n_n130) & (x12x)) + ((i_9_) & (n_n528) & (n_n509) & (!n_n130) & (x12x)) + ((i_9_) & (n_n528) & (n_n509) & (n_n130) & (x12x)));
	assign x16724x = (((!n_n5112) & (!n_n5110) & (!n_n5114) & (!n_n5116) & (n_n5115)) + ((!n_n5112) & (!n_n5110) & (!n_n5114) & (n_n5116) & (!n_n5115)) + ((!n_n5112) & (!n_n5110) & (!n_n5114) & (n_n5116) & (n_n5115)) + ((!n_n5112) & (!n_n5110) & (n_n5114) & (!n_n5116) & (!n_n5115)) + ((!n_n5112) & (!n_n5110) & (n_n5114) & (!n_n5116) & (n_n5115)) + ((!n_n5112) & (!n_n5110) & (n_n5114) & (n_n5116) & (!n_n5115)) + ((!n_n5112) & (!n_n5110) & (n_n5114) & (n_n5116) & (n_n5115)) + ((!n_n5112) & (n_n5110) & (!n_n5114) & (!n_n5116) & (!n_n5115)) + ((!n_n5112) & (n_n5110) & (!n_n5114) & (!n_n5116) & (n_n5115)) + ((!n_n5112) & (n_n5110) & (!n_n5114) & (n_n5116) & (!n_n5115)) + ((!n_n5112) & (n_n5110) & (!n_n5114) & (n_n5116) & (n_n5115)) + ((!n_n5112) & (n_n5110) & (n_n5114) & (!n_n5116) & (!n_n5115)) + ((!n_n5112) & (n_n5110) & (n_n5114) & (!n_n5116) & (n_n5115)) + ((!n_n5112) & (n_n5110) & (n_n5114) & (n_n5116) & (!n_n5115)) + ((!n_n5112) & (n_n5110) & (n_n5114) & (n_n5116) & (n_n5115)) + ((n_n5112) & (!n_n5110) & (!n_n5114) & (!n_n5116) & (!n_n5115)) + ((n_n5112) & (!n_n5110) & (!n_n5114) & (!n_n5116) & (n_n5115)) + ((n_n5112) & (!n_n5110) & (!n_n5114) & (n_n5116) & (!n_n5115)) + ((n_n5112) & (!n_n5110) & (!n_n5114) & (n_n5116) & (n_n5115)) + ((n_n5112) & (!n_n5110) & (n_n5114) & (!n_n5116) & (!n_n5115)) + ((n_n5112) & (!n_n5110) & (n_n5114) & (!n_n5116) & (n_n5115)) + ((n_n5112) & (!n_n5110) & (n_n5114) & (n_n5116) & (!n_n5115)) + ((n_n5112) & (!n_n5110) & (n_n5114) & (n_n5116) & (n_n5115)) + ((n_n5112) & (n_n5110) & (!n_n5114) & (!n_n5116) & (!n_n5115)) + ((n_n5112) & (n_n5110) & (!n_n5114) & (!n_n5116) & (n_n5115)) + ((n_n5112) & (n_n5110) & (!n_n5114) & (n_n5116) & (!n_n5115)) + ((n_n5112) & (n_n5110) & (!n_n5114) & (n_n5116) & (n_n5115)) + ((n_n5112) & (n_n5110) & (n_n5114) & (!n_n5116) & (!n_n5115)) + ((n_n5112) & (n_n5110) & (n_n5114) & (!n_n5116) & (n_n5115)) + ((n_n5112) & (n_n5110) & (n_n5114) & (n_n5116) & (!n_n5115)) + ((n_n5112) & (n_n5110) & (n_n5114) & (n_n5116) & (n_n5115)));
	assign n_n2209 = (((!n_n5111) & (!n_n5113) & (!n_n5118) & (!n_n5119) & (x16724x)) + ((!n_n5111) & (!n_n5113) & (!n_n5118) & (n_n5119) & (!x16724x)) + ((!n_n5111) & (!n_n5113) & (!n_n5118) & (n_n5119) & (x16724x)) + ((!n_n5111) & (!n_n5113) & (n_n5118) & (!n_n5119) & (!x16724x)) + ((!n_n5111) & (!n_n5113) & (n_n5118) & (!n_n5119) & (x16724x)) + ((!n_n5111) & (!n_n5113) & (n_n5118) & (n_n5119) & (!x16724x)) + ((!n_n5111) & (!n_n5113) & (n_n5118) & (n_n5119) & (x16724x)) + ((!n_n5111) & (n_n5113) & (!n_n5118) & (!n_n5119) & (!x16724x)) + ((!n_n5111) & (n_n5113) & (!n_n5118) & (!n_n5119) & (x16724x)) + ((!n_n5111) & (n_n5113) & (!n_n5118) & (n_n5119) & (!x16724x)) + ((!n_n5111) & (n_n5113) & (!n_n5118) & (n_n5119) & (x16724x)) + ((!n_n5111) & (n_n5113) & (n_n5118) & (!n_n5119) & (!x16724x)) + ((!n_n5111) & (n_n5113) & (n_n5118) & (!n_n5119) & (x16724x)) + ((!n_n5111) & (n_n5113) & (n_n5118) & (n_n5119) & (!x16724x)) + ((!n_n5111) & (n_n5113) & (n_n5118) & (n_n5119) & (x16724x)) + ((n_n5111) & (!n_n5113) & (!n_n5118) & (!n_n5119) & (!x16724x)) + ((n_n5111) & (!n_n5113) & (!n_n5118) & (!n_n5119) & (x16724x)) + ((n_n5111) & (!n_n5113) & (!n_n5118) & (n_n5119) & (!x16724x)) + ((n_n5111) & (!n_n5113) & (!n_n5118) & (n_n5119) & (x16724x)) + ((n_n5111) & (!n_n5113) & (n_n5118) & (!n_n5119) & (!x16724x)) + ((n_n5111) & (!n_n5113) & (n_n5118) & (!n_n5119) & (x16724x)) + ((n_n5111) & (!n_n5113) & (n_n5118) & (n_n5119) & (!x16724x)) + ((n_n5111) & (!n_n5113) & (n_n5118) & (n_n5119) & (x16724x)) + ((n_n5111) & (n_n5113) & (!n_n5118) & (!n_n5119) & (!x16724x)) + ((n_n5111) & (n_n5113) & (!n_n5118) & (!n_n5119) & (x16724x)) + ((n_n5111) & (n_n5113) & (!n_n5118) & (n_n5119) & (!x16724x)) + ((n_n5111) & (n_n5113) & (!n_n5118) & (n_n5119) & (x16724x)) + ((n_n5111) & (n_n5113) & (n_n5118) & (!n_n5119) & (!x16724x)) + ((n_n5111) & (n_n5113) & (n_n5118) & (!n_n5119) & (x16724x)) + ((n_n5111) & (n_n5113) & (n_n5118) & (n_n5119) & (!x16724x)) + ((n_n5111) & (n_n5113) & (n_n5118) & (n_n5119) & (x16724x)));
	assign n_n4893 = (((!i_9_) & (n_n260) & (n_n491) & (n_n530)));
	assign x154x = (((!i_9_) & (n_n482) & (n_n532) & (n_n260)) + ((i_9_) & (n_n482) & (n_n532) & (n_n260)));
	assign x16785x = (((!n_n4865) & (!n_n4905) & (!n_n4893) & (x154x)) + ((!n_n4865) & (!n_n4905) & (n_n4893) & (!x154x)) + ((!n_n4865) & (!n_n4905) & (n_n4893) & (x154x)) + ((!n_n4865) & (n_n4905) & (!n_n4893) & (!x154x)) + ((!n_n4865) & (n_n4905) & (!n_n4893) & (x154x)) + ((!n_n4865) & (n_n4905) & (n_n4893) & (!x154x)) + ((!n_n4865) & (n_n4905) & (n_n4893) & (x154x)) + ((n_n4865) & (!n_n4905) & (!n_n4893) & (!x154x)) + ((n_n4865) & (!n_n4905) & (!n_n4893) & (x154x)) + ((n_n4865) & (!n_n4905) & (n_n4893) & (!x154x)) + ((n_n4865) & (!n_n4905) & (n_n4893) & (x154x)) + ((n_n4865) & (n_n4905) & (!n_n4893) & (!x154x)) + ((n_n4865) & (n_n4905) & (!n_n4893) & (x154x)) + ((n_n4865) & (n_n4905) & (n_n4893) & (!x154x)) + ((n_n4865) & (n_n4905) & (n_n4893) & (x154x)));
	assign n_n2095 = (((!n_n4902) & (!n_n4856) & (!n_n4854) & (!n_n4894) & (x16785x)) + ((!n_n4902) & (!n_n4856) & (!n_n4854) & (n_n4894) & (!x16785x)) + ((!n_n4902) & (!n_n4856) & (!n_n4854) & (n_n4894) & (x16785x)) + ((!n_n4902) & (!n_n4856) & (n_n4854) & (!n_n4894) & (!x16785x)) + ((!n_n4902) & (!n_n4856) & (n_n4854) & (!n_n4894) & (x16785x)) + ((!n_n4902) & (!n_n4856) & (n_n4854) & (n_n4894) & (!x16785x)) + ((!n_n4902) & (!n_n4856) & (n_n4854) & (n_n4894) & (x16785x)) + ((!n_n4902) & (n_n4856) & (!n_n4854) & (!n_n4894) & (!x16785x)) + ((!n_n4902) & (n_n4856) & (!n_n4854) & (!n_n4894) & (x16785x)) + ((!n_n4902) & (n_n4856) & (!n_n4854) & (n_n4894) & (!x16785x)) + ((!n_n4902) & (n_n4856) & (!n_n4854) & (n_n4894) & (x16785x)) + ((!n_n4902) & (n_n4856) & (n_n4854) & (!n_n4894) & (!x16785x)) + ((!n_n4902) & (n_n4856) & (n_n4854) & (!n_n4894) & (x16785x)) + ((!n_n4902) & (n_n4856) & (n_n4854) & (n_n4894) & (!x16785x)) + ((!n_n4902) & (n_n4856) & (n_n4854) & (n_n4894) & (x16785x)) + ((n_n4902) & (!n_n4856) & (!n_n4854) & (!n_n4894) & (!x16785x)) + ((n_n4902) & (!n_n4856) & (!n_n4854) & (!n_n4894) & (x16785x)) + ((n_n4902) & (!n_n4856) & (!n_n4854) & (n_n4894) & (!x16785x)) + ((n_n4902) & (!n_n4856) & (!n_n4854) & (n_n4894) & (x16785x)) + ((n_n4902) & (!n_n4856) & (n_n4854) & (!n_n4894) & (!x16785x)) + ((n_n4902) & (!n_n4856) & (n_n4854) & (!n_n4894) & (x16785x)) + ((n_n4902) & (!n_n4856) & (n_n4854) & (n_n4894) & (!x16785x)) + ((n_n4902) & (!n_n4856) & (n_n4854) & (n_n4894) & (x16785x)) + ((n_n4902) & (n_n4856) & (!n_n4854) & (!n_n4894) & (!x16785x)) + ((n_n4902) & (n_n4856) & (!n_n4854) & (!n_n4894) & (x16785x)) + ((n_n4902) & (n_n4856) & (!n_n4854) & (n_n4894) & (!x16785x)) + ((n_n4902) & (n_n4856) & (!n_n4854) & (n_n4894) & (x16785x)) + ((n_n4902) & (n_n4856) & (n_n4854) & (!n_n4894) & (!x16785x)) + ((n_n4902) & (n_n4856) & (n_n4854) & (!n_n4894) & (x16785x)) + ((n_n4902) & (n_n4856) & (n_n4854) & (n_n4894) & (!x16785x)) + ((n_n4902) & (n_n4856) & (n_n4854) & (n_n4894) & (x16785x)));
	assign n_n5168 = (((i_7_) & (i_8_) & (!i_6_) & (n_n482) & (x12x)));
	assign x126x = (((!n_n520) & (n_n130) & (!x12x) & (x20x) & (n_n500)) + ((!n_n520) & (n_n130) & (x12x) & (x20x) & (n_n500)) + ((n_n520) & (!n_n130) & (x12x) & (!x20x) & (n_n500)) + ((n_n520) & (!n_n130) & (x12x) & (x20x) & (n_n500)) + ((n_n520) & (n_n130) & (!x12x) & (x20x) & (n_n500)) + ((n_n520) & (n_n130) & (x12x) & (!x20x) & (n_n500)) + ((n_n520) & (n_n130) & (x12x) & (x20x) & (n_n500)));
	assign x16804x = (((!n_n4975) & (!n_n4991) & (!n_n5000) & (!n_n4973) & (n_n4957)) + ((!n_n4975) & (!n_n4991) & (!n_n5000) & (n_n4973) & (!n_n4957)) + ((!n_n4975) & (!n_n4991) & (!n_n5000) & (n_n4973) & (n_n4957)) + ((!n_n4975) & (!n_n4991) & (n_n5000) & (!n_n4973) & (!n_n4957)) + ((!n_n4975) & (!n_n4991) & (n_n5000) & (!n_n4973) & (n_n4957)) + ((!n_n4975) & (!n_n4991) & (n_n5000) & (n_n4973) & (!n_n4957)) + ((!n_n4975) & (!n_n4991) & (n_n5000) & (n_n4973) & (n_n4957)) + ((!n_n4975) & (n_n4991) & (!n_n5000) & (!n_n4973) & (!n_n4957)) + ((!n_n4975) & (n_n4991) & (!n_n5000) & (!n_n4973) & (n_n4957)) + ((!n_n4975) & (n_n4991) & (!n_n5000) & (n_n4973) & (!n_n4957)) + ((!n_n4975) & (n_n4991) & (!n_n5000) & (n_n4973) & (n_n4957)) + ((!n_n4975) & (n_n4991) & (n_n5000) & (!n_n4973) & (!n_n4957)) + ((!n_n4975) & (n_n4991) & (n_n5000) & (!n_n4973) & (n_n4957)) + ((!n_n4975) & (n_n4991) & (n_n5000) & (n_n4973) & (!n_n4957)) + ((!n_n4975) & (n_n4991) & (n_n5000) & (n_n4973) & (n_n4957)) + ((n_n4975) & (!n_n4991) & (!n_n5000) & (!n_n4973) & (!n_n4957)) + ((n_n4975) & (!n_n4991) & (!n_n5000) & (!n_n4973) & (n_n4957)) + ((n_n4975) & (!n_n4991) & (!n_n5000) & (n_n4973) & (!n_n4957)) + ((n_n4975) & (!n_n4991) & (!n_n5000) & (n_n4973) & (n_n4957)) + ((n_n4975) & (!n_n4991) & (n_n5000) & (!n_n4973) & (!n_n4957)) + ((n_n4975) & (!n_n4991) & (n_n5000) & (!n_n4973) & (n_n4957)) + ((n_n4975) & (!n_n4991) & (n_n5000) & (n_n4973) & (!n_n4957)) + ((n_n4975) & (!n_n4991) & (n_n5000) & (n_n4973) & (n_n4957)) + ((n_n4975) & (n_n4991) & (!n_n5000) & (!n_n4973) & (!n_n4957)) + ((n_n4975) & (n_n4991) & (!n_n5000) & (!n_n4973) & (n_n4957)) + ((n_n4975) & (n_n4991) & (!n_n5000) & (n_n4973) & (!n_n4957)) + ((n_n4975) & (n_n4991) & (!n_n5000) & (n_n4973) & (n_n4957)) + ((n_n4975) & (n_n4991) & (n_n5000) & (!n_n4973) & (!n_n4957)) + ((n_n4975) & (n_n4991) & (n_n5000) & (!n_n4973) & (n_n4957)) + ((n_n4975) & (n_n4991) & (n_n5000) & (n_n4973) & (!n_n4957)) + ((n_n4975) & (n_n4991) & (n_n5000) & (n_n4973) & (n_n4957)));
	assign n_n4709 = (((!i_1_) & (!i_2_) & (i_0_) & (n_n535) & (x20x)));
	assign x14962x = (((!i_9_) & (n_n524) & (n_n260) & (n_n464)) + ((i_9_) & (n_n524) & (n_n260) & (n_n464)));
	assign n_n4603 = (((!i_9_) & (n_n390) & (n_n532) & (n_n509)));
	assign n_n2037 = (((!x10x) & (!n_n534) & (!n_n509) & (!n_n530) & (n_n4603)) + ((!x10x) & (!n_n534) & (!n_n509) & (n_n530) & (n_n4603)) + ((!x10x) & (!n_n534) & (n_n509) & (!n_n530) & (n_n4603)) + ((!x10x) & (!n_n534) & (n_n509) & (n_n530) & (n_n4603)) + ((!x10x) & (n_n534) & (!n_n509) & (!n_n530) & (n_n4603)) + ((!x10x) & (n_n534) & (!n_n509) & (n_n530) & (n_n4603)) + ((!x10x) & (n_n534) & (n_n509) & (!n_n530) & (n_n4603)) + ((!x10x) & (n_n534) & (n_n509) & (n_n530) & (n_n4603)) + ((x10x) & (!n_n534) & (!n_n509) & (!n_n530) & (n_n4603)) + ((x10x) & (!n_n534) & (!n_n509) & (n_n530) & (n_n4603)) + ((x10x) & (!n_n534) & (n_n509) & (!n_n530) & (n_n4603)) + ((x10x) & (!n_n534) & (n_n509) & (n_n530) & (!n_n4603)) + ((x10x) & (!n_n534) & (n_n509) & (n_n530) & (n_n4603)) + ((x10x) & (n_n534) & (!n_n509) & (!n_n530) & (n_n4603)) + ((x10x) & (n_n534) & (!n_n509) & (n_n530) & (n_n4603)) + ((x10x) & (n_n534) & (n_n509) & (!n_n530) & (!n_n4603)) + ((x10x) & (n_n534) & (n_n509) & (!n_n530) & (n_n4603)) + ((x10x) & (n_n534) & (n_n509) & (n_n530) & (!n_n4603)) + ((x10x) & (n_n534) & (n_n509) & (n_n530) & (n_n4603)));
	assign x12311x = (((!x120x) & (!n_n5058) & (!n_n5067) & (n_n5061)) + ((!x120x) & (!n_n5058) & (n_n5067) & (!n_n5061)) + ((!x120x) & (!n_n5058) & (n_n5067) & (n_n5061)) + ((!x120x) & (n_n5058) & (!n_n5067) & (!n_n5061)) + ((!x120x) & (n_n5058) & (!n_n5067) & (n_n5061)) + ((!x120x) & (n_n5058) & (n_n5067) & (!n_n5061)) + ((!x120x) & (n_n5058) & (n_n5067) & (n_n5061)) + ((x120x) & (!n_n5058) & (!n_n5067) & (!n_n5061)) + ((x120x) & (!n_n5058) & (!n_n5067) & (n_n5061)) + ((x120x) & (!n_n5058) & (n_n5067) & (!n_n5061)) + ((x120x) & (!n_n5058) & (n_n5067) & (n_n5061)) + ((x120x) & (n_n5058) & (!n_n5067) & (!n_n5061)) + ((x120x) & (n_n5058) & (!n_n5067) & (n_n5061)) + ((x120x) & (n_n5058) & (n_n5067) & (!n_n5061)) + ((x120x) & (n_n5058) & (n_n5067) & (n_n5061)));
	assign n_n5159 = (((i_5_) & (!i_3_) & (i_4_) & (n_n130) & (x23x)));
	assign x195x = (((n_n491) & (!n_n520) & (n_n130) & (!x12x) & (x23x)) + ((n_n491) & (!n_n520) & (n_n130) & (x12x) & (x23x)) + ((n_n491) & (n_n520) & (!n_n130) & (x12x) & (!x23x)) + ((n_n491) & (n_n520) & (!n_n130) & (x12x) & (x23x)) + ((n_n491) & (n_n520) & (n_n130) & (!x12x) & (x23x)) + ((n_n491) & (n_n520) & (n_n130) & (x12x) & (!x23x)) + ((n_n491) & (n_n520) & (n_n130) & (x12x) & (x23x)));
	assign x358x = (((!i_9_) & (n_n524) & (n_n491) & (!n_n130) & (x12x)) + ((!i_9_) & (n_n524) & (n_n491) & (n_n130) & (!x12x)) + ((!i_9_) & (n_n524) & (n_n491) & (n_n130) & (x12x)) + ((i_9_) & (n_n524) & (n_n491) & (!n_n130) & (x12x)) + ((i_9_) & (n_n524) & (n_n491) & (n_n130) & (x12x)));
	assign n_n5151 = (((!i_9_) & (n_n528) & (n_n491) & (n_n130)));
	assign x406x = (((!i_9_) & (n_n528) & (n_n491) & (!n_n130) & (x12x)) + ((!i_9_) & (n_n528) & (n_n491) & (n_n130) & (!x12x)) + ((!i_9_) & (n_n528) & (n_n491) & (n_n130) & (x12x)) + ((i_9_) & (n_n528) & (n_n491) & (!n_n130) & (x12x)) + ((i_9_) & (n_n528) & (n_n491) & (n_n130) & (x12x)));
	assign x12261x = (((!x21x) & (!n_n491) & (!n_n130) & (!n_n5154) & (x406x)) + ((!x21x) & (!n_n491) & (!n_n130) & (n_n5154) & (!x406x)) + ((!x21x) & (!n_n491) & (!n_n130) & (n_n5154) & (x406x)) + ((!x21x) & (!n_n491) & (n_n130) & (!n_n5154) & (x406x)) + ((!x21x) & (!n_n491) & (n_n130) & (n_n5154) & (!x406x)) + ((!x21x) & (!n_n491) & (n_n130) & (n_n5154) & (x406x)) + ((!x21x) & (n_n491) & (!n_n130) & (!n_n5154) & (x406x)) + ((!x21x) & (n_n491) & (!n_n130) & (n_n5154) & (!x406x)) + ((!x21x) & (n_n491) & (!n_n130) & (n_n5154) & (x406x)) + ((!x21x) & (n_n491) & (n_n130) & (!n_n5154) & (x406x)) + ((!x21x) & (n_n491) & (n_n130) & (n_n5154) & (!x406x)) + ((!x21x) & (n_n491) & (n_n130) & (n_n5154) & (x406x)) + ((x21x) & (!n_n491) & (!n_n130) & (!n_n5154) & (x406x)) + ((x21x) & (!n_n491) & (!n_n130) & (n_n5154) & (!x406x)) + ((x21x) & (!n_n491) & (!n_n130) & (n_n5154) & (x406x)) + ((x21x) & (!n_n491) & (n_n130) & (!n_n5154) & (x406x)) + ((x21x) & (!n_n491) & (n_n130) & (n_n5154) & (!x406x)) + ((x21x) & (!n_n491) & (n_n130) & (n_n5154) & (x406x)) + ((x21x) & (n_n491) & (!n_n130) & (!n_n5154) & (x406x)) + ((x21x) & (n_n491) & (!n_n130) & (n_n5154) & (!x406x)) + ((x21x) & (n_n491) & (!n_n130) & (n_n5154) & (x406x)) + ((x21x) & (n_n491) & (n_n130) & (!n_n5154) & (!x406x)) + ((x21x) & (n_n491) & (n_n130) & (!n_n5154) & (x406x)) + ((x21x) & (n_n491) & (n_n130) & (n_n5154) & (!x406x)) + ((x21x) & (n_n491) & (n_n130) & (n_n5154) & (x406x)));
	assign n_n1443 = (((!n_n5157) & (!n_n5149) & (!n_n5152) & (!x195x) & (x12261x)) + ((!n_n5157) & (!n_n5149) & (!n_n5152) & (x195x) & (!x12261x)) + ((!n_n5157) & (!n_n5149) & (!n_n5152) & (x195x) & (x12261x)) + ((!n_n5157) & (!n_n5149) & (n_n5152) & (!x195x) & (!x12261x)) + ((!n_n5157) & (!n_n5149) & (n_n5152) & (!x195x) & (x12261x)) + ((!n_n5157) & (!n_n5149) & (n_n5152) & (x195x) & (!x12261x)) + ((!n_n5157) & (!n_n5149) & (n_n5152) & (x195x) & (x12261x)) + ((!n_n5157) & (n_n5149) & (!n_n5152) & (!x195x) & (!x12261x)) + ((!n_n5157) & (n_n5149) & (!n_n5152) & (!x195x) & (x12261x)) + ((!n_n5157) & (n_n5149) & (!n_n5152) & (x195x) & (!x12261x)) + ((!n_n5157) & (n_n5149) & (!n_n5152) & (x195x) & (x12261x)) + ((!n_n5157) & (n_n5149) & (n_n5152) & (!x195x) & (!x12261x)) + ((!n_n5157) & (n_n5149) & (n_n5152) & (!x195x) & (x12261x)) + ((!n_n5157) & (n_n5149) & (n_n5152) & (x195x) & (!x12261x)) + ((!n_n5157) & (n_n5149) & (n_n5152) & (x195x) & (x12261x)) + ((n_n5157) & (!n_n5149) & (!n_n5152) & (!x195x) & (!x12261x)) + ((n_n5157) & (!n_n5149) & (!n_n5152) & (!x195x) & (x12261x)) + ((n_n5157) & (!n_n5149) & (!n_n5152) & (x195x) & (!x12261x)) + ((n_n5157) & (!n_n5149) & (!n_n5152) & (x195x) & (x12261x)) + ((n_n5157) & (!n_n5149) & (n_n5152) & (!x195x) & (!x12261x)) + ((n_n5157) & (!n_n5149) & (n_n5152) & (!x195x) & (x12261x)) + ((n_n5157) & (!n_n5149) & (n_n5152) & (x195x) & (!x12261x)) + ((n_n5157) & (!n_n5149) & (n_n5152) & (x195x) & (x12261x)) + ((n_n5157) & (n_n5149) & (!n_n5152) & (!x195x) & (!x12261x)) + ((n_n5157) & (n_n5149) & (!n_n5152) & (!x195x) & (x12261x)) + ((n_n5157) & (n_n5149) & (!n_n5152) & (x195x) & (!x12261x)) + ((n_n5157) & (n_n5149) & (!n_n5152) & (x195x) & (x12261x)) + ((n_n5157) & (n_n5149) & (n_n5152) & (!x195x) & (!x12261x)) + ((n_n5157) & (n_n5149) & (n_n5152) & (!x195x) & (x12261x)) + ((n_n5157) & (n_n5149) & (n_n5152) & (x195x) & (!x12261x)) + ((n_n5157) & (n_n5149) & (n_n5152) & (x195x) & (x12261x)));
	assign n_n5288 = (((!i_5_) & (!i_3_) & (i_4_) & (x19x) & (n_n534)));
	assign n_n5292 = (((!i_5_) & (!i_3_) & (i_4_) & (x19x) & (n_n530)));
	assign x208x = (((!i_9_) & (!n_n482) & (!n_n532) & (!n_n65) & (n_n5292)) + ((!i_9_) & (!n_n482) & (!n_n532) & (n_n65) & (n_n5292)) + ((!i_9_) & (!n_n482) & (n_n532) & (!n_n65) & (n_n5292)) + ((!i_9_) & (!n_n482) & (n_n532) & (n_n65) & (n_n5292)) + ((!i_9_) & (n_n482) & (!n_n532) & (!n_n65) & (n_n5292)) + ((!i_9_) & (n_n482) & (!n_n532) & (n_n65) & (n_n5292)) + ((!i_9_) & (n_n482) & (n_n532) & (!n_n65) & (n_n5292)) + ((!i_9_) & (n_n482) & (n_n532) & (n_n65) & (!n_n5292)) + ((!i_9_) & (n_n482) & (n_n532) & (n_n65) & (n_n5292)) + ((i_9_) & (!n_n482) & (!n_n532) & (!n_n65) & (n_n5292)) + ((i_9_) & (!n_n482) & (!n_n532) & (n_n65) & (n_n5292)) + ((i_9_) & (!n_n482) & (n_n532) & (!n_n65) & (n_n5292)) + ((i_9_) & (!n_n482) & (n_n532) & (n_n65) & (n_n5292)) + ((i_9_) & (n_n482) & (!n_n532) & (!n_n65) & (n_n5292)) + ((i_9_) & (n_n482) & (!n_n532) & (n_n65) & (n_n5292)) + ((i_9_) & (n_n482) & (n_n532) & (!n_n65) & (n_n5292)) + ((i_9_) & (n_n482) & (n_n532) & (n_n65) & (n_n5292)));
	assign n_n5298 = (((i_7_) & (!i_8_) & (!i_6_) & (x19x) & (n_n482)));
	assign x22205x = (((!x592x) & (!n_n5293) & (!n_n5297) & (!x11x) & (!n_n5298)) + ((!x592x) & (!n_n5293) & (!n_n5297) & (x11x) & (!n_n5298)) + ((x592x) & (!n_n5293) & (!n_n5297) & (!x11x) & (!n_n5298)));
	assign n_n1432 = (((!n_n5290) & (!n_n5289) & (!n_n5288) & (!x208x) & (!x22205x)) + ((!n_n5290) & (!n_n5289) & (!n_n5288) & (x208x) & (!x22205x)) + ((!n_n5290) & (!n_n5289) & (!n_n5288) & (x208x) & (x22205x)) + ((!n_n5290) & (!n_n5289) & (n_n5288) & (!x208x) & (!x22205x)) + ((!n_n5290) & (!n_n5289) & (n_n5288) & (!x208x) & (x22205x)) + ((!n_n5290) & (!n_n5289) & (n_n5288) & (x208x) & (!x22205x)) + ((!n_n5290) & (!n_n5289) & (n_n5288) & (x208x) & (x22205x)) + ((!n_n5290) & (n_n5289) & (!n_n5288) & (!x208x) & (!x22205x)) + ((!n_n5290) & (n_n5289) & (!n_n5288) & (!x208x) & (x22205x)) + ((!n_n5290) & (n_n5289) & (!n_n5288) & (x208x) & (!x22205x)) + ((!n_n5290) & (n_n5289) & (!n_n5288) & (x208x) & (x22205x)) + ((!n_n5290) & (n_n5289) & (n_n5288) & (!x208x) & (!x22205x)) + ((!n_n5290) & (n_n5289) & (n_n5288) & (!x208x) & (x22205x)) + ((!n_n5290) & (n_n5289) & (n_n5288) & (x208x) & (!x22205x)) + ((!n_n5290) & (n_n5289) & (n_n5288) & (x208x) & (x22205x)) + ((n_n5290) & (!n_n5289) & (!n_n5288) & (!x208x) & (!x22205x)) + ((n_n5290) & (!n_n5289) & (!n_n5288) & (!x208x) & (x22205x)) + ((n_n5290) & (!n_n5289) & (!n_n5288) & (x208x) & (!x22205x)) + ((n_n5290) & (!n_n5289) & (!n_n5288) & (x208x) & (x22205x)) + ((n_n5290) & (!n_n5289) & (n_n5288) & (!x208x) & (!x22205x)) + ((n_n5290) & (!n_n5289) & (n_n5288) & (!x208x) & (x22205x)) + ((n_n5290) & (!n_n5289) & (n_n5288) & (x208x) & (!x22205x)) + ((n_n5290) & (!n_n5289) & (n_n5288) & (x208x) & (x22205x)) + ((n_n5290) & (n_n5289) & (!n_n5288) & (!x208x) & (!x22205x)) + ((n_n5290) & (n_n5289) & (!n_n5288) & (!x208x) & (x22205x)) + ((n_n5290) & (n_n5289) & (!n_n5288) & (x208x) & (!x22205x)) + ((n_n5290) & (n_n5289) & (!n_n5288) & (x208x) & (x22205x)) + ((n_n5290) & (n_n5289) & (n_n5288) & (!x208x) & (!x22205x)) + ((n_n5290) & (n_n5289) & (n_n5288) & (!x208x) & (x22205x)) + ((n_n5290) & (n_n5289) & (n_n5288) & (x208x) & (!x22205x)) + ((n_n5290) & (n_n5289) & (n_n5288) & (x208x) & (x22205x)));
	assign x12117x = (((!x492x) & (!x18x) & (!n_n5022) & (!n_n5043) & (n_n5045)) + ((!x492x) & (!x18x) & (!n_n5022) & (n_n5043) & (!n_n5045)) + ((!x492x) & (!x18x) & (!n_n5022) & (n_n5043) & (n_n5045)) + ((!x492x) & (!x18x) & (n_n5022) & (!n_n5043) & (!n_n5045)) + ((!x492x) & (!x18x) & (n_n5022) & (!n_n5043) & (n_n5045)) + ((!x492x) & (!x18x) & (n_n5022) & (n_n5043) & (!n_n5045)) + ((!x492x) & (!x18x) & (n_n5022) & (n_n5043) & (n_n5045)) + ((!x492x) & (x18x) & (!n_n5022) & (!n_n5043) & (n_n5045)) + ((!x492x) & (x18x) & (!n_n5022) & (n_n5043) & (!n_n5045)) + ((!x492x) & (x18x) & (!n_n5022) & (n_n5043) & (n_n5045)) + ((!x492x) & (x18x) & (n_n5022) & (!n_n5043) & (!n_n5045)) + ((!x492x) & (x18x) & (n_n5022) & (!n_n5043) & (n_n5045)) + ((!x492x) & (x18x) & (n_n5022) & (n_n5043) & (!n_n5045)) + ((!x492x) & (x18x) & (n_n5022) & (n_n5043) & (n_n5045)) + ((x492x) & (!x18x) & (!n_n5022) & (!n_n5043) & (n_n5045)) + ((x492x) & (!x18x) & (!n_n5022) & (n_n5043) & (!n_n5045)) + ((x492x) & (!x18x) & (!n_n5022) & (n_n5043) & (n_n5045)) + ((x492x) & (!x18x) & (n_n5022) & (!n_n5043) & (!n_n5045)) + ((x492x) & (!x18x) & (n_n5022) & (!n_n5043) & (n_n5045)) + ((x492x) & (!x18x) & (n_n5022) & (n_n5043) & (!n_n5045)) + ((x492x) & (!x18x) & (n_n5022) & (n_n5043) & (n_n5045)) + ((x492x) & (x18x) & (!n_n5022) & (!n_n5043) & (!n_n5045)) + ((x492x) & (x18x) & (!n_n5022) & (!n_n5043) & (n_n5045)) + ((x492x) & (x18x) & (!n_n5022) & (n_n5043) & (!n_n5045)) + ((x492x) & (x18x) & (!n_n5022) & (n_n5043) & (n_n5045)) + ((x492x) & (x18x) & (n_n5022) & (!n_n5043) & (!n_n5045)) + ((x492x) & (x18x) & (n_n5022) & (!n_n5043) & (n_n5045)) + ((x492x) & (x18x) & (n_n5022) & (n_n5043) & (!n_n5045)) + ((x492x) & (x18x) & (n_n5022) & (n_n5043) & (n_n5045)));
	assign x12118x = (((!n_n5025) & (!n_n5057) & (!n_n5048) & (!n_n5053) & (n_n5009)) + ((!n_n5025) & (!n_n5057) & (!n_n5048) & (n_n5053) & (!n_n5009)) + ((!n_n5025) & (!n_n5057) & (!n_n5048) & (n_n5053) & (n_n5009)) + ((!n_n5025) & (!n_n5057) & (n_n5048) & (!n_n5053) & (!n_n5009)) + ((!n_n5025) & (!n_n5057) & (n_n5048) & (!n_n5053) & (n_n5009)) + ((!n_n5025) & (!n_n5057) & (n_n5048) & (n_n5053) & (!n_n5009)) + ((!n_n5025) & (!n_n5057) & (n_n5048) & (n_n5053) & (n_n5009)) + ((!n_n5025) & (n_n5057) & (!n_n5048) & (!n_n5053) & (!n_n5009)) + ((!n_n5025) & (n_n5057) & (!n_n5048) & (!n_n5053) & (n_n5009)) + ((!n_n5025) & (n_n5057) & (!n_n5048) & (n_n5053) & (!n_n5009)) + ((!n_n5025) & (n_n5057) & (!n_n5048) & (n_n5053) & (n_n5009)) + ((!n_n5025) & (n_n5057) & (n_n5048) & (!n_n5053) & (!n_n5009)) + ((!n_n5025) & (n_n5057) & (n_n5048) & (!n_n5053) & (n_n5009)) + ((!n_n5025) & (n_n5057) & (n_n5048) & (n_n5053) & (!n_n5009)) + ((!n_n5025) & (n_n5057) & (n_n5048) & (n_n5053) & (n_n5009)) + ((n_n5025) & (!n_n5057) & (!n_n5048) & (!n_n5053) & (!n_n5009)) + ((n_n5025) & (!n_n5057) & (!n_n5048) & (!n_n5053) & (n_n5009)) + ((n_n5025) & (!n_n5057) & (!n_n5048) & (n_n5053) & (!n_n5009)) + ((n_n5025) & (!n_n5057) & (!n_n5048) & (n_n5053) & (n_n5009)) + ((n_n5025) & (!n_n5057) & (n_n5048) & (!n_n5053) & (!n_n5009)) + ((n_n5025) & (!n_n5057) & (n_n5048) & (!n_n5053) & (n_n5009)) + ((n_n5025) & (!n_n5057) & (n_n5048) & (n_n5053) & (!n_n5009)) + ((n_n5025) & (!n_n5057) & (n_n5048) & (n_n5053) & (n_n5009)) + ((n_n5025) & (n_n5057) & (!n_n5048) & (!n_n5053) & (!n_n5009)) + ((n_n5025) & (n_n5057) & (!n_n5048) & (!n_n5053) & (n_n5009)) + ((n_n5025) & (n_n5057) & (!n_n5048) & (n_n5053) & (!n_n5009)) + ((n_n5025) & (n_n5057) & (!n_n5048) & (n_n5053) & (n_n5009)) + ((n_n5025) & (n_n5057) & (n_n5048) & (!n_n5053) & (!n_n5009)) + ((n_n5025) & (n_n5057) & (n_n5048) & (!n_n5053) & (n_n5009)) + ((n_n5025) & (n_n5057) & (n_n5048) & (n_n5053) & (!n_n5009)) + ((n_n5025) & (n_n5057) & (n_n5048) & (n_n5053) & (n_n5009)));
	assign n_n4954 = (((i_9_) & (n_n532) & (n_n535) & (n_n195)));
	assign x12124x = (((!n_n4971) & (!x68x) & (!n_n4972) & (n_n4954)) + ((!n_n4971) & (!x68x) & (n_n4972) & (!n_n4954)) + ((!n_n4971) & (!x68x) & (n_n4972) & (n_n4954)) + ((!n_n4971) & (x68x) & (!n_n4972) & (!n_n4954)) + ((!n_n4971) & (x68x) & (!n_n4972) & (n_n4954)) + ((!n_n4971) & (x68x) & (n_n4972) & (!n_n4954)) + ((!n_n4971) & (x68x) & (n_n4972) & (n_n4954)) + ((n_n4971) & (!x68x) & (!n_n4972) & (!n_n4954)) + ((n_n4971) & (!x68x) & (!n_n4972) & (n_n4954)) + ((n_n4971) & (!x68x) & (n_n4972) & (!n_n4954)) + ((n_n4971) & (!x68x) & (n_n4972) & (n_n4954)) + ((n_n4971) & (x68x) & (!n_n4972) & (!n_n4954)) + ((n_n4971) & (x68x) & (!n_n4972) & (n_n4954)) + ((n_n4971) & (x68x) & (n_n4972) & (!n_n4954)) + ((n_n4971) & (x68x) & (n_n4972) & (n_n4954)));
	assign n_n1333 = (((!n_n4987) & (!n_n4980) & (!n_n5005) & (!n_n4974) & (x12124x)) + ((!n_n4987) & (!n_n4980) & (!n_n5005) & (n_n4974) & (!x12124x)) + ((!n_n4987) & (!n_n4980) & (!n_n5005) & (n_n4974) & (x12124x)) + ((!n_n4987) & (!n_n4980) & (n_n5005) & (!n_n4974) & (!x12124x)) + ((!n_n4987) & (!n_n4980) & (n_n5005) & (!n_n4974) & (x12124x)) + ((!n_n4987) & (!n_n4980) & (n_n5005) & (n_n4974) & (!x12124x)) + ((!n_n4987) & (!n_n4980) & (n_n5005) & (n_n4974) & (x12124x)) + ((!n_n4987) & (n_n4980) & (!n_n5005) & (!n_n4974) & (!x12124x)) + ((!n_n4987) & (n_n4980) & (!n_n5005) & (!n_n4974) & (x12124x)) + ((!n_n4987) & (n_n4980) & (!n_n5005) & (n_n4974) & (!x12124x)) + ((!n_n4987) & (n_n4980) & (!n_n5005) & (n_n4974) & (x12124x)) + ((!n_n4987) & (n_n4980) & (n_n5005) & (!n_n4974) & (!x12124x)) + ((!n_n4987) & (n_n4980) & (n_n5005) & (!n_n4974) & (x12124x)) + ((!n_n4987) & (n_n4980) & (n_n5005) & (n_n4974) & (!x12124x)) + ((!n_n4987) & (n_n4980) & (n_n5005) & (n_n4974) & (x12124x)) + ((n_n4987) & (!n_n4980) & (!n_n5005) & (!n_n4974) & (!x12124x)) + ((n_n4987) & (!n_n4980) & (!n_n5005) & (!n_n4974) & (x12124x)) + ((n_n4987) & (!n_n4980) & (!n_n5005) & (n_n4974) & (!x12124x)) + ((n_n4987) & (!n_n4980) & (!n_n5005) & (n_n4974) & (x12124x)) + ((n_n4987) & (!n_n4980) & (n_n5005) & (!n_n4974) & (!x12124x)) + ((n_n4987) & (!n_n4980) & (n_n5005) & (!n_n4974) & (x12124x)) + ((n_n4987) & (!n_n4980) & (n_n5005) & (n_n4974) & (!x12124x)) + ((n_n4987) & (!n_n4980) & (n_n5005) & (n_n4974) & (x12124x)) + ((n_n4987) & (n_n4980) & (!n_n5005) & (!n_n4974) & (!x12124x)) + ((n_n4987) & (n_n4980) & (!n_n5005) & (!n_n4974) & (x12124x)) + ((n_n4987) & (n_n4980) & (!n_n5005) & (n_n4974) & (!x12124x)) + ((n_n4987) & (n_n4980) & (!n_n5005) & (n_n4974) & (x12124x)) + ((n_n4987) & (n_n4980) & (n_n5005) & (!n_n4974) & (!x12124x)) + ((n_n4987) & (n_n4980) & (n_n5005) & (!n_n4974) & (x12124x)) + ((n_n4987) & (n_n4980) & (n_n5005) & (n_n4974) & (!x12124x)) + ((n_n4987) & (n_n4980) & (n_n5005) & (n_n4974) & (x12124x)));
	assign n_n4626 = (((i_9_) & (n_n524) & (n_n390) & (n_n500)));
	assign n_n4627 = (((!i_9_) & (n_n524) & (n_n390) & (n_n500)));
	assign n_n4660 = (((i_9_) & (n_n482) & (n_n390) & (n_n522)));
	assign n_n4955 = (((!i_9_) & (n_n532) & (n_n535) & (n_n195)));
	assign n_n5138 = (((i_7_) & (!i_8_) & (!i_6_) & (x12x) & (n_n500)));
	assign n_n5309 = (((!i_9_) & (n_n473) & (n_n530) & (n_n65)));
	assign n_n1128 = (((!i_9_) & (!n_n473) & (!n_n530) & (n_n5310) & (!n_n65)) + ((!i_9_) & (!n_n473) & (!n_n530) & (n_n5310) & (n_n65)) + ((!i_9_) & (!n_n473) & (n_n530) & (n_n5310) & (!n_n65)) + ((!i_9_) & (!n_n473) & (n_n530) & (n_n5310) & (n_n65)) + ((!i_9_) & (n_n473) & (!n_n530) & (n_n5310) & (!n_n65)) + ((!i_9_) & (n_n473) & (!n_n530) & (n_n5310) & (n_n65)) + ((!i_9_) & (n_n473) & (n_n530) & (!n_n5310) & (n_n65)) + ((!i_9_) & (n_n473) & (n_n530) & (n_n5310) & (!n_n65)) + ((!i_9_) & (n_n473) & (n_n530) & (n_n5310) & (n_n65)) + ((i_9_) & (!n_n473) & (!n_n530) & (n_n5310) & (!n_n65)) + ((i_9_) & (!n_n473) & (!n_n530) & (n_n5310) & (n_n65)) + ((i_9_) & (!n_n473) & (n_n530) & (n_n5310) & (!n_n65)) + ((i_9_) & (!n_n473) & (n_n530) & (n_n5310) & (n_n65)) + ((i_9_) & (n_n473) & (!n_n530) & (n_n5310) & (!n_n65)) + ((i_9_) & (n_n473) & (!n_n530) & (n_n5310) & (n_n65)) + ((i_9_) & (n_n473) & (n_n530) & (!n_n5310) & (n_n65)) + ((i_9_) & (n_n473) & (n_n530) & (n_n5310) & (!n_n65)) + ((i_9_) & (n_n473) & (n_n530) & (n_n5310) & (n_n65)));
	assign x420x = (((!i_9_) & (n_n536) & (!n_n526) & (n_n528) & (n_n491)) + ((!i_9_) & (n_n536) & (n_n526) & (!n_n528) & (n_n491)) + ((!i_9_) & (n_n536) & (n_n526) & (n_n528) & (n_n491)));
	assign x11592x = (((!n_n4380) & (!n_n4379) & (!n_n4388) & (!n_n4386) & (n_n4387)) + ((!n_n4380) & (!n_n4379) & (!n_n4388) & (n_n4386) & (!n_n4387)) + ((!n_n4380) & (!n_n4379) & (!n_n4388) & (n_n4386) & (n_n4387)) + ((!n_n4380) & (!n_n4379) & (n_n4388) & (!n_n4386) & (!n_n4387)) + ((!n_n4380) & (!n_n4379) & (n_n4388) & (!n_n4386) & (n_n4387)) + ((!n_n4380) & (!n_n4379) & (n_n4388) & (n_n4386) & (!n_n4387)) + ((!n_n4380) & (!n_n4379) & (n_n4388) & (n_n4386) & (n_n4387)) + ((!n_n4380) & (n_n4379) & (!n_n4388) & (!n_n4386) & (!n_n4387)) + ((!n_n4380) & (n_n4379) & (!n_n4388) & (!n_n4386) & (n_n4387)) + ((!n_n4380) & (n_n4379) & (!n_n4388) & (n_n4386) & (!n_n4387)) + ((!n_n4380) & (n_n4379) & (!n_n4388) & (n_n4386) & (n_n4387)) + ((!n_n4380) & (n_n4379) & (n_n4388) & (!n_n4386) & (!n_n4387)) + ((!n_n4380) & (n_n4379) & (n_n4388) & (!n_n4386) & (n_n4387)) + ((!n_n4380) & (n_n4379) & (n_n4388) & (n_n4386) & (!n_n4387)) + ((!n_n4380) & (n_n4379) & (n_n4388) & (n_n4386) & (n_n4387)) + ((n_n4380) & (!n_n4379) & (!n_n4388) & (!n_n4386) & (!n_n4387)) + ((n_n4380) & (!n_n4379) & (!n_n4388) & (!n_n4386) & (n_n4387)) + ((n_n4380) & (!n_n4379) & (!n_n4388) & (n_n4386) & (!n_n4387)) + ((n_n4380) & (!n_n4379) & (!n_n4388) & (n_n4386) & (n_n4387)) + ((n_n4380) & (!n_n4379) & (n_n4388) & (!n_n4386) & (!n_n4387)) + ((n_n4380) & (!n_n4379) & (n_n4388) & (!n_n4386) & (n_n4387)) + ((n_n4380) & (!n_n4379) & (n_n4388) & (n_n4386) & (!n_n4387)) + ((n_n4380) & (!n_n4379) & (n_n4388) & (n_n4386) & (n_n4387)) + ((n_n4380) & (n_n4379) & (!n_n4388) & (!n_n4386) & (!n_n4387)) + ((n_n4380) & (n_n4379) & (!n_n4388) & (!n_n4386) & (n_n4387)) + ((n_n4380) & (n_n4379) & (!n_n4388) & (n_n4386) & (!n_n4387)) + ((n_n4380) & (n_n4379) & (!n_n4388) & (n_n4386) & (n_n4387)) + ((n_n4380) & (n_n4379) & (n_n4388) & (!n_n4386) & (!n_n4387)) + ((n_n4380) & (n_n4379) & (n_n4388) & (!n_n4386) & (n_n4387)) + ((n_n4380) & (n_n4379) & (n_n4388) & (n_n4386) & (!n_n4387)) + ((n_n4380) & (n_n4379) & (n_n4388) & (n_n4386) & (n_n4387)));
	assign n_n1117 = (((!n_n4383) & (!n_n4389) & (!n_n4381) & (!n_n4385) & (x11592x)) + ((!n_n4383) & (!n_n4389) & (!n_n4381) & (n_n4385) & (!x11592x)) + ((!n_n4383) & (!n_n4389) & (!n_n4381) & (n_n4385) & (x11592x)) + ((!n_n4383) & (!n_n4389) & (n_n4381) & (!n_n4385) & (!x11592x)) + ((!n_n4383) & (!n_n4389) & (n_n4381) & (!n_n4385) & (x11592x)) + ((!n_n4383) & (!n_n4389) & (n_n4381) & (n_n4385) & (!x11592x)) + ((!n_n4383) & (!n_n4389) & (n_n4381) & (n_n4385) & (x11592x)) + ((!n_n4383) & (n_n4389) & (!n_n4381) & (!n_n4385) & (!x11592x)) + ((!n_n4383) & (n_n4389) & (!n_n4381) & (!n_n4385) & (x11592x)) + ((!n_n4383) & (n_n4389) & (!n_n4381) & (n_n4385) & (!x11592x)) + ((!n_n4383) & (n_n4389) & (!n_n4381) & (n_n4385) & (x11592x)) + ((!n_n4383) & (n_n4389) & (n_n4381) & (!n_n4385) & (!x11592x)) + ((!n_n4383) & (n_n4389) & (n_n4381) & (!n_n4385) & (x11592x)) + ((!n_n4383) & (n_n4389) & (n_n4381) & (n_n4385) & (!x11592x)) + ((!n_n4383) & (n_n4389) & (n_n4381) & (n_n4385) & (x11592x)) + ((n_n4383) & (!n_n4389) & (!n_n4381) & (!n_n4385) & (!x11592x)) + ((n_n4383) & (!n_n4389) & (!n_n4381) & (!n_n4385) & (x11592x)) + ((n_n4383) & (!n_n4389) & (!n_n4381) & (n_n4385) & (!x11592x)) + ((n_n4383) & (!n_n4389) & (!n_n4381) & (n_n4385) & (x11592x)) + ((n_n4383) & (!n_n4389) & (n_n4381) & (!n_n4385) & (!x11592x)) + ((n_n4383) & (!n_n4389) & (n_n4381) & (!n_n4385) & (x11592x)) + ((n_n4383) & (!n_n4389) & (n_n4381) & (n_n4385) & (!x11592x)) + ((n_n4383) & (!n_n4389) & (n_n4381) & (n_n4385) & (x11592x)) + ((n_n4383) & (n_n4389) & (!n_n4381) & (!n_n4385) & (!x11592x)) + ((n_n4383) & (n_n4389) & (!n_n4381) & (!n_n4385) & (x11592x)) + ((n_n4383) & (n_n4389) & (!n_n4381) & (n_n4385) & (!x11592x)) + ((n_n4383) & (n_n4389) & (!n_n4381) & (n_n4385) & (x11592x)) + ((n_n4383) & (n_n4389) & (n_n4381) & (!n_n4385) & (!x11592x)) + ((n_n4383) & (n_n4389) & (n_n4381) & (!n_n4385) & (x11592x)) + ((n_n4383) & (n_n4389) & (n_n4381) & (n_n4385) & (!x11592x)) + ((n_n4383) & (n_n4389) & (n_n4381) & (n_n4385) & (x11592x)));
	assign x11505x = (((!i_9_) & (n_n524) & (n_n518) & (n_n455)) + ((i_9_) & (n_n524) & (n_n518) & (n_n455)));
	assign x22169x = (((!n_n4617) & (!n_n4613) & (!n_n4612) & (!n_n4611)));
	assign n_n1099 = (((!n_n4618) & (!n_n4619) & (!n_n4232) & (!x22169x)) + ((!n_n4618) & (!n_n4619) & (n_n4232) & (!x22169x)) + ((!n_n4618) & (!n_n4619) & (n_n4232) & (x22169x)) + ((!n_n4618) & (n_n4619) & (!n_n4232) & (!x22169x)) + ((!n_n4618) & (n_n4619) & (!n_n4232) & (x22169x)) + ((!n_n4618) & (n_n4619) & (n_n4232) & (!x22169x)) + ((!n_n4618) & (n_n4619) & (n_n4232) & (x22169x)) + ((n_n4618) & (!n_n4619) & (!n_n4232) & (!x22169x)) + ((n_n4618) & (!n_n4619) & (!n_n4232) & (x22169x)) + ((n_n4618) & (!n_n4619) & (n_n4232) & (!x22169x)) + ((n_n4618) & (!n_n4619) & (n_n4232) & (x22169x)) + ((n_n4618) & (n_n4619) & (!n_n4232) & (!x22169x)) + ((n_n4618) & (n_n4619) & (!n_n4232) & (x22169x)) + ((n_n4618) & (n_n4619) & (n_n4232) & (!x22169x)) + ((n_n4618) & (n_n4619) & (n_n4232) & (x22169x)));
	assign x111x = (((!i_9_) & (n_n524) & (!n_n522) & (n_n491) & (n_n195)) + ((!i_9_) & (n_n524) & (n_n522) & (n_n491) & (n_n195)) + ((i_9_) & (!n_n524) & (n_n522) & (n_n491) & (n_n195)) + ((i_9_) & (n_n524) & (n_n522) & (n_n491) & (n_n195)));
	assign x458x = (((!n_n491) & (!n_n195) & (!x20x) & (x50x)) + ((!n_n491) & (!n_n195) & (x20x) & (x50x)) + ((!n_n491) & (n_n195) & (!x20x) & (x50x)) + ((!n_n491) & (n_n195) & (x20x) & (x50x)) + ((n_n491) & (!n_n195) & (!x20x) & (x50x)) + ((n_n491) & (!n_n195) & (x20x) & (x50x)) + ((n_n491) & (n_n195) & (!x20x) & (x50x)) + ((n_n491) & (n_n195) & (x20x) & (!x50x)) + ((n_n491) & (n_n195) & (x20x) & (x50x)));
	assign n_n1066 = (((!n_n5026) & (!n_n5022) & (!x296x) & (!x111x) & (x458x)) + ((!n_n5026) & (!n_n5022) & (!x296x) & (x111x) & (!x458x)) + ((!n_n5026) & (!n_n5022) & (!x296x) & (x111x) & (x458x)) + ((!n_n5026) & (!n_n5022) & (x296x) & (!x111x) & (!x458x)) + ((!n_n5026) & (!n_n5022) & (x296x) & (!x111x) & (x458x)) + ((!n_n5026) & (!n_n5022) & (x296x) & (x111x) & (!x458x)) + ((!n_n5026) & (!n_n5022) & (x296x) & (x111x) & (x458x)) + ((!n_n5026) & (n_n5022) & (!x296x) & (!x111x) & (!x458x)) + ((!n_n5026) & (n_n5022) & (!x296x) & (!x111x) & (x458x)) + ((!n_n5026) & (n_n5022) & (!x296x) & (x111x) & (!x458x)) + ((!n_n5026) & (n_n5022) & (!x296x) & (x111x) & (x458x)) + ((!n_n5026) & (n_n5022) & (x296x) & (!x111x) & (!x458x)) + ((!n_n5026) & (n_n5022) & (x296x) & (!x111x) & (x458x)) + ((!n_n5026) & (n_n5022) & (x296x) & (x111x) & (!x458x)) + ((!n_n5026) & (n_n5022) & (x296x) & (x111x) & (x458x)) + ((n_n5026) & (!n_n5022) & (!x296x) & (!x111x) & (!x458x)) + ((n_n5026) & (!n_n5022) & (!x296x) & (!x111x) & (x458x)) + ((n_n5026) & (!n_n5022) & (!x296x) & (x111x) & (!x458x)) + ((n_n5026) & (!n_n5022) & (!x296x) & (x111x) & (x458x)) + ((n_n5026) & (!n_n5022) & (x296x) & (!x111x) & (!x458x)) + ((n_n5026) & (!n_n5022) & (x296x) & (!x111x) & (x458x)) + ((n_n5026) & (!n_n5022) & (x296x) & (x111x) & (!x458x)) + ((n_n5026) & (!n_n5022) & (x296x) & (x111x) & (x458x)) + ((n_n5026) & (n_n5022) & (!x296x) & (!x111x) & (!x458x)) + ((n_n5026) & (n_n5022) & (!x296x) & (!x111x) & (x458x)) + ((n_n5026) & (n_n5022) & (!x296x) & (x111x) & (!x458x)) + ((n_n5026) & (n_n5022) & (!x296x) & (x111x) & (x458x)) + ((n_n5026) & (n_n5022) & (x296x) & (!x111x) & (!x458x)) + ((n_n5026) & (n_n5022) & (x296x) & (!x111x) & (x458x)) + ((n_n5026) & (n_n5022) & (x296x) & (x111x) & (!x458x)) + ((n_n5026) & (n_n5022) & (x296x) & (x111x) & (x458x)));
	assign n_n4745 = (((!i_9_) & (n_n534) & (n_n325) & (n_n500)));
	assign x11842x = (((!n_n4751) & (!n_n4750) & (!n_n4748) & (!n_n4747) & (n_n4745)) + ((!n_n4751) & (!n_n4750) & (!n_n4748) & (n_n4747) & (!n_n4745)) + ((!n_n4751) & (!n_n4750) & (!n_n4748) & (n_n4747) & (n_n4745)) + ((!n_n4751) & (!n_n4750) & (n_n4748) & (!n_n4747) & (!n_n4745)) + ((!n_n4751) & (!n_n4750) & (n_n4748) & (!n_n4747) & (n_n4745)) + ((!n_n4751) & (!n_n4750) & (n_n4748) & (n_n4747) & (!n_n4745)) + ((!n_n4751) & (!n_n4750) & (n_n4748) & (n_n4747) & (n_n4745)) + ((!n_n4751) & (n_n4750) & (!n_n4748) & (!n_n4747) & (!n_n4745)) + ((!n_n4751) & (n_n4750) & (!n_n4748) & (!n_n4747) & (n_n4745)) + ((!n_n4751) & (n_n4750) & (!n_n4748) & (n_n4747) & (!n_n4745)) + ((!n_n4751) & (n_n4750) & (!n_n4748) & (n_n4747) & (n_n4745)) + ((!n_n4751) & (n_n4750) & (n_n4748) & (!n_n4747) & (!n_n4745)) + ((!n_n4751) & (n_n4750) & (n_n4748) & (!n_n4747) & (n_n4745)) + ((!n_n4751) & (n_n4750) & (n_n4748) & (n_n4747) & (!n_n4745)) + ((!n_n4751) & (n_n4750) & (n_n4748) & (n_n4747) & (n_n4745)) + ((n_n4751) & (!n_n4750) & (!n_n4748) & (!n_n4747) & (!n_n4745)) + ((n_n4751) & (!n_n4750) & (!n_n4748) & (!n_n4747) & (n_n4745)) + ((n_n4751) & (!n_n4750) & (!n_n4748) & (n_n4747) & (!n_n4745)) + ((n_n4751) & (!n_n4750) & (!n_n4748) & (n_n4747) & (n_n4745)) + ((n_n4751) & (!n_n4750) & (n_n4748) & (!n_n4747) & (!n_n4745)) + ((n_n4751) & (!n_n4750) & (n_n4748) & (!n_n4747) & (n_n4745)) + ((n_n4751) & (!n_n4750) & (n_n4748) & (n_n4747) & (!n_n4745)) + ((n_n4751) & (!n_n4750) & (n_n4748) & (n_n4747) & (n_n4745)) + ((n_n4751) & (n_n4750) & (!n_n4748) & (!n_n4747) & (!n_n4745)) + ((n_n4751) & (n_n4750) & (!n_n4748) & (!n_n4747) & (n_n4745)) + ((n_n4751) & (n_n4750) & (!n_n4748) & (n_n4747) & (!n_n4745)) + ((n_n4751) & (n_n4750) & (!n_n4748) & (n_n4747) & (n_n4745)) + ((n_n4751) & (n_n4750) & (n_n4748) & (!n_n4747) & (!n_n4745)) + ((n_n4751) & (n_n4750) & (n_n4748) & (!n_n4747) & (n_n4745)) + ((n_n4751) & (n_n4750) & (n_n4748) & (n_n4747) & (!n_n4745)) + ((n_n4751) & (n_n4750) & (n_n4748) & (n_n4747) & (n_n4745)));
	assign n_n1088 = (((!n_n4754) & (!n_n4753) & (!x47x) & (x11842x)) + ((!n_n4754) & (!n_n4753) & (x47x) & (!x11842x)) + ((!n_n4754) & (!n_n4753) & (x47x) & (x11842x)) + ((!n_n4754) & (n_n4753) & (!x47x) & (!x11842x)) + ((!n_n4754) & (n_n4753) & (!x47x) & (x11842x)) + ((!n_n4754) & (n_n4753) & (x47x) & (!x11842x)) + ((!n_n4754) & (n_n4753) & (x47x) & (x11842x)) + ((n_n4754) & (!n_n4753) & (!x47x) & (!x11842x)) + ((n_n4754) & (!n_n4753) & (!x47x) & (x11842x)) + ((n_n4754) & (!n_n4753) & (x47x) & (!x11842x)) + ((n_n4754) & (!n_n4753) & (x47x) & (x11842x)) + ((n_n4754) & (n_n4753) & (!x47x) & (!x11842x)) + ((n_n4754) & (n_n4753) & (!x47x) & (x11842x)) + ((n_n4754) & (n_n4753) & (x47x) & (!x11842x)) + ((n_n4754) & (n_n4753) & (x47x) & (x11842x)));
	assign n_n4736 = (((i_9_) & (n_n526) & (n_n509) & (n_n325)));
	assign x39x = (((!i_9_) & (!n_n524) & (n_n518) & (n_n526) & (n_n325)) + ((!i_9_) & (n_n524) & (n_n518) & (n_n526) & (n_n325)) + ((i_9_) & (n_n524) & (n_n518) & (!n_n526) & (n_n325)) + ((i_9_) & (n_n524) & (n_n518) & (n_n526) & (n_n325)));
	assign x457x = (((!i_9_) & (!n_n524) & (n_n518) & (n_n526) & (n_n325)) + ((!i_9_) & (n_n524) & (n_n518) & (n_n526) & (n_n325)) + ((i_9_) & (!n_n524) & (n_n518) & (n_n526) & (n_n325)) + ((i_9_) & (n_n524) & (n_n518) & (!n_n526) & (n_n325)) + ((i_9_) & (n_n524) & (n_n518) & (n_n526) & (n_n325)));
	assign x22159x = (((!x483x) & (!x23x) & (!n_n4728) & (!n_n4730) & (!n_n4733)) + ((!x483x) & (x23x) & (!n_n4728) & (!n_n4730) & (!n_n4733)) + ((x483x) & (!x23x) & (!n_n4728) & (!n_n4730) & (!n_n4733)));
	assign x11851x = (((!n_n4720) & (!x95x) & (!n_n4736) & (!x39x) & (!x22159x)) + ((!n_n4720) & (!x95x) & (!n_n4736) & (x39x) & (!x22159x)) + ((!n_n4720) & (!x95x) & (!n_n4736) & (x39x) & (x22159x)) + ((!n_n4720) & (!x95x) & (n_n4736) & (!x39x) & (!x22159x)) + ((!n_n4720) & (!x95x) & (n_n4736) & (!x39x) & (x22159x)) + ((!n_n4720) & (!x95x) & (n_n4736) & (x39x) & (!x22159x)) + ((!n_n4720) & (!x95x) & (n_n4736) & (x39x) & (x22159x)) + ((!n_n4720) & (x95x) & (!n_n4736) & (!x39x) & (!x22159x)) + ((!n_n4720) & (x95x) & (!n_n4736) & (!x39x) & (x22159x)) + ((!n_n4720) & (x95x) & (!n_n4736) & (x39x) & (!x22159x)) + ((!n_n4720) & (x95x) & (!n_n4736) & (x39x) & (x22159x)) + ((!n_n4720) & (x95x) & (n_n4736) & (!x39x) & (!x22159x)) + ((!n_n4720) & (x95x) & (n_n4736) & (!x39x) & (x22159x)) + ((!n_n4720) & (x95x) & (n_n4736) & (x39x) & (!x22159x)) + ((!n_n4720) & (x95x) & (n_n4736) & (x39x) & (x22159x)) + ((n_n4720) & (!x95x) & (!n_n4736) & (!x39x) & (!x22159x)) + ((n_n4720) & (!x95x) & (!n_n4736) & (!x39x) & (x22159x)) + ((n_n4720) & (!x95x) & (!n_n4736) & (x39x) & (!x22159x)) + ((n_n4720) & (!x95x) & (!n_n4736) & (x39x) & (x22159x)) + ((n_n4720) & (!x95x) & (n_n4736) & (!x39x) & (!x22159x)) + ((n_n4720) & (!x95x) & (n_n4736) & (!x39x) & (x22159x)) + ((n_n4720) & (!x95x) & (n_n4736) & (x39x) & (!x22159x)) + ((n_n4720) & (!x95x) & (n_n4736) & (x39x) & (x22159x)) + ((n_n4720) & (x95x) & (!n_n4736) & (!x39x) & (!x22159x)) + ((n_n4720) & (x95x) & (!n_n4736) & (!x39x) & (x22159x)) + ((n_n4720) & (x95x) & (!n_n4736) & (x39x) & (!x22159x)) + ((n_n4720) & (x95x) & (!n_n4736) & (x39x) & (x22159x)) + ((n_n4720) & (x95x) & (n_n4736) & (!x39x) & (!x22159x)) + ((n_n4720) & (x95x) & (n_n4736) & (!x39x) & (x22159x)) + ((n_n4720) & (x95x) & (n_n4736) & (x39x) & (!x22159x)) + ((n_n4720) & (x95x) & (n_n4736) & (x39x) & (x22159x)));
	assign n_n5160 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n534) & (x12x)));
	assign x11900x = (((!n_n5152) & (!n_n5159) & (!x406x) & (n_n5160)) + ((!n_n5152) & (!n_n5159) & (x406x) & (!n_n5160)) + ((!n_n5152) & (!n_n5159) & (x406x) & (n_n5160)) + ((!n_n5152) & (n_n5159) & (!x406x) & (!n_n5160)) + ((!n_n5152) & (n_n5159) & (!x406x) & (n_n5160)) + ((!n_n5152) & (n_n5159) & (x406x) & (!n_n5160)) + ((!n_n5152) & (n_n5159) & (x406x) & (n_n5160)) + ((n_n5152) & (!n_n5159) & (!x406x) & (!n_n5160)) + ((n_n5152) & (!n_n5159) & (!x406x) & (n_n5160)) + ((n_n5152) & (!n_n5159) & (x406x) & (!n_n5160)) + ((n_n5152) & (!n_n5159) & (x406x) & (n_n5160)) + ((n_n5152) & (n_n5159) & (!x406x) & (!n_n5160)) + ((n_n5152) & (n_n5159) & (!x406x) & (n_n5160)) + ((n_n5152) & (n_n5159) & (x406x) & (!n_n5160)) + ((n_n5152) & (n_n5159) & (x406x) & (n_n5160)));
	assign n_n1057 = (((!n_n5156) & (!n_n5162) & (!n_n5157) & (!n_n5154) & (x11900x)) + ((!n_n5156) & (!n_n5162) & (!n_n5157) & (n_n5154) & (!x11900x)) + ((!n_n5156) & (!n_n5162) & (!n_n5157) & (n_n5154) & (x11900x)) + ((!n_n5156) & (!n_n5162) & (n_n5157) & (!n_n5154) & (!x11900x)) + ((!n_n5156) & (!n_n5162) & (n_n5157) & (!n_n5154) & (x11900x)) + ((!n_n5156) & (!n_n5162) & (n_n5157) & (n_n5154) & (!x11900x)) + ((!n_n5156) & (!n_n5162) & (n_n5157) & (n_n5154) & (x11900x)) + ((!n_n5156) & (n_n5162) & (!n_n5157) & (!n_n5154) & (!x11900x)) + ((!n_n5156) & (n_n5162) & (!n_n5157) & (!n_n5154) & (x11900x)) + ((!n_n5156) & (n_n5162) & (!n_n5157) & (n_n5154) & (!x11900x)) + ((!n_n5156) & (n_n5162) & (!n_n5157) & (n_n5154) & (x11900x)) + ((!n_n5156) & (n_n5162) & (n_n5157) & (!n_n5154) & (!x11900x)) + ((!n_n5156) & (n_n5162) & (n_n5157) & (!n_n5154) & (x11900x)) + ((!n_n5156) & (n_n5162) & (n_n5157) & (n_n5154) & (!x11900x)) + ((!n_n5156) & (n_n5162) & (n_n5157) & (n_n5154) & (x11900x)) + ((n_n5156) & (!n_n5162) & (!n_n5157) & (!n_n5154) & (!x11900x)) + ((n_n5156) & (!n_n5162) & (!n_n5157) & (!n_n5154) & (x11900x)) + ((n_n5156) & (!n_n5162) & (!n_n5157) & (n_n5154) & (!x11900x)) + ((n_n5156) & (!n_n5162) & (!n_n5157) & (n_n5154) & (x11900x)) + ((n_n5156) & (!n_n5162) & (n_n5157) & (!n_n5154) & (!x11900x)) + ((n_n5156) & (!n_n5162) & (n_n5157) & (!n_n5154) & (x11900x)) + ((n_n5156) & (!n_n5162) & (n_n5157) & (n_n5154) & (!x11900x)) + ((n_n5156) & (!n_n5162) & (n_n5157) & (n_n5154) & (x11900x)) + ((n_n5156) & (n_n5162) & (!n_n5157) & (!n_n5154) & (!x11900x)) + ((n_n5156) & (n_n5162) & (!n_n5157) & (!n_n5154) & (x11900x)) + ((n_n5156) & (n_n5162) & (!n_n5157) & (n_n5154) & (!x11900x)) + ((n_n5156) & (n_n5162) & (!n_n5157) & (n_n5154) & (x11900x)) + ((n_n5156) & (n_n5162) & (n_n5157) & (!n_n5154) & (!x11900x)) + ((n_n5156) & (n_n5162) & (n_n5157) & (!n_n5154) & (x11900x)) + ((n_n5156) & (n_n5162) & (n_n5157) & (n_n5154) & (!x11900x)) + ((n_n5156) & (n_n5162) & (n_n5157) & (n_n5154) & (x11900x)));
	assign n_n5169 = (((!i_9_) & (n_n526) & (n_n482) & (n_n130)));
	assign x33x = (((!i_9_) & (n_n482) & (!n_n130) & (x12x) & (n_n530)) + ((!i_9_) & (n_n482) & (n_n130) & (!x12x) & (n_n530)) + ((!i_9_) & (n_n482) & (n_n130) & (x12x) & (n_n530)) + ((i_9_) & (n_n482) & (!n_n130) & (x12x) & (n_n530)) + ((i_9_) & (n_n482) & (n_n130) & (x12x) & (n_n530)));
	assign n_n5170 = (((i_7_) & (!i_8_) & (!i_6_) & (n_n482) & (x12x)));
	assign x113x = (((!i_9_) & (n_n526) & (n_n473) & (!n_n130) & (x12x)) + ((!i_9_) & (n_n526) & (n_n473) & (n_n130) & (!x12x)) + ((!i_9_) & (n_n526) & (n_n473) & (n_n130) & (x12x)) + ((i_9_) & (n_n526) & (n_n473) & (!n_n130) & (x12x)) + ((i_9_) & (n_n526) & (n_n473) & (n_n130) & (x12x)));
	assign x254x = (((!i_9_) & (n_n482) & (n_n528) & (!n_n130) & (x12x)) + ((!i_9_) & (n_n482) & (n_n528) & (n_n130) & (!x12x)) + ((!i_9_) & (n_n482) & (n_n528) & (n_n130) & (x12x)) + ((i_9_) & (n_n482) & (n_n528) & (!n_n130) & (x12x)) + ((i_9_) & (n_n482) & (n_n528) & (n_n130) & (x12x)));
	assign n_n5176 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n534) & (x12x)));
	assign x22182x = (((!n_n5174) & (!n_n5181) & (!n_n5173) & (!n_n5175) & (!n_n5176)));
	assign x11908x = (((!n_n3399) & (!n_n5163) & (!n_n5169) & (!x22182x)) + ((!n_n3399) & (!n_n5163) & (n_n5169) & (!x22182x)) + ((!n_n3399) & (!n_n5163) & (n_n5169) & (x22182x)) + ((!n_n3399) & (n_n5163) & (!n_n5169) & (!x22182x)) + ((!n_n3399) & (n_n5163) & (!n_n5169) & (x22182x)) + ((!n_n3399) & (n_n5163) & (n_n5169) & (!x22182x)) + ((!n_n3399) & (n_n5163) & (n_n5169) & (x22182x)) + ((n_n3399) & (!n_n5163) & (!n_n5169) & (!x22182x)) + ((n_n3399) & (!n_n5163) & (!n_n5169) & (x22182x)) + ((n_n3399) & (!n_n5163) & (n_n5169) & (!x22182x)) + ((n_n3399) & (!n_n5163) & (n_n5169) & (x22182x)) + ((n_n3399) & (n_n5163) & (!n_n5169) & (!x22182x)) + ((n_n3399) & (n_n5163) & (!n_n5169) & (x22182x)) + ((n_n3399) & (n_n5163) & (n_n5169) & (!x22182x)) + ((n_n3399) & (n_n5163) & (n_n5169) & (x22182x)));
	assign x11907x = (((!n_n5171) & (!x33x) & (!n_n5170) & (!x113x) & (x254x)) + ((!n_n5171) & (!x33x) & (!n_n5170) & (x113x) & (!x254x)) + ((!n_n5171) & (!x33x) & (!n_n5170) & (x113x) & (x254x)) + ((!n_n5171) & (!x33x) & (n_n5170) & (!x113x) & (!x254x)) + ((!n_n5171) & (!x33x) & (n_n5170) & (!x113x) & (x254x)) + ((!n_n5171) & (!x33x) & (n_n5170) & (x113x) & (!x254x)) + ((!n_n5171) & (!x33x) & (n_n5170) & (x113x) & (x254x)) + ((!n_n5171) & (x33x) & (!n_n5170) & (!x113x) & (!x254x)) + ((!n_n5171) & (x33x) & (!n_n5170) & (!x113x) & (x254x)) + ((!n_n5171) & (x33x) & (!n_n5170) & (x113x) & (!x254x)) + ((!n_n5171) & (x33x) & (!n_n5170) & (x113x) & (x254x)) + ((!n_n5171) & (x33x) & (n_n5170) & (!x113x) & (!x254x)) + ((!n_n5171) & (x33x) & (n_n5170) & (!x113x) & (x254x)) + ((!n_n5171) & (x33x) & (n_n5170) & (x113x) & (!x254x)) + ((!n_n5171) & (x33x) & (n_n5170) & (x113x) & (x254x)) + ((n_n5171) & (!x33x) & (!n_n5170) & (!x113x) & (!x254x)) + ((n_n5171) & (!x33x) & (!n_n5170) & (!x113x) & (x254x)) + ((n_n5171) & (!x33x) & (!n_n5170) & (x113x) & (!x254x)) + ((n_n5171) & (!x33x) & (!n_n5170) & (x113x) & (x254x)) + ((n_n5171) & (!x33x) & (n_n5170) & (!x113x) & (!x254x)) + ((n_n5171) & (!x33x) & (n_n5170) & (!x113x) & (x254x)) + ((n_n5171) & (!x33x) & (n_n5170) & (x113x) & (!x254x)) + ((n_n5171) & (!x33x) & (n_n5170) & (x113x) & (x254x)) + ((n_n5171) & (x33x) & (!n_n5170) & (!x113x) & (!x254x)) + ((n_n5171) & (x33x) & (!n_n5170) & (!x113x) & (x254x)) + ((n_n5171) & (x33x) & (!n_n5170) & (x113x) & (!x254x)) + ((n_n5171) & (x33x) & (!n_n5170) & (x113x) & (x254x)) + ((n_n5171) & (x33x) & (n_n5170) & (!x113x) & (!x254x)) + ((n_n5171) & (x33x) & (n_n5170) & (!x113x) & (x254x)) + ((n_n5171) & (x33x) & (n_n5170) & (x113x) & (!x254x)) + ((n_n5171) & (x33x) & (n_n5170) & (x113x) & (x254x)));
	assign n_n4663 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n390) & (x23x)));
	assign n_n4698 = (((i_9_) & (n_n532) & (n_n325) & (n_n535)));
	assign n_n4705 = (((!i_9_) & (n_n526) & (n_n325) & (n_n535)));
	assign n_n4805 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n325) & (x20x)));
	assign n_n4944 = (((i_9_) & (n_n526) & (n_n260) & (n_n464)));
	assign n_n5199 = (((!i_9_) & (n_n528) & (n_n130) & (n_n464)));
	assign n_n5260 = (((!i_5_) & (i_3_) & (!i_4_) & (x19x) & (n_n530)));
	assign n_n5272 = (((i_7_) & (i_8_) & (i_6_) & (x19x) & (n_n491)));
	assign n_n4501 = (((i_1_) & (!i_2_) & (i_0_) & (x20x) & (n_n500)));
	assign n_n4684 = (((i_9_) & (n_n390) & (n_n530) & (n_n464)));
	assign x426x = (((!i_9_) & (n_n390) & (n_n532) & (!n_n530) & (n_n464)) + ((!i_9_) & (n_n390) & (n_n532) & (n_n530) & (n_n464)) + ((i_9_) & (n_n390) & (!n_n532) & (n_n530) & (n_n464)) + ((i_9_) & (n_n390) & (n_n532) & (n_n530) & (n_n464)));
	assign n_n5221 = (((i_5_) & (i_3_) & (i_4_) & (x20x) & (n_n65)));
	assign n_n5220 = (((i_5_) & (i_3_) & (i_4_) & (x19x) & (n_n522)));
	assign n_n834 = (((!i_9_) & (!n_n524) & (n_n518) & (n_n526) & (n_n260)) + ((!i_9_) & (n_n524) & (n_n518) & (n_n526) & (n_n260)) + ((i_9_) & (!n_n524) & (n_n518) & (n_n526) & (n_n260)) + ((i_9_) & (n_n524) & (n_n518) & (!n_n526) & (n_n260)) + ((i_9_) & (n_n524) & (n_n518) & (n_n526) & (n_n260)));
	assign n_n1970 = (((!i_9_) & (!n_n532) & (n_n535) & (n_n195) & (n_n530)) + ((!i_9_) & (n_n532) & (n_n535) & (n_n195) & (!n_n530)) + ((!i_9_) & (n_n532) & (n_n535) & (n_n195) & (n_n530)) + ((i_9_) & (!n_n532) & (n_n535) & (n_n195) & (n_n530)) + ((i_9_) & (n_n532) & (n_n535) & (n_n195) & (n_n530)));
	assign n_n5134 = (((!i_7_) & (!i_8_) & (i_6_) & (x12x) & (n_n500)));
	assign n_n5125 = (((i_5_) & (i_3_) & (!i_4_) & (n_n130) & (x20x)));
	assign n_n5140 = (((!i_7_) & (i_8_) & (!i_6_) & (x12x) & (n_n500)));
	assign n_n5143 = (((!i_1_) & (i_2_) & (!i_0_) & (x23x) & (n_n500)));
	assign x13284x = (((!n_n5150) & (!n_n5149) & (!n_n5148) & (!n_n5140) & (n_n5143)) + ((!n_n5150) & (!n_n5149) & (!n_n5148) & (n_n5140) & (!n_n5143)) + ((!n_n5150) & (!n_n5149) & (!n_n5148) & (n_n5140) & (n_n5143)) + ((!n_n5150) & (!n_n5149) & (n_n5148) & (!n_n5140) & (!n_n5143)) + ((!n_n5150) & (!n_n5149) & (n_n5148) & (!n_n5140) & (n_n5143)) + ((!n_n5150) & (!n_n5149) & (n_n5148) & (n_n5140) & (!n_n5143)) + ((!n_n5150) & (!n_n5149) & (n_n5148) & (n_n5140) & (n_n5143)) + ((!n_n5150) & (n_n5149) & (!n_n5148) & (!n_n5140) & (!n_n5143)) + ((!n_n5150) & (n_n5149) & (!n_n5148) & (!n_n5140) & (n_n5143)) + ((!n_n5150) & (n_n5149) & (!n_n5148) & (n_n5140) & (!n_n5143)) + ((!n_n5150) & (n_n5149) & (!n_n5148) & (n_n5140) & (n_n5143)) + ((!n_n5150) & (n_n5149) & (n_n5148) & (!n_n5140) & (!n_n5143)) + ((!n_n5150) & (n_n5149) & (n_n5148) & (!n_n5140) & (n_n5143)) + ((!n_n5150) & (n_n5149) & (n_n5148) & (n_n5140) & (!n_n5143)) + ((!n_n5150) & (n_n5149) & (n_n5148) & (n_n5140) & (n_n5143)) + ((n_n5150) & (!n_n5149) & (!n_n5148) & (!n_n5140) & (!n_n5143)) + ((n_n5150) & (!n_n5149) & (!n_n5148) & (!n_n5140) & (n_n5143)) + ((n_n5150) & (!n_n5149) & (!n_n5148) & (n_n5140) & (!n_n5143)) + ((n_n5150) & (!n_n5149) & (!n_n5148) & (n_n5140) & (n_n5143)) + ((n_n5150) & (!n_n5149) & (n_n5148) & (!n_n5140) & (!n_n5143)) + ((n_n5150) & (!n_n5149) & (n_n5148) & (!n_n5140) & (n_n5143)) + ((n_n5150) & (!n_n5149) & (n_n5148) & (n_n5140) & (!n_n5143)) + ((n_n5150) & (!n_n5149) & (n_n5148) & (n_n5140) & (n_n5143)) + ((n_n5150) & (n_n5149) & (!n_n5148) & (!n_n5140) & (!n_n5143)) + ((n_n5150) & (n_n5149) & (!n_n5148) & (!n_n5140) & (n_n5143)) + ((n_n5150) & (n_n5149) & (!n_n5148) & (n_n5140) & (!n_n5143)) + ((n_n5150) & (n_n5149) & (!n_n5148) & (n_n5140) & (n_n5143)) + ((n_n5150) & (n_n5149) & (n_n5148) & (!n_n5140) & (!n_n5143)) + ((n_n5150) & (n_n5149) & (n_n5148) & (!n_n5140) & (n_n5143)) + ((n_n5150) & (n_n5149) & (n_n5148) & (n_n5140) & (!n_n5143)) + ((n_n5150) & (n_n5149) & (n_n5148) & (n_n5140) & (n_n5143)));
	assign n_n4039 = (((!n_n5142) & (!n_n5146) & (!n_n5135) & (!n_n5147) & (x13284x)) + ((!n_n5142) & (!n_n5146) & (!n_n5135) & (n_n5147) & (!x13284x)) + ((!n_n5142) & (!n_n5146) & (!n_n5135) & (n_n5147) & (x13284x)) + ((!n_n5142) & (!n_n5146) & (n_n5135) & (!n_n5147) & (!x13284x)) + ((!n_n5142) & (!n_n5146) & (n_n5135) & (!n_n5147) & (x13284x)) + ((!n_n5142) & (!n_n5146) & (n_n5135) & (n_n5147) & (!x13284x)) + ((!n_n5142) & (!n_n5146) & (n_n5135) & (n_n5147) & (x13284x)) + ((!n_n5142) & (n_n5146) & (!n_n5135) & (!n_n5147) & (!x13284x)) + ((!n_n5142) & (n_n5146) & (!n_n5135) & (!n_n5147) & (x13284x)) + ((!n_n5142) & (n_n5146) & (!n_n5135) & (n_n5147) & (!x13284x)) + ((!n_n5142) & (n_n5146) & (!n_n5135) & (n_n5147) & (x13284x)) + ((!n_n5142) & (n_n5146) & (n_n5135) & (!n_n5147) & (!x13284x)) + ((!n_n5142) & (n_n5146) & (n_n5135) & (!n_n5147) & (x13284x)) + ((!n_n5142) & (n_n5146) & (n_n5135) & (n_n5147) & (!x13284x)) + ((!n_n5142) & (n_n5146) & (n_n5135) & (n_n5147) & (x13284x)) + ((n_n5142) & (!n_n5146) & (!n_n5135) & (!n_n5147) & (!x13284x)) + ((n_n5142) & (!n_n5146) & (!n_n5135) & (!n_n5147) & (x13284x)) + ((n_n5142) & (!n_n5146) & (!n_n5135) & (n_n5147) & (!x13284x)) + ((n_n5142) & (!n_n5146) & (!n_n5135) & (n_n5147) & (x13284x)) + ((n_n5142) & (!n_n5146) & (n_n5135) & (!n_n5147) & (!x13284x)) + ((n_n5142) & (!n_n5146) & (n_n5135) & (!n_n5147) & (x13284x)) + ((n_n5142) & (!n_n5146) & (n_n5135) & (n_n5147) & (!x13284x)) + ((n_n5142) & (!n_n5146) & (n_n5135) & (n_n5147) & (x13284x)) + ((n_n5142) & (n_n5146) & (!n_n5135) & (!n_n5147) & (!x13284x)) + ((n_n5142) & (n_n5146) & (!n_n5135) & (!n_n5147) & (x13284x)) + ((n_n5142) & (n_n5146) & (!n_n5135) & (n_n5147) & (!x13284x)) + ((n_n5142) & (n_n5146) & (!n_n5135) & (n_n5147) & (x13284x)) + ((n_n5142) & (n_n5146) & (n_n5135) & (!n_n5147) & (!x13284x)) + ((n_n5142) & (n_n5146) & (n_n5135) & (!n_n5147) & (x13284x)) + ((n_n5142) & (n_n5146) & (n_n5135) & (n_n5147) & (!x13284x)) + ((n_n5142) & (n_n5146) & (n_n5135) & (n_n5147) & (x13284x)));
	assign x22202x = (((!n_n5161) & (!n_n5157) & (!n_n5159) & (!n_n5160)));
	assign n_n4038 = (((!n_n5152) & (!n_n5153) & (!x358x) & (!n_n5151) & (!x22202x)) + ((!n_n5152) & (!n_n5153) & (!x358x) & (n_n5151) & (!x22202x)) + ((!n_n5152) & (!n_n5153) & (!x358x) & (n_n5151) & (x22202x)) + ((!n_n5152) & (!n_n5153) & (x358x) & (!n_n5151) & (!x22202x)) + ((!n_n5152) & (!n_n5153) & (x358x) & (!n_n5151) & (x22202x)) + ((!n_n5152) & (!n_n5153) & (x358x) & (n_n5151) & (!x22202x)) + ((!n_n5152) & (!n_n5153) & (x358x) & (n_n5151) & (x22202x)) + ((!n_n5152) & (n_n5153) & (!x358x) & (!n_n5151) & (!x22202x)) + ((!n_n5152) & (n_n5153) & (!x358x) & (!n_n5151) & (x22202x)) + ((!n_n5152) & (n_n5153) & (!x358x) & (n_n5151) & (!x22202x)) + ((!n_n5152) & (n_n5153) & (!x358x) & (n_n5151) & (x22202x)) + ((!n_n5152) & (n_n5153) & (x358x) & (!n_n5151) & (!x22202x)) + ((!n_n5152) & (n_n5153) & (x358x) & (!n_n5151) & (x22202x)) + ((!n_n5152) & (n_n5153) & (x358x) & (n_n5151) & (!x22202x)) + ((!n_n5152) & (n_n5153) & (x358x) & (n_n5151) & (x22202x)) + ((n_n5152) & (!n_n5153) & (!x358x) & (!n_n5151) & (!x22202x)) + ((n_n5152) & (!n_n5153) & (!x358x) & (!n_n5151) & (x22202x)) + ((n_n5152) & (!n_n5153) & (!x358x) & (n_n5151) & (!x22202x)) + ((n_n5152) & (!n_n5153) & (!x358x) & (n_n5151) & (x22202x)) + ((n_n5152) & (!n_n5153) & (x358x) & (!n_n5151) & (!x22202x)) + ((n_n5152) & (!n_n5153) & (x358x) & (!n_n5151) & (x22202x)) + ((n_n5152) & (!n_n5153) & (x358x) & (n_n5151) & (!x22202x)) + ((n_n5152) & (!n_n5153) & (x358x) & (n_n5151) & (x22202x)) + ((n_n5152) & (n_n5153) & (!x358x) & (!n_n5151) & (!x22202x)) + ((n_n5152) & (n_n5153) & (!x358x) & (!n_n5151) & (x22202x)) + ((n_n5152) & (n_n5153) & (!x358x) & (n_n5151) & (!x22202x)) + ((n_n5152) & (n_n5153) & (!x358x) & (n_n5151) & (x22202x)) + ((n_n5152) & (n_n5153) & (x358x) & (!n_n5151) & (!x22202x)) + ((n_n5152) & (n_n5153) & (x358x) & (!n_n5151) & (x22202x)) + ((n_n5152) & (n_n5153) & (x358x) & (n_n5151) & (!x22202x)) + ((n_n5152) & (n_n5153) & (x358x) & (n_n5151) & (x22202x)));
	assign n_n5196 = (((!i_7_) & (i_8_) & (i_6_) & (x12x) & (n_n464)));
	assign x13302x = (((!n_n534) & (!x12x) & (!n_n464) & (!n_n5195) & (n_n2670)) + ((!n_n534) & (!x12x) & (!n_n464) & (n_n5195) & (!n_n2670)) + ((!n_n534) & (!x12x) & (!n_n464) & (n_n5195) & (n_n2670)) + ((!n_n534) & (!x12x) & (n_n464) & (!n_n5195) & (n_n2670)) + ((!n_n534) & (!x12x) & (n_n464) & (n_n5195) & (!n_n2670)) + ((!n_n534) & (!x12x) & (n_n464) & (n_n5195) & (n_n2670)) + ((!n_n534) & (x12x) & (!n_n464) & (!n_n5195) & (n_n2670)) + ((!n_n534) & (x12x) & (!n_n464) & (n_n5195) & (!n_n2670)) + ((!n_n534) & (x12x) & (!n_n464) & (n_n5195) & (n_n2670)) + ((!n_n534) & (x12x) & (n_n464) & (!n_n5195) & (n_n2670)) + ((!n_n534) & (x12x) & (n_n464) & (n_n5195) & (!n_n2670)) + ((!n_n534) & (x12x) & (n_n464) & (n_n5195) & (n_n2670)) + ((n_n534) & (!x12x) & (!n_n464) & (!n_n5195) & (n_n2670)) + ((n_n534) & (!x12x) & (!n_n464) & (n_n5195) & (!n_n2670)) + ((n_n534) & (!x12x) & (!n_n464) & (n_n5195) & (n_n2670)) + ((n_n534) & (!x12x) & (n_n464) & (!n_n5195) & (n_n2670)) + ((n_n534) & (!x12x) & (n_n464) & (n_n5195) & (!n_n2670)) + ((n_n534) & (!x12x) & (n_n464) & (n_n5195) & (n_n2670)) + ((n_n534) & (x12x) & (!n_n464) & (!n_n5195) & (n_n2670)) + ((n_n534) & (x12x) & (!n_n464) & (n_n5195) & (!n_n2670)) + ((n_n534) & (x12x) & (!n_n464) & (n_n5195) & (n_n2670)) + ((n_n534) & (x12x) & (n_n464) & (!n_n5195) & (!n_n2670)) + ((n_n534) & (x12x) & (n_n464) & (!n_n5195) & (n_n2670)) + ((n_n534) & (x12x) & (n_n464) & (n_n5195) & (!n_n2670)) + ((n_n534) & (x12x) & (n_n464) & (n_n5195) & (n_n2670)));
	assign x13303x = (((!n_n5187) & (!n_n5189) & (!n_n5188) & (!n_n5196) & (x13302x)) + ((!n_n5187) & (!n_n5189) & (!n_n5188) & (n_n5196) & (!x13302x)) + ((!n_n5187) & (!n_n5189) & (!n_n5188) & (n_n5196) & (x13302x)) + ((!n_n5187) & (!n_n5189) & (n_n5188) & (!n_n5196) & (!x13302x)) + ((!n_n5187) & (!n_n5189) & (n_n5188) & (!n_n5196) & (x13302x)) + ((!n_n5187) & (!n_n5189) & (n_n5188) & (n_n5196) & (!x13302x)) + ((!n_n5187) & (!n_n5189) & (n_n5188) & (n_n5196) & (x13302x)) + ((!n_n5187) & (n_n5189) & (!n_n5188) & (!n_n5196) & (!x13302x)) + ((!n_n5187) & (n_n5189) & (!n_n5188) & (!n_n5196) & (x13302x)) + ((!n_n5187) & (n_n5189) & (!n_n5188) & (n_n5196) & (!x13302x)) + ((!n_n5187) & (n_n5189) & (!n_n5188) & (n_n5196) & (x13302x)) + ((!n_n5187) & (n_n5189) & (n_n5188) & (!n_n5196) & (!x13302x)) + ((!n_n5187) & (n_n5189) & (n_n5188) & (!n_n5196) & (x13302x)) + ((!n_n5187) & (n_n5189) & (n_n5188) & (n_n5196) & (!x13302x)) + ((!n_n5187) & (n_n5189) & (n_n5188) & (n_n5196) & (x13302x)) + ((n_n5187) & (!n_n5189) & (!n_n5188) & (!n_n5196) & (!x13302x)) + ((n_n5187) & (!n_n5189) & (!n_n5188) & (!n_n5196) & (x13302x)) + ((n_n5187) & (!n_n5189) & (!n_n5188) & (n_n5196) & (!x13302x)) + ((n_n5187) & (!n_n5189) & (!n_n5188) & (n_n5196) & (x13302x)) + ((n_n5187) & (!n_n5189) & (n_n5188) & (!n_n5196) & (!x13302x)) + ((n_n5187) & (!n_n5189) & (n_n5188) & (!n_n5196) & (x13302x)) + ((n_n5187) & (!n_n5189) & (n_n5188) & (n_n5196) & (!x13302x)) + ((n_n5187) & (!n_n5189) & (n_n5188) & (n_n5196) & (x13302x)) + ((n_n5187) & (n_n5189) & (!n_n5188) & (!n_n5196) & (!x13302x)) + ((n_n5187) & (n_n5189) & (!n_n5188) & (!n_n5196) & (x13302x)) + ((n_n5187) & (n_n5189) & (!n_n5188) & (n_n5196) & (!x13302x)) + ((n_n5187) & (n_n5189) & (!n_n5188) & (n_n5196) & (x13302x)) + ((n_n5187) & (n_n5189) & (n_n5188) & (!n_n5196) & (!x13302x)) + ((n_n5187) & (n_n5189) & (n_n5188) & (!n_n5196) & (x13302x)) + ((n_n5187) & (n_n5189) & (n_n5188) & (n_n5196) & (!x13302x)) + ((n_n5187) & (n_n5189) & (n_n5188) & (n_n5196) & (x13302x)));
	assign x144x = (((!n_n524) & (!n_n535) & (!x12x) & (!n_n4148) & (x13306x)) + ((!n_n524) & (!n_n535) & (!x12x) & (n_n4148) & (!x13306x)) + ((!n_n524) & (!n_n535) & (!x12x) & (n_n4148) & (x13306x)) + ((!n_n524) & (!n_n535) & (x12x) & (!n_n4148) & (x13306x)) + ((!n_n524) & (!n_n535) & (x12x) & (n_n4148) & (!x13306x)) + ((!n_n524) & (!n_n535) & (x12x) & (n_n4148) & (x13306x)) + ((!n_n524) & (n_n535) & (!x12x) & (!n_n4148) & (x13306x)) + ((!n_n524) & (n_n535) & (!x12x) & (n_n4148) & (!x13306x)) + ((!n_n524) & (n_n535) & (!x12x) & (n_n4148) & (x13306x)) + ((!n_n524) & (n_n535) & (x12x) & (!n_n4148) & (x13306x)) + ((!n_n524) & (n_n535) & (x12x) & (n_n4148) & (!x13306x)) + ((!n_n524) & (n_n535) & (x12x) & (n_n4148) & (x13306x)) + ((n_n524) & (!n_n535) & (!x12x) & (!n_n4148) & (x13306x)) + ((n_n524) & (!n_n535) & (!x12x) & (n_n4148) & (!x13306x)) + ((n_n524) & (!n_n535) & (!x12x) & (n_n4148) & (x13306x)) + ((n_n524) & (!n_n535) & (x12x) & (!n_n4148) & (x13306x)) + ((n_n524) & (!n_n535) & (x12x) & (n_n4148) & (!x13306x)) + ((n_n524) & (!n_n535) & (x12x) & (n_n4148) & (x13306x)) + ((n_n524) & (n_n535) & (!x12x) & (!n_n4148) & (x13306x)) + ((n_n524) & (n_n535) & (!x12x) & (n_n4148) & (!x13306x)) + ((n_n524) & (n_n535) & (!x12x) & (n_n4148) & (x13306x)) + ((n_n524) & (n_n535) & (x12x) & (!n_n4148) & (!x13306x)) + ((n_n524) & (n_n535) & (x12x) & (!n_n4148) & (x13306x)) + ((n_n524) & (n_n535) & (x12x) & (n_n4148) & (!x13306x)) + ((n_n524) & (n_n535) & (x12x) & (n_n4148) & (x13306x)));
	assign x13317x = (((!n_n5086) & (!n_n5087) & (!n_n5095) & (!n_n5106) & (x144x)) + ((!n_n5086) & (!n_n5087) & (!n_n5095) & (n_n5106) & (!x144x)) + ((!n_n5086) & (!n_n5087) & (!n_n5095) & (n_n5106) & (x144x)) + ((!n_n5086) & (!n_n5087) & (n_n5095) & (!n_n5106) & (!x144x)) + ((!n_n5086) & (!n_n5087) & (n_n5095) & (!n_n5106) & (x144x)) + ((!n_n5086) & (!n_n5087) & (n_n5095) & (n_n5106) & (!x144x)) + ((!n_n5086) & (!n_n5087) & (n_n5095) & (n_n5106) & (x144x)) + ((!n_n5086) & (n_n5087) & (!n_n5095) & (!n_n5106) & (!x144x)) + ((!n_n5086) & (n_n5087) & (!n_n5095) & (!n_n5106) & (x144x)) + ((!n_n5086) & (n_n5087) & (!n_n5095) & (n_n5106) & (!x144x)) + ((!n_n5086) & (n_n5087) & (!n_n5095) & (n_n5106) & (x144x)) + ((!n_n5086) & (n_n5087) & (n_n5095) & (!n_n5106) & (!x144x)) + ((!n_n5086) & (n_n5087) & (n_n5095) & (!n_n5106) & (x144x)) + ((!n_n5086) & (n_n5087) & (n_n5095) & (n_n5106) & (!x144x)) + ((!n_n5086) & (n_n5087) & (n_n5095) & (n_n5106) & (x144x)) + ((n_n5086) & (!n_n5087) & (!n_n5095) & (!n_n5106) & (!x144x)) + ((n_n5086) & (!n_n5087) & (!n_n5095) & (!n_n5106) & (x144x)) + ((n_n5086) & (!n_n5087) & (!n_n5095) & (n_n5106) & (!x144x)) + ((n_n5086) & (!n_n5087) & (!n_n5095) & (n_n5106) & (x144x)) + ((n_n5086) & (!n_n5087) & (n_n5095) & (!n_n5106) & (!x144x)) + ((n_n5086) & (!n_n5087) & (n_n5095) & (!n_n5106) & (x144x)) + ((n_n5086) & (!n_n5087) & (n_n5095) & (n_n5106) & (!x144x)) + ((n_n5086) & (!n_n5087) & (n_n5095) & (n_n5106) & (x144x)) + ((n_n5086) & (n_n5087) & (!n_n5095) & (!n_n5106) & (!x144x)) + ((n_n5086) & (n_n5087) & (!n_n5095) & (!n_n5106) & (x144x)) + ((n_n5086) & (n_n5087) & (!n_n5095) & (n_n5106) & (!x144x)) + ((n_n5086) & (n_n5087) & (!n_n5095) & (n_n5106) & (x144x)) + ((n_n5086) & (n_n5087) & (n_n5095) & (!n_n5106) & (!x144x)) + ((n_n5086) & (n_n5087) & (n_n5095) & (!n_n5106) & (x144x)) + ((n_n5086) & (n_n5087) & (n_n5095) & (n_n5106) & (!x144x)) + ((n_n5086) & (n_n5087) & (n_n5095) & (n_n5106) & (x144x)));
	assign n_n4041 = (((!n_n5111) & (!n_n5110) & (!n_n5113) & (!n_n4144) & (x11915x)) + ((!n_n5111) & (!n_n5110) & (!n_n5113) & (n_n4144) & (!x11915x)) + ((!n_n5111) & (!n_n5110) & (!n_n5113) & (n_n4144) & (x11915x)) + ((!n_n5111) & (!n_n5110) & (n_n5113) & (!n_n4144) & (!x11915x)) + ((!n_n5111) & (!n_n5110) & (n_n5113) & (!n_n4144) & (x11915x)) + ((!n_n5111) & (!n_n5110) & (n_n5113) & (n_n4144) & (!x11915x)) + ((!n_n5111) & (!n_n5110) & (n_n5113) & (n_n4144) & (x11915x)) + ((!n_n5111) & (n_n5110) & (!n_n5113) & (!n_n4144) & (!x11915x)) + ((!n_n5111) & (n_n5110) & (!n_n5113) & (!n_n4144) & (x11915x)) + ((!n_n5111) & (n_n5110) & (!n_n5113) & (n_n4144) & (!x11915x)) + ((!n_n5111) & (n_n5110) & (!n_n5113) & (n_n4144) & (x11915x)) + ((!n_n5111) & (n_n5110) & (n_n5113) & (!n_n4144) & (!x11915x)) + ((!n_n5111) & (n_n5110) & (n_n5113) & (!n_n4144) & (x11915x)) + ((!n_n5111) & (n_n5110) & (n_n5113) & (n_n4144) & (!x11915x)) + ((!n_n5111) & (n_n5110) & (n_n5113) & (n_n4144) & (x11915x)) + ((n_n5111) & (!n_n5110) & (!n_n5113) & (!n_n4144) & (!x11915x)) + ((n_n5111) & (!n_n5110) & (!n_n5113) & (!n_n4144) & (x11915x)) + ((n_n5111) & (!n_n5110) & (!n_n5113) & (n_n4144) & (!x11915x)) + ((n_n5111) & (!n_n5110) & (!n_n5113) & (n_n4144) & (x11915x)) + ((n_n5111) & (!n_n5110) & (n_n5113) & (!n_n4144) & (!x11915x)) + ((n_n5111) & (!n_n5110) & (n_n5113) & (!n_n4144) & (x11915x)) + ((n_n5111) & (!n_n5110) & (n_n5113) & (n_n4144) & (!x11915x)) + ((n_n5111) & (!n_n5110) & (n_n5113) & (n_n4144) & (x11915x)) + ((n_n5111) & (n_n5110) & (!n_n5113) & (!n_n4144) & (!x11915x)) + ((n_n5111) & (n_n5110) & (!n_n5113) & (!n_n4144) & (x11915x)) + ((n_n5111) & (n_n5110) & (!n_n5113) & (n_n4144) & (!x11915x)) + ((n_n5111) & (n_n5110) & (!n_n5113) & (n_n4144) & (x11915x)) + ((n_n5111) & (n_n5110) & (n_n5113) & (!n_n4144) & (!x11915x)) + ((n_n5111) & (n_n5110) & (n_n5113) & (!n_n4144) & (x11915x)) + ((n_n5111) & (n_n5110) & (n_n5113) & (n_n4144) & (!x11915x)) + ((n_n5111) & (n_n5110) & (n_n5113) & (n_n4144) & (x11915x)));
	assign x279x = (((!i_9_) & (n_n518) & (n_n534) & (!n_n130) & (x12x)) + ((!i_9_) & (n_n518) & (n_n534) & (n_n130) & (!x12x)) + ((!i_9_) & (n_n518) & (n_n534) & (n_n130) & (x12x)) + ((i_9_) & (n_n518) & (n_n534) & (!n_n130) & (x12x)) + ((i_9_) & (n_n518) & (n_n534) & (n_n130) & (x12x)));
	assign x13314x = (((!n_n5099) & (!n_n5085) & (!n_n5100) & (n_n5098)) + ((!n_n5099) & (!n_n5085) & (n_n5100) & (!n_n5098)) + ((!n_n5099) & (!n_n5085) & (n_n5100) & (n_n5098)) + ((!n_n5099) & (n_n5085) & (!n_n5100) & (!n_n5098)) + ((!n_n5099) & (n_n5085) & (!n_n5100) & (n_n5098)) + ((!n_n5099) & (n_n5085) & (n_n5100) & (!n_n5098)) + ((!n_n5099) & (n_n5085) & (n_n5100) & (n_n5098)) + ((n_n5099) & (!n_n5085) & (!n_n5100) & (!n_n5098)) + ((n_n5099) & (!n_n5085) & (!n_n5100) & (n_n5098)) + ((n_n5099) & (!n_n5085) & (n_n5100) & (!n_n5098)) + ((n_n5099) & (!n_n5085) & (n_n5100) & (n_n5098)) + ((n_n5099) & (n_n5085) & (!n_n5100) & (!n_n5098)) + ((n_n5099) & (n_n5085) & (!n_n5100) & (n_n5098)) + ((n_n5099) & (n_n5085) & (n_n5100) & (!n_n5098)) + ((n_n5099) & (n_n5085) & (n_n5100) & (n_n5098)));
	assign n_n4002 = (((!x289x) & (!x13317x) & (!n_n4041) & (!x279x) & (x13314x)) + ((!x289x) & (!x13317x) & (!n_n4041) & (x279x) & (!x13314x)) + ((!x289x) & (!x13317x) & (!n_n4041) & (x279x) & (x13314x)) + ((!x289x) & (!x13317x) & (n_n4041) & (!x279x) & (!x13314x)) + ((!x289x) & (!x13317x) & (n_n4041) & (!x279x) & (x13314x)) + ((!x289x) & (!x13317x) & (n_n4041) & (x279x) & (!x13314x)) + ((!x289x) & (!x13317x) & (n_n4041) & (x279x) & (x13314x)) + ((!x289x) & (x13317x) & (!n_n4041) & (!x279x) & (!x13314x)) + ((!x289x) & (x13317x) & (!n_n4041) & (!x279x) & (x13314x)) + ((!x289x) & (x13317x) & (!n_n4041) & (x279x) & (!x13314x)) + ((!x289x) & (x13317x) & (!n_n4041) & (x279x) & (x13314x)) + ((!x289x) & (x13317x) & (n_n4041) & (!x279x) & (!x13314x)) + ((!x289x) & (x13317x) & (n_n4041) & (!x279x) & (x13314x)) + ((!x289x) & (x13317x) & (n_n4041) & (x279x) & (!x13314x)) + ((!x289x) & (x13317x) & (n_n4041) & (x279x) & (x13314x)) + ((x289x) & (!x13317x) & (!n_n4041) & (!x279x) & (!x13314x)) + ((x289x) & (!x13317x) & (!n_n4041) & (!x279x) & (x13314x)) + ((x289x) & (!x13317x) & (!n_n4041) & (x279x) & (!x13314x)) + ((x289x) & (!x13317x) & (!n_n4041) & (x279x) & (x13314x)) + ((x289x) & (!x13317x) & (n_n4041) & (!x279x) & (!x13314x)) + ((x289x) & (!x13317x) & (n_n4041) & (!x279x) & (x13314x)) + ((x289x) & (!x13317x) & (n_n4041) & (x279x) & (!x13314x)) + ((x289x) & (!x13317x) & (n_n4041) & (x279x) & (x13314x)) + ((x289x) & (x13317x) & (!n_n4041) & (!x279x) & (!x13314x)) + ((x289x) & (x13317x) & (!n_n4041) & (!x279x) & (x13314x)) + ((x289x) & (x13317x) & (!n_n4041) & (x279x) & (!x13314x)) + ((x289x) & (x13317x) & (!n_n4041) & (x279x) & (x13314x)) + ((x289x) & (x13317x) & (n_n4041) & (!x279x) & (!x13314x)) + ((x289x) & (x13317x) & (n_n4041) & (!x279x) & (x13314x)) + ((x289x) & (x13317x) & (n_n4041) & (x279x) & (!x13314x)) + ((x289x) & (x13317x) & (n_n4041) & (x279x) & (x13314x)));
	assign n_n5126 = (((i_5_) & (i_3_) & (!i_4_) & (n_n520) & (x12x)));
	assign x13322x = (((!n_n5130) & (!n_n5124) & (!n_n5127) & (n_n5126)) + ((!n_n5130) & (!n_n5124) & (n_n5127) & (!n_n5126)) + ((!n_n5130) & (!n_n5124) & (n_n5127) & (n_n5126)) + ((!n_n5130) & (n_n5124) & (!n_n5127) & (!n_n5126)) + ((!n_n5130) & (n_n5124) & (!n_n5127) & (n_n5126)) + ((!n_n5130) & (n_n5124) & (n_n5127) & (!n_n5126)) + ((!n_n5130) & (n_n5124) & (n_n5127) & (n_n5126)) + ((n_n5130) & (!n_n5124) & (!n_n5127) & (!n_n5126)) + ((n_n5130) & (!n_n5124) & (!n_n5127) & (n_n5126)) + ((n_n5130) & (!n_n5124) & (n_n5127) & (!n_n5126)) + ((n_n5130) & (!n_n5124) & (n_n5127) & (n_n5126)) + ((n_n5130) & (n_n5124) & (!n_n5127) & (!n_n5126)) + ((n_n5130) & (n_n5124) & (!n_n5127) & (n_n5126)) + ((n_n5130) & (n_n5124) & (n_n5127) & (!n_n5126)) + ((n_n5130) & (n_n5124) & (n_n5127) & (n_n5126)));
	assign x13323x = (((!n_n5121) & (!n_n5122) & (!n_n5118) & (!n_n5134) & (n_n5125)) + ((!n_n5121) & (!n_n5122) & (!n_n5118) & (n_n5134) & (!n_n5125)) + ((!n_n5121) & (!n_n5122) & (!n_n5118) & (n_n5134) & (n_n5125)) + ((!n_n5121) & (!n_n5122) & (n_n5118) & (!n_n5134) & (!n_n5125)) + ((!n_n5121) & (!n_n5122) & (n_n5118) & (!n_n5134) & (n_n5125)) + ((!n_n5121) & (!n_n5122) & (n_n5118) & (n_n5134) & (!n_n5125)) + ((!n_n5121) & (!n_n5122) & (n_n5118) & (n_n5134) & (n_n5125)) + ((!n_n5121) & (n_n5122) & (!n_n5118) & (!n_n5134) & (!n_n5125)) + ((!n_n5121) & (n_n5122) & (!n_n5118) & (!n_n5134) & (n_n5125)) + ((!n_n5121) & (n_n5122) & (!n_n5118) & (n_n5134) & (!n_n5125)) + ((!n_n5121) & (n_n5122) & (!n_n5118) & (n_n5134) & (n_n5125)) + ((!n_n5121) & (n_n5122) & (n_n5118) & (!n_n5134) & (!n_n5125)) + ((!n_n5121) & (n_n5122) & (n_n5118) & (!n_n5134) & (n_n5125)) + ((!n_n5121) & (n_n5122) & (n_n5118) & (n_n5134) & (!n_n5125)) + ((!n_n5121) & (n_n5122) & (n_n5118) & (n_n5134) & (n_n5125)) + ((n_n5121) & (!n_n5122) & (!n_n5118) & (!n_n5134) & (!n_n5125)) + ((n_n5121) & (!n_n5122) & (!n_n5118) & (!n_n5134) & (n_n5125)) + ((n_n5121) & (!n_n5122) & (!n_n5118) & (n_n5134) & (!n_n5125)) + ((n_n5121) & (!n_n5122) & (!n_n5118) & (n_n5134) & (n_n5125)) + ((n_n5121) & (!n_n5122) & (n_n5118) & (!n_n5134) & (!n_n5125)) + ((n_n5121) & (!n_n5122) & (n_n5118) & (!n_n5134) & (n_n5125)) + ((n_n5121) & (!n_n5122) & (n_n5118) & (n_n5134) & (!n_n5125)) + ((n_n5121) & (!n_n5122) & (n_n5118) & (n_n5134) & (n_n5125)) + ((n_n5121) & (n_n5122) & (!n_n5118) & (!n_n5134) & (!n_n5125)) + ((n_n5121) & (n_n5122) & (!n_n5118) & (!n_n5134) & (n_n5125)) + ((n_n5121) & (n_n5122) & (!n_n5118) & (n_n5134) & (!n_n5125)) + ((n_n5121) & (n_n5122) & (!n_n5118) & (n_n5134) & (n_n5125)) + ((n_n5121) & (n_n5122) & (n_n5118) & (!n_n5134) & (!n_n5125)) + ((n_n5121) & (n_n5122) & (n_n5118) & (!n_n5134) & (n_n5125)) + ((n_n5121) & (n_n5122) & (n_n5118) & (n_n5134) & (!n_n5125)) + ((n_n5121) & (n_n5122) & (n_n5118) & (n_n5134) & (n_n5125)));
	assign x13326x = (((!n_n4039) & (!n_n4038) & (!x13322x) & (x13323x)) + ((!n_n4039) & (!n_n4038) & (x13322x) & (!x13323x)) + ((!n_n4039) & (!n_n4038) & (x13322x) & (x13323x)) + ((!n_n4039) & (n_n4038) & (!x13322x) & (!x13323x)) + ((!n_n4039) & (n_n4038) & (!x13322x) & (x13323x)) + ((!n_n4039) & (n_n4038) & (x13322x) & (!x13323x)) + ((!n_n4039) & (n_n4038) & (x13322x) & (x13323x)) + ((n_n4039) & (!n_n4038) & (!x13322x) & (!x13323x)) + ((n_n4039) & (!n_n4038) & (!x13322x) & (x13323x)) + ((n_n4039) & (!n_n4038) & (x13322x) & (!x13323x)) + ((n_n4039) & (!n_n4038) & (x13322x) & (x13323x)) + ((n_n4039) & (n_n4038) & (!x13322x) & (!x13323x)) + ((n_n4039) & (n_n4038) & (!x13322x) & (x13323x)) + ((n_n4039) & (n_n4038) & (x13322x) & (!x13323x)) + ((n_n4039) & (n_n4038) & (x13322x) & (x13323x)));
	assign n_n4036 = (((!n_n5174) & (!n_n5184) & (!n_n5185) & (!n_n5183) & (x13293x)) + ((!n_n5174) & (!n_n5184) & (!n_n5185) & (n_n5183) & (!x13293x)) + ((!n_n5174) & (!n_n5184) & (!n_n5185) & (n_n5183) & (x13293x)) + ((!n_n5174) & (!n_n5184) & (n_n5185) & (!n_n5183) & (!x13293x)) + ((!n_n5174) & (!n_n5184) & (n_n5185) & (!n_n5183) & (x13293x)) + ((!n_n5174) & (!n_n5184) & (n_n5185) & (n_n5183) & (!x13293x)) + ((!n_n5174) & (!n_n5184) & (n_n5185) & (n_n5183) & (x13293x)) + ((!n_n5174) & (n_n5184) & (!n_n5185) & (!n_n5183) & (!x13293x)) + ((!n_n5174) & (n_n5184) & (!n_n5185) & (!n_n5183) & (x13293x)) + ((!n_n5174) & (n_n5184) & (!n_n5185) & (n_n5183) & (!x13293x)) + ((!n_n5174) & (n_n5184) & (!n_n5185) & (n_n5183) & (x13293x)) + ((!n_n5174) & (n_n5184) & (n_n5185) & (!n_n5183) & (!x13293x)) + ((!n_n5174) & (n_n5184) & (n_n5185) & (!n_n5183) & (x13293x)) + ((!n_n5174) & (n_n5184) & (n_n5185) & (n_n5183) & (!x13293x)) + ((!n_n5174) & (n_n5184) & (n_n5185) & (n_n5183) & (x13293x)) + ((n_n5174) & (!n_n5184) & (!n_n5185) & (!n_n5183) & (!x13293x)) + ((n_n5174) & (!n_n5184) & (!n_n5185) & (!n_n5183) & (x13293x)) + ((n_n5174) & (!n_n5184) & (!n_n5185) & (n_n5183) & (!x13293x)) + ((n_n5174) & (!n_n5184) & (!n_n5185) & (n_n5183) & (x13293x)) + ((n_n5174) & (!n_n5184) & (n_n5185) & (!n_n5183) & (!x13293x)) + ((n_n5174) & (!n_n5184) & (n_n5185) & (!n_n5183) & (x13293x)) + ((n_n5174) & (!n_n5184) & (n_n5185) & (n_n5183) & (!x13293x)) + ((n_n5174) & (!n_n5184) & (n_n5185) & (n_n5183) & (x13293x)) + ((n_n5174) & (n_n5184) & (!n_n5185) & (!n_n5183) & (!x13293x)) + ((n_n5174) & (n_n5184) & (!n_n5185) & (!n_n5183) & (x13293x)) + ((n_n5174) & (n_n5184) & (!n_n5185) & (n_n5183) & (!x13293x)) + ((n_n5174) & (n_n5184) & (!n_n5185) & (n_n5183) & (x13293x)) + ((n_n5174) & (n_n5184) & (n_n5185) & (!n_n5183) & (!x13293x)) + ((n_n5174) & (n_n5184) & (n_n5185) & (!n_n5183) & (x13293x)) + ((n_n5174) & (n_n5184) & (n_n5185) & (n_n5183) & (!x13293x)) + ((n_n5174) & (n_n5184) & (n_n5185) & (n_n5183) & (x13293x)));
	assign n_n4037 = (((!n_n5162) & (!n_n5168) & (!n_n5169) & (!x33x) & (x13296x)) + ((!n_n5162) & (!n_n5168) & (!n_n5169) & (x33x) & (!x13296x)) + ((!n_n5162) & (!n_n5168) & (!n_n5169) & (x33x) & (x13296x)) + ((!n_n5162) & (!n_n5168) & (n_n5169) & (!x33x) & (!x13296x)) + ((!n_n5162) & (!n_n5168) & (n_n5169) & (!x33x) & (x13296x)) + ((!n_n5162) & (!n_n5168) & (n_n5169) & (x33x) & (!x13296x)) + ((!n_n5162) & (!n_n5168) & (n_n5169) & (x33x) & (x13296x)) + ((!n_n5162) & (n_n5168) & (!n_n5169) & (!x33x) & (!x13296x)) + ((!n_n5162) & (n_n5168) & (!n_n5169) & (!x33x) & (x13296x)) + ((!n_n5162) & (n_n5168) & (!n_n5169) & (x33x) & (!x13296x)) + ((!n_n5162) & (n_n5168) & (!n_n5169) & (x33x) & (x13296x)) + ((!n_n5162) & (n_n5168) & (n_n5169) & (!x33x) & (!x13296x)) + ((!n_n5162) & (n_n5168) & (n_n5169) & (!x33x) & (x13296x)) + ((!n_n5162) & (n_n5168) & (n_n5169) & (x33x) & (!x13296x)) + ((!n_n5162) & (n_n5168) & (n_n5169) & (x33x) & (x13296x)) + ((n_n5162) & (!n_n5168) & (!n_n5169) & (!x33x) & (!x13296x)) + ((n_n5162) & (!n_n5168) & (!n_n5169) & (!x33x) & (x13296x)) + ((n_n5162) & (!n_n5168) & (!n_n5169) & (x33x) & (!x13296x)) + ((n_n5162) & (!n_n5168) & (!n_n5169) & (x33x) & (x13296x)) + ((n_n5162) & (!n_n5168) & (n_n5169) & (!x33x) & (!x13296x)) + ((n_n5162) & (!n_n5168) & (n_n5169) & (!x33x) & (x13296x)) + ((n_n5162) & (!n_n5168) & (n_n5169) & (x33x) & (!x13296x)) + ((n_n5162) & (!n_n5168) & (n_n5169) & (x33x) & (x13296x)) + ((n_n5162) & (n_n5168) & (!n_n5169) & (!x33x) & (!x13296x)) + ((n_n5162) & (n_n5168) & (!n_n5169) & (!x33x) & (x13296x)) + ((n_n5162) & (n_n5168) & (!n_n5169) & (x33x) & (!x13296x)) + ((n_n5162) & (n_n5168) & (!n_n5169) & (x33x) & (x13296x)) + ((n_n5162) & (n_n5168) & (n_n5169) & (!x33x) & (!x13296x)) + ((n_n5162) & (n_n5168) & (n_n5169) & (!x33x) & (x13296x)) + ((n_n5162) & (n_n5168) & (n_n5169) & (x33x) & (!x13296x)) + ((n_n5162) & (n_n5168) & (n_n5169) & (x33x) & (x13296x)));
	assign x325x = (((!i_9_) & (!n_n473) & (!n_n534) & (!n_n65) & (n_n5306)) + ((!i_9_) & (!n_n473) & (!n_n534) & (n_n65) & (n_n5306)) + ((!i_9_) & (!n_n473) & (n_n534) & (!n_n65) & (n_n5306)) + ((!i_9_) & (!n_n473) & (n_n534) & (n_n65) & (n_n5306)) + ((!i_9_) & (n_n473) & (!n_n534) & (!n_n65) & (n_n5306)) + ((!i_9_) & (n_n473) & (!n_n534) & (n_n65) & (n_n5306)) + ((!i_9_) & (n_n473) & (n_n534) & (!n_n65) & (n_n5306)) + ((!i_9_) & (n_n473) & (n_n534) & (n_n65) & (!n_n5306)) + ((!i_9_) & (n_n473) & (n_n534) & (n_n65) & (n_n5306)) + ((i_9_) & (!n_n473) & (!n_n534) & (!n_n65) & (n_n5306)) + ((i_9_) & (!n_n473) & (!n_n534) & (n_n65) & (n_n5306)) + ((i_9_) & (!n_n473) & (n_n534) & (!n_n65) & (n_n5306)) + ((i_9_) & (!n_n473) & (n_n534) & (n_n65) & (n_n5306)) + ((i_9_) & (n_n473) & (!n_n534) & (!n_n65) & (n_n5306)) + ((i_9_) & (n_n473) & (!n_n534) & (n_n65) & (n_n5306)) + ((i_9_) & (n_n473) & (n_n534) & (!n_n65) & (n_n5306)) + ((i_9_) & (n_n473) & (n_n534) & (n_n65) & (n_n5306)));
	assign n_n4026 = (((!n_n5303) & (!n_n1128) & (!x63x) & (!x325x) & (n_n5304)) + ((!n_n5303) & (!n_n1128) & (!x63x) & (x325x) & (!n_n5304)) + ((!n_n5303) & (!n_n1128) & (!x63x) & (x325x) & (n_n5304)) + ((!n_n5303) & (!n_n1128) & (x63x) & (!x325x) & (!n_n5304)) + ((!n_n5303) & (!n_n1128) & (x63x) & (!x325x) & (n_n5304)) + ((!n_n5303) & (!n_n1128) & (x63x) & (x325x) & (!n_n5304)) + ((!n_n5303) & (!n_n1128) & (x63x) & (x325x) & (n_n5304)) + ((!n_n5303) & (n_n1128) & (!x63x) & (!x325x) & (!n_n5304)) + ((!n_n5303) & (n_n1128) & (!x63x) & (!x325x) & (n_n5304)) + ((!n_n5303) & (n_n1128) & (!x63x) & (x325x) & (!n_n5304)) + ((!n_n5303) & (n_n1128) & (!x63x) & (x325x) & (n_n5304)) + ((!n_n5303) & (n_n1128) & (x63x) & (!x325x) & (!n_n5304)) + ((!n_n5303) & (n_n1128) & (x63x) & (!x325x) & (n_n5304)) + ((!n_n5303) & (n_n1128) & (x63x) & (x325x) & (!n_n5304)) + ((!n_n5303) & (n_n1128) & (x63x) & (x325x) & (n_n5304)) + ((n_n5303) & (!n_n1128) & (!x63x) & (!x325x) & (!n_n5304)) + ((n_n5303) & (!n_n1128) & (!x63x) & (!x325x) & (n_n5304)) + ((n_n5303) & (!n_n1128) & (!x63x) & (x325x) & (!n_n5304)) + ((n_n5303) & (!n_n1128) & (!x63x) & (x325x) & (n_n5304)) + ((n_n5303) & (!n_n1128) & (x63x) & (!x325x) & (!n_n5304)) + ((n_n5303) & (!n_n1128) & (x63x) & (!x325x) & (n_n5304)) + ((n_n5303) & (!n_n1128) & (x63x) & (x325x) & (!n_n5304)) + ((n_n5303) & (!n_n1128) & (x63x) & (x325x) & (n_n5304)) + ((n_n5303) & (n_n1128) & (!x63x) & (!x325x) & (!n_n5304)) + ((n_n5303) & (n_n1128) & (!x63x) & (!x325x) & (n_n5304)) + ((n_n5303) & (n_n1128) & (!x63x) & (x325x) & (!n_n5304)) + ((n_n5303) & (n_n1128) & (!x63x) & (x325x) & (n_n5304)) + ((n_n5303) & (n_n1128) & (x63x) & (!x325x) & (!n_n5304)) + ((n_n5303) & (n_n1128) & (x63x) & (!x325x) & (n_n5304)) + ((n_n5303) & (n_n1128) & (x63x) & (x325x) & (!n_n5304)) + ((n_n5303) & (n_n1128) & (x63x) & (x325x) & (n_n5304)));
	assign x217x = (((!i_9_) & (!n_n528) & (!n_n491) & (!n_n65) & (n_n5280)) + ((!i_9_) & (!n_n528) & (!n_n491) & (n_n65) & (n_n5280)) + ((!i_9_) & (!n_n528) & (n_n491) & (!n_n65) & (n_n5280)) + ((!i_9_) & (!n_n528) & (n_n491) & (n_n65) & (n_n5280)) + ((!i_9_) & (n_n528) & (!n_n491) & (!n_n65) & (n_n5280)) + ((!i_9_) & (n_n528) & (!n_n491) & (n_n65) & (n_n5280)) + ((!i_9_) & (n_n528) & (n_n491) & (!n_n65) & (n_n5280)) + ((!i_9_) & (n_n528) & (n_n491) & (n_n65) & (!n_n5280)) + ((!i_9_) & (n_n528) & (n_n491) & (n_n65) & (n_n5280)) + ((i_9_) & (!n_n528) & (!n_n491) & (!n_n65) & (n_n5280)) + ((i_9_) & (!n_n528) & (!n_n491) & (n_n65) & (n_n5280)) + ((i_9_) & (!n_n528) & (n_n491) & (!n_n65) & (n_n5280)) + ((i_9_) & (!n_n528) & (n_n491) & (n_n65) & (n_n5280)) + ((i_9_) & (n_n528) & (!n_n491) & (!n_n65) & (n_n5280)) + ((i_9_) & (n_n528) & (!n_n491) & (n_n65) & (n_n5280)) + ((i_9_) & (n_n528) & (n_n491) & (!n_n65) & (n_n5280)) + ((i_9_) & (n_n528) & (n_n491) & (n_n65) & (n_n5280)));
	assign x333x = (((!i_9_) & (!x19x) & (n_n532) & (n_n491) & (n_n65)) + ((!i_9_) & (x19x) & (n_n532) & (n_n491) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n532) & (n_n491) & (n_n65)) + ((i_9_) & (x19x) & (n_n532) & (n_n491) & (!n_n65)) + ((i_9_) & (x19x) & (n_n532) & (n_n491) & (n_n65)));
	assign x13332x = (((!x15x) & (!x21x) & (!n_n491) & (!n_n65) & (n_n5282)) + ((!x15x) & (!x21x) & (!n_n491) & (n_n65) & (n_n5282)) + ((!x15x) & (!x21x) & (n_n491) & (!n_n65) & (n_n5282)) + ((!x15x) & (!x21x) & (n_n491) & (n_n65) & (n_n5282)) + ((!x15x) & (x21x) & (!n_n491) & (!n_n65) & (n_n5282)) + ((!x15x) & (x21x) & (!n_n491) & (n_n65) & (n_n5282)) + ((!x15x) & (x21x) & (n_n491) & (!n_n65) & (n_n5282)) + ((!x15x) & (x21x) & (n_n491) & (n_n65) & (!n_n5282)) + ((!x15x) & (x21x) & (n_n491) & (n_n65) & (n_n5282)) + ((x15x) & (!x21x) & (!n_n491) & (!n_n65) & (n_n5282)) + ((x15x) & (!x21x) & (!n_n491) & (n_n65) & (n_n5282)) + ((x15x) & (!x21x) & (n_n491) & (!n_n65) & (n_n5282)) + ((x15x) & (!x21x) & (n_n491) & (n_n65) & (!n_n5282)) + ((x15x) & (!x21x) & (n_n491) & (n_n65) & (n_n5282)) + ((x15x) & (x21x) & (!n_n491) & (!n_n65) & (n_n5282)) + ((x15x) & (x21x) & (!n_n491) & (n_n65) & (n_n5282)) + ((x15x) & (x21x) & (n_n491) & (!n_n65) & (n_n5282)) + ((x15x) & (x21x) & (n_n491) & (n_n65) & (!n_n5282)) + ((x15x) & (x21x) & (n_n491) & (n_n65) & (n_n5282)));
	assign n_n4028 = (((!n_n5276) & (!n_n5281) & (!x217x) & (!x333x) & (x13332x)) + ((!n_n5276) & (!n_n5281) & (!x217x) & (x333x) & (!x13332x)) + ((!n_n5276) & (!n_n5281) & (!x217x) & (x333x) & (x13332x)) + ((!n_n5276) & (!n_n5281) & (x217x) & (!x333x) & (!x13332x)) + ((!n_n5276) & (!n_n5281) & (x217x) & (!x333x) & (x13332x)) + ((!n_n5276) & (!n_n5281) & (x217x) & (x333x) & (!x13332x)) + ((!n_n5276) & (!n_n5281) & (x217x) & (x333x) & (x13332x)) + ((!n_n5276) & (n_n5281) & (!x217x) & (!x333x) & (!x13332x)) + ((!n_n5276) & (n_n5281) & (!x217x) & (!x333x) & (x13332x)) + ((!n_n5276) & (n_n5281) & (!x217x) & (x333x) & (!x13332x)) + ((!n_n5276) & (n_n5281) & (!x217x) & (x333x) & (x13332x)) + ((!n_n5276) & (n_n5281) & (x217x) & (!x333x) & (!x13332x)) + ((!n_n5276) & (n_n5281) & (x217x) & (!x333x) & (x13332x)) + ((!n_n5276) & (n_n5281) & (x217x) & (x333x) & (!x13332x)) + ((!n_n5276) & (n_n5281) & (x217x) & (x333x) & (x13332x)) + ((n_n5276) & (!n_n5281) & (!x217x) & (!x333x) & (!x13332x)) + ((n_n5276) & (!n_n5281) & (!x217x) & (!x333x) & (x13332x)) + ((n_n5276) & (!n_n5281) & (!x217x) & (x333x) & (!x13332x)) + ((n_n5276) & (!n_n5281) & (!x217x) & (x333x) & (x13332x)) + ((n_n5276) & (!n_n5281) & (x217x) & (!x333x) & (!x13332x)) + ((n_n5276) & (!n_n5281) & (x217x) & (!x333x) & (x13332x)) + ((n_n5276) & (!n_n5281) & (x217x) & (x333x) & (!x13332x)) + ((n_n5276) & (!n_n5281) & (x217x) & (x333x) & (x13332x)) + ((n_n5276) & (n_n5281) & (!x217x) & (!x333x) & (!x13332x)) + ((n_n5276) & (n_n5281) & (!x217x) & (!x333x) & (x13332x)) + ((n_n5276) & (n_n5281) & (!x217x) & (x333x) & (!x13332x)) + ((n_n5276) & (n_n5281) & (!x217x) & (x333x) & (x13332x)) + ((n_n5276) & (n_n5281) & (x217x) & (!x333x) & (!x13332x)) + ((n_n5276) & (n_n5281) & (x217x) & (!x333x) & (x13332x)) + ((n_n5276) & (n_n5281) & (x217x) & (x333x) & (!x13332x)) + ((n_n5276) & (n_n5281) & (x217x) & (x333x) & (x13332x)));
	assign x77x = (((!x19x) & (!n_n522) & (x20x) & (n_n500) & (n_n65)) + ((!x19x) & (n_n522) & (x20x) & (n_n500) & (n_n65)) + ((x19x) & (!n_n522) & (x20x) & (n_n500) & (n_n65)) + ((x19x) & (n_n522) & (!x20x) & (n_n500) & (!n_n65)) + ((x19x) & (n_n522) & (!x20x) & (n_n500) & (n_n65)) + ((x19x) & (n_n522) & (x20x) & (n_n500) & (!n_n65)) + ((x19x) & (n_n522) & (x20x) & (n_n500) & (n_n65)));
	assign x205x = (((!i_9_) & (!x19x) & (n_n526) & (n_n500) & (n_n65)) + ((!i_9_) & (x19x) & (n_n526) & (n_n500) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n526) & (n_n500) & (n_n65)) + ((i_9_) & (x19x) & (n_n526) & (n_n500) & (!n_n65)) + ((i_9_) & (x19x) & (n_n526) & (n_n500) & (n_n65)));
	assign x22187x = (((!x19x) & (!n_n524) & (!n_n520) & (!n_n500) & (!n_n5271)) + ((!x19x) & (!n_n524) & (!n_n520) & (n_n500) & (!n_n5271)) + ((!x19x) & (!n_n524) & (n_n520) & (!n_n500) & (!n_n5271)) + ((!x19x) & (!n_n524) & (n_n520) & (n_n500) & (!n_n5271)) + ((!x19x) & (n_n524) & (!n_n520) & (!n_n500) & (!n_n5271)) + ((!x19x) & (n_n524) & (!n_n520) & (n_n500) & (!n_n5271)) + ((!x19x) & (n_n524) & (n_n520) & (!n_n500) & (!n_n5271)) + ((!x19x) & (n_n524) & (n_n520) & (n_n500) & (!n_n5271)) + ((x19x) & (!n_n524) & (!n_n520) & (!n_n500) & (!n_n5271)) + ((x19x) & (!n_n524) & (!n_n520) & (n_n500) & (!n_n5271)) + ((x19x) & (!n_n524) & (n_n520) & (!n_n500) & (!n_n5271)) + ((x19x) & (n_n524) & (!n_n520) & (!n_n500) & (!n_n5271)) + ((x19x) & (n_n524) & (n_n520) & (!n_n500) & (!n_n5271)));
	assign x13348x = (((!n_n5273) & (!n_n5272) & (!x77x) & (!x205x) & (!x22187x)) + ((!n_n5273) & (!n_n5272) & (!x77x) & (x205x) & (!x22187x)) + ((!n_n5273) & (!n_n5272) & (!x77x) & (x205x) & (x22187x)) + ((!n_n5273) & (!n_n5272) & (x77x) & (!x205x) & (!x22187x)) + ((!n_n5273) & (!n_n5272) & (x77x) & (!x205x) & (x22187x)) + ((!n_n5273) & (!n_n5272) & (x77x) & (x205x) & (!x22187x)) + ((!n_n5273) & (!n_n5272) & (x77x) & (x205x) & (x22187x)) + ((!n_n5273) & (n_n5272) & (!x77x) & (!x205x) & (!x22187x)) + ((!n_n5273) & (n_n5272) & (!x77x) & (!x205x) & (x22187x)) + ((!n_n5273) & (n_n5272) & (!x77x) & (x205x) & (!x22187x)) + ((!n_n5273) & (n_n5272) & (!x77x) & (x205x) & (x22187x)) + ((!n_n5273) & (n_n5272) & (x77x) & (!x205x) & (!x22187x)) + ((!n_n5273) & (n_n5272) & (x77x) & (!x205x) & (x22187x)) + ((!n_n5273) & (n_n5272) & (x77x) & (x205x) & (!x22187x)) + ((!n_n5273) & (n_n5272) & (x77x) & (x205x) & (x22187x)) + ((n_n5273) & (!n_n5272) & (!x77x) & (!x205x) & (!x22187x)) + ((n_n5273) & (!n_n5272) & (!x77x) & (!x205x) & (x22187x)) + ((n_n5273) & (!n_n5272) & (!x77x) & (x205x) & (!x22187x)) + ((n_n5273) & (!n_n5272) & (!x77x) & (x205x) & (x22187x)) + ((n_n5273) & (!n_n5272) & (x77x) & (!x205x) & (!x22187x)) + ((n_n5273) & (!n_n5272) & (x77x) & (!x205x) & (x22187x)) + ((n_n5273) & (!n_n5272) & (x77x) & (x205x) & (!x22187x)) + ((n_n5273) & (!n_n5272) & (x77x) & (x205x) & (x22187x)) + ((n_n5273) & (n_n5272) & (!x77x) & (!x205x) & (!x22187x)) + ((n_n5273) & (n_n5272) & (!x77x) & (!x205x) & (x22187x)) + ((n_n5273) & (n_n5272) & (!x77x) & (x205x) & (!x22187x)) + ((n_n5273) & (n_n5272) & (!x77x) & (x205x) & (x22187x)) + ((n_n5273) & (n_n5272) & (x77x) & (!x205x) & (!x22187x)) + ((n_n5273) & (n_n5272) & (x77x) & (!x205x) & (x22187x)) + ((n_n5273) & (n_n5272) & (x77x) & (x205x) & (!x22187x)) + ((n_n5273) & (n_n5272) & (x77x) & (x205x) & (x22187x)));
	assign x13338x = (((!n_n5258) & (!n_n5251) & (!n_n5254) & (n_n5253)) + ((!n_n5258) & (!n_n5251) & (n_n5254) & (!n_n5253)) + ((!n_n5258) & (!n_n5251) & (n_n5254) & (n_n5253)) + ((!n_n5258) & (n_n5251) & (!n_n5254) & (!n_n5253)) + ((!n_n5258) & (n_n5251) & (!n_n5254) & (n_n5253)) + ((!n_n5258) & (n_n5251) & (n_n5254) & (!n_n5253)) + ((!n_n5258) & (n_n5251) & (n_n5254) & (n_n5253)) + ((n_n5258) & (!n_n5251) & (!n_n5254) & (!n_n5253)) + ((n_n5258) & (!n_n5251) & (!n_n5254) & (n_n5253)) + ((n_n5258) & (!n_n5251) & (n_n5254) & (!n_n5253)) + ((n_n5258) & (!n_n5251) & (n_n5254) & (n_n5253)) + ((n_n5258) & (n_n5251) & (!n_n5254) & (!n_n5253)) + ((n_n5258) & (n_n5251) & (!n_n5254) & (n_n5253)) + ((n_n5258) & (n_n5251) & (n_n5254) & (!n_n5253)) + ((n_n5258) & (n_n5251) & (n_n5254) & (n_n5253)));
	assign x13339x = (((!n_n5262) & (!n_n5252) & (!n_n5261) & (!n_n5256) & (n_n5259)) + ((!n_n5262) & (!n_n5252) & (!n_n5261) & (n_n5256) & (!n_n5259)) + ((!n_n5262) & (!n_n5252) & (!n_n5261) & (n_n5256) & (n_n5259)) + ((!n_n5262) & (!n_n5252) & (n_n5261) & (!n_n5256) & (!n_n5259)) + ((!n_n5262) & (!n_n5252) & (n_n5261) & (!n_n5256) & (n_n5259)) + ((!n_n5262) & (!n_n5252) & (n_n5261) & (n_n5256) & (!n_n5259)) + ((!n_n5262) & (!n_n5252) & (n_n5261) & (n_n5256) & (n_n5259)) + ((!n_n5262) & (n_n5252) & (!n_n5261) & (!n_n5256) & (!n_n5259)) + ((!n_n5262) & (n_n5252) & (!n_n5261) & (!n_n5256) & (n_n5259)) + ((!n_n5262) & (n_n5252) & (!n_n5261) & (n_n5256) & (!n_n5259)) + ((!n_n5262) & (n_n5252) & (!n_n5261) & (n_n5256) & (n_n5259)) + ((!n_n5262) & (n_n5252) & (n_n5261) & (!n_n5256) & (!n_n5259)) + ((!n_n5262) & (n_n5252) & (n_n5261) & (!n_n5256) & (n_n5259)) + ((!n_n5262) & (n_n5252) & (n_n5261) & (n_n5256) & (!n_n5259)) + ((!n_n5262) & (n_n5252) & (n_n5261) & (n_n5256) & (n_n5259)) + ((n_n5262) & (!n_n5252) & (!n_n5261) & (!n_n5256) & (!n_n5259)) + ((n_n5262) & (!n_n5252) & (!n_n5261) & (!n_n5256) & (n_n5259)) + ((n_n5262) & (!n_n5252) & (!n_n5261) & (n_n5256) & (!n_n5259)) + ((n_n5262) & (!n_n5252) & (!n_n5261) & (n_n5256) & (n_n5259)) + ((n_n5262) & (!n_n5252) & (n_n5261) & (!n_n5256) & (!n_n5259)) + ((n_n5262) & (!n_n5252) & (n_n5261) & (!n_n5256) & (n_n5259)) + ((n_n5262) & (!n_n5252) & (n_n5261) & (n_n5256) & (!n_n5259)) + ((n_n5262) & (!n_n5252) & (n_n5261) & (n_n5256) & (n_n5259)) + ((n_n5262) & (n_n5252) & (!n_n5261) & (!n_n5256) & (!n_n5259)) + ((n_n5262) & (n_n5252) & (!n_n5261) & (!n_n5256) & (n_n5259)) + ((n_n5262) & (n_n5252) & (!n_n5261) & (n_n5256) & (!n_n5259)) + ((n_n5262) & (n_n5252) & (!n_n5261) & (n_n5256) & (n_n5259)) + ((n_n5262) & (n_n5252) & (n_n5261) & (!n_n5256) & (!n_n5259)) + ((n_n5262) & (n_n5252) & (n_n5261) & (!n_n5256) & (n_n5259)) + ((n_n5262) & (n_n5252) & (n_n5261) & (n_n5256) & (!n_n5259)) + ((n_n5262) & (n_n5252) & (n_n5261) & (n_n5256) & (n_n5259)));
	assign n_n4031 = (((!n_n5244) & (!n_n5247) & (!n_n5246) & (!n_n5243) & (x13343x)) + ((!n_n5244) & (!n_n5247) & (!n_n5246) & (n_n5243) & (!x13343x)) + ((!n_n5244) & (!n_n5247) & (!n_n5246) & (n_n5243) & (x13343x)) + ((!n_n5244) & (!n_n5247) & (n_n5246) & (!n_n5243) & (!x13343x)) + ((!n_n5244) & (!n_n5247) & (n_n5246) & (!n_n5243) & (x13343x)) + ((!n_n5244) & (!n_n5247) & (n_n5246) & (n_n5243) & (!x13343x)) + ((!n_n5244) & (!n_n5247) & (n_n5246) & (n_n5243) & (x13343x)) + ((!n_n5244) & (n_n5247) & (!n_n5246) & (!n_n5243) & (!x13343x)) + ((!n_n5244) & (n_n5247) & (!n_n5246) & (!n_n5243) & (x13343x)) + ((!n_n5244) & (n_n5247) & (!n_n5246) & (n_n5243) & (!x13343x)) + ((!n_n5244) & (n_n5247) & (!n_n5246) & (n_n5243) & (x13343x)) + ((!n_n5244) & (n_n5247) & (n_n5246) & (!n_n5243) & (!x13343x)) + ((!n_n5244) & (n_n5247) & (n_n5246) & (!n_n5243) & (x13343x)) + ((!n_n5244) & (n_n5247) & (n_n5246) & (n_n5243) & (!x13343x)) + ((!n_n5244) & (n_n5247) & (n_n5246) & (n_n5243) & (x13343x)) + ((n_n5244) & (!n_n5247) & (!n_n5246) & (!n_n5243) & (!x13343x)) + ((n_n5244) & (!n_n5247) & (!n_n5246) & (!n_n5243) & (x13343x)) + ((n_n5244) & (!n_n5247) & (!n_n5246) & (n_n5243) & (!x13343x)) + ((n_n5244) & (!n_n5247) & (!n_n5246) & (n_n5243) & (x13343x)) + ((n_n5244) & (!n_n5247) & (n_n5246) & (!n_n5243) & (!x13343x)) + ((n_n5244) & (!n_n5247) & (n_n5246) & (!n_n5243) & (x13343x)) + ((n_n5244) & (!n_n5247) & (n_n5246) & (n_n5243) & (!x13343x)) + ((n_n5244) & (!n_n5247) & (n_n5246) & (n_n5243) & (x13343x)) + ((n_n5244) & (n_n5247) & (!n_n5246) & (!n_n5243) & (!x13343x)) + ((n_n5244) & (n_n5247) & (!n_n5246) & (!n_n5243) & (x13343x)) + ((n_n5244) & (n_n5247) & (!n_n5246) & (n_n5243) & (!x13343x)) + ((n_n5244) & (n_n5247) & (!n_n5246) & (n_n5243) & (x13343x)) + ((n_n5244) & (n_n5247) & (n_n5246) & (!n_n5243) & (!x13343x)) + ((n_n5244) & (n_n5247) & (n_n5246) & (!n_n5243) & (x13343x)) + ((n_n5244) & (n_n5247) & (n_n5246) & (n_n5243) & (!x13343x)) + ((n_n5244) & (n_n5247) & (n_n5246) & (n_n5243) & (x13343x)));
	assign n_n3998 = (((!x13348x) & (!x13338x) & (!x13339x) & (n_n4031)) + ((!x13348x) & (!x13338x) & (x13339x) & (!n_n4031)) + ((!x13348x) & (!x13338x) & (x13339x) & (n_n4031)) + ((!x13348x) & (x13338x) & (!x13339x) & (!n_n4031)) + ((!x13348x) & (x13338x) & (!x13339x) & (n_n4031)) + ((!x13348x) & (x13338x) & (x13339x) & (!n_n4031)) + ((!x13348x) & (x13338x) & (x13339x) & (n_n4031)) + ((x13348x) & (!x13338x) & (!x13339x) & (!n_n4031)) + ((x13348x) & (!x13338x) & (!x13339x) & (n_n4031)) + ((x13348x) & (!x13338x) & (x13339x) & (!n_n4031)) + ((x13348x) & (!x13338x) & (x13339x) & (n_n4031)) + ((x13348x) & (x13338x) & (!x13339x) & (!n_n4031)) + ((x13348x) & (x13338x) & (!x13339x) & (n_n4031)) + ((x13348x) & (x13338x) & (x13339x) & (!n_n4031)) + ((x13348x) & (x13338x) & (x13339x) & (n_n4031)));
	assign n_n1530 = (((!i_9_) & (!n_n518) & (!n_n534) & (!n_n65) & (n_n5226)) + ((!i_9_) & (!n_n518) & (!n_n534) & (n_n65) & (n_n5226)) + ((!i_9_) & (!n_n518) & (n_n534) & (!n_n65) & (n_n5226)) + ((!i_9_) & (!n_n518) & (n_n534) & (n_n65) & (n_n5226)) + ((!i_9_) & (n_n518) & (!n_n534) & (!n_n65) & (n_n5226)) + ((!i_9_) & (n_n518) & (!n_n534) & (n_n65) & (n_n5226)) + ((!i_9_) & (n_n518) & (n_n534) & (!n_n65) & (n_n5226)) + ((!i_9_) & (n_n518) & (n_n534) & (n_n65) & (!n_n5226)) + ((!i_9_) & (n_n518) & (n_n534) & (n_n65) & (n_n5226)) + ((i_9_) & (!n_n518) & (!n_n534) & (!n_n65) & (n_n5226)) + ((i_9_) & (!n_n518) & (!n_n534) & (n_n65) & (n_n5226)) + ((i_9_) & (!n_n518) & (n_n534) & (!n_n65) & (n_n5226)) + ((i_9_) & (!n_n518) & (n_n534) & (n_n65) & (n_n5226)) + ((i_9_) & (n_n518) & (!n_n534) & (!n_n65) & (n_n5226)) + ((i_9_) & (n_n518) & (!n_n534) & (n_n65) & (n_n5226)) + ((i_9_) & (n_n518) & (n_n534) & (!n_n65) & (n_n5226)) + ((i_9_) & (n_n518) & (n_n534) & (n_n65) & (!n_n5226)) + ((i_9_) & (n_n518) & (n_n534) & (n_n65) & (n_n5226)));
	assign n_n2290 = (((!i_9_) & (!n_n528) & (!n_n535) & (!n_n65) & (n_n5218)) + ((!i_9_) & (!n_n528) & (!n_n535) & (n_n65) & (n_n5218)) + ((!i_9_) & (!n_n528) & (n_n535) & (!n_n65) & (n_n5218)) + ((!i_9_) & (!n_n528) & (n_n535) & (n_n65) & (n_n5218)) + ((!i_9_) & (n_n528) & (!n_n535) & (!n_n65) & (n_n5218)) + ((!i_9_) & (n_n528) & (!n_n535) & (n_n65) & (n_n5218)) + ((!i_9_) & (n_n528) & (n_n535) & (!n_n65) & (n_n5218)) + ((!i_9_) & (n_n528) & (n_n535) & (n_n65) & (!n_n5218)) + ((!i_9_) & (n_n528) & (n_n535) & (n_n65) & (n_n5218)) + ((i_9_) & (!n_n528) & (!n_n535) & (!n_n65) & (n_n5218)) + ((i_9_) & (!n_n528) & (!n_n535) & (n_n65) & (n_n5218)) + ((i_9_) & (!n_n528) & (n_n535) & (!n_n65) & (n_n5218)) + ((i_9_) & (!n_n528) & (n_n535) & (n_n65) & (n_n5218)) + ((i_9_) & (n_n528) & (!n_n535) & (!n_n65) & (n_n5218)) + ((i_9_) & (n_n528) & (!n_n535) & (n_n65) & (n_n5218)) + ((i_9_) & (n_n528) & (n_n535) & (!n_n65) & (n_n5218)) + ((i_9_) & (n_n528) & (n_n535) & (n_n65) & (!n_n5218)) + ((i_9_) & (n_n528) & (n_n535) & (n_n65) & (n_n5218)));
	assign n_n4032 = (((!n_n5237) & (!n_n5235) & (!x181x) & (!x13351x) & (x13353x)) + ((!n_n5237) & (!n_n5235) & (!x181x) & (x13351x) & (!x13353x)) + ((!n_n5237) & (!n_n5235) & (!x181x) & (x13351x) & (x13353x)) + ((!n_n5237) & (!n_n5235) & (x181x) & (!x13351x) & (!x13353x)) + ((!n_n5237) & (!n_n5235) & (x181x) & (!x13351x) & (x13353x)) + ((!n_n5237) & (!n_n5235) & (x181x) & (x13351x) & (!x13353x)) + ((!n_n5237) & (!n_n5235) & (x181x) & (x13351x) & (x13353x)) + ((!n_n5237) & (n_n5235) & (!x181x) & (!x13351x) & (!x13353x)) + ((!n_n5237) & (n_n5235) & (!x181x) & (!x13351x) & (x13353x)) + ((!n_n5237) & (n_n5235) & (!x181x) & (x13351x) & (!x13353x)) + ((!n_n5237) & (n_n5235) & (!x181x) & (x13351x) & (x13353x)) + ((!n_n5237) & (n_n5235) & (x181x) & (!x13351x) & (!x13353x)) + ((!n_n5237) & (n_n5235) & (x181x) & (!x13351x) & (x13353x)) + ((!n_n5237) & (n_n5235) & (x181x) & (x13351x) & (!x13353x)) + ((!n_n5237) & (n_n5235) & (x181x) & (x13351x) & (x13353x)) + ((n_n5237) & (!n_n5235) & (!x181x) & (!x13351x) & (!x13353x)) + ((n_n5237) & (!n_n5235) & (!x181x) & (!x13351x) & (x13353x)) + ((n_n5237) & (!n_n5235) & (!x181x) & (x13351x) & (!x13353x)) + ((n_n5237) & (!n_n5235) & (!x181x) & (x13351x) & (x13353x)) + ((n_n5237) & (!n_n5235) & (x181x) & (!x13351x) & (!x13353x)) + ((n_n5237) & (!n_n5235) & (x181x) & (!x13351x) & (x13353x)) + ((n_n5237) & (!n_n5235) & (x181x) & (x13351x) & (!x13353x)) + ((n_n5237) & (!n_n5235) & (x181x) & (x13351x) & (x13353x)) + ((n_n5237) & (n_n5235) & (!x181x) & (!x13351x) & (!x13353x)) + ((n_n5237) & (n_n5235) & (!x181x) & (!x13351x) & (x13353x)) + ((n_n5237) & (n_n5235) & (!x181x) & (x13351x) & (!x13353x)) + ((n_n5237) & (n_n5235) & (!x181x) & (x13351x) & (x13353x)) + ((n_n5237) & (n_n5235) & (x181x) & (!x13351x) & (!x13353x)) + ((n_n5237) & (n_n5235) & (x181x) & (!x13351x) & (x13353x)) + ((n_n5237) & (n_n5235) & (x181x) & (x13351x) & (!x13353x)) + ((n_n5237) & (n_n5235) & (x181x) & (x13351x) & (x13353x)));
	assign x13361x = (((!n_n5220) & (!n_n5203) & (!n_n5205) & (n_n5211)) + ((!n_n5220) & (!n_n5203) & (n_n5205) & (!n_n5211)) + ((!n_n5220) & (!n_n5203) & (n_n5205) & (n_n5211)) + ((!n_n5220) & (n_n5203) & (!n_n5205) & (!n_n5211)) + ((!n_n5220) & (n_n5203) & (!n_n5205) & (n_n5211)) + ((!n_n5220) & (n_n5203) & (n_n5205) & (!n_n5211)) + ((!n_n5220) & (n_n5203) & (n_n5205) & (n_n5211)) + ((n_n5220) & (!n_n5203) & (!n_n5205) & (!n_n5211)) + ((n_n5220) & (!n_n5203) & (!n_n5205) & (n_n5211)) + ((n_n5220) & (!n_n5203) & (n_n5205) & (!n_n5211)) + ((n_n5220) & (!n_n5203) & (n_n5205) & (n_n5211)) + ((n_n5220) & (n_n5203) & (!n_n5205) & (!n_n5211)) + ((n_n5220) & (n_n5203) & (!n_n5205) & (n_n5211)) + ((n_n5220) & (n_n5203) & (n_n5205) & (!n_n5211)) + ((n_n5220) & (n_n5203) & (n_n5205) & (n_n5211)));
	assign x13363x = (((!n_n5204) & (!n_n5201) & (!x223x) & (!x384x) & (x450x)) + ((!n_n5204) & (!n_n5201) & (!x223x) & (x384x) & (!x450x)) + ((!n_n5204) & (!n_n5201) & (!x223x) & (x384x) & (x450x)) + ((!n_n5204) & (!n_n5201) & (x223x) & (!x384x) & (!x450x)) + ((!n_n5204) & (!n_n5201) & (x223x) & (!x384x) & (x450x)) + ((!n_n5204) & (!n_n5201) & (x223x) & (x384x) & (!x450x)) + ((!n_n5204) & (!n_n5201) & (x223x) & (x384x) & (x450x)) + ((!n_n5204) & (n_n5201) & (!x223x) & (!x384x) & (!x450x)) + ((!n_n5204) & (n_n5201) & (!x223x) & (!x384x) & (x450x)) + ((!n_n5204) & (n_n5201) & (!x223x) & (x384x) & (!x450x)) + ((!n_n5204) & (n_n5201) & (!x223x) & (x384x) & (x450x)) + ((!n_n5204) & (n_n5201) & (x223x) & (!x384x) & (!x450x)) + ((!n_n5204) & (n_n5201) & (x223x) & (!x384x) & (x450x)) + ((!n_n5204) & (n_n5201) & (x223x) & (x384x) & (!x450x)) + ((!n_n5204) & (n_n5201) & (x223x) & (x384x) & (x450x)) + ((n_n5204) & (!n_n5201) & (!x223x) & (!x384x) & (!x450x)) + ((n_n5204) & (!n_n5201) & (!x223x) & (!x384x) & (x450x)) + ((n_n5204) & (!n_n5201) & (!x223x) & (x384x) & (!x450x)) + ((n_n5204) & (!n_n5201) & (!x223x) & (x384x) & (x450x)) + ((n_n5204) & (!n_n5201) & (x223x) & (!x384x) & (!x450x)) + ((n_n5204) & (!n_n5201) & (x223x) & (!x384x) & (x450x)) + ((n_n5204) & (!n_n5201) & (x223x) & (x384x) & (!x450x)) + ((n_n5204) & (!n_n5201) & (x223x) & (x384x) & (x450x)) + ((n_n5204) & (n_n5201) & (!x223x) & (!x384x) & (!x450x)) + ((n_n5204) & (n_n5201) & (!x223x) & (!x384x) & (x450x)) + ((n_n5204) & (n_n5201) & (!x223x) & (x384x) & (!x450x)) + ((n_n5204) & (n_n5201) & (!x223x) & (x384x) & (x450x)) + ((n_n5204) & (n_n5201) & (x223x) & (!x384x) & (!x450x)) + ((n_n5204) & (n_n5201) & (x223x) & (!x384x) & (x450x)) + ((n_n5204) & (n_n5201) & (x223x) & (x384x) & (!x450x)) + ((n_n5204) & (n_n5201) & (x223x) & (x384x) & (x450x)));
	assign n_n3999 = (((!n_n1530) & (!n_n2290) & (!n_n4032) & (!x13361x) & (x13363x)) + ((!n_n1530) & (!n_n2290) & (!n_n4032) & (x13361x) & (!x13363x)) + ((!n_n1530) & (!n_n2290) & (!n_n4032) & (x13361x) & (x13363x)) + ((!n_n1530) & (!n_n2290) & (n_n4032) & (!x13361x) & (!x13363x)) + ((!n_n1530) & (!n_n2290) & (n_n4032) & (!x13361x) & (x13363x)) + ((!n_n1530) & (!n_n2290) & (n_n4032) & (x13361x) & (!x13363x)) + ((!n_n1530) & (!n_n2290) & (n_n4032) & (x13361x) & (x13363x)) + ((!n_n1530) & (n_n2290) & (!n_n4032) & (!x13361x) & (!x13363x)) + ((!n_n1530) & (n_n2290) & (!n_n4032) & (!x13361x) & (x13363x)) + ((!n_n1530) & (n_n2290) & (!n_n4032) & (x13361x) & (!x13363x)) + ((!n_n1530) & (n_n2290) & (!n_n4032) & (x13361x) & (x13363x)) + ((!n_n1530) & (n_n2290) & (n_n4032) & (!x13361x) & (!x13363x)) + ((!n_n1530) & (n_n2290) & (n_n4032) & (!x13361x) & (x13363x)) + ((!n_n1530) & (n_n2290) & (n_n4032) & (x13361x) & (!x13363x)) + ((!n_n1530) & (n_n2290) & (n_n4032) & (x13361x) & (x13363x)) + ((n_n1530) & (!n_n2290) & (!n_n4032) & (!x13361x) & (!x13363x)) + ((n_n1530) & (!n_n2290) & (!n_n4032) & (!x13361x) & (x13363x)) + ((n_n1530) & (!n_n2290) & (!n_n4032) & (x13361x) & (!x13363x)) + ((n_n1530) & (!n_n2290) & (!n_n4032) & (x13361x) & (x13363x)) + ((n_n1530) & (!n_n2290) & (n_n4032) & (!x13361x) & (!x13363x)) + ((n_n1530) & (!n_n2290) & (n_n4032) & (!x13361x) & (x13363x)) + ((n_n1530) & (!n_n2290) & (n_n4032) & (x13361x) & (!x13363x)) + ((n_n1530) & (!n_n2290) & (n_n4032) & (x13361x) & (x13363x)) + ((n_n1530) & (n_n2290) & (!n_n4032) & (!x13361x) & (!x13363x)) + ((n_n1530) & (n_n2290) & (!n_n4032) & (!x13361x) & (x13363x)) + ((n_n1530) & (n_n2290) & (!n_n4032) & (x13361x) & (!x13363x)) + ((n_n1530) & (n_n2290) & (!n_n4032) & (x13361x) & (x13363x)) + ((n_n1530) & (n_n2290) & (n_n4032) & (!x13361x) & (!x13363x)) + ((n_n1530) & (n_n2290) & (n_n4032) & (!x13361x) & (x13363x)) + ((n_n1530) & (n_n2290) & (n_n4032) & (x13361x) & (!x13363x)) + ((n_n1530) & (n_n2290) & (n_n4032) & (x13361x) & (x13363x)));
	assign n_n5285 = (((i_5_) & (!i_3_) & (i_4_) & (x20x) & (n_n65)));
	assign x441x = (((!x19x) & (!n_n522) & (n_n491) & (x20x) & (n_n65)) + ((!x19x) & (n_n522) & (n_n491) & (x20x) & (n_n65)) + ((x19x) & (!n_n522) & (n_n491) & (x20x) & (n_n65)) + ((x19x) & (n_n522) & (n_n491) & (!x20x) & (!n_n65)) + ((x19x) & (n_n522) & (n_n491) & (!x20x) & (n_n65)) + ((x19x) & (n_n522) & (n_n491) & (x20x) & (!n_n65)) + ((x19x) & (n_n522) & (n_n491) & (x20x) & (n_n65)));
	assign x13370x = (((!x592x) & (!x21x) & (!n_n5294) & (!n_n5287) & (n_n5288)) + ((!x592x) & (!x21x) & (!n_n5294) & (n_n5287) & (!n_n5288)) + ((!x592x) & (!x21x) & (!n_n5294) & (n_n5287) & (n_n5288)) + ((!x592x) & (!x21x) & (n_n5294) & (!n_n5287) & (!n_n5288)) + ((!x592x) & (!x21x) & (n_n5294) & (!n_n5287) & (n_n5288)) + ((!x592x) & (!x21x) & (n_n5294) & (n_n5287) & (!n_n5288)) + ((!x592x) & (!x21x) & (n_n5294) & (n_n5287) & (n_n5288)) + ((!x592x) & (x21x) & (!n_n5294) & (!n_n5287) & (n_n5288)) + ((!x592x) & (x21x) & (!n_n5294) & (n_n5287) & (!n_n5288)) + ((!x592x) & (x21x) & (!n_n5294) & (n_n5287) & (n_n5288)) + ((!x592x) & (x21x) & (n_n5294) & (!n_n5287) & (!n_n5288)) + ((!x592x) & (x21x) & (n_n5294) & (!n_n5287) & (n_n5288)) + ((!x592x) & (x21x) & (n_n5294) & (n_n5287) & (!n_n5288)) + ((!x592x) & (x21x) & (n_n5294) & (n_n5287) & (n_n5288)) + ((x592x) & (!x21x) & (!n_n5294) & (!n_n5287) & (n_n5288)) + ((x592x) & (!x21x) & (!n_n5294) & (n_n5287) & (!n_n5288)) + ((x592x) & (!x21x) & (!n_n5294) & (n_n5287) & (n_n5288)) + ((x592x) & (!x21x) & (n_n5294) & (!n_n5287) & (!n_n5288)) + ((x592x) & (!x21x) & (n_n5294) & (!n_n5287) & (n_n5288)) + ((x592x) & (!x21x) & (n_n5294) & (n_n5287) & (!n_n5288)) + ((x592x) & (!x21x) & (n_n5294) & (n_n5287) & (n_n5288)) + ((x592x) & (x21x) & (!n_n5294) & (!n_n5287) & (!n_n5288)) + ((x592x) & (x21x) & (!n_n5294) & (!n_n5287) & (n_n5288)) + ((x592x) & (x21x) & (!n_n5294) & (n_n5287) & (!n_n5288)) + ((x592x) & (x21x) & (!n_n5294) & (n_n5287) & (n_n5288)) + ((x592x) & (x21x) & (n_n5294) & (!n_n5287) & (!n_n5288)) + ((x592x) & (x21x) & (n_n5294) & (!n_n5287) & (n_n5288)) + ((x592x) & (x21x) & (n_n5294) & (n_n5287) & (!n_n5288)) + ((x592x) & (x21x) & (n_n5294) & (n_n5287) & (n_n5288)));
	assign x13371x = (((!x592x) & (!x24x) & (!n_n5290) & (!n_n5292) & (x441x)) + ((!x592x) & (!x24x) & (!n_n5290) & (n_n5292) & (!x441x)) + ((!x592x) & (!x24x) & (!n_n5290) & (n_n5292) & (x441x)) + ((!x592x) & (!x24x) & (n_n5290) & (!n_n5292) & (!x441x)) + ((!x592x) & (!x24x) & (n_n5290) & (!n_n5292) & (x441x)) + ((!x592x) & (!x24x) & (n_n5290) & (n_n5292) & (!x441x)) + ((!x592x) & (!x24x) & (n_n5290) & (n_n5292) & (x441x)) + ((!x592x) & (x24x) & (!n_n5290) & (!n_n5292) & (x441x)) + ((!x592x) & (x24x) & (!n_n5290) & (n_n5292) & (!x441x)) + ((!x592x) & (x24x) & (!n_n5290) & (n_n5292) & (x441x)) + ((!x592x) & (x24x) & (n_n5290) & (!n_n5292) & (!x441x)) + ((!x592x) & (x24x) & (n_n5290) & (!n_n5292) & (x441x)) + ((!x592x) & (x24x) & (n_n5290) & (n_n5292) & (!x441x)) + ((!x592x) & (x24x) & (n_n5290) & (n_n5292) & (x441x)) + ((x592x) & (!x24x) & (!n_n5290) & (!n_n5292) & (x441x)) + ((x592x) & (!x24x) & (!n_n5290) & (n_n5292) & (!x441x)) + ((x592x) & (!x24x) & (!n_n5290) & (n_n5292) & (x441x)) + ((x592x) & (!x24x) & (n_n5290) & (!n_n5292) & (!x441x)) + ((x592x) & (!x24x) & (n_n5290) & (!n_n5292) & (x441x)) + ((x592x) & (!x24x) & (n_n5290) & (n_n5292) & (!x441x)) + ((x592x) & (!x24x) & (n_n5290) & (n_n5292) & (x441x)) + ((x592x) & (x24x) & (!n_n5290) & (!n_n5292) & (!x441x)) + ((x592x) & (x24x) & (!n_n5290) & (!n_n5292) & (x441x)) + ((x592x) & (x24x) & (!n_n5290) & (n_n5292) & (!x441x)) + ((x592x) & (x24x) & (!n_n5290) & (n_n5292) & (x441x)) + ((x592x) & (x24x) & (n_n5290) & (!n_n5292) & (!x441x)) + ((x592x) & (x24x) & (n_n5290) & (!n_n5292) & (x441x)) + ((x592x) & (x24x) & (n_n5290) & (n_n5292) & (!x441x)) + ((x592x) & (x24x) & (n_n5290) & (n_n5292) & (x441x)));
	assign x13374x = (((!n_n4026) & (!n_n4028) & (!x13370x) & (x13371x)) + ((!n_n4026) & (!n_n4028) & (x13370x) & (!x13371x)) + ((!n_n4026) & (!n_n4028) & (x13370x) & (x13371x)) + ((!n_n4026) & (n_n4028) & (!x13370x) & (!x13371x)) + ((!n_n4026) & (n_n4028) & (!x13370x) & (x13371x)) + ((!n_n4026) & (n_n4028) & (x13370x) & (!x13371x)) + ((!n_n4026) & (n_n4028) & (x13370x) & (x13371x)) + ((n_n4026) & (!n_n4028) & (!x13370x) & (!x13371x)) + ((n_n4026) & (!n_n4028) & (!x13370x) & (x13371x)) + ((n_n4026) & (!n_n4028) & (x13370x) & (!x13371x)) + ((n_n4026) & (!n_n4028) & (x13370x) & (x13371x)) + ((n_n4026) & (n_n4028) & (!x13370x) & (!x13371x)) + ((n_n4026) & (n_n4028) & (!x13370x) & (x13371x)) + ((n_n4026) & (n_n4028) & (x13370x) & (!x13371x)) + ((n_n4026) & (n_n4028) & (x13370x) & (x13371x)));
	assign x343x = (((!i_7_) & (i_8_) & (!i_6_) & (x18x) & (n_n500)) + ((i_7_) & (!i_8_) & (!i_6_) & (x18x) & (n_n500)));
	assign x13383x = (((!i_9_) & (!n_n526) & (n_n528) & (n_n195) & (n_n500)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n195) & (n_n500)) + ((i_9_) & (!n_n526) & (n_n528) & (n_n195) & (n_n500)) + ((i_9_) & (n_n526) & (!n_n528) & (n_n195) & (n_n500)) + ((i_9_) & (n_n526) & (n_n528) & (n_n195) & (n_n500)));
	assign n_n4050 = (((!n_n5004) & (!x393x) & (!n_n5013) & (!x343x) & (x13383x)) + ((!n_n5004) & (!x393x) & (!n_n5013) & (x343x) & (!x13383x)) + ((!n_n5004) & (!x393x) & (!n_n5013) & (x343x) & (x13383x)) + ((!n_n5004) & (!x393x) & (n_n5013) & (!x343x) & (!x13383x)) + ((!n_n5004) & (!x393x) & (n_n5013) & (!x343x) & (x13383x)) + ((!n_n5004) & (!x393x) & (n_n5013) & (x343x) & (!x13383x)) + ((!n_n5004) & (!x393x) & (n_n5013) & (x343x) & (x13383x)) + ((!n_n5004) & (x393x) & (!n_n5013) & (!x343x) & (!x13383x)) + ((!n_n5004) & (x393x) & (!n_n5013) & (!x343x) & (x13383x)) + ((!n_n5004) & (x393x) & (!n_n5013) & (x343x) & (!x13383x)) + ((!n_n5004) & (x393x) & (!n_n5013) & (x343x) & (x13383x)) + ((!n_n5004) & (x393x) & (n_n5013) & (!x343x) & (!x13383x)) + ((!n_n5004) & (x393x) & (n_n5013) & (!x343x) & (x13383x)) + ((!n_n5004) & (x393x) & (n_n5013) & (x343x) & (!x13383x)) + ((!n_n5004) & (x393x) & (n_n5013) & (x343x) & (x13383x)) + ((n_n5004) & (!x393x) & (!n_n5013) & (!x343x) & (!x13383x)) + ((n_n5004) & (!x393x) & (!n_n5013) & (!x343x) & (x13383x)) + ((n_n5004) & (!x393x) & (!n_n5013) & (x343x) & (!x13383x)) + ((n_n5004) & (!x393x) & (!n_n5013) & (x343x) & (x13383x)) + ((n_n5004) & (!x393x) & (n_n5013) & (!x343x) & (!x13383x)) + ((n_n5004) & (!x393x) & (n_n5013) & (!x343x) & (x13383x)) + ((n_n5004) & (!x393x) & (n_n5013) & (x343x) & (!x13383x)) + ((n_n5004) & (!x393x) & (n_n5013) & (x343x) & (x13383x)) + ((n_n5004) & (x393x) & (!n_n5013) & (!x343x) & (!x13383x)) + ((n_n5004) & (x393x) & (!n_n5013) & (!x343x) & (x13383x)) + ((n_n5004) & (x393x) & (!n_n5013) & (x343x) & (!x13383x)) + ((n_n5004) & (x393x) & (!n_n5013) & (x343x) & (x13383x)) + ((n_n5004) & (x393x) & (n_n5013) & (!x343x) & (!x13383x)) + ((n_n5004) & (x393x) & (n_n5013) & (!x343x) & (x13383x)) + ((n_n5004) & (x393x) & (n_n5013) & (x343x) & (!x13383x)) + ((n_n5004) & (x393x) & (n_n5013) & (x343x) & (x13383x)));
	assign x90x = (((!n_n5076) & (!n_n5075) & (!n_n5078) & (!n_n5077) & (n_n5080)) + ((!n_n5076) & (!n_n5075) & (!n_n5078) & (n_n5077) & (!n_n5080)) + ((!n_n5076) & (!n_n5075) & (!n_n5078) & (n_n5077) & (n_n5080)) + ((!n_n5076) & (!n_n5075) & (n_n5078) & (!n_n5077) & (!n_n5080)) + ((!n_n5076) & (!n_n5075) & (n_n5078) & (!n_n5077) & (n_n5080)) + ((!n_n5076) & (!n_n5075) & (n_n5078) & (n_n5077) & (!n_n5080)) + ((!n_n5076) & (!n_n5075) & (n_n5078) & (n_n5077) & (n_n5080)) + ((!n_n5076) & (n_n5075) & (!n_n5078) & (!n_n5077) & (!n_n5080)) + ((!n_n5076) & (n_n5075) & (!n_n5078) & (!n_n5077) & (n_n5080)) + ((!n_n5076) & (n_n5075) & (!n_n5078) & (n_n5077) & (!n_n5080)) + ((!n_n5076) & (n_n5075) & (!n_n5078) & (n_n5077) & (n_n5080)) + ((!n_n5076) & (n_n5075) & (n_n5078) & (!n_n5077) & (!n_n5080)) + ((!n_n5076) & (n_n5075) & (n_n5078) & (!n_n5077) & (n_n5080)) + ((!n_n5076) & (n_n5075) & (n_n5078) & (n_n5077) & (!n_n5080)) + ((!n_n5076) & (n_n5075) & (n_n5078) & (n_n5077) & (n_n5080)) + ((n_n5076) & (!n_n5075) & (!n_n5078) & (!n_n5077) & (!n_n5080)) + ((n_n5076) & (!n_n5075) & (!n_n5078) & (!n_n5077) & (n_n5080)) + ((n_n5076) & (!n_n5075) & (!n_n5078) & (n_n5077) & (!n_n5080)) + ((n_n5076) & (!n_n5075) & (!n_n5078) & (n_n5077) & (n_n5080)) + ((n_n5076) & (!n_n5075) & (n_n5078) & (!n_n5077) & (!n_n5080)) + ((n_n5076) & (!n_n5075) & (n_n5078) & (!n_n5077) & (n_n5080)) + ((n_n5076) & (!n_n5075) & (n_n5078) & (n_n5077) & (!n_n5080)) + ((n_n5076) & (!n_n5075) & (n_n5078) & (n_n5077) & (n_n5080)) + ((n_n5076) & (n_n5075) & (!n_n5078) & (!n_n5077) & (!n_n5080)) + ((n_n5076) & (n_n5075) & (!n_n5078) & (!n_n5077) & (n_n5080)) + ((n_n5076) & (n_n5075) & (!n_n5078) & (n_n5077) & (!n_n5080)) + ((n_n5076) & (n_n5075) & (!n_n5078) & (n_n5077) & (n_n5080)) + ((n_n5076) & (n_n5075) & (n_n5078) & (!n_n5077) & (!n_n5080)) + ((n_n5076) & (n_n5075) & (n_n5078) & (!n_n5077) & (n_n5080)) + ((n_n5076) & (n_n5075) & (n_n5078) & (n_n5077) & (!n_n5080)) + ((n_n5076) & (n_n5075) & (n_n5078) & (n_n5077) & (n_n5080)));
	assign x404x = (((!i_9_) & (!n_n534) & (!n_n535) & (!n_n130) & (n_n5082)) + ((!i_9_) & (!n_n534) & (!n_n535) & (n_n130) & (n_n5082)) + ((!i_9_) & (!n_n534) & (n_n535) & (!n_n130) & (n_n5082)) + ((!i_9_) & (!n_n534) & (n_n535) & (n_n130) & (n_n5082)) + ((!i_9_) & (n_n534) & (!n_n535) & (!n_n130) & (n_n5082)) + ((!i_9_) & (n_n534) & (!n_n535) & (n_n130) & (n_n5082)) + ((!i_9_) & (n_n534) & (n_n535) & (!n_n130) & (n_n5082)) + ((!i_9_) & (n_n534) & (n_n535) & (n_n130) & (!n_n5082)) + ((!i_9_) & (n_n534) & (n_n535) & (n_n130) & (n_n5082)) + ((i_9_) & (!n_n534) & (!n_n535) & (!n_n130) & (n_n5082)) + ((i_9_) & (!n_n534) & (!n_n535) & (n_n130) & (n_n5082)) + ((i_9_) & (!n_n534) & (n_n535) & (!n_n130) & (n_n5082)) + ((i_9_) & (!n_n534) & (n_n535) & (n_n130) & (n_n5082)) + ((i_9_) & (n_n534) & (!n_n535) & (!n_n130) & (n_n5082)) + ((i_9_) & (n_n534) & (!n_n535) & (n_n130) & (n_n5082)) + ((i_9_) & (n_n534) & (n_n535) & (!n_n130) & (n_n5082)) + ((i_9_) & (n_n534) & (n_n535) & (n_n130) & (n_n5082)));
	assign x13396x = (((!n_n5057) & (!n_n5058) & (!n_n5067) & (!x160x) & (x275x)) + ((!n_n5057) & (!n_n5058) & (!n_n5067) & (x160x) & (!x275x)) + ((!n_n5057) & (!n_n5058) & (!n_n5067) & (x160x) & (x275x)) + ((!n_n5057) & (!n_n5058) & (n_n5067) & (!x160x) & (!x275x)) + ((!n_n5057) & (!n_n5058) & (n_n5067) & (!x160x) & (x275x)) + ((!n_n5057) & (!n_n5058) & (n_n5067) & (x160x) & (!x275x)) + ((!n_n5057) & (!n_n5058) & (n_n5067) & (x160x) & (x275x)) + ((!n_n5057) & (n_n5058) & (!n_n5067) & (!x160x) & (!x275x)) + ((!n_n5057) & (n_n5058) & (!n_n5067) & (!x160x) & (x275x)) + ((!n_n5057) & (n_n5058) & (!n_n5067) & (x160x) & (!x275x)) + ((!n_n5057) & (n_n5058) & (!n_n5067) & (x160x) & (x275x)) + ((!n_n5057) & (n_n5058) & (n_n5067) & (!x160x) & (!x275x)) + ((!n_n5057) & (n_n5058) & (n_n5067) & (!x160x) & (x275x)) + ((!n_n5057) & (n_n5058) & (n_n5067) & (x160x) & (!x275x)) + ((!n_n5057) & (n_n5058) & (n_n5067) & (x160x) & (x275x)) + ((n_n5057) & (!n_n5058) & (!n_n5067) & (!x160x) & (!x275x)) + ((n_n5057) & (!n_n5058) & (!n_n5067) & (!x160x) & (x275x)) + ((n_n5057) & (!n_n5058) & (!n_n5067) & (x160x) & (!x275x)) + ((n_n5057) & (!n_n5058) & (!n_n5067) & (x160x) & (x275x)) + ((n_n5057) & (!n_n5058) & (n_n5067) & (!x160x) & (!x275x)) + ((n_n5057) & (!n_n5058) & (n_n5067) & (!x160x) & (x275x)) + ((n_n5057) & (!n_n5058) & (n_n5067) & (x160x) & (!x275x)) + ((n_n5057) & (!n_n5058) & (n_n5067) & (x160x) & (x275x)) + ((n_n5057) & (n_n5058) & (!n_n5067) & (!x160x) & (!x275x)) + ((n_n5057) & (n_n5058) & (!n_n5067) & (!x160x) & (x275x)) + ((n_n5057) & (n_n5058) & (!n_n5067) & (x160x) & (!x275x)) + ((n_n5057) & (n_n5058) & (!n_n5067) & (x160x) & (x275x)) + ((n_n5057) & (n_n5058) & (n_n5067) & (!x160x) & (!x275x)) + ((n_n5057) & (n_n5058) & (n_n5067) & (!x160x) & (x275x)) + ((n_n5057) & (n_n5058) & (n_n5067) & (x160x) & (!x275x)) + ((n_n5057) & (n_n5058) & (n_n5067) & (x160x) & (x275x)));
	assign x13398x = (((!n_n5084) & (!n_n5079) & (!x90x) & (!x404x) & (x13396x)) + ((!n_n5084) & (!n_n5079) & (!x90x) & (x404x) & (!x13396x)) + ((!n_n5084) & (!n_n5079) & (!x90x) & (x404x) & (x13396x)) + ((!n_n5084) & (!n_n5079) & (x90x) & (!x404x) & (!x13396x)) + ((!n_n5084) & (!n_n5079) & (x90x) & (!x404x) & (x13396x)) + ((!n_n5084) & (!n_n5079) & (x90x) & (x404x) & (!x13396x)) + ((!n_n5084) & (!n_n5079) & (x90x) & (x404x) & (x13396x)) + ((!n_n5084) & (n_n5079) & (!x90x) & (!x404x) & (!x13396x)) + ((!n_n5084) & (n_n5079) & (!x90x) & (!x404x) & (x13396x)) + ((!n_n5084) & (n_n5079) & (!x90x) & (x404x) & (!x13396x)) + ((!n_n5084) & (n_n5079) & (!x90x) & (x404x) & (x13396x)) + ((!n_n5084) & (n_n5079) & (x90x) & (!x404x) & (!x13396x)) + ((!n_n5084) & (n_n5079) & (x90x) & (!x404x) & (x13396x)) + ((!n_n5084) & (n_n5079) & (x90x) & (x404x) & (!x13396x)) + ((!n_n5084) & (n_n5079) & (x90x) & (x404x) & (x13396x)) + ((n_n5084) & (!n_n5079) & (!x90x) & (!x404x) & (!x13396x)) + ((n_n5084) & (!n_n5079) & (!x90x) & (!x404x) & (x13396x)) + ((n_n5084) & (!n_n5079) & (!x90x) & (x404x) & (!x13396x)) + ((n_n5084) & (!n_n5079) & (!x90x) & (x404x) & (x13396x)) + ((n_n5084) & (!n_n5079) & (x90x) & (!x404x) & (!x13396x)) + ((n_n5084) & (!n_n5079) & (x90x) & (!x404x) & (x13396x)) + ((n_n5084) & (!n_n5079) & (x90x) & (x404x) & (!x13396x)) + ((n_n5084) & (!n_n5079) & (x90x) & (x404x) & (x13396x)) + ((n_n5084) & (n_n5079) & (!x90x) & (!x404x) & (!x13396x)) + ((n_n5084) & (n_n5079) & (!x90x) & (!x404x) & (x13396x)) + ((n_n5084) & (n_n5079) & (!x90x) & (x404x) & (!x13396x)) + ((n_n5084) & (n_n5079) & (!x90x) & (x404x) & (x13396x)) + ((n_n5084) & (n_n5079) & (x90x) & (!x404x) & (!x13396x)) + ((n_n5084) & (n_n5079) & (x90x) & (!x404x) & (x13396x)) + ((n_n5084) & (n_n5079) & (x90x) & (x404x) & (!x13396x)) + ((n_n5084) & (n_n5079) & (x90x) & (x404x) & (x13396x)));
	assign n_n1952 = (((!i_9_) & (!n_n528) & (n_n195) & (n_n530) & (n_n464)) + ((!i_9_) & (n_n528) & (n_n195) & (!n_n530) & (n_n464)) + ((!i_9_) & (n_n528) & (n_n195) & (n_n530) & (n_n464)) + ((i_9_) & (n_n528) & (n_n195) & (!n_n530) & (n_n464)) + ((i_9_) & (n_n528) & (n_n195) & (n_n530) & (n_n464)));
	assign n_n789 = (((!i_9_) & (!n_n534) & (!n_n195) & (!n_n464) & (n_n5063)) + ((!i_9_) & (!n_n534) & (!n_n195) & (n_n464) & (n_n5063)) + ((!i_9_) & (!n_n534) & (n_n195) & (!n_n464) & (n_n5063)) + ((!i_9_) & (!n_n534) & (n_n195) & (n_n464) & (n_n5063)) + ((!i_9_) & (n_n534) & (!n_n195) & (!n_n464) & (n_n5063)) + ((!i_9_) & (n_n534) & (!n_n195) & (n_n464) & (n_n5063)) + ((!i_9_) & (n_n534) & (n_n195) & (!n_n464) & (n_n5063)) + ((!i_9_) & (n_n534) & (n_n195) & (n_n464) & (!n_n5063)) + ((!i_9_) & (n_n534) & (n_n195) & (n_n464) & (n_n5063)) + ((i_9_) & (!n_n534) & (!n_n195) & (!n_n464) & (n_n5063)) + ((i_9_) & (!n_n534) & (!n_n195) & (n_n464) & (n_n5063)) + ((i_9_) & (!n_n534) & (n_n195) & (!n_n464) & (n_n5063)) + ((i_9_) & (!n_n534) & (n_n195) & (n_n464) & (n_n5063)) + ((i_9_) & (n_n534) & (!n_n195) & (!n_n464) & (n_n5063)) + ((i_9_) & (n_n534) & (!n_n195) & (n_n464) & (n_n5063)) + ((i_9_) & (n_n534) & (n_n195) & (!n_n464) & (n_n5063)) + ((i_9_) & (n_n534) & (n_n195) & (n_n464) & (!n_n5063)) + ((i_9_) & (n_n534) & (n_n195) & (n_n464) & (n_n5063)));
	assign x13394x = (((!x21x) & (!x11x) & (!n_n473) & (!n_n195) & (n_n4152)) + ((!x21x) & (!x11x) & (!n_n473) & (n_n195) & (n_n4152)) + ((!x21x) & (!x11x) & (n_n473) & (!n_n195) & (n_n4152)) + ((!x21x) & (!x11x) & (n_n473) & (n_n195) & (n_n4152)) + ((!x21x) & (x11x) & (!n_n473) & (!n_n195) & (n_n4152)) + ((!x21x) & (x11x) & (!n_n473) & (n_n195) & (n_n4152)) + ((!x21x) & (x11x) & (n_n473) & (!n_n195) & (n_n4152)) + ((!x21x) & (x11x) & (n_n473) & (n_n195) & (!n_n4152)) + ((!x21x) & (x11x) & (n_n473) & (n_n195) & (n_n4152)) + ((x21x) & (!x11x) & (!n_n473) & (!n_n195) & (n_n4152)) + ((x21x) & (!x11x) & (!n_n473) & (n_n195) & (n_n4152)) + ((x21x) & (!x11x) & (n_n473) & (!n_n195) & (n_n4152)) + ((x21x) & (!x11x) & (n_n473) & (n_n195) & (!n_n4152)) + ((x21x) & (!x11x) & (n_n473) & (n_n195) & (n_n4152)) + ((x21x) & (x11x) & (!n_n473) & (!n_n195) & (n_n4152)) + ((x21x) & (x11x) & (!n_n473) & (n_n195) & (n_n4152)) + ((x21x) & (x11x) & (n_n473) & (!n_n195) & (n_n4152)) + ((x21x) & (x11x) & (n_n473) & (n_n195) & (!n_n4152)) + ((x21x) & (x11x) & (n_n473) & (n_n195) & (n_n4152)));
	assign n_n4003 = (((!x13398x) & (!n_n1952) & (!n_n789) & (x13394x)) + ((!x13398x) & (!n_n1952) & (n_n789) & (!x13394x)) + ((!x13398x) & (!n_n1952) & (n_n789) & (x13394x)) + ((!x13398x) & (n_n1952) & (!n_n789) & (!x13394x)) + ((!x13398x) & (n_n1952) & (!n_n789) & (x13394x)) + ((!x13398x) & (n_n1952) & (n_n789) & (!x13394x)) + ((!x13398x) & (n_n1952) & (n_n789) & (x13394x)) + ((x13398x) & (!n_n1952) & (!n_n789) & (!x13394x)) + ((x13398x) & (!n_n1952) & (!n_n789) & (x13394x)) + ((x13398x) & (!n_n1952) & (n_n789) & (!x13394x)) + ((x13398x) & (!n_n1952) & (n_n789) & (x13394x)) + ((x13398x) & (n_n1952) & (!n_n789) & (!x13394x)) + ((x13398x) & (n_n1952) & (!n_n789) & (x13394x)) + ((x13398x) & (n_n1952) & (n_n789) & (!x13394x)) + ((x13398x) & (n_n1952) & (n_n789) & (x13394x)));
	assign x13414x = (((!n_n3424) & (!n_n5018) & (!n_n5014) & (!n_n5019) & (n_n4161)) + ((!n_n3424) & (!n_n5018) & (!n_n5014) & (n_n5019) & (!n_n4161)) + ((!n_n3424) & (!n_n5018) & (!n_n5014) & (n_n5019) & (n_n4161)) + ((!n_n3424) & (!n_n5018) & (n_n5014) & (!n_n5019) & (!n_n4161)) + ((!n_n3424) & (!n_n5018) & (n_n5014) & (!n_n5019) & (n_n4161)) + ((!n_n3424) & (!n_n5018) & (n_n5014) & (n_n5019) & (!n_n4161)) + ((!n_n3424) & (!n_n5018) & (n_n5014) & (n_n5019) & (n_n4161)) + ((!n_n3424) & (n_n5018) & (!n_n5014) & (!n_n5019) & (!n_n4161)) + ((!n_n3424) & (n_n5018) & (!n_n5014) & (!n_n5019) & (n_n4161)) + ((!n_n3424) & (n_n5018) & (!n_n5014) & (n_n5019) & (!n_n4161)) + ((!n_n3424) & (n_n5018) & (!n_n5014) & (n_n5019) & (n_n4161)) + ((!n_n3424) & (n_n5018) & (n_n5014) & (!n_n5019) & (!n_n4161)) + ((!n_n3424) & (n_n5018) & (n_n5014) & (!n_n5019) & (n_n4161)) + ((!n_n3424) & (n_n5018) & (n_n5014) & (n_n5019) & (!n_n4161)) + ((!n_n3424) & (n_n5018) & (n_n5014) & (n_n5019) & (n_n4161)) + ((n_n3424) & (!n_n5018) & (!n_n5014) & (!n_n5019) & (!n_n4161)) + ((n_n3424) & (!n_n5018) & (!n_n5014) & (!n_n5019) & (n_n4161)) + ((n_n3424) & (!n_n5018) & (!n_n5014) & (n_n5019) & (!n_n4161)) + ((n_n3424) & (!n_n5018) & (!n_n5014) & (n_n5019) & (n_n4161)) + ((n_n3424) & (!n_n5018) & (n_n5014) & (!n_n5019) & (!n_n4161)) + ((n_n3424) & (!n_n5018) & (n_n5014) & (!n_n5019) & (n_n4161)) + ((n_n3424) & (!n_n5018) & (n_n5014) & (n_n5019) & (!n_n4161)) + ((n_n3424) & (!n_n5018) & (n_n5014) & (n_n5019) & (n_n4161)) + ((n_n3424) & (n_n5018) & (!n_n5014) & (!n_n5019) & (!n_n4161)) + ((n_n3424) & (n_n5018) & (!n_n5014) & (!n_n5019) & (n_n4161)) + ((n_n3424) & (n_n5018) & (!n_n5014) & (n_n5019) & (!n_n4161)) + ((n_n3424) & (n_n5018) & (!n_n5014) & (n_n5019) & (n_n4161)) + ((n_n3424) & (n_n5018) & (n_n5014) & (!n_n5019) & (!n_n4161)) + ((n_n3424) & (n_n5018) & (n_n5014) & (!n_n5019) & (n_n4161)) + ((n_n3424) & (n_n5018) & (n_n5014) & (n_n5019) & (!n_n4161)) + ((n_n3424) & (n_n5018) & (n_n5014) & (n_n5019) & (n_n4161)));
	assign n_n4047 = (((!n_n5050) & (!n_n5054) & (!n_n5048) & (!n_n5049) & (x13405x)) + ((!n_n5050) & (!n_n5054) & (!n_n5048) & (n_n5049) & (!x13405x)) + ((!n_n5050) & (!n_n5054) & (!n_n5048) & (n_n5049) & (x13405x)) + ((!n_n5050) & (!n_n5054) & (n_n5048) & (!n_n5049) & (!x13405x)) + ((!n_n5050) & (!n_n5054) & (n_n5048) & (!n_n5049) & (x13405x)) + ((!n_n5050) & (!n_n5054) & (n_n5048) & (n_n5049) & (!x13405x)) + ((!n_n5050) & (!n_n5054) & (n_n5048) & (n_n5049) & (x13405x)) + ((!n_n5050) & (n_n5054) & (!n_n5048) & (!n_n5049) & (!x13405x)) + ((!n_n5050) & (n_n5054) & (!n_n5048) & (!n_n5049) & (x13405x)) + ((!n_n5050) & (n_n5054) & (!n_n5048) & (n_n5049) & (!x13405x)) + ((!n_n5050) & (n_n5054) & (!n_n5048) & (n_n5049) & (x13405x)) + ((!n_n5050) & (n_n5054) & (n_n5048) & (!n_n5049) & (!x13405x)) + ((!n_n5050) & (n_n5054) & (n_n5048) & (!n_n5049) & (x13405x)) + ((!n_n5050) & (n_n5054) & (n_n5048) & (n_n5049) & (!x13405x)) + ((!n_n5050) & (n_n5054) & (n_n5048) & (n_n5049) & (x13405x)) + ((n_n5050) & (!n_n5054) & (!n_n5048) & (!n_n5049) & (!x13405x)) + ((n_n5050) & (!n_n5054) & (!n_n5048) & (!n_n5049) & (x13405x)) + ((n_n5050) & (!n_n5054) & (!n_n5048) & (n_n5049) & (!x13405x)) + ((n_n5050) & (!n_n5054) & (!n_n5048) & (n_n5049) & (x13405x)) + ((n_n5050) & (!n_n5054) & (n_n5048) & (!n_n5049) & (!x13405x)) + ((n_n5050) & (!n_n5054) & (n_n5048) & (!n_n5049) & (x13405x)) + ((n_n5050) & (!n_n5054) & (n_n5048) & (n_n5049) & (!x13405x)) + ((n_n5050) & (!n_n5054) & (n_n5048) & (n_n5049) & (x13405x)) + ((n_n5050) & (n_n5054) & (!n_n5048) & (!n_n5049) & (!x13405x)) + ((n_n5050) & (n_n5054) & (!n_n5048) & (!n_n5049) & (x13405x)) + ((n_n5050) & (n_n5054) & (!n_n5048) & (n_n5049) & (!x13405x)) + ((n_n5050) & (n_n5054) & (!n_n5048) & (n_n5049) & (x13405x)) + ((n_n5050) & (n_n5054) & (n_n5048) & (!n_n5049) & (!x13405x)) + ((n_n5050) & (n_n5054) & (n_n5048) & (!n_n5049) & (x13405x)) + ((n_n5050) & (n_n5054) & (n_n5048) & (n_n5049) & (!x13405x)) + ((n_n5050) & (n_n5054) & (n_n5048) & (n_n5049) & (x13405x)));
	assign n_n4048 = (((!x50x) & (!n_n5042) & (!n_n5043) & (!n_n5029) & (!x22124x)) + ((!x50x) & (!n_n5042) & (!n_n5043) & (n_n5029) & (!x22124x)) + ((!x50x) & (!n_n5042) & (!n_n5043) & (n_n5029) & (x22124x)) + ((!x50x) & (!n_n5042) & (n_n5043) & (!n_n5029) & (!x22124x)) + ((!x50x) & (!n_n5042) & (n_n5043) & (!n_n5029) & (x22124x)) + ((!x50x) & (!n_n5042) & (n_n5043) & (n_n5029) & (!x22124x)) + ((!x50x) & (!n_n5042) & (n_n5043) & (n_n5029) & (x22124x)) + ((!x50x) & (n_n5042) & (!n_n5043) & (!n_n5029) & (!x22124x)) + ((!x50x) & (n_n5042) & (!n_n5043) & (!n_n5029) & (x22124x)) + ((!x50x) & (n_n5042) & (!n_n5043) & (n_n5029) & (!x22124x)) + ((!x50x) & (n_n5042) & (!n_n5043) & (n_n5029) & (x22124x)) + ((!x50x) & (n_n5042) & (n_n5043) & (!n_n5029) & (!x22124x)) + ((!x50x) & (n_n5042) & (n_n5043) & (!n_n5029) & (x22124x)) + ((!x50x) & (n_n5042) & (n_n5043) & (n_n5029) & (!x22124x)) + ((!x50x) & (n_n5042) & (n_n5043) & (n_n5029) & (x22124x)) + ((x50x) & (!n_n5042) & (!n_n5043) & (!n_n5029) & (!x22124x)) + ((x50x) & (!n_n5042) & (!n_n5043) & (!n_n5029) & (x22124x)) + ((x50x) & (!n_n5042) & (!n_n5043) & (n_n5029) & (!x22124x)) + ((x50x) & (!n_n5042) & (!n_n5043) & (n_n5029) & (x22124x)) + ((x50x) & (!n_n5042) & (n_n5043) & (!n_n5029) & (!x22124x)) + ((x50x) & (!n_n5042) & (n_n5043) & (!n_n5029) & (x22124x)) + ((x50x) & (!n_n5042) & (n_n5043) & (n_n5029) & (!x22124x)) + ((x50x) & (!n_n5042) & (n_n5043) & (n_n5029) & (x22124x)) + ((x50x) & (n_n5042) & (!n_n5043) & (!n_n5029) & (!x22124x)) + ((x50x) & (n_n5042) & (!n_n5043) & (!n_n5029) & (x22124x)) + ((x50x) & (n_n5042) & (!n_n5043) & (n_n5029) & (!x22124x)) + ((x50x) & (n_n5042) & (!n_n5043) & (n_n5029) & (x22124x)) + ((x50x) & (n_n5042) & (n_n5043) & (!n_n5029) & (!x22124x)) + ((x50x) & (n_n5042) & (n_n5043) & (!n_n5029) & (x22124x)) + ((x50x) & (n_n5042) & (n_n5043) & (n_n5029) & (!x22124x)) + ((x50x) & (n_n5042) & (n_n5043) & (n_n5029) & (x22124x)));
	assign n_n4004 = (((!x13414x) & (!n_n4047) & (n_n4048)) + ((!x13414x) & (n_n4047) & (!n_n4048)) + ((!x13414x) & (n_n4047) & (n_n4048)) + ((x13414x) & (!n_n4047) & (!n_n4048)) + ((x13414x) & (!n_n4047) & (n_n4048)) + ((x13414x) & (n_n4047) & (!n_n4048)) + ((x13414x) & (n_n4047) & (n_n4048)));
	assign x13421x = (((!n_n4982) & (!n_n4981) & (!n_n4979) & (!n_n4978) & (x13420x)) + ((!n_n4982) & (!n_n4981) & (!n_n4979) & (n_n4978) & (!x13420x)) + ((!n_n4982) & (!n_n4981) & (!n_n4979) & (n_n4978) & (x13420x)) + ((!n_n4982) & (!n_n4981) & (n_n4979) & (!n_n4978) & (!x13420x)) + ((!n_n4982) & (!n_n4981) & (n_n4979) & (!n_n4978) & (x13420x)) + ((!n_n4982) & (!n_n4981) & (n_n4979) & (n_n4978) & (!x13420x)) + ((!n_n4982) & (!n_n4981) & (n_n4979) & (n_n4978) & (x13420x)) + ((!n_n4982) & (n_n4981) & (!n_n4979) & (!n_n4978) & (!x13420x)) + ((!n_n4982) & (n_n4981) & (!n_n4979) & (!n_n4978) & (x13420x)) + ((!n_n4982) & (n_n4981) & (!n_n4979) & (n_n4978) & (!x13420x)) + ((!n_n4982) & (n_n4981) & (!n_n4979) & (n_n4978) & (x13420x)) + ((!n_n4982) & (n_n4981) & (n_n4979) & (!n_n4978) & (!x13420x)) + ((!n_n4982) & (n_n4981) & (n_n4979) & (!n_n4978) & (x13420x)) + ((!n_n4982) & (n_n4981) & (n_n4979) & (n_n4978) & (!x13420x)) + ((!n_n4982) & (n_n4981) & (n_n4979) & (n_n4978) & (x13420x)) + ((n_n4982) & (!n_n4981) & (!n_n4979) & (!n_n4978) & (!x13420x)) + ((n_n4982) & (!n_n4981) & (!n_n4979) & (!n_n4978) & (x13420x)) + ((n_n4982) & (!n_n4981) & (!n_n4979) & (n_n4978) & (!x13420x)) + ((n_n4982) & (!n_n4981) & (!n_n4979) & (n_n4978) & (x13420x)) + ((n_n4982) & (!n_n4981) & (n_n4979) & (!n_n4978) & (!x13420x)) + ((n_n4982) & (!n_n4981) & (n_n4979) & (!n_n4978) & (x13420x)) + ((n_n4982) & (!n_n4981) & (n_n4979) & (n_n4978) & (!x13420x)) + ((n_n4982) & (!n_n4981) & (n_n4979) & (n_n4978) & (x13420x)) + ((n_n4982) & (n_n4981) & (!n_n4979) & (!n_n4978) & (!x13420x)) + ((n_n4982) & (n_n4981) & (!n_n4979) & (!n_n4978) & (x13420x)) + ((n_n4982) & (n_n4981) & (!n_n4979) & (n_n4978) & (!x13420x)) + ((n_n4982) & (n_n4981) & (!n_n4979) & (n_n4978) & (x13420x)) + ((n_n4982) & (n_n4981) & (n_n4979) & (!n_n4978) & (!x13420x)) + ((n_n4982) & (n_n4981) & (n_n4979) & (!n_n4978) & (x13420x)) + ((n_n4982) & (n_n4981) & (n_n4979) & (n_n4978) & (!x13420x)) + ((n_n4982) & (n_n4981) & (n_n4979) & (n_n4978) & (x13420x)));
	assign n_n4650 = (((i_9_) & (n_n482) & (n_n390) & (n_n532)));
	assign x14659x = (((!n_n5050) & (!n_n5054) & (!n_n5048) & (n_n5047)) + ((!n_n5050) & (!n_n5054) & (n_n5048) & (!n_n5047)) + ((!n_n5050) & (!n_n5054) & (n_n5048) & (n_n5047)) + ((!n_n5050) & (n_n5054) & (!n_n5048) & (!n_n5047)) + ((!n_n5050) & (n_n5054) & (!n_n5048) & (n_n5047)) + ((!n_n5050) & (n_n5054) & (n_n5048) & (!n_n5047)) + ((!n_n5050) & (n_n5054) & (n_n5048) & (n_n5047)) + ((n_n5050) & (!n_n5054) & (!n_n5048) & (!n_n5047)) + ((n_n5050) & (!n_n5054) & (!n_n5048) & (n_n5047)) + ((n_n5050) & (!n_n5054) & (n_n5048) & (!n_n5047)) + ((n_n5050) & (!n_n5054) & (n_n5048) & (n_n5047)) + ((n_n5050) & (n_n5054) & (!n_n5048) & (!n_n5047)) + ((n_n5050) & (n_n5054) & (!n_n5048) & (n_n5047)) + ((n_n5050) & (n_n5054) & (n_n5048) & (!n_n5047)) + ((n_n5050) & (n_n5054) & (n_n5048) & (n_n5047)));
	assign x14660x = (((!n_n5055) & (!n_n5045) & (!n_n5056) & (!n_n5053) & (n_n5051)) + ((!n_n5055) & (!n_n5045) & (!n_n5056) & (n_n5053) & (!n_n5051)) + ((!n_n5055) & (!n_n5045) & (!n_n5056) & (n_n5053) & (n_n5051)) + ((!n_n5055) & (!n_n5045) & (n_n5056) & (!n_n5053) & (!n_n5051)) + ((!n_n5055) & (!n_n5045) & (n_n5056) & (!n_n5053) & (n_n5051)) + ((!n_n5055) & (!n_n5045) & (n_n5056) & (n_n5053) & (!n_n5051)) + ((!n_n5055) & (!n_n5045) & (n_n5056) & (n_n5053) & (n_n5051)) + ((!n_n5055) & (n_n5045) & (!n_n5056) & (!n_n5053) & (!n_n5051)) + ((!n_n5055) & (n_n5045) & (!n_n5056) & (!n_n5053) & (n_n5051)) + ((!n_n5055) & (n_n5045) & (!n_n5056) & (n_n5053) & (!n_n5051)) + ((!n_n5055) & (n_n5045) & (!n_n5056) & (n_n5053) & (n_n5051)) + ((!n_n5055) & (n_n5045) & (n_n5056) & (!n_n5053) & (!n_n5051)) + ((!n_n5055) & (n_n5045) & (n_n5056) & (!n_n5053) & (n_n5051)) + ((!n_n5055) & (n_n5045) & (n_n5056) & (n_n5053) & (!n_n5051)) + ((!n_n5055) & (n_n5045) & (n_n5056) & (n_n5053) & (n_n5051)) + ((n_n5055) & (!n_n5045) & (!n_n5056) & (!n_n5053) & (!n_n5051)) + ((n_n5055) & (!n_n5045) & (!n_n5056) & (!n_n5053) & (n_n5051)) + ((n_n5055) & (!n_n5045) & (!n_n5056) & (n_n5053) & (!n_n5051)) + ((n_n5055) & (!n_n5045) & (!n_n5056) & (n_n5053) & (n_n5051)) + ((n_n5055) & (!n_n5045) & (n_n5056) & (!n_n5053) & (!n_n5051)) + ((n_n5055) & (!n_n5045) & (n_n5056) & (!n_n5053) & (n_n5051)) + ((n_n5055) & (!n_n5045) & (n_n5056) & (n_n5053) & (!n_n5051)) + ((n_n5055) & (!n_n5045) & (n_n5056) & (n_n5053) & (n_n5051)) + ((n_n5055) & (n_n5045) & (!n_n5056) & (!n_n5053) & (!n_n5051)) + ((n_n5055) & (n_n5045) & (!n_n5056) & (!n_n5053) & (n_n5051)) + ((n_n5055) & (n_n5045) & (!n_n5056) & (n_n5053) & (!n_n5051)) + ((n_n5055) & (n_n5045) & (!n_n5056) & (n_n5053) & (n_n5051)) + ((n_n5055) & (n_n5045) & (n_n5056) & (!n_n5053) & (!n_n5051)) + ((n_n5055) & (n_n5045) & (n_n5056) & (!n_n5053) & (n_n5051)) + ((n_n5055) & (n_n5045) & (n_n5056) & (n_n5053) & (!n_n5051)) + ((n_n5055) & (n_n5045) & (n_n5056) & (n_n5053) & (n_n5051)));
	assign x253x = (((!i_9_) & (n_n482) & (n_n534) & (n_n195)) + ((i_9_) & (n_n482) & (n_n534) & (n_n195)));
	assign x14665x = (((!n_n524) & (!n_n482) & (!x18x) & (!n_n5025) & (x97x)) + ((!n_n524) & (!n_n482) & (!x18x) & (n_n5025) & (!x97x)) + ((!n_n524) & (!n_n482) & (!x18x) & (n_n5025) & (x97x)) + ((!n_n524) & (!n_n482) & (x18x) & (!n_n5025) & (x97x)) + ((!n_n524) & (!n_n482) & (x18x) & (n_n5025) & (!x97x)) + ((!n_n524) & (!n_n482) & (x18x) & (n_n5025) & (x97x)) + ((!n_n524) & (n_n482) & (!x18x) & (!n_n5025) & (x97x)) + ((!n_n524) & (n_n482) & (!x18x) & (n_n5025) & (!x97x)) + ((!n_n524) & (n_n482) & (!x18x) & (n_n5025) & (x97x)) + ((!n_n524) & (n_n482) & (x18x) & (!n_n5025) & (x97x)) + ((!n_n524) & (n_n482) & (x18x) & (n_n5025) & (!x97x)) + ((!n_n524) & (n_n482) & (x18x) & (n_n5025) & (x97x)) + ((n_n524) & (!n_n482) & (!x18x) & (!n_n5025) & (x97x)) + ((n_n524) & (!n_n482) & (!x18x) & (n_n5025) & (!x97x)) + ((n_n524) & (!n_n482) & (!x18x) & (n_n5025) & (x97x)) + ((n_n524) & (!n_n482) & (x18x) & (!n_n5025) & (x97x)) + ((n_n524) & (!n_n482) & (x18x) & (n_n5025) & (!x97x)) + ((n_n524) & (!n_n482) & (x18x) & (n_n5025) & (x97x)) + ((n_n524) & (n_n482) & (!x18x) & (!n_n5025) & (x97x)) + ((n_n524) & (n_n482) & (!x18x) & (n_n5025) & (!x97x)) + ((n_n524) & (n_n482) & (!x18x) & (n_n5025) & (x97x)) + ((n_n524) & (n_n482) & (x18x) & (!n_n5025) & (!x97x)) + ((n_n524) & (n_n482) & (x18x) & (!n_n5025) & (x97x)) + ((n_n524) & (n_n482) & (x18x) & (n_n5025) & (!x97x)) + ((n_n524) & (n_n482) & (x18x) & (n_n5025) & (x97x)));
	assign x14666x = (((!n_n5038) & (!n_n5035) & (!n_n5037) & (!n_n5039) & (x153x)) + ((!n_n5038) & (!n_n5035) & (!n_n5037) & (n_n5039) & (!x153x)) + ((!n_n5038) & (!n_n5035) & (!n_n5037) & (n_n5039) & (x153x)) + ((!n_n5038) & (!n_n5035) & (n_n5037) & (!n_n5039) & (!x153x)) + ((!n_n5038) & (!n_n5035) & (n_n5037) & (!n_n5039) & (x153x)) + ((!n_n5038) & (!n_n5035) & (n_n5037) & (n_n5039) & (!x153x)) + ((!n_n5038) & (!n_n5035) & (n_n5037) & (n_n5039) & (x153x)) + ((!n_n5038) & (n_n5035) & (!n_n5037) & (!n_n5039) & (!x153x)) + ((!n_n5038) & (n_n5035) & (!n_n5037) & (!n_n5039) & (x153x)) + ((!n_n5038) & (n_n5035) & (!n_n5037) & (n_n5039) & (!x153x)) + ((!n_n5038) & (n_n5035) & (!n_n5037) & (n_n5039) & (x153x)) + ((!n_n5038) & (n_n5035) & (n_n5037) & (!n_n5039) & (!x153x)) + ((!n_n5038) & (n_n5035) & (n_n5037) & (!n_n5039) & (x153x)) + ((!n_n5038) & (n_n5035) & (n_n5037) & (n_n5039) & (!x153x)) + ((!n_n5038) & (n_n5035) & (n_n5037) & (n_n5039) & (x153x)) + ((n_n5038) & (!n_n5035) & (!n_n5037) & (!n_n5039) & (!x153x)) + ((n_n5038) & (!n_n5035) & (!n_n5037) & (!n_n5039) & (x153x)) + ((n_n5038) & (!n_n5035) & (!n_n5037) & (n_n5039) & (!x153x)) + ((n_n5038) & (!n_n5035) & (!n_n5037) & (n_n5039) & (x153x)) + ((n_n5038) & (!n_n5035) & (n_n5037) & (!n_n5039) & (!x153x)) + ((n_n5038) & (!n_n5035) & (n_n5037) & (!n_n5039) & (x153x)) + ((n_n5038) & (!n_n5035) & (n_n5037) & (n_n5039) & (!x153x)) + ((n_n5038) & (!n_n5035) & (n_n5037) & (n_n5039) & (x153x)) + ((n_n5038) & (n_n5035) & (!n_n5037) & (!n_n5039) & (!x153x)) + ((n_n5038) & (n_n5035) & (!n_n5037) & (!n_n5039) & (x153x)) + ((n_n5038) & (n_n5035) & (!n_n5037) & (n_n5039) & (!x153x)) + ((n_n5038) & (n_n5035) & (!n_n5037) & (n_n5039) & (x153x)) + ((n_n5038) & (n_n5035) & (n_n5037) & (!n_n5039) & (!x153x)) + ((n_n5038) & (n_n5035) & (n_n5037) & (!n_n5039) & (x153x)) + ((n_n5038) & (n_n5035) & (n_n5037) & (n_n5039) & (!x153x)) + ((n_n5038) & (n_n5035) & (n_n5037) & (n_n5039) & (x153x)));
	assign x125x = (((!i_9_) & (!n_n532) & (n_n534) & (n_n491) & (n_n130)) + ((!i_9_) & (n_n532) & (!n_n534) & (n_n491) & (n_n130)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n491) & (n_n130)));
	assign n_n5197 = (((!i_9_) & (n_n130) & (n_n530) & (n_n464)));
	assign n_n5205 = (((!i_1_) & (i_2_) & (!i_0_) & (x20x) & (n_n464)));
	assign n_n5211 = (((!i_9_) & (n_n532) & (n_n535) & (n_n65)));
	assign n_n5071 = (((!i_9_) & (n_n528) & (n_n195) & (n_n464)));
	assign n_n5226 = (((!i_5_) & (i_3_) & (i_4_) & (x19x) & (n_n532)));
	assign n_n5218 = (((i_7_) & (!i_8_) & (!i_6_) & (x19x) & (n_n535)));
	assign n_n5256 = (((i_7_) & (i_8_) & (i_6_) & (x19x) & (n_n500)));
	assign n_n5257 = (((!i_9_) & (n_n534) & (n_n500) & (n_n65)));
	assign n_n5283 = (((!i_9_) & (n_n524) & (n_n491) & (n_n65)));
	assign n_n5250 = (((i_7_) & (!i_8_) & (!i_6_) & (x19x) & (n_n509)));
	assign n_n3412 = (((!n_n524) & (!n_n518) & (!n_n526) & (!x12x) & (n_n5105)) + ((!n_n524) & (!n_n518) & (!n_n526) & (x12x) & (n_n5105)) + ((!n_n524) & (!n_n518) & (n_n526) & (!x12x) & (n_n5105)) + ((!n_n524) & (!n_n518) & (n_n526) & (x12x) & (n_n5105)) + ((!n_n524) & (n_n518) & (!n_n526) & (!x12x) & (n_n5105)) + ((!n_n524) & (n_n518) & (!n_n526) & (x12x) & (n_n5105)) + ((!n_n524) & (n_n518) & (n_n526) & (!x12x) & (n_n5105)) + ((!n_n524) & (n_n518) & (n_n526) & (x12x) & (!n_n5105)) + ((!n_n524) & (n_n518) & (n_n526) & (x12x) & (n_n5105)) + ((n_n524) & (!n_n518) & (!n_n526) & (!x12x) & (n_n5105)) + ((n_n524) & (!n_n518) & (!n_n526) & (x12x) & (n_n5105)) + ((n_n524) & (!n_n518) & (n_n526) & (!x12x) & (n_n5105)) + ((n_n524) & (!n_n518) & (n_n526) & (x12x) & (n_n5105)) + ((n_n524) & (n_n518) & (!n_n526) & (!x12x) & (n_n5105)) + ((n_n524) & (n_n518) & (!n_n526) & (x12x) & (!n_n5105)) + ((n_n524) & (n_n518) & (!n_n526) & (x12x) & (n_n5105)) + ((n_n524) & (n_n518) & (n_n526) & (!x12x) & (n_n5105)) + ((n_n524) & (n_n518) & (n_n526) & (x12x) & (!n_n5105)) + ((n_n524) & (n_n518) & (n_n526) & (x12x) & (n_n5105)));
	assign x191x = (((!i_9_) & (!n_n526) & (n_n482) & (n_n528) & (n_n325)) + ((!i_9_) & (n_n526) & (n_n482) & (n_n528) & (n_n325)) + ((i_9_) & (n_n526) & (n_n482) & (!n_n528) & (n_n325)) + ((i_9_) & (n_n526) & (n_n482) & (n_n528) & (n_n325)));
	assign x13789x = (((!n_n4782) & (!x131x) & (!n_n4789) & (n_n4788)) + ((!n_n4782) & (!x131x) & (n_n4789) & (!n_n4788)) + ((!n_n4782) & (!x131x) & (n_n4789) & (n_n4788)) + ((!n_n4782) & (x131x) & (!n_n4789) & (!n_n4788)) + ((!n_n4782) & (x131x) & (!n_n4789) & (n_n4788)) + ((!n_n4782) & (x131x) & (n_n4789) & (!n_n4788)) + ((!n_n4782) & (x131x) & (n_n4789) & (n_n4788)) + ((n_n4782) & (!x131x) & (!n_n4789) & (!n_n4788)) + ((n_n4782) & (!x131x) & (!n_n4789) & (n_n4788)) + ((n_n4782) & (!x131x) & (n_n4789) & (!n_n4788)) + ((n_n4782) & (!x131x) & (n_n4789) & (n_n4788)) + ((n_n4782) & (x131x) & (!n_n4789) & (!n_n4788)) + ((n_n4782) & (x131x) & (!n_n4789) & (n_n4788)) + ((n_n4782) & (x131x) & (n_n4789) & (!n_n4788)) + ((n_n4782) & (x131x) & (n_n4789) & (n_n4788)));
	assign n_n3333 = (((!n_n4784) & (!n_n4790) & (!n_n4791) & (!n_n4783) & (x13789x)) + ((!n_n4784) & (!n_n4790) & (!n_n4791) & (n_n4783) & (!x13789x)) + ((!n_n4784) & (!n_n4790) & (!n_n4791) & (n_n4783) & (x13789x)) + ((!n_n4784) & (!n_n4790) & (n_n4791) & (!n_n4783) & (!x13789x)) + ((!n_n4784) & (!n_n4790) & (n_n4791) & (!n_n4783) & (x13789x)) + ((!n_n4784) & (!n_n4790) & (n_n4791) & (n_n4783) & (!x13789x)) + ((!n_n4784) & (!n_n4790) & (n_n4791) & (n_n4783) & (x13789x)) + ((!n_n4784) & (n_n4790) & (!n_n4791) & (!n_n4783) & (!x13789x)) + ((!n_n4784) & (n_n4790) & (!n_n4791) & (!n_n4783) & (x13789x)) + ((!n_n4784) & (n_n4790) & (!n_n4791) & (n_n4783) & (!x13789x)) + ((!n_n4784) & (n_n4790) & (!n_n4791) & (n_n4783) & (x13789x)) + ((!n_n4784) & (n_n4790) & (n_n4791) & (!n_n4783) & (!x13789x)) + ((!n_n4784) & (n_n4790) & (n_n4791) & (!n_n4783) & (x13789x)) + ((!n_n4784) & (n_n4790) & (n_n4791) & (n_n4783) & (!x13789x)) + ((!n_n4784) & (n_n4790) & (n_n4791) & (n_n4783) & (x13789x)) + ((n_n4784) & (!n_n4790) & (!n_n4791) & (!n_n4783) & (!x13789x)) + ((n_n4784) & (!n_n4790) & (!n_n4791) & (!n_n4783) & (x13789x)) + ((n_n4784) & (!n_n4790) & (!n_n4791) & (n_n4783) & (!x13789x)) + ((n_n4784) & (!n_n4790) & (!n_n4791) & (n_n4783) & (x13789x)) + ((n_n4784) & (!n_n4790) & (n_n4791) & (!n_n4783) & (!x13789x)) + ((n_n4784) & (!n_n4790) & (n_n4791) & (!n_n4783) & (x13789x)) + ((n_n4784) & (!n_n4790) & (n_n4791) & (n_n4783) & (!x13789x)) + ((n_n4784) & (!n_n4790) & (n_n4791) & (n_n4783) & (x13789x)) + ((n_n4784) & (n_n4790) & (!n_n4791) & (!n_n4783) & (!x13789x)) + ((n_n4784) & (n_n4790) & (!n_n4791) & (!n_n4783) & (x13789x)) + ((n_n4784) & (n_n4790) & (!n_n4791) & (n_n4783) & (!x13789x)) + ((n_n4784) & (n_n4790) & (!n_n4791) & (n_n4783) & (x13789x)) + ((n_n4784) & (n_n4790) & (n_n4791) & (!n_n4783) & (!x13789x)) + ((n_n4784) & (n_n4790) & (n_n4791) & (!n_n4783) & (x13789x)) + ((n_n4784) & (n_n4790) & (n_n4791) & (n_n4783) & (!x13789x)) + ((n_n4784) & (n_n4790) & (n_n4791) & (n_n4783) & (x13789x)));
	assign x13994x = (((!i_9_) & (!n_n534) & (n_n491) & (n_n195) & (n_n530)) + ((!i_9_) & (n_n534) & (n_n491) & (n_n195) & (n_n530)) + ((i_9_) & (n_n534) & (n_n491) & (n_n195) & (!n_n530)) + ((i_9_) & (n_n534) & (n_n491) & (n_n195) & (n_n530)));
	assign n_n3315 = (((!n_n5018) & (!n_n5015) & (!x298x) & (!n_n4161) & (x13994x)) + ((!n_n5018) & (!n_n5015) & (!x298x) & (n_n4161) & (!x13994x)) + ((!n_n5018) & (!n_n5015) & (!x298x) & (n_n4161) & (x13994x)) + ((!n_n5018) & (!n_n5015) & (x298x) & (!n_n4161) & (!x13994x)) + ((!n_n5018) & (!n_n5015) & (x298x) & (!n_n4161) & (x13994x)) + ((!n_n5018) & (!n_n5015) & (x298x) & (n_n4161) & (!x13994x)) + ((!n_n5018) & (!n_n5015) & (x298x) & (n_n4161) & (x13994x)) + ((!n_n5018) & (n_n5015) & (!x298x) & (!n_n4161) & (!x13994x)) + ((!n_n5018) & (n_n5015) & (!x298x) & (!n_n4161) & (x13994x)) + ((!n_n5018) & (n_n5015) & (!x298x) & (n_n4161) & (!x13994x)) + ((!n_n5018) & (n_n5015) & (!x298x) & (n_n4161) & (x13994x)) + ((!n_n5018) & (n_n5015) & (x298x) & (!n_n4161) & (!x13994x)) + ((!n_n5018) & (n_n5015) & (x298x) & (!n_n4161) & (x13994x)) + ((!n_n5018) & (n_n5015) & (x298x) & (n_n4161) & (!x13994x)) + ((!n_n5018) & (n_n5015) & (x298x) & (n_n4161) & (x13994x)) + ((n_n5018) & (!n_n5015) & (!x298x) & (!n_n4161) & (!x13994x)) + ((n_n5018) & (!n_n5015) & (!x298x) & (!n_n4161) & (x13994x)) + ((n_n5018) & (!n_n5015) & (!x298x) & (n_n4161) & (!x13994x)) + ((n_n5018) & (!n_n5015) & (!x298x) & (n_n4161) & (x13994x)) + ((n_n5018) & (!n_n5015) & (x298x) & (!n_n4161) & (!x13994x)) + ((n_n5018) & (!n_n5015) & (x298x) & (!n_n4161) & (x13994x)) + ((n_n5018) & (!n_n5015) & (x298x) & (n_n4161) & (!x13994x)) + ((n_n5018) & (!n_n5015) & (x298x) & (n_n4161) & (x13994x)) + ((n_n5018) & (n_n5015) & (!x298x) & (!n_n4161) & (!x13994x)) + ((n_n5018) & (n_n5015) & (!x298x) & (!n_n4161) & (x13994x)) + ((n_n5018) & (n_n5015) & (!x298x) & (n_n4161) & (!x13994x)) + ((n_n5018) & (n_n5015) & (!x298x) & (n_n4161) & (x13994x)) + ((n_n5018) & (n_n5015) & (x298x) & (!n_n4161) & (!x13994x)) + ((n_n5018) & (n_n5015) & (x298x) & (!n_n4161) & (x13994x)) + ((n_n5018) & (n_n5015) & (x298x) & (n_n4161) & (!x13994x)) + ((n_n5018) & (n_n5015) & (x298x) & (n_n4161) & (x13994x)));
	assign n_n3771 = (((!x15x) & (!n_n130) & (!n_n500) & (!n_n5137) & (n_n5136)) + ((!x15x) & (!n_n130) & (!n_n500) & (n_n5137) & (!n_n5136)) + ((!x15x) & (!n_n130) & (!n_n500) & (n_n5137) & (n_n5136)) + ((!x15x) & (!n_n130) & (n_n500) & (!n_n5137) & (n_n5136)) + ((!x15x) & (!n_n130) & (n_n500) & (n_n5137) & (!n_n5136)) + ((!x15x) & (!n_n130) & (n_n500) & (n_n5137) & (n_n5136)) + ((!x15x) & (n_n130) & (!n_n500) & (!n_n5137) & (n_n5136)) + ((!x15x) & (n_n130) & (!n_n500) & (n_n5137) & (!n_n5136)) + ((!x15x) & (n_n130) & (!n_n500) & (n_n5137) & (n_n5136)) + ((!x15x) & (n_n130) & (n_n500) & (!n_n5137) & (n_n5136)) + ((!x15x) & (n_n130) & (n_n500) & (n_n5137) & (!n_n5136)) + ((!x15x) & (n_n130) & (n_n500) & (n_n5137) & (n_n5136)) + ((x15x) & (!n_n130) & (!n_n500) & (!n_n5137) & (n_n5136)) + ((x15x) & (!n_n130) & (!n_n500) & (n_n5137) & (!n_n5136)) + ((x15x) & (!n_n130) & (!n_n500) & (n_n5137) & (n_n5136)) + ((x15x) & (!n_n130) & (n_n500) & (!n_n5137) & (n_n5136)) + ((x15x) & (!n_n130) & (n_n500) & (n_n5137) & (!n_n5136)) + ((x15x) & (!n_n130) & (n_n500) & (n_n5137) & (n_n5136)) + ((x15x) & (n_n130) & (!n_n500) & (!n_n5137) & (n_n5136)) + ((x15x) & (n_n130) & (!n_n500) & (n_n5137) & (!n_n5136)) + ((x15x) & (n_n130) & (!n_n500) & (n_n5137) & (n_n5136)) + ((x15x) & (n_n130) & (n_n500) & (!n_n5137) & (!n_n5136)) + ((x15x) & (n_n130) & (n_n500) & (!n_n5137) & (n_n5136)) + ((x15x) & (n_n130) & (n_n500) & (n_n5137) & (!n_n5136)) + ((x15x) & (n_n130) & (n_n500) & (n_n5137) & (n_n5136)));
	assign n_n4654 = (((i_9_) & (n_n482) & (n_n528) & (n_n390)));
	assign x140x = (((!i_9_) & (n_n482) & (n_n390) & (n_n532)) + ((i_9_) & (n_n482) & (n_n390) & (n_n532)));
	assign n_n4657 = (((!i_9_) & (n_n526) & (n_n482) & (n_n390)));
	assign x13887x = (((!i_9_) & (!n_n526) & (n_n482) & (n_n390) & (n_n532)) + ((!i_9_) & (n_n526) & (n_n482) & (n_n390) & (!n_n532)) + ((!i_9_) & (n_n526) & (n_n482) & (n_n390) & (n_n532)) + ((i_9_) & (!n_n526) & (n_n482) & (n_n390) & (n_n532)) + ((i_9_) & (n_n526) & (n_n482) & (n_n390) & (!n_n532)) + ((i_9_) & (n_n526) & (n_n482) & (n_n390) & (n_n532)));
	assign n_n2987 = (((!n_n4649) & (!x311x) & (!n_n4655) & (!n_n4654) & (x13887x)) + ((!n_n4649) & (!x311x) & (!n_n4655) & (n_n4654) & (!x13887x)) + ((!n_n4649) & (!x311x) & (!n_n4655) & (n_n4654) & (x13887x)) + ((!n_n4649) & (!x311x) & (n_n4655) & (!n_n4654) & (!x13887x)) + ((!n_n4649) & (!x311x) & (n_n4655) & (!n_n4654) & (x13887x)) + ((!n_n4649) & (!x311x) & (n_n4655) & (n_n4654) & (!x13887x)) + ((!n_n4649) & (!x311x) & (n_n4655) & (n_n4654) & (x13887x)) + ((!n_n4649) & (x311x) & (!n_n4655) & (!n_n4654) & (!x13887x)) + ((!n_n4649) & (x311x) & (!n_n4655) & (!n_n4654) & (x13887x)) + ((!n_n4649) & (x311x) & (!n_n4655) & (n_n4654) & (!x13887x)) + ((!n_n4649) & (x311x) & (!n_n4655) & (n_n4654) & (x13887x)) + ((!n_n4649) & (x311x) & (n_n4655) & (!n_n4654) & (!x13887x)) + ((!n_n4649) & (x311x) & (n_n4655) & (!n_n4654) & (x13887x)) + ((!n_n4649) & (x311x) & (n_n4655) & (n_n4654) & (!x13887x)) + ((!n_n4649) & (x311x) & (n_n4655) & (n_n4654) & (x13887x)) + ((n_n4649) & (!x311x) & (!n_n4655) & (!n_n4654) & (!x13887x)) + ((n_n4649) & (!x311x) & (!n_n4655) & (!n_n4654) & (x13887x)) + ((n_n4649) & (!x311x) & (!n_n4655) & (n_n4654) & (!x13887x)) + ((n_n4649) & (!x311x) & (!n_n4655) & (n_n4654) & (x13887x)) + ((n_n4649) & (!x311x) & (n_n4655) & (!n_n4654) & (!x13887x)) + ((n_n4649) & (!x311x) & (n_n4655) & (!n_n4654) & (x13887x)) + ((n_n4649) & (!x311x) & (n_n4655) & (n_n4654) & (!x13887x)) + ((n_n4649) & (!x311x) & (n_n4655) & (n_n4654) & (x13887x)) + ((n_n4649) & (x311x) & (!n_n4655) & (!n_n4654) & (!x13887x)) + ((n_n4649) & (x311x) & (!n_n4655) & (!n_n4654) & (x13887x)) + ((n_n4649) & (x311x) & (!n_n4655) & (n_n4654) & (!x13887x)) + ((n_n4649) & (x311x) & (!n_n4655) & (n_n4654) & (x13887x)) + ((n_n4649) & (x311x) & (n_n4655) & (!n_n4654) & (!x13887x)) + ((n_n4649) & (x311x) & (n_n4655) & (!n_n4654) & (x13887x)) + ((n_n4649) & (x311x) & (n_n4655) & (n_n4654) & (!x13887x)) + ((n_n4649) & (x311x) & (n_n4655) & (n_n4654) & (x13887x)));
	assign n_n4665 = (((!i_9_) & (n_n390) & (n_n473) & (n_n534)));
	assign x72x = (((!i_9_) & (!n_n524) & (n_n482) & (n_n390) & (x20x)) + ((!i_9_) & (n_n524) & (n_n482) & (n_n390) & (!x20x)) + ((!i_9_) & (n_n524) & (n_n482) & (n_n390) & (x20x)) + ((i_9_) & (!n_n524) & (n_n482) & (n_n390) & (x20x)) + ((i_9_) & (n_n524) & (n_n482) & (n_n390) & (x20x)));
	assign x11854x = (((!i_9_) & (!n_n524) & (n_n390) & (n_n473) & (x20x)) + ((!i_9_) & (n_n524) & (n_n390) & (n_n473) & (x20x)) + ((i_9_) & (!n_n524) & (n_n390) & (n_n473) & (x20x)) + ((i_9_) & (n_n524) & (n_n390) & (n_n473) & (!x20x)) + ((i_9_) & (n_n524) & (n_n390) & (n_n473) & (x20x)));
	assign x192x = (((!n_n4675) & (!n_n4676) & (!n_n4679) & (!n_n4678) & (x11854x)) + ((!n_n4675) & (!n_n4676) & (!n_n4679) & (n_n4678) & (!x11854x)) + ((!n_n4675) & (!n_n4676) & (!n_n4679) & (n_n4678) & (x11854x)) + ((!n_n4675) & (!n_n4676) & (n_n4679) & (!n_n4678) & (!x11854x)) + ((!n_n4675) & (!n_n4676) & (n_n4679) & (!n_n4678) & (x11854x)) + ((!n_n4675) & (!n_n4676) & (n_n4679) & (n_n4678) & (!x11854x)) + ((!n_n4675) & (!n_n4676) & (n_n4679) & (n_n4678) & (x11854x)) + ((!n_n4675) & (n_n4676) & (!n_n4679) & (!n_n4678) & (!x11854x)) + ((!n_n4675) & (n_n4676) & (!n_n4679) & (!n_n4678) & (x11854x)) + ((!n_n4675) & (n_n4676) & (!n_n4679) & (n_n4678) & (!x11854x)) + ((!n_n4675) & (n_n4676) & (!n_n4679) & (n_n4678) & (x11854x)) + ((!n_n4675) & (n_n4676) & (n_n4679) & (!n_n4678) & (!x11854x)) + ((!n_n4675) & (n_n4676) & (n_n4679) & (!n_n4678) & (x11854x)) + ((!n_n4675) & (n_n4676) & (n_n4679) & (n_n4678) & (!x11854x)) + ((!n_n4675) & (n_n4676) & (n_n4679) & (n_n4678) & (x11854x)) + ((n_n4675) & (!n_n4676) & (!n_n4679) & (!n_n4678) & (!x11854x)) + ((n_n4675) & (!n_n4676) & (!n_n4679) & (!n_n4678) & (x11854x)) + ((n_n4675) & (!n_n4676) & (!n_n4679) & (n_n4678) & (!x11854x)) + ((n_n4675) & (!n_n4676) & (!n_n4679) & (n_n4678) & (x11854x)) + ((n_n4675) & (!n_n4676) & (n_n4679) & (!n_n4678) & (!x11854x)) + ((n_n4675) & (!n_n4676) & (n_n4679) & (!n_n4678) & (x11854x)) + ((n_n4675) & (!n_n4676) & (n_n4679) & (n_n4678) & (!x11854x)) + ((n_n4675) & (!n_n4676) & (n_n4679) & (n_n4678) & (x11854x)) + ((n_n4675) & (n_n4676) & (!n_n4679) & (!n_n4678) & (!x11854x)) + ((n_n4675) & (n_n4676) & (!n_n4679) & (!n_n4678) & (x11854x)) + ((n_n4675) & (n_n4676) & (!n_n4679) & (n_n4678) & (!x11854x)) + ((n_n4675) & (n_n4676) & (!n_n4679) & (n_n4678) & (x11854x)) + ((n_n4675) & (n_n4676) & (n_n4679) & (!n_n4678) & (!x11854x)) + ((n_n4675) & (n_n4676) & (n_n4679) & (!n_n4678) & (x11854x)) + ((n_n4675) & (n_n4676) & (n_n4679) & (n_n4678) & (!x11854x)) + ((n_n4675) & (n_n4676) & (n_n4679) & (n_n4678) & (x11854x)));
	assign x193x = (((!i_9_) & (!n_n526) & (n_n528) & (n_n390) & (n_n473)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n390) & (n_n473)) + ((i_9_) & (n_n526) & (!n_n528) & (n_n390) & (n_n473)) + ((i_9_) & (n_n526) & (n_n528) & (n_n390) & (n_n473)));
	assign n_n4680 = (((i_9_) & (n_n390) & (n_n534) & (n_n464)));
	assign x13893x = (((!n_n4673) & (!n_n4658) & (!n_n4684) & (n_n4665)) + ((!n_n4673) & (!n_n4658) & (n_n4684) & (!n_n4665)) + ((!n_n4673) & (!n_n4658) & (n_n4684) & (n_n4665)) + ((!n_n4673) & (n_n4658) & (!n_n4684) & (!n_n4665)) + ((!n_n4673) & (n_n4658) & (!n_n4684) & (n_n4665)) + ((!n_n4673) & (n_n4658) & (n_n4684) & (!n_n4665)) + ((!n_n4673) & (n_n4658) & (n_n4684) & (n_n4665)) + ((n_n4673) & (!n_n4658) & (!n_n4684) & (!n_n4665)) + ((n_n4673) & (!n_n4658) & (!n_n4684) & (n_n4665)) + ((n_n4673) & (!n_n4658) & (n_n4684) & (!n_n4665)) + ((n_n4673) & (!n_n4658) & (n_n4684) & (n_n4665)) + ((n_n4673) & (n_n4658) & (!n_n4684) & (!n_n4665)) + ((n_n4673) & (n_n4658) & (!n_n4684) & (n_n4665)) + ((n_n4673) & (n_n4658) & (n_n4684) & (!n_n4665)) + ((n_n4673) & (n_n4658) & (n_n4684) & (n_n4665)));
	assign x13894x = (((!n_n4681) & (!x338x) & (!x72x) & (!x193x) & (n_n4680)) + ((!n_n4681) & (!x338x) & (!x72x) & (x193x) & (!n_n4680)) + ((!n_n4681) & (!x338x) & (!x72x) & (x193x) & (n_n4680)) + ((!n_n4681) & (!x338x) & (x72x) & (!x193x) & (!n_n4680)) + ((!n_n4681) & (!x338x) & (x72x) & (!x193x) & (n_n4680)) + ((!n_n4681) & (!x338x) & (x72x) & (x193x) & (!n_n4680)) + ((!n_n4681) & (!x338x) & (x72x) & (x193x) & (n_n4680)) + ((!n_n4681) & (x338x) & (!x72x) & (!x193x) & (!n_n4680)) + ((!n_n4681) & (x338x) & (!x72x) & (!x193x) & (n_n4680)) + ((!n_n4681) & (x338x) & (!x72x) & (x193x) & (!n_n4680)) + ((!n_n4681) & (x338x) & (!x72x) & (x193x) & (n_n4680)) + ((!n_n4681) & (x338x) & (x72x) & (!x193x) & (!n_n4680)) + ((!n_n4681) & (x338x) & (x72x) & (!x193x) & (n_n4680)) + ((!n_n4681) & (x338x) & (x72x) & (x193x) & (!n_n4680)) + ((!n_n4681) & (x338x) & (x72x) & (x193x) & (n_n4680)) + ((n_n4681) & (!x338x) & (!x72x) & (!x193x) & (!n_n4680)) + ((n_n4681) & (!x338x) & (!x72x) & (!x193x) & (n_n4680)) + ((n_n4681) & (!x338x) & (!x72x) & (x193x) & (!n_n4680)) + ((n_n4681) & (!x338x) & (!x72x) & (x193x) & (n_n4680)) + ((n_n4681) & (!x338x) & (x72x) & (!x193x) & (!n_n4680)) + ((n_n4681) & (!x338x) & (x72x) & (!x193x) & (n_n4680)) + ((n_n4681) & (!x338x) & (x72x) & (x193x) & (!n_n4680)) + ((n_n4681) & (!x338x) & (x72x) & (x193x) & (n_n4680)) + ((n_n4681) & (x338x) & (!x72x) & (!x193x) & (!n_n4680)) + ((n_n4681) & (x338x) & (!x72x) & (!x193x) & (n_n4680)) + ((n_n4681) & (x338x) & (!x72x) & (x193x) & (!n_n4680)) + ((n_n4681) & (x338x) & (!x72x) & (x193x) & (n_n4680)) + ((n_n4681) & (x338x) & (x72x) & (!x193x) & (!n_n4680)) + ((n_n4681) & (x338x) & (x72x) & (!x193x) & (n_n4680)) + ((n_n4681) & (x338x) & (x72x) & (x193x) & (!n_n4680)) + ((n_n4681) & (x338x) & (x72x) & (x193x) & (n_n4680)));
	assign n_n3280 = (((!n_n2987) & (!x192x) & (!x13893x) & (x13894x)) + ((!n_n2987) & (!x192x) & (x13893x) & (!x13894x)) + ((!n_n2987) & (!x192x) & (x13893x) & (x13894x)) + ((!n_n2987) & (x192x) & (!x13893x) & (!x13894x)) + ((!n_n2987) & (x192x) & (!x13893x) & (x13894x)) + ((!n_n2987) & (x192x) & (x13893x) & (!x13894x)) + ((!n_n2987) & (x192x) & (x13893x) & (x13894x)) + ((n_n2987) & (!x192x) & (!x13893x) & (!x13894x)) + ((n_n2987) & (!x192x) & (!x13893x) & (x13894x)) + ((n_n2987) & (!x192x) & (x13893x) & (!x13894x)) + ((n_n2987) & (!x192x) & (x13893x) & (x13894x)) + ((n_n2987) & (x192x) & (!x13893x) & (!x13894x)) + ((n_n2987) & (x192x) & (!x13893x) & (x13894x)) + ((n_n2987) & (x192x) & (x13893x) & (!x13894x)) + ((n_n2987) & (x192x) & (x13893x) & (x13894x)));
	assign x41x = (((!i_9_) & (!n_n528) & (n_n509) & (n_n195) & (n_n530)) + ((!i_9_) & (n_n528) & (n_n509) & (n_n195) & (!n_n530)) + ((!i_9_) & (n_n528) & (n_n509) & (n_n195) & (n_n530)) + ((i_9_) & (n_n528) & (n_n509) & (n_n195) & (!n_n530)) + ((i_9_) & (n_n528) & (n_n509) & (n_n195) & (n_n530)));
	assign x248x = (((!i_9_) & (!n_n524) & (n_n509) & (n_n195) & (x20x)) + ((!i_9_) & (n_n524) & (n_n509) & (n_n195) & (!x20x)) + ((!i_9_) & (n_n524) & (n_n509) & (n_n195) & (x20x)) + ((i_9_) & (!n_n524) & (n_n509) & (n_n195) & (x20x)) + ((i_9_) & (n_n524) & (n_n509) & (n_n195) & (x20x)));
	assign n_n3317 = (((!n_n4998) & (!x103x) & (!n_n4993) & (!x41x) & (x248x)) + ((!n_n4998) & (!x103x) & (!n_n4993) & (x41x) & (!x248x)) + ((!n_n4998) & (!x103x) & (!n_n4993) & (x41x) & (x248x)) + ((!n_n4998) & (!x103x) & (n_n4993) & (!x41x) & (!x248x)) + ((!n_n4998) & (!x103x) & (n_n4993) & (!x41x) & (x248x)) + ((!n_n4998) & (!x103x) & (n_n4993) & (x41x) & (!x248x)) + ((!n_n4998) & (!x103x) & (n_n4993) & (x41x) & (x248x)) + ((!n_n4998) & (x103x) & (!n_n4993) & (!x41x) & (!x248x)) + ((!n_n4998) & (x103x) & (!n_n4993) & (!x41x) & (x248x)) + ((!n_n4998) & (x103x) & (!n_n4993) & (x41x) & (!x248x)) + ((!n_n4998) & (x103x) & (!n_n4993) & (x41x) & (x248x)) + ((!n_n4998) & (x103x) & (n_n4993) & (!x41x) & (!x248x)) + ((!n_n4998) & (x103x) & (n_n4993) & (!x41x) & (x248x)) + ((!n_n4998) & (x103x) & (n_n4993) & (x41x) & (!x248x)) + ((!n_n4998) & (x103x) & (n_n4993) & (x41x) & (x248x)) + ((n_n4998) & (!x103x) & (!n_n4993) & (!x41x) & (!x248x)) + ((n_n4998) & (!x103x) & (!n_n4993) & (!x41x) & (x248x)) + ((n_n4998) & (!x103x) & (!n_n4993) & (x41x) & (!x248x)) + ((n_n4998) & (!x103x) & (!n_n4993) & (x41x) & (x248x)) + ((n_n4998) & (!x103x) & (n_n4993) & (!x41x) & (!x248x)) + ((n_n4998) & (!x103x) & (n_n4993) & (!x41x) & (x248x)) + ((n_n4998) & (!x103x) & (n_n4993) & (x41x) & (!x248x)) + ((n_n4998) & (!x103x) & (n_n4993) & (x41x) & (x248x)) + ((n_n4998) & (x103x) & (!n_n4993) & (!x41x) & (!x248x)) + ((n_n4998) & (x103x) & (!n_n4993) & (!x41x) & (x248x)) + ((n_n4998) & (x103x) & (!n_n4993) & (x41x) & (!x248x)) + ((n_n4998) & (x103x) & (!n_n4993) & (x41x) & (x248x)) + ((n_n4998) & (x103x) & (n_n4993) & (!x41x) & (!x248x)) + ((n_n4998) & (x103x) & (n_n4993) & (!x41x) & (x248x)) + ((n_n4998) & (x103x) & (n_n4993) & (x41x) & (!x248x)) + ((n_n4998) & (x103x) & (n_n4993) & (x41x) & (x248x)));
	assign n_n4273 = (((!n_n536) & (!x23x) & (!n_n500) & (x423x)) + ((!n_n536) & (!x23x) & (n_n500) & (x423x)) + ((!n_n536) & (x23x) & (!n_n500) & (x423x)) + ((!n_n536) & (x23x) & (n_n500) & (x423x)) + ((n_n536) & (!x23x) & (!n_n500) & (x423x)) + ((n_n536) & (!x23x) & (n_n500) & (x423x)) + ((n_n536) & (x23x) & (!n_n500) & (x423x)) + ((n_n536) & (x23x) & (n_n500) & (!x423x)) + ((n_n536) & (x23x) & (n_n500) & (x423x)));
	assign x22113x = (((!n_n4361) & (!n_n4360) & (!n_n4357) & (!n_n4356)));
	assign n_n3367 = (((!n_n4358) & (!n_n4353) & (!n_n4354) & (!x399x) & (!x22113x)) + ((!n_n4358) & (!n_n4353) & (!n_n4354) & (x399x) & (!x22113x)) + ((!n_n4358) & (!n_n4353) & (!n_n4354) & (x399x) & (x22113x)) + ((!n_n4358) & (!n_n4353) & (n_n4354) & (!x399x) & (!x22113x)) + ((!n_n4358) & (!n_n4353) & (n_n4354) & (!x399x) & (x22113x)) + ((!n_n4358) & (!n_n4353) & (n_n4354) & (x399x) & (!x22113x)) + ((!n_n4358) & (!n_n4353) & (n_n4354) & (x399x) & (x22113x)) + ((!n_n4358) & (n_n4353) & (!n_n4354) & (!x399x) & (!x22113x)) + ((!n_n4358) & (n_n4353) & (!n_n4354) & (!x399x) & (x22113x)) + ((!n_n4358) & (n_n4353) & (!n_n4354) & (x399x) & (!x22113x)) + ((!n_n4358) & (n_n4353) & (!n_n4354) & (x399x) & (x22113x)) + ((!n_n4358) & (n_n4353) & (n_n4354) & (!x399x) & (!x22113x)) + ((!n_n4358) & (n_n4353) & (n_n4354) & (!x399x) & (x22113x)) + ((!n_n4358) & (n_n4353) & (n_n4354) & (x399x) & (!x22113x)) + ((!n_n4358) & (n_n4353) & (n_n4354) & (x399x) & (x22113x)) + ((n_n4358) & (!n_n4353) & (!n_n4354) & (!x399x) & (!x22113x)) + ((n_n4358) & (!n_n4353) & (!n_n4354) & (!x399x) & (x22113x)) + ((n_n4358) & (!n_n4353) & (!n_n4354) & (x399x) & (!x22113x)) + ((n_n4358) & (!n_n4353) & (!n_n4354) & (x399x) & (x22113x)) + ((n_n4358) & (!n_n4353) & (n_n4354) & (!x399x) & (!x22113x)) + ((n_n4358) & (!n_n4353) & (n_n4354) & (!x399x) & (x22113x)) + ((n_n4358) & (!n_n4353) & (n_n4354) & (x399x) & (!x22113x)) + ((n_n4358) & (!n_n4353) & (n_n4354) & (x399x) & (x22113x)) + ((n_n4358) & (n_n4353) & (!n_n4354) & (!x399x) & (!x22113x)) + ((n_n4358) & (n_n4353) & (!n_n4354) & (!x399x) & (x22113x)) + ((n_n4358) & (n_n4353) & (!n_n4354) & (x399x) & (!x22113x)) + ((n_n4358) & (n_n4353) & (!n_n4354) & (x399x) & (x22113x)) + ((n_n4358) & (n_n4353) & (n_n4354) & (!x399x) & (!x22113x)) + ((n_n4358) & (n_n4353) & (n_n4354) & (!x399x) & (x22113x)) + ((n_n4358) & (n_n4353) & (n_n4354) & (x399x) & (!x22113x)) + ((n_n4358) & (n_n4353) & (n_n4354) & (x399x) & (x22113x)));
	assign x301x = (((!i_9_) & (n_n536) & (!n_n520) & (x20x) & (n_n500)) + ((!i_9_) & (n_n536) & (n_n520) & (x20x) & (n_n500)) + ((i_9_) & (n_n536) & (!n_n520) & (x20x) & (n_n500)) + ((i_9_) & (n_n536) & (n_n520) & (!x20x) & (n_n500)) + ((i_9_) & (n_n536) & (n_n520) & (x20x) & (n_n500)));
	assign x14163x = (((!n_n4371) & (!n_n3533) & (!n_n1308) & (!n_n4370) & (n_n4273)) + ((!n_n4371) & (!n_n3533) & (!n_n1308) & (n_n4370) & (!n_n4273)) + ((!n_n4371) & (!n_n3533) & (!n_n1308) & (n_n4370) & (n_n4273)) + ((!n_n4371) & (!n_n3533) & (n_n1308) & (!n_n4370) & (!n_n4273)) + ((!n_n4371) & (!n_n3533) & (n_n1308) & (!n_n4370) & (n_n4273)) + ((!n_n4371) & (!n_n3533) & (n_n1308) & (n_n4370) & (!n_n4273)) + ((!n_n4371) & (!n_n3533) & (n_n1308) & (n_n4370) & (n_n4273)) + ((!n_n4371) & (n_n3533) & (!n_n1308) & (!n_n4370) & (!n_n4273)) + ((!n_n4371) & (n_n3533) & (!n_n1308) & (!n_n4370) & (n_n4273)) + ((!n_n4371) & (n_n3533) & (!n_n1308) & (n_n4370) & (!n_n4273)) + ((!n_n4371) & (n_n3533) & (!n_n1308) & (n_n4370) & (n_n4273)) + ((!n_n4371) & (n_n3533) & (n_n1308) & (!n_n4370) & (!n_n4273)) + ((!n_n4371) & (n_n3533) & (n_n1308) & (!n_n4370) & (n_n4273)) + ((!n_n4371) & (n_n3533) & (n_n1308) & (n_n4370) & (!n_n4273)) + ((!n_n4371) & (n_n3533) & (n_n1308) & (n_n4370) & (n_n4273)) + ((n_n4371) & (!n_n3533) & (!n_n1308) & (!n_n4370) & (!n_n4273)) + ((n_n4371) & (!n_n3533) & (!n_n1308) & (!n_n4370) & (n_n4273)) + ((n_n4371) & (!n_n3533) & (!n_n1308) & (n_n4370) & (!n_n4273)) + ((n_n4371) & (!n_n3533) & (!n_n1308) & (n_n4370) & (n_n4273)) + ((n_n4371) & (!n_n3533) & (n_n1308) & (!n_n4370) & (!n_n4273)) + ((n_n4371) & (!n_n3533) & (n_n1308) & (!n_n4370) & (n_n4273)) + ((n_n4371) & (!n_n3533) & (n_n1308) & (n_n4370) & (!n_n4273)) + ((n_n4371) & (!n_n3533) & (n_n1308) & (n_n4370) & (n_n4273)) + ((n_n4371) & (n_n3533) & (!n_n1308) & (!n_n4370) & (!n_n4273)) + ((n_n4371) & (n_n3533) & (!n_n1308) & (!n_n4370) & (n_n4273)) + ((n_n4371) & (n_n3533) & (!n_n1308) & (n_n4370) & (!n_n4273)) + ((n_n4371) & (n_n3533) & (!n_n1308) & (n_n4370) & (n_n4273)) + ((n_n4371) & (n_n3533) & (n_n1308) & (!n_n4370) & (!n_n4273)) + ((n_n4371) & (n_n3533) & (n_n1308) & (!n_n4370) & (n_n4273)) + ((n_n4371) & (n_n3533) & (n_n1308) & (n_n4370) & (!n_n4273)) + ((n_n4371) & (n_n3533) & (n_n1308) & (n_n4370) & (n_n4273)));
	assign x14159x = (((!n_n4382) & (!n_n4383) & (!n_n4380) & (n_n4372)) + ((!n_n4382) & (!n_n4383) & (n_n4380) & (!n_n4372)) + ((!n_n4382) & (!n_n4383) & (n_n4380) & (n_n4372)) + ((!n_n4382) & (n_n4383) & (!n_n4380) & (!n_n4372)) + ((!n_n4382) & (n_n4383) & (!n_n4380) & (n_n4372)) + ((!n_n4382) & (n_n4383) & (n_n4380) & (!n_n4372)) + ((!n_n4382) & (n_n4383) & (n_n4380) & (n_n4372)) + ((n_n4382) & (!n_n4383) & (!n_n4380) & (!n_n4372)) + ((n_n4382) & (!n_n4383) & (!n_n4380) & (n_n4372)) + ((n_n4382) & (!n_n4383) & (n_n4380) & (!n_n4372)) + ((n_n4382) & (!n_n4383) & (n_n4380) & (n_n4372)) + ((n_n4382) & (n_n4383) & (!n_n4380) & (!n_n4372)) + ((n_n4382) & (n_n4383) & (!n_n4380) & (n_n4372)) + ((n_n4382) & (n_n4383) & (n_n4380) & (!n_n4372)) + ((n_n4382) & (n_n4383) & (n_n4380) & (n_n4372)));
	assign n_n3288 = (((!n_n4368) & (!n_n3367) & (!x301x) & (!x14163x) & (x14159x)) + ((!n_n4368) & (!n_n3367) & (!x301x) & (x14163x) & (!x14159x)) + ((!n_n4368) & (!n_n3367) & (!x301x) & (x14163x) & (x14159x)) + ((!n_n4368) & (!n_n3367) & (x301x) & (!x14163x) & (!x14159x)) + ((!n_n4368) & (!n_n3367) & (x301x) & (!x14163x) & (x14159x)) + ((!n_n4368) & (!n_n3367) & (x301x) & (x14163x) & (!x14159x)) + ((!n_n4368) & (!n_n3367) & (x301x) & (x14163x) & (x14159x)) + ((!n_n4368) & (n_n3367) & (!x301x) & (!x14163x) & (!x14159x)) + ((!n_n4368) & (n_n3367) & (!x301x) & (!x14163x) & (x14159x)) + ((!n_n4368) & (n_n3367) & (!x301x) & (x14163x) & (!x14159x)) + ((!n_n4368) & (n_n3367) & (!x301x) & (x14163x) & (x14159x)) + ((!n_n4368) & (n_n3367) & (x301x) & (!x14163x) & (!x14159x)) + ((!n_n4368) & (n_n3367) & (x301x) & (!x14163x) & (x14159x)) + ((!n_n4368) & (n_n3367) & (x301x) & (x14163x) & (!x14159x)) + ((!n_n4368) & (n_n3367) & (x301x) & (x14163x) & (x14159x)) + ((n_n4368) & (!n_n3367) & (!x301x) & (!x14163x) & (!x14159x)) + ((n_n4368) & (!n_n3367) & (!x301x) & (!x14163x) & (x14159x)) + ((n_n4368) & (!n_n3367) & (!x301x) & (x14163x) & (!x14159x)) + ((n_n4368) & (!n_n3367) & (!x301x) & (x14163x) & (x14159x)) + ((n_n4368) & (!n_n3367) & (x301x) & (!x14163x) & (!x14159x)) + ((n_n4368) & (!n_n3367) & (x301x) & (!x14163x) & (x14159x)) + ((n_n4368) & (!n_n3367) & (x301x) & (x14163x) & (!x14159x)) + ((n_n4368) & (!n_n3367) & (x301x) & (x14163x) & (x14159x)) + ((n_n4368) & (n_n3367) & (!x301x) & (!x14163x) & (!x14159x)) + ((n_n4368) & (n_n3367) & (!x301x) & (!x14163x) & (x14159x)) + ((n_n4368) & (n_n3367) & (!x301x) & (x14163x) & (!x14159x)) + ((n_n4368) & (n_n3367) & (!x301x) & (x14163x) & (x14159x)) + ((n_n4368) & (n_n3367) & (x301x) & (!x14163x) & (!x14159x)) + ((n_n4368) & (n_n3367) & (x301x) & (!x14163x) & (x14159x)) + ((n_n4368) & (n_n3367) & (x301x) & (x14163x) & (!x14159x)) + ((n_n4368) & (n_n3367) & (x301x) & (x14163x) & (x14159x)));
	assign x14170x = (((!n_n4407) & (!n_n4404) & (!n_n4405) & (!n_n4406) & (n_n4398)) + ((!n_n4407) & (!n_n4404) & (!n_n4405) & (n_n4406) & (!n_n4398)) + ((!n_n4407) & (!n_n4404) & (!n_n4405) & (n_n4406) & (n_n4398)) + ((!n_n4407) & (!n_n4404) & (n_n4405) & (!n_n4406) & (!n_n4398)) + ((!n_n4407) & (!n_n4404) & (n_n4405) & (!n_n4406) & (n_n4398)) + ((!n_n4407) & (!n_n4404) & (n_n4405) & (n_n4406) & (!n_n4398)) + ((!n_n4407) & (!n_n4404) & (n_n4405) & (n_n4406) & (n_n4398)) + ((!n_n4407) & (n_n4404) & (!n_n4405) & (!n_n4406) & (!n_n4398)) + ((!n_n4407) & (n_n4404) & (!n_n4405) & (!n_n4406) & (n_n4398)) + ((!n_n4407) & (n_n4404) & (!n_n4405) & (n_n4406) & (!n_n4398)) + ((!n_n4407) & (n_n4404) & (!n_n4405) & (n_n4406) & (n_n4398)) + ((!n_n4407) & (n_n4404) & (n_n4405) & (!n_n4406) & (!n_n4398)) + ((!n_n4407) & (n_n4404) & (n_n4405) & (!n_n4406) & (n_n4398)) + ((!n_n4407) & (n_n4404) & (n_n4405) & (n_n4406) & (!n_n4398)) + ((!n_n4407) & (n_n4404) & (n_n4405) & (n_n4406) & (n_n4398)) + ((n_n4407) & (!n_n4404) & (!n_n4405) & (!n_n4406) & (!n_n4398)) + ((n_n4407) & (!n_n4404) & (!n_n4405) & (!n_n4406) & (n_n4398)) + ((n_n4407) & (!n_n4404) & (!n_n4405) & (n_n4406) & (!n_n4398)) + ((n_n4407) & (!n_n4404) & (!n_n4405) & (n_n4406) & (n_n4398)) + ((n_n4407) & (!n_n4404) & (n_n4405) & (!n_n4406) & (!n_n4398)) + ((n_n4407) & (!n_n4404) & (n_n4405) & (!n_n4406) & (n_n4398)) + ((n_n4407) & (!n_n4404) & (n_n4405) & (n_n4406) & (!n_n4398)) + ((n_n4407) & (!n_n4404) & (n_n4405) & (n_n4406) & (n_n4398)) + ((n_n4407) & (n_n4404) & (!n_n4405) & (!n_n4406) & (!n_n4398)) + ((n_n4407) & (n_n4404) & (!n_n4405) & (!n_n4406) & (n_n4398)) + ((n_n4407) & (n_n4404) & (!n_n4405) & (n_n4406) & (!n_n4398)) + ((n_n4407) & (n_n4404) & (!n_n4405) & (n_n4406) & (n_n4398)) + ((n_n4407) & (n_n4404) & (n_n4405) & (!n_n4406) & (!n_n4398)) + ((n_n4407) & (n_n4404) & (n_n4405) & (!n_n4406) & (n_n4398)) + ((n_n4407) & (n_n4404) & (n_n4405) & (n_n4406) & (!n_n4398)) + ((n_n4407) & (n_n4404) & (n_n4405) & (n_n4406) & (n_n4398)));
	assign n_n3363 = (((!n_n4403) & (!n_n4400) & (!n_n4396) & (!n_n4399) & (x14170x)) + ((!n_n4403) & (!n_n4400) & (!n_n4396) & (n_n4399) & (!x14170x)) + ((!n_n4403) & (!n_n4400) & (!n_n4396) & (n_n4399) & (x14170x)) + ((!n_n4403) & (!n_n4400) & (n_n4396) & (!n_n4399) & (!x14170x)) + ((!n_n4403) & (!n_n4400) & (n_n4396) & (!n_n4399) & (x14170x)) + ((!n_n4403) & (!n_n4400) & (n_n4396) & (n_n4399) & (!x14170x)) + ((!n_n4403) & (!n_n4400) & (n_n4396) & (n_n4399) & (x14170x)) + ((!n_n4403) & (n_n4400) & (!n_n4396) & (!n_n4399) & (!x14170x)) + ((!n_n4403) & (n_n4400) & (!n_n4396) & (!n_n4399) & (x14170x)) + ((!n_n4403) & (n_n4400) & (!n_n4396) & (n_n4399) & (!x14170x)) + ((!n_n4403) & (n_n4400) & (!n_n4396) & (n_n4399) & (x14170x)) + ((!n_n4403) & (n_n4400) & (n_n4396) & (!n_n4399) & (!x14170x)) + ((!n_n4403) & (n_n4400) & (n_n4396) & (!n_n4399) & (x14170x)) + ((!n_n4403) & (n_n4400) & (n_n4396) & (n_n4399) & (!x14170x)) + ((!n_n4403) & (n_n4400) & (n_n4396) & (n_n4399) & (x14170x)) + ((n_n4403) & (!n_n4400) & (!n_n4396) & (!n_n4399) & (!x14170x)) + ((n_n4403) & (!n_n4400) & (!n_n4396) & (!n_n4399) & (x14170x)) + ((n_n4403) & (!n_n4400) & (!n_n4396) & (n_n4399) & (!x14170x)) + ((n_n4403) & (!n_n4400) & (!n_n4396) & (n_n4399) & (x14170x)) + ((n_n4403) & (!n_n4400) & (n_n4396) & (!n_n4399) & (!x14170x)) + ((n_n4403) & (!n_n4400) & (n_n4396) & (!n_n4399) & (x14170x)) + ((n_n4403) & (!n_n4400) & (n_n4396) & (n_n4399) & (!x14170x)) + ((n_n4403) & (!n_n4400) & (n_n4396) & (n_n4399) & (x14170x)) + ((n_n4403) & (n_n4400) & (!n_n4396) & (!n_n4399) & (!x14170x)) + ((n_n4403) & (n_n4400) & (!n_n4396) & (!n_n4399) & (x14170x)) + ((n_n4403) & (n_n4400) & (!n_n4396) & (n_n4399) & (!x14170x)) + ((n_n4403) & (n_n4400) & (!n_n4396) & (n_n4399) & (x14170x)) + ((n_n4403) & (n_n4400) & (n_n4396) & (!n_n4399) & (!x14170x)) + ((n_n4403) & (n_n4400) & (n_n4396) & (!n_n4399) & (x14170x)) + ((n_n4403) & (n_n4400) & (n_n4396) & (n_n4399) & (!x14170x)) + ((n_n4403) & (n_n4400) & (n_n4396) & (n_n4399) & (x14170x)));
	assign x14175x = (((!n_n4415) & (!n_n4408) & (!n_n4414) & (!n_n4411) & (n_n4412)) + ((!n_n4415) & (!n_n4408) & (!n_n4414) & (n_n4411) & (!n_n4412)) + ((!n_n4415) & (!n_n4408) & (!n_n4414) & (n_n4411) & (n_n4412)) + ((!n_n4415) & (!n_n4408) & (n_n4414) & (!n_n4411) & (!n_n4412)) + ((!n_n4415) & (!n_n4408) & (n_n4414) & (!n_n4411) & (n_n4412)) + ((!n_n4415) & (!n_n4408) & (n_n4414) & (n_n4411) & (!n_n4412)) + ((!n_n4415) & (!n_n4408) & (n_n4414) & (n_n4411) & (n_n4412)) + ((!n_n4415) & (n_n4408) & (!n_n4414) & (!n_n4411) & (!n_n4412)) + ((!n_n4415) & (n_n4408) & (!n_n4414) & (!n_n4411) & (n_n4412)) + ((!n_n4415) & (n_n4408) & (!n_n4414) & (n_n4411) & (!n_n4412)) + ((!n_n4415) & (n_n4408) & (!n_n4414) & (n_n4411) & (n_n4412)) + ((!n_n4415) & (n_n4408) & (n_n4414) & (!n_n4411) & (!n_n4412)) + ((!n_n4415) & (n_n4408) & (n_n4414) & (!n_n4411) & (n_n4412)) + ((!n_n4415) & (n_n4408) & (n_n4414) & (n_n4411) & (!n_n4412)) + ((!n_n4415) & (n_n4408) & (n_n4414) & (n_n4411) & (n_n4412)) + ((n_n4415) & (!n_n4408) & (!n_n4414) & (!n_n4411) & (!n_n4412)) + ((n_n4415) & (!n_n4408) & (!n_n4414) & (!n_n4411) & (n_n4412)) + ((n_n4415) & (!n_n4408) & (!n_n4414) & (n_n4411) & (!n_n4412)) + ((n_n4415) & (!n_n4408) & (!n_n4414) & (n_n4411) & (n_n4412)) + ((n_n4415) & (!n_n4408) & (n_n4414) & (!n_n4411) & (!n_n4412)) + ((n_n4415) & (!n_n4408) & (n_n4414) & (!n_n4411) & (n_n4412)) + ((n_n4415) & (!n_n4408) & (n_n4414) & (n_n4411) & (!n_n4412)) + ((n_n4415) & (!n_n4408) & (n_n4414) & (n_n4411) & (n_n4412)) + ((n_n4415) & (n_n4408) & (!n_n4414) & (!n_n4411) & (!n_n4412)) + ((n_n4415) & (n_n4408) & (!n_n4414) & (!n_n4411) & (n_n4412)) + ((n_n4415) & (n_n4408) & (!n_n4414) & (n_n4411) & (!n_n4412)) + ((n_n4415) & (n_n4408) & (!n_n4414) & (n_n4411) & (n_n4412)) + ((n_n4415) & (n_n4408) & (n_n4414) & (!n_n4411) & (!n_n4412)) + ((n_n4415) & (n_n4408) & (n_n4414) & (!n_n4411) & (n_n4412)) + ((n_n4415) & (n_n4408) & (n_n4414) & (n_n4411) & (!n_n4412)) + ((n_n4415) & (n_n4408) & (n_n4414) & (n_n4411) & (n_n4412)));
	assign x79x = (((!i_9_) & (n_n536) & (n_n524) & (n_n473)) + ((i_9_) & (n_n536) & (n_n524) & (n_n473)));
	assign n_n3362 = (((!n_n4413) & (!n_n4417) & (!x14175x) & (x79x)) + ((!n_n4413) & (!n_n4417) & (x14175x) & (!x79x)) + ((!n_n4413) & (!n_n4417) & (x14175x) & (x79x)) + ((!n_n4413) & (n_n4417) & (!x14175x) & (!x79x)) + ((!n_n4413) & (n_n4417) & (!x14175x) & (x79x)) + ((!n_n4413) & (n_n4417) & (x14175x) & (!x79x)) + ((!n_n4413) & (n_n4417) & (x14175x) & (x79x)) + ((n_n4413) & (!n_n4417) & (!x14175x) & (!x79x)) + ((n_n4413) & (!n_n4417) & (!x14175x) & (x79x)) + ((n_n4413) & (!n_n4417) & (x14175x) & (!x79x)) + ((n_n4413) & (!n_n4417) & (x14175x) & (x79x)) + ((n_n4413) & (n_n4417) & (!x14175x) & (!x79x)) + ((n_n4413) & (n_n4417) & (!x14175x) & (x79x)) + ((n_n4413) & (n_n4417) & (x14175x) & (!x79x)) + ((n_n4413) & (n_n4417) & (x14175x) & (x79x)));
	assign x14179x = (((!i_9_) & (!n_n536) & (!n_n482) & (!n_n532) & (n_n2435)) + ((!i_9_) & (!n_n536) & (!n_n482) & (n_n532) & (n_n2435)) + ((!i_9_) & (!n_n536) & (n_n482) & (!n_n532) & (n_n2435)) + ((!i_9_) & (!n_n536) & (n_n482) & (n_n532) & (n_n2435)) + ((!i_9_) & (n_n536) & (!n_n482) & (!n_n532) & (n_n2435)) + ((!i_9_) & (n_n536) & (!n_n482) & (n_n532) & (n_n2435)) + ((!i_9_) & (n_n536) & (n_n482) & (!n_n532) & (n_n2435)) + ((!i_9_) & (n_n536) & (n_n482) & (n_n532) & (!n_n2435)) + ((!i_9_) & (n_n536) & (n_n482) & (n_n532) & (n_n2435)) + ((i_9_) & (!n_n536) & (!n_n482) & (!n_n532) & (n_n2435)) + ((i_9_) & (!n_n536) & (!n_n482) & (n_n532) & (n_n2435)) + ((i_9_) & (!n_n536) & (n_n482) & (!n_n532) & (n_n2435)) + ((i_9_) & (!n_n536) & (n_n482) & (n_n532) & (n_n2435)) + ((i_9_) & (n_n536) & (!n_n482) & (!n_n532) & (n_n2435)) + ((i_9_) & (n_n536) & (!n_n482) & (n_n532) & (n_n2435)) + ((i_9_) & (n_n536) & (n_n482) & (!n_n532) & (n_n2435)) + ((i_9_) & (n_n536) & (n_n482) & (n_n532) & (!n_n2435)) + ((i_9_) & (n_n536) & (n_n482) & (n_n532) & (n_n2435)));
	assign x14180x = (((!n_n4392) & (!n_n4384) & (!n_n4386) & (!n_n4387) & (x14179x)) + ((!n_n4392) & (!n_n4384) & (!n_n4386) & (n_n4387) & (!x14179x)) + ((!n_n4392) & (!n_n4384) & (!n_n4386) & (n_n4387) & (x14179x)) + ((!n_n4392) & (!n_n4384) & (n_n4386) & (!n_n4387) & (!x14179x)) + ((!n_n4392) & (!n_n4384) & (n_n4386) & (!n_n4387) & (x14179x)) + ((!n_n4392) & (!n_n4384) & (n_n4386) & (n_n4387) & (!x14179x)) + ((!n_n4392) & (!n_n4384) & (n_n4386) & (n_n4387) & (x14179x)) + ((!n_n4392) & (n_n4384) & (!n_n4386) & (!n_n4387) & (!x14179x)) + ((!n_n4392) & (n_n4384) & (!n_n4386) & (!n_n4387) & (x14179x)) + ((!n_n4392) & (n_n4384) & (!n_n4386) & (n_n4387) & (!x14179x)) + ((!n_n4392) & (n_n4384) & (!n_n4386) & (n_n4387) & (x14179x)) + ((!n_n4392) & (n_n4384) & (n_n4386) & (!n_n4387) & (!x14179x)) + ((!n_n4392) & (n_n4384) & (n_n4386) & (!n_n4387) & (x14179x)) + ((!n_n4392) & (n_n4384) & (n_n4386) & (n_n4387) & (!x14179x)) + ((!n_n4392) & (n_n4384) & (n_n4386) & (n_n4387) & (x14179x)) + ((n_n4392) & (!n_n4384) & (!n_n4386) & (!n_n4387) & (!x14179x)) + ((n_n4392) & (!n_n4384) & (!n_n4386) & (!n_n4387) & (x14179x)) + ((n_n4392) & (!n_n4384) & (!n_n4386) & (n_n4387) & (!x14179x)) + ((n_n4392) & (!n_n4384) & (!n_n4386) & (n_n4387) & (x14179x)) + ((n_n4392) & (!n_n4384) & (n_n4386) & (!n_n4387) & (!x14179x)) + ((n_n4392) & (!n_n4384) & (n_n4386) & (!n_n4387) & (x14179x)) + ((n_n4392) & (!n_n4384) & (n_n4386) & (n_n4387) & (!x14179x)) + ((n_n4392) & (!n_n4384) & (n_n4386) & (n_n4387) & (x14179x)) + ((n_n4392) & (n_n4384) & (!n_n4386) & (!n_n4387) & (!x14179x)) + ((n_n4392) & (n_n4384) & (!n_n4386) & (!n_n4387) & (x14179x)) + ((n_n4392) & (n_n4384) & (!n_n4386) & (n_n4387) & (!x14179x)) + ((n_n4392) & (n_n4384) & (!n_n4386) & (n_n4387) & (x14179x)) + ((n_n4392) & (n_n4384) & (n_n4386) & (!n_n4387) & (!x14179x)) + ((n_n4392) & (n_n4384) & (n_n4386) & (!n_n4387) & (x14179x)) + ((n_n4392) & (n_n4384) & (n_n4386) & (n_n4387) & (!x14179x)) + ((n_n4392) & (n_n4384) & (n_n4386) & (n_n4387) & (x14179x)));
	assign n_n3287 = (((!n_n3363) & (!n_n3362) & (x14180x)) + ((!n_n3363) & (n_n3362) & (!x14180x)) + ((!n_n3363) & (n_n3362) & (x14180x)) + ((n_n3363) & (!n_n3362) & (!x14180x)) + ((n_n3363) & (!n_n3362) & (x14180x)) + ((n_n3363) & (n_n3362) & (!x14180x)) + ((n_n3363) & (n_n3362) & (x14180x)));
	assign n_n4279 = (((!i_9_) & (n_n536) & (n_n518) & (!n_n532) & (n_n534)) + ((!i_9_) & (n_n536) & (n_n518) & (n_n532) & (n_n534)) + ((i_9_) & (n_n536) & (n_n518) & (!n_n532) & (n_n534)) + ((i_9_) & (n_n536) & (n_n518) & (n_n532) & (!n_n534)) + ((i_9_) & (n_n536) & (n_n518) & (n_n532) & (n_n534)));
	assign x106x = (((n_n536) & (n_n535) & (!x20x) & (x23x)) + ((n_n536) & (n_n535) & (x20x) & (!x23x)) + ((n_n536) & (n_n535) & (x20x) & (x23x)));
	assign n_n3369 = (((!n_n4324) & (!x198x) & (!n_n4335) & (!n_n4279) & (x106x)) + ((!n_n4324) & (!x198x) & (!n_n4335) & (n_n4279) & (!x106x)) + ((!n_n4324) & (!x198x) & (!n_n4335) & (n_n4279) & (x106x)) + ((!n_n4324) & (!x198x) & (n_n4335) & (!n_n4279) & (!x106x)) + ((!n_n4324) & (!x198x) & (n_n4335) & (!n_n4279) & (x106x)) + ((!n_n4324) & (!x198x) & (n_n4335) & (n_n4279) & (!x106x)) + ((!n_n4324) & (!x198x) & (n_n4335) & (n_n4279) & (x106x)) + ((!n_n4324) & (x198x) & (!n_n4335) & (!n_n4279) & (!x106x)) + ((!n_n4324) & (x198x) & (!n_n4335) & (!n_n4279) & (x106x)) + ((!n_n4324) & (x198x) & (!n_n4335) & (n_n4279) & (!x106x)) + ((!n_n4324) & (x198x) & (!n_n4335) & (n_n4279) & (x106x)) + ((!n_n4324) & (x198x) & (n_n4335) & (!n_n4279) & (!x106x)) + ((!n_n4324) & (x198x) & (n_n4335) & (!n_n4279) & (x106x)) + ((!n_n4324) & (x198x) & (n_n4335) & (n_n4279) & (!x106x)) + ((!n_n4324) & (x198x) & (n_n4335) & (n_n4279) & (x106x)) + ((n_n4324) & (!x198x) & (!n_n4335) & (!n_n4279) & (!x106x)) + ((n_n4324) & (!x198x) & (!n_n4335) & (!n_n4279) & (x106x)) + ((n_n4324) & (!x198x) & (!n_n4335) & (n_n4279) & (!x106x)) + ((n_n4324) & (!x198x) & (!n_n4335) & (n_n4279) & (x106x)) + ((n_n4324) & (!x198x) & (n_n4335) & (!n_n4279) & (!x106x)) + ((n_n4324) & (!x198x) & (n_n4335) & (!n_n4279) & (x106x)) + ((n_n4324) & (!x198x) & (n_n4335) & (n_n4279) & (!x106x)) + ((n_n4324) & (!x198x) & (n_n4335) & (n_n4279) & (x106x)) + ((n_n4324) & (x198x) & (!n_n4335) & (!n_n4279) & (!x106x)) + ((n_n4324) & (x198x) & (!n_n4335) & (!n_n4279) & (x106x)) + ((n_n4324) & (x198x) & (!n_n4335) & (n_n4279) & (!x106x)) + ((n_n4324) & (x198x) & (!n_n4335) & (n_n4279) & (x106x)) + ((n_n4324) & (x198x) & (n_n4335) & (!n_n4279) & (!x106x)) + ((n_n4324) & (x198x) & (n_n4335) & (!n_n4279) & (x106x)) + ((n_n4324) & (x198x) & (n_n4335) & (n_n4279) & (!x106x)) + ((n_n4324) & (x198x) & (n_n4335) & (n_n4279) & (x106x)));
	assign x14186x = (((!i_9_) & (n_n536) & (!n_n532) & (n_n535) & (n_n530)) + ((!i_9_) & (n_n536) & (n_n532) & (n_n535) & (!n_n530)) + ((!i_9_) & (n_n536) & (n_n532) & (n_n535) & (n_n530)) + ((i_9_) & (n_n536) & (!n_n532) & (n_n535) & (n_n530)) + ((i_9_) & (n_n536) & (n_n532) & (n_n535) & (n_n530)));
	assign x363x = (((!n_n4318) & (!n_n4321) & (!n_n4322) & (n_n4323)) + ((!n_n4318) & (!n_n4321) & (n_n4322) & (!n_n4323)) + ((!n_n4318) & (!n_n4321) & (n_n4322) & (n_n4323)) + ((!n_n4318) & (n_n4321) & (!n_n4322) & (!n_n4323)) + ((!n_n4318) & (n_n4321) & (!n_n4322) & (n_n4323)) + ((!n_n4318) & (n_n4321) & (n_n4322) & (!n_n4323)) + ((!n_n4318) & (n_n4321) & (n_n4322) & (n_n4323)) + ((n_n4318) & (!n_n4321) & (!n_n4322) & (!n_n4323)) + ((n_n4318) & (!n_n4321) & (!n_n4322) & (n_n4323)) + ((n_n4318) & (!n_n4321) & (n_n4322) & (!n_n4323)) + ((n_n4318) & (!n_n4321) & (n_n4322) & (n_n4323)) + ((n_n4318) & (n_n4321) & (!n_n4322) & (!n_n4323)) + ((n_n4318) & (n_n4321) & (!n_n4322) & (n_n4323)) + ((n_n4318) & (n_n4321) & (n_n4322) & (!n_n4323)) + ((n_n4318) & (n_n4321) & (n_n4322) & (n_n4323)));
	assign n_n3370 = (((!n_n4319) & (!n_n4320) & (!x14186x) & (x363x)) + ((!n_n4319) & (!n_n4320) & (x14186x) & (!x363x)) + ((!n_n4319) & (!n_n4320) & (x14186x) & (x363x)) + ((!n_n4319) & (n_n4320) & (!x14186x) & (!x363x)) + ((!n_n4319) & (n_n4320) & (!x14186x) & (x363x)) + ((!n_n4319) & (n_n4320) & (x14186x) & (!x363x)) + ((!n_n4319) & (n_n4320) & (x14186x) & (x363x)) + ((n_n4319) & (!n_n4320) & (!x14186x) & (!x363x)) + ((n_n4319) & (!n_n4320) & (!x14186x) & (x363x)) + ((n_n4319) & (!n_n4320) & (x14186x) & (!x363x)) + ((n_n4319) & (!n_n4320) & (x14186x) & (x363x)) + ((n_n4319) & (n_n4320) & (!x14186x) & (!x363x)) + ((n_n4319) & (n_n4320) & (!x14186x) & (x363x)) + ((n_n4319) & (n_n4320) & (x14186x) & (!x363x)) + ((n_n4319) & (n_n4320) & (x14186x) & (x363x)));
	assign x156x = (((!i_9_) & (n_n536) & (n_n518) & (!n_n520) & (x23x)) + ((!i_9_) & (n_n536) & (n_n518) & (n_n520) & (x23x)) + ((i_9_) & (n_n536) & (n_n518) & (!n_n520) & (x23x)) + ((i_9_) & (n_n536) & (n_n518) & (n_n520) & (!x23x)) + ((i_9_) & (n_n536) & (n_n518) & (n_n520) & (x23x)));
	assign x14193x = (((!n_n4343) & (!n_n4342) & (!x67x) & (!n_n4348) & (!x22112x)) + ((!n_n4343) & (!n_n4342) & (!x67x) & (n_n4348) & (!x22112x)) + ((!n_n4343) & (!n_n4342) & (!x67x) & (n_n4348) & (x22112x)) + ((!n_n4343) & (!n_n4342) & (x67x) & (!n_n4348) & (!x22112x)) + ((!n_n4343) & (!n_n4342) & (x67x) & (!n_n4348) & (x22112x)) + ((!n_n4343) & (!n_n4342) & (x67x) & (n_n4348) & (!x22112x)) + ((!n_n4343) & (!n_n4342) & (x67x) & (n_n4348) & (x22112x)) + ((!n_n4343) & (n_n4342) & (!x67x) & (!n_n4348) & (!x22112x)) + ((!n_n4343) & (n_n4342) & (!x67x) & (!n_n4348) & (x22112x)) + ((!n_n4343) & (n_n4342) & (!x67x) & (n_n4348) & (!x22112x)) + ((!n_n4343) & (n_n4342) & (!x67x) & (n_n4348) & (x22112x)) + ((!n_n4343) & (n_n4342) & (x67x) & (!n_n4348) & (!x22112x)) + ((!n_n4343) & (n_n4342) & (x67x) & (!n_n4348) & (x22112x)) + ((!n_n4343) & (n_n4342) & (x67x) & (n_n4348) & (!x22112x)) + ((!n_n4343) & (n_n4342) & (x67x) & (n_n4348) & (x22112x)) + ((n_n4343) & (!n_n4342) & (!x67x) & (!n_n4348) & (!x22112x)) + ((n_n4343) & (!n_n4342) & (!x67x) & (!n_n4348) & (x22112x)) + ((n_n4343) & (!n_n4342) & (!x67x) & (n_n4348) & (!x22112x)) + ((n_n4343) & (!n_n4342) & (!x67x) & (n_n4348) & (x22112x)) + ((n_n4343) & (!n_n4342) & (x67x) & (!n_n4348) & (!x22112x)) + ((n_n4343) & (!n_n4342) & (x67x) & (!n_n4348) & (x22112x)) + ((n_n4343) & (!n_n4342) & (x67x) & (n_n4348) & (!x22112x)) + ((n_n4343) & (!n_n4342) & (x67x) & (n_n4348) & (x22112x)) + ((n_n4343) & (n_n4342) & (!x67x) & (!n_n4348) & (!x22112x)) + ((n_n4343) & (n_n4342) & (!x67x) & (!n_n4348) & (x22112x)) + ((n_n4343) & (n_n4342) & (!x67x) & (n_n4348) & (!x22112x)) + ((n_n4343) & (n_n4342) & (!x67x) & (n_n4348) & (x22112x)) + ((n_n4343) & (n_n4342) & (x67x) & (!n_n4348) & (!x22112x)) + ((n_n4343) & (n_n4342) & (x67x) & (!n_n4348) & (x22112x)) + ((n_n4343) & (n_n4342) & (x67x) & (n_n4348) & (!x22112x)) + ((n_n4343) & (n_n4342) & (x67x) & (n_n4348) & (x22112x)));
	assign n_n3262 = (((!n_n3288) & (!n_n3287) & (!n_n3369) & (!n_n3370) & (x14193x)) + ((!n_n3288) & (!n_n3287) & (!n_n3369) & (n_n3370) & (!x14193x)) + ((!n_n3288) & (!n_n3287) & (!n_n3369) & (n_n3370) & (x14193x)) + ((!n_n3288) & (!n_n3287) & (n_n3369) & (!n_n3370) & (!x14193x)) + ((!n_n3288) & (!n_n3287) & (n_n3369) & (!n_n3370) & (x14193x)) + ((!n_n3288) & (!n_n3287) & (n_n3369) & (n_n3370) & (!x14193x)) + ((!n_n3288) & (!n_n3287) & (n_n3369) & (n_n3370) & (x14193x)) + ((!n_n3288) & (n_n3287) & (!n_n3369) & (!n_n3370) & (!x14193x)) + ((!n_n3288) & (n_n3287) & (!n_n3369) & (!n_n3370) & (x14193x)) + ((!n_n3288) & (n_n3287) & (!n_n3369) & (n_n3370) & (!x14193x)) + ((!n_n3288) & (n_n3287) & (!n_n3369) & (n_n3370) & (x14193x)) + ((!n_n3288) & (n_n3287) & (n_n3369) & (!n_n3370) & (!x14193x)) + ((!n_n3288) & (n_n3287) & (n_n3369) & (!n_n3370) & (x14193x)) + ((!n_n3288) & (n_n3287) & (n_n3369) & (n_n3370) & (!x14193x)) + ((!n_n3288) & (n_n3287) & (n_n3369) & (n_n3370) & (x14193x)) + ((n_n3288) & (!n_n3287) & (!n_n3369) & (!n_n3370) & (!x14193x)) + ((n_n3288) & (!n_n3287) & (!n_n3369) & (!n_n3370) & (x14193x)) + ((n_n3288) & (!n_n3287) & (!n_n3369) & (n_n3370) & (!x14193x)) + ((n_n3288) & (!n_n3287) & (!n_n3369) & (n_n3370) & (x14193x)) + ((n_n3288) & (!n_n3287) & (n_n3369) & (!n_n3370) & (!x14193x)) + ((n_n3288) & (!n_n3287) & (n_n3369) & (!n_n3370) & (x14193x)) + ((n_n3288) & (!n_n3287) & (n_n3369) & (n_n3370) & (!x14193x)) + ((n_n3288) & (!n_n3287) & (n_n3369) & (n_n3370) & (x14193x)) + ((n_n3288) & (n_n3287) & (!n_n3369) & (!n_n3370) & (!x14193x)) + ((n_n3288) & (n_n3287) & (!n_n3369) & (!n_n3370) & (x14193x)) + ((n_n3288) & (n_n3287) & (!n_n3369) & (n_n3370) & (!x14193x)) + ((n_n3288) & (n_n3287) & (!n_n3369) & (n_n3370) & (x14193x)) + ((n_n3288) & (n_n3287) & (n_n3369) & (!n_n3370) & (!x14193x)) + ((n_n3288) & (n_n3287) & (n_n3369) & (!n_n3370) & (x14193x)) + ((n_n3288) & (n_n3287) & (n_n3369) & (n_n3370) & (!x14193x)) + ((n_n3288) & (n_n3287) & (n_n3369) & (n_n3370) & (x14193x)));
	assign n_n4896 = (((i_9_) & (n_n526) & (n_n260) & (n_n491)));
	assign n_n4328 = (((i_9_) & (n_n536) & (n_n518) & (n_n534)));
	assign n_n4585 = (((!i_9_) & (n_n518) & (n_n390) & (n_n534)));
	assign x15489x = (((!x108x) & (!n_n4595) & (!n_n4592) & (n_n4603)) + ((!x108x) & (!n_n4595) & (n_n4592) & (!n_n4603)) + ((!x108x) & (!n_n4595) & (n_n4592) & (n_n4603)) + ((!x108x) & (n_n4595) & (!n_n4592) & (!n_n4603)) + ((!x108x) & (n_n4595) & (!n_n4592) & (n_n4603)) + ((!x108x) & (n_n4595) & (n_n4592) & (!n_n4603)) + ((!x108x) & (n_n4595) & (n_n4592) & (n_n4603)) + ((x108x) & (!n_n4595) & (!n_n4592) & (!n_n4603)) + ((x108x) & (!n_n4595) & (!n_n4592) & (n_n4603)) + ((x108x) & (!n_n4595) & (n_n4592) & (!n_n4603)) + ((x108x) & (!n_n4595) & (n_n4592) & (n_n4603)) + ((x108x) & (n_n4595) & (!n_n4592) & (!n_n4603)) + ((x108x) & (n_n4595) & (!n_n4592) & (n_n4603)) + ((x108x) & (n_n4595) & (n_n4592) & (!n_n4603)) + ((x108x) & (n_n4595) & (n_n4592) & (n_n4603)));
	assign x15602x = (((!n_n5050) & (!n_n5054) & (!n_n5046) & (n_n5049)) + ((!n_n5050) & (!n_n5054) & (n_n5046) & (!n_n5049)) + ((!n_n5050) & (!n_n5054) & (n_n5046) & (n_n5049)) + ((!n_n5050) & (n_n5054) & (!n_n5046) & (!n_n5049)) + ((!n_n5050) & (n_n5054) & (!n_n5046) & (n_n5049)) + ((!n_n5050) & (n_n5054) & (n_n5046) & (!n_n5049)) + ((!n_n5050) & (n_n5054) & (n_n5046) & (n_n5049)) + ((n_n5050) & (!n_n5054) & (!n_n5046) & (!n_n5049)) + ((n_n5050) & (!n_n5054) & (!n_n5046) & (n_n5049)) + ((n_n5050) & (!n_n5054) & (n_n5046) & (!n_n5049)) + ((n_n5050) & (!n_n5054) & (n_n5046) & (n_n5049)) + ((n_n5050) & (n_n5054) & (!n_n5046) & (!n_n5049)) + ((n_n5050) & (n_n5054) & (!n_n5046) & (n_n5049)) + ((n_n5050) & (n_n5054) & (n_n5046) & (!n_n5049)) + ((n_n5050) & (n_n5054) & (n_n5046) & (n_n5049)));
	assign x15603x = (((!n_n5055) & (!n_n5056) & (!n_n5052) & (!n_n5047) & (n_n5051)) + ((!n_n5055) & (!n_n5056) & (!n_n5052) & (n_n5047) & (!n_n5051)) + ((!n_n5055) & (!n_n5056) & (!n_n5052) & (n_n5047) & (n_n5051)) + ((!n_n5055) & (!n_n5056) & (n_n5052) & (!n_n5047) & (!n_n5051)) + ((!n_n5055) & (!n_n5056) & (n_n5052) & (!n_n5047) & (n_n5051)) + ((!n_n5055) & (!n_n5056) & (n_n5052) & (n_n5047) & (!n_n5051)) + ((!n_n5055) & (!n_n5056) & (n_n5052) & (n_n5047) & (n_n5051)) + ((!n_n5055) & (n_n5056) & (!n_n5052) & (!n_n5047) & (!n_n5051)) + ((!n_n5055) & (n_n5056) & (!n_n5052) & (!n_n5047) & (n_n5051)) + ((!n_n5055) & (n_n5056) & (!n_n5052) & (n_n5047) & (!n_n5051)) + ((!n_n5055) & (n_n5056) & (!n_n5052) & (n_n5047) & (n_n5051)) + ((!n_n5055) & (n_n5056) & (n_n5052) & (!n_n5047) & (!n_n5051)) + ((!n_n5055) & (n_n5056) & (n_n5052) & (!n_n5047) & (n_n5051)) + ((!n_n5055) & (n_n5056) & (n_n5052) & (n_n5047) & (!n_n5051)) + ((!n_n5055) & (n_n5056) & (n_n5052) & (n_n5047) & (n_n5051)) + ((n_n5055) & (!n_n5056) & (!n_n5052) & (!n_n5047) & (!n_n5051)) + ((n_n5055) & (!n_n5056) & (!n_n5052) & (!n_n5047) & (n_n5051)) + ((n_n5055) & (!n_n5056) & (!n_n5052) & (n_n5047) & (!n_n5051)) + ((n_n5055) & (!n_n5056) & (!n_n5052) & (n_n5047) & (n_n5051)) + ((n_n5055) & (!n_n5056) & (n_n5052) & (!n_n5047) & (!n_n5051)) + ((n_n5055) & (!n_n5056) & (n_n5052) & (!n_n5047) & (n_n5051)) + ((n_n5055) & (!n_n5056) & (n_n5052) & (n_n5047) & (!n_n5051)) + ((n_n5055) & (!n_n5056) & (n_n5052) & (n_n5047) & (n_n5051)) + ((n_n5055) & (n_n5056) & (!n_n5052) & (!n_n5047) & (!n_n5051)) + ((n_n5055) & (n_n5056) & (!n_n5052) & (!n_n5047) & (n_n5051)) + ((n_n5055) & (n_n5056) & (!n_n5052) & (n_n5047) & (!n_n5051)) + ((n_n5055) & (n_n5056) & (!n_n5052) & (n_n5047) & (n_n5051)) + ((n_n5055) & (n_n5056) & (n_n5052) & (!n_n5047) & (!n_n5051)) + ((n_n5055) & (n_n5056) & (n_n5052) & (!n_n5047) & (n_n5051)) + ((n_n5055) & (n_n5056) & (n_n5052) & (n_n5047) & (!n_n5051)) + ((n_n5055) & (n_n5056) & (n_n5052) & (n_n5047) & (n_n5051)));
	assign n_n5235 = (((!i_9_) & (n_n524) & (n_n518) & (n_n65)));
	assign n_n5234 = (((i_7_) & (!i_8_) & (!i_6_) & (x19x) & (n_n518)));
	assign n_n5286 = (((i_5_) & (!i_3_) & (i_4_) & (x19x) & (n_n520)));
	assign x227x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n260) & (n_n491)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n260) & (n_n491)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n260) & (n_n491)) + ((i_9_) & (n_n524) & (n_n526) & (n_n260) & (n_n491)));
	assign n_n3810 = (((!i_9_) & (!n_n524) & (n_n526) & (n_n260) & (n_n491)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n260) & (n_n491)) + ((i_9_) & (!n_n524) & (n_n526) & (n_n260) & (n_n491)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n260) & (n_n491)) + ((i_9_) & (n_n524) & (n_n526) & (n_n260) & (n_n491)));
	assign x16447x = (((!i_9_) & (n_n482) & (!n_n528) & (n_n260) & (n_n530)) + ((!i_9_) & (n_n482) & (n_n528) & (n_n260) & (!n_n530)) + ((!i_9_) & (n_n482) & (n_n528) & (n_n260) & (n_n530)));
	assign n_n2304 = (((!x15x) & (!n_n130) & (!n_n500) & (!n_n5130) & (n_n5134)) + ((!x15x) & (!n_n130) & (!n_n500) & (n_n5130) & (!n_n5134)) + ((!x15x) & (!n_n130) & (!n_n500) & (n_n5130) & (n_n5134)) + ((!x15x) & (!n_n130) & (n_n500) & (!n_n5130) & (n_n5134)) + ((!x15x) & (!n_n130) & (n_n500) & (n_n5130) & (!n_n5134)) + ((!x15x) & (!n_n130) & (n_n500) & (n_n5130) & (n_n5134)) + ((!x15x) & (n_n130) & (!n_n500) & (!n_n5130) & (n_n5134)) + ((!x15x) & (n_n130) & (!n_n500) & (n_n5130) & (!n_n5134)) + ((!x15x) & (n_n130) & (!n_n500) & (n_n5130) & (n_n5134)) + ((!x15x) & (n_n130) & (n_n500) & (!n_n5130) & (n_n5134)) + ((!x15x) & (n_n130) & (n_n500) & (n_n5130) & (!n_n5134)) + ((!x15x) & (n_n130) & (n_n500) & (n_n5130) & (n_n5134)) + ((x15x) & (!n_n130) & (!n_n500) & (!n_n5130) & (n_n5134)) + ((x15x) & (!n_n130) & (!n_n500) & (n_n5130) & (!n_n5134)) + ((x15x) & (!n_n130) & (!n_n500) & (n_n5130) & (n_n5134)) + ((x15x) & (!n_n130) & (n_n500) & (!n_n5130) & (n_n5134)) + ((x15x) & (!n_n130) & (n_n500) & (n_n5130) & (!n_n5134)) + ((x15x) & (!n_n130) & (n_n500) & (n_n5130) & (n_n5134)) + ((x15x) & (n_n130) & (!n_n500) & (!n_n5130) & (n_n5134)) + ((x15x) & (n_n130) & (!n_n500) & (n_n5130) & (!n_n5134)) + ((x15x) & (n_n130) & (!n_n500) & (n_n5130) & (n_n5134)) + ((x15x) & (n_n130) & (n_n500) & (!n_n5130) & (!n_n5134)) + ((x15x) & (n_n130) & (n_n500) & (!n_n5130) & (n_n5134)) + ((x15x) & (n_n130) & (n_n500) & (n_n5130) & (!n_n5134)) + ((x15x) & (n_n130) & (n_n500) & (n_n5130) & (n_n5134)));
	assign n_n5253 = (((i_5_) & (i_3_) & (!i_4_) & (x20x) & (n_n65)));
	assign n_n1139 = (((!n_n509) & (!x20x) & (!x23x) & (!n_n65) & (n_n5256)) + ((!n_n509) & (!x20x) & (!x23x) & (n_n65) & (n_n5256)) + ((!n_n509) & (!x20x) & (x23x) & (!n_n65) & (n_n5256)) + ((!n_n509) & (!x20x) & (x23x) & (n_n65) & (n_n5256)) + ((!n_n509) & (x20x) & (!x23x) & (!n_n65) & (n_n5256)) + ((!n_n509) & (x20x) & (!x23x) & (n_n65) & (n_n5256)) + ((!n_n509) & (x20x) & (x23x) & (!n_n65) & (n_n5256)) + ((!n_n509) & (x20x) & (x23x) & (n_n65) & (n_n5256)) + ((n_n509) & (!x20x) & (!x23x) & (!n_n65) & (n_n5256)) + ((n_n509) & (!x20x) & (!x23x) & (n_n65) & (n_n5256)) + ((n_n509) & (!x20x) & (x23x) & (!n_n65) & (n_n5256)) + ((n_n509) & (!x20x) & (x23x) & (n_n65) & (!n_n5256)) + ((n_n509) & (!x20x) & (x23x) & (n_n65) & (n_n5256)) + ((n_n509) & (x20x) & (!x23x) & (!n_n65) & (n_n5256)) + ((n_n509) & (x20x) & (!x23x) & (n_n65) & (!n_n5256)) + ((n_n509) & (x20x) & (!x23x) & (n_n65) & (n_n5256)) + ((n_n509) & (x20x) & (x23x) & (!n_n65) & (n_n5256)) + ((n_n509) & (x20x) & (x23x) & (n_n65) & (!n_n5256)) + ((n_n509) & (x20x) & (x23x) & (n_n65) & (n_n5256)));
	assign n_n3031 = (((!x19x) & (!n_n524) & (!n_n509) & (!n_n522) & (n_n5251)) + ((!x19x) & (!n_n524) & (!n_n509) & (n_n522) & (n_n5251)) + ((!x19x) & (!n_n524) & (n_n509) & (!n_n522) & (n_n5251)) + ((!x19x) & (!n_n524) & (n_n509) & (n_n522) & (n_n5251)) + ((!x19x) & (n_n524) & (!n_n509) & (!n_n522) & (n_n5251)) + ((!x19x) & (n_n524) & (!n_n509) & (n_n522) & (n_n5251)) + ((!x19x) & (n_n524) & (n_n509) & (!n_n522) & (n_n5251)) + ((!x19x) & (n_n524) & (n_n509) & (n_n522) & (n_n5251)) + ((x19x) & (!n_n524) & (!n_n509) & (!n_n522) & (n_n5251)) + ((x19x) & (!n_n524) & (!n_n509) & (n_n522) & (n_n5251)) + ((x19x) & (!n_n524) & (n_n509) & (!n_n522) & (n_n5251)) + ((x19x) & (!n_n524) & (n_n509) & (n_n522) & (!n_n5251)) + ((x19x) & (!n_n524) & (n_n509) & (n_n522) & (n_n5251)) + ((x19x) & (n_n524) & (!n_n509) & (!n_n522) & (n_n5251)) + ((x19x) & (n_n524) & (!n_n509) & (n_n522) & (n_n5251)) + ((x19x) & (n_n524) & (n_n509) & (!n_n522) & (!n_n5251)) + ((x19x) & (n_n524) & (n_n509) & (!n_n522) & (n_n5251)) + ((x19x) & (n_n524) & (n_n509) & (n_n522) & (!n_n5251)) + ((x19x) & (n_n524) & (n_n509) & (n_n522) & (n_n5251)));
	assign x83x = (((!i_9_) & (n_n536) & (n_n473) & (n_n532) & (!n_n530)) + ((!i_9_) & (n_n536) & (n_n473) & (n_n532) & (n_n530)) + ((i_9_) & (n_n536) & (n_n473) & (!n_n532) & (n_n530)) + ((i_9_) & (n_n536) & (n_n473) & (n_n532) & (n_n530)));
	assign x427x = (((!i_9_) & (n_n536) & (n_n473) & (!n_n532) & (n_n534)) + ((!i_9_) & (n_n536) & (n_n473) & (n_n532) & (n_n534)) + ((i_9_) & (n_n536) & (n_n473) & (n_n532) & (!n_n534)) + ((i_9_) & (n_n536) & (n_n473) & (n_n532) & (n_n534)));
	assign x16666x = (((!n_n5158) & (!n_n5149) & (!n_n5148) & (!n_n5152) & (n_n5140)) + ((!n_n5158) & (!n_n5149) & (!n_n5148) & (n_n5152) & (!n_n5140)) + ((!n_n5158) & (!n_n5149) & (!n_n5148) & (n_n5152) & (n_n5140)) + ((!n_n5158) & (!n_n5149) & (n_n5148) & (!n_n5152) & (!n_n5140)) + ((!n_n5158) & (!n_n5149) & (n_n5148) & (!n_n5152) & (n_n5140)) + ((!n_n5158) & (!n_n5149) & (n_n5148) & (n_n5152) & (!n_n5140)) + ((!n_n5158) & (!n_n5149) & (n_n5148) & (n_n5152) & (n_n5140)) + ((!n_n5158) & (n_n5149) & (!n_n5148) & (!n_n5152) & (!n_n5140)) + ((!n_n5158) & (n_n5149) & (!n_n5148) & (!n_n5152) & (n_n5140)) + ((!n_n5158) & (n_n5149) & (!n_n5148) & (n_n5152) & (!n_n5140)) + ((!n_n5158) & (n_n5149) & (!n_n5148) & (n_n5152) & (n_n5140)) + ((!n_n5158) & (n_n5149) & (n_n5148) & (!n_n5152) & (!n_n5140)) + ((!n_n5158) & (n_n5149) & (n_n5148) & (!n_n5152) & (n_n5140)) + ((!n_n5158) & (n_n5149) & (n_n5148) & (n_n5152) & (!n_n5140)) + ((!n_n5158) & (n_n5149) & (n_n5148) & (n_n5152) & (n_n5140)) + ((n_n5158) & (!n_n5149) & (!n_n5148) & (!n_n5152) & (!n_n5140)) + ((n_n5158) & (!n_n5149) & (!n_n5148) & (!n_n5152) & (n_n5140)) + ((n_n5158) & (!n_n5149) & (!n_n5148) & (n_n5152) & (!n_n5140)) + ((n_n5158) & (!n_n5149) & (!n_n5148) & (n_n5152) & (n_n5140)) + ((n_n5158) & (!n_n5149) & (n_n5148) & (!n_n5152) & (!n_n5140)) + ((n_n5158) & (!n_n5149) & (n_n5148) & (!n_n5152) & (n_n5140)) + ((n_n5158) & (!n_n5149) & (n_n5148) & (n_n5152) & (!n_n5140)) + ((n_n5158) & (!n_n5149) & (n_n5148) & (n_n5152) & (n_n5140)) + ((n_n5158) & (n_n5149) & (!n_n5148) & (!n_n5152) & (!n_n5140)) + ((n_n5158) & (n_n5149) & (!n_n5148) & (!n_n5152) & (n_n5140)) + ((n_n5158) & (n_n5149) & (!n_n5148) & (n_n5152) & (!n_n5140)) + ((n_n5158) & (n_n5149) & (!n_n5148) & (n_n5152) & (n_n5140)) + ((n_n5158) & (n_n5149) & (n_n5148) & (!n_n5152) & (!n_n5140)) + ((n_n5158) & (n_n5149) & (n_n5148) & (!n_n5152) & (n_n5140)) + ((n_n5158) & (n_n5149) & (n_n5148) & (n_n5152) & (!n_n5140)) + ((n_n5158) & (n_n5149) & (n_n5148) & (n_n5152) & (n_n5140)));
	assign x22179x = (((!n_n5174) & (!n_n5179) & (!n_n5178) & (!n_n5175) & (!x332x)));
	assign n_n2205 = (((!n_n5171) & (!n_n5181) & (!n_n5177) & (!x22179x)) + ((!n_n5171) & (!n_n5181) & (n_n5177) & (!x22179x)) + ((!n_n5171) & (!n_n5181) & (n_n5177) & (x22179x)) + ((!n_n5171) & (n_n5181) & (!n_n5177) & (!x22179x)) + ((!n_n5171) & (n_n5181) & (!n_n5177) & (x22179x)) + ((!n_n5171) & (n_n5181) & (n_n5177) & (!x22179x)) + ((!n_n5171) & (n_n5181) & (n_n5177) & (x22179x)) + ((n_n5171) & (!n_n5181) & (!n_n5177) & (!x22179x)) + ((n_n5171) & (!n_n5181) & (!n_n5177) & (x22179x)) + ((n_n5171) & (!n_n5181) & (n_n5177) & (!x22179x)) + ((n_n5171) & (!n_n5181) & (n_n5177) & (x22179x)) + ((n_n5171) & (n_n5181) & (!n_n5177) & (!x22179x)) + ((n_n5171) & (n_n5181) & (!n_n5177) & (x22179x)) + ((n_n5171) & (n_n5181) & (n_n5177) & (!x22179x)) + ((n_n5171) & (n_n5181) & (n_n5177) & (x22179x)));
	assign n_n5203 = (((!i_9_) & (n_n524) & (n_n130) & (n_n464)));
	assign x22217x = (((!x223x) & (!n_n5195) & (!n_n5197) & (!n_n5208)));
	assign x16682x = (((!n_n5212) & (!n_n5203) & (!n_n2290) & (!x22217x)) + ((!n_n5212) & (!n_n5203) & (n_n2290) & (!x22217x)) + ((!n_n5212) & (!n_n5203) & (n_n2290) & (x22217x)) + ((!n_n5212) & (n_n5203) & (!n_n2290) & (!x22217x)) + ((!n_n5212) & (n_n5203) & (!n_n2290) & (x22217x)) + ((!n_n5212) & (n_n5203) & (n_n2290) & (!x22217x)) + ((!n_n5212) & (n_n5203) & (n_n2290) & (x22217x)) + ((n_n5212) & (!n_n5203) & (!n_n2290) & (!x22217x)) + ((n_n5212) & (!n_n5203) & (!n_n2290) & (x22217x)) + ((n_n5212) & (!n_n5203) & (n_n2290) & (!x22217x)) + ((n_n5212) & (!n_n5203) & (n_n2290) & (x22217x)) + ((n_n5212) & (n_n5203) & (!n_n2290) & (!x22217x)) + ((n_n5212) & (n_n5203) & (!n_n2290) & (x22217x)) + ((n_n5212) & (n_n5203) & (n_n2290) & (!x22217x)) + ((n_n5212) & (n_n5203) & (n_n2290) & (x22217x)));
	assign n_n2204 = (((!n_n5186) & (!n_n5187) & (!n_n5188) & (!x113x) & (!x22199x)) + ((!n_n5186) & (!n_n5187) & (!n_n5188) & (x113x) & (!x22199x)) + ((!n_n5186) & (!n_n5187) & (!n_n5188) & (x113x) & (x22199x)) + ((!n_n5186) & (!n_n5187) & (n_n5188) & (!x113x) & (!x22199x)) + ((!n_n5186) & (!n_n5187) & (n_n5188) & (!x113x) & (x22199x)) + ((!n_n5186) & (!n_n5187) & (n_n5188) & (x113x) & (!x22199x)) + ((!n_n5186) & (!n_n5187) & (n_n5188) & (x113x) & (x22199x)) + ((!n_n5186) & (n_n5187) & (!n_n5188) & (!x113x) & (!x22199x)) + ((!n_n5186) & (n_n5187) & (!n_n5188) & (!x113x) & (x22199x)) + ((!n_n5186) & (n_n5187) & (!n_n5188) & (x113x) & (!x22199x)) + ((!n_n5186) & (n_n5187) & (!n_n5188) & (x113x) & (x22199x)) + ((!n_n5186) & (n_n5187) & (n_n5188) & (!x113x) & (!x22199x)) + ((!n_n5186) & (n_n5187) & (n_n5188) & (!x113x) & (x22199x)) + ((!n_n5186) & (n_n5187) & (n_n5188) & (x113x) & (!x22199x)) + ((!n_n5186) & (n_n5187) & (n_n5188) & (x113x) & (x22199x)) + ((n_n5186) & (!n_n5187) & (!n_n5188) & (!x113x) & (!x22199x)) + ((n_n5186) & (!n_n5187) & (!n_n5188) & (!x113x) & (x22199x)) + ((n_n5186) & (!n_n5187) & (!n_n5188) & (x113x) & (!x22199x)) + ((n_n5186) & (!n_n5187) & (!n_n5188) & (x113x) & (x22199x)) + ((n_n5186) & (!n_n5187) & (n_n5188) & (!x113x) & (!x22199x)) + ((n_n5186) & (!n_n5187) & (n_n5188) & (!x113x) & (x22199x)) + ((n_n5186) & (!n_n5187) & (n_n5188) & (x113x) & (!x22199x)) + ((n_n5186) & (!n_n5187) & (n_n5188) & (x113x) & (x22199x)) + ((n_n5186) & (n_n5187) & (!n_n5188) & (!x113x) & (!x22199x)) + ((n_n5186) & (n_n5187) & (!n_n5188) & (!x113x) & (x22199x)) + ((n_n5186) & (n_n5187) & (!n_n5188) & (x113x) & (!x22199x)) + ((n_n5186) & (n_n5187) & (!n_n5188) & (x113x) & (x22199x)) + ((n_n5186) & (n_n5187) & (n_n5188) & (!x113x) & (!x22199x)) + ((n_n5186) & (n_n5187) & (n_n5188) & (!x113x) & (x22199x)) + ((n_n5186) & (n_n5187) & (n_n5188) & (x113x) & (!x22199x)) + ((n_n5186) & (n_n5187) & (n_n5188) & (x113x) & (x22199x)));
	assign x16681x = (((!n_n5204) & (!n_n5205) & (!x454x) & (!x36x) & (x451x)) + ((!n_n5204) & (!n_n5205) & (!x454x) & (x36x) & (!x451x)) + ((!n_n5204) & (!n_n5205) & (!x454x) & (x36x) & (x451x)) + ((!n_n5204) & (!n_n5205) & (x454x) & (!x36x) & (!x451x)) + ((!n_n5204) & (!n_n5205) & (x454x) & (!x36x) & (x451x)) + ((!n_n5204) & (!n_n5205) & (x454x) & (x36x) & (!x451x)) + ((!n_n5204) & (!n_n5205) & (x454x) & (x36x) & (x451x)) + ((!n_n5204) & (n_n5205) & (!x454x) & (!x36x) & (!x451x)) + ((!n_n5204) & (n_n5205) & (!x454x) & (!x36x) & (x451x)) + ((!n_n5204) & (n_n5205) & (!x454x) & (x36x) & (!x451x)) + ((!n_n5204) & (n_n5205) & (!x454x) & (x36x) & (x451x)) + ((!n_n5204) & (n_n5205) & (x454x) & (!x36x) & (!x451x)) + ((!n_n5204) & (n_n5205) & (x454x) & (!x36x) & (x451x)) + ((!n_n5204) & (n_n5205) & (x454x) & (x36x) & (!x451x)) + ((!n_n5204) & (n_n5205) & (x454x) & (x36x) & (x451x)) + ((n_n5204) & (!n_n5205) & (!x454x) & (!x36x) & (!x451x)) + ((n_n5204) & (!n_n5205) & (!x454x) & (!x36x) & (x451x)) + ((n_n5204) & (!n_n5205) & (!x454x) & (x36x) & (!x451x)) + ((n_n5204) & (!n_n5205) & (!x454x) & (x36x) & (x451x)) + ((n_n5204) & (!n_n5205) & (x454x) & (!x36x) & (!x451x)) + ((n_n5204) & (!n_n5205) & (x454x) & (!x36x) & (x451x)) + ((n_n5204) & (!n_n5205) & (x454x) & (x36x) & (!x451x)) + ((n_n5204) & (!n_n5205) & (x454x) & (x36x) & (x451x)) + ((n_n5204) & (n_n5205) & (!x454x) & (!x36x) & (!x451x)) + ((n_n5204) & (n_n5205) & (!x454x) & (!x36x) & (x451x)) + ((n_n5204) & (n_n5205) & (!x454x) & (x36x) & (!x451x)) + ((n_n5204) & (n_n5205) & (!x454x) & (x36x) & (x451x)) + ((n_n5204) & (n_n5205) & (x454x) & (!x36x) & (!x451x)) + ((n_n5204) & (n_n5205) & (x454x) & (!x36x) & (x451x)) + ((n_n5204) & (n_n5205) & (x454x) & (x36x) & (!x451x)) + ((n_n5204) & (n_n5205) & (x454x) & (x36x) & (x451x)));
	assign x16695x = (((!n_n5232) & (!n_n5237) & (!x62x) & (!x181x) & (x183x)) + ((!n_n5232) & (!n_n5237) & (!x62x) & (x181x) & (!x183x)) + ((!n_n5232) & (!n_n5237) & (!x62x) & (x181x) & (x183x)) + ((!n_n5232) & (!n_n5237) & (x62x) & (!x181x) & (!x183x)) + ((!n_n5232) & (!n_n5237) & (x62x) & (!x181x) & (x183x)) + ((!n_n5232) & (!n_n5237) & (x62x) & (x181x) & (!x183x)) + ((!n_n5232) & (!n_n5237) & (x62x) & (x181x) & (x183x)) + ((!n_n5232) & (n_n5237) & (!x62x) & (!x181x) & (!x183x)) + ((!n_n5232) & (n_n5237) & (!x62x) & (!x181x) & (x183x)) + ((!n_n5232) & (n_n5237) & (!x62x) & (x181x) & (!x183x)) + ((!n_n5232) & (n_n5237) & (!x62x) & (x181x) & (x183x)) + ((!n_n5232) & (n_n5237) & (x62x) & (!x181x) & (!x183x)) + ((!n_n5232) & (n_n5237) & (x62x) & (!x181x) & (x183x)) + ((!n_n5232) & (n_n5237) & (x62x) & (x181x) & (!x183x)) + ((!n_n5232) & (n_n5237) & (x62x) & (x181x) & (x183x)) + ((n_n5232) & (!n_n5237) & (!x62x) & (!x181x) & (!x183x)) + ((n_n5232) & (!n_n5237) & (!x62x) & (!x181x) & (x183x)) + ((n_n5232) & (!n_n5237) & (!x62x) & (x181x) & (!x183x)) + ((n_n5232) & (!n_n5237) & (!x62x) & (x181x) & (x183x)) + ((n_n5232) & (!n_n5237) & (x62x) & (!x181x) & (!x183x)) + ((n_n5232) & (!n_n5237) & (x62x) & (!x181x) & (x183x)) + ((n_n5232) & (!n_n5237) & (x62x) & (x181x) & (!x183x)) + ((n_n5232) & (!n_n5237) & (x62x) & (x181x) & (x183x)) + ((n_n5232) & (n_n5237) & (!x62x) & (!x181x) & (!x183x)) + ((n_n5232) & (n_n5237) & (!x62x) & (!x181x) & (x183x)) + ((n_n5232) & (n_n5237) & (!x62x) & (x181x) & (!x183x)) + ((n_n5232) & (n_n5237) & (!x62x) & (x181x) & (x183x)) + ((n_n5232) & (n_n5237) & (x62x) & (!x181x) & (!x183x)) + ((n_n5232) & (n_n5237) & (x62x) & (!x181x) & (x183x)) + ((n_n5232) & (n_n5237) & (x62x) & (x181x) & (!x183x)) + ((n_n5232) & (n_n5237) & (x62x) & (x181x) & (x183x)));
	assign x16697x = (((!n_n5247) & (!n_n5246) & (!x319x) & (!x16687x) & (x16695x)) + ((!n_n5247) & (!n_n5246) & (!x319x) & (x16687x) & (!x16695x)) + ((!n_n5247) & (!n_n5246) & (!x319x) & (x16687x) & (x16695x)) + ((!n_n5247) & (!n_n5246) & (x319x) & (!x16687x) & (!x16695x)) + ((!n_n5247) & (!n_n5246) & (x319x) & (!x16687x) & (x16695x)) + ((!n_n5247) & (!n_n5246) & (x319x) & (x16687x) & (!x16695x)) + ((!n_n5247) & (!n_n5246) & (x319x) & (x16687x) & (x16695x)) + ((!n_n5247) & (n_n5246) & (!x319x) & (!x16687x) & (!x16695x)) + ((!n_n5247) & (n_n5246) & (!x319x) & (!x16687x) & (x16695x)) + ((!n_n5247) & (n_n5246) & (!x319x) & (x16687x) & (!x16695x)) + ((!n_n5247) & (n_n5246) & (!x319x) & (x16687x) & (x16695x)) + ((!n_n5247) & (n_n5246) & (x319x) & (!x16687x) & (!x16695x)) + ((!n_n5247) & (n_n5246) & (x319x) & (!x16687x) & (x16695x)) + ((!n_n5247) & (n_n5246) & (x319x) & (x16687x) & (!x16695x)) + ((!n_n5247) & (n_n5246) & (x319x) & (x16687x) & (x16695x)) + ((n_n5247) & (!n_n5246) & (!x319x) & (!x16687x) & (!x16695x)) + ((n_n5247) & (!n_n5246) & (!x319x) & (!x16687x) & (x16695x)) + ((n_n5247) & (!n_n5246) & (!x319x) & (x16687x) & (!x16695x)) + ((n_n5247) & (!n_n5246) & (!x319x) & (x16687x) & (x16695x)) + ((n_n5247) & (!n_n5246) & (x319x) & (!x16687x) & (!x16695x)) + ((n_n5247) & (!n_n5246) & (x319x) & (!x16687x) & (x16695x)) + ((n_n5247) & (!n_n5246) & (x319x) & (x16687x) & (!x16695x)) + ((n_n5247) & (!n_n5246) & (x319x) & (x16687x) & (x16695x)) + ((n_n5247) & (n_n5246) & (!x319x) & (!x16687x) & (!x16695x)) + ((n_n5247) & (n_n5246) & (!x319x) & (!x16687x) & (x16695x)) + ((n_n5247) & (n_n5246) & (!x319x) & (x16687x) & (!x16695x)) + ((n_n5247) & (n_n5246) & (!x319x) & (x16687x) & (x16695x)) + ((n_n5247) & (n_n5246) & (x319x) & (!x16687x) & (!x16695x)) + ((n_n5247) & (n_n5246) & (x319x) & (!x16687x) & (x16695x)) + ((n_n5247) & (n_n5246) & (x319x) & (x16687x) & (!x16695x)) + ((n_n5247) & (n_n5246) & (x319x) & (x16687x) & (x16695x)));
	assign x16693x = (((!n_n5260) & (!n_n5226) & (!n_n5235) & (n_n5234)) + ((!n_n5260) & (!n_n5226) & (n_n5235) & (!n_n5234)) + ((!n_n5260) & (!n_n5226) & (n_n5235) & (n_n5234)) + ((!n_n5260) & (n_n5226) & (!n_n5235) & (!n_n5234)) + ((!n_n5260) & (n_n5226) & (!n_n5235) & (n_n5234)) + ((!n_n5260) & (n_n5226) & (n_n5235) & (!n_n5234)) + ((!n_n5260) & (n_n5226) & (n_n5235) & (n_n5234)) + ((n_n5260) & (!n_n5226) & (!n_n5235) & (!n_n5234)) + ((n_n5260) & (!n_n5226) & (!n_n5235) & (n_n5234)) + ((n_n5260) & (!n_n5226) & (n_n5235) & (!n_n5234)) + ((n_n5260) & (!n_n5226) & (n_n5235) & (n_n5234)) + ((n_n5260) & (n_n5226) & (!n_n5235) & (!n_n5234)) + ((n_n5260) & (n_n5226) & (!n_n5235) & (n_n5234)) + ((n_n5260) & (n_n5226) & (n_n5235) & (!n_n5234)) + ((n_n5260) & (n_n5226) & (n_n5235) & (n_n5234)));
	assign x16703x = (((!n_n5161) & (!n_n5160) & (!x33x) & (!n_n5170) & (!x22059x)) + ((!n_n5161) & (!n_n5160) & (!x33x) & (n_n5170) & (!x22059x)) + ((!n_n5161) & (!n_n5160) & (!x33x) & (n_n5170) & (x22059x)) + ((!n_n5161) & (!n_n5160) & (x33x) & (!n_n5170) & (!x22059x)) + ((!n_n5161) & (!n_n5160) & (x33x) & (!n_n5170) & (x22059x)) + ((!n_n5161) & (!n_n5160) & (x33x) & (n_n5170) & (!x22059x)) + ((!n_n5161) & (!n_n5160) & (x33x) & (n_n5170) & (x22059x)) + ((!n_n5161) & (n_n5160) & (!x33x) & (!n_n5170) & (!x22059x)) + ((!n_n5161) & (n_n5160) & (!x33x) & (!n_n5170) & (x22059x)) + ((!n_n5161) & (n_n5160) & (!x33x) & (n_n5170) & (!x22059x)) + ((!n_n5161) & (n_n5160) & (!x33x) & (n_n5170) & (x22059x)) + ((!n_n5161) & (n_n5160) & (x33x) & (!n_n5170) & (!x22059x)) + ((!n_n5161) & (n_n5160) & (x33x) & (!n_n5170) & (x22059x)) + ((!n_n5161) & (n_n5160) & (x33x) & (n_n5170) & (!x22059x)) + ((!n_n5161) & (n_n5160) & (x33x) & (n_n5170) & (x22059x)) + ((n_n5161) & (!n_n5160) & (!x33x) & (!n_n5170) & (!x22059x)) + ((n_n5161) & (!n_n5160) & (!x33x) & (!n_n5170) & (x22059x)) + ((n_n5161) & (!n_n5160) & (!x33x) & (n_n5170) & (!x22059x)) + ((n_n5161) & (!n_n5160) & (!x33x) & (n_n5170) & (x22059x)) + ((n_n5161) & (!n_n5160) & (x33x) & (!n_n5170) & (!x22059x)) + ((n_n5161) & (!n_n5160) & (x33x) & (!n_n5170) & (x22059x)) + ((n_n5161) & (!n_n5160) & (x33x) & (n_n5170) & (!x22059x)) + ((n_n5161) & (!n_n5160) & (x33x) & (n_n5170) & (x22059x)) + ((n_n5161) & (n_n5160) & (!x33x) & (!n_n5170) & (!x22059x)) + ((n_n5161) & (n_n5160) & (!x33x) & (!n_n5170) & (x22059x)) + ((n_n5161) & (n_n5160) & (!x33x) & (n_n5170) & (!x22059x)) + ((n_n5161) & (n_n5160) & (!x33x) & (n_n5170) & (x22059x)) + ((n_n5161) & (n_n5160) & (x33x) & (!n_n5170) & (!x22059x)) + ((n_n5161) & (n_n5160) & (x33x) & (!n_n5170) & (x22059x)) + ((n_n5161) & (n_n5160) & (x33x) & (n_n5170) & (!x22059x)) + ((n_n5161) & (n_n5160) & (x33x) & (n_n5170) & (x22059x)));
	assign x16715x = (((!n_n4152) & (!n_n5079) & (!n_n5083) & (x144x)) + ((!n_n4152) & (!n_n5079) & (n_n5083) & (!x144x)) + ((!n_n4152) & (!n_n5079) & (n_n5083) & (x144x)) + ((!n_n4152) & (n_n5079) & (!n_n5083) & (!x144x)) + ((!n_n4152) & (n_n5079) & (!n_n5083) & (x144x)) + ((!n_n4152) & (n_n5079) & (n_n5083) & (!x144x)) + ((!n_n4152) & (n_n5079) & (n_n5083) & (x144x)) + ((n_n4152) & (!n_n5079) & (!n_n5083) & (!x144x)) + ((n_n4152) & (!n_n5079) & (!n_n5083) & (x144x)) + ((n_n4152) & (!n_n5079) & (n_n5083) & (!x144x)) + ((n_n4152) & (!n_n5079) & (n_n5083) & (x144x)) + ((n_n4152) & (n_n5079) & (!n_n5083) & (!x144x)) + ((n_n4152) & (n_n5079) & (!n_n5083) & (x144x)) + ((n_n4152) & (n_n5079) & (n_n5083) & (!x144x)) + ((n_n4152) & (n_n5079) & (n_n5083) & (x144x)));
	assign x16711x = (((!n_n5064) & (!n_n5081) & (!n_n5087) & (n_n5082)) + ((!n_n5064) & (!n_n5081) & (n_n5087) & (!n_n5082)) + ((!n_n5064) & (!n_n5081) & (n_n5087) & (n_n5082)) + ((!n_n5064) & (n_n5081) & (!n_n5087) & (!n_n5082)) + ((!n_n5064) & (n_n5081) & (!n_n5087) & (n_n5082)) + ((!n_n5064) & (n_n5081) & (n_n5087) & (!n_n5082)) + ((!n_n5064) & (n_n5081) & (n_n5087) & (n_n5082)) + ((n_n5064) & (!n_n5081) & (!n_n5087) & (!n_n5082)) + ((n_n5064) & (!n_n5081) & (!n_n5087) & (n_n5082)) + ((n_n5064) & (!n_n5081) & (n_n5087) & (!n_n5082)) + ((n_n5064) & (!n_n5081) & (n_n5087) & (n_n5082)) + ((n_n5064) & (n_n5081) & (!n_n5087) & (!n_n5082)) + ((n_n5064) & (n_n5081) & (!n_n5087) & (n_n5082)) + ((n_n5064) & (n_n5081) & (n_n5087) & (!n_n5082)) + ((n_n5064) & (n_n5081) & (n_n5087) & (n_n5082)));
	assign x16713x = (((!n_n5085) & (!x344x) & (!n_n5084) & (!n_n5068) & (x159x)) + ((!n_n5085) & (!x344x) & (!n_n5084) & (n_n5068) & (!x159x)) + ((!n_n5085) & (!x344x) & (!n_n5084) & (n_n5068) & (x159x)) + ((!n_n5085) & (!x344x) & (n_n5084) & (!n_n5068) & (!x159x)) + ((!n_n5085) & (!x344x) & (n_n5084) & (!n_n5068) & (x159x)) + ((!n_n5085) & (!x344x) & (n_n5084) & (n_n5068) & (!x159x)) + ((!n_n5085) & (!x344x) & (n_n5084) & (n_n5068) & (x159x)) + ((!n_n5085) & (x344x) & (!n_n5084) & (!n_n5068) & (!x159x)) + ((!n_n5085) & (x344x) & (!n_n5084) & (!n_n5068) & (x159x)) + ((!n_n5085) & (x344x) & (!n_n5084) & (n_n5068) & (!x159x)) + ((!n_n5085) & (x344x) & (!n_n5084) & (n_n5068) & (x159x)) + ((!n_n5085) & (x344x) & (n_n5084) & (!n_n5068) & (!x159x)) + ((!n_n5085) & (x344x) & (n_n5084) & (!n_n5068) & (x159x)) + ((!n_n5085) & (x344x) & (n_n5084) & (n_n5068) & (!x159x)) + ((!n_n5085) & (x344x) & (n_n5084) & (n_n5068) & (x159x)) + ((n_n5085) & (!x344x) & (!n_n5084) & (!n_n5068) & (!x159x)) + ((n_n5085) & (!x344x) & (!n_n5084) & (!n_n5068) & (x159x)) + ((n_n5085) & (!x344x) & (!n_n5084) & (n_n5068) & (!x159x)) + ((n_n5085) & (!x344x) & (!n_n5084) & (n_n5068) & (x159x)) + ((n_n5085) & (!x344x) & (n_n5084) & (!n_n5068) & (!x159x)) + ((n_n5085) & (!x344x) & (n_n5084) & (!n_n5068) & (x159x)) + ((n_n5085) & (!x344x) & (n_n5084) & (n_n5068) & (!x159x)) + ((n_n5085) & (!x344x) & (n_n5084) & (n_n5068) & (x159x)) + ((n_n5085) & (x344x) & (!n_n5084) & (!n_n5068) & (!x159x)) + ((n_n5085) & (x344x) & (!n_n5084) & (!n_n5068) & (x159x)) + ((n_n5085) & (x344x) & (!n_n5084) & (n_n5068) & (!x159x)) + ((n_n5085) & (x344x) & (!n_n5084) & (n_n5068) & (x159x)) + ((n_n5085) & (x344x) & (n_n5084) & (!n_n5068) & (!x159x)) + ((n_n5085) & (x344x) & (n_n5084) & (!n_n5068) & (x159x)) + ((n_n5085) & (x344x) & (n_n5084) & (n_n5068) & (!x159x)) + ((n_n5085) & (x344x) & (n_n5084) & (n_n5068) & (x159x)));
	assign x16728x = (((!n_n5136) & (!n_n5127) & (!n_n5128) & (n_n5135)) + ((!n_n5136) & (!n_n5127) & (n_n5128) & (!n_n5135)) + ((!n_n5136) & (!n_n5127) & (n_n5128) & (n_n5135)) + ((!n_n5136) & (n_n5127) & (!n_n5128) & (!n_n5135)) + ((!n_n5136) & (n_n5127) & (!n_n5128) & (n_n5135)) + ((!n_n5136) & (n_n5127) & (n_n5128) & (!n_n5135)) + ((!n_n5136) & (n_n5127) & (n_n5128) & (n_n5135)) + ((n_n5136) & (!n_n5127) & (!n_n5128) & (!n_n5135)) + ((n_n5136) & (!n_n5127) & (!n_n5128) & (n_n5135)) + ((n_n5136) & (!n_n5127) & (n_n5128) & (!n_n5135)) + ((n_n5136) & (!n_n5127) & (n_n5128) & (n_n5135)) + ((n_n5136) & (n_n5127) & (!n_n5128) & (!n_n5135)) + ((n_n5136) & (n_n5127) & (!n_n5128) & (n_n5135)) + ((n_n5136) & (n_n5127) & (n_n5128) & (!n_n5135)) + ((n_n5136) & (n_n5127) & (n_n5128) & (n_n5135)));
	assign x16729x = (((!x21x) & (!n_n130) & (!n_n500) & (!n_n5125) & (n_n2304)) + ((!x21x) & (!n_n130) & (!n_n500) & (n_n5125) & (!n_n2304)) + ((!x21x) & (!n_n130) & (!n_n500) & (n_n5125) & (n_n2304)) + ((!x21x) & (!n_n130) & (n_n500) & (!n_n5125) & (n_n2304)) + ((!x21x) & (!n_n130) & (n_n500) & (n_n5125) & (!n_n2304)) + ((!x21x) & (!n_n130) & (n_n500) & (n_n5125) & (n_n2304)) + ((!x21x) & (n_n130) & (!n_n500) & (!n_n5125) & (n_n2304)) + ((!x21x) & (n_n130) & (!n_n500) & (n_n5125) & (!n_n2304)) + ((!x21x) & (n_n130) & (!n_n500) & (n_n5125) & (n_n2304)) + ((!x21x) & (n_n130) & (n_n500) & (!n_n5125) & (n_n2304)) + ((!x21x) & (n_n130) & (n_n500) & (n_n5125) & (!n_n2304)) + ((!x21x) & (n_n130) & (n_n500) & (n_n5125) & (n_n2304)) + ((x21x) & (!n_n130) & (!n_n500) & (!n_n5125) & (n_n2304)) + ((x21x) & (!n_n130) & (!n_n500) & (n_n5125) & (!n_n2304)) + ((x21x) & (!n_n130) & (!n_n500) & (n_n5125) & (n_n2304)) + ((x21x) & (!n_n130) & (n_n500) & (!n_n5125) & (n_n2304)) + ((x21x) & (!n_n130) & (n_n500) & (n_n5125) & (!n_n2304)) + ((x21x) & (!n_n130) & (n_n500) & (n_n5125) & (n_n2304)) + ((x21x) & (n_n130) & (!n_n500) & (!n_n5125) & (n_n2304)) + ((x21x) & (n_n130) & (!n_n500) & (n_n5125) & (!n_n2304)) + ((x21x) & (n_n130) & (!n_n500) & (n_n5125) & (n_n2304)) + ((x21x) & (n_n130) & (n_n500) & (!n_n5125) & (!n_n2304)) + ((x21x) & (n_n130) & (n_n500) & (!n_n5125) & (n_n2304)) + ((x21x) & (n_n130) & (n_n500) & (n_n5125) & (!n_n2304)) + ((x21x) & (n_n130) & (n_n500) & (n_n5125) & (n_n2304)));
	assign x22221x = (((!n_n5060) & (!n_n5055) & (!n_n5057) & (!n_n5058)));
	assign x22225x = (((!n_n5274) & (!n_n5266) & (!n_n5285) & (!x14542x)));
	assign x16758x = (((!n_n5275) & (!n_n5281) & (!n_n5261) & (!x217x) & (!x22225x)) + ((!n_n5275) & (!n_n5281) & (!n_n5261) & (x217x) & (!x22225x)) + ((!n_n5275) & (!n_n5281) & (!n_n5261) & (x217x) & (x22225x)) + ((!n_n5275) & (!n_n5281) & (n_n5261) & (!x217x) & (!x22225x)) + ((!n_n5275) & (!n_n5281) & (n_n5261) & (!x217x) & (x22225x)) + ((!n_n5275) & (!n_n5281) & (n_n5261) & (x217x) & (!x22225x)) + ((!n_n5275) & (!n_n5281) & (n_n5261) & (x217x) & (x22225x)) + ((!n_n5275) & (n_n5281) & (!n_n5261) & (!x217x) & (!x22225x)) + ((!n_n5275) & (n_n5281) & (!n_n5261) & (!x217x) & (x22225x)) + ((!n_n5275) & (n_n5281) & (!n_n5261) & (x217x) & (!x22225x)) + ((!n_n5275) & (n_n5281) & (!n_n5261) & (x217x) & (x22225x)) + ((!n_n5275) & (n_n5281) & (n_n5261) & (!x217x) & (!x22225x)) + ((!n_n5275) & (n_n5281) & (n_n5261) & (!x217x) & (x22225x)) + ((!n_n5275) & (n_n5281) & (n_n5261) & (x217x) & (!x22225x)) + ((!n_n5275) & (n_n5281) & (n_n5261) & (x217x) & (x22225x)) + ((n_n5275) & (!n_n5281) & (!n_n5261) & (!x217x) & (!x22225x)) + ((n_n5275) & (!n_n5281) & (!n_n5261) & (!x217x) & (x22225x)) + ((n_n5275) & (!n_n5281) & (!n_n5261) & (x217x) & (!x22225x)) + ((n_n5275) & (!n_n5281) & (!n_n5261) & (x217x) & (x22225x)) + ((n_n5275) & (!n_n5281) & (n_n5261) & (!x217x) & (!x22225x)) + ((n_n5275) & (!n_n5281) & (n_n5261) & (!x217x) & (x22225x)) + ((n_n5275) & (!n_n5281) & (n_n5261) & (x217x) & (!x22225x)) + ((n_n5275) & (!n_n5281) & (n_n5261) & (x217x) & (x22225x)) + ((n_n5275) & (n_n5281) & (!n_n5261) & (!x217x) & (!x22225x)) + ((n_n5275) & (n_n5281) & (!n_n5261) & (!x217x) & (x22225x)) + ((n_n5275) & (n_n5281) & (!n_n5261) & (x217x) & (!x22225x)) + ((n_n5275) & (n_n5281) & (!n_n5261) & (x217x) & (x22225x)) + ((n_n5275) & (n_n5281) & (n_n5261) & (!x217x) & (!x22225x)) + ((n_n5275) & (n_n5281) & (n_n5261) & (!x217x) & (x22225x)) + ((n_n5275) & (n_n5281) & (n_n5261) & (x217x) & (!x22225x)) + ((n_n5275) & (n_n5281) & (n_n5261) & (x217x) & (x22225x)));
	assign n_n2196 = (((!n_n5293) & (!n_n5296) & (!n_n5297) & (!n_n5298) & (x16750x)) + ((!n_n5293) & (!n_n5296) & (!n_n5297) & (n_n5298) & (!x16750x)) + ((!n_n5293) & (!n_n5296) & (!n_n5297) & (n_n5298) & (x16750x)) + ((!n_n5293) & (!n_n5296) & (n_n5297) & (!n_n5298) & (!x16750x)) + ((!n_n5293) & (!n_n5296) & (n_n5297) & (!n_n5298) & (x16750x)) + ((!n_n5293) & (!n_n5296) & (n_n5297) & (n_n5298) & (!x16750x)) + ((!n_n5293) & (!n_n5296) & (n_n5297) & (n_n5298) & (x16750x)) + ((!n_n5293) & (n_n5296) & (!n_n5297) & (!n_n5298) & (!x16750x)) + ((!n_n5293) & (n_n5296) & (!n_n5297) & (!n_n5298) & (x16750x)) + ((!n_n5293) & (n_n5296) & (!n_n5297) & (n_n5298) & (!x16750x)) + ((!n_n5293) & (n_n5296) & (!n_n5297) & (n_n5298) & (x16750x)) + ((!n_n5293) & (n_n5296) & (n_n5297) & (!n_n5298) & (!x16750x)) + ((!n_n5293) & (n_n5296) & (n_n5297) & (!n_n5298) & (x16750x)) + ((!n_n5293) & (n_n5296) & (n_n5297) & (n_n5298) & (!x16750x)) + ((!n_n5293) & (n_n5296) & (n_n5297) & (n_n5298) & (x16750x)) + ((n_n5293) & (!n_n5296) & (!n_n5297) & (!n_n5298) & (!x16750x)) + ((n_n5293) & (!n_n5296) & (!n_n5297) & (!n_n5298) & (x16750x)) + ((n_n5293) & (!n_n5296) & (!n_n5297) & (n_n5298) & (!x16750x)) + ((n_n5293) & (!n_n5296) & (!n_n5297) & (n_n5298) & (x16750x)) + ((n_n5293) & (!n_n5296) & (n_n5297) & (!n_n5298) & (!x16750x)) + ((n_n5293) & (!n_n5296) & (n_n5297) & (!n_n5298) & (x16750x)) + ((n_n5293) & (!n_n5296) & (n_n5297) & (n_n5298) & (!x16750x)) + ((n_n5293) & (!n_n5296) & (n_n5297) & (n_n5298) & (x16750x)) + ((n_n5293) & (n_n5296) & (!n_n5297) & (!n_n5298) & (!x16750x)) + ((n_n5293) & (n_n5296) & (!n_n5297) & (!n_n5298) & (x16750x)) + ((n_n5293) & (n_n5296) & (!n_n5297) & (n_n5298) & (!x16750x)) + ((n_n5293) & (n_n5296) & (!n_n5297) & (n_n5298) & (x16750x)) + ((n_n5293) & (n_n5296) & (n_n5297) & (!n_n5298) & (!x16750x)) + ((n_n5293) & (n_n5296) & (n_n5297) & (!n_n5298) & (x16750x)) + ((n_n5293) & (n_n5296) & (n_n5297) & (n_n5298) & (!x16750x)) + ((n_n5293) & (n_n5296) & (n_n5297) & (n_n5298) & (x16750x)));
	assign x16757x = (((!n_n5273) & (!n_n5272) & (!x205x) & (!x419x) & (x438x)) + ((!n_n5273) & (!n_n5272) & (!x205x) & (x419x) & (!x438x)) + ((!n_n5273) & (!n_n5272) & (!x205x) & (x419x) & (x438x)) + ((!n_n5273) & (!n_n5272) & (x205x) & (!x419x) & (!x438x)) + ((!n_n5273) & (!n_n5272) & (x205x) & (!x419x) & (x438x)) + ((!n_n5273) & (!n_n5272) & (x205x) & (x419x) & (!x438x)) + ((!n_n5273) & (!n_n5272) & (x205x) & (x419x) & (x438x)) + ((!n_n5273) & (n_n5272) & (!x205x) & (!x419x) & (!x438x)) + ((!n_n5273) & (n_n5272) & (!x205x) & (!x419x) & (x438x)) + ((!n_n5273) & (n_n5272) & (!x205x) & (x419x) & (!x438x)) + ((!n_n5273) & (n_n5272) & (!x205x) & (x419x) & (x438x)) + ((!n_n5273) & (n_n5272) & (x205x) & (!x419x) & (!x438x)) + ((!n_n5273) & (n_n5272) & (x205x) & (!x419x) & (x438x)) + ((!n_n5273) & (n_n5272) & (x205x) & (x419x) & (!x438x)) + ((!n_n5273) & (n_n5272) & (x205x) & (x419x) & (x438x)) + ((n_n5273) & (!n_n5272) & (!x205x) & (!x419x) & (!x438x)) + ((n_n5273) & (!n_n5272) & (!x205x) & (!x419x) & (x438x)) + ((n_n5273) & (!n_n5272) & (!x205x) & (x419x) & (!x438x)) + ((n_n5273) & (!n_n5272) & (!x205x) & (x419x) & (x438x)) + ((n_n5273) & (!n_n5272) & (x205x) & (!x419x) & (!x438x)) + ((n_n5273) & (!n_n5272) & (x205x) & (!x419x) & (x438x)) + ((n_n5273) & (!n_n5272) & (x205x) & (x419x) & (!x438x)) + ((n_n5273) & (!n_n5272) & (x205x) & (x419x) & (x438x)) + ((n_n5273) & (n_n5272) & (!x205x) & (!x419x) & (!x438x)) + ((n_n5273) & (n_n5272) & (!x205x) & (!x419x) & (x438x)) + ((n_n5273) & (n_n5272) & (!x205x) & (x419x) & (!x438x)) + ((n_n5273) & (n_n5272) & (!x205x) & (x419x) & (x438x)) + ((n_n5273) & (n_n5272) & (x205x) & (!x419x) & (!x438x)) + ((n_n5273) & (n_n5272) & (x205x) & (!x419x) & (x438x)) + ((n_n5273) & (n_n5272) & (x205x) & (x419x) & (!x438x)) + ((n_n5273) & (n_n5272) & (x205x) & (x419x) & (x438x)));
	assign n_n5334 = (((!i_7_) & (!i_8_) & (!i_6_) & (x19x) & (n_n464)));
	assign n_n5333 = (((!i_5_) & (!i_3_) & (!i_4_) & (x20x) & (n_n65)));
	assign n_n4813 = (((!i_9_) & (n_n325) & (n_n530) & (n_n464)));
	assign n_n4815 = (((!i_9_) & (n_n528) & (n_n325) & (n_n464)));
	assign x16812x = (((!n_n4827) & (!n_n4816) & (!n_n4833) & (n_n4813)) + ((!n_n4827) & (!n_n4816) & (n_n4833) & (!n_n4813)) + ((!n_n4827) & (!n_n4816) & (n_n4833) & (n_n4813)) + ((!n_n4827) & (n_n4816) & (!n_n4833) & (!n_n4813)) + ((!n_n4827) & (n_n4816) & (!n_n4833) & (n_n4813)) + ((!n_n4827) & (n_n4816) & (n_n4833) & (!n_n4813)) + ((!n_n4827) & (n_n4816) & (n_n4833) & (n_n4813)) + ((n_n4827) & (!n_n4816) & (!n_n4833) & (!n_n4813)) + ((n_n4827) & (!n_n4816) & (!n_n4833) & (n_n4813)) + ((n_n4827) & (!n_n4816) & (n_n4833) & (!n_n4813)) + ((n_n4827) & (!n_n4816) & (n_n4833) & (n_n4813)) + ((n_n4827) & (n_n4816) & (!n_n4833) & (!n_n4813)) + ((n_n4827) & (n_n4816) & (!n_n4833) & (n_n4813)) + ((n_n4827) & (n_n4816) & (n_n4833) & (!n_n4813)) + ((n_n4827) & (n_n4816) & (n_n4833) & (n_n4813)));
	assign x16813x = (((!n_n4847) & (!n_n4817) & (!n_n4838) & (!n_n4815) & (x85x)) + ((!n_n4847) & (!n_n4817) & (!n_n4838) & (n_n4815) & (!x85x)) + ((!n_n4847) & (!n_n4817) & (!n_n4838) & (n_n4815) & (x85x)) + ((!n_n4847) & (!n_n4817) & (n_n4838) & (!n_n4815) & (!x85x)) + ((!n_n4847) & (!n_n4817) & (n_n4838) & (!n_n4815) & (x85x)) + ((!n_n4847) & (!n_n4817) & (n_n4838) & (n_n4815) & (!x85x)) + ((!n_n4847) & (!n_n4817) & (n_n4838) & (n_n4815) & (x85x)) + ((!n_n4847) & (n_n4817) & (!n_n4838) & (!n_n4815) & (!x85x)) + ((!n_n4847) & (n_n4817) & (!n_n4838) & (!n_n4815) & (x85x)) + ((!n_n4847) & (n_n4817) & (!n_n4838) & (n_n4815) & (!x85x)) + ((!n_n4847) & (n_n4817) & (!n_n4838) & (n_n4815) & (x85x)) + ((!n_n4847) & (n_n4817) & (n_n4838) & (!n_n4815) & (!x85x)) + ((!n_n4847) & (n_n4817) & (n_n4838) & (!n_n4815) & (x85x)) + ((!n_n4847) & (n_n4817) & (n_n4838) & (n_n4815) & (!x85x)) + ((!n_n4847) & (n_n4817) & (n_n4838) & (n_n4815) & (x85x)) + ((n_n4847) & (!n_n4817) & (!n_n4838) & (!n_n4815) & (!x85x)) + ((n_n4847) & (!n_n4817) & (!n_n4838) & (!n_n4815) & (x85x)) + ((n_n4847) & (!n_n4817) & (!n_n4838) & (n_n4815) & (!x85x)) + ((n_n4847) & (!n_n4817) & (!n_n4838) & (n_n4815) & (x85x)) + ((n_n4847) & (!n_n4817) & (n_n4838) & (!n_n4815) & (!x85x)) + ((n_n4847) & (!n_n4817) & (n_n4838) & (!n_n4815) & (x85x)) + ((n_n4847) & (!n_n4817) & (n_n4838) & (n_n4815) & (!x85x)) + ((n_n4847) & (!n_n4817) & (n_n4838) & (n_n4815) & (x85x)) + ((n_n4847) & (n_n4817) & (!n_n4838) & (!n_n4815) & (!x85x)) + ((n_n4847) & (n_n4817) & (!n_n4838) & (!n_n4815) & (x85x)) + ((n_n4847) & (n_n4817) & (!n_n4838) & (n_n4815) & (!x85x)) + ((n_n4847) & (n_n4817) & (!n_n4838) & (n_n4815) & (x85x)) + ((n_n4847) & (n_n4817) & (n_n4838) & (!n_n4815) & (!x85x)) + ((n_n4847) & (n_n4817) & (n_n4838) & (!n_n4815) & (x85x)) + ((n_n4847) & (n_n4817) & (n_n4838) & (n_n4815) & (!x85x)) + ((n_n4847) & (n_n4817) & (n_n4838) & (n_n4815) & (x85x)));
	assign n_n4715 = (((!i_9_) & (n_n518) & (n_n532) & (n_n325)));
	assign n_n5225 = (((!i_9_) & (n_n518) & (n_n534) & (n_n65)));
	assign n_n5224 = (((!i_5_) & (i_3_) & (i_4_) & (x19x) & (n_n534)));
	assign x12316x = (((!n_n5046) & (!n_n5044) & (!n_n5049) & (!n_n5052) & (n_n5039)) + ((!n_n5046) & (!n_n5044) & (!n_n5049) & (n_n5052) & (!n_n5039)) + ((!n_n5046) & (!n_n5044) & (!n_n5049) & (n_n5052) & (n_n5039)) + ((!n_n5046) & (!n_n5044) & (n_n5049) & (!n_n5052) & (!n_n5039)) + ((!n_n5046) & (!n_n5044) & (n_n5049) & (!n_n5052) & (n_n5039)) + ((!n_n5046) & (!n_n5044) & (n_n5049) & (n_n5052) & (!n_n5039)) + ((!n_n5046) & (!n_n5044) & (n_n5049) & (n_n5052) & (n_n5039)) + ((!n_n5046) & (n_n5044) & (!n_n5049) & (!n_n5052) & (!n_n5039)) + ((!n_n5046) & (n_n5044) & (!n_n5049) & (!n_n5052) & (n_n5039)) + ((!n_n5046) & (n_n5044) & (!n_n5049) & (n_n5052) & (!n_n5039)) + ((!n_n5046) & (n_n5044) & (!n_n5049) & (n_n5052) & (n_n5039)) + ((!n_n5046) & (n_n5044) & (n_n5049) & (!n_n5052) & (!n_n5039)) + ((!n_n5046) & (n_n5044) & (n_n5049) & (!n_n5052) & (n_n5039)) + ((!n_n5046) & (n_n5044) & (n_n5049) & (n_n5052) & (!n_n5039)) + ((!n_n5046) & (n_n5044) & (n_n5049) & (n_n5052) & (n_n5039)) + ((n_n5046) & (!n_n5044) & (!n_n5049) & (!n_n5052) & (!n_n5039)) + ((n_n5046) & (!n_n5044) & (!n_n5049) & (!n_n5052) & (n_n5039)) + ((n_n5046) & (!n_n5044) & (!n_n5049) & (n_n5052) & (!n_n5039)) + ((n_n5046) & (!n_n5044) & (!n_n5049) & (n_n5052) & (n_n5039)) + ((n_n5046) & (!n_n5044) & (n_n5049) & (!n_n5052) & (!n_n5039)) + ((n_n5046) & (!n_n5044) & (n_n5049) & (!n_n5052) & (n_n5039)) + ((n_n5046) & (!n_n5044) & (n_n5049) & (n_n5052) & (!n_n5039)) + ((n_n5046) & (!n_n5044) & (n_n5049) & (n_n5052) & (n_n5039)) + ((n_n5046) & (n_n5044) & (!n_n5049) & (!n_n5052) & (!n_n5039)) + ((n_n5046) & (n_n5044) & (!n_n5049) & (!n_n5052) & (n_n5039)) + ((n_n5046) & (n_n5044) & (!n_n5049) & (n_n5052) & (!n_n5039)) + ((n_n5046) & (n_n5044) & (!n_n5049) & (n_n5052) & (n_n5039)) + ((n_n5046) & (n_n5044) & (n_n5049) & (!n_n5052) & (!n_n5039)) + ((n_n5046) & (n_n5044) & (n_n5049) & (!n_n5052) & (n_n5039)) + ((n_n5046) & (n_n5044) & (n_n5049) & (n_n5052) & (!n_n5039)) + ((n_n5046) & (n_n5044) & (n_n5049) & (n_n5052) & (n_n5039)));
	assign x12287x = (((!n_n5161) & (!n_n5168) & (!n_n5160) & (n_n5169)) + ((!n_n5161) & (!n_n5168) & (n_n5160) & (!n_n5169)) + ((!n_n5161) & (!n_n5168) & (n_n5160) & (n_n5169)) + ((!n_n5161) & (n_n5168) & (!n_n5160) & (!n_n5169)) + ((!n_n5161) & (n_n5168) & (!n_n5160) & (n_n5169)) + ((!n_n5161) & (n_n5168) & (n_n5160) & (!n_n5169)) + ((!n_n5161) & (n_n5168) & (n_n5160) & (n_n5169)) + ((n_n5161) & (!n_n5168) & (!n_n5160) & (!n_n5169)) + ((n_n5161) & (!n_n5168) & (!n_n5160) & (n_n5169)) + ((n_n5161) & (!n_n5168) & (n_n5160) & (!n_n5169)) + ((n_n5161) & (!n_n5168) & (n_n5160) & (n_n5169)) + ((n_n5161) & (n_n5168) & (!n_n5160) & (!n_n5169)) + ((n_n5161) & (n_n5168) & (!n_n5160) & (n_n5169)) + ((n_n5161) & (n_n5168) & (n_n5160) & (!n_n5169)) + ((n_n5161) & (n_n5168) & (n_n5160) & (n_n5169)));
	assign n_n1442 = (((!n_n5167) & (!n_n5166) & (!n_n5163) & (!x33x) & (x12287x)) + ((!n_n5167) & (!n_n5166) & (!n_n5163) & (x33x) & (!x12287x)) + ((!n_n5167) & (!n_n5166) & (!n_n5163) & (x33x) & (x12287x)) + ((!n_n5167) & (!n_n5166) & (n_n5163) & (!x33x) & (!x12287x)) + ((!n_n5167) & (!n_n5166) & (n_n5163) & (!x33x) & (x12287x)) + ((!n_n5167) & (!n_n5166) & (n_n5163) & (x33x) & (!x12287x)) + ((!n_n5167) & (!n_n5166) & (n_n5163) & (x33x) & (x12287x)) + ((!n_n5167) & (n_n5166) & (!n_n5163) & (!x33x) & (!x12287x)) + ((!n_n5167) & (n_n5166) & (!n_n5163) & (!x33x) & (x12287x)) + ((!n_n5167) & (n_n5166) & (!n_n5163) & (x33x) & (!x12287x)) + ((!n_n5167) & (n_n5166) & (!n_n5163) & (x33x) & (x12287x)) + ((!n_n5167) & (n_n5166) & (n_n5163) & (!x33x) & (!x12287x)) + ((!n_n5167) & (n_n5166) & (n_n5163) & (!x33x) & (x12287x)) + ((!n_n5167) & (n_n5166) & (n_n5163) & (x33x) & (!x12287x)) + ((!n_n5167) & (n_n5166) & (n_n5163) & (x33x) & (x12287x)) + ((n_n5167) & (!n_n5166) & (!n_n5163) & (!x33x) & (!x12287x)) + ((n_n5167) & (!n_n5166) & (!n_n5163) & (!x33x) & (x12287x)) + ((n_n5167) & (!n_n5166) & (!n_n5163) & (x33x) & (!x12287x)) + ((n_n5167) & (!n_n5166) & (!n_n5163) & (x33x) & (x12287x)) + ((n_n5167) & (!n_n5166) & (n_n5163) & (!x33x) & (!x12287x)) + ((n_n5167) & (!n_n5166) & (n_n5163) & (!x33x) & (x12287x)) + ((n_n5167) & (!n_n5166) & (n_n5163) & (x33x) & (!x12287x)) + ((n_n5167) & (!n_n5166) & (n_n5163) & (x33x) & (x12287x)) + ((n_n5167) & (n_n5166) & (!n_n5163) & (!x33x) & (!x12287x)) + ((n_n5167) & (n_n5166) & (!n_n5163) & (!x33x) & (x12287x)) + ((n_n5167) & (n_n5166) & (!n_n5163) & (x33x) & (!x12287x)) + ((n_n5167) & (n_n5166) & (!n_n5163) & (x33x) & (x12287x)) + ((n_n5167) & (n_n5166) & (n_n5163) & (!x33x) & (!x12287x)) + ((n_n5167) & (n_n5166) & (n_n5163) & (!x33x) & (x12287x)) + ((n_n5167) & (n_n5166) & (n_n5163) & (x33x) & (!x12287x)) + ((n_n5167) & (n_n5166) & (n_n5163) & (x33x) & (x12287x)));
	assign n_n5279 = (((!i_9_) & (n_n528) & (n_n491) & (n_n65)));
	assign n_n3382 = (((!x15x) & (!x11x) & (!n_n491) & (!n_n65) & (n_n5278)) + ((!x15x) & (!x11x) & (!n_n491) & (n_n65) & (n_n5278)) + ((!x15x) & (!x11x) & (n_n491) & (!n_n65) & (n_n5278)) + ((!x15x) & (!x11x) & (n_n491) & (n_n65) & (n_n5278)) + ((!x15x) & (x11x) & (!n_n491) & (!n_n65) & (n_n5278)) + ((!x15x) & (x11x) & (!n_n491) & (n_n65) & (n_n5278)) + ((!x15x) & (x11x) & (n_n491) & (!n_n65) & (n_n5278)) + ((!x15x) & (x11x) & (n_n491) & (n_n65) & (!n_n5278)) + ((!x15x) & (x11x) & (n_n491) & (n_n65) & (n_n5278)) + ((x15x) & (!x11x) & (!n_n491) & (!n_n65) & (n_n5278)) + ((x15x) & (!x11x) & (!n_n491) & (n_n65) & (n_n5278)) + ((x15x) & (!x11x) & (n_n491) & (!n_n65) & (n_n5278)) + ((x15x) & (!x11x) & (n_n491) & (n_n65) & (!n_n5278)) + ((x15x) & (!x11x) & (n_n491) & (n_n65) & (n_n5278)) + ((x15x) & (x11x) & (!n_n491) & (!n_n65) & (n_n5278)) + ((x15x) & (x11x) & (!n_n491) & (n_n65) & (n_n5278)) + ((x15x) & (x11x) & (n_n491) & (!n_n65) & (n_n5278)) + ((x15x) & (x11x) & (n_n491) & (n_n65) & (!n_n5278)) + ((x15x) & (x11x) & (n_n491) & (n_n65) & (n_n5278)));
	assign n_n4716 = (((i_9_) & (n_n518) & (n_n325) & (n_n530)));
	assign n_n1162 = (((!i_9_) & (!n_n528) & (!n_n130) & (!n_n500) & (n_n5136)) + ((!i_9_) & (!n_n528) & (!n_n130) & (n_n500) & (n_n5136)) + ((!i_9_) & (!n_n528) & (n_n130) & (!n_n500) & (n_n5136)) + ((!i_9_) & (!n_n528) & (n_n130) & (n_n500) & (n_n5136)) + ((!i_9_) & (n_n528) & (!n_n130) & (!n_n500) & (n_n5136)) + ((!i_9_) & (n_n528) & (!n_n130) & (n_n500) & (n_n5136)) + ((!i_9_) & (n_n528) & (n_n130) & (!n_n500) & (n_n5136)) + ((!i_9_) & (n_n528) & (n_n130) & (n_n500) & (!n_n5136)) + ((!i_9_) & (n_n528) & (n_n130) & (n_n500) & (n_n5136)) + ((i_9_) & (!n_n528) & (!n_n130) & (!n_n500) & (n_n5136)) + ((i_9_) & (!n_n528) & (!n_n130) & (n_n500) & (n_n5136)) + ((i_9_) & (!n_n528) & (n_n130) & (!n_n500) & (n_n5136)) + ((i_9_) & (!n_n528) & (n_n130) & (n_n500) & (n_n5136)) + ((i_9_) & (n_n528) & (!n_n130) & (!n_n500) & (n_n5136)) + ((i_9_) & (n_n528) & (!n_n130) & (n_n500) & (n_n5136)) + ((i_9_) & (n_n528) & (n_n130) & (!n_n500) & (n_n5136)) + ((i_9_) & (n_n528) & (n_n130) & (n_n500) & (!n_n5136)) + ((i_9_) & (n_n528) & (n_n130) & (n_n500) & (n_n5136)));
	assign x11563x = (((!n_n4596) & (!n_n4608) & (!n_n4606) & (!n_n4610) & (n_n4600)) + ((!n_n4596) & (!n_n4608) & (!n_n4606) & (n_n4610) & (!n_n4600)) + ((!n_n4596) & (!n_n4608) & (!n_n4606) & (n_n4610) & (n_n4600)) + ((!n_n4596) & (!n_n4608) & (n_n4606) & (!n_n4610) & (!n_n4600)) + ((!n_n4596) & (!n_n4608) & (n_n4606) & (!n_n4610) & (n_n4600)) + ((!n_n4596) & (!n_n4608) & (n_n4606) & (n_n4610) & (!n_n4600)) + ((!n_n4596) & (!n_n4608) & (n_n4606) & (n_n4610) & (n_n4600)) + ((!n_n4596) & (n_n4608) & (!n_n4606) & (!n_n4610) & (!n_n4600)) + ((!n_n4596) & (n_n4608) & (!n_n4606) & (!n_n4610) & (n_n4600)) + ((!n_n4596) & (n_n4608) & (!n_n4606) & (n_n4610) & (!n_n4600)) + ((!n_n4596) & (n_n4608) & (!n_n4606) & (n_n4610) & (n_n4600)) + ((!n_n4596) & (n_n4608) & (n_n4606) & (!n_n4610) & (!n_n4600)) + ((!n_n4596) & (n_n4608) & (n_n4606) & (!n_n4610) & (n_n4600)) + ((!n_n4596) & (n_n4608) & (n_n4606) & (n_n4610) & (!n_n4600)) + ((!n_n4596) & (n_n4608) & (n_n4606) & (n_n4610) & (n_n4600)) + ((n_n4596) & (!n_n4608) & (!n_n4606) & (!n_n4610) & (!n_n4600)) + ((n_n4596) & (!n_n4608) & (!n_n4606) & (!n_n4610) & (n_n4600)) + ((n_n4596) & (!n_n4608) & (!n_n4606) & (n_n4610) & (!n_n4600)) + ((n_n4596) & (!n_n4608) & (!n_n4606) & (n_n4610) & (n_n4600)) + ((n_n4596) & (!n_n4608) & (n_n4606) & (!n_n4610) & (!n_n4600)) + ((n_n4596) & (!n_n4608) & (n_n4606) & (!n_n4610) & (n_n4600)) + ((n_n4596) & (!n_n4608) & (n_n4606) & (n_n4610) & (!n_n4600)) + ((n_n4596) & (!n_n4608) & (n_n4606) & (n_n4610) & (n_n4600)) + ((n_n4596) & (n_n4608) & (!n_n4606) & (!n_n4610) & (!n_n4600)) + ((n_n4596) & (n_n4608) & (!n_n4606) & (!n_n4610) & (n_n4600)) + ((n_n4596) & (n_n4608) & (!n_n4606) & (n_n4610) & (!n_n4600)) + ((n_n4596) & (n_n4608) & (!n_n4606) & (n_n4610) & (n_n4600)) + ((n_n4596) & (n_n4608) & (n_n4606) & (!n_n4610) & (!n_n4600)) + ((n_n4596) & (n_n4608) & (n_n4606) & (!n_n4610) & (n_n4600)) + ((n_n4596) & (n_n4608) & (n_n4606) & (n_n4610) & (!n_n4600)) + ((n_n4596) & (n_n4608) & (n_n4606) & (n_n4610) & (n_n4600)));
	assign n_n1100 = (((!x23x) & (!x583x) & (!n_n4598) & (!x256x) & (x11563x)) + ((!x23x) & (!x583x) & (!n_n4598) & (x256x) & (!x11563x)) + ((!x23x) & (!x583x) & (!n_n4598) & (x256x) & (x11563x)) + ((!x23x) & (!x583x) & (n_n4598) & (!x256x) & (!x11563x)) + ((!x23x) & (!x583x) & (n_n4598) & (!x256x) & (x11563x)) + ((!x23x) & (!x583x) & (n_n4598) & (x256x) & (!x11563x)) + ((!x23x) & (!x583x) & (n_n4598) & (x256x) & (x11563x)) + ((!x23x) & (x583x) & (!n_n4598) & (!x256x) & (x11563x)) + ((!x23x) & (x583x) & (!n_n4598) & (x256x) & (!x11563x)) + ((!x23x) & (x583x) & (!n_n4598) & (x256x) & (x11563x)) + ((!x23x) & (x583x) & (n_n4598) & (!x256x) & (!x11563x)) + ((!x23x) & (x583x) & (n_n4598) & (!x256x) & (x11563x)) + ((!x23x) & (x583x) & (n_n4598) & (x256x) & (!x11563x)) + ((!x23x) & (x583x) & (n_n4598) & (x256x) & (x11563x)) + ((x23x) & (!x583x) & (!n_n4598) & (!x256x) & (x11563x)) + ((x23x) & (!x583x) & (!n_n4598) & (x256x) & (!x11563x)) + ((x23x) & (!x583x) & (!n_n4598) & (x256x) & (x11563x)) + ((x23x) & (!x583x) & (n_n4598) & (!x256x) & (!x11563x)) + ((x23x) & (!x583x) & (n_n4598) & (!x256x) & (x11563x)) + ((x23x) & (!x583x) & (n_n4598) & (x256x) & (!x11563x)) + ((x23x) & (!x583x) & (n_n4598) & (x256x) & (x11563x)) + ((x23x) & (x583x) & (!n_n4598) & (!x256x) & (!x11563x)) + ((x23x) & (x583x) & (!n_n4598) & (!x256x) & (x11563x)) + ((x23x) & (x583x) & (!n_n4598) & (x256x) & (!x11563x)) + ((x23x) & (x583x) & (!n_n4598) & (x256x) & (x11563x)) + ((x23x) & (x583x) & (n_n4598) & (!x256x) & (!x11563x)) + ((x23x) & (x583x) & (n_n4598) & (!x256x) & (x11563x)) + ((x23x) & (x583x) & (n_n4598) & (x256x) & (!x11563x)) + ((x23x) & (x583x) & (n_n4598) & (x256x) & (x11563x)));
	assign x71x = (((!i_9_) & (n_n524) & (n_n473) & (n_n325) & (!n_n522)) + ((!i_9_) & (n_n524) & (n_n473) & (n_n325) & (n_n522)) + ((i_9_) & (!n_n524) & (n_n473) & (n_n325) & (n_n522)) + ((i_9_) & (n_n524) & (n_n473) & (n_n325) & (n_n522)));
	assign x11913x = (((!x15x) & (!n_n130) & (!n_n500) & (!n_n5128) & (n_n1162)) + ((!x15x) & (!n_n130) & (!n_n500) & (n_n5128) & (!n_n1162)) + ((!x15x) & (!n_n130) & (!n_n500) & (n_n5128) & (n_n1162)) + ((!x15x) & (!n_n130) & (n_n500) & (!n_n5128) & (n_n1162)) + ((!x15x) & (!n_n130) & (n_n500) & (n_n5128) & (!n_n1162)) + ((!x15x) & (!n_n130) & (n_n500) & (n_n5128) & (n_n1162)) + ((!x15x) & (n_n130) & (!n_n500) & (!n_n5128) & (n_n1162)) + ((!x15x) & (n_n130) & (!n_n500) & (n_n5128) & (!n_n1162)) + ((!x15x) & (n_n130) & (!n_n500) & (n_n5128) & (n_n1162)) + ((!x15x) & (n_n130) & (n_n500) & (!n_n5128) & (n_n1162)) + ((!x15x) & (n_n130) & (n_n500) & (n_n5128) & (!n_n1162)) + ((!x15x) & (n_n130) & (n_n500) & (n_n5128) & (n_n1162)) + ((x15x) & (!n_n130) & (!n_n500) & (!n_n5128) & (n_n1162)) + ((x15x) & (!n_n130) & (!n_n500) & (n_n5128) & (!n_n1162)) + ((x15x) & (!n_n130) & (!n_n500) & (n_n5128) & (n_n1162)) + ((x15x) & (!n_n130) & (n_n500) & (!n_n5128) & (n_n1162)) + ((x15x) & (!n_n130) & (n_n500) & (n_n5128) & (!n_n1162)) + ((x15x) & (!n_n130) & (n_n500) & (n_n5128) & (n_n1162)) + ((x15x) & (n_n130) & (!n_n500) & (!n_n5128) & (n_n1162)) + ((x15x) & (n_n130) & (!n_n500) & (n_n5128) & (!n_n1162)) + ((x15x) & (n_n130) & (!n_n500) & (n_n5128) & (n_n1162)) + ((x15x) & (n_n130) & (n_n500) & (!n_n5128) & (!n_n1162)) + ((x15x) & (n_n130) & (n_n500) & (!n_n5128) & (n_n1162)) + ((x15x) & (n_n130) & (n_n500) & (n_n5128) & (!n_n1162)) + ((x15x) & (n_n130) & (n_n500) & (n_n5128) & (n_n1162)));
	assign n_n1059 = (((!n_n5124) & (!n_n5126) & (!x155x) & (x11913x)) + ((!n_n5124) & (!n_n5126) & (x155x) & (!x11913x)) + ((!n_n5124) & (!n_n5126) & (x155x) & (x11913x)) + ((!n_n5124) & (n_n5126) & (!x155x) & (!x11913x)) + ((!n_n5124) & (n_n5126) & (!x155x) & (x11913x)) + ((!n_n5124) & (n_n5126) & (x155x) & (!x11913x)) + ((!n_n5124) & (n_n5126) & (x155x) & (x11913x)) + ((n_n5124) & (!n_n5126) & (!x155x) & (!x11913x)) + ((n_n5124) & (!n_n5126) & (!x155x) & (x11913x)) + ((n_n5124) & (!n_n5126) & (x155x) & (!x11913x)) + ((n_n5124) & (!n_n5126) & (x155x) & (x11913x)) + ((n_n5124) & (n_n5126) & (!x155x) & (!x11913x)) + ((n_n5124) & (n_n5126) & (!x155x) & (x11913x)) + ((n_n5124) & (n_n5126) & (x155x) & (!x11913x)) + ((n_n5124) & (n_n5126) & (x155x) & (x11913x)));
	assign x11915x = (((!n_n532) & (!n_n509) & (!x12x) & (!n_n530) & (n_n5115)) + ((!n_n532) & (!n_n509) & (!x12x) & (n_n530) & (n_n5115)) + ((!n_n532) & (!n_n509) & (x12x) & (!n_n530) & (n_n5115)) + ((!n_n532) & (!n_n509) & (x12x) & (n_n530) & (n_n5115)) + ((!n_n532) & (n_n509) & (!x12x) & (!n_n530) & (n_n5115)) + ((!n_n532) & (n_n509) & (!x12x) & (n_n530) & (n_n5115)) + ((!n_n532) & (n_n509) & (x12x) & (!n_n530) & (n_n5115)) + ((!n_n532) & (n_n509) & (x12x) & (n_n530) & (!n_n5115)) + ((!n_n532) & (n_n509) & (x12x) & (n_n530) & (n_n5115)) + ((n_n532) & (!n_n509) & (!x12x) & (!n_n530) & (n_n5115)) + ((n_n532) & (!n_n509) & (!x12x) & (n_n530) & (n_n5115)) + ((n_n532) & (!n_n509) & (x12x) & (!n_n530) & (n_n5115)) + ((n_n532) & (!n_n509) & (x12x) & (n_n530) & (n_n5115)) + ((n_n532) & (n_n509) & (!x12x) & (!n_n530) & (n_n5115)) + ((n_n532) & (n_n509) & (!x12x) & (n_n530) & (n_n5115)) + ((n_n532) & (n_n509) & (x12x) & (!n_n530) & (!n_n5115)) + ((n_n532) & (n_n509) & (x12x) & (!n_n530) & (n_n5115)) + ((n_n532) & (n_n509) & (x12x) & (n_n530) & (!n_n5115)) + ((n_n532) & (n_n509) & (x12x) & (n_n530) & (n_n5115)));
	assign x28x = (((!n_n5111) & (!n_n5110) & (!n_n5114) & (!n_n5116) & (n_n5115)) + ((!n_n5111) & (!n_n5110) & (!n_n5114) & (n_n5116) & (!n_n5115)) + ((!n_n5111) & (!n_n5110) & (!n_n5114) & (n_n5116) & (n_n5115)) + ((!n_n5111) & (!n_n5110) & (n_n5114) & (!n_n5116) & (!n_n5115)) + ((!n_n5111) & (!n_n5110) & (n_n5114) & (!n_n5116) & (n_n5115)) + ((!n_n5111) & (!n_n5110) & (n_n5114) & (n_n5116) & (!n_n5115)) + ((!n_n5111) & (!n_n5110) & (n_n5114) & (n_n5116) & (n_n5115)) + ((!n_n5111) & (n_n5110) & (!n_n5114) & (!n_n5116) & (!n_n5115)) + ((!n_n5111) & (n_n5110) & (!n_n5114) & (!n_n5116) & (n_n5115)) + ((!n_n5111) & (n_n5110) & (!n_n5114) & (n_n5116) & (!n_n5115)) + ((!n_n5111) & (n_n5110) & (!n_n5114) & (n_n5116) & (n_n5115)) + ((!n_n5111) & (n_n5110) & (n_n5114) & (!n_n5116) & (!n_n5115)) + ((!n_n5111) & (n_n5110) & (n_n5114) & (!n_n5116) & (n_n5115)) + ((!n_n5111) & (n_n5110) & (n_n5114) & (n_n5116) & (!n_n5115)) + ((!n_n5111) & (n_n5110) & (n_n5114) & (n_n5116) & (n_n5115)) + ((n_n5111) & (!n_n5110) & (!n_n5114) & (!n_n5116) & (!n_n5115)) + ((n_n5111) & (!n_n5110) & (!n_n5114) & (!n_n5116) & (n_n5115)) + ((n_n5111) & (!n_n5110) & (!n_n5114) & (n_n5116) & (!n_n5115)) + ((n_n5111) & (!n_n5110) & (!n_n5114) & (n_n5116) & (n_n5115)) + ((n_n5111) & (!n_n5110) & (n_n5114) & (!n_n5116) & (!n_n5115)) + ((n_n5111) & (!n_n5110) & (n_n5114) & (!n_n5116) & (n_n5115)) + ((n_n5111) & (!n_n5110) & (n_n5114) & (n_n5116) & (!n_n5115)) + ((n_n5111) & (!n_n5110) & (n_n5114) & (n_n5116) & (n_n5115)) + ((n_n5111) & (n_n5110) & (!n_n5114) & (!n_n5116) & (!n_n5115)) + ((n_n5111) & (n_n5110) & (!n_n5114) & (!n_n5116) & (n_n5115)) + ((n_n5111) & (n_n5110) & (!n_n5114) & (n_n5116) & (!n_n5115)) + ((n_n5111) & (n_n5110) & (!n_n5114) & (n_n5116) & (n_n5115)) + ((n_n5111) & (n_n5110) & (n_n5114) & (!n_n5116) & (!n_n5115)) + ((n_n5111) & (n_n5110) & (n_n5114) & (!n_n5116) & (n_n5115)) + ((n_n5111) & (n_n5110) & (n_n5114) & (n_n5116) & (!n_n5115)) + ((n_n5111) & (n_n5110) & (n_n5114) & (n_n5116) & (n_n5115)));
	assign n_n1060 = (((!n_n5112) & (!n_n5120) & (!n_n5117) & (!n_n5121) & (x28x)) + ((!n_n5112) & (!n_n5120) & (!n_n5117) & (n_n5121) & (!x28x)) + ((!n_n5112) & (!n_n5120) & (!n_n5117) & (n_n5121) & (x28x)) + ((!n_n5112) & (!n_n5120) & (n_n5117) & (!n_n5121) & (!x28x)) + ((!n_n5112) & (!n_n5120) & (n_n5117) & (!n_n5121) & (x28x)) + ((!n_n5112) & (!n_n5120) & (n_n5117) & (n_n5121) & (!x28x)) + ((!n_n5112) & (!n_n5120) & (n_n5117) & (n_n5121) & (x28x)) + ((!n_n5112) & (n_n5120) & (!n_n5117) & (!n_n5121) & (!x28x)) + ((!n_n5112) & (n_n5120) & (!n_n5117) & (!n_n5121) & (x28x)) + ((!n_n5112) & (n_n5120) & (!n_n5117) & (n_n5121) & (!x28x)) + ((!n_n5112) & (n_n5120) & (!n_n5117) & (n_n5121) & (x28x)) + ((!n_n5112) & (n_n5120) & (n_n5117) & (!n_n5121) & (!x28x)) + ((!n_n5112) & (n_n5120) & (n_n5117) & (!n_n5121) & (x28x)) + ((!n_n5112) & (n_n5120) & (n_n5117) & (n_n5121) & (!x28x)) + ((!n_n5112) & (n_n5120) & (n_n5117) & (n_n5121) & (x28x)) + ((n_n5112) & (!n_n5120) & (!n_n5117) & (!n_n5121) & (!x28x)) + ((n_n5112) & (!n_n5120) & (!n_n5117) & (!n_n5121) & (x28x)) + ((n_n5112) & (!n_n5120) & (!n_n5117) & (n_n5121) & (!x28x)) + ((n_n5112) & (!n_n5120) & (!n_n5117) & (n_n5121) & (x28x)) + ((n_n5112) & (!n_n5120) & (n_n5117) & (!n_n5121) & (!x28x)) + ((n_n5112) & (!n_n5120) & (n_n5117) & (!n_n5121) & (x28x)) + ((n_n5112) & (!n_n5120) & (n_n5117) & (n_n5121) & (!x28x)) + ((n_n5112) & (!n_n5120) & (n_n5117) & (n_n5121) & (x28x)) + ((n_n5112) & (n_n5120) & (!n_n5117) & (!n_n5121) & (!x28x)) + ((n_n5112) & (n_n5120) & (!n_n5117) & (!n_n5121) & (x28x)) + ((n_n5112) & (n_n5120) & (!n_n5117) & (n_n5121) & (!x28x)) + ((n_n5112) & (n_n5120) & (!n_n5117) & (n_n5121) & (x28x)) + ((n_n5112) & (n_n5120) & (n_n5117) & (!n_n5121) & (!x28x)) + ((n_n5112) & (n_n5120) & (n_n5117) & (!n_n5121) & (x28x)) + ((n_n5112) & (n_n5120) & (n_n5117) & (n_n5121) & (!x28x)) + ((n_n5112) & (n_n5120) & (n_n5117) & (n_n5121) & (x28x)));
	assign n_n4446 = (((i_9_) & (n_n455) & (n_n528) & (n_n535)));
	assign n_n4961 = (((!i_9_) & (n_n526) & (n_n535) & (n_n195)));
	assign n_n5194 = (((i_7_) & (!i_8_) & (i_6_) & (x12x) & (n_n464)));
	assign n_n5259 = (((!i_9_) & (n_n532) & (n_n500) & (n_n65)));
	assign n_n5265 = (((!i_9_) & (n_n526) & (n_n500) & (n_n65)));
	assign n_n5271 = (((!i_5_) & (i_3_) & (!i_4_) & (x23x) & (n_n65)));
	assign n_n4537 = (((!i_9_) & (n_n455) & (n_n473) & (n_n534)));
	assign x11532x = (((!i_9_) & (n_n455) & (n_n473) & (n_n532)) + ((i_9_) & (n_n455) & (n_n473) & (n_n532)));
	assign n_n1648 = (((!x21x) & (!n_n390) & (!x20x) & (!n_n500) & (n_n4628)) + ((!x21x) & (!n_n390) & (!x20x) & (n_n500) & (n_n4628)) + ((!x21x) & (!n_n390) & (x20x) & (!n_n500) & (n_n4628)) + ((!x21x) & (!n_n390) & (x20x) & (n_n500) & (n_n4628)) + ((!x21x) & (n_n390) & (!x20x) & (!n_n500) & (n_n4628)) + ((!x21x) & (n_n390) & (!x20x) & (n_n500) & (n_n4628)) + ((!x21x) & (n_n390) & (x20x) & (!n_n500) & (n_n4628)) + ((!x21x) & (n_n390) & (x20x) & (n_n500) & (!n_n4628)) + ((!x21x) & (n_n390) & (x20x) & (n_n500) & (n_n4628)) + ((x21x) & (!n_n390) & (!x20x) & (!n_n500) & (n_n4628)) + ((x21x) & (!n_n390) & (!x20x) & (n_n500) & (n_n4628)) + ((x21x) & (!n_n390) & (x20x) & (!n_n500) & (n_n4628)) + ((x21x) & (!n_n390) & (x20x) & (n_n500) & (n_n4628)) + ((x21x) & (n_n390) & (!x20x) & (!n_n500) & (n_n4628)) + ((x21x) & (n_n390) & (!x20x) & (n_n500) & (!n_n4628)) + ((x21x) & (n_n390) & (!x20x) & (n_n500) & (n_n4628)) + ((x21x) & (n_n390) & (x20x) & (!n_n500) & (n_n4628)) + ((x21x) & (n_n390) & (x20x) & (n_n500) & (!n_n4628)) + ((x21x) & (n_n390) & (x20x) & (n_n500) & (n_n4628)));
	assign x13204x = (((!n_n4911) & (!n_n4912) & (!n_n4914) & (!n_n4917) & (n_n4915)) + ((!n_n4911) & (!n_n4912) & (!n_n4914) & (n_n4917) & (!n_n4915)) + ((!n_n4911) & (!n_n4912) & (!n_n4914) & (n_n4917) & (n_n4915)) + ((!n_n4911) & (!n_n4912) & (n_n4914) & (!n_n4917) & (!n_n4915)) + ((!n_n4911) & (!n_n4912) & (n_n4914) & (!n_n4917) & (n_n4915)) + ((!n_n4911) & (!n_n4912) & (n_n4914) & (n_n4917) & (!n_n4915)) + ((!n_n4911) & (!n_n4912) & (n_n4914) & (n_n4917) & (n_n4915)) + ((!n_n4911) & (n_n4912) & (!n_n4914) & (!n_n4917) & (!n_n4915)) + ((!n_n4911) & (n_n4912) & (!n_n4914) & (!n_n4917) & (n_n4915)) + ((!n_n4911) & (n_n4912) & (!n_n4914) & (n_n4917) & (!n_n4915)) + ((!n_n4911) & (n_n4912) & (!n_n4914) & (n_n4917) & (n_n4915)) + ((!n_n4911) & (n_n4912) & (n_n4914) & (!n_n4917) & (!n_n4915)) + ((!n_n4911) & (n_n4912) & (n_n4914) & (!n_n4917) & (n_n4915)) + ((!n_n4911) & (n_n4912) & (n_n4914) & (n_n4917) & (!n_n4915)) + ((!n_n4911) & (n_n4912) & (n_n4914) & (n_n4917) & (n_n4915)) + ((n_n4911) & (!n_n4912) & (!n_n4914) & (!n_n4917) & (!n_n4915)) + ((n_n4911) & (!n_n4912) & (!n_n4914) & (!n_n4917) & (n_n4915)) + ((n_n4911) & (!n_n4912) & (!n_n4914) & (n_n4917) & (!n_n4915)) + ((n_n4911) & (!n_n4912) & (!n_n4914) & (n_n4917) & (n_n4915)) + ((n_n4911) & (!n_n4912) & (n_n4914) & (!n_n4917) & (!n_n4915)) + ((n_n4911) & (!n_n4912) & (n_n4914) & (!n_n4917) & (n_n4915)) + ((n_n4911) & (!n_n4912) & (n_n4914) & (n_n4917) & (!n_n4915)) + ((n_n4911) & (!n_n4912) & (n_n4914) & (n_n4917) & (n_n4915)) + ((n_n4911) & (n_n4912) & (!n_n4914) & (!n_n4917) & (!n_n4915)) + ((n_n4911) & (n_n4912) & (!n_n4914) & (!n_n4917) & (n_n4915)) + ((n_n4911) & (n_n4912) & (!n_n4914) & (n_n4917) & (!n_n4915)) + ((n_n4911) & (n_n4912) & (!n_n4914) & (n_n4917) & (n_n4915)) + ((n_n4911) & (n_n4912) & (n_n4914) & (!n_n4917) & (!n_n4915)) + ((n_n4911) & (n_n4912) & (n_n4914) & (!n_n4917) & (n_n4915)) + ((n_n4911) & (n_n4912) & (n_n4914) & (n_n4917) & (!n_n4915)) + ((n_n4911) & (n_n4912) & (n_n4914) & (n_n4917) & (n_n4915)));
	assign x13405x = (((!n_n5044) & (!n_n5045) & (!n_n5053) & (!n_n5052) & (n_n5051)) + ((!n_n5044) & (!n_n5045) & (!n_n5053) & (n_n5052) & (!n_n5051)) + ((!n_n5044) & (!n_n5045) & (!n_n5053) & (n_n5052) & (n_n5051)) + ((!n_n5044) & (!n_n5045) & (n_n5053) & (!n_n5052) & (!n_n5051)) + ((!n_n5044) & (!n_n5045) & (n_n5053) & (!n_n5052) & (n_n5051)) + ((!n_n5044) & (!n_n5045) & (n_n5053) & (n_n5052) & (!n_n5051)) + ((!n_n5044) & (!n_n5045) & (n_n5053) & (n_n5052) & (n_n5051)) + ((!n_n5044) & (n_n5045) & (!n_n5053) & (!n_n5052) & (!n_n5051)) + ((!n_n5044) & (n_n5045) & (!n_n5053) & (!n_n5052) & (n_n5051)) + ((!n_n5044) & (n_n5045) & (!n_n5053) & (n_n5052) & (!n_n5051)) + ((!n_n5044) & (n_n5045) & (!n_n5053) & (n_n5052) & (n_n5051)) + ((!n_n5044) & (n_n5045) & (n_n5053) & (!n_n5052) & (!n_n5051)) + ((!n_n5044) & (n_n5045) & (n_n5053) & (!n_n5052) & (n_n5051)) + ((!n_n5044) & (n_n5045) & (n_n5053) & (n_n5052) & (!n_n5051)) + ((!n_n5044) & (n_n5045) & (n_n5053) & (n_n5052) & (n_n5051)) + ((n_n5044) & (!n_n5045) & (!n_n5053) & (!n_n5052) & (!n_n5051)) + ((n_n5044) & (!n_n5045) & (!n_n5053) & (!n_n5052) & (n_n5051)) + ((n_n5044) & (!n_n5045) & (!n_n5053) & (n_n5052) & (!n_n5051)) + ((n_n5044) & (!n_n5045) & (!n_n5053) & (n_n5052) & (n_n5051)) + ((n_n5044) & (!n_n5045) & (n_n5053) & (!n_n5052) & (!n_n5051)) + ((n_n5044) & (!n_n5045) & (n_n5053) & (!n_n5052) & (n_n5051)) + ((n_n5044) & (!n_n5045) & (n_n5053) & (n_n5052) & (!n_n5051)) + ((n_n5044) & (!n_n5045) & (n_n5053) & (n_n5052) & (n_n5051)) + ((n_n5044) & (n_n5045) & (!n_n5053) & (!n_n5052) & (!n_n5051)) + ((n_n5044) & (n_n5045) & (!n_n5053) & (!n_n5052) & (n_n5051)) + ((n_n5044) & (n_n5045) & (!n_n5053) & (n_n5052) & (!n_n5051)) + ((n_n5044) & (n_n5045) & (!n_n5053) & (n_n5052) & (n_n5051)) + ((n_n5044) & (n_n5045) & (n_n5053) & (!n_n5052) & (!n_n5051)) + ((n_n5044) & (n_n5045) & (n_n5053) & (!n_n5052) & (n_n5051)) + ((n_n5044) & (n_n5045) & (n_n5053) & (n_n5052) & (!n_n5051)) + ((n_n5044) & (n_n5045) & (n_n5053) & (n_n5052) & (n_n5051)));
	assign x22123x = (((!x25x) & (!x496x) & (!n_n4423) & (!x84x) & (!n_n4428)) + ((!x25x) & (x496x) & (!n_n4423) & (!x84x) & (!n_n4428)) + ((x25x) & (!x496x) & (!n_n4423) & (!x84x) & (!n_n4428)));
	assign x13438x = (((!n_n4430) & (!n_n4424) & (!n_n4421) & (!n_n4429) & (!x22123x)) + ((!n_n4430) & (!n_n4424) & (!n_n4421) & (n_n4429) & (!x22123x)) + ((!n_n4430) & (!n_n4424) & (!n_n4421) & (n_n4429) & (x22123x)) + ((!n_n4430) & (!n_n4424) & (n_n4421) & (!n_n4429) & (!x22123x)) + ((!n_n4430) & (!n_n4424) & (n_n4421) & (!n_n4429) & (x22123x)) + ((!n_n4430) & (!n_n4424) & (n_n4421) & (n_n4429) & (!x22123x)) + ((!n_n4430) & (!n_n4424) & (n_n4421) & (n_n4429) & (x22123x)) + ((!n_n4430) & (n_n4424) & (!n_n4421) & (!n_n4429) & (!x22123x)) + ((!n_n4430) & (n_n4424) & (!n_n4421) & (!n_n4429) & (x22123x)) + ((!n_n4430) & (n_n4424) & (!n_n4421) & (n_n4429) & (!x22123x)) + ((!n_n4430) & (n_n4424) & (!n_n4421) & (n_n4429) & (x22123x)) + ((!n_n4430) & (n_n4424) & (n_n4421) & (!n_n4429) & (!x22123x)) + ((!n_n4430) & (n_n4424) & (n_n4421) & (!n_n4429) & (x22123x)) + ((!n_n4430) & (n_n4424) & (n_n4421) & (n_n4429) & (!x22123x)) + ((!n_n4430) & (n_n4424) & (n_n4421) & (n_n4429) & (x22123x)) + ((n_n4430) & (!n_n4424) & (!n_n4421) & (!n_n4429) & (!x22123x)) + ((n_n4430) & (!n_n4424) & (!n_n4421) & (!n_n4429) & (x22123x)) + ((n_n4430) & (!n_n4424) & (!n_n4421) & (n_n4429) & (!x22123x)) + ((n_n4430) & (!n_n4424) & (!n_n4421) & (n_n4429) & (x22123x)) + ((n_n4430) & (!n_n4424) & (n_n4421) & (!n_n4429) & (!x22123x)) + ((n_n4430) & (!n_n4424) & (n_n4421) & (!n_n4429) & (x22123x)) + ((n_n4430) & (!n_n4424) & (n_n4421) & (n_n4429) & (!x22123x)) + ((n_n4430) & (!n_n4424) & (n_n4421) & (n_n4429) & (x22123x)) + ((n_n4430) & (n_n4424) & (!n_n4421) & (!n_n4429) & (!x22123x)) + ((n_n4430) & (n_n4424) & (!n_n4421) & (!n_n4429) & (x22123x)) + ((n_n4430) & (n_n4424) & (!n_n4421) & (n_n4429) & (!x22123x)) + ((n_n4430) & (n_n4424) & (!n_n4421) & (n_n4429) & (x22123x)) + ((n_n4430) & (n_n4424) & (n_n4421) & (!n_n4429) & (!x22123x)) + ((n_n4430) & (n_n4424) & (n_n4421) & (!n_n4429) & (x22123x)) + ((n_n4430) & (n_n4424) & (n_n4421) & (n_n4429) & (!x22123x)) + ((n_n4430) & (n_n4424) & (n_n4421) & (n_n4429) & (x22123x)));
	assign n_n4094 = (((!x323x) & (!n_n4441) & (!n_n4449) & (!x470x) & (x421x)) + ((!x323x) & (!n_n4441) & (!n_n4449) & (x470x) & (!x421x)) + ((!x323x) & (!n_n4441) & (!n_n4449) & (x470x) & (x421x)) + ((!x323x) & (!n_n4441) & (n_n4449) & (!x470x) & (!x421x)) + ((!x323x) & (!n_n4441) & (n_n4449) & (!x470x) & (x421x)) + ((!x323x) & (!n_n4441) & (n_n4449) & (x470x) & (!x421x)) + ((!x323x) & (!n_n4441) & (n_n4449) & (x470x) & (x421x)) + ((!x323x) & (n_n4441) & (!n_n4449) & (!x470x) & (!x421x)) + ((!x323x) & (n_n4441) & (!n_n4449) & (!x470x) & (x421x)) + ((!x323x) & (n_n4441) & (!n_n4449) & (x470x) & (!x421x)) + ((!x323x) & (n_n4441) & (!n_n4449) & (x470x) & (x421x)) + ((!x323x) & (n_n4441) & (n_n4449) & (!x470x) & (!x421x)) + ((!x323x) & (n_n4441) & (n_n4449) & (!x470x) & (x421x)) + ((!x323x) & (n_n4441) & (n_n4449) & (x470x) & (!x421x)) + ((!x323x) & (n_n4441) & (n_n4449) & (x470x) & (x421x)) + ((x323x) & (!n_n4441) & (!n_n4449) & (!x470x) & (!x421x)) + ((x323x) & (!n_n4441) & (!n_n4449) & (!x470x) & (x421x)) + ((x323x) & (!n_n4441) & (!n_n4449) & (x470x) & (!x421x)) + ((x323x) & (!n_n4441) & (!n_n4449) & (x470x) & (x421x)) + ((x323x) & (!n_n4441) & (n_n4449) & (!x470x) & (!x421x)) + ((x323x) & (!n_n4441) & (n_n4449) & (!x470x) & (x421x)) + ((x323x) & (!n_n4441) & (n_n4449) & (x470x) & (!x421x)) + ((x323x) & (!n_n4441) & (n_n4449) & (x470x) & (x421x)) + ((x323x) & (n_n4441) & (!n_n4449) & (!x470x) & (!x421x)) + ((x323x) & (n_n4441) & (!n_n4449) & (!x470x) & (x421x)) + ((x323x) & (n_n4441) & (!n_n4449) & (x470x) & (!x421x)) + ((x323x) & (n_n4441) & (!n_n4449) & (x470x) & (x421x)) + ((x323x) & (n_n4441) & (n_n4449) & (!x470x) & (!x421x)) + ((x323x) & (n_n4441) & (n_n4449) & (!x470x) & (x421x)) + ((x323x) & (n_n4441) & (n_n4449) & (x470x) & (!x421x)) + ((x323x) & (n_n4441) & (n_n4449) & (x470x) & (x421x)));
	assign n_n4020 = (((!n_n4095) & (!x13438x) & (n_n4094)) + ((!n_n4095) & (x13438x) & (!n_n4094)) + ((!n_n4095) & (x13438x) & (n_n4094)) + ((n_n4095) & (!x13438x) & (!n_n4094)) + ((n_n4095) & (!x13438x) & (n_n4094)) + ((n_n4095) & (x13438x) & (!n_n4094)) + ((n_n4095) & (x13438x) & (n_n4094)));
	assign x13471x = (((!n_n4560) & (!n_n4569) & (!x471x) & (x91x)) + ((!n_n4560) & (!n_n4569) & (x471x) & (!x91x)) + ((!n_n4560) & (!n_n4569) & (x471x) & (x91x)) + ((!n_n4560) & (n_n4569) & (!x471x) & (!x91x)) + ((!n_n4560) & (n_n4569) & (!x471x) & (x91x)) + ((!n_n4560) & (n_n4569) & (x471x) & (!x91x)) + ((!n_n4560) & (n_n4569) & (x471x) & (x91x)) + ((n_n4560) & (!n_n4569) & (!x471x) & (!x91x)) + ((n_n4560) & (!n_n4569) & (!x471x) & (x91x)) + ((n_n4560) & (!n_n4569) & (x471x) & (!x91x)) + ((n_n4560) & (!n_n4569) & (x471x) & (x91x)) + ((n_n4560) & (n_n4569) & (!x471x) & (!x91x)) + ((n_n4560) & (n_n4569) & (!x471x) & (x91x)) + ((n_n4560) & (n_n4569) & (x471x) & (!x91x)) + ((n_n4560) & (n_n4569) & (x471x) & (x91x)));
	assign n_n4086 = (((!n_n4554) & (!n_n4541) & (!n_n4545) & (!x13091x) & (!x22207x)) + ((!n_n4554) & (!n_n4541) & (!n_n4545) & (x13091x) & (!x22207x)) + ((!n_n4554) & (!n_n4541) & (!n_n4545) & (x13091x) & (x22207x)) + ((!n_n4554) & (!n_n4541) & (n_n4545) & (!x13091x) & (!x22207x)) + ((!n_n4554) & (!n_n4541) & (n_n4545) & (!x13091x) & (x22207x)) + ((!n_n4554) & (!n_n4541) & (n_n4545) & (x13091x) & (!x22207x)) + ((!n_n4554) & (!n_n4541) & (n_n4545) & (x13091x) & (x22207x)) + ((!n_n4554) & (n_n4541) & (!n_n4545) & (!x13091x) & (!x22207x)) + ((!n_n4554) & (n_n4541) & (!n_n4545) & (!x13091x) & (x22207x)) + ((!n_n4554) & (n_n4541) & (!n_n4545) & (x13091x) & (!x22207x)) + ((!n_n4554) & (n_n4541) & (!n_n4545) & (x13091x) & (x22207x)) + ((!n_n4554) & (n_n4541) & (n_n4545) & (!x13091x) & (!x22207x)) + ((!n_n4554) & (n_n4541) & (n_n4545) & (!x13091x) & (x22207x)) + ((!n_n4554) & (n_n4541) & (n_n4545) & (x13091x) & (!x22207x)) + ((!n_n4554) & (n_n4541) & (n_n4545) & (x13091x) & (x22207x)) + ((n_n4554) & (!n_n4541) & (!n_n4545) & (!x13091x) & (!x22207x)) + ((n_n4554) & (!n_n4541) & (!n_n4545) & (!x13091x) & (x22207x)) + ((n_n4554) & (!n_n4541) & (!n_n4545) & (x13091x) & (!x22207x)) + ((n_n4554) & (!n_n4541) & (!n_n4545) & (x13091x) & (x22207x)) + ((n_n4554) & (!n_n4541) & (n_n4545) & (!x13091x) & (!x22207x)) + ((n_n4554) & (!n_n4541) & (n_n4545) & (!x13091x) & (x22207x)) + ((n_n4554) & (!n_n4541) & (n_n4545) & (x13091x) & (!x22207x)) + ((n_n4554) & (!n_n4541) & (n_n4545) & (x13091x) & (x22207x)) + ((n_n4554) & (n_n4541) & (!n_n4545) & (!x13091x) & (!x22207x)) + ((n_n4554) & (n_n4541) & (!n_n4545) & (!x13091x) & (x22207x)) + ((n_n4554) & (n_n4541) & (!n_n4545) & (x13091x) & (!x22207x)) + ((n_n4554) & (n_n4541) & (!n_n4545) & (x13091x) & (x22207x)) + ((n_n4554) & (n_n4541) & (n_n4545) & (!x13091x) & (!x22207x)) + ((n_n4554) & (n_n4541) & (n_n4545) & (!x13091x) & (x22207x)) + ((n_n4554) & (n_n4541) & (n_n4545) & (x13091x) & (!x22207x)) + ((n_n4554) & (n_n4541) & (n_n4545) & (x13091x) & (x22207x)));
	assign x13480x = (((!n_n4533) & (!n_n4536) & (!n_n4243) & (!x379x) & (x13477x)) + ((!n_n4533) & (!n_n4536) & (!n_n4243) & (x379x) & (!x13477x)) + ((!n_n4533) & (!n_n4536) & (!n_n4243) & (x379x) & (x13477x)) + ((!n_n4533) & (!n_n4536) & (n_n4243) & (!x379x) & (!x13477x)) + ((!n_n4533) & (!n_n4536) & (n_n4243) & (!x379x) & (x13477x)) + ((!n_n4533) & (!n_n4536) & (n_n4243) & (x379x) & (!x13477x)) + ((!n_n4533) & (!n_n4536) & (n_n4243) & (x379x) & (x13477x)) + ((!n_n4533) & (n_n4536) & (!n_n4243) & (!x379x) & (!x13477x)) + ((!n_n4533) & (n_n4536) & (!n_n4243) & (!x379x) & (x13477x)) + ((!n_n4533) & (n_n4536) & (!n_n4243) & (x379x) & (!x13477x)) + ((!n_n4533) & (n_n4536) & (!n_n4243) & (x379x) & (x13477x)) + ((!n_n4533) & (n_n4536) & (n_n4243) & (!x379x) & (!x13477x)) + ((!n_n4533) & (n_n4536) & (n_n4243) & (!x379x) & (x13477x)) + ((!n_n4533) & (n_n4536) & (n_n4243) & (x379x) & (!x13477x)) + ((!n_n4533) & (n_n4536) & (n_n4243) & (x379x) & (x13477x)) + ((n_n4533) & (!n_n4536) & (!n_n4243) & (!x379x) & (!x13477x)) + ((n_n4533) & (!n_n4536) & (!n_n4243) & (!x379x) & (x13477x)) + ((n_n4533) & (!n_n4536) & (!n_n4243) & (x379x) & (!x13477x)) + ((n_n4533) & (!n_n4536) & (!n_n4243) & (x379x) & (x13477x)) + ((n_n4533) & (!n_n4536) & (n_n4243) & (!x379x) & (!x13477x)) + ((n_n4533) & (!n_n4536) & (n_n4243) & (!x379x) & (x13477x)) + ((n_n4533) & (!n_n4536) & (n_n4243) & (x379x) & (!x13477x)) + ((n_n4533) & (!n_n4536) & (n_n4243) & (x379x) & (x13477x)) + ((n_n4533) & (n_n4536) & (!n_n4243) & (!x379x) & (!x13477x)) + ((n_n4533) & (n_n4536) & (!n_n4243) & (!x379x) & (x13477x)) + ((n_n4533) & (n_n4536) & (!n_n4243) & (x379x) & (!x13477x)) + ((n_n4533) & (n_n4536) & (!n_n4243) & (x379x) & (x13477x)) + ((n_n4533) & (n_n4536) & (n_n4243) & (!x379x) & (!x13477x)) + ((n_n4533) & (n_n4536) & (n_n4243) & (!x379x) & (x13477x)) + ((n_n4533) & (n_n4536) & (n_n4243) & (x379x) & (!x13477x)) + ((n_n4533) & (n_n4536) & (n_n4243) & (x379x) & (x13477x)));
	assign x13482x = (((!x455x) & (!x13471x) & (!n_n4086) & (!x222x) & (x13480x)) + ((!x455x) & (!x13471x) & (!n_n4086) & (x222x) & (!x13480x)) + ((!x455x) & (!x13471x) & (!n_n4086) & (x222x) & (x13480x)) + ((!x455x) & (!x13471x) & (n_n4086) & (!x222x) & (!x13480x)) + ((!x455x) & (!x13471x) & (n_n4086) & (!x222x) & (x13480x)) + ((!x455x) & (!x13471x) & (n_n4086) & (x222x) & (!x13480x)) + ((!x455x) & (!x13471x) & (n_n4086) & (x222x) & (x13480x)) + ((!x455x) & (x13471x) & (!n_n4086) & (!x222x) & (!x13480x)) + ((!x455x) & (x13471x) & (!n_n4086) & (!x222x) & (x13480x)) + ((!x455x) & (x13471x) & (!n_n4086) & (x222x) & (!x13480x)) + ((!x455x) & (x13471x) & (!n_n4086) & (x222x) & (x13480x)) + ((!x455x) & (x13471x) & (n_n4086) & (!x222x) & (!x13480x)) + ((!x455x) & (x13471x) & (n_n4086) & (!x222x) & (x13480x)) + ((!x455x) & (x13471x) & (n_n4086) & (x222x) & (!x13480x)) + ((!x455x) & (x13471x) & (n_n4086) & (x222x) & (x13480x)) + ((x455x) & (!x13471x) & (!n_n4086) & (!x222x) & (!x13480x)) + ((x455x) & (!x13471x) & (!n_n4086) & (!x222x) & (x13480x)) + ((x455x) & (!x13471x) & (!n_n4086) & (x222x) & (!x13480x)) + ((x455x) & (!x13471x) & (!n_n4086) & (x222x) & (x13480x)) + ((x455x) & (!x13471x) & (n_n4086) & (!x222x) & (!x13480x)) + ((x455x) & (!x13471x) & (n_n4086) & (!x222x) & (x13480x)) + ((x455x) & (!x13471x) & (n_n4086) & (x222x) & (!x13480x)) + ((x455x) & (!x13471x) & (n_n4086) & (x222x) & (x13480x)) + ((x455x) & (x13471x) & (!n_n4086) & (!x222x) & (!x13480x)) + ((x455x) & (x13471x) & (!n_n4086) & (!x222x) & (x13480x)) + ((x455x) & (x13471x) & (!n_n4086) & (x222x) & (!x13480x)) + ((x455x) & (x13471x) & (!n_n4086) & (x222x) & (x13480x)) + ((x455x) & (x13471x) & (n_n4086) & (!x222x) & (!x13480x)) + ((x455x) & (x13471x) & (n_n4086) & (!x222x) & (x13480x)) + ((x455x) & (x13471x) & (n_n4086) & (x222x) & (!x13480x)) + ((x455x) & (x13471x) & (n_n4086) & (x222x) & (x13480x)));
	assign n_n4016 = (((!n_n4083) & (!n_n4082) & (!x13450x) & (x13451x)) + ((!n_n4083) & (!n_n4082) & (x13450x) & (!x13451x)) + ((!n_n4083) & (!n_n4082) & (x13450x) & (x13451x)) + ((!n_n4083) & (n_n4082) & (!x13450x) & (!x13451x)) + ((!n_n4083) & (n_n4082) & (!x13450x) & (x13451x)) + ((!n_n4083) & (n_n4082) & (x13450x) & (!x13451x)) + ((!n_n4083) & (n_n4082) & (x13450x) & (x13451x)) + ((n_n4083) & (!n_n4082) & (!x13450x) & (!x13451x)) + ((n_n4083) & (!n_n4082) & (!x13450x) & (x13451x)) + ((n_n4083) & (!n_n4082) & (x13450x) & (!x13451x)) + ((n_n4083) & (!n_n4082) & (x13450x) & (x13451x)) + ((n_n4083) & (n_n4082) & (!x13450x) & (!x13451x)) + ((n_n4083) & (n_n4082) & (!x13450x) & (x13451x)) + ((n_n4083) & (n_n4082) & (x13450x) & (!x13451x)) + ((n_n4083) & (n_n4082) & (x13450x) & (x13451x)));
	assign n_n4015 = (((!n_n4232) & (!n_n1648) & (!n_n4079) & (!x13464x) & (x13466x)) + ((!n_n4232) & (!n_n1648) & (!n_n4079) & (x13464x) & (!x13466x)) + ((!n_n4232) & (!n_n1648) & (!n_n4079) & (x13464x) & (x13466x)) + ((!n_n4232) & (!n_n1648) & (n_n4079) & (!x13464x) & (!x13466x)) + ((!n_n4232) & (!n_n1648) & (n_n4079) & (!x13464x) & (x13466x)) + ((!n_n4232) & (!n_n1648) & (n_n4079) & (x13464x) & (!x13466x)) + ((!n_n4232) & (!n_n1648) & (n_n4079) & (x13464x) & (x13466x)) + ((!n_n4232) & (n_n1648) & (!n_n4079) & (!x13464x) & (!x13466x)) + ((!n_n4232) & (n_n1648) & (!n_n4079) & (!x13464x) & (x13466x)) + ((!n_n4232) & (n_n1648) & (!n_n4079) & (x13464x) & (!x13466x)) + ((!n_n4232) & (n_n1648) & (!n_n4079) & (x13464x) & (x13466x)) + ((!n_n4232) & (n_n1648) & (n_n4079) & (!x13464x) & (!x13466x)) + ((!n_n4232) & (n_n1648) & (n_n4079) & (!x13464x) & (x13466x)) + ((!n_n4232) & (n_n1648) & (n_n4079) & (x13464x) & (!x13466x)) + ((!n_n4232) & (n_n1648) & (n_n4079) & (x13464x) & (x13466x)) + ((n_n4232) & (!n_n1648) & (!n_n4079) & (!x13464x) & (!x13466x)) + ((n_n4232) & (!n_n1648) & (!n_n4079) & (!x13464x) & (x13466x)) + ((n_n4232) & (!n_n1648) & (!n_n4079) & (x13464x) & (!x13466x)) + ((n_n4232) & (!n_n1648) & (!n_n4079) & (x13464x) & (x13466x)) + ((n_n4232) & (!n_n1648) & (n_n4079) & (!x13464x) & (!x13466x)) + ((n_n4232) & (!n_n1648) & (n_n4079) & (!x13464x) & (x13466x)) + ((n_n4232) & (!n_n1648) & (n_n4079) & (x13464x) & (!x13466x)) + ((n_n4232) & (!n_n1648) & (n_n4079) & (x13464x) & (x13466x)) + ((n_n4232) & (n_n1648) & (!n_n4079) & (!x13464x) & (!x13466x)) + ((n_n4232) & (n_n1648) & (!n_n4079) & (!x13464x) & (x13466x)) + ((n_n4232) & (n_n1648) & (!n_n4079) & (x13464x) & (!x13466x)) + ((n_n4232) & (n_n1648) & (!n_n4079) & (x13464x) & (x13466x)) + ((n_n4232) & (n_n1648) & (n_n4079) & (!x13464x) & (!x13466x)) + ((n_n4232) & (n_n1648) & (n_n4079) & (!x13464x) & (x13466x)) + ((n_n4232) & (n_n1648) & (n_n4079) & (x13464x) & (!x13466x)) + ((n_n4232) & (n_n1648) & (n_n4079) & (x13464x) & (x13466x)));
	assign x13487x = (((!n_n524) & (!x13x) & (!n_n509) & (!n_n4489) & (x199x)) + ((!n_n524) & (!x13x) & (!n_n509) & (n_n4489) & (!x199x)) + ((!n_n524) & (!x13x) & (!n_n509) & (n_n4489) & (x199x)) + ((!n_n524) & (!x13x) & (n_n509) & (!n_n4489) & (x199x)) + ((!n_n524) & (!x13x) & (n_n509) & (n_n4489) & (!x199x)) + ((!n_n524) & (!x13x) & (n_n509) & (n_n4489) & (x199x)) + ((!n_n524) & (x13x) & (!n_n509) & (!n_n4489) & (x199x)) + ((!n_n524) & (x13x) & (!n_n509) & (n_n4489) & (!x199x)) + ((!n_n524) & (x13x) & (!n_n509) & (n_n4489) & (x199x)) + ((!n_n524) & (x13x) & (n_n509) & (!n_n4489) & (x199x)) + ((!n_n524) & (x13x) & (n_n509) & (n_n4489) & (!x199x)) + ((!n_n524) & (x13x) & (n_n509) & (n_n4489) & (x199x)) + ((n_n524) & (!x13x) & (!n_n509) & (!n_n4489) & (x199x)) + ((n_n524) & (!x13x) & (!n_n509) & (n_n4489) & (!x199x)) + ((n_n524) & (!x13x) & (!n_n509) & (n_n4489) & (x199x)) + ((n_n524) & (!x13x) & (n_n509) & (!n_n4489) & (x199x)) + ((n_n524) & (!x13x) & (n_n509) & (n_n4489) & (!x199x)) + ((n_n524) & (!x13x) & (n_n509) & (n_n4489) & (x199x)) + ((n_n524) & (x13x) & (!n_n509) & (!n_n4489) & (x199x)) + ((n_n524) & (x13x) & (!n_n509) & (n_n4489) & (!x199x)) + ((n_n524) & (x13x) & (!n_n509) & (n_n4489) & (x199x)) + ((n_n524) & (x13x) & (n_n509) & (!n_n4489) & (!x199x)) + ((n_n524) & (x13x) & (n_n509) & (!n_n4489) & (x199x)) + ((n_n524) & (x13x) & (n_n509) & (n_n4489) & (!x199x)) + ((n_n524) & (x13x) & (n_n509) & (n_n4489) & (x199x)));
	assign x13488x = (((!n_n4487) & (!n_n4478) & (!x70x) & (n_n4486)) + ((!n_n4487) & (!n_n4478) & (x70x) & (!n_n4486)) + ((!n_n4487) & (!n_n4478) & (x70x) & (n_n4486)) + ((!n_n4487) & (n_n4478) & (!x70x) & (!n_n4486)) + ((!n_n4487) & (n_n4478) & (!x70x) & (n_n4486)) + ((!n_n4487) & (n_n4478) & (x70x) & (!n_n4486)) + ((!n_n4487) & (n_n4478) & (x70x) & (n_n4486)) + ((n_n4487) & (!n_n4478) & (!x70x) & (!n_n4486)) + ((n_n4487) & (!n_n4478) & (!x70x) & (n_n4486)) + ((n_n4487) & (!n_n4478) & (x70x) & (!n_n4486)) + ((n_n4487) & (!n_n4478) & (x70x) & (n_n4486)) + ((n_n4487) & (n_n4478) & (!x70x) & (!n_n4486)) + ((n_n4487) & (n_n4478) & (!x70x) & (n_n4486)) + ((n_n4487) & (n_n4478) & (x70x) & (!n_n4486)) + ((n_n4487) & (n_n4478) & (x70x) & (n_n4486)));
	assign x13501x = (((!n_n4512) & (!n_n4247) & (!n_n4246) & (!n_n3152) & (n_n4503)) + ((!n_n4512) & (!n_n4247) & (!n_n4246) & (n_n3152) & (!n_n4503)) + ((!n_n4512) & (!n_n4247) & (!n_n4246) & (n_n3152) & (n_n4503)) + ((!n_n4512) & (!n_n4247) & (n_n4246) & (!n_n3152) & (!n_n4503)) + ((!n_n4512) & (!n_n4247) & (n_n4246) & (!n_n3152) & (n_n4503)) + ((!n_n4512) & (!n_n4247) & (n_n4246) & (n_n3152) & (!n_n4503)) + ((!n_n4512) & (!n_n4247) & (n_n4246) & (n_n3152) & (n_n4503)) + ((!n_n4512) & (n_n4247) & (!n_n4246) & (!n_n3152) & (!n_n4503)) + ((!n_n4512) & (n_n4247) & (!n_n4246) & (!n_n3152) & (n_n4503)) + ((!n_n4512) & (n_n4247) & (!n_n4246) & (n_n3152) & (!n_n4503)) + ((!n_n4512) & (n_n4247) & (!n_n4246) & (n_n3152) & (n_n4503)) + ((!n_n4512) & (n_n4247) & (n_n4246) & (!n_n3152) & (!n_n4503)) + ((!n_n4512) & (n_n4247) & (n_n4246) & (!n_n3152) & (n_n4503)) + ((!n_n4512) & (n_n4247) & (n_n4246) & (n_n3152) & (!n_n4503)) + ((!n_n4512) & (n_n4247) & (n_n4246) & (n_n3152) & (n_n4503)) + ((n_n4512) & (!n_n4247) & (!n_n4246) & (!n_n3152) & (!n_n4503)) + ((n_n4512) & (!n_n4247) & (!n_n4246) & (!n_n3152) & (n_n4503)) + ((n_n4512) & (!n_n4247) & (!n_n4246) & (n_n3152) & (!n_n4503)) + ((n_n4512) & (!n_n4247) & (!n_n4246) & (n_n3152) & (n_n4503)) + ((n_n4512) & (!n_n4247) & (n_n4246) & (!n_n3152) & (!n_n4503)) + ((n_n4512) & (!n_n4247) & (n_n4246) & (!n_n3152) & (n_n4503)) + ((n_n4512) & (!n_n4247) & (n_n4246) & (n_n3152) & (!n_n4503)) + ((n_n4512) & (!n_n4247) & (n_n4246) & (n_n3152) & (n_n4503)) + ((n_n4512) & (n_n4247) & (!n_n4246) & (!n_n3152) & (!n_n4503)) + ((n_n4512) & (n_n4247) & (!n_n4246) & (!n_n3152) & (n_n4503)) + ((n_n4512) & (n_n4247) & (!n_n4246) & (n_n3152) & (!n_n4503)) + ((n_n4512) & (n_n4247) & (!n_n4246) & (n_n3152) & (n_n4503)) + ((n_n4512) & (n_n4247) & (n_n4246) & (!n_n3152) & (!n_n4503)) + ((n_n4512) & (n_n4247) & (n_n4246) & (!n_n3152) & (n_n4503)) + ((n_n4512) & (n_n4247) & (n_n4246) & (n_n3152) & (!n_n4503)) + ((n_n4512) & (n_n4247) & (n_n4246) & (n_n3152) & (n_n4503)));
	assign x13503x = (((!i_9_) & (!n_n524) & (n_n518) & (n_n455) & (x23x)) + ((!i_9_) & (n_n524) & (n_n518) & (n_n455) & (!x23x)) + ((!i_9_) & (n_n524) & (n_n518) & (n_n455) & (x23x)) + ((i_9_) & (!n_n524) & (n_n518) & (n_n455) & (x23x)) + ((i_9_) & (n_n524) & (n_n518) & (n_n455) & (x23x)));
	assign n_n4092 = (((!x147x) & (!n_n4468) & (!n_n4254) & (!n_n4469) & (x13503x)) + ((!x147x) & (!n_n4468) & (!n_n4254) & (n_n4469) & (!x13503x)) + ((!x147x) & (!n_n4468) & (!n_n4254) & (n_n4469) & (x13503x)) + ((!x147x) & (!n_n4468) & (n_n4254) & (!n_n4469) & (!x13503x)) + ((!x147x) & (!n_n4468) & (n_n4254) & (!n_n4469) & (x13503x)) + ((!x147x) & (!n_n4468) & (n_n4254) & (n_n4469) & (!x13503x)) + ((!x147x) & (!n_n4468) & (n_n4254) & (n_n4469) & (x13503x)) + ((!x147x) & (n_n4468) & (!n_n4254) & (!n_n4469) & (!x13503x)) + ((!x147x) & (n_n4468) & (!n_n4254) & (!n_n4469) & (x13503x)) + ((!x147x) & (n_n4468) & (!n_n4254) & (n_n4469) & (!x13503x)) + ((!x147x) & (n_n4468) & (!n_n4254) & (n_n4469) & (x13503x)) + ((!x147x) & (n_n4468) & (n_n4254) & (!n_n4469) & (!x13503x)) + ((!x147x) & (n_n4468) & (n_n4254) & (!n_n4469) & (x13503x)) + ((!x147x) & (n_n4468) & (n_n4254) & (n_n4469) & (!x13503x)) + ((!x147x) & (n_n4468) & (n_n4254) & (n_n4469) & (x13503x)) + ((x147x) & (!n_n4468) & (!n_n4254) & (!n_n4469) & (!x13503x)) + ((x147x) & (!n_n4468) & (!n_n4254) & (!n_n4469) & (x13503x)) + ((x147x) & (!n_n4468) & (!n_n4254) & (n_n4469) & (!x13503x)) + ((x147x) & (!n_n4468) & (!n_n4254) & (n_n4469) & (x13503x)) + ((x147x) & (!n_n4468) & (n_n4254) & (!n_n4469) & (!x13503x)) + ((x147x) & (!n_n4468) & (n_n4254) & (!n_n4469) & (x13503x)) + ((x147x) & (!n_n4468) & (n_n4254) & (n_n4469) & (!x13503x)) + ((x147x) & (!n_n4468) & (n_n4254) & (n_n4469) & (x13503x)) + ((x147x) & (n_n4468) & (!n_n4254) & (!n_n4469) & (!x13503x)) + ((x147x) & (n_n4468) & (!n_n4254) & (!n_n4469) & (x13503x)) + ((x147x) & (n_n4468) & (!n_n4254) & (n_n4469) & (!x13503x)) + ((x147x) & (n_n4468) & (!n_n4254) & (n_n4469) & (x13503x)) + ((x147x) & (n_n4468) & (n_n4254) & (!n_n4469) & (!x13503x)) + ((x147x) & (n_n4468) & (n_n4254) & (!n_n4469) & (x13503x)) + ((x147x) & (n_n4468) & (n_n4254) & (n_n4469) & (!x13503x)) + ((x147x) & (n_n4468) & (n_n4254) & (n_n4469) & (x13503x)));
	assign n_n4023 = (((!x283x) & (!n_n4103) & (!x363x) & (!x443x) & (x13519x)) + ((!x283x) & (!n_n4103) & (!x363x) & (x443x) & (!x13519x)) + ((!x283x) & (!n_n4103) & (!x363x) & (x443x) & (x13519x)) + ((!x283x) & (!n_n4103) & (x363x) & (!x443x) & (!x13519x)) + ((!x283x) & (!n_n4103) & (x363x) & (!x443x) & (x13519x)) + ((!x283x) & (!n_n4103) & (x363x) & (x443x) & (!x13519x)) + ((!x283x) & (!n_n4103) & (x363x) & (x443x) & (x13519x)) + ((!x283x) & (n_n4103) & (!x363x) & (!x443x) & (!x13519x)) + ((!x283x) & (n_n4103) & (!x363x) & (!x443x) & (x13519x)) + ((!x283x) & (n_n4103) & (!x363x) & (x443x) & (!x13519x)) + ((!x283x) & (n_n4103) & (!x363x) & (x443x) & (x13519x)) + ((!x283x) & (n_n4103) & (x363x) & (!x443x) & (!x13519x)) + ((!x283x) & (n_n4103) & (x363x) & (!x443x) & (x13519x)) + ((!x283x) & (n_n4103) & (x363x) & (x443x) & (!x13519x)) + ((!x283x) & (n_n4103) & (x363x) & (x443x) & (x13519x)) + ((x283x) & (!n_n4103) & (!x363x) & (!x443x) & (!x13519x)) + ((x283x) & (!n_n4103) & (!x363x) & (!x443x) & (x13519x)) + ((x283x) & (!n_n4103) & (!x363x) & (x443x) & (!x13519x)) + ((x283x) & (!n_n4103) & (!x363x) & (x443x) & (x13519x)) + ((x283x) & (!n_n4103) & (x363x) & (!x443x) & (!x13519x)) + ((x283x) & (!n_n4103) & (x363x) & (!x443x) & (x13519x)) + ((x283x) & (!n_n4103) & (x363x) & (x443x) & (!x13519x)) + ((x283x) & (!n_n4103) & (x363x) & (x443x) & (x13519x)) + ((x283x) & (n_n4103) & (!x363x) & (!x443x) & (!x13519x)) + ((x283x) & (n_n4103) & (!x363x) & (!x443x) & (x13519x)) + ((x283x) & (n_n4103) & (!x363x) & (x443x) & (!x13519x)) + ((x283x) & (n_n4103) & (!x363x) & (x443x) & (x13519x)) + ((x283x) & (n_n4103) & (x363x) & (!x443x) & (!x13519x)) + ((x283x) & (n_n4103) & (x363x) & (!x443x) & (x13519x)) + ((x283x) & (n_n4103) & (x363x) & (x443x) & (!x13519x)) + ((x283x) & (n_n4103) & (x363x) & (x443x) & (x13519x)));
	assign n_n4100 = (((!n_n4372) & (!x423x) & (!n_n4375) & (!x301x) & (x27x)) + ((!n_n4372) & (!x423x) & (!n_n4375) & (x301x) & (!x27x)) + ((!n_n4372) & (!x423x) & (!n_n4375) & (x301x) & (x27x)) + ((!n_n4372) & (!x423x) & (n_n4375) & (!x301x) & (!x27x)) + ((!n_n4372) & (!x423x) & (n_n4375) & (!x301x) & (x27x)) + ((!n_n4372) & (!x423x) & (n_n4375) & (x301x) & (!x27x)) + ((!n_n4372) & (!x423x) & (n_n4375) & (x301x) & (x27x)) + ((!n_n4372) & (x423x) & (!n_n4375) & (!x301x) & (!x27x)) + ((!n_n4372) & (x423x) & (!n_n4375) & (!x301x) & (x27x)) + ((!n_n4372) & (x423x) & (!n_n4375) & (x301x) & (!x27x)) + ((!n_n4372) & (x423x) & (!n_n4375) & (x301x) & (x27x)) + ((!n_n4372) & (x423x) & (n_n4375) & (!x301x) & (!x27x)) + ((!n_n4372) & (x423x) & (n_n4375) & (!x301x) & (x27x)) + ((!n_n4372) & (x423x) & (n_n4375) & (x301x) & (!x27x)) + ((!n_n4372) & (x423x) & (n_n4375) & (x301x) & (x27x)) + ((n_n4372) & (!x423x) & (!n_n4375) & (!x301x) & (!x27x)) + ((n_n4372) & (!x423x) & (!n_n4375) & (!x301x) & (x27x)) + ((n_n4372) & (!x423x) & (!n_n4375) & (x301x) & (!x27x)) + ((n_n4372) & (!x423x) & (!n_n4375) & (x301x) & (x27x)) + ((n_n4372) & (!x423x) & (n_n4375) & (!x301x) & (!x27x)) + ((n_n4372) & (!x423x) & (n_n4375) & (!x301x) & (x27x)) + ((n_n4372) & (!x423x) & (n_n4375) & (x301x) & (!x27x)) + ((n_n4372) & (!x423x) & (n_n4375) & (x301x) & (x27x)) + ((n_n4372) & (x423x) & (!n_n4375) & (!x301x) & (!x27x)) + ((n_n4372) & (x423x) & (!n_n4375) & (!x301x) & (x27x)) + ((n_n4372) & (x423x) & (!n_n4375) & (x301x) & (!x27x)) + ((n_n4372) & (x423x) & (!n_n4375) & (x301x) & (x27x)) + ((n_n4372) & (x423x) & (n_n4375) & (!x301x) & (!x27x)) + ((n_n4372) & (x423x) & (n_n4375) & (!x301x) & (x27x)) + ((n_n4372) & (x423x) & (n_n4375) & (x301x) & (!x27x)) + ((n_n4372) & (x423x) & (n_n4375) & (x301x) & (x27x)));
	assign n_n4102 = (((!n_n4357) & (!n_n4353) & (!n_n1002) & (!x74x) & (x398x)) + ((!n_n4357) & (!n_n4353) & (!n_n1002) & (x74x) & (!x398x)) + ((!n_n4357) & (!n_n4353) & (!n_n1002) & (x74x) & (x398x)) + ((!n_n4357) & (!n_n4353) & (n_n1002) & (!x74x) & (!x398x)) + ((!n_n4357) & (!n_n4353) & (n_n1002) & (!x74x) & (x398x)) + ((!n_n4357) & (!n_n4353) & (n_n1002) & (x74x) & (!x398x)) + ((!n_n4357) & (!n_n4353) & (n_n1002) & (x74x) & (x398x)) + ((!n_n4357) & (n_n4353) & (!n_n1002) & (!x74x) & (!x398x)) + ((!n_n4357) & (n_n4353) & (!n_n1002) & (!x74x) & (x398x)) + ((!n_n4357) & (n_n4353) & (!n_n1002) & (x74x) & (!x398x)) + ((!n_n4357) & (n_n4353) & (!n_n1002) & (x74x) & (x398x)) + ((!n_n4357) & (n_n4353) & (n_n1002) & (!x74x) & (!x398x)) + ((!n_n4357) & (n_n4353) & (n_n1002) & (!x74x) & (x398x)) + ((!n_n4357) & (n_n4353) & (n_n1002) & (x74x) & (!x398x)) + ((!n_n4357) & (n_n4353) & (n_n1002) & (x74x) & (x398x)) + ((n_n4357) & (!n_n4353) & (!n_n1002) & (!x74x) & (!x398x)) + ((n_n4357) & (!n_n4353) & (!n_n1002) & (!x74x) & (x398x)) + ((n_n4357) & (!n_n4353) & (!n_n1002) & (x74x) & (!x398x)) + ((n_n4357) & (!n_n4353) & (!n_n1002) & (x74x) & (x398x)) + ((n_n4357) & (!n_n4353) & (n_n1002) & (!x74x) & (!x398x)) + ((n_n4357) & (!n_n4353) & (n_n1002) & (!x74x) & (x398x)) + ((n_n4357) & (!n_n4353) & (n_n1002) & (x74x) & (!x398x)) + ((n_n4357) & (!n_n4353) & (n_n1002) & (x74x) & (x398x)) + ((n_n4357) & (n_n4353) & (!n_n1002) & (!x74x) & (!x398x)) + ((n_n4357) & (n_n4353) & (!n_n1002) & (!x74x) & (x398x)) + ((n_n4357) & (n_n4353) & (!n_n1002) & (x74x) & (!x398x)) + ((n_n4357) & (n_n4353) & (!n_n1002) & (x74x) & (x398x)) + ((n_n4357) & (n_n4353) & (n_n1002) & (!x74x) & (!x398x)) + ((n_n4357) & (n_n4353) & (n_n1002) & (!x74x) & (x398x)) + ((n_n4357) & (n_n4353) & (n_n1002) & (x74x) & (!x398x)) + ((n_n4357) & (n_n4353) & (n_n1002) & (x74x) & (x398x)));
	assign n_n4021 = (((!x425x) & (!x420x) & (!n_n4097) & (!x13533x) & (x13539x)) + ((!x425x) & (!x420x) & (!n_n4097) & (x13533x) & (!x13539x)) + ((!x425x) & (!x420x) & (!n_n4097) & (x13533x) & (x13539x)) + ((!x425x) & (!x420x) & (n_n4097) & (!x13533x) & (!x13539x)) + ((!x425x) & (!x420x) & (n_n4097) & (!x13533x) & (x13539x)) + ((!x425x) & (!x420x) & (n_n4097) & (x13533x) & (!x13539x)) + ((!x425x) & (!x420x) & (n_n4097) & (x13533x) & (x13539x)) + ((!x425x) & (x420x) & (!n_n4097) & (!x13533x) & (!x13539x)) + ((!x425x) & (x420x) & (!n_n4097) & (!x13533x) & (x13539x)) + ((!x425x) & (x420x) & (!n_n4097) & (x13533x) & (!x13539x)) + ((!x425x) & (x420x) & (!n_n4097) & (x13533x) & (x13539x)) + ((!x425x) & (x420x) & (n_n4097) & (!x13533x) & (!x13539x)) + ((!x425x) & (x420x) & (n_n4097) & (!x13533x) & (x13539x)) + ((!x425x) & (x420x) & (n_n4097) & (x13533x) & (!x13539x)) + ((!x425x) & (x420x) & (n_n4097) & (x13533x) & (x13539x)) + ((x425x) & (!x420x) & (!n_n4097) & (!x13533x) & (!x13539x)) + ((x425x) & (!x420x) & (!n_n4097) & (!x13533x) & (x13539x)) + ((x425x) & (!x420x) & (!n_n4097) & (x13533x) & (!x13539x)) + ((x425x) & (!x420x) & (!n_n4097) & (x13533x) & (x13539x)) + ((x425x) & (!x420x) & (n_n4097) & (!x13533x) & (!x13539x)) + ((x425x) & (!x420x) & (n_n4097) & (!x13533x) & (x13539x)) + ((x425x) & (!x420x) & (n_n4097) & (x13533x) & (!x13539x)) + ((x425x) & (!x420x) & (n_n4097) & (x13533x) & (x13539x)) + ((x425x) & (x420x) & (!n_n4097) & (!x13533x) & (!x13539x)) + ((x425x) & (x420x) & (!n_n4097) & (!x13533x) & (x13539x)) + ((x425x) & (x420x) & (!n_n4097) & (x13533x) & (!x13539x)) + ((x425x) & (x420x) & (!n_n4097) & (x13533x) & (x13539x)) + ((x425x) & (x420x) & (n_n4097) & (!x13533x) & (!x13539x)) + ((x425x) & (x420x) & (n_n4097) & (!x13533x) & (x13539x)) + ((x425x) & (x420x) & (n_n4097) & (x13533x) & (!x13539x)) + ((x425x) & (x420x) & (n_n4097) & (x13533x) & (x13539x)));
	assign x13545x = (((!n_n4369) & (!n_n4361) & (!n_n4359) & (!n_n4367) & (x13544x)) + ((!n_n4369) & (!n_n4361) & (!n_n4359) & (n_n4367) & (!x13544x)) + ((!n_n4369) & (!n_n4361) & (!n_n4359) & (n_n4367) & (x13544x)) + ((!n_n4369) & (!n_n4361) & (n_n4359) & (!n_n4367) & (!x13544x)) + ((!n_n4369) & (!n_n4361) & (n_n4359) & (!n_n4367) & (x13544x)) + ((!n_n4369) & (!n_n4361) & (n_n4359) & (n_n4367) & (!x13544x)) + ((!n_n4369) & (!n_n4361) & (n_n4359) & (n_n4367) & (x13544x)) + ((!n_n4369) & (n_n4361) & (!n_n4359) & (!n_n4367) & (!x13544x)) + ((!n_n4369) & (n_n4361) & (!n_n4359) & (!n_n4367) & (x13544x)) + ((!n_n4369) & (n_n4361) & (!n_n4359) & (n_n4367) & (!x13544x)) + ((!n_n4369) & (n_n4361) & (!n_n4359) & (n_n4367) & (x13544x)) + ((!n_n4369) & (n_n4361) & (n_n4359) & (!n_n4367) & (!x13544x)) + ((!n_n4369) & (n_n4361) & (n_n4359) & (!n_n4367) & (x13544x)) + ((!n_n4369) & (n_n4361) & (n_n4359) & (n_n4367) & (!x13544x)) + ((!n_n4369) & (n_n4361) & (n_n4359) & (n_n4367) & (x13544x)) + ((n_n4369) & (!n_n4361) & (!n_n4359) & (!n_n4367) & (!x13544x)) + ((n_n4369) & (!n_n4361) & (!n_n4359) & (!n_n4367) & (x13544x)) + ((n_n4369) & (!n_n4361) & (!n_n4359) & (n_n4367) & (!x13544x)) + ((n_n4369) & (!n_n4361) & (!n_n4359) & (n_n4367) & (x13544x)) + ((n_n4369) & (!n_n4361) & (n_n4359) & (!n_n4367) & (!x13544x)) + ((n_n4369) & (!n_n4361) & (n_n4359) & (!n_n4367) & (x13544x)) + ((n_n4369) & (!n_n4361) & (n_n4359) & (n_n4367) & (!x13544x)) + ((n_n4369) & (!n_n4361) & (n_n4359) & (n_n4367) & (x13544x)) + ((n_n4369) & (n_n4361) & (!n_n4359) & (!n_n4367) & (!x13544x)) + ((n_n4369) & (n_n4361) & (!n_n4359) & (!n_n4367) & (x13544x)) + ((n_n4369) & (n_n4361) & (!n_n4359) & (n_n4367) & (!x13544x)) + ((n_n4369) & (n_n4361) & (!n_n4359) & (n_n4367) & (x13544x)) + ((n_n4369) & (n_n4361) & (n_n4359) & (!n_n4367) & (!x13544x)) + ((n_n4369) & (n_n4361) & (n_n4359) & (!n_n4367) & (x13544x)) + ((n_n4369) & (n_n4361) & (n_n4359) & (n_n4367) & (!x13544x)) + ((n_n4369) & (n_n4361) & (n_n4359) & (n_n4367) & (x13544x)));
	assign x55x = (((!i_9_) & (n_n518) & (n_n455) & (!n_n528) & (n_n530)) + ((!i_9_) & (n_n518) & (n_n455) & (n_n528) & (n_n530)) + ((i_9_) & (n_n518) & (n_n455) & (!n_n528) & (n_n530)) + ((i_9_) & (n_n518) & (n_n455) & (n_n528) & (!n_n530)) + ((i_9_) & (n_n518) & (n_n455) & (n_n528) & (n_n530)));
	assign n_n4090 = (((!n_n4494) & (!n_n4495) & (!x163x) & (!n_n4493) & (!x22122x)) + ((!n_n4494) & (!n_n4495) & (!x163x) & (n_n4493) & (!x22122x)) + ((!n_n4494) & (!n_n4495) & (!x163x) & (n_n4493) & (x22122x)) + ((!n_n4494) & (!n_n4495) & (x163x) & (!n_n4493) & (!x22122x)) + ((!n_n4494) & (!n_n4495) & (x163x) & (!n_n4493) & (x22122x)) + ((!n_n4494) & (!n_n4495) & (x163x) & (n_n4493) & (!x22122x)) + ((!n_n4494) & (!n_n4495) & (x163x) & (n_n4493) & (x22122x)) + ((!n_n4494) & (n_n4495) & (!x163x) & (!n_n4493) & (!x22122x)) + ((!n_n4494) & (n_n4495) & (!x163x) & (!n_n4493) & (x22122x)) + ((!n_n4494) & (n_n4495) & (!x163x) & (n_n4493) & (!x22122x)) + ((!n_n4494) & (n_n4495) & (!x163x) & (n_n4493) & (x22122x)) + ((!n_n4494) & (n_n4495) & (x163x) & (!n_n4493) & (!x22122x)) + ((!n_n4494) & (n_n4495) & (x163x) & (!n_n4493) & (x22122x)) + ((!n_n4494) & (n_n4495) & (x163x) & (n_n4493) & (!x22122x)) + ((!n_n4494) & (n_n4495) & (x163x) & (n_n4493) & (x22122x)) + ((n_n4494) & (!n_n4495) & (!x163x) & (!n_n4493) & (!x22122x)) + ((n_n4494) & (!n_n4495) & (!x163x) & (!n_n4493) & (x22122x)) + ((n_n4494) & (!n_n4495) & (!x163x) & (n_n4493) & (!x22122x)) + ((n_n4494) & (!n_n4495) & (!x163x) & (n_n4493) & (x22122x)) + ((n_n4494) & (!n_n4495) & (x163x) & (!n_n4493) & (!x22122x)) + ((n_n4494) & (!n_n4495) & (x163x) & (!n_n4493) & (x22122x)) + ((n_n4494) & (!n_n4495) & (x163x) & (n_n4493) & (!x22122x)) + ((n_n4494) & (!n_n4495) & (x163x) & (n_n4493) & (x22122x)) + ((n_n4494) & (n_n4495) & (!x163x) & (!n_n4493) & (!x22122x)) + ((n_n4494) & (n_n4495) & (!x163x) & (!n_n4493) & (x22122x)) + ((n_n4494) & (n_n4495) & (!x163x) & (n_n4493) & (!x22122x)) + ((n_n4494) & (n_n4495) & (!x163x) & (n_n4493) & (x22122x)) + ((n_n4494) & (n_n4495) & (x163x) & (!n_n4493) & (!x22122x)) + ((n_n4494) & (n_n4495) & (x163x) & (!n_n4493) & (x22122x)) + ((n_n4494) & (n_n4495) & (x163x) & (n_n4493) & (!x22122x)) + ((n_n4494) & (n_n4495) & (x163x) & (n_n4493) & (x22122x)));
	assign x13500x = (((!x13x) & (!x572x) & (!x189x) & (!x308x) & (x162x)) + ((!x13x) & (!x572x) & (!x189x) & (x308x) & (!x162x)) + ((!x13x) & (!x572x) & (!x189x) & (x308x) & (x162x)) + ((!x13x) & (!x572x) & (x189x) & (!x308x) & (!x162x)) + ((!x13x) & (!x572x) & (x189x) & (!x308x) & (x162x)) + ((!x13x) & (!x572x) & (x189x) & (x308x) & (!x162x)) + ((!x13x) & (!x572x) & (x189x) & (x308x) & (x162x)) + ((!x13x) & (x572x) & (!x189x) & (!x308x) & (x162x)) + ((!x13x) & (x572x) & (!x189x) & (x308x) & (!x162x)) + ((!x13x) & (x572x) & (!x189x) & (x308x) & (x162x)) + ((!x13x) & (x572x) & (x189x) & (!x308x) & (!x162x)) + ((!x13x) & (x572x) & (x189x) & (!x308x) & (x162x)) + ((!x13x) & (x572x) & (x189x) & (x308x) & (!x162x)) + ((!x13x) & (x572x) & (x189x) & (x308x) & (x162x)) + ((x13x) & (!x572x) & (!x189x) & (!x308x) & (x162x)) + ((x13x) & (!x572x) & (!x189x) & (x308x) & (!x162x)) + ((x13x) & (!x572x) & (!x189x) & (x308x) & (x162x)) + ((x13x) & (!x572x) & (x189x) & (!x308x) & (!x162x)) + ((x13x) & (!x572x) & (x189x) & (!x308x) & (x162x)) + ((x13x) & (!x572x) & (x189x) & (x308x) & (!x162x)) + ((x13x) & (!x572x) & (x189x) & (x308x) & (x162x)) + ((x13x) & (x572x) & (!x189x) & (!x308x) & (!x162x)) + ((x13x) & (x572x) & (!x189x) & (!x308x) & (x162x)) + ((x13x) & (x572x) & (!x189x) & (x308x) & (!x162x)) + ((x13x) & (x572x) & (!x189x) & (x308x) & (x162x)) + ((x13x) & (x572x) & (x189x) & (!x308x) & (!x162x)) + ((x13x) & (x572x) & (x189x) & (!x308x) & (x162x)) + ((x13x) & (x572x) & (x189x) & (x308x) & (!x162x)) + ((x13x) & (x572x) & (x189x) & (x308x) & (x162x)));
	assign x13553x = (((!x13487x) & (!x13488x) & (!n_n4092) & (x13551x)) + ((!x13487x) & (!x13488x) & (n_n4092) & (!x13551x)) + ((!x13487x) & (!x13488x) & (n_n4092) & (x13551x)) + ((!x13487x) & (x13488x) & (!n_n4092) & (!x13551x)) + ((!x13487x) & (x13488x) & (!n_n4092) & (x13551x)) + ((!x13487x) & (x13488x) & (n_n4092) & (!x13551x)) + ((!x13487x) & (x13488x) & (n_n4092) & (x13551x)) + ((x13487x) & (!x13488x) & (!n_n4092) & (!x13551x)) + ((x13487x) & (!x13488x) & (!n_n4092) & (x13551x)) + ((x13487x) & (!x13488x) & (n_n4092) & (!x13551x)) + ((x13487x) & (!x13488x) & (n_n4092) & (x13551x)) + ((x13487x) & (x13488x) & (!n_n4092) & (!x13551x)) + ((x13487x) & (x13488x) & (!n_n4092) & (x13551x)) + ((x13487x) & (x13488x) & (n_n4092) & (!x13551x)) + ((x13487x) & (x13488x) & (n_n4092) & (x13551x)));
	assign n_n4701 = (((!i_9_) & (n_n325) & (n_n535) & (n_n530)));
	assign x14393x = (((!n_n4615) & (!n_n4618) & (!n_n4629) & (n_n4630)) + ((!n_n4615) & (!n_n4618) & (n_n4629) & (!n_n4630)) + ((!n_n4615) & (!n_n4618) & (n_n4629) & (n_n4630)) + ((!n_n4615) & (n_n4618) & (!n_n4629) & (!n_n4630)) + ((!n_n4615) & (n_n4618) & (!n_n4629) & (n_n4630)) + ((!n_n4615) & (n_n4618) & (n_n4629) & (!n_n4630)) + ((!n_n4615) & (n_n4618) & (n_n4629) & (n_n4630)) + ((n_n4615) & (!n_n4618) & (!n_n4629) & (!n_n4630)) + ((n_n4615) & (!n_n4618) & (!n_n4629) & (n_n4630)) + ((n_n4615) & (!n_n4618) & (n_n4629) & (!n_n4630)) + ((n_n4615) & (!n_n4618) & (n_n4629) & (n_n4630)) + ((n_n4615) & (n_n4618) & (!n_n4629) & (!n_n4630)) + ((n_n4615) & (n_n4618) & (!n_n4629) & (n_n4630)) + ((n_n4615) & (n_n4618) & (n_n4629) & (!n_n4630)) + ((n_n4615) & (n_n4618) & (n_n4629) & (n_n4630)));
	assign x14394x = (((!n_n4625) & (!n_n4621) & (!n_n4622) & (!x75x) & (n_n4620)) + ((!n_n4625) & (!n_n4621) & (!n_n4622) & (x75x) & (!n_n4620)) + ((!n_n4625) & (!n_n4621) & (!n_n4622) & (x75x) & (n_n4620)) + ((!n_n4625) & (!n_n4621) & (n_n4622) & (!x75x) & (!n_n4620)) + ((!n_n4625) & (!n_n4621) & (n_n4622) & (!x75x) & (n_n4620)) + ((!n_n4625) & (!n_n4621) & (n_n4622) & (x75x) & (!n_n4620)) + ((!n_n4625) & (!n_n4621) & (n_n4622) & (x75x) & (n_n4620)) + ((!n_n4625) & (n_n4621) & (!n_n4622) & (!x75x) & (!n_n4620)) + ((!n_n4625) & (n_n4621) & (!n_n4622) & (!x75x) & (n_n4620)) + ((!n_n4625) & (n_n4621) & (!n_n4622) & (x75x) & (!n_n4620)) + ((!n_n4625) & (n_n4621) & (!n_n4622) & (x75x) & (n_n4620)) + ((!n_n4625) & (n_n4621) & (n_n4622) & (!x75x) & (!n_n4620)) + ((!n_n4625) & (n_n4621) & (n_n4622) & (!x75x) & (n_n4620)) + ((!n_n4625) & (n_n4621) & (n_n4622) & (x75x) & (!n_n4620)) + ((!n_n4625) & (n_n4621) & (n_n4622) & (x75x) & (n_n4620)) + ((n_n4625) & (!n_n4621) & (!n_n4622) & (!x75x) & (!n_n4620)) + ((n_n4625) & (!n_n4621) & (!n_n4622) & (!x75x) & (n_n4620)) + ((n_n4625) & (!n_n4621) & (!n_n4622) & (x75x) & (!n_n4620)) + ((n_n4625) & (!n_n4621) & (!n_n4622) & (x75x) & (n_n4620)) + ((n_n4625) & (!n_n4621) & (n_n4622) & (!x75x) & (!n_n4620)) + ((n_n4625) & (!n_n4621) & (n_n4622) & (!x75x) & (n_n4620)) + ((n_n4625) & (!n_n4621) & (n_n4622) & (x75x) & (!n_n4620)) + ((n_n4625) & (!n_n4621) & (n_n4622) & (x75x) & (n_n4620)) + ((n_n4625) & (n_n4621) & (!n_n4622) & (!x75x) & (!n_n4620)) + ((n_n4625) & (n_n4621) & (!n_n4622) & (!x75x) & (n_n4620)) + ((n_n4625) & (n_n4621) & (!n_n4622) & (x75x) & (!n_n4620)) + ((n_n4625) & (n_n4621) & (!n_n4622) & (x75x) & (n_n4620)) + ((n_n4625) & (n_n4621) & (n_n4622) & (!x75x) & (!n_n4620)) + ((n_n4625) & (n_n4621) & (n_n4622) & (!x75x) & (n_n4620)) + ((n_n4625) & (n_n4621) & (n_n4622) & (x75x) & (!n_n4620)) + ((n_n4625) & (n_n4621) & (n_n4622) & (x75x) & (n_n4620)));
	assign x431x = (((!i_9_) & (n_n482) & (n_n528) & (n_n390)) + ((i_9_) & (n_n482) & (n_n528) & (n_n390)));
	assign n_n2761 = (((!n_n390) & (!n_n491) & (!x20x) & (!x23x) & (n_n4648)) + ((!n_n390) & (!n_n491) & (!x20x) & (x23x) & (n_n4648)) + ((!n_n390) & (!n_n491) & (x20x) & (!x23x) & (n_n4648)) + ((!n_n390) & (!n_n491) & (x20x) & (x23x) & (n_n4648)) + ((!n_n390) & (n_n491) & (!x20x) & (!x23x) & (n_n4648)) + ((!n_n390) & (n_n491) & (!x20x) & (x23x) & (n_n4648)) + ((!n_n390) & (n_n491) & (x20x) & (!x23x) & (n_n4648)) + ((!n_n390) & (n_n491) & (x20x) & (x23x) & (n_n4648)) + ((n_n390) & (!n_n491) & (!x20x) & (!x23x) & (n_n4648)) + ((n_n390) & (!n_n491) & (!x20x) & (x23x) & (n_n4648)) + ((n_n390) & (!n_n491) & (x20x) & (!x23x) & (n_n4648)) + ((n_n390) & (!n_n491) & (x20x) & (x23x) & (n_n4648)) + ((n_n390) & (n_n491) & (!x20x) & (!x23x) & (n_n4648)) + ((n_n390) & (n_n491) & (!x20x) & (x23x) & (!n_n4648)) + ((n_n390) & (n_n491) & (!x20x) & (x23x) & (n_n4648)) + ((n_n390) & (n_n491) & (x20x) & (!x23x) & (!n_n4648)) + ((n_n390) & (n_n491) & (x20x) & (!x23x) & (n_n4648)) + ((n_n390) & (n_n491) & (x20x) & (x23x) & (!n_n4648)) + ((n_n390) & (n_n491) & (x20x) & (x23x) & (n_n4648)));
	assign n_n3714 = (((!n_n4652) & (!n_n4656) & (!x140x) & (!x431x) & (n_n2761)) + ((!n_n4652) & (!n_n4656) & (!x140x) & (x431x) & (!n_n2761)) + ((!n_n4652) & (!n_n4656) & (!x140x) & (x431x) & (n_n2761)) + ((!n_n4652) & (!n_n4656) & (x140x) & (!x431x) & (!n_n2761)) + ((!n_n4652) & (!n_n4656) & (x140x) & (!x431x) & (n_n2761)) + ((!n_n4652) & (!n_n4656) & (x140x) & (x431x) & (!n_n2761)) + ((!n_n4652) & (!n_n4656) & (x140x) & (x431x) & (n_n2761)) + ((!n_n4652) & (n_n4656) & (!x140x) & (!x431x) & (!n_n2761)) + ((!n_n4652) & (n_n4656) & (!x140x) & (!x431x) & (n_n2761)) + ((!n_n4652) & (n_n4656) & (!x140x) & (x431x) & (!n_n2761)) + ((!n_n4652) & (n_n4656) & (!x140x) & (x431x) & (n_n2761)) + ((!n_n4652) & (n_n4656) & (x140x) & (!x431x) & (!n_n2761)) + ((!n_n4652) & (n_n4656) & (x140x) & (!x431x) & (n_n2761)) + ((!n_n4652) & (n_n4656) & (x140x) & (x431x) & (!n_n2761)) + ((!n_n4652) & (n_n4656) & (x140x) & (x431x) & (n_n2761)) + ((n_n4652) & (!n_n4656) & (!x140x) & (!x431x) & (!n_n2761)) + ((n_n4652) & (!n_n4656) & (!x140x) & (!x431x) & (n_n2761)) + ((n_n4652) & (!n_n4656) & (!x140x) & (x431x) & (!n_n2761)) + ((n_n4652) & (!n_n4656) & (!x140x) & (x431x) & (n_n2761)) + ((n_n4652) & (!n_n4656) & (x140x) & (!x431x) & (!n_n2761)) + ((n_n4652) & (!n_n4656) & (x140x) & (!x431x) & (n_n2761)) + ((n_n4652) & (!n_n4656) & (x140x) & (x431x) & (!n_n2761)) + ((n_n4652) & (!n_n4656) & (x140x) & (x431x) & (n_n2761)) + ((n_n4652) & (n_n4656) & (!x140x) & (!x431x) & (!n_n2761)) + ((n_n4652) & (n_n4656) & (!x140x) & (!x431x) & (n_n2761)) + ((n_n4652) & (n_n4656) & (!x140x) & (x431x) & (!n_n2761)) + ((n_n4652) & (n_n4656) & (!x140x) & (x431x) & (n_n2761)) + ((n_n4652) & (n_n4656) & (x140x) & (!x431x) & (!n_n2761)) + ((n_n4652) & (n_n4656) & (x140x) & (!x431x) & (n_n2761)) + ((n_n4652) & (n_n4656) & (x140x) & (x431x) & (!n_n2761)) + ((n_n4652) & (n_n4656) & (x140x) & (x431x) & (n_n2761)));
	assign x119x = (((!i_9_) & (!n_n390) & (!n_n532) & (!n_n491) & (n_n4631)) + ((!i_9_) & (!n_n390) & (!n_n532) & (n_n491) & (n_n4631)) + ((!i_9_) & (!n_n390) & (n_n532) & (!n_n491) & (n_n4631)) + ((!i_9_) & (!n_n390) & (n_n532) & (n_n491) & (n_n4631)) + ((!i_9_) & (n_n390) & (!n_n532) & (!n_n491) & (n_n4631)) + ((!i_9_) & (n_n390) & (!n_n532) & (n_n491) & (n_n4631)) + ((!i_9_) & (n_n390) & (n_n532) & (!n_n491) & (n_n4631)) + ((!i_9_) & (n_n390) & (n_n532) & (n_n491) & (n_n4631)) + ((i_9_) & (!n_n390) & (!n_n532) & (!n_n491) & (n_n4631)) + ((i_9_) & (!n_n390) & (!n_n532) & (n_n491) & (n_n4631)) + ((i_9_) & (!n_n390) & (n_n532) & (!n_n491) & (n_n4631)) + ((i_9_) & (!n_n390) & (n_n532) & (n_n491) & (n_n4631)) + ((i_9_) & (n_n390) & (!n_n532) & (!n_n491) & (n_n4631)) + ((i_9_) & (n_n390) & (!n_n532) & (n_n491) & (n_n4631)) + ((i_9_) & (n_n390) & (n_n532) & (!n_n491) & (n_n4631)) + ((i_9_) & (n_n390) & (n_n532) & (n_n491) & (!n_n4631)) + ((i_9_) & (n_n390) & (n_n532) & (n_n491) & (n_n4631)));
	assign x14403x = (((!x492x) & (!x10x) & (!n_n4641) & (!n_n4639) & (n_n4640)) + ((!x492x) & (!x10x) & (!n_n4641) & (n_n4639) & (!n_n4640)) + ((!x492x) & (!x10x) & (!n_n4641) & (n_n4639) & (n_n4640)) + ((!x492x) & (!x10x) & (n_n4641) & (!n_n4639) & (!n_n4640)) + ((!x492x) & (!x10x) & (n_n4641) & (!n_n4639) & (n_n4640)) + ((!x492x) & (!x10x) & (n_n4641) & (n_n4639) & (!n_n4640)) + ((!x492x) & (!x10x) & (n_n4641) & (n_n4639) & (n_n4640)) + ((!x492x) & (x10x) & (!n_n4641) & (!n_n4639) & (n_n4640)) + ((!x492x) & (x10x) & (!n_n4641) & (n_n4639) & (!n_n4640)) + ((!x492x) & (x10x) & (!n_n4641) & (n_n4639) & (n_n4640)) + ((!x492x) & (x10x) & (n_n4641) & (!n_n4639) & (!n_n4640)) + ((!x492x) & (x10x) & (n_n4641) & (!n_n4639) & (n_n4640)) + ((!x492x) & (x10x) & (n_n4641) & (n_n4639) & (!n_n4640)) + ((!x492x) & (x10x) & (n_n4641) & (n_n4639) & (n_n4640)) + ((x492x) & (!x10x) & (!n_n4641) & (!n_n4639) & (n_n4640)) + ((x492x) & (!x10x) & (!n_n4641) & (n_n4639) & (!n_n4640)) + ((x492x) & (!x10x) & (!n_n4641) & (n_n4639) & (n_n4640)) + ((x492x) & (!x10x) & (n_n4641) & (!n_n4639) & (!n_n4640)) + ((x492x) & (!x10x) & (n_n4641) & (!n_n4639) & (n_n4640)) + ((x492x) & (!x10x) & (n_n4641) & (n_n4639) & (!n_n4640)) + ((x492x) & (!x10x) & (n_n4641) & (n_n4639) & (n_n4640)) + ((x492x) & (x10x) & (!n_n4641) & (!n_n4639) & (!n_n4640)) + ((x492x) & (x10x) & (!n_n4641) & (!n_n4639) & (n_n4640)) + ((x492x) & (x10x) & (!n_n4641) & (n_n4639) & (!n_n4640)) + ((x492x) & (x10x) & (!n_n4641) & (n_n4639) & (n_n4640)) + ((x492x) & (x10x) & (n_n4641) & (!n_n4639) & (!n_n4640)) + ((x492x) & (x10x) & (n_n4641) & (!n_n4639) & (n_n4640)) + ((x492x) & (x10x) & (n_n4641) & (n_n4639) & (!n_n4640)) + ((x492x) & (x10x) & (n_n4641) & (n_n4639) & (n_n4640)));
	assign x14404x = (((!n_n4634) & (!n_n4643) & (!n_n4642) & (!n_n4631) & (n_n4635)) + ((!n_n4634) & (!n_n4643) & (!n_n4642) & (n_n4631) & (!n_n4635)) + ((!n_n4634) & (!n_n4643) & (!n_n4642) & (n_n4631) & (n_n4635)) + ((!n_n4634) & (!n_n4643) & (n_n4642) & (!n_n4631) & (!n_n4635)) + ((!n_n4634) & (!n_n4643) & (n_n4642) & (!n_n4631) & (n_n4635)) + ((!n_n4634) & (!n_n4643) & (n_n4642) & (n_n4631) & (!n_n4635)) + ((!n_n4634) & (!n_n4643) & (n_n4642) & (n_n4631) & (n_n4635)) + ((!n_n4634) & (n_n4643) & (!n_n4642) & (!n_n4631) & (!n_n4635)) + ((!n_n4634) & (n_n4643) & (!n_n4642) & (!n_n4631) & (n_n4635)) + ((!n_n4634) & (n_n4643) & (!n_n4642) & (n_n4631) & (!n_n4635)) + ((!n_n4634) & (n_n4643) & (!n_n4642) & (n_n4631) & (n_n4635)) + ((!n_n4634) & (n_n4643) & (n_n4642) & (!n_n4631) & (!n_n4635)) + ((!n_n4634) & (n_n4643) & (n_n4642) & (!n_n4631) & (n_n4635)) + ((!n_n4634) & (n_n4643) & (n_n4642) & (n_n4631) & (!n_n4635)) + ((!n_n4634) & (n_n4643) & (n_n4642) & (n_n4631) & (n_n4635)) + ((n_n4634) & (!n_n4643) & (!n_n4642) & (!n_n4631) & (!n_n4635)) + ((n_n4634) & (!n_n4643) & (!n_n4642) & (!n_n4631) & (n_n4635)) + ((n_n4634) & (!n_n4643) & (!n_n4642) & (n_n4631) & (!n_n4635)) + ((n_n4634) & (!n_n4643) & (!n_n4642) & (n_n4631) & (n_n4635)) + ((n_n4634) & (!n_n4643) & (n_n4642) & (!n_n4631) & (!n_n4635)) + ((n_n4634) & (!n_n4643) & (n_n4642) & (!n_n4631) & (n_n4635)) + ((n_n4634) & (!n_n4643) & (n_n4642) & (n_n4631) & (!n_n4635)) + ((n_n4634) & (!n_n4643) & (n_n4642) & (n_n4631) & (n_n4635)) + ((n_n4634) & (n_n4643) & (!n_n4642) & (!n_n4631) & (!n_n4635)) + ((n_n4634) & (n_n4643) & (!n_n4642) & (!n_n4631) & (n_n4635)) + ((n_n4634) & (n_n4643) & (!n_n4642) & (n_n4631) & (!n_n4635)) + ((n_n4634) & (n_n4643) & (!n_n4642) & (n_n4631) & (n_n4635)) + ((n_n4634) & (n_n4643) & (n_n4642) & (!n_n4631) & (!n_n4635)) + ((n_n4634) & (n_n4643) & (n_n4642) & (!n_n4631) & (n_n4635)) + ((n_n4634) & (n_n4643) & (n_n4642) & (n_n4631) & (!n_n4635)) + ((n_n4634) & (n_n4643) & (n_n4642) & (n_n4631) & (n_n4635)));
	assign n_n3650 = (((!x14393x) & (!x14394x) & (!n_n3714) & (!x14403x) & (x14404x)) + ((!x14393x) & (!x14394x) & (!n_n3714) & (x14403x) & (!x14404x)) + ((!x14393x) & (!x14394x) & (!n_n3714) & (x14403x) & (x14404x)) + ((!x14393x) & (!x14394x) & (n_n3714) & (!x14403x) & (!x14404x)) + ((!x14393x) & (!x14394x) & (n_n3714) & (!x14403x) & (x14404x)) + ((!x14393x) & (!x14394x) & (n_n3714) & (x14403x) & (!x14404x)) + ((!x14393x) & (!x14394x) & (n_n3714) & (x14403x) & (x14404x)) + ((!x14393x) & (x14394x) & (!n_n3714) & (!x14403x) & (!x14404x)) + ((!x14393x) & (x14394x) & (!n_n3714) & (!x14403x) & (x14404x)) + ((!x14393x) & (x14394x) & (!n_n3714) & (x14403x) & (!x14404x)) + ((!x14393x) & (x14394x) & (!n_n3714) & (x14403x) & (x14404x)) + ((!x14393x) & (x14394x) & (n_n3714) & (!x14403x) & (!x14404x)) + ((!x14393x) & (x14394x) & (n_n3714) & (!x14403x) & (x14404x)) + ((!x14393x) & (x14394x) & (n_n3714) & (x14403x) & (!x14404x)) + ((!x14393x) & (x14394x) & (n_n3714) & (x14403x) & (x14404x)) + ((x14393x) & (!x14394x) & (!n_n3714) & (!x14403x) & (!x14404x)) + ((x14393x) & (!x14394x) & (!n_n3714) & (!x14403x) & (x14404x)) + ((x14393x) & (!x14394x) & (!n_n3714) & (x14403x) & (!x14404x)) + ((x14393x) & (!x14394x) & (!n_n3714) & (x14403x) & (x14404x)) + ((x14393x) & (!x14394x) & (n_n3714) & (!x14403x) & (!x14404x)) + ((x14393x) & (!x14394x) & (n_n3714) & (!x14403x) & (x14404x)) + ((x14393x) & (!x14394x) & (n_n3714) & (x14403x) & (!x14404x)) + ((x14393x) & (!x14394x) & (n_n3714) & (x14403x) & (x14404x)) + ((x14393x) & (x14394x) & (!n_n3714) & (!x14403x) & (!x14404x)) + ((x14393x) & (x14394x) & (!n_n3714) & (!x14403x) & (x14404x)) + ((x14393x) & (x14394x) & (!n_n3714) & (x14403x) & (!x14404x)) + ((x14393x) & (x14394x) & (!n_n3714) & (x14403x) & (x14404x)) + ((x14393x) & (x14394x) & (n_n3714) & (!x14403x) & (!x14404x)) + ((x14393x) & (x14394x) & (n_n3714) & (!x14403x) & (x14404x)) + ((x14393x) & (x14394x) & (n_n3714) & (x14403x) & (!x14404x)) + ((x14393x) & (x14394x) & (n_n3714) & (x14403x) & (x14404x)));
	assign n_n4550 = (((i_9_) & (n_n455) & (n_n473) & (n_n520)));
	assign n_n3870 = (((!i_9_) & (n_n524) & (n_n455) & (!n_n522) & (n_n464)) + ((!i_9_) & (n_n524) & (n_n455) & (n_n522) & (n_n464)) + ((i_9_) & (!n_n524) & (n_n455) & (n_n522) & (n_n464)) + ((i_9_) & (n_n524) & (n_n455) & (!n_n522) & (n_n464)) + ((i_9_) & (n_n524) & (n_n455) & (n_n522) & (n_n464)));
	assign x22214x = (((!n_n4539) & (!n_n4536) & (!n_n4545) & (!x13091x)));
	assign n_n3722 = (((!n_n4540) & (!n_n4541) & (!n_n4543) & (!n_n4537) & (!x22214x)) + ((!n_n4540) & (!n_n4541) & (!n_n4543) & (n_n4537) & (!x22214x)) + ((!n_n4540) & (!n_n4541) & (!n_n4543) & (n_n4537) & (x22214x)) + ((!n_n4540) & (!n_n4541) & (n_n4543) & (!n_n4537) & (!x22214x)) + ((!n_n4540) & (!n_n4541) & (n_n4543) & (!n_n4537) & (x22214x)) + ((!n_n4540) & (!n_n4541) & (n_n4543) & (n_n4537) & (!x22214x)) + ((!n_n4540) & (!n_n4541) & (n_n4543) & (n_n4537) & (x22214x)) + ((!n_n4540) & (n_n4541) & (!n_n4543) & (!n_n4537) & (!x22214x)) + ((!n_n4540) & (n_n4541) & (!n_n4543) & (!n_n4537) & (x22214x)) + ((!n_n4540) & (n_n4541) & (!n_n4543) & (n_n4537) & (!x22214x)) + ((!n_n4540) & (n_n4541) & (!n_n4543) & (n_n4537) & (x22214x)) + ((!n_n4540) & (n_n4541) & (n_n4543) & (!n_n4537) & (!x22214x)) + ((!n_n4540) & (n_n4541) & (n_n4543) & (!n_n4537) & (x22214x)) + ((!n_n4540) & (n_n4541) & (n_n4543) & (n_n4537) & (!x22214x)) + ((!n_n4540) & (n_n4541) & (n_n4543) & (n_n4537) & (x22214x)) + ((n_n4540) & (!n_n4541) & (!n_n4543) & (!n_n4537) & (!x22214x)) + ((n_n4540) & (!n_n4541) & (!n_n4543) & (!n_n4537) & (x22214x)) + ((n_n4540) & (!n_n4541) & (!n_n4543) & (n_n4537) & (!x22214x)) + ((n_n4540) & (!n_n4541) & (!n_n4543) & (n_n4537) & (x22214x)) + ((n_n4540) & (!n_n4541) & (n_n4543) & (!n_n4537) & (!x22214x)) + ((n_n4540) & (!n_n4541) & (n_n4543) & (!n_n4537) & (x22214x)) + ((n_n4540) & (!n_n4541) & (n_n4543) & (n_n4537) & (!x22214x)) + ((n_n4540) & (!n_n4541) & (n_n4543) & (n_n4537) & (x22214x)) + ((n_n4540) & (n_n4541) & (!n_n4543) & (!n_n4537) & (!x22214x)) + ((n_n4540) & (n_n4541) & (!n_n4543) & (!n_n4537) & (x22214x)) + ((n_n4540) & (n_n4541) & (!n_n4543) & (n_n4537) & (!x22214x)) + ((n_n4540) & (n_n4541) & (!n_n4543) & (n_n4537) & (x22214x)) + ((n_n4540) & (n_n4541) & (n_n4543) & (!n_n4537) & (!x22214x)) + ((n_n4540) & (n_n4541) & (n_n4543) & (!n_n4537) & (x22214x)) + ((n_n4540) & (n_n4541) & (n_n4543) & (n_n4537) & (!x22214x)) + ((n_n4540) & (n_n4541) & (n_n4543) & (n_n4537) & (x22214x)));
	assign x91x = (((i_9_) & (n_n455) & (n_n520) & (n_n464)));
	assign x214x = (((!i_9_) & (n_n455) & (!n_n528) & (n_n530) & (n_n464)) + ((!i_9_) & (n_n455) & (n_n528) & (n_n530) & (n_n464)) + ((i_9_) & (n_n455) & (n_n528) & (!n_n530) & (n_n464)) + ((i_9_) & (n_n455) & (n_n528) & (n_n530) & (n_n464)));
	assign x14416x = (((!x13x) & (!x506x) & (!n_n4569) & (!n_n4556) & (x91x)) + ((!x13x) & (!x506x) & (!n_n4569) & (n_n4556) & (!x91x)) + ((!x13x) & (!x506x) & (!n_n4569) & (n_n4556) & (x91x)) + ((!x13x) & (!x506x) & (n_n4569) & (!n_n4556) & (!x91x)) + ((!x13x) & (!x506x) & (n_n4569) & (!n_n4556) & (x91x)) + ((!x13x) & (!x506x) & (n_n4569) & (n_n4556) & (!x91x)) + ((!x13x) & (!x506x) & (n_n4569) & (n_n4556) & (x91x)) + ((!x13x) & (x506x) & (!n_n4569) & (!n_n4556) & (x91x)) + ((!x13x) & (x506x) & (!n_n4569) & (n_n4556) & (!x91x)) + ((!x13x) & (x506x) & (!n_n4569) & (n_n4556) & (x91x)) + ((!x13x) & (x506x) & (n_n4569) & (!n_n4556) & (!x91x)) + ((!x13x) & (x506x) & (n_n4569) & (!n_n4556) & (x91x)) + ((!x13x) & (x506x) & (n_n4569) & (n_n4556) & (!x91x)) + ((!x13x) & (x506x) & (n_n4569) & (n_n4556) & (x91x)) + ((x13x) & (!x506x) & (!n_n4569) & (!n_n4556) & (x91x)) + ((x13x) & (!x506x) & (!n_n4569) & (n_n4556) & (!x91x)) + ((x13x) & (!x506x) & (!n_n4569) & (n_n4556) & (x91x)) + ((x13x) & (!x506x) & (n_n4569) & (!n_n4556) & (!x91x)) + ((x13x) & (!x506x) & (n_n4569) & (!n_n4556) & (x91x)) + ((x13x) & (!x506x) & (n_n4569) & (n_n4556) & (!x91x)) + ((x13x) & (!x506x) & (n_n4569) & (n_n4556) & (x91x)) + ((x13x) & (x506x) & (!n_n4569) & (!n_n4556) & (!x91x)) + ((x13x) & (x506x) & (!n_n4569) & (!n_n4556) & (x91x)) + ((x13x) & (x506x) & (!n_n4569) & (n_n4556) & (!x91x)) + ((x13x) & (x506x) & (!n_n4569) & (n_n4556) & (x91x)) + ((x13x) & (x506x) & (n_n4569) & (!n_n4556) & (!x91x)) + ((x13x) & (x506x) & (n_n4569) & (!n_n4556) & (x91x)) + ((x13x) & (x506x) & (n_n4569) & (n_n4556) & (!x91x)) + ((x13x) & (x506x) & (n_n4569) & (n_n4556) & (x91x)));
	assign x14418x = (((!n_n4571) & (!n_n4560) & (!x212x) & (!x214x) & (x430x)) + ((!n_n4571) & (!n_n4560) & (!x212x) & (x214x) & (!x430x)) + ((!n_n4571) & (!n_n4560) & (!x212x) & (x214x) & (x430x)) + ((!n_n4571) & (!n_n4560) & (x212x) & (!x214x) & (!x430x)) + ((!n_n4571) & (!n_n4560) & (x212x) & (!x214x) & (x430x)) + ((!n_n4571) & (!n_n4560) & (x212x) & (x214x) & (!x430x)) + ((!n_n4571) & (!n_n4560) & (x212x) & (x214x) & (x430x)) + ((!n_n4571) & (n_n4560) & (!x212x) & (!x214x) & (!x430x)) + ((!n_n4571) & (n_n4560) & (!x212x) & (!x214x) & (x430x)) + ((!n_n4571) & (n_n4560) & (!x212x) & (x214x) & (!x430x)) + ((!n_n4571) & (n_n4560) & (!x212x) & (x214x) & (x430x)) + ((!n_n4571) & (n_n4560) & (x212x) & (!x214x) & (!x430x)) + ((!n_n4571) & (n_n4560) & (x212x) & (!x214x) & (x430x)) + ((!n_n4571) & (n_n4560) & (x212x) & (x214x) & (!x430x)) + ((!n_n4571) & (n_n4560) & (x212x) & (x214x) & (x430x)) + ((n_n4571) & (!n_n4560) & (!x212x) & (!x214x) & (!x430x)) + ((n_n4571) & (!n_n4560) & (!x212x) & (!x214x) & (x430x)) + ((n_n4571) & (!n_n4560) & (!x212x) & (x214x) & (!x430x)) + ((n_n4571) & (!n_n4560) & (!x212x) & (x214x) & (x430x)) + ((n_n4571) & (!n_n4560) & (x212x) & (!x214x) & (!x430x)) + ((n_n4571) & (!n_n4560) & (x212x) & (!x214x) & (x430x)) + ((n_n4571) & (!n_n4560) & (x212x) & (x214x) & (!x430x)) + ((n_n4571) & (!n_n4560) & (x212x) & (x214x) & (x430x)) + ((n_n4571) & (n_n4560) & (!x212x) & (!x214x) & (!x430x)) + ((n_n4571) & (n_n4560) & (!x212x) & (!x214x) & (x430x)) + ((n_n4571) & (n_n4560) & (!x212x) & (x214x) & (!x430x)) + ((n_n4571) & (n_n4560) & (!x212x) & (x214x) & (x430x)) + ((n_n4571) & (n_n4560) & (x212x) & (!x214x) & (!x430x)) + ((n_n4571) & (n_n4560) & (x212x) & (!x214x) & (x430x)) + ((n_n4571) & (n_n4560) & (x212x) & (x214x) & (!x430x)) + ((n_n4571) & (n_n4560) & (x212x) & (x214x) & (x430x)));
	assign n_n3652 = (((!n_n3871) & (!n_n3870) & (!n_n3722) & (!x14416x) & (x14418x)) + ((!n_n3871) & (!n_n3870) & (!n_n3722) & (x14416x) & (!x14418x)) + ((!n_n3871) & (!n_n3870) & (!n_n3722) & (x14416x) & (x14418x)) + ((!n_n3871) & (!n_n3870) & (n_n3722) & (!x14416x) & (!x14418x)) + ((!n_n3871) & (!n_n3870) & (n_n3722) & (!x14416x) & (x14418x)) + ((!n_n3871) & (!n_n3870) & (n_n3722) & (x14416x) & (!x14418x)) + ((!n_n3871) & (!n_n3870) & (n_n3722) & (x14416x) & (x14418x)) + ((!n_n3871) & (n_n3870) & (!n_n3722) & (!x14416x) & (!x14418x)) + ((!n_n3871) & (n_n3870) & (!n_n3722) & (!x14416x) & (x14418x)) + ((!n_n3871) & (n_n3870) & (!n_n3722) & (x14416x) & (!x14418x)) + ((!n_n3871) & (n_n3870) & (!n_n3722) & (x14416x) & (x14418x)) + ((!n_n3871) & (n_n3870) & (n_n3722) & (!x14416x) & (!x14418x)) + ((!n_n3871) & (n_n3870) & (n_n3722) & (!x14416x) & (x14418x)) + ((!n_n3871) & (n_n3870) & (n_n3722) & (x14416x) & (!x14418x)) + ((!n_n3871) & (n_n3870) & (n_n3722) & (x14416x) & (x14418x)) + ((n_n3871) & (!n_n3870) & (!n_n3722) & (!x14416x) & (!x14418x)) + ((n_n3871) & (!n_n3870) & (!n_n3722) & (!x14416x) & (x14418x)) + ((n_n3871) & (!n_n3870) & (!n_n3722) & (x14416x) & (!x14418x)) + ((n_n3871) & (!n_n3870) & (!n_n3722) & (x14416x) & (x14418x)) + ((n_n3871) & (!n_n3870) & (n_n3722) & (!x14416x) & (!x14418x)) + ((n_n3871) & (!n_n3870) & (n_n3722) & (!x14416x) & (x14418x)) + ((n_n3871) & (!n_n3870) & (n_n3722) & (x14416x) & (!x14418x)) + ((n_n3871) & (!n_n3870) & (n_n3722) & (x14416x) & (x14418x)) + ((n_n3871) & (n_n3870) & (!n_n3722) & (!x14416x) & (!x14418x)) + ((n_n3871) & (n_n3870) & (!n_n3722) & (!x14416x) & (x14418x)) + ((n_n3871) & (n_n3870) & (!n_n3722) & (x14416x) & (!x14418x)) + ((n_n3871) & (n_n3870) & (!n_n3722) & (x14416x) & (x14418x)) + ((n_n3871) & (n_n3870) & (n_n3722) & (!x14416x) & (!x14418x)) + ((n_n3871) & (n_n3870) & (n_n3722) & (!x14416x) & (x14418x)) + ((n_n3871) & (n_n3870) & (n_n3722) & (x14416x) & (!x14418x)) + ((n_n3871) & (n_n3870) & (n_n3722) & (x14416x) & (x14418x)));
	assign x14424x = (((!x20x) & (!x583x) & (!n_n4596) & (!x172x) & (n_n4588)) + ((!x20x) & (!x583x) & (!n_n4596) & (x172x) & (!n_n4588)) + ((!x20x) & (!x583x) & (!n_n4596) & (x172x) & (n_n4588)) + ((!x20x) & (!x583x) & (n_n4596) & (!x172x) & (!n_n4588)) + ((!x20x) & (!x583x) & (n_n4596) & (!x172x) & (n_n4588)) + ((!x20x) & (!x583x) & (n_n4596) & (x172x) & (!n_n4588)) + ((!x20x) & (!x583x) & (n_n4596) & (x172x) & (n_n4588)) + ((!x20x) & (x583x) & (!n_n4596) & (!x172x) & (n_n4588)) + ((!x20x) & (x583x) & (!n_n4596) & (x172x) & (!n_n4588)) + ((!x20x) & (x583x) & (!n_n4596) & (x172x) & (n_n4588)) + ((!x20x) & (x583x) & (n_n4596) & (!x172x) & (!n_n4588)) + ((!x20x) & (x583x) & (n_n4596) & (!x172x) & (n_n4588)) + ((!x20x) & (x583x) & (n_n4596) & (x172x) & (!n_n4588)) + ((!x20x) & (x583x) & (n_n4596) & (x172x) & (n_n4588)) + ((x20x) & (!x583x) & (!n_n4596) & (!x172x) & (n_n4588)) + ((x20x) & (!x583x) & (!n_n4596) & (x172x) & (!n_n4588)) + ((x20x) & (!x583x) & (!n_n4596) & (x172x) & (n_n4588)) + ((x20x) & (!x583x) & (n_n4596) & (!x172x) & (!n_n4588)) + ((x20x) & (!x583x) & (n_n4596) & (!x172x) & (n_n4588)) + ((x20x) & (!x583x) & (n_n4596) & (x172x) & (!n_n4588)) + ((x20x) & (!x583x) & (n_n4596) & (x172x) & (n_n4588)) + ((x20x) & (x583x) & (!n_n4596) & (!x172x) & (!n_n4588)) + ((x20x) & (x583x) & (!n_n4596) & (!x172x) & (n_n4588)) + ((x20x) & (x583x) & (!n_n4596) & (x172x) & (!n_n4588)) + ((x20x) & (x583x) & (!n_n4596) & (x172x) & (n_n4588)) + ((x20x) & (x583x) & (n_n4596) & (!x172x) & (!n_n4588)) + ((x20x) & (x583x) & (n_n4596) & (!x172x) & (n_n4588)) + ((x20x) & (x583x) & (n_n4596) & (x172x) & (!n_n4588)) + ((x20x) & (x583x) & (n_n4596) & (x172x) & (n_n4588)));
	assign x14429x = (((!n_n4587) & (!n_n4586) & (!n_n4574) & (!n_n4572) & (n_n4583)) + ((!n_n4587) & (!n_n4586) & (!n_n4574) & (n_n4572) & (!n_n4583)) + ((!n_n4587) & (!n_n4586) & (!n_n4574) & (n_n4572) & (n_n4583)) + ((!n_n4587) & (!n_n4586) & (n_n4574) & (!n_n4572) & (!n_n4583)) + ((!n_n4587) & (!n_n4586) & (n_n4574) & (!n_n4572) & (n_n4583)) + ((!n_n4587) & (!n_n4586) & (n_n4574) & (n_n4572) & (!n_n4583)) + ((!n_n4587) & (!n_n4586) & (n_n4574) & (n_n4572) & (n_n4583)) + ((!n_n4587) & (n_n4586) & (!n_n4574) & (!n_n4572) & (!n_n4583)) + ((!n_n4587) & (n_n4586) & (!n_n4574) & (!n_n4572) & (n_n4583)) + ((!n_n4587) & (n_n4586) & (!n_n4574) & (n_n4572) & (!n_n4583)) + ((!n_n4587) & (n_n4586) & (!n_n4574) & (n_n4572) & (n_n4583)) + ((!n_n4587) & (n_n4586) & (n_n4574) & (!n_n4572) & (!n_n4583)) + ((!n_n4587) & (n_n4586) & (n_n4574) & (!n_n4572) & (n_n4583)) + ((!n_n4587) & (n_n4586) & (n_n4574) & (n_n4572) & (!n_n4583)) + ((!n_n4587) & (n_n4586) & (n_n4574) & (n_n4572) & (n_n4583)) + ((n_n4587) & (!n_n4586) & (!n_n4574) & (!n_n4572) & (!n_n4583)) + ((n_n4587) & (!n_n4586) & (!n_n4574) & (!n_n4572) & (n_n4583)) + ((n_n4587) & (!n_n4586) & (!n_n4574) & (n_n4572) & (!n_n4583)) + ((n_n4587) & (!n_n4586) & (!n_n4574) & (n_n4572) & (n_n4583)) + ((n_n4587) & (!n_n4586) & (n_n4574) & (!n_n4572) & (!n_n4583)) + ((n_n4587) & (!n_n4586) & (n_n4574) & (!n_n4572) & (n_n4583)) + ((n_n4587) & (!n_n4586) & (n_n4574) & (n_n4572) & (!n_n4583)) + ((n_n4587) & (!n_n4586) & (n_n4574) & (n_n4572) & (n_n4583)) + ((n_n4587) & (n_n4586) & (!n_n4574) & (!n_n4572) & (!n_n4583)) + ((n_n4587) & (n_n4586) & (!n_n4574) & (!n_n4572) & (n_n4583)) + ((n_n4587) & (n_n4586) & (!n_n4574) & (n_n4572) & (!n_n4583)) + ((n_n4587) & (n_n4586) & (!n_n4574) & (n_n4572) & (n_n4583)) + ((n_n4587) & (n_n4586) & (n_n4574) & (!n_n4572) & (!n_n4583)) + ((n_n4587) & (n_n4586) & (n_n4574) & (!n_n4572) & (n_n4583)) + ((n_n4587) & (n_n4586) & (n_n4574) & (n_n4572) & (!n_n4583)) + ((n_n4587) & (n_n4586) & (n_n4574) & (n_n4572) & (n_n4583)));
	assign n_n3719 = (((!n_n4578) & (!n_n4575) & (!n_n4577) & (!n_n4576) & (x14429x)) + ((!n_n4578) & (!n_n4575) & (!n_n4577) & (n_n4576) & (!x14429x)) + ((!n_n4578) & (!n_n4575) & (!n_n4577) & (n_n4576) & (x14429x)) + ((!n_n4578) & (!n_n4575) & (n_n4577) & (!n_n4576) & (!x14429x)) + ((!n_n4578) & (!n_n4575) & (n_n4577) & (!n_n4576) & (x14429x)) + ((!n_n4578) & (!n_n4575) & (n_n4577) & (n_n4576) & (!x14429x)) + ((!n_n4578) & (!n_n4575) & (n_n4577) & (n_n4576) & (x14429x)) + ((!n_n4578) & (n_n4575) & (!n_n4577) & (!n_n4576) & (!x14429x)) + ((!n_n4578) & (n_n4575) & (!n_n4577) & (!n_n4576) & (x14429x)) + ((!n_n4578) & (n_n4575) & (!n_n4577) & (n_n4576) & (!x14429x)) + ((!n_n4578) & (n_n4575) & (!n_n4577) & (n_n4576) & (x14429x)) + ((!n_n4578) & (n_n4575) & (n_n4577) & (!n_n4576) & (!x14429x)) + ((!n_n4578) & (n_n4575) & (n_n4577) & (!n_n4576) & (x14429x)) + ((!n_n4578) & (n_n4575) & (n_n4577) & (n_n4576) & (!x14429x)) + ((!n_n4578) & (n_n4575) & (n_n4577) & (n_n4576) & (x14429x)) + ((n_n4578) & (!n_n4575) & (!n_n4577) & (!n_n4576) & (!x14429x)) + ((n_n4578) & (!n_n4575) & (!n_n4577) & (!n_n4576) & (x14429x)) + ((n_n4578) & (!n_n4575) & (!n_n4577) & (n_n4576) & (!x14429x)) + ((n_n4578) & (!n_n4575) & (!n_n4577) & (n_n4576) & (x14429x)) + ((n_n4578) & (!n_n4575) & (n_n4577) & (!n_n4576) & (!x14429x)) + ((n_n4578) & (!n_n4575) & (n_n4577) & (!n_n4576) & (x14429x)) + ((n_n4578) & (!n_n4575) & (n_n4577) & (n_n4576) & (!x14429x)) + ((n_n4578) & (!n_n4575) & (n_n4577) & (n_n4576) & (x14429x)) + ((n_n4578) & (n_n4575) & (!n_n4577) & (!n_n4576) & (!x14429x)) + ((n_n4578) & (n_n4575) & (!n_n4577) & (!n_n4576) & (x14429x)) + ((n_n4578) & (n_n4575) & (!n_n4577) & (n_n4576) & (!x14429x)) + ((n_n4578) & (n_n4575) & (!n_n4577) & (n_n4576) & (x14429x)) + ((n_n4578) & (n_n4575) & (n_n4577) & (!n_n4576) & (!x14429x)) + ((n_n4578) & (n_n4575) & (n_n4577) & (!n_n4576) & (x14429x)) + ((n_n4578) & (n_n4575) & (n_n4577) & (n_n4576) & (!x14429x)) + ((n_n4578) & (n_n4575) & (n_n4577) & (n_n4576) & (x14429x)));
	assign x46x = (((!i_9_) & (!n_n524) & (n_n518) & (n_n526) & (n_n390)) + ((!i_9_) & (n_n524) & (n_n518) & (n_n526) & (n_n390)) + ((i_9_) & (n_n524) & (n_n518) & (!n_n526) & (n_n390)) + ((i_9_) & (n_n524) & (n_n518) & (n_n526) & (n_n390)));
	assign x14434x = (((!n_n4609) & (!n_n4614) & (!n_n2037) & (!x22168x)) + ((!n_n4609) & (!n_n4614) & (n_n2037) & (!x22168x)) + ((!n_n4609) & (!n_n4614) & (n_n2037) & (x22168x)) + ((!n_n4609) & (n_n4614) & (!n_n2037) & (!x22168x)) + ((!n_n4609) & (n_n4614) & (!n_n2037) & (x22168x)) + ((!n_n4609) & (n_n4614) & (n_n2037) & (!x22168x)) + ((!n_n4609) & (n_n4614) & (n_n2037) & (x22168x)) + ((n_n4609) & (!n_n4614) & (!n_n2037) & (!x22168x)) + ((n_n4609) & (!n_n4614) & (!n_n2037) & (x22168x)) + ((n_n4609) & (!n_n4614) & (n_n2037) & (!x22168x)) + ((n_n4609) & (!n_n4614) & (n_n2037) & (x22168x)) + ((n_n4609) & (n_n4614) & (!n_n2037) & (!x22168x)) + ((n_n4609) & (n_n4614) & (!n_n2037) & (x22168x)) + ((n_n4609) & (n_n4614) & (n_n2037) & (!x22168x)) + ((n_n4609) & (n_n4614) & (n_n2037) & (x22168x)));
	assign x14436x = (((!x45x) & (!x14424x) & (!n_n3719) & (!x46x) & (x14434x)) + ((!x45x) & (!x14424x) & (!n_n3719) & (x46x) & (!x14434x)) + ((!x45x) & (!x14424x) & (!n_n3719) & (x46x) & (x14434x)) + ((!x45x) & (!x14424x) & (n_n3719) & (!x46x) & (!x14434x)) + ((!x45x) & (!x14424x) & (n_n3719) & (!x46x) & (x14434x)) + ((!x45x) & (!x14424x) & (n_n3719) & (x46x) & (!x14434x)) + ((!x45x) & (!x14424x) & (n_n3719) & (x46x) & (x14434x)) + ((!x45x) & (x14424x) & (!n_n3719) & (!x46x) & (!x14434x)) + ((!x45x) & (x14424x) & (!n_n3719) & (!x46x) & (x14434x)) + ((!x45x) & (x14424x) & (!n_n3719) & (x46x) & (!x14434x)) + ((!x45x) & (x14424x) & (!n_n3719) & (x46x) & (x14434x)) + ((!x45x) & (x14424x) & (n_n3719) & (!x46x) & (!x14434x)) + ((!x45x) & (x14424x) & (n_n3719) & (!x46x) & (x14434x)) + ((!x45x) & (x14424x) & (n_n3719) & (x46x) & (!x14434x)) + ((!x45x) & (x14424x) & (n_n3719) & (x46x) & (x14434x)) + ((x45x) & (!x14424x) & (!n_n3719) & (!x46x) & (!x14434x)) + ((x45x) & (!x14424x) & (!n_n3719) & (!x46x) & (x14434x)) + ((x45x) & (!x14424x) & (!n_n3719) & (x46x) & (!x14434x)) + ((x45x) & (!x14424x) & (!n_n3719) & (x46x) & (x14434x)) + ((x45x) & (!x14424x) & (n_n3719) & (!x46x) & (!x14434x)) + ((x45x) & (!x14424x) & (n_n3719) & (!x46x) & (x14434x)) + ((x45x) & (!x14424x) & (n_n3719) & (x46x) & (!x14434x)) + ((x45x) & (!x14424x) & (n_n3719) & (x46x) & (x14434x)) + ((x45x) & (x14424x) & (!n_n3719) & (!x46x) & (!x14434x)) + ((x45x) & (x14424x) & (!n_n3719) & (!x46x) & (x14434x)) + ((x45x) & (x14424x) & (!n_n3719) & (x46x) & (!x14434x)) + ((x45x) & (x14424x) & (!n_n3719) & (x46x) & (x14434x)) + ((x45x) & (x14424x) & (n_n3719) & (!x46x) & (!x14434x)) + ((x45x) & (x14424x) & (n_n3719) & (!x46x) & (x14434x)) + ((x45x) & (x14424x) & (n_n3719) & (x46x) & (!x14434x)) + ((x45x) & (x14424x) & (n_n3719) & (x46x) & (x14434x)));
	assign n_n3461 = (((!i_9_) & (!n_n526) & (n_n528) & (n_n260) & (n_n535)) + ((!i_9_) & (n_n526) & (!n_n528) & (n_n260) & (n_n535)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n260) & (n_n535)) + ((i_9_) & (n_n526) & (!n_n528) & (n_n260) & (n_n535)) + ((i_9_) & (n_n526) & (n_n528) & (n_n260) & (n_n535)));
	assign n_n3329 = (((!n_n3460) & (!n_n4838) & (!n_n4841) & (!n_n4840) & (n_n3461)) + ((!n_n3460) & (!n_n4838) & (!n_n4841) & (n_n4840) & (!n_n3461)) + ((!n_n3460) & (!n_n4838) & (!n_n4841) & (n_n4840) & (n_n3461)) + ((!n_n3460) & (!n_n4838) & (n_n4841) & (!n_n4840) & (!n_n3461)) + ((!n_n3460) & (!n_n4838) & (n_n4841) & (!n_n4840) & (n_n3461)) + ((!n_n3460) & (!n_n4838) & (n_n4841) & (n_n4840) & (!n_n3461)) + ((!n_n3460) & (!n_n4838) & (n_n4841) & (n_n4840) & (n_n3461)) + ((!n_n3460) & (n_n4838) & (!n_n4841) & (!n_n4840) & (!n_n3461)) + ((!n_n3460) & (n_n4838) & (!n_n4841) & (!n_n4840) & (n_n3461)) + ((!n_n3460) & (n_n4838) & (!n_n4841) & (n_n4840) & (!n_n3461)) + ((!n_n3460) & (n_n4838) & (!n_n4841) & (n_n4840) & (n_n3461)) + ((!n_n3460) & (n_n4838) & (n_n4841) & (!n_n4840) & (!n_n3461)) + ((!n_n3460) & (n_n4838) & (n_n4841) & (!n_n4840) & (n_n3461)) + ((!n_n3460) & (n_n4838) & (n_n4841) & (n_n4840) & (!n_n3461)) + ((!n_n3460) & (n_n4838) & (n_n4841) & (n_n4840) & (n_n3461)) + ((n_n3460) & (!n_n4838) & (!n_n4841) & (!n_n4840) & (!n_n3461)) + ((n_n3460) & (!n_n4838) & (!n_n4841) & (!n_n4840) & (n_n3461)) + ((n_n3460) & (!n_n4838) & (!n_n4841) & (n_n4840) & (!n_n3461)) + ((n_n3460) & (!n_n4838) & (!n_n4841) & (n_n4840) & (n_n3461)) + ((n_n3460) & (!n_n4838) & (n_n4841) & (!n_n4840) & (!n_n3461)) + ((n_n3460) & (!n_n4838) & (n_n4841) & (!n_n4840) & (n_n3461)) + ((n_n3460) & (!n_n4838) & (n_n4841) & (n_n4840) & (!n_n3461)) + ((n_n3460) & (!n_n4838) & (n_n4841) & (n_n4840) & (n_n3461)) + ((n_n3460) & (n_n4838) & (!n_n4841) & (!n_n4840) & (!n_n3461)) + ((n_n3460) & (n_n4838) & (!n_n4841) & (!n_n4840) & (n_n3461)) + ((n_n3460) & (n_n4838) & (!n_n4841) & (n_n4840) & (!n_n3461)) + ((n_n3460) & (n_n4838) & (!n_n4841) & (n_n4840) & (n_n3461)) + ((n_n3460) & (n_n4838) & (n_n4841) & (!n_n4840) & (!n_n3461)) + ((n_n3460) & (n_n4838) & (n_n4841) & (!n_n4840) & (n_n3461)) + ((n_n3460) & (n_n4838) & (n_n4841) & (n_n4840) & (!n_n3461)) + ((n_n3460) & (n_n4838) & (n_n4841) & (n_n4840) & (n_n3461)));
	assign x13924x = (((!n_n509) & (!n_n522) & (!x12x) & (!n_n5127) & (x155x)) + ((!n_n509) & (!n_n522) & (!x12x) & (n_n5127) & (!x155x)) + ((!n_n509) & (!n_n522) & (!x12x) & (n_n5127) & (x155x)) + ((!n_n509) & (!n_n522) & (x12x) & (!n_n5127) & (x155x)) + ((!n_n509) & (!n_n522) & (x12x) & (n_n5127) & (!x155x)) + ((!n_n509) & (!n_n522) & (x12x) & (n_n5127) & (x155x)) + ((!n_n509) & (n_n522) & (!x12x) & (!n_n5127) & (x155x)) + ((!n_n509) & (n_n522) & (!x12x) & (n_n5127) & (!x155x)) + ((!n_n509) & (n_n522) & (!x12x) & (n_n5127) & (x155x)) + ((!n_n509) & (n_n522) & (x12x) & (!n_n5127) & (x155x)) + ((!n_n509) & (n_n522) & (x12x) & (n_n5127) & (!x155x)) + ((!n_n509) & (n_n522) & (x12x) & (n_n5127) & (x155x)) + ((n_n509) & (!n_n522) & (!x12x) & (!n_n5127) & (x155x)) + ((n_n509) & (!n_n522) & (!x12x) & (n_n5127) & (!x155x)) + ((n_n509) & (!n_n522) & (!x12x) & (n_n5127) & (x155x)) + ((n_n509) & (!n_n522) & (x12x) & (!n_n5127) & (x155x)) + ((n_n509) & (!n_n522) & (x12x) & (n_n5127) & (!x155x)) + ((n_n509) & (!n_n522) & (x12x) & (n_n5127) & (x155x)) + ((n_n509) & (n_n522) & (!x12x) & (!n_n5127) & (x155x)) + ((n_n509) & (n_n522) & (!x12x) & (n_n5127) & (!x155x)) + ((n_n509) & (n_n522) & (!x12x) & (n_n5127) & (x155x)) + ((n_n509) & (n_n522) & (x12x) & (!n_n5127) & (!x155x)) + ((n_n509) & (n_n522) & (x12x) & (!n_n5127) & (x155x)) + ((n_n509) & (n_n522) & (x12x) & (n_n5127) & (!x155x)) + ((n_n509) & (n_n522) & (x12x) & (n_n5127) & (x155x)));
	assign x13925x = (((!n_n5121) & (!n_n5122) & (!n_n5128) & (!n_n5125) & (n_n5126)) + ((!n_n5121) & (!n_n5122) & (!n_n5128) & (n_n5125) & (!n_n5126)) + ((!n_n5121) & (!n_n5122) & (!n_n5128) & (n_n5125) & (n_n5126)) + ((!n_n5121) & (!n_n5122) & (n_n5128) & (!n_n5125) & (!n_n5126)) + ((!n_n5121) & (!n_n5122) & (n_n5128) & (!n_n5125) & (n_n5126)) + ((!n_n5121) & (!n_n5122) & (n_n5128) & (n_n5125) & (!n_n5126)) + ((!n_n5121) & (!n_n5122) & (n_n5128) & (n_n5125) & (n_n5126)) + ((!n_n5121) & (n_n5122) & (!n_n5128) & (!n_n5125) & (!n_n5126)) + ((!n_n5121) & (n_n5122) & (!n_n5128) & (!n_n5125) & (n_n5126)) + ((!n_n5121) & (n_n5122) & (!n_n5128) & (n_n5125) & (!n_n5126)) + ((!n_n5121) & (n_n5122) & (!n_n5128) & (n_n5125) & (n_n5126)) + ((!n_n5121) & (n_n5122) & (n_n5128) & (!n_n5125) & (!n_n5126)) + ((!n_n5121) & (n_n5122) & (n_n5128) & (!n_n5125) & (n_n5126)) + ((!n_n5121) & (n_n5122) & (n_n5128) & (n_n5125) & (!n_n5126)) + ((!n_n5121) & (n_n5122) & (n_n5128) & (n_n5125) & (n_n5126)) + ((n_n5121) & (!n_n5122) & (!n_n5128) & (!n_n5125) & (!n_n5126)) + ((n_n5121) & (!n_n5122) & (!n_n5128) & (!n_n5125) & (n_n5126)) + ((n_n5121) & (!n_n5122) & (!n_n5128) & (n_n5125) & (!n_n5126)) + ((n_n5121) & (!n_n5122) & (!n_n5128) & (n_n5125) & (n_n5126)) + ((n_n5121) & (!n_n5122) & (n_n5128) & (!n_n5125) & (!n_n5126)) + ((n_n5121) & (!n_n5122) & (n_n5128) & (!n_n5125) & (n_n5126)) + ((n_n5121) & (!n_n5122) & (n_n5128) & (n_n5125) & (!n_n5126)) + ((n_n5121) & (!n_n5122) & (n_n5128) & (n_n5125) & (n_n5126)) + ((n_n5121) & (n_n5122) & (!n_n5128) & (!n_n5125) & (!n_n5126)) + ((n_n5121) & (n_n5122) & (!n_n5128) & (!n_n5125) & (n_n5126)) + ((n_n5121) & (n_n5122) & (!n_n5128) & (n_n5125) & (!n_n5126)) + ((n_n5121) & (n_n5122) & (!n_n5128) & (n_n5125) & (n_n5126)) + ((n_n5121) & (n_n5122) & (n_n5128) & (!n_n5125) & (!n_n5126)) + ((n_n5121) & (n_n5122) & (n_n5128) & (!n_n5125) & (n_n5126)) + ((n_n5121) & (n_n5122) & (n_n5128) & (n_n5125) & (!n_n5126)) + ((n_n5121) & (n_n5122) & (n_n5128) & (n_n5125) & (n_n5126)));
	assign x13793x = (((!n_n325) & (!x23x) & (!n_n500) & (!n_n2130) & (n_n4764)) + ((!n_n325) & (!x23x) & (!n_n500) & (n_n2130) & (!n_n4764)) + ((!n_n325) & (!x23x) & (!n_n500) & (n_n2130) & (n_n4764)) + ((!n_n325) & (!x23x) & (n_n500) & (!n_n2130) & (n_n4764)) + ((!n_n325) & (!x23x) & (n_n500) & (n_n2130) & (!n_n4764)) + ((!n_n325) & (!x23x) & (n_n500) & (n_n2130) & (n_n4764)) + ((!n_n325) & (x23x) & (!n_n500) & (!n_n2130) & (n_n4764)) + ((!n_n325) & (x23x) & (!n_n500) & (n_n2130) & (!n_n4764)) + ((!n_n325) & (x23x) & (!n_n500) & (n_n2130) & (n_n4764)) + ((!n_n325) & (x23x) & (n_n500) & (!n_n2130) & (n_n4764)) + ((!n_n325) & (x23x) & (n_n500) & (n_n2130) & (!n_n4764)) + ((!n_n325) & (x23x) & (n_n500) & (n_n2130) & (n_n4764)) + ((n_n325) & (!x23x) & (!n_n500) & (!n_n2130) & (n_n4764)) + ((n_n325) & (!x23x) & (!n_n500) & (n_n2130) & (!n_n4764)) + ((n_n325) & (!x23x) & (!n_n500) & (n_n2130) & (n_n4764)) + ((n_n325) & (!x23x) & (n_n500) & (!n_n2130) & (n_n4764)) + ((n_n325) & (!x23x) & (n_n500) & (n_n2130) & (!n_n4764)) + ((n_n325) & (!x23x) & (n_n500) & (n_n2130) & (n_n4764)) + ((n_n325) & (x23x) & (!n_n500) & (!n_n2130) & (n_n4764)) + ((n_n325) & (x23x) & (!n_n500) & (n_n2130) & (!n_n4764)) + ((n_n325) & (x23x) & (!n_n500) & (n_n2130) & (n_n4764)) + ((n_n325) & (x23x) & (n_n500) & (!n_n2130) & (!n_n4764)) + ((n_n325) & (x23x) & (n_n500) & (!n_n2130) & (n_n4764)) + ((n_n325) & (x23x) & (n_n500) & (n_n2130) & (!n_n4764)) + ((n_n325) & (x23x) & (n_n500) & (n_n2130) & (n_n4764)));
	assign x13795x = (((!n_n4761) & (!n_n4762) & (!n_n4765) & (!x164x) & (x370x)) + ((!n_n4761) & (!n_n4762) & (!n_n4765) & (x164x) & (!x370x)) + ((!n_n4761) & (!n_n4762) & (!n_n4765) & (x164x) & (x370x)) + ((!n_n4761) & (!n_n4762) & (n_n4765) & (!x164x) & (!x370x)) + ((!n_n4761) & (!n_n4762) & (n_n4765) & (!x164x) & (x370x)) + ((!n_n4761) & (!n_n4762) & (n_n4765) & (x164x) & (!x370x)) + ((!n_n4761) & (!n_n4762) & (n_n4765) & (x164x) & (x370x)) + ((!n_n4761) & (n_n4762) & (!n_n4765) & (!x164x) & (!x370x)) + ((!n_n4761) & (n_n4762) & (!n_n4765) & (!x164x) & (x370x)) + ((!n_n4761) & (n_n4762) & (!n_n4765) & (x164x) & (!x370x)) + ((!n_n4761) & (n_n4762) & (!n_n4765) & (x164x) & (x370x)) + ((!n_n4761) & (n_n4762) & (n_n4765) & (!x164x) & (!x370x)) + ((!n_n4761) & (n_n4762) & (n_n4765) & (!x164x) & (x370x)) + ((!n_n4761) & (n_n4762) & (n_n4765) & (x164x) & (!x370x)) + ((!n_n4761) & (n_n4762) & (n_n4765) & (x164x) & (x370x)) + ((n_n4761) & (!n_n4762) & (!n_n4765) & (!x164x) & (!x370x)) + ((n_n4761) & (!n_n4762) & (!n_n4765) & (!x164x) & (x370x)) + ((n_n4761) & (!n_n4762) & (!n_n4765) & (x164x) & (!x370x)) + ((n_n4761) & (!n_n4762) & (!n_n4765) & (x164x) & (x370x)) + ((n_n4761) & (!n_n4762) & (n_n4765) & (!x164x) & (!x370x)) + ((n_n4761) & (!n_n4762) & (n_n4765) & (!x164x) & (x370x)) + ((n_n4761) & (!n_n4762) & (n_n4765) & (x164x) & (!x370x)) + ((n_n4761) & (!n_n4762) & (n_n4765) & (x164x) & (x370x)) + ((n_n4761) & (n_n4762) & (!n_n4765) & (!x164x) & (!x370x)) + ((n_n4761) & (n_n4762) & (!n_n4765) & (!x164x) & (x370x)) + ((n_n4761) & (n_n4762) & (!n_n4765) & (x164x) & (!x370x)) + ((n_n4761) & (n_n4762) & (!n_n4765) & (x164x) & (x370x)) + ((n_n4761) & (n_n4762) & (n_n4765) & (!x164x) & (!x370x)) + ((n_n4761) & (n_n4762) & (n_n4765) & (!x164x) & (x370x)) + ((n_n4761) & (n_n4762) & (n_n4765) & (x164x) & (!x370x)) + ((n_n4761) & (n_n4762) & (n_n4765) & (x164x) & (x370x)));
	assign n_n3277 = (((!n_n4204) & (!n_n3469) & (!n_n3333) & (!x13793x) & (x13795x)) + ((!n_n4204) & (!n_n3469) & (!n_n3333) & (x13793x) & (!x13795x)) + ((!n_n4204) & (!n_n3469) & (!n_n3333) & (x13793x) & (x13795x)) + ((!n_n4204) & (!n_n3469) & (n_n3333) & (!x13793x) & (!x13795x)) + ((!n_n4204) & (!n_n3469) & (n_n3333) & (!x13793x) & (x13795x)) + ((!n_n4204) & (!n_n3469) & (n_n3333) & (x13793x) & (!x13795x)) + ((!n_n4204) & (!n_n3469) & (n_n3333) & (x13793x) & (x13795x)) + ((!n_n4204) & (n_n3469) & (!n_n3333) & (!x13793x) & (!x13795x)) + ((!n_n4204) & (n_n3469) & (!n_n3333) & (!x13793x) & (x13795x)) + ((!n_n4204) & (n_n3469) & (!n_n3333) & (x13793x) & (!x13795x)) + ((!n_n4204) & (n_n3469) & (!n_n3333) & (x13793x) & (x13795x)) + ((!n_n4204) & (n_n3469) & (n_n3333) & (!x13793x) & (!x13795x)) + ((!n_n4204) & (n_n3469) & (n_n3333) & (!x13793x) & (x13795x)) + ((!n_n4204) & (n_n3469) & (n_n3333) & (x13793x) & (!x13795x)) + ((!n_n4204) & (n_n3469) & (n_n3333) & (x13793x) & (x13795x)) + ((n_n4204) & (!n_n3469) & (!n_n3333) & (!x13793x) & (!x13795x)) + ((n_n4204) & (!n_n3469) & (!n_n3333) & (!x13793x) & (x13795x)) + ((n_n4204) & (!n_n3469) & (!n_n3333) & (x13793x) & (!x13795x)) + ((n_n4204) & (!n_n3469) & (!n_n3333) & (x13793x) & (x13795x)) + ((n_n4204) & (!n_n3469) & (n_n3333) & (!x13793x) & (!x13795x)) + ((n_n4204) & (!n_n3469) & (n_n3333) & (!x13793x) & (x13795x)) + ((n_n4204) & (!n_n3469) & (n_n3333) & (x13793x) & (!x13795x)) + ((n_n4204) & (!n_n3469) & (n_n3333) & (x13793x) & (x13795x)) + ((n_n4204) & (n_n3469) & (!n_n3333) & (!x13793x) & (!x13795x)) + ((n_n4204) & (n_n3469) & (!n_n3333) & (!x13793x) & (x13795x)) + ((n_n4204) & (n_n3469) & (!n_n3333) & (x13793x) & (!x13795x)) + ((n_n4204) & (n_n3469) & (!n_n3333) & (x13793x) & (x13795x)) + ((n_n4204) & (n_n3469) & (n_n3333) & (!x13793x) & (!x13795x)) + ((n_n4204) & (n_n3469) & (n_n3333) & (!x13793x) & (x13795x)) + ((n_n4204) & (n_n3469) & (n_n3333) & (x13793x) & (!x13795x)) + ((n_n4204) & (n_n3469) & (n_n3333) & (x13793x) & (x13795x)));
	assign n_n4808 = (((i_9_) & (n_n534) & (n_n325) & (n_n464)));
	assign x380x = (((!i_7_) & (!i_8_) & (i_6_) & (n_n473) & (x14x)) + ((!i_7_) & (i_8_) & (i_6_) & (n_n473) & (x14x)));
	assign x381x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n473) & (n_n325)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n473) & (n_n325)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n473) & (n_n325)) + ((i_9_) & (n_n524) & (n_n526) & (n_n473) & (n_n325)));
	assign x13799x = (((!i_9_) & (n_n473) & (!n_n532) & (n_n534) & (n_n325)) + ((!i_9_) & (n_n473) & (n_n532) & (!n_n534) & (n_n325)) + ((!i_9_) & (n_n473) & (n_n532) & (n_n534) & (n_n325)) + ((i_9_) & (n_n473) & (!n_n532) & (n_n534) & (n_n325)) + ((i_9_) & (n_n473) & (n_n532) & (n_n534) & (n_n325)));
	assign n_n3332 = (((!n_n4800) & (!n_n4794) & (!x380x) & (!x381x) & (x13799x)) + ((!n_n4800) & (!n_n4794) & (!x380x) & (x381x) & (!x13799x)) + ((!n_n4800) & (!n_n4794) & (!x380x) & (x381x) & (x13799x)) + ((!n_n4800) & (!n_n4794) & (x380x) & (!x381x) & (!x13799x)) + ((!n_n4800) & (!n_n4794) & (x380x) & (!x381x) & (x13799x)) + ((!n_n4800) & (!n_n4794) & (x380x) & (x381x) & (!x13799x)) + ((!n_n4800) & (!n_n4794) & (x380x) & (x381x) & (x13799x)) + ((!n_n4800) & (n_n4794) & (!x380x) & (!x381x) & (!x13799x)) + ((!n_n4800) & (n_n4794) & (!x380x) & (!x381x) & (x13799x)) + ((!n_n4800) & (n_n4794) & (!x380x) & (x381x) & (!x13799x)) + ((!n_n4800) & (n_n4794) & (!x380x) & (x381x) & (x13799x)) + ((!n_n4800) & (n_n4794) & (x380x) & (!x381x) & (!x13799x)) + ((!n_n4800) & (n_n4794) & (x380x) & (!x381x) & (x13799x)) + ((!n_n4800) & (n_n4794) & (x380x) & (x381x) & (!x13799x)) + ((!n_n4800) & (n_n4794) & (x380x) & (x381x) & (x13799x)) + ((n_n4800) & (!n_n4794) & (!x380x) & (!x381x) & (!x13799x)) + ((n_n4800) & (!n_n4794) & (!x380x) & (!x381x) & (x13799x)) + ((n_n4800) & (!n_n4794) & (!x380x) & (x381x) & (!x13799x)) + ((n_n4800) & (!n_n4794) & (!x380x) & (x381x) & (x13799x)) + ((n_n4800) & (!n_n4794) & (x380x) & (!x381x) & (!x13799x)) + ((n_n4800) & (!n_n4794) & (x380x) & (!x381x) & (x13799x)) + ((n_n4800) & (!n_n4794) & (x380x) & (x381x) & (!x13799x)) + ((n_n4800) & (!n_n4794) & (x380x) & (x381x) & (x13799x)) + ((n_n4800) & (n_n4794) & (!x380x) & (!x381x) & (!x13799x)) + ((n_n4800) & (n_n4794) & (!x380x) & (!x381x) & (x13799x)) + ((n_n4800) & (n_n4794) & (!x380x) & (x381x) & (!x13799x)) + ((n_n4800) & (n_n4794) & (!x380x) & (x381x) & (x13799x)) + ((n_n4800) & (n_n4794) & (x380x) & (!x381x) & (!x13799x)) + ((n_n4800) & (n_n4794) & (x380x) & (!x381x) & (x13799x)) + ((n_n4800) & (n_n4794) & (x380x) & (x381x) & (!x13799x)) + ((n_n4800) & (n_n4794) & (x380x) & (x381x) & (x13799x)));
	assign x13805x = (((!n_n4827) & (!n_n4825) & (!n_n4826) & (!n_n4822) & (n_n4815)) + ((!n_n4827) & (!n_n4825) & (!n_n4826) & (n_n4822) & (!n_n4815)) + ((!n_n4827) & (!n_n4825) & (!n_n4826) & (n_n4822) & (n_n4815)) + ((!n_n4827) & (!n_n4825) & (n_n4826) & (!n_n4822) & (!n_n4815)) + ((!n_n4827) & (!n_n4825) & (n_n4826) & (!n_n4822) & (n_n4815)) + ((!n_n4827) & (!n_n4825) & (n_n4826) & (n_n4822) & (!n_n4815)) + ((!n_n4827) & (!n_n4825) & (n_n4826) & (n_n4822) & (n_n4815)) + ((!n_n4827) & (n_n4825) & (!n_n4826) & (!n_n4822) & (!n_n4815)) + ((!n_n4827) & (n_n4825) & (!n_n4826) & (!n_n4822) & (n_n4815)) + ((!n_n4827) & (n_n4825) & (!n_n4826) & (n_n4822) & (!n_n4815)) + ((!n_n4827) & (n_n4825) & (!n_n4826) & (n_n4822) & (n_n4815)) + ((!n_n4827) & (n_n4825) & (n_n4826) & (!n_n4822) & (!n_n4815)) + ((!n_n4827) & (n_n4825) & (n_n4826) & (!n_n4822) & (n_n4815)) + ((!n_n4827) & (n_n4825) & (n_n4826) & (n_n4822) & (!n_n4815)) + ((!n_n4827) & (n_n4825) & (n_n4826) & (n_n4822) & (n_n4815)) + ((n_n4827) & (!n_n4825) & (!n_n4826) & (!n_n4822) & (!n_n4815)) + ((n_n4827) & (!n_n4825) & (!n_n4826) & (!n_n4822) & (n_n4815)) + ((n_n4827) & (!n_n4825) & (!n_n4826) & (n_n4822) & (!n_n4815)) + ((n_n4827) & (!n_n4825) & (!n_n4826) & (n_n4822) & (n_n4815)) + ((n_n4827) & (!n_n4825) & (n_n4826) & (!n_n4822) & (!n_n4815)) + ((n_n4827) & (!n_n4825) & (n_n4826) & (!n_n4822) & (n_n4815)) + ((n_n4827) & (!n_n4825) & (n_n4826) & (n_n4822) & (!n_n4815)) + ((n_n4827) & (!n_n4825) & (n_n4826) & (n_n4822) & (n_n4815)) + ((n_n4827) & (n_n4825) & (!n_n4826) & (!n_n4822) & (!n_n4815)) + ((n_n4827) & (n_n4825) & (!n_n4826) & (!n_n4822) & (n_n4815)) + ((n_n4827) & (n_n4825) & (!n_n4826) & (n_n4822) & (!n_n4815)) + ((n_n4827) & (n_n4825) & (!n_n4826) & (n_n4822) & (n_n4815)) + ((n_n4827) & (n_n4825) & (n_n4826) & (!n_n4822) & (!n_n4815)) + ((n_n4827) & (n_n4825) & (n_n4826) & (!n_n4822) & (n_n4815)) + ((n_n4827) & (n_n4825) & (n_n4826) & (n_n4822) & (!n_n4815)) + ((n_n4827) & (n_n4825) & (n_n4826) & (n_n4822) & (n_n4815)));
	assign x22116x = (((!n_n4856) & (!n_n4850) & (!n_n4843) & (!n_n4845)));
	assign x13820x = (((!x102x) & (!n_n4852) & (!n_n4846) & (!n_n4848) & (!x22116x)) + ((!x102x) & (!n_n4852) & (!n_n4846) & (n_n4848) & (!x22116x)) + ((!x102x) & (!n_n4852) & (!n_n4846) & (n_n4848) & (x22116x)) + ((!x102x) & (!n_n4852) & (n_n4846) & (!n_n4848) & (!x22116x)) + ((!x102x) & (!n_n4852) & (n_n4846) & (!n_n4848) & (x22116x)) + ((!x102x) & (!n_n4852) & (n_n4846) & (n_n4848) & (!x22116x)) + ((!x102x) & (!n_n4852) & (n_n4846) & (n_n4848) & (x22116x)) + ((!x102x) & (n_n4852) & (!n_n4846) & (!n_n4848) & (!x22116x)) + ((!x102x) & (n_n4852) & (!n_n4846) & (!n_n4848) & (x22116x)) + ((!x102x) & (n_n4852) & (!n_n4846) & (n_n4848) & (!x22116x)) + ((!x102x) & (n_n4852) & (!n_n4846) & (n_n4848) & (x22116x)) + ((!x102x) & (n_n4852) & (n_n4846) & (!n_n4848) & (!x22116x)) + ((!x102x) & (n_n4852) & (n_n4846) & (!n_n4848) & (x22116x)) + ((!x102x) & (n_n4852) & (n_n4846) & (n_n4848) & (!x22116x)) + ((!x102x) & (n_n4852) & (n_n4846) & (n_n4848) & (x22116x)) + ((x102x) & (!n_n4852) & (!n_n4846) & (!n_n4848) & (!x22116x)) + ((x102x) & (!n_n4852) & (!n_n4846) & (!n_n4848) & (x22116x)) + ((x102x) & (!n_n4852) & (!n_n4846) & (n_n4848) & (!x22116x)) + ((x102x) & (!n_n4852) & (!n_n4846) & (n_n4848) & (x22116x)) + ((x102x) & (!n_n4852) & (n_n4846) & (!n_n4848) & (!x22116x)) + ((x102x) & (!n_n4852) & (n_n4846) & (!n_n4848) & (x22116x)) + ((x102x) & (!n_n4852) & (n_n4846) & (n_n4848) & (!x22116x)) + ((x102x) & (!n_n4852) & (n_n4846) & (n_n4848) & (x22116x)) + ((x102x) & (n_n4852) & (!n_n4846) & (!n_n4848) & (!x22116x)) + ((x102x) & (n_n4852) & (!n_n4846) & (!n_n4848) & (x22116x)) + ((x102x) & (n_n4852) & (!n_n4846) & (n_n4848) & (!x22116x)) + ((x102x) & (n_n4852) & (!n_n4846) & (n_n4848) & (x22116x)) + ((x102x) & (n_n4852) & (n_n4846) & (!n_n4848) & (!x22116x)) + ((x102x) & (n_n4852) & (n_n4846) & (!n_n4848) & (x22116x)) + ((x102x) & (n_n4852) & (n_n4846) & (n_n4848) & (!x22116x)) + ((x102x) & (n_n4852) & (n_n4846) & (n_n4848) & (x22116x)));
	assign n_n3327 = (((!n_n4857) & (!x40x) & (!x245x) & (!n_n4860) & (n_n1988)) + ((!n_n4857) & (!x40x) & (!x245x) & (n_n4860) & (!n_n1988)) + ((!n_n4857) & (!x40x) & (!x245x) & (n_n4860) & (n_n1988)) + ((!n_n4857) & (!x40x) & (x245x) & (!n_n4860) & (!n_n1988)) + ((!n_n4857) & (!x40x) & (x245x) & (!n_n4860) & (n_n1988)) + ((!n_n4857) & (!x40x) & (x245x) & (n_n4860) & (!n_n1988)) + ((!n_n4857) & (!x40x) & (x245x) & (n_n4860) & (n_n1988)) + ((!n_n4857) & (x40x) & (!x245x) & (!n_n4860) & (!n_n1988)) + ((!n_n4857) & (x40x) & (!x245x) & (!n_n4860) & (n_n1988)) + ((!n_n4857) & (x40x) & (!x245x) & (n_n4860) & (!n_n1988)) + ((!n_n4857) & (x40x) & (!x245x) & (n_n4860) & (n_n1988)) + ((!n_n4857) & (x40x) & (x245x) & (!n_n4860) & (!n_n1988)) + ((!n_n4857) & (x40x) & (x245x) & (!n_n4860) & (n_n1988)) + ((!n_n4857) & (x40x) & (x245x) & (n_n4860) & (!n_n1988)) + ((!n_n4857) & (x40x) & (x245x) & (n_n4860) & (n_n1988)) + ((n_n4857) & (!x40x) & (!x245x) & (!n_n4860) & (!n_n1988)) + ((n_n4857) & (!x40x) & (!x245x) & (!n_n4860) & (n_n1988)) + ((n_n4857) & (!x40x) & (!x245x) & (n_n4860) & (!n_n1988)) + ((n_n4857) & (!x40x) & (!x245x) & (n_n4860) & (n_n1988)) + ((n_n4857) & (!x40x) & (x245x) & (!n_n4860) & (!n_n1988)) + ((n_n4857) & (!x40x) & (x245x) & (!n_n4860) & (n_n1988)) + ((n_n4857) & (!x40x) & (x245x) & (n_n4860) & (!n_n1988)) + ((n_n4857) & (!x40x) & (x245x) & (n_n4860) & (n_n1988)) + ((n_n4857) & (x40x) & (!x245x) & (!n_n4860) & (!n_n1988)) + ((n_n4857) & (x40x) & (!x245x) & (!n_n4860) & (n_n1988)) + ((n_n4857) & (x40x) & (!x245x) & (n_n4860) & (!n_n1988)) + ((n_n4857) & (x40x) & (!x245x) & (n_n4860) & (n_n1988)) + ((n_n4857) & (x40x) & (x245x) & (!n_n4860) & (!n_n1988)) + ((n_n4857) & (x40x) & (x245x) & (!n_n4860) & (n_n1988)) + ((n_n4857) & (x40x) & (x245x) & (n_n4860) & (!n_n1988)) + ((n_n4857) & (x40x) & (x245x) & (n_n4860) & (n_n1988)));
	assign n_n3275 = (((!n_n3329) & (!x13820x) & (n_n3327)) + ((!n_n3329) & (x13820x) & (!n_n3327)) + ((!n_n3329) & (x13820x) & (n_n3327)) + ((n_n3329) & (!x13820x) & (!n_n3327)) + ((n_n3329) & (!x13820x) & (n_n3327)) + ((n_n3329) & (x13820x) & (!n_n3327)) + ((n_n3329) & (x13820x) & (n_n3327)));
	assign x13825x = (((!n_n4807) & (!x439x) & (!n_n4808) & (!n_n4196) & (x395x)) + ((!n_n4807) & (!x439x) & (!n_n4808) & (n_n4196) & (!x395x)) + ((!n_n4807) & (!x439x) & (!n_n4808) & (n_n4196) & (x395x)) + ((!n_n4807) & (!x439x) & (n_n4808) & (!n_n4196) & (!x395x)) + ((!n_n4807) & (!x439x) & (n_n4808) & (!n_n4196) & (x395x)) + ((!n_n4807) & (!x439x) & (n_n4808) & (n_n4196) & (!x395x)) + ((!n_n4807) & (!x439x) & (n_n4808) & (n_n4196) & (x395x)) + ((!n_n4807) & (x439x) & (!n_n4808) & (!n_n4196) & (!x395x)) + ((!n_n4807) & (x439x) & (!n_n4808) & (!n_n4196) & (x395x)) + ((!n_n4807) & (x439x) & (!n_n4808) & (n_n4196) & (!x395x)) + ((!n_n4807) & (x439x) & (!n_n4808) & (n_n4196) & (x395x)) + ((!n_n4807) & (x439x) & (n_n4808) & (!n_n4196) & (!x395x)) + ((!n_n4807) & (x439x) & (n_n4808) & (!n_n4196) & (x395x)) + ((!n_n4807) & (x439x) & (n_n4808) & (n_n4196) & (!x395x)) + ((!n_n4807) & (x439x) & (n_n4808) & (n_n4196) & (x395x)) + ((n_n4807) & (!x439x) & (!n_n4808) & (!n_n4196) & (!x395x)) + ((n_n4807) & (!x439x) & (!n_n4808) & (!n_n4196) & (x395x)) + ((n_n4807) & (!x439x) & (!n_n4808) & (n_n4196) & (!x395x)) + ((n_n4807) & (!x439x) & (!n_n4808) & (n_n4196) & (x395x)) + ((n_n4807) & (!x439x) & (n_n4808) & (!n_n4196) & (!x395x)) + ((n_n4807) & (!x439x) & (n_n4808) & (!n_n4196) & (x395x)) + ((n_n4807) & (!x439x) & (n_n4808) & (n_n4196) & (!x395x)) + ((n_n4807) & (!x439x) & (n_n4808) & (n_n4196) & (x395x)) + ((n_n4807) & (x439x) & (!n_n4808) & (!n_n4196) & (!x395x)) + ((n_n4807) & (x439x) & (!n_n4808) & (!n_n4196) & (x395x)) + ((n_n4807) & (x439x) & (!n_n4808) & (n_n4196) & (!x395x)) + ((n_n4807) & (x439x) & (!n_n4808) & (n_n4196) & (x395x)) + ((n_n4807) & (x439x) & (n_n4808) & (!n_n4196) & (!x395x)) + ((n_n4807) & (x439x) & (n_n4808) & (!n_n4196) & (x395x)) + ((n_n4807) & (x439x) & (n_n4808) & (n_n4196) & (!x395x)) + ((n_n4807) & (x439x) & (n_n4808) & (n_n4196) & (x395x)));
	assign x13827x = (((!x38x) & (!x186x) & (!n_n3332) & (!x13805x) & (x13825x)) + ((!x38x) & (!x186x) & (!n_n3332) & (x13805x) & (!x13825x)) + ((!x38x) & (!x186x) & (!n_n3332) & (x13805x) & (x13825x)) + ((!x38x) & (!x186x) & (n_n3332) & (!x13805x) & (!x13825x)) + ((!x38x) & (!x186x) & (n_n3332) & (!x13805x) & (x13825x)) + ((!x38x) & (!x186x) & (n_n3332) & (x13805x) & (!x13825x)) + ((!x38x) & (!x186x) & (n_n3332) & (x13805x) & (x13825x)) + ((!x38x) & (x186x) & (!n_n3332) & (!x13805x) & (!x13825x)) + ((!x38x) & (x186x) & (!n_n3332) & (!x13805x) & (x13825x)) + ((!x38x) & (x186x) & (!n_n3332) & (x13805x) & (!x13825x)) + ((!x38x) & (x186x) & (!n_n3332) & (x13805x) & (x13825x)) + ((!x38x) & (x186x) & (n_n3332) & (!x13805x) & (!x13825x)) + ((!x38x) & (x186x) & (n_n3332) & (!x13805x) & (x13825x)) + ((!x38x) & (x186x) & (n_n3332) & (x13805x) & (!x13825x)) + ((!x38x) & (x186x) & (n_n3332) & (x13805x) & (x13825x)) + ((x38x) & (!x186x) & (!n_n3332) & (!x13805x) & (!x13825x)) + ((x38x) & (!x186x) & (!n_n3332) & (!x13805x) & (x13825x)) + ((x38x) & (!x186x) & (!n_n3332) & (x13805x) & (!x13825x)) + ((x38x) & (!x186x) & (!n_n3332) & (x13805x) & (x13825x)) + ((x38x) & (!x186x) & (n_n3332) & (!x13805x) & (!x13825x)) + ((x38x) & (!x186x) & (n_n3332) & (!x13805x) & (x13825x)) + ((x38x) & (!x186x) & (n_n3332) & (x13805x) & (!x13825x)) + ((x38x) & (!x186x) & (n_n3332) & (x13805x) & (x13825x)) + ((x38x) & (x186x) & (!n_n3332) & (!x13805x) & (!x13825x)) + ((x38x) & (x186x) & (!n_n3332) & (!x13805x) & (x13825x)) + ((x38x) & (x186x) & (!n_n3332) & (x13805x) & (!x13825x)) + ((x38x) & (x186x) & (!n_n3332) & (x13805x) & (x13825x)) + ((x38x) & (x186x) & (n_n3332) & (!x13805x) & (!x13825x)) + ((x38x) & (x186x) & (n_n3332) & (!x13805x) & (x13825x)) + ((x38x) & (x186x) & (n_n3332) & (x13805x) & (!x13825x)) + ((x38x) & (x186x) & (n_n3332) & (x13805x) & (x13825x)));
	assign x13857x = (((!n_n4909) & (!n_n4894) & (!n_n4905) & (n_n4889)) + ((!n_n4909) & (!n_n4894) & (n_n4905) & (!n_n4889)) + ((!n_n4909) & (!n_n4894) & (n_n4905) & (n_n4889)) + ((!n_n4909) & (n_n4894) & (!n_n4905) & (!n_n4889)) + ((!n_n4909) & (n_n4894) & (!n_n4905) & (n_n4889)) + ((!n_n4909) & (n_n4894) & (n_n4905) & (!n_n4889)) + ((!n_n4909) & (n_n4894) & (n_n4905) & (n_n4889)) + ((n_n4909) & (!n_n4894) & (!n_n4905) & (!n_n4889)) + ((n_n4909) & (!n_n4894) & (!n_n4905) & (n_n4889)) + ((n_n4909) & (!n_n4894) & (n_n4905) & (!n_n4889)) + ((n_n4909) & (!n_n4894) & (n_n4905) & (n_n4889)) + ((n_n4909) & (n_n4894) & (!n_n4905) & (!n_n4889)) + ((n_n4909) & (n_n4894) & (!n_n4905) & (n_n4889)) + ((n_n4909) & (n_n4894) & (n_n4905) & (!n_n4889)) + ((n_n4909) & (n_n4894) & (n_n4905) & (n_n4889)));
	assign x22119x = (((!n_n4902) & (!n_n4907) & (!x353x) & (!x227x) & (!x49x)));
	assign n_n3274 = (((!n_n3450) & (!n_n3451) & (!n_n3326) & (!x13857x) & (!x22119x)) + ((!n_n3450) & (!n_n3451) & (!n_n3326) & (x13857x) & (!x22119x)) + ((!n_n3450) & (!n_n3451) & (!n_n3326) & (x13857x) & (x22119x)) + ((!n_n3450) & (!n_n3451) & (n_n3326) & (!x13857x) & (!x22119x)) + ((!n_n3450) & (!n_n3451) & (n_n3326) & (!x13857x) & (x22119x)) + ((!n_n3450) & (!n_n3451) & (n_n3326) & (x13857x) & (!x22119x)) + ((!n_n3450) & (!n_n3451) & (n_n3326) & (x13857x) & (x22119x)) + ((!n_n3450) & (n_n3451) & (!n_n3326) & (!x13857x) & (!x22119x)) + ((!n_n3450) & (n_n3451) & (!n_n3326) & (!x13857x) & (x22119x)) + ((!n_n3450) & (n_n3451) & (!n_n3326) & (x13857x) & (!x22119x)) + ((!n_n3450) & (n_n3451) & (!n_n3326) & (x13857x) & (x22119x)) + ((!n_n3450) & (n_n3451) & (n_n3326) & (!x13857x) & (!x22119x)) + ((!n_n3450) & (n_n3451) & (n_n3326) & (!x13857x) & (x22119x)) + ((!n_n3450) & (n_n3451) & (n_n3326) & (x13857x) & (!x22119x)) + ((!n_n3450) & (n_n3451) & (n_n3326) & (x13857x) & (x22119x)) + ((n_n3450) & (!n_n3451) & (!n_n3326) & (!x13857x) & (!x22119x)) + ((n_n3450) & (!n_n3451) & (!n_n3326) & (!x13857x) & (x22119x)) + ((n_n3450) & (!n_n3451) & (!n_n3326) & (x13857x) & (!x22119x)) + ((n_n3450) & (!n_n3451) & (!n_n3326) & (x13857x) & (x22119x)) + ((n_n3450) & (!n_n3451) & (n_n3326) & (!x13857x) & (!x22119x)) + ((n_n3450) & (!n_n3451) & (n_n3326) & (!x13857x) & (x22119x)) + ((n_n3450) & (!n_n3451) & (n_n3326) & (x13857x) & (!x22119x)) + ((n_n3450) & (!n_n3451) & (n_n3326) & (x13857x) & (x22119x)) + ((n_n3450) & (n_n3451) & (!n_n3326) & (!x13857x) & (!x22119x)) + ((n_n3450) & (n_n3451) & (!n_n3326) & (!x13857x) & (x22119x)) + ((n_n3450) & (n_n3451) & (!n_n3326) & (x13857x) & (!x22119x)) + ((n_n3450) & (n_n3451) & (!n_n3326) & (x13857x) & (x22119x)) + ((n_n3450) & (n_n3451) & (n_n3326) & (!x13857x) & (!x22119x)) + ((n_n3450) & (n_n3451) & (n_n3326) & (!x13857x) & (x22119x)) + ((n_n3450) & (n_n3451) & (n_n3326) & (x13857x) & (!x22119x)) + ((n_n3450) & (n_n3451) & (n_n3326) & (x13857x) & (x22119x)));
	assign x22118x = (((!x17x) & (!n_n4927) & (!x502x) & (!n_n4934) & (!n_n4933)) + ((!x17x) & (!n_n4927) & (x502x) & (!n_n4934) & (!n_n4933)) + ((x17x) & (!n_n4927) & (!x502x) & (!n_n4934) & (!n_n4933)));
	assign n_n3322 = (((!n_n4926) & (!n_n4925) & (!x31x) & (!n_n4931) & (!x22118x)) + ((!n_n4926) & (!n_n4925) & (!x31x) & (n_n4931) & (!x22118x)) + ((!n_n4926) & (!n_n4925) & (!x31x) & (n_n4931) & (x22118x)) + ((!n_n4926) & (!n_n4925) & (x31x) & (!n_n4931) & (!x22118x)) + ((!n_n4926) & (!n_n4925) & (x31x) & (!n_n4931) & (x22118x)) + ((!n_n4926) & (!n_n4925) & (x31x) & (n_n4931) & (!x22118x)) + ((!n_n4926) & (!n_n4925) & (x31x) & (n_n4931) & (x22118x)) + ((!n_n4926) & (n_n4925) & (!x31x) & (!n_n4931) & (!x22118x)) + ((!n_n4926) & (n_n4925) & (!x31x) & (!n_n4931) & (x22118x)) + ((!n_n4926) & (n_n4925) & (!x31x) & (n_n4931) & (!x22118x)) + ((!n_n4926) & (n_n4925) & (!x31x) & (n_n4931) & (x22118x)) + ((!n_n4926) & (n_n4925) & (x31x) & (!n_n4931) & (!x22118x)) + ((!n_n4926) & (n_n4925) & (x31x) & (!n_n4931) & (x22118x)) + ((!n_n4926) & (n_n4925) & (x31x) & (n_n4931) & (!x22118x)) + ((!n_n4926) & (n_n4925) & (x31x) & (n_n4931) & (x22118x)) + ((n_n4926) & (!n_n4925) & (!x31x) & (!n_n4931) & (!x22118x)) + ((n_n4926) & (!n_n4925) & (!x31x) & (!n_n4931) & (x22118x)) + ((n_n4926) & (!n_n4925) & (!x31x) & (n_n4931) & (!x22118x)) + ((n_n4926) & (!n_n4925) & (!x31x) & (n_n4931) & (x22118x)) + ((n_n4926) & (!n_n4925) & (x31x) & (!n_n4931) & (!x22118x)) + ((n_n4926) & (!n_n4925) & (x31x) & (!n_n4931) & (x22118x)) + ((n_n4926) & (!n_n4925) & (x31x) & (n_n4931) & (!x22118x)) + ((n_n4926) & (!n_n4925) & (x31x) & (n_n4931) & (x22118x)) + ((n_n4926) & (n_n4925) & (!x31x) & (!n_n4931) & (!x22118x)) + ((n_n4926) & (n_n4925) & (!x31x) & (!n_n4931) & (x22118x)) + ((n_n4926) & (n_n4925) & (!x31x) & (n_n4931) & (!x22118x)) + ((n_n4926) & (n_n4925) & (!x31x) & (n_n4931) & (x22118x)) + ((n_n4926) & (n_n4925) & (x31x) & (!n_n4931) & (!x22118x)) + ((n_n4926) & (n_n4925) & (x31x) & (!n_n4931) & (x22118x)) + ((n_n4926) & (n_n4925) & (x31x) & (n_n4931) & (!x22118x)) + ((n_n4926) & (n_n4925) & (x31x) & (n_n4931) & (x22118x)));
	assign n_n4910 = (((i_9_) & (n_n482) & (n_n528) & (n_n260)));
	assign x13868x = (((!i_9_) & (n_n482) & (n_n528) & (n_n260) & (!n_n522)) + ((!i_9_) & (n_n482) & (n_n528) & (n_n260) & (n_n522)) + ((i_9_) & (n_n482) & (!n_n528) & (n_n260) & (n_n522)) + ((i_9_) & (n_n482) & (n_n528) & (n_n260) & (n_n522)));
	assign x138x = (((!n_n4918) & (!n_n4919) & (!n_n4917) & (!n_n4910) & (x13868x)) + ((!n_n4918) & (!n_n4919) & (!n_n4917) & (n_n4910) & (!x13868x)) + ((!n_n4918) & (!n_n4919) & (!n_n4917) & (n_n4910) & (x13868x)) + ((!n_n4918) & (!n_n4919) & (n_n4917) & (!n_n4910) & (!x13868x)) + ((!n_n4918) & (!n_n4919) & (n_n4917) & (!n_n4910) & (x13868x)) + ((!n_n4918) & (!n_n4919) & (n_n4917) & (n_n4910) & (!x13868x)) + ((!n_n4918) & (!n_n4919) & (n_n4917) & (n_n4910) & (x13868x)) + ((!n_n4918) & (n_n4919) & (!n_n4917) & (!n_n4910) & (!x13868x)) + ((!n_n4918) & (n_n4919) & (!n_n4917) & (!n_n4910) & (x13868x)) + ((!n_n4918) & (n_n4919) & (!n_n4917) & (n_n4910) & (!x13868x)) + ((!n_n4918) & (n_n4919) & (!n_n4917) & (n_n4910) & (x13868x)) + ((!n_n4918) & (n_n4919) & (n_n4917) & (!n_n4910) & (!x13868x)) + ((!n_n4918) & (n_n4919) & (n_n4917) & (!n_n4910) & (x13868x)) + ((!n_n4918) & (n_n4919) & (n_n4917) & (n_n4910) & (!x13868x)) + ((!n_n4918) & (n_n4919) & (n_n4917) & (n_n4910) & (x13868x)) + ((n_n4918) & (!n_n4919) & (!n_n4917) & (!n_n4910) & (!x13868x)) + ((n_n4918) & (!n_n4919) & (!n_n4917) & (!n_n4910) & (x13868x)) + ((n_n4918) & (!n_n4919) & (!n_n4917) & (n_n4910) & (!x13868x)) + ((n_n4918) & (!n_n4919) & (!n_n4917) & (n_n4910) & (x13868x)) + ((n_n4918) & (!n_n4919) & (n_n4917) & (!n_n4910) & (!x13868x)) + ((n_n4918) & (!n_n4919) & (n_n4917) & (!n_n4910) & (x13868x)) + ((n_n4918) & (!n_n4919) & (n_n4917) & (n_n4910) & (!x13868x)) + ((n_n4918) & (!n_n4919) & (n_n4917) & (n_n4910) & (x13868x)) + ((n_n4918) & (n_n4919) & (!n_n4917) & (!n_n4910) & (!x13868x)) + ((n_n4918) & (n_n4919) & (!n_n4917) & (!n_n4910) & (x13868x)) + ((n_n4918) & (n_n4919) & (!n_n4917) & (n_n4910) & (!x13868x)) + ((n_n4918) & (n_n4919) & (!n_n4917) & (n_n4910) & (x13868x)) + ((n_n4918) & (n_n4919) & (n_n4917) & (!n_n4910) & (!x13868x)) + ((n_n4918) & (n_n4919) & (n_n4917) & (!n_n4910) & (x13868x)) + ((n_n4918) & (n_n4919) & (n_n4917) & (n_n4910) & (!x13868x)) + ((n_n4918) & (n_n4919) & (n_n4917) & (n_n4910) & (x13868x)));
	assign x331x = (((!i_9_) & (!n_n532) & (n_n534) & (n_n260) & (n_n464)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n260) & (n_n464)) + ((i_9_) & (n_n532) & (!n_n534) & (n_n260) & (n_n464)) + ((i_9_) & (n_n532) & (n_n534) & (n_n260) & (n_n464)));
	assign x13875x = (((!n_n4923) & (!n_n4924) & (!n_n4937) & (!n_n4938) & (x58x)) + ((!n_n4923) & (!n_n4924) & (!n_n4937) & (n_n4938) & (!x58x)) + ((!n_n4923) & (!n_n4924) & (!n_n4937) & (n_n4938) & (x58x)) + ((!n_n4923) & (!n_n4924) & (n_n4937) & (!n_n4938) & (!x58x)) + ((!n_n4923) & (!n_n4924) & (n_n4937) & (!n_n4938) & (x58x)) + ((!n_n4923) & (!n_n4924) & (n_n4937) & (n_n4938) & (!x58x)) + ((!n_n4923) & (!n_n4924) & (n_n4937) & (n_n4938) & (x58x)) + ((!n_n4923) & (n_n4924) & (!n_n4937) & (!n_n4938) & (!x58x)) + ((!n_n4923) & (n_n4924) & (!n_n4937) & (!n_n4938) & (x58x)) + ((!n_n4923) & (n_n4924) & (!n_n4937) & (n_n4938) & (!x58x)) + ((!n_n4923) & (n_n4924) & (!n_n4937) & (n_n4938) & (x58x)) + ((!n_n4923) & (n_n4924) & (n_n4937) & (!n_n4938) & (!x58x)) + ((!n_n4923) & (n_n4924) & (n_n4937) & (!n_n4938) & (x58x)) + ((!n_n4923) & (n_n4924) & (n_n4937) & (n_n4938) & (!x58x)) + ((!n_n4923) & (n_n4924) & (n_n4937) & (n_n4938) & (x58x)) + ((n_n4923) & (!n_n4924) & (!n_n4937) & (!n_n4938) & (!x58x)) + ((n_n4923) & (!n_n4924) & (!n_n4937) & (!n_n4938) & (x58x)) + ((n_n4923) & (!n_n4924) & (!n_n4937) & (n_n4938) & (!x58x)) + ((n_n4923) & (!n_n4924) & (!n_n4937) & (n_n4938) & (x58x)) + ((n_n4923) & (!n_n4924) & (n_n4937) & (!n_n4938) & (!x58x)) + ((n_n4923) & (!n_n4924) & (n_n4937) & (!n_n4938) & (x58x)) + ((n_n4923) & (!n_n4924) & (n_n4937) & (n_n4938) & (!x58x)) + ((n_n4923) & (!n_n4924) & (n_n4937) & (n_n4938) & (x58x)) + ((n_n4923) & (n_n4924) & (!n_n4937) & (!n_n4938) & (!x58x)) + ((n_n4923) & (n_n4924) & (!n_n4937) & (!n_n4938) & (x58x)) + ((n_n4923) & (n_n4924) & (!n_n4937) & (n_n4938) & (!x58x)) + ((n_n4923) & (n_n4924) & (!n_n4937) & (n_n4938) & (x58x)) + ((n_n4923) & (n_n4924) & (n_n4937) & (!n_n4938) & (!x58x)) + ((n_n4923) & (n_n4924) & (n_n4937) & (!n_n4938) & (x58x)) + ((n_n4923) & (n_n4924) & (n_n4937) & (n_n4938) & (!x58x)) + ((n_n4923) & (n_n4924) & (n_n4937) & (n_n4938) & (x58x)));
	assign x13876x = (((!n_n4921) & (!n_n4935) & (!n_n2710) & (x138x)) + ((!n_n4921) & (!n_n4935) & (n_n2710) & (!x138x)) + ((!n_n4921) & (!n_n4935) & (n_n2710) & (x138x)) + ((!n_n4921) & (n_n4935) & (!n_n2710) & (!x138x)) + ((!n_n4921) & (n_n4935) & (!n_n2710) & (x138x)) + ((!n_n4921) & (n_n4935) & (n_n2710) & (!x138x)) + ((!n_n4921) & (n_n4935) & (n_n2710) & (x138x)) + ((n_n4921) & (!n_n4935) & (!n_n2710) & (!x138x)) + ((n_n4921) & (!n_n4935) & (!n_n2710) & (x138x)) + ((n_n4921) & (!n_n4935) & (n_n2710) & (!x138x)) + ((n_n4921) & (!n_n4935) & (n_n2710) & (x138x)) + ((n_n4921) & (n_n4935) & (!n_n2710) & (!x138x)) + ((n_n4921) & (n_n4935) & (!n_n2710) & (x138x)) + ((n_n4921) & (n_n4935) & (n_n2710) & (!x138x)) + ((n_n4921) & (n_n4935) & (n_n2710) & (x138x)));
	assign n_n3124 = (((!i_9_) & (n_n524) & (n_n325) & (n_n535) & (!n_n522)) + ((!i_9_) & (n_n524) & (n_n325) & (n_n535) & (n_n522)) + ((i_9_) & (!n_n524) & (n_n325) & (n_n535) & (n_n522)) + ((i_9_) & (n_n524) & (n_n325) & (n_n535) & (!n_n522)) + ((i_9_) & (n_n524) & (n_n325) & (n_n535) & (n_n522)));
	assign x13910x = (((!n_n4711) & (!n_n4719) & (!x457x) & (!n_n3124) & (n_n2378)) + ((!n_n4711) & (!n_n4719) & (!x457x) & (n_n3124) & (!n_n2378)) + ((!n_n4711) & (!n_n4719) & (!x457x) & (n_n3124) & (n_n2378)) + ((!n_n4711) & (!n_n4719) & (x457x) & (!n_n3124) & (!n_n2378)) + ((!n_n4711) & (!n_n4719) & (x457x) & (!n_n3124) & (n_n2378)) + ((!n_n4711) & (!n_n4719) & (x457x) & (n_n3124) & (!n_n2378)) + ((!n_n4711) & (!n_n4719) & (x457x) & (n_n3124) & (n_n2378)) + ((!n_n4711) & (n_n4719) & (!x457x) & (!n_n3124) & (!n_n2378)) + ((!n_n4711) & (n_n4719) & (!x457x) & (!n_n3124) & (n_n2378)) + ((!n_n4711) & (n_n4719) & (!x457x) & (n_n3124) & (!n_n2378)) + ((!n_n4711) & (n_n4719) & (!x457x) & (n_n3124) & (n_n2378)) + ((!n_n4711) & (n_n4719) & (x457x) & (!n_n3124) & (!n_n2378)) + ((!n_n4711) & (n_n4719) & (x457x) & (!n_n3124) & (n_n2378)) + ((!n_n4711) & (n_n4719) & (x457x) & (n_n3124) & (!n_n2378)) + ((!n_n4711) & (n_n4719) & (x457x) & (n_n3124) & (n_n2378)) + ((n_n4711) & (!n_n4719) & (!x457x) & (!n_n3124) & (!n_n2378)) + ((n_n4711) & (!n_n4719) & (!x457x) & (!n_n3124) & (n_n2378)) + ((n_n4711) & (!n_n4719) & (!x457x) & (n_n3124) & (!n_n2378)) + ((n_n4711) & (!n_n4719) & (!x457x) & (n_n3124) & (n_n2378)) + ((n_n4711) & (!n_n4719) & (x457x) & (!n_n3124) & (!n_n2378)) + ((n_n4711) & (!n_n4719) & (x457x) & (!n_n3124) & (n_n2378)) + ((n_n4711) & (!n_n4719) & (x457x) & (n_n3124) & (!n_n2378)) + ((n_n4711) & (!n_n4719) & (x457x) & (n_n3124) & (n_n2378)) + ((n_n4711) & (n_n4719) & (!x457x) & (!n_n3124) & (!n_n2378)) + ((n_n4711) & (n_n4719) & (!x457x) & (!n_n3124) & (n_n2378)) + ((n_n4711) & (n_n4719) & (!x457x) & (n_n3124) & (!n_n2378)) + ((n_n4711) & (n_n4719) & (!x457x) & (n_n3124) & (n_n2378)) + ((n_n4711) & (n_n4719) & (x457x) & (!n_n3124) & (!n_n2378)) + ((n_n4711) & (n_n4719) & (x457x) & (!n_n3124) & (n_n2378)) + ((n_n4711) & (n_n4719) & (x457x) & (n_n3124) & (!n_n2378)) + ((n_n4711) & (n_n4719) & (x457x) & (n_n3124) & (n_n2378)));
	assign x442x = (((!i_9_) & (n_n325) & (n_n535) & (n_n530)) + ((i_9_) & (n_n325) & (n_n535) & (n_n530)));
	assign x13903x = (((!n_n4688) & (!n_n4691) & (!n_n4686) & (!n_n4694) & (n_n4693)) + ((!n_n4688) & (!n_n4691) & (!n_n4686) & (n_n4694) & (!n_n4693)) + ((!n_n4688) & (!n_n4691) & (!n_n4686) & (n_n4694) & (n_n4693)) + ((!n_n4688) & (!n_n4691) & (n_n4686) & (!n_n4694) & (!n_n4693)) + ((!n_n4688) & (!n_n4691) & (n_n4686) & (!n_n4694) & (n_n4693)) + ((!n_n4688) & (!n_n4691) & (n_n4686) & (n_n4694) & (!n_n4693)) + ((!n_n4688) & (!n_n4691) & (n_n4686) & (n_n4694) & (n_n4693)) + ((!n_n4688) & (n_n4691) & (!n_n4686) & (!n_n4694) & (!n_n4693)) + ((!n_n4688) & (n_n4691) & (!n_n4686) & (!n_n4694) & (n_n4693)) + ((!n_n4688) & (n_n4691) & (!n_n4686) & (n_n4694) & (!n_n4693)) + ((!n_n4688) & (n_n4691) & (!n_n4686) & (n_n4694) & (n_n4693)) + ((!n_n4688) & (n_n4691) & (n_n4686) & (!n_n4694) & (!n_n4693)) + ((!n_n4688) & (n_n4691) & (n_n4686) & (!n_n4694) & (n_n4693)) + ((!n_n4688) & (n_n4691) & (n_n4686) & (n_n4694) & (!n_n4693)) + ((!n_n4688) & (n_n4691) & (n_n4686) & (n_n4694) & (n_n4693)) + ((n_n4688) & (!n_n4691) & (!n_n4686) & (!n_n4694) & (!n_n4693)) + ((n_n4688) & (!n_n4691) & (!n_n4686) & (!n_n4694) & (n_n4693)) + ((n_n4688) & (!n_n4691) & (!n_n4686) & (n_n4694) & (!n_n4693)) + ((n_n4688) & (!n_n4691) & (!n_n4686) & (n_n4694) & (n_n4693)) + ((n_n4688) & (!n_n4691) & (n_n4686) & (!n_n4694) & (!n_n4693)) + ((n_n4688) & (!n_n4691) & (n_n4686) & (!n_n4694) & (n_n4693)) + ((n_n4688) & (!n_n4691) & (n_n4686) & (n_n4694) & (!n_n4693)) + ((n_n4688) & (!n_n4691) & (n_n4686) & (n_n4694) & (n_n4693)) + ((n_n4688) & (n_n4691) & (!n_n4686) & (!n_n4694) & (!n_n4693)) + ((n_n4688) & (n_n4691) & (!n_n4686) & (!n_n4694) & (n_n4693)) + ((n_n4688) & (n_n4691) & (!n_n4686) & (n_n4694) & (!n_n4693)) + ((n_n4688) & (n_n4691) & (!n_n4686) & (n_n4694) & (n_n4693)) + ((n_n4688) & (n_n4691) & (n_n4686) & (!n_n4694) & (!n_n4693)) + ((n_n4688) & (n_n4691) & (n_n4686) & (!n_n4694) & (n_n4693)) + ((n_n4688) & (n_n4691) & (n_n4686) & (n_n4694) & (!n_n4693)) + ((n_n4688) & (n_n4691) & (n_n4686) & (n_n4694) & (n_n4693)));
	assign x13899x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n390) & (n_n464)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n390) & (n_n464)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n390) & (n_n464)) + ((i_9_) & (n_n524) & (n_n526) & (n_n390) & (n_n464)));
	assign x13909x = (((!x241x) & (!n_n4712) & (!n_n4714) & (!n_n4716) & (x30x)) + ((!x241x) & (!n_n4712) & (!n_n4714) & (n_n4716) & (!x30x)) + ((!x241x) & (!n_n4712) & (!n_n4714) & (n_n4716) & (x30x)) + ((!x241x) & (!n_n4712) & (n_n4714) & (!n_n4716) & (!x30x)) + ((!x241x) & (!n_n4712) & (n_n4714) & (!n_n4716) & (x30x)) + ((!x241x) & (!n_n4712) & (n_n4714) & (n_n4716) & (!x30x)) + ((!x241x) & (!n_n4712) & (n_n4714) & (n_n4716) & (x30x)) + ((!x241x) & (n_n4712) & (!n_n4714) & (!n_n4716) & (!x30x)) + ((!x241x) & (n_n4712) & (!n_n4714) & (!n_n4716) & (x30x)) + ((!x241x) & (n_n4712) & (!n_n4714) & (n_n4716) & (!x30x)) + ((!x241x) & (n_n4712) & (!n_n4714) & (n_n4716) & (x30x)) + ((!x241x) & (n_n4712) & (n_n4714) & (!n_n4716) & (!x30x)) + ((!x241x) & (n_n4712) & (n_n4714) & (!n_n4716) & (x30x)) + ((!x241x) & (n_n4712) & (n_n4714) & (n_n4716) & (!x30x)) + ((!x241x) & (n_n4712) & (n_n4714) & (n_n4716) & (x30x)) + ((x241x) & (!n_n4712) & (!n_n4714) & (!n_n4716) & (!x30x)) + ((x241x) & (!n_n4712) & (!n_n4714) & (!n_n4716) & (x30x)) + ((x241x) & (!n_n4712) & (!n_n4714) & (n_n4716) & (!x30x)) + ((x241x) & (!n_n4712) & (!n_n4714) & (n_n4716) & (x30x)) + ((x241x) & (!n_n4712) & (n_n4714) & (!n_n4716) & (!x30x)) + ((x241x) & (!n_n4712) & (n_n4714) & (!n_n4716) & (x30x)) + ((x241x) & (!n_n4712) & (n_n4714) & (n_n4716) & (!x30x)) + ((x241x) & (!n_n4712) & (n_n4714) & (n_n4716) & (x30x)) + ((x241x) & (n_n4712) & (!n_n4714) & (!n_n4716) & (!x30x)) + ((x241x) & (n_n4712) & (!n_n4714) & (!n_n4716) & (x30x)) + ((x241x) & (n_n4712) & (!n_n4714) & (n_n4716) & (!x30x)) + ((x241x) & (n_n4712) & (!n_n4714) & (n_n4716) & (x30x)) + ((x241x) & (n_n4712) & (n_n4714) & (!n_n4716) & (!x30x)) + ((x241x) & (n_n4712) & (n_n4714) & (!n_n4716) & (x30x)) + ((x241x) & (n_n4712) & (n_n4714) & (n_n4716) & (!x30x)) + ((x241x) & (n_n4712) & (n_n4714) & (n_n4716) & (x30x)));
	assign n_n3279 = (((!x13910x) & (!x442x) & (!x13903x) & (!x13899x) & (x13909x)) + ((!x13910x) & (!x442x) & (!x13903x) & (x13899x) & (!x13909x)) + ((!x13910x) & (!x442x) & (!x13903x) & (x13899x) & (x13909x)) + ((!x13910x) & (!x442x) & (x13903x) & (!x13899x) & (!x13909x)) + ((!x13910x) & (!x442x) & (x13903x) & (!x13899x) & (x13909x)) + ((!x13910x) & (!x442x) & (x13903x) & (x13899x) & (!x13909x)) + ((!x13910x) & (!x442x) & (x13903x) & (x13899x) & (x13909x)) + ((!x13910x) & (x442x) & (!x13903x) & (!x13899x) & (!x13909x)) + ((!x13910x) & (x442x) & (!x13903x) & (!x13899x) & (x13909x)) + ((!x13910x) & (x442x) & (!x13903x) & (x13899x) & (!x13909x)) + ((!x13910x) & (x442x) & (!x13903x) & (x13899x) & (x13909x)) + ((!x13910x) & (x442x) & (x13903x) & (!x13899x) & (!x13909x)) + ((!x13910x) & (x442x) & (x13903x) & (!x13899x) & (x13909x)) + ((!x13910x) & (x442x) & (x13903x) & (x13899x) & (!x13909x)) + ((!x13910x) & (x442x) & (x13903x) & (x13899x) & (x13909x)) + ((x13910x) & (!x442x) & (!x13903x) & (!x13899x) & (!x13909x)) + ((x13910x) & (!x442x) & (!x13903x) & (!x13899x) & (x13909x)) + ((x13910x) & (!x442x) & (!x13903x) & (x13899x) & (!x13909x)) + ((x13910x) & (!x442x) & (!x13903x) & (x13899x) & (x13909x)) + ((x13910x) & (!x442x) & (x13903x) & (!x13899x) & (!x13909x)) + ((x13910x) & (!x442x) & (x13903x) & (!x13899x) & (x13909x)) + ((x13910x) & (!x442x) & (x13903x) & (x13899x) & (!x13909x)) + ((x13910x) & (!x442x) & (x13903x) & (x13899x) & (x13909x)) + ((x13910x) & (x442x) & (!x13903x) & (!x13899x) & (!x13909x)) + ((x13910x) & (x442x) & (!x13903x) & (!x13899x) & (x13909x)) + ((x13910x) & (x442x) & (!x13903x) & (x13899x) & (!x13909x)) + ((x13910x) & (x442x) & (!x13903x) & (x13899x) & (x13909x)) + ((x13910x) & (x442x) & (x13903x) & (!x13899x) & (!x13909x)) + ((x13910x) & (x442x) & (x13903x) & (!x13899x) & (x13909x)) + ((x13910x) & (x442x) & (x13903x) & (x13899x) & (!x13909x)) + ((x13910x) & (x442x) & (x13903x) & (x13899x) & (x13909x)));
	assign x456x = (((!x21x) & (!x483x) & (!x20x) & (!x373x) & (x94x)) + ((!x21x) & (!x483x) & (!x20x) & (x373x) & (!x94x)) + ((!x21x) & (!x483x) & (!x20x) & (x373x) & (x94x)) + ((!x21x) & (!x483x) & (x20x) & (!x373x) & (x94x)) + ((!x21x) & (!x483x) & (x20x) & (x373x) & (!x94x)) + ((!x21x) & (!x483x) & (x20x) & (x373x) & (x94x)) + ((!x21x) & (x483x) & (!x20x) & (!x373x) & (x94x)) + ((!x21x) & (x483x) & (!x20x) & (x373x) & (!x94x)) + ((!x21x) & (x483x) & (!x20x) & (x373x) & (x94x)) + ((!x21x) & (x483x) & (x20x) & (!x373x) & (!x94x)) + ((!x21x) & (x483x) & (x20x) & (!x373x) & (x94x)) + ((!x21x) & (x483x) & (x20x) & (x373x) & (!x94x)) + ((!x21x) & (x483x) & (x20x) & (x373x) & (x94x)) + ((x21x) & (!x483x) & (!x20x) & (!x373x) & (x94x)) + ((x21x) & (!x483x) & (!x20x) & (x373x) & (!x94x)) + ((x21x) & (!x483x) & (!x20x) & (x373x) & (x94x)) + ((x21x) & (!x483x) & (x20x) & (!x373x) & (x94x)) + ((x21x) & (!x483x) & (x20x) & (x373x) & (!x94x)) + ((x21x) & (!x483x) & (x20x) & (x373x) & (x94x)) + ((x21x) & (x483x) & (!x20x) & (!x373x) & (!x94x)) + ((x21x) & (x483x) & (!x20x) & (!x373x) & (x94x)) + ((x21x) & (x483x) & (!x20x) & (x373x) & (!x94x)) + ((x21x) & (x483x) & (!x20x) & (x373x) & (x94x)) + ((x21x) & (x483x) & (x20x) & (!x373x) & (!x94x)) + ((x21x) & (x483x) & (x20x) & (!x373x) & (x94x)) + ((x21x) & (x483x) & (x20x) & (x373x) & (!x94x)) + ((x21x) & (x483x) & (x20x) & (x373x) & (x94x)));
	assign x13916x = (((!x25x) & (!x483x) & (!x101x) & (!x244x) & (x73x)) + ((!x25x) & (!x483x) & (!x101x) & (x244x) & (!x73x)) + ((!x25x) & (!x483x) & (!x101x) & (x244x) & (x73x)) + ((!x25x) & (!x483x) & (x101x) & (!x244x) & (!x73x)) + ((!x25x) & (!x483x) & (x101x) & (!x244x) & (x73x)) + ((!x25x) & (!x483x) & (x101x) & (x244x) & (!x73x)) + ((!x25x) & (!x483x) & (x101x) & (x244x) & (x73x)) + ((!x25x) & (x483x) & (!x101x) & (!x244x) & (x73x)) + ((!x25x) & (x483x) & (!x101x) & (x244x) & (!x73x)) + ((!x25x) & (x483x) & (!x101x) & (x244x) & (x73x)) + ((!x25x) & (x483x) & (x101x) & (!x244x) & (!x73x)) + ((!x25x) & (x483x) & (x101x) & (!x244x) & (x73x)) + ((!x25x) & (x483x) & (x101x) & (x244x) & (!x73x)) + ((!x25x) & (x483x) & (x101x) & (x244x) & (x73x)) + ((x25x) & (!x483x) & (!x101x) & (!x244x) & (x73x)) + ((x25x) & (!x483x) & (!x101x) & (x244x) & (!x73x)) + ((x25x) & (!x483x) & (!x101x) & (x244x) & (x73x)) + ((x25x) & (!x483x) & (x101x) & (!x244x) & (!x73x)) + ((x25x) & (!x483x) & (x101x) & (!x244x) & (x73x)) + ((x25x) & (!x483x) & (x101x) & (x244x) & (!x73x)) + ((x25x) & (!x483x) & (x101x) & (x244x) & (x73x)) + ((x25x) & (x483x) & (!x101x) & (!x244x) & (!x73x)) + ((x25x) & (x483x) & (!x101x) & (!x244x) & (x73x)) + ((x25x) & (x483x) & (!x101x) & (x244x) & (!x73x)) + ((x25x) & (x483x) & (!x101x) & (x244x) & (x73x)) + ((x25x) & (x483x) & (x101x) & (!x244x) & (!x73x)) + ((x25x) & (x483x) & (x101x) & (!x244x) & (x73x)) + ((x25x) & (x483x) & (x101x) & (x244x) & (!x73x)) + ((x25x) & (x483x) & (x101x) & (x244x) & (x73x)));
	assign x13917x = (((!n_n4727) & (!x95x) & (!n_n4733) & (!n_n4736) & (x456x)) + ((!n_n4727) & (!x95x) & (!n_n4733) & (n_n4736) & (!x456x)) + ((!n_n4727) & (!x95x) & (!n_n4733) & (n_n4736) & (x456x)) + ((!n_n4727) & (!x95x) & (n_n4733) & (!n_n4736) & (!x456x)) + ((!n_n4727) & (!x95x) & (n_n4733) & (!n_n4736) & (x456x)) + ((!n_n4727) & (!x95x) & (n_n4733) & (n_n4736) & (!x456x)) + ((!n_n4727) & (!x95x) & (n_n4733) & (n_n4736) & (x456x)) + ((!n_n4727) & (x95x) & (!n_n4733) & (!n_n4736) & (!x456x)) + ((!n_n4727) & (x95x) & (!n_n4733) & (!n_n4736) & (x456x)) + ((!n_n4727) & (x95x) & (!n_n4733) & (n_n4736) & (!x456x)) + ((!n_n4727) & (x95x) & (!n_n4733) & (n_n4736) & (x456x)) + ((!n_n4727) & (x95x) & (n_n4733) & (!n_n4736) & (!x456x)) + ((!n_n4727) & (x95x) & (n_n4733) & (!n_n4736) & (x456x)) + ((!n_n4727) & (x95x) & (n_n4733) & (n_n4736) & (!x456x)) + ((!n_n4727) & (x95x) & (n_n4733) & (n_n4736) & (x456x)) + ((n_n4727) & (!x95x) & (!n_n4733) & (!n_n4736) & (!x456x)) + ((n_n4727) & (!x95x) & (!n_n4733) & (!n_n4736) & (x456x)) + ((n_n4727) & (!x95x) & (!n_n4733) & (n_n4736) & (!x456x)) + ((n_n4727) & (!x95x) & (!n_n4733) & (n_n4736) & (x456x)) + ((n_n4727) & (!x95x) & (n_n4733) & (!n_n4736) & (!x456x)) + ((n_n4727) & (!x95x) & (n_n4733) & (!n_n4736) & (x456x)) + ((n_n4727) & (!x95x) & (n_n4733) & (n_n4736) & (!x456x)) + ((n_n4727) & (!x95x) & (n_n4733) & (n_n4736) & (x456x)) + ((n_n4727) & (x95x) & (!n_n4733) & (!n_n4736) & (!x456x)) + ((n_n4727) & (x95x) & (!n_n4733) & (!n_n4736) & (x456x)) + ((n_n4727) & (x95x) & (!n_n4733) & (n_n4736) & (!x456x)) + ((n_n4727) & (x95x) & (!n_n4733) & (n_n4736) & (x456x)) + ((n_n4727) & (x95x) & (n_n4733) & (!n_n4736) & (!x456x)) + ((n_n4727) & (x95x) & (n_n4733) & (!n_n4736) & (x456x)) + ((n_n4727) & (x95x) & (n_n4733) & (n_n4736) & (!x456x)) + ((n_n4727) & (x95x) & (n_n4733) & (n_n4736) & (x456x)));
	assign n_n4723 = (((!i_9_) & (n_n524) & (n_n518) & (n_n325)));
	assign x357x = (((!i_9_) & (!n_n390) & (!n_n534) & (!n_n491) & (n_n4630)) + ((!i_9_) & (!n_n390) & (!n_n534) & (n_n491) & (n_n4630)) + ((!i_9_) & (!n_n390) & (n_n534) & (!n_n491) & (n_n4630)) + ((!i_9_) & (!n_n390) & (n_n534) & (n_n491) & (n_n4630)) + ((!i_9_) & (n_n390) & (!n_n534) & (!n_n491) & (n_n4630)) + ((!i_9_) & (n_n390) & (!n_n534) & (n_n491) & (n_n4630)) + ((!i_9_) & (n_n390) & (n_n534) & (!n_n491) & (n_n4630)) + ((!i_9_) & (n_n390) & (n_n534) & (n_n491) & (!n_n4630)) + ((!i_9_) & (n_n390) & (n_n534) & (n_n491) & (n_n4630)) + ((i_9_) & (!n_n390) & (!n_n534) & (!n_n491) & (n_n4630)) + ((i_9_) & (!n_n390) & (!n_n534) & (n_n491) & (n_n4630)) + ((i_9_) & (!n_n390) & (n_n534) & (!n_n491) & (n_n4630)) + ((i_9_) & (!n_n390) & (n_n534) & (n_n491) & (n_n4630)) + ((i_9_) & (n_n390) & (!n_n534) & (!n_n491) & (n_n4630)) + ((i_9_) & (n_n390) & (!n_n534) & (n_n491) & (n_n4630)) + ((i_9_) & (n_n390) & (n_n534) & (!n_n491) & (n_n4630)) + ((i_9_) & (n_n390) & (n_n534) & (n_n491) & (n_n4630)));
	assign n_n3125 = (((!i_9_) & (!n_n532) & (n_n534) & (n_n325) & (n_n535)) + ((!i_9_) & (n_n532) & (!n_n534) & (n_n325) & (n_n535)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n325) & (n_n535)) + ((i_9_) & (!n_n532) & (n_n534) & (n_n325) & (n_n535)) + ((i_9_) & (n_n532) & (n_n534) & (n_n325) & (n_n535)));
	assign n_n4520 = (((i_9_) & (n_n482) & (n_n455) & (n_n534)));
	assign n_n5008 = (((i_9_) & (n_n526) & (n_n195) & (n_n500)));
	assign x22081x = (((!n_n4494) & (!n_n4495) & (!n_n4497) & (!n_n4500)));
	assign x13454x = (((!i_9_) & (n_n526) & (n_n390) & (n_n491)) + ((i_9_) & (n_n526) & (n_n390) & (n_n491)));
	assign x15754x = (((!i_9_) & (!n_n526) & (n_n482) & (n_n534) & (n_n325)) + ((!i_9_) & (n_n526) & (n_n482) & (!n_n534) & (n_n325)) + ((!i_9_) & (n_n526) & (n_n482) & (n_n534) & (n_n325)));
	assign x15757x = (((!n_n4782) & (!n_n4781) & (!n_n4775) & (x15754x)) + ((!n_n4782) & (!n_n4781) & (n_n4775) & (!x15754x)) + ((!n_n4782) & (!n_n4781) & (n_n4775) & (x15754x)) + ((!n_n4782) & (n_n4781) & (!n_n4775) & (!x15754x)) + ((!n_n4782) & (n_n4781) & (!n_n4775) & (x15754x)) + ((!n_n4782) & (n_n4781) & (n_n4775) & (!x15754x)) + ((!n_n4782) & (n_n4781) & (n_n4775) & (x15754x)) + ((n_n4782) & (!n_n4781) & (!n_n4775) & (!x15754x)) + ((n_n4782) & (!n_n4781) & (!n_n4775) & (x15754x)) + ((n_n4782) & (!n_n4781) & (n_n4775) & (!x15754x)) + ((n_n4782) & (!n_n4781) & (n_n4775) & (x15754x)) + ((n_n4782) & (n_n4781) & (!n_n4775) & (!x15754x)) + ((n_n4782) & (n_n4781) & (!n_n4775) & (x15754x)) + ((n_n4782) & (n_n4781) & (n_n4775) & (!x15754x)) + ((n_n4782) & (n_n4781) & (n_n4775) & (x15754x)));
	assign n_n2977 = (((!n_n4784) & (!n_n4779) & (!n_n4786) & (!n_n4783) & (x15757x)) + ((!n_n4784) & (!n_n4779) & (!n_n4786) & (n_n4783) & (!x15757x)) + ((!n_n4784) & (!n_n4779) & (!n_n4786) & (n_n4783) & (x15757x)) + ((!n_n4784) & (!n_n4779) & (n_n4786) & (!n_n4783) & (!x15757x)) + ((!n_n4784) & (!n_n4779) & (n_n4786) & (!n_n4783) & (x15757x)) + ((!n_n4784) & (!n_n4779) & (n_n4786) & (n_n4783) & (!x15757x)) + ((!n_n4784) & (!n_n4779) & (n_n4786) & (n_n4783) & (x15757x)) + ((!n_n4784) & (n_n4779) & (!n_n4786) & (!n_n4783) & (!x15757x)) + ((!n_n4784) & (n_n4779) & (!n_n4786) & (!n_n4783) & (x15757x)) + ((!n_n4784) & (n_n4779) & (!n_n4786) & (n_n4783) & (!x15757x)) + ((!n_n4784) & (n_n4779) & (!n_n4786) & (n_n4783) & (x15757x)) + ((!n_n4784) & (n_n4779) & (n_n4786) & (!n_n4783) & (!x15757x)) + ((!n_n4784) & (n_n4779) & (n_n4786) & (!n_n4783) & (x15757x)) + ((!n_n4784) & (n_n4779) & (n_n4786) & (n_n4783) & (!x15757x)) + ((!n_n4784) & (n_n4779) & (n_n4786) & (n_n4783) & (x15757x)) + ((n_n4784) & (!n_n4779) & (!n_n4786) & (!n_n4783) & (!x15757x)) + ((n_n4784) & (!n_n4779) & (!n_n4786) & (!n_n4783) & (x15757x)) + ((n_n4784) & (!n_n4779) & (!n_n4786) & (n_n4783) & (!x15757x)) + ((n_n4784) & (!n_n4779) & (!n_n4786) & (n_n4783) & (x15757x)) + ((n_n4784) & (!n_n4779) & (n_n4786) & (!n_n4783) & (!x15757x)) + ((n_n4784) & (!n_n4779) & (n_n4786) & (!n_n4783) & (x15757x)) + ((n_n4784) & (!n_n4779) & (n_n4786) & (n_n4783) & (!x15757x)) + ((n_n4784) & (!n_n4779) & (n_n4786) & (n_n4783) & (x15757x)) + ((n_n4784) & (n_n4779) & (!n_n4786) & (!n_n4783) & (!x15757x)) + ((n_n4784) & (n_n4779) & (!n_n4786) & (!n_n4783) & (x15757x)) + ((n_n4784) & (n_n4779) & (!n_n4786) & (n_n4783) & (!x15757x)) + ((n_n4784) & (n_n4779) & (!n_n4786) & (n_n4783) & (x15757x)) + ((n_n4784) & (n_n4779) & (n_n4786) & (!n_n4783) & (!x15757x)) + ((n_n4784) & (n_n4779) & (n_n4786) & (!n_n4783) & (x15757x)) + ((n_n4784) & (n_n4779) & (n_n4786) & (n_n4783) & (!x15757x)) + ((n_n4784) & (n_n4779) & (n_n4786) & (n_n4783) & (x15757x)));
	assign x22172x = (((!n_n4926) & (!n_n4928) & (!n_n4925) & (!n_n4922)));
	assign n_n2966 = (((!n_n4920) & (!n_n4930) & (!n_n4919) & (!x382x) & (!x22172x)) + ((!n_n4920) & (!n_n4930) & (!n_n4919) & (x382x) & (!x22172x)) + ((!n_n4920) & (!n_n4930) & (!n_n4919) & (x382x) & (x22172x)) + ((!n_n4920) & (!n_n4930) & (n_n4919) & (!x382x) & (!x22172x)) + ((!n_n4920) & (!n_n4930) & (n_n4919) & (!x382x) & (x22172x)) + ((!n_n4920) & (!n_n4930) & (n_n4919) & (x382x) & (!x22172x)) + ((!n_n4920) & (!n_n4930) & (n_n4919) & (x382x) & (x22172x)) + ((!n_n4920) & (n_n4930) & (!n_n4919) & (!x382x) & (!x22172x)) + ((!n_n4920) & (n_n4930) & (!n_n4919) & (!x382x) & (x22172x)) + ((!n_n4920) & (n_n4930) & (!n_n4919) & (x382x) & (!x22172x)) + ((!n_n4920) & (n_n4930) & (!n_n4919) & (x382x) & (x22172x)) + ((!n_n4920) & (n_n4930) & (n_n4919) & (!x382x) & (!x22172x)) + ((!n_n4920) & (n_n4930) & (n_n4919) & (!x382x) & (x22172x)) + ((!n_n4920) & (n_n4930) & (n_n4919) & (x382x) & (!x22172x)) + ((!n_n4920) & (n_n4930) & (n_n4919) & (x382x) & (x22172x)) + ((n_n4920) & (!n_n4930) & (!n_n4919) & (!x382x) & (!x22172x)) + ((n_n4920) & (!n_n4930) & (!n_n4919) & (!x382x) & (x22172x)) + ((n_n4920) & (!n_n4930) & (!n_n4919) & (x382x) & (!x22172x)) + ((n_n4920) & (!n_n4930) & (!n_n4919) & (x382x) & (x22172x)) + ((n_n4920) & (!n_n4930) & (n_n4919) & (!x382x) & (!x22172x)) + ((n_n4920) & (!n_n4930) & (n_n4919) & (!x382x) & (x22172x)) + ((n_n4920) & (!n_n4930) & (n_n4919) & (x382x) & (!x22172x)) + ((n_n4920) & (!n_n4930) & (n_n4919) & (x382x) & (x22172x)) + ((n_n4920) & (n_n4930) & (!n_n4919) & (!x382x) & (!x22172x)) + ((n_n4920) & (n_n4930) & (!n_n4919) & (!x382x) & (x22172x)) + ((n_n4920) & (n_n4930) & (!n_n4919) & (x382x) & (!x22172x)) + ((n_n4920) & (n_n4930) & (!n_n4919) & (x382x) & (x22172x)) + ((n_n4920) & (n_n4930) & (n_n4919) & (!x382x) & (!x22172x)) + ((n_n4920) & (n_n4930) & (n_n4919) & (!x382x) & (x22172x)) + ((n_n4920) & (n_n4930) & (n_n4919) & (x382x) & (!x22172x)) + ((n_n4920) & (n_n4930) & (n_n4919) & (x382x) & (x22172x)));
	assign n_n5317 = (((i_5_) & (!i_3_) & (!i_4_) & (x20x) & (n_n65)));
	assign n_n2803 = (((!n_n536) & (!n_n473) & (!x20x) & (x215x)) + ((!n_n536) & (!n_n473) & (x20x) & (x215x)) + ((!n_n536) & (n_n473) & (!x20x) & (x215x)) + ((!n_n536) & (n_n473) & (x20x) & (x215x)) + ((n_n536) & (!n_n473) & (!x20x) & (x215x)) + ((n_n536) & (!n_n473) & (x20x) & (x215x)) + ((n_n536) & (n_n473) & (!x20x) & (x215x)) + ((n_n536) & (n_n473) & (x20x) & (!x215x)) + ((n_n536) & (n_n473) & (x20x) & (x215x)));
	assign x304x = (((!i_7_) & (i_8_) & (!i_6_) & (x17x) & (n_n535)) + ((i_7_) & (!i_8_) & (!i_6_) & (x17x) & (n_n535)));
	assign x22216x = (((!n_n5254) & (!n_n5256) & (!n_n5253) & (!n_n3031) & (!n_n5257)));
	assign n_n2568 = (((!x19x) & (!n_n532) & (!n_n500) & (!n_n5255) & (!x22216x)) + ((!x19x) & (!n_n532) & (!n_n500) & (n_n5255) & (!x22216x)) + ((!x19x) & (!n_n532) & (!n_n500) & (n_n5255) & (x22216x)) + ((!x19x) & (!n_n532) & (n_n500) & (!n_n5255) & (!x22216x)) + ((!x19x) & (!n_n532) & (n_n500) & (n_n5255) & (!x22216x)) + ((!x19x) & (!n_n532) & (n_n500) & (n_n5255) & (x22216x)) + ((!x19x) & (n_n532) & (!n_n500) & (!n_n5255) & (!x22216x)) + ((!x19x) & (n_n532) & (!n_n500) & (n_n5255) & (!x22216x)) + ((!x19x) & (n_n532) & (!n_n500) & (n_n5255) & (x22216x)) + ((!x19x) & (n_n532) & (n_n500) & (!n_n5255) & (!x22216x)) + ((!x19x) & (n_n532) & (n_n500) & (n_n5255) & (!x22216x)) + ((!x19x) & (n_n532) & (n_n500) & (n_n5255) & (x22216x)) + ((x19x) & (!n_n532) & (!n_n500) & (!n_n5255) & (!x22216x)) + ((x19x) & (!n_n532) & (!n_n500) & (n_n5255) & (!x22216x)) + ((x19x) & (!n_n532) & (!n_n500) & (n_n5255) & (x22216x)) + ((x19x) & (!n_n532) & (n_n500) & (!n_n5255) & (!x22216x)) + ((x19x) & (!n_n532) & (n_n500) & (n_n5255) & (!x22216x)) + ((x19x) & (!n_n532) & (n_n500) & (n_n5255) & (x22216x)) + ((x19x) & (n_n532) & (!n_n500) & (!n_n5255) & (!x22216x)) + ((x19x) & (n_n532) & (!n_n500) & (n_n5255) & (!x22216x)) + ((x19x) & (n_n532) & (!n_n500) & (n_n5255) & (x22216x)) + ((x19x) & (n_n532) & (n_n500) & (!n_n5255) & (!x22216x)) + ((x19x) & (n_n532) & (n_n500) & (!n_n5255) & (x22216x)) + ((x19x) & (n_n532) & (n_n500) & (n_n5255) & (!x22216x)) + ((x19x) & (n_n532) & (n_n500) & (n_n5255) & (x22216x)));
	assign x146x = (((!x19x) & (x24x) & (n_n509) & (!n_n530) & (n_n65)) + ((!x19x) & (x24x) & (n_n509) & (n_n530) & (n_n65)) + ((x19x) & (!x24x) & (n_n509) & (n_n530) & (!n_n65)) + ((x19x) & (!x24x) & (n_n509) & (n_n530) & (n_n65)) + ((x19x) & (x24x) & (n_n509) & (!n_n530) & (n_n65)) + ((x19x) & (x24x) & (n_n509) & (n_n530) & (!n_n65)) + ((x19x) & (x24x) & (n_n509) & (n_n530) & (n_n65)));
	assign x320x = (((n_n518) & (!x20x) & (x23x) & (n_n65)) + ((n_n518) & (x20x) & (!x23x) & (n_n65)) + ((n_n518) & (x20x) & (x23x) & (n_n65)));
	assign x15177x = (((!x19x) & (!n_n528) & (!n_n532) & (!n_n509) & (n_n5247)) + ((!x19x) & (!n_n528) & (!n_n532) & (n_n509) & (n_n5247)) + ((!x19x) & (!n_n528) & (n_n532) & (!n_n509) & (n_n5247)) + ((!x19x) & (!n_n528) & (n_n532) & (n_n509) & (n_n5247)) + ((!x19x) & (n_n528) & (!n_n532) & (!n_n509) & (n_n5247)) + ((!x19x) & (n_n528) & (!n_n532) & (n_n509) & (n_n5247)) + ((!x19x) & (n_n528) & (n_n532) & (!n_n509) & (n_n5247)) + ((!x19x) & (n_n528) & (n_n532) & (n_n509) & (n_n5247)) + ((x19x) & (!n_n528) & (!n_n532) & (!n_n509) & (n_n5247)) + ((x19x) & (!n_n528) & (!n_n532) & (n_n509) & (n_n5247)) + ((x19x) & (!n_n528) & (n_n532) & (!n_n509) & (n_n5247)) + ((x19x) & (!n_n528) & (n_n532) & (n_n509) & (!n_n5247)) + ((x19x) & (!n_n528) & (n_n532) & (n_n509) & (n_n5247)) + ((x19x) & (n_n528) & (!n_n532) & (!n_n509) & (n_n5247)) + ((x19x) & (n_n528) & (!n_n532) & (n_n509) & (!n_n5247)) + ((x19x) & (n_n528) & (!n_n532) & (n_n509) & (n_n5247)) + ((x19x) & (n_n528) & (n_n532) & (!n_n509) & (n_n5247)) + ((x19x) & (n_n528) & (n_n532) & (n_n509) & (!n_n5247)) + ((x19x) & (n_n528) & (n_n532) & (n_n509) & (n_n5247)));
	assign n_n2569 = (((!n_n5238) & (!n_n5249) & (!x146x) & (!x320x) & (x15177x)) + ((!n_n5238) & (!n_n5249) & (!x146x) & (x320x) & (!x15177x)) + ((!n_n5238) & (!n_n5249) & (!x146x) & (x320x) & (x15177x)) + ((!n_n5238) & (!n_n5249) & (x146x) & (!x320x) & (!x15177x)) + ((!n_n5238) & (!n_n5249) & (x146x) & (!x320x) & (x15177x)) + ((!n_n5238) & (!n_n5249) & (x146x) & (x320x) & (!x15177x)) + ((!n_n5238) & (!n_n5249) & (x146x) & (x320x) & (x15177x)) + ((!n_n5238) & (n_n5249) & (!x146x) & (!x320x) & (!x15177x)) + ((!n_n5238) & (n_n5249) & (!x146x) & (!x320x) & (x15177x)) + ((!n_n5238) & (n_n5249) & (!x146x) & (x320x) & (!x15177x)) + ((!n_n5238) & (n_n5249) & (!x146x) & (x320x) & (x15177x)) + ((!n_n5238) & (n_n5249) & (x146x) & (!x320x) & (!x15177x)) + ((!n_n5238) & (n_n5249) & (x146x) & (!x320x) & (x15177x)) + ((!n_n5238) & (n_n5249) & (x146x) & (x320x) & (!x15177x)) + ((!n_n5238) & (n_n5249) & (x146x) & (x320x) & (x15177x)) + ((n_n5238) & (!n_n5249) & (!x146x) & (!x320x) & (!x15177x)) + ((n_n5238) & (!n_n5249) & (!x146x) & (!x320x) & (x15177x)) + ((n_n5238) & (!n_n5249) & (!x146x) & (x320x) & (!x15177x)) + ((n_n5238) & (!n_n5249) & (!x146x) & (x320x) & (x15177x)) + ((n_n5238) & (!n_n5249) & (x146x) & (!x320x) & (!x15177x)) + ((n_n5238) & (!n_n5249) & (x146x) & (!x320x) & (x15177x)) + ((n_n5238) & (!n_n5249) & (x146x) & (x320x) & (!x15177x)) + ((n_n5238) & (!n_n5249) & (x146x) & (x320x) & (x15177x)) + ((n_n5238) & (n_n5249) & (!x146x) & (!x320x) & (!x15177x)) + ((n_n5238) & (n_n5249) & (!x146x) & (!x320x) & (x15177x)) + ((n_n5238) & (n_n5249) & (!x146x) & (x320x) & (!x15177x)) + ((n_n5238) & (n_n5249) & (!x146x) & (x320x) & (x15177x)) + ((n_n5238) & (n_n5249) & (x146x) & (!x320x) & (!x15177x)) + ((n_n5238) & (n_n5249) & (x146x) & (!x320x) & (x15177x)) + ((n_n5238) & (n_n5249) & (x146x) & (x320x) & (!x15177x)) + ((n_n5238) & (n_n5249) & (x146x) & (x320x) & (x15177x)));
	assign n_n5264 = (((i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n500)));
	assign x334x = (((!i_9_) & (!x19x) & (n_n524) & (n_n500) & (n_n65)) + ((!i_9_) & (x19x) & (n_n524) & (n_n500) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n524) & (n_n500) & (n_n65)) + ((i_9_) & (x19x) & (n_n524) & (n_n500) & (!n_n65)) + ((i_9_) & (x19x) & (n_n524) & (n_n500) & (n_n65)));
	assign x22185x = (((!x19x) & (!n_n526) & (!n_n520) & (!n_n500) & (!n_n5265)) + ((!x19x) & (!n_n526) & (!n_n520) & (n_n500) & (!n_n5265)) + ((!x19x) & (!n_n526) & (n_n520) & (!n_n500) & (!n_n5265)) + ((!x19x) & (!n_n526) & (n_n520) & (n_n500) & (!n_n5265)) + ((!x19x) & (n_n526) & (!n_n520) & (!n_n500) & (!n_n5265)) + ((!x19x) & (n_n526) & (!n_n520) & (n_n500) & (!n_n5265)) + ((!x19x) & (n_n526) & (n_n520) & (!n_n500) & (!n_n5265)) + ((!x19x) & (n_n526) & (n_n520) & (n_n500) & (!n_n5265)) + ((x19x) & (!n_n526) & (!n_n520) & (!n_n500) & (!n_n5265)) + ((x19x) & (!n_n526) & (!n_n520) & (n_n500) & (!n_n5265)) + ((x19x) & (!n_n526) & (n_n520) & (!n_n500) & (!n_n5265)) + ((x19x) & (n_n526) & (!n_n520) & (!n_n500) & (!n_n5265)) + ((x19x) & (n_n526) & (n_n520) & (!n_n500) & (!n_n5265)));
	assign x15184x = (((!n_n5262) & (!n_n5259) & (!x77x) & (!x334x) & (!x22185x)) + ((!n_n5262) & (!n_n5259) & (!x77x) & (x334x) & (!x22185x)) + ((!n_n5262) & (!n_n5259) & (!x77x) & (x334x) & (x22185x)) + ((!n_n5262) & (!n_n5259) & (x77x) & (!x334x) & (!x22185x)) + ((!n_n5262) & (!n_n5259) & (x77x) & (!x334x) & (x22185x)) + ((!n_n5262) & (!n_n5259) & (x77x) & (x334x) & (!x22185x)) + ((!n_n5262) & (!n_n5259) & (x77x) & (x334x) & (x22185x)) + ((!n_n5262) & (n_n5259) & (!x77x) & (!x334x) & (!x22185x)) + ((!n_n5262) & (n_n5259) & (!x77x) & (!x334x) & (x22185x)) + ((!n_n5262) & (n_n5259) & (!x77x) & (x334x) & (!x22185x)) + ((!n_n5262) & (n_n5259) & (!x77x) & (x334x) & (x22185x)) + ((!n_n5262) & (n_n5259) & (x77x) & (!x334x) & (!x22185x)) + ((!n_n5262) & (n_n5259) & (x77x) & (!x334x) & (x22185x)) + ((!n_n5262) & (n_n5259) & (x77x) & (x334x) & (!x22185x)) + ((!n_n5262) & (n_n5259) & (x77x) & (x334x) & (x22185x)) + ((n_n5262) & (!n_n5259) & (!x77x) & (!x334x) & (!x22185x)) + ((n_n5262) & (!n_n5259) & (!x77x) & (!x334x) & (x22185x)) + ((n_n5262) & (!n_n5259) & (!x77x) & (x334x) & (!x22185x)) + ((n_n5262) & (!n_n5259) & (!x77x) & (x334x) & (x22185x)) + ((n_n5262) & (!n_n5259) & (x77x) & (!x334x) & (!x22185x)) + ((n_n5262) & (!n_n5259) & (x77x) & (!x334x) & (x22185x)) + ((n_n5262) & (!n_n5259) & (x77x) & (x334x) & (!x22185x)) + ((n_n5262) & (!n_n5259) & (x77x) & (x334x) & (x22185x)) + ((n_n5262) & (n_n5259) & (!x77x) & (!x334x) & (!x22185x)) + ((n_n5262) & (n_n5259) & (!x77x) & (!x334x) & (x22185x)) + ((n_n5262) & (n_n5259) & (!x77x) & (x334x) & (!x22185x)) + ((n_n5262) & (n_n5259) & (!x77x) & (x334x) & (x22185x)) + ((n_n5262) & (n_n5259) & (x77x) & (!x334x) & (!x22185x)) + ((n_n5262) & (n_n5259) & (x77x) & (!x334x) & (x22185x)) + ((n_n5262) & (n_n5259) & (x77x) & (x334x) & (!x22185x)) + ((n_n5262) & (n_n5259) & (x77x) & (x334x) & (x22185x)));
	assign x267x = (((!x19x) & (!x506x) & (!x502x) & (!x115x) & (n_n5315)) + ((!x19x) & (!x506x) & (!x502x) & (x115x) & (!n_n5315)) + ((!x19x) & (!x506x) & (!x502x) & (x115x) & (n_n5315)) + ((!x19x) & (!x506x) & (x502x) & (!x115x) & (n_n5315)) + ((!x19x) & (!x506x) & (x502x) & (x115x) & (!n_n5315)) + ((!x19x) & (!x506x) & (x502x) & (x115x) & (n_n5315)) + ((!x19x) & (x506x) & (!x502x) & (!x115x) & (n_n5315)) + ((!x19x) & (x506x) & (!x502x) & (x115x) & (!n_n5315)) + ((!x19x) & (x506x) & (!x502x) & (x115x) & (n_n5315)) + ((!x19x) & (x506x) & (x502x) & (!x115x) & (n_n5315)) + ((!x19x) & (x506x) & (x502x) & (x115x) & (!n_n5315)) + ((!x19x) & (x506x) & (x502x) & (x115x) & (n_n5315)) + ((x19x) & (!x506x) & (!x502x) & (!x115x) & (n_n5315)) + ((x19x) & (!x506x) & (!x502x) & (x115x) & (!n_n5315)) + ((x19x) & (!x506x) & (!x502x) & (x115x) & (n_n5315)) + ((x19x) & (!x506x) & (x502x) & (!x115x) & (!n_n5315)) + ((x19x) & (!x506x) & (x502x) & (!x115x) & (n_n5315)) + ((x19x) & (!x506x) & (x502x) & (x115x) & (!n_n5315)) + ((x19x) & (!x506x) & (x502x) & (x115x) & (n_n5315)) + ((x19x) & (x506x) & (!x502x) & (!x115x) & (!n_n5315)) + ((x19x) & (x506x) & (!x502x) & (!x115x) & (n_n5315)) + ((x19x) & (x506x) & (!x502x) & (x115x) & (!n_n5315)) + ((x19x) & (x506x) & (!x502x) & (x115x) & (n_n5315)) + ((x19x) & (x506x) & (x502x) & (!x115x) & (!n_n5315)) + ((x19x) & (x506x) & (x502x) & (!x115x) & (n_n5315)) + ((x19x) & (x506x) & (x502x) & (x115x) & (!n_n5315)) + ((x19x) & (x506x) & (x502x) & (x115x) & (n_n5315)));
	assign x15191x = (((!n_n5321) & (!n_n5319) & (!n_n5332) & (!n_n5334) & (x267x)) + ((!n_n5321) & (!n_n5319) & (!n_n5332) & (n_n5334) & (!x267x)) + ((!n_n5321) & (!n_n5319) & (!n_n5332) & (n_n5334) & (x267x)) + ((!n_n5321) & (!n_n5319) & (n_n5332) & (!n_n5334) & (!x267x)) + ((!n_n5321) & (!n_n5319) & (n_n5332) & (!n_n5334) & (x267x)) + ((!n_n5321) & (!n_n5319) & (n_n5332) & (n_n5334) & (!x267x)) + ((!n_n5321) & (!n_n5319) & (n_n5332) & (n_n5334) & (x267x)) + ((!n_n5321) & (n_n5319) & (!n_n5332) & (!n_n5334) & (!x267x)) + ((!n_n5321) & (n_n5319) & (!n_n5332) & (!n_n5334) & (x267x)) + ((!n_n5321) & (n_n5319) & (!n_n5332) & (n_n5334) & (!x267x)) + ((!n_n5321) & (n_n5319) & (!n_n5332) & (n_n5334) & (x267x)) + ((!n_n5321) & (n_n5319) & (n_n5332) & (!n_n5334) & (!x267x)) + ((!n_n5321) & (n_n5319) & (n_n5332) & (!n_n5334) & (x267x)) + ((!n_n5321) & (n_n5319) & (n_n5332) & (n_n5334) & (!x267x)) + ((!n_n5321) & (n_n5319) & (n_n5332) & (n_n5334) & (x267x)) + ((n_n5321) & (!n_n5319) & (!n_n5332) & (!n_n5334) & (!x267x)) + ((n_n5321) & (!n_n5319) & (!n_n5332) & (!n_n5334) & (x267x)) + ((n_n5321) & (!n_n5319) & (!n_n5332) & (n_n5334) & (!x267x)) + ((n_n5321) & (!n_n5319) & (!n_n5332) & (n_n5334) & (x267x)) + ((n_n5321) & (!n_n5319) & (n_n5332) & (!n_n5334) & (!x267x)) + ((n_n5321) & (!n_n5319) & (n_n5332) & (!n_n5334) & (x267x)) + ((n_n5321) & (!n_n5319) & (n_n5332) & (n_n5334) & (!x267x)) + ((n_n5321) & (!n_n5319) & (n_n5332) & (n_n5334) & (x267x)) + ((n_n5321) & (n_n5319) & (!n_n5332) & (!n_n5334) & (!x267x)) + ((n_n5321) & (n_n5319) & (!n_n5332) & (!n_n5334) & (x267x)) + ((n_n5321) & (n_n5319) & (!n_n5332) & (n_n5334) & (!x267x)) + ((n_n5321) & (n_n5319) & (!n_n5332) & (n_n5334) & (x267x)) + ((n_n5321) & (n_n5319) & (n_n5332) & (!n_n5334) & (!x267x)) + ((n_n5321) & (n_n5319) & (n_n5332) & (!n_n5334) & (x267x)) + ((n_n5321) & (n_n5319) & (n_n5332) & (n_n5334) & (!x267x)) + ((n_n5321) & (n_n5319) & (n_n5332) & (n_n5334) & (x267x)));
	assign x22188x = (((!x19x) & (!n_n5331) & (!x516x) & (!n_n5322) & (!n_n5328)) + ((!x19x) & (!n_n5331) & (x516x) & (!n_n5322) & (!n_n5328)) + ((x19x) & (!n_n5331) & (!x516x) & (!n_n5322) & (!n_n5328)));
	assign x15192x = (((!n_n5312) & (!n_n2643) & (!n_n3019) & (!x22188x)) + ((!n_n5312) & (!n_n2643) & (n_n3019) & (!x22188x)) + ((!n_n5312) & (!n_n2643) & (n_n3019) & (x22188x)) + ((!n_n5312) & (n_n2643) & (!n_n3019) & (!x22188x)) + ((!n_n5312) & (n_n2643) & (!n_n3019) & (x22188x)) + ((!n_n5312) & (n_n2643) & (n_n3019) & (!x22188x)) + ((!n_n5312) & (n_n2643) & (n_n3019) & (x22188x)) + ((n_n5312) & (!n_n2643) & (!n_n3019) & (!x22188x)) + ((n_n5312) & (!n_n2643) & (!n_n3019) & (x22188x)) + ((n_n5312) & (!n_n2643) & (n_n3019) & (!x22188x)) + ((n_n5312) & (!n_n2643) & (n_n3019) & (x22188x)) + ((n_n5312) & (n_n2643) & (!n_n3019) & (!x22188x)) + ((n_n5312) & (n_n2643) & (!n_n3019) & (x22188x)) + ((n_n5312) & (n_n2643) & (n_n3019) & (!x22188x)) + ((n_n5312) & (n_n2643) & (n_n3019) & (x22188x)));
	assign x15196x = (((!n_n5305) & (!n_n5297) & (!n_n5302) & (!n_n5295) & (n_n5298)) + ((!n_n5305) & (!n_n5297) & (!n_n5302) & (n_n5295) & (!n_n5298)) + ((!n_n5305) & (!n_n5297) & (!n_n5302) & (n_n5295) & (n_n5298)) + ((!n_n5305) & (!n_n5297) & (n_n5302) & (!n_n5295) & (!n_n5298)) + ((!n_n5305) & (!n_n5297) & (n_n5302) & (!n_n5295) & (n_n5298)) + ((!n_n5305) & (!n_n5297) & (n_n5302) & (n_n5295) & (!n_n5298)) + ((!n_n5305) & (!n_n5297) & (n_n5302) & (n_n5295) & (n_n5298)) + ((!n_n5305) & (n_n5297) & (!n_n5302) & (!n_n5295) & (!n_n5298)) + ((!n_n5305) & (n_n5297) & (!n_n5302) & (!n_n5295) & (n_n5298)) + ((!n_n5305) & (n_n5297) & (!n_n5302) & (n_n5295) & (!n_n5298)) + ((!n_n5305) & (n_n5297) & (!n_n5302) & (n_n5295) & (n_n5298)) + ((!n_n5305) & (n_n5297) & (n_n5302) & (!n_n5295) & (!n_n5298)) + ((!n_n5305) & (n_n5297) & (n_n5302) & (!n_n5295) & (n_n5298)) + ((!n_n5305) & (n_n5297) & (n_n5302) & (n_n5295) & (!n_n5298)) + ((!n_n5305) & (n_n5297) & (n_n5302) & (n_n5295) & (n_n5298)) + ((n_n5305) & (!n_n5297) & (!n_n5302) & (!n_n5295) & (!n_n5298)) + ((n_n5305) & (!n_n5297) & (!n_n5302) & (!n_n5295) & (n_n5298)) + ((n_n5305) & (!n_n5297) & (!n_n5302) & (n_n5295) & (!n_n5298)) + ((n_n5305) & (!n_n5297) & (!n_n5302) & (n_n5295) & (n_n5298)) + ((n_n5305) & (!n_n5297) & (n_n5302) & (!n_n5295) & (!n_n5298)) + ((n_n5305) & (!n_n5297) & (n_n5302) & (!n_n5295) & (n_n5298)) + ((n_n5305) & (!n_n5297) & (n_n5302) & (n_n5295) & (!n_n5298)) + ((n_n5305) & (!n_n5297) & (n_n5302) & (n_n5295) & (n_n5298)) + ((n_n5305) & (n_n5297) & (!n_n5302) & (!n_n5295) & (!n_n5298)) + ((n_n5305) & (n_n5297) & (!n_n5302) & (!n_n5295) & (n_n5298)) + ((n_n5305) & (n_n5297) & (!n_n5302) & (n_n5295) & (!n_n5298)) + ((n_n5305) & (n_n5297) & (!n_n5302) & (n_n5295) & (n_n5298)) + ((n_n5305) & (n_n5297) & (n_n5302) & (!n_n5295) & (!n_n5298)) + ((n_n5305) & (n_n5297) & (n_n5302) & (!n_n5295) & (n_n5298)) + ((n_n5305) & (n_n5297) & (n_n5302) & (n_n5295) & (!n_n5298)) + ((n_n5305) & (n_n5297) & (n_n5302) & (n_n5295) & (n_n5298)));
	assign n_n2651 = (((!x11x) & (!n_n491) & (!n_n65) & (!n_n5281) & (n_n5280)) + ((!x11x) & (!n_n491) & (!n_n65) & (n_n5281) & (!n_n5280)) + ((!x11x) & (!n_n491) & (!n_n65) & (n_n5281) & (n_n5280)) + ((!x11x) & (!n_n491) & (n_n65) & (!n_n5281) & (n_n5280)) + ((!x11x) & (!n_n491) & (n_n65) & (n_n5281) & (!n_n5280)) + ((!x11x) & (!n_n491) & (n_n65) & (n_n5281) & (n_n5280)) + ((!x11x) & (n_n491) & (!n_n65) & (!n_n5281) & (n_n5280)) + ((!x11x) & (n_n491) & (!n_n65) & (n_n5281) & (!n_n5280)) + ((!x11x) & (n_n491) & (!n_n65) & (n_n5281) & (n_n5280)) + ((!x11x) & (n_n491) & (n_n65) & (!n_n5281) & (n_n5280)) + ((!x11x) & (n_n491) & (n_n65) & (n_n5281) & (!n_n5280)) + ((!x11x) & (n_n491) & (n_n65) & (n_n5281) & (n_n5280)) + ((x11x) & (!n_n491) & (!n_n65) & (!n_n5281) & (n_n5280)) + ((x11x) & (!n_n491) & (!n_n65) & (n_n5281) & (!n_n5280)) + ((x11x) & (!n_n491) & (!n_n65) & (n_n5281) & (n_n5280)) + ((x11x) & (!n_n491) & (n_n65) & (!n_n5281) & (n_n5280)) + ((x11x) & (!n_n491) & (n_n65) & (n_n5281) & (!n_n5280)) + ((x11x) & (!n_n491) & (n_n65) & (n_n5281) & (n_n5280)) + ((x11x) & (n_n491) & (!n_n65) & (!n_n5281) & (n_n5280)) + ((x11x) & (n_n491) & (!n_n65) & (n_n5281) & (!n_n5280)) + ((x11x) & (n_n491) & (!n_n65) & (n_n5281) & (n_n5280)) + ((x11x) & (n_n491) & (n_n65) & (!n_n5281) & (!n_n5280)) + ((x11x) & (n_n491) & (n_n65) & (!n_n5281) & (n_n5280)) + ((x11x) & (n_n491) & (n_n65) & (n_n5281) & (!n_n5280)) + ((x11x) & (n_n491) & (n_n65) & (n_n5281) & (n_n5280)));
	assign x203x = (((!i_9_) & (!x19x) & (n_n534) & (n_n491) & (n_n65)) + ((!i_9_) & (x19x) & (n_n534) & (n_n491) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n534) & (n_n491) & (n_n65)) + ((i_9_) & (x19x) & (n_n534) & (n_n491) & (!n_n65)) + ((i_9_) & (x19x) & (n_n534) & (n_n491) & (n_n65)));
	assign x438x = (((!i_9_) & (!x19x) & (n_n491) & (n_n530) & (n_n65)) + ((!i_9_) & (x19x) & (n_n491) & (n_n530) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n491) & (n_n530) & (n_n65)) + ((i_9_) & (x19x) & (n_n491) & (n_n530) & (!n_n65)) + ((i_9_) & (x19x) & (n_n491) & (n_n530) & (n_n65)));
	assign n_n2566 = (((!n_n5274) & (!n_n5271) & (!n_n2651) & (!x203x) & (x438x)) + ((!n_n5274) & (!n_n5271) & (!n_n2651) & (x203x) & (!x438x)) + ((!n_n5274) & (!n_n5271) & (!n_n2651) & (x203x) & (x438x)) + ((!n_n5274) & (!n_n5271) & (n_n2651) & (!x203x) & (!x438x)) + ((!n_n5274) & (!n_n5271) & (n_n2651) & (!x203x) & (x438x)) + ((!n_n5274) & (!n_n5271) & (n_n2651) & (x203x) & (!x438x)) + ((!n_n5274) & (!n_n5271) & (n_n2651) & (x203x) & (x438x)) + ((!n_n5274) & (n_n5271) & (!n_n2651) & (!x203x) & (!x438x)) + ((!n_n5274) & (n_n5271) & (!n_n2651) & (!x203x) & (x438x)) + ((!n_n5274) & (n_n5271) & (!n_n2651) & (x203x) & (!x438x)) + ((!n_n5274) & (n_n5271) & (!n_n2651) & (x203x) & (x438x)) + ((!n_n5274) & (n_n5271) & (n_n2651) & (!x203x) & (!x438x)) + ((!n_n5274) & (n_n5271) & (n_n2651) & (!x203x) & (x438x)) + ((!n_n5274) & (n_n5271) & (n_n2651) & (x203x) & (!x438x)) + ((!n_n5274) & (n_n5271) & (n_n2651) & (x203x) & (x438x)) + ((n_n5274) & (!n_n5271) & (!n_n2651) & (!x203x) & (!x438x)) + ((n_n5274) & (!n_n5271) & (!n_n2651) & (!x203x) & (x438x)) + ((n_n5274) & (!n_n5271) & (!n_n2651) & (x203x) & (!x438x)) + ((n_n5274) & (!n_n5271) & (!n_n2651) & (x203x) & (x438x)) + ((n_n5274) & (!n_n5271) & (n_n2651) & (!x203x) & (!x438x)) + ((n_n5274) & (!n_n5271) & (n_n2651) & (!x203x) & (x438x)) + ((n_n5274) & (!n_n5271) & (n_n2651) & (x203x) & (!x438x)) + ((n_n5274) & (!n_n5271) & (n_n2651) & (x203x) & (x438x)) + ((n_n5274) & (n_n5271) & (!n_n2651) & (!x203x) & (!x438x)) + ((n_n5274) & (n_n5271) & (!n_n2651) & (!x203x) & (x438x)) + ((n_n5274) & (n_n5271) & (!n_n2651) & (x203x) & (!x438x)) + ((n_n5274) & (n_n5271) & (!n_n2651) & (x203x) & (x438x)) + ((n_n5274) & (n_n5271) & (n_n2651) & (!x203x) & (!x438x)) + ((n_n5274) & (n_n5271) & (n_n2651) & (!x203x) & (x438x)) + ((n_n5274) & (n_n5271) & (n_n2651) & (x203x) & (!x438x)) + ((n_n5274) & (n_n5271) & (n_n2651) & (x203x) & (x438x)));
	assign x197x = (((!x15x) & (x19x) & (n_n482) & (n_n528) & (!n_n65)) + ((!x15x) & (x19x) & (n_n482) & (n_n528) & (n_n65)) + ((x15x) & (!x19x) & (n_n482) & (!n_n528) & (n_n65)) + ((x15x) & (!x19x) & (n_n482) & (n_n528) & (n_n65)) + ((x15x) & (x19x) & (n_n482) & (!n_n528) & (n_n65)) + ((x15x) & (x19x) & (n_n482) & (n_n528) & (!n_n65)) + ((x15x) & (x19x) & (n_n482) & (n_n528) & (n_n65)));
	assign x207x = (((x19x) & (!n_n482) & (!n_n534) & (n_n491) & (n_n520)) + ((x19x) & (!n_n482) & (n_n534) & (n_n491) & (n_n520)) + ((x19x) & (n_n482) & (!n_n534) & (n_n491) & (n_n520)) + ((x19x) & (n_n482) & (n_n534) & (!n_n491) & (!n_n520)) + ((x19x) & (n_n482) & (n_n534) & (!n_n491) & (n_n520)) + ((x19x) & (n_n482) & (n_n534) & (n_n491) & (!n_n520)) + ((x19x) & (n_n482) & (n_n534) & (n_n491) & (n_n520)));
	assign n_n5282 = (((i_7_) & (!i_8_) & (!i_6_) & (x19x) & (n_n491)));
	assign x218x = (((!i_9_) & (!x19x) & (n_n524) & (n_n491) & (n_n65)) + ((!i_9_) & (x19x) & (n_n524) & (n_n491) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n524) & (n_n491) & (n_n65)) + ((i_9_) & (x19x) & (n_n524) & (n_n491) & (!n_n65)) + ((i_9_) & (x19x) & (n_n524) & (n_n491) & (n_n65)));
	assign x15203x = (((!x592x) & (!x24x) & (!n_n5290) & (!n_n5285) & (x197x)) + ((!x592x) & (!x24x) & (!n_n5290) & (n_n5285) & (!x197x)) + ((!x592x) & (!x24x) & (!n_n5290) & (n_n5285) & (x197x)) + ((!x592x) & (!x24x) & (n_n5290) & (!n_n5285) & (!x197x)) + ((!x592x) & (!x24x) & (n_n5290) & (!n_n5285) & (x197x)) + ((!x592x) & (!x24x) & (n_n5290) & (n_n5285) & (!x197x)) + ((!x592x) & (!x24x) & (n_n5290) & (n_n5285) & (x197x)) + ((!x592x) & (x24x) & (!n_n5290) & (!n_n5285) & (x197x)) + ((!x592x) & (x24x) & (!n_n5290) & (n_n5285) & (!x197x)) + ((!x592x) & (x24x) & (!n_n5290) & (n_n5285) & (x197x)) + ((!x592x) & (x24x) & (n_n5290) & (!n_n5285) & (!x197x)) + ((!x592x) & (x24x) & (n_n5290) & (!n_n5285) & (x197x)) + ((!x592x) & (x24x) & (n_n5290) & (n_n5285) & (!x197x)) + ((!x592x) & (x24x) & (n_n5290) & (n_n5285) & (x197x)) + ((x592x) & (!x24x) & (!n_n5290) & (!n_n5285) & (x197x)) + ((x592x) & (!x24x) & (!n_n5290) & (n_n5285) & (!x197x)) + ((x592x) & (!x24x) & (!n_n5290) & (n_n5285) & (x197x)) + ((x592x) & (!x24x) & (n_n5290) & (!n_n5285) & (!x197x)) + ((x592x) & (!x24x) & (n_n5290) & (!n_n5285) & (x197x)) + ((x592x) & (!x24x) & (n_n5290) & (n_n5285) & (!x197x)) + ((x592x) & (!x24x) & (n_n5290) & (n_n5285) & (x197x)) + ((x592x) & (x24x) & (!n_n5290) & (!n_n5285) & (!x197x)) + ((x592x) & (x24x) & (!n_n5290) & (!n_n5285) & (x197x)) + ((x592x) & (x24x) & (!n_n5290) & (n_n5285) & (!x197x)) + ((x592x) & (x24x) & (!n_n5290) & (n_n5285) & (x197x)) + ((x592x) & (x24x) & (n_n5290) & (!n_n5285) & (!x197x)) + ((x592x) & (x24x) & (n_n5290) & (!n_n5285) & (x197x)) + ((x592x) & (x24x) & (n_n5290) & (n_n5285) & (!x197x)) + ((x592x) & (x24x) & (n_n5290) & (n_n5285) & (x197x)));
	assign x15206x = (((!x15191x) & (!x15192x) & (!x207x) & (!x218x) & (x15203x)) + ((!x15191x) & (!x15192x) & (!x207x) & (x218x) & (!x15203x)) + ((!x15191x) & (!x15192x) & (!x207x) & (x218x) & (x15203x)) + ((!x15191x) & (!x15192x) & (x207x) & (!x218x) & (!x15203x)) + ((!x15191x) & (!x15192x) & (x207x) & (!x218x) & (x15203x)) + ((!x15191x) & (!x15192x) & (x207x) & (x218x) & (!x15203x)) + ((!x15191x) & (!x15192x) & (x207x) & (x218x) & (x15203x)) + ((!x15191x) & (x15192x) & (!x207x) & (!x218x) & (!x15203x)) + ((!x15191x) & (x15192x) & (!x207x) & (!x218x) & (x15203x)) + ((!x15191x) & (x15192x) & (!x207x) & (x218x) & (!x15203x)) + ((!x15191x) & (x15192x) & (!x207x) & (x218x) & (x15203x)) + ((!x15191x) & (x15192x) & (x207x) & (!x218x) & (!x15203x)) + ((!x15191x) & (x15192x) & (x207x) & (!x218x) & (x15203x)) + ((!x15191x) & (x15192x) & (x207x) & (x218x) & (!x15203x)) + ((!x15191x) & (x15192x) & (x207x) & (x218x) & (x15203x)) + ((x15191x) & (!x15192x) & (!x207x) & (!x218x) & (!x15203x)) + ((x15191x) & (!x15192x) & (!x207x) & (!x218x) & (x15203x)) + ((x15191x) & (!x15192x) & (!x207x) & (x218x) & (!x15203x)) + ((x15191x) & (!x15192x) & (!x207x) & (x218x) & (x15203x)) + ((x15191x) & (!x15192x) & (x207x) & (!x218x) & (!x15203x)) + ((x15191x) & (!x15192x) & (x207x) & (!x218x) & (x15203x)) + ((x15191x) & (!x15192x) & (x207x) & (x218x) & (!x15203x)) + ((x15191x) & (!x15192x) & (x207x) & (x218x) & (x15203x)) + ((x15191x) & (x15192x) & (!x207x) & (!x218x) & (!x15203x)) + ((x15191x) & (x15192x) & (!x207x) & (!x218x) & (x15203x)) + ((x15191x) & (x15192x) & (!x207x) & (x218x) & (!x15203x)) + ((x15191x) & (x15192x) & (!x207x) & (x218x) & (x15203x)) + ((x15191x) & (x15192x) & (x207x) & (!x218x) & (!x15203x)) + ((x15191x) & (x15192x) & (x207x) & (!x218x) & (x15203x)) + ((x15191x) & (x15192x) & (x207x) & (x218x) & (!x15203x)) + ((x15191x) & (x15192x) & (x207x) & (x218x) & (x15203x)));
	assign x15205x = (((!n_n5303) & (!x15196x) & (!n_n2566) & (!x63x) & (n_n5304)) + ((!n_n5303) & (!x15196x) & (!n_n2566) & (x63x) & (!n_n5304)) + ((!n_n5303) & (!x15196x) & (!n_n2566) & (x63x) & (n_n5304)) + ((!n_n5303) & (!x15196x) & (n_n2566) & (!x63x) & (!n_n5304)) + ((!n_n5303) & (!x15196x) & (n_n2566) & (!x63x) & (n_n5304)) + ((!n_n5303) & (!x15196x) & (n_n2566) & (x63x) & (!n_n5304)) + ((!n_n5303) & (!x15196x) & (n_n2566) & (x63x) & (n_n5304)) + ((!n_n5303) & (x15196x) & (!n_n2566) & (!x63x) & (!n_n5304)) + ((!n_n5303) & (x15196x) & (!n_n2566) & (!x63x) & (n_n5304)) + ((!n_n5303) & (x15196x) & (!n_n2566) & (x63x) & (!n_n5304)) + ((!n_n5303) & (x15196x) & (!n_n2566) & (x63x) & (n_n5304)) + ((!n_n5303) & (x15196x) & (n_n2566) & (!x63x) & (!n_n5304)) + ((!n_n5303) & (x15196x) & (n_n2566) & (!x63x) & (n_n5304)) + ((!n_n5303) & (x15196x) & (n_n2566) & (x63x) & (!n_n5304)) + ((!n_n5303) & (x15196x) & (n_n2566) & (x63x) & (n_n5304)) + ((n_n5303) & (!x15196x) & (!n_n2566) & (!x63x) & (!n_n5304)) + ((n_n5303) & (!x15196x) & (!n_n2566) & (!x63x) & (n_n5304)) + ((n_n5303) & (!x15196x) & (!n_n2566) & (x63x) & (!n_n5304)) + ((n_n5303) & (!x15196x) & (!n_n2566) & (x63x) & (n_n5304)) + ((n_n5303) & (!x15196x) & (n_n2566) & (!x63x) & (!n_n5304)) + ((n_n5303) & (!x15196x) & (n_n2566) & (!x63x) & (n_n5304)) + ((n_n5303) & (!x15196x) & (n_n2566) & (x63x) & (!n_n5304)) + ((n_n5303) & (!x15196x) & (n_n2566) & (x63x) & (n_n5304)) + ((n_n5303) & (x15196x) & (!n_n2566) & (!x63x) & (!n_n5304)) + ((n_n5303) & (x15196x) & (!n_n2566) & (!x63x) & (n_n5304)) + ((n_n5303) & (x15196x) & (!n_n2566) & (x63x) & (!n_n5304)) + ((n_n5303) & (x15196x) & (!n_n2566) & (x63x) & (n_n5304)) + ((n_n5303) & (x15196x) & (n_n2566) & (!x63x) & (!n_n5304)) + ((n_n5303) & (x15196x) & (n_n2566) & (!x63x) & (n_n5304)) + ((n_n5303) & (x15196x) & (n_n2566) & (x63x) & (!n_n5304)) + ((n_n5303) & (x15196x) & (n_n2566) & (x63x) & (n_n5304)));
	assign n_n5227 = (((!i_9_) & (n_n518) & (n_n532) & (n_n65)));
	assign x385x = (((!i_9_) & (!x19x) & (n_n518) & (n_n532) & (n_n65)) + ((!i_9_) & (x19x) & (n_n518) & (n_n532) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n518) & (n_n532) & (n_n65)) + ((i_9_) & (x19x) & (n_n518) & (n_n532) & (!n_n65)) + ((i_9_) & (x19x) & (n_n518) & (n_n532) & (n_n65)));
	assign x16750x = (((!x592x) & (!x21x) & (!x11x) & (!n_n5294) & (x208x)) + ((!x592x) & (!x21x) & (!x11x) & (n_n5294) & (!x208x)) + ((!x592x) & (!x21x) & (!x11x) & (n_n5294) & (x208x)) + ((!x592x) & (!x21x) & (x11x) & (!n_n5294) & (x208x)) + ((!x592x) & (!x21x) & (x11x) & (n_n5294) & (!x208x)) + ((!x592x) & (!x21x) & (x11x) & (n_n5294) & (x208x)) + ((!x592x) & (x21x) & (!x11x) & (!n_n5294) & (x208x)) + ((!x592x) & (x21x) & (!x11x) & (n_n5294) & (!x208x)) + ((!x592x) & (x21x) & (!x11x) & (n_n5294) & (x208x)) + ((!x592x) & (x21x) & (x11x) & (!n_n5294) & (x208x)) + ((!x592x) & (x21x) & (x11x) & (n_n5294) & (!x208x)) + ((!x592x) & (x21x) & (x11x) & (n_n5294) & (x208x)) + ((x592x) & (!x21x) & (!x11x) & (!n_n5294) & (x208x)) + ((x592x) & (!x21x) & (!x11x) & (n_n5294) & (!x208x)) + ((x592x) & (!x21x) & (!x11x) & (n_n5294) & (x208x)) + ((x592x) & (!x21x) & (x11x) & (!n_n5294) & (!x208x)) + ((x592x) & (!x21x) & (x11x) & (!n_n5294) & (x208x)) + ((x592x) & (!x21x) & (x11x) & (n_n5294) & (!x208x)) + ((x592x) & (!x21x) & (x11x) & (n_n5294) & (x208x)) + ((x592x) & (x21x) & (!x11x) & (!n_n5294) & (!x208x)) + ((x592x) & (x21x) & (!x11x) & (!n_n5294) & (x208x)) + ((x592x) & (x21x) & (!x11x) & (n_n5294) & (!x208x)) + ((x592x) & (x21x) & (!x11x) & (n_n5294) & (x208x)) + ((x592x) & (x21x) & (x11x) & (!n_n5294) & (!x208x)) + ((x592x) & (x21x) & (x11x) & (!n_n5294) & (x208x)) + ((x592x) & (x21x) & (x11x) & (n_n5294) & (!x208x)) + ((x592x) & (x21x) & (x11x) & (n_n5294) & (x208x)));
	assign x332x = (((n_n482) & (!n_n522) & (n_n130) & (!x12x) & (x20x)) + ((n_n482) & (!n_n522) & (n_n130) & (x12x) & (x20x)) + ((n_n482) & (n_n522) & (!n_n130) & (x12x) & (!x20x)) + ((n_n482) & (n_n522) & (!n_n130) & (x12x) & (x20x)) + ((n_n482) & (n_n522) & (n_n130) & (!x12x) & (x20x)) + ((n_n482) & (n_n522) & (n_n130) & (x12x) & (!x20x)) + ((n_n482) & (n_n522) & (n_n130) & (x12x) & (x20x)));
	assign n_n5080 = (((i_7_) & (i_8_) & (i_6_) & (n_n535) & (x12x)));
	assign x13306x = (((!i_9_) & (n_n526) & (n_n535) & (!n_n130) & (x12x)) + ((!i_9_) & (n_n526) & (n_n535) & (n_n130) & (!x12x)) + ((!i_9_) & (n_n526) & (n_n535) & (n_n130) & (x12x)) + ((i_9_) & (n_n526) & (n_n535) & (!n_n130) & (x12x)) + ((i_9_) & (n_n526) & (n_n535) & (n_n130) & (x12x)));
	assign x410x = (((!i_9_) & (n_n536) & (n_n518) & (!n_n532) & (n_n534)) + ((!i_9_) & (n_n536) & (n_n518) & (n_n532) & (n_n534)) + ((i_9_) & (n_n536) & (n_n518) & (n_n532) & (!n_n534)) + ((i_9_) & (n_n536) & (n_n518) & (n_n532) & (n_n534)));
	assign n_n5219 = (((!i_9_) & (n_n524) & (n_n535) & (n_n65)));
	assign n_n1521 = (((!x19x) & (!n_n520) & (!n_n500) & (!n_n5272) & (n_n5271)) + ((!x19x) & (!n_n520) & (!n_n500) & (n_n5272) & (!n_n5271)) + ((!x19x) & (!n_n520) & (!n_n500) & (n_n5272) & (n_n5271)) + ((!x19x) & (!n_n520) & (n_n500) & (!n_n5272) & (n_n5271)) + ((!x19x) & (!n_n520) & (n_n500) & (n_n5272) & (!n_n5271)) + ((!x19x) & (!n_n520) & (n_n500) & (n_n5272) & (n_n5271)) + ((!x19x) & (n_n520) & (!n_n500) & (!n_n5272) & (n_n5271)) + ((!x19x) & (n_n520) & (!n_n500) & (n_n5272) & (!n_n5271)) + ((!x19x) & (n_n520) & (!n_n500) & (n_n5272) & (n_n5271)) + ((!x19x) & (n_n520) & (n_n500) & (!n_n5272) & (n_n5271)) + ((!x19x) & (n_n520) & (n_n500) & (n_n5272) & (!n_n5271)) + ((!x19x) & (n_n520) & (n_n500) & (n_n5272) & (n_n5271)) + ((x19x) & (!n_n520) & (!n_n500) & (!n_n5272) & (n_n5271)) + ((x19x) & (!n_n520) & (!n_n500) & (n_n5272) & (!n_n5271)) + ((x19x) & (!n_n520) & (!n_n500) & (n_n5272) & (n_n5271)) + ((x19x) & (!n_n520) & (n_n500) & (!n_n5272) & (n_n5271)) + ((x19x) & (!n_n520) & (n_n500) & (n_n5272) & (!n_n5271)) + ((x19x) & (!n_n520) & (n_n500) & (n_n5272) & (n_n5271)) + ((x19x) & (n_n520) & (!n_n500) & (!n_n5272) & (n_n5271)) + ((x19x) & (n_n520) & (!n_n500) & (n_n5272) & (!n_n5271)) + ((x19x) & (n_n520) & (!n_n500) & (n_n5272) & (n_n5271)) + ((x19x) & (n_n520) & (n_n500) & (!n_n5272) & (!n_n5271)) + ((x19x) & (n_n520) & (n_n500) & (!n_n5272) & (n_n5271)) + ((x19x) & (n_n520) & (n_n500) & (n_n5272) & (!n_n5271)) + ((x19x) & (n_n520) & (n_n500) & (n_n5272) & (n_n5271)));
	assign n_n4529 = (((!i_9_) & (n_n526) & (n_n482) & (n_n455)));
	assign x328x = (((!i_9_) & (n_n536) & (n_n473) & (n_n530)) + ((i_9_) & (n_n536) & (n_n473) & (n_n530)));
	assign x22151x = (((!n_n4403) & (!n_n4407) & (!n_n4406) & (!n_n4408)));
	assign n_n1115 = (((!n_n4415) & (!n_n4404) & (!n_n4411) & (!x328x) & (!x22151x)) + ((!n_n4415) & (!n_n4404) & (!n_n4411) & (x328x) & (!x22151x)) + ((!n_n4415) & (!n_n4404) & (!n_n4411) & (x328x) & (x22151x)) + ((!n_n4415) & (!n_n4404) & (n_n4411) & (!x328x) & (!x22151x)) + ((!n_n4415) & (!n_n4404) & (n_n4411) & (!x328x) & (x22151x)) + ((!n_n4415) & (!n_n4404) & (n_n4411) & (x328x) & (!x22151x)) + ((!n_n4415) & (!n_n4404) & (n_n4411) & (x328x) & (x22151x)) + ((!n_n4415) & (n_n4404) & (!n_n4411) & (!x328x) & (!x22151x)) + ((!n_n4415) & (n_n4404) & (!n_n4411) & (!x328x) & (x22151x)) + ((!n_n4415) & (n_n4404) & (!n_n4411) & (x328x) & (!x22151x)) + ((!n_n4415) & (n_n4404) & (!n_n4411) & (x328x) & (x22151x)) + ((!n_n4415) & (n_n4404) & (n_n4411) & (!x328x) & (!x22151x)) + ((!n_n4415) & (n_n4404) & (n_n4411) & (!x328x) & (x22151x)) + ((!n_n4415) & (n_n4404) & (n_n4411) & (x328x) & (!x22151x)) + ((!n_n4415) & (n_n4404) & (n_n4411) & (x328x) & (x22151x)) + ((n_n4415) & (!n_n4404) & (!n_n4411) & (!x328x) & (!x22151x)) + ((n_n4415) & (!n_n4404) & (!n_n4411) & (!x328x) & (x22151x)) + ((n_n4415) & (!n_n4404) & (!n_n4411) & (x328x) & (!x22151x)) + ((n_n4415) & (!n_n4404) & (!n_n4411) & (x328x) & (x22151x)) + ((n_n4415) & (!n_n4404) & (n_n4411) & (!x328x) & (!x22151x)) + ((n_n4415) & (!n_n4404) & (n_n4411) & (!x328x) & (x22151x)) + ((n_n4415) & (!n_n4404) & (n_n4411) & (x328x) & (!x22151x)) + ((n_n4415) & (!n_n4404) & (n_n4411) & (x328x) & (x22151x)) + ((n_n4415) & (n_n4404) & (!n_n4411) & (!x328x) & (!x22151x)) + ((n_n4415) & (n_n4404) & (!n_n4411) & (!x328x) & (x22151x)) + ((n_n4415) & (n_n4404) & (!n_n4411) & (x328x) & (!x22151x)) + ((n_n4415) & (n_n4404) & (!n_n4411) & (x328x) & (x22151x)) + ((n_n4415) & (n_n4404) & (n_n4411) & (!x328x) & (!x22151x)) + ((n_n4415) & (n_n4404) & (n_n4411) & (!x328x) & (x22151x)) + ((n_n4415) & (n_n4404) & (n_n4411) & (x328x) & (!x22151x)) + ((n_n4415) & (n_n4404) & (n_n4411) & (x328x) & (x22151x)));
	assign x22161x = (((!n_n4547) & (!n_n4544) & (!n_n4543) & (!n_n4545)));
	assign n_n4692 = (((i_9_) & (n_n390) & (n_n522) & (n_n464)));
	assign x86x = (((!i_9_) & (!n_n534) & (!n_n325) & (!n_n535) & (n_n4695)) + ((!i_9_) & (!n_n534) & (!n_n325) & (n_n535) & (n_n4695)) + ((!i_9_) & (!n_n534) & (n_n325) & (!n_n535) & (n_n4695)) + ((!i_9_) & (!n_n534) & (n_n325) & (n_n535) & (n_n4695)) + ((!i_9_) & (n_n534) & (!n_n325) & (!n_n535) & (n_n4695)) + ((!i_9_) & (n_n534) & (!n_n325) & (n_n535) & (n_n4695)) + ((!i_9_) & (n_n534) & (n_n325) & (!n_n535) & (n_n4695)) + ((!i_9_) & (n_n534) & (n_n325) & (n_n535) & (n_n4695)) + ((i_9_) & (!n_n534) & (!n_n325) & (!n_n535) & (n_n4695)) + ((i_9_) & (!n_n534) & (!n_n325) & (n_n535) & (n_n4695)) + ((i_9_) & (!n_n534) & (n_n325) & (!n_n535) & (n_n4695)) + ((i_9_) & (!n_n534) & (n_n325) & (n_n535) & (n_n4695)) + ((i_9_) & (n_n534) & (!n_n325) & (!n_n535) & (n_n4695)) + ((i_9_) & (n_n534) & (!n_n325) & (n_n535) & (n_n4695)) + ((i_9_) & (n_n534) & (n_n325) & (!n_n535) & (n_n4695)) + ((i_9_) & (n_n534) & (n_n325) & (n_n535) & (!n_n4695)) + ((i_9_) & (n_n534) & (n_n325) & (n_n535) & (n_n4695)));
	assign x219x = (((!i_9_) & (!n_n528) & (n_n390) & (n_n530) & (n_n464)) + ((!i_9_) & (n_n528) & (n_n390) & (n_n530) & (n_n464)) + ((i_9_) & (n_n528) & (n_n390) & (!n_n530) & (n_n464)) + ((i_9_) & (n_n528) & (n_n390) & (n_n530) & (n_n464)));
	assign n_n1093 = (((!n_n4683) & (!n_n3849) & (!n_n4692) & (!x86x) & (x219x)) + ((!n_n4683) & (!n_n3849) & (!n_n4692) & (x86x) & (!x219x)) + ((!n_n4683) & (!n_n3849) & (!n_n4692) & (x86x) & (x219x)) + ((!n_n4683) & (!n_n3849) & (n_n4692) & (!x86x) & (!x219x)) + ((!n_n4683) & (!n_n3849) & (n_n4692) & (!x86x) & (x219x)) + ((!n_n4683) & (!n_n3849) & (n_n4692) & (x86x) & (!x219x)) + ((!n_n4683) & (!n_n3849) & (n_n4692) & (x86x) & (x219x)) + ((!n_n4683) & (n_n3849) & (!n_n4692) & (!x86x) & (!x219x)) + ((!n_n4683) & (n_n3849) & (!n_n4692) & (!x86x) & (x219x)) + ((!n_n4683) & (n_n3849) & (!n_n4692) & (x86x) & (!x219x)) + ((!n_n4683) & (n_n3849) & (!n_n4692) & (x86x) & (x219x)) + ((!n_n4683) & (n_n3849) & (n_n4692) & (!x86x) & (!x219x)) + ((!n_n4683) & (n_n3849) & (n_n4692) & (!x86x) & (x219x)) + ((!n_n4683) & (n_n3849) & (n_n4692) & (x86x) & (!x219x)) + ((!n_n4683) & (n_n3849) & (n_n4692) & (x86x) & (x219x)) + ((n_n4683) & (!n_n3849) & (!n_n4692) & (!x86x) & (!x219x)) + ((n_n4683) & (!n_n3849) & (!n_n4692) & (!x86x) & (x219x)) + ((n_n4683) & (!n_n3849) & (!n_n4692) & (x86x) & (!x219x)) + ((n_n4683) & (!n_n3849) & (!n_n4692) & (x86x) & (x219x)) + ((n_n4683) & (!n_n3849) & (n_n4692) & (!x86x) & (!x219x)) + ((n_n4683) & (!n_n3849) & (n_n4692) & (!x86x) & (x219x)) + ((n_n4683) & (!n_n3849) & (n_n4692) & (x86x) & (!x219x)) + ((n_n4683) & (!n_n3849) & (n_n4692) & (x86x) & (x219x)) + ((n_n4683) & (n_n3849) & (!n_n4692) & (!x86x) & (!x219x)) + ((n_n4683) & (n_n3849) & (!n_n4692) & (!x86x) & (x219x)) + ((n_n4683) & (n_n3849) & (!n_n4692) & (x86x) & (!x219x)) + ((n_n4683) & (n_n3849) & (!n_n4692) & (x86x) & (x219x)) + ((n_n4683) & (n_n3849) & (n_n4692) & (!x86x) & (!x219x)) + ((n_n4683) & (n_n3849) & (n_n4692) & (!x86x) & (x219x)) + ((n_n4683) & (n_n3849) & (n_n4692) & (x86x) & (!x219x)) + ((n_n4683) & (n_n3849) & (n_n4692) & (x86x) & (x219x)));
	assign x299x = (((!i_9_) & (n_n195) & (n_n500) & (n_n530)) + ((i_9_) & (n_n195) & (n_n500) & (n_n530)));
	assign x11980x = (((!i_9_) & (!n_n528) & (n_n534) & (n_n195) & (n_n500)) + ((!i_9_) & (n_n528) & (n_n534) & (n_n195) & (n_n500)) + ((i_9_) & (!n_n528) & (n_n534) & (n_n195) & (n_n500)) + ((i_9_) & (n_n528) & (!n_n534) & (n_n195) & (n_n500)) + ((i_9_) & (n_n528) & (n_n534) & (n_n195) & (n_n500)));
	assign n_n1068 = (((!n_n4994) & (!n_n5003) & (!x248x) & (!x299x) & (x11980x)) + ((!n_n4994) & (!n_n5003) & (!x248x) & (x299x) & (!x11980x)) + ((!n_n4994) & (!n_n5003) & (!x248x) & (x299x) & (x11980x)) + ((!n_n4994) & (!n_n5003) & (x248x) & (!x299x) & (!x11980x)) + ((!n_n4994) & (!n_n5003) & (x248x) & (!x299x) & (x11980x)) + ((!n_n4994) & (!n_n5003) & (x248x) & (x299x) & (!x11980x)) + ((!n_n4994) & (!n_n5003) & (x248x) & (x299x) & (x11980x)) + ((!n_n4994) & (n_n5003) & (!x248x) & (!x299x) & (!x11980x)) + ((!n_n4994) & (n_n5003) & (!x248x) & (!x299x) & (x11980x)) + ((!n_n4994) & (n_n5003) & (!x248x) & (x299x) & (!x11980x)) + ((!n_n4994) & (n_n5003) & (!x248x) & (x299x) & (x11980x)) + ((!n_n4994) & (n_n5003) & (x248x) & (!x299x) & (!x11980x)) + ((!n_n4994) & (n_n5003) & (x248x) & (!x299x) & (x11980x)) + ((!n_n4994) & (n_n5003) & (x248x) & (x299x) & (!x11980x)) + ((!n_n4994) & (n_n5003) & (x248x) & (x299x) & (x11980x)) + ((n_n4994) & (!n_n5003) & (!x248x) & (!x299x) & (!x11980x)) + ((n_n4994) & (!n_n5003) & (!x248x) & (!x299x) & (x11980x)) + ((n_n4994) & (!n_n5003) & (!x248x) & (x299x) & (!x11980x)) + ((n_n4994) & (!n_n5003) & (!x248x) & (x299x) & (x11980x)) + ((n_n4994) & (!n_n5003) & (x248x) & (!x299x) & (!x11980x)) + ((n_n4994) & (!n_n5003) & (x248x) & (!x299x) & (x11980x)) + ((n_n4994) & (!n_n5003) & (x248x) & (x299x) & (!x11980x)) + ((n_n4994) & (!n_n5003) & (x248x) & (x299x) & (x11980x)) + ((n_n4994) & (n_n5003) & (!x248x) & (!x299x) & (!x11980x)) + ((n_n4994) & (n_n5003) & (!x248x) & (!x299x) & (x11980x)) + ((n_n4994) & (n_n5003) & (!x248x) & (x299x) & (!x11980x)) + ((n_n4994) & (n_n5003) & (!x248x) & (x299x) & (x11980x)) + ((n_n4994) & (n_n5003) & (x248x) & (!x299x) & (!x11980x)) + ((n_n4994) & (n_n5003) & (x248x) & (!x299x) & (x11980x)) + ((n_n4994) & (n_n5003) & (x248x) & (x299x) & (!x11980x)) + ((n_n4994) & (n_n5003) & (x248x) & (x299x) & (x11980x)));
	assign x62x = (((!i_9_) & (!x19x) & (n_n532) & (n_n500) & (n_n65)) + ((!i_9_) & (x19x) & (n_n532) & (n_n500) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n532) & (n_n500) & (n_n65)) + ((i_9_) & (x19x) & (n_n532) & (n_n500) & (!n_n65)) + ((i_9_) & (x19x) & (n_n532) & (n_n500) & (n_n65)));
	assign x409x = (((!i_9_) & (!x19x) & (n_n500) & (n_n530) & (n_n65)) + ((!i_9_) & (x19x) & (n_n500) & (n_n530) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n500) & (n_n530) & (n_n65)) + ((i_9_) & (x19x) & (n_n500) & (n_n530) & (!n_n65)) + ((i_9_) & (x19x) & (n_n500) & (n_n530) & (n_n65)));
	assign x11925x = (((!x11x) & (!x24x) & (!n_n500) & (!n_n65) & (n_n5258)) + ((!x11x) & (!x24x) & (!n_n500) & (n_n65) & (n_n5258)) + ((!x11x) & (!x24x) & (n_n500) & (!n_n65) & (n_n5258)) + ((!x11x) & (!x24x) & (n_n500) & (n_n65) & (n_n5258)) + ((!x11x) & (x24x) & (!n_n500) & (!n_n65) & (n_n5258)) + ((!x11x) & (x24x) & (!n_n500) & (n_n65) & (n_n5258)) + ((!x11x) & (x24x) & (n_n500) & (!n_n65) & (n_n5258)) + ((!x11x) & (x24x) & (n_n500) & (n_n65) & (!n_n5258)) + ((!x11x) & (x24x) & (n_n500) & (n_n65) & (n_n5258)) + ((x11x) & (!x24x) & (!n_n500) & (!n_n65) & (n_n5258)) + ((x11x) & (!x24x) & (!n_n500) & (n_n65) & (n_n5258)) + ((x11x) & (!x24x) & (n_n500) & (!n_n65) & (n_n5258)) + ((x11x) & (!x24x) & (n_n500) & (n_n65) & (!n_n5258)) + ((x11x) & (!x24x) & (n_n500) & (n_n65) & (n_n5258)) + ((x11x) & (x24x) & (!n_n500) & (!n_n65) & (n_n5258)) + ((x11x) & (x24x) & (!n_n500) & (n_n65) & (n_n5258)) + ((x11x) & (x24x) & (n_n500) & (!n_n65) & (n_n5258)) + ((x11x) & (x24x) & (n_n500) & (n_n65) & (!n_n5258)) + ((x11x) & (x24x) & (n_n500) & (n_n65) & (n_n5258)));
	assign x22193x = (((!x20x) & (!n_n500) & (!n_n65) & (!n_n5266) & (!n_n5264)) + ((!x20x) & (!n_n500) & (n_n65) & (!n_n5266) & (!n_n5264)) + ((!x20x) & (n_n500) & (!n_n65) & (!n_n5266) & (!n_n5264)) + ((!x20x) & (n_n500) & (n_n65) & (!n_n5266) & (!n_n5264)) + ((x20x) & (!n_n500) & (!n_n65) & (!n_n5266) & (!n_n5264)) + ((x20x) & (!n_n500) & (n_n65) & (!n_n5266) & (!n_n5264)) + ((x20x) & (n_n500) & (!n_n65) & (!n_n5266) & (!n_n5264)));
	assign n_n1049 = (((!n_n5261) & (!n_n5260) & (!n_n5257) & (!x11925x) & (!x22193x)) + ((!n_n5261) & (!n_n5260) & (!n_n5257) & (x11925x) & (!x22193x)) + ((!n_n5261) & (!n_n5260) & (!n_n5257) & (x11925x) & (x22193x)) + ((!n_n5261) & (!n_n5260) & (n_n5257) & (!x11925x) & (!x22193x)) + ((!n_n5261) & (!n_n5260) & (n_n5257) & (!x11925x) & (x22193x)) + ((!n_n5261) & (!n_n5260) & (n_n5257) & (x11925x) & (!x22193x)) + ((!n_n5261) & (!n_n5260) & (n_n5257) & (x11925x) & (x22193x)) + ((!n_n5261) & (n_n5260) & (!n_n5257) & (!x11925x) & (!x22193x)) + ((!n_n5261) & (n_n5260) & (!n_n5257) & (!x11925x) & (x22193x)) + ((!n_n5261) & (n_n5260) & (!n_n5257) & (x11925x) & (!x22193x)) + ((!n_n5261) & (n_n5260) & (!n_n5257) & (x11925x) & (x22193x)) + ((!n_n5261) & (n_n5260) & (n_n5257) & (!x11925x) & (!x22193x)) + ((!n_n5261) & (n_n5260) & (n_n5257) & (!x11925x) & (x22193x)) + ((!n_n5261) & (n_n5260) & (n_n5257) & (x11925x) & (!x22193x)) + ((!n_n5261) & (n_n5260) & (n_n5257) & (x11925x) & (x22193x)) + ((n_n5261) & (!n_n5260) & (!n_n5257) & (!x11925x) & (!x22193x)) + ((n_n5261) & (!n_n5260) & (!n_n5257) & (!x11925x) & (x22193x)) + ((n_n5261) & (!n_n5260) & (!n_n5257) & (x11925x) & (!x22193x)) + ((n_n5261) & (!n_n5260) & (!n_n5257) & (x11925x) & (x22193x)) + ((n_n5261) & (!n_n5260) & (n_n5257) & (!x11925x) & (!x22193x)) + ((n_n5261) & (!n_n5260) & (n_n5257) & (!x11925x) & (x22193x)) + ((n_n5261) & (!n_n5260) & (n_n5257) & (x11925x) & (!x22193x)) + ((n_n5261) & (!n_n5260) & (n_n5257) & (x11925x) & (x22193x)) + ((n_n5261) & (n_n5260) & (!n_n5257) & (!x11925x) & (!x22193x)) + ((n_n5261) & (n_n5260) & (!n_n5257) & (!x11925x) & (x22193x)) + ((n_n5261) & (n_n5260) & (!n_n5257) & (x11925x) & (!x22193x)) + ((n_n5261) & (n_n5260) & (!n_n5257) & (x11925x) & (x22193x)) + ((n_n5261) & (n_n5260) & (n_n5257) & (!x11925x) & (!x22193x)) + ((n_n5261) & (n_n5260) & (n_n5257) & (!x11925x) & (x22193x)) + ((n_n5261) & (n_n5260) & (n_n5257) & (x11925x) & (!x22193x)) + ((n_n5261) & (n_n5260) & (n_n5257) & (x11925x) & (x22193x)));
	assign n_n1047 = (((!n_n5287) & (!x441x) & (!x207x) & (!n_n5283) & (n_n2651)) + ((!n_n5287) & (!x441x) & (!x207x) & (n_n5283) & (!n_n2651)) + ((!n_n5287) & (!x441x) & (!x207x) & (n_n5283) & (n_n2651)) + ((!n_n5287) & (!x441x) & (x207x) & (!n_n5283) & (!n_n2651)) + ((!n_n5287) & (!x441x) & (x207x) & (!n_n5283) & (n_n2651)) + ((!n_n5287) & (!x441x) & (x207x) & (n_n5283) & (!n_n2651)) + ((!n_n5287) & (!x441x) & (x207x) & (n_n5283) & (n_n2651)) + ((!n_n5287) & (x441x) & (!x207x) & (!n_n5283) & (!n_n2651)) + ((!n_n5287) & (x441x) & (!x207x) & (!n_n5283) & (n_n2651)) + ((!n_n5287) & (x441x) & (!x207x) & (n_n5283) & (!n_n2651)) + ((!n_n5287) & (x441x) & (!x207x) & (n_n5283) & (n_n2651)) + ((!n_n5287) & (x441x) & (x207x) & (!n_n5283) & (!n_n2651)) + ((!n_n5287) & (x441x) & (x207x) & (!n_n5283) & (n_n2651)) + ((!n_n5287) & (x441x) & (x207x) & (n_n5283) & (!n_n2651)) + ((!n_n5287) & (x441x) & (x207x) & (n_n5283) & (n_n2651)) + ((n_n5287) & (!x441x) & (!x207x) & (!n_n5283) & (!n_n2651)) + ((n_n5287) & (!x441x) & (!x207x) & (!n_n5283) & (n_n2651)) + ((n_n5287) & (!x441x) & (!x207x) & (n_n5283) & (!n_n2651)) + ((n_n5287) & (!x441x) & (!x207x) & (n_n5283) & (n_n2651)) + ((n_n5287) & (!x441x) & (x207x) & (!n_n5283) & (!n_n2651)) + ((n_n5287) & (!x441x) & (x207x) & (!n_n5283) & (n_n2651)) + ((n_n5287) & (!x441x) & (x207x) & (n_n5283) & (!n_n2651)) + ((n_n5287) & (!x441x) & (x207x) & (n_n5283) & (n_n2651)) + ((n_n5287) & (x441x) & (!x207x) & (!n_n5283) & (!n_n2651)) + ((n_n5287) & (x441x) & (!x207x) & (!n_n5283) & (n_n2651)) + ((n_n5287) & (x441x) & (!x207x) & (n_n5283) & (!n_n2651)) + ((n_n5287) & (x441x) & (!x207x) & (n_n5283) & (n_n2651)) + ((n_n5287) & (x441x) & (x207x) & (!n_n5283) & (!n_n2651)) + ((n_n5287) & (x441x) & (x207x) & (!n_n5283) & (n_n2651)) + ((n_n5287) & (x441x) & (x207x) & (n_n5283) & (!n_n2651)) + ((n_n5287) & (x441x) & (x207x) & (n_n5283) & (n_n2651)));
	assign n_n1048 = (((!n_n5273) & (!n_n5278) & (!n_n1521) & (!x438x) & (x333x)) + ((!n_n5273) & (!n_n5278) & (!n_n1521) & (x438x) & (!x333x)) + ((!n_n5273) & (!n_n5278) & (!n_n1521) & (x438x) & (x333x)) + ((!n_n5273) & (!n_n5278) & (n_n1521) & (!x438x) & (!x333x)) + ((!n_n5273) & (!n_n5278) & (n_n1521) & (!x438x) & (x333x)) + ((!n_n5273) & (!n_n5278) & (n_n1521) & (x438x) & (!x333x)) + ((!n_n5273) & (!n_n5278) & (n_n1521) & (x438x) & (x333x)) + ((!n_n5273) & (n_n5278) & (!n_n1521) & (!x438x) & (!x333x)) + ((!n_n5273) & (n_n5278) & (!n_n1521) & (!x438x) & (x333x)) + ((!n_n5273) & (n_n5278) & (!n_n1521) & (x438x) & (!x333x)) + ((!n_n5273) & (n_n5278) & (!n_n1521) & (x438x) & (x333x)) + ((!n_n5273) & (n_n5278) & (n_n1521) & (!x438x) & (!x333x)) + ((!n_n5273) & (n_n5278) & (n_n1521) & (!x438x) & (x333x)) + ((!n_n5273) & (n_n5278) & (n_n1521) & (x438x) & (!x333x)) + ((!n_n5273) & (n_n5278) & (n_n1521) & (x438x) & (x333x)) + ((n_n5273) & (!n_n5278) & (!n_n1521) & (!x438x) & (!x333x)) + ((n_n5273) & (!n_n5278) & (!n_n1521) & (!x438x) & (x333x)) + ((n_n5273) & (!n_n5278) & (!n_n1521) & (x438x) & (!x333x)) + ((n_n5273) & (!n_n5278) & (!n_n1521) & (x438x) & (x333x)) + ((n_n5273) & (!n_n5278) & (n_n1521) & (!x438x) & (!x333x)) + ((n_n5273) & (!n_n5278) & (n_n1521) & (!x438x) & (x333x)) + ((n_n5273) & (!n_n5278) & (n_n1521) & (x438x) & (!x333x)) + ((n_n5273) & (!n_n5278) & (n_n1521) & (x438x) & (x333x)) + ((n_n5273) & (n_n5278) & (!n_n1521) & (!x438x) & (!x333x)) + ((n_n5273) & (n_n5278) & (!n_n1521) & (!x438x) & (x333x)) + ((n_n5273) & (n_n5278) & (!n_n1521) & (x438x) & (!x333x)) + ((n_n5273) & (n_n5278) & (!n_n1521) & (x438x) & (x333x)) + ((n_n5273) & (n_n5278) & (n_n1521) & (!x438x) & (!x333x)) + ((n_n5273) & (n_n5278) & (n_n1521) & (!x438x) & (x333x)) + ((n_n5273) & (n_n5278) & (n_n1521) & (x438x) & (!x333x)) + ((n_n5273) & (n_n5278) & (n_n1521) & (x438x) & (x333x)));
	assign x200x = (((i_7_) & (!i_8_) & (!i_6_) & (x19x) & (n_n482)) + ((i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n482)));
	assign x22156x = (((!x592x) & (!n_n5293) & (!x24x) & (!n_n5294) & (!x63x)) + ((!x592x) & (!n_n5293) & (x24x) & (!n_n5294) & (!x63x)) + ((x592x) & (!n_n5293) & (!x24x) & (!n_n5294) & (!x63x)));
	assign x11940x = (((!x592x) & (!x21x) & (!n_n5290) & (!x200x) & (!x22156x)) + ((!x592x) & (!x21x) & (!n_n5290) & (x200x) & (!x22156x)) + ((!x592x) & (!x21x) & (!n_n5290) & (x200x) & (x22156x)) + ((!x592x) & (!x21x) & (n_n5290) & (!x200x) & (!x22156x)) + ((!x592x) & (!x21x) & (n_n5290) & (!x200x) & (x22156x)) + ((!x592x) & (!x21x) & (n_n5290) & (x200x) & (!x22156x)) + ((!x592x) & (!x21x) & (n_n5290) & (x200x) & (x22156x)) + ((!x592x) & (x21x) & (!n_n5290) & (!x200x) & (!x22156x)) + ((!x592x) & (x21x) & (!n_n5290) & (x200x) & (!x22156x)) + ((!x592x) & (x21x) & (!n_n5290) & (x200x) & (x22156x)) + ((!x592x) & (x21x) & (n_n5290) & (!x200x) & (!x22156x)) + ((!x592x) & (x21x) & (n_n5290) & (!x200x) & (x22156x)) + ((!x592x) & (x21x) & (n_n5290) & (x200x) & (!x22156x)) + ((!x592x) & (x21x) & (n_n5290) & (x200x) & (x22156x)) + ((x592x) & (!x21x) & (!n_n5290) & (!x200x) & (!x22156x)) + ((x592x) & (!x21x) & (!n_n5290) & (x200x) & (!x22156x)) + ((x592x) & (!x21x) & (!n_n5290) & (x200x) & (x22156x)) + ((x592x) & (!x21x) & (n_n5290) & (!x200x) & (!x22156x)) + ((x592x) & (!x21x) & (n_n5290) & (!x200x) & (x22156x)) + ((x592x) & (!x21x) & (n_n5290) & (x200x) & (!x22156x)) + ((x592x) & (!x21x) & (n_n5290) & (x200x) & (x22156x)) + ((x592x) & (x21x) & (!n_n5290) & (!x200x) & (!x22156x)) + ((x592x) & (x21x) & (!n_n5290) & (!x200x) & (x22156x)) + ((x592x) & (x21x) & (!n_n5290) & (x200x) & (!x22156x)) + ((x592x) & (x21x) & (!n_n5290) & (x200x) & (x22156x)) + ((x592x) & (x21x) & (n_n5290) & (!x200x) & (!x22156x)) + ((x592x) & (x21x) & (n_n5290) & (!x200x) & (x22156x)) + ((x592x) & (x21x) & (n_n5290) & (x200x) & (!x22156x)) + ((x592x) & (x21x) & (n_n5290) & (x200x) & (x22156x)));
	assign n_n1017 = (((!n_n1047) & (!n_n1048) & (x11940x)) + ((!n_n1047) & (n_n1048) & (!x11940x)) + ((!n_n1047) & (n_n1048) & (x11940x)) + ((n_n1047) & (!n_n1048) & (!x11940x)) + ((n_n1047) & (!n_n1048) & (x11940x)) + ((n_n1047) & (n_n1048) & (!x11940x)) + ((n_n1047) & (n_n1048) & (x11940x)));
	assign n_n1045 = (((!x459x) & (!n_n5311) & (!n_n5303) & (!n_n1128) & (x325x)) + ((!x459x) & (!n_n5311) & (!n_n5303) & (n_n1128) & (!x325x)) + ((!x459x) & (!n_n5311) & (!n_n5303) & (n_n1128) & (x325x)) + ((!x459x) & (!n_n5311) & (n_n5303) & (!n_n1128) & (!x325x)) + ((!x459x) & (!n_n5311) & (n_n5303) & (!n_n1128) & (x325x)) + ((!x459x) & (!n_n5311) & (n_n5303) & (n_n1128) & (!x325x)) + ((!x459x) & (!n_n5311) & (n_n5303) & (n_n1128) & (x325x)) + ((!x459x) & (n_n5311) & (!n_n5303) & (!n_n1128) & (!x325x)) + ((!x459x) & (n_n5311) & (!n_n5303) & (!n_n1128) & (x325x)) + ((!x459x) & (n_n5311) & (!n_n5303) & (n_n1128) & (!x325x)) + ((!x459x) & (n_n5311) & (!n_n5303) & (n_n1128) & (x325x)) + ((!x459x) & (n_n5311) & (n_n5303) & (!n_n1128) & (!x325x)) + ((!x459x) & (n_n5311) & (n_n5303) & (!n_n1128) & (x325x)) + ((!x459x) & (n_n5311) & (n_n5303) & (n_n1128) & (!x325x)) + ((!x459x) & (n_n5311) & (n_n5303) & (n_n1128) & (x325x)) + ((x459x) & (!n_n5311) & (!n_n5303) & (!n_n1128) & (!x325x)) + ((x459x) & (!n_n5311) & (!n_n5303) & (!n_n1128) & (x325x)) + ((x459x) & (!n_n5311) & (!n_n5303) & (n_n1128) & (!x325x)) + ((x459x) & (!n_n5311) & (!n_n5303) & (n_n1128) & (x325x)) + ((x459x) & (!n_n5311) & (n_n5303) & (!n_n1128) & (!x325x)) + ((x459x) & (!n_n5311) & (n_n5303) & (!n_n1128) & (x325x)) + ((x459x) & (!n_n5311) & (n_n5303) & (n_n1128) & (!x325x)) + ((x459x) & (!n_n5311) & (n_n5303) & (n_n1128) & (x325x)) + ((x459x) & (n_n5311) & (!n_n5303) & (!n_n1128) & (!x325x)) + ((x459x) & (n_n5311) & (!n_n5303) & (!n_n1128) & (x325x)) + ((x459x) & (n_n5311) & (!n_n5303) & (n_n1128) & (!x325x)) + ((x459x) & (n_n5311) & (!n_n5303) & (n_n1128) & (x325x)) + ((x459x) & (n_n5311) & (n_n5303) & (!n_n1128) & (!x325x)) + ((x459x) & (n_n5311) & (n_n5303) & (!n_n1128) & (x325x)) + ((x459x) & (n_n5311) & (n_n5303) & (n_n1128) & (!x325x)) + ((x459x) & (n_n5311) & (n_n5303) & (n_n1128) & (x325x)));
	assign n_n1900 = (((!i_9_) & (!n_n532) & (n_n534) & (n_n464) & (n_n65)) + ((!i_9_) & (n_n532) & (!n_n534) & (n_n464) & (n_n65)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n464) & (n_n65)) + ((i_9_) & (n_n532) & (!n_n534) & (n_n464) & (n_n65)) + ((i_9_) & (n_n532) & (n_n534) & (n_n464) & (n_n65)));
	assign x175x = (((!i_9_) & (!x19x) & (n_n530) & (n_n464) & (n_n65)) + ((!i_9_) & (x19x) & (n_n530) & (n_n464) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n530) & (n_n464) & (n_n65)) + ((i_9_) & (x19x) & (n_n530) & (n_n464) & (!n_n65)) + ((i_9_) & (x19x) & (n_n530) & (n_n464) & (n_n65)));
	assign x11950x = (((!i_9_) & (!n_n528) & (!n_n464) & (!n_n65) & (x175x)) + ((!i_9_) & (!n_n528) & (!n_n464) & (n_n65) & (x175x)) + ((!i_9_) & (!n_n528) & (n_n464) & (!n_n65) & (x175x)) + ((!i_9_) & (!n_n528) & (n_n464) & (n_n65) & (x175x)) + ((!i_9_) & (n_n528) & (!n_n464) & (!n_n65) & (x175x)) + ((!i_9_) & (n_n528) & (!n_n464) & (n_n65) & (x175x)) + ((!i_9_) & (n_n528) & (n_n464) & (!n_n65) & (x175x)) + ((!i_9_) & (n_n528) & (n_n464) & (n_n65) & (!x175x)) + ((!i_9_) & (n_n528) & (n_n464) & (n_n65) & (x175x)) + ((i_9_) & (!n_n528) & (!n_n464) & (!n_n65) & (x175x)) + ((i_9_) & (!n_n528) & (!n_n464) & (n_n65) & (x175x)) + ((i_9_) & (!n_n528) & (n_n464) & (!n_n65) & (x175x)) + ((i_9_) & (!n_n528) & (n_n464) & (n_n65) & (x175x)) + ((i_9_) & (n_n528) & (!n_n464) & (!n_n65) & (x175x)) + ((i_9_) & (n_n528) & (!n_n464) & (n_n65) & (x175x)) + ((i_9_) & (n_n528) & (n_n464) & (!n_n65) & (x175x)) + ((i_9_) & (n_n528) & (n_n464) & (n_n65) & (!x175x)) + ((i_9_) & (n_n528) & (n_n464) & (n_n65) & (x175x)));
	assign x22189x = (((!x19x) & (!n_n5331) & (!x516x) & (!n_n5319) & (!n_n5333)) + ((!x19x) & (!n_n5331) & (x516x) & (!n_n5319) & (!n_n5333)) + ((x19x) & (!n_n5331) & (!x516x) & (!n_n5319) & (!n_n5333)));
	assign x11953x = (((!n_n1900) & (!x115x) & (!x11950x) & (!x22189x)) + ((!n_n1900) & (!x115x) & (x11950x) & (!x22189x)) + ((!n_n1900) & (!x115x) & (x11950x) & (x22189x)) + ((!n_n1900) & (x115x) & (!x11950x) & (!x22189x)) + ((!n_n1900) & (x115x) & (!x11950x) & (x22189x)) + ((!n_n1900) & (x115x) & (x11950x) & (!x22189x)) + ((!n_n1900) & (x115x) & (x11950x) & (x22189x)) + ((n_n1900) & (!x115x) & (!x11950x) & (!x22189x)) + ((n_n1900) & (!x115x) & (!x11950x) & (x22189x)) + ((n_n1900) & (!x115x) & (x11950x) & (!x22189x)) + ((n_n1900) & (!x115x) & (x11950x) & (x22189x)) + ((n_n1900) & (x115x) & (!x11950x) & (!x22189x)) + ((n_n1900) & (x115x) & (!x11950x) & (x22189x)) + ((n_n1900) & (x115x) & (x11950x) & (!x22189x)) + ((n_n1900) & (x115x) & (x11950x) & (x22189x)));
	assign x11960x = (((!n_n5240) & (!n_n5238) & (!n_n5241) & (!n_n5243) & (x11959x)) + ((!n_n5240) & (!n_n5238) & (!n_n5241) & (n_n5243) & (!x11959x)) + ((!n_n5240) & (!n_n5238) & (!n_n5241) & (n_n5243) & (x11959x)) + ((!n_n5240) & (!n_n5238) & (n_n5241) & (!n_n5243) & (!x11959x)) + ((!n_n5240) & (!n_n5238) & (n_n5241) & (!n_n5243) & (x11959x)) + ((!n_n5240) & (!n_n5238) & (n_n5241) & (n_n5243) & (!x11959x)) + ((!n_n5240) & (!n_n5238) & (n_n5241) & (n_n5243) & (x11959x)) + ((!n_n5240) & (n_n5238) & (!n_n5241) & (!n_n5243) & (!x11959x)) + ((!n_n5240) & (n_n5238) & (!n_n5241) & (!n_n5243) & (x11959x)) + ((!n_n5240) & (n_n5238) & (!n_n5241) & (n_n5243) & (!x11959x)) + ((!n_n5240) & (n_n5238) & (!n_n5241) & (n_n5243) & (x11959x)) + ((!n_n5240) & (n_n5238) & (n_n5241) & (!n_n5243) & (!x11959x)) + ((!n_n5240) & (n_n5238) & (n_n5241) & (!n_n5243) & (x11959x)) + ((!n_n5240) & (n_n5238) & (n_n5241) & (n_n5243) & (!x11959x)) + ((!n_n5240) & (n_n5238) & (n_n5241) & (n_n5243) & (x11959x)) + ((n_n5240) & (!n_n5238) & (!n_n5241) & (!n_n5243) & (!x11959x)) + ((n_n5240) & (!n_n5238) & (!n_n5241) & (!n_n5243) & (x11959x)) + ((n_n5240) & (!n_n5238) & (!n_n5241) & (n_n5243) & (!x11959x)) + ((n_n5240) & (!n_n5238) & (!n_n5241) & (n_n5243) & (x11959x)) + ((n_n5240) & (!n_n5238) & (n_n5241) & (!n_n5243) & (!x11959x)) + ((n_n5240) & (!n_n5238) & (n_n5241) & (!n_n5243) & (x11959x)) + ((n_n5240) & (!n_n5238) & (n_n5241) & (n_n5243) & (!x11959x)) + ((n_n5240) & (!n_n5238) & (n_n5241) & (n_n5243) & (x11959x)) + ((n_n5240) & (n_n5238) & (!n_n5241) & (!n_n5243) & (!x11959x)) + ((n_n5240) & (n_n5238) & (!n_n5241) & (!n_n5243) & (x11959x)) + ((n_n5240) & (n_n5238) & (!n_n5241) & (n_n5243) & (!x11959x)) + ((n_n5240) & (n_n5238) & (!n_n5241) & (n_n5243) & (x11959x)) + ((n_n5240) & (n_n5238) & (n_n5241) & (!n_n5243) & (!x11959x)) + ((n_n5240) & (n_n5238) & (n_n5241) & (!n_n5243) & (x11959x)) + ((n_n5240) & (n_n5238) & (n_n5241) & (n_n5243) & (!x11959x)) + ((n_n5240) & (n_n5238) & (n_n5241) & (n_n5243) & (x11959x)));
	assign x11961x = (((!n_n5252) & (!n_n5250) & (!n_n1049) & (!x22192x)) + ((!n_n5252) & (!n_n5250) & (n_n1049) & (!x22192x)) + ((!n_n5252) & (!n_n5250) & (n_n1049) & (x22192x)) + ((!n_n5252) & (n_n5250) & (!n_n1049) & (!x22192x)) + ((!n_n5252) & (n_n5250) & (!n_n1049) & (x22192x)) + ((!n_n5252) & (n_n5250) & (n_n1049) & (!x22192x)) + ((!n_n5252) & (n_n5250) & (n_n1049) & (x22192x)) + ((n_n5252) & (!n_n5250) & (!n_n1049) & (!x22192x)) + ((n_n5252) & (!n_n5250) & (!n_n1049) & (x22192x)) + ((n_n5252) & (!n_n5250) & (n_n1049) & (!x22192x)) + ((n_n5252) & (!n_n5250) & (n_n1049) & (x22192x)) + ((n_n5252) & (n_n5250) & (!n_n1049) & (!x22192x)) + ((n_n5252) & (n_n5250) & (!n_n1049) & (x22192x)) + ((n_n5252) & (n_n5250) & (n_n1049) & (!x22192x)) + ((n_n5252) & (n_n5250) & (n_n1049) & (x22192x)));
	assign x12621x = (((!n_n4668) & (!n_n4670) & (!n_n4672) & (!n_n4692) & (n_n4686)) + ((!n_n4668) & (!n_n4670) & (!n_n4672) & (n_n4692) & (!n_n4686)) + ((!n_n4668) & (!n_n4670) & (!n_n4672) & (n_n4692) & (n_n4686)) + ((!n_n4668) & (!n_n4670) & (n_n4672) & (!n_n4692) & (!n_n4686)) + ((!n_n4668) & (!n_n4670) & (n_n4672) & (!n_n4692) & (n_n4686)) + ((!n_n4668) & (!n_n4670) & (n_n4672) & (n_n4692) & (!n_n4686)) + ((!n_n4668) & (!n_n4670) & (n_n4672) & (n_n4692) & (n_n4686)) + ((!n_n4668) & (n_n4670) & (!n_n4672) & (!n_n4692) & (!n_n4686)) + ((!n_n4668) & (n_n4670) & (!n_n4672) & (!n_n4692) & (n_n4686)) + ((!n_n4668) & (n_n4670) & (!n_n4672) & (n_n4692) & (!n_n4686)) + ((!n_n4668) & (n_n4670) & (!n_n4672) & (n_n4692) & (n_n4686)) + ((!n_n4668) & (n_n4670) & (n_n4672) & (!n_n4692) & (!n_n4686)) + ((!n_n4668) & (n_n4670) & (n_n4672) & (!n_n4692) & (n_n4686)) + ((!n_n4668) & (n_n4670) & (n_n4672) & (n_n4692) & (!n_n4686)) + ((!n_n4668) & (n_n4670) & (n_n4672) & (n_n4692) & (n_n4686)) + ((n_n4668) & (!n_n4670) & (!n_n4672) & (!n_n4692) & (!n_n4686)) + ((n_n4668) & (!n_n4670) & (!n_n4672) & (!n_n4692) & (n_n4686)) + ((n_n4668) & (!n_n4670) & (!n_n4672) & (n_n4692) & (!n_n4686)) + ((n_n4668) & (!n_n4670) & (!n_n4672) & (n_n4692) & (n_n4686)) + ((n_n4668) & (!n_n4670) & (n_n4672) & (!n_n4692) & (!n_n4686)) + ((n_n4668) & (!n_n4670) & (n_n4672) & (!n_n4692) & (n_n4686)) + ((n_n4668) & (!n_n4670) & (n_n4672) & (n_n4692) & (!n_n4686)) + ((n_n4668) & (!n_n4670) & (n_n4672) & (n_n4692) & (n_n4686)) + ((n_n4668) & (n_n4670) & (!n_n4672) & (!n_n4692) & (!n_n4686)) + ((n_n4668) & (n_n4670) & (!n_n4672) & (!n_n4692) & (n_n4686)) + ((n_n4668) & (n_n4670) & (!n_n4672) & (n_n4692) & (!n_n4686)) + ((n_n4668) & (n_n4670) & (!n_n4672) & (n_n4692) & (n_n4686)) + ((n_n4668) & (n_n4670) & (n_n4672) & (!n_n4692) & (!n_n4686)) + ((n_n4668) & (n_n4670) & (n_n4672) & (!n_n4692) & (n_n4686)) + ((n_n4668) & (n_n4670) & (n_n4672) & (n_n4692) & (!n_n4686)) + ((n_n4668) & (n_n4670) & (n_n4672) & (n_n4692) & (n_n4686)));
	assign x22136x = (((!n_n5258) & (!n_n5212) & (!n_n5266) & (!n_n5236)));
	assign n_n546 = (((!n_n5262) & (!n_n5235) & (!n_n5259) & (!x320x) & (!x22136x)) + ((!n_n5262) & (!n_n5235) & (!n_n5259) & (x320x) & (!x22136x)) + ((!n_n5262) & (!n_n5235) & (!n_n5259) & (x320x) & (x22136x)) + ((!n_n5262) & (!n_n5235) & (n_n5259) & (!x320x) & (!x22136x)) + ((!n_n5262) & (!n_n5235) & (n_n5259) & (!x320x) & (x22136x)) + ((!n_n5262) & (!n_n5235) & (n_n5259) & (x320x) & (!x22136x)) + ((!n_n5262) & (!n_n5235) & (n_n5259) & (x320x) & (x22136x)) + ((!n_n5262) & (n_n5235) & (!n_n5259) & (!x320x) & (!x22136x)) + ((!n_n5262) & (n_n5235) & (!n_n5259) & (!x320x) & (x22136x)) + ((!n_n5262) & (n_n5235) & (!n_n5259) & (x320x) & (!x22136x)) + ((!n_n5262) & (n_n5235) & (!n_n5259) & (x320x) & (x22136x)) + ((!n_n5262) & (n_n5235) & (n_n5259) & (!x320x) & (!x22136x)) + ((!n_n5262) & (n_n5235) & (n_n5259) & (!x320x) & (x22136x)) + ((!n_n5262) & (n_n5235) & (n_n5259) & (x320x) & (!x22136x)) + ((!n_n5262) & (n_n5235) & (n_n5259) & (x320x) & (x22136x)) + ((n_n5262) & (!n_n5235) & (!n_n5259) & (!x320x) & (!x22136x)) + ((n_n5262) & (!n_n5235) & (!n_n5259) & (!x320x) & (x22136x)) + ((n_n5262) & (!n_n5235) & (!n_n5259) & (x320x) & (!x22136x)) + ((n_n5262) & (!n_n5235) & (!n_n5259) & (x320x) & (x22136x)) + ((n_n5262) & (!n_n5235) & (n_n5259) & (!x320x) & (!x22136x)) + ((n_n5262) & (!n_n5235) & (n_n5259) & (!x320x) & (x22136x)) + ((n_n5262) & (!n_n5235) & (n_n5259) & (x320x) & (!x22136x)) + ((n_n5262) & (!n_n5235) & (n_n5259) & (x320x) & (x22136x)) + ((n_n5262) & (n_n5235) & (!n_n5259) & (!x320x) & (!x22136x)) + ((n_n5262) & (n_n5235) & (!n_n5259) & (!x320x) & (x22136x)) + ((n_n5262) & (n_n5235) & (!n_n5259) & (x320x) & (!x22136x)) + ((n_n5262) & (n_n5235) & (!n_n5259) & (x320x) & (x22136x)) + ((n_n5262) & (n_n5235) & (n_n5259) & (!x320x) & (!x22136x)) + ((n_n5262) & (n_n5235) & (n_n5259) & (!x320x) & (x22136x)) + ((n_n5262) & (n_n5235) & (n_n5259) & (x320x) & (!x22136x)) + ((n_n5262) & (n_n5235) & (n_n5259) & (x320x) & (x22136x)));
	assign n_n5210 = (((i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n535)));
	assign x13568x = (((!x268x) & (!n_n5313) & (!n_n5335) & (!n_n5334) & (x267x)) + ((!x268x) & (!n_n5313) & (!n_n5335) & (n_n5334) & (!x267x)) + ((!x268x) & (!n_n5313) & (!n_n5335) & (n_n5334) & (x267x)) + ((!x268x) & (!n_n5313) & (n_n5335) & (!n_n5334) & (!x267x)) + ((!x268x) & (!n_n5313) & (n_n5335) & (!n_n5334) & (x267x)) + ((!x268x) & (!n_n5313) & (n_n5335) & (n_n5334) & (!x267x)) + ((!x268x) & (!n_n5313) & (n_n5335) & (n_n5334) & (x267x)) + ((!x268x) & (n_n5313) & (!n_n5335) & (!n_n5334) & (!x267x)) + ((!x268x) & (n_n5313) & (!n_n5335) & (!n_n5334) & (x267x)) + ((!x268x) & (n_n5313) & (!n_n5335) & (n_n5334) & (!x267x)) + ((!x268x) & (n_n5313) & (!n_n5335) & (n_n5334) & (x267x)) + ((!x268x) & (n_n5313) & (n_n5335) & (!n_n5334) & (!x267x)) + ((!x268x) & (n_n5313) & (n_n5335) & (!n_n5334) & (x267x)) + ((!x268x) & (n_n5313) & (n_n5335) & (n_n5334) & (!x267x)) + ((!x268x) & (n_n5313) & (n_n5335) & (n_n5334) & (x267x)) + ((x268x) & (!n_n5313) & (!n_n5335) & (!n_n5334) & (!x267x)) + ((x268x) & (!n_n5313) & (!n_n5335) & (!n_n5334) & (x267x)) + ((x268x) & (!n_n5313) & (!n_n5335) & (n_n5334) & (!x267x)) + ((x268x) & (!n_n5313) & (!n_n5335) & (n_n5334) & (x267x)) + ((x268x) & (!n_n5313) & (n_n5335) & (!n_n5334) & (!x267x)) + ((x268x) & (!n_n5313) & (n_n5335) & (!n_n5334) & (x267x)) + ((x268x) & (!n_n5313) & (n_n5335) & (n_n5334) & (!x267x)) + ((x268x) & (!n_n5313) & (n_n5335) & (n_n5334) & (x267x)) + ((x268x) & (n_n5313) & (!n_n5335) & (!n_n5334) & (!x267x)) + ((x268x) & (n_n5313) & (!n_n5335) & (!n_n5334) & (x267x)) + ((x268x) & (n_n5313) & (!n_n5335) & (n_n5334) & (!x267x)) + ((x268x) & (n_n5313) & (!n_n5335) & (n_n5334) & (x267x)) + ((x268x) & (n_n5313) & (n_n5335) & (!n_n5334) & (!x267x)) + ((x268x) & (n_n5313) & (n_n5335) & (!n_n5334) & (x267x)) + ((x268x) & (n_n5313) & (n_n5335) & (n_n5334) & (!x267x)) + ((x268x) & (n_n5313) & (n_n5335) & (n_n5334) & (x267x)));
	assign x13565x = (((!n_n5322) & (!n_n5329) & (!n_n5327) & (n_n5328)) + ((!n_n5322) & (!n_n5329) & (n_n5327) & (!n_n5328)) + ((!n_n5322) & (!n_n5329) & (n_n5327) & (n_n5328)) + ((!n_n5322) & (n_n5329) & (!n_n5327) & (!n_n5328)) + ((!n_n5322) & (n_n5329) & (!n_n5327) & (n_n5328)) + ((!n_n5322) & (n_n5329) & (n_n5327) & (!n_n5328)) + ((!n_n5322) & (n_n5329) & (n_n5327) & (n_n5328)) + ((n_n5322) & (!n_n5329) & (!n_n5327) & (!n_n5328)) + ((n_n5322) & (!n_n5329) & (!n_n5327) & (n_n5328)) + ((n_n5322) & (!n_n5329) & (n_n5327) & (!n_n5328)) + ((n_n5322) & (!n_n5329) & (n_n5327) & (n_n5328)) + ((n_n5322) & (n_n5329) & (!n_n5327) & (!n_n5328)) + ((n_n5322) & (n_n5329) & (!n_n5327) & (n_n5328)) + ((n_n5322) & (n_n5329) & (n_n5327) & (!n_n5328)) + ((n_n5322) & (n_n5329) & (n_n5327) & (n_n5328)));
	assign n_n3996 = (((!n_n5320) & (!n_n5326) & (!x175x) & (!x13568x) & (x13565x)) + ((!n_n5320) & (!n_n5326) & (!x175x) & (x13568x) & (!x13565x)) + ((!n_n5320) & (!n_n5326) & (!x175x) & (x13568x) & (x13565x)) + ((!n_n5320) & (!n_n5326) & (x175x) & (!x13568x) & (!x13565x)) + ((!n_n5320) & (!n_n5326) & (x175x) & (!x13568x) & (x13565x)) + ((!n_n5320) & (!n_n5326) & (x175x) & (x13568x) & (!x13565x)) + ((!n_n5320) & (!n_n5326) & (x175x) & (x13568x) & (x13565x)) + ((!n_n5320) & (n_n5326) & (!x175x) & (!x13568x) & (!x13565x)) + ((!n_n5320) & (n_n5326) & (!x175x) & (!x13568x) & (x13565x)) + ((!n_n5320) & (n_n5326) & (!x175x) & (x13568x) & (!x13565x)) + ((!n_n5320) & (n_n5326) & (!x175x) & (x13568x) & (x13565x)) + ((!n_n5320) & (n_n5326) & (x175x) & (!x13568x) & (!x13565x)) + ((!n_n5320) & (n_n5326) & (x175x) & (!x13568x) & (x13565x)) + ((!n_n5320) & (n_n5326) & (x175x) & (x13568x) & (!x13565x)) + ((!n_n5320) & (n_n5326) & (x175x) & (x13568x) & (x13565x)) + ((n_n5320) & (!n_n5326) & (!x175x) & (!x13568x) & (!x13565x)) + ((n_n5320) & (!n_n5326) & (!x175x) & (!x13568x) & (x13565x)) + ((n_n5320) & (!n_n5326) & (!x175x) & (x13568x) & (!x13565x)) + ((n_n5320) & (!n_n5326) & (!x175x) & (x13568x) & (x13565x)) + ((n_n5320) & (!n_n5326) & (x175x) & (!x13568x) & (!x13565x)) + ((n_n5320) & (!n_n5326) & (x175x) & (!x13568x) & (x13565x)) + ((n_n5320) & (!n_n5326) & (x175x) & (x13568x) & (!x13565x)) + ((n_n5320) & (!n_n5326) & (x175x) & (x13568x) & (x13565x)) + ((n_n5320) & (n_n5326) & (!x175x) & (!x13568x) & (!x13565x)) + ((n_n5320) & (n_n5326) & (!x175x) & (!x13568x) & (x13565x)) + ((n_n5320) & (n_n5326) & (!x175x) & (x13568x) & (!x13565x)) + ((n_n5320) & (n_n5326) & (!x175x) & (x13568x) & (x13565x)) + ((n_n5320) & (n_n5326) & (x175x) & (!x13568x) & (!x13565x)) + ((n_n5320) & (n_n5326) & (x175x) & (!x13568x) & (x13565x)) + ((n_n5320) & (n_n5326) & (x175x) & (x13568x) & (!x13565x)) + ((n_n5320) & (n_n5326) & (x175x) & (x13568x) & (x13565x)));
	assign x13091x = (((!i_9_) & (n_n524) & (n_n455) & (n_n473)) + ((i_9_) & (n_n524) & (n_n455) & (n_n473)));
	assign x13457x = (((!i_9_) & (n_n482) & (n_n390) & (!n_n532) & (n_n534)) + ((!i_9_) & (n_n482) & (n_n390) & (n_n532) & (!n_n534)) + ((!i_9_) & (n_n482) & (n_n390) & (n_n532) & (n_n534)) + ((i_9_) & (n_n482) & (n_n390) & (!n_n532) & (n_n534)) + ((i_9_) & (n_n482) & (n_n390) & (n_n532) & (!n_n534)) + ((i_9_) & (n_n482) & (n_n390) & (n_n532) & (n_n534)));
	assign n_n4079 = (((!n_n4643) & (!n_n4642) & (!n_n4652) & (!x13454x) & (x13457x)) + ((!n_n4643) & (!n_n4642) & (!n_n4652) & (x13454x) & (!x13457x)) + ((!n_n4643) & (!n_n4642) & (!n_n4652) & (x13454x) & (x13457x)) + ((!n_n4643) & (!n_n4642) & (n_n4652) & (!x13454x) & (!x13457x)) + ((!n_n4643) & (!n_n4642) & (n_n4652) & (!x13454x) & (x13457x)) + ((!n_n4643) & (!n_n4642) & (n_n4652) & (x13454x) & (!x13457x)) + ((!n_n4643) & (!n_n4642) & (n_n4652) & (x13454x) & (x13457x)) + ((!n_n4643) & (n_n4642) & (!n_n4652) & (!x13454x) & (!x13457x)) + ((!n_n4643) & (n_n4642) & (!n_n4652) & (!x13454x) & (x13457x)) + ((!n_n4643) & (n_n4642) & (!n_n4652) & (x13454x) & (!x13457x)) + ((!n_n4643) & (n_n4642) & (!n_n4652) & (x13454x) & (x13457x)) + ((!n_n4643) & (n_n4642) & (n_n4652) & (!x13454x) & (!x13457x)) + ((!n_n4643) & (n_n4642) & (n_n4652) & (!x13454x) & (x13457x)) + ((!n_n4643) & (n_n4642) & (n_n4652) & (x13454x) & (!x13457x)) + ((!n_n4643) & (n_n4642) & (n_n4652) & (x13454x) & (x13457x)) + ((n_n4643) & (!n_n4642) & (!n_n4652) & (!x13454x) & (!x13457x)) + ((n_n4643) & (!n_n4642) & (!n_n4652) & (!x13454x) & (x13457x)) + ((n_n4643) & (!n_n4642) & (!n_n4652) & (x13454x) & (!x13457x)) + ((n_n4643) & (!n_n4642) & (!n_n4652) & (x13454x) & (x13457x)) + ((n_n4643) & (!n_n4642) & (n_n4652) & (!x13454x) & (!x13457x)) + ((n_n4643) & (!n_n4642) & (n_n4652) & (!x13454x) & (x13457x)) + ((n_n4643) & (!n_n4642) & (n_n4652) & (x13454x) & (!x13457x)) + ((n_n4643) & (!n_n4642) & (n_n4652) & (x13454x) & (x13457x)) + ((n_n4643) & (n_n4642) & (!n_n4652) & (!x13454x) & (!x13457x)) + ((n_n4643) & (n_n4642) & (!n_n4652) & (!x13454x) & (x13457x)) + ((n_n4643) & (n_n4642) & (!n_n4652) & (x13454x) & (!x13457x)) + ((n_n4643) & (n_n4642) & (!n_n4652) & (x13454x) & (x13457x)) + ((n_n4643) & (n_n4642) & (n_n4652) & (!x13454x) & (!x13457x)) + ((n_n4643) & (n_n4642) & (n_n4652) & (!x13454x) & (x13457x)) + ((n_n4643) & (n_n4642) & (n_n4652) & (x13454x) & (!x13457x)) + ((n_n4643) & (n_n4642) & (n_n4652) & (x13454x) & (x13457x)));
	assign x22124x = (((!n_n5038) & (!n_n5040) & (!n_n5034) & (!n_n5041)));
	assign n_n4527 = (((!i_9_) & (n_n482) & (n_n455) & (n_n528)));
	assign n_n4713 = (((!i_9_) & (n_n518) & (n_n534) & (n_n325)));
	assign n_n4722 = (((i_9_) & (n_n524) & (n_n518) & (n_n325)));
	assign x242x = (((!i_9_) & (n_n518) & (!n_n526) & (n_n528) & (n_n325)) + ((!i_9_) & (n_n518) & (n_n526) & (n_n528) & (n_n325)) + ((i_9_) & (n_n518) & (n_n526) & (!n_n528) & (n_n325)) + ((i_9_) & (n_n518) & (n_n526) & (n_n528) & (n_n325)));
	assign x22103x = (((!n_n4718) & (!n_n4726) & (!n_n4715) & (!n_n4716)));
	assign n_n3708 = (((!n_n4724) & (!n_n4723) & (!n_n4722) & (!x242x) & (!x22103x)) + ((!n_n4724) & (!n_n4723) & (!n_n4722) & (x242x) & (!x22103x)) + ((!n_n4724) & (!n_n4723) & (!n_n4722) & (x242x) & (x22103x)) + ((!n_n4724) & (!n_n4723) & (n_n4722) & (!x242x) & (!x22103x)) + ((!n_n4724) & (!n_n4723) & (n_n4722) & (!x242x) & (x22103x)) + ((!n_n4724) & (!n_n4723) & (n_n4722) & (x242x) & (!x22103x)) + ((!n_n4724) & (!n_n4723) & (n_n4722) & (x242x) & (x22103x)) + ((!n_n4724) & (n_n4723) & (!n_n4722) & (!x242x) & (!x22103x)) + ((!n_n4724) & (n_n4723) & (!n_n4722) & (!x242x) & (x22103x)) + ((!n_n4724) & (n_n4723) & (!n_n4722) & (x242x) & (!x22103x)) + ((!n_n4724) & (n_n4723) & (!n_n4722) & (x242x) & (x22103x)) + ((!n_n4724) & (n_n4723) & (n_n4722) & (!x242x) & (!x22103x)) + ((!n_n4724) & (n_n4723) & (n_n4722) & (!x242x) & (x22103x)) + ((!n_n4724) & (n_n4723) & (n_n4722) & (x242x) & (!x22103x)) + ((!n_n4724) & (n_n4723) & (n_n4722) & (x242x) & (x22103x)) + ((n_n4724) & (!n_n4723) & (!n_n4722) & (!x242x) & (!x22103x)) + ((n_n4724) & (!n_n4723) & (!n_n4722) & (!x242x) & (x22103x)) + ((n_n4724) & (!n_n4723) & (!n_n4722) & (x242x) & (!x22103x)) + ((n_n4724) & (!n_n4723) & (!n_n4722) & (x242x) & (x22103x)) + ((n_n4724) & (!n_n4723) & (n_n4722) & (!x242x) & (!x22103x)) + ((n_n4724) & (!n_n4723) & (n_n4722) & (!x242x) & (x22103x)) + ((n_n4724) & (!n_n4723) & (n_n4722) & (x242x) & (!x22103x)) + ((n_n4724) & (!n_n4723) & (n_n4722) & (x242x) & (x22103x)) + ((n_n4724) & (n_n4723) & (!n_n4722) & (!x242x) & (!x22103x)) + ((n_n4724) & (n_n4723) & (!n_n4722) & (!x242x) & (x22103x)) + ((n_n4724) & (n_n4723) & (!n_n4722) & (x242x) & (!x22103x)) + ((n_n4724) & (n_n4723) & (!n_n4722) & (x242x) & (x22103x)) + ((n_n4724) & (n_n4723) & (n_n4722) & (!x242x) & (!x22103x)) + ((n_n4724) & (n_n4723) & (n_n4722) & (!x242x) & (x22103x)) + ((n_n4724) & (n_n4723) & (n_n4722) & (x242x) & (!x22103x)) + ((n_n4724) & (n_n4723) & (n_n4722) & (x242x) & (x22103x)));
	assign x221x = (((!i_9_) & (n_n532) & (n_n325) & (n_n535)) + ((i_9_) & (n_n532) & (n_n325) & (n_n535)));
	assign n_n3710 = (((!n_n4696) & (!n_n4702) & (!x221x) & (!x442x) & (n_n3848)) + ((!n_n4696) & (!n_n4702) & (!x221x) & (x442x) & (!n_n3848)) + ((!n_n4696) & (!n_n4702) & (!x221x) & (x442x) & (n_n3848)) + ((!n_n4696) & (!n_n4702) & (x221x) & (!x442x) & (!n_n3848)) + ((!n_n4696) & (!n_n4702) & (x221x) & (!x442x) & (n_n3848)) + ((!n_n4696) & (!n_n4702) & (x221x) & (x442x) & (!n_n3848)) + ((!n_n4696) & (!n_n4702) & (x221x) & (x442x) & (n_n3848)) + ((!n_n4696) & (n_n4702) & (!x221x) & (!x442x) & (!n_n3848)) + ((!n_n4696) & (n_n4702) & (!x221x) & (!x442x) & (n_n3848)) + ((!n_n4696) & (n_n4702) & (!x221x) & (x442x) & (!n_n3848)) + ((!n_n4696) & (n_n4702) & (!x221x) & (x442x) & (n_n3848)) + ((!n_n4696) & (n_n4702) & (x221x) & (!x442x) & (!n_n3848)) + ((!n_n4696) & (n_n4702) & (x221x) & (!x442x) & (n_n3848)) + ((!n_n4696) & (n_n4702) & (x221x) & (x442x) & (!n_n3848)) + ((!n_n4696) & (n_n4702) & (x221x) & (x442x) & (n_n3848)) + ((n_n4696) & (!n_n4702) & (!x221x) & (!x442x) & (!n_n3848)) + ((n_n4696) & (!n_n4702) & (!x221x) & (!x442x) & (n_n3848)) + ((n_n4696) & (!n_n4702) & (!x221x) & (x442x) & (!n_n3848)) + ((n_n4696) & (!n_n4702) & (!x221x) & (x442x) & (n_n3848)) + ((n_n4696) & (!n_n4702) & (x221x) & (!x442x) & (!n_n3848)) + ((n_n4696) & (!n_n4702) & (x221x) & (!x442x) & (n_n3848)) + ((n_n4696) & (!n_n4702) & (x221x) & (x442x) & (!n_n3848)) + ((n_n4696) & (!n_n4702) & (x221x) & (x442x) & (n_n3848)) + ((n_n4696) & (n_n4702) & (!x221x) & (!x442x) & (!n_n3848)) + ((n_n4696) & (n_n4702) & (!x221x) & (!x442x) & (n_n3848)) + ((n_n4696) & (n_n4702) & (!x221x) & (x442x) & (!n_n3848)) + ((n_n4696) & (n_n4702) & (!x221x) & (x442x) & (n_n3848)) + ((n_n4696) & (n_n4702) & (x221x) & (!x442x) & (!n_n3848)) + ((n_n4696) & (n_n4702) & (x221x) & (!x442x) & (n_n3848)) + ((n_n4696) & (n_n4702) & (x221x) & (x442x) & (!n_n3848)) + ((n_n4696) & (n_n4702) & (x221x) & (x442x) & (n_n3848)));
	assign x367x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n325) & (n_n535)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n325) & (n_n535)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n325) & (n_n535)) + ((i_9_) & (n_n524) & (n_n526) & (n_n325) & (n_n535)));
	assign x22102x = (((!n_n4704) & (!n_n4711) & (!n_n4710) & (!n_n4707)));
	assign x14357x = (((!n_n4712) & (!n_n4714) & (!n_n4713) & (!x367x) & (!x22102x)) + ((!n_n4712) & (!n_n4714) & (!n_n4713) & (x367x) & (!x22102x)) + ((!n_n4712) & (!n_n4714) & (!n_n4713) & (x367x) & (x22102x)) + ((!n_n4712) & (!n_n4714) & (n_n4713) & (!x367x) & (!x22102x)) + ((!n_n4712) & (!n_n4714) & (n_n4713) & (!x367x) & (x22102x)) + ((!n_n4712) & (!n_n4714) & (n_n4713) & (x367x) & (!x22102x)) + ((!n_n4712) & (!n_n4714) & (n_n4713) & (x367x) & (x22102x)) + ((!n_n4712) & (n_n4714) & (!n_n4713) & (!x367x) & (!x22102x)) + ((!n_n4712) & (n_n4714) & (!n_n4713) & (!x367x) & (x22102x)) + ((!n_n4712) & (n_n4714) & (!n_n4713) & (x367x) & (!x22102x)) + ((!n_n4712) & (n_n4714) & (!n_n4713) & (x367x) & (x22102x)) + ((!n_n4712) & (n_n4714) & (n_n4713) & (!x367x) & (!x22102x)) + ((!n_n4712) & (n_n4714) & (n_n4713) & (!x367x) & (x22102x)) + ((!n_n4712) & (n_n4714) & (n_n4713) & (x367x) & (!x22102x)) + ((!n_n4712) & (n_n4714) & (n_n4713) & (x367x) & (x22102x)) + ((n_n4712) & (!n_n4714) & (!n_n4713) & (!x367x) & (!x22102x)) + ((n_n4712) & (!n_n4714) & (!n_n4713) & (!x367x) & (x22102x)) + ((n_n4712) & (!n_n4714) & (!n_n4713) & (x367x) & (!x22102x)) + ((n_n4712) & (!n_n4714) & (!n_n4713) & (x367x) & (x22102x)) + ((n_n4712) & (!n_n4714) & (n_n4713) & (!x367x) & (!x22102x)) + ((n_n4712) & (!n_n4714) & (n_n4713) & (!x367x) & (x22102x)) + ((n_n4712) & (!n_n4714) & (n_n4713) & (x367x) & (!x22102x)) + ((n_n4712) & (!n_n4714) & (n_n4713) & (x367x) & (x22102x)) + ((n_n4712) & (n_n4714) & (!n_n4713) & (!x367x) & (!x22102x)) + ((n_n4712) & (n_n4714) & (!n_n4713) & (!x367x) & (x22102x)) + ((n_n4712) & (n_n4714) & (!n_n4713) & (x367x) & (!x22102x)) + ((n_n4712) & (n_n4714) & (!n_n4713) & (x367x) & (x22102x)) + ((n_n4712) & (n_n4714) & (n_n4713) & (!x367x) & (!x22102x)) + ((n_n4712) & (n_n4714) & (n_n4713) & (!x367x) & (x22102x)) + ((n_n4712) & (n_n4714) & (n_n4713) & (x367x) & (!x22102x)) + ((n_n4712) & (n_n4714) & (n_n4713) & (x367x) & (x22102x)));
	assign x14362x = (((!n_n4676) & (!n_n4681) & (!n_n4679) & (!n_n4672) & (n_n4680)) + ((!n_n4676) & (!n_n4681) & (!n_n4679) & (n_n4672) & (!n_n4680)) + ((!n_n4676) & (!n_n4681) & (!n_n4679) & (n_n4672) & (n_n4680)) + ((!n_n4676) & (!n_n4681) & (n_n4679) & (!n_n4672) & (!n_n4680)) + ((!n_n4676) & (!n_n4681) & (n_n4679) & (!n_n4672) & (n_n4680)) + ((!n_n4676) & (!n_n4681) & (n_n4679) & (n_n4672) & (!n_n4680)) + ((!n_n4676) & (!n_n4681) & (n_n4679) & (n_n4672) & (n_n4680)) + ((!n_n4676) & (n_n4681) & (!n_n4679) & (!n_n4672) & (!n_n4680)) + ((!n_n4676) & (n_n4681) & (!n_n4679) & (!n_n4672) & (n_n4680)) + ((!n_n4676) & (n_n4681) & (!n_n4679) & (n_n4672) & (!n_n4680)) + ((!n_n4676) & (n_n4681) & (!n_n4679) & (n_n4672) & (n_n4680)) + ((!n_n4676) & (n_n4681) & (n_n4679) & (!n_n4672) & (!n_n4680)) + ((!n_n4676) & (n_n4681) & (n_n4679) & (!n_n4672) & (n_n4680)) + ((!n_n4676) & (n_n4681) & (n_n4679) & (n_n4672) & (!n_n4680)) + ((!n_n4676) & (n_n4681) & (n_n4679) & (n_n4672) & (n_n4680)) + ((n_n4676) & (!n_n4681) & (!n_n4679) & (!n_n4672) & (!n_n4680)) + ((n_n4676) & (!n_n4681) & (!n_n4679) & (!n_n4672) & (n_n4680)) + ((n_n4676) & (!n_n4681) & (!n_n4679) & (n_n4672) & (!n_n4680)) + ((n_n4676) & (!n_n4681) & (!n_n4679) & (n_n4672) & (n_n4680)) + ((n_n4676) & (!n_n4681) & (n_n4679) & (!n_n4672) & (!n_n4680)) + ((n_n4676) & (!n_n4681) & (n_n4679) & (!n_n4672) & (n_n4680)) + ((n_n4676) & (!n_n4681) & (n_n4679) & (n_n4672) & (!n_n4680)) + ((n_n4676) & (!n_n4681) & (n_n4679) & (n_n4672) & (n_n4680)) + ((n_n4676) & (n_n4681) & (!n_n4679) & (!n_n4672) & (!n_n4680)) + ((n_n4676) & (n_n4681) & (!n_n4679) & (!n_n4672) & (n_n4680)) + ((n_n4676) & (n_n4681) & (!n_n4679) & (n_n4672) & (!n_n4680)) + ((n_n4676) & (n_n4681) & (!n_n4679) & (n_n4672) & (n_n4680)) + ((n_n4676) & (n_n4681) & (n_n4679) & (!n_n4672) & (!n_n4680)) + ((n_n4676) & (n_n4681) & (n_n4679) & (!n_n4672) & (n_n4680)) + ((n_n4676) & (n_n4681) & (n_n4679) & (n_n4672) & (!n_n4680)) + ((n_n4676) & (n_n4681) & (n_n4679) & (n_n4672) & (n_n4680)));
	assign n_n3711 = (((!x81x) & (!x426x) & (!n_n4688) & (!n_n3849) & (x219x)) + ((!x81x) & (!x426x) & (!n_n4688) & (n_n3849) & (!x219x)) + ((!x81x) & (!x426x) & (!n_n4688) & (n_n3849) & (x219x)) + ((!x81x) & (!x426x) & (n_n4688) & (!n_n3849) & (!x219x)) + ((!x81x) & (!x426x) & (n_n4688) & (!n_n3849) & (x219x)) + ((!x81x) & (!x426x) & (n_n4688) & (n_n3849) & (!x219x)) + ((!x81x) & (!x426x) & (n_n4688) & (n_n3849) & (x219x)) + ((!x81x) & (x426x) & (!n_n4688) & (!n_n3849) & (!x219x)) + ((!x81x) & (x426x) & (!n_n4688) & (!n_n3849) & (x219x)) + ((!x81x) & (x426x) & (!n_n4688) & (n_n3849) & (!x219x)) + ((!x81x) & (x426x) & (!n_n4688) & (n_n3849) & (x219x)) + ((!x81x) & (x426x) & (n_n4688) & (!n_n3849) & (!x219x)) + ((!x81x) & (x426x) & (n_n4688) & (!n_n3849) & (x219x)) + ((!x81x) & (x426x) & (n_n4688) & (n_n3849) & (!x219x)) + ((!x81x) & (x426x) & (n_n4688) & (n_n3849) & (x219x)) + ((x81x) & (!x426x) & (!n_n4688) & (!n_n3849) & (!x219x)) + ((x81x) & (!x426x) & (!n_n4688) & (!n_n3849) & (x219x)) + ((x81x) & (!x426x) & (!n_n4688) & (n_n3849) & (!x219x)) + ((x81x) & (!x426x) & (!n_n4688) & (n_n3849) & (x219x)) + ((x81x) & (!x426x) & (n_n4688) & (!n_n3849) & (!x219x)) + ((x81x) & (!x426x) & (n_n4688) & (!n_n3849) & (x219x)) + ((x81x) & (!x426x) & (n_n4688) & (n_n3849) & (!x219x)) + ((x81x) & (!x426x) & (n_n4688) & (n_n3849) & (x219x)) + ((x81x) & (x426x) & (!n_n4688) & (!n_n3849) & (!x219x)) + ((x81x) & (x426x) & (!n_n4688) & (!n_n3849) & (x219x)) + ((x81x) & (x426x) & (!n_n4688) & (n_n3849) & (!x219x)) + ((x81x) & (x426x) & (!n_n4688) & (n_n3849) & (x219x)) + ((x81x) & (x426x) & (n_n4688) & (!n_n3849) & (!x219x)) + ((x81x) & (x426x) & (n_n4688) & (!n_n3849) & (x219x)) + ((x81x) & (x426x) & (n_n4688) & (n_n3849) & (!x219x)) + ((x81x) & (x426x) & (n_n4688) & (n_n3849) & (x219x)));
	assign x22101x = (((!n_n4666) & (!n_n4667) & (!n_n4664) & (!n_n4669)));
	assign x14371x = (((!n_n4662) & (!n_n4663) & (!n_n4657) & (!x72x) & (!x22101x)) + ((!n_n4662) & (!n_n4663) & (!n_n4657) & (x72x) & (!x22101x)) + ((!n_n4662) & (!n_n4663) & (!n_n4657) & (x72x) & (x22101x)) + ((!n_n4662) & (!n_n4663) & (n_n4657) & (!x72x) & (!x22101x)) + ((!n_n4662) & (!n_n4663) & (n_n4657) & (!x72x) & (x22101x)) + ((!n_n4662) & (!n_n4663) & (n_n4657) & (x72x) & (!x22101x)) + ((!n_n4662) & (!n_n4663) & (n_n4657) & (x72x) & (x22101x)) + ((!n_n4662) & (n_n4663) & (!n_n4657) & (!x72x) & (!x22101x)) + ((!n_n4662) & (n_n4663) & (!n_n4657) & (!x72x) & (x22101x)) + ((!n_n4662) & (n_n4663) & (!n_n4657) & (x72x) & (!x22101x)) + ((!n_n4662) & (n_n4663) & (!n_n4657) & (x72x) & (x22101x)) + ((!n_n4662) & (n_n4663) & (n_n4657) & (!x72x) & (!x22101x)) + ((!n_n4662) & (n_n4663) & (n_n4657) & (!x72x) & (x22101x)) + ((!n_n4662) & (n_n4663) & (n_n4657) & (x72x) & (!x22101x)) + ((!n_n4662) & (n_n4663) & (n_n4657) & (x72x) & (x22101x)) + ((n_n4662) & (!n_n4663) & (!n_n4657) & (!x72x) & (!x22101x)) + ((n_n4662) & (!n_n4663) & (!n_n4657) & (!x72x) & (x22101x)) + ((n_n4662) & (!n_n4663) & (!n_n4657) & (x72x) & (!x22101x)) + ((n_n4662) & (!n_n4663) & (!n_n4657) & (x72x) & (x22101x)) + ((n_n4662) & (!n_n4663) & (n_n4657) & (!x72x) & (!x22101x)) + ((n_n4662) & (!n_n4663) & (n_n4657) & (!x72x) & (x22101x)) + ((n_n4662) & (!n_n4663) & (n_n4657) & (x72x) & (!x22101x)) + ((n_n4662) & (!n_n4663) & (n_n4657) & (x72x) & (x22101x)) + ((n_n4662) & (n_n4663) & (!n_n4657) & (!x72x) & (!x22101x)) + ((n_n4662) & (n_n4663) & (!n_n4657) & (!x72x) & (x22101x)) + ((n_n4662) & (n_n4663) & (!n_n4657) & (x72x) & (!x22101x)) + ((n_n4662) & (n_n4663) & (!n_n4657) & (x72x) & (x22101x)) + ((n_n4662) & (n_n4663) & (n_n4657) & (!x72x) & (!x22101x)) + ((n_n4662) & (n_n4663) & (n_n4657) & (!x72x) & (x22101x)) + ((n_n4662) & (n_n4663) & (n_n4657) & (x72x) & (!x22101x)) + ((n_n4662) & (n_n4663) & (n_n4657) & (x72x) & (x22101x)));
	assign x80x = (((!i_9_) & (!n_n524) & (n_n390) & (n_n473) & (x20x)) + ((!i_9_) & (n_n524) & (n_n390) & (n_n473) & (!x20x)) + ((!i_9_) & (n_n524) & (n_n390) & (n_n473) & (x20x)) + ((i_9_) & (!n_n524) & (n_n390) & (n_n473) & (x20x)) + ((i_9_) & (n_n524) & (n_n390) & (n_n473) & (x20x)));
	assign n_n3649 = (((!x14362x) & (!n_n3711) & (!x14371x) & (!x80x) & (x339x)) + ((!x14362x) & (!n_n3711) & (!x14371x) & (x80x) & (!x339x)) + ((!x14362x) & (!n_n3711) & (!x14371x) & (x80x) & (x339x)) + ((!x14362x) & (!n_n3711) & (x14371x) & (!x80x) & (!x339x)) + ((!x14362x) & (!n_n3711) & (x14371x) & (!x80x) & (x339x)) + ((!x14362x) & (!n_n3711) & (x14371x) & (x80x) & (!x339x)) + ((!x14362x) & (!n_n3711) & (x14371x) & (x80x) & (x339x)) + ((!x14362x) & (n_n3711) & (!x14371x) & (!x80x) & (!x339x)) + ((!x14362x) & (n_n3711) & (!x14371x) & (!x80x) & (x339x)) + ((!x14362x) & (n_n3711) & (!x14371x) & (x80x) & (!x339x)) + ((!x14362x) & (n_n3711) & (!x14371x) & (x80x) & (x339x)) + ((!x14362x) & (n_n3711) & (x14371x) & (!x80x) & (!x339x)) + ((!x14362x) & (n_n3711) & (x14371x) & (!x80x) & (x339x)) + ((!x14362x) & (n_n3711) & (x14371x) & (x80x) & (!x339x)) + ((!x14362x) & (n_n3711) & (x14371x) & (x80x) & (x339x)) + ((x14362x) & (!n_n3711) & (!x14371x) & (!x80x) & (!x339x)) + ((x14362x) & (!n_n3711) & (!x14371x) & (!x80x) & (x339x)) + ((x14362x) & (!n_n3711) & (!x14371x) & (x80x) & (!x339x)) + ((x14362x) & (!n_n3711) & (!x14371x) & (x80x) & (x339x)) + ((x14362x) & (!n_n3711) & (x14371x) & (!x80x) & (!x339x)) + ((x14362x) & (!n_n3711) & (x14371x) & (!x80x) & (x339x)) + ((x14362x) & (!n_n3711) & (x14371x) & (x80x) & (!x339x)) + ((x14362x) & (!n_n3711) & (x14371x) & (x80x) & (x339x)) + ((x14362x) & (n_n3711) & (!x14371x) & (!x80x) & (!x339x)) + ((x14362x) & (n_n3711) & (!x14371x) & (!x80x) & (x339x)) + ((x14362x) & (n_n3711) & (!x14371x) & (x80x) & (!x339x)) + ((x14362x) & (n_n3711) & (!x14371x) & (x80x) & (x339x)) + ((x14362x) & (n_n3711) & (x14371x) & (!x80x) & (!x339x)) + ((x14362x) & (n_n3711) & (x14371x) & (!x80x) & (x339x)) + ((x14362x) & (n_n3711) & (x14371x) & (x80x) & (!x339x)) + ((x14362x) & (n_n3711) & (x14371x) & (x80x) & (x339x)));
	assign x22104x = (((!x21x) & (!x483x) & (!n_n4737) & (!n_n4732) & (!n_n4740)) + ((!x21x) & (x483x) & (!n_n4737) & (!n_n4732) & (!n_n4740)) + ((x21x) & (!x483x) & (!n_n4737) & (!n_n4732) & (!n_n4740)));
	assign x376x = (((!x21x) & (!n_n455) & (!n_n509) & (!x23x) & (n_n4484)) + ((!x21x) & (!n_n455) & (!n_n509) & (x23x) & (n_n4484)) + ((!x21x) & (!n_n455) & (n_n509) & (!x23x) & (n_n4484)) + ((!x21x) & (!n_n455) & (n_n509) & (x23x) & (n_n4484)) + ((!x21x) & (n_n455) & (!n_n509) & (!x23x) & (n_n4484)) + ((!x21x) & (n_n455) & (!n_n509) & (x23x) & (n_n4484)) + ((!x21x) & (n_n455) & (n_n509) & (!x23x) & (n_n4484)) + ((!x21x) & (n_n455) & (n_n509) & (x23x) & (!n_n4484)) + ((!x21x) & (n_n455) & (n_n509) & (x23x) & (n_n4484)) + ((x21x) & (!n_n455) & (!n_n509) & (!x23x) & (n_n4484)) + ((x21x) & (!n_n455) & (!n_n509) & (x23x) & (n_n4484)) + ((x21x) & (!n_n455) & (n_n509) & (!x23x) & (n_n4484)) + ((x21x) & (!n_n455) & (n_n509) & (x23x) & (n_n4484)) + ((x21x) & (n_n455) & (!n_n509) & (!x23x) & (n_n4484)) + ((x21x) & (n_n455) & (!n_n509) & (x23x) & (n_n4484)) + ((x21x) & (n_n455) & (n_n509) & (!x23x) & (!n_n4484)) + ((x21x) & (n_n455) & (n_n509) & (!x23x) & (n_n4484)) + ((x21x) & (n_n455) & (n_n509) & (x23x) & (!n_n4484)) + ((x21x) & (n_n455) & (n_n509) & (x23x) & (n_n4484)));
	assign n_n3727 = (((!n_n4482) & (!n_n4478) & (!x78x) & (!x199x) & (x376x)) + ((!n_n4482) & (!n_n4478) & (!x78x) & (x199x) & (!x376x)) + ((!n_n4482) & (!n_n4478) & (!x78x) & (x199x) & (x376x)) + ((!n_n4482) & (!n_n4478) & (x78x) & (!x199x) & (!x376x)) + ((!n_n4482) & (!n_n4478) & (x78x) & (!x199x) & (x376x)) + ((!n_n4482) & (!n_n4478) & (x78x) & (x199x) & (!x376x)) + ((!n_n4482) & (!n_n4478) & (x78x) & (x199x) & (x376x)) + ((!n_n4482) & (n_n4478) & (!x78x) & (!x199x) & (!x376x)) + ((!n_n4482) & (n_n4478) & (!x78x) & (!x199x) & (x376x)) + ((!n_n4482) & (n_n4478) & (!x78x) & (x199x) & (!x376x)) + ((!n_n4482) & (n_n4478) & (!x78x) & (x199x) & (x376x)) + ((!n_n4482) & (n_n4478) & (x78x) & (!x199x) & (!x376x)) + ((!n_n4482) & (n_n4478) & (x78x) & (!x199x) & (x376x)) + ((!n_n4482) & (n_n4478) & (x78x) & (x199x) & (!x376x)) + ((!n_n4482) & (n_n4478) & (x78x) & (x199x) & (x376x)) + ((n_n4482) & (!n_n4478) & (!x78x) & (!x199x) & (!x376x)) + ((n_n4482) & (!n_n4478) & (!x78x) & (!x199x) & (x376x)) + ((n_n4482) & (!n_n4478) & (!x78x) & (x199x) & (!x376x)) + ((n_n4482) & (!n_n4478) & (!x78x) & (x199x) & (x376x)) + ((n_n4482) & (!n_n4478) & (x78x) & (!x199x) & (!x376x)) + ((n_n4482) & (!n_n4478) & (x78x) & (!x199x) & (x376x)) + ((n_n4482) & (!n_n4478) & (x78x) & (x199x) & (!x376x)) + ((n_n4482) & (!n_n4478) & (x78x) & (x199x) & (x376x)) + ((n_n4482) & (n_n4478) & (!x78x) & (!x199x) & (!x376x)) + ((n_n4482) & (n_n4478) & (!x78x) & (!x199x) & (x376x)) + ((n_n4482) & (n_n4478) & (!x78x) & (x199x) & (!x376x)) + ((n_n4482) & (n_n4478) & (!x78x) & (x199x) & (x376x)) + ((n_n4482) & (n_n4478) & (x78x) & (!x199x) & (!x376x)) + ((n_n4482) & (n_n4478) & (x78x) & (!x199x) & (x376x)) + ((n_n4482) & (n_n4478) & (x78x) & (x199x) & (!x376x)) + ((n_n4482) & (n_n4478) & (x78x) & (x199x) & (x376x)));
	assign x14442x = (((!i_9_) & (n_n455) & (n_n528) & (n_n500)) + ((i_9_) & (n_n455) & (n_n528) & (n_n500)));
	assign n_n3726 = (((!n_n3883) & (!n_n4500) & (!n_n4496) & (!x163x) & (x14442x)) + ((!n_n3883) & (!n_n4500) & (!n_n4496) & (x163x) & (!x14442x)) + ((!n_n3883) & (!n_n4500) & (!n_n4496) & (x163x) & (x14442x)) + ((!n_n3883) & (!n_n4500) & (n_n4496) & (!x163x) & (!x14442x)) + ((!n_n3883) & (!n_n4500) & (n_n4496) & (!x163x) & (x14442x)) + ((!n_n3883) & (!n_n4500) & (n_n4496) & (x163x) & (!x14442x)) + ((!n_n3883) & (!n_n4500) & (n_n4496) & (x163x) & (x14442x)) + ((!n_n3883) & (n_n4500) & (!n_n4496) & (!x163x) & (!x14442x)) + ((!n_n3883) & (n_n4500) & (!n_n4496) & (!x163x) & (x14442x)) + ((!n_n3883) & (n_n4500) & (!n_n4496) & (x163x) & (!x14442x)) + ((!n_n3883) & (n_n4500) & (!n_n4496) & (x163x) & (x14442x)) + ((!n_n3883) & (n_n4500) & (n_n4496) & (!x163x) & (!x14442x)) + ((!n_n3883) & (n_n4500) & (n_n4496) & (!x163x) & (x14442x)) + ((!n_n3883) & (n_n4500) & (n_n4496) & (x163x) & (!x14442x)) + ((!n_n3883) & (n_n4500) & (n_n4496) & (x163x) & (x14442x)) + ((n_n3883) & (!n_n4500) & (!n_n4496) & (!x163x) & (!x14442x)) + ((n_n3883) & (!n_n4500) & (!n_n4496) & (!x163x) & (x14442x)) + ((n_n3883) & (!n_n4500) & (!n_n4496) & (x163x) & (!x14442x)) + ((n_n3883) & (!n_n4500) & (!n_n4496) & (x163x) & (x14442x)) + ((n_n3883) & (!n_n4500) & (n_n4496) & (!x163x) & (!x14442x)) + ((n_n3883) & (!n_n4500) & (n_n4496) & (!x163x) & (x14442x)) + ((n_n3883) & (!n_n4500) & (n_n4496) & (x163x) & (!x14442x)) + ((n_n3883) & (!n_n4500) & (n_n4496) & (x163x) & (x14442x)) + ((n_n3883) & (n_n4500) & (!n_n4496) & (!x163x) & (!x14442x)) + ((n_n3883) & (n_n4500) & (!n_n4496) & (!x163x) & (x14442x)) + ((n_n3883) & (n_n4500) & (!n_n4496) & (x163x) & (!x14442x)) + ((n_n3883) & (n_n4500) & (!n_n4496) & (x163x) & (x14442x)) + ((n_n3883) & (n_n4500) & (n_n4496) & (!x163x) & (!x14442x)) + ((n_n3883) & (n_n4500) & (n_n4496) & (!x163x) & (x14442x)) + ((n_n3883) & (n_n4500) & (n_n4496) & (x163x) & (!x14442x)) + ((n_n3883) & (n_n4500) & (n_n4496) & (x163x) & (x14442x)));
	assign x14448x = (((!x25x) & (!n_n482) & (!n_n455) & (!x24x) & (x130x)) + ((!x25x) & (!n_n482) & (!n_n455) & (x24x) & (x130x)) + ((!x25x) & (!n_n482) & (n_n455) & (!x24x) & (x130x)) + ((!x25x) & (!n_n482) & (n_n455) & (x24x) & (x130x)) + ((!x25x) & (n_n482) & (!n_n455) & (!x24x) & (x130x)) + ((!x25x) & (n_n482) & (!n_n455) & (x24x) & (x130x)) + ((!x25x) & (n_n482) & (n_n455) & (!x24x) & (x130x)) + ((!x25x) & (n_n482) & (n_n455) & (x24x) & (!x130x)) + ((!x25x) & (n_n482) & (n_n455) & (x24x) & (x130x)) + ((x25x) & (!n_n482) & (!n_n455) & (!x24x) & (x130x)) + ((x25x) & (!n_n482) & (!n_n455) & (x24x) & (x130x)) + ((x25x) & (!n_n482) & (n_n455) & (!x24x) & (x130x)) + ((x25x) & (!n_n482) & (n_n455) & (x24x) & (x130x)) + ((x25x) & (n_n482) & (!n_n455) & (!x24x) & (x130x)) + ((x25x) & (n_n482) & (!n_n455) & (x24x) & (x130x)) + ((x25x) & (n_n482) & (n_n455) & (!x24x) & (!x130x)) + ((x25x) & (n_n482) & (n_n455) & (!x24x) & (x130x)) + ((x25x) & (n_n482) & (n_n455) & (x24x) & (!x130x)) + ((x25x) & (n_n482) & (n_n455) & (x24x) & (x130x)));
	assign x14449x = (((!n_n4524) & (!n_n4518) & (!n_n4517) & (x307x)) + ((!n_n4524) & (!n_n4518) & (n_n4517) & (!x307x)) + ((!n_n4524) & (!n_n4518) & (n_n4517) & (x307x)) + ((!n_n4524) & (n_n4518) & (!n_n4517) & (!x307x)) + ((!n_n4524) & (n_n4518) & (!n_n4517) & (x307x)) + ((!n_n4524) & (n_n4518) & (n_n4517) & (!x307x)) + ((!n_n4524) & (n_n4518) & (n_n4517) & (x307x)) + ((n_n4524) & (!n_n4518) & (!n_n4517) & (!x307x)) + ((n_n4524) & (!n_n4518) & (!n_n4517) & (x307x)) + ((n_n4524) & (!n_n4518) & (n_n4517) & (!x307x)) + ((n_n4524) & (!n_n4518) & (n_n4517) & (x307x)) + ((n_n4524) & (n_n4518) & (!n_n4517) & (!x307x)) + ((n_n4524) & (n_n4518) & (!n_n4517) & (x307x)) + ((n_n4524) & (n_n4518) & (n_n4517) & (!x307x)) + ((n_n4524) & (n_n4518) & (n_n4517) & (x307x)));
	assign x14455x = (((!n_n4531) & (!n_n4507) & (!n_n4510) & (n_n4501)) + ((!n_n4531) & (!n_n4507) & (n_n4510) & (!n_n4501)) + ((!n_n4531) & (!n_n4507) & (n_n4510) & (n_n4501)) + ((!n_n4531) & (n_n4507) & (!n_n4510) & (!n_n4501)) + ((!n_n4531) & (n_n4507) & (!n_n4510) & (n_n4501)) + ((!n_n4531) & (n_n4507) & (n_n4510) & (!n_n4501)) + ((!n_n4531) & (n_n4507) & (n_n4510) & (n_n4501)) + ((n_n4531) & (!n_n4507) & (!n_n4510) & (!n_n4501)) + ((n_n4531) & (!n_n4507) & (!n_n4510) & (n_n4501)) + ((n_n4531) & (!n_n4507) & (n_n4510) & (!n_n4501)) + ((n_n4531) & (!n_n4507) & (n_n4510) & (n_n4501)) + ((n_n4531) & (n_n4507) & (!n_n4510) & (!n_n4501)) + ((n_n4531) & (n_n4507) & (!n_n4510) & (n_n4501)) + ((n_n4531) & (n_n4507) & (n_n4510) & (!n_n4501)) + ((n_n4531) & (n_n4507) & (n_n4510) & (n_n4501)));
	assign x14456x = (((!n_n4506) & (!n_n4505) & (!n_n4529) & (n_n3875)) + ((!n_n4506) & (!n_n4505) & (n_n4529) & (!n_n3875)) + ((!n_n4506) & (!n_n4505) & (n_n4529) & (n_n3875)) + ((!n_n4506) & (n_n4505) & (!n_n4529) & (!n_n3875)) + ((!n_n4506) & (n_n4505) & (!n_n4529) & (n_n3875)) + ((!n_n4506) & (n_n4505) & (n_n4529) & (!n_n3875)) + ((!n_n4506) & (n_n4505) & (n_n4529) & (n_n3875)) + ((n_n4506) & (!n_n4505) & (!n_n4529) & (!n_n3875)) + ((n_n4506) & (!n_n4505) & (!n_n4529) & (n_n3875)) + ((n_n4506) & (!n_n4505) & (n_n4529) & (!n_n3875)) + ((n_n4506) & (!n_n4505) & (n_n4529) & (n_n3875)) + ((n_n4506) & (n_n4505) & (!n_n4529) & (!n_n3875)) + ((n_n4506) & (n_n4505) & (!n_n4529) & (n_n3875)) + ((n_n4506) & (n_n4505) & (n_n4529) & (!n_n3875)) + ((n_n4506) & (n_n4505) & (n_n4529) & (n_n3875)));
	assign x14457x = (((!n_n4504) & (!n_n4503) & (!x129x) & (!x378x) & (x379x)) + ((!n_n4504) & (!n_n4503) & (!x129x) & (x378x) & (!x379x)) + ((!n_n4504) & (!n_n4503) & (!x129x) & (x378x) & (x379x)) + ((!n_n4504) & (!n_n4503) & (x129x) & (!x378x) & (!x379x)) + ((!n_n4504) & (!n_n4503) & (x129x) & (!x378x) & (x379x)) + ((!n_n4504) & (!n_n4503) & (x129x) & (x378x) & (!x379x)) + ((!n_n4504) & (!n_n4503) & (x129x) & (x378x) & (x379x)) + ((!n_n4504) & (n_n4503) & (!x129x) & (!x378x) & (!x379x)) + ((!n_n4504) & (n_n4503) & (!x129x) & (!x378x) & (x379x)) + ((!n_n4504) & (n_n4503) & (!x129x) & (x378x) & (!x379x)) + ((!n_n4504) & (n_n4503) & (!x129x) & (x378x) & (x379x)) + ((!n_n4504) & (n_n4503) & (x129x) & (!x378x) & (!x379x)) + ((!n_n4504) & (n_n4503) & (x129x) & (!x378x) & (x379x)) + ((!n_n4504) & (n_n4503) & (x129x) & (x378x) & (!x379x)) + ((!n_n4504) & (n_n4503) & (x129x) & (x378x) & (x379x)) + ((n_n4504) & (!n_n4503) & (!x129x) & (!x378x) & (!x379x)) + ((n_n4504) & (!n_n4503) & (!x129x) & (!x378x) & (x379x)) + ((n_n4504) & (!n_n4503) & (!x129x) & (x378x) & (!x379x)) + ((n_n4504) & (!n_n4503) & (!x129x) & (x378x) & (x379x)) + ((n_n4504) & (!n_n4503) & (x129x) & (!x378x) & (!x379x)) + ((n_n4504) & (!n_n4503) & (x129x) & (!x378x) & (x379x)) + ((n_n4504) & (!n_n4503) & (x129x) & (x378x) & (!x379x)) + ((n_n4504) & (!n_n4503) & (x129x) & (x378x) & (x379x)) + ((n_n4504) & (n_n4503) & (!x129x) & (!x378x) & (!x379x)) + ((n_n4504) & (n_n4503) & (!x129x) & (!x378x) & (x379x)) + ((n_n4504) & (n_n4503) & (!x129x) & (x378x) & (!x379x)) + ((n_n4504) & (n_n4503) & (!x129x) & (x378x) & (x379x)) + ((n_n4504) & (n_n4503) & (x129x) & (!x378x) & (!x379x)) + ((n_n4504) & (n_n4503) & (x129x) & (!x378x) & (x379x)) + ((n_n4504) & (n_n4503) & (x129x) & (x378x) & (!x379x)) + ((n_n4504) & (n_n4503) & (x129x) & (x378x) & (x379x)));
	assign n_n3737 = (((!n_n4359) & (!n_n4365) & (!n_n4360) & (!n_n4352) & (x14467x)) + ((!n_n4359) & (!n_n4365) & (!n_n4360) & (n_n4352) & (!x14467x)) + ((!n_n4359) & (!n_n4365) & (!n_n4360) & (n_n4352) & (x14467x)) + ((!n_n4359) & (!n_n4365) & (n_n4360) & (!n_n4352) & (!x14467x)) + ((!n_n4359) & (!n_n4365) & (n_n4360) & (!n_n4352) & (x14467x)) + ((!n_n4359) & (!n_n4365) & (n_n4360) & (n_n4352) & (!x14467x)) + ((!n_n4359) & (!n_n4365) & (n_n4360) & (n_n4352) & (x14467x)) + ((!n_n4359) & (n_n4365) & (!n_n4360) & (!n_n4352) & (!x14467x)) + ((!n_n4359) & (n_n4365) & (!n_n4360) & (!n_n4352) & (x14467x)) + ((!n_n4359) & (n_n4365) & (!n_n4360) & (n_n4352) & (!x14467x)) + ((!n_n4359) & (n_n4365) & (!n_n4360) & (n_n4352) & (x14467x)) + ((!n_n4359) & (n_n4365) & (n_n4360) & (!n_n4352) & (!x14467x)) + ((!n_n4359) & (n_n4365) & (n_n4360) & (!n_n4352) & (x14467x)) + ((!n_n4359) & (n_n4365) & (n_n4360) & (n_n4352) & (!x14467x)) + ((!n_n4359) & (n_n4365) & (n_n4360) & (n_n4352) & (x14467x)) + ((n_n4359) & (!n_n4365) & (!n_n4360) & (!n_n4352) & (!x14467x)) + ((n_n4359) & (!n_n4365) & (!n_n4360) & (!n_n4352) & (x14467x)) + ((n_n4359) & (!n_n4365) & (!n_n4360) & (n_n4352) & (!x14467x)) + ((n_n4359) & (!n_n4365) & (!n_n4360) & (n_n4352) & (x14467x)) + ((n_n4359) & (!n_n4365) & (n_n4360) & (!n_n4352) & (!x14467x)) + ((n_n4359) & (!n_n4365) & (n_n4360) & (!n_n4352) & (x14467x)) + ((n_n4359) & (!n_n4365) & (n_n4360) & (n_n4352) & (!x14467x)) + ((n_n4359) & (!n_n4365) & (n_n4360) & (n_n4352) & (x14467x)) + ((n_n4359) & (n_n4365) & (!n_n4360) & (!n_n4352) & (!x14467x)) + ((n_n4359) & (n_n4365) & (!n_n4360) & (!n_n4352) & (x14467x)) + ((n_n4359) & (n_n4365) & (!n_n4360) & (n_n4352) & (!x14467x)) + ((n_n4359) & (n_n4365) & (!n_n4360) & (n_n4352) & (x14467x)) + ((n_n4359) & (n_n4365) & (n_n4360) & (!n_n4352) & (!x14467x)) + ((n_n4359) & (n_n4365) & (n_n4360) & (!n_n4352) & (x14467x)) + ((n_n4359) & (n_n4365) & (n_n4360) & (n_n4352) & (!x14467x)) + ((n_n4359) & (n_n4365) & (n_n4360) & (n_n4352) & (x14467x)));
	assign n_n3736 = (((!n_n4369) & (!n_n4373) & (!x64x) & (x14472x)) + ((!n_n4369) & (!n_n4373) & (x64x) & (!x14472x)) + ((!n_n4369) & (!n_n4373) & (x64x) & (x14472x)) + ((!n_n4369) & (n_n4373) & (!x64x) & (!x14472x)) + ((!n_n4369) & (n_n4373) & (!x64x) & (x14472x)) + ((!n_n4369) & (n_n4373) & (x64x) & (!x14472x)) + ((!n_n4369) & (n_n4373) & (x64x) & (x14472x)) + ((n_n4369) & (!n_n4373) & (!x64x) & (!x14472x)) + ((n_n4369) & (!n_n4373) & (!x64x) & (x14472x)) + ((n_n4369) & (!n_n4373) & (x64x) & (!x14472x)) + ((n_n4369) & (!n_n4373) & (x64x) & (x14472x)) + ((n_n4369) & (n_n4373) & (!x64x) & (!x14472x)) + ((n_n4369) & (n_n4373) & (!x64x) & (x14472x)) + ((n_n4369) & (n_n4373) & (x64x) & (!x14472x)) + ((n_n4369) & (n_n4373) & (x64x) & (x14472x)));
	assign x14511x = (((!n_n4382) & (!n_n3903) & (!x14460x) & (!n_n4377) & (x281x)) + ((!n_n4382) & (!n_n3903) & (!x14460x) & (n_n4377) & (!x281x)) + ((!n_n4382) & (!n_n3903) & (!x14460x) & (n_n4377) & (x281x)) + ((!n_n4382) & (!n_n3903) & (x14460x) & (!n_n4377) & (!x281x)) + ((!n_n4382) & (!n_n3903) & (x14460x) & (!n_n4377) & (x281x)) + ((!n_n4382) & (!n_n3903) & (x14460x) & (n_n4377) & (!x281x)) + ((!n_n4382) & (!n_n3903) & (x14460x) & (n_n4377) & (x281x)) + ((!n_n4382) & (n_n3903) & (!x14460x) & (!n_n4377) & (!x281x)) + ((!n_n4382) & (n_n3903) & (!x14460x) & (!n_n4377) & (x281x)) + ((!n_n4382) & (n_n3903) & (!x14460x) & (n_n4377) & (!x281x)) + ((!n_n4382) & (n_n3903) & (!x14460x) & (n_n4377) & (x281x)) + ((!n_n4382) & (n_n3903) & (x14460x) & (!n_n4377) & (!x281x)) + ((!n_n4382) & (n_n3903) & (x14460x) & (!n_n4377) & (x281x)) + ((!n_n4382) & (n_n3903) & (x14460x) & (n_n4377) & (!x281x)) + ((!n_n4382) & (n_n3903) & (x14460x) & (n_n4377) & (x281x)) + ((n_n4382) & (!n_n3903) & (!x14460x) & (!n_n4377) & (!x281x)) + ((n_n4382) & (!n_n3903) & (!x14460x) & (!n_n4377) & (x281x)) + ((n_n4382) & (!n_n3903) & (!x14460x) & (n_n4377) & (!x281x)) + ((n_n4382) & (!n_n3903) & (!x14460x) & (n_n4377) & (x281x)) + ((n_n4382) & (!n_n3903) & (x14460x) & (!n_n4377) & (!x281x)) + ((n_n4382) & (!n_n3903) & (x14460x) & (!n_n4377) & (x281x)) + ((n_n4382) & (!n_n3903) & (x14460x) & (n_n4377) & (!x281x)) + ((n_n4382) & (!n_n3903) & (x14460x) & (n_n4377) & (x281x)) + ((n_n4382) & (n_n3903) & (!x14460x) & (!n_n4377) & (!x281x)) + ((n_n4382) & (n_n3903) & (!x14460x) & (!n_n4377) & (x281x)) + ((n_n4382) & (n_n3903) & (!x14460x) & (n_n4377) & (!x281x)) + ((n_n4382) & (n_n3903) & (!x14460x) & (n_n4377) & (x281x)) + ((n_n4382) & (n_n3903) & (x14460x) & (!n_n4377) & (!x281x)) + ((n_n4382) & (n_n3903) & (x14460x) & (!n_n4377) & (x281x)) + ((n_n4382) & (n_n3903) & (x14460x) & (n_n4377) & (!x281x)) + ((n_n4382) & (n_n3903) & (x14460x) & (n_n4377) & (x281x)));
	assign x14513x = (((!n_n3737) & (!n_n3736) & (x14511x)) + ((!n_n3737) & (n_n3736) & (!x14511x)) + ((!n_n3737) & (n_n3736) & (x14511x)) + ((n_n3737) & (!n_n3736) & (!x14511x)) + ((n_n3737) & (!n_n3736) & (x14511x)) + ((n_n3737) & (n_n3736) & (!x14511x)) + ((n_n3737) & (n_n3736) & (x14511x)));
	assign n_n3658 = (((!n_n2443) & (!n_n2445) & (!n_n3740) & (!x14486x) & (x14488x)) + ((!n_n2443) & (!n_n2445) & (!n_n3740) & (x14486x) & (!x14488x)) + ((!n_n2443) & (!n_n2445) & (!n_n3740) & (x14486x) & (x14488x)) + ((!n_n2443) & (!n_n2445) & (n_n3740) & (!x14486x) & (!x14488x)) + ((!n_n2443) & (!n_n2445) & (n_n3740) & (!x14486x) & (x14488x)) + ((!n_n2443) & (!n_n2445) & (n_n3740) & (x14486x) & (!x14488x)) + ((!n_n2443) & (!n_n2445) & (n_n3740) & (x14486x) & (x14488x)) + ((!n_n2443) & (n_n2445) & (!n_n3740) & (!x14486x) & (!x14488x)) + ((!n_n2443) & (n_n2445) & (!n_n3740) & (!x14486x) & (x14488x)) + ((!n_n2443) & (n_n2445) & (!n_n3740) & (x14486x) & (!x14488x)) + ((!n_n2443) & (n_n2445) & (!n_n3740) & (x14486x) & (x14488x)) + ((!n_n2443) & (n_n2445) & (n_n3740) & (!x14486x) & (!x14488x)) + ((!n_n2443) & (n_n2445) & (n_n3740) & (!x14486x) & (x14488x)) + ((!n_n2443) & (n_n2445) & (n_n3740) & (x14486x) & (!x14488x)) + ((!n_n2443) & (n_n2445) & (n_n3740) & (x14486x) & (x14488x)) + ((n_n2443) & (!n_n2445) & (!n_n3740) & (!x14486x) & (!x14488x)) + ((n_n2443) & (!n_n2445) & (!n_n3740) & (!x14486x) & (x14488x)) + ((n_n2443) & (!n_n2445) & (!n_n3740) & (x14486x) & (!x14488x)) + ((n_n2443) & (!n_n2445) & (!n_n3740) & (x14486x) & (x14488x)) + ((n_n2443) & (!n_n2445) & (n_n3740) & (!x14486x) & (!x14488x)) + ((n_n2443) & (!n_n2445) & (n_n3740) & (!x14486x) & (x14488x)) + ((n_n2443) & (!n_n2445) & (n_n3740) & (x14486x) & (!x14488x)) + ((n_n2443) & (!n_n2445) & (n_n3740) & (x14486x) & (x14488x)) + ((n_n2443) & (n_n2445) & (!n_n3740) & (!x14486x) & (!x14488x)) + ((n_n2443) & (n_n2445) & (!n_n3740) & (!x14486x) & (x14488x)) + ((n_n2443) & (n_n2445) & (!n_n3740) & (x14486x) & (!x14488x)) + ((n_n2443) & (n_n2445) & (!n_n3740) & (x14486x) & (x14488x)) + ((n_n2443) & (n_n2445) & (n_n3740) & (!x14486x) & (!x14488x)) + ((n_n2443) & (n_n2445) & (n_n3740) & (!x14486x) & (x14488x)) + ((n_n2443) & (n_n2445) & (n_n3740) & (x14486x) & (!x14488x)) + ((n_n2443) & (n_n2445) & (n_n3740) & (x14486x) & (x14488x)));
	assign x14507x = (((!n_n4400) & (!n_n4407) & (!n_n4405) & (!n_n4398) & (x14506x)) + ((!n_n4400) & (!n_n4407) & (!n_n4405) & (n_n4398) & (!x14506x)) + ((!n_n4400) & (!n_n4407) & (!n_n4405) & (n_n4398) & (x14506x)) + ((!n_n4400) & (!n_n4407) & (n_n4405) & (!n_n4398) & (!x14506x)) + ((!n_n4400) & (!n_n4407) & (n_n4405) & (!n_n4398) & (x14506x)) + ((!n_n4400) & (!n_n4407) & (n_n4405) & (n_n4398) & (!x14506x)) + ((!n_n4400) & (!n_n4407) & (n_n4405) & (n_n4398) & (x14506x)) + ((!n_n4400) & (n_n4407) & (!n_n4405) & (!n_n4398) & (!x14506x)) + ((!n_n4400) & (n_n4407) & (!n_n4405) & (!n_n4398) & (x14506x)) + ((!n_n4400) & (n_n4407) & (!n_n4405) & (n_n4398) & (!x14506x)) + ((!n_n4400) & (n_n4407) & (!n_n4405) & (n_n4398) & (x14506x)) + ((!n_n4400) & (n_n4407) & (n_n4405) & (!n_n4398) & (!x14506x)) + ((!n_n4400) & (n_n4407) & (n_n4405) & (!n_n4398) & (x14506x)) + ((!n_n4400) & (n_n4407) & (n_n4405) & (n_n4398) & (!x14506x)) + ((!n_n4400) & (n_n4407) & (n_n4405) & (n_n4398) & (x14506x)) + ((n_n4400) & (!n_n4407) & (!n_n4405) & (!n_n4398) & (!x14506x)) + ((n_n4400) & (!n_n4407) & (!n_n4405) & (!n_n4398) & (x14506x)) + ((n_n4400) & (!n_n4407) & (!n_n4405) & (n_n4398) & (!x14506x)) + ((n_n4400) & (!n_n4407) & (!n_n4405) & (n_n4398) & (x14506x)) + ((n_n4400) & (!n_n4407) & (n_n4405) & (!n_n4398) & (!x14506x)) + ((n_n4400) & (!n_n4407) & (n_n4405) & (!n_n4398) & (x14506x)) + ((n_n4400) & (!n_n4407) & (n_n4405) & (n_n4398) & (!x14506x)) + ((n_n4400) & (!n_n4407) & (n_n4405) & (n_n4398) & (x14506x)) + ((n_n4400) & (n_n4407) & (!n_n4405) & (!n_n4398) & (!x14506x)) + ((n_n4400) & (n_n4407) & (!n_n4405) & (!n_n4398) & (x14506x)) + ((n_n4400) & (n_n4407) & (!n_n4405) & (n_n4398) & (!x14506x)) + ((n_n4400) & (n_n4407) & (!n_n4405) & (n_n4398) & (x14506x)) + ((n_n4400) & (n_n4407) & (n_n4405) & (!n_n4398) & (!x14506x)) + ((n_n4400) & (n_n4407) & (n_n4405) & (!n_n4398) & (x14506x)) + ((n_n4400) & (n_n4407) & (n_n4405) & (n_n4398) & (!x14506x)) + ((n_n4400) & (n_n4407) & (n_n4405) & (n_n4398) & (x14506x)));
	assign n_n3732 = (((!n_n4415) & (!n_n4414) & (!x14494x) & (!x22108x)) + ((!n_n4415) & (!n_n4414) & (x14494x) & (!x22108x)) + ((!n_n4415) & (!n_n4414) & (x14494x) & (x22108x)) + ((!n_n4415) & (n_n4414) & (!x14494x) & (!x22108x)) + ((!n_n4415) & (n_n4414) & (!x14494x) & (x22108x)) + ((!n_n4415) & (n_n4414) & (x14494x) & (!x22108x)) + ((!n_n4415) & (n_n4414) & (x14494x) & (x22108x)) + ((n_n4415) & (!n_n4414) & (!x14494x) & (!x22108x)) + ((n_n4415) & (!n_n4414) & (!x14494x) & (x22108x)) + ((n_n4415) & (!n_n4414) & (x14494x) & (!x22108x)) + ((n_n4415) & (!n_n4414) & (x14494x) & (x22108x)) + ((n_n4415) & (n_n4414) & (!x14494x) & (!x22108x)) + ((n_n4415) & (n_n4414) & (!x14494x) & (x22108x)) + ((n_n4415) & (n_n4414) & (x14494x) & (!x22108x)) + ((n_n4415) & (n_n4414) & (x14494x) & (x22108x)));
	assign n_n3734 = (((!n_n4391) & (!n_n4397) & (!x216x) & (!n_n1693) & (x360x)) + ((!n_n4391) & (!n_n4397) & (!x216x) & (n_n1693) & (!x360x)) + ((!n_n4391) & (!n_n4397) & (!x216x) & (n_n1693) & (x360x)) + ((!n_n4391) & (!n_n4397) & (x216x) & (!n_n1693) & (!x360x)) + ((!n_n4391) & (!n_n4397) & (x216x) & (!n_n1693) & (x360x)) + ((!n_n4391) & (!n_n4397) & (x216x) & (n_n1693) & (!x360x)) + ((!n_n4391) & (!n_n4397) & (x216x) & (n_n1693) & (x360x)) + ((!n_n4391) & (n_n4397) & (!x216x) & (!n_n1693) & (!x360x)) + ((!n_n4391) & (n_n4397) & (!x216x) & (!n_n1693) & (x360x)) + ((!n_n4391) & (n_n4397) & (!x216x) & (n_n1693) & (!x360x)) + ((!n_n4391) & (n_n4397) & (!x216x) & (n_n1693) & (x360x)) + ((!n_n4391) & (n_n4397) & (x216x) & (!n_n1693) & (!x360x)) + ((!n_n4391) & (n_n4397) & (x216x) & (!n_n1693) & (x360x)) + ((!n_n4391) & (n_n4397) & (x216x) & (n_n1693) & (!x360x)) + ((!n_n4391) & (n_n4397) & (x216x) & (n_n1693) & (x360x)) + ((n_n4391) & (!n_n4397) & (!x216x) & (!n_n1693) & (!x360x)) + ((n_n4391) & (!n_n4397) & (!x216x) & (!n_n1693) & (x360x)) + ((n_n4391) & (!n_n4397) & (!x216x) & (n_n1693) & (!x360x)) + ((n_n4391) & (!n_n4397) & (!x216x) & (n_n1693) & (x360x)) + ((n_n4391) & (!n_n4397) & (x216x) & (!n_n1693) & (!x360x)) + ((n_n4391) & (!n_n4397) & (x216x) & (!n_n1693) & (x360x)) + ((n_n4391) & (!n_n4397) & (x216x) & (n_n1693) & (!x360x)) + ((n_n4391) & (!n_n4397) & (x216x) & (n_n1693) & (x360x)) + ((n_n4391) & (n_n4397) & (!x216x) & (!n_n1693) & (!x360x)) + ((n_n4391) & (n_n4397) & (!x216x) & (!n_n1693) & (x360x)) + ((n_n4391) & (n_n4397) & (!x216x) & (n_n1693) & (!x360x)) + ((n_n4391) & (n_n4397) & (!x216x) & (n_n1693) & (x360x)) + ((n_n4391) & (n_n4397) & (x216x) & (!n_n1693) & (!x360x)) + ((n_n4391) & (n_n4397) & (x216x) & (!n_n1693) & (x360x)) + ((n_n4391) & (n_n4397) & (x216x) & (n_n1693) & (!x360x)) + ((n_n4391) & (n_n4397) & (x216x) & (n_n1693) & (x360x)));
	assign x22165x = (((!x20x) & (!n_n4447) & (!x496x) & (!n_n4443) & (!x14527x)) + ((!x20x) & (!n_n4447) & (x496x) & (!n_n4443) & (!x14527x)) + ((x20x) & (!n_n4447) & (!x496x) & (!n_n4443) & (!x14527x)));
	assign x322x = (((!i_9_) & (!n_n524) & (n_n518) & (n_n455) & (n_n528)) + ((!i_9_) & (n_n524) & (n_n518) & (n_n455) & (n_n528)) + ((i_9_) & (n_n524) & (n_n518) & (n_n455) & (!n_n528)) + ((i_9_) & (n_n524) & (n_n518) & (n_n455) & (n_n528)));
	assign n_n5144 = (((i_7_) & (i_8_) & (i_6_) & (n_n491) & (x12x)));
	assign x13929x = (((!n_n5111) & (!n_n5112) & (!n_n5114) & (n_n5116)) + ((!n_n5111) & (!n_n5112) & (n_n5114) & (!n_n5116)) + ((!n_n5111) & (!n_n5112) & (n_n5114) & (n_n5116)) + ((!n_n5111) & (n_n5112) & (!n_n5114) & (!n_n5116)) + ((!n_n5111) & (n_n5112) & (!n_n5114) & (n_n5116)) + ((!n_n5111) & (n_n5112) & (n_n5114) & (!n_n5116)) + ((!n_n5111) & (n_n5112) & (n_n5114) & (n_n5116)) + ((n_n5111) & (!n_n5112) & (!n_n5114) & (!n_n5116)) + ((n_n5111) & (!n_n5112) & (!n_n5114) & (n_n5116)) + ((n_n5111) & (!n_n5112) & (n_n5114) & (!n_n5116)) + ((n_n5111) & (!n_n5112) & (n_n5114) & (n_n5116)) + ((n_n5111) & (n_n5112) & (!n_n5114) & (!n_n5116)) + ((n_n5111) & (n_n5112) & (!n_n5114) & (n_n5116)) + ((n_n5111) & (n_n5112) & (n_n5114) & (!n_n5116)) + ((n_n5111) & (n_n5112) & (n_n5114) & (n_n5116)));
	assign x13930x = (((!n_n5109) & (!n_n5113) & (!n_n5120) & (!n_n5117) & (n_n5119)) + ((!n_n5109) & (!n_n5113) & (!n_n5120) & (n_n5117) & (!n_n5119)) + ((!n_n5109) & (!n_n5113) & (!n_n5120) & (n_n5117) & (n_n5119)) + ((!n_n5109) & (!n_n5113) & (n_n5120) & (!n_n5117) & (!n_n5119)) + ((!n_n5109) & (!n_n5113) & (n_n5120) & (!n_n5117) & (n_n5119)) + ((!n_n5109) & (!n_n5113) & (n_n5120) & (n_n5117) & (!n_n5119)) + ((!n_n5109) & (!n_n5113) & (n_n5120) & (n_n5117) & (n_n5119)) + ((!n_n5109) & (n_n5113) & (!n_n5120) & (!n_n5117) & (!n_n5119)) + ((!n_n5109) & (n_n5113) & (!n_n5120) & (!n_n5117) & (n_n5119)) + ((!n_n5109) & (n_n5113) & (!n_n5120) & (n_n5117) & (!n_n5119)) + ((!n_n5109) & (n_n5113) & (!n_n5120) & (n_n5117) & (n_n5119)) + ((!n_n5109) & (n_n5113) & (n_n5120) & (!n_n5117) & (!n_n5119)) + ((!n_n5109) & (n_n5113) & (n_n5120) & (!n_n5117) & (n_n5119)) + ((!n_n5109) & (n_n5113) & (n_n5120) & (n_n5117) & (!n_n5119)) + ((!n_n5109) & (n_n5113) & (n_n5120) & (n_n5117) & (n_n5119)) + ((n_n5109) & (!n_n5113) & (!n_n5120) & (!n_n5117) & (!n_n5119)) + ((n_n5109) & (!n_n5113) & (!n_n5120) & (!n_n5117) & (n_n5119)) + ((n_n5109) & (!n_n5113) & (!n_n5120) & (n_n5117) & (!n_n5119)) + ((n_n5109) & (!n_n5113) & (!n_n5120) & (n_n5117) & (n_n5119)) + ((n_n5109) & (!n_n5113) & (n_n5120) & (!n_n5117) & (!n_n5119)) + ((n_n5109) & (!n_n5113) & (n_n5120) & (!n_n5117) & (n_n5119)) + ((n_n5109) & (!n_n5113) & (n_n5120) & (n_n5117) & (!n_n5119)) + ((n_n5109) & (!n_n5113) & (n_n5120) & (n_n5117) & (n_n5119)) + ((n_n5109) & (n_n5113) & (!n_n5120) & (!n_n5117) & (!n_n5119)) + ((n_n5109) & (n_n5113) & (!n_n5120) & (!n_n5117) & (n_n5119)) + ((n_n5109) & (n_n5113) & (!n_n5120) & (n_n5117) & (!n_n5119)) + ((n_n5109) & (n_n5113) & (!n_n5120) & (n_n5117) & (n_n5119)) + ((n_n5109) & (n_n5113) & (n_n5120) & (!n_n5117) & (!n_n5119)) + ((n_n5109) & (n_n5113) & (n_n5120) & (!n_n5117) & (n_n5119)) + ((n_n5109) & (n_n5113) & (n_n5120) & (n_n5117) & (!n_n5119)) + ((n_n5109) & (n_n5113) & (n_n5120) & (n_n5117) & (n_n5119)));
	assign x13947x = (((!n_n5330) & (!n_n2274) & (!n_n5329) & (!n_n2643) & (n_n5328)) + ((!n_n5330) & (!n_n2274) & (!n_n5329) & (n_n2643) & (!n_n5328)) + ((!n_n5330) & (!n_n2274) & (!n_n5329) & (n_n2643) & (n_n5328)) + ((!n_n5330) & (!n_n2274) & (n_n5329) & (!n_n2643) & (!n_n5328)) + ((!n_n5330) & (!n_n2274) & (n_n5329) & (!n_n2643) & (n_n5328)) + ((!n_n5330) & (!n_n2274) & (n_n5329) & (n_n2643) & (!n_n5328)) + ((!n_n5330) & (!n_n2274) & (n_n5329) & (n_n2643) & (n_n5328)) + ((!n_n5330) & (n_n2274) & (!n_n5329) & (!n_n2643) & (!n_n5328)) + ((!n_n5330) & (n_n2274) & (!n_n5329) & (!n_n2643) & (n_n5328)) + ((!n_n5330) & (n_n2274) & (!n_n5329) & (n_n2643) & (!n_n5328)) + ((!n_n5330) & (n_n2274) & (!n_n5329) & (n_n2643) & (n_n5328)) + ((!n_n5330) & (n_n2274) & (n_n5329) & (!n_n2643) & (!n_n5328)) + ((!n_n5330) & (n_n2274) & (n_n5329) & (!n_n2643) & (n_n5328)) + ((!n_n5330) & (n_n2274) & (n_n5329) & (n_n2643) & (!n_n5328)) + ((!n_n5330) & (n_n2274) & (n_n5329) & (n_n2643) & (n_n5328)) + ((n_n5330) & (!n_n2274) & (!n_n5329) & (!n_n2643) & (!n_n5328)) + ((n_n5330) & (!n_n2274) & (!n_n5329) & (!n_n2643) & (n_n5328)) + ((n_n5330) & (!n_n2274) & (!n_n5329) & (n_n2643) & (!n_n5328)) + ((n_n5330) & (!n_n2274) & (!n_n5329) & (n_n2643) & (n_n5328)) + ((n_n5330) & (!n_n2274) & (n_n5329) & (!n_n2643) & (!n_n5328)) + ((n_n5330) & (!n_n2274) & (n_n5329) & (!n_n2643) & (n_n5328)) + ((n_n5330) & (!n_n2274) & (n_n5329) & (n_n2643) & (!n_n5328)) + ((n_n5330) & (!n_n2274) & (n_n5329) & (n_n2643) & (n_n5328)) + ((n_n5330) & (n_n2274) & (!n_n5329) & (!n_n2643) & (!n_n5328)) + ((n_n5330) & (n_n2274) & (!n_n5329) & (!n_n2643) & (n_n5328)) + ((n_n5330) & (n_n2274) & (!n_n5329) & (n_n2643) & (!n_n5328)) + ((n_n5330) & (n_n2274) & (!n_n5329) & (n_n2643) & (n_n5328)) + ((n_n5330) & (n_n2274) & (n_n5329) & (!n_n2643) & (!n_n5328)) + ((n_n5330) & (n_n2274) & (n_n5329) & (!n_n2643) & (n_n5328)) + ((n_n5330) & (n_n2274) & (n_n5329) & (n_n2643) & (!n_n5328)) + ((n_n5330) & (n_n2274) & (n_n5329) & (n_n2643) & (n_n5328)));
	assign n_n3299 = (((!n_n5222) & (!n_n5225) & (!x384x) & (!x181x) & (x13950x)) + ((!n_n5222) & (!n_n5225) & (!x384x) & (x181x) & (!x13950x)) + ((!n_n5222) & (!n_n5225) & (!x384x) & (x181x) & (x13950x)) + ((!n_n5222) & (!n_n5225) & (x384x) & (!x181x) & (!x13950x)) + ((!n_n5222) & (!n_n5225) & (x384x) & (!x181x) & (x13950x)) + ((!n_n5222) & (!n_n5225) & (x384x) & (x181x) & (!x13950x)) + ((!n_n5222) & (!n_n5225) & (x384x) & (x181x) & (x13950x)) + ((!n_n5222) & (n_n5225) & (!x384x) & (!x181x) & (!x13950x)) + ((!n_n5222) & (n_n5225) & (!x384x) & (!x181x) & (x13950x)) + ((!n_n5222) & (n_n5225) & (!x384x) & (x181x) & (!x13950x)) + ((!n_n5222) & (n_n5225) & (!x384x) & (x181x) & (x13950x)) + ((!n_n5222) & (n_n5225) & (x384x) & (!x181x) & (!x13950x)) + ((!n_n5222) & (n_n5225) & (x384x) & (!x181x) & (x13950x)) + ((!n_n5222) & (n_n5225) & (x384x) & (x181x) & (!x13950x)) + ((!n_n5222) & (n_n5225) & (x384x) & (x181x) & (x13950x)) + ((n_n5222) & (!n_n5225) & (!x384x) & (!x181x) & (!x13950x)) + ((n_n5222) & (!n_n5225) & (!x384x) & (!x181x) & (x13950x)) + ((n_n5222) & (!n_n5225) & (!x384x) & (x181x) & (!x13950x)) + ((n_n5222) & (!n_n5225) & (!x384x) & (x181x) & (x13950x)) + ((n_n5222) & (!n_n5225) & (x384x) & (!x181x) & (!x13950x)) + ((n_n5222) & (!n_n5225) & (x384x) & (!x181x) & (x13950x)) + ((n_n5222) & (!n_n5225) & (x384x) & (x181x) & (!x13950x)) + ((n_n5222) & (!n_n5225) & (x384x) & (x181x) & (x13950x)) + ((n_n5222) & (n_n5225) & (!x384x) & (!x181x) & (!x13950x)) + ((n_n5222) & (n_n5225) & (!x384x) & (!x181x) & (x13950x)) + ((n_n5222) & (n_n5225) & (!x384x) & (x181x) & (!x13950x)) + ((n_n5222) & (n_n5225) & (!x384x) & (x181x) & (x13950x)) + ((n_n5222) & (n_n5225) & (x384x) & (!x181x) & (!x13950x)) + ((n_n5222) & (n_n5225) & (x384x) & (!x181x) & (x13950x)) + ((n_n5222) & (n_n5225) & (x384x) & (x181x) & (!x13950x)) + ((n_n5222) & (n_n5225) & (x384x) & (x181x) & (x13950x)));
	assign n_n3297 = (((!n_n5247) & (!n_n5250) & (!x446x) & (!n_n3385) & (x434x)) + ((!n_n5247) & (!n_n5250) & (!x446x) & (n_n3385) & (!x434x)) + ((!n_n5247) & (!n_n5250) & (!x446x) & (n_n3385) & (x434x)) + ((!n_n5247) & (!n_n5250) & (x446x) & (!n_n3385) & (!x434x)) + ((!n_n5247) & (!n_n5250) & (x446x) & (!n_n3385) & (x434x)) + ((!n_n5247) & (!n_n5250) & (x446x) & (n_n3385) & (!x434x)) + ((!n_n5247) & (!n_n5250) & (x446x) & (n_n3385) & (x434x)) + ((!n_n5247) & (n_n5250) & (!x446x) & (!n_n3385) & (!x434x)) + ((!n_n5247) & (n_n5250) & (!x446x) & (!n_n3385) & (x434x)) + ((!n_n5247) & (n_n5250) & (!x446x) & (n_n3385) & (!x434x)) + ((!n_n5247) & (n_n5250) & (!x446x) & (n_n3385) & (x434x)) + ((!n_n5247) & (n_n5250) & (x446x) & (!n_n3385) & (!x434x)) + ((!n_n5247) & (n_n5250) & (x446x) & (!n_n3385) & (x434x)) + ((!n_n5247) & (n_n5250) & (x446x) & (n_n3385) & (!x434x)) + ((!n_n5247) & (n_n5250) & (x446x) & (n_n3385) & (x434x)) + ((n_n5247) & (!n_n5250) & (!x446x) & (!n_n3385) & (!x434x)) + ((n_n5247) & (!n_n5250) & (!x446x) & (!n_n3385) & (x434x)) + ((n_n5247) & (!n_n5250) & (!x446x) & (n_n3385) & (!x434x)) + ((n_n5247) & (!n_n5250) & (!x446x) & (n_n3385) & (x434x)) + ((n_n5247) & (!n_n5250) & (x446x) & (!n_n3385) & (!x434x)) + ((n_n5247) & (!n_n5250) & (x446x) & (!n_n3385) & (x434x)) + ((n_n5247) & (!n_n5250) & (x446x) & (n_n3385) & (!x434x)) + ((n_n5247) & (!n_n5250) & (x446x) & (n_n3385) & (x434x)) + ((n_n5247) & (n_n5250) & (!x446x) & (!n_n3385) & (!x434x)) + ((n_n5247) & (n_n5250) & (!x446x) & (!n_n3385) & (x434x)) + ((n_n5247) & (n_n5250) & (!x446x) & (n_n3385) & (!x434x)) + ((n_n5247) & (n_n5250) & (!x446x) & (n_n3385) & (x434x)) + ((n_n5247) & (n_n5250) & (x446x) & (!n_n3385) & (!x434x)) + ((n_n5247) & (n_n5250) & (x446x) & (!n_n3385) & (x434x)) + ((n_n5247) & (n_n5250) & (x446x) & (n_n3385) & (!x434x)) + ((n_n5247) & (n_n5250) & (x446x) & (n_n3385) & (x434x)));
	assign x13959x = (((!n_n5241) & (!n_n5232) & (!n_n5236) & (n_n5237)) + ((!n_n5241) & (!n_n5232) & (n_n5236) & (!n_n5237)) + ((!n_n5241) & (!n_n5232) & (n_n5236) & (n_n5237)) + ((!n_n5241) & (n_n5232) & (!n_n5236) & (!n_n5237)) + ((!n_n5241) & (n_n5232) & (!n_n5236) & (n_n5237)) + ((!n_n5241) & (n_n5232) & (n_n5236) & (!n_n5237)) + ((!n_n5241) & (n_n5232) & (n_n5236) & (n_n5237)) + ((n_n5241) & (!n_n5232) & (!n_n5236) & (!n_n5237)) + ((n_n5241) & (!n_n5232) & (!n_n5236) & (n_n5237)) + ((n_n5241) & (!n_n5232) & (n_n5236) & (!n_n5237)) + ((n_n5241) & (!n_n5232) & (n_n5236) & (n_n5237)) + ((n_n5241) & (n_n5232) & (!n_n5236) & (!n_n5237)) + ((n_n5241) & (n_n5232) & (!n_n5236) & (n_n5237)) + ((n_n5241) & (n_n5232) & (n_n5236) & (!n_n5237)) + ((n_n5241) & (n_n5232) & (n_n5236) & (n_n5237)));
	assign x13960x = (((!n_n5244) & (!n_n5246) & (!n_n5243) & (!n_n5235) & (n_n5234)) + ((!n_n5244) & (!n_n5246) & (!n_n5243) & (n_n5235) & (!n_n5234)) + ((!n_n5244) & (!n_n5246) & (!n_n5243) & (n_n5235) & (n_n5234)) + ((!n_n5244) & (!n_n5246) & (n_n5243) & (!n_n5235) & (!n_n5234)) + ((!n_n5244) & (!n_n5246) & (n_n5243) & (!n_n5235) & (n_n5234)) + ((!n_n5244) & (!n_n5246) & (n_n5243) & (n_n5235) & (!n_n5234)) + ((!n_n5244) & (!n_n5246) & (n_n5243) & (n_n5235) & (n_n5234)) + ((!n_n5244) & (n_n5246) & (!n_n5243) & (!n_n5235) & (!n_n5234)) + ((!n_n5244) & (n_n5246) & (!n_n5243) & (!n_n5235) & (n_n5234)) + ((!n_n5244) & (n_n5246) & (!n_n5243) & (n_n5235) & (!n_n5234)) + ((!n_n5244) & (n_n5246) & (!n_n5243) & (n_n5235) & (n_n5234)) + ((!n_n5244) & (n_n5246) & (n_n5243) & (!n_n5235) & (!n_n5234)) + ((!n_n5244) & (n_n5246) & (n_n5243) & (!n_n5235) & (n_n5234)) + ((!n_n5244) & (n_n5246) & (n_n5243) & (n_n5235) & (!n_n5234)) + ((!n_n5244) & (n_n5246) & (n_n5243) & (n_n5235) & (n_n5234)) + ((n_n5244) & (!n_n5246) & (!n_n5243) & (!n_n5235) & (!n_n5234)) + ((n_n5244) & (!n_n5246) & (!n_n5243) & (!n_n5235) & (n_n5234)) + ((n_n5244) & (!n_n5246) & (!n_n5243) & (n_n5235) & (!n_n5234)) + ((n_n5244) & (!n_n5246) & (!n_n5243) & (n_n5235) & (n_n5234)) + ((n_n5244) & (!n_n5246) & (n_n5243) & (!n_n5235) & (!n_n5234)) + ((n_n5244) & (!n_n5246) & (n_n5243) & (!n_n5235) & (n_n5234)) + ((n_n5244) & (!n_n5246) & (n_n5243) & (n_n5235) & (!n_n5234)) + ((n_n5244) & (!n_n5246) & (n_n5243) & (n_n5235) & (n_n5234)) + ((n_n5244) & (n_n5246) & (!n_n5243) & (!n_n5235) & (!n_n5234)) + ((n_n5244) & (n_n5246) & (!n_n5243) & (!n_n5235) & (n_n5234)) + ((n_n5244) & (n_n5246) & (!n_n5243) & (n_n5235) & (!n_n5234)) + ((n_n5244) & (n_n5246) & (!n_n5243) & (n_n5235) & (n_n5234)) + ((n_n5244) & (n_n5246) & (n_n5243) & (!n_n5235) & (!n_n5234)) + ((n_n5244) & (n_n5246) & (n_n5243) & (!n_n5235) & (n_n5234)) + ((n_n5244) & (n_n5246) & (n_n5243) & (n_n5235) & (!n_n5234)) + ((n_n5244) & (n_n5246) & (n_n5243) & (n_n5235) & (n_n5234)));
	assign n_n3265 = (((!n_n3299) & (!n_n3297) & (!x13959x) & (x13960x)) + ((!n_n3299) & (!n_n3297) & (x13959x) & (!x13960x)) + ((!n_n3299) & (!n_n3297) & (x13959x) & (x13960x)) + ((!n_n3299) & (n_n3297) & (!x13959x) & (!x13960x)) + ((!n_n3299) & (n_n3297) & (!x13959x) & (x13960x)) + ((!n_n3299) & (n_n3297) & (x13959x) & (!x13960x)) + ((!n_n3299) & (n_n3297) & (x13959x) & (x13960x)) + ((n_n3299) & (!n_n3297) & (!x13959x) & (!x13960x)) + ((n_n3299) & (!n_n3297) & (!x13959x) & (x13960x)) + ((n_n3299) & (!n_n3297) & (x13959x) & (!x13960x)) + ((n_n3299) & (!n_n3297) & (x13959x) & (x13960x)) + ((n_n3299) & (n_n3297) & (!x13959x) & (!x13960x)) + ((n_n3299) & (n_n3297) & (!x13959x) & (x13960x)) + ((n_n3299) & (n_n3297) & (x13959x) & (!x13960x)) + ((n_n3299) & (n_n3297) & (x13959x) & (x13960x)));
	assign x419x = (((!x19x) & (!n_n520) & (x20x) & (n_n500) & (n_n65)) + ((!x19x) & (n_n520) & (x20x) & (n_n500) & (n_n65)) + ((x19x) & (!n_n520) & (x20x) & (n_n500) & (n_n65)) + ((x19x) & (n_n520) & (!x20x) & (n_n500) & (!n_n65)) + ((x19x) & (n_n520) & (!x20x) & (n_n500) & (n_n65)) + ((x19x) & (n_n520) & (x20x) & (n_n500) & (!n_n65)) + ((x19x) & (n_n520) & (x20x) & (n_n500) & (n_n65)));
	assign x13963x = (((!i_9_) & (!x19x) & (n_n524) & (n_n500) & (n_n65)) + ((!i_9_) & (x19x) & (n_n524) & (n_n500) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n524) & (n_n500) & (n_n65)) + ((i_9_) & (x19x) & (n_n524) & (n_n500) & (!n_n65)) + ((i_9_) & (x19x) & (n_n524) & (n_n500) & (n_n65)));
	assign x13965x = (((!x11x) & (!x24x) & (!n_n500) & (!n_n65) & (n_n5258)) + ((!x11x) & (!x24x) & (!n_n500) & (n_n65) & (n_n5258)) + ((!x11x) & (!x24x) & (n_n500) & (!n_n65) & (n_n5258)) + ((!x11x) & (!x24x) & (n_n500) & (n_n65) & (n_n5258)) + ((!x11x) & (x24x) & (!n_n500) & (!n_n65) & (n_n5258)) + ((!x11x) & (x24x) & (!n_n500) & (n_n65) & (n_n5258)) + ((!x11x) & (x24x) & (n_n500) & (!n_n65) & (n_n5258)) + ((!x11x) & (x24x) & (n_n500) & (n_n65) & (!n_n5258)) + ((!x11x) & (x24x) & (n_n500) & (n_n65) & (n_n5258)) + ((x11x) & (!x24x) & (!n_n500) & (!n_n65) & (n_n5258)) + ((x11x) & (!x24x) & (!n_n500) & (n_n65) & (n_n5258)) + ((x11x) & (!x24x) & (n_n500) & (!n_n65) & (n_n5258)) + ((x11x) & (!x24x) & (n_n500) & (n_n65) & (!n_n5258)) + ((x11x) & (!x24x) & (n_n500) & (n_n65) & (n_n5258)) + ((x11x) & (x24x) & (!n_n500) & (!n_n65) & (n_n5258)) + ((x11x) & (x24x) & (!n_n500) & (n_n65) & (n_n5258)) + ((x11x) & (x24x) & (n_n500) & (!n_n65) & (n_n5258)) + ((x11x) & (x24x) & (n_n500) & (n_n65) & (!n_n5258)) + ((x11x) & (x24x) & (n_n500) & (n_n65) & (n_n5258)));
	assign n_n3296 = (((!n_n5262) & (!n_n5260) & (!x419x) & (!x13963x) & (x13965x)) + ((!n_n5262) & (!n_n5260) & (!x419x) & (x13963x) & (!x13965x)) + ((!n_n5262) & (!n_n5260) & (!x419x) & (x13963x) & (x13965x)) + ((!n_n5262) & (!n_n5260) & (x419x) & (!x13963x) & (!x13965x)) + ((!n_n5262) & (!n_n5260) & (x419x) & (!x13963x) & (x13965x)) + ((!n_n5262) & (!n_n5260) & (x419x) & (x13963x) & (!x13965x)) + ((!n_n5262) & (!n_n5260) & (x419x) & (x13963x) & (x13965x)) + ((!n_n5262) & (n_n5260) & (!x419x) & (!x13963x) & (!x13965x)) + ((!n_n5262) & (n_n5260) & (!x419x) & (!x13963x) & (x13965x)) + ((!n_n5262) & (n_n5260) & (!x419x) & (x13963x) & (!x13965x)) + ((!n_n5262) & (n_n5260) & (!x419x) & (x13963x) & (x13965x)) + ((!n_n5262) & (n_n5260) & (x419x) & (!x13963x) & (!x13965x)) + ((!n_n5262) & (n_n5260) & (x419x) & (!x13963x) & (x13965x)) + ((!n_n5262) & (n_n5260) & (x419x) & (x13963x) & (!x13965x)) + ((!n_n5262) & (n_n5260) & (x419x) & (x13963x) & (x13965x)) + ((n_n5262) & (!n_n5260) & (!x419x) & (!x13963x) & (!x13965x)) + ((n_n5262) & (!n_n5260) & (!x419x) & (!x13963x) & (x13965x)) + ((n_n5262) & (!n_n5260) & (!x419x) & (x13963x) & (!x13965x)) + ((n_n5262) & (!n_n5260) & (!x419x) & (x13963x) & (x13965x)) + ((n_n5262) & (!n_n5260) & (x419x) & (!x13963x) & (!x13965x)) + ((n_n5262) & (!n_n5260) & (x419x) & (!x13963x) & (x13965x)) + ((n_n5262) & (!n_n5260) & (x419x) & (x13963x) & (!x13965x)) + ((n_n5262) & (!n_n5260) & (x419x) & (x13963x) & (x13965x)) + ((n_n5262) & (n_n5260) & (!x419x) & (!x13963x) & (!x13965x)) + ((n_n5262) & (n_n5260) & (!x419x) & (!x13963x) & (x13965x)) + ((n_n5262) & (n_n5260) & (!x419x) & (x13963x) & (!x13965x)) + ((n_n5262) & (n_n5260) & (!x419x) & (x13963x) & (x13965x)) + ((n_n5262) & (n_n5260) & (x419x) & (!x13963x) & (!x13965x)) + ((n_n5262) & (n_n5260) & (x419x) & (!x13963x) & (x13965x)) + ((n_n5262) & (n_n5260) & (x419x) & (x13963x) & (!x13965x)) + ((n_n5262) & (n_n5260) & (x419x) & (x13963x) & (x13965x)));
	assign x12372x = (((!i_9_) & (!n_n532) & (n_n534) & (n_n491) & (n_n65)) + ((!i_9_) & (n_n532) & (!n_n534) & (n_n491) & (n_n65)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n491) & (n_n65)));
	assign x204x = (((!x19x) & (!n_n491) & (!n_n530) & (!n_n3382) & (x12372x)) + ((!x19x) & (!n_n491) & (!n_n530) & (n_n3382) & (!x12372x)) + ((!x19x) & (!n_n491) & (!n_n530) & (n_n3382) & (x12372x)) + ((!x19x) & (!n_n491) & (n_n530) & (!n_n3382) & (x12372x)) + ((!x19x) & (!n_n491) & (n_n530) & (n_n3382) & (!x12372x)) + ((!x19x) & (!n_n491) & (n_n530) & (n_n3382) & (x12372x)) + ((!x19x) & (n_n491) & (!n_n530) & (!n_n3382) & (x12372x)) + ((!x19x) & (n_n491) & (!n_n530) & (n_n3382) & (!x12372x)) + ((!x19x) & (n_n491) & (!n_n530) & (n_n3382) & (x12372x)) + ((!x19x) & (n_n491) & (n_n530) & (!n_n3382) & (x12372x)) + ((!x19x) & (n_n491) & (n_n530) & (n_n3382) & (!x12372x)) + ((!x19x) & (n_n491) & (n_n530) & (n_n3382) & (x12372x)) + ((x19x) & (!n_n491) & (!n_n530) & (!n_n3382) & (x12372x)) + ((x19x) & (!n_n491) & (!n_n530) & (n_n3382) & (!x12372x)) + ((x19x) & (!n_n491) & (!n_n530) & (n_n3382) & (x12372x)) + ((x19x) & (!n_n491) & (n_n530) & (!n_n3382) & (x12372x)) + ((x19x) & (!n_n491) & (n_n530) & (n_n3382) & (!x12372x)) + ((x19x) & (!n_n491) & (n_n530) & (n_n3382) & (x12372x)) + ((x19x) & (n_n491) & (!n_n530) & (!n_n3382) & (x12372x)) + ((x19x) & (n_n491) & (!n_n530) & (n_n3382) & (!x12372x)) + ((x19x) & (n_n491) & (!n_n530) & (n_n3382) & (x12372x)) + ((x19x) & (n_n491) & (n_n530) & (!n_n3382) & (!x12372x)) + ((x19x) & (n_n491) & (n_n530) & (!n_n3382) & (x12372x)) + ((x19x) & (n_n491) & (n_n530) & (n_n3382) & (!x12372x)) + ((x19x) & (n_n491) & (n_n530) & (n_n3382) & (x12372x)));
	assign n_n5280 = (((i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n491)));
	assign x13974x = (((!x592x) & (!x11x) & (!n_n5294) & (!x441x) & (x13973x)) + ((!x592x) & (!x11x) & (!n_n5294) & (x441x) & (!x13973x)) + ((!x592x) & (!x11x) & (!n_n5294) & (x441x) & (x13973x)) + ((!x592x) & (!x11x) & (n_n5294) & (!x441x) & (!x13973x)) + ((!x592x) & (!x11x) & (n_n5294) & (!x441x) & (x13973x)) + ((!x592x) & (!x11x) & (n_n5294) & (x441x) & (!x13973x)) + ((!x592x) & (!x11x) & (n_n5294) & (x441x) & (x13973x)) + ((!x592x) & (x11x) & (!n_n5294) & (!x441x) & (x13973x)) + ((!x592x) & (x11x) & (!n_n5294) & (x441x) & (!x13973x)) + ((!x592x) & (x11x) & (!n_n5294) & (x441x) & (x13973x)) + ((!x592x) & (x11x) & (n_n5294) & (!x441x) & (!x13973x)) + ((!x592x) & (x11x) & (n_n5294) & (!x441x) & (x13973x)) + ((!x592x) & (x11x) & (n_n5294) & (x441x) & (!x13973x)) + ((!x592x) & (x11x) & (n_n5294) & (x441x) & (x13973x)) + ((x592x) & (!x11x) & (!n_n5294) & (!x441x) & (x13973x)) + ((x592x) & (!x11x) & (!n_n5294) & (x441x) & (!x13973x)) + ((x592x) & (!x11x) & (!n_n5294) & (x441x) & (x13973x)) + ((x592x) & (!x11x) & (n_n5294) & (!x441x) & (!x13973x)) + ((x592x) & (!x11x) & (n_n5294) & (!x441x) & (x13973x)) + ((x592x) & (!x11x) & (n_n5294) & (x441x) & (!x13973x)) + ((x592x) & (!x11x) & (n_n5294) & (x441x) & (x13973x)) + ((x592x) & (x11x) & (!n_n5294) & (!x441x) & (!x13973x)) + ((x592x) & (x11x) & (!n_n5294) & (!x441x) & (x13973x)) + ((x592x) & (x11x) & (!n_n5294) & (x441x) & (!x13973x)) + ((x592x) & (x11x) & (!n_n5294) & (x441x) & (x13973x)) + ((x592x) & (x11x) & (n_n5294) & (!x441x) & (!x13973x)) + ((x592x) & (x11x) & (n_n5294) & (!x441x) & (x13973x)) + ((x592x) & (x11x) & (n_n5294) & (x441x) & (!x13973x)) + ((x592x) & (x11x) & (n_n5294) & (x441x) & (x13973x)));
	assign x13976x = (((!x218x) & (!n_n3296) & (!x204x) & (!n_n5280) & (x13974x)) + ((!x218x) & (!n_n3296) & (!x204x) & (n_n5280) & (!x13974x)) + ((!x218x) & (!n_n3296) & (!x204x) & (n_n5280) & (x13974x)) + ((!x218x) & (!n_n3296) & (x204x) & (!n_n5280) & (!x13974x)) + ((!x218x) & (!n_n3296) & (x204x) & (!n_n5280) & (x13974x)) + ((!x218x) & (!n_n3296) & (x204x) & (n_n5280) & (!x13974x)) + ((!x218x) & (!n_n3296) & (x204x) & (n_n5280) & (x13974x)) + ((!x218x) & (n_n3296) & (!x204x) & (!n_n5280) & (!x13974x)) + ((!x218x) & (n_n3296) & (!x204x) & (!n_n5280) & (x13974x)) + ((!x218x) & (n_n3296) & (!x204x) & (n_n5280) & (!x13974x)) + ((!x218x) & (n_n3296) & (!x204x) & (n_n5280) & (x13974x)) + ((!x218x) & (n_n3296) & (x204x) & (!n_n5280) & (!x13974x)) + ((!x218x) & (n_n3296) & (x204x) & (!n_n5280) & (x13974x)) + ((!x218x) & (n_n3296) & (x204x) & (n_n5280) & (!x13974x)) + ((!x218x) & (n_n3296) & (x204x) & (n_n5280) & (x13974x)) + ((x218x) & (!n_n3296) & (!x204x) & (!n_n5280) & (!x13974x)) + ((x218x) & (!n_n3296) & (!x204x) & (!n_n5280) & (x13974x)) + ((x218x) & (!n_n3296) & (!x204x) & (n_n5280) & (!x13974x)) + ((x218x) & (!n_n3296) & (!x204x) & (n_n5280) & (x13974x)) + ((x218x) & (!n_n3296) & (x204x) & (!n_n5280) & (!x13974x)) + ((x218x) & (!n_n3296) & (x204x) & (!n_n5280) & (x13974x)) + ((x218x) & (!n_n3296) & (x204x) & (n_n5280) & (!x13974x)) + ((x218x) & (!n_n3296) & (x204x) & (n_n5280) & (x13974x)) + ((x218x) & (n_n3296) & (!x204x) & (!n_n5280) & (!x13974x)) + ((x218x) & (n_n3296) & (!x204x) & (!n_n5280) & (x13974x)) + ((x218x) & (n_n3296) & (!x204x) & (n_n5280) & (!x13974x)) + ((x218x) & (n_n3296) & (!x204x) & (n_n5280) & (x13974x)) + ((x218x) & (n_n3296) & (x204x) & (!n_n5280) & (!x13974x)) + ((x218x) & (n_n3296) & (x204x) & (!n_n5280) & (x13974x)) + ((x218x) & (n_n3296) & (x204x) & (n_n5280) & (!x13974x)) + ((x218x) & (n_n3296) & (x204x) & (n_n5280) & (x13974x)));
	assign n_n3293 = (((!n_n5297) & (!n_n5299) & (!n_n5306) & (!n_n5309) & (x13943x)) + ((!n_n5297) & (!n_n5299) & (!n_n5306) & (n_n5309) & (!x13943x)) + ((!n_n5297) & (!n_n5299) & (!n_n5306) & (n_n5309) & (x13943x)) + ((!n_n5297) & (!n_n5299) & (n_n5306) & (!n_n5309) & (!x13943x)) + ((!n_n5297) & (!n_n5299) & (n_n5306) & (!n_n5309) & (x13943x)) + ((!n_n5297) & (!n_n5299) & (n_n5306) & (n_n5309) & (!x13943x)) + ((!n_n5297) & (!n_n5299) & (n_n5306) & (n_n5309) & (x13943x)) + ((!n_n5297) & (n_n5299) & (!n_n5306) & (!n_n5309) & (!x13943x)) + ((!n_n5297) & (n_n5299) & (!n_n5306) & (!n_n5309) & (x13943x)) + ((!n_n5297) & (n_n5299) & (!n_n5306) & (n_n5309) & (!x13943x)) + ((!n_n5297) & (n_n5299) & (!n_n5306) & (n_n5309) & (x13943x)) + ((!n_n5297) & (n_n5299) & (n_n5306) & (!n_n5309) & (!x13943x)) + ((!n_n5297) & (n_n5299) & (n_n5306) & (!n_n5309) & (x13943x)) + ((!n_n5297) & (n_n5299) & (n_n5306) & (n_n5309) & (!x13943x)) + ((!n_n5297) & (n_n5299) & (n_n5306) & (n_n5309) & (x13943x)) + ((n_n5297) & (!n_n5299) & (!n_n5306) & (!n_n5309) & (!x13943x)) + ((n_n5297) & (!n_n5299) & (!n_n5306) & (!n_n5309) & (x13943x)) + ((n_n5297) & (!n_n5299) & (!n_n5306) & (n_n5309) & (!x13943x)) + ((n_n5297) & (!n_n5299) & (!n_n5306) & (n_n5309) & (x13943x)) + ((n_n5297) & (!n_n5299) & (n_n5306) & (!n_n5309) & (!x13943x)) + ((n_n5297) & (!n_n5299) & (n_n5306) & (!n_n5309) & (x13943x)) + ((n_n5297) & (!n_n5299) & (n_n5306) & (n_n5309) & (!x13943x)) + ((n_n5297) & (!n_n5299) & (n_n5306) & (n_n5309) & (x13943x)) + ((n_n5297) & (n_n5299) & (!n_n5306) & (!n_n5309) & (!x13943x)) + ((n_n5297) & (n_n5299) & (!n_n5306) & (!n_n5309) & (x13943x)) + ((n_n5297) & (n_n5299) & (!n_n5306) & (n_n5309) & (!x13943x)) + ((n_n5297) & (n_n5299) & (!n_n5306) & (n_n5309) & (x13943x)) + ((n_n5297) & (n_n5299) & (n_n5306) & (!n_n5309) & (!x13943x)) + ((n_n5297) & (n_n5299) & (n_n5306) & (!n_n5309) & (x13943x)) + ((n_n5297) & (n_n5299) & (n_n5306) & (n_n5309) & (!x13943x)) + ((n_n5297) & (n_n5299) & (n_n5306) & (n_n5309) & (x13943x)));
	assign n_n3254 = (((!n_n3292) & (!x13947x) & (!n_n3265) & (!x13976x) & (n_n3293)) + ((!n_n3292) & (!x13947x) & (!n_n3265) & (x13976x) & (!n_n3293)) + ((!n_n3292) & (!x13947x) & (!n_n3265) & (x13976x) & (n_n3293)) + ((!n_n3292) & (!x13947x) & (n_n3265) & (!x13976x) & (!n_n3293)) + ((!n_n3292) & (!x13947x) & (n_n3265) & (!x13976x) & (n_n3293)) + ((!n_n3292) & (!x13947x) & (n_n3265) & (x13976x) & (!n_n3293)) + ((!n_n3292) & (!x13947x) & (n_n3265) & (x13976x) & (n_n3293)) + ((!n_n3292) & (x13947x) & (!n_n3265) & (!x13976x) & (!n_n3293)) + ((!n_n3292) & (x13947x) & (!n_n3265) & (!x13976x) & (n_n3293)) + ((!n_n3292) & (x13947x) & (!n_n3265) & (x13976x) & (!n_n3293)) + ((!n_n3292) & (x13947x) & (!n_n3265) & (x13976x) & (n_n3293)) + ((!n_n3292) & (x13947x) & (n_n3265) & (!x13976x) & (!n_n3293)) + ((!n_n3292) & (x13947x) & (n_n3265) & (!x13976x) & (n_n3293)) + ((!n_n3292) & (x13947x) & (n_n3265) & (x13976x) & (!n_n3293)) + ((!n_n3292) & (x13947x) & (n_n3265) & (x13976x) & (n_n3293)) + ((n_n3292) & (!x13947x) & (!n_n3265) & (!x13976x) & (!n_n3293)) + ((n_n3292) & (!x13947x) & (!n_n3265) & (!x13976x) & (n_n3293)) + ((n_n3292) & (!x13947x) & (!n_n3265) & (x13976x) & (!n_n3293)) + ((n_n3292) & (!x13947x) & (!n_n3265) & (x13976x) & (n_n3293)) + ((n_n3292) & (!x13947x) & (n_n3265) & (!x13976x) & (!n_n3293)) + ((n_n3292) & (!x13947x) & (n_n3265) & (!x13976x) & (n_n3293)) + ((n_n3292) & (!x13947x) & (n_n3265) & (x13976x) & (!n_n3293)) + ((n_n3292) & (!x13947x) & (n_n3265) & (x13976x) & (n_n3293)) + ((n_n3292) & (x13947x) & (!n_n3265) & (!x13976x) & (!n_n3293)) + ((n_n3292) & (x13947x) & (!n_n3265) & (!x13976x) & (n_n3293)) + ((n_n3292) & (x13947x) & (!n_n3265) & (x13976x) & (!n_n3293)) + ((n_n3292) & (x13947x) & (!n_n3265) & (x13976x) & (n_n3293)) + ((n_n3292) & (x13947x) & (n_n3265) & (!x13976x) & (!n_n3293)) + ((n_n3292) & (x13947x) & (n_n3265) & (!x13976x) & (n_n3293)) + ((n_n3292) & (x13947x) & (n_n3265) & (x13976x) & (!n_n3293)) + ((n_n3292) & (x13947x) & (n_n3265) & (x13976x) & (n_n3293)));
	assign n_n1167 = (((!i_9_) & (!n_n518) & (!n_n528) & (!n_n130) & (n_n5100)) + ((!i_9_) & (!n_n518) & (!n_n528) & (n_n130) & (n_n5100)) + ((!i_9_) & (!n_n518) & (n_n528) & (!n_n130) & (n_n5100)) + ((!i_9_) & (!n_n518) & (n_n528) & (n_n130) & (n_n5100)) + ((!i_9_) & (n_n518) & (!n_n528) & (!n_n130) & (n_n5100)) + ((!i_9_) & (n_n518) & (!n_n528) & (n_n130) & (n_n5100)) + ((!i_9_) & (n_n518) & (n_n528) & (!n_n130) & (n_n5100)) + ((!i_9_) & (n_n518) & (n_n528) & (n_n130) & (!n_n5100)) + ((!i_9_) & (n_n518) & (n_n528) & (n_n130) & (n_n5100)) + ((i_9_) & (!n_n518) & (!n_n528) & (!n_n130) & (n_n5100)) + ((i_9_) & (!n_n518) & (!n_n528) & (n_n130) & (n_n5100)) + ((i_9_) & (!n_n518) & (n_n528) & (!n_n130) & (n_n5100)) + ((i_9_) & (!n_n518) & (n_n528) & (n_n130) & (n_n5100)) + ((i_9_) & (n_n518) & (!n_n528) & (!n_n130) & (n_n5100)) + ((i_9_) & (n_n518) & (!n_n528) & (n_n130) & (n_n5100)) + ((i_9_) & (n_n518) & (n_n528) & (!n_n130) & (n_n5100)) + ((i_9_) & (n_n518) & (n_n528) & (n_n130) & (!n_n5100)) + ((i_9_) & (n_n518) & (n_n528) & (n_n130) & (n_n5100)));
	assign n_n783 = (((!n_n535) & (!n_n522) & (!n_n520) & (!x12x) & (n_n5093)) + ((!n_n535) & (!n_n522) & (!n_n520) & (x12x) & (n_n5093)) + ((!n_n535) & (!n_n522) & (n_n520) & (!x12x) & (n_n5093)) + ((!n_n535) & (!n_n522) & (n_n520) & (x12x) & (n_n5093)) + ((!n_n535) & (n_n522) & (!n_n520) & (!x12x) & (n_n5093)) + ((!n_n535) & (n_n522) & (!n_n520) & (x12x) & (n_n5093)) + ((!n_n535) & (n_n522) & (n_n520) & (!x12x) & (n_n5093)) + ((!n_n535) & (n_n522) & (n_n520) & (x12x) & (n_n5093)) + ((n_n535) & (!n_n522) & (!n_n520) & (!x12x) & (n_n5093)) + ((n_n535) & (!n_n522) & (!n_n520) & (x12x) & (n_n5093)) + ((n_n535) & (!n_n522) & (n_n520) & (!x12x) & (n_n5093)) + ((n_n535) & (!n_n522) & (n_n520) & (x12x) & (!n_n5093)) + ((n_n535) & (!n_n522) & (n_n520) & (x12x) & (n_n5093)) + ((n_n535) & (n_n522) & (!n_n520) & (!x12x) & (n_n5093)) + ((n_n535) & (n_n522) & (!n_n520) & (x12x) & (!n_n5093)) + ((n_n535) & (n_n522) & (!n_n520) & (x12x) & (n_n5093)) + ((n_n535) & (n_n522) & (n_n520) & (!x12x) & (n_n5093)) + ((n_n535) & (n_n522) & (n_n520) & (x12x) & (!n_n5093)) + ((n_n535) & (n_n522) & (n_n520) & (x12x) & (n_n5093)));
	assign x14015x = (((!n_n5086) & (!n_n5087) & (!n_n3412) & (!n_n1167) & (n_n783)) + ((!n_n5086) & (!n_n5087) & (!n_n3412) & (n_n1167) & (!n_n783)) + ((!n_n5086) & (!n_n5087) & (!n_n3412) & (n_n1167) & (n_n783)) + ((!n_n5086) & (!n_n5087) & (n_n3412) & (!n_n1167) & (!n_n783)) + ((!n_n5086) & (!n_n5087) & (n_n3412) & (!n_n1167) & (n_n783)) + ((!n_n5086) & (!n_n5087) & (n_n3412) & (n_n1167) & (!n_n783)) + ((!n_n5086) & (!n_n5087) & (n_n3412) & (n_n1167) & (n_n783)) + ((!n_n5086) & (n_n5087) & (!n_n3412) & (!n_n1167) & (!n_n783)) + ((!n_n5086) & (n_n5087) & (!n_n3412) & (!n_n1167) & (n_n783)) + ((!n_n5086) & (n_n5087) & (!n_n3412) & (n_n1167) & (!n_n783)) + ((!n_n5086) & (n_n5087) & (!n_n3412) & (n_n1167) & (n_n783)) + ((!n_n5086) & (n_n5087) & (n_n3412) & (!n_n1167) & (!n_n783)) + ((!n_n5086) & (n_n5087) & (n_n3412) & (!n_n1167) & (n_n783)) + ((!n_n5086) & (n_n5087) & (n_n3412) & (n_n1167) & (!n_n783)) + ((!n_n5086) & (n_n5087) & (n_n3412) & (n_n1167) & (n_n783)) + ((n_n5086) & (!n_n5087) & (!n_n3412) & (!n_n1167) & (!n_n783)) + ((n_n5086) & (!n_n5087) & (!n_n3412) & (!n_n1167) & (n_n783)) + ((n_n5086) & (!n_n5087) & (!n_n3412) & (n_n1167) & (!n_n783)) + ((n_n5086) & (!n_n5087) & (!n_n3412) & (n_n1167) & (n_n783)) + ((n_n5086) & (!n_n5087) & (n_n3412) & (!n_n1167) & (!n_n783)) + ((n_n5086) & (!n_n5087) & (n_n3412) & (!n_n1167) & (n_n783)) + ((n_n5086) & (!n_n5087) & (n_n3412) & (n_n1167) & (!n_n783)) + ((n_n5086) & (!n_n5087) & (n_n3412) & (n_n1167) & (n_n783)) + ((n_n5086) & (n_n5087) & (!n_n3412) & (!n_n1167) & (!n_n783)) + ((n_n5086) & (n_n5087) & (!n_n3412) & (!n_n1167) & (n_n783)) + ((n_n5086) & (n_n5087) & (!n_n3412) & (n_n1167) & (!n_n783)) + ((n_n5086) & (n_n5087) & (!n_n3412) & (n_n1167) & (n_n783)) + ((n_n5086) & (n_n5087) & (n_n3412) & (!n_n1167) & (!n_n783)) + ((n_n5086) & (n_n5087) & (n_n3412) & (!n_n1167) & (n_n783)) + ((n_n5086) & (n_n5087) & (n_n3412) & (n_n1167) & (!n_n783)) + ((n_n5086) & (n_n5087) & (n_n3412) & (n_n1167) & (n_n783)));
	assign x14006x = (((!x18x) & (!x516x) & (!n_n5081) & (!n_n5069) & (n_n5076)) + ((!x18x) & (!x516x) & (!n_n5081) & (n_n5069) & (!n_n5076)) + ((!x18x) & (!x516x) & (!n_n5081) & (n_n5069) & (n_n5076)) + ((!x18x) & (!x516x) & (n_n5081) & (!n_n5069) & (!n_n5076)) + ((!x18x) & (!x516x) & (n_n5081) & (!n_n5069) & (n_n5076)) + ((!x18x) & (!x516x) & (n_n5081) & (n_n5069) & (!n_n5076)) + ((!x18x) & (!x516x) & (n_n5081) & (n_n5069) & (n_n5076)) + ((!x18x) & (x516x) & (!n_n5081) & (!n_n5069) & (n_n5076)) + ((!x18x) & (x516x) & (!n_n5081) & (n_n5069) & (!n_n5076)) + ((!x18x) & (x516x) & (!n_n5081) & (n_n5069) & (n_n5076)) + ((!x18x) & (x516x) & (n_n5081) & (!n_n5069) & (!n_n5076)) + ((!x18x) & (x516x) & (n_n5081) & (!n_n5069) & (n_n5076)) + ((!x18x) & (x516x) & (n_n5081) & (n_n5069) & (!n_n5076)) + ((!x18x) & (x516x) & (n_n5081) & (n_n5069) & (n_n5076)) + ((x18x) & (!x516x) & (!n_n5081) & (!n_n5069) & (n_n5076)) + ((x18x) & (!x516x) & (!n_n5081) & (n_n5069) & (!n_n5076)) + ((x18x) & (!x516x) & (!n_n5081) & (n_n5069) & (n_n5076)) + ((x18x) & (!x516x) & (n_n5081) & (!n_n5069) & (!n_n5076)) + ((x18x) & (!x516x) & (n_n5081) & (!n_n5069) & (n_n5076)) + ((x18x) & (!x516x) & (n_n5081) & (n_n5069) & (!n_n5076)) + ((x18x) & (!x516x) & (n_n5081) & (n_n5069) & (n_n5076)) + ((x18x) & (x516x) & (!n_n5081) & (!n_n5069) & (!n_n5076)) + ((x18x) & (x516x) & (!n_n5081) & (!n_n5069) & (n_n5076)) + ((x18x) & (x516x) & (!n_n5081) & (n_n5069) & (!n_n5076)) + ((x18x) & (x516x) & (!n_n5081) & (n_n5069) & (n_n5076)) + ((x18x) & (x516x) & (n_n5081) & (!n_n5069) & (!n_n5076)) + ((x18x) & (x516x) & (n_n5081) & (!n_n5069) & (n_n5076)) + ((x18x) & (x516x) & (n_n5081) & (n_n5069) & (!n_n5076)) + ((x18x) & (x516x) & (n_n5081) & (n_n5069) & (n_n5076)));
	assign x14007x = (((!n_n5083) & (!x160x) & (!n_n5077) & (n_n5071)) + ((!n_n5083) & (!x160x) & (n_n5077) & (!n_n5071)) + ((!n_n5083) & (!x160x) & (n_n5077) & (n_n5071)) + ((!n_n5083) & (x160x) & (!n_n5077) & (!n_n5071)) + ((!n_n5083) & (x160x) & (!n_n5077) & (n_n5071)) + ((!n_n5083) & (x160x) & (n_n5077) & (!n_n5071)) + ((!n_n5083) & (x160x) & (n_n5077) & (n_n5071)) + ((n_n5083) & (!x160x) & (!n_n5077) & (!n_n5071)) + ((n_n5083) & (!x160x) & (!n_n5077) & (n_n5071)) + ((n_n5083) & (!x160x) & (n_n5077) & (!n_n5071)) + ((n_n5083) & (!x160x) & (n_n5077) & (n_n5071)) + ((n_n5083) & (x160x) & (!n_n5077) & (!n_n5071)) + ((n_n5083) & (x160x) & (!n_n5077) & (n_n5071)) + ((n_n5083) & (x160x) & (n_n5077) & (!n_n5071)) + ((n_n5083) & (x160x) & (n_n5077) & (n_n5071)));
	assign x14014x = (((!n_n5097) & (!n_n5089) & (!x34x) & (!n_n5084) & (x232x)) + ((!n_n5097) & (!n_n5089) & (!x34x) & (n_n5084) & (!x232x)) + ((!n_n5097) & (!n_n5089) & (!x34x) & (n_n5084) & (x232x)) + ((!n_n5097) & (!n_n5089) & (x34x) & (!n_n5084) & (!x232x)) + ((!n_n5097) & (!n_n5089) & (x34x) & (!n_n5084) & (x232x)) + ((!n_n5097) & (!n_n5089) & (x34x) & (n_n5084) & (!x232x)) + ((!n_n5097) & (!n_n5089) & (x34x) & (n_n5084) & (x232x)) + ((!n_n5097) & (n_n5089) & (!x34x) & (!n_n5084) & (!x232x)) + ((!n_n5097) & (n_n5089) & (!x34x) & (!n_n5084) & (x232x)) + ((!n_n5097) & (n_n5089) & (!x34x) & (n_n5084) & (!x232x)) + ((!n_n5097) & (n_n5089) & (!x34x) & (n_n5084) & (x232x)) + ((!n_n5097) & (n_n5089) & (x34x) & (!n_n5084) & (!x232x)) + ((!n_n5097) & (n_n5089) & (x34x) & (!n_n5084) & (x232x)) + ((!n_n5097) & (n_n5089) & (x34x) & (n_n5084) & (!x232x)) + ((!n_n5097) & (n_n5089) & (x34x) & (n_n5084) & (x232x)) + ((n_n5097) & (!n_n5089) & (!x34x) & (!n_n5084) & (!x232x)) + ((n_n5097) & (!n_n5089) & (!x34x) & (!n_n5084) & (x232x)) + ((n_n5097) & (!n_n5089) & (!x34x) & (n_n5084) & (!x232x)) + ((n_n5097) & (!n_n5089) & (!x34x) & (n_n5084) & (x232x)) + ((n_n5097) & (!n_n5089) & (x34x) & (!n_n5084) & (!x232x)) + ((n_n5097) & (!n_n5089) & (x34x) & (!n_n5084) & (x232x)) + ((n_n5097) & (!n_n5089) & (x34x) & (n_n5084) & (!x232x)) + ((n_n5097) & (!n_n5089) & (x34x) & (n_n5084) & (x232x)) + ((n_n5097) & (n_n5089) & (!x34x) & (!n_n5084) & (!x232x)) + ((n_n5097) & (n_n5089) & (!x34x) & (!n_n5084) & (x232x)) + ((n_n5097) & (n_n5089) & (!x34x) & (n_n5084) & (!x232x)) + ((n_n5097) & (n_n5089) & (!x34x) & (n_n5084) & (x232x)) + ((n_n5097) & (n_n5089) & (x34x) & (!n_n5084) & (!x232x)) + ((n_n5097) & (n_n5089) & (x34x) & (!n_n5084) & (x232x)) + ((n_n5097) & (n_n5089) & (x34x) & (n_n5084) & (!x232x)) + ((n_n5097) & (n_n5089) & (x34x) & (n_n5084) & (x232x)));
	assign n_n3269 = (((!x14015x) & (!x14006x) & (!x14007x) & (x14014x)) + ((!x14015x) & (!x14006x) & (x14007x) & (!x14014x)) + ((!x14015x) & (!x14006x) & (x14007x) & (x14014x)) + ((!x14015x) & (x14006x) & (!x14007x) & (!x14014x)) + ((!x14015x) & (x14006x) & (!x14007x) & (x14014x)) + ((!x14015x) & (x14006x) & (x14007x) & (!x14014x)) + ((!x14015x) & (x14006x) & (x14007x) & (x14014x)) + ((x14015x) & (!x14006x) & (!x14007x) & (!x14014x)) + ((x14015x) & (!x14006x) & (!x14007x) & (x14014x)) + ((x14015x) & (!x14006x) & (x14007x) & (!x14014x)) + ((x14015x) & (!x14006x) & (x14007x) & (x14014x)) + ((x14015x) & (x14006x) & (!x14007x) & (!x14014x)) + ((x14015x) & (x14006x) & (!x14007x) & (x14014x)) + ((x14015x) & (x14006x) & (x14007x) & (!x14014x)) + ((x14015x) & (x14006x) & (x14007x) & (x14014x)));
	assign x14022x = (((!n_n5005) & (!n_n5003) & (!n_n5010) & (!n_n5011) & (x14021x)) + ((!n_n5005) & (!n_n5003) & (!n_n5010) & (n_n5011) & (!x14021x)) + ((!n_n5005) & (!n_n5003) & (!n_n5010) & (n_n5011) & (x14021x)) + ((!n_n5005) & (!n_n5003) & (n_n5010) & (!n_n5011) & (!x14021x)) + ((!n_n5005) & (!n_n5003) & (n_n5010) & (!n_n5011) & (x14021x)) + ((!n_n5005) & (!n_n5003) & (n_n5010) & (n_n5011) & (!x14021x)) + ((!n_n5005) & (!n_n5003) & (n_n5010) & (n_n5011) & (x14021x)) + ((!n_n5005) & (n_n5003) & (!n_n5010) & (!n_n5011) & (!x14021x)) + ((!n_n5005) & (n_n5003) & (!n_n5010) & (!n_n5011) & (x14021x)) + ((!n_n5005) & (n_n5003) & (!n_n5010) & (n_n5011) & (!x14021x)) + ((!n_n5005) & (n_n5003) & (!n_n5010) & (n_n5011) & (x14021x)) + ((!n_n5005) & (n_n5003) & (n_n5010) & (!n_n5011) & (!x14021x)) + ((!n_n5005) & (n_n5003) & (n_n5010) & (!n_n5011) & (x14021x)) + ((!n_n5005) & (n_n5003) & (n_n5010) & (n_n5011) & (!x14021x)) + ((!n_n5005) & (n_n5003) & (n_n5010) & (n_n5011) & (x14021x)) + ((n_n5005) & (!n_n5003) & (!n_n5010) & (!n_n5011) & (!x14021x)) + ((n_n5005) & (!n_n5003) & (!n_n5010) & (!n_n5011) & (x14021x)) + ((n_n5005) & (!n_n5003) & (!n_n5010) & (n_n5011) & (!x14021x)) + ((n_n5005) & (!n_n5003) & (!n_n5010) & (n_n5011) & (x14021x)) + ((n_n5005) & (!n_n5003) & (n_n5010) & (!n_n5011) & (!x14021x)) + ((n_n5005) & (!n_n5003) & (n_n5010) & (!n_n5011) & (x14021x)) + ((n_n5005) & (!n_n5003) & (n_n5010) & (n_n5011) & (!x14021x)) + ((n_n5005) & (!n_n5003) & (n_n5010) & (n_n5011) & (x14021x)) + ((n_n5005) & (n_n5003) & (!n_n5010) & (!n_n5011) & (!x14021x)) + ((n_n5005) & (n_n5003) & (!n_n5010) & (!n_n5011) & (x14021x)) + ((n_n5005) & (n_n5003) & (!n_n5010) & (n_n5011) & (!x14021x)) + ((n_n5005) & (n_n5003) & (!n_n5010) & (n_n5011) & (x14021x)) + ((n_n5005) & (n_n5003) & (n_n5010) & (!n_n5011) & (!x14021x)) + ((n_n5005) & (n_n5003) & (n_n5010) & (!n_n5011) & (x14021x)) + ((n_n5005) & (n_n5003) & (n_n5010) & (n_n5011) & (!x14021x)) + ((n_n5005) & (n_n5003) & (n_n5010) & (n_n5011) & (x14021x)));
	assign n_n3256 = (((!n_n3270) & (!n_n3315) & (!n_n3317) & (!n_n3269) & (x14022x)) + ((!n_n3270) & (!n_n3315) & (!n_n3317) & (n_n3269) & (!x14022x)) + ((!n_n3270) & (!n_n3315) & (!n_n3317) & (n_n3269) & (x14022x)) + ((!n_n3270) & (!n_n3315) & (n_n3317) & (!n_n3269) & (!x14022x)) + ((!n_n3270) & (!n_n3315) & (n_n3317) & (!n_n3269) & (x14022x)) + ((!n_n3270) & (!n_n3315) & (n_n3317) & (n_n3269) & (!x14022x)) + ((!n_n3270) & (!n_n3315) & (n_n3317) & (n_n3269) & (x14022x)) + ((!n_n3270) & (n_n3315) & (!n_n3317) & (!n_n3269) & (!x14022x)) + ((!n_n3270) & (n_n3315) & (!n_n3317) & (!n_n3269) & (x14022x)) + ((!n_n3270) & (n_n3315) & (!n_n3317) & (n_n3269) & (!x14022x)) + ((!n_n3270) & (n_n3315) & (!n_n3317) & (n_n3269) & (x14022x)) + ((!n_n3270) & (n_n3315) & (n_n3317) & (!n_n3269) & (!x14022x)) + ((!n_n3270) & (n_n3315) & (n_n3317) & (!n_n3269) & (x14022x)) + ((!n_n3270) & (n_n3315) & (n_n3317) & (n_n3269) & (!x14022x)) + ((!n_n3270) & (n_n3315) & (n_n3317) & (n_n3269) & (x14022x)) + ((n_n3270) & (!n_n3315) & (!n_n3317) & (!n_n3269) & (!x14022x)) + ((n_n3270) & (!n_n3315) & (!n_n3317) & (!n_n3269) & (x14022x)) + ((n_n3270) & (!n_n3315) & (!n_n3317) & (n_n3269) & (!x14022x)) + ((n_n3270) & (!n_n3315) & (!n_n3317) & (n_n3269) & (x14022x)) + ((n_n3270) & (!n_n3315) & (n_n3317) & (!n_n3269) & (!x14022x)) + ((n_n3270) & (!n_n3315) & (n_n3317) & (!n_n3269) & (x14022x)) + ((n_n3270) & (!n_n3315) & (n_n3317) & (n_n3269) & (!x14022x)) + ((n_n3270) & (!n_n3315) & (n_n3317) & (n_n3269) & (x14022x)) + ((n_n3270) & (n_n3315) & (!n_n3317) & (!n_n3269) & (!x14022x)) + ((n_n3270) & (n_n3315) & (!n_n3317) & (!n_n3269) & (x14022x)) + ((n_n3270) & (n_n3315) & (!n_n3317) & (n_n3269) & (!x14022x)) + ((n_n3270) & (n_n3315) & (!n_n3317) & (n_n3269) & (x14022x)) + ((n_n3270) & (n_n3315) & (n_n3317) & (!n_n3269) & (!x14022x)) + ((n_n3270) & (n_n3315) & (n_n3317) & (!n_n3269) & (x14022x)) + ((n_n3270) & (n_n3315) & (n_n3317) & (n_n3269) & (!x14022x)) + ((n_n3270) & (n_n3315) & (n_n3317) & (n_n3269) & (x14022x)));
	assign x14040x = (((!n_n5164) & (!n_n5162) & (!n_n5175) & (!n_n5177) & (n_n5176)) + ((!n_n5164) & (!n_n5162) & (!n_n5175) & (n_n5177) & (!n_n5176)) + ((!n_n5164) & (!n_n5162) & (!n_n5175) & (n_n5177) & (n_n5176)) + ((!n_n5164) & (!n_n5162) & (n_n5175) & (!n_n5177) & (!n_n5176)) + ((!n_n5164) & (!n_n5162) & (n_n5175) & (!n_n5177) & (n_n5176)) + ((!n_n5164) & (!n_n5162) & (n_n5175) & (n_n5177) & (!n_n5176)) + ((!n_n5164) & (!n_n5162) & (n_n5175) & (n_n5177) & (n_n5176)) + ((!n_n5164) & (n_n5162) & (!n_n5175) & (!n_n5177) & (!n_n5176)) + ((!n_n5164) & (n_n5162) & (!n_n5175) & (!n_n5177) & (n_n5176)) + ((!n_n5164) & (n_n5162) & (!n_n5175) & (n_n5177) & (!n_n5176)) + ((!n_n5164) & (n_n5162) & (!n_n5175) & (n_n5177) & (n_n5176)) + ((!n_n5164) & (n_n5162) & (n_n5175) & (!n_n5177) & (!n_n5176)) + ((!n_n5164) & (n_n5162) & (n_n5175) & (!n_n5177) & (n_n5176)) + ((!n_n5164) & (n_n5162) & (n_n5175) & (n_n5177) & (!n_n5176)) + ((!n_n5164) & (n_n5162) & (n_n5175) & (n_n5177) & (n_n5176)) + ((n_n5164) & (!n_n5162) & (!n_n5175) & (!n_n5177) & (!n_n5176)) + ((n_n5164) & (!n_n5162) & (!n_n5175) & (!n_n5177) & (n_n5176)) + ((n_n5164) & (!n_n5162) & (!n_n5175) & (n_n5177) & (!n_n5176)) + ((n_n5164) & (!n_n5162) & (!n_n5175) & (n_n5177) & (n_n5176)) + ((n_n5164) & (!n_n5162) & (n_n5175) & (!n_n5177) & (!n_n5176)) + ((n_n5164) & (!n_n5162) & (n_n5175) & (!n_n5177) & (n_n5176)) + ((n_n5164) & (!n_n5162) & (n_n5175) & (n_n5177) & (!n_n5176)) + ((n_n5164) & (!n_n5162) & (n_n5175) & (n_n5177) & (n_n5176)) + ((n_n5164) & (n_n5162) & (!n_n5175) & (!n_n5177) & (!n_n5176)) + ((n_n5164) & (n_n5162) & (!n_n5175) & (!n_n5177) & (n_n5176)) + ((n_n5164) & (n_n5162) & (!n_n5175) & (n_n5177) & (!n_n5176)) + ((n_n5164) & (n_n5162) & (!n_n5175) & (n_n5177) & (n_n5176)) + ((n_n5164) & (n_n5162) & (n_n5175) & (!n_n5177) & (!n_n5176)) + ((n_n5164) & (n_n5162) & (n_n5175) & (!n_n5177) & (n_n5176)) + ((n_n5164) & (n_n5162) & (n_n5175) & (n_n5177) & (!n_n5176)) + ((n_n5164) & (n_n5162) & (n_n5175) & (n_n5177) & (n_n5176)));
	assign x14041x = (((!n_n5171) & (!n_n5174) & (!n_n5167) & (!n_n5161) & (x14040x)) + ((!n_n5171) & (!n_n5174) & (!n_n5167) & (n_n5161) & (!x14040x)) + ((!n_n5171) & (!n_n5174) & (!n_n5167) & (n_n5161) & (x14040x)) + ((!n_n5171) & (!n_n5174) & (n_n5167) & (!n_n5161) & (!x14040x)) + ((!n_n5171) & (!n_n5174) & (n_n5167) & (!n_n5161) & (x14040x)) + ((!n_n5171) & (!n_n5174) & (n_n5167) & (n_n5161) & (!x14040x)) + ((!n_n5171) & (!n_n5174) & (n_n5167) & (n_n5161) & (x14040x)) + ((!n_n5171) & (n_n5174) & (!n_n5167) & (!n_n5161) & (!x14040x)) + ((!n_n5171) & (n_n5174) & (!n_n5167) & (!n_n5161) & (x14040x)) + ((!n_n5171) & (n_n5174) & (!n_n5167) & (n_n5161) & (!x14040x)) + ((!n_n5171) & (n_n5174) & (!n_n5167) & (n_n5161) & (x14040x)) + ((!n_n5171) & (n_n5174) & (n_n5167) & (!n_n5161) & (!x14040x)) + ((!n_n5171) & (n_n5174) & (n_n5167) & (!n_n5161) & (x14040x)) + ((!n_n5171) & (n_n5174) & (n_n5167) & (n_n5161) & (!x14040x)) + ((!n_n5171) & (n_n5174) & (n_n5167) & (n_n5161) & (x14040x)) + ((n_n5171) & (!n_n5174) & (!n_n5167) & (!n_n5161) & (!x14040x)) + ((n_n5171) & (!n_n5174) & (!n_n5167) & (!n_n5161) & (x14040x)) + ((n_n5171) & (!n_n5174) & (!n_n5167) & (n_n5161) & (!x14040x)) + ((n_n5171) & (!n_n5174) & (!n_n5167) & (n_n5161) & (x14040x)) + ((n_n5171) & (!n_n5174) & (n_n5167) & (!n_n5161) & (!x14040x)) + ((n_n5171) & (!n_n5174) & (n_n5167) & (!n_n5161) & (x14040x)) + ((n_n5171) & (!n_n5174) & (n_n5167) & (n_n5161) & (!x14040x)) + ((n_n5171) & (!n_n5174) & (n_n5167) & (n_n5161) & (x14040x)) + ((n_n5171) & (n_n5174) & (!n_n5167) & (!n_n5161) & (!x14040x)) + ((n_n5171) & (n_n5174) & (!n_n5167) & (!n_n5161) & (x14040x)) + ((n_n5171) & (n_n5174) & (!n_n5167) & (n_n5161) & (!x14040x)) + ((n_n5171) & (n_n5174) & (!n_n5167) & (n_n5161) & (x14040x)) + ((n_n5171) & (n_n5174) & (n_n5167) & (!n_n5161) & (!x14040x)) + ((n_n5171) & (n_n5174) & (n_n5167) & (!n_n5161) & (x14040x)) + ((n_n5171) & (n_n5174) & (n_n5167) & (n_n5161) & (!x14040x)) + ((n_n5171) & (n_n5174) & (n_n5167) & (n_n5161) & (x14040x)));
	assign n_n3267 = (((!n_n3303) & (!n_n3305) & (x14041x)) + ((!n_n3303) & (n_n3305) & (!x14041x)) + ((!n_n3303) & (n_n3305) & (x14041x)) + ((n_n3303) & (!n_n3305) & (!x14041x)) + ((n_n3303) & (!n_n3305) & (x14041x)) + ((n_n3303) & (n_n3305) & (!x14041x)) + ((n_n3303) & (n_n3305) & (x14041x)));
	assign x14056x = (((!n_n528) & (!x12x) & (!n_n464) & (!n_n5197) & (x14054x)) + ((!n_n528) & (!x12x) & (!n_n464) & (n_n5197) & (!x14054x)) + ((!n_n528) & (!x12x) & (!n_n464) & (n_n5197) & (x14054x)) + ((!n_n528) & (!x12x) & (n_n464) & (!n_n5197) & (x14054x)) + ((!n_n528) & (!x12x) & (n_n464) & (n_n5197) & (!x14054x)) + ((!n_n528) & (!x12x) & (n_n464) & (n_n5197) & (x14054x)) + ((!n_n528) & (x12x) & (!n_n464) & (!n_n5197) & (x14054x)) + ((!n_n528) & (x12x) & (!n_n464) & (n_n5197) & (!x14054x)) + ((!n_n528) & (x12x) & (!n_n464) & (n_n5197) & (x14054x)) + ((!n_n528) & (x12x) & (n_n464) & (!n_n5197) & (x14054x)) + ((!n_n528) & (x12x) & (n_n464) & (n_n5197) & (!x14054x)) + ((!n_n528) & (x12x) & (n_n464) & (n_n5197) & (x14054x)) + ((n_n528) & (!x12x) & (!n_n464) & (!n_n5197) & (x14054x)) + ((n_n528) & (!x12x) & (!n_n464) & (n_n5197) & (!x14054x)) + ((n_n528) & (!x12x) & (!n_n464) & (n_n5197) & (x14054x)) + ((n_n528) & (!x12x) & (n_n464) & (!n_n5197) & (x14054x)) + ((n_n528) & (!x12x) & (n_n464) & (n_n5197) & (!x14054x)) + ((n_n528) & (!x12x) & (n_n464) & (n_n5197) & (x14054x)) + ((n_n528) & (x12x) & (!n_n464) & (!n_n5197) & (x14054x)) + ((n_n528) & (x12x) & (!n_n464) & (n_n5197) & (!x14054x)) + ((n_n528) & (x12x) & (!n_n464) & (n_n5197) & (x14054x)) + ((n_n528) & (x12x) & (n_n464) & (!n_n5197) & (!x14054x)) + ((n_n528) & (x12x) & (n_n464) & (!n_n5197) & (x14054x)) + ((n_n528) & (x12x) & (n_n464) & (n_n5197) & (!x14054x)) + ((n_n528) & (x12x) & (n_n464) & (n_n5197) & (x14054x)));
	assign x14057x = (((!n_n5193) & (!n_n5189) & (!n_n5188) & (!n_n5199) & (x14056x)) + ((!n_n5193) & (!n_n5189) & (!n_n5188) & (n_n5199) & (!x14056x)) + ((!n_n5193) & (!n_n5189) & (!n_n5188) & (n_n5199) & (x14056x)) + ((!n_n5193) & (!n_n5189) & (n_n5188) & (!n_n5199) & (!x14056x)) + ((!n_n5193) & (!n_n5189) & (n_n5188) & (!n_n5199) & (x14056x)) + ((!n_n5193) & (!n_n5189) & (n_n5188) & (n_n5199) & (!x14056x)) + ((!n_n5193) & (!n_n5189) & (n_n5188) & (n_n5199) & (x14056x)) + ((!n_n5193) & (n_n5189) & (!n_n5188) & (!n_n5199) & (!x14056x)) + ((!n_n5193) & (n_n5189) & (!n_n5188) & (!n_n5199) & (x14056x)) + ((!n_n5193) & (n_n5189) & (!n_n5188) & (n_n5199) & (!x14056x)) + ((!n_n5193) & (n_n5189) & (!n_n5188) & (n_n5199) & (x14056x)) + ((!n_n5193) & (n_n5189) & (n_n5188) & (!n_n5199) & (!x14056x)) + ((!n_n5193) & (n_n5189) & (n_n5188) & (!n_n5199) & (x14056x)) + ((!n_n5193) & (n_n5189) & (n_n5188) & (n_n5199) & (!x14056x)) + ((!n_n5193) & (n_n5189) & (n_n5188) & (n_n5199) & (x14056x)) + ((n_n5193) & (!n_n5189) & (!n_n5188) & (!n_n5199) & (!x14056x)) + ((n_n5193) & (!n_n5189) & (!n_n5188) & (!n_n5199) & (x14056x)) + ((n_n5193) & (!n_n5189) & (!n_n5188) & (n_n5199) & (!x14056x)) + ((n_n5193) & (!n_n5189) & (!n_n5188) & (n_n5199) & (x14056x)) + ((n_n5193) & (!n_n5189) & (n_n5188) & (!n_n5199) & (!x14056x)) + ((n_n5193) & (!n_n5189) & (n_n5188) & (!n_n5199) & (x14056x)) + ((n_n5193) & (!n_n5189) & (n_n5188) & (n_n5199) & (!x14056x)) + ((n_n5193) & (!n_n5189) & (n_n5188) & (n_n5199) & (x14056x)) + ((n_n5193) & (n_n5189) & (!n_n5188) & (!n_n5199) & (!x14056x)) + ((n_n5193) & (n_n5189) & (!n_n5188) & (!n_n5199) & (x14056x)) + ((n_n5193) & (n_n5189) & (!n_n5188) & (n_n5199) & (!x14056x)) + ((n_n5193) & (n_n5189) & (!n_n5188) & (n_n5199) & (x14056x)) + ((n_n5193) & (n_n5189) & (n_n5188) & (!n_n5199) & (!x14056x)) + ((n_n5193) & (n_n5189) & (n_n5188) & (!n_n5199) & (x14056x)) + ((n_n5193) & (n_n5189) & (n_n5188) & (n_n5199) & (!x14056x)) + ((n_n5193) & (n_n5189) & (n_n5188) & (n_n5199) & (x14056x)));
	assign x211x = (((!n_n522) & (n_n130) & (!x12x) & (x20x) & (n_n500)) + ((!n_n522) & (n_n130) & (x12x) & (x20x) & (n_n500)) + ((n_n522) & (!n_n130) & (x12x) & (!x20x) & (n_n500)) + ((n_n522) & (!n_n130) & (x12x) & (x20x) & (n_n500)) + ((n_n522) & (n_n130) & (!x12x) & (x20x) & (n_n500)) + ((n_n522) & (n_n130) & (x12x) & (!x20x) & (n_n500)) + ((n_n522) & (n_n130) & (x12x) & (x20x) & (n_n500)));
	assign n_n3300 = (((!n_n5212) & (!x449x) & (!n_n2665) & (!x223x) & (n_n5211)) + ((!n_n5212) & (!x449x) & (!n_n2665) & (x223x) & (!n_n5211)) + ((!n_n5212) & (!x449x) & (!n_n2665) & (x223x) & (n_n5211)) + ((!n_n5212) & (!x449x) & (n_n2665) & (!x223x) & (!n_n5211)) + ((!n_n5212) & (!x449x) & (n_n2665) & (!x223x) & (n_n5211)) + ((!n_n5212) & (!x449x) & (n_n2665) & (x223x) & (!n_n5211)) + ((!n_n5212) & (!x449x) & (n_n2665) & (x223x) & (n_n5211)) + ((!n_n5212) & (x449x) & (!n_n2665) & (!x223x) & (!n_n5211)) + ((!n_n5212) & (x449x) & (!n_n2665) & (!x223x) & (n_n5211)) + ((!n_n5212) & (x449x) & (!n_n2665) & (x223x) & (!n_n5211)) + ((!n_n5212) & (x449x) & (!n_n2665) & (x223x) & (n_n5211)) + ((!n_n5212) & (x449x) & (n_n2665) & (!x223x) & (!n_n5211)) + ((!n_n5212) & (x449x) & (n_n2665) & (!x223x) & (n_n5211)) + ((!n_n5212) & (x449x) & (n_n2665) & (x223x) & (!n_n5211)) + ((!n_n5212) & (x449x) & (n_n2665) & (x223x) & (n_n5211)) + ((n_n5212) & (!x449x) & (!n_n2665) & (!x223x) & (!n_n5211)) + ((n_n5212) & (!x449x) & (!n_n2665) & (!x223x) & (n_n5211)) + ((n_n5212) & (!x449x) & (!n_n2665) & (x223x) & (!n_n5211)) + ((n_n5212) & (!x449x) & (!n_n2665) & (x223x) & (n_n5211)) + ((n_n5212) & (!x449x) & (n_n2665) & (!x223x) & (!n_n5211)) + ((n_n5212) & (!x449x) & (n_n2665) & (!x223x) & (n_n5211)) + ((n_n5212) & (!x449x) & (n_n2665) & (x223x) & (!n_n5211)) + ((n_n5212) & (!x449x) & (n_n2665) & (x223x) & (n_n5211)) + ((n_n5212) & (x449x) & (!n_n2665) & (!x223x) & (!n_n5211)) + ((n_n5212) & (x449x) & (!n_n2665) & (!x223x) & (n_n5211)) + ((n_n5212) & (x449x) & (!n_n2665) & (x223x) & (!n_n5211)) + ((n_n5212) & (x449x) & (!n_n2665) & (x223x) & (n_n5211)) + ((n_n5212) & (x449x) & (n_n2665) & (!x223x) & (!n_n5211)) + ((n_n5212) & (x449x) & (n_n2665) & (!x223x) & (n_n5211)) + ((n_n5212) & (x449x) & (n_n2665) & (x223x) & (!n_n5211)) + ((n_n5212) & (x449x) & (n_n2665) & (x223x) & (n_n5211)));
	assign n_n3301 = (((!n_n5203) & (!x220x) & (!x36x) & (!x450x) & (x14047x)) + ((!n_n5203) & (!x220x) & (!x36x) & (x450x) & (!x14047x)) + ((!n_n5203) & (!x220x) & (!x36x) & (x450x) & (x14047x)) + ((!n_n5203) & (!x220x) & (x36x) & (!x450x) & (!x14047x)) + ((!n_n5203) & (!x220x) & (x36x) & (!x450x) & (x14047x)) + ((!n_n5203) & (!x220x) & (x36x) & (x450x) & (!x14047x)) + ((!n_n5203) & (!x220x) & (x36x) & (x450x) & (x14047x)) + ((!n_n5203) & (x220x) & (!x36x) & (!x450x) & (!x14047x)) + ((!n_n5203) & (x220x) & (!x36x) & (!x450x) & (x14047x)) + ((!n_n5203) & (x220x) & (!x36x) & (x450x) & (!x14047x)) + ((!n_n5203) & (x220x) & (!x36x) & (x450x) & (x14047x)) + ((!n_n5203) & (x220x) & (x36x) & (!x450x) & (!x14047x)) + ((!n_n5203) & (x220x) & (x36x) & (!x450x) & (x14047x)) + ((!n_n5203) & (x220x) & (x36x) & (x450x) & (!x14047x)) + ((!n_n5203) & (x220x) & (x36x) & (x450x) & (x14047x)) + ((n_n5203) & (!x220x) & (!x36x) & (!x450x) & (!x14047x)) + ((n_n5203) & (!x220x) & (!x36x) & (!x450x) & (x14047x)) + ((n_n5203) & (!x220x) & (!x36x) & (x450x) & (!x14047x)) + ((n_n5203) & (!x220x) & (!x36x) & (x450x) & (x14047x)) + ((n_n5203) & (!x220x) & (x36x) & (!x450x) & (!x14047x)) + ((n_n5203) & (!x220x) & (x36x) & (!x450x) & (x14047x)) + ((n_n5203) & (!x220x) & (x36x) & (x450x) & (!x14047x)) + ((n_n5203) & (!x220x) & (x36x) & (x450x) & (x14047x)) + ((n_n5203) & (x220x) & (!x36x) & (!x450x) & (!x14047x)) + ((n_n5203) & (x220x) & (!x36x) & (!x450x) & (x14047x)) + ((n_n5203) & (x220x) & (!x36x) & (x450x) & (!x14047x)) + ((n_n5203) & (x220x) & (!x36x) & (x450x) & (x14047x)) + ((n_n5203) & (x220x) & (x36x) & (!x450x) & (!x14047x)) + ((n_n5203) & (x220x) & (x36x) & (!x450x) & (x14047x)) + ((n_n5203) & (x220x) & (x36x) & (x450x) & (!x14047x)) + ((n_n5203) & (x220x) & (x36x) & (x450x) & (x14047x)));
	assign x14065x = (((!x13924x) & (!x13925x) & (!x13929x) & (!x13930x) & (x14063x)) + ((!x13924x) & (!x13925x) & (!x13929x) & (x13930x) & (!x14063x)) + ((!x13924x) & (!x13925x) & (!x13929x) & (x13930x) & (x14063x)) + ((!x13924x) & (!x13925x) & (x13929x) & (!x13930x) & (!x14063x)) + ((!x13924x) & (!x13925x) & (x13929x) & (!x13930x) & (x14063x)) + ((!x13924x) & (!x13925x) & (x13929x) & (x13930x) & (!x14063x)) + ((!x13924x) & (!x13925x) & (x13929x) & (x13930x) & (x14063x)) + ((!x13924x) & (x13925x) & (!x13929x) & (!x13930x) & (!x14063x)) + ((!x13924x) & (x13925x) & (!x13929x) & (!x13930x) & (x14063x)) + ((!x13924x) & (x13925x) & (!x13929x) & (x13930x) & (!x14063x)) + ((!x13924x) & (x13925x) & (!x13929x) & (x13930x) & (x14063x)) + ((!x13924x) & (x13925x) & (x13929x) & (!x13930x) & (!x14063x)) + ((!x13924x) & (x13925x) & (x13929x) & (!x13930x) & (x14063x)) + ((!x13924x) & (x13925x) & (x13929x) & (x13930x) & (!x14063x)) + ((!x13924x) & (x13925x) & (x13929x) & (x13930x) & (x14063x)) + ((x13924x) & (!x13925x) & (!x13929x) & (!x13930x) & (!x14063x)) + ((x13924x) & (!x13925x) & (!x13929x) & (!x13930x) & (x14063x)) + ((x13924x) & (!x13925x) & (!x13929x) & (x13930x) & (!x14063x)) + ((x13924x) & (!x13925x) & (!x13929x) & (x13930x) & (x14063x)) + ((x13924x) & (!x13925x) & (x13929x) & (!x13930x) & (!x14063x)) + ((x13924x) & (!x13925x) & (x13929x) & (!x13930x) & (x14063x)) + ((x13924x) & (!x13925x) & (x13929x) & (x13930x) & (!x14063x)) + ((x13924x) & (!x13925x) & (x13929x) & (x13930x) & (x14063x)) + ((x13924x) & (x13925x) & (!x13929x) & (!x13930x) & (!x14063x)) + ((x13924x) & (x13925x) & (!x13929x) & (!x13930x) & (x14063x)) + ((x13924x) & (x13925x) & (!x13929x) & (x13930x) & (!x14063x)) + ((x13924x) & (x13925x) & (!x13929x) & (x13930x) & (x14063x)) + ((x13924x) & (x13925x) & (x13929x) & (!x13930x) & (!x14063x)) + ((x13924x) & (x13925x) & (x13929x) & (!x13930x) & (x14063x)) + ((x13924x) & (x13925x) & (x13929x) & (x13930x) & (!x14063x)) + ((x13924x) & (x13925x) & (x13929x) & (x13930x) & (x14063x)));
	assign x14067x = (((!n_n3267) & (!x14057x) & (!n_n3300) & (!n_n3301) & (x14065x)) + ((!n_n3267) & (!x14057x) & (!n_n3300) & (n_n3301) & (!x14065x)) + ((!n_n3267) & (!x14057x) & (!n_n3300) & (n_n3301) & (x14065x)) + ((!n_n3267) & (!x14057x) & (n_n3300) & (!n_n3301) & (!x14065x)) + ((!n_n3267) & (!x14057x) & (n_n3300) & (!n_n3301) & (x14065x)) + ((!n_n3267) & (!x14057x) & (n_n3300) & (n_n3301) & (!x14065x)) + ((!n_n3267) & (!x14057x) & (n_n3300) & (n_n3301) & (x14065x)) + ((!n_n3267) & (x14057x) & (!n_n3300) & (!n_n3301) & (!x14065x)) + ((!n_n3267) & (x14057x) & (!n_n3300) & (!n_n3301) & (x14065x)) + ((!n_n3267) & (x14057x) & (!n_n3300) & (n_n3301) & (!x14065x)) + ((!n_n3267) & (x14057x) & (!n_n3300) & (n_n3301) & (x14065x)) + ((!n_n3267) & (x14057x) & (n_n3300) & (!n_n3301) & (!x14065x)) + ((!n_n3267) & (x14057x) & (n_n3300) & (!n_n3301) & (x14065x)) + ((!n_n3267) & (x14057x) & (n_n3300) & (n_n3301) & (!x14065x)) + ((!n_n3267) & (x14057x) & (n_n3300) & (n_n3301) & (x14065x)) + ((n_n3267) & (!x14057x) & (!n_n3300) & (!n_n3301) & (!x14065x)) + ((n_n3267) & (!x14057x) & (!n_n3300) & (!n_n3301) & (x14065x)) + ((n_n3267) & (!x14057x) & (!n_n3300) & (n_n3301) & (!x14065x)) + ((n_n3267) & (!x14057x) & (!n_n3300) & (n_n3301) & (x14065x)) + ((n_n3267) & (!x14057x) & (n_n3300) & (!n_n3301) & (!x14065x)) + ((n_n3267) & (!x14057x) & (n_n3300) & (!n_n3301) & (x14065x)) + ((n_n3267) & (!x14057x) & (n_n3300) & (n_n3301) & (!x14065x)) + ((n_n3267) & (!x14057x) & (n_n3300) & (n_n3301) & (x14065x)) + ((n_n3267) & (x14057x) & (!n_n3300) & (!n_n3301) & (!x14065x)) + ((n_n3267) & (x14057x) & (!n_n3300) & (!n_n3301) & (x14065x)) + ((n_n3267) & (x14057x) & (!n_n3300) & (n_n3301) & (!x14065x)) + ((n_n3267) & (x14057x) & (!n_n3300) & (n_n3301) & (x14065x)) + ((n_n3267) & (x14057x) & (n_n3300) & (!n_n3301) & (!x14065x)) + ((n_n3267) & (x14057x) & (n_n3300) & (!n_n3301) & (x14065x)) + ((n_n3267) & (x14057x) & (n_n3300) & (n_n3301) & (!x14065x)) + ((n_n3267) & (x14057x) & (n_n3300) & (n_n3301) & (x14065x)));
	assign n_n4334 = (((i_9_) & (n_n536) & (n_n518) & (n_n528)));
	assign n_n3509 = (((!i_9_) & (n_n455) & (!n_n528) & (n_n491) & (n_n530)) + ((!i_9_) & (n_n455) & (n_n528) & (n_n491) & (n_n530)) + ((i_9_) & (n_n455) & (!n_n528) & (n_n491) & (n_n530)) + ((i_9_) & (n_n455) & (n_n528) & (n_n491) & (!n_n530)) + ((i_9_) & (n_n455) & (n_n528) & (n_n491) & (n_n530)));
	assign n_n1646 = (((!x25x) & (!x15x) & (x11x) & (n_n390) & (n_n491)) + ((!x25x) & (x15x) & (!x11x) & (n_n390) & (n_n491)) + ((!x25x) & (x15x) & (x11x) & (n_n390) & (n_n491)) + ((x25x) & (!x15x) & (!x11x) & (n_n390) & (n_n491)) + ((x25x) & (!x15x) & (x11x) & (n_n390) & (n_n491)) + ((x25x) & (x15x) & (!x11x) & (n_n390) & (n_n491)) + ((x25x) & (x15x) & (x11x) & (n_n390) & (n_n491)));
	assign x158x = (((!i_9_) & (n_n473) & (n_n534) & (n_n325)) + ((i_9_) & (n_n473) & (n_n534) & (n_n325)));
	assign x15791x = (((!n_n4790) & (!n_n4791) & (!n_n4787) & (!n_n4795) & (n_n4799)) + ((!n_n4790) & (!n_n4791) & (!n_n4787) & (n_n4795) & (!n_n4799)) + ((!n_n4790) & (!n_n4791) & (!n_n4787) & (n_n4795) & (n_n4799)) + ((!n_n4790) & (!n_n4791) & (n_n4787) & (!n_n4795) & (!n_n4799)) + ((!n_n4790) & (!n_n4791) & (n_n4787) & (!n_n4795) & (n_n4799)) + ((!n_n4790) & (!n_n4791) & (n_n4787) & (n_n4795) & (!n_n4799)) + ((!n_n4790) & (!n_n4791) & (n_n4787) & (n_n4795) & (n_n4799)) + ((!n_n4790) & (n_n4791) & (!n_n4787) & (!n_n4795) & (!n_n4799)) + ((!n_n4790) & (n_n4791) & (!n_n4787) & (!n_n4795) & (n_n4799)) + ((!n_n4790) & (n_n4791) & (!n_n4787) & (n_n4795) & (!n_n4799)) + ((!n_n4790) & (n_n4791) & (!n_n4787) & (n_n4795) & (n_n4799)) + ((!n_n4790) & (n_n4791) & (n_n4787) & (!n_n4795) & (!n_n4799)) + ((!n_n4790) & (n_n4791) & (n_n4787) & (!n_n4795) & (n_n4799)) + ((!n_n4790) & (n_n4791) & (n_n4787) & (n_n4795) & (!n_n4799)) + ((!n_n4790) & (n_n4791) & (n_n4787) & (n_n4795) & (n_n4799)) + ((n_n4790) & (!n_n4791) & (!n_n4787) & (!n_n4795) & (!n_n4799)) + ((n_n4790) & (!n_n4791) & (!n_n4787) & (!n_n4795) & (n_n4799)) + ((n_n4790) & (!n_n4791) & (!n_n4787) & (n_n4795) & (!n_n4799)) + ((n_n4790) & (!n_n4791) & (!n_n4787) & (n_n4795) & (n_n4799)) + ((n_n4790) & (!n_n4791) & (n_n4787) & (!n_n4795) & (!n_n4799)) + ((n_n4790) & (!n_n4791) & (n_n4787) & (!n_n4795) & (n_n4799)) + ((n_n4790) & (!n_n4791) & (n_n4787) & (n_n4795) & (!n_n4799)) + ((n_n4790) & (!n_n4791) & (n_n4787) & (n_n4795) & (n_n4799)) + ((n_n4790) & (n_n4791) & (!n_n4787) & (!n_n4795) & (!n_n4799)) + ((n_n4790) & (n_n4791) & (!n_n4787) & (!n_n4795) & (n_n4799)) + ((n_n4790) & (n_n4791) & (!n_n4787) & (n_n4795) & (!n_n4799)) + ((n_n4790) & (n_n4791) & (!n_n4787) & (n_n4795) & (n_n4799)) + ((n_n4790) & (n_n4791) & (n_n4787) & (!n_n4795) & (!n_n4799)) + ((n_n4790) & (n_n4791) & (n_n4787) & (!n_n4795) & (n_n4799)) + ((n_n4790) & (n_n4791) & (n_n4787) & (n_n4795) & (!n_n4799)) + ((n_n4790) & (n_n4791) & (n_n4787) & (n_n4795) & (n_n4799)));
	assign x48x = (((!i_9_) & (!n_n532) & (n_n534) & (n_n260) & (n_n491)) + ((!i_9_) & (n_n532) & (!n_n534) & (n_n260) & (n_n491)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n260) & (n_n491)) + ((i_9_) & (n_n532) & (!n_n534) & (n_n260) & (n_n491)) + ((i_9_) & (n_n532) & (n_n534) & (n_n260) & (n_n491)));
	assign x383x = (((!x25x) & (x19x) & (n_n518) & (n_n530) & (!n_n65)) + ((!x25x) & (x19x) & (n_n518) & (n_n530) & (n_n65)) + ((x25x) & (!x19x) & (n_n518) & (!n_n530) & (n_n65)) + ((x25x) & (!x19x) & (n_n518) & (n_n530) & (n_n65)) + ((x25x) & (x19x) & (n_n518) & (!n_n530) & (n_n65)) + ((x25x) & (x19x) & (n_n518) & (n_n530) & (!n_n65)) + ((x25x) & (x19x) & (n_n518) & (n_n530) & (n_n65)));
	assign x15208x = (((!i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n518)) + ((!i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n518)));
	assign x15210x = (((!n_n518) & (!x11x) & (!n_n65) & (!n_n5232) & (n_n5233)) + ((!n_n518) & (!x11x) & (!n_n65) & (n_n5232) & (!n_n5233)) + ((!n_n518) & (!x11x) & (!n_n65) & (n_n5232) & (n_n5233)) + ((!n_n518) & (!x11x) & (n_n65) & (!n_n5232) & (n_n5233)) + ((!n_n518) & (!x11x) & (n_n65) & (n_n5232) & (!n_n5233)) + ((!n_n518) & (!x11x) & (n_n65) & (n_n5232) & (n_n5233)) + ((!n_n518) & (x11x) & (!n_n65) & (!n_n5232) & (n_n5233)) + ((!n_n518) & (x11x) & (!n_n65) & (n_n5232) & (!n_n5233)) + ((!n_n518) & (x11x) & (!n_n65) & (n_n5232) & (n_n5233)) + ((!n_n518) & (x11x) & (n_n65) & (!n_n5232) & (n_n5233)) + ((!n_n518) & (x11x) & (n_n65) & (n_n5232) & (!n_n5233)) + ((!n_n518) & (x11x) & (n_n65) & (n_n5232) & (n_n5233)) + ((n_n518) & (!x11x) & (!n_n65) & (!n_n5232) & (n_n5233)) + ((n_n518) & (!x11x) & (!n_n65) & (n_n5232) & (!n_n5233)) + ((n_n518) & (!x11x) & (!n_n65) & (n_n5232) & (n_n5233)) + ((n_n518) & (!x11x) & (n_n65) & (!n_n5232) & (n_n5233)) + ((n_n518) & (!x11x) & (n_n65) & (n_n5232) & (!n_n5233)) + ((n_n518) & (!x11x) & (n_n65) & (n_n5232) & (n_n5233)) + ((n_n518) & (x11x) & (!n_n65) & (!n_n5232) & (n_n5233)) + ((n_n518) & (x11x) & (!n_n65) & (n_n5232) & (!n_n5233)) + ((n_n518) & (x11x) & (!n_n65) & (n_n5232) & (n_n5233)) + ((n_n518) & (x11x) & (n_n65) & (!n_n5232) & (!n_n5233)) + ((n_n518) & (x11x) & (n_n65) & (!n_n5232) & (n_n5233)) + ((n_n518) & (x11x) & (n_n65) & (n_n5232) & (!n_n5233)) + ((n_n518) & (x11x) & (n_n65) & (n_n5232) & (n_n5233)));
	assign n_n2570 = (((!n_n5229) & (!n_n5224) & (!x383x) & (!x15208x) & (x15210x)) + ((!n_n5229) & (!n_n5224) & (!x383x) & (x15208x) & (!x15210x)) + ((!n_n5229) & (!n_n5224) & (!x383x) & (x15208x) & (x15210x)) + ((!n_n5229) & (!n_n5224) & (x383x) & (!x15208x) & (!x15210x)) + ((!n_n5229) & (!n_n5224) & (x383x) & (!x15208x) & (x15210x)) + ((!n_n5229) & (!n_n5224) & (x383x) & (x15208x) & (!x15210x)) + ((!n_n5229) & (!n_n5224) & (x383x) & (x15208x) & (x15210x)) + ((!n_n5229) & (n_n5224) & (!x383x) & (!x15208x) & (!x15210x)) + ((!n_n5229) & (n_n5224) & (!x383x) & (!x15208x) & (x15210x)) + ((!n_n5229) & (n_n5224) & (!x383x) & (x15208x) & (!x15210x)) + ((!n_n5229) & (n_n5224) & (!x383x) & (x15208x) & (x15210x)) + ((!n_n5229) & (n_n5224) & (x383x) & (!x15208x) & (!x15210x)) + ((!n_n5229) & (n_n5224) & (x383x) & (!x15208x) & (x15210x)) + ((!n_n5229) & (n_n5224) & (x383x) & (x15208x) & (!x15210x)) + ((!n_n5229) & (n_n5224) & (x383x) & (x15208x) & (x15210x)) + ((n_n5229) & (!n_n5224) & (!x383x) & (!x15208x) & (!x15210x)) + ((n_n5229) & (!n_n5224) & (!x383x) & (!x15208x) & (x15210x)) + ((n_n5229) & (!n_n5224) & (!x383x) & (x15208x) & (!x15210x)) + ((n_n5229) & (!n_n5224) & (!x383x) & (x15208x) & (x15210x)) + ((n_n5229) & (!n_n5224) & (x383x) & (!x15208x) & (!x15210x)) + ((n_n5229) & (!n_n5224) & (x383x) & (!x15208x) & (x15210x)) + ((n_n5229) & (!n_n5224) & (x383x) & (x15208x) & (!x15210x)) + ((n_n5229) & (!n_n5224) & (x383x) & (x15208x) & (x15210x)) + ((n_n5229) & (n_n5224) & (!x383x) & (!x15208x) & (!x15210x)) + ((n_n5229) & (n_n5224) & (!x383x) & (!x15208x) & (x15210x)) + ((n_n5229) & (n_n5224) & (!x383x) & (x15208x) & (!x15210x)) + ((n_n5229) & (n_n5224) & (!x383x) & (x15208x) & (x15210x)) + ((n_n5229) & (n_n5224) & (x383x) & (!x15208x) & (!x15210x)) + ((n_n5229) & (n_n5224) & (x383x) & (!x15208x) & (x15210x)) + ((n_n5229) & (n_n5224) & (x383x) & (x15208x) & (!x15210x)) + ((n_n5229) & (n_n5224) & (x383x) & (x15208x) & (x15210x)));
	assign n_n5215 = (((!i_9_) & (n_n528) & (n_n535) & (n_n65)));
	assign n_n2665 = (((!i_9_) & (!n_n524) & (!n_n535) & (!n_n65) & (n_n5220)) + ((!i_9_) & (!n_n524) & (!n_n535) & (n_n65) & (n_n5220)) + ((!i_9_) & (!n_n524) & (n_n535) & (!n_n65) & (n_n5220)) + ((!i_9_) & (!n_n524) & (n_n535) & (n_n65) & (n_n5220)) + ((!i_9_) & (n_n524) & (!n_n535) & (!n_n65) & (n_n5220)) + ((!i_9_) & (n_n524) & (!n_n535) & (n_n65) & (n_n5220)) + ((!i_9_) & (n_n524) & (n_n535) & (!n_n65) & (n_n5220)) + ((!i_9_) & (n_n524) & (n_n535) & (n_n65) & (!n_n5220)) + ((!i_9_) & (n_n524) & (n_n535) & (n_n65) & (n_n5220)) + ((i_9_) & (!n_n524) & (!n_n535) & (!n_n65) & (n_n5220)) + ((i_9_) & (!n_n524) & (!n_n535) & (n_n65) & (n_n5220)) + ((i_9_) & (!n_n524) & (n_n535) & (!n_n65) & (n_n5220)) + ((i_9_) & (!n_n524) & (n_n535) & (n_n65) & (n_n5220)) + ((i_9_) & (n_n524) & (!n_n535) & (!n_n65) & (n_n5220)) + ((i_9_) & (n_n524) & (!n_n535) & (n_n65) & (n_n5220)) + ((i_9_) & (n_n524) & (n_n535) & (!n_n65) & (n_n5220)) + ((i_9_) & (n_n524) & (n_n535) & (n_n65) & (!n_n5220)) + ((i_9_) & (n_n524) & (n_n535) & (n_n65) & (n_n5220)));
	assign x220x = (((!n_n522) & (n_n130) & (!x12x) & (x20x) & (n_n464)) + ((!n_n522) & (n_n130) & (x12x) & (x20x) & (n_n464)) + ((n_n522) & (!n_n130) & (x12x) & (!x20x) & (n_n464)) + ((n_n522) & (!n_n130) & (x12x) & (x20x) & (n_n464)) + ((n_n522) & (n_n130) & (!x12x) & (x20x) & (n_n464)) + ((n_n522) & (n_n130) & (x12x) & (!x20x) & (n_n464)) + ((n_n522) & (n_n130) & (x12x) & (x20x) & (n_n464)));
	assign n_n5209 = (((!i_9_) & (n_n534) & (n_n535) & (n_n65)));
	assign x223x = (((!x25x) & (x19x) & (n_n532) & (n_n535) & (!n_n65)) + ((!x25x) & (x19x) & (n_n532) & (n_n535) & (n_n65)) + ((x25x) & (!x19x) & (!n_n532) & (n_n535) & (n_n65)) + ((x25x) & (!x19x) & (n_n532) & (n_n535) & (n_n65)) + ((x25x) & (x19x) & (!n_n532) & (n_n535) & (n_n65)) + ((x25x) & (x19x) & (n_n532) & (n_n535) & (!n_n65)) + ((x25x) & (x19x) & (n_n532) & (n_n535) & (n_n65)));
	assign x384x = (((n_n535) & (!x20x) & (x23x) & (n_n65)) + ((n_n535) & (x20x) & (!x23x) & (n_n65)) + ((n_n535) & (x20x) & (x23x) & (n_n65)));
	assign n_n5213 = (((!i_9_) & (n_n535) & (n_n530) & (n_n65)));
	assign x454x = (((!i_9_) & (!n_n532) & (n_n535) & (n_n530) & (n_n65)) + ((!i_9_) & (n_n532) & (n_n535) & (!n_n530) & (n_n65)) + ((!i_9_) & (n_n532) & (n_n535) & (n_n530) & (n_n65)));
	assign x22095x = (((!n_n5206) & (!n_n5216) & (!n_n5222) & (!n_n5217) & (!n_n5215)));
	assign x15221x = (((!n_n5214) & (!n_n5207) & (!n_n2665) & (!x22095x)) + ((!n_n5214) & (!n_n5207) & (n_n2665) & (!x22095x)) + ((!n_n5214) & (!n_n5207) & (n_n2665) & (x22095x)) + ((!n_n5214) & (n_n5207) & (!n_n2665) & (!x22095x)) + ((!n_n5214) & (n_n5207) & (!n_n2665) & (x22095x)) + ((!n_n5214) & (n_n5207) & (n_n2665) & (!x22095x)) + ((!n_n5214) & (n_n5207) & (n_n2665) & (x22095x)) + ((n_n5214) & (!n_n5207) & (!n_n2665) & (!x22095x)) + ((n_n5214) & (!n_n5207) & (!n_n2665) & (x22095x)) + ((n_n5214) & (!n_n5207) & (n_n2665) & (!x22095x)) + ((n_n5214) & (!n_n5207) & (n_n2665) & (x22095x)) + ((n_n5214) & (n_n5207) & (!n_n2665) & (!x22095x)) + ((n_n5214) & (n_n5207) & (!n_n2665) & (x22095x)) + ((n_n5214) & (n_n5207) & (n_n2665) & (!x22095x)) + ((n_n5214) & (n_n5207) & (n_n2665) & (x22095x)));
	assign x15220x = (((!n_n5204) & (!n_n5205) & (!x223x) & (!x384x) & (x454x)) + ((!n_n5204) & (!n_n5205) & (!x223x) & (x384x) & (!x454x)) + ((!n_n5204) & (!n_n5205) & (!x223x) & (x384x) & (x454x)) + ((!n_n5204) & (!n_n5205) & (x223x) & (!x384x) & (!x454x)) + ((!n_n5204) & (!n_n5205) & (x223x) & (!x384x) & (x454x)) + ((!n_n5204) & (!n_n5205) & (x223x) & (x384x) & (!x454x)) + ((!n_n5204) & (!n_n5205) & (x223x) & (x384x) & (x454x)) + ((!n_n5204) & (n_n5205) & (!x223x) & (!x384x) & (!x454x)) + ((!n_n5204) & (n_n5205) & (!x223x) & (!x384x) & (x454x)) + ((!n_n5204) & (n_n5205) & (!x223x) & (x384x) & (!x454x)) + ((!n_n5204) & (n_n5205) & (!x223x) & (x384x) & (x454x)) + ((!n_n5204) & (n_n5205) & (x223x) & (!x384x) & (!x454x)) + ((!n_n5204) & (n_n5205) & (x223x) & (!x384x) & (x454x)) + ((!n_n5204) & (n_n5205) & (x223x) & (x384x) & (!x454x)) + ((!n_n5204) & (n_n5205) & (x223x) & (x384x) & (x454x)) + ((n_n5204) & (!n_n5205) & (!x223x) & (!x384x) & (!x454x)) + ((n_n5204) & (!n_n5205) & (!x223x) & (!x384x) & (x454x)) + ((n_n5204) & (!n_n5205) & (!x223x) & (x384x) & (!x454x)) + ((n_n5204) & (!n_n5205) & (!x223x) & (x384x) & (x454x)) + ((n_n5204) & (!n_n5205) & (x223x) & (!x384x) & (!x454x)) + ((n_n5204) & (!n_n5205) & (x223x) & (!x384x) & (x454x)) + ((n_n5204) & (!n_n5205) & (x223x) & (x384x) & (!x454x)) + ((n_n5204) & (!n_n5205) & (x223x) & (x384x) & (x454x)) + ((n_n5204) & (n_n5205) & (!x223x) & (!x384x) & (!x454x)) + ((n_n5204) & (n_n5205) & (!x223x) & (!x384x) & (x454x)) + ((n_n5204) & (n_n5205) & (!x223x) & (x384x) & (!x454x)) + ((n_n5204) & (n_n5205) & (!x223x) & (x384x) & (x454x)) + ((n_n5204) & (n_n5205) & (x223x) & (!x384x) & (!x454x)) + ((n_n5204) & (n_n5205) & (x223x) & (!x384x) & (x454x)) + ((n_n5204) & (n_n5205) & (x223x) & (x384x) & (!x454x)) + ((n_n5204) & (n_n5205) & (x223x) & (x384x) & (x454x)));
	assign n_n4534 = (((i_9_) & (n_n482) & (n_n455) & (n_n520)));
	assign x15061x = (((!n_n4547) & (!n_n4539) & (!n_n4544) & (n_n4538)) + ((!n_n4547) & (!n_n4539) & (n_n4544) & (!n_n4538)) + ((!n_n4547) & (!n_n4539) & (n_n4544) & (n_n4538)) + ((!n_n4547) & (n_n4539) & (!n_n4544) & (!n_n4538)) + ((!n_n4547) & (n_n4539) & (!n_n4544) & (n_n4538)) + ((!n_n4547) & (n_n4539) & (n_n4544) & (!n_n4538)) + ((!n_n4547) & (n_n4539) & (n_n4544) & (n_n4538)) + ((n_n4547) & (!n_n4539) & (!n_n4544) & (!n_n4538)) + ((n_n4547) & (!n_n4539) & (!n_n4544) & (n_n4538)) + ((n_n4547) & (!n_n4539) & (n_n4544) & (!n_n4538)) + ((n_n4547) & (!n_n4539) & (n_n4544) & (n_n4538)) + ((n_n4547) & (n_n4539) & (!n_n4544) & (!n_n4538)) + ((n_n4547) & (n_n4539) & (!n_n4544) & (n_n4538)) + ((n_n4547) & (n_n4539) & (n_n4544) & (!n_n4538)) + ((n_n4547) & (n_n4539) & (n_n4544) & (n_n4538)));
	assign x15062x = (((!n_n4535) & (!n_n4536) & (!n_n4541) & (!n_n4543) & (n_n4537)) + ((!n_n4535) & (!n_n4536) & (!n_n4541) & (n_n4543) & (!n_n4537)) + ((!n_n4535) & (!n_n4536) & (!n_n4541) & (n_n4543) & (n_n4537)) + ((!n_n4535) & (!n_n4536) & (n_n4541) & (!n_n4543) & (!n_n4537)) + ((!n_n4535) & (!n_n4536) & (n_n4541) & (!n_n4543) & (n_n4537)) + ((!n_n4535) & (!n_n4536) & (n_n4541) & (n_n4543) & (!n_n4537)) + ((!n_n4535) & (!n_n4536) & (n_n4541) & (n_n4543) & (n_n4537)) + ((!n_n4535) & (n_n4536) & (!n_n4541) & (!n_n4543) & (!n_n4537)) + ((!n_n4535) & (n_n4536) & (!n_n4541) & (!n_n4543) & (n_n4537)) + ((!n_n4535) & (n_n4536) & (!n_n4541) & (n_n4543) & (!n_n4537)) + ((!n_n4535) & (n_n4536) & (!n_n4541) & (n_n4543) & (n_n4537)) + ((!n_n4535) & (n_n4536) & (n_n4541) & (!n_n4543) & (!n_n4537)) + ((!n_n4535) & (n_n4536) & (n_n4541) & (!n_n4543) & (n_n4537)) + ((!n_n4535) & (n_n4536) & (n_n4541) & (n_n4543) & (!n_n4537)) + ((!n_n4535) & (n_n4536) & (n_n4541) & (n_n4543) & (n_n4537)) + ((n_n4535) & (!n_n4536) & (!n_n4541) & (!n_n4543) & (!n_n4537)) + ((n_n4535) & (!n_n4536) & (!n_n4541) & (!n_n4543) & (n_n4537)) + ((n_n4535) & (!n_n4536) & (!n_n4541) & (n_n4543) & (!n_n4537)) + ((n_n4535) & (!n_n4536) & (!n_n4541) & (n_n4543) & (n_n4537)) + ((n_n4535) & (!n_n4536) & (n_n4541) & (!n_n4543) & (!n_n4537)) + ((n_n4535) & (!n_n4536) & (n_n4541) & (!n_n4543) & (n_n4537)) + ((n_n4535) & (!n_n4536) & (n_n4541) & (n_n4543) & (!n_n4537)) + ((n_n4535) & (!n_n4536) & (n_n4541) & (n_n4543) & (n_n4537)) + ((n_n4535) & (n_n4536) & (!n_n4541) & (!n_n4543) & (!n_n4537)) + ((n_n4535) & (n_n4536) & (!n_n4541) & (!n_n4543) & (n_n4537)) + ((n_n4535) & (n_n4536) & (!n_n4541) & (n_n4543) & (!n_n4537)) + ((n_n4535) & (n_n4536) & (!n_n4541) & (n_n4543) & (n_n4537)) + ((n_n4535) & (n_n4536) & (n_n4541) & (!n_n4543) & (!n_n4537)) + ((n_n4535) & (n_n4536) & (n_n4541) & (!n_n4543) & (n_n4537)) + ((n_n4535) & (n_n4536) & (n_n4541) & (n_n4543) & (!n_n4537)) + ((n_n4535) & (n_n4536) & (n_n4541) & (n_n4543) & (n_n4537)));
	assign x15074x = (((!n_n536) & (!x23x) & (!n_n464) & (!n_n4443) & (n_n910)) + ((!n_n536) & (!x23x) & (!n_n464) & (n_n4443) & (!n_n910)) + ((!n_n536) & (!x23x) & (!n_n464) & (n_n4443) & (n_n910)) + ((!n_n536) & (!x23x) & (n_n464) & (!n_n4443) & (n_n910)) + ((!n_n536) & (!x23x) & (n_n464) & (n_n4443) & (!n_n910)) + ((!n_n536) & (!x23x) & (n_n464) & (n_n4443) & (n_n910)) + ((!n_n536) & (x23x) & (!n_n464) & (!n_n4443) & (n_n910)) + ((!n_n536) & (x23x) & (!n_n464) & (n_n4443) & (!n_n910)) + ((!n_n536) & (x23x) & (!n_n464) & (n_n4443) & (n_n910)) + ((!n_n536) & (x23x) & (n_n464) & (!n_n4443) & (n_n910)) + ((!n_n536) & (x23x) & (n_n464) & (n_n4443) & (!n_n910)) + ((!n_n536) & (x23x) & (n_n464) & (n_n4443) & (n_n910)) + ((n_n536) & (!x23x) & (!n_n464) & (!n_n4443) & (n_n910)) + ((n_n536) & (!x23x) & (!n_n464) & (n_n4443) & (!n_n910)) + ((n_n536) & (!x23x) & (!n_n464) & (n_n4443) & (n_n910)) + ((n_n536) & (!x23x) & (n_n464) & (!n_n4443) & (n_n910)) + ((n_n536) & (!x23x) & (n_n464) & (n_n4443) & (!n_n910)) + ((n_n536) & (!x23x) & (n_n464) & (n_n4443) & (n_n910)) + ((n_n536) & (x23x) & (!n_n464) & (!n_n4443) & (n_n910)) + ((n_n536) & (x23x) & (!n_n464) & (n_n4443) & (!n_n910)) + ((n_n536) & (x23x) & (!n_n464) & (n_n4443) & (n_n910)) + ((n_n536) & (x23x) & (n_n464) & (!n_n4443) & (!n_n910)) + ((n_n536) & (x23x) & (n_n464) & (!n_n4443) & (n_n910)) + ((n_n536) & (x23x) & (n_n464) & (n_n4443) & (!n_n910)) + ((n_n536) & (x23x) & (n_n464) & (n_n4443) & (n_n910)));
	assign x15075x = (((!x236x) & (!n_n4445) & (!n_n4441) & (x15074x)) + ((!x236x) & (!n_n4445) & (n_n4441) & (!x15074x)) + ((!x236x) & (!n_n4445) & (n_n4441) & (x15074x)) + ((!x236x) & (n_n4445) & (!n_n4441) & (!x15074x)) + ((!x236x) & (n_n4445) & (!n_n4441) & (x15074x)) + ((!x236x) & (n_n4445) & (n_n4441) & (!x15074x)) + ((!x236x) & (n_n4445) & (n_n4441) & (x15074x)) + ((x236x) & (!n_n4445) & (!n_n4441) & (!x15074x)) + ((x236x) & (!n_n4445) & (!n_n4441) & (x15074x)) + ((x236x) & (!n_n4445) & (n_n4441) & (!x15074x)) + ((x236x) & (!n_n4445) & (n_n4441) & (x15074x)) + ((x236x) & (n_n4445) & (!n_n4441) & (!x15074x)) + ((x236x) & (n_n4445) & (!n_n4441) & (x15074x)) + ((x236x) & (n_n4445) & (n_n4441) & (!x15074x)) + ((x236x) & (n_n4445) & (n_n4441) & (x15074x)));
	assign x128x = (((!i_9_) & (n_n455) & (n_n535) & (!n_n520) & (x23x)) + ((!i_9_) & (n_n455) & (n_n535) & (n_n520) & (x23x)) + ((i_9_) & (n_n455) & (n_n535) & (!n_n520) & (x23x)) + ((i_9_) & (n_n455) & (n_n535) & (n_n520) & (!x23x)) + ((i_9_) & (n_n455) & (n_n535) & (n_n520) & (x23x)));
	assign x291x = (((!i_9_) & (n_n518) & (n_n455) & (!n_n532) & (n_n530)) + ((!i_9_) & (n_n518) & (n_n455) & (n_n532) & (!n_n530)) + ((!i_9_) & (n_n518) & (n_n455) & (n_n532) & (n_n530)));
	assign x15066x = (((!x368x) & (!n_n4456) & (!n_n4458) & (n_n4446)) + ((!x368x) & (!n_n4456) & (n_n4458) & (!n_n4446)) + ((!x368x) & (!n_n4456) & (n_n4458) & (n_n4446)) + ((!x368x) & (n_n4456) & (!n_n4458) & (!n_n4446)) + ((!x368x) & (n_n4456) & (!n_n4458) & (n_n4446)) + ((!x368x) & (n_n4456) & (n_n4458) & (!n_n4446)) + ((!x368x) & (n_n4456) & (n_n4458) & (n_n4446)) + ((x368x) & (!n_n4456) & (!n_n4458) & (!n_n4446)) + ((x368x) & (!n_n4456) & (!n_n4458) & (n_n4446)) + ((x368x) & (!n_n4456) & (n_n4458) & (!n_n4446)) + ((x368x) & (!n_n4456) & (n_n4458) & (n_n4446)) + ((x368x) & (n_n4456) & (!n_n4458) & (!n_n4446)) + ((x368x) & (n_n4456) & (!n_n4458) & (n_n4446)) + ((x368x) & (n_n4456) & (n_n4458) & (!n_n4446)) + ((x368x) & (n_n4456) & (n_n4458) & (n_n4446)));
	assign n_n2630 = (((!n_n4466) & (!x412x) & (!n_n4465) & (!n_n4462) & (!x22224x)) + ((!n_n4466) & (!x412x) & (!n_n4465) & (n_n4462) & (!x22224x)) + ((!n_n4466) & (!x412x) & (!n_n4465) & (n_n4462) & (x22224x)) + ((!n_n4466) & (!x412x) & (n_n4465) & (!n_n4462) & (!x22224x)) + ((!n_n4466) & (!x412x) & (n_n4465) & (!n_n4462) & (x22224x)) + ((!n_n4466) & (!x412x) & (n_n4465) & (n_n4462) & (!x22224x)) + ((!n_n4466) & (!x412x) & (n_n4465) & (n_n4462) & (x22224x)) + ((!n_n4466) & (x412x) & (!n_n4465) & (!n_n4462) & (!x22224x)) + ((!n_n4466) & (x412x) & (!n_n4465) & (!n_n4462) & (x22224x)) + ((!n_n4466) & (x412x) & (!n_n4465) & (n_n4462) & (!x22224x)) + ((!n_n4466) & (x412x) & (!n_n4465) & (n_n4462) & (x22224x)) + ((!n_n4466) & (x412x) & (n_n4465) & (!n_n4462) & (!x22224x)) + ((!n_n4466) & (x412x) & (n_n4465) & (!n_n4462) & (x22224x)) + ((!n_n4466) & (x412x) & (n_n4465) & (n_n4462) & (!x22224x)) + ((!n_n4466) & (x412x) & (n_n4465) & (n_n4462) & (x22224x)) + ((n_n4466) & (!x412x) & (!n_n4465) & (!n_n4462) & (!x22224x)) + ((n_n4466) & (!x412x) & (!n_n4465) & (!n_n4462) & (x22224x)) + ((n_n4466) & (!x412x) & (!n_n4465) & (n_n4462) & (!x22224x)) + ((n_n4466) & (!x412x) & (!n_n4465) & (n_n4462) & (x22224x)) + ((n_n4466) & (!x412x) & (n_n4465) & (!n_n4462) & (!x22224x)) + ((n_n4466) & (!x412x) & (n_n4465) & (!n_n4462) & (x22224x)) + ((n_n4466) & (!x412x) & (n_n4465) & (n_n4462) & (!x22224x)) + ((n_n4466) & (!x412x) & (n_n4465) & (n_n4462) & (x22224x)) + ((n_n4466) & (x412x) & (!n_n4465) & (!n_n4462) & (!x22224x)) + ((n_n4466) & (x412x) & (!n_n4465) & (!n_n4462) & (x22224x)) + ((n_n4466) & (x412x) & (!n_n4465) & (n_n4462) & (!x22224x)) + ((n_n4466) & (x412x) & (!n_n4465) & (n_n4462) & (x22224x)) + ((n_n4466) & (x412x) & (n_n4465) & (!n_n4462) & (!x22224x)) + ((n_n4466) & (x412x) & (n_n4465) & (!n_n4462) & (x22224x)) + ((n_n4466) & (x412x) & (n_n4465) & (n_n4462) & (!x22224x)) + ((n_n4466) & (x412x) & (n_n4465) & (n_n4462) & (x22224x)));
	assign n_n2558 = (((!x15075x) & (!x128x) & (!x291x) & (!x15066x) & (n_n2630)) + ((!x15075x) & (!x128x) & (!x291x) & (x15066x) & (!n_n2630)) + ((!x15075x) & (!x128x) & (!x291x) & (x15066x) & (n_n2630)) + ((!x15075x) & (!x128x) & (x291x) & (!x15066x) & (!n_n2630)) + ((!x15075x) & (!x128x) & (x291x) & (!x15066x) & (n_n2630)) + ((!x15075x) & (!x128x) & (x291x) & (x15066x) & (!n_n2630)) + ((!x15075x) & (!x128x) & (x291x) & (x15066x) & (n_n2630)) + ((!x15075x) & (x128x) & (!x291x) & (!x15066x) & (!n_n2630)) + ((!x15075x) & (x128x) & (!x291x) & (!x15066x) & (n_n2630)) + ((!x15075x) & (x128x) & (!x291x) & (x15066x) & (!n_n2630)) + ((!x15075x) & (x128x) & (!x291x) & (x15066x) & (n_n2630)) + ((!x15075x) & (x128x) & (x291x) & (!x15066x) & (!n_n2630)) + ((!x15075x) & (x128x) & (x291x) & (!x15066x) & (n_n2630)) + ((!x15075x) & (x128x) & (x291x) & (x15066x) & (!n_n2630)) + ((!x15075x) & (x128x) & (x291x) & (x15066x) & (n_n2630)) + ((x15075x) & (!x128x) & (!x291x) & (!x15066x) & (!n_n2630)) + ((x15075x) & (!x128x) & (!x291x) & (!x15066x) & (n_n2630)) + ((x15075x) & (!x128x) & (!x291x) & (x15066x) & (!n_n2630)) + ((x15075x) & (!x128x) & (!x291x) & (x15066x) & (n_n2630)) + ((x15075x) & (!x128x) & (x291x) & (!x15066x) & (!n_n2630)) + ((x15075x) & (!x128x) & (x291x) & (!x15066x) & (n_n2630)) + ((x15075x) & (!x128x) & (x291x) & (x15066x) & (!n_n2630)) + ((x15075x) & (!x128x) & (x291x) & (x15066x) & (n_n2630)) + ((x15075x) & (x128x) & (!x291x) & (!x15066x) & (!n_n2630)) + ((x15075x) & (x128x) & (!x291x) & (!x15066x) & (n_n2630)) + ((x15075x) & (x128x) & (!x291x) & (x15066x) & (!n_n2630)) + ((x15075x) & (x128x) & (!x291x) & (x15066x) & (n_n2630)) + ((x15075x) & (x128x) & (x291x) & (!x15066x) & (!n_n2630)) + ((x15075x) & (x128x) & (x291x) & (!x15066x) & (n_n2630)) + ((x15075x) & (x128x) & (x291x) & (x15066x) & (!n_n2630)) + ((x15075x) & (x128x) & (x291x) & (x15066x) & (n_n2630)));
	assign x307x = (((!n_n455) & (!n_n491) & (!x23x) & (n_n4520)) + ((!n_n455) & (!n_n491) & (x23x) & (n_n4520)) + ((!n_n455) & (n_n491) & (!x23x) & (n_n4520)) + ((!n_n455) & (n_n491) & (x23x) & (n_n4520)) + ((n_n455) & (!n_n491) & (!x23x) & (n_n4520)) + ((n_n455) & (!n_n491) & (x23x) & (n_n4520)) + ((n_n455) & (n_n491) & (!x23x) & (n_n4520)) + ((n_n455) & (n_n491) & (x23x) & (!n_n4520)) + ((n_n455) & (n_n491) & (x23x) & (n_n4520)));
	assign x15080x = (((!n_n524) & (!n_n526) & (!x13x) & (!n_n491) & (x307x)) + ((!n_n524) & (!n_n526) & (!x13x) & (n_n491) & (x307x)) + ((!n_n524) & (!n_n526) & (x13x) & (!n_n491) & (x307x)) + ((!n_n524) & (!n_n526) & (x13x) & (n_n491) & (x307x)) + ((!n_n524) & (n_n526) & (!x13x) & (!n_n491) & (x307x)) + ((!n_n524) & (n_n526) & (!x13x) & (n_n491) & (x307x)) + ((!n_n524) & (n_n526) & (x13x) & (!n_n491) & (x307x)) + ((!n_n524) & (n_n526) & (x13x) & (n_n491) & (!x307x)) + ((!n_n524) & (n_n526) & (x13x) & (n_n491) & (x307x)) + ((n_n524) & (!n_n526) & (!x13x) & (!n_n491) & (x307x)) + ((n_n524) & (!n_n526) & (!x13x) & (n_n491) & (x307x)) + ((n_n524) & (!n_n526) & (x13x) & (!n_n491) & (x307x)) + ((n_n524) & (!n_n526) & (x13x) & (n_n491) & (!x307x)) + ((n_n524) & (!n_n526) & (x13x) & (n_n491) & (x307x)) + ((n_n524) & (n_n526) & (!x13x) & (!n_n491) & (x307x)) + ((n_n524) & (n_n526) & (!x13x) & (n_n491) & (x307x)) + ((n_n524) & (n_n526) & (x13x) & (!n_n491) & (x307x)) + ((n_n524) & (n_n526) & (x13x) & (n_n491) & (!x307x)) + ((n_n524) & (n_n526) & (x13x) & (n_n491) & (x307x)));
	assign x15081x = (((!x130x) & (!n_n4521) & (!n_n4511) & (n_n4518)) + ((!x130x) & (!n_n4521) & (n_n4511) & (!n_n4518)) + ((!x130x) & (!n_n4521) & (n_n4511) & (n_n4518)) + ((!x130x) & (n_n4521) & (!n_n4511) & (!n_n4518)) + ((!x130x) & (n_n4521) & (!n_n4511) & (n_n4518)) + ((!x130x) & (n_n4521) & (n_n4511) & (!n_n4518)) + ((!x130x) & (n_n4521) & (n_n4511) & (n_n4518)) + ((x130x) & (!n_n4521) & (!n_n4511) & (!n_n4518)) + ((x130x) & (!n_n4521) & (!n_n4511) & (n_n4518)) + ((x130x) & (!n_n4521) & (n_n4511) & (!n_n4518)) + ((x130x) & (!n_n4521) & (n_n4511) & (n_n4518)) + ((x130x) & (n_n4521) & (!n_n4511) & (!n_n4518)) + ((x130x) & (n_n4521) & (!n_n4511) & (n_n4518)) + ((x130x) & (n_n4521) & (n_n4511) & (!n_n4518)) + ((x130x) & (n_n4521) & (n_n4511) & (n_n4518)));
	assign n_n1677 = (((!n_n455) & (!n_n509) & (!x23x) & (!n_n4488) & (n_n4486)) + ((!n_n455) & (!n_n509) & (!x23x) & (n_n4488) & (!n_n4486)) + ((!n_n455) & (!n_n509) & (!x23x) & (n_n4488) & (n_n4486)) + ((!n_n455) & (!n_n509) & (x23x) & (!n_n4488) & (n_n4486)) + ((!n_n455) & (!n_n509) & (x23x) & (n_n4488) & (!n_n4486)) + ((!n_n455) & (!n_n509) & (x23x) & (n_n4488) & (n_n4486)) + ((!n_n455) & (n_n509) & (!x23x) & (!n_n4488) & (n_n4486)) + ((!n_n455) & (n_n509) & (!x23x) & (n_n4488) & (!n_n4486)) + ((!n_n455) & (n_n509) & (!x23x) & (n_n4488) & (n_n4486)) + ((!n_n455) & (n_n509) & (x23x) & (!n_n4488) & (n_n4486)) + ((!n_n455) & (n_n509) & (x23x) & (n_n4488) & (!n_n4486)) + ((!n_n455) & (n_n509) & (x23x) & (n_n4488) & (n_n4486)) + ((n_n455) & (!n_n509) & (!x23x) & (!n_n4488) & (n_n4486)) + ((n_n455) & (!n_n509) & (!x23x) & (n_n4488) & (!n_n4486)) + ((n_n455) & (!n_n509) & (!x23x) & (n_n4488) & (n_n4486)) + ((n_n455) & (!n_n509) & (x23x) & (!n_n4488) & (n_n4486)) + ((n_n455) & (!n_n509) & (x23x) & (n_n4488) & (!n_n4486)) + ((n_n455) & (!n_n509) & (x23x) & (n_n4488) & (n_n4486)) + ((n_n455) & (n_n509) & (!x23x) & (!n_n4488) & (n_n4486)) + ((n_n455) & (n_n509) & (!x23x) & (n_n4488) & (!n_n4486)) + ((n_n455) & (n_n509) & (!x23x) & (n_n4488) & (n_n4486)) + ((n_n455) & (n_n509) & (x23x) & (!n_n4488) & (!n_n4486)) + ((n_n455) & (n_n509) & (x23x) & (!n_n4488) & (n_n4486)) + ((n_n455) & (n_n509) & (x23x) & (n_n4488) & (!n_n4486)) + ((n_n455) & (n_n509) & (x23x) & (n_n4488) & (n_n4486)));
	assign n_n2629 = (((!x70x) & (!n_n3515) & (!n_n4474) & (!n_n4484) & (x15082x)) + ((!x70x) & (!n_n3515) & (!n_n4474) & (n_n4484) & (!x15082x)) + ((!x70x) & (!n_n3515) & (!n_n4474) & (n_n4484) & (x15082x)) + ((!x70x) & (!n_n3515) & (n_n4474) & (!n_n4484) & (!x15082x)) + ((!x70x) & (!n_n3515) & (n_n4474) & (!n_n4484) & (x15082x)) + ((!x70x) & (!n_n3515) & (n_n4474) & (n_n4484) & (!x15082x)) + ((!x70x) & (!n_n3515) & (n_n4474) & (n_n4484) & (x15082x)) + ((!x70x) & (n_n3515) & (!n_n4474) & (!n_n4484) & (!x15082x)) + ((!x70x) & (n_n3515) & (!n_n4474) & (!n_n4484) & (x15082x)) + ((!x70x) & (n_n3515) & (!n_n4474) & (n_n4484) & (!x15082x)) + ((!x70x) & (n_n3515) & (!n_n4474) & (n_n4484) & (x15082x)) + ((!x70x) & (n_n3515) & (n_n4474) & (!n_n4484) & (!x15082x)) + ((!x70x) & (n_n3515) & (n_n4474) & (!n_n4484) & (x15082x)) + ((!x70x) & (n_n3515) & (n_n4474) & (n_n4484) & (!x15082x)) + ((!x70x) & (n_n3515) & (n_n4474) & (n_n4484) & (x15082x)) + ((x70x) & (!n_n3515) & (!n_n4474) & (!n_n4484) & (!x15082x)) + ((x70x) & (!n_n3515) & (!n_n4474) & (!n_n4484) & (x15082x)) + ((x70x) & (!n_n3515) & (!n_n4474) & (n_n4484) & (!x15082x)) + ((x70x) & (!n_n3515) & (!n_n4474) & (n_n4484) & (x15082x)) + ((x70x) & (!n_n3515) & (n_n4474) & (!n_n4484) & (!x15082x)) + ((x70x) & (!n_n3515) & (n_n4474) & (!n_n4484) & (x15082x)) + ((x70x) & (!n_n3515) & (n_n4474) & (n_n4484) & (!x15082x)) + ((x70x) & (!n_n3515) & (n_n4474) & (n_n4484) & (x15082x)) + ((x70x) & (n_n3515) & (!n_n4474) & (!n_n4484) & (!x15082x)) + ((x70x) & (n_n3515) & (!n_n4474) & (!n_n4484) & (x15082x)) + ((x70x) & (n_n3515) & (!n_n4474) & (n_n4484) & (!x15082x)) + ((x70x) & (n_n3515) & (!n_n4474) & (n_n4484) & (x15082x)) + ((x70x) & (n_n3515) & (n_n4474) & (!n_n4484) & (!x15082x)) + ((x70x) & (n_n3515) & (n_n4474) & (!n_n4484) & (x15082x)) + ((x70x) & (n_n3515) & (n_n4474) & (n_n4484) & (!x15082x)) + ((x70x) & (n_n3515) & (n_n4474) & (n_n4484) & (x15082x)));
	assign x15091x = (((!n_n4505) & (!n_n4492) & (!n_n4507) & (n_n4501)) + ((!n_n4505) & (!n_n4492) & (n_n4507) & (!n_n4501)) + ((!n_n4505) & (!n_n4492) & (n_n4507) & (n_n4501)) + ((!n_n4505) & (n_n4492) & (!n_n4507) & (!n_n4501)) + ((!n_n4505) & (n_n4492) & (!n_n4507) & (n_n4501)) + ((!n_n4505) & (n_n4492) & (n_n4507) & (!n_n4501)) + ((!n_n4505) & (n_n4492) & (n_n4507) & (n_n4501)) + ((n_n4505) & (!n_n4492) & (!n_n4507) & (!n_n4501)) + ((n_n4505) & (!n_n4492) & (!n_n4507) & (n_n4501)) + ((n_n4505) & (!n_n4492) & (n_n4507) & (!n_n4501)) + ((n_n4505) & (!n_n4492) & (n_n4507) & (n_n4501)) + ((n_n4505) & (n_n4492) & (!n_n4507) & (!n_n4501)) + ((n_n4505) & (n_n4492) & (!n_n4507) & (n_n4501)) + ((n_n4505) & (n_n4492) & (n_n4507) & (!n_n4501)) + ((n_n4505) & (n_n4492) & (n_n4507) & (n_n4501)));
	assign x15093x = (((!n_n4497) & (!x428x) & (!x65x) & (!n_n4502) & (x347x)) + ((!n_n4497) & (!x428x) & (!x65x) & (n_n4502) & (!x347x)) + ((!n_n4497) & (!x428x) & (!x65x) & (n_n4502) & (x347x)) + ((!n_n4497) & (!x428x) & (x65x) & (!n_n4502) & (!x347x)) + ((!n_n4497) & (!x428x) & (x65x) & (!n_n4502) & (x347x)) + ((!n_n4497) & (!x428x) & (x65x) & (n_n4502) & (!x347x)) + ((!n_n4497) & (!x428x) & (x65x) & (n_n4502) & (x347x)) + ((!n_n4497) & (x428x) & (!x65x) & (!n_n4502) & (!x347x)) + ((!n_n4497) & (x428x) & (!x65x) & (!n_n4502) & (x347x)) + ((!n_n4497) & (x428x) & (!x65x) & (n_n4502) & (!x347x)) + ((!n_n4497) & (x428x) & (!x65x) & (n_n4502) & (x347x)) + ((!n_n4497) & (x428x) & (x65x) & (!n_n4502) & (!x347x)) + ((!n_n4497) & (x428x) & (x65x) & (!n_n4502) & (x347x)) + ((!n_n4497) & (x428x) & (x65x) & (n_n4502) & (!x347x)) + ((!n_n4497) & (x428x) & (x65x) & (n_n4502) & (x347x)) + ((n_n4497) & (!x428x) & (!x65x) & (!n_n4502) & (!x347x)) + ((n_n4497) & (!x428x) & (!x65x) & (!n_n4502) & (x347x)) + ((n_n4497) & (!x428x) & (!x65x) & (n_n4502) & (!x347x)) + ((n_n4497) & (!x428x) & (!x65x) & (n_n4502) & (x347x)) + ((n_n4497) & (!x428x) & (x65x) & (!n_n4502) & (!x347x)) + ((n_n4497) & (!x428x) & (x65x) & (!n_n4502) & (x347x)) + ((n_n4497) & (!x428x) & (x65x) & (n_n4502) & (!x347x)) + ((n_n4497) & (!x428x) & (x65x) & (n_n4502) & (x347x)) + ((n_n4497) & (x428x) & (!x65x) & (!n_n4502) & (!x347x)) + ((n_n4497) & (x428x) & (!x65x) & (!n_n4502) & (x347x)) + ((n_n4497) & (x428x) & (!x65x) & (n_n4502) & (!x347x)) + ((n_n4497) & (x428x) & (!x65x) & (n_n4502) & (x347x)) + ((n_n4497) & (x428x) & (x65x) & (!n_n4502) & (!x347x)) + ((n_n4497) & (x428x) & (x65x) & (!n_n4502) & (x347x)) + ((n_n4497) & (x428x) & (x65x) & (n_n4502) & (!x347x)) + ((n_n4497) & (x428x) & (x65x) & (n_n4502) & (x347x)));
	assign n_n2557 = (((!n_n3509) & (!n_n1677) & (!n_n2629) & (!x15091x) & (x15093x)) + ((!n_n3509) & (!n_n1677) & (!n_n2629) & (x15091x) & (!x15093x)) + ((!n_n3509) & (!n_n1677) & (!n_n2629) & (x15091x) & (x15093x)) + ((!n_n3509) & (!n_n1677) & (n_n2629) & (!x15091x) & (!x15093x)) + ((!n_n3509) & (!n_n1677) & (n_n2629) & (!x15091x) & (x15093x)) + ((!n_n3509) & (!n_n1677) & (n_n2629) & (x15091x) & (!x15093x)) + ((!n_n3509) & (!n_n1677) & (n_n2629) & (x15091x) & (x15093x)) + ((!n_n3509) & (n_n1677) & (!n_n2629) & (!x15091x) & (!x15093x)) + ((!n_n3509) & (n_n1677) & (!n_n2629) & (!x15091x) & (x15093x)) + ((!n_n3509) & (n_n1677) & (!n_n2629) & (x15091x) & (!x15093x)) + ((!n_n3509) & (n_n1677) & (!n_n2629) & (x15091x) & (x15093x)) + ((!n_n3509) & (n_n1677) & (n_n2629) & (!x15091x) & (!x15093x)) + ((!n_n3509) & (n_n1677) & (n_n2629) & (!x15091x) & (x15093x)) + ((!n_n3509) & (n_n1677) & (n_n2629) & (x15091x) & (!x15093x)) + ((!n_n3509) & (n_n1677) & (n_n2629) & (x15091x) & (x15093x)) + ((n_n3509) & (!n_n1677) & (!n_n2629) & (!x15091x) & (!x15093x)) + ((n_n3509) & (!n_n1677) & (!n_n2629) & (!x15091x) & (x15093x)) + ((n_n3509) & (!n_n1677) & (!n_n2629) & (x15091x) & (!x15093x)) + ((n_n3509) & (!n_n1677) & (!n_n2629) & (x15091x) & (x15093x)) + ((n_n3509) & (!n_n1677) & (n_n2629) & (!x15091x) & (!x15093x)) + ((n_n3509) & (!n_n1677) & (n_n2629) & (!x15091x) & (x15093x)) + ((n_n3509) & (!n_n1677) & (n_n2629) & (x15091x) & (!x15093x)) + ((n_n3509) & (!n_n1677) & (n_n2629) & (x15091x) & (x15093x)) + ((n_n3509) & (n_n1677) & (!n_n2629) & (!x15091x) & (!x15093x)) + ((n_n3509) & (n_n1677) & (!n_n2629) & (!x15091x) & (x15093x)) + ((n_n3509) & (n_n1677) & (!n_n2629) & (x15091x) & (!x15093x)) + ((n_n3509) & (n_n1677) & (!n_n2629) & (x15091x) & (x15093x)) + ((n_n3509) & (n_n1677) & (n_n2629) & (!x15091x) & (!x15093x)) + ((n_n3509) & (n_n1677) & (n_n2629) & (!x15091x) & (x15093x)) + ((n_n3509) & (n_n1677) & (n_n2629) & (x15091x) & (!x15093x)) + ((n_n3509) & (n_n1677) & (n_n2629) & (x15091x) & (x15093x)));
	assign x178x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n482) & (n_n455)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n482) & (n_n455)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n482) & (n_n455)) + ((i_9_) & (n_n524) & (n_n526) & (n_n482) & (n_n455)));
	assign x15101x = (((!n_n4532) & (!n_n4528) & (!x178x) & (!x15096x) & (x15098x)) + ((!n_n4532) & (!n_n4528) & (!x178x) & (x15096x) & (!x15098x)) + ((!n_n4532) & (!n_n4528) & (!x178x) & (x15096x) & (x15098x)) + ((!n_n4532) & (!n_n4528) & (x178x) & (!x15096x) & (!x15098x)) + ((!n_n4532) & (!n_n4528) & (x178x) & (!x15096x) & (x15098x)) + ((!n_n4532) & (!n_n4528) & (x178x) & (x15096x) & (!x15098x)) + ((!n_n4532) & (!n_n4528) & (x178x) & (x15096x) & (x15098x)) + ((!n_n4532) & (n_n4528) & (!x178x) & (!x15096x) & (!x15098x)) + ((!n_n4532) & (n_n4528) & (!x178x) & (!x15096x) & (x15098x)) + ((!n_n4532) & (n_n4528) & (!x178x) & (x15096x) & (!x15098x)) + ((!n_n4532) & (n_n4528) & (!x178x) & (x15096x) & (x15098x)) + ((!n_n4532) & (n_n4528) & (x178x) & (!x15096x) & (!x15098x)) + ((!n_n4532) & (n_n4528) & (x178x) & (!x15096x) & (x15098x)) + ((!n_n4532) & (n_n4528) & (x178x) & (x15096x) & (!x15098x)) + ((!n_n4532) & (n_n4528) & (x178x) & (x15096x) & (x15098x)) + ((n_n4532) & (!n_n4528) & (!x178x) & (!x15096x) & (!x15098x)) + ((n_n4532) & (!n_n4528) & (!x178x) & (!x15096x) & (x15098x)) + ((n_n4532) & (!n_n4528) & (!x178x) & (x15096x) & (!x15098x)) + ((n_n4532) & (!n_n4528) & (!x178x) & (x15096x) & (x15098x)) + ((n_n4532) & (!n_n4528) & (x178x) & (!x15096x) & (!x15098x)) + ((n_n4532) & (!n_n4528) & (x178x) & (!x15096x) & (x15098x)) + ((n_n4532) & (!n_n4528) & (x178x) & (x15096x) & (!x15098x)) + ((n_n4532) & (!n_n4528) & (x178x) & (x15096x) & (x15098x)) + ((n_n4532) & (n_n4528) & (!x178x) & (!x15096x) & (!x15098x)) + ((n_n4532) & (n_n4528) & (!x178x) & (!x15096x) & (x15098x)) + ((n_n4532) & (n_n4528) & (!x178x) & (x15096x) & (!x15098x)) + ((n_n4532) & (n_n4528) & (!x178x) & (x15096x) & (x15098x)) + ((n_n4532) & (n_n4528) & (x178x) & (!x15096x) & (!x15098x)) + ((n_n4532) & (n_n4528) & (x178x) & (!x15096x) & (x15098x)) + ((n_n4532) & (n_n4528) & (x178x) & (x15096x) & (!x15098x)) + ((n_n4532) & (n_n4528) & (x178x) & (x15096x) & (x15098x)));
	assign x15103x = (((!x15061x) & (!x15062x) & (!x15080x) & (!x15081x) & (x15101x)) + ((!x15061x) & (!x15062x) & (!x15080x) & (x15081x) & (!x15101x)) + ((!x15061x) & (!x15062x) & (!x15080x) & (x15081x) & (x15101x)) + ((!x15061x) & (!x15062x) & (x15080x) & (!x15081x) & (!x15101x)) + ((!x15061x) & (!x15062x) & (x15080x) & (!x15081x) & (x15101x)) + ((!x15061x) & (!x15062x) & (x15080x) & (x15081x) & (!x15101x)) + ((!x15061x) & (!x15062x) & (x15080x) & (x15081x) & (x15101x)) + ((!x15061x) & (x15062x) & (!x15080x) & (!x15081x) & (!x15101x)) + ((!x15061x) & (x15062x) & (!x15080x) & (!x15081x) & (x15101x)) + ((!x15061x) & (x15062x) & (!x15080x) & (x15081x) & (!x15101x)) + ((!x15061x) & (x15062x) & (!x15080x) & (x15081x) & (x15101x)) + ((!x15061x) & (x15062x) & (x15080x) & (!x15081x) & (!x15101x)) + ((!x15061x) & (x15062x) & (x15080x) & (!x15081x) & (x15101x)) + ((!x15061x) & (x15062x) & (x15080x) & (x15081x) & (!x15101x)) + ((!x15061x) & (x15062x) & (x15080x) & (x15081x) & (x15101x)) + ((x15061x) & (!x15062x) & (!x15080x) & (!x15081x) & (!x15101x)) + ((x15061x) & (!x15062x) & (!x15080x) & (!x15081x) & (x15101x)) + ((x15061x) & (!x15062x) & (!x15080x) & (x15081x) & (!x15101x)) + ((x15061x) & (!x15062x) & (!x15080x) & (x15081x) & (x15101x)) + ((x15061x) & (!x15062x) & (x15080x) & (!x15081x) & (!x15101x)) + ((x15061x) & (!x15062x) & (x15080x) & (!x15081x) & (x15101x)) + ((x15061x) & (!x15062x) & (x15080x) & (x15081x) & (!x15101x)) + ((x15061x) & (!x15062x) & (x15080x) & (x15081x) & (x15101x)) + ((x15061x) & (x15062x) & (!x15080x) & (!x15081x) & (!x15101x)) + ((x15061x) & (x15062x) & (!x15080x) & (!x15081x) & (x15101x)) + ((x15061x) & (x15062x) & (!x15080x) & (x15081x) & (!x15101x)) + ((x15061x) & (x15062x) & (!x15080x) & (x15081x) & (x15101x)) + ((x15061x) & (x15062x) & (x15080x) & (!x15081x) & (!x15101x)) + ((x15061x) & (x15062x) & (x15080x) & (!x15081x) & (x15101x)) + ((x15061x) & (x15062x) & (x15080x) & (x15081x) & (!x15101x)) + ((x15061x) & (x15062x) & (x15080x) & (x15081x) & (x15101x)));
	assign n_n2619 = (((!x108x) & (!x45x) & (!n_n4603) & (!x22097x)) + ((!x108x) & (!x45x) & (n_n4603) & (!x22097x)) + ((!x108x) & (!x45x) & (n_n4603) & (x22097x)) + ((!x108x) & (x45x) & (!n_n4603) & (!x22097x)) + ((!x108x) & (x45x) & (!n_n4603) & (x22097x)) + ((!x108x) & (x45x) & (n_n4603) & (!x22097x)) + ((!x108x) & (x45x) & (n_n4603) & (x22097x)) + ((x108x) & (!x45x) & (!n_n4603) & (!x22097x)) + ((x108x) & (!x45x) & (!n_n4603) & (x22097x)) + ((x108x) & (!x45x) & (n_n4603) & (!x22097x)) + ((x108x) & (!x45x) & (n_n4603) & (x22097x)) + ((x108x) & (x45x) & (!n_n4603) & (!x22097x)) + ((x108x) & (x45x) & (!n_n4603) & (x22097x)) + ((x108x) & (x45x) & (n_n4603) & (!x22097x)) + ((x108x) & (x45x) & (n_n4603) & (x22097x)));
	assign n_n2618 = (((!n_n4617) & (!n_n4610) & (!x51x) & (!x22167x)) + ((!n_n4617) & (!n_n4610) & (x51x) & (!x22167x)) + ((!n_n4617) & (!n_n4610) & (x51x) & (x22167x)) + ((!n_n4617) & (n_n4610) & (!x51x) & (!x22167x)) + ((!n_n4617) & (n_n4610) & (!x51x) & (x22167x)) + ((!n_n4617) & (n_n4610) & (x51x) & (!x22167x)) + ((!n_n4617) & (n_n4610) & (x51x) & (x22167x)) + ((n_n4617) & (!n_n4610) & (!x51x) & (!x22167x)) + ((n_n4617) & (!n_n4610) & (!x51x) & (x22167x)) + ((n_n4617) & (!n_n4610) & (x51x) & (!x22167x)) + ((n_n4617) & (!n_n4610) & (x51x) & (x22167x)) + ((n_n4617) & (n_n4610) & (!x51x) & (!x22167x)) + ((n_n4617) & (n_n4610) & (!x51x) & (x22167x)) + ((n_n4617) & (n_n4610) & (x51x) & (!x22167x)) + ((n_n4617) & (n_n4610) & (x51x) & (x22167x)));
	assign x15119x = (((!n_n4594) & (!n_n4586) & (!n_n4588) & (n_n4583)) + ((!n_n4594) & (!n_n4586) & (n_n4588) & (!n_n4583)) + ((!n_n4594) & (!n_n4586) & (n_n4588) & (n_n4583)) + ((!n_n4594) & (n_n4586) & (!n_n4588) & (!n_n4583)) + ((!n_n4594) & (n_n4586) & (!n_n4588) & (n_n4583)) + ((!n_n4594) & (n_n4586) & (n_n4588) & (!n_n4583)) + ((!n_n4594) & (n_n4586) & (n_n4588) & (n_n4583)) + ((n_n4594) & (!n_n4586) & (!n_n4588) & (!n_n4583)) + ((n_n4594) & (!n_n4586) & (!n_n4588) & (n_n4583)) + ((n_n4594) & (!n_n4586) & (n_n4588) & (!n_n4583)) + ((n_n4594) & (!n_n4586) & (n_n4588) & (n_n4583)) + ((n_n4594) & (n_n4586) & (!n_n4588) & (!n_n4583)) + ((n_n4594) & (n_n4586) & (!n_n4588) & (n_n4583)) + ((n_n4594) & (n_n4586) & (n_n4588) & (!n_n4583)) + ((n_n4594) & (n_n4586) & (n_n4588) & (n_n4583)));
	assign x15120x = (((!n_n4597) & (!n_n4595) & (!n_n4590) & (!n_n4591) & (n_n4585)) + ((!n_n4597) & (!n_n4595) & (!n_n4590) & (n_n4591) & (!n_n4585)) + ((!n_n4597) & (!n_n4595) & (!n_n4590) & (n_n4591) & (n_n4585)) + ((!n_n4597) & (!n_n4595) & (n_n4590) & (!n_n4591) & (!n_n4585)) + ((!n_n4597) & (!n_n4595) & (n_n4590) & (!n_n4591) & (n_n4585)) + ((!n_n4597) & (!n_n4595) & (n_n4590) & (n_n4591) & (!n_n4585)) + ((!n_n4597) & (!n_n4595) & (n_n4590) & (n_n4591) & (n_n4585)) + ((!n_n4597) & (n_n4595) & (!n_n4590) & (!n_n4591) & (!n_n4585)) + ((!n_n4597) & (n_n4595) & (!n_n4590) & (!n_n4591) & (n_n4585)) + ((!n_n4597) & (n_n4595) & (!n_n4590) & (n_n4591) & (!n_n4585)) + ((!n_n4597) & (n_n4595) & (!n_n4590) & (n_n4591) & (n_n4585)) + ((!n_n4597) & (n_n4595) & (n_n4590) & (!n_n4591) & (!n_n4585)) + ((!n_n4597) & (n_n4595) & (n_n4590) & (!n_n4591) & (n_n4585)) + ((!n_n4597) & (n_n4595) & (n_n4590) & (n_n4591) & (!n_n4585)) + ((!n_n4597) & (n_n4595) & (n_n4590) & (n_n4591) & (n_n4585)) + ((n_n4597) & (!n_n4595) & (!n_n4590) & (!n_n4591) & (!n_n4585)) + ((n_n4597) & (!n_n4595) & (!n_n4590) & (!n_n4591) & (n_n4585)) + ((n_n4597) & (!n_n4595) & (!n_n4590) & (n_n4591) & (!n_n4585)) + ((n_n4597) & (!n_n4595) & (!n_n4590) & (n_n4591) & (n_n4585)) + ((n_n4597) & (!n_n4595) & (n_n4590) & (!n_n4591) & (!n_n4585)) + ((n_n4597) & (!n_n4595) & (n_n4590) & (!n_n4591) & (n_n4585)) + ((n_n4597) & (!n_n4595) & (n_n4590) & (n_n4591) & (!n_n4585)) + ((n_n4597) & (!n_n4595) & (n_n4590) & (n_n4591) & (n_n4585)) + ((n_n4597) & (n_n4595) & (!n_n4590) & (!n_n4591) & (!n_n4585)) + ((n_n4597) & (n_n4595) & (!n_n4590) & (!n_n4591) & (n_n4585)) + ((n_n4597) & (n_n4595) & (!n_n4590) & (n_n4591) & (!n_n4585)) + ((n_n4597) & (n_n4595) & (!n_n4590) & (n_n4591) & (n_n4585)) + ((n_n4597) & (n_n4595) & (n_n4590) & (!n_n4591) & (!n_n4585)) + ((n_n4597) & (n_n4595) & (n_n4590) & (!n_n4591) & (n_n4585)) + ((n_n4597) & (n_n4595) & (n_n4590) & (n_n4591) & (!n_n4585)) + ((n_n4597) & (n_n4595) & (n_n4590) & (n_n4591) & (n_n4585)));
	assign n_n2554 = (((!n_n2619) & (!n_n2618) & (!x15119x) & (x15120x)) + ((!n_n2619) & (!n_n2618) & (x15119x) & (!x15120x)) + ((!n_n2619) & (!n_n2618) & (x15119x) & (x15120x)) + ((!n_n2619) & (n_n2618) & (!x15119x) & (!x15120x)) + ((!n_n2619) & (n_n2618) & (!x15119x) & (x15120x)) + ((!n_n2619) & (n_n2618) & (x15119x) & (!x15120x)) + ((!n_n2619) & (n_n2618) & (x15119x) & (x15120x)) + ((n_n2619) & (!n_n2618) & (!x15119x) & (!x15120x)) + ((n_n2619) & (!n_n2618) & (!x15119x) & (x15120x)) + ((n_n2619) & (!n_n2618) & (x15119x) & (!x15120x)) + ((n_n2619) & (!n_n2618) & (x15119x) & (x15120x)) + ((n_n2619) & (n_n2618) & (!x15119x) & (!x15120x)) + ((n_n2619) & (n_n2618) & (!x15119x) & (x15120x)) + ((n_n2619) & (n_n2618) & (x15119x) & (!x15120x)) + ((n_n2619) & (n_n2618) & (x15119x) & (x15120x)));
	assign x238x = (((!i_9_) & (!n_n528) & (n_n390) & (n_n535) & (n_n530)) + ((!i_9_) & (n_n528) & (n_n390) & (n_n535) & (!n_n530)) + ((!i_9_) & (n_n528) & (n_n390) & (n_n535) & (n_n530)));
	assign x15126x = (((!n_n4578) & (!n_n4574) & (!n_n4580) & (x238x)) + ((!n_n4578) & (!n_n4574) & (n_n4580) & (!x238x)) + ((!n_n4578) & (!n_n4574) & (n_n4580) & (x238x)) + ((!n_n4578) & (n_n4574) & (!n_n4580) & (!x238x)) + ((!n_n4578) & (n_n4574) & (!n_n4580) & (x238x)) + ((!n_n4578) & (n_n4574) & (n_n4580) & (!x238x)) + ((!n_n4578) & (n_n4574) & (n_n4580) & (x238x)) + ((n_n4578) & (!n_n4574) & (!n_n4580) & (!x238x)) + ((n_n4578) & (!n_n4574) & (!n_n4580) & (x238x)) + ((n_n4578) & (!n_n4574) & (n_n4580) & (!x238x)) + ((n_n4578) & (!n_n4574) & (n_n4580) & (x238x)) + ((n_n4578) & (n_n4574) & (!n_n4580) & (!x238x)) + ((n_n4578) & (n_n4574) & (!n_n4580) & (x238x)) + ((n_n4578) & (n_n4574) & (n_n4580) & (!x238x)) + ((n_n4578) & (n_n4574) & (n_n4580) & (x238x)));
	assign n_n2621 = (((!n_n4582) & (!n_n4577) & (!n_n4576) & (!n_n4581) & (x15126x)) + ((!n_n4582) & (!n_n4577) & (!n_n4576) & (n_n4581) & (!x15126x)) + ((!n_n4582) & (!n_n4577) & (!n_n4576) & (n_n4581) & (x15126x)) + ((!n_n4582) & (!n_n4577) & (n_n4576) & (!n_n4581) & (!x15126x)) + ((!n_n4582) & (!n_n4577) & (n_n4576) & (!n_n4581) & (x15126x)) + ((!n_n4582) & (!n_n4577) & (n_n4576) & (n_n4581) & (!x15126x)) + ((!n_n4582) & (!n_n4577) & (n_n4576) & (n_n4581) & (x15126x)) + ((!n_n4582) & (n_n4577) & (!n_n4576) & (!n_n4581) & (!x15126x)) + ((!n_n4582) & (n_n4577) & (!n_n4576) & (!n_n4581) & (x15126x)) + ((!n_n4582) & (n_n4577) & (!n_n4576) & (n_n4581) & (!x15126x)) + ((!n_n4582) & (n_n4577) & (!n_n4576) & (n_n4581) & (x15126x)) + ((!n_n4582) & (n_n4577) & (n_n4576) & (!n_n4581) & (!x15126x)) + ((!n_n4582) & (n_n4577) & (n_n4576) & (!n_n4581) & (x15126x)) + ((!n_n4582) & (n_n4577) & (n_n4576) & (n_n4581) & (!x15126x)) + ((!n_n4582) & (n_n4577) & (n_n4576) & (n_n4581) & (x15126x)) + ((n_n4582) & (!n_n4577) & (!n_n4576) & (!n_n4581) & (!x15126x)) + ((n_n4582) & (!n_n4577) & (!n_n4576) & (!n_n4581) & (x15126x)) + ((n_n4582) & (!n_n4577) & (!n_n4576) & (n_n4581) & (!x15126x)) + ((n_n4582) & (!n_n4577) & (!n_n4576) & (n_n4581) & (x15126x)) + ((n_n4582) & (!n_n4577) & (n_n4576) & (!n_n4581) & (!x15126x)) + ((n_n4582) & (!n_n4577) & (n_n4576) & (!n_n4581) & (x15126x)) + ((n_n4582) & (!n_n4577) & (n_n4576) & (n_n4581) & (!x15126x)) + ((n_n4582) & (!n_n4577) & (n_n4576) & (n_n4581) & (x15126x)) + ((n_n4582) & (n_n4577) & (!n_n4576) & (!n_n4581) & (!x15126x)) + ((n_n4582) & (n_n4577) & (!n_n4576) & (!n_n4581) & (x15126x)) + ((n_n4582) & (n_n4577) & (!n_n4576) & (n_n4581) & (!x15126x)) + ((n_n4582) & (n_n4577) & (!n_n4576) & (n_n4581) & (x15126x)) + ((n_n4582) & (n_n4577) & (n_n4576) & (!n_n4581) & (!x15126x)) + ((n_n4582) & (n_n4577) & (n_n4576) & (!n_n4581) & (x15126x)) + ((n_n4582) & (n_n4577) & (n_n4576) & (n_n4581) & (!x15126x)) + ((n_n4582) & (n_n4577) & (n_n4576) & (n_n4581) & (x15126x)));
	assign n_n2615 = (((!n_n4659) & (!n_n4661) & (!n_n4657) & (!x431x) & (!x22096x)) + ((!n_n4659) & (!n_n4661) & (!n_n4657) & (x431x) & (!x22096x)) + ((!n_n4659) & (!n_n4661) & (!n_n4657) & (x431x) & (x22096x)) + ((!n_n4659) & (!n_n4661) & (n_n4657) & (!x431x) & (!x22096x)) + ((!n_n4659) & (!n_n4661) & (n_n4657) & (!x431x) & (x22096x)) + ((!n_n4659) & (!n_n4661) & (n_n4657) & (x431x) & (!x22096x)) + ((!n_n4659) & (!n_n4661) & (n_n4657) & (x431x) & (x22096x)) + ((!n_n4659) & (n_n4661) & (!n_n4657) & (!x431x) & (!x22096x)) + ((!n_n4659) & (n_n4661) & (!n_n4657) & (!x431x) & (x22096x)) + ((!n_n4659) & (n_n4661) & (!n_n4657) & (x431x) & (!x22096x)) + ((!n_n4659) & (n_n4661) & (!n_n4657) & (x431x) & (x22096x)) + ((!n_n4659) & (n_n4661) & (n_n4657) & (!x431x) & (!x22096x)) + ((!n_n4659) & (n_n4661) & (n_n4657) & (!x431x) & (x22096x)) + ((!n_n4659) & (n_n4661) & (n_n4657) & (x431x) & (!x22096x)) + ((!n_n4659) & (n_n4661) & (n_n4657) & (x431x) & (x22096x)) + ((n_n4659) & (!n_n4661) & (!n_n4657) & (!x431x) & (!x22096x)) + ((n_n4659) & (!n_n4661) & (!n_n4657) & (!x431x) & (x22096x)) + ((n_n4659) & (!n_n4661) & (!n_n4657) & (x431x) & (!x22096x)) + ((n_n4659) & (!n_n4661) & (!n_n4657) & (x431x) & (x22096x)) + ((n_n4659) & (!n_n4661) & (n_n4657) & (!x431x) & (!x22096x)) + ((n_n4659) & (!n_n4661) & (n_n4657) & (!x431x) & (x22096x)) + ((n_n4659) & (!n_n4661) & (n_n4657) & (x431x) & (!x22096x)) + ((n_n4659) & (!n_n4661) & (n_n4657) & (x431x) & (x22096x)) + ((n_n4659) & (n_n4661) & (!n_n4657) & (!x431x) & (!x22096x)) + ((n_n4659) & (n_n4661) & (!n_n4657) & (!x431x) & (x22096x)) + ((n_n4659) & (n_n4661) & (!n_n4657) & (x431x) & (!x22096x)) + ((n_n4659) & (n_n4661) & (!n_n4657) & (x431x) & (x22096x)) + ((n_n4659) & (n_n4661) & (n_n4657) & (!x431x) & (!x22096x)) + ((n_n4659) & (n_n4661) & (n_n4657) & (!x431x) & (x22096x)) + ((n_n4659) & (n_n4661) & (n_n4657) & (x431x) & (!x22096x)) + ((n_n4659) & (n_n4661) & (n_n4657) & (x431x) & (x22096x)));
	assign n_n2030 = (((!i_9_) & (!n_n526) & (n_n528) & (n_n390) & (n_n491)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n390) & (n_n491)) + ((i_9_) & (!n_n526) & (n_n528) & (n_n390) & (n_n491)) + ((i_9_) & (n_n526) & (!n_n528) & (n_n390) & (n_n491)) + ((i_9_) & (n_n526) & (n_n528) & (n_n390) & (n_n491)));
	assign x15137x = (((!n_n4634) & (!n_n4642) & (!n_n4635) & (n_n4623)) + ((!n_n4634) & (!n_n4642) & (n_n4635) & (!n_n4623)) + ((!n_n4634) & (!n_n4642) & (n_n4635) & (n_n4623)) + ((!n_n4634) & (n_n4642) & (!n_n4635) & (!n_n4623)) + ((!n_n4634) & (n_n4642) & (!n_n4635) & (n_n4623)) + ((!n_n4634) & (n_n4642) & (n_n4635) & (!n_n4623)) + ((!n_n4634) & (n_n4642) & (n_n4635) & (n_n4623)) + ((n_n4634) & (!n_n4642) & (!n_n4635) & (!n_n4623)) + ((n_n4634) & (!n_n4642) & (!n_n4635) & (n_n4623)) + ((n_n4634) & (!n_n4642) & (n_n4635) & (!n_n4623)) + ((n_n4634) & (!n_n4642) & (n_n4635) & (n_n4623)) + ((n_n4634) & (n_n4642) & (!n_n4635) & (!n_n4623)) + ((n_n4634) & (n_n4642) & (!n_n4635) & (n_n4623)) + ((n_n4634) & (n_n4642) & (n_n4635) & (!n_n4623)) + ((n_n4634) & (n_n4642) & (n_n4635) & (n_n4623)));
	assign x15139x = (((!n_n4641) & (!x26x) & (!n_n4643) & (!x357x) & (x190x)) + ((!n_n4641) & (!x26x) & (!n_n4643) & (x357x) & (!x190x)) + ((!n_n4641) & (!x26x) & (!n_n4643) & (x357x) & (x190x)) + ((!n_n4641) & (!x26x) & (n_n4643) & (!x357x) & (!x190x)) + ((!n_n4641) & (!x26x) & (n_n4643) & (!x357x) & (x190x)) + ((!n_n4641) & (!x26x) & (n_n4643) & (x357x) & (!x190x)) + ((!n_n4641) & (!x26x) & (n_n4643) & (x357x) & (x190x)) + ((!n_n4641) & (x26x) & (!n_n4643) & (!x357x) & (!x190x)) + ((!n_n4641) & (x26x) & (!n_n4643) & (!x357x) & (x190x)) + ((!n_n4641) & (x26x) & (!n_n4643) & (x357x) & (!x190x)) + ((!n_n4641) & (x26x) & (!n_n4643) & (x357x) & (x190x)) + ((!n_n4641) & (x26x) & (n_n4643) & (!x357x) & (!x190x)) + ((!n_n4641) & (x26x) & (n_n4643) & (!x357x) & (x190x)) + ((!n_n4641) & (x26x) & (n_n4643) & (x357x) & (!x190x)) + ((!n_n4641) & (x26x) & (n_n4643) & (x357x) & (x190x)) + ((n_n4641) & (!x26x) & (!n_n4643) & (!x357x) & (!x190x)) + ((n_n4641) & (!x26x) & (!n_n4643) & (!x357x) & (x190x)) + ((n_n4641) & (!x26x) & (!n_n4643) & (x357x) & (!x190x)) + ((n_n4641) & (!x26x) & (!n_n4643) & (x357x) & (x190x)) + ((n_n4641) & (!x26x) & (n_n4643) & (!x357x) & (!x190x)) + ((n_n4641) & (!x26x) & (n_n4643) & (!x357x) & (x190x)) + ((n_n4641) & (!x26x) & (n_n4643) & (x357x) & (!x190x)) + ((n_n4641) & (!x26x) & (n_n4643) & (x357x) & (x190x)) + ((n_n4641) & (x26x) & (!n_n4643) & (!x357x) & (!x190x)) + ((n_n4641) & (x26x) & (!n_n4643) & (!x357x) & (x190x)) + ((n_n4641) & (x26x) & (!n_n4643) & (x357x) & (!x190x)) + ((n_n4641) & (x26x) & (!n_n4643) & (x357x) & (x190x)) + ((n_n4641) & (x26x) & (n_n4643) & (!x357x) & (!x190x)) + ((n_n4641) & (x26x) & (n_n4643) & (!x357x) & (x190x)) + ((n_n4641) & (x26x) & (n_n4643) & (x357x) & (!x190x)) + ((n_n4641) & (x26x) & (n_n4643) & (x357x) & (x190x)));
	assign n_n2553 = (((!n_n2615) & (!n_n2761) & (!n_n2030) & (!x15137x) & (x15139x)) + ((!n_n2615) & (!n_n2761) & (!n_n2030) & (x15137x) & (!x15139x)) + ((!n_n2615) & (!n_n2761) & (!n_n2030) & (x15137x) & (x15139x)) + ((!n_n2615) & (!n_n2761) & (n_n2030) & (!x15137x) & (!x15139x)) + ((!n_n2615) & (!n_n2761) & (n_n2030) & (!x15137x) & (x15139x)) + ((!n_n2615) & (!n_n2761) & (n_n2030) & (x15137x) & (!x15139x)) + ((!n_n2615) & (!n_n2761) & (n_n2030) & (x15137x) & (x15139x)) + ((!n_n2615) & (n_n2761) & (!n_n2030) & (!x15137x) & (!x15139x)) + ((!n_n2615) & (n_n2761) & (!n_n2030) & (!x15137x) & (x15139x)) + ((!n_n2615) & (n_n2761) & (!n_n2030) & (x15137x) & (!x15139x)) + ((!n_n2615) & (n_n2761) & (!n_n2030) & (x15137x) & (x15139x)) + ((!n_n2615) & (n_n2761) & (n_n2030) & (!x15137x) & (!x15139x)) + ((!n_n2615) & (n_n2761) & (n_n2030) & (!x15137x) & (x15139x)) + ((!n_n2615) & (n_n2761) & (n_n2030) & (x15137x) & (!x15139x)) + ((!n_n2615) & (n_n2761) & (n_n2030) & (x15137x) & (x15139x)) + ((n_n2615) & (!n_n2761) & (!n_n2030) & (!x15137x) & (!x15139x)) + ((n_n2615) & (!n_n2761) & (!n_n2030) & (!x15137x) & (x15139x)) + ((n_n2615) & (!n_n2761) & (!n_n2030) & (x15137x) & (!x15139x)) + ((n_n2615) & (!n_n2761) & (!n_n2030) & (x15137x) & (x15139x)) + ((n_n2615) & (!n_n2761) & (n_n2030) & (!x15137x) & (!x15139x)) + ((n_n2615) & (!n_n2761) & (n_n2030) & (!x15137x) & (x15139x)) + ((n_n2615) & (!n_n2761) & (n_n2030) & (x15137x) & (!x15139x)) + ((n_n2615) & (!n_n2761) & (n_n2030) & (x15137x) & (x15139x)) + ((n_n2615) & (n_n2761) & (!n_n2030) & (!x15137x) & (!x15139x)) + ((n_n2615) & (n_n2761) & (!n_n2030) & (!x15137x) & (x15139x)) + ((n_n2615) & (n_n2761) & (!n_n2030) & (x15137x) & (!x15139x)) + ((n_n2615) & (n_n2761) & (!n_n2030) & (x15137x) & (x15139x)) + ((n_n2615) & (n_n2761) & (n_n2030) & (!x15137x) & (!x15139x)) + ((n_n2615) & (n_n2761) & (n_n2030) & (!x15137x) & (x15139x)) + ((n_n2615) & (n_n2761) & (n_n2030) & (x15137x) & (!x15139x)) + ((n_n2615) & (n_n2761) & (n_n2030) & (x15137x) & (x15139x)));
	assign x82x = (((!i_9_) & (n_n455) & (!n_n532) & (n_n534) & (n_n464)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n534) & (n_n464)) + ((i_9_) & (n_n455) & (!n_n532) & (n_n534) & (n_n464)) + ((i_9_) & (n_n455) & (n_n532) & (!n_n534) & (n_n464)) + ((i_9_) & (n_n455) & (n_n532) & (n_n534) & (n_n464)));
	assign x224x = (((!n_n4562) & (!x471x) & (!x91x) & (x222x)) + ((!n_n4562) & (!x471x) & (x91x) & (!x222x)) + ((!n_n4562) & (!x471x) & (x91x) & (x222x)) + ((!n_n4562) & (x471x) & (!x91x) & (!x222x)) + ((!n_n4562) & (x471x) & (!x91x) & (x222x)) + ((!n_n4562) & (x471x) & (x91x) & (!x222x)) + ((!n_n4562) & (x471x) & (x91x) & (x222x)) + ((n_n4562) & (!x471x) & (!x91x) & (!x222x)) + ((n_n4562) & (!x471x) & (!x91x) & (x222x)) + ((n_n4562) & (!x471x) & (x91x) & (!x222x)) + ((n_n4562) & (!x471x) & (x91x) & (x222x)) + ((n_n4562) & (x471x) & (!x91x) & (!x222x)) + ((n_n4562) & (x471x) & (!x91x) & (x222x)) + ((n_n4562) & (x471x) & (x91x) & (!x222x)) + ((n_n4562) & (x471x) & (x91x) & (x222x)));
	assign x15146x = (((!x10x) & (!n_n535) & (!n_n530) & (!n_n4555) & (x82x)) + ((!x10x) & (!n_n535) & (!n_n530) & (n_n4555) & (!x82x)) + ((!x10x) & (!n_n535) & (!n_n530) & (n_n4555) & (x82x)) + ((!x10x) & (!n_n535) & (n_n530) & (!n_n4555) & (x82x)) + ((!x10x) & (!n_n535) & (n_n530) & (n_n4555) & (!x82x)) + ((!x10x) & (!n_n535) & (n_n530) & (n_n4555) & (x82x)) + ((!x10x) & (n_n535) & (!n_n530) & (!n_n4555) & (x82x)) + ((!x10x) & (n_n535) & (!n_n530) & (n_n4555) & (!x82x)) + ((!x10x) & (n_n535) & (!n_n530) & (n_n4555) & (x82x)) + ((!x10x) & (n_n535) & (n_n530) & (!n_n4555) & (x82x)) + ((!x10x) & (n_n535) & (n_n530) & (n_n4555) & (!x82x)) + ((!x10x) & (n_n535) & (n_n530) & (n_n4555) & (x82x)) + ((x10x) & (!n_n535) & (!n_n530) & (!n_n4555) & (x82x)) + ((x10x) & (!n_n535) & (!n_n530) & (n_n4555) & (!x82x)) + ((x10x) & (!n_n535) & (!n_n530) & (n_n4555) & (x82x)) + ((x10x) & (!n_n535) & (n_n530) & (!n_n4555) & (x82x)) + ((x10x) & (!n_n535) & (n_n530) & (n_n4555) & (!x82x)) + ((x10x) & (!n_n535) & (n_n530) & (n_n4555) & (x82x)) + ((x10x) & (n_n535) & (!n_n530) & (!n_n4555) & (x82x)) + ((x10x) & (n_n535) & (!n_n530) & (n_n4555) & (!x82x)) + ((x10x) & (n_n535) & (!n_n530) & (n_n4555) & (x82x)) + ((x10x) & (n_n535) & (n_n530) & (!n_n4555) & (!x82x)) + ((x10x) & (n_n535) & (n_n530) & (!n_n4555) & (x82x)) + ((x10x) & (n_n535) & (n_n530) & (n_n4555) & (!x82x)) + ((x10x) & (n_n535) & (n_n530) & (n_n4555) & (x82x)));
	assign x15147x = (((!n_n4560) & (!n_n4561) & (!x212x) & (!n_n4551) & (x121x)) + ((!n_n4560) & (!n_n4561) & (!x212x) & (n_n4551) & (!x121x)) + ((!n_n4560) & (!n_n4561) & (!x212x) & (n_n4551) & (x121x)) + ((!n_n4560) & (!n_n4561) & (x212x) & (!n_n4551) & (!x121x)) + ((!n_n4560) & (!n_n4561) & (x212x) & (!n_n4551) & (x121x)) + ((!n_n4560) & (!n_n4561) & (x212x) & (n_n4551) & (!x121x)) + ((!n_n4560) & (!n_n4561) & (x212x) & (n_n4551) & (x121x)) + ((!n_n4560) & (n_n4561) & (!x212x) & (!n_n4551) & (!x121x)) + ((!n_n4560) & (n_n4561) & (!x212x) & (!n_n4551) & (x121x)) + ((!n_n4560) & (n_n4561) & (!x212x) & (n_n4551) & (!x121x)) + ((!n_n4560) & (n_n4561) & (!x212x) & (n_n4551) & (x121x)) + ((!n_n4560) & (n_n4561) & (x212x) & (!n_n4551) & (!x121x)) + ((!n_n4560) & (n_n4561) & (x212x) & (!n_n4551) & (x121x)) + ((!n_n4560) & (n_n4561) & (x212x) & (n_n4551) & (!x121x)) + ((!n_n4560) & (n_n4561) & (x212x) & (n_n4551) & (x121x)) + ((n_n4560) & (!n_n4561) & (!x212x) & (!n_n4551) & (!x121x)) + ((n_n4560) & (!n_n4561) & (!x212x) & (!n_n4551) & (x121x)) + ((n_n4560) & (!n_n4561) & (!x212x) & (n_n4551) & (!x121x)) + ((n_n4560) & (!n_n4561) & (!x212x) & (n_n4551) & (x121x)) + ((n_n4560) & (!n_n4561) & (x212x) & (!n_n4551) & (!x121x)) + ((n_n4560) & (!n_n4561) & (x212x) & (!n_n4551) & (x121x)) + ((n_n4560) & (!n_n4561) & (x212x) & (n_n4551) & (!x121x)) + ((n_n4560) & (!n_n4561) & (x212x) & (n_n4551) & (x121x)) + ((n_n4560) & (n_n4561) & (!x212x) & (!n_n4551) & (!x121x)) + ((n_n4560) & (n_n4561) & (!x212x) & (!n_n4551) & (x121x)) + ((n_n4560) & (n_n4561) & (!x212x) & (n_n4551) & (!x121x)) + ((n_n4560) & (n_n4561) & (!x212x) & (n_n4551) & (x121x)) + ((n_n4560) & (n_n4561) & (x212x) & (!n_n4551) & (!x121x)) + ((n_n4560) & (n_n4561) & (x212x) & (!n_n4551) & (x121x)) + ((n_n4560) & (n_n4561) & (x212x) & (n_n4551) & (!x121x)) + ((n_n4560) & (n_n4561) & (x212x) & (n_n4551) & (x121x)));
	assign x15150x = (((!n_n2621) & (!x224x) & (!x15146x) & (x15147x)) + ((!n_n2621) & (!x224x) & (x15146x) & (!x15147x)) + ((!n_n2621) & (!x224x) & (x15146x) & (x15147x)) + ((!n_n2621) & (x224x) & (!x15146x) & (!x15147x)) + ((!n_n2621) & (x224x) & (!x15146x) & (x15147x)) + ((!n_n2621) & (x224x) & (x15146x) & (!x15147x)) + ((!n_n2621) & (x224x) & (x15146x) & (x15147x)) + ((n_n2621) & (!x224x) & (!x15146x) & (!x15147x)) + ((n_n2621) & (!x224x) & (!x15146x) & (x15147x)) + ((n_n2621) & (!x224x) & (x15146x) & (!x15147x)) + ((n_n2621) & (!x224x) & (x15146x) & (x15147x)) + ((n_n2621) & (x224x) & (!x15146x) & (!x15147x)) + ((n_n2621) & (x224x) & (!x15146x) & (x15147x)) + ((n_n2621) & (x224x) & (x15146x) & (!x15147x)) + ((n_n2621) & (x224x) & (x15146x) & (x15147x)));
	assign x469x = (((!i_9_) & (n_n536) & (!n_n524) & (n_n518) & (n_n526)) + ((!i_9_) & (n_n536) & (n_n524) & (n_n518) & (!n_n526)) + ((!i_9_) & (n_n536) & (n_n524) & (n_n518) & (n_n526)) + ((i_9_) & (n_n536) & (n_n524) & (n_n518) & (!n_n526)) + ((i_9_) & (n_n536) & (n_n524) & (n_n518) & (n_n526)));
	assign x15152x = (((!i_9_) & (n_n536) & (n_n518) & (!n_n526) & (n_n534)) + ((!i_9_) & (n_n536) & (n_n518) & (n_n526) & (n_n534)) + ((i_9_) & (n_n536) & (n_n518) & (n_n526) & (!n_n534)) + ((i_9_) & (n_n536) & (n_n518) & (n_n526) & (n_n534)));
	assign n_n2640 = (((!x198x) & (!n_n4335) & (!n_n4334) & (!x469x) & (x15152x)) + ((!x198x) & (!n_n4335) & (!n_n4334) & (x469x) & (!x15152x)) + ((!x198x) & (!n_n4335) & (!n_n4334) & (x469x) & (x15152x)) + ((!x198x) & (!n_n4335) & (n_n4334) & (!x469x) & (!x15152x)) + ((!x198x) & (!n_n4335) & (n_n4334) & (!x469x) & (x15152x)) + ((!x198x) & (!n_n4335) & (n_n4334) & (x469x) & (!x15152x)) + ((!x198x) & (!n_n4335) & (n_n4334) & (x469x) & (x15152x)) + ((!x198x) & (n_n4335) & (!n_n4334) & (!x469x) & (!x15152x)) + ((!x198x) & (n_n4335) & (!n_n4334) & (!x469x) & (x15152x)) + ((!x198x) & (n_n4335) & (!n_n4334) & (x469x) & (!x15152x)) + ((!x198x) & (n_n4335) & (!n_n4334) & (x469x) & (x15152x)) + ((!x198x) & (n_n4335) & (n_n4334) & (!x469x) & (!x15152x)) + ((!x198x) & (n_n4335) & (n_n4334) & (!x469x) & (x15152x)) + ((!x198x) & (n_n4335) & (n_n4334) & (x469x) & (!x15152x)) + ((!x198x) & (n_n4335) & (n_n4334) & (x469x) & (x15152x)) + ((x198x) & (!n_n4335) & (!n_n4334) & (!x469x) & (!x15152x)) + ((x198x) & (!n_n4335) & (!n_n4334) & (!x469x) & (x15152x)) + ((x198x) & (!n_n4335) & (!n_n4334) & (x469x) & (!x15152x)) + ((x198x) & (!n_n4335) & (!n_n4334) & (x469x) & (x15152x)) + ((x198x) & (!n_n4335) & (n_n4334) & (!x469x) & (!x15152x)) + ((x198x) & (!n_n4335) & (n_n4334) & (!x469x) & (x15152x)) + ((x198x) & (!n_n4335) & (n_n4334) & (x469x) & (!x15152x)) + ((x198x) & (!n_n4335) & (n_n4334) & (x469x) & (x15152x)) + ((x198x) & (n_n4335) & (!n_n4334) & (!x469x) & (!x15152x)) + ((x198x) & (n_n4335) & (!n_n4334) & (!x469x) & (x15152x)) + ((x198x) & (n_n4335) & (!n_n4334) & (x469x) & (!x15152x)) + ((x198x) & (n_n4335) & (!n_n4334) & (x469x) & (x15152x)) + ((x198x) & (n_n4335) & (n_n4334) & (!x469x) & (!x15152x)) + ((x198x) & (n_n4335) & (n_n4334) & (!x469x) & (x15152x)) + ((x198x) & (n_n4335) & (n_n4334) & (x469x) & (!x15152x)) + ((x198x) & (n_n4335) & (n_n4334) & (x469x) & (x15152x)));
	assign n_n4322 = (((i_9_) & (n_n536) & (n_n524) & (n_n535)));
	assign x22098x = (((!n_n4324) & (!n_n4319) & (!n_n4326) & (!n_n4321)));
	assign n_n2641 = (((!n_n4325) & (!n_n4327) & (!x283x) & (!n_n4322) & (!x22098x)) + ((!n_n4325) & (!n_n4327) & (!x283x) & (n_n4322) & (!x22098x)) + ((!n_n4325) & (!n_n4327) & (!x283x) & (n_n4322) & (x22098x)) + ((!n_n4325) & (!n_n4327) & (x283x) & (!n_n4322) & (!x22098x)) + ((!n_n4325) & (!n_n4327) & (x283x) & (!n_n4322) & (x22098x)) + ((!n_n4325) & (!n_n4327) & (x283x) & (n_n4322) & (!x22098x)) + ((!n_n4325) & (!n_n4327) & (x283x) & (n_n4322) & (x22098x)) + ((!n_n4325) & (n_n4327) & (!x283x) & (!n_n4322) & (!x22098x)) + ((!n_n4325) & (n_n4327) & (!x283x) & (!n_n4322) & (x22098x)) + ((!n_n4325) & (n_n4327) & (!x283x) & (n_n4322) & (!x22098x)) + ((!n_n4325) & (n_n4327) & (!x283x) & (n_n4322) & (x22098x)) + ((!n_n4325) & (n_n4327) & (x283x) & (!n_n4322) & (!x22098x)) + ((!n_n4325) & (n_n4327) & (x283x) & (!n_n4322) & (x22098x)) + ((!n_n4325) & (n_n4327) & (x283x) & (n_n4322) & (!x22098x)) + ((!n_n4325) & (n_n4327) & (x283x) & (n_n4322) & (x22098x)) + ((n_n4325) & (!n_n4327) & (!x283x) & (!n_n4322) & (!x22098x)) + ((n_n4325) & (!n_n4327) & (!x283x) & (!n_n4322) & (x22098x)) + ((n_n4325) & (!n_n4327) & (!x283x) & (n_n4322) & (!x22098x)) + ((n_n4325) & (!n_n4327) & (!x283x) & (n_n4322) & (x22098x)) + ((n_n4325) & (!n_n4327) & (x283x) & (!n_n4322) & (!x22098x)) + ((n_n4325) & (!n_n4327) & (x283x) & (!n_n4322) & (x22098x)) + ((n_n4325) & (!n_n4327) & (x283x) & (n_n4322) & (!x22098x)) + ((n_n4325) & (!n_n4327) & (x283x) & (n_n4322) & (x22098x)) + ((n_n4325) & (n_n4327) & (!x283x) & (!n_n4322) & (!x22098x)) + ((n_n4325) & (n_n4327) & (!x283x) & (!n_n4322) & (x22098x)) + ((n_n4325) & (n_n4327) & (!x283x) & (n_n4322) & (!x22098x)) + ((n_n4325) & (n_n4327) & (!x283x) & (n_n4322) & (x22098x)) + ((n_n4325) & (n_n4327) & (x283x) & (!n_n4322) & (!x22098x)) + ((n_n4325) & (n_n4327) & (x283x) & (!n_n4322) & (x22098x)) + ((n_n4325) & (n_n4327) & (x283x) & (n_n4322) & (!x22098x)) + ((n_n4325) & (n_n4327) & (x283x) & (n_n4322) & (x22098x)));
	assign x337x = (((!i_9_) & (n_n536) & (!n_n532) & (n_n534) & (n_n509)) + ((!i_9_) & (n_n536) & (n_n532) & (n_n534) & (n_n509)) + ((i_9_) & (n_n536) & (n_n532) & (!n_n534) & (n_n509)) + ((i_9_) & (n_n536) & (n_n532) & (n_n534) & (n_n509)));
	assign n_n5248 = (((i_7_) & (i_8_) & (!i_6_) & (x19x) & (n_n509)));
	assign n_n5192 = (((i_7_) & (i_8_) & (i_6_) & (x12x) & (n_n464)));
	assign x22199x = (((!x12x) & (!n_n5183) & (!x506x) & (!n_n5191) & (!n_n5192)) + ((!x12x) & (!n_n5183) & (x506x) & (!n_n5191) & (!n_n5192)) + ((x12x) & (!n_n5183) & (!x506x) & (!n_n5191) & (!n_n5192)));
	assign n_n5195 = (((!i_9_) & (n_n532) & (n_n130) & (n_n464)));
	assign n_n5208 = (((i_7_) & (i_8_) & (i_6_) & (x19x) & (n_n535)));
	assign x36x = (((!n_n524) & (!x12x) & (!n_n464) & (n_n5201)) + ((!n_n524) & (!x12x) & (n_n464) & (n_n5201)) + ((!n_n524) & (x12x) & (!n_n464) & (n_n5201)) + ((!n_n524) & (x12x) & (n_n464) & (n_n5201)) + ((n_n524) & (!x12x) & (!n_n464) & (n_n5201)) + ((n_n524) & (!x12x) & (n_n464) & (n_n5201)) + ((n_n524) & (x12x) & (!n_n464) & (n_n5201)) + ((n_n524) & (x12x) & (n_n464) & (!n_n5201)) + ((n_n524) & (x12x) & (n_n464) & (n_n5201)));
	assign x451x = (((!i_7_) & (i_8_) & (i_6_) & (x12x) & (n_n464)) + ((i_7_) & (!i_8_) & (i_6_) & (x12x) & (n_n464)));
	assign x22065x = (((!n_n4998) & (!n_n4999) & (!n_n4994) & (!n_n5004)));
	assign x133x = (((!i_9_) & (n_n532) & (n_n509) & (n_n195) & (!n_n530)) + ((!i_9_) & (n_n532) & (n_n509) & (n_n195) & (n_n530)) + ((i_9_) & (!n_n532) & (n_n509) & (n_n195) & (n_n530)) + ((i_9_) & (n_n532) & (n_n509) & (n_n195) & (n_n530)));
	assign n_n1532 = (((!i_9_) & (!n_n535) & (!n_n530) & (!n_n65) & (x223x)) + ((!i_9_) & (!n_n535) & (!n_n530) & (n_n65) & (x223x)) + ((!i_9_) & (!n_n535) & (n_n530) & (!n_n65) & (x223x)) + ((!i_9_) & (!n_n535) & (n_n530) & (n_n65) & (x223x)) + ((!i_9_) & (n_n535) & (!n_n530) & (!n_n65) & (x223x)) + ((!i_9_) & (n_n535) & (!n_n530) & (n_n65) & (x223x)) + ((!i_9_) & (n_n535) & (n_n530) & (!n_n65) & (x223x)) + ((!i_9_) & (n_n535) & (n_n530) & (n_n65) & (!x223x)) + ((!i_9_) & (n_n535) & (n_n530) & (n_n65) & (x223x)) + ((i_9_) & (!n_n535) & (!n_n530) & (!n_n65) & (x223x)) + ((i_9_) & (!n_n535) & (!n_n530) & (n_n65) & (x223x)) + ((i_9_) & (!n_n535) & (n_n530) & (!n_n65) & (x223x)) + ((i_9_) & (!n_n535) & (n_n530) & (n_n65) & (x223x)) + ((i_9_) & (n_n535) & (!n_n530) & (!n_n65) & (x223x)) + ((i_9_) & (n_n535) & (!n_n530) & (n_n65) & (x223x)) + ((i_9_) & (n_n535) & (n_n530) & (!n_n65) & (x223x)) + ((i_9_) & (n_n535) & (n_n530) & (n_n65) & (x223x)));
	assign x12265x = (((!n_n520) & (!x12x) & (!n_n500) & (!n_n5143) & (x211x)) + ((!n_n520) & (!x12x) & (!n_n500) & (n_n5143) & (!x211x)) + ((!n_n520) & (!x12x) & (!n_n500) & (n_n5143) & (x211x)) + ((!n_n520) & (!x12x) & (n_n500) & (!n_n5143) & (x211x)) + ((!n_n520) & (!x12x) & (n_n500) & (n_n5143) & (!x211x)) + ((!n_n520) & (!x12x) & (n_n500) & (n_n5143) & (x211x)) + ((!n_n520) & (x12x) & (!n_n500) & (!n_n5143) & (x211x)) + ((!n_n520) & (x12x) & (!n_n500) & (n_n5143) & (!x211x)) + ((!n_n520) & (x12x) & (!n_n500) & (n_n5143) & (x211x)) + ((!n_n520) & (x12x) & (n_n500) & (!n_n5143) & (x211x)) + ((!n_n520) & (x12x) & (n_n500) & (n_n5143) & (!x211x)) + ((!n_n520) & (x12x) & (n_n500) & (n_n5143) & (x211x)) + ((n_n520) & (!x12x) & (!n_n500) & (!n_n5143) & (x211x)) + ((n_n520) & (!x12x) & (!n_n500) & (n_n5143) & (!x211x)) + ((n_n520) & (!x12x) & (!n_n500) & (n_n5143) & (x211x)) + ((n_n520) & (!x12x) & (n_n500) & (!n_n5143) & (x211x)) + ((n_n520) & (!x12x) & (n_n500) & (n_n5143) & (!x211x)) + ((n_n520) & (!x12x) & (n_n500) & (n_n5143) & (x211x)) + ((n_n520) & (x12x) & (!n_n500) & (!n_n5143) & (x211x)) + ((n_n520) & (x12x) & (!n_n500) & (n_n5143) & (!x211x)) + ((n_n520) & (x12x) & (!n_n500) & (n_n5143) & (x211x)) + ((n_n520) & (x12x) & (n_n500) & (!n_n5143) & (!x211x)) + ((n_n520) & (x12x) & (n_n500) & (!n_n5143) & (x211x)) + ((n_n520) & (x12x) & (n_n500) & (n_n5143) & (!x211x)) + ((n_n520) & (x12x) & (n_n500) & (n_n5143) & (x211x)));
	assign n_n1444 = (((!n_n5135) & (!n_n5148) & (!x125x) & (!n_n5144) & (x12265x)) + ((!n_n5135) & (!n_n5148) & (!x125x) & (n_n5144) & (!x12265x)) + ((!n_n5135) & (!n_n5148) & (!x125x) & (n_n5144) & (x12265x)) + ((!n_n5135) & (!n_n5148) & (x125x) & (!n_n5144) & (!x12265x)) + ((!n_n5135) & (!n_n5148) & (x125x) & (!n_n5144) & (x12265x)) + ((!n_n5135) & (!n_n5148) & (x125x) & (n_n5144) & (!x12265x)) + ((!n_n5135) & (!n_n5148) & (x125x) & (n_n5144) & (x12265x)) + ((!n_n5135) & (n_n5148) & (!x125x) & (!n_n5144) & (!x12265x)) + ((!n_n5135) & (n_n5148) & (!x125x) & (!n_n5144) & (x12265x)) + ((!n_n5135) & (n_n5148) & (!x125x) & (n_n5144) & (!x12265x)) + ((!n_n5135) & (n_n5148) & (!x125x) & (n_n5144) & (x12265x)) + ((!n_n5135) & (n_n5148) & (x125x) & (!n_n5144) & (!x12265x)) + ((!n_n5135) & (n_n5148) & (x125x) & (!n_n5144) & (x12265x)) + ((!n_n5135) & (n_n5148) & (x125x) & (n_n5144) & (!x12265x)) + ((!n_n5135) & (n_n5148) & (x125x) & (n_n5144) & (x12265x)) + ((n_n5135) & (!n_n5148) & (!x125x) & (!n_n5144) & (!x12265x)) + ((n_n5135) & (!n_n5148) & (!x125x) & (!n_n5144) & (x12265x)) + ((n_n5135) & (!n_n5148) & (!x125x) & (n_n5144) & (!x12265x)) + ((n_n5135) & (!n_n5148) & (!x125x) & (n_n5144) & (x12265x)) + ((n_n5135) & (!n_n5148) & (x125x) & (!n_n5144) & (!x12265x)) + ((n_n5135) & (!n_n5148) & (x125x) & (!n_n5144) & (x12265x)) + ((n_n5135) & (!n_n5148) & (x125x) & (n_n5144) & (!x12265x)) + ((n_n5135) & (!n_n5148) & (x125x) & (n_n5144) & (x12265x)) + ((n_n5135) & (n_n5148) & (!x125x) & (!n_n5144) & (!x12265x)) + ((n_n5135) & (n_n5148) & (!x125x) & (!n_n5144) & (x12265x)) + ((n_n5135) & (n_n5148) & (!x125x) & (n_n5144) & (!x12265x)) + ((n_n5135) & (n_n5148) & (!x125x) & (n_n5144) & (x12265x)) + ((n_n5135) & (n_n5148) & (x125x) & (!n_n5144) & (!x12265x)) + ((n_n5135) & (n_n5148) & (x125x) & (!n_n5144) & (x12265x)) + ((n_n5135) & (n_n5148) & (x125x) & (n_n5144) & (!x12265x)) + ((n_n5135) & (n_n5148) & (x125x) & (n_n5144) & (x12265x)));
	assign x446x = (((!i_9_) & (!x19x) & (n_n526) & (n_n509) & (n_n65)) + ((!i_9_) & (x19x) & (n_n526) & (n_n509) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n526) & (n_n509) & (n_n65)) + ((i_9_) & (x19x) & (n_n526) & (n_n509) & (!n_n65)) + ((i_9_) & (x19x) & (n_n526) & (n_n509) & (n_n65)));
	assign x12349x = (((!n_n5247) & (!n_n5251) & (!n_n5252) & (!n_n5250) & (n_n5257)) + ((!n_n5247) & (!n_n5251) & (!n_n5252) & (n_n5250) & (!n_n5257)) + ((!n_n5247) & (!n_n5251) & (!n_n5252) & (n_n5250) & (n_n5257)) + ((!n_n5247) & (!n_n5251) & (n_n5252) & (!n_n5250) & (!n_n5257)) + ((!n_n5247) & (!n_n5251) & (n_n5252) & (!n_n5250) & (n_n5257)) + ((!n_n5247) & (!n_n5251) & (n_n5252) & (n_n5250) & (!n_n5257)) + ((!n_n5247) & (!n_n5251) & (n_n5252) & (n_n5250) & (n_n5257)) + ((!n_n5247) & (n_n5251) & (!n_n5252) & (!n_n5250) & (!n_n5257)) + ((!n_n5247) & (n_n5251) & (!n_n5252) & (!n_n5250) & (n_n5257)) + ((!n_n5247) & (n_n5251) & (!n_n5252) & (n_n5250) & (!n_n5257)) + ((!n_n5247) & (n_n5251) & (!n_n5252) & (n_n5250) & (n_n5257)) + ((!n_n5247) & (n_n5251) & (n_n5252) & (!n_n5250) & (!n_n5257)) + ((!n_n5247) & (n_n5251) & (n_n5252) & (!n_n5250) & (n_n5257)) + ((!n_n5247) & (n_n5251) & (n_n5252) & (n_n5250) & (!n_n5257)) + ((!n_n5247) & (n_n5251) & (n_n5252) & (n_n5250) & (n_n5257)) + ((n_n5247) & (!n_n5251) & (!n_n5252) & (!n_n5250) & (!n_n5257)) + ((n_n5247) & (!n_n5251) & (!n_n5252) & (!n_n5250) & (n_n5257)) + ((n_n5247) & (!n_n5251) & (!n_n5252) & (n_n5250) & (!n_n5257)) + ((n_n5247) & (!n_n5251) & (!n_n5252) & (n_n5250) & (n_n5257)) + ((n_n5247) & (!n_n5251) & (n_n5252) & (!n_n5250) & (!n_n5257)) + ((n_n5247) & (!n_n5251) & (n_n5252) & (!n_n5250) & (n_n5257)) + ((n_n5247) & (!n_n5251) & (n_n5252) & (n_n5250) & (!n_n5257)) + ((n_n5247) & (!n_n5251) & (n_n5252) & (n_n5250) & (n_n5257)) + ((n_n5247) & (n_n5251) & (!n_n5252) & (!n_n5250) & (!n_n5257)) + ((n_n5247) & (n_n5251) & (!n_n5252) & (!n_n5250) & (n_n5257)) + ((n_n5247) & (n_n5251) & (!n_n5252) & (n_n5250) & (!n_n5257)) + ((n_n5247) & (n_n5251) & (!n_n5252) & (n_n5250) & (n_n5257)) + ((n_n5247) & (n_n5251) & (n_n5252) & (!n_n5250) & (!n_n5257)) + ((n_n5247) & (n_n5251) & (n_n5252) & (!n_n5250) & (n_n5257)) + ((n_n5247) & (n_n5251) & (n_n5252) & (n_n5250) & (!n_n5257)) + ((n_n5247) & (n_n5251) & (n_n5252) & (n_n5250) & (n_n5257)));
	assign n_n1435 = (((!n_n5254) & (!n_n5249) & (!n_n5259) & (!n_n5248) & (x12349x)) + ((!n_n5254) & (!n_n5249) & (!n_n5259) & (n_n5248) & (!x12349x)) + ((!n_n5254) & (!n_n5249) & (!n_n5259) & (n_n5248) & (x12349x)) + ((!n_n5254) & (!n_n5249) & (n_n5259) & (!n_n5248) & (!x12349x)) + ((!n_n5254) & (!n_n5249) & (n_n5259) & (!n_n5248) & (x12349x)) + ((!n_n5254) & (!n_n5249) & (n_n5259) & (n_n5248) & (!x12349x)) + ((!n_n5254) & (!n_n5249) & (n_n5259) & (n_n5248) & (x12349x)) + ((!n_n5254) & (n_n5249) & (!n_n5259) & (!n_n5248) & (!x12349x)) + ((!n_n5254) & (n_n5249) & (!n_n5259) & (!n_n5248) & (x12349x)) + ((!n_n5254) & (n_n5249) & (!n_n5259) & (n_n5248) & (!x12349x)) + ((!n_n5254) & (n_n5249) & (!n_n5259) & (n_n5248) & (x12349x)) + ((!n_n5254) & (n_n5249) & (n_n5259) & (!n_n5248) & (!x12349x)) + ((!n_n5254) & (n_n5249) & (n_n5259) & (!n_n5248) & (x12349x)) + ((!n_n5254) & (n_n5249) & (n_n5259) & (n_n5248) & (!x12349x)) + ((!n_n5254) & (n_n5249) & (n_n5259) & (n_n5248) & (x12349x)) + ((n_n5254) & (!n_n5249) & (!n_n5259) & (!n_n5248) & (!x12349x)) + ((n_n5254) & (!n_n5249) & (!n_n5259) & (!n_n5248) & (x12349x)) + ((n_n5254) & (!n_n5249) & (!n_n5259) & (n_n5248) & (!x12349x)) + ((n_n5254) & (!n_n5249) & (!n_n5259) & (n_n5248) & (x12349x)) + ((n_n5254) & (!n_n5249) & (n_n5259) & (!n_n5248) & (!x12349x)) + ((n_n5254) & (!n_n5249) & (n_n5259) & (!n_n5248) & (x12349x)) + ((n_n5254) & (!n_n5249) & (n_n5259) & (n_n5248) & (!x12349x)) + ((n_n5254) & (!n_n5249) & (n_n5259) & (n_n5248) & (x12349x)) + ((n_n5254) & (n_n5249) & (!n_n5259) & (!n_n5248) & (!x12349x)) + ((n_n5254) & (n_n5249) & (!n_n5259) & (!n_n5248) & (x12349x)) + ((n_n5254) & (n_n5249) & (!n_n5259) & (n_n5248) & (!x12349x)) + ((n_n5254) & (n_n5249) & (!n_n5259) & (n_n5248) & (x12349x)) + ((n_n5254) & (n_n5249) & (n_n5259) & (!n_n5248) & (!x12349x)) + ((n_n5254) & (n_n5249) & (n_n5259) & (!n_n5248) & (x12349x)) + ((n_n5254) & (n_n5249) & (n_n5259) & (n_n5248) & (!x12349x)) + ((n_n5254) & (n_n5249) & (n_n5259) & (n_n5248) & (x12349x)));
	assign x11542x = (((!n_n455) & (!x24x) & (!n_n464) & (!n_n4556) & (x82x)) + ((!n_n455) & (!x24x) & (!n_n464) & (n_n4556) & (!x82x)) + ((!n_n455) & (!x24x) & (!n_n464) & (n_n4556) & (x82x)) + ((!n_n455) & (!x24x) & (n_n464) & (!n_n4556) & (x82x)) + ((!n_n455) & (!x24x) & (n_n464) & (n_n4556) & (!x82x)) + ((!n_n455) & (!x24x) & (n_n464) & (n_n4556) & (x82x)) + ((!n_n455) & (x24x) & (!n_n464) & (!n_n4556) & (x82x)) + ((!n_n455) & (x24x) & (!n_n464) & (n_n4556) & (!x82x)) + ((!n_n455) & (x24x) & (!n_n464) & (n_n4556) & (x82x)) + ((!n_n455) & (x24x) & (n_n464) & (!n_n4556) & (x82x)) + ((!n_n455) & (x24x) & (n_n464) & (n_n4556) & (!x82x)) + ((!n_n455) & (x24x) & (n_n464) & (n_n4556) & (x82x)) + ((n_n455) & (!x24x) & (!n_n464) & (!n_n4556) & (x82x)) + ((n_n455) & (!x24x) & (!n_n464) & (n_n4556) & (!x82x)) + ((n_n455) & (!x24x) & (!n_n464) & (n_n4556) & (x82x)) + ((n_n455) & (!x24x) & (n_n464) & (!n_n4556) & (x82x)) + ((n_n455) & (!x24x) & (n_n464) & (n_n4556) & (!x82x)) + ((n_n455) & (!x24x) & (n_n464) & (n_n4556) & (x82x)) + ((n_n455) & (x24x) & (!n_n464) & (!n_n4556) & (x82x)) + ((n_n455) & (x24x) & (!n_n464) & (n_n4556) & (!x82x)) + ((n_n455) & (x24x) & (!n_n464) & (n_n4556) & (x82x)) + ((n_n455) & (x24x) & (n_n464) & (!n_n4556) & (!x82x)) + ((n_n455) & (x24x) & (n_n464) & (!n_n4556) & (x82x)) + ((n_n455) & (x24x) & (n_n464) & (n_n4556) & (!x82x)) + ((n_n455) & (x24x) & (n_n464) & (n_n4556) & (x82x)));
	assign n_n1636 = (((!i_9_) & (n_n390) & (!n_n532) & (n_n534) & (n_n464)) + ((!i_9_) & (n_n390) & (n_n532) & (n_n534) & (n_n464)) + ((i_9_) & (n_n390) & (!n_n532) & (n_n534) & (n_n464)) + ((i_9_) & (n_n390) & (n_n532) & (!n_n534) & (n_n464)) + ((i_9_) & (n_n390) & (n_n532) & (n_n534) & (n_n464)));
	assign x22152x = (((!n_n5014) & (!n_n5015) & (!n_n5007) & (!n_n5012) & (!n_n5009)));
	assign n_n1067 = (((!n_n5017) & (!n_n5019) & (!n_n5020) & (!n_n5010) & (!x22152x)) + ((!n_n5017) & (!n_n5019) & (!n_n5020) & (n_n5010) & (!x22152x)) + ((!n_n5017) & (!n_n5019) & (!n_n5020) & (n_n5010) & (x22152x)) + ((!n_n5017) & (!n_n5019) & (n_n5020) & (!n_n5010) & (!x22152x)) + ((!n_n5017) & (!n_n5019) & (n_n5020) & (!n_n5010) & (x22152x)) + ((!n_n5017) & (!n_n5019) & (n_n5020) & (n_n5010) & (!x22152x)) + ((!n_n5017) & (!n_n5019) & (n_n5020) & (n_n5010) & (x22152x)) + ((!n_n5017) & (n_n5019) & (!n_n5020) & (!n_n5010) & (!x22152x)) + ((!n_n5017) & (n_n5019) & (!n_n5020) & (!n_n5010) & (x22152x)) + ((!n_n5017) & (n_n5019) & (!n_n5020) & (n_n5010) & (!x22152x)) + ((!n_n5017) & (n_n5019) & (!n_n5020) & (n_n5010) & (x22152x)) + ((!n_n5017) & (n_n5019) & (n_n5020) & (!n_n5010) & (!x22152x)) + ((!n_n5017) & (n_n5019) & (n_n5020) & (!n_n5010) & (x22152x)) + ((!n_n5017) & (n_n5019) & (n_n5020) & (n_n5010) & (!x22152x)) + ((!n_n5017) & (n_n5019) & (n_n5020) & (n_n5010) & (x22152x)) + ((n_n5017) & (!n_n5019) & (!n_n5020) & (!n_n5010) & (!x22152x)) + ((n_n5017) & (!n_n5019) & (!n_n5020) & (!n_n5010) & (x22152x)) + ((n_n5017) & (!n_n5019) & (!n_n5020) & (n_n5010) & (!x22152x)) + ((n_n5017) & (!n_n5019) & (!n_n5020) & (n_n5010) & (x22152x)) + ((n_n5017) & (!n_n5019) & (n_n5020) & (!n_n5010) & (!x22152x)) + ((n_n5017) & (!n_n5019) & (n_n5020) & (!n_n5010) & (x22152x)) + ((n_n5017) & (!n_n5019) & (n_n5020) & (n_n5010) & (!x22152x)) + ((n_n5017) & (!n_n5019) & (n_n5020) & (n_n5010) & (x22152x)) + ((n_n5017) & (n_n5019) & (!n_n5020) & (!n_n5010) & (!x22152x)) + ((n_n5017) & (n_n5019) & (!n_n5020) & (!n_n5010) & (x22152x)) + ((n_n5017) & (n_n5019) & (!n_n5020) & (n_n5010) & (!x22152x)) + ((n_n5017) & (n_n5019) & (!n_n5020) & (n_n5010) & (x22152x)) + ((n_n5017) & (n_n5019) & (n_n5020) & (!n_n5010) & (!x22152x)) + ((n_n5017) & (n_n5019) & (n_n5020) & (!n_n5010) & (x22152x)) + ((n_n5017) & (n_n5019) & (n_n5020) & (n_n5010) & (!x22152x)) + ((n_n5017) & (n_n5019) & (n_n5020) & (n_n5010) & (x22152x)));
	assign x181x = (((!i_9_) & (!x19x) & (n_n518) & (n_n530) & (n_n65)) + ((!i_9_) & (x19x) & (n_n518) & (n_n530) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n518) & (n_n530) & (n_n65)) + ((i_9_) & (x19x) & (n_n518) & (n_n530) & (!n_n65)) + ((i_9_) & (x19x) & (n_n518) & (n_n530) & (n_n65)));
	assign x22157x = (((!n_n5212) & (!n_n5220) & (!n_n5226) & (!n_n5225)));
	assign x453x = (((!i_9_) & (!n_n532) & (n_n534) & (n_n130) & (n_n464)) + ((!i_9_) & (n_n532) & (!n_n534) & (n_n130) & (n_n464)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n130) & (n_n464)));
	assign n_n1927 = (((!n_n532) & (!x12x) & (!n_n464) & (x453x)) + ((!n_n532) & (!x12x) & (n_n464) & (x453x)) + ((!n_n532) & (x12x) & (!n_n464) & (x453x)) + ((!n_n532) & (x12x) & (n_n464) & (x453x)) + ((n_n532) & (!x12x) & (!n_n464) & (x453x)) + ((n_n532) & (!x12x) & (n_n464) & (x453x)) + ((n_n532) & (x12x) & (!n_n464) & (x453x)) + ((n_n532) & (x12x) & (n_n464) & (!x453x)) + ((n_n532) & (x12x) & (n_n464) & (x453x)));
	assign x188x = (((n_n473) & (!n_n520) & (n_n130) & (!x12x) & (x20x)) + ((n_n473) & (!n_n520) & (n_n130) & (x12x) & (x20x)) + ((n_n473) & (n_n520) & (!n_n130) & (x12x) & (!x20x)) + ((n_n473) & (n_n520) & (!n_n130) & (x12x) & (x20x)) + ((n_n473) & (n_n520) & (n_n130) & (!x12x) & (x20x)) + ((n_n473) & (n_n520) & (n_n130) & (x12x) & (!x20x)) + ((n_n473) & (n_n520) & (n_n130) & (x12x) & (x20x)));
	assign x452x = (((!i_7_) & (!i_8_) & (i_6_) & (x12x) & (n_n464)) + ((!i_7_) & (i_8_) & (i_6_) & (x12x) & (n_n464)));
	assign x11976x = (((!n_n5204) & (!n_n5210) & (!n_n5205) & (!n_n5211) & (n_n5208)) + ((!n_n5204) & (!n_n5210) & (!n_n5205) & (n_n5211) & (!n_n5208)) + ((!n_n5204) & (!n_n5210) & (!n_n5205) & (n_n5211) & (n_n5208)) + ((!n_n5204) & (!n_n5210) & (n_n5205) & (!n_n5211) & (!n_n5208)) + ((!n_n5204) & (!n_n5210) & (n_n5205) & (!n_n5211) & (n_n5208)) + ((!n_n5204) & (!n_n5210) & (n_n5205) & (n_n5211) & (!n_n5208)) + ((!n_n5204) & (!n_n5210) & (n_n5205) & (n_n5211) & (n_n5208)) + ((!n_n5204) & (n_n5210) & (!n_n5205) & (!n_n5211) & (!n_n5208)) + ((!n_n5204) & (n_n5210) & (!n_n5205) & (!n_n5211) & (n_n5208)) + ((!n_n5204) & (n_n5210) & (!n_n5205) & (n_n5211) & (!n_n5208)) + ((!n_n5204) & (n_n5210) & (!n_n5205) & (n_n5211) & (n_n5208)) + ((!n_n5204) & (n_n5210) & (n_n5205) & (!n_n5211) & (!n_n5208)) + ((!n_n5204) & (n_n5210) & (n_n5205) & (!n_n5211) & (n_n5208)) + ((!n_n5204) & (n_n5210) & (n_n5205) & (n_n5211) & (!n_n5208)) + ((!n_n5204) & (n_n5210) & (n_n5205) & (n_n5211) & (n_n5208)) + ((n_n5204) & (!n_n5210) & (!n_n5205) & (!n_n5211) & (!n_n5208)) + ((n_n5204) & (!n_n5210) & (!n_n5205) & (!n_n5211) & (n_n5208)) + ((n_n5204) & (!n_n5210) & (!n_n5205) & (n_n5211) & (!n_n5208)) + ((n_n5204) & (!n_n5210) & (!n_n5205) & (n_n5211) & (n_n5208)) + ((n_n5204) & (!n_n5210) & (n_n5205) & (!n_n5211) & (!n_n5208)) + ((n_n5204) & (!n_n5210) & (n_n5205) & (!n_n5211) & (n_n5208)) + ((n_n5204) & (!n_n5210) & (n_n5205) & (n_n5211) & (!n_n5208)) + ((n_n5204) & (!n_n5210) & (n_n5205) & (n_n5211) & (n_n5208)) + ((n_n5204) & (n_n5210) & (!n_n5205) & (!n_n5211) & (!n_n5208)) + ((n_n5204) & (n_n5210) & (!n_n5205) & (!n_n5211) & (n_n5208)) + ((n_n5204) & (n_n5210) & (!n_n5205) & (n_n5211) & (!n_n5208)) + ((n_n5204) & (n_n5210) & (!n_n5205) & (n_n5211) & (n_n5208)) + ((n_n5204) & (n_n5210) & (n_n5205) & (!n_n5211) & (!n_n5208)) + ((n_n5204) & (n_n5210) & (n_n5205) & (!n_n5211) & (n_n5208)) + ((n_n5204) & (n_n5210) & (n_n5205) & (n_n5211) & (!n_n5208)) + ((n_n5204) & (n_n5210) & (n_n5205) & (n_n5211) & (n_n5208)));
	assign x22164x = (((!n_n4432) & (!n_n4438) & (!x236x) & (!n_n4435)));
	assign x22162x = (((!n_n4521) & (!n_n4504) & (!n_n4517) & (!n_n4497)));
	assign n_n1111 = (((!n_n4459) & (!n_n4461) & (!x147x) & (!n_n4462) & (!x22166x)) + ((!n_n4459) & (!n_n4461) & (!x147x) & (n_n4462) & (!x22166x)) + ((!n_n4459) & (!n_n4461) & (!x147x) & (n_n4462) & (x22166x)) + ((!n_n4459) & (!n_n4461) & (x147x) & (!n_n4462) & (!x22166x)) + ((!n_n4459) & (!n_n4461) & (x147x) & (!n_n4462) & (x22166x)) + ((!n_n4459) & (!n_n4461) & (x147x) & (n_n4462) & (!x22166x)) + ((!n_n4459) & (!n_n4461) & (x147x) & (n_n4462) & (x22166x)) + ((!n_n4459) & (n_n4461) & (!x147x) & (!n_n4462) & (!x22166x)) + ((!n_n4459) & (n_n4461) & (!x147x) & (!n_n4462) & (x22166x)) + ((!n_n4459) & (n_n4461) & (!x147x) & (n_n4462) & (!x22166x)) + ((!n_n4459) & (n_n4461) & (!x147x) & (n_n4462) & (x22166x)) + ((!n_n4459) & (n_n4461) & (x147x) & (!n_n4462) & (!x22166x)) + ((!n_n4459) & (n_n4461) & (x147x) & (!n_n4462) & (x22166x)) + ((!n_n4459) & (n_n4461) & (x147x) & (n_n4462) & (!x22166x)) + ((!n_n4459) & (n_n4461) & (x147x) & (n_n4462) & (x22166x)) + ((n_n4459) & (!n_n4461) & (!x147x) & (!n_n4462) & (!x22166x)) + ((n_n4459) & (!n_n4461) & (!x147x) & (!n_n4462) & (x22166x)) + ((n_n4459) & (!n_n4461) & (!x147x) & (n_n4462) & (!x22166x)) + ((n_n4459) & (!n_n4461) & (!x147x) & (n_n4462) & (x22166x)) + ((n_n4459) & (!n_n4461) & (x147x) & (!n_n4462) & (!x22166x)) + ((n_n4459) & (!n_n4461) & (x147x) & (!n_n4462) & (x22166x)) + ((n_n4459) & (!n_n4461) & (x147x) & (n_n4462) & (!x22166x)) + ((n_n4459) & (!n_n4461) & (x147x) & (n_n4462) & (x22166x)) + ((n_n4459) & (n_n4461) & (!x147x) & (!n_n4462) & (!x22166x)) + ((n_n4459) & (n_n4461) & (!x147x) & (!n_n4462) & (x22166x)) + ((n_n4459) & (n_n4461) & (!x147x) & (n_n4462) & (!x22166x)) + ((n_n4459) & (n_n4461) & (!x147x) & (n_n4462) & (x22166x)) + ((n_n4459) & (n_n4461) & (x147x) & (!n_n4462) & (!x22166x)) + ((n_n4459) & (n_n4461) & (x147x) & (!n_n4462) & (x22166x)) + ((n_n4459) & (n_n4461) & (x147x) & (n_n4462) & (!x22166x)) + ((n_n4459) & (n_n4461) & (x147x) & (n_n4462) & (x22166x)));
	assign x11516x = (((!n_n4473) & (!n_n4471) & (!n_n4472) & (n_n4487)) + ((!n_n4473) & (!n_n4471) & (n_n4472) & (!n_n4487)) + ((!n_n4473) & (!n_n4471) & (n_n4472) & (n_n4487)) + ((!n_n4473) & (n_n4471) & (!n_n4472) & (!n_n4487)) + ((!n_n4473) & (n_n4471) & (!n_n4472) & (n_n4487)) + ((!n_n4473) & (n_n4471) & (n_n4472) & (!n_n4487)) + ((!n_n4473) & (n_n4471) & (n_n4472) & (n_n4487)) + ((n_n4473) & (!n_n4471) & (!n_n4472) & (!n_n4487)) + ((n_n4473) & (!n_n4471) & (!n_n4472) & (n_n4487)) + ((n_n4473) & (!n_n4471) & (n_n4472) & (!n_n4487)) + ((n_n4473) & (!n_n4471) & (n_n4472) & (n_n4487)) + ((n_n4473) & (n_n4471) & (!n_n4472) & (!n_n4487)) + ((n_n4473) & (n_n4471) & (!n_n4472) & (n_n4487)) + ((n_n4473) & (n_n4471) & (n_n4472) & (!n_n4487)) + ((n_n4473) & (n_n4471) & (n_n4472) & (n_n4487)));
	assign x11517x = (((!n_n4470) & (!n_n4475) & (!n_n4469) & (!n_n4465) & (x11505x)) + ((!n_n4470) & (!n_n4475) & (!n_n4469) & (n_n4465) & (!x11505x)) + ((!n_n4470) & (!n_n4475) & (!n_n4469) & (n_n4465) & (x11505x)) + ((!n_n4470) & (!n_n4475) & (n_n4469) & (!n_n4465) & (!x11505x)) + ((!n_n4470) & (!n_n4475) & (n_n4469) & (!n_n4465) & (x11505x)) + ((!n_n4470) & (!n_n4475) & (n_n4469) & (n_n4465) & (!x11505x)) + ((!n_n4470) & (!n_n4475) & (n_n4469) & (n_n4465) & (x11505x)) + ((!n_n4470) & (n_n4475) & (!n_n4469) & (!n_n4465) & (!x11505x)) + ((!n_n4470) & (n_n4475) & (!n_n4469) & (!n_n4465) & (x11505x)) + ((!n_n4470) & (n_n4475) & (!n_n4469) & (n_n4465) & (!x11505x)) + ((!n_n4470) & (n_n4475) & (!n_n4469) & (n_n4465) & (x11505x)) + ((!n_n4470) & (n_n4475) & (n_n4469) & (!n_n4465) & (!x11505x)) + ((!n_n4470) & (n_n4475) & (n_n4469) & (!n_n4465) & (x11505x)) + ((!n_n4470) & (n_n4475) & (n_n4469) & (n_n4465) & (!x11505x)) + ((!n_n4470) & (n_n4475) & (n_n4469) & (n_n4465) & (x11505x)) + ((n_n4470) & (!n_n4475) & (!n_n4469) & (!n_n4465) & (!x11505x)) + ((n_n4470) & (!n_n4475) & (!n_n4469) & (!n_n4465) & (x11505x)) + ((n_n4470) & (!n_n4475) & (!n_n4469) & (n_n4465) & (!x11505x)) + ((n_n4470) & (!n_n4475) & (!n_n4469) & (n_n4465) & (x11505x)) + ((n_n4470) & (!n_n4475) & (n_n4469) & (!n_n4465) & (!x11505x)) + ((n_n4470) & (!n_n4475) & (n_n4469) & (!n_n4465) & (x11505x)) + ((n_n4470) & (!n_n4475) & (n_n4469) & (n_n4465) & (!x11505x)) + ((n_n4470) & (!n_n4475) & (n_n4469) & (n_n4465) & (x11505x)) + ((n_n4470) & (n_n4475) & (!n_n4469) & (!n_n4465) & (!x11505x)) + ((n_n4470) & (n_n4475) & (!n_n4469) & (!n_n4465) & (x11505x)) + ((n_n4470) & (n_n4475) & (!n_n4469) & (n_n4465) & (!x11505x)) + ((n_n4470) & (n_n4475) & (!n_n4469) & (n_n4465) & (x11505x)) + ((n_n4470) & (n_n4475) & (n_n4469) & (!n_n4465) & (!x11505x)) + ((n_n4470) & (n_n4475) & (n_n4469) & (!n_n4465) & (x11505x)) + ((n_n4470) & (n_n4475) & (n_n4469) & (n_n4465) & (!x11505x)) + ((n_n4470) & (n_n4475) & (n_n4469) & (n_n4465) & (x11505x)));
	assign x11555x = (((!n_n4637) & (!n_n4648) & (!n_n4628) & (n_n4635)) + ((!n_n4637) & (!n_n4648) & (n_n4628) & (!n_n4635)) + ((!n_n4637) & (!n_n4648) & (n_n4628) & (n_n4635)) + ((!n_n4637) & (n_n4648) & (!n_n4628) & (!n_n4635)) + ((!n_n4637) & (n_n4648) & (!n_n4628) & (n_n4635)) + ((!n_n4637) & (n_n4648) & (n_n4628) & (!n_n4635)) + ((!n_n4637) & (n_n4648) & (n_n4628) & (n_n4635)) + ((n_n4637) & (!n_n4648) & (!n_n4628) & (!n_n4635)) + ((n_n4637) & (!n_n4648) & (!n_n4628) & (n_n4635)) + ((n_n4637) & (!n_n4648) & (n_n4628) & (!n_n4635)) + ((n_n4637) & (!n_n4648) & (n_n4628) & (n_n4635)) + ((n_n4637) & (n_n4648) & (!n_n4628) & (!n_n4635)) + ((n_n4637) & (n_n4648) & (!n_n4628) & (n_n4635)) + ((n_n4637) & (n_n4648) & (n_n4628) & (!n_n4635)) + ((n_n4637) & (n_n4648) & (n_n4628) & (n_n4635)));
	assign x11556x = (((!n_n4621) & (!x309x) & (!n_n4622) & (!x75x) & (n_n4626)) + ((!n_n4621) & (!x309x) & (!n_n4622) & (x75x) & (!n_n4626)) + ((!n_n4621) & (!x309x) & (!n_n4622) & (x75x) & (n_n4626)) + ((!n_n4621) & (!x309x) & (n_n4622) & (!x75x) & (!n_n4626)) + ((!n_n4621) & (!x309x) & (n_n4622) & (!x75x) & (n_n4626)) + ((!n_n4621) & (!x309x) & (n_n4622) & (x75x) & (!n_n4626)) + ((!n_n4621) & (!x309x) & (n_n4622) & (x75x) & (n_n4626)) + ((!n_n4621) & (x309x) & (!n_n4622) & (!x75x) & (!n_n4626)) + ((!n_n4621) & (x309x) & (!n_n4622) & (!x75x) & (n_n4626)) + ((!n_n4621) & (x309x) & (!n_n4622) & (x75x) & (!n_n4626)) + ((!n_n4621) & (x309x) & (!n_n4622) & (x75x) & (n_n4626)) + ((!n_n4621) & (x309x) & (n_n4622) & (!x75x) & (!n_n4626)) + ((!n_n4621) & (x309x) & (n_n4622) & (!x75x) & (n_n4626)) + ((!n_n4621) & (x309x) & (n_n4622) & (x75x) & (!n_n4626)) + ((!n_n4621) & (x309x) & (n_n4622) & (x75x) & (n_n4626)) + ((n_n4621) & (!x309x) & (!n_n4622) & (!x75x) & (!n_n4626)) + ((n_n4621) & (!x309x) & (!n_n4622) & (!x75x) & (n_n4626)) + ((n_n4621) & (!x309x) & (!n_n4622) & (x75x) & (!n_n4626)) + ((n_n4621) & (!x309x) & (!n_n4622) & (x75x) & (n_n4626)) + ((n_n4621) & (!x309x) & (n_n4622) & (!x75x) & (!n_n4626)) + ((n_n4621) & (!x309x) & (n_n4622) & (!x75x) & (n_n4626)) + ((n_n4621) & (!x309x) & (n_n4622) & (x75x) & (!n_n4626)) + ((n_n4621) & (!x309x) & (n_n4622) & (x75x) & (n_n4626)) + ((n_n4621) & (x309x) & (!n_n4622) & (!x75x) & (!n_n4626)) + ((n_n4621) & (x309x) & (!n_n4622) & (!x75x) & (n_n4626)) + ((n_n4621) & (x309x) & (!n_n4622) & (x75x) & (!n_n4626)) + ((n_n4621) & (x309x) & (!n_n4622) & (x75x) & (n_n4626)) + ((n_n4621) & (x309x) & (n_n4622) & (!x75x) & (!n_n4626)) + ((n_n4621) & (x309x) & (n_n4622) & (!x75x) & (n_n4626)) + ((n_n4621) & (x309x) & (n_n4622) & (x75x) & (!n_n4626)) + ((n_n4621) & (x309x) & (n_n4622) & (x75x) & (n_n4626)));
	assign x11557x = (((!x348x) & (!n_n4629) & (!n_n4630) & (!x119x) & (x190x)) + ((!x348x) & (!n_n4629) & (!n_n4630) & (x119x) & (!x190x)) + ((!x348x) & (!n_n4629) & (!n_n4630) & (x119x) & (x190x)) + ((!x348x) & (!n_n4629) & (n_n4630) & (!x119x) & (!x190x)) + ((!x348x) & (!n_n4629) & (n_n4630) & (!x119x) & (x190x)) + ((!x348x) & (!n_n4629) & (n_n4630) & (x119x) & (!x190x)) + ((!x348x) & (!n_n4629) & (n_n4630) & (x119x) & (x190x)) + ((!x348x) & (n_n4629) & (!n_n4630) & (!x119x) & (!x190x)) + ((!x348x) & (n_n4629) & (!n_n4630) & (!x119x) & (x190x)) + ((!x348x) & (n_n4629) & (!n_n4630) & (x119x) & (!x190x)) + ((!x348x) & (n_n4629) & (!n_n4630) & (x119x) & (x190x)) + ((!x348x) & (n_n4629) & (n_n4630) & (!x119x) & (!x190x)) + ((!x348x) & (n_n4629) & (n_n4630) & (!x119x) & (x190x)) + ((!x348x) & (n_n4629) & (n_n4630) & (x119x) & (!x190x)) + ((!x348x) & (n_n4629) & (n_n4630) & (x119x) & (x190x)) + ((x348x) & (!n_n4629) & (!n_n4630) & (!x119x) & (!x190x)) + ((x348x) & (!n_n4629) & (!n_n4630) & (!x119x) & (x190x)) + ((x348x) & (!n_n4629) & (!n_n4630) & (x119x) & (!x190x)) + ((x348x) & (!n_n4629) & (!n_n4630) & (x119x) & (x190x)) + ((x348x) & (!n_n4629) & (n_n4630) & (!x119x) & (!x190x)) + ((x348x) & (!n_n4629) & (n_n4630) & (!x119x) & (x190x)) + ((x348x) & (!n_n4629) & (n_n4630) & (x119x) & (!x190x)) + ((x348x) & (!n_n4629) & (n_n4630) & (x119x) & (x190x)) + ((x348x) & (n_n4629) & (!n_n4630) & (!x119x) & (!x190x)) + ((x348x) & (n_n4629) & (!n_n4630) & (!x119x) & (x190x)) + ((x348x) & (n_n4629) & (!n_n4630) & (x119x) & (!x190x)) + ((x348x) & (n_n4629) & (!n_n4630) & (x119x) & (x190x)) + ((x348x) & (n_n4629) & (n_n4630) & (!x119x) & (!x190x)) + ((x348x) & (n_n4629) & (n_n4630) & (!x119x) & (x190x)) + ((x348x) & (n_n4629) & (n_n4630) & (x119x) & (!x190x)) + ((x348x) & (n_n4629) & (n_n4630) & (x119x) & (x190x)));
	assign x11572x = (((!n_n4591) & (!n_n4592) & (!n_n4579) & (n_n4583)) + ((!n_n4591) & (!n_n4592) & (n_n4579) & (!n_n4583)) + ((!n_n4591) & (!n_n4592) & (n_n4579) & (n_n4583)) + ((!n_n4591) & (n_n4592) & (!n_n4579) & (!n_n4583)) + ((!n_n4591) & (n_n4592) & (!n_n4579) & (n_n4583)) + ((!n_n4591) & (n_n4592) & (n_n4579) & (!n_n4583)) + ((!n_n4591) & (n_n4592) & (n_n4579) & (n_n4583)) + ((n_n4591) & (!n_n4592) & (!n_n4579) & (!n_n4583)) + ((n_n4591) & (!n_n4592) & (!n_n4579) & (n_n4583)) + ((n_n4591) & (!n_n4592) & (n_n4579) & (!n_n4583)) + ((n_n4591) & (!n_n4592) & (n_n4579) & (n_n4583)) + ((n_n4591) & (n_n4592) & (!n_n4579) & (!n_n4583)) + ((n_n4591) & (n_n4592) & (!n_n4579) & (n_n4583)) + ((n_n4591) & (n_n4592) & (n_n4579) & (!n_n4583)) + ((n_n4591) & (n_n4592) & (n_n4579) & (n_n4583)));
	assign x11573x = (((!n_n4593) & (!n_n4594) & (!x365x) & (x11571x)) + ((!n_n4593) & (!n_n4594) & (x365x) & (!x11571x)) + ((!n_n4593) & (!n_n4594) & (x365x) & (x11571x)) + ((!n_n4593) & (n_n4594) & (!x365x) & (!x11571x)) + ((!n_n4593) & (n_n4594) & (!x365x) & (x11571x)) + ((!n_n4593) & (n_n4594) & (x365x) & (!x11571x)) + ((!n_n4593) & (n_n4594) & (x365x) & (x11571x)) + ((n_n4593) & (!n_n4594) & (!x365x) & (!x11571x)) + ((n_n4593) & (!n_n4594) & (!x365x) & (x11571x)) + ((n_n4593) & (!n_n4594) & (x365x) & (!x11571x)) + ((n_n4593) & (!n_n4594) & (x365x) & (x11571x)) + ((n_n4593) & (n_n4594) & (!x365x) & (!x11571x)) + ((n_n4593) & (n_n4594) & (!x365x) & (x11571x)) + ((n_n4593) & (n_n4594) & (x365x) & (!x11571x)) + ((n_n4593) & (n_n4594) & (x365x) & (x11571x)));
	assign x284x = (((!i_9_) & (n_n536) & (!n_n532) & (n_n534) & (n_n535)) + ((!i_9_) & (n_n536) & (n_n532) & (n_n534) & (n_n535)) + ((i_9_) & (n_n536) & (!n_n532) & (n_n534) & (n_n535)) + ((i_9_) & (n_n536) & (n_n532) & (!n_n534) & (n_n535)) + ((i_9_) & (n_n536) & (n_n532) & (n_n534) & (n_n535)));
	assign x11587x = (((!n_n536) & (!x24x) & (!n_n535) & (!n_n4321) & (x284x)) + ((!n_n536) & (!x24x) & (!n_n535) & (n_n4321) & (!x284x)) + ((!n_n536) & (!x24x) & (!n_n535) & (n_n4321) & (x284x)) + ((!n_n536) & (!x24x) & (n_n535) & (!n_n4321) & (x284x)) + ((!n_n536) & (!x24x) & (n_n535) & (n_n4321) & (!x284x)) + ((!n_n536) & (!x24x) & (n_n535) & (n_n4321) & (x284x)) + ((!n_n536) & (x24x) & (!n_n535) & (!n_n4321) & (x284x)) + ((!n_n536) & (x24x) & (!n_n535) & (n_n4321) & (!x284x)) + ((!n_n536) & (x24x) & (!n_n535) & (n_n4321) & (x284x)) + ((!n_n536) & (x24x) & (n_n535) & (!n_n4321) & (x284x)) + ((!n_n536) & (x24x) & (n_n535) & (n_n4321) & (!x284x)) + ((!n_n536) & (x24x) & (n_n535) & (n_n4321) & (x284x)) + ((n_n536) & (!x24x) & (!n_n535) & (!n_n4321) & (x284x)) + ((n_n536) & (!x24x) & (!n_n535) & (n_n4321) & (!x284x)) + ((n_n536) & (!x24x) & (!n_n535) & (n_n4321) & (x284x)) + ((n_n536) & (!x24x) & (n_n535) & (!n_n4321) & (x284x)) + ((n_n536) & (!x24x) & (n_n535) & (n_n4321) & (!x284x)) + ((n_n536) & (!x24x) & (n_n535) & (n_n4321) & (x284x)) + ((n_n536) & (x24x) & (!n_n535) & (!n_n4321) & (x284x)) + ((n_n536) & (x24x) & (!n_n535) & (n_n4321) & (!x284x)) + ((n_n536) & (x24x) & (!n_n535) & (n_n4321) & (x284x)) + ((n_n536) & (x24x) & (n_n535) & (!n_n4321) & (!x284x)) + ((n_n536) & (x24x) & (n_n535) & (!n_n4321) & (x284x)) + ((n_n536) & (x24x) & (n_n535) & (n_n4321) & (!x284x)) + ((n_n536) & (x24x) & (n_n535) & (n_n4321) & (x284x)));
	assign x11603x = (((!n_n4401) & (!n_n4393) & (!n_n4391) & (!n_n4397) & (n_n4402)) + ((!n_n4401) & (!n_n4393) & (!n_n4391) & (n_n4397) & (!n_n4402)) + ((!n_n4401) & (!n_n4393) & (!n_n4391) & (n_n4397) & (n_n4402)) + ((!n_n4401) & (!n_n4393) & (n_n4391) & (!n_n4397) & (!n_n4402)) + ((!n_n4401) & (!n_n4393) & (n_n4391) & (!n_n4397) & (n_n4402)) + ((!n_n4401) & (!n_n4393) & (n_n4391) & (n_n4397) & (!n_n4402)) + ((!n_n4401) & (!n_n4393) & (n_n4391) & (n_n4397) & (n_n4402)) + ((!n_n4401) & (n_n4393) & (!n_n4391) & (!n_n4397) & (!n_n4402)) + ((!n_n4401) & (n_n4393) & (!n_n4391) & (!n_n4397) & (n_n4402)) + ((!n_n4401) & (n_n4393) & (!n_n4391) & (n_n4397) & (!n_n4402)) + ((!n_n4401) & (n_n4393) & (!n_n4391) & (n_n4397) & (n_n4402)) + ((!n_n4401) & (n_n4393) & (n_n4391) & (!n_n4397) & (!n_n4402)) + ((!n_n4401) & (n_n4393) & (n_n4391) & (!n_n4397) & (n_n4402)) + ((!n_n4401) & (n_n4393) & (n_n4391) & (n_n4397) & (!n_n4402)) + ((!n_n4401) & (n_n4393) & (n_n4391) & (n_n4397) & (n_n4402)) + ((n_n4401) & (!n_n4393) & (!n_n4391) & (!n_n4397) & (!n_n4402)) + ((n_n4401) & (!n_n4393) & (!n_n4391) & (!n_n4397) & (n_n4402)) + ((n_n4401) & (!n_n4393) & (!n_n4391) & (n_n4397) & (!n_n4402)) + ((n_n4401) & (!n_n4393) & (!n_n4391) & (n_n4397) & (n_n4402)) + ((n_n4401) & (!n_n4393) & (n_n4391) & (!n_n4397) & (!n_n4402)) + ((n_n4401) & (!n_n4393) & (n_n4391) & (!n_n4397) & (n_n4402)) + ((n_n4401) & (!n_n4393) & (n_n4391) & (n_n4397) & (!n_n4402)) + ((n_n4401) & (!n_n4393) & (n_n4391) & (n_n4397) & (n_n4402)) + ((n_n4401) & (n_n4393) & (!n_n4391) & (!n_n4397) & (!n_n4402)) + ((n_n4401) & (n_n4393) & (!n_n4391) & (!n_n4397) & (n_n4402)) + ((n_n4401) & (n_n4393) & (!n_n4391) & (n_n4397) & (!n_n4402)) + ((n_n4401) & (n_n4393) & (!n_n4391) & (n_n4397) & (n_n4402)) + ((n_n4401) & (n_n4393) & (n_n4391) & (!n_n4397) & (!n_n4402)) + ((n_n4401) & (n_n4393) & (n_n4391) & (!n_n4397) & (n_n4402)) + ((n_n4401) & (n_n4393) & (n_n4391) & (n_n4397) & (!n_n4402)) + ((n_n4401) & (n_n4393) & (n_n4391) & (n_n4397) & (n_n4402)));
	assign x11604x = (((!n_n4400) & (!n_n4392) & (!n_n4396) & (!n_n4399) & (x11603x)) + ((!n_n4400) & (!n_n4392) & (!n_n4396) & (n_n4399) & (!x11603x)) + ((!n_n4400) & (!n_n4392) & (!n_n4396) & (n_n4399) & (x11603x)) + ((!n_n4400) & (!n_n4392) & (n_n4396) & (!n_n4399) & (!x11603x)) + ((!n_n4400) & (!n_n4392) & (n_n4396) & (!n_n4399) & (x11603x)) + ((!n_n4400) & (!n_n4392) & (n_n4396) & (n_n4399) & (!x11603x)) + ((!n_n4400) & (!n_n4392) & (n_n4396) & (n_n4399) & (x11603x)) + ((!n_n4400) & (n_n4392) & (!n_n4396) & (!n_n4399) & (!x11603x)) + ((!n_n4400) & (n_n4392) & (!n_n4396) & (!n_n4399) & (x11603x)) + ((!n_n4400) & (n_n4392) & (!n_n4396) & (n_n4399) & (!x11603x)) + ((!n_n4400) & (n_n4392) & (!n_n4396) & (n_n4399) & (x11603x)) + ((!n_n4400) & (n_n4392) & (n_n4396) & (!n_n4399) & (!x11603x)) + ((!n_n4400) & (n_n4392) & (n_n4396) & (!n_n4399) & (x11603x)) + ((!n_n4400) & (n_n4392) & (n_n4396) & (n_n4399) & (!x11603x)) + ((!n_n4400) & (n_n4392) & (n_n4396) & (n_n4399) & (x11603x)) + ((n_n4400) & (!n_n4392) & (!n_n4396) & (!n_n4399) & (!x11603x)) + ((n_n4400) & (!n_n4392) & (!n_n4396) & (!n_n4399) & (x11603x)) + ((n_n4400) & (!n_n4392) & (!n_n4396) & (n_n4399) & (!x11603x)) + ((n_n4400) & (!n_n4392) & (!n_n4396) & (n_n4399) & (x11603x)) + ((n_n4400) & (!n_n4392) & (n_n4396) & (!n_n4399) & (!x11603x)) + ((n_n4400) & (!n_n4392) & (n_n4396) & (!n_n4399) & (x11603x)) + ((n_n4400) & (!n_n4392) & (n_n4396) & (n_n4399) & (!x11603x)) + ((n_n4400) & (!n_n4392) & (n_n4396) & (n_n4399) & (x11603x)) + ((n_n4400) & (n_n4392) & (!n_n4396) & (!n_n4399) & (!x11603x)) + ((n_n4400) & (n_n4392) & (!n_n4396) & (!n_n4399) & (x11603x)) + ((n_n4400) & (n_n4392) & (!n_n4396) & (n_n4399) & (!x11603x)) + ((n_n4400) & (n_n4392) & (!n_n4396) & (n_n4399) & (x11603x)) + ((n_n4400) & (n_n4392) & (n_n4396) & (!n_n4399) & (!x11603x)) + ((n_n4400) & (n_n4392) & (n_n4396) & (!n_n4399) & (x11603x)) + ((n_n4400) & (n_n4392) & (n_n4396) & (n_n4399) & (!x11603x)) + ((n_n4400) & (n_n4392) & (n_n4396) & (n_n4399) & (x11603x)));
	assign x11618x = (((!n_n3533) & (!n_n1308) & (!n_n4360) & (!x282x) & (n_n4375)) + ((!n_n3533) & (!n_n1308) & (!n_n4360) & (x282x) & (!n_n4375)) + ((!n_n3533) & (!n_n1308) & (!n_n4360) & (x282x) & (n_n4375)) + ((!n_n3533) & (!n_n1308) & (n_n4360) & (!x282x) & (!n_n4375)) + ((!n_n3533) & (!n_n1308) & (n_n4360) & (!x282x) & (n_n4375)) + ((!n_n3533) & (!n_n1308) & (n_n4360) & (x282x) & (!n_n4375)) + ((!n_n3533) & (!n_n1308) & (n_n4360) & (x282x) & (n_n4375)) + ((!n_n3533) & (n_n1308) & (!n_n4360) & (!x282x) & (!n_n4375)) + ((!n_n3533) & (n_n1308) & (!n_n4360) & (!x282x) & (n_n4375)) + ((!n_n3533) & (n_n1308) & (!n_n4360) & (x282x) & (!n_n4375)) + ((!n_n3533) & (n_n1308) & (!n_n4360) & (x282x) & (n_n4375)) + ((!n_n3533) & (n_n1308) & (n_n4360) & (!x282x) & (!n_n4375)) + ((!n_n3533) & (n_n1308) & (n_n4360) & (!x282x) & (n_n4375)) + ((!n_n3533) & (n_n1308) & (n_n4360) & (x282x) & (!n_n4375)) + ((!n_n3533) & (n_n1308) & (n_n4360) & (x282x) & (n_n4375)) + ((n_n3533) & (!n_n1308) & (!n_n4360) & (!x282x) & (!n_n4375)) + ((n_n3533) & (!n_n1308) & (!n_n4360) & (!x282x) & (n_n4375)) + ((n_n3533) & (!n_n1308) & (!n_n4360) & (x282x) & (!n_n4375)) + ((n_n3533) & (!n_n1308) & (!n_n4360) & (x282x) & (n_n4375)) + ((n_n3533) & (!n_n1308) & (n_n4360) & (!x282x) & (!n_n4375)) + ((n_n3533) & (!n_n1308) & (n_n4360) & (!x282x) & (n_n4375)) + ((n_n3533) & (!n_n1308) & (n_n4360) & (x282x) & (!n_n4375)) + ((n_n3533) & (!n_n1308) & (n_n4360) & (x282x) & (n_n4375)) + ((n_n3533) & (n_n1308) & (!n_n4360) & (!x282x) & (!n_n4375)) + ((n_n3533) & (n_n1308) & (!n_n4360) & (!x282x) & (n_n4375)) + ((n_n3533) & (n_n1308) & (!n_n4360) & (x282x) & (!n_n4375)) + ((n_n3533) & (n_n1308) & (!n_n4360) & (x282x) & (n_n4375)) + ((n_n3533) & (n_n1308) & (n_n4360) & (!x282x) & (!n_n4375)) + ((n_n3533) & (n_n1308) & (n_n4360) & (!x282x) & (n_n4375)) + ((n_n3533) & (n_n1308) & (n_n4360) & (x282x) & (!n_n4375)) + ((n_n3533) & (n_n1308) & (n_n4360) & (x282x) & (n_n4375)));
	assign x161x = (((!i_9_) & (!n_n536) & (!n_n534) & (!n_n500) & (n_n4359)) + ((!i_9_) & (!n_n536) & (!n_n534) & (n_n500) & (n_n4359)) + ((!i_9_) & (!n_n536) & (n_n534) & (!n_n500) & (n_n4359)) + ((!i_9_) & (!n_n536) & (n_n534) & (n_n500) & (n_n4359)) + ((!i_9_) & (n_n536) & (!n_n534) & (!n_n500) & (n_n4359)) + ((!i_9_) & (n_n536) & (!n_n534) & (n_n500) & (n_n4359)) + ((!i_9_) & (n_n536) & (n_n534) & (!n_n500) & (n_n4359)) + ((!i_9_) & (n_n536) & (n_n534) & (n_n500) & (!n_n4359)) + ((!i_9_) & (n_n536) & (n_n534) & (n_n500) & (n_n4359)) + ((i_9_) & (!n_n536) & (!n_n534) & (!n_n500) & (n_n4359)) + ((i_9_) & (!n_n536) & (!n_n534) & (n_n500) & (n_n4359)) + ((i_9_) & (!n_n536) & (n_n534) & (!n_n500) & (n_n4359)) + ((i_9_) & (!n_n536) & (n_n534) & (n_n500) & (n_n4359)) + ((i_9_) & (n_n536) & (!n_n534) & (!n_n500) & (n_n4359)) + ((i_9_) & (n_n536) & (!n_n534) & (n_n500) & (n_n4359)) + ((i_9_) & (n_n536) & (n_n534) & (!n_n500) & (n_n4359)) + ((i_9_) & (n_n536) & (n_n534) & (n_n500) & (n_n4359)));
	assign x11620x = (((!i_9_) & (n_n536) & (n_n524) & (n_n518)) + ((i_9_) & (n_n536) & (n_n524) & (n_n518)));
	assign x22150x = (((!n_n4345) & (!n_n4343) & (!n_n4341) & (!n_n4342)));
	assign x12640x = (((!n_n5183) & (!n_n5204) & (!n_n5182) & (n_n5173)) + ((!n_n5183) & (!n_n5204) & (n_n5182) & (!n_n5173)) + ((!n_n5183) & (!n_n5204) & (n_n5182) & (n_n5173)) + ((!n_n5183) & (n_n5204) & (!n_n5182) & (!n_n5173)) + ((!n_n5183) & (n_n5204) & (!n_n5182) & (n_n5173)) + ((!n_n5183) & (n_n5204) & (n_n5182) & (!n_n5173)) + ((!n_n5183) & (n_n5204) & (n_n5182) & (n_n5173)) + ((n_n5183) & (!n_n5204) & (!n_n5182) & (!n_n5173)) + ((n_n5183) & (!n_n5204) & (!n_n5182) & (n_n5173)) + ((n_n5183) & (!n_n5204) & (n_n5182) & (!n_n5173)) + ((n_n5183) & (!n_n5204) & (n_n5182) & (n_n5173)) + ((n_n5183) & (n_n5204) & (!n_n5182) & (!n_n5173)) + ((n_n5183) & (n_n5204) & (!n_n5182) & (n_n5173)) + ((n_n5183) & (n_n5204) & (n_n5182) & (!n_n5173)) + ((n_n5183) & (n_n5204) & (n_n5182) & (n_n5173)));
	assign x12641x = (((!n_n5179) & (!n_n5178) & (!n_n5166) & (!n_n5168) & (n_n5211)) + ((!n_n5179) & (!n_n5178) & (!n_n5166) & (n_n5168) & (!n_n5211)) + ((!n_n5179) & (!n_n5178) & (!n_n5166) & (n_n5168) & (n_n5211)) + ((!n_n5179) & (!n_n5178) & (n_n5166) & (!n_n5168) & (!n_n5211)) + ((!n_n5179) & (!n_n5178) & (n_n5166) & (!n_n5168) & (n_n5211)) + ((!n_n5179) & (!n_n5178) & (n_n5166) & (n_n5168) & (!n_n5211)) + ((!n_n5179) & (!n_n5178) & (n_n5166) & (n_n5168) & (n_n5211)) + ((!n_n5179) & (n_n5178) & (!n_n5166) & (!n_n5168) & (!n_n5211)) + ((!n_n5179) & (n_n5178) & (!n_n5166) & (!n_n5168) & (n_n5211)) + ((!n_n5179) & (n_n5178) & (!n_n5166) & (n_n5168) & (!n_n5211)) + ((!n_n5179) & (n_n5178) & (!n_n5166) & (n_n5168) & (n_n5211)) + ((!n_n5179) & (n_n5178) & (n_n5166) & (!n_n5168) & (!n_n5211)) + ((!n_n5179) & (n_n5178) & (n_n5166) & (!n_n5168) & (n_n5211)) + ((!n_n5179) & (n_n5178) & (n_n5166) & (n_n5168) & (!n_n5211)) + ((!n_n5179) & (n_n5178) & (n_n5166) & (n_n5168) & (n_n5211)) + ((n_n5179) & (!n_n5178) & (!n_n5166) & (!n_n5168) & (!n_n5211)) + ((n_n5179) & (!n_n5178) & (!n_n5166) & (!n_n5168) & (n_n5211)) + ((n_n5179) & (!n_n5178) & (!n_n5166) & (n_n5168) & (!n_n5211)) + ((n_n5179) & (!n_n5178) & (!n_n5166) & (n_n5168) & (n_n5211)) + ((n_n5179) & (!n_n5178) & (n_n5166) & (!n_n5168) & (!n_n5211)) + ((n_n5179) & (!n_n5178) & (n_n5166) & (!n_n5168) & (n_n5211)) + ((n_n5179) & (!n_n5178) & (n_n5166) & (n_n5168) & (!n_n5211)) + ((n_n5179) & (!n_n5178) & (n_n5166) & (n_n5168) & (n_n5211)) + ((n_n5179) & (n_n5178) & (!n_n5166) & (!n_n5168) & (!n_n5211)) + ((n_n5179) & (n_n5178) & (!n_n5166) & (!n_n5168) & (n_n5211)) + ((n_n5179) & (n_n5178) & (!n_n5166) & (n_n5168) & (!n_n5211)) + ((n_n5179) & (n_n5178) & (!n_n5166) & (n_n5168) & (n_n5211)) + ((n_n5179) & (n_n5178) & (n_n5166) & (!n_n5168) & (!n_n5211)) + ((n_n5179) & (n_n5178) & (n_n5166) & (!n_n5168) & (n_n5211)) + ((n_n5179) & (n_n5178) & (n_n5166) & (n_n5168) & (!n_n5211)) + ((n_n5179) & (n_n5178) & (n_n5166) & (n_n5168) & (n_n5211)));
	assign x312x = (((!i_9_) & (!n_n524) & (n_n482) & (n_n390) & (n_n530)) + ((!i_9_) & (n_n524) & (n_n482) & (n_n390) & (n_n530)) + ((i_9_) & (n_n524) & (n_n482) & (n_n390) & (!n_n530)) + ((i_9_) & (n_n524) & (n_n482) & (n_n390) & (n_n530)));
	assign x22126x = (((!n_n4666) & (!n_n4667) & (!n_n4664) & (!n_n4662)));
	assign x330x = (((!i_9_) & (n_n528) & (n_n260) & (n_n500)) + ((i_9_) & (n_n528) & (n_n260) & (n_n500)));
	assign n_n1988 = (((!i_9_) & (!n_n524) & (n_n509) & (n_n260) & (x20x)) + ((!i_9_) & (n_n524) & (n_n509) & (n_n260) & (!x20x)) + ((!i_9_) & (n_n524) & (n_n509) & (n_n260) & (x20x)) + ((i_9_) & (!n_n524) & (n_n509) & (n_n260) & (x20x)) + ((i_9_) & (n_n524) & (n_n509) & (n_n260) & (!x20x)) + ((i_9_) & (n_n524) & (n_n509) & (n_n260) & (x20x)));
	assign x162x = (((!i_9_) & (n_n455) & (!n_n520) & (x20x) & (n_n500)) + ((!i_9_) & (n_n455) & (n_n520) & (x20x) & (n_n500)) + ((i_9_) & (n_n455) & (!n_n520) & (x20x) & (n_n500)) + ((i_9_) & (n_n455) & (n_n520) & (!x20x) & (n_n500)) + ((i_9_) & (n_n455) & (n_n520) & (x20x) & (n_n500)));
	assign n_n897 = (((!i_9_) & (!n_n524) & (n_n526) & (n_n455) & (n_n500)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n455) & (n_n500)) + ((i_9_) & (!n_n524) & (n_n526) & (n_n455) & (n_n500)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n455) & (n_n500)) + ((i_9_) & (n_n524) & (n_n526) & (n_n455) & (n_n500)));
	assign n_n3355 = (((!x66x) & (!n_n4500) & (!n_n4493) & (!x162x) & (n_n897)) + ((!x66x) & (!n_n4500) & (!n_n4493) & (x162x) & (!n_n897)) + ((!x66x) & (!n_n4500) & (!n_n4493) & (x162x) & (n_n897)) + ((!x66x) & (!n_n4500) & (n_n4493) & (!x162x) & (!n_n897)) + ((!x66x) & (!n_n4500) & (n_n4493) & (!x162x) & (n_n897)) + ((!x66x) & (!n_n4500) & (n_n4493) & (x162x) & (!n_n897)) + ((!x66x) & (!n_n4500) & (n_n4493) & (x162x) & (n_n897)) + ((!x66x) & (n_n4500) & (!n_n4493) & (!x162x) & (!n_n897)) + ((!x66x) & (n_n4500) & (!n_n4493) & (!x162x) & (n_n897)) + ((!x66x) & (n_n4500) & (!n_n4493) & (x162x) & (!n_n897)) + ((!x66x) & (n_n4500) & (!n_n4493) & (x162x) & (n_n897)) + ((!x66x) & (n_n4500) & (n_n4493) & (!x162x) & (!n_n897)) + ((!x66x) & (n_n4500) & (n_n4493) & (!x162x) & (n_n897)) + ((!x66x) & (n_n4500) & (n_n4493) & (x162x) & (!n_n897)) + ((!x66x) & (n_n4500) & (n_n4493) & (x162x) & (n_n897)) + ((x66x) & (!n_n4500) & (!n_n4493) & (!x162x) & (!n_n897)) + ((x66x) & (!n_n4500) & (!n_n4493) & (!x162x) & (n_n897)) + ((x66x) & (!n_n4500) & (!n_n4493) & (x162x) & (!n_n897)) + ((x66x) & (!n_n4500) & (!n_n4493) & (x162x) & (n_n897)) + ((x66x) & (!n_n4500) & (n_n4493) & (!x162x) & (!n_n897)) + ((x66x) & (!n_n4500) & (n_n4493) & (!x162x) & (n_n897)) + ((x66x) & (!n_n4500) & (n_n4493) & (x162x) & (!n_n897)) + ((x66x) & (!n_n4500) & (n_n4493) & (x162x) & (n_n897)) + ((x66x) & (n_n4500) & (!n_n4493) & (!x162x) & (!n_n897)) + ((x66x) & (n_n4500) & (!n_n4493) & (!x162x) & (n_n897)) + ((x66x) & (n_n4500) & (!n_n4493) & (x162x) & (!n_n897)) + ((x66x) & (n_n4500) & (!n_n4493) & (x162x) & (n_n897)) + ((x66x) & (n_n4500) & (n_n4493) & (!x162x) & (!n_n897)) + ((x66x) & (n_n4500) & (n_n4493) & (!x162x) & (n_n897)) + ((x66x) & (n_n4500) & (n_n4493) & (x162x) & (!n_n897)) + ((x66x) & (n_n4500) & (n_n4493) & (x162x) & (n_n897)));
	assign n_n3354 = (((!n_n4511) & (!n_n4503) & (!x189x) & (!x129x) & (n_n3509)) + ((!n_n4511) & (!n_n4503) & (!x189x) & (x129x) & (!n_n3509)) + ((!n_n4511) & (!n_n4503) & (!x189x) & (x129x) & (n_n3509)) + ((!n_n4511) & (!n_n4503) & (x189x) & (!x129x) & (!n_n3509)) + ((!n_n4511) & (!n_n4503) & (x189x) & (!x129x) & (n_n3509)) + ((!n_n4511) & (!n_n4503) & (x189x) & (x129x) & (!n_n3509)) + ((!n_n4511) & (!n_n4503) & (x189x) & (x129x) & (n_n3509)) + ((!n_n4511) & (n_n4503) & (!x189x) & (!x129x) & (!n_n3509)) + ((!n_n4511) & (n_n4503) & (!x189x) & (!x129x) & (n_n3509)) + ((!n_n4511) & (n_n4503) & (!x189x) & (x129x) & (!n_n3509)) + ((!n_n4511) & (n_n4503) & (!x189x) & (x129x) & (n_n3509)) + ((!n_n4511) & (n_n4503) & (x189x) & (!x129x) & (!n_n3509)) + ((!n_n4511) & (n_n4503) & (x189x) & (!x129x) & (n_n3509)) + ((!n_n4511) & (n_n4503) & (x189x) & (x129x) & (!n_n3509)) + ((!n_n4511) & (n_n4503) & (x189x) & (x129x) & (n_n3509)) + ((n_n4511) & (!n_n4503) & (!x189x) & (!x129x) & (!n_n3509)) + ((n_n4511) & (!n_n4503) & (!x189x) & (!x129x) & (n_n3509)) + ((n_n4511) & (!n_n4503) & (!x189x) & (x129x) & (!n_n3509)) + ((n_n4511) & (!n_n4503) & (!x189x) & (x129x) & (n_n3509)) + ((n_n4511) & (!n_n4503) & (x189x) & (!x129x) & (!n_n3509)) + ((n_n4511) & (!n_n4503) & (x189x) & (!x129x) & (n_n3509)) + ((n_n4511) & (!n_n4503) & (x189x) & (x129x) & (!n_n3509)) + ((n_n4511) & (!n_n4503) & (x189x) & (x129x) & (n_n3509)) + ((n_n4511) & (n_n4503) & (!x189x) & (!x129x) & (!n_n3509)) + ((n_n4511) & (n_n4503) & (!x189x) & (!x129x) & (n_n3509)) + ((n_n4511) & (n_n4503) & (!x189x) & (x129x) & (!n_n3509)) + ((n_n4511) & (n_n4503) & (!x189x) & (x129x) & (n_n3509)) + ((n_n4511) & (n_n4503) & (x189x) & (!x129x) & (!n_n3509)) + ((n_n4511) & (n_n4503) & (x189x) & (!x129x) & (n_n3509)) + ((n_n4511) & (n_n4503) & (x189x) & (x129x) & (!n_n3509)) + ((n_n4511) & (n_n4503) & (x189x) & (x129x) & (n_n3509)));
	assign x14207x = (((!n_n4247) & (!n_n4521) & (!n_n4246) & (!n_n4517) & (n_n4520)) + ((!n_n4247) & (!n_n4521) & (!n_n4246) & (n_n4517) & (!n_n4520)) + ((!n_n4247) & (!n_n4521) & (!n_n4246) & (n_n4517) & (n_n4520)) + ((!n_n4247) & (!n_n4521) & (n_n4246) & (!n_n4517) & (!n_n4520)) + ((!n_n4247) & (!n_n4521) & (n_n4246) & (!n_n4517) & (n_n4520)) + ((!n_n4247) & (!n_n4521) & (n_n4246) & (n_n4517) & (!n_n4520)) + ((!n_n4247) & (!n_n4521) & (n_n4246) & (n_n4517) & (n_n4520)) + ((!n_n4247) & (n_n4521) & (!n_n4246) & (!n_n4517) & (!n_n4520)) + ((!n_n4247) & (n_n4521) & (!n_n4246) & (!n_n4517) & (n_n4520)) + ((!n_n4247) & (n_n4521) & (!n_n4246) & (n_n4517) & (!n_n4520)) + ((!n_n4247) & (n_n4521) & (!n_n4246) & (n_n4517) & (n_n4520)) + ((!n_n4247) & (n_n4521) & (n_n4246) & (!n_n4517) & (!n_n4520)) + ((!n_n4247) & (n_n4521) & (n_n4246) & (!n_n4517) & (n_n4520)) + ((!n_n4247) & (n_n4521) & (n_n4246) & (n_n4517) & (!n_n4520)) + ((!n_n4247) & (n_n4521) & (n_n4246) & (n_n4517) & (n_n4520)) + ((n_n4247) & (!n_n4521) & (!n_n4246) & (!n_n4517) & (!n_n4520)) + ((n_n4247) & (!n_n4521) & (!n_n4246) & (!n_n4517) & (n_n4520)) + ((n_n4247) & (!n_n4521) & (!n_n4246) & (n_n4517) & (!n_n4520)) + ((n_n4247) & (!n_n4521) & (!n_n4246) & (n_n4517) & (n_n4520)) + ((n_n4247) & (!n_n4521) & (n_n4246) & (!n_n4517) & (!n_n4520)) + ((n_n4247) & (!n_n4521) & (n_n4246) & (!n_n4517) & (n_n4520)) + ((n_n4247) & (!n_n4521) & (n_n4246) & (n_n4517) & (!n_n4520)) + ((n_n4247) & (!n_n4521) & (n_n4246) & (n_n4517) & (n_n4520)) + ((n_n4247) & (n_n4521) & (!n_n4246) & (!n_n4517) & (!n_n4520)) + ((n_n4247) & (n_n4521) & (!n_n4246) & (!n_n4517) & (n_n4520)) + ((n_n4247) & (n_n4521) & (!n_n4246) & (n_n4517) & (!n_n4520)) + ((n_n4247) & (n_n4521) & (!n_n4246) & (n_n4517) & (n_n4520)) + ((n_n4247) & (n_n4521) & (n_n4246) & (!n_n4517) & (!n_n4520)) + ((n_n4247) & (n_n4521) & (n_n4246) & (!n_n4517) & (n_n4520)) + ((n_n4247) & (n_n4521) & (n_n4246) & (n_n4517) & (!n_n4520)) + ((n_n4247) & (n_n4521) & (n_n4246) & (n_n4517) & (n_n4520)));
	assign x14211x = (((!n_n3285) & (!n_n3286) & (!n_n3355) & (!n_n3354) & (x14207x)) + ((!n_n3285) & (!n_n3286) & (!n_n3355) & (n_n3354) & (!x14207x)) + ((!n_n3285) & (!n_n3286) & (!n_n3355) & (n_n3354) & (x14207x)) + ((!n_n3285) & (!n_n3286) & (n_n3355) & (!n_n3354) & (!x14207x)) + ((!n_n3285) & (!n_n3286) & (n_n3355) & (!n_n3354) & (x14207x)) + ((!n_n3285) & (!n_n3286) & (n_n3355) & (n_n3354) & (!x14207x)) + ((!n_n3285) & (!n_n3286) & (n_n3355) & (n_n3354) & (x14207x)) + ((!n_n3285) & (n_n3286) & (!n_n3355) & (!n_n3354) & (!x14207x)) + ((!n_n3285) & (n_n3286) & (!n_n3355) & (!n_n3354) & (x14207x)) + ((!n_n3285) & (n_n3286) & (!n_n3355) & (n_n3354) & (!x14207x)) + ((!n_n3285) & (n_n3286) & (!n_n3355) & (n_n3354) & (x14207x)) + ((!n_n3285) & (n_n3286) & (n_n3355) & (!n_n3354) & (!x14207x)) + ((!n_n3285) & (n_n3286) & (n_n3355) & (!n_n3354) & (x14207x)) + ((!n_n3285) & (n_n3286) & (n_n3355) & (n_n3354) & (!x14207x)) + ((!n_n3285) & (n_n3286) & (n_n3355) & (n_n3354) & (x14207x)) + ((n_n3285) & (!n_n3286) & (!n_n3355) & (!n_n3354) & (!x14207x)) + ((n_n3285) & (!n_n3286) & (!n_n3355) & (!n_n3354) & (x14207x)) + ((n_n3285) & (!n_n3286) & (!n_n3355) & (n_n3354) & (!x14207x)) + ((n_n3285) & (!n_n3286) & (!n_n3355) & (n_n3354) & (x14207x)) + ((n_n3285) & (!n_n3286) & (n_n3355) & (!n_n3354) & (!x14207x)) + ((n_n3285) & (!n_n3286) & (n_n3355) & (!n_n3354) & (x14207x)) + ((n_n3285) & (!n_n3286) & (n_n3355) & (n_n3354) & (!x14207x)) + ((n_n3285) & (!n_n3286) & (n_n3355) & (n_n3354) & (x14207x)) + ((n_n3285) & (n_n3286) & (!n_n3355) & (!n_n3354) & (!x14207x)) + ((n_n3285) & (n_n3286) & (!n_n3355) & (!n_n3354) & (x14207x)) + ((n_n3285) & (n_n3286) & (!n_n3355) & (n_n3354) & (!x14207x)) + ((n_n3285) & (n_n3286) & (!n_n3355) & (n_n3354) & (x14207x)) + ((n_n3285) & (n_n3286) & (n_n3355) & (!n_n3354) & (!x14207x)) + ((n_n3285) & (n_n3286) & (n_n3355) & (!n_n3354) & (x14207x)) + ((n_n3285) & (n_n3286) & (n_n3355) & (n_n3354) & (!x14207x)) + ((n_n3285) & (n_n3286) & (n_n3355) & (n_n3354) & (x14207x)));
	assign n_n2997 = (((!n_n4515) & (!x170x) & (!n_n3152) & (!x129x) & (n_n4520)) + ((!n_n4515) & (!x170x) & (!n_n3152) & (x129x) & (!n_n4520)) + ((!n_n4515) & (!x170x) & (!n_n3152) & (x129x) & (n_n4520)) + ((!n_n4515) & (!x170x) & (n_n3152) & (!x129x) & (!n_n4520)) + ((!n_n4515) & (!x170x) & (n_n3152) & (!x129x) & (n_n4520)) + ((!n_n4515) & (!x170x) & (n_n3152) & (x129x) & (!n_n4520)) + ((!n_n4515) & (!x170x) & (n_n3152) & (x129x) & (n_n4520)) + ((!n_n4515) & (x170x) & (!n_n3152) & (!x129x) & (!n_n4520)) + ((!n_n4515) & (x170x) & (!n_n3152) & (!x129x) & (n_n4520)) + ((!n_n4515) & (x170x) & (!n_n3152) & (x129x) & (!n_n4520)) + ((!n_n4515) & (x170x) & (!n_n3152) & (x129x) & (n_n4520)) + ((!n_n4515) & (x170x) & (n_n3152) & (!x129x) & (!n_n4520)) + ((!n_n4515) & (x170x) & (n_n3152) & (!x129x) & (n_n4520)) + ((!n_n4515) & (x170x) & (n_n3152) & (x129x) & (!n_n4520)) + ((!n_n4515) & (x170x) & (n_n3152) & (x129x) & (n_n4520)) + ((n_n4515) & (!x170x) & (!n_n3152) & (!x129x) & (!n_n4520)) + ((n_n4515) & (!x170x) & (!n_n3152) & (!x129x) & (n_n4520)) + ((n_n4515) & (!x170x) & (!n_n3152) & (x129x) & (!n_n4520)) + ((n_n4515) & (!x170x) & (!n_n3152) & (x129x) & (n_n4520)) + ((n_n4515) & (!x170x) & (n_n3152) & (!x129x) & (!n_n4520)) + ((n_n4515) & (!x170x) & (n_n3152) & (!x129x) & (n_n4520)) + ((n_n4515) & (!x170x) & (n_n3152) & (x129x) & (!n_n4520)) + ((n_n4515) & (!x170x) & (n_n3152) & (x129x) & (n_n4520)) + ((n_n4515) & (x170x) & (!n_n3152) & (!x129x) & (!n_n4520)) + ((n_n4515) & (x170x) & (!n_n3152) & (!x129x) & (n_n4520)) + ((n_n4515) & (x170x) & (!n_n3152) & (x129x) & (!n_n4520)) + ((n_n4515) & (x170x) & (!n_n3152) & (x129x) & (n_n4520)) + ((n_n4515) & (x170x) & (n_n3152) & (!x129x) & (!n_n4520)) + ((n_n4515) & (x170x) & (n_n3152) & (!x129x) & (n_n4520)) + ((n_n4515) & (x170x) & (n_n3152) & (x129x) & (!n_n4520)) + ((n_n4515) & (x170x) & (n_n3152) & (x129x) & (n_n4520)));
	assign x15758x = (((!i_9_) & (n_n325) & (!n_n520) & (x23x) & (n_n500)) + ((!i_9_) & (n_n325) & (n_n520) & (x23x) & (n_n500)) + ((i_9_) & (n_n325) & (!n_n520) & (x23x) & (n_n500)) + ((i_9_) & (n_n325) & (n_n520) & (!x23x) & (n_n500)) + ((i_9_) & (n_n325) & (n_n520) & (x23x) & (n_n500)));
	assign n_n2979 = (((!x109x) & (!x69x) & (!n_n4752) & (!x258x) & (x15758x)) + ((!x109x) & (!x69x) & (!n_n4752) & (x258x) & (!x15758x)) + ((!x109x) & (!x69x) & (!n_n4752) & (x258x) & (x15758x)) + ((!x109x) & (!x69x) & (n_n4752) & (!x258x) & (!x15758x)) + ((!x109x) & (!x69x) & (n_n4752) & (!x258x) & (x15758x)) + ((!x109x) & (!x69x) & (n_n4752) & (x258x) & (!x15758x)) + ((!x109x) & (!x69x) & (n_n4752) & (x258x) & (x15758x)) + ((!x109x) & (x69x) & (!n_n4752) & (!x258x) & (!x15758x)) + ((!x109x) & (x69x) & (!n_n4752) & (!x258x) & (x15758x)) + ((!x109x) & (x69x) & (!n_n4752) & (x258x) & (!x15758x)) + ((!x109x) & (x69x) & (!n_n4752) & (x258x) & (x15758x)) + ((!x109x) & (x69x) & (n_n4752) & (!x258x) & (!x15758x)) + ((!x109x) & (x69x) & (n_n4752) & (!x258x) & (x15758x)) + ((!x109x) & (x69x) & (n_n4752) & (x258x) & (!x15758x)) + ((!x109x) & (x69x) & (n_n4752) & (x258x) & (x15758x)) + ((x109x) & (!x69x) & (!n_n4752) & (!x258x) & (!x15758x)) + ((x109x) & (!x69x) & (!n_n4752) & (!x258x) & (x15758x)) + ((x109x) & (!x69x) & (!n_n4752) & (x258x) & (!x15758x)) + ((x109x) & (!x69x) & (!n_n4752) & (x258x) & (x15758x)) + ((x109x) & (!x69x) & (n_n4752) & (!x258x) & (!x15758x)) + ((x109x) & (!x69x) & (n_n4752) & (!x258x) & (x15758x)) + ((x109x) & (!x69x) & (n_n4752) & (x258x) & (!x15758x)) + ((x109x) & (!x69x) & (n_n4752) & (x258x) & (x15758x)) + ((x109x) & (x69x) & (!n_n4752) & (!x258x) & (!x15758x)) + ((x109x) & (x69x) & (!n_n4752) & (!x258x) & (x15758x)) + ((x109x) & (x69x) & (!n_n4752) & (x258x) & (!x15758x)) + ((x109x) & (x69x) & (!n_n4752) & (x258x) & (x15758x)) + ((x109x) & (x69x) & (n_n4752) & (!x258x) & (!x15758x)) + ((x109x) & (x69x) & (n_n4752) & (!x258x) & (x15758x)) + ((x109x) & (x69x) & (n_n4752) & (x258x) & (!x15758x)) + ((x109x) & (x69x) & (n_n4752) & (x258x) & (x15758x)));
	assign n_n2968 = (((!n_n4903) & (!x96x) & (!n_n4896) & (!x48x) & (x49x)) + ((!n_n4903) & (!x96x) & (!n_n4896) & (x48x) & (!x49x)) + ((!n_n4903) & (!x96x) & (!n_n4896) & (x48x) & (x49x)) + ((!n_n4903) & (!x96x) & (n_n4896) & (!x48x) & (!x49x)) + ((!n_n4903) & (!x96x) & (n_n4896) & (!x48x) & (x49x)) + ((!n_n4903) & (!x96x) & (n_n4896) & (x48x) & (!x49x)) + ((!n_n4903) & (!x96x) & (n_n4896) & (x48x) & (x49x)) + ((!n_n4903) & (x96x) & (!n_n4896) & (!x48x) & (!x49x)) + ((!n_n4903) & (x96x) & (!n_n4896) & (!x48x) & (x49x)) + ((!n_n4903) & (x96x) & (!n_n4896) & (x48x) & (!x49x)) + ((!n_n4903) & (x96x) & (!n_n4896) & (x48x) & (x49x)) + ((!n_n4903) & (x96x) & (n_n4896) & (!x48x) & (!x49x)) + ((!n_n4903) & (x96x) & (n_n4896) & (!x48x) & (x49x)) + ((!n_n4903) & (x96x) & (n_n4896) & (x48x) & (!x49x)) + ((!n_n4903) & (x96x) & (n_n4896) & (x48x) & (x49x)) + ((n_n4903) & (!x96x) & (!n_n4896) & (!x48x) & (!x49x)) + ((n_n4903) & (!x96x) & (!n_n4896) & (!x48x) & (x49x)) + ((n_n4903) & (!x96x) & (!n_n4896) & (x48x) & (!x49x)) + ((n_n4903) & (!x96x) & (!n_n4896) & (x48x) & (x49x)) + ((n_n4903) & (!x96x) & (n_n4896) & (!x48x) & (!x49x)) + ((n_n4903) & (!x96x) & (n_n4896) & (!x48x) & (x49x)) + ((n_n4903) & (!x96x) & (n_n4896) & (x48x) & (!x49x)) + ((n_n4903) & (!x96x) & (n_n4896) & (x48x) & (x49x)) + ((n_n4903) & (x96x) & (!n_n4896) & (!x48x) & (!x49x)) + ((n_n4903) & (x96x) & (!n_n4896) & (!x48x) & (x49x)) + ((n_n4903) & (x96x) & (!n_n4896) & (x48x) & (!x49x)) + ((n_n4903) & (x96x) & (!n_n4896) & (x48x) & (x49x)) + ((n_n4903) & (x96x) & (n_n4896) & (!x48x) & (!x49x)) + ((n_n4903) & (x96x) & (n_n4896) & (!x48x) & (x49x)) + ((n_n4903) & (x96x) & (n_n4896) & (x48x) & (!x49x)) + ((n_n4903) & (x96x) & (n_n4896) & (x48x) & (x49x)));
	assign n_n3037 = (((!i_9_) & (!n_n528) & (!n_n535) & (!n_n65) & (n_n5216)) + ((!i_9_) & (!n_n528) & (!n_n535) & (n_n65) & (n_n5216)) + ((!i_9_) & (!n_n528) & (n_n535) & (!n_n65) & (n_n5216)) + ((!i_9_) & (!n_n528) & (n_n535) & (n_n65) & (n_n5216)) + ((!i_9_) & (n_n528) & (!n_n535) & (!n_n65) & (n_n5216)) + ((!i_9_) & (n_n528) & (!n_n535) & (n_n65) & (n_n5216)) + ((!i_9_) & (n_n528) & (n_n535) & (!n_n65) & (n_n5216)) + ((!i_9_) & (n_n528) & (n_n535) & (n_n65) & (!n_n5216)) + ((!i_9_) & (n_n528) & (n_n535) & (n_n65) & (n_n5216)) + ((i_9_) & (!n_n528) & (!n_n535) & (!n_n65) & (n_n5216)) + ((i_9_) & (!n_n528) & (!n_n535) & (n_n65) & (n_n5216)) + ((i_9_) & (!n_n528) & (n_n535) & (!n_n65) & (n_n5216)) + ((i_9_) & (!n_n528) & (n_n535) & (n_n65) & (n_n5216)) + ((i_9_) & (n_n528) & (!n_n535) & (!n_n65) & (n_n5216)) + ((i_9_) & (n_n528) & (!n_n535) & (n_n65) & (n_n5216)) + ((i_9_) & (n_n528) & (n_n535) & (!n_n65) & (n_n5216)) + ((i_9_) & (n_n528) & (n_n535) & (n_n65) & (!n_n5216)) + ((i_9_) & (n_n528) & (n_n535) & (n_n65) & (n_n5216)));
	assign x15554x = (((!n_n5200) & (!n_n5206) & (!n_n5207) & (n_n5208)) + ((!n_n5200) & (!n_n5206) & (n_n5207) & (!n_n5208)) + ((!n_n5200) & (!n_n5206) & (n_n5207) & (n_n5208)) + ((!n_n5200) & (n_n5206) & (!n_n5207) & (!n_n5208)) + ((!n_n5200) & (n_n5206) & (!n_n5207) & (n_n5208)) + ((!n_n5200) & (n_n5206) & (n_n5207) & (!n_n5208)) + ((!n_n5200) & (n_n5206) & (n_n5207) & (n_n5208)) + ((n_n5200) & (!n_n5206) & (!n_n5207) & (!n_n5208)) + ((n_n5200) & (!n_n5206) & (!n_n5207) & (n_n5208)) + ((n_n5200) & (!n_n5206) & (n_n5207) & (!n_n5208)) + ((n_n5200) & (!n_n5206) & (n_n5207) & (n_n5208)) + ((n_n5200) & (n_n5206) & (!n_n5207) & (!n_n5208)) + ((n_n5200) & (n_n5206) & (!n_n5207) & (n_n5208)) + ((n_n5200) & (n_n5206) & (n_n5207) & (!n_n5208)) + ((n_n5200) & (n_n5206) & (n_n5207) & (n_n5208)));
	assign x15555x = (((!x12x) & (!x516x) & (!n_n5199) & (!x220x) & (n_n5209)) + ((!x12x) & (!x516x) & (!n_n5199) & (x220x) & (!n_n5209)) + ((!x12x) & (!x516x) & (!n_n5199) & (x220x) & (n_n5209)) + ((!x12x) & (!x516x) & (n_n5199) & (!x220x) & (!n_n5209)) + ((!x12x) & (!x516x) & (n_n5199) & (!x220x) & (n_n5209)) + ((!x12x) & (!x516x) & (n_n5199) & (x220x) & (!n_n5209)) + ((!x12x) & (!x516x) & (n_n5199) & (x220x) & (n_n5209)) + ((!x12x) & (x516x) & (!n_n5199) & (!x220x) & (n_n5209)) + ((!x12x) & (x516x) & (!n_n5199) & (x220x) & (!n_n5209)) + ((!x12x) & (x516x) & (!n_n5199) & (x220x) & (n_n5209)) + ((!x12x) & (x516x) & (n_n5199) & (!x220x) & (!n_n5209)) + ((!x12x) & (x516x) & (n_n5199) & (!x220x) & (n_n5209)) + ((!x12x) & (x516x) & (n_n5199) & (x220x) & (!n_n5209)) + ((!x12x) & (x516x) & (n_n5199) & (x220x) & (n_n5209)) + ((x12x) & (!x516x) & (!n_n5199) & (!x220x) & (n_n5209)) + ((x12x) & (!x516x) & (!n_n5199) & (x220x) & (!n_n5209)) + ((x12x) & (!x516x) & (!n_n5199) & (x220x) & (n_n5209)) + ((x12x) & (!x516x) & (n_n5199) & (!x220x) & (!n_n5209)) + ((x12x) & (!x516x) & (n_n5199) & (!x220x) & (n_n5209)) + ((x12x) & (!x516x) & (n_n5199) & (x220x) & (!n_n5209)) + ((x12x) & (!x516x) & (n_n5199) & (x220x) & (n_n5209)) + ((x12x) & (x516x) & (!n_n5199) & (!x220x) & (!n_n5209)) + ((x12x) & (x516x) & (!n_n5199) & (!x220x) & (n_n5209)) + ((x12x) & (x516x) & (!n_n5199) & (x220x) & (!n_n5209)) + ((x12x) & (x516x) & (!n_n5199) & (x220x) & (n_n5209)) + ((x12x) & (x516x) & (n_n5199) & (!x220x) & (!n_n5209)) + ((x12x) & (x516x) & (n_n5199) & (!x220x) & (n_n5209)) + ((x12x) & (x516x) & (n_n5199) & (x220x) & (!n_n5209)) + ((x12x) & (x516x) & (n_n5199) & (x220x) & (n_n5209)));
	assign x183x = (((!i_9_) & (!n_n524) & (n_n535) & (x20x) & (n_n65)) + ((!i_9_) & (n_n524) & (n_n535) & (!x20x) & (n_n65)) + ((!i_9_) & (n_n524) & (n_n535) & (x20x) & (n_n65)) + ((i_9_) & (!n_n524) & (n_n535) & (x20x) & (n_n65)) + ((i_9_) & (n_n524) & (n_n535) & (x20x) & (n_n65)));
	assign x15562x = (((!n_n528) & (!x12x) & (!x112x) & (!n_n464) & (n_n3037)) + ((!n_n528) & (!x12x) & (!x112x) & (n_n464) & (n_n3037)) + ((!n_n528) & (!x12x) & (x112x) & (!n_n464) & (!n_n3037)) + ((!n_n528) & (!x12x) & (x112x) & (!n_n464) & (n_n3037)) + ((!n_n528) & (!x12x) & (x112x) & (n_n464) & (!n_n3037)) + ((!n_n528) & (!x12x) & (x112x) & (n_n464) & (n_n3037)) + ((!n_n528) & (x12x) & (!x112x) & (!n_n464) & (n_n3037)) + ((!n_n528) & (x12x) & (!x112x) & (n_n464) & (n_n3037)) + ((!n_n528) & (x12x) & (x112x) & (!n_n464) & (!n_n3037)) + ((!n_n528) & (x12x) & (x112x) & (!n_n464) & (n_n3037)) + ((!n_n528) & (x12x) & (x112x) & (n_n464) & (!n_n3037)) + ((!n_n528) & (x12x) & (x112x) & (n_n464) & (n_n3037)) + ((n_n528) & (!x12x) & (!x112x) & (!n_n464) & (n_n3037)) + ((n_n528) & (!x12x) & (!x112x) & (n_n464) & (n_n3037)) + ((n_n528) & (!x12x) & (x112x) & (!n_n464) & (!n_n3037)) + ((n_n528) & (!x12x) & (x112x) & (!n_n464) & (n_n3037)) + ((n_n528) & (!x12x) & (x112x) & (n_n464) & (!n_n3037)) + ((n_n528) & (!x12x) & (x112x) & (n_n464) & (n_n3037)) + ((n_n528) & (x12x) & (!x112x) & (!n_n464) & (n_n3037)) + ((n_n528) & (x12x) & (!x112x) & (n_n464) & (!n_n3037)) + ((n_n528) & (x12x) & (!x112x) & (n_n464) & (n_n3037)) + ((n_n528) & (x12x) & (x112x) & (!n_n464) & (!n_n3037)) + ((n_n528) & (x12x) & (x112x) & (!n_n464) & (n_n3037)) + ((n_n528) & (x12x) & (x112x) & (n_n464) & (!n_n3037)) + ((n_n528) & (x12x) & (x112x) & (n_n464) & (n_n3037)));
	assign x15564x = (((!n_n5183) & (!n_n5188) & (!n_n5220) & (!n_n5210) & (x15562x)) + ((!n_n5183) & (!n_n5188) & (!n_n5220) & (n_n5210) & (!x15562x)) + ((!n_n5183) & (!n_n5188) & (!n_n5220) & (n_n5210) & (x15562x)) + ((!n_n5183) & (!n_n5188) & (n_n5220) & (!n_n5210) & (!x15562x)) + ((!n_n5183) & (!n_n5188) & (n_n5220) & (!n_n5210) & (x15562x)) + ((!n_n5183) & (!n_n5188) & (n_n5220) & (n_n5210) & (!x15562x)) + ((!n_n5183) & (!n_n5188) & (n_n5220) & (n_n5210) & (x15562x)) + ((!n_n5183) & (n_n5188) & (!n_n5220) & (!n_n5210) & (!x15562x)) + ((!n_n5183) & (n_n5188) & (!n_n5220) & (!n_n5210) & (x15562x)) + ((!n_n5183) & (n_n5188) & (!n_n5220) & (n_n5210) & (!x15562x)) + ((!n_n5183) & (n_n5188) & (!n_n5220) & (n_n5210) & (x15562x)) + ((!n_n5183) & (n_n5188) & (n_n5220) & (!n_n5210) & (!x15562x)) + ((!n_n5183) & (n_n5188) & (n_n5220) & (!n_n5210) & (x15562x)) + ((!n_n5183) & (n_n5188) & (n_n5220) & (n_n5210) & (!x15562x)) + ((!n_n5183) & (n_n5188) & (n_n5220) & (n_n5210) & (x15562x)) + ((n_n5183) & (!n_n5188) & (!n_n5220) & (!n_n5210) & (!x15562x)) + ((n_n5183) & (!n_n5188) & (!n_n5220) & (!n_n5210) & (x15562x)) + ((n_n5183) & (!n_n5188) & (!n_n5220) & (n_n5210) & (!x15562x)) + ((n_n5183) & (!n_n5188) & (!n_n5220) & (n_n5210) & (x15562x)) + ((n_n5183) & (!n_n5188) & (n_n5220) & (!n_n5210) & (!x15562x)) + ((n_n5183) & (!n_n5188) & (n_n5220) & (!n_n5210) & (x15562x)) + ((n_n5183) & (!n_n5188) & (n_n5220) & (n_n5210) & (!x15562x)) + ((n_n5183) & (!n_n5188) & (n_n5220) & (n_n5210) & (x15562x)) + ((n_n5183) & (n_n5188) & (!n_n5220) & (!n_n5210) & (!x15562x)) + ((n_n5183) & (n_n5188) & (!n_n5220) & (!n_n5210) & (x15562x)) + ((n_n5183) & (n_n5188) & (!n_n5220) & (n_n5210) & (!x15562x)) + ((n_n5183) & (n_n5188) & (!n_n5220) & (n_n5210) & (x15562x)) + ((n_n5183) & (n_n5188) & (n_n5220) & (!n_n5210) & (!x15562x)) + ((n_n5183) & (n_n5188) & (n_n5220) & (!n_n5210) & (x15562x)) + ((n_n5183) & (n_n5188) & (n_n5220) & (n_n5210) & (!x15562x)) + ((n_n5183) & (n_n5188) & (n_n5220) & (n_n5210) & (x15562x)));
	assign x15563x = (((!n_n5191) & (!x454x) & (!n_n5192) & (!x453x) & (x183x)) + ((!n_n5191) & (!x454x) & (!n_n5192) & (x453x) & (!x183x)) + ((!n_n5191) & (!x454x) & (!n_n5192) & (x453x) & (x183x)) + ((!n_n5191) & (!x454x) & (n_n5192) & (!x453x) & (!x183x)) + ((!n_n5191) & (!x454x) & (n_n5192) & (!x453x) & (x183x)) + ((!n_n5191) & (!x454x) & (n_n5192) & (x453x) & (!x183x)) + ((!n_n5191) & (!x454x) & (n_n5192) & (x453x) & (x183x)) + ((!n_n5191) & (x454x) & (!n_n5192) & (!x453x) & (!x183x)) + ((!n_n5191) & (x454x) & (!n_n5192) & (!x453x) & (x183x)) + ((!n_n5191) & (x454x) & (!n_n5192) & (x453x) & (!x183x)) + ((!n_n5191) & (x454x) & (!n_n5192) & (x453x) & (x183x)) + ((!n_n5191) & (x454x) & (n_n5192) & (!x453x) & (!x183x)) + ((!n_n5191) & (x454x) & (n_n5192) & (!x453x) & (x183x)) + ((!n_n5191) & (x454x) & (n_n5192) & (x453x) & (!x183x)) + ((!n_n5191) & (x454x) & (n_n5192) & (x453x) & (x183x)) + ((n_n5191) & (!x454x) & (!n_n5192) & (!x453x) & (!x183x)) + ((n_n5191) & (!x454x) & (!n_n5192) & (!x453x) & (x183x)) + ((n_n5191) & (!x454x) & (!n_n5192) & (x453x) & (!x183x)) + ((n_n5191) & (!x454x) & (!n_n5192) & (x453x) & (x183x)) + ((n_n5191) & (!x454x) & (n_n5192) & (!x453x) & (!x183x)) + ((n_n5191) & (!x454x) & (n_n5192) & (!x453x) & (x183x)) + ((n_n5191) & (!x454x) & (n_n5192) & (x453x) & (!x183x)) + ((n_n5191) & (!x454x) & (n_n5192) & (x453x) & (x183x)) + ((n_n5191) & (x454x) & (!n_n5192) & (!x453x) & (!x183x)) + ((n_n5191) & (x454x) & (!n_n5192) & (!x453x) & (x183x)) + ((n_n5191) & (x454x) & (!n_n5192) & (x453x) & (!x183x)) + ((n_n5191) & (x454x) & (!n_n5192) & (x453x) & (x183x)) + ((n_n5191) & (x454x) & (n_n5192) & (!x453x) & (!x183x)) + ((n_n5191) & (x454x) & (n_n5192) & (!x453x) & (x183x)) + ((n_n5191) & (x454x) & (n_n5192) & (x453x) & (!x183x)) + ((n_n5191) & (x454x) & (n_n5192) & (x453x) & (x183x)));
	assign x22085x = (((!n_n5223) & (!n_n5229) & (!n_n5228) & (!n_n5225)));
	assign n_n2943 = (((!n_n5232) & (!n_n5233) & (!n_n5224) & (!x385x) & (!x22085x)) + ((!n_n5232) & (!n_n5233) & (!n_n5224) & (x385x) & (!x22085x)) + ((!n_n5232) & (!n_n5233) & (!n_n5224) & (x385x) & (x22085x)) + ((!n_n5232) & (!n_n5233) & (n_n5224) & (!x385x) & (!x22085x)) + ((!n_n5232) & (!n_n5233) & (n_n5224) & (!x385x) & (x22085x)) + ((!n_n5232) & (!n_n5233) & (n_n5224) & (x385x) & (!x22085x)) + ((!n_n5232) & (!n_n5233) & (n_n5224) & (x385x) & (x22085x)) + ((!n_n5232) & (n_n5233) & (!n_n5224) & (!x385x) & (!x22085x)) + ((!n_n5232) & (n_n5233) & (!n_n5224) & (!x385x) & (x22085x)) + ((!n_n5232) & (n_n5233) & (!n_n5224) & (x385x) & (!x22085x)) + ((!n_n5232) & (n_n5233) & (!n_n5224) & (x385x) & (x22085x)) + ((!n_n5232) & (n_n5233) & (n_n5224) & (!x385x) & (!x22085x)) + ((!n_n5232) & (n_n5233) & (n_n5224) & (!x385x) & (x22085x)) + ((!n_n5232) & (n_n5233) & (n_n5224) & (x385x) & (!x22085x)) + ((!n_n5232) & (n_n5233) & (n_n5224) & (x385x) & (x22085x)) + ((n_n5232) & (!n_n5233) & (!n_n5224) & (!x385x) & (!x22085x)) + ((n_n5232) & (!n_n5233) & (!n_n5224) & (!x385x) & (x22085x)) + ((n_n5232) & (!n_n5233) & (!n_n5224) & (x385x) & (!x22085x)) + ((n_n5232) & (!n_n5233) & (!n_n5224) & (x385x) & (x22085x)) + ((n_n5232) & (!n_n5233) & (n_n5224) & (!x385x) & (!x22085x)) + ((n_n5232) & (!n_n5233) & (n_n5224) & (!x385x) & (x22085x)) + ((n_n5232) & (!n_n5233) & (n_n5224) & (x385x) & (!x22085x)) + ((n_n5232) & (!n_n5233) & (n_n5224) & (x385x) & (x22085x)) + ((n_n5232) & (n_n5233) & (!n_n5224) & (!x385x) & (!x22085x)) + ((n_n5232) & (n_n5233) & (!n_n5224) & (!x385x) & (x22085x)) + ((n_n5232) & (n_n5233) & (!n_n5224) & (x385x) & (!x22085x)) + ((n_n5232) & (n_n5233) & (!n_n5224) & (x385x) & (x22085x)) + ((n_n5232) & (n_n5233) & (n_n5224) & (!x385x) & (!x22085x)) + ((n_n5232) & (n_n5233) & (n_n5224) & (!x385x) & (x22085x)) + ((n_n5232) & (n_n5233) & (n_n5224) & (x385x) & (!x22085x)) + ((n_n5232) & (n_n5233) & (n_n5224) & (x385x) & (x22085x)));
	assign n_n3385 = (((!n_n509) & (!x23x) & (!n_n65) & (!n_n5256) & (n_n5257)) + ((!n_n509) & (!x23x) & (!n_n65) & (n_n5256) & (!n_n5257)) + ((!n_n509) & (!x23x) & (!n_n65) & (n_n5256) & (n_n5257)) + ((!n_n509) & (!x23x) & (n_n65) & (!n_n5256) & (n_n5257)) + ((!n_n509) & (!x23x) & (n_n65) & (n_n5256) & (!n_n5257)) + ((!n_n509) & (!x23x) & (n_n65) & (n_n5256) & (n_n5257)) + ((!n_n509) & (x23x) & (!n_n65) & (!n_n5256) & (n_n5257)) + ((!n_n509) & (x23x) & (!n_n65) & (n_n5256) & (!n_n5257)) + ((!n_n509) & (x23x) & (!n_n65) & (n_n5256) & (n_n5257)) + ((!n_n509) & (x23x) & (n_n65) & (!n_n5256) & (n_n5257)) + ((!n_n509) & (x23x) & (n_n65) & (n_n5256) & (!n_n5257)) + ((!n_n509) & (x23x) & (n_n65) & (n_n5256) & (n_n5257)) + ((n_n509) & (!x23x) & (!n_n65) & (!n_n5256) & (n_n5257)) + ((n_n509) & (!x23x) & (!n_n65) & (n_n5256) & (!n_n5257)) + ((n_n509) & (!x23x) & (!n_n65) & (n_n5256) & (n_n5257)) + ((n_n509) & (!x23x) & (n_n65) & (!n_n5256) & (n_n5257)) + ((n_n509) & (!x23x) & (n_n65) & (n_n5256) & (!n_n5257)) + ((n_n509) & (!x23x) & (n_n65) & (n_n5256) & (n_n5257)) + ((n_n509) & (x23x) & (!n_n65) & (!n_n5256) & (n_n5257)) + ((n_n509) & (x23x) & (!n_n65) & (n_n5256) & (!n_n5257)) + ((n_n509) & (x23x) & (!n_n65) & (n_n5256) & (n_n5257)) + ((n_n509) & (x23x) & (n_n65) & (!n_n5256) & (!n_n5257)) + ((n_n509) & (x23x) & (n_n65) & (!n_n5256) & (n_n5257)) + ((n_n509) & (x23x) & (n_n65) & (n_n5256) & (!n_n5257)) + ((n_n509) & (x23x) & (n_n65) & (n_n5256) & (n_n5257)));
	assign x15575x = (((!n_n5241) & (!n_n5246) & (!n_n5262) & (n_n5234)) + ((!n_n5241) & (!n_n5246) & (n_n5262) & (!n_n5234)) + ((!n_n5241) & (!n_n5246) & (n_n5262) & (n_n5234)) + ((!n_n5241) & (n_n5246) & (!n_n5262) & (!n_n5234)) + ((!n_n5241) & (n_n5246) & (!n_n5262) & (n_n5234)) + ((!n_n5241) & (n_n5246) & (n_n5262) & (!n_n5234)) + ((!n_n5241) & (n_n5246) & (n_n5262) & (n_n5234)) + ((n_n5241) & (!n_n5246) & (!n_n5262) & (!n_n5234)) + ((n_n5241) & (!n_n5246) & (!n_n5262) & (n_n5234)) + ((n_n5241) & (!n_n5246) & (n_n5262) & (!n_n5234)) + ((n_n5241) & (!n_n5246) & (n_n5262) & (n_n5234)) + ((n_n5241) & (n_n5246) & (!n_n5262) & (!n_n5234)) + ((n_n5241) & (n_n5246) & (!n_n5262) & (n_n5234)) + ((n_n5241) & (n_n5246) & (n_n5262) & (!n_n5234)) + ((n_n5241) & (n_n5246) & (n_n5262) & (n_n5234)));
	assign x15577x = (((!n_n5239) & (!n_n5240) & (!x146x) & (!x62x) & (x446x)) + ((!n_n5239) & (!n_n5240) & (!x146x) & (x62x) & (!x446x)) + ((!n_n5239) & (!n_n5240) & (!x146x) & (x62x) & (x446x)) + ((!n_n5239) & (!n_n5240) & (x146x) & (!x62x) & (!x446x)) + ((!n_n5239) & (!n_n5240) & (x146x) & (!x62x) & (x446x)) + ((!n_n5239) & (!n_n5240) & (x146x) & (x62x) & (!x446x)) + ((!n_n5239) & (!n_n5240) & (x146x) & (x62x) & (x446x)) + ((!n_n5239) & (n_n5240) & (!x146x) & (!x62x) & (!x446x)) + ((!n_n5239) & (n_n5240) & (!x146x) & (!x62x) & (x446x)) + ((!n_n5239) & (n_n5240) & (!x146x) & (x62x) & (!x446x)) + ((!n_n5239) & (n_n5240) & (!x146x) & (x62x) & (x446x)) + ((!n_n5239) & (n_n5240) & (x146x) & (!x62x) & (!x446x)) + ((!n_n5239) & (n_n5240) & (x146x) & (!x62x) & (x446x)) + ((!n_n5239) & (n_n5240) & (x146x) & (x62x) & (!x446x)) + ((!n_n5239) & (n_n5240) & (x146x) & (x62x) & (x446x)) + ((n_n5239) & (!n_n5240) & (!x146x) & (!x62x) & (!x446x)) + ((n_n5239) & (!n_n5240) & (!x146x) & (!x62x) & (x446x)) + ((n_n5239) & (!n_n5240) & (!x146x) & (x62x) & (!x446x)) + ((n_n5239) & (!n_n5240) & (!x146x) & (x62x) & (x446x)) + ((n_n5239) & (!n_n5240) & (x146x) & (!x62x) & (!x446x)) + ((n_n5239) & (!n_n5240) & (x146x) & (!x62x) & (x446x)) + ((n_n5239) & (!n_n5240) & (x146x) & (x62x) & (!x446x)) + ((n_n5239) & (!n_n5240) & (x146x) & (x62x) & (x446x)) + ((n_n5239) & (n_n5240) & (!x146x) & (!x62x) & (!x446x)) + ((n_n5239) & (n_n5240) & (!x146x) & (!x62x) & (x446x)) + ((n_n5239) & (n_n5240) & (!x146x) & (x62x) & (!x446x)) + ((n_n5239) & (n_n5240) & (!x146x) & (x62x) & (x446x)) + ((n_n5239) & (n_n5240) & (x146x) & (!x62x) & (!x446x)) + ((n_n5239) & (n_n5240) & (x146x) & (!x62x) & (x446x)) + ((n_n5239) & (n_n5240) & (x146x) & (x62x) & (!x446x)) + ((n_n5239) & (n_n5240) & (x146x) & (x62x) & (x446x)));
	assign n_n2948 = (((!n_n5167) & (!n_n5163) & (!n_n5172) & (x466x)) + ((!n_n5167) & (!n_n5163) & (n_n5172) & (!x466x)) + ((!n_n5167) & (!n_n5163) & (n_n5172) & (x466x)) + ((!n_n5167) & (n_n5163) & (!n_n5172) & (!x466x)) + ((!n_n5167) & (n_n5163) & (!n_n5172) & (x466x)) + ((!n_n5167) & (n_n5163) & (n_n5172) & (!x466x)) + ((!n_n5167) & (n_n5163) & (n_n5172) & (x466x)) + ((n_n5167) & (!n_n5163) & (!n_n5172) & (!x466x)) + ((n_n5167) & (!n_n5163) & (!n_n5172) & (x466x)) + ((n_n5167) & (!n_n5163) & (n_n5172) & (!x466x)) + ((n_n5167) & (!n_n5163) & (n_n5172) & (x466x)) + ((n_n5167) & (n_n5163) & (!n_n5172) & (!x466x)) + ((n_n5167) & (n_n5163) & (!n_n5172) & (x466x)) + ((n_n5167) & (n_n5163) & (n_n5172) & (!x466x)) + ((n_n5167) & (n_n5163) & (n_n5172) & (x466x)));
	assign x22183x = (((!x21x) & (!n_n130) & (!n_n500) & (!x76x) & (!n_n5151)) + ((!x21x) & (!n_n130) & (n_n500) & (!x76x) & (!n_n5151)) + ((!x21x) & (n_n130) & (!n_n500) & (!x76x) & (!n_n5151)) + ((!x21x) & (n_n130) & (n_n500) & (!x76x) & (!n_n5151)) + ((x21x) & (!n_n130) & (!n_n500) & (!x76x) & (!n_n5151)) + ((x21x) & (!n_n130) & (n_n500) & (!x76x) & (!n_n5151)) + ((x21x) & (n_n130) & (!n_n500) & (!x76x) & (!n_n5151)));
	assign n_n2949 = (((!n_n5146) & (!n_n5152) & (!n_n5153) & (!x126x) & (!x22183x)) + ((!n_n5146) & (!n_n5152) & (!n_n5153) & (x126x) & (!x22183x)) + ((!n_n5146) & (!n_n5152) & (!n_n5153) & (x126x) & (x22183x)) + ((!n_n5146) & (!n_n5152) & (n_n5153) & (!x126x) & (!x22183x)) + ((!n_n5146) & (!n_n5152) & (n_n5153) & (!x126x) & (x22183x)) + ((!n_n5146) & (!n_n5152) & (n_n5153) & (x126x) & (!x22183x)) + ((!n_n5146) & (!n_n5152) & (n_n5153) & (x126x) & (x22183x)) + ((!n_n5146) & (n_n5152) & (!n_n5153) & (!x126x) & (!x22183x)) + ((!n_n5146) & (n_n5152) & (!n_n5153) & (!x126x) & (x22183x)) + ((!n_n5146) & (n_n5152) & (!n_n5153) & (x126x) & (!x22183x)) + ((!n_n5146) & (n_n5152) & (!n_n5153) & (x126x) & (x22183x)) + ((!n_n5146) & (n_n5152) & (n_n5153) & (!x126x) & (!x22183x)) + ((!n_n5146) & (n_n5152) & (n_n5153) & (!x126x) & (x22183x)) + ((!n_n5146) & (n_n5152) & (n_n5153) & (x126x) & (!x22183x)) + ((!n_n5146) & (n_n5152) & (n_n5153) & (x126x) & (x22183x)) + ((n_n5146) & (!n_n5152) & (!n_n5153) & (!x126x) & (!x22183x)) + ((n_n5146) & (!n_n5152) & (!n_n5153) & (!x126x) & (x22183x)) + ((n_n5146) & (!n_n5152) & (!n_n5153) & (x126x) & (!x22183x)) + ((n_n5146) & (!n_n5152) & (!n_n5153) & (x126x) & (x22183x)) + ((n_n5146) & (!n_n5152) & (n_n5153) & (!x126x) & (!x22183x)) + ((n_n5146) & (!n_n5152) & (n_n5153) & (!x126x) & (x22183x)) + ((n_n5146) & (!n_n5152) & (n_n5153) & (x126x) & (!x22183x)) + ((n_n5146) & (!n_n5152) & (n_n5153) & (x126x) & (x22183x)) + ((n_n5146) & (n_n5152) & (!n_n5153) & (!x126x) & (!x22183x)) + ((n_n5146) & (n_n5152) & (!n_n5153) & (!x126x) & (x22183x)) + ((n_n5146) & (n_n5152) & (!n_n5153) & (x126x) & (!x22183x)) + ((n_n5146) & (n_n5152) & (!n_n5153) & (x126x) & (x22183x)) + ((n_n5146) & (n_n5152) & (n_n5153) & (!x126x) & (!x22183x)) + ((n_n5146) & (n_n5152) & (n_n5153) & (!x126x) & (x22183x)) + ((n_n5146) & (n_n5152) & (n_n5153) & (x126x) & (!x22183x)) + ((n_n5146) & (n_n5152) & (n_n5153) & (x126x) & (x22183x)));
	assign x22180x = (((!n_n5174) & (!n_n5175) & (!n_n5177) & (!n_n4129) & (!n_n5176)));
	assign x22091x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x10x) & (!n_n473)) + ((!i_7_) & (!i_8_) & (!i_6_) & (!x10x) & (n_n473)) + ((!i_7_) & (!i_8_) & (!i_6_) & (x10x) & (!n_n473)) + ((!i_7_) & (!i_8_) & (!i_6_) & (x10x) & (n_n473)) + ((!i_7_) & (!i_8_) & (i_6_) & (!x10x) & (!n_n473)) + ((!i_7_) & (!i_8_) & (i_6_) & (!x10x) & (n_n473)) + ((!i_7_) & (!i_8_) & (i_6_) & (x10x) & (!n_n473)) + ((!i_7_) & (i_8_) & (!i_6_) & (!x10x) & (!n_n473)) + ((!i_7_) & (i_8_) & (!i_6_) & (!x10x) & (n_n473)) + ((!i_7_) & (i_8_) & (!i_6_) & (x10x) & (!n_n473)) + ((!i_7_) & (i_8_) & (i_6_) & (!x10x) & (!n_n473)) + ((!i_7_) & (i_8_) & (i_6_) & (!x10x) & (n_n473)) + ((!i_7_) & (i_8_) & (i_6_) & (x10x) & (!n_n473)) + ((!i_7_) & (i_8_) & (i_6_) & (x10x) & (n_n473)) + ((i_7_) & (!i_8_) & (!i_6_) & (!x10x) & (!n_n473)) + ((i_7_) & (!i_8_) & (!i_6_) & (!x10x) & (n_n473)) + ((i_7_) & (!i_8_) & (!i_6_) & (x10x) & (!n_n473)) + ((i_7_) & (!i_8_) & (i_6_) & (!x10x) & (!n_n473)) + ((i_7_) & (!i_8_) & (i_6_) & (!x10x) & (n_n473)) + ((i_7_) & (!i_8_) & (i_6_) & (x10x) & (!n_n473)) + ((i_7_) & (i_8_) & (!i_6_) & (!x10x) & (!n_n473)) + ((i_7_) & (i_8_) & (!i_6_) & (!x10x) & (n_n473)) + ((i_7_) & (i_8_) & (!i_6_) & (x10x) & (!n_n473)) + ((i_7_) & (i_8_) & (!i_6_) & (x10x) & (n_n473)) + ((i_7_) & (i_8_) & (i_6_) & (!x10x) & (!n_n473)) + ((i_7_) & (i_8_) & (i_6_) & (!x10x) & (n_n473)) + ((i_7_) & (i_8_) & (i_6_) & (x10x) & (!n_n473)) + ((i_7_) & (i_8_) & (i_6_) & (x10x) & (n_n473)));
	assign x14953x = (((!i_7_) & (!i_8_) & (!i_6_) & (x17x) & (n_n491)) + ((!i_7_) & (i_8_) & (!i_6_) & (x17x) & (n_n491)) + ((i_7_) & (i_8_) & (!i_6_) & (x17x) & (n_n491)));
	assign x14955x = (((!n_n482) & (!n_n532) & (!x17x) & (!n_n4905) & (x14953x)) + ((!n_n482) & (!n_n532) & (!x17x) & (n_n4905) & (!x14953x)) + ((!n_n482) & (!n_n532) & (!x17x) & (n_n4905) & (x14953x)) + ((!n_n482) & (!n_n532) & (x17x) & (!n_n4905) & (x14953x)) + ((!n_n482) & (!n_n532) & (x17x) & (n_n4905) & (!x14953x)) + ((!n_n482) & (!n_n532) & (x17x) & (n_n4905) & (x14953x)) + ((!n_n482) & (n_n532) & (!x17x) & (!n_n4905) & (x14953x)) + ((!n_n482) & (n_n532) & (!x17x) & (n_n4905) & (!x14953x)) + ((!n_n482) & (n_n532) & (!x17x) & (n_n4905) & (x14953x)) + ((!n_n482) & (n_n532) & (x17x) & (!n_n4905) & (x14953x)) + ((!n_n482) & (n_n532) & (x17x) & (n_n4905) & (!x14953x)) + ((!n_n482) & (n_n532) & (x17x) & (n_n4905) & (x14953x)) + ((n_n482) & (!n_n532) & (!x17x) & (!n_n4905) & (x14953x)) + ((n_n482) & (!n_n532) & (!x17x) & (n_n4905) & (!x14953x)) + ((n_n482) & (!n_n532) & (!x17x) & (n_n4905) & (x14953x)) + ((n_n482) & (!n_n532) & (x17x) & (!n_n4905) & (x14953x)) + ((n_n482) & (!n_n532) & (x17x) & (n_n4905) & (!x14953x)) + ((n_n482) & (!n_n532) & (x17x) & (n_n4905) & (x14953x)) + ((n_n482) & (n_n532) & (!x17x) & (!n_n4905) & (x14953x)) + ((n_n482) & (n_n532) & (!x17x) & (n_n4905) & (!x14953x)) + ((n_n482) & (n_n532) & (!x17x) & (n_n4905) & (x14953x)) + ((n_n482) & (n_n532) & (x17x) & (!n_n4905) & (!x14953x)) + ((n_n482) & (n_n532) & (x17x) & (!n_n4905) & (x14953x)) + ((n_n482) & (n_n532) & (x17x) & (n_n4905) & (!x14953x)) + ((n_n482) & (n_n532) & (x17x) & (n_n4905) & (x14953x)));
	assign n_n2718 = (((!i_9_) & (n_n482) & (!n_n528) & (n_n260) & (n_n530)) + ((!i_9_) & (n_n482) & (n_n528) & (n_n260) & (!n_n530)) + ((!i_9_) & (n_n482) & (n_n528) & (n_n260) & (n_n530)) + ((i_9_) & (n_n482) & (n_n528) & (n_n260) & (!n_n530)) + ((i_9_) & (n_n482) & (n_n528) & (n_n260) & (n_n530)));
	assign x22094x = (((!n_n5050) & (!n_n5060) & (!n_n5057) & (!n_n5061)));
	assign n_n2584 = (((!n_n5055) & (!n_n5058) & (!n_n5056) & (!x166x) & (!x22094x)) + ((!n_n5055) & (!n_n5058) & (!n_n5056) & (x166x) & (!x22094x)) + ((!n_n5055) & (!n_n5058) & (!n_n5056) & (x166x) & (x22094x)) + ((!n_n5055) & (!n_n5058) & (n_n5056) & (!x166x) & (!x22094x)) + ((!n_n5055) & (!n_n5058) & (n_n5056) & (!x166x) & (x22094x)) + ((!n_n5055) & (!n_n5058) & (n_n5056) & (x166x) & (!x22094x)) + ((!n_n5055) & (!n_n5058) & (n_n5056) & (x166x) & (x22094x)) + ((!n_n5055) & (n_n5058) & (!n_n5056) & (!x166x) & (!x22094x)) + ((!n_n5055) & (n_n5058) & (!n_n5056) & (!x166x) & (x22094x)) + ((!n_n5055) & (n_n5058) & (!n_n5056) & (x166x) & (!x22094x)) + ((!n_n5055) & (n_n5058) & (!n_n5056) & (x166x) & (x22094x)) + ((!n_n5055) & (n_n5058) & (n_n5056) & (!x166x) & (!x22094x)) + ((!n_n5055) & (n_n5058) & (n_n5056) & (!x166x) & (x22094x)) + ((!n_n5055) & (n_n5058) & (n_n5056) & (x166x) & (!x22094x)) + ((!n_n5055) & (n_n5058) & (n_n5056) & (x166x) & (x22094x)) + ((n_n5055) & (!n_n5058) & (!n_n5056) & (!x166x) & (!x22094x)) + ((n_n5055) & (!n_n5058) & (!n_n5056) & (!x166x) & (x22094x)) + ((n_n5055) & (!n_n5058) & (!n_n5056) & (x166x) & (!x22094x)) + ((n_n5055) & (!n_n5058) & (!n_n5056) & (x166x) & (x22094x)) + ((n_n5055) & (!n_n5058) & (n_n5056) & (!x166x) & (!x22094x)) + ((n_n5055) & (!n_n5058) & (n_n5056) & (!x166x) & (x22094x)) + ((n_n5055) & (!n_n5058) & (n_n5056) & (x166x) & (!x22094x)) + ((n_n5055) & (!n_n5058) & (n_n5056) & (x166x) & (x22094x)) + ((n_n5055) & (n_n5058) & (!n_n5056) & (!x166x) & (!x22094x)) + ((n_n5055) & (n_n5058) & (!n_n5056) & (!x166x) & (x22094x)) + ((n_n5055) & (n_n5058) & (!n_n5056) & (x166x) & (!x22094x)) + ((n_n5055) & (n_n5058) & (!n_n5056) & (x166x) & (x22094x)) + ((n_n5055) & (n_n5058) & (n_n5056) & (!x166x) & (!x22094x)) + ((n_n5055) & (n_n5058) & (n_n5056) & (!x166x) & (x22094x)) + ((n_n5055) & (n_n5058) & (n_n5056) & (x166x) & (!x22094x)) + ((n_n5055) & (n_n5058) & (n_n5056) & (x166x) & (x22094x)));
	assign x15232x = (((!n_n524) & (!n_n535) & (!x12x) & (!n_n4152) & (n_n5065)) + ((!n_n524) & (!n_n535) & (!x12x) & (n_n4152) & (!n_n5065)) + ((!n_n524) & (!n_n535) & (!x12x) & (n_n4152) & (n_n5065)) + ((!n_n524) & (!n_n535) & (x12x) & (!n_n4152) & (n_n5065)) + ((!n_n524) & (!n_n535) & (x12x) & (n_n4152) & (!n_n5065)) + ((!n_n524) & (!n_n535) & (x12x) & (n_n4152) & (n_n5065)) + ((!n_n524) & (n_n535) & (!x12x) & (!n_n4152) & (n_n5065)) + ((!n_n524) & (n_n535) & (!x12x) & (n_n4152) & (!n_n5065)) + ((!n_n524) & (n_n535) & (!x12x) & (n_n4152) & (n_n5065)) + ((!n_n524) & (n_n535) & (x12x) & (!n_n4152) & (n_n5065)) + ((!n_n524) & (n_n535) & (x12x) & (n_n4152) & (!n_n5065)) + ((!n_n524) & (n_n535) & (x12x) & (n_n4152) & (n_n5065)) + ((n_n524) & (!n_n535) & (!x12x) & (!n_n4152) & (n_n5065)) + ((n_n524) & (!n_n535) & (!x12x) & (n_n4152) & (!n_n5065)) + ((n_n524) & (!n_n535) & (!x12x) & (n_n4152) & (n_n5065)) + ((n_n524) & (!n_n535) & (x12x) & (!n_n4152) & (n_n5065)) + ((n_n524) & (!n_n535) & (x12x) & (n_n4152) & (!n_n5065)) + ((n_n524) & (!n_n535) & (x12x) & (n_n4152) & (n_n5065)) + ((n_n524) & (n_n535) & (!x12x) & (!n_n4152) & (n_n5065)) + ((n_n524) & (n_n535) & (!x12x) & (n_n4152) & (!n_n5065)) + ((n_n524) & (n_n535) & (!x12x) & (n_n4152) & (n_n5065)) + ((n_n524) & (n_n535) & (x12x) & (!n_n4152) & (!n_n5065)) + ((n_n524) & (n_n535) & (x12x) & (!n_n4152) & (n_n5065)) + ((n_n524) & (n_n535) & (x12x) & (n_n4152) & (!n_n5065)) + ((n_n524) & (n_n535) & (x12x) & (n_n4152) & (n_n5065)));
	assign x22093x = (((!x344x) & (!n_n5070) & (!n_n5082) & (!x123x) & (!x159x)));
	assign x15239x = (((!n_n5129) & (!n_n5124) & (!n_n5122) & (n_n5128)) + ((!n_n5129) & (!n_n5124) & (n_n5122) & (!n_n5128)) + ((!n_n5129) & (!n_n5124) & (n_n5122) & (n_n5128)) + ((!n_n5129) & (n_n5124) & (!n_n5122) & (!n_n5128)) + ((!n_n5129) & (n_n5124) & (!n_n5122) & (n_n5128)) + ((!n_n5129) & (n_n5124) & (n_n5122) & (!n_n5128)) + ((!n_n5129) & (n_n5124) & (n_n5122) & (n_n5128)) + ((n_n5129) & (!n_n5124) & (!n_n5122) & (!n_n5128)) + ((n_n5129) & (!n_n5124) & (!n_n5122) & (n_n5128)) + ((n_n5129) & (!n_n5124) & (n_n5122) & (!n_n5128)) + ((n_n5129) & (!n_n5124) & (n_n5122) & (n_n5128)) + ((n_n5129) & (n_n5124) & (!n_n5122) & (!n_n5128)) + ((n_n5129) & (n_n5124) & (!n_n5122) & (n_n5128)) + ((n_n5129) & (n_n5124) & (n_n5122) & (!n_n5128)) + ((n_n5129) & (n_n5124) & (n_n5122) & (n_n5128)));
	assign x15240x = (((!n_n5120) & (!n_n5117) & (!n_n5119) & (!n_n5125) & (n_n5126)) + ((!n_n5120) & (!n_n5117) & (!n_n5119) & (n_n5125) & (!n_n5126)) + ((!n_n5120) & (!n_n5117) & (!n_n5119) & (n_n5125) & (n_n5126)) + ((!n_n5120) & (!n_n5117) & (n_n5119) & (!n_n5125) & (!n_n5126)) + ((!n_n5120) & (!n_n5117) & (n_n5119) & (!n_n5125) & (n_n5126)) + ((!n_n5120) & (!n_n5117) & (n_n5119) & (n_n5125) & (!n_n5126)) + ((!n_n5120) & (!n_n5117) & (n_n5119) & (n_n5125) & (n_n5126)) + ((!n_n5120) & (n_n5117) & (!n_n5119) & (!n_n5125) & (!n_n5126)) + ((!n_n5120) & (n_n5117) & (!n_n5119) & (!n_n5125) & (n_n5126)) + ((!n_n5120) & (n_n5117) & (!n_n5119) & (n_n5125) & (!n_n5126)) + ((!n_n5120) & (n_n5117) & (!n_n5119) & (n_n5125) & (n_n5126)) + ((!n_n5120) & (n_n5117) & (n_n5119) & (!n_n5125) & (!n_n5126)) + ((!n_n5120) & (n_n5117) & (n_n5119) & (!n_n5125) & (n_n5126)) + ((!n_n5120) & (n_n5117) & (n_n5119) & (n_n5125) & (!n_n5126)) + ((!n_n5120) & (n_n5117) & (n_n5119) & (n_n5125) & (n_n5126)) + ((n_n5120) & (!n_n5117) & (!n_n5119) & (!n_n5125) & (!n_n5126)) + ((n_n5120) & (!n_n5117) & (!n_n5119) & (!n_n5125) & (n_n5126)) + ((n_n5120) & (!n_n5117) & (!n_n5119) & (n_n5125) & (!n_n5126)) + ((n_n5120) & (!n_n5117) & (!n_n5119) & (n_n5125) & (n_n5126)) + ((n_n5120) & (!n_n5117) & (n_n5119) & (!n_n5125) & (!n_n5126)) + ((n_n5120) & (!n_n5117) & (n_n5119) & (!n_n5125) & (n_n5126)) + ((n_n5120) & (!n_n5117) & (n_n5119) & (n_n5125) & (!n_n5126)) + ((n_n5120) & (!n_n5117) & (n_n5119) & (n_n5125) & (n_n5126)) + ((n_n5120) & (n_n5117) & (!n_n5119) & (!n_n5125) & (!n_n5126)) + ((n_n5120) & (n_n5117) & (!n_n5119) & (!n_n5125) & (n_n5126)) + ((n_n5120) & (n_n5117) & (!n_n5119) & (n_n5125) & (!n_n5126)) + ((n_n5120) & (n_n5117) & (!n_n5119) & (n_n5125) & (n_n5126)) + ((n_n5120) & (n_n5117) & (n_n5119) & (!n_n5125) & (!n_n5126)) + ((n_n5120) & (n_n5117) & (n_n5119) & (!n_n5125) & (n_n5126)) + ((n_n5120) & (n_n5117) & (n_n5119) & (n_n5125) & (!n_n5126)) + ((n_n5120) & (n_n5117) & (n_n5119) & (n_n5125) & (n_n5126)));
	assign x88x = (((i_5_) & (i_3_) & (i_4_) & (n_n520) & (x12x)));
	assign x15249x = (((!n_n4148) & (!n_n5108) & (!x28x) & (x88x)) + ((!n_n4148) & (!n_n5108) & (x28x) & (!x88x)) + ((!n_n4148) & (!n_n5108) & (x28x) & (x88x)) + ((!n_n4148) & (n_n5108) & (!x28x) & (!x88x)) + ((!n_n4148) & (n_n5108) & (!x28x) & (x88x)) + ((!n_n4148) & (n_n5108) & (x28x) & (!x88x)) + ((!n_n4148) & (n_n5108) & (x28x) & (x88x)) + ((n_n4148) & (!n_n5108) & (!x28x) & (!x88x)) + ((n_n4148) & (!n_n5108) & (!x28x) & (x88x)) + ((n_n4148) & (!n_n5108) & (x28x) & (!x88x)) + ((n_n4148) & (!n_n5108) & (x28x) & (x88x)) + ((n_n4148) & (n_n5108) & (!x28x) & (!x88x)) + ((n_n4148) & (n_n5108) & (!x28x) & (x88x)) + ((n_n4148) & (n_n5108) & (x28x) & (!x88x)) + ((n_n4148) & (n_n5108) & (x28x) & (x88x)));
	assign x15248x = (((!n_n5096) & (!n_n5099) & (!n_n5101) & (!n_n5107) & (x15246x)) + ((!n_n5096) & (!n_n5099) & (!n_n5101) & (n_n5107) & (!x15246x)) + ((!n_n5096) & (!n_n5099) & (!n_n5101) & (n_n5107) & (x15246x)) + ((!n_n5096) & (!n_n5099) & (n_n5101) & (!n_n5107) & (!x15246x)) + ((!n_n5096) & (!n_n5099) & (n_n5101) & (!n_n5107) & (x15246x)) + ((!n_n5096) & (!n_n5099) & (n_n5101) & (n_n5107) & (!x15246x)) + ((!n_n5096) & (!n_n5099) & (n_n5101) & (n_n5107) & (x15246x)) + ((!n_n5096) & (n_n5099) & (!n_n5101) & (!n_n5107) & (!x15246x)) + ((!n_n5096) & (n_n5099) & (!n_n5101) & (!n_n5107) & (x15246x)) + ((!n_n5096) & (n_n5099) & (!n_n5101) & (n_n5107) & (!x15246x)) + ((!n_n5096) & (n_n5099) & (!n_n5101) & (n_n5107) & (x15246x)) + ((!n_n5096) & (n_n5099) & (n_n5101) & (!n_n5107) & (!x15246x)) + ((!n_n5096) & (n_n5099) & (n_n5101) & (!n_n5107) & (x15246x)) + ((!n_n5096) & (n_n5099) & (n_n5101) & (n_n5107) & (!x15246x)) + ((!n_n5096) & (n_n5099) & (n_n5101) & (n_n5107) & (x15246x)) + ((n_n5096) & (!n_n5099) & (!n_n5101) & (!n_n5107) & (!x15246x)) + ((n_n5096) & (!n_n5099) & (!n_n5101) & (!n_n5107) & (x15246x)) + ((n_n5096) & (!n_n5099) & (!n_n5101) & (n_n5107) & (!x15246x)) + ((n_n5096) & (!n_n5099) & (!n_n5101) & (n_n5107) & (x15246x)) + ((n_n5096) & (!n_n5099) & (n_n5101) & (!n_n5107) & (!x15246x)) + ((n_n5096) & (!n_n5099) & (n_n5101) & (!n_n5107) & (x15246x)) + ((n_n5096) & (!n_n5099) & (n_n5101) & (n_n5107) & (!x15246x)) + ((n_n5096) & (!n_n5099) & (n_n5101) & (n_n5107) & (x15246x)) + ((n_n5096) & (n_n5099) & (!n_n5101) & (!n_n5107) & (!x15246x)) + ((n_n5096) & (n_n5099) & (!n_n5101) & (!n_n5107) & (x15246x)) + ((n_n5096) & (n_n5099) & (!n_n5101) & (n_n5107) & (!x15246x)) + ((n_n5096) & (n_n5099) & (!n_n5101) & (n_n5107) & (x15246x)) + ((n_n5096) & (n_n5099) & (n_n5101) & (!n_n5107) & (!x15246x)) + ((n_n5096) & (n_n5099) & (n_n5101) & (!n_n5107) & (x15246x)) + ((n_n5096) & (n_n5099) & (n_n5101) & (n_n5107) & (!x15246x)) + ((n_n5096) & (n_n5099) & (n_n5101) & (n_n5107) & (x15246x)));
	assign x15254x = (((!n_n482) & (!x18x) & (!n_n530) & (!n_n5049) & (x253x)) + ((!n_n482) & (!x18x) & (!n_n530) & (n_n5049) & (!x253x)) + ((!n_n482) & (!x18x) & (!n_n530) & (n_n5049) & (x253x)) + ((!n_n482) & (!x18x) & (n_n530) & (!n_n5049) & (x253x)) + ((!n_n482) & (!x18x) & (n_n530) & (n_n5049) & (!x253x)) + ((!n_n482) & (!x18x) & (n_n530) & (n_n5049) & (x253x)) + ((!n_n482) & (x18x) & (!n_n530) & (!n_n5049) & (x253x)) + ((!n_n482) & (x18x) & (!n_n530) & (n_n5049) & (!x253x)) + ((!n_n482) & (x18x) & (!n_n530) & (n_n5049) & (x253x)) + ((!n_n482) & (x18x) & (n_n530) & (!n_n5049) & (x253x)) + ((!n_n482) & (x18x) & (n_n530) & (n_n5049) & (!x253x)) + ((!n_n482) & (x18x) & (n_n530) & (n_n5049) & (x253x)) + ((n_n482) & (!x18x) & (!n_n530) & (!n_n5049) & (x253x)) + ((n_n482) & (!x18x) & (!n_n530) & (n_n5049) & (!x253x)) + ((n_n482) & (!x18x) & (!n_n530) & (n_n5049) & (x253x)) + ((n_n482) & (!x18x) & (n_n530) & (!n_n5049) & (x253x)) + ((n_n482) & (!x18x) & (n_n530) & (n_n5049) & (!x253x)) + ((n_n482) & (!x18x) & (n_n530) & (n_n5049) & (x253x)) + ((n_n482) & (x18x) & (!n_n530) & (!n_n5049) & (x253x)) + ((n_n482) & (x18x) & (!n_n530) & (n_n5049) & (!x253x)) + ((n_n482) & (x18x) & (!n_n530) & (n_n5049) & (x253x)) + ((n_n482) & (x18x) & (n_n530) & (!n_n5049) & (!x253x)) + ((n_n482) & (x18x) & (n_n530) & (!n_n5049) & (x253x)) + ((n_n482) & (x18x) & (n_n530) & (n_n5049) & (!x253x)) + ((n_n482) & (x18x) & (n_n530) & (n_n5049) & (x253x)));
	assign x15255x = (((!n_n5046) & (!n_n5044) & (!n_n5037) & (!n_n5043) & (n_n5039)) + ((!n_n5046) & (!n_n5044) & (!n_n5037) & (n_n5043) & (!n_n5039)) + ((!n_n5046) & (!n_n5044) & (!n_n5037) & (n_n5043) & (n_n5039)) + ((!n_n5046) & (!n_n5044) & (n_n5037) & (!n_n5043) & (!n_n5039)) + ((!n_n5046) & (!n_n5044) & (n_n5037) & (!n_n5043) & (n_n5039)) + ((!n_n5046) & (!n_n5044) & (n_n5037) & (n_n5043) & (!n_n5039)) + ((!n_n5046) & (!n_n5044) & (n_n5037) & (n_n5043) & (n_n5039)) + ((!n_n5046) & (n_n5044) & (!n_n5037) & (!n_n5043) & (!n_n5039)) + ((!n_n5046) & (n_n5044) & (!n_n5037) & (!n_n5043) & (n_n5039)) + ((!n_n5046) & (n_n5044) & (!n_n5037) & (n_n5043) & (!n_n5039)) + ((!n_n5046) & (n_n5044) & (!n_n5037) & (n_n5043) & (n_n5039)) + ((!n_n5046) & (n_n5044) & (n_n5037) & (!n_n5043) & (!n_n5039)) + ((!n_n5046) & (n_n5044) & (n_n5037) & (!n_n5043) & (n_n5039)) + ((!n_n5046) & (n_n5044) & (n_n5037) & (n_n5043) & (!n_n5039)) + ((!n_n5046) & (n_n5044) & (n_n5037) & (n_n5043) & (n_n5039)) + ((n_n5046) & (!n_n5044) & (!n_n5037) & (!n_n5043) & (!n_n5039)) + ((n_n5046) & (!n_n5044) & (!n_n5037) & (!n_n5043) & (n_n5039)) + ((n_n5046) & (!n_n5044) & (!n_n5037) & (n_n5043) & (!n_n5039)) + ((n_n5046) & (!n_n5044) & (!n_n5037) & (n_n5043) & (n_n5039)) + ((n_n5046) & (!n_n5044) & (n_n5037) & (!n_n5043) & (!n_n5039)) + ((n_n5046) & (!n_n5044) & (n_n5037) & (!n_n5043) & (n_n5039)) + ((n_n5046) & (!n_n5044) & (n_n5037) & (n_n5043) & (!n_n5039)) + ((n_n5046) & (!n_n5044) & (n_n5037) & (n_n5043) & (n_n5039)) + ((n_n5046) & (n_n5044) & (!n_n5037) & (!n_n5043) & (!n_n5039)) + ((n_n5046) & (n_n5044) & (!n_n5037) & (!n_n5043) & (n_n5039)) + ((n_n5046) & (n_n5044) & (!n_n5037) & (n_n5043) & (!n_n5039)) + ((n_n5046) & (n_n5044) & (!n_n5037) & (n_n5043) & (n_n5039)) + ((n_n5046) & (n_n5044) & (n_n5037) & (!n_n5043) & (!n_n5039)) + ((n_n5046) & (n_n5044) & (n_n5037) & (!n_n5043) & (n_n5039)) + ((n_n5046) & (n_n5044) & (n_n5037) & (n_n5043) & (!n_n5039)) + ((n_n5046) & (n_n5044) & (n_n5037) & (n_n5043) & (n_n5039)));
	assign x265x = (((!i_9_) & (n_n526) & (n_n491) & (n_n195)) + ((i_9_) & (n_n526) & (n_n491) & (n_n195)));
	assign n_n2586 = (((!n_n5026) & (!n_n5023) & (!x111x) & (!x458x) & (x265x)) + ((!n_n5026) & (!n_n5023) & (!x111x) & (x458x) & (!x265x)) + ((!n_n5026) & (!n_n5023) & (!x111x) & (x458x) & (x265x)) + ((!n_n5026) & (!n_n5023) & (x111x) & (!x458x) & (!x265x)) + ((!n_n5026) & (!n_n5023) & (x111x) & (!x458x) & (x265x)) + ((!n_n5026) & (!n_n5023) & (x111x) & (x458x) & (!x265x)) + ((!n_n5026) & (!n_n5023) & (x111x) & (x458x) & (x265x)) + ((!n_n5026) & (n_n5023) & (!x111x) & (!x458x) & (!x265x)) + ((!n_n5026) & (n_n5023) & (!x111x) & (!x458x) & (x265x)) + ((!n_n5026) & (n_n5023) & (!x111x) & (x458x) & (!x265x)) + ((!n_n5026) & (n_n5023) & (!x111x) & (x458x) & (x265x)) + ((!n_n5026) & (n_n5023) & (x111x) & (!x458x) & (!x265x)) + ((!n_n5026) & (n_n5023) & (x111x) & (!x458x) & (x265x)) + ((!n_n5026) & (n_n5023) & (x111x) & (x458x) & (!x265x)) + ((!n_n5026) & (n_n5023) & (x111x) & (x458x) & (x265x)) + ((n_n5026) & (!n_n5023) & (!x111x) & (!x458x) & (!x265x)) + ((n_n5026) & (!n_n5023) & (!x111x) & (!x458x) & (x265x)) + ((n_n5026) & (!n_n5023) & (!x111x) & (x458x) & (!x265x)) + ((n_n5026) & (!n_n5023) & (!x111x) & (x458x) & (x265x)) + ((n_n5026) & (!n_n5023) & (x111x) & (!x458x) & (!x265x)) + ((n_n5026) & (!n_n5023) & (x111x) & (!x458x) & (x265x)) + ((n_n5026) & (!n_n5023) & (x111x) & (x458x) & (!x265x)) + ((n_n5026) & (!n_n5023) & (x111x) & (x458x) & (x265x)) + ((n_n5026) & (n_n5023) & (!x111x) & (!x458x) & (!x265x)) + ((n_n5026) & (n_n5023) & (!x111x) & (!x458x) & (x265x)) + ((n_n5026) & (n_n5023) & (!x111x) & (x458x) & (!x265x)) + ((n_n5026) & (n_n5023) & (!x111x) & (x458x) & (x265x)) + ((n_n5026) & (n_n5023) & (x111x) & (!x458x) & (!x265x)) + ((n_n5026) & (n_n5023) & (x111x) & (!x458x) & (x265x)) + ((n_n5026) & (n_n5023) & (x111x) & (x458x) & (!x265x)) + ((n_n5026) & (n_n5023) & (x111x) & (x458x) & (x265x)));
	assign x297x = (((!i_9_) & (!n_n534) & (n_n491) & (n_n195) & (n_n530)) + ((!i_9_) & (n_n534) & (n_n491) & (n_n195) & (!n_n530)) + ((!i_9_) & (n_n534) & (n_n491) & (n_n195) & (n_n530)));
	assign x394x = (((!i_9_) & (n_n526) & (n_n195) & (n_n500)) + ((i_9_) & (n_n526) & (n_n195) & (n_n500)));
	assign x15262x = (((!n_n5022) & (!n_n5011) & (!n_n3427) & (!x297x) & (x394x)) + ((!n_n5022) & (!n_n5011) & (!n_n3427) & (x297x) & (!x394x)) + ((!n_n5022) & (!n_n5011) & (!n_n3427) & (x297x) & (x394x)) + ((!n_n5022) & (!n_n5011) & (n_n3427) & (!x297x) & (!x394x)) + ((!n_n5022) & (!n_n5011) & (n_n3427) & (!x297x) & (x394x)) + ((!n_n5022) & (!n_n5011) & (n_n3427) & (x297x) & (!x394x)) + ((!n_n5022) & (!n_n5011) & (n_n3427) & (x297x) & (x394x)) + ((!n_n5022) & (n_n5011) & (!n_n3427) & (!x297x) & (!x394x)) + ((!n_n5022) & (n_n5011) & (!n_n3427) & (!x297x) & (x394x)) + ((!n_n5022) & (n_n5011) & (!n_n3427) & (x297x) & (!x394x)) + ((!n_n5022) & (n_n5011) & (!n_n3427) & (x297x) & (x394x)) + ((!n_n5022) & (n_n5011) & (n_n3427) & (!x297x) & (!x394x)) + ((!n_n5022) & (n_n5011) & (n_n3427) & (!x297x) & (x394x)) + ((!n_n5022) & (n_n5011) & (n_n3427) & (x297x) & (!x394x)) + ((!n_n5022) & (n_n5011) & (n_n3427) & (x297x) & (x394x)) + ((n_n5022) & (!n_n5011) & (!n_n3427) & (!x297x) & (!x394x)) + ((n_n5022) & (!n_n5011) & (!n_n3427) & (!x297x) & (x394x)) + ((n_n5022) & (!n_n5011) & (!n_n3427) & (x297x) & (!x394x)) + ((n_n5022) & (!n_n5011) & (!n_n3427) & (x297x) & (x394x)) + ((n_n5022) & (!n_n5011) & (n_n3427) & (!x297x) & (!x394x)) + ((n_n5022) & (!n_n5011) & (n_n3427) & (!x297x) & (x394x)) + ((n_n5022) & (!n_n5011) & (n_n3427) & (x297x) & (!x394x)) + ((n_n5022) & (!n_n5011) & (n_n3427) & (x297x) & (x394x)) + ((n_n5022) & (n_n5011) & (!n_n3427) & (!x297x) & (!x394x)) + ((n_n5022) & (n_n5011) & (!n_n3427) & (!x297x) & (x394x)) + ((n_n5022) & (n_n5011) & (!n_n3427) & (x297x) & (!x394x)) + ((n_n5022) & (n_n5011) & (!n_n3427) & (x297x) & (x394x)) + ((n_n5022) & (n_n5011) & (n_n3427) & (!x297x) & (!x394x)) + ((n_n5022) & (n_n5011) & (n_n3427) & (!x297x) & (x394x)) + ((n_n5022) & (n_n5011) & (n_n3427) & (x297x) & (!x394x)) + ((n_n5022) & (n_n5011) & (n_n3427) & (x297x) & (x394x)));
	assign x361x = (((!i_9_) & (n_n482) & (n_n455) & (n_n530)) + ((i_9_) & (n_n482) & (n_n455) & (n_n530)));
	assign x378x = (((!i_9_) & (n_n482) & (n_n455) & (n_n528)) + ((i_9_) & (n_n482) & (n_n455) & (n_n528)));
	assign x14542x = (((!i_9_) & (!x19x) & (n_n491) & (n_n520) & (n_n65)) + ((!i_9_) & (x19x) & (n_n491) & (n_n520) & (!n_n65)) + ((!i_9_) & (x19x) & (n_n491) & (n_n520) & (n_n65)) + ((i_9_) & (x19x) & (n_n491) & (n_n520) & (!n_n65)) + ((i_9_) & (x19x) & (n_n491) & (n_n520) & (n_n65)));
	assign n_n801 = (((!n_n528) & (!x18x) & (!n_n500) & (!n_n530) & (n_n5003)) + ((!n_n528) & (!x18x) & (!n_n500) & (n_n530) & (n_n5003)) + ((!n_n528) & (!x18x) & (n_n500) & (!n_n530) & (n_n5003)) + ((!n_n528) & (!x18x) & (n_n500) & (n_n530) & (n_n5003)) + ((!n_n528) & (x18x) & (!n_n500) & (!n_n530) & (n_n5003)) + ((!n_n528) & (x18x) & (!n_n500) & (n_n530) & (n_n5003)) + ((!n_n528) & (x18x) & (n_n500) & (!n_n530) & (n_n5003)) + ((!n_n528) & (x18x) & (n_n500) & (n_n530) & (!n_n5003)) + ((!n_n528) & (x18x) & (n_n500) & (n_n530) & (n_n5003)) + ((n_n528) & (!x18x) & (!n_n500) & (!n_n530) & (n_n5003)) + ((n_n528) & (!x18x) & (!n_n500) & (n_n530) & (n_n5003)) + ((n_n528) & (!x18x) & (n_n500) & (!n_n530) & (n_n5003)) + ((n_n528) & (!x18x) & (n_n500) & (n_n530) & (n_n5003)) + ((n_n528) & (x18x) & (!n_n500) & (!n_n530) & (n_n5003)) + ((n_n528) & (x18x) & (!n_n500) & (n_n530) & (n_n5003)) + ((n_n528) & (x18x) & (n_n500) & (!n_n530) & (!n_n5003)) + ((n_n528) & (x18x) & (n_n500) & (!n_n530) & (n_n5003)) + ((n_n528) & (x18x) & (n_n500) & (n_n530) & (!n_n5003)) + ((n_n528) & (x18x) & (n_n500) & (n_n530) & (n_n5003)));
	assign x405x = (((!i_9_) & (!n_n524) & (n_n522) & (n_n195) & (n_n500)) + ((!i_9_) & (n_n524) & (!n_n522) & (n_n195) & (n_n500)) + ((!i_9_) & (n_n524) & (n_n522) & (n_n195) & (n_n500)) + ((i_9_) & (!n_n524) & (n_n522) & (n_n195) & (n_n500)) + ((i_9_) & (n_n524) & (!n_n522) & (n_n195) & (n_n500)) + ((i_9_) & (n_n524) & (n_n522) & (n_n195) & (n_n500)));
	assign n_n1454 = (((!n_n5007) & (!n_n5008) & (!n_n801) & (x405x)) + ((!n_n5007) & (!n_n5008) & (n_n801) & (!x405x)) + ((!n_n5007) & (!n_n5008) & (n_n801) & (x405x)) + ((!n_n5007) & (n_n5008) & (!n_n801) & (!x405x)) + ((!n_n5007) & (n_n5008) & (!n_n801) & (x405x)) + ((!n_n5007) & (n_n5008) & (n_n801) & (!x405x)) + ((!n_n5007) & (n_n5008) & (n_n801) & (x405x)) + ((n_n5007) & (!n_n5008) & (!n_n801) & (!x405x)) + ((n_n5007) & (!n_n5008) & (!n_n801) & (x405x)) + ((n_n5007) & (!n_n5008) & (n_n801) & (!x405x)) + ((n_n5007) & (!n_n5008) & (n_n801) & (x405x)) + ((n_n5007) & (n_n5008) & (!n_n801) & (!x405x)) + ((n_n5007) & (n_n5008) & (!n_n801) & (x405x)) + ((n_n5007) & (n_n5008) & (n_n801) & (!x405x)) + ((n_n5007) & (n_n5008) & (n_n801) & (x405x)));
	assign x12354x = (((!n_n5241) & (!n_n5242) & (!n_n5246) & (!n_n5243) & (n_n5235)) + ((!n_n5241) & (!n_n5242) & (!n_n5246) & (n_n5243) & (!n_n5235)) + ((!n_n5241) & (!n_n5242) & (!n_n5246) & (n_n5243) & (n_n5235)) + ((!n_n5241) & (!n_n5242) & (n_n5246) & (!n_n5243) & (!n_n5235)) + ((!n_n5241) & (!n_n5242) & (n_n5246) & (!n_n5243) & (n_n5235)) + ((!n_n5241) & (!n_n5242) & (n_n5246) & (n_n5243) & (!n_n5235)) + ((!n_n5241) & (!n_n5242) & (n_n5246) & (n_n5243) & (n_n5235)) + ((!n_n5241) & (n_n5242) & (!n_n5246) & (!n_n5243) & (!n_n5235)) + ((!n_n5241) & (n_n5242) & (!n_n5246) & (!n_n5243) & (n_n5235)) + ((!n_n5241) & (n_n5242) & (!n_n5246) & (n_n5243) & (!n_n5235)) + ((!n_n5241) & (n_n5242) & (!n_n5246) & (n_n5243) & (n_n5235)) + ((!n_n5241) & (n_n5242) & (n_n5246) & (!n_n5243) & (!n_n5235)) + ((!n_n5241) & (n_n5242) & (n_n5246) & (!n_n5243) & (n_n5235)) + ((!n_n5241) & (n_n5242) & (n_n5246) & (n_n5243) & (!n_n5235)) + ((!n_n5241) & (n_n5242) & (n_n5246) & (n_n5243) & (n_n5235)) + ((n_n5241) & (!n_n5242) & (!n_n5246) & (!n_n5243) & (!n_n5235)) + ((n_n5241) & (!n_n5242) & (!n_n5246) & (!n_n5243) & (n_n5235)) + ((n_n5241) & (!n_n5242) & (!n_n5246) & (n_n5243) & (!n_n5235)) + ((n_n5241) & (!n_n5242) & (!n_n5246) & (n_n5243) & (n_n5235)) + ((n_n5241) & (!n_n5242) & (n_n5246) & (!n_n5243) & (!n_n5235)) + ((n_n5241) & (!n_n5242) & (n_n5246) & (!n_n5243) & (n_n5235)) + ((n_n5241) & (!n_n5242) & (n_n5246) & (n_n5243) & (!n_n5235)) + ((n_n5241) & (!n_n5242) & (n_n5246) & (n_n5243) & (n_n5235)) + ((n_n5241) & (n_n5242) & (!n_n5246) & (!n_n5243) & (!n_n5235)) + ((n_n5241) & (n_n5242) & (!n_n5246) & (!n_n5243) & (n_n5235)) + ((n_n5241) & (n_n5242) & (!n_n5246) & (n_n5243) & (!n_n5235)) + ((n_n5241) & (n_n5242) & (!n_n5246) & (n_n5243) & (n_n5235)) + ((n_n5241) & (n_n5242) & (n_n5246) & (!n_n5243) & (!n_n5235)) + ((n_n5241) & (n_n5242) & (n_n5246) & (!n_n5243) & (n_n5235)) + ((n_n5241) & (n_n5242) & (n_n5246) & (n_n5243) & (!n_n5235)) + ((n_n5241) & (n_n5242) & (n_n5246) & (n_n5243) & (n_n5235)));
	assign n_n1436 = (((!n_n5239) & (!n_n5240) & (!n_n5245) & (!n_n5237) & (x12354x)) + ((!n_n5239) & (!n_n5240) & (!n_n5245) & (n_n5237) & (!x12354x)) + ((!n_n5239) & (!n_n5240) & (!n_n5245) & (n_n5237) & (x12354x)) + ((!n_n5239) & (!n_n5240) & (n_n5245) & (!n_n5237) & (!x12354x)) + ((!n_n5239) & (!n_n5240) & (n_n5245) & (!n_n5237) & (x12354x)) + ((!n_n5239) & (!n_n5240) & (n_n5245) & (n_n5237) & (!x12354x)) + ((!n_n5239) & (!n_n5240) & (n_n5245) & (n_n5237) & (x12354x)) + ((!n_n5239) & (n_n5240) & (!n_n5245) & (!n_n5237) & (!x12354x)) + ((!n_n5239) & (n_n5240) & (!n_n5245) & (!n_n5237) & (x12354x)) + ((!n_n5239) & (n_n5240) & (!n_n5245) & (n_n5237) & (!x12354x)) + ((!n_n5239) & (n_n5240) & (!n_n5245) & (n_n5237) & (x12354x)) + ((!n_n5239) & (n_n5240) & (n_n5245) & (!n_n5237) & (!x12354x)) + ((!n_n5239) & (n_n5240) & (n_n5245) & (!n_n5237) & (x12354x)) + ((!n_n5239) & (n_n5240) & (n_n5245) & (n_n5237) & (!x12354x)) + ((!n_n5239) & (n_n5240) & (n_n5245) & (n_n5237) & (x12354x)) + ((n_n5239) & (!n_n5240) & (!n_n5245) & (!n_n5237) & (!x12354x)) + ((n_n5239) & (!n_n5240) & (!n_n5245) & (!n_n5237) & (x12354x)) + ((n_n5239) & (!n_n5240) & (!n_n5245) & (n_n5237) & (!x12354x)) + ((n_n5239) & (!n_n5240) & (!n_n5245) & (n_n5237) & (x12354x)) + ((n_n5239) & (!n_n5240) & (n_n5245) & (!n_n5237) & (!x12354x)) + ((n_n5239) & (!n_n5240) & (n_n5245) & (!n_n5237) & (x12354x)) + ((n_n5239) & (!n_n5240) & (n_n5245) & (n_n5237) & (!x12354x)) + ((n_n5239) & (!n_n5240) & (n_n5245) & (n_n5237) & (x12354x)) + ((n_n5239) & (n_n5240) & (!n_n5245) & (!n_n5237) & (!x12354x)) + ((n_n5239) & (n_n5240) & (!n_n5245) & (!n_n5237) & (x12354x)) + ((n_n5239) & (n_n5240) & (!n_n5245) & (n_n5237) & (!x12354x)) + ((n_n5239) & (n_n5240) & (!n_n5245) & (n_n5237) & (x12354x)) + ((n_n5239) & (n_n5240) & (n_n5245) & (!n_n5237) & (!x12354x)) + ((n_n5239) & (n_n5240) & (n_n5245) & (!n_n5237) & (x12354x)) + ((n_n5239) & (n_n5240) & (n_n5245) & (n_n5237) & (!x12354x)) + ((n_n5239) & (n_n5240) & (n_n5245) & (n_n5237) & (x12354x)));
	assign x225x = (((!i_9_) & (n_n390) & (n_n473) & (n_n534)) + ((i_9_) & (n_n390) & (n_n473) & (n_n534)));
	assign x432x = (((!n_n4661) & (!n_n4660) & (!n_n4663) & (x225x)) + ((!n_n4661) & (!n_n4660) & (n_n4663) & (!x225x)) + ((!n_n4661) & (!n_n4660) & (n_n4663) & (x225x)) + ((!n_n4661) & (n_n4660) & (!n_n4663) & (!x225x)) + ((!n_n4661) & (n_n4660) & (!n_n4663) & (x225x)) + ((!n_n4661) & (n_n4660) & (n_n4663) & (!x225x)) + ((!n_n4661) & (n_n4660) & (n_n4663) & (x225x)) + ((n_n4661) & (!n_n4660) & (!n_n4663) & (!x225x)) + ((n_n4661) & (!n_n4660) & (!n_n4663) & (x225x)) + ((n_n4661) & (!n_n4660) & (n_n4663) & (!x225x)) + ((n_n4661) & (!n_n4660) & (n_n4663) & (x225x)) + ((n_n4661) & (n_n4660) & (!n_n4663) & (!x225x)) + ((n_n4661) & (n_n4660) & (!n_n4663) & (x225x)) + ((n_n4661) & (n_n4660) & (n_n4663) & (!x225x)) + ((n_n4661) & (n_n4660) & (n_n4663) & (x225x)));
	assign x11859x = (((!n_n4669) & (!n_n4673) & (!n_n4668) & (n_n4662)) + ((!n_n4669) & (!n_n4673) & (n_n4668) & (!n_n4662)) + ((!n_n4669) & (!n_n4673) & (n_n4668) & (n_n4662)) + ((!n_n4669) & (n_n4673) & (!n_n4668) & (!n_n4662)) + ((!n_n4669) & (n_n4673) & (!n_n4668) & (n_n4662)) + ((!n_n4669) & (n_n4673) & (n_n4668) & (!n_n4662)) + ((!n_n4669) & (n_n4673) & (n_n4668) & (n_n4662)) + ((n_n4669) & (!n_n4673) & (!n_n4668) & (!n_n4662)) + ((n_n4669) & (!n_n4673) & (!n_n4668) & (n_n4662)) + ((n_n4669) & (!n_n4673) & (n_n4668) & (!n_n4662)) + ((n_n4669) & (!n_n4673) & (n_n4668) & (n_n4662)) + ((n_n4669) & (n_n4673) & (!n_n4668) & (!n_n4662)) + ((n_n4669) & (n_n4673) & (!n_n4668) & (n_n4662)) + ((n_n4669) & (n_n4673) & (n_n4668) & (!n_n4662)) + ((n_n4669) & (n_n4673) & (n_n4668) & (n_n4662)));
	assign x22154x = (((!n_n5038) & (!n_n5034) & (!n_n5035) & (!n_n5036)));
	assign x12003x = (((!n_n5041) & (!n_n5043) & (!n_n5039) & (!x253x) & (!x22154x)) + ((!n_n5041) & (!n_n5043) & (!n_n5039) & (x253x) & (!x22154x)) + ((!n_n5041) & (!n_n5043) & (!n_n5039) & (x253x) & (x22154x)) + ((!n_n5041) & (!n_n5043) & (n_n5039) & (!x253x) & (!x22154x)) + ((!n_n5041) & (!n_n5043) & (n_n5039) & (!x253x) & (x22154x)) + ((!n_n5041) & (!n_n5043) & (n_n5039) & (x253x) & (!x22154x)) + ((!n_n5041) & (!n_n5043) & (n_n5039) & (x253x) & (x22154x)) + ((!n_n5041) & (n_n5043) & (!n_n5039) & (!x253x) & (!x22154x)) + ((!n_n5041) & (n_n5043) & (!n_n5039) & (!x253x) & (x22154x)) + ((!n_n5041) & (n_n5043) & (!n_n5039) & (x253x) & (!x22154x)) + ((!n_n5041) & (n_n5043) & (!n_n5039) & (x253x) & (x22154x)) + ((!n_n5041) & (n_n5043) & (n_n5039) & (!x253x) & (!x22154x)) + ((!n_n5041) & (n_n5043) & (n_n5039) & (!x253x) & (x22154x)) + ((!n_n5041) & (n_n5043) & (n_n5039) & (x253x) & (!x22154x)) + ((!n_n5041) & (n_n5043) & (n_n5039) & (x253x) & (x22154x)) + ((n_n5041) & (!n_n5043) & (!n_n5039) & (!x253x) & (!x22154x)) + ((n_n5041) & (!n_n5043) & (!n_n5039) & (!x253x) & (x22154x)) + ((n_n5041) & (!n_n5043) & (!n_n5039) & (x253x) & (!x22154x)) + ((n_n5041) & (!n_n5043) & (!n_n5039) & (x253x) & (x22154x)) + ((n_n5041) & (!n_n5043) & (n_n5039) & (!x253x) & (!x22154x)) + ((n_n5041) & (!n_n5043) & (n_n5039) & (!x253x) & (x22154x)) + ((n_n5041) & (!n_n5043) & (n_n5039) & (x253x) & (!x22154x)) + ((n_n5041) & (!n_n5043) & (n_n5039) & (x253x) & (x22154x)) + ((n_n5041) & (n_n5043) & (!n_n5039) & (!x253x) & (!x22154x)) + ((n_n5041) & (n_n5043) & (!n_n5039) & (!x253x) & (x22154x)) + ((n_n5041) & (n_n5043) & (!n_n5039) & (x253x) & (!x22154x)) + ((n_n5041) & (n_n5043) & (!n_n5039) & (x253x) & (x22154x)) + ((n_n5041) & (n_n5043) & (n_n5039) & (!x253x) & (!x22154x)) + ((n_n5041) & (n_n5043) & (n_n5039) & (!x253x) & (x22154x)) + ((n_n5041) & (n_n5043) & (n_n5039) & (x253x) & (!x22154x)) + ((n_n5041) & (n_n5043) & (n_n5039) & (x253x) & (x22154x)));
	assign n_n1023 = (((!n_n1064) & (!n_n1066) & (x12003x)) + ((!n_n1064) & (n_n1066) & (!x12003x)) + ((!n_n1064) & (n_n1066) & (x12003x)) + ((n_n1064) & (!n_n1066) & (!x12003x)) + ((n_n1064) & (!n_n1066) & (x12003x)) + ((n_n1064) & (n_n1066) & (!x12003x)) + ((n_n1064) & (n_n1066) & (x12003x)));
	assign x22194x = (((!n_n5096) & (!n_n5099) & (!n_n5098) & (!n_n5105) & (!n_n1167)));
	assign n_n1061 = (((!n_n518) & (!x21x) & (!n_n130) & (!x20x) & (!x22194x)) + ((!n_n518) & (!x21x) & (!n_n130) & (x20x) & (!x22194x)) + ((!n_n518) & (!x21x) & (n_n130) & (!x20x) & (!x22194x)) + ((!n_n518) & (!x21x) & (n_n130) & (x20x) & (!x22194x)) + ((!n_n518) & (x21x) & (!n_n130) & (!x20x) & (!x22194x)) + ((!n_n518) & (x21x) & (!n_n130) & (x20x) & (!x22194x)) + ((!n_n518) & (x21x) & (n_n130) & (!x20x) & (!x22194x)) + ((!n_n518) & (x21x) & (n_n130) & (x20x) & (!x22194x)) + ((n_n518) & (!x21x) & (!n_n130) & (!x20x) & (!x22194x)) + ((n_n518) & (!x21x) & (!n_n130) & (x20x) & (!x22194x)) + ((n_n518) & (!x21x) & (n_n130) & (!x20x) & (!x22194x)) + ((n_n518) & (!x21x) & (n_n130) & (x20x) & (!x22194x)) + ((n_n518) & (!x21x) & (n_n130) & (x20x) & (x22194x)) + ((n_n518) & (x21x) & (!n_n130) & (!x20x) & (!x22194x)) + ((n_n518) & (x21x) & (!n_n130) & (x20x) & (!x22194x)) + ((n_n518) & (x21x) & (n_n130) & (!x20x) & (!x22194x)) + ((n_n518) & (x21x) & (n_n130) & (!x20x) & (x22194x)) + ((n_n518) & (x21x) & (n_n130) & (x20x) & (!x22194x)) + ((n_n518) & (x21x) & (n_n130) & (x20x) & (x22194x)));
	assign x22153x = (((!n_n5091) & (!n_n5089) & (!n_n5095) & (!n_n5084) & (!n_n5090)));
	assign n_n1062 = (((!n_n5081) & (!n_n5082) & (!n_n5078) & (!n_n5083) & (!x22153x)) + ((!n_n5081) & (!n_n5082) & (!n_n5078) & (n_n5083) & (!x22153x)) + ((!n_n5081) & (!n_n5082) & (!n_n5078) & (n_n5083) & (x22153x)) + ((!n_n5081) & (!n_n5082) & (n_n5078) & (!n_n5083) & (!x22153x)) + ((!n_n5081) & (!n_n5082) & (n_n5078) & (!n_n5083) & (x22153x)) + ((!n_n5081) & (!n_n5082) & (n_n5078) & (n_n5083) & (!x22153x)) + ((!n_n5081) & (!n_n5082) & (n_n5078) & (n_n5083) & (x22153x)) + ((!n_n5081) & (n_n5082) & (!n_n5078) & (!n_n5083) & (!x22153x)) + ((!n_n5081) & (n_n5082) & (!n_n5078) & (!n_n5083) & (x22153x)) + ((!n_n5081) & (n_n5082) & (!n_n5078) & (n_n5083) & (!x22153x)) + ((!n_n5081) & (n_n5082) & (!n_n5078) & (n_n5083) & (x22153x)) + ((!n_n5081) & (n_n5082) & (n_n5078) & (!n_n5083) & (!x22153x)) + ((!n_n5081) & (n_n5082) & (n_n5078) & (!n_n5083) & (x22153x)) + ((!n_n5081) & (n_n5082) & (n_n5078) & (n_n5083) & (!x22153x)) + ((!n_n5081) & (n_n5082) & (n_n5078) & (n_n5083) & (x22153x)) + ((n_n5081) & (!n_n5082) & (!n_n5078) & (!n_n5083) & (!x22153x)) + ((n_n5081) & (!n_n5082) & (!n_n5078) & (!n_n5083) & (x22153x)) + ((n_n5081) & (!n_n5082) & (!n_n5078) & (n_n5083) & (!x22153x)) + ((n_n5081) & (!n_n5082) & (!n_n5078) & (n_n5083) & (x22153x)) + ((n_n5081) & (!n_n5082) & (n_n5078) & (!n_n5083) & (!x22153x)) + ((n_n5081) & (!n_n5082) & (n_n5078) & (!n_n5083) & (x22153x)) + ((n_n5081) & (!n_n5082) & (n_n5078) & (n_n5083) & (!x22153x)) + ((n_n5081) & (!n_n5082) & (n_n5078) & (n_n5083) & (x22153x)) + ((n_n5081) & (n_n5082) & (!n_n5078) & (!n_n5083) & (!x22153x)) + ((n_n5081) & (n_n5082) & (!n_n5078) & (!n_n5083) & (x22153x)) + ((n_n5081) & (n_n5082) & (!n_n5078) & (n_n5083) & (!x22153x)) + ((n_n5081) & (n_n5082) & (!n_n5078) & (n_n5083) & (x22153x)) + ((n_n5081) & (n_n5082) & (n_n5078) & (!n_n5083) & (!x22153x)) + ((n_n5081) & (n_n5082) & (n_n5078) & (!n_n5083) & (x22153x)) + ((n_n5081) & (n_n5082) & (n_n5078) & (n_n5083) & (!x22153x)) + ((n_n5081) & (n_n5082) & (n_n5078) & (n_n5083) & (x22153x)));
	assign x12019x = (((!n_n532) & (!x18x) & (!n_n464) & (!n_n5069) & (n_n4152)) + ((!n_n532) & (!x18x) & (!n_n464) & (n_n5069) & (!n_n4152)) + ((!n_n532) & (!x18x) & (!n_n464) & (n_n5069) & (n_n4152)) + ((!n_n532) & (!x18x) & (n_n464) & (!n_n5069) & (n_n4152)) + ((!n_n532) & (!x18x) & (n_n464) & (n_n5069) & (!n_n4152)) + ((!n_n532) & (!x18x) & (n_n464) & (n_n5069) & (n_n4152)) + ((!n_n532) & (x18x) & (!n_n464) & (!n_n5069) & (n_n4152)) + ((!n_n532) & (x18x) & (!n_n464) & (n_n5069) & (!n_n4152)) + ((!n_n532) & (x18x) & (!n_n464) & (n_n5069) & (n_n4152)) + ((!n_n532) & (x18x) & (n_n464) & (!n_n5069) & (n_n4152)) + ((!n_n532) & (x18x) & (n_n464) & (n_n5069) & (!n_n4152)) + ((!n_n532) & (x18x) & (n_n464) & (n_n5069) & (n_n4152)) + ((n_n532) & (!x18x) & (!n_n464) & (!n_n5069) & (n_n4152)) + ((n_n532) & (!x18x) & (!n_n464) & (n_n5069) & (!n_n4152)) + ((n_n532) & (!x18x) & (!n_n464) & (n_n5069) & (n_n4152)) + ((n_n532) & (!x18x) & (n_n464) & (!n_n5069) & (n_n4152)) + ((n_n532) & (!x18x) & (n_n464) & (n_n5069) & (!n_n4152)) + ((n_n532) & (!x18x) & (n_n464) & (n_n5069) & (n_n4152)) + ((n_n532) & (x18x) & (!n_n464) & (!n_n5069) & (n_n4152)) + ((n_n532) & (x18x) & (!n_n464) & (n_n5069) & (!n_n4152)) + ((n_n532) & (x18x) & (!n_n464) & (n_n5069) & (n_n4152)) + ((n_n532) & (x18x) & (n_n464) & (!n_n5069) & (!n_n4152)) + ((n_n532) & (x18x) & (n_n464) & (!n_n5069) & (n_n4152)) + ((n_n532) & (x18x) & (n_n464) & (n_n5069) & (!n_n4152)) + ((n_n532) & (x18x) & (n_n464) & (n_n5069) & (n_n4152)));
	assign x12020x = (((!n_n5060) & (!x120x) & (!n_n5067) & (x12019x)) + ((!n_n5060) & (!x120x) & (n_n5067) & (!x12019x)) + ((!n_n5060) & (!x120x) & (n_n5067) & (x12019x)) + ((!n_n5060) & (x120x) & (!n_n5067) & (!x12019x)) + ((!n_n5060) & (x120x) & (!n_n5067) & (x12019x)) + ((!n_n5060) & (x120x) & (n_n5067) & (!x12019x)) + ((!n_n5060) & (x120x) & (n_n5067) & (x12019x)) + ((n_n5060) & (!x120x) & (!n_n5067) & (!x12019x)) + ((n_n5060) & (!x120x) & (!n_n5067) & (x12019x)) + ((n_n5060) & (!x120x) & (n_n5067) & (!x12019x)) + ((n_n5060) & (!x120x) & (n_n5067) & (x12019x)) + ((n_n5060) & (x120x) & (!n_n5067) & (!x12019x)) + ((n_n5060) & (x120x) & (!n_n5067) & (x12019x)) + ((n_n5060) & (x120x) & (n_n5067) & (!x12019x)) + ((n_n5060) & (x120x) & (n_n5067) & (x12019x)));
	assign x104x = (((!i_9_) & (n_n526) & (n_n509) & (n_n195)) + ((i_9_) & (n_n526) & (n_n509) & (n_n195)));
	assign x12025x = (((!n_n4990) & (!n_n4982) & (!n_n4983) & (!n_n4985) & (n_n4984)) + ((!n_n4990) & (!n_n4982) & (!n_n4983) & (n_n4985) & (!n_n4984)) + ((!n_n4990) & (!n_n4982) & (!n_n4983) & (n_n4985) & (n_n4984)) + ((!n_n4990) & (!n_n4982) & (n_n4983) & (!n_n4985) & (!n_n4984)) + ((!n_n4990) & (!n_n4982) & (n_n4983) & (!n_n4985) & (n_n4984)) + ((!n_n4990) & (!n_n4982) & (n_n4983) & (n_n4985) & (!n_n4984)) + ((!n_n4990) & (!n_n4982) & (n_n4983) & (n_n4985) & (n_n4984)) + ((!n_n4990) & (n_n4982) & (!n_n4983) & (!n_n4985) & (!n_n4984)) + ((!n_n4990) & (n_n4982) & (!n_n4983) & (!n_n4985) & (n_n4984)) + ((!n_n4990) & (n_n4982) & (!n_n4983) & (n_n4985) & (!n_n4984)) + ((!n_n4990) & (n_n4982) & (!n_n4983) & (n_n4985) & (n_n4984)) + ((!n_n4990) & (n_n4982) & (n_n4983) & (!n_n4985) & (!n_n4984)) + ((!n_n4990) & (n_n4982) & (n_n4983) & (!n_n4985) & (n_n4984)) + ((!n_n4990) & (n_n4982) & (n_n4983) & (n_n4985) & (!n_n4984)) + ((!n_n4990) & (n_n4982) & (n_n4983) & (n_n4985) & (n_n4984)) + ((n_n4990) & (!n_n4982) & (!n_n4983) & (!n_n4985) & (!n_n4984)) + ((n_n4990) & (!n_n4982) & (!n_n4983) & (!n_n4985) & (n_n4984)) + ((n_n4990) & (!n_n4982) & (!n_n4983) & (n_n4985) & (!n_n4984)) + ((n_n4990) & (!n_n4982) & (!n_n4983) & (n_n4985) & (n_n4984)) + ((n_n4990) & (!n_n4982) & (n_n4983) & (!n_n4985) & (!n_n4984)) + ((n_n4990) & (!n_n4982) & (n_n4983) & (!n_n4985) & (n_n4984)) + ((n_n4990) & (!n_n4982) & (n_n4983) & (n_n4985) & (!n_n4984)) + ((n_n4990) & (!n_n4982) & (n_n4983) & (n_n4985) & (n_n4984)) + ((n_n4990) & (n_n4982) & (!n_n4983) & (!n_n4985) & (!n_n4984)) + ((n_n4990) & (n_n4982) & (!n_n4983) & (!n_n4985) & (n_n4984)) + ((n_n4990) & (n_n4982) & (!n_n4983) & (n_n4985) & (!n_n4984)) + ((n_n4990) & (n_n4982) & (!n_n4983) & (n_n4985) & (n_n4984)) + ((n_n4990) & (n_n4982) & (n_n4983) & (!n_n4985) & (!n_n4984)) + ((n_n4990) & (n_n4982) & (n_n4983) & (!n_n4985) & (n_n4984)) + ((n_n4990) & (n_n4982) & (n_n4983) & (n_n4985) & (!n_n4984)) + ((n_n4990) & (n_n4982) & (n_n4983) & (n_n4985) & (n_n4984)));
	assign x12028x = (((!n_n1068) & (!x133x) & (!n_n1067) & (!x104x) & (x12025x)) + ((!n_n1068) & (!x133x) & (!n_n1067) & (x104x) & (!x12025x)) + ((!n_n1068) & (!x133x) & (!n_n1067) & (x104x) & (x12025x)) + ((!n_n1068) & (!x133x) & (n_n1067) & (!x104x) & (!x12025x)) + ((!n_n1068) & (!x133x) & (n_n1067) & (!x104x) & (x12025x)) + ((!n_n1068) & (!x133x) & (n_n1067) & (x104x) & (!x12025x)) + ((!n_n1068) & (!x133x) & (n_n1067) & (x104x) & (x12025x)) + ((!n_n1068) & (x133x) & (!n_n1067) & (!x104x) & (!x12025x)) + ((!n_n1068) & (x133x) & (!n_n1067) & (!x104x) & (x12025x)) + ((!n_n1068) & (x133x) & (!n_n1067) & (x104x) & (!x12025x)) + ((!n_n1068) & (x133x) & (!n_n1067) & (x104x) & (x12025x)) + ((!n_n1068) & (x133x) & (n_n1067) & (!x104x) & (!x12025x)) + ((!n_n1068) & (x133x) & (n_n1067) & (!x104x) & (x12025x)) + ((!n_n1068) & (x133x) & (n_n1067) & (x104x) & (!x12025x)) + ((!n_n1068) & (x133x) & (n_n1067) & (x104x) & (x12025x)) + ((n_n1068) & (!x133x) & (!n_n1067) & (!x104x) & (!x12025x)) + ((n_n1068) & (!x133x) & (!n_n1067) & (!x104x) & (x12025x)) + ((n_n1068) & (!x133x) & (!n_n1067) & (x104x) & (!x12025x)) + ((n_n1068) & (!x133x) & (!n_n1067) & (x104x) & (x12025x)) + ((n_n1068) & (!x133x) & (n_n1067) & (!x104x) & (!x12025x)) + ((n_n1068) & (!x133x) & (n_n1067) & (!x104x) & (x12025x)) + ((n_n1068) & (!x133x) & (n_n1067) & (x104x) & (!x12025x)) + ((n_n1068) & (!x133x) & (n_n1067) & (x104x) & (x12025x)) + ((n_n1068) & (x133x) & (!n_n1067) & (!x104x) & (!x12025x)) + ((n_n1068) & (x133x) & (!n_n1067) & (!x104x) & (x12025x)) + ((n_n1068) & (x133x) & (!n_n1067) & (x104x) & (!x12025x)) + ((n_n1068) & (x133x) & (!n_n1067) & (x104x) & (x12025x)) + ((n_n1068) & (x133x) & (n_n1067) & (!x104x) & (!x12025x)) + ((n_n1068) & (x133x) & (n_n1067) & (!x104x) & (x12025x)) + ((n_n1068) & (x133x) & (n_n1067) & (x104x) & (!x12025x)) + ((n_n1068) & (x133x) & (n_n1067) & (x104x) & (x12025x)));
	assign n_n4323 = (((!i_9_) & (n_n536) & (n_n524) & (n_n535)));
	assign x13003x = (((!i_7_) & (i_8_) & (!i_6_) & (x13x) & (n_n535)) + ((i_7_) & (i_8_) & (!i_6_) & (x13x) & (n_n535)));
	assign n_n727 = (((!n_n4447) & (!x368x) & (!x32x) & (!x128x) & (x13003x)) + ((!n_n4447) & (!x368x) & (!x32x) & (x128x) & (!x13003x)) + ((!n_n4447) & (!x368x) & (!x32x) & (x128x) & (x13003x)) + ((!n_n4447) & (!x368x) & (x32x) & (!x128x) & (!x13003x)) + ((!n_n4447) & (!x368x) & (x32x) & (!x128x) & (x13003x)) + ((!n_n4447) & (!x368x) & (x32x) & (x128x) & (!x13003x)) + ((!n_n4447) & (!x368x) & (x32x) & (x128x) & (x13003x)) + ((!n_n4447) & (x368x) & (!x32x) & (!x128x) & (!x13003x)) + ((!n_n4447) & (x368x) & (!x32x) & (!x128x) & (x13003x)) + ((!n_n4447) & (x368x) & (!x32x) & (x128x) & (!x13003x)) + ((!n_n4447) & (x368x) & (!x32x) & (x128x) & (x13003x)) + ((!n_n4447) & (x368x) & (x32x) & (!x128x) & (!x13003x)) + ((!n_n4447) & (x368x) & (x32x) & (!x128x) & (x13003x)) + ((!n_n4447) & (x368x) & (x32x) & (x128x) & (!x13003x)) + ((!n_n4447) & (x368x) & (x32x) & (x128x) & (x13003x)) + ((n_n4447) & (!x368x) & (!x32x) & (!x128x) & (!x13003x)) + ((n_n4447) & (!x368x) & (!x32x) & (!x128x) & (x13003x)) + ((n_n4447) & (!x368x) & (!x32x) & (x128x) & (!x13003x)) + ((n_n4447) & (!x368x) & (!x32x) & (x128x) & (x13003x)) + ((n_n4447) & (!x368x) & (x32x) & (!x128x) & (!x13003x)) + ((n_n4447) & (!x368x) & (x32x) & (!x128x) & (x13003x)) + ((n_n4447) & (!x368x) & (x32x) & (x128x) & (!x13003x)) + ((n_n4447) & (!x368x) & (x32x) & (x128x) & (x13003x)) + ((n_n4447) & (x368x) & (!x32x) & (!x128x) & (!x13003x)) + ((n_n4447) & (x368x) & (!x32x) & (!x128x) & (x13003x)) + ((n_n4447) & (x368x) & (!x32x) & (x128x) & (!x13003x)) + ((n_n4447) & (x368x) & (!x32x) & (x128x) & (x13003x)) + ((n_n4447) & (x368x) & (x32x) & (!x128x) & (!x13003x)) + ((n_n4447) & (x368x) & (x32x) & (!x128x) & (x13003x)) + ((n_n4447) & (x368x) & (x32x) & (x128x) & (!x13003x)) + ((n_n4447) & (x368x) & (x32x) & (x128x) & (x13003x)));
	assign n_n910 = (((!i_9_) & (n_n536) & (!n_n524) & (n_n526) & (n_n464)) + ((!i_9_) & (n_n536) & (n_n524) & (!n_n526) & (n_n464)) + ((!i_9_) & (n_n536) & (n_n524) & (n_n526) & (n_n464)) + ((i_9_) & (n_n536) & (n_n524) & (!n_n526) & (n_n464)) + ((i_9_) & (n_n536) & (n_n524) & (n_n526) & (n_n464)));
	assign x13010x = (((!i_9_) & (n_n536) & (n_n532) & (!n_n530) & (n_n464)) + ((!i_9_) & (n_n536) & (n_n532) & (n_n530) & (n_n464)) + ((i_9_) & (n_n536) & (!n_n532) & (n_n530) & (n_n464)) + ((i_9_) & (n_n536) & (n_n532) & (n_n530) & (n_n464)));
	assign x13016x = (((!n_n4436) & (!n_n4443) & (!n_n2803) & (!n_n910) & (x13010x)) + ((!n_n4436) & (!n_n4443) & (!n_n2803) & (n_n910) & (!x13010x)) + ((!n_n4436) & (!n_n4443) & (!n_n2803) & (n_n910) & (x13010x)) + ((!n_n4436) & (!n_n4443) & (n_n2803) & (!n_n910) & (!x13010x)) + ((!n_n4436) & (!n_n4443) & (n_n2803) & (!n_n910) & (x13010x)) + ((!n_n4436) & (!n_n4443) & (n_n2803) & (n_n910) & (!x13010x)) + ((!n_n4436) & (!n_n4443) & (n_n2803) & (n_n910) & (x13010x)) + ((!n_n4436) & (n_n4443) & (!n_n2803) & (!n_n910) & (!x13010x)) + ((!n_n4436) & (n_n4443) & (!n_n2803) & (!n_n910) & (x13010x)) + ((!n_n4436) & (n_n4443) & (!n_n2803) & (n_n910) & (!x13010x)) + ((!n_n4436) & (n_n4443) & (!n_n2803) & (n_n910) & (x13010x)) + ((!n_n4436) & (n_n4443) & (n_n2803) & (!n_n910) & (!x13010x)) + ((!n_n4436) & (n_n4443) & (n_n2803) & (!n_n910) & (x13010x)) + ((!n_n4436) & (n_n4443) & (n_n2803) & (n_n910) & (!x13010x)) + ((!n_n4436) & (n_n4443) & (n_n2803) & (n_n910) & (x13010x)) + ((n_n4436) & (!n_n4443) & (!n_n2803) & (!n_n910) & (!x13010x)) + ((n_n4436) & (!n_n4443) & (!n_n2803) & (!n_n910) & (x13010x)) + ((n_n4436) & (!n_n4443) & (!n_n2803) & (n_n910) & (!x13010x)) + ((n_n4436) & (!n_n4443) & (!n_n2803) & (n_n910) & (x13010x)) + ((n_n4436) & (!n_n4443) & (n_n2803) & (!n_n910) & (!x13010x)) + ((n_n4436) & (!n_n4443) & (n_n2803) & (!n_n910) & (x13010x)) + ((n_n4436) & (!n_n4443) & (n_n2803) & (n_n910) & (!x13010x)) + ((n_n4436) & (!n_n4443) & (n_n2803) & (n_n910) & (x13010x)) + ((n_n4436) & (n_n4443) & (!n_n2803) & (!n_n910) & (!x13010x)) + ((n_n4436) & (n_n4443) & (!n_n2803) & (!n_n910) & (x13010x)) + ((n_n4436) & (n_n4443) & (!n_n2803) & (n_n910) & (!x13010x)) + ((n_n4436) & (n_n4443) & (!n_n2803) & (n_n910) & (x13010x)) + ((n_n4436) & (n_n4443) & (n_n2803) & (!n_n910) & (!x13010x)) + ((n_n4436) & (n_n4443) & (n_n2803) & (!n_n910) & (x13010x)) + ((n_n4436) & (n_n4443) & (n_n2803) & (n_n910) & (!x13010x)) + ((n_n4436) & (n_n4443) & (n_n2803) & (n_n910) & (x13010x)));
	assign x12729x = (((!n_n4869) & (!n_n4878) & (!n_n4879) & (n_n4876)) + ((!n_n4869) & (!n_n4878) & (n_n4879) & (!n_n4876)) + ((!n_n4869) & (!n_n4878) & (n_n4879) & (n_n4876)) + ((!n_n4869) & (n_n4878) & (!n_n4879) & (!n_n4876)) + ((!n_n4869) & (n_n4878) & (!n_n4879) & (n_n4876)) + ((!n_n4869) & (n_n4878) & (n_n4879) & (!n_n4876)) + ((!n_n4869) & (n_n4878) & (n_n4879) & (n_n4876)) + ((n_n4869) & (!n_n4878) & (!n_n4879) & (!n_n4876)) + ((n_n4869) & (!n_n4878) & (!n_n4879) & (n_n4876)) + ((n_n4869) & (!n_n4878) & (n_n4879) & (!n_n4876)) + ((n_n4869) & (!n_n4878) & (n_n4879) & (n_n4876)) + ((n_n4869) & (n_n4878) & (!n_n4879) & (!n_n4876)) + ((n_n4869) & (n_n4878) & (!n_n4879) & (n_n4876)) + ((n_n4869) & (n_n4878) & (n_n4879) & (!n_n4876)) + ((n_n4869) & (n_n4878) & (n_n4879) & (n_n4876)));
	assign x12730x = (((!x295x) & (!n_n4875) & (!n_n4871) & (n_n4874)) + ((!x295x) & (!n_n4875) & (n_n4871) & (!n_n4874)) + ((!x295x) & (!n_n4875) & (n_n4871) & (n_n4874)) + ((!x295x) & (n_n4875) & (!n_n4871) & (!n_n4874)) + ((!x295x) & (n_n4875) & (!n_n4871) & (n_n4874)) + ((!x295x) & (n_n4875) & (n_n4871) & (!n_n4874)) + ((!x295x) & (n_n4875) & (n_n4871) & (n_n4874)) + ((x295x) & (!n_n4875) & (!n_n4871) & (!n_n4874)) + ((x295x) & (!n_n4875) & (!n_n4871) & (n_n4874)) + ((x295x) & (!n_n4875) & (n_n4871) & (!n_n4874)) + ((x295x) & (!n_n4875) & (n_n4871) & (n_n4874)) + ((x295x) & (n_n4875) & (!n_n4871) & (!n_n4874)) + ((x295x) & (n_n4875) & (!n_n4871) & (n_n4874)) + ((x295x) & (n_n4875) & (n_n4871) & (!n_n4874)) + ((x295x) & (n_n4875) & (n_n4871) & (n_n4874)));
	assign x12736x = (((!n_n4863) & (!n_n4853) & (!n_n4861) & (!n_n4852) & (n_n4851)) + ((!n_n4863) & (!n_n4853) & (!n_n4861) & (n_n4852) & (!n_n4851)) + ((!n_n4863) & (!n_n4853) & (!n_n4861) & (n_n4852) & (n_n4851)) + ((!n_n4863) & (!n_n4853) & (n_n4861) & (!n_n4852) & (!n_n4851)) + ((!n_n4863) & (!n_n4853) & (n_n4861) & (!n_n4852) & (n_n4851)) + ((!n_n4863) & (!n_n4853) & (n_n4861) & (n_n4852) & (!n_n4851)) + ((!n_n4863) & (!n_n4853) & (n_n4861) & (n_n4852) & (n_n4851)) + ((!n_n4863) & (n_n4853) & (!n_n4861) & (!n_n4852) & (!n_n4851)) + ((!n_n4863) & (n_n4853) & (!n_n4861) & (!n_n4852) & (n_n4851)) + ((!n_n4863) & (n_n4853) & (!n_n4861) & (n_n4852) & (!n_n4851)) + ((!n_n4863) & (n_n4853) & (!n_n4861) & (n_n4852) & (n_n4851)) + ((!n_n4863) & (n_n4853) & (n_n4861) & (!n_n4852) & (!n_n4851)) + ((!n_n4863) & (n_n4853) & (n_n4861) & (!n_n4852) & (n_n4851)) + ((!n_n4863) & (n_n4853) & (n_n4861) & (n_n4852) & (!n_n4851)) + ((!n_n4863) & (n_n4853) & (n_n4861) & (n_n4852) & (n_n4851)) + ((n_n4863) & (!n_n4853) & (!n_n4861) & (!n_n4852) & (!n_n4851)) + ((n_n4863) & (!n_n4853) & (!n_n4861) & (!n_n4852) & (n_n4851)) + ((n_n4863) & (!n_n4853) & (!n_n4861) & (n_n4852) & (!n_n4851)) + ((n_n4863) & (!n_n4853) & (!n_n4861) & (n_n4852) & (n_n4851)) + ((n_n4863) & (!n_n4853) & (n_n4861) & (!n_n4852) & (!n_n4851)) + ((n_n4863) & (!n_n4853) & (n_n4861) & (!n_n4852) & (n_n4851)) + ((n_n4863) & (!n_n4853) & (n_n4861) & (n_n4852) & (!n_n4851)) + ((n_n4863) & (!n_n4853) & (n_n4861) & (n_n4852) & (n_n4851)) + ((n_n4863) & (n_n4853) & (!n_n4861) & (!n_n4852) & (!n_n4851)) + ((n_n4863) & (n_n4853) & (!n_n4861) & (!n_n4852) & (n_n4851)) + ((n_n4863) & (n_n4853) & (!n_n4861) & (n_n4852) & (!n_n4851)) + ((n_n4863) & (n_n4853) & (!n_n4861) & (n_n4852) & (n_n4851)) + ((n_n4863) & (n_n4853) & (n_n4861) & (!n_n4852) & (!n_n4851)) + ((n_n4863) & (n_n4853) & (n_n4861) & (!n_n4852) & (n_n4851)) + ((n_n4863) & (n_n4853) & (n_n4861) & (n_n4852) & (!n_n4851)) + ((n_n4863) & (n_n4853) & (n_n4861) & (n_n4852) & (n_n4851)));
	assign n_n696 = (((!n_n4857) & (!n_n4862) & (!n_n4860) & (!n_n4864) & (x12736x)) + ((!n_n4857) & (!n_n4862) & (!n_n4860) & (n_n4864) & (!x12736x)) + ((!n_n4857) & (!n_n4862) & (!n_n4860) & (n_n4864) & (x12736x)) + ((!n_n4857) & (!n_n4862) & (n_n4860) & (!n_n4864) & (!x12736x)) + ((!n_n4857) & (!n_n4862) & (n_n4860) & (!n_n4864) & (x12736x)) + ((!n_n4857) & (!n_n4862) & (n_n4860) & (n_n4864) & (!x12736x)) + ((!n_n4857) & (!n_n4862) & (n_n4860) & (n_n4864) & (x12736x)) + ((!n_n4857) & (n_n4862) & (!n_n4860) & (!n_n4864) & (!x12736x)) + ((!n_n4857) & (n_n4862) & (!n_n4860) & (!n_n4864) & (x12736x)) + ((!n_n4857) & (n_n4862) & (!n_n4860) & (n_n4864) & (!x12736x)) + ((!n_n4857) & (n_n4862) & (!n_n4860) & (n_n4864) & (x12736x)) + ((!n_n4857) & (n_n4862) & (n_n4860) & (!n_n4864) & (!x12736x)) + ((!n_n4857) & (n_n4862) & (n_n4860) & (!n_n4864) & (x12736x)) + ((!n_n4857) & (n_n4862) & (n_n4860) & (n_n4864) & (!x12736x)) + ((!n_n4857) & (n_n4862) & (n_n4860) & (n_n4864) & (x12736x)) + ((n_n4857) & (!n_n4862) & (!n_n4860) & (!n_n4864) & (!x12736x)) + ((n_n4857) & (!n_n4862) & (!n_n4860) & (!n_n4864) & (x12736x)) + ((n_n4857) & (!n_n4862) & (!n_n4860) & (n_n4864) & (!x12736x)) + ((n_n4857) & (!n_n4862) & (!n_n4860) & (n_n4864) & (x12736x)) + ((n_n4857) & (!n_n4862) & (n_n4860) & (!n_n4864) & (!x12736x)) + ((n_n4857) & (!n_n4862) & (n_n4860) & (!n_n4864) & (x12736x)) + ((n_n4857) & (!n_n4862) & (n_n4860) & (n_n4864) & (!x12736x)) + ((n_n4857) & (!n_n4862) & (n_n4860) & (n_n4864) & (x12736x)) + ((n_n4857) & (n_n4862) & (!n_n4860) & (!n_n4864) & (!x12736x)) + ((n_n4857) & (n_n4862) & (!n_n4860) & (!n_n4864) & (x12736x)) + ((n_n4857) & (n_n4862) & (!n_n4860) & (n_n4864) & (!x12736x)) + ((n_n4857) & (n_n4862) & (!n_n4860) & (n_n4864) & (x12736x)) + ((n_n4857) & (n_n4862) & (n_n4860) & (!n_n4864) & (!x12736x)) + ((n_n4857) & (n_n4862) & (n_n4860) & (!n_n4864) & (x12736x)) + ((n_n4857) & (n_n4862) & (n_n4860) & (n_n4864) & (!x12736x)) + ((n_n4857) & (n_n4862) & (n_n4860) & (n_n4864) & (x12736x)));
	assign x12597x = (((!n_n4597) & (!n_n4601) & (!n_n4631) & (!n_n4592) & (n_n4585)) + ((!n_n4597) & (!n_n4601) & (!n_n4631) & (n_n4592) & (!n_n4585)) + ((!n_n4597) & (!n_n4601) & (!n_n4631) & (n_n4592) & (n_n4585)) + ((!n_n4597) & (!n_n4601) & (n_n4631) & (!n_n4592) & (!n_n4585)) + ((!n_n4597) & (!n_n4601) & (n_n4631) & (!n_n4592) & (n_n4585)) + ((!n_n4597) & (!n_n4601) & (n_n4631) & (n_n4592) & (!n_n4585)) + ((!n_n4597) & (!n_n4601) & (n_n4631) & (n_n4592) & (n_n4585)) + ((!n_n4597) & (n_n4601) & (!n_n4631) & (!n_n4592) & (!n_n4585)) + ((!n_n4597) & (n_n4601) & (!n_n4631) & (!n_n4592) & (n_n4585)) + ((!n_n4597) & (n_n4601) & (!n_n4631) & (n_n4592) & (!n_n4585)) + ((!n_n4597) & (n_n4601) & (!n_n4631) & (n_n4592) & (n_n4585)) + ((!n_n4597) & (n_n4601) & (n_n4631) & (!n_n4592) & (!n_n4585)) + ((!n_n4597) & (n_n4601) & (n_n4631) & (!n_n4592) & (n_n4585)) + ((!n_n4597) & (n_n4601) & (n_n4631) & (n_n4592) & (!n_n4585)) + ((!n_n4597) & (n_n4601) & (n_n4631) & (n_n4592) & (n_n4585)) + ((n_n4597) & (!n_n4601) & (!n_n4631) & (!n_n4592) & (!n_n4585)) + ((n_n4597) & (!n_n4601) & (!n_n4631) & (!n_n4592) & (n_n4585)) + ((n_n4597) & (!n_n4601) & (!n_n4631) & (n_n4592) & (!n_n4585)) + ((n_n4597) & (!n_n4601) & (!n_n4631) & (n_n4592) & (n_n4585)) + ((n_n4597) & (!n_n4601) & (n_n4631) & (!n_n4592) & (!n_n4585)) + ((n_n4597) & (!n_n4601) & (n_n4631) & (!n_n4592) & (n_n4585)) + ((n_n4597) & (!n_n4601) & (n_n4631) & (n_n4592) & (!n_n4585)) + ((n_n4597) & (!n_n4601) & (n_n4631) & (n_n4592) & (n_n4585)) + ((n_n4597) & (n_n4601) & (!n_n4631) & (!n_n4592) & (!n_n4585)) + ((n_n4597) & (n_n4601) & (!n_n4631) & (!n_n4592) & (n_n4585)) + ((n_n4597) & (n_n4601) & (!n_n4631) & (n_n4592) & (!n_n4585)) + ((n_n4597) & (n_n4601) & (!n_n4631) & (n_n4592) & (n_n4585)) + ((n_n4597) & (n_n4601) & (n_n4631) & (!n_n4592) & (!n_n4585)) + ((n_n4597) & (n_n4601) & (n_n4631) & (!n_n4592) & (n_n4585)) + ((n_n4597) & (n_n4601) & (n_n4631) & (n_n4592) & (!n_n4585)) + ((n_n4597) & (n_n4601) & (n_n4631) & (n_n4592) & (n_n4585)));
	assign x379x = (((!i_7_) & (i_8_) & (!i_6_) & (n_n482) & (x13x)) + ((i_7_) & (!i_8_) & (!i_6_) & (n_n482) & (x13x)));
	assign x15445x = (((!n_n482) & (!x13x) & (!n_n528) & (!n_n4533) & (x379x)) + ((!n_n482) & (!x13x) & (!n_n528) & (n_n4533) & (!x379x)) + ((!n_n482) & (!x13x) & (!n_n528) & (n_n4533) & (x379x)) + ((!n_n482) & (!x13x) & (n_n528) & (!n_n4533) & (x379x)) + ((!n_n482) & (!x13x) & (n_n528) & (n_n4533) & (!x379x)) + ((!n_n482) & (!x13x) & (n_n528) & (n_n4533) & (x379x)) + ((!n_n482) & (x13x) & (!n_n528) & (!n_n4533) & (x379x)) + ((!n_n482) & (x13x) & (!n_n528) & (n_n4533) & (!x379x)) + ((!n_n482) & (x13x) & (!n_n528) & (n_n4533) & (x379x)) + ((!n_n482) & (x13x) & (n_n528) & (!n_n4533) & (x379x)) + ((!n_n482) & (x13x) & (n_n528) & (n_n4533) & (!x379x)) + ((!n_n482) & (x13x) & (n_n528) & (n_n4533) & (x379x)) + ((n_n482) & (!x13x) & (!n_n528) & (!n_n4533) & (x379x)) + ((n_n482) & (!x13x) & (!n_n528) & (n_n4533) & (!x379x)) + ((n_n482) & (!x13x) & (!n_n528) & (n_n4533) & (x379x)) + ((n_n482) & (!x13x) & (n_n528) & (!n_n4533) & (x379x)) + ((n_n482) & (!x13x) & (n_n528) & (n_n4533) & (!x379x)) + ((n_n482) & (!x13x) & (n_n528) & (n_n4533) & (x379x)) + ((n_n482) & (x13x) & (!n_n528) & (!n_n4533) & (x379x)) + ((n_n482) & (x13x) & (!n_n528) & (n_n4533) & (!x379x)) + ((n_n482) & (x13x) & (!n_n528) & (n_n4533) & (x379x)) + ((n_n482) & (x13x) & (n_n528) & (!n_n4533) & (!x379x)) + ((n_n482) & (x13x) & (n_n528) & (!n_n4533) & (x379x)) + ((n_n482) & (x13x) & (n_n528) & (n_n4533) & (!x379x)) + ((n_n482) & (x13x) & (n_n528) & (n_n4533) & (x379x)));
	assign x15446x = (((!n_n4524) & (!n_n4535) & (!n_n4536) & (!n_n4537) & (n_n4529)) + ((!n_n4524) & (!n_n4535) & (!n_n4536) & (n_n4537) & (!n_n4529)) + ((!n_n4524) & (!n_n4535) & (!n_n4536) & (n_n4537) & (n_n4529)) + ((!n_n4524) & (!n_n4535) & (n_n4536) & (!n_n4537) & (!n_n4529)) + ((!n_n4524) & (!n_n4535) & (n_n4536) & (!n_n4537) & (n_n4529)) + ((!n_n4524) & (!n_n4535) & (n_n4536) & (n_n4537) & (!n_n4529)) + ((!n_n4524) & (!n_n4535) & (n_n4536) & (n_n4537) & (n_n4529)) + ((!n_n4524) & (n_n4535) & (!n_n4536) & (!n_n4537) & (!n_n4529)) + ((!n_n4524) & (n_n4535) & (!n_n4536) & (!n_n4537) & (n_n4529)) + ((!n_n4524) & (n_n4535) & (!n_n4536) & (n_n4537) & (!n_n4529)) + ((!n_n4524) & (n_n4535) & (!n_n4536) & (n_n4537) & (n_n4529)) + ((!n_n4524) & (n_n4535) & (n_n4536) & (!n_n4537) & (!n_n4529)) + ((!n_n4524) & (n_n4535) & (n_n4536) & (!n_n4537) & (n_n4529)) + ((!n_n4524) & (n_n4535) & (n_n4536) & (n_n4537) & (!n_n4529)) + ((!n_n4524) & (n_n4535) & (n_n4536) & (n_n4537) & (n_n4529)) + ((n_n4524) & (!n_n4535) & (!n_n4536) & (!n_n4537) & (!n_n4529)) + ((n_n4524) & (!n_n4535) & (!n_n4536) & (!n_n4537) & (n_n4529)) + ((n_n4524) & (!n_n4535) & (!n_n4536) & (n_n4537) & (!n_n4529)) + ((n_n4524) & (!n_n4535) & (!n_n4536) & (n_n4537) & (n_n4529)) + ((n_n4524) & (!n_n4535) & (n_n4536) & (!n_n4537) & (!n_n4529)) + ((n_n4524) & (!n_n4535) & (n_n4536) & (!n_n4537) & (n_n4529)) + ((n_n4524) & (!n_n4535) & (n_n4536) & (n_n4537) & (!n_n4529)) + ((n_n4524) & (!n_n4535) & (n_n4536) & (n_n4537) & (n_n4529)) + ((n_n4524) & (n_n4535) & (!n_n4536) & (!n_n4537) & (!n_n4529)) + ((n_n4524) & (n_n4535) & (!n_n4536) & (!n_n4537) & (n_n4529)) + ((n_n4524) & (n_n4535) & (!n_n4536) & (n_n4537) & (!n_n4529)) + ((n_n4524) & (n_n4535) & (!n_n4536) & (n_n4537) & (n_n4529)) + ((n_n4524) & (n_n4535) & (n_n4536) & (!n_n4537) & (!n_n4529)) + ((n_n4524) & (n_n4535) & (n_n4536) & (!n_n4537) & (n_n4529)) + ((n_n4524) & (n_n4535) & (n_n4536) & (n_n4537) & (!n_n4529)) + ((n_n4524) & (n_n4535) & (n_n4536) & (n_n4537) & (n_n4529)));
	assign x22096x = (((!n_n4651) & (!n_n4649) & (!n_n4652) & (!n_n4663)));
	assign x210x = (((!i_9_) & (!n_n526) & (n_n528) & (n_n535) & (n_n195)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n535) & (n_n195)) + ((i_9_) & (n_n526) & (!n_n528) & (n_n535) & (n_n195)) + ((i_9_) & (n_n526) & (n_n528) & (n_n535) & (n_n195)));
	assign x60x = (((!n_n482) & (!x23x) & (!n_n65) & (n_n5304)) + ((!n_n482) & (!x23x) & (n_n65) & (n_n5304)) + ((!n_n482) & (x23x) & (!n_n65) & (n_n5304)) + ((!n_n482) & (x23x) & (n_n65) & (n_n5304)) + ((n_n482) & (!x23x) & (!n_n65) & (n_n5304)) + ((n_n482) & (!x23x) & (n_n65) & (n_n5304)) + ((n_n482) & (x23x) & (!n_n65) & (n_n5304)) + ((n_n482) & (x23x) & (n_n65) & (!n_n5304)) + ((n_n482) & (x23x) & (n_n65) & (n_n5304)));
	assign n_n2670 = (((!i_9_) & (!n_n528) & (!n_n130) & (!n_n464) & (n_n5200)) + ((!i_9_) & (!n_n528) & (!n_n130) & (n_n464) & (n_n5200)) + ((!i_9_) & (!n_n528) & (n_n130) & (!n_n464) & (n_n5200)) + ((!i_9_) & (!n_n528) & (n_n130) & (n_n464) & (n_n5200)) + ((!i_9_) & (n_n528) & (!n_n130) & (!n_n464) & (n_n5200)) + ((!i_9_) & (n_n528) & (!n_n130) & (n_n464) & (n_n5200)) + ((!i_9_) & (n_n528) & (n_n130) & (!n_n464) & (n_n5200)) + ((!i_9_) & (n_n528) & (n_n130) & (n_n464) & (!n_n5200)) + ((!i_9_) & (n_n528) & (n_n130) & (n_n464) & (n_n5200)) + ((i_9_) & (!n_n528) & (!n_n130) & (!n_n464) & (n_n5200)) + ((i_9_) & (!n_n528) & (!n_n130) & (n_n464) & (n_n5200)) + ((i_9_) & (!n_n528) & (n_n130) & (!n_n464) & (n_n5200)) + ((i_9_) & (!n_n528) & (n_n130) & (n_n464) & (n_n5200)) + ((i_9_) & (n_n528) & (!n_n130) & (!n_n464) & (n_n5200)) + ((i_9_) & (n_n528) & (!n_n130) & (n_n464) & (n_n5200)) + ((i_9_) & (n_n528) & (n_n130) & (!n_n464) & (n_n5200)) + ((i_9_) & (n_n528) & (n_n130) & (n_n464) & (!n_n5200)) + ((i_9_) & (n_n528) & (n_n130) & (n_n464) & (n_n5200)));
	assign x15269x = (((!n_n5181) & (!n_n5185) & (!n_n5191) & (n_n5192)) + ((!n_n5181) & (!n_n5185) & (n_n5191) & (!n_n5192)) + ((!n_n5181) & (!n_n5185) & (n_n5191) & (n_n5192)) + ((!n_n5181) & (n_n5185) & (!n_n5191) & (!n_n5192)) + ((!n_n5181) & (n_n5185) & (!n_n5191) & (n_n5192)) + ((!n_n5181) & (n_n5185) & (n_n5191) & (!n_n5192)) + ((!n_n5181) & (n_n5185) & (n_n5191) & (n_n5192)) + ((n_n5181) & (!n_n5185) & (!n_n5191) & (!n_n5192)) + ((n_n5181) & (!n_n5185) & (!n_n5191) & (n_n5192)) + ((n_n5181) & (!n_n5185) & (n_n5191) & (!n_n5192)) + ((n_n5181) & (!n_n5185) & (n_n5191) & (n_n5192)) + ((n_n5181) & (n_n5185) & (!n_n5191) & (!n_n5192)) + ((n_n5181) & (n_n5185) & (!n_n5191) & (n_n5192)) + ((n_n5181) & (n_n5185) & (n_n5191) & (!n_n5192)) + ((n_n5181) & (n_n5185) & (n_n5191) & (n_n5192)));
	assign x15268x = (((!n_n524) & (!n_n473) & (!n_n520) & (!x12x) & (n_n5187)) + ((!n_n524) & (!n_n473) & (!n_n520) & (x12x) & (n_n5187)) + ((!n_n524) & (!n_n473) & (n_n520) & (!x12x) & (n_n5187)) + ((!n_n524) & (!n_n473) & (n_n520) & (x12x) & (n_n5187)) + ((!n_n524) & (n_n473) & (!n_n520) & (!x12x) & (n_n5187)) + ((!n_n524) & (n_n473) & (!n_n520) & (x12x) & (n_n5187)) + ((!n_n524) & (n_n473) & (n_n520) & (!x12x) & (n_n5187)) + ((!n_n524) & (n_n473) & (n_n520) & (x12x) & (!n_n5187)) + ((!n_n524) & (n_n473) & (n_n520) & (x12x) & (n_n5187)) + ((n_n524) & (!n_n473) & (!n_n520) & (!x12x) & (n_n5187)) + ((n_n524) & (!n_n473) & (!n_n520) & (x12x) & (n_n5187)) + ((n_n524) & (!n_n473) & (n_n520) & (!x12x) & (n_n5187)) + ((n_n524) & (!n_n473) & (n_n520) & (x12x) & (n_n5187)) + ((n_n524) & (n_n473) & (!n_n520) & (!x12x) & (n_n5187)) + ((n_n524) & (n_n473) & (!n_n520) & (x12x) & (!n_n5187)) + ((n_n524) & (n_n473) & (!n_n520) & (x12x) & (n_n5187)) + ((n_n524) & (n_n473) & (n_n520) & (!x12x) & (n_n5187)) + ((n_n524) & (n_n473) & (n_n520) & (x12x) & (!n_n5187)) + ((n_n524) & (n_n473) & (n_n520) & (x12x) & (n_n5187)));
	assign x15270x = (((!x25x) & (!n_n130) & (!n_n464) & (!n_n5182) & (x15268x)) + ((!x25x) & (!n_n130) & (!n_n464) & (n_n5182) & (!x15268x)) + ((!x25x) & (!n_n130) & (!n_n464) & (n_n5182) & (x15268x)) + ((!x25x) & (!n_n130) & (n_n464) & (!n_n5182) & (x15268x)) + ((!x25x) & (!n_n130) & (n_n464) & (n_n5182) & (!x15268x)) + ((!x25x) & (!n_n130) & (n_n464) & (n_n5182) & (x15268x)) + ((!x25x) & (n_n130) & (!n_n464) & (!n_n5182) & (x15268x)) + ((!x25x) & (n_n130) & (!n_n464) & (n_n5182) & (!x15268x)) + ((!x25x) & (n_n130) & (!n_n464) & (n_n5182) & (x15268x)) + ((!x25x) & (n_n130) & (n_n464) & (!n_n5182) & (x15268x)) + ((!x25x) & (n_n130) & (n_n464) & (n_n5182) & (!x15268x)) + ((!x25x) & (n_n130) & (n_n464) & (n_n5182) & (x15268x)) + ((x25x) & (!n_n130) & (!n_n464) & (!n_n5182) & (x15268x)) + ((x25x) & (!n_n130) & (!n_n464) & (n_n5182) & (!x15268x)) + ((x25x) & (!n_n130) & (!n_n464) & (n_n5182) & (x15268x)) + ((x25x) & (!n_n130) & (n_n464) & (!n_n5182) & (x15268x)) + ((x25x) & (!n_n130) & (n_n464) & (n_n5182) & (!x15268x)) + ((x25x) & (!n_n130) & (n_n464) & (n_n5182) & (x15268x)) + ((x25x) & (n_n130) & (!n_n464) & (!n_n5182) & (x15268x)) + ((x25x) & (n_n130) & (!n_n464) & (n_n5182) & (!x15268x)) + ((x25x) & (n_n130) & (!n_n464) & (n_n5182) & (x15268x)) + ((x25x) & (n_n130) & (n_n464) & (!n_n5182) & (!x15268x)) + ((x25x) & (n_n130) & (n_n464) & (!n_n5182) & (x15268x)) + ((x25x) & (n_n130) & (n_n464) & (n_n5182) & (!x15268x)) + ((x25x) & (n_n130) & (n_n464) & (n_n5182) & (x15268x)));
	assign x152x = (((!x25x) & (n_n482) & (!n_n473) & (n_n130) & (x23x)) + ((!x25x) & (n_n482) & (n_n473) & (n_n130) & (x23x)) + ((x25x) & (!n_n482) & (n_n473) & (n_n130) & (!x23x)) + ((x25x) & (!n_n482) & (n_n473) & (n_n130) & (x23x)) + ((x25x) & (n_n482) & (!n_n473) & (n_n130) & (x23x)) + ((x25x) & (n_n482) & (n_n473) & (n_n130) & (!x23x)) + ((x25x) & (n_n482) & (n_n473) & (n_n130) & (x23x)));
	assign x15271x = (((!x21x) & (n_n482) & (n_n130) & (x20x) & (!n_n464)) + ((!x21x) & (n_n482) & (n_n130) & (x20x) & (n_n464)) + ((x21x) & (!n_n482) & (n_n130) & (!x20x) & (n_n464)) + ((x21x) & (!n_n482) & (n_n130) & (x20x) & (n_n464)) + ((x21x) & (n_n482) & (n_n130) & (!x20x) & (n_n464)) + ((x21x) & (n_n482) & (n_n130) & (x20x) & (!n_n464)) + ((x21x) & (n_n482) & (n_n130) & (x20x) & (n_n464)));
	assign x15278x = (((!n_n3399) & (!n_n5176) & (!n_n5197) & (!n_n2670) & (x15271x)) + ((!n_n3399) & (!n_n5176) & (!n_n5197) & (n_n2670) & (!x15271x)) + ((!n_n3399) & (!n_n5176) & (!n_n5197) & (n_n2670) & (x15271x)) + ((!n_n3399) & (!n_n5176) & (n_n5197) & (!n_n2670) & (!x15271x)) + ((!n_n3399) & (!n_n5176) & (n_n5197) & (!n_n2670) & (x15271x)) + ((!n_n3399) & (!n_n5176) & (n_n5197) & (n_n2670) & (!x15271x)) + ((!n_n3399) & (!n_n5176) & (n_n5197) & (n_n2670) & (x15271x)) + ((!n_n3399) & (n_n5176) & (!n_n5197) & (!n_n2670) & (!x15271x)) + ((!n_n3399) & (n_n5176) & (!n_n5197) & (!n_n2670) & (x15271x)) + ((!n_n3399) & (n_n5176) & (!n_n5197) & (n_n2670) & (!x15271x)) + ((!n_n3399) & (n_n5176) & (!n_n5197) & (n_n2670) & (x15271x)) + ((!n_n3399) & (n_n5176) & (n_n5197) & (!n_n2670) & (!x15271x)) + ((!n_n3399) & (n_n5176) & (n_n5197) & (!n_n2670) & (x15271x)) + ((!n_n3399) & (n_n5176) & (n_n5197) & (n_n2670) & (!x15271x)) + ((!n_n3399) & (n_n5176) & (n_n5197) & (n_n2670) & (x15271x)) + ((n_n3399) & (!n_n5176) & (!n_n5197) & (!n_n2670) & (!x15271x)) + ((n_n3399) & (!n_n5176) & (!n_n5197) & (!n_n2670) & (x15271x)) + ((n_n3399) & (!n_n5176) & (!n_n5197) & (n_n2670) & (!x15271x)) + ((n_n3399) & (!n_n5176) & (!n_n5197) & (n_n2670) & (x15271x)) + ((n_n3399) & (!n_n5176) & (n_n5197) & (!n_n2670) & (!x15271x)) + ((n_n3399) & (!n_n5176) & (n_n5197) & (!n_n2670) & (x15271x)) + ((n_n3399) & (!n_n5176) & (n_n5197) & (n_n2670) & (!x15271x)) + ((n_n3399) & (!n_n5176) & (n_n5197) & (n_n2670) & (x15271x)) + ((n_n3399) & (n_n5176) & (!n_n5197) & (!n_n2670) & (!x15271x)) + ((n_n3399) & (n_n5176) & (!n_n5197) & (!n_n2670) & (x15271x)) + ((n_n3399) & (n_n5176) & (!n_n5197) & (n_n2670) & (!x15271x)) + ((n_n3399) & (n_n5176) & (!n_n5197) & (n_n2670) & (x15271x)) + ((n_n3399) & (n_n5176) & (n_n5197) & (!n_n2670) & (!x15271x)) + ((n_n3399) & (n_n5176) & (n_n5197) & (!n_n2670) & (x15271x)) + ((n_n3399) & (n_n5176) & (n_n5197) & (n_n2670) & (!x15271x)) + ((n_n3399) & (n_n5176) & (n_n5197) & (n_n2670) & (x15271x)));
	assign x15277x = (((!n_n5168) & (!n_n5169) & (!x36x) & (!x451x) & (x152x)) + ((!n_n5168) & (!n_n5169) & (!x36x) & (x451x) & (!x152x)) + ((!n_n5168) & (!n_n5169) & (!x36x) & (x451x) & (x152x)) + ((!n_n5168) & (!n_n5169) & (x36x) & (!x451x) & (!x152x)) + ((!n_n5168) & (!n_n5169) & (x36x) & (!x451x) & (x152x)) + ((!n_n5168) & (!n_n5169) & (x36x) & (x451x) & (!x152x)) + ((!n_n5168) & (!n_n5169) & (x36x) & (x451x) & (x152x)) + ((!n_n5168) & (n_n5169) & (!x36x) & (!x451x) & (!x152x)) + ((!n_n5168) & (n_n5169) & (!x36x) & (!x451x) & (x152x)) + ((!n_n5168) & (n_n5169) & (!x36x) & (x451x) & (!x152x)) + ((!n_n5168) & (n_n5169) & (!x36x) & (x451x) & (x152x)) + ((!n_n5168) & (n_n5169) & (x36x) & (!x451x) & (!x152x)) + ((!n_n5168) & (n_n5169) & (x36x) & (!x451x) & (x152x)) + ((!n_n5168) & (n_n5169) & (x36x) & (x451x) & (!x152x)) + ((!n_n5168) & (n_n5169) & (x36x) & (x451x) & (x152x)) + ((n_n5168) & (!n_n5169) & (!x36x) & (!x451x) & (!x152x)) + ((n_n5168) & (!n_n5169) & (!x36x) & (!x451x) & (x152x)) + ((n_n5168) & (!n_n5169) & (!x36x) & (x451x) & (!x152x)) + ((n_n5168) & (!n_n5169) & (!x36x) & (x451x) & (x152x)) + ((n_n5168) & (!n_n5169) & (x36x) & (!x451x) & (!x152x)) + ((n_n5168) & (!n_n5169) & (x36x) & (!x451x) & (x152x)) + ((n_n5168) & (!n_n5169) & (x36x) & (x451x) & (!x152x)) + ((n_n5168) & (!n_n5169) & (x36x) & (x451x) & (x152x)) + ((n_n5168) & (n_n5169) & (!x36x) & (!x451x) & (!x152x)) + ((n_n5168) & (n_n5169) & (!x36x) & (!x451x) & (x152x)) + ((n_n5168) & (n_n5169) & (!x36x) & (x451x) & (!x152x)) + ((n_n5168) & (n_n5169) & (!x36x) & (x451x) & (x152x)) + ((n_n5168) & (n_n5169) & (x36x) & (!x451x) & (!x152x)) + ((n_n5168) & (n_n5169) & (x36x) & (!x451x) & (x152x)) + ((n_n5168) & (n_n5169) & (x36x) & (x451x) & (!x152x)) + ((n_n5168) & (n_n5169) & (x36x) & (x451x) & (x152x)));
	assign x276x = (((!i_9_) & (n_n524) & (n_n390) & (n_n535)) + ((i_9_) & (n_n524) & (n_n390) & (n_n535)));
	assign n_n1446 = (((!n_n5115) & (!n_n4144) & (!n_n5117) & (!x127x) & (x414x)) + ((!n_n5115) & (!n_n4144) & (!n_n5117) & (x127x) & (!x414x)) + ((!n_n5115) & (!n_n4144) & (!n_n5117) & (x127x) & (x414x)) + ((!n_n5115) & (!n_n4144) & (n_n5117) & (!x127x) & (!x414x)) + ((!n_n5115) & (!n_n4144) & (n_n5117) & (!x127x) & (x414x)) + ((!n_n5115) & (!n_n4144) & (n_n5117) & (x127x) & (!x414x)) + ((!n_n5115) & (!n_n4144) & (n_n5117) & (x127x) & (x414x)) + ((!n_n5115) & (n_n4144) & (!n_n5117) & (!x127x) & (!x414x)) + ((!n_n5115) & (n_n4144) & (!n_n5117) & (!x127x) & (x414x)) + ((!n_n5115) & (n_n4144) & (!n_n5117) & (x127x) & (!x414x)) + ((!n_n5115) & (n_n4144) & (!n_n5117) & (x127x) & (x414x)) + ((!n_n5115) & (n_n4144) & (n_n5117) & (!x127x) & (!x414x)) + ((!n_n5115) & (n_n4144) & (n_n5117) & (!x127x) & (x414x)) + ((!n_n5115) & (n_n4144) & (n_n5117) & (x127x) & (!x414x)) + ((!n_n5115) & (n_n4144) & (n_n5117) & (x127x) & (x414x)) + ((n_n5115) & (!n_n4144) & (!n_n5117) & (!x127x) & (!x414x)) + ((n_n5115) & (!n_n4144) & (!n_n5117) & (!x127x) & (x414x)) + ((n_n5115) & (!n_n4144) & (!n_n5117) & (x127x) & (!x414x)) + ((n_n5115) & (!n_n4144) & (!n_n5117) & (x127x) & (x414x)) + ((n_n5115) & (!n_n4144) & (n_n5117) & (!x127x) & (!x414x)) + ((n_n5115) & (!n_n4144) & (n_n5117) & (!x127x) & (x414x)) + ((n_n5115) & (!n_n4144) & (n_n5117) & (x127x) & (!x414x)) + ((n_n5115) & (!n_n4144) & (n_n5117) & (x127x) & (x414x)) + ((n_n5115) & (n_n4144) & (!n_n5117) & (!x127x) & (!x414x)) + ((n_n5115) & (n_n4144) & (!n_n5117) & (!x127x) & (x414x)) + ((n_n5115) & (n_n4144) & (!n_n5117) & (x127x) & (!x414x)) + ((n_n5115) & (n_n4144) & (!n_n5117) & (x127x) & (x414x)) + ((n_n5115) & (n_n4144) & (n_n5117) & (!x127x) & (!x414x)) + ((n_n5115) & (n_n4144) & (n_n5117) & (!x127x) & (x414x)) + ((n_n5115) & (n_n4144) & (n_n5117) & (x127x) & (!x414x)) + ((n_n5115) & (n_n4144) & (n_n5117) & (x127x) & (x414x)));
	assign x364x = (((!i_9_) & (n_n536) & (n_n535) & (n_n530)) + ((i_9_) & (n_n536) & (n_n535) & (n_n530)));
	assign x139x = (((!i_9_) & (n_n390) & (n_n491) & (!n_n520) & (x23x)) + ((!i_9_) & (n_n390) & (n_n491) & (n_n520) & (x23x)) + ((i_9_) & (n_n390) & (n_n491) & (!n_n520) & (x23x)) + ((i_9_) & (n_n390) & (n_n491) & (n_n520) & (!x23x)) + ((i_9_) & (n_n390) & (n_n491) & (n_n520) & (x23x)));
	assign x22149x = (((!x492x) & (!x10x) & (!n_n4607) & (!n_n4641) & (!n_n4638)) + ((!x492x) & (x10x) & (!n_n4607) & (!n_n4641) & (!n_n4638)) + ((x492x) & (!x10x) & (!n_n4607) & (!n_n4641) & (!n_n4638)));
	assign n_n954 = (((!n_n4605) & (!n_n4632) & (!n_n4633) & (!x139x) & (!x22149x)) + ((!n_n4605) & (!n_n4632) & (!n_n4633) & (x139x) & (!x22149x)) + ((!n_n4605) & (!n_n4632) & (!n_n4633) & (x139x) & (x22149x)) + ((!n_n4605) & (!n_n4632) & (n_n4633) & (!x139x) & (!x22149x)) + ((!n_n4605) & (!n_n4632) & (n_n4633) & (!x139x) & (x22149x)) + ((!n_n4605) & (!n_n4632) & (n_n4633) & (x139x) & (!x22149x)) + ((!n_n4605) & (!n_n4632) & (n_n4633) & (x139x) & (x22149x)) + ((!n_n4605) & (n_n4632) & (!n_n4633) & (!x139x) & (!x22149x)) + ((!n_n4605) & (n_n4632) & (!n_n4633) & (!x139x) & (x22149x)) + ((!n_n4605) & (n_n4632) & (!n_n4633) & (x139x) & (!x22149x)) + ((!n_n4605) & (n_n4632) & (!n_n4633) & (x139x) & (x22149x)) + ((!n_n4605) & (n_n4632) & (n_n4633) & (!x139x) & (!x22149x)) + ((!n_n4605) & (n_n4632) & (n_n4633) & (!x139x) & (x22149x)) + ((!n_n4605) & (n_n4632) & (n_n4633) & (x139x) & (!x22149x)) + ((!n_n4605) & (n_n4632) & (n_n4633) & (x139x) & (x22149x)) + ((n_n4605) & (!n_n4632) & (!n_n4633) & (!x139x) & (!x22149x)) + ((n_n4605) & (!n_n4632) & (!n_n4633) & (!x139x) & (x22149x)) + ((n_n4605) & (!n_n4632) & (!n_n4633) & (x139x) & (!x22149x)) + ((n_n4605) & (!n_n4632) & (!n_n4633) & (x139x) & (x22149x)) + ((n_n4605) & (!n_n4632) & (n_n4633) & (!x139x) & (!x22149x)) + ((n_n4605) & (!n_n4632) & (n_n4633) & (!x139x) & (x22149x)) + ((n_n4605) & (!n_n4632) & (n_n4633) & (x139x) & (!x22149x)) + ((n_n4605) & (!n_n4632) & (n_n4633) & (x139x) & (x22149x)) + ((n_n4605) & (n_n4632) & (!n_n4633) & (!x139x) & (!x22149x)) + ((n_n4605) & (n_n4632) & (!n_n4633) & (!x139x) & (x22149x)) + ((n_n4605) & (n_n4632) & (!n_n4633) & (x139x) & (!x22149x)) + ((n_n4605) & (n_n4632) & (!n_n4633) & (x139x) & (x22149x)) + ((n_n4605) & (n_n4632) & (n_n4633) & (!x139x) & (!x22149x)) + ((n_n4605) & (n_n4632) & (n_n4633) & (!x139x) & (x22149x)) + ((n_n4605) & (n_n4632) & (n_n4633) & (x139x) & (!x22149x)) + ((n_n4605) & (n_n4632) & (n_n4633) & (x139x) & (x22149x)));
	assign x11647x = (((!n_n390) & (!n_n473) & (!x24x) & (!n_n4703) & (x312x)) + ((!n_n390) & (!n_n473) & (!x24x) & (n_n4703) & (!x312x)) + ((!n_n390) & (!n_n473) & (!x24x) & (n_n4703) & (x312x)) + ((!n_n390) & (!n_n473) & (x24x) & (!n_n4703) & (x312x)) + ((!n_n390) & (!n_n473) & (x24x) & (n_n4703) & (!x312x)) + ((!n_n390) & (!n_n473) & (x24x) & (n_n4703) & (x312x)) + ((!n_n390) & (n_n473) & (!x24x) & (!n_n4703) & (x312x)) + ((!n_n390) & (n_n473) & (!x24x) & (n_n4703) & (!x312x)) + ((!n_n390) & (n_n473) & (!x24x) & (n_n4703) & (x312x)) + ((!n_n390) & (n_n473) & (x24x) & (!n_n4703) & (x312x)) + ((!n_n390) & (n_n473) & (x24x) & (n_n4703) & (!x312x)) + ((!n_n390) & (n_n473) & (x24x) & (n_n4703) & (x312x)) + ((n_n390) & (!n_n473) & (!x24x) & (!n_n4703) & (x312x)) + ((n_n390) & (!n_n473) & (!x24x) & (n_n4703) & (!x312x)) + ((n_n390) & (!n_n473) & (!x24x) & (n_n4703) & (x312x)) + ((n_n390) & (!n_n473) & (x24x) & (!n_n4703) & (x312x)) + ((n_n390) & (!n_n473) & (x24x) & (n_n4703) & (!x312x)) + ((n_n390) & (!n_n473) & (x24x) & (n_n4703) & (x312x)) + ((n_n390) & (n_n473) & (!x24x) & (!n_n4703) & (x312x)) + ((n_n390) & (n_n473) & (!x24x) & (n_n4703) & (!x312x)) + ((n_n390) & (n_n473) & (!x24x) & (n_n4703) & (x312x)) + ((n_n390) & (n_n473) & (x24x) & (!n_n4703) & (!x312x)) + ((n_n390) & (n_n473) & (x24x) & (!n_n4703) & (x312x)) + ((n_n390) & (n_n473) & (x24x) & (n_n4703) & (!x312x)) + ((n_n390) & (n_n473) & (x24x) & (n_n4703) & (x312x)));
	assign x11648x = (((!n_n4671) & (!n_n4684) & (!n_n4672) & (!n_n4708) & (n_n4723)) + ((!n_n4671) & (!n_n4684) & (!n_n4672) & (n_n4708) & (!n_n4723)) + ((!n_n4671) & (!n_n4684) & (!n_n4672) & (n_n4708) & (n_n4723)) + ((!n_n4671) & (!n_n4684) & (n_n4672) & (!n_n4708) & (!n_n4723)) + ((!n_n4671) & (!n_n4684) & (n_n4672) & (!n_n4708) & (n_n4723)) + ((!n_n4671) & (!n_n4684) & (n_n4672) & (n_n4708) & (!n_n4723)) + ((!n_n4671) & (!n_n4684) & (n_n4672) & (n_n4708) & (n_n4723)) + ((!n_n4671) & (n_n4684) & (!n_n4672) & (!n_n4708) & (!n_n4723)) + ((!n_n4671) & (n_n4684) & (!n_n4672) & (!n_n4708) & (n_n4723)) + ((!n_n4671) & (n_n4684) & (!n_n4672) & (n_n4708) & (!n_n4723)) + ((!n_n4671) & (n_n4684) & (!n_n4672) & (n_n4708) & (n_n4723)) + ((!n_n4671) & (n_n4684) & (n_n4672) & (!n_n4708) & (!n_n4723)) + ((!n_n4671) & (n_n4684) & (n_n4672) & (!n_n4708) & (n_n4723)) + ((!n_n4671) & (n_n4684) & (n_n4672) & (n_n4708) & (!n_n4723)) + ((!n_n4671) & (n_n4684) & (n_n4672) & (n_n4708) & (n_n4723)) + ((n_n4671) & (!n_n4684) & (!n_n4672) & (!n_n4708) & (!n_n4723)) + ((n_n4671) & (!n_n4684) & (!n_n4672) & (!n_n4708) & (n_n4723)) + ((n_n4671) & (!n_n4684) & (!n_n4672) & (n_n4708) & (!n_n4723)) + ((n_n4671) & (!n_n4684) & (!n_n4672) & (n_n4708) & (n_n4723)) + ((n_n4671) & (!n_n4684) & (n_n4672) & (!n_n4708) & (!n_n4723)) + ((n_n4671) & (!n_n4684) & (n_n4672) & (!n_n4708) & (n_n4723)) + ((n_n4671) & (!n_n4684) & (n_n4672) & (n_n4708) & (!n_n4723)) + ((n_n4671) & (!n_n4684) & (n_n4672) & (n_n4708) & (n_n4723)) + ((n_n4671) & (n_n4684) & (!n_n4672) & (!n_n4708) & (!n_n4723)) + ((n_n4671) & (n_n4684) & (!n_n4672) & (!n_n4708) & (n_n4723)) + ((n_n4671) & (n_n4684) & (!n_n4672) & (n_n4708) & (!n_n4723)) + ((n_n4671) & (n_n4684) & (!n_n4672) & (n_n4708) & (n_n4723)) + ((n_n4671) & (n_n4684) & (n_n4672) & (!n_n4708) & (!n_n4723)) + ((n_n4671) & (n_n4684) & (n_n4672) & (!n_n4708) & (n_n4723)) + ((n_n4671) & (n_n4684) & (n_n4672) & (n_n4708) & (!n_n4723)) + ((n_n4671) & (n_n4684) & (n_n4672) & (n_n4708) & (n_n4723)));
	assign x11653x = (((!n_n4601) & (!n_n4571) & (!n_n4587) & (n_n4584)) + ((!n_n4601) & (!n_n4571) & (n_n4587) & (!n_n4584)) + ((!n_n4601) & (!n_n4571) & (n_n4587) & (n_n4584)) + ((!n_n4601) & (n_n4571) & (!n_n4587) & (!n_n4584)) + ((!n_n4601) & (n_n4571) & (!n_n4587) & (n_n4584)) + ((!n_n4601) & (n_n4571) & (n_n4587) & (!n_n4584)) + ((!n_n4601) & (n_n4571) & (n_n4587) & (n_n4584)) + ((n_n4601) & (!n_n4571) & (!n_n4587) & (!n_n4584)) + ((n_n4601) & (!n_n4571) & (!n_n4587) & (n_n4584)) + ((n_n4601) & (!n_n4571) & (n_n4587) & (!n_n4584)) + ((n_n4601) & (!n_n4571) & (n_n4587) & (n_n4584)) + ((n_n4601) & (n_n4571) & (!n_n4587) & (!n_n4584)) + ((n_n4601) & (n_n4571) & (!n_n4587) & (n_n4584)) + ((n_n4601) & (n_n4571) & (n_n4587) & (!n_n4584)) + ((n_n4601) & (n_n4571) & (n_n4587) & (n_n4584)));
	assign x11654x = (((!n_n4577) & (!n_n4576) & (!n_n4574) & (!n_n4550) & (n_n4527)) + ((!n_n4577) & (!n_n4576) & (!n_n4574) & (n_n4550) & (!n_n4527)) + ((!n_n4577) & (!n_n4576) & (!n_n4574) & (n_n4550) & (n_n4527)) + ((!n_n4577) & (!n_n4576) & (n_n4574) & (!n_n4550) & (!n_n4527)) + ((!n_n4577) & (!n_n4576) & (n_n4574) & (!n_n4550) & (n_n4527)) + ((!n_n4577) & (!n_n4576) & (n_n4574) & (n_n4550) & (!n_n4527)) + ((!n_n4577) & (!n_n4576) & (n_n4574) & (n_n4550) & (n_n4527)) + ((!n_n4577) & (n_n4576) & (!n_n4574) & (!n_n4550) & (!n_n4527)) + ((!n_n4577) & (n_n4576) & (!n_n4574) & (!n_n4550) & (n_n4527)) + ((!n_n4577) & (n_n4576) & (!n_n4574) & (n_n4550) & (!n_n4527)) + ((!n_n4577) & (n_n4576) & (!n_n4574) & (n_n4550) & (n_n4527)) + ((!n_n4577) & (n_n4576) & (n_n4574) & (!n_n4550) & (!n_n4527)) + ((!n_n4577) & (n_n4576) & (n_n4574) & (!n_n4550) & (n_n4527)) + ((!n_n4577) & (n_n4576) & (n_n4574) & (n_n4550) & (!n_n4527)) + ((!n_n4577) & (n_n4576) & (n_n4574) & (n_n4550) & (n_n4527)) + ((n_n4577) & (!n_n4576) & (!n_n4574) & (!n_n4550) & (!n_n4527)) + ((n_n4577) & (!n_n4576) & (!n_n4574) & (!n_n4550) & (n_n4527)) + ((n_n4577) & (!n_n4576) & (!n_n4574) & (n_n4550) & (!n_n4527)) + ((n_n4577) & (!n_n4576) & (!n_n4574) & (n_n4550) & (n_n4527)) + ((n_n4577) & (!n_n4576) & (n_n4574) & (!n_n4550) & (!n_n4527)) + ((n_n4577) & (!n_n4576) & (n_n4574) & (!n_n4550) & (n_n4527)) + ((n_n4577) & (!n_n4576) & (n_n4574) & (n_n4550) & (!n_n4527)) + ((n_n4577) & (!n_n4576) & (n_n4574) & (n_n4550) & (n_n4527)) + ((n_n4577) & (n_n4576) & (!n_n4574) & (!n_n4550) & (!n_n4527)) + ((n_n4577) & (n_n4576) & (!n_n4574) & (!n_n4550) & (n_n4527)) + ((n_n4577) & (n_n4576) & (!n_n4574) & (n_n4550) & (!n_n4527)) + ((n_n4577) & (n_n4576) & (!n_n4574) & (n_n4550) & (n_n4527)) + ((n_n4577) & (n_n4576) & (n_n4574) & (!n_n4550) & (!n_n4527)) + ((n_n4577) & (n_n4576) & (n_n4574) & (!n_n4550) & (n_n4527)) + ((n_n4577) & (n_n4576) & (n_n4574) & (n_n4550) & (!n_n4527)) + ((n_n4577) & (n_n4576) & (n_n4574) & (n_n4550) & (n_n4527)));
	assign n_n942 = (((!n_n954) & (!x11647x) & (!x11648x) & (!x11653x) & (x11654x)) + ((!n_n954) & (!x11647x) & (!x11648x) & (x11653x) & (!x11654x)) + ((!n_n954) & (!x11647x) & (!x11648x) & (x11653x) & (x11654x)) + ((!n_n954) & (!x11647x) & (x11648x) & (!x11653x) & (!x11654x)) + ((!n_n954) & (!x11647x) & (x11648x) & (!x11653x) & (x11654x)) + ((!n_n954) & (!x11647x) & (x11648x) & (x11653x) & (!x11654x)) + ((!n_n954) & (!x11647x) & (x11648x) & (x11653x) & (x11654x)) + ((!n_n954) & (x11647x) & (!x11648x) & (!x11653x) & (!x11654x)) + ((!n_n954) & (x11647x) & (!x11648x) & (!x11653x) & (x11654x)) + ((!n_n954) & (x11647x) & (!x11648x) & (x11653x) & (!x11654x)) + ((!n_n954) & (x11647x) & (!x11648x) & (x11653x) & (x11654x)) + ((!n_n954) & (x11647x) & (x11648x) & (!x11653x) & (!x11654x)) + ((!n_n954) & (x11647x) & (x11648x) & (!x11653x) & (x11654x)) + ((!n_n954) & (x11647x) & (x11648x) & (x11653x) & (!x11654x)) + ((!n_n954) & (x11647x) & (x11648x) & (x11653x) & (x11654x)) + ((n_n954) & (!x11647x) & (!x11648x) & (!x11653x) & (!x11654x)) + ((n_n954) & (!x11647x) & (!x11648x) & (!x11653x) & (x11654x)) + ((n_n954) & (!x11647x) & (!x11648x) & (x11653x) & (!x11654x)) + ((n_n954) & (!x11647x) & (!x11648x) & (x11653x) & (x11654x)) + ((n_n954) & (!x11647x) & (x11648x) & (!x11653x) & (!x11654x)) + ((n_n954) & (!x11647x) & (x11648x) & (!x11653x) & (x11654x)) + ((n_n954) & (!x11647x) & (x11648x) & (x11653x) & (!x11654x)) + ((n_n954) & (!x11647x) & (x11648x) & (x11653x) & (x11654x)) + ((n_n954) & (x11647x) & (!x11648x) & (!x11653x) & (!x11654x)) + ((n_n954) & (x11647x) & (!x11648x) & (!x11653x) & (x11654x)) + ((n_n954) & (x11647x) & (!x11648x) & (x11653x) & (!x11654x)) + ((n_n954) & (x11647x) & (!x11648x) & (x11653x) & (x11654x)) + ((n_n954) & (x11647x) & (x11648x) & (!x11653x) & (!x11654x)) + ((n_n954) & (x11647x) & (x11648x) & (!x11653x) & (x11654x)) + ((n_n954) & (x11647x) & (x11648x) & (x11653x) & (!x11654x)) + ((n_n954) & (x11647x) & (x11648x) & (x11653x) & (x11654x)));
	assign n_n725 = (((!n_n4470) & (!n_n4472) & (!n_n3515) & (!n_n901) & (n_n4476)) + ((!n_n4470) & (!n_n4472) & (!n_n3515) & (n_n901) & (!n_n4476)) + ((!n_n4470) & (!n_n4472) & (!n_n3515) & (n_n901) & (n_n4476)) + ((!n_n4470) & (!n_n4472) & (n_n3515) & (!n_n901) & (!n_n4476)) + ((!n_n4470) & (!n_n4472) & (n_n3515) & (!n_n901) & (n_n4476)) + ((!n_n4470) & (!n_n4472) & (n_n3515) & (n_n901) & (!n_n4476)) + ((!n_n4470) & (!n_n4472) & (n_n3515) & (n_n901) & (n_n4476)) + ((!n_n4470) & (n_n4472) & (!n_n3515) & (!n_n901) & (!n_n4476)) + ((!n_n4470) & (n_n4472) & (!n_n3515) & (!n_n901) & (n_n4476)) + ((!n_n4470) & (n_n4472) & (!n_n3515) & (n_n901) & (!n_n4476)) + ((!n_n4470) & (n_n4472) & (!n_n3515) & (n_n901) & (n_n4476)) + ((!n_n4470) & (n_n4472) & (n_n3515) & (!n_n901) & (!n_n4476)) + ((!n_n4470) & (n_n4472) & (n_n3515) & (!n_n901) & (n_n4476)) + ((!n_n4470) & (n_n4472) & (n_n3515) & (n_n901) & (!n_n4476)) + ((!n_n4470) & (n_n4472) & (n_n3515) & (n_n901) & (n_n4476)) + ((n_n4470) & (!n_n4472) & (!n_n3515) & (!n_n901) & (!n_n4476)) + ((n_n4470) & (!n_n4472) & (!n_n3515) & (!n_n901) & (n_n4476)) + ((n_n4470) & (!n_n4472) & (!n_n3515) & (n_n901) & (!n_n4476)) + ((n_n4470) & (!n_n4472) & (!n_n3515) & (n_n901) & (n_n4476)) + ((n_n4470) & (!n_n4472) & (n_n3515) & (!n_n901) & (!n_n4476)) + ((n_n4470) & (!n_n4472) & (n_n3515) & (!n_n901) & (n_n4476)) + ((n_n4470) & (!n_n4472) & (n_n3515) & (n_n901) & (!n_n4476)) + ((n_n4470) & (!n_n4472) & (n_n3515) & (n_n901) & (n_n4476)) + ((n_n4470) & (n_n4472) & (!n_n3515) & (!n_n901) & (!n_n4476)) + ((n_n4470) & (n_n4472) & (!n_n3515) & (!n_n901) & (n_n4476)) + ((n_n4470) & (n_n4472) & (!n_n3515) & (n_n901) & (!n_n4476)) + ((n_n4470) & (n_n4472) & (!n_n3515) & (n_n901) & (n_n4476)) + ((n_n4470) & (n_n4472) & (n_n3515) & (!n_n901) & (!n_n4476)) + ((n_n4470) & (n_n4472) & (n_n3515) & (!n_n901) & (n_n4476)) + ((n_n4470) & (n_n4472) & (n_n3515) & (n_n901) & (!n_n4476)) + ((n_n4470) & (n_n4472) & (n_n3515) & (n_n901) & (n_n4476)));
	assign x13025x = (((!x25x) & (!n_n455) & (!x24x) & (!n_n500) & (x70x)) + ((!x25x) & (!n_n455) & (!x24x) & (n_n500) & (x70x)) + ((!x25x) & (!n_n455) & (x24x) & (!n_n500) & (x70x)) + ((!x25x) & (!n_n455) & (x24x) & (n_n500) & (x70x)) + ((!x25x) & (n_n455) & (!x24x) & (!n_n500) & (x70x)) + ((!x25x) & (n_n455) & (!x24x) & (n_n500) & (x70x)) + ((!x25x) & (n_n455) & (x24x) & (!n_n500) & (x70x)) + ((!x25x) & (n_n455) & (x24x) & (n_n500) & (!x70x)) + ((!x25x) & (n_n455) & (x24x) & (n_n500) & (x70x)) + ((x25x) & (!n_n455) & (!x24x) & (!n_n500) & (x70x)) + ((x25x) & (!n_n455) & (!x24x) & (n_n500) & (x70x)) + ((x25x) & (!n_n455) & (x24x) & (!n_n500) & (x70x)) + ((x25x) & (!n_n455) & (x24x) & (n_n500) & (x70x)) + ((x25x) & (n_n455) & (!x24x) & (!n_n500) & (x70x)) + ((x25x) & (n_n455) & (!x24x) & (n_n500) & (!x70x)) + ((x25x) & (n_n455) & (!x24x) & (n_n500) & (x70x)) + ((x25x) & (n_n455) & (x24x) & (!n_n500) & (x70x)) + ((x25x) & (n_n455) & (x24x) & (n_n500) & (!x70x)) + ((x25x) & (n_n455) & (x24x) & (n_n500) & (x70x)));
	assign x13026x = (((!n_n4494) & (!n_n4495) & (!n_n4487) & (!n_n4492) & (n_n4486)) + ((!n_n4494) & (!n_n4495) & (!n_n4487) & (n_n4492) & (!n_n4486)) + ((!n_n4494) & (!n_n4495) & (!n_n4487) & (n_n4492) & (n_n4486)) + ((!n_n4494) & (!n_n4495) & (n_n4487) & (!n_n4492) & (!n_n4486)) + ((!n_n4494) & (!n_n4495) & (n_n4487) & (!n_n4492) & (n_n4486)) + ((!n_n4494) & (!n_n4495) & (n_n4487) & (n_n4492) & (!n_n4486)) + ((!n_n4494) & (!n_n4495) & (n_n4487) & (n_n4492) & (n_n4486)) + ((!n_n4494) & (n_n4495) & (!n_n4487) & (!n_n4492) & (!n_n4486)) + ((!n_n4494) & (n_n4495) & (!n_n4487) & (!n_n4492) & (n_n4486)) + ((!n_n4494) & (n_n4495) & (!n_n4487) & (n_n4492) & (!n_n4486)) + ((!n_n4494) & (n_n4495) & (!n_n4487) & (n_n4492) & (n_n4486)) + ((!n_n4494) & (n_n4495) & (n_n4487) & (!n_n4492) & (!n_n4486)) + ((!n_n4494) & (n_n4495) & (n_n4487) & (!n_n4492) & (n_n4486)) + ((!n_n4494) & (n_n4495) & (n_n4487) & (n_n4492) & (!n_n4486)) + ((!n_n4494) & (n_n4495) & (n_n4487) & (n_n4492) & (n_n4486)) + ((n_n4494) & (!n_n4495) & (!n_n4487) & (!n_n4492) & (!n_n4486)) + ((n_n4494) & (!n_n4495) & (!n_n4487) & (!n_n4492) & (n_n4486)) + ((n_n4494) & (!n_n4495) & (!n_n4487) & (n_n4492) & (!n_n4486)) + ((n_n4494) & (!n_n4495) & (!n_n4487) & (n_n4492) & (n_n4486)) + ((n_n4494) & (!n_n4495) & (n_n4487) & (!n_n4492) & (!n_n4486)) + ((n_n4494) & (!n_n4495) & (n_n4487) & (!n_n4492) & (n_n4486)) + ((n_n4494) & (!n_n4495) & (n_n4487) & (n_n4492) & (!n_n4486)) + ((n_n4494) & (!n_n4495) & (n_n4487) & (n_n4492) & (n_n4486)) + ((n_n4494) & (n_n4495) & (!n_n4487) & (!n_n4492) & (!n_n4486)) + ((n_n4494) & (n_n4495) & (!n_n4487) & (!n_n4492) & (n_n4486)) + ((n_n4494) & (n_n4495) & (!n_n4487) & (n_n4492) & (!n_n4486)) + ((n_n4494) & (n_n4495) & (!n_n4487) & (n_n4492) & (n_n4486)) + ((n_n4494) & (n_n4495) & (n_n4487) & (!n_n4492) & (!n_n4486)) + ((n_n4494) & (n_n4495) & (n_n4487) & (!n_n4492) & (n_n4486)) + ((n_n4494) & (n_n4495) & (n_n4487) & (n_n4492) & (!n_n4486)) + ((n_n4494) & (n_n4495) & (n_n4487) & (n_n4492) & (n_n4486)));
	assign x22171x = (((!x552x) & (!x20x) & (!x23x) & (!n_n4833) & (!x12741x)) + ((!x552x) & (!x20x) & (x23x) & (!n_n4833) & (!x12741x)) + ((!x552x) & (x20x) & (!x23x) & (!n_n4833) & (!x12741x)) + ((!x552x) & (x20x) & (x23x) & (!n_n4833) & (!x12741x)) + ((x552x) & (!x20x) & (!x23x) & (!n_n4833) & (!x12741x)));
	assign n_n698 = (((!x21x) & (!x552x) & (!n_n4832) & (!n_n4828) & (!x22171x)) + ((!x21x) & (!x552x) & (!n_n4832) & (n_n4828) & (!x22171x)) + ((!x21x) & (!x552x) & (!n_n4832) & (n_n4828) & (x22171x)) + ((!x21x) & (!x552x) & (n_n4832) & (!n_n4828) & (!x22171x)) + ((!x21x) & (!x552x) & (n_n4832) & (!n_n4828) & (x22171x)) + ((!x21x) & (!x552x) & (n_n4832) & (n_n4828) & (!x22171x)) + ((!x21x) & (!x552x) & (n_n4832) & (n_n4828) & (x22171x)) + ((!x21x) & (x552x) & (!n_n4832) & (!n_n4828) & (!x22171x)) + ((!x21x) & (x552x) & (!n_n4832) & (n_n4828) & (!x22171x)) + ((!x21x) & (x552x) & (!n_n4832) & (n_n4828) & (x22171x)) + ((!x21x) & (x552x) & (n_n4832) & (!n_n4828) & (!x22171x)) + ((!x21x) & (x552x) & (n_n4832) & (!n_n4828) & (x22171x)) + ((!x21x) & (x552x) & (n_n4832) & (n_n4828) & (!x22171x)) + ((!x21x) & (x552x) & (n_n4832) & (n_n4828) & (x22171x)) + ((x21x) & (!x552x) & (!n_n4832) & (!n_n4828) & (!x22171x)) + ((x21x) & (!x552x) & (!n_n4832) & (n_n4828) & (!x22171x)) + ((x21x) & (!x552x) & (!n_n4832) & (n_n4828) & (x22171x)) + ((x21x) & (!x552x) & (n_n4832) & (!n_n4828) & (!x22171x)) + ((x21x) & (!x552x) & (n_n4832) & (!n_n4828) & (x22171x)) + ((x21x) & (!x552x) & (n_n4832) & (n_n4828) & (!x22171x)) + ((x21x) & (!x552x) & (n_n4832) & (n_n4828) & (x22171x)) + ((x21x) & (x552x) & (!n_n4832) & (!n_n4828) & (!x22171x)) + ((x21x) & (x552x) & (!n_n4832) & (!n_n4828) & (x22171x)) + ((x21x) & (x552x) & (!n_n4832) & (n_n4828) & (!x22171x)) + ((x21x) & (x552x) & (!n_n4832) & (n_n4828) & (x22171x)) + ((x21x) & (x552x) & (n_n4832) & (!n_n4828) & (!x22171x)) + ((x21x) & (x552x) & (n_n4832) & (!n_n4828) & (x22171x)) + ((x21x) & (x552x) & (n_n4832) & (n_n4828) & (!x22171x)) + ((x21x) & (x552x) & (n_n4832) & (n_n4828) & (x22171x)));
	assign x52x = (((!i_9_) & (n_n518) & (n_n528) & (n_n260)) + ((i_9_) & (n_n518) & (n_n528) & (n_n260)));
	assign x150x = (((!i_9_) & (!i_7_) & (!i_8_) & (!i_6_) & (x530x)) + ((!i_9_) & (i_7_) & (i_8_) & (!i_6_) & (x530x)));
	assign x326x = (((!i_9_) & (n_n532) & (!n_n534) & (n_n260) & (n_n535)) + ((!i_9_) & (n_n532) & (n_n534) & (n_n260) & (n_n535)) + ((i_9_) & (!n_n532) & (n_n534) & (n_n260) & (n_n535)) + ((i_9_) & (n_n532) & (n_n534) & (n_n260) & (n_n535)));
	assign x12745x = (((!i_7_) & (i_8_) & (i_6_) & (n_n518) & (x17x)) + ((i_7_) & (i_8_) & (i_6_) & (n_n518) & (x17x)));
	assign x12752x = (((!n_n4826) & (!n_n4822) & (!n_n834) & (!n_n4196) & (x12745x)) + ((!n_n4826) & (!n_n4822) & (!n_n834) & (n_n4196) & (!x12745x)) + ((!n_n4826) & (!n_n4822) & (!n_n834) & (n_n4196) & (x12745x)) + ((!n_n4826) & (!n_n4822) & (n_n834) & (!n_n4196) & (!x12745x)) + ((!n_n4826) & (!n_n4822) & (n_n834) & (!n_n4196) & (x12745x)) + ((!n_n4826) & (!n_n4822) & (n_n834) & (n_n4196) & (!x12745x)) + ((!n_n4826) & (!n_n4822) & (n_n834) & (n_n4196) & (x12745x)) + ((!n_n4826) & (n_n4822) & (!n_n834) & (!n_n4196) & (!x12745x)) + ((!n_n4826) & (n_n4822) & (!n_n834) & (!n_n4196) & (x12745x)) + ((!n_n4826) & (n_n4822) & (!n_n834) & (n_n4196) & (!x12745x)) + ((!n_n4826) & (n_n4822) & (!n_n834) & (n_n4196) & (x12745x)) + ((!n_n4826) & (n_n4822) & (n_n834) & (!n_n4196) & (!x12745x)) + ((!n_n4826) & (n_n4822) & (n_n834) & (!n_n4196) & (x12745x)) + ((!n_n4826) & (n_n4822) & (n_n834) & (n_n4196) & (!x12745x)) + ((!n_n4826) & (n_n4822) & (n_n834) & (n_n4196) & (x12745x)) + ((n_n4826) & (!n_n4822) & (!n_n834) & (!n_n4196) & (!x12745x)) + ((n_n4826) & (!n_n4822) & (!n_n834) & (!n_n4196) & (x12745x)) + ((n_n4826) & (!n_n4822) & (!n_n834) & (n_n4196) & (!x12745x)) + ((n_n4826) & (!n_n4822) & (!n_n834) & (n_n4196) & (x12745x)) + ((n_n4826) & (!n_n4822) & (n_n834) & (!n_n4196) & (!x12745x)) + ((n_n4826) & (!n_n4822) & (n_n834) & (!n_n4196) & (x12745x)) + ((n_n4826) & (!n_n4822) & (n_n834) & (n_n4196) & (!x12745x)) + ((n_n4826) & (!n_n4822) & (n_n834) & (n_n4196) & (x12745x)) + ((n_n4826) & (n_n4822) & (!n_n834) & (!n_n4196) & (!x12745x)) + ((n_n4826) & (n_n4822) & (!n_n834) & (!n_n4196) & (x12745x)) + ((n_n4826) & (n_n4822) & (!n_n834) & (n_n4196) & (!x12745x)) + ((n_n4826) & (n_n4822) & (!n_n834) & (n_n4196) & (x12745x)) + ((n_n4826) & (n_n4822) & (n_n834) & (!n_n4196) & (!x12745x)) + ((n_n4826) & (n_n4822) & (n_n834) & (!n_n4196) & (x12745x)) + ((n_n4826) & (n_n4822) & (n_n834) & (n_n4196) & (!x12745x)) + ((n_n4826) & (n_n4822) & (n_n834) & (n_n4196) & (x12745x)));
	assign x12656x = (((!n_n5089) & (!n_n5098) & (!n_n5105) & (n_n5103)) + ((!n_n5089) & (!n_n5098) & (n_n5105) & (!n_n5103)) + ((!n_n5089) & (!n_n5098) & (n_n5105) & (n_n5103)) + ((!n_n5089) & (n_n5098) & (!n_n5105) & (!n_n5103)) + ((!n_n5089) & (n_n5098) & (!n_n5105) & (n_n5103)) + ((!n_n5089) & (n_n5098) & (n_n5105) & (!n_n5103)) + ((!n_n5089) & (n_n5098) & (n_n5105) & (n_n5103)) + ((n_n5089) & (!n_n5098) & (!n_n5105) & (!n_n5103)) + ((n_n5089) & (!n_n5098) & (!n_n5105) & (n_n5103)) + ((n_n5089) & (!n_n5098) & (n_n5105) & (!n_n5103)) + ((n_n5089) & (!n_n5098) & (n_n5105) & (n_n5103)) + ((n_n5089) & (n_n5098) & (!n_n5105) & (!n_n5103)) + ((n_n5089) & (n_n5098) & (!n_n5105) & (n_n5103)) + ((n_n5089) & (n_n5098) & (n_n5105) & (!n_n5103)) + ((n_n5089) & (n_n5098) & (n_n5105) & (n_n5103)));
	assign x12657x = (((!n_n5096) & (!n_n5100) & (!n_n5104) & (!n_n5078) & (n_n5090)) + ((!n_n5096) & (!n_n5100) & (!n_n5104) & (n_n5078) & (!n_n5090)) + ((!n_n5096) & (!n_n5100) & (!n_n5104) & (n_n5078) & (n_n5090)) + ((!n_n5096) & (!n_n5100) & (n_n5104) & (!n_n5078) & (!n_n5090)) + ((!n_n5096) & (!n_n5100) & (n_n5104) & (!n_n5078) & (n_n5090)) + ((!n_n5096) & (!n_n5100) & (n_n5104) & (n_n5078) & (!n_n5090)) + ((!n_n5096) & (!n_n5100) & (n_n5104) & (n_n5078) & (n_n5090)) + ((!n_n5096) & (n_n5100) & (!n_n5104) & (!n_n5078) & (!n_n5090)) + ((!n_n5096) & (n_n5100) & (!n_n5104) & (!n_n5078) & (n_n5090)) + ((!n_n5096) & (n_n5100) & (!n_n5104) & (n_n5078) & (!n_n5090)) + ((!n_n5096) & (n_n5100) & (!n_n5104) & (n_n5078) & (n_n5090)) + ((!n_n5096) & (n_n5100) & (n_n5104) & (!n_n5078) & (!n_n5090)) + ((!n_n5096) & (n_n5100) & (n_n5104) & (!n_n5078) & (n_n5090)) + ((!n_n5096) & (n_n5100) & (n_n5104) & (n_n5078) & (!n_n5090)) + ((!n_n5096) & (n_n5100) & (n_n5104) & (n_n5078) & (n_n5090)) + ((n_n5096) & (!n_n5100) & (!n_n5104) & (!n_n5078) & (!n_n5090)) + ((n_n5096) & (!n_n5100) & (!n_n5104) & (!n_n5078) & (n_n5090)) + ((n_n5096) & (!n_n5100) & (!n_n5104) & (n_n5078) & (!n_n5090)) + ((n_n5096) & (!n_n5100) & (!n_n5104) & (n_n5078) & (n_n5090)) + ((n_n5096) & (!n_n5100) & (n_n5104) & (!n_n5078) & (!n_n5090)) + ((n_n5096) & (!n_n5100) & (n_n5104) & (!n_n5078) & (n_n5090)) + ((n_n5096) & (!n_n5100) & (n_n5104) & (n_n5078) & (!n_n5090)) + ((n_n5096) & (!n_n5100) & (n_n5104) & (n_n5078) & (n_n5090)) + ((n_n5096) & (n_n5100) & (!n_n5104) & (!n_n5078) & (!n_n5090)) + ((n_n5096) & (n_n5100) & (!n_n5104) & (!n_n5078) & (n_n5090)) + ((n_n5096) & (n_n5100) & (!n_n5104) & (n_n5078) & (!n_n5090)) + ((n_n5096) & (n_n5100) & (!n_n5104) & (n_n5078) & (n_n5090)) + ((n_n5096) & (n_n5100) & (n_n5104) & (!n_n5078) & (!n_n5090)) + ((n_n5096) & (n_n5100) & (n_n5104) & (!n_n5078) & (n_n5090)) + ((n_n5096) & (n_n5100) & (n_n5104) & (n_n5078) & (!n_n5090)) + ((n_n5096) & (n_n5100) & (n_n5104) & (n_n5078) & (n_n5090)));
	assign x53x = (((!i_9_) & (n_n536) & (n_n524) & (n_n518)) + ((i_9_) & (n_n536) & (n_n524) & (n_n518)));
	assign n_n4103 = (((!n_n4344) & (!n_n4345) & (!x67x) & (!x156x) & (x469x)) + ((!n_n4344) & (!n_n4345) & (!x67x) & (x156x) & (!x469x)) + ((!n_n4344) & (!n_n4345) & (!x67x) & (x156x) & (x469x)) + ((!n_n4344) & (!n_n4345) & (x67x) & (!x156x) & (!x469x)) + ((!n_n4344) & (!n_n4345) & (x67x) & (!x156x) & (x469x)) + ((!n_n4344) & (!n_n4345) & (x67x) & (x156x) & (!x469x)) + ((!n_n4344) & (!n_n4345) & (x67x) & (x156x) & (x469x)) + ((!n_n4344) & (n_n4345) & (!x67x) & (!x156x) & (!x469x)) + ((!n_n4344) & (n_n4345) & (!x67x) & (!x156x) & (x469x)) + ((!n_n4344) & (n_n4345) & (!x67x) & (x156x) & (!x469x)) + ((!n_n4344) & (n_n4345) & (!x67x) & (x156x) & (x469x)) + ((!n_n4344) & (n_n4345) & (x67x) & (!x156x) & (!x469x)) + ((!n_n4344) & (n_n4345) & (x67x) & (!x156x) & (x469x)) + ((!n_n4344) & (n_n4345) & (x67x) & (x156x) & (!x469x)) + ((!n_n4344) & (n_n4345) & (x67x) & (x156x) & (x469x)) + ((n_n4344) & (!n_n4345) & (!x67x) & (!x156x) & (!x469x)) + ((n_n4344) & (!n_n4345) & (!x67x) & (!x156x) & (x469x)) + ((n_n4344) & (!n_n4345) & (!x67x) & (x156x) & (!x469x)) + ((n_n4344) & (!n_n4345) & (!x67x) & (x156x) & (x469x)) + ((n_n4344) & (!n_n4345) & (x67x) & (!x156x) & (!x469x)) + ((n_n4344) & (!n_n4345) & (x67x) & (!x156x) & (x469x)) + ((n_n4344) & (!n_n4345) & (x67x) & (x156x) & (!x469x)) + ((n_n4344) & (!n_n4345) & (x67x) & (x156x) & (x469x)) + ((n_n4344) & (n_n4345) & (!x67x) & (!x156x) & (!x469x)) + ((n_n4344) & (n_n4345) & (!x67x) & (!x156x) & (x469x)) + ((n_n4344) & (n_n4345) & (!x67x) & (x156x) & (!x469x)) + ((n_n4344) & (n_n4345) & (!x67x) & (x156x) & (x469x)) + ((n_n4344) & (n_n4345) & (x67x) & (!x156x) & (!x469x)) + ((n_n4344) & (n_n4345) & (x67x) & (!x156x) & (x469x)) + ((n_n4344) & (n_n4345) & (x67x) & (x156x) & (!x469x)) + ((n_n4344) & (n_n4345) & (x67x) & (x156x) & (x469x)));
	assign x443x = (((!i_9_) & (n_n536) & (n_n518) & (!n_n528) & (n_n530)) + ((!i_9_) & (n_n536) & (n_n518) & (n_n528) & (n_n530)) + ((i_9_) & (n_n536) & (n_n518) & (n_n528) & (!n_n530)) + ((i_9_) & (n_n536) & (n_n518) & (n_n528) & (n_n530)));
	assign x13513x = (((i_9_) & (n_n536) & (!n_n518) & (n_n526) & (n_n535)) + ((i_9_) & (n_n536) & (n_n518) & (n_n526) & (!n_n535)) + ((i_9_) & (n_n536) & (n_n518) & (n_n526) & (n_n535)));
	assign x13519x = (((!n_n2446) & (!n_n4279) & (!n_n4316) & (!n_n4313) & (x13513x)) + ((!n_n2446) & (!n_n4279) & (!n_n4316) & (n_n4313) & (!x13513x)) + ((!n_n2446) & (!n_n4279) & (!n_n4316) & (n_n4313) & (x13513x)) + ((!n_n2446) & (!n_n4279) & (n_n4316) & (!n_n4313) & (!x13513x)) + ((!n_n2446) & (!n_n4279) & (n_n4316) & (!n_n4313) & (x13513x)) + ((!n_n2446) & (!n_n4279) & (n_n4316) & (n_n4313) & (!x13513x)) + ((!n_n2446) & (!n_n4279) & (n_n4316) & (n_n4313) & (x13513x)) + ((!n_n2446) & (n_n4279) & (!n_n4316) & (!n_n4313) & (!x13513x)) + ((!n_n2446) & (n_n4279) & (!n_n4316) & (!n_n4313) & (x13513x)) + ((!n_n2446) & (n_n4279) & (!n_n4316) & (n_n4313) & (!x13513x)) + ((!n_n2446) & (n_n4279) & (!n_n4316) & (n_n4313) & (x13513x)) + ((!n_n2446) & (n_n4279) & (n_n4316) & (!n_n4313) & (!x13513x)) + ((!n_n2446) & (n_n4279) & (n_n4316) & (!n_n4313) & (x13513x)) + ((!n_n2446) & (n_n4279) & (n_n4316) & (n_n4313) & (!x13513x)) + ((!n_n2446) & (n_n4279) & (n_n4316) & (n_n4313) & (x13513x)) + ((n_n2446) & (!n_n4279) & (!n_n4316) & (!n_n4313) & (!x13513x)) + ((n_n2446) & (!n_n4279) & (!n_n4316) & (!n_n4313) & (x13513x)) + ((n_n2446) & (!n_n4279) & (!n_n4316) & (n_n4313) & (!x13513x)) + ((n_n2446) & (!n_n4279) & (!n_n4316) & (n_n4313) & (x13513x)) + ((n_n2446) & (!n_n4279) & (n_n4316) & (!n_n4313) & (!x13513x)) + ((n_n2446) & (!n_n4279) & (n_n4316) & (!n_n4313) & (x13513x)) + ((n_n2446) & (!n_n4279) & (n_n4316) & (n_n4313) & (!x13513x)) + ((n_n2446) & (!n_n4279) & (n_n4316) & (n_n4313) & (x13513x)) + ((n_n2446) & (n_n4279) & (!n_n4316) & (!n_n4313) & (!x13513x)) + ((n_n2446) & (n_n4279) & (!n_n4316) & (!n_n4313) & (x13513x)) + ((n_n2446) & (n_n4279) & (!n_n4316) & (n_n4313) & (!x13513x)) + ((n_n2446) & (n_n4279) & (!n_n4316) & (n_n4313) & (x13513x)) + ((n_n2446) & (n_n4279) & (n_n4316) & (!n_n4313) & (!x13513x)) + ((n_n2446) & (n_n4279) & (n_n4316) & (!n_n4313) & (x13513x)) + ((n_n2446) & (n_n4279) & (n_n4316) & (n_n4313) & (!x13513x)) + ((n_n2446) & (n_n4279) & (n_n4316) & (n_n4313) & (x13513x)));
	assign x407x = (((!i_9_) & (n_n532) & (n_n491) & (!n_n130) & (x12x)) + ((!i_9_) & (n_n532) & (n_n491) & (n_n130) & (!x12x)) + ((!i_9_) & (n_n532) & (n_n491) & (n_n130) & (x12x)) + ((i_9_) & (n_n532) & (n_n491) & (!n_n130) & (x12x)) + ((i_9_) & (n_n532) & (n_n491) & (n_n130) & (x12x)));
	assign n_n814 = (((!i_9_) & (!n_n524) & (n_n526) & (n_n260) & (n_n464)) + ((!i_9_) & (n_n524) & (!n_n526) & (n_n260) & (n_n464)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n260) & (n_n464)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n260) & (n_n464)) + ((i_9_) & (n_n524) & (n_n526) & (n_n260) & (n_n464)));
	assign x137x = (((!n_n4975) & (!n_n4973) & (!n_n4971) & (!x228x) & (n_n4972)) + ((!n_n4975) & (!n_n4973) & (!n_n4971) & (x228x) & (!n_n4972)) + ((!n_n4975) & (!n_n4973) & (!n_n4971) & (x228x) & (n_n4972)) + ((!n_n4975) & (!n_n4973) & (n_n4971) & (!x228x) & (!n_n4972)) + ((!n_n4975) & (!n_n4973) & (n_n4971) & (!x228x) & (n_n4972)) + ((!n_n4975) & (!n_n4973) & (n_n4971) & (x228x) & (!n_n4972)) + ((!n_n4975) & (!n_n4973) & (n_n4971) & (x228x) & (n_n4972)) + ((!n_n4975) & (n_n4973) & (!n_n4971) & (!x228x) & (!n_n4972)) + ((!n_n4975) & (n_n4973) & (!n_n4971) & (!x228x) & (n_n4972)) + ((!n_n4975) & (n_n4973) & (!n_n4971) & (x228x) & (!n_n4972)) + ((!n_n4975) & (n_n4973) & (!n_n4971) & (x228x) & (n_n4972)) + ((!n_n4975) & (n_n4973) & (n_n4971) & (!x228x) & (!n_n4972)) + ((!n_n4975) & (n_n4973) & (n_n4971) & (!x228x) & (n_n4972)) + ((!n_n4975) & (n_n4973) & (n_n4971) & (x228x) & (!n_n4972)) + ((!n_n4975) & (n_n4973) & (n_n4971) & (x228x) & (n_n4972)) + ((n_n4975) & (!n_n4973) & (!n_n4971) & (!x228x) & (!n_n4972)) + ((n_n4975) & (!n_n4973) & (!n_n4971) & (!x228x) & (n_n4972)) + ((n_n4975) & (!n_n4973) & (!n_n4971) & (x228x) & (!n_n4972)) + ((n_n4975) & (!n_n4973) & (!n_n4971) & (x228x) & (n_n4972)) + ((n_n4975) & (!n_n4973) & (n_n4971) & (!x228x) & (!n_n4972)) + ((n_n4975) & (!n_n4973) & (n_n4971) & (!x228x) & (n_n4972)) + ((n_n4975) & (!n_n4973) & (n_n4971) & (x228x) & (!n_n4972)) + ((n_n4975) & (!n_n4973) & (n_n4971) & (x228x) & (n_n4972)) + ((n_n4975) & (n_n4973) & (!n_n4971) & (!x228x) & (!n_n4972)) + ((n_n4975) & (n_n4973) & (!n_n4971) & (!x228x) & (n_n4972)) + ((n_n4975) & (n_n4973) & (!n_n4971) & (x228x) & (!n_n4972)) + ((n_n4975) & (n_n4973) & (!n_n4971) & (x228x) & (n_n4972)) + ((n_n4975) & (n_n4973) & (n_n4971) & (!x228x) & (!n_n4972)) + ((n_n4975) & (n_n4973) & (n_n4971) & (!x228x) & (n_n4972)) + ((n_n4975) & (n_n4973) & (n_n4971) & (x228x) & (!n_n4972)) + ((n_n4975) & (n_n4973) & (n_n4971) & (x228x) & (n_n4972)));
	assign x141x = (((i_7_) & (!i_8_) & (i_6_) & (n_n535) & (x18x)) + ((i_7_) & (i_8_) & (i_6_) & (n_n535) & (x18x)));
	assign x317x = (((n_n260) & (!x20x) & (x23x) & (n_n464)) + ((n_n260) & (x20x) & (!x23x) & (n_n464)) + ((n_n260) & (x20x) & (x23x) & (n_n464)));
	assign n_n2973 = (((!n_n4828) & (!n_n4821) & (!x38x) & (!n_n3461) & (x326x)) + ((!n_n4828) & (!n_n4821) & (!x38x) & (n_n3461) & (!x326x)) + ((!n_n4828) & (!n_n4821) & (!x38x) & (n_n3461) & (x326x)) + ((!n_n4828) & (!n_n4821) & (x38x) & (!n_n3461) & (!x326x)) + ((!n_n4828) & (!n_n4821) & (x38x) & (!n_n3461) & (x326x)) + ((!n_n4828) & (!n_n4821) & (x38x) & (n_n3461) & (!x326x)) + ((!n_n4828) & (!n_n4821) & (x38x) & (n_n3461) & (x326x)) + ((!n_n4828) & (n_n4821) & (!x38x) & (!n_n3461) & (!x326x)) + ((!n_n4828) & (n_n4821) & (!x38x) & (!n_n3461) & (x326x)) + ((!n_n4828) & (n_n4821) & (!x38x) & (n_n3461) & (!x326x)) + ((!n_n4828) & (n_n4821) & (!x38x) & (n_n3461) & (x326x)) + ((!n_n4828) & (n_n4821) & (x38x) & (!n_n3461) & (!x326x)) + ((!n_n4828) & (n_n4821) & (x38x) & (!n_n3461) & (x326x)) + ((!n_n4828) & (n_n4821) & (x38x) & (n_n3461) & (!x326x)) + ((!n_n4828) & (n_n4821) & (x38x) & (n_n3461) & (x326x)) + ((n_n4828) & (!n_n4821) & (!x38x) & (!n_n3461) & (!x326x)) + ((n_n4828) & (!n_n4821) & (!x38x) & (!n_n3461) & (x326x)) + ((n_n4828) & (!n_n4821) & (!x38x) & (n_n3461) & (!x326x)) + ((n_n4828) & (!n_n4821) & (!x38x) & (n_n3461) & (x326x)) + ((n_n4828) & (!n_n4821) & (x38x) & (!n_n3461) & (!x326x)) + ((n_n4828) & (!n_n4821) & (x38x) & (!n_n3461) & (x326x)) + ((n_n4828) & (!n_n4821) & (x38x) & (n_n3461) & (!x326x)) + ((n_n4828) & (!n_n4821) & (x38x) & (n_n3461) & (x326x)) + ((n_n4828) & (n_n4821) & (!x38x) & (!n_n3461) & (!x326x)) + ((n_n4828) & (n_n4821) & (!x38x) & (!n_n3461) & (x326x)) + ((n_n4828) & (n_n4821) & (!x38x) & (n_n3461) & (!x326x)) + ((n_n4828) & (n_n4821) & (!x38x) & (n_n3461) & (x326x)) + ((n_n4828) & (n_n4821) & (x38x) & (!n_n3461) & (!x326x)) + ((n_n4828) & (n_n4821) & (x38x) & (!n_n3461) & (x326x)) + ((n_n4828) & (n_n4821) & (x38x) & (n_n3461) & (!x326x)) + ((n_n4828) & (n_n4821) & (x38x) & (n_n3461) & (x326x)));
	assign x375x = (((!i_9_) & (n_n524) & (n_n518) & (n_n260)) + ((i_9_) & (n_n524) & (n_n518) & (n_n260)));
	assign x15693x = (((!n_n4855) & (!n_n4849) & (!n_n4853) & (n_n4842)) + ((!n_n4855) & (!n_n4849) & (n_n4853) & (!n_n4842)) + ((!n_n4855) & (!n_n4849) & (n_n4853) & (n_n4842)) + ((!n_n4855) & (n_n4849) & (!n_n4853) & (!n_n4842)) + ((!n_n4855) & (n_n4849) & (!n_n4853) & (n_n4842)) + ((!n_n4855) & (n_n4849) & (n_n4853) & (!n_n4842)) + ((!n_n4855) & (n_n4849) & (n_n4853) & (n_n4842)) + ((n_n4855) & (!n_n4849) & (!n_n4853) & (!n_n4842)) + ((n_n4855) & (!n_n4849) & (!n_n4853) & (n_n4842)) + ((n_n4855) & (!n_n4849) & (n_n4853) & (!n_n4842)) + ((n_n4855) & (!n_n4849) & (n_n4853) & (n_n4842)) + ((n_n4855) & (n_n4849) & (!n_n4853) & (!n_n4842)) + ((n_n4855) & (n_n4849) & (!n_n4853) & (n_n4842)) + ((n_n4855) & (n_n4849) & (n_n4853) & (!n_n4842)) + ((n_n4855) & (n_n4849) & (n_n4853) & (n_n4842)));
	assign x15695x = (((!n_n4857) & (!n_n4856) & (!x176x) & (!x52x) & (x375x)) + ((!n_n4857) & (!n_n4856) & (!x176x) & (x52x) & (!x375x)) + ((!n_n4857) & (!n_n4856) & (!x176x) & (x52x) & (x375x)) + ((!n_n4857) & (!n_n4856) & (x176x) & (!x52x) & (!x375x)) + ((!n_n4857) & (!n_n4856) & (x176x) & (!x52x) & (x375x)) + ((!n_n4857) & (!n_n4856) & (x176x) & (x52x) & (!x375x)) + ((!n_n4857) & (!n_n4856) & (x176x) & (x52x) & (x375x)) + ((!n_n4857) & (n_n4856) & (!x176x) & (!x52x) & (!x375x)) + ((!n_n4857) & (n_n4856) & (!x176x) & (!x52x) & (x375x)) + ((!n_n4857) & (n_n4856) & (!x176x) & (x52x) & (!x375x)) + ((!n_n4857) & (n_n4856) & (!x176x) & (x52x) & (x375x)) + ((!n_n4857) & (n_n4856) & (x176x) & (!x52x) & (!x375x)) + ((!n_n4857) & (n_n4856) & (x176x) & (!x52x) & (x375x)) + ((!n_n4857) & (n_n4856) & (x176x) & (x52x) & (!x375x)) + ((!n_n4857) & (n_n4856) & (x176x) & (x52x) & (x375x)) + ((n_n4857) & (!n_n4856) & (!x176x) & (!x52x) & (!x375x)) + ((n_n4857) & (!n_n4856) & (!x176x) & (!x52x) & (x375x)) + ((n_n4857) & (!n_n4856) & (!x176x) & (x52x) & (!x375x)) + ((n_n4857) & (!n_n4856) & (!x176x) & (x52x) & (x375x)) + ((n_n4857) & (!n_n4856) & (x176x) & (!x52x) & (!x375x)) + ((n_n4857) & (!n_n4856) & (x176x) & (!x52x) & (x375x)) + ((n_n4857) & (!n_n4856) & (x176x) & (x52x) & (!x375x)) + ((n_n4857) & (!n_n4856) & (x176x) & (x52x) & (x375x)) + ((n_n4857) & (n_n4856) & (!x176x) & (!x52x) & (!x375x)) + ((n_n4857) & (n_n4856) & (!x176x) & (!x52x) & (x375x)) + ((n_n4857) & (n_n4856) & (!x176x) & (x52x) & (!x375x)) + ((n_n4857) & (n_n4856) & (!x176x) & (x52x) & (x375x)) + ((n_n4857) & (n_n4856) & (x176x) & (!x52x) & (!x375x)) + ((n_n4857) & (n_n4856) & (x176x) & (!x52x) & (x375x)) + ((n_n4857) & (n_n4856) & (x176x) & (x52x) & (!x375x)) + ((n_n4857) & (n_n4856) & (x176x) & (x52x) & (x375x)));
	assign x16632x = (((!n_n4628) & (!n_n4621) & (!n_n4619) & (!n_n4620) & (n_n4626)) + ((!n_n4628) & (!n_n4621) & (!n_n4619) & (n_n4620) & (!n_n4626)) + ((!n_n4628) & (!n_n4621) & (!n_n4619) & (n_n4620) & (n_n4626)) + ((!n_n4628) & (!n_n4621) & (n_n4619) & (!n_n4620) & (!n_n4626)) + ((!n_n4628) & (!n_n4621) & (n_n4619) & (!n_n4620) & (n_n4626)) + ((!n_n4628) & (!n_n4621) & (n_n4619) & (n_n4620) & (!n_n4626)) + ((!n_n4628) & (!n_n4621) & (n_n4619) & (n_n4620) & (n_n4626)) + ((!n_n4628) & (n_n4621) & (!n_n4619) & (!n_n4620) & (!n_n4626)) + ((!n_n4628) & (n_n4621) & (!n_n4619) & (!n_n4620) & (n_n4626)) + ((!n_n4628) & (n_n4621) & (!n_n4619) & (n_n4620) & (!n_n4626)) + ((!n_n4628) & (n_n4621) & (!n_n4619) & (n_n4620) & (n_n4626)) + ((!n_n4628) & (n_n4621) & (n_n4619) & (!n_n4620) & (!n_n4626)) + ((!n_n4628) & (n_n4621) & (n_n4619) & (!n_n4620) & (n_n4626)) + ((!n_n4628) & (n_n4621) & (n_n4619) & (n_n4620) & (!n_n4626)) + ((!n_n4628) & (n_n4621) & (n_n4619) & (n_n4620) & (n_n4626)) + ((n_n4628) & (!n_n4621) & (!n_n4619) & (!n_n4620) & (!n_n4626)) + ((n_n4628) & (!n_n4621) & (!n_n4619) & (!n_n4620) & (n_n4626)) + ((n_n4628) & (!n_n4621) & (!n_n4619) & (n_n4620) & (!n_n4626)) + ((n_n4628) & (!n_n4621) & (!n_n4619) & (n_n4620) & (n_n4626)) + ((n_n4628) & (!n_n4621) & (n_n4619) & (!n_n4620) & (!n_n4626)) + ((n_n4628) & (!n_n4621) & (n_n4619) & (!n_n4620) & (n_n4626)) + ((n_n4628) & (!n_n4621) & (n_n4619) & (n_n4620) & (!n_n4626)) + ((n_n4628) & (!n_n4621) & (n_n4619) & (n_n4620) & (n_n4626)) + ((n_n4628) & (n_n4621) & (!n_n4619) & (!n_n4620) & (!n_n4626)) + ((n_n4628) & (n_n4621) & (!n_n4619) & (!n_n4620) & (n_n4626)) + ((n_n4628) & (n_n4621) & (!n_n4619) & (n_n4620) & (!n_n4626)) + ((n_n4628) & (n_n4621) & (!n_n4619) & (n_n4620) & (n_n4626)) + ((n_n4628) & (n_n4621) & (n_n4619) & (!n_n4620) & (!n_n4626)) + ((n_n4628) & (n_n4621) & (n_n4619) & (!n_n4620) & (n_n4626)) + ((n_n4628) & (n_n4621) & (n_n4619) & (n_n4620) & (!n_n4626)) + ((n_n4628) & (n_n4621) & (n_n4619) & (n_n4620) & (n_n4626)));
	assign x190x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n390) & (n_n500)) + ((!i_9_) & (n_n524) & (!n_n526) & (n_n390) & (n_n500)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n390) & (n_n500)));
	assign x271x = (((!i_9_) & (!n_n528) & (n_n390) & (n_n491) & (n_n530)) + ((!i_9_) & (n_n528) & (n_n390) & (n_n491) & (n_n530)) + ((i_9_) & (n_n528) & (n_n390) & (n_n491) & (!n_n530)) + ((i_9_) & (n_n528) & (n_n390) & (n_n491) & (n_n530)));
	assign x12497x = (((!i_9_) & (n_n455) & (!n_n528) & (n_n473) & (n_n530)) + ((!i_9_) & (n_n455) & (n_n528) & (n_n473) & (!n_n530)) + ((!i_9_) & (n_n455) & (n_n528) & (n_n473) & (n_n530)) + ((i_9_) & (n_n455) & (!n_n528) & (n_n473) & (n_n530)) + ((i_9_) & (n_n455) & (n_n528) & (n_n473) & (!n_n530)) + ((i_9_) & (n_n455) & (n_n528) & (n_n473) & (n_n530)));
	assign n_n1491 = (((!n_n4547) & (!n_n4538) & (!x212x) & (!n_n4545) & (x12497x)) + ((!n_n4547) & (!n_n4538) & (!x212x) & (n_n4545) & (!x12497x)) + ((!n_n4547) & (!n_n4538) & (!x212x) & (n_n4545) & (x12497x)) + ((!n_n4547) & (!n_n4538) & (x212x) & (!n_n4545) & (!x12497x)) + ((!n_n4547) & (!n_n4538) & (x212x) & (!n_n4545) & (x12497x)) + ((!n_n4547) & (!n_n4538) & (x212x) & (n_n4545) & (!x12497x)) + ((!n_n4547) & (!n_n4538) & (x212x) & (n_n4545) & (x12497x)) + ((!n_n4547) & (n_n4538) & (!x212x) & (!n_n4545) & (!x12497x)) + ((!n_n4547) & (n_n4538) & (!x212x) & (!n_n4545) & (x12497x)) + ((!n_n4547) & (n_n4538) & (!x212x) & (n_n4545) & (!x12497x)) + ((!n_n4547) & (n_n4538) & (!x212x) & (n_n4545) & (x12497x)) + ((!n_n4547) & (n_n4538) & (x212x) & (!n_n4545) & (!x12497x)) + ((!n_n4547) & (n_n4538) & (x212x) & (!n_n4545) & (x12497x)) + ((!n_n4547) & (n_n4538) & (x212x) & (n_n4545) & (!x12497x)) + ((!n_n4547) & (n_n4538) & (x212x) & (n_n4545) & (x12497x)) + ((n_n4547) & (!n_n4538) & (!x212x) & (!n_n4545) & (!x12497x)) + ((n_n4547) & (!n_n4538) & (!x212x) & (!n_n4545) & (x12497x)) + ((n_n4547) & (!n_n4538) & (!x212x) & (n_n4545) & (!x12497x)) + ((n_n4547) & (!n_n4538) & (!x212x) & (n_n4545) & (x12497x)) + ((n_n4547) & (!n_n4538) & (x212x) & (!n_n4545) & (!x12497x)) + ((n_n4547) & (!n_n4538) & (x212x) & (!n_n4545) & (x12497x)) + ((n_n4547) & (!n_n4538) & (x212x) & (n_n4545) & (!x12497x)) + ((n_n4547) & (!n_n4538) & (x212x) & (n_n4545) & (x12497x)) + ((n_n4547) & (n_n4538) & (!x212x) & (!n_n4545) & (!x12497x)) + ((n_n4547) & (n_n4538) & (!x212x) & (!n_n4545) & (x12497x)) + ((n_n4547) & (n_n4538) & (!x212x) & (n_n4545) & (!x12497x)) + ((n_n4547) & (n_n4538) & (!x212x) & (n_n4545) & (x12497x)) + ((n_n4547) & (n_n4538) & (x212x) & (!n_n4545) & (!x12497x)) + ((n_n4547) & (n_n4538) & (x212x) & (!n_n4545) & (x12497x)) + ((n_n4547) & (n_n4538) & (x212x) & (n_n4545) & (!x12497x)) + ((n_n4547) & (n_n4538) & (x212x) & (n_n4545) & (x12497x)));
	assign x417x = (((!i_9_) & (n_n390) & (n_n473) & (!n_n520) & (x23x)) + ((!i_9_) & (n_n390) & (n_n473) & (n_n520) & (x23x)) + ((i_9_) & (n_n390) & (n_n473) & (!n_n520) & (x23x)) + ((i_9_) & (n_n390) & (n_n473) & (n_n520) & (!x23x)) + ((i_9_) & (n_n390) & (n_n473) & (n_n520) & (x23x)));
	assign x12418x = (((!i_9_) & (n_n526) & (!n_n528) & (n_n390) & (n_n473)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n390) & (n_n473)) + ((i_9_) & (!n_n526) & (n_n528) & (n_n390) & (n_n473)) + ((i_9_) & (n_n526) & (n_n528) & (n_n390) & (n_n473)));
	assign x12446x = (((!n_n4379) & (!n_n4378) & (!n_n4365) & (!n_n4374) & (n_n4370)) + ((!n_n4379) & (!n_n4378) & (!n_n4365) & (n_n4374) & (!n_n4370)) + ((!n_n4379) & (!n_n4378) & (!n_n4365) & (n_n4374) & (n_n4370)) + ((!n_n4379) & (!n_n4378) & (n_n4365) & (!n_n4374) & (!n_n4370)) + ((!n_n4379) & (!n_n4378) & (n_n4365) & (!n_n4374) & (n_n4370)) + ((!n_n4379) & (!n_n4378) & (n_n4365) & (n_n4374) & (!n_n4370)) + ((!n_n4379) & (!n_n4378) & (n_n4365) & (n_n4374) & (n_n4370)) + ((!n_n4379) & (n_n4378) & (!n_n4365) & (!n_n4374) & (!n_n4370)) + ((!n_n4379) & (n_n4378) & (!n_n4365) & (!n_n4374) & (n_n4370)) + ((!n_n4379) & (n_n4378) & (!n_n4365) & (n_n4374) & (!n_n4370)) + ((!n_n4379) & (n_n4378) & (!n_n4365) & (n_n4374) & (n_n4370)) + ((!n_n4379) & (n_n4378) & (n_n4365) & (!n_n4374) & (!n_n4370)) + ((!n_n4379) & (n_n4378) & (n_n4365) & (!n_n4374) & (n_n4370)) + ((!n_n4379) & (n_n4378) & (n_n4365) & (n_n4374) & (!n_n4370)) + ((!n_n4379) & (n_n4378) & (n_n4365) & (n_n4374) & (n_n4370)) + ((n_n4379) & (!n_n4378) & (!n_n4365) & (!n_n4374) & (!n_n4370)) + ((n_n4379) & (!n_n4378) & (!n_n4365) & (!n_n4374) & (n_n4370)) + ((n_n4379) & (!n_n4378) & (!n_n4365) & (n_n4374) & (!n_n4370)) + ((n_n4379) & (!n_n4378) & (!n_n4365) & (n_n4374) & (n_n4370)) + ((n_n4379) & (!n_n4378) & (n_n4365) & (!n_n4374) & (!n_n4370)) + ((n_n4379) & (!n_n4378) & (n_n4365) & (!n_n4374) & (n_n4370)) + ((n_n4379) & (!n_n4378) & (n_n4365) & (n_n4374) & (!n_n4370)) + ((n_n4379) & (!n_n4378) & (n_n4365) & (n_n4374) & (n_n4370)) + ((n_n4379) & (n_n4378) & (!n_n4365) & (!n_n4374) & (!n_n4370)) + ((n_n4379) & (n_n4378) & (!n_n4365) & (!n_n4374) & (n_n4370)) + ((n_n4379) & (n_n4378) & (!n_n4365) & (n_n4374) & (!n_n4370)) + ((n_n4379) & (n_n4378) & (!n_n4365) & (n_n4374) & (n_n4370)) + ((n_n4379) & (n_n4378) & (n_n4365) & (!n_n4374) & (!n_n4370)) + ((n_n4379) & (n_n4378) & (n_n4365) & (!n_n4374) & (n_n4370)) + ((n_n4379) & (n_n4378) & (n_n4365) & (n_n4374) & (!n_n4370)) + ((n_n4379) & (n_n4378) & (n_n4365) & (n_n4374) & (n_n4370)));
	assign n_n1504 = (((!n_n4373) & (!n_n4371) & (!x64x) & (x12446x)) + ((!n_n4373) & (!n_n4371) & (x64x) & (!x12446x)) + ((!n_n4373) & (!n_n4371) & (x64x) & (x12446x)) + ((!n_n4373) & (n_n4371) & (!x64x) & (!x12446x)) + ((!n_n4373) & (n_n4371) & (!x64x) & (x12446x)) + ((!n_n4373) & (n_n4371) & (x64x) & (!x12446x)) + ((!n_n4373) & (n_n4371) & (x64x) & (x12446x)) + ((n_n4373) & (!n_n4371) & (!x64x) & (!x12446x)) + ((n_n4373) & (!n_n4371) & (!x64x) & (x12446x)) + ((n_n4373) & (!n_n4371) & (x64x) & (!x12446x)) + ((n_n4373) & (!n_n4371) & (x64x) & (x12446x)) + ((n_n4373) & (n_n4371) & (!x64x) & (!x12446x)) + ((n_n4373) & (n_n4371) & (!x64x) & (x12446x)) + ((n_n4373) & (n_n4371) & (x64x) & (!x12446x)) + ((n_n4373) & (n_n4371) & (x64x) & (x12446x)));
	assign x12447x = (((!i_9_) & (n_n536) & (n_n526) & (n_n491)) + ((i_9_) & (n_n536) & (n_n526) & (n_n491)));
	assign n_n1693 = (((!n_n536) & (!x21x) & (!n_n491) & (!n_n4388) & (n_n4390)) + ((!n_n536) & (!x21x) & (!n_n491) & (n_n4388) & (!n_n4390)) + ((!n_n536) & (!x21x) & (!n_n491) & (n_n4388) & (n_n4390)) + ((!n_n536) & (!x21x) & (n_n491) & (!n_n4388) & (n_n4390)) + ((!n_n536) & (!x21x) & (n_n491) & (n_n4388) & (!n_n4390)) + ((!n_n536) & (!x21x) & (n_n491) & (n_n4388) & (n_n4390)) + ((!n_n536) & (x21x) & (!n_n491) & (!n_n4388) & (n_n4390)) + ((!n_n536) & (x21x) & (!n_n491) & (n_n4388) & (!n_n4390)) + ((!n_n536) & (x21x) & (!n_n491) & (n_n4388) & (n_n4390)) + ((!n_n536) & (x21x) & (n_n491) & (!n_n4388) & (n_n4390)) + ((!n_n536) & (x21x) & (n_n491) & (n_n4388) & (!n_n4390)) + ((!n_n536) & (x21x) & (n_n491) & (n_n4388) & (n_n4390)) + ((n_n536) & (!x21x) & (!n_n491) & (!n_n4388) & (n_n4390)) + ((n_n536) & (!x21x) & (!n_n491) & (n_n4388) & (!n_n4390)) + ((n_n536) & (!x21x) & (!n_n491) & (n_n4388) & (n_n4390)) + ((n_n536) & (!x21x) & (n_n491) & (!n_n4388) & (n_n4390)) + ((n_n536) & (!x21x) & (n_n491) & (n_n4388) & (!n_n4390)) + ((n_n536) & (!x21x) & (n_n491) & (n_n4388) & (n_n4390)) + ((n_n536) & (x21x) & (!n_n491) & (!n_n4388) & (n_n4390)) + ((n_n536) & (x21x) & (!n_n491) & (n_n4388) & (!n_n4390)) + ((n_n536) & (x21x) & (!n_n491) & (n_n4388) & (n_n4390)) + ((n_n536) & (x21x) & (n_n491) & (!n_n4388) & (!n_n4390)) + ((n_n536) & (x21x) & (n_n491) & (!n_n4388) & (n_n4390)) + ((n_n536) & (x21x) & (n_n491) & (n_n4388) & (!n_n4390)) + ((n_n536) & (x21x) & (n_n491) & (n_n4388) & (n_n4390)));
	assign x27x = (((!i_9_) & (n_n536) & (!n_n528) & (n_n491) & (n_n530)) + ((!i_9_) & (n_n536) & (n_n528) & (n_n491) & (n_n530)) + ((i_9_) & (n_n536) & (!n_n528) & (n_n491) & (n_n530)) + ((i_9_) & (n_n536) & (n_n528) & (n_n491) & (!n_n530)) + ((i_9_) & (n_n536) & (n_n528) & (n_n491) & (n_n530)));
	assign x12452x = (((!x25x) & (!n_n536) & (!n_n500) & (!n_n3533) & (n_n4348)) + ((!x25x) & (!n_n536) & (!n_n500) & (n_n3533) & (!n_n4348)) + ((!x25x) & (!n_n536) & (!n_n500) & (n_n3533) & (n_n4348)) + ((!x25x) & (!n_n536) & (n_n500) & (!n_n3533) & (n_n4348)) + ((!x25x) & (!n_n536) & (n_n500) & (n_n3533) & (!n_n4348)) + ((!x25x) & (!n_n536) & (n_n500) & (n_n3533) & (n_n4348)) + ((!x25x) & (n_n536) & (!n_n500) & (!n_n3533) & (n_n4348)) + ((!x25x) & (n_n536) & (!n_n500) & (n_n3533) & (!n_n4348)) + ((!x25x) & (n_n536) & (!n_n500) & (n_n3533) & (n_n4348)) + ((!x25x) & (n_n536) & (n_n500) & (!n_n3533) & (n_n4348)) + ((!x25x) & (n_n536) & (n_n500) & (n_n3533) & (!n_n4348)) + ((!x25x) & (n_n536) & (n_n500) & (n_n3533) & (n_n4348)) + ((x25x) & (!n_n536) & (!n_n500) & (!n_n3533) & (n_n4348)) + ((x25x) & (!n_n536) & (!n_n500) & (n_n3533) & (!n_n4348)) + ((x25x) & (!n_n536) & (!n_n500) & (n_n3533) & (n_n4348)) + ((x25x) & (!n_n536) & (n_n500) & (!n_n3533) & (n_n4348)) + ((x25x) & (!n_n536) & (n_n500) & (n_n3533) & (!n_n4348)) + ((x25x) & (!n_n536) & (n_n500) & (n_n3533) & (n_n4348)) + ((x25x) & (n_n536) & (!n_n500) & (!n_n3533) & (n_n4348)) + ((x25x) & (n_n536) & (!n_n500) & (n_n3533) & (!n_n4348)) + ((x25x) & (n_n536) & (!n_n500) & (n_n3533) & (n_n4348)) + ((x25x) & (n_n536) & (n_n500) & (!n_n3533) & (!n_n4348)) + ((x25x) & (n_n536) & (n_n500) & (!n_n3533) & (n_n4348)) + ((x25x) & (n_n536) & (n_n500) & (n_n3533) & (!n_n4348)) + ((x25x) & (n_n536) & (n_n500) & (n_n3533) & (n_n4348)));
	assign x12454x = (((!n_n4357) & (!n_n4358) & (!n_n4356) & (!n_n4355) & (x27x)) + ((!n_n4357) & (!n_n4358) & (!n_n4356) & (n_n4355) & (!x27x)) + ((!n_n4357) & (!n_n4358) & (!n_n4356) & (n_n4355) & (x27x)) + ((!n_n4357) & (!n_n4358) & (n_n4356) & (!n_n4355) & (!x27x)) + ((!n_n4357) & (!n_n4358) & (n_n4356) & (!n_n4355) & (x27x)) + ((!n_n4357) & (!n_n4358) & (n_n4356) & (n_n4355) & (!x27x)) + ((!n_n4357) & (!n_n4358) & (n_n4356) & (n_n4355) & (x27x)) + ((!n_n4357) & (n_n4358) & (!n_n4356) & (!n_n4355) & (!x27x)) + ((!n_n4357) & (n_n4358) & (!n_n4356) & (!n_n4355) & (x27x)) + ((!n_n4357) & (n_n4358) & (!n_n4356) & (n_n4355) & (!x27x)) + ((!n_n4357) & (n_n4358) & (!n_n4356) & (n_n4355) & (x27x)) + ((!n_n4357) & (n_n4358) & (n_n4356) & (!n_n4355) & (!x27x)) + ((!n_n4357) & (n_n4358) & (n_n4356) & (!n_n4355) & (x27x)) + ((!n_n4357) & (n_n4358) & (n_n4356) & (n_n4355) & (!x27x)) + ((!n_n4357) & (n_n4358) & (n_n4356) & (n_n4355) & (x27x)) + ((n_n4357) & (!n_n4358) & (!n_n4356) & (!n_n4355) & (!x27x)) + ((n_n4357) & (!n_n4358) & (!n_n4356) & (!n_n4355) & (x27x)) + ((n_n4357) & (!n_n4358) & (!n_n4356) & (n_n4355) & (!x27x)) + ((n_n4357) & (!n_n4358) & (!n_n4356) & (n_n4355) & (x27x)) + ((n_n4357) & (!n_n4358) & (n_n4356) & (!n_n4355) & (!x27x)) + ((n_n4357) & (!n_n4358) & (n_n4356) & (!n_n4355) & (x27x)) + ((n_n4357) & (!n_n4358) & (n_n4356) & (n_n4355) & (!x27x)) + ((n_n4357) & (!n_n4358) & (n_n4356) & (n_n4355) & (x27x)) + ((n_n4357) & (n_n4358) & (!n_n4356) & (!n_n4355) & (!x27x)) + ((n_n4357) & (n_n4358) & (!n_n4356) & (!n_n4355) & (x27x)) + ((n_n4357) & (n_n4358) & (!n_n4356) & (n_n4355) & (!x27x)) + ((n_n4357) & (n_n4358) & (!n_n4356) & (n_n4355) & (x27x)) + ((n_n4357) & (n_n4358) & (n_n4356) & (!n_n4355) & (!x27x)) + ((n_n4357) & (n_n4358) & (n_n4356) & (!n_n4355) & (x27x)) + ((n_n4357) & (n_n4358) & (n_n4356) & (n_n4355) & (!x27x)) + ((n_n4357) & (n_n4358) & (n_n4356) & (n_n4355) & (x27x)));
	assign x22147x = (((!n_n4784) & (!n_n4791) & (!n_n4787) & (!n_n4789)));
	assign x12269x = (((!i_9_) & (!n_n524) & (n_n130) & (n_n530) & (n_n464)) + ((!i_9_) & (n_n524) & (n_n130) & (!n_n530) & (n_n464)) + ((!i_9_) & (n_n524) & (n_n130) & (n_n530) & (n_n464)));
	assign x12270x = (((!i_7_) & (!i_8_) & (i_6_) & (x12x) & (n_n464)) + ((!i_7_) & (i_8_) & (i_6_) & (x12x) & (n_n464)) + ((i_7_) & (i_8_) & (i_6_) & (x12x) & (n_n464)));
	assign n_n1439 = (((!n_n5201) & (!n_n5199) & (!x453x) & (!x12269x) & (x12270x)) + ((!n_n5201) & (!n_n5199) & (!x453x) & (x12269x) & (!x12270x)) + ((!n_n5201) & (!n_n5199) & (!x453x) & (x12269x) & (x12270x)) + ((!n_n5201) & (!n_n5199) & (x453x) & (!x12269x) & (!x12270x)) + ((!n_n5201) & (!n_n5199) & (x453x) & (!x12269x) & (x12270x)) + ((!n_n5201) & (!n_n5199) & (x453x) & (x12269x) & (!x12270x)) + ((!n_n5201) & (!n_n5199) & (x453x) & (x12269x) & (x12270x)) + ((!n_n5201) & (n_n5199) & (!x453x) & (!x12269x) & (!x12270x)) + ((!n_n5201) & (n_n5199) & (!x453x) & (!x12269x) & (x12270x)) + ((!n_n5201) & (n_n5199) & (!x453x) & (x12269x) & (!x12270x)) + ((!n_n5201) & (n_n5199) & (!x453x) & (x12269x) & (x12270x)) + ((!n_n5201) & (n_n5199) & (x453x) & (!x12269x) & (!x12270x)) + ((!n_n5201) & (n_n5199) & (x453x) & (!x12269x) & (x12270x)) + ((!n_n5201) & (n_n5199) & (x453x) & (x12269x) & (!x12270x)) + ((!n_n5201) & (n_n5199) & (x453x) & (x12269x) & (x12270x)) + ((n_n5201) & (!n_n5199) & (!x453x) & (!x12269x) & (!x12270x)) + ((n_n5201) & (!n_n5199) & (!x453x) & (!x12269x) & (x12270x)) + ((n_n5201) & (!n_n5199) & (!x453x) & (x12269x) & (!x12270x)) + ((n_n5201) & (!n_n5199) & (!x453x) & (x12269x) & (x12270x)) + ((n_n5201) & (!n_n5199) & (x453x) & (!x12269x) & (!x12270x)) + ((n_n5201) & (!n_n5199) & (x453x) & (!x12269x) & (x12270x)) + ((n_n5201) & (!n_n5199) & (x453x) & (x12269x) & (!x12270x)) + ((n_n5201) & (!n_n5199) & (x453x) & (x12269x) & (x12270x)) + ((n_n5201) & (n_n5199) & (!x453x) & (!x12269x) & (!x12270x)) + ((n_n5201) & (n_n5199) & (!x453x) & (!x12269x) & (x12270x)) + ((n_n5201) & (n_n5199) & (!x453x) & (x12269x) & (!x12270x)) + ((n_n5201) & (n_n5199) & (!x453x) & (x12269x) & (x12270x)) + ((n_n5201) & (n_n5199) & (x453x) & (!x12269x) & (!x12270x)) + ((n_n5201) & (n_n5199) & (x453x) & (!x12269x) & (x12270x)) + ((n_n5201) & (n_n5199) & (x453x) & (x12269x) & (!x12270x)) + ((n_n5201) & (n_n5199) & (x453x) & (x12269x) & (x12270x)));
	assign x450x = (((!n_n130) & (!x23x) & (!n_n464) & (n_n5208)) + ((!n_n130) & (!x23x) & (n_n464) & (n_n5208)) + ((!n_n130) & (x23x) & (!n_n464) & (n_n5208)) + ((!n_n130) & (x23x) & (n_n464) & (n_n5208)) + ((n_n130) & (!x23x) & (!n_n464) & (n_n5208)) + ((n_n130) & (!x23x) & (n_n464) & (n_n5208)) + ((n_n130) & (x23x) & (!n_n464) & (n_n5208)) + ((n_n130) & (x23x) & (n_n464) & (!n_n5208)) + ((n_n130) & (x23x) & (n_n464) & (n_n5208)));
	assign x12278x = (((!n_n5230) & (!n_n5223) & (!n_n5233) & (n_n5220)) + ((!n_n5230) & (!n_n5223) & (n_n5233) & (!n_n5220)) + ((!n_n5230) & (!n_n5223) & (n_n5233) & (n_n5220)) + ((!n_n5230) & (n_n5223) & (!n_n5233) & (!n_n5220)) + ((!n_n5230) & (n_n5223) & (!n_n5233) & (n_n5220)) + ((!n_n5230) & (n_n5223) & (n_n5233) & (!n_n5220)) + ((!n_n5230) & (n_n5223) & (n_n5233) & (n_n5220)) + ((n_n5230) & (!n_n5223) & (!n_n5233) & (!n_n5220)) + ((n_n5230) & (!n_n5223) & (!n_n5233) & (n_n5220)) + ((n_n5230) & (!n_n5223) & (n_n5233) & (!n_n5220)) + ((n_n5230) & (!n_n5223) & (n_n5233) & (n_n5220)) + ((n_n5230) & (n_n5223) & (!n_n5233) & (!n_n5220)) + ((n_n5230) & (n_n5223) & (!n_n5233) & (n_n5220)) + ((n_n5230) & (n_n5223) & (n_n5233) & (!n_n5220)) + ((n_n5230) & (n_n5223) & (n_n5233) & (n_n5220)));
	assign x12280x = (((!n_n5217) & (!n_n5218) & (!n_n5215) & (!x223x) & (n_n5213)) + ((!n_n5217) & (!n_n5218) & (!n_n5215) & (x223x) & (!n_n5213)) + ((!n_n5217) & (!n_n5218) & (!n_n5215) & (x223x) & (n_n5213)) + ((!n_n5217) & (!n_n5218) & (n_n5215) & (!x223x) & (!n_n5213)) + ((!n_n5217) & (!n_n5218) & (n_n5215) & (!x223x) & (n_n5213)) + ((!n_n5217) & (!n_n5218) & (n_n5215) & (x223x) & (!n_n5213)) + ((!n_n5217) & (!n_n5218) & (n_n5215) & (x223x) & (n_n5213)) + ((!n_n5217) & (n_n5218) & (!n_n5215) & (!x223x) & (!n_n5213)) + ((!n_n5217) & (n_n5218) & (!n_n5215) & (!x223x) & (n_n5213)) + ((!n_n5217) & (n_n5218) & (!n_n5215) & (x223x) & (!n_n5213)) + ((!n_n5217) & (n_n5218) & (!n_n5215) & (x223x) & (n_n5213)) + ((!n_n5217) & (n_n5218) & (n_n5215) & (!x223x) & (!n_n5213)) + ((!n_n5217) & (n_n5218) & (n_n5215) & (!x223x) & (n_n5213)) + ((!n_n5217) & (n_n5218) & (n_n5215) & (x223x) & (!n_n5213)) + ((!n_n5217) & (n_n5218) & (n_n5215) & (x223x) & (n_n5213)) + ((n_n5217) & (!n_n5218) & (!n_n5215) & (!x223x) & (!n_n5213)) + ((n_n5217) & (!n_n5218) & (!n_n5215) & (!x223x) & (n_n5213)) + ((n_n5217) & (!n_n5218) & (!n_n5215) & (x223x) & (!n_n5213)) + ((n_n5217) & (!n_n5218) & (!n_n5215) & (x223x) & (n_n5213)) + ((n_n5217) & (!n_n5218) & (n_n5215) & (!x223x) & (!n_n5213)) + ((n_n5217) & (!n_n5218) & (n_n5215) & (!x223x) & (n_n5213)) + ((n_n5217) & (!n_n5218) & (n_n5215) & (x223x) & (!n_n5213)) + ((n_n5217) & (!n_n5218) & (n_n5215) & (x223x) & (n_n5213)) + ((n_n5217) & (n_n5218) & (!n_n5215) & (!x223x) & (!n_n5213)) + ((n_n5217) & (n_n5218) & (!n_n5215) & (!x223x) & (n_n5213)) + ((n_n5217) & (n_n5218) & (!n_n5215) & (x223x) & (!n_n5213)) + ((n_n5217) & (n_n5218) & (!n_n5215) & (x223x) & (n_n5213)) + ((n_n5217) & (n_n5218) & (n_n5215) & (!x223x) & (!n_n5213)) + ((n_n5217) & (n_n5218) & (n_n5215) & (!x223x) & (n_n5213)) + ((n_n5217) & (n_n5218) & (n_n5215) & (x223x) & (!n_n5213)) + ((n_n5217) & (n_n5218) & (n_n5215) & (x223x) & (n_n5213)));
	assign x22145x = (((!n_n5234) & (!n_n1530) & (!n_n5219) & (!n_n5205) & (!x450x)));
	assign n_n1405 = (((!n_n1439) & (!x12278x) & (!x12280x) & (!x22145x)) + ((!n_n1439) & (!x12278x) & (x12280x) & (!x22145x)) + ((!n_n1439) & (!x12278x) & (x12280x) & (x22145x)) + ((!n_n1439) & (x12278x) & (!x12280x) & (!x22145x)) + ((!n_n1439) & (x12278x) & (!x12280x) & (x22145x)) + ((!n_n1439) & (x12278x) & (x12280x) & (!x22145x)) + ((!n_n1439) & (x12278x) & (x12280x) & (x22145x)) + ((n_n1439) & (!x12278x) & (!x12280x) & (!x22145x)) + ((n_n1439) & (!x12278x) & (!x12280x) & (x22145x)) + ((n_n1439) & (!x12278x) & (x12280x) & (!x22145x)) + ((n_n1439) & (!x12278x) & (x12280x) & (x22145x)) + ((n_n1439) & (x12278x) & (!x12280x) & (!x22145x)) + ((n_n1439) & (x12278x) & (!x12280x) & (x22145x)) + ((n_n1439) & (x12278x) & (x12280x) & (!x22145x)) + ((n_n1439) & (x12278x) & (x12280x) & (x22145x)));
	assign x22181x = (((!n_n5171) & (!n_n5174) & (!n_n5186) & (!n_n5175) & (!n_n5176)));
	assign x12296x = (((!n_n5187) & (!n_n5177) & (!n_n4129) & (!x22181x)) + ((!n_n5187) & (!n_n5177) & (n_n4129) & (!x22181x)) + ((!n_n5187) & (!n_n5177) & (n_n4129) & (x22181x)) + ((!n_n5187) & (n_n5177) & (!n_n4129) & (!x22181x)) + ((!n_n5187) & (n_n5177) & (!n_n4129) & (x22181x)) + ((!n_n5187) & (n_n5177) & (n_n4129) & (!x22181x)) + ((!n_n5187) & (n_n5177) & (n_n4129) & (x22181x)) + ((n_n5187) & (!n_n5177) & (!n_n4129) & (!x22181x)) + ((n_n5187) & (!n_n5177) & (!n_n4129) & (x22181x)) + ((n_n5187) & (!n_n5177) & (n_n4129) & (!x22181x)) + ((n_n5187) & (!n_n5177) & (n_n4129) & (x22181x)) + ((n_n5187) & (n_n5177) & (!n_n4129) & (!x22181x)) + ((n_n5187) & (n_n5177) & (!n_n4129) & (x22181x)) + ((n_n5187) & (n_n5177) & (n_n4129) & (!x22181x)) + ((n_n5187) & (n_n5177) & (n_n4129) & (x22181x)));
	assign x286x = (((!i_9_) & (!n_n524) & (n_n509) & (n_n130) & (x20x)) + ((!i_9_) & (n_n524) & (n_n509) & (n_n130) & (!x20x)) + ((!i_9_) & (n_n524) & (n_n509) & (n_n130) & (x20x)) + ((i_9_) & (!n_n524) & (n_n509) & (n_n130) & (x20x)) + ((i_9_) & (n_n524) & (n_n509) & (n_n130) & (x20x)));
	assign x12301x = (((!n_n5130) & (!n_n5123) & (!n_n5120) & (n_n5125)) + ((!n_n5130) & (!n_n5123) & (n_n5120) & (!n_n5125)) + ((!n_n5130) & (!n_n5123) & (n_n5120) & (n_n5125)) + ((!n_n5130) & (n_n5123) & (!n_n5120) & (!n_n5125)) + ((!n_n5130) & (n_n5123) & (!n_n5120) & (n_n5125)) + ((!n_n5130) & (n_n5123) & (n_n5120) & (!n_n5125)) + ((!n_n5130) & (n_n5123) & (n_n5120) & (n_n5125)) + ((n_n5130) & (!n_n5123) & (!n_n5120) & (!n_n5125)) + ((n_n5130) & (!n_n5123) & (!n_n5120) & (n_n5125)) + ((n_n5130) & (!n_n5123) & (n_n5120) & (!n_n5125)) + ((n_n5130) & (!n_n5123) & (n_n5120) & (n_n5125)) + ((n_n5130) & (n_n5123) & (!n_n5120) & (!n_n5125)) + ((n_n5130) & (n_n5123) & (!n_n5120) & (n_n5125)) + ((n_n5130) & (n_n5123) & (n_n5120) & (!n_n5125)) + ((n_n5130) & (n_n5123) & (n_n5120) & (n_n5125)));
	assign x12302x = (((!n_n5127) & (!n_n5121) & (!n_n5122) & (!n_n5132) & (n_n5128)) + ((!n_n5127) & (!n_n5121) & (!n_n5122) & (n_n5132) & (!n_n5128)) + ((!n_n5127) & (!n_n5121) & (!n_n5122) & (n_n5132) & (n_n5128)) + ((!n_n5127) & (!n_n5121) & (n_n5122) & (!n_n5132) & (!n_n5128)) + ((!n_n5127) & (!n_n5121) & (n_n5122) & (!n_n5132) & (n_n5128)) + ((!n_n5127) & (!n_n5121) & (n_n5122) & (n_n5132) & (!n_n5128)) + ((!n_n5127) & (!n_n5121) & (n_n5122) & (n_n5132) & (n_n5128)) + ((!n_n5127) & (n_n5121) & (!n_n5122) & (!n_n5132) & (!n_n5128)) + ((!n_n5127) & (n_n5121) & (!n_n5122) & (!n_n5132) & (n_n5128)) + ((!n_n5127) & (n_n5121) & (!n_n5122) & (n_n5132) & (!n_n5128)) + ((!n_n5127) & (n_n5121) & (!n_n5122) & (n_n5132) & (n_n5128)) + ((!n_n5127) & (n_n5121) & (n_n5122) & (!n_n5132) & (!n_n5128)) + ((!n_n5127) & (n_n5121) & (n_n5122) & (!n_n5132) & (n_n5128)) + ((!n_n5127) & (n_n5121) & (n_n5122) & (n_n5132) & (!n_n5128)) + ((!n_n5127) & (n_n5121) & (n_n5122) & (n_n5132) & (n_n5128)) + ((n_n5127) & (!n_n5121) & (!n_n5122) & (!n_n5132) & (!n_n5128)) + ((n_n5127) & (!n_n5121) & (!n_n5122) & (!n_n5132) & (n_n5128)) + ((n_n5127) & (!n_n5121) & (!n_n5122) & (n_n5132) & (!n_n5128)) + ((n_n5127) & (!n_n5121) & (!n_n5122) & (n_n5132) & (n_n5128)) + ((n_n5127) & (!n_n5121) & (n_n5122) & (!n_n5132) & (!n_n5128)) + ((n_n5127) & (!n_n5121) & (n_n5122) & (!n_n5132) & (n_n5128)) + ((n_n5127) & (!n_n5121) & (n_n5122) & (n_n5132) & (!n_n5128)) + ((n_n5127) & (!n_n5121) & (n_n5122) & (n_n5132) & (n_n5128)) + ((n_n5127) & (n_n5121) & (!n_n5122) & (!n_n5132) & (!n_n5128)) + ((n_n5127) & (n_n5121) & (!n_n5122) & (!n_n5132) & (n_n5128)) + ((n_n5127) & (n_n5121) & (!n_n5122) & (n_n5132) & (!n_n5128)) + ((n_n5127) & (n_n5121) & (!n_n5122) & (n_n5132) & (n_n5128)) + ((n_n5127) & (n_n5121) & (n_n5122) & (!n_n5132) & (!n_n5128)) + ((n_n5127) & (n_n5121) & (n_n5122) & (!n_n5132) & (n_n5128)) + ((n_n5127) & (n_n5121) & (n_n5122) & (n_n5132) & (!n_n5128)) + ((n_n5127) & (n_n5121) & (n_n5122) & (n_n5132) & (n_n5128)));
	assign x12305x = (((!n_n1443) & (!n_n1444) & (!x12301x) & (x12302x)) + ((!n_n1443) & (!n_n1444) & (x12301x) & (!x12302x)) + ((!n_n1443) & (!n_n1444) & (x12301x) & (x12302x)) + ((!n_n1443) & (n_n1444) & (!x12301x) & (!x12302x)) + ((!n_n1443) & (n_n1444) & (!x12301x) & (x12302x)) + ((!n_n1443) & (n_n1444) & (x12301x) & (!x12302x)) + ((!n_n1443) & (n_n1444) & (x12301x) & (x12302x)) + ((n_n1443) & (!n_n1444) & (!x12301x) & (!x12302x)) + ((n_n1443) & (!n_n1444) & (!x12301x) & (x12302x)) + ((n_n1443) & (!n_n1444) & (x12301x) & (!x12302x)) + ((n_n1443) & (!n_n1444) & (x12301x) & (x12302x)) + ((n_n1443) & (n_n1444) & (!x12301x) & (!x12302x)) + ((n_n1443) & (n_n1444) & (!x12301x) & (x12302x)) + ((n_n1443) & (n_n1444) & (x12301x) & (!x12302x)) + ((n_n1443) & (n_n1444) & (x12301x) & (x12302x)));
	assign x12295x = (((!n_n5179) & (!n_n5178) & (!x113x) & (!x332x) & (x188x)) + ((!n_n5179) & (!n_n5178) & (!x113x) & (x332x) & (!x188x)) + ((!n_n5179) & (!n_n5178) & (!x113x) & (x332x) & (x188x)) + ((!n_n5179) & (!n_n5178) & (x113x) & (!x332x) & (!x188x)) + ((!n_n5179) & (!n_n5178) & (x113x) & (!x332x) & (x188x)) + ((!n_n5179) & (!n_n5178) & (x113x) & (x332x) & (!x188x)) + ((!n_n5179) & (!n_n5178) & (x113x) & (x332x) & (x188x)) + ((!n_n5179) & (n_n5178) & (!x113x) & (!x332x) & (!x188x)) + ((!n_n5179) & (n_n5178) & (!x113x) & (!x332x) & (x188x)) + ((!n_n5179) & (n_n5178) & (!x113x) & (x332x) & (!x188x)) + ((!n_n5179) & (n_n5178) & (!x113x) & (x332x) & (x188x)) + ((!n_n5179) & (n_n5178) & (x113x) & (!x332x) & (!x188x)) + ((!n_n5179) & (n_n5178) & (x113x) & (!x332x) & (x188x)) + ((!n_n5179) & (n_n5178) & (x113x) & (x332x) & (!x188x)) + ((!n_n5179) & (n_n5178) & (x113x) & (x332x) & (x188x)) + ((n_n5179) & (!n_n5178) & (!x113x) & (!x332x) & (!x188x)) + ((n_n5179) & (!n_n5178) & (!x113x) & (!x332x) & (x188x)) + ((n_n5179) & (!n_n5178) & (!x113x) & (x332x) & (!x188x)) + ((n_n5179) & (!n_n5178) & (!x113x) & (x332x) & (x188x)) + ((n_n5179) & (!n_n5178) & (x113x) & (!x332x) & (!x188x)) + ((n_n5179) & (!n_n5178) & (x113x) & (!x332x) & (x188x)) + ((n_n5179) & (!n_n5178) & (x113x) & (x332x) & (!x188x)) + ((n_n5179) & (!n_n5178) & (x113x) & (x332x) & (x188x)) + ((n_n5179) & (n_n5178) & (!x113x) & (!x332x) & (!x188x)) + ((n_n5179) & (n_n5178) & (!x113x) & (!x332x) & (x188x)) + ((n_n5179) & (n_n5178) & (!x113x) & (x332x) & (!x188x)) + ((n_n5179) & (n_n5178) & (!x113x) & (x332x) & (x188x)) + ((n_n5179) & (n_n5178) & (x113x) & (!x332x) & (!x188x)) + ((n_n5179) & (n_n5178) & (x113x) & (!x332x) & (x188x)) + ((n_n5179) & (n_n5178) & (x113x) & (x332x) & (!x188x)) + ((n_n5179) & (n_n5178) & (x113x) & (x332x) & (x188x)));
	assign x22144x = (((!n_n4430) & (!n_n4404) & (!n_n4409) & (!n_n4417)));
	assign n_n1341 = (((!n_n4420) & (!n_n4407) & (!x84x) & (!n_n4410) & (!x22144x)) + ((!n_n4420) & (!n_n4407) & (!x84x) & (n_n4410) & (!x22144x)) + ((!n_n4420) & (!n_n4407) & (!x84x) & (n_n4410) & (x22144x)) + ((!n_n4420) & (!n_n4407) & (x84x) & (!n_n4410) & (!x22144x)) + ((!n_n4420) & (!n_n4407) & (x84x) & (!n_n4410) & (x22144x)) + ((!n_n4420) & (!n_n4407) & (x84x) & (n_n4410) & (!x22144x)) + ((!n_n4420) & (!n_n4407) & (x84x) & (n_n4410) & (x22144x)) + ((!n_n4420) & (n_n4407) & (!x84x) & (!n_n4410) & (!x22144x)) + ((!n_n4420) & (n_n4407) & (!x84x) & (!n_n4410) & (x22144x)) + ((!n_n4420) & (n_n4407) & (!x84x) & (n_n4410) & (!x22144x)) + ((!n_n4420) & (n_n4407) & (!x84x) & (n_n4410) & (x22144x)) + ((!n_n4420) & (n_n4407) & (x84x) & (!n_n4410) & (!x22144x)) + ((!n_n4420) & (n_n4407) & (x84x) & (!n_n4410) & (x22144x)) + ((!n_n4420) & (n_n4407) & (x84x) & (n_n4410) & (!x22144x)) + ((!n_n4420) & (n_n4407) & (x84x) & (n_n4410) & (x22144x)) + ((n_n4420) & (!n_n4407) & (!x84x) & (!n_n4410) & (!x22144x)) + ((n_n4420) & (!n_n4407) & (!x84x) & (!n_n4410) & (x22144x)) + ((n_n4420) & (!n_n4407) & (!x84x) & (n_n4410) & (!x22144x)) + ((n_n4420) & (!n_n4407) & (!x84x) & (n_n4410) & (x22144x)) + ((n_n4420) & (!n_n4407) & (x84x) & (!n_n4410) & (!x22144x)) + ((n_n4420) & (!n_n4407) & (x84x) & (!n_n4410) & (x22144x)) + ((n_n4420) & (!n_n4407) & (x84x) & (n_n4410) & (!x22144x)) + ((n_n4420) & (!n_n4407) & (x84x) & (n_n4410) & (x22144x)) + ((n_n4420) & (n_n4407) & (!x84x) & (!n_n4410) & (!x22144x)) + ((n_n4420) & (n_n4407) & (!x84x) & (!n_n4410) & (x22144x)) + ((n_n4420) & (n_n4407) & (!x84x) & (n_n4410) & (!x22144x)) + ((n_n4420) & (n_n4407) & (!x84x) & (n_n4410) & (x22144x)) + ((n_n4420) & (n_n4407) & (x84x) & (!n_n4410) & (!x22144x)) + ((n_n4420) & (n_n4407) & (x84x) & (!n_n4410) & (x22144x)) + ((n_n4420) & (n_n4407) & (x84x) & (n_n4410) & (!x22144x)) + ((n_n4420) & (n_n4407) & (x84x) & (n_n4410) & (x22144x)));
	assign x12141x = (((!x25x) & (!n_n536) & (!n_n509) & (!n_n4340) & (x399x)) + ((!x25x) & (!n_n536) & (!n_n509) & (n_n4340) & (!x399x)) + ((!x25x) & (!n_n536) & (!n_n509) & (n_n4340) & (x399x)) + ((!x25x) & (!n_n536) & (n_n509) & (!n_n4340) & (x399x)) + ((!x25x) & (!n_n536) & (n_n509) & (n_n4340) & (!x399x)) + ((!x25x) & (!n_n536) & (n_n509) & (n_n4340) & (x399x)) + ((!x25x) & (n_n536) & (!n_n509) & (!n_n4340) & (x399x)) + ((!x25x) & (n_n536) & (!n_n509) & (n_n4340) & (!x399x)) + ((!x25x) & (n_n536) & (!n_n509) & (n_n4340) & (x399x)) + ((!x25x) & (n_n536) & (n_n509) & (!n_n4340) & (x399x)) + ((!x25x) & (n_n536) & (n_n509) & (n_n4340) & (!x399x)) + ((!x25x) & (n_n536) & (n_n509) & (n_n4340) & (x399x)) + ((x25x) & (!n_n536) & (!n_n509) & (!n_n4340) & (x399x)) + ((x25x) & (!n_n536) & (!n_n509) & (n_n4340) & (!x399x)) + ((x25x) & (!n_n536) & (!n_n509) & (n_n4340) & (x399x)) + ((x25x) & (!n_n536) & (n_n509) & (!n_n4340) & (x399x)) + ((x25x) & (!n_n536) & (n_n509) & (n_n4340) & (!x399x)) + ((x25x) & (!n_n536) & (n_n509) & (n_n4340) & (x399x)) + ((x25x) & (n_n536) & (!n_n509) & (!n_n4340) & (x399x)) + ((x25x) & (n_n536) & (!n_n509) & (n_n4340) & (!x399x)) + ((x25x) & (n_n536) & (!n_n509) & (n_n4340) & (x399x)) + ((x25x) & (n_n536) & (n_n509) & (!n_n4340) & (!x399x)) + ((x25x) & (n_n536) & (n_n509) & (!n_n4340) & (x399x)) + ((x25x) & (n_n536) & (n_n509) & (n_n4340) & (!x399x)) + ((x25x) & (n_n536) & (n_n509) & (n_n4340) & (x399x)));
	assign x12142x = (((!n_n4343) & (!n_n4312) & (!n_n4326) & (!n_n4342) & (n_n4331)) + ((!n_n4343) & (!n_n4312) & (!n_n4326) & (n_n4342) & (!n_n4331)) + ((!n_n4343) & (!n_n4312) & (!n_n4326) & (n_n4342) & (n_n4331)) + ((!n_n4343) & (!n_n4312) & (n_n4326) & (!n_n4342) & (!n_n4331)) + ((!n_n4343) & (!n_n4312) & (n_n4326) & (!n_n4342) & (n_n4331)) + ((!n_n4343) & (!n_n4312) & (n_n4326) & (n_n4342) & (!n_n4331)) + ((!n_n4343) & (!n_n4312) & (n_n4326) & (n_n4342) & (n_n4331)) + ((!n_n4343) & (n_n4312) & (!n_n4326) & (!n_n4342) & (!n_n4331)) + ((!n_n4343) & (n_n4312) & (!n_n4326) & (!n_n4342) & (n_n4331)) + ((!n_n4343) & (n_n4312) & (!n_n4326) & (n_n4342) & (!n_n4331)) + ((!n_n4343) & (n_n4312) & (!n_n4326) & (n_n4342) & (n_n4331)) + ((!n_n4343) & (n_n4312) & (n_n4326) & (!n_n4342) & (!n_n4331)) + ((!n_n4343) & (n_n4312) & (n_n4326) & (!n_n4342) & (n_n4331)) + ((!n_n4343) & (n_n4312) & (n_n4326) & (n_n4342) & (!n_n4331)) + ((!n_n4343) & (n_n4312) & (n_n4326) & (n_n4342) & (n_n4331)) + ((n_n4343) & (!n_n4312) & (!n_n4326) & (!n_n4342) & (!n_n4331)) + ((n_n4343) & (!n_n4312) & (!n_n4326) & (!n_n4342) & (n_n4331)) + ((n_n4343) & (!n_n4312) & (!n_n4326) & (n_n4342) & (!n_n4331)) + ((n_n4343) & (!n_n4312) & (!n_n4326) & (n_n4342) & (n_n4331)) + ((n_n4343) & (!n_n4312) & (n_n4326) & (!n_n4342) & (!n_n4331)) + ((n_n4343) & (!n_n4312) & (n_n4326) & (!n_n4342) & (n_n4331)) + ((n_n4343) & (!n_n4312) & (n_n4326) & (n_n4342) & (!n_n4331)) + ((n_n4343) & (!n_n4312) & (n_n4326) & (n_n4342) & (n_n4331)) + ((n_n4343) & (n_n4312) & (!n_n4326) & (!n_n4342) & (!n_n4331)) + ((n_n4343) & (n_n4312) & (!n_n4326) & (!n_n4342) & (n_n4331)) + ((n_n4343) & (n_n4312) & (!n_n4326) & (n_n4342) & (!n_n4331)) + ((n_n4343) & (n_n4312) & (!n_n4326) & (n_n4342) & (n_n4331)) + ((n_n4343) & (n_n4312) & (n_n4326) & (!n_n4342) & (!n_n4331)) + ((n_n4343) & (n_n4312) & (n_n4326) & (!n_n4342) & (n_n4331)) + ((n_n4343) & (n_n4312) & (n_n4326) & (n_n4342) & (!n_n4331)) + ((n_n4343) & (n_n4312) & (n_n4326) & (n_n4342) & (n_n4331)));
	assign x11675x = (((!n_n4781) & (!n_n4797) & (!n_n4801) & (n_n4778)) + ((!n_n4781) & (!n_n4797) & (n_n4801) & (!n_n4778)) + ((!n_n4781) & (!n_n4797) & (n_n4801) & (n_n4778)) + ((!n_n4781) & (n_n4797) & (!n_n4801) & (!n_n4778)) + ((!n_n4781) & (n_n4797) & (!n_n4801) & (n_n4778)) + ((!n_n4781) & (n_n4797) & (n_n4801) & (!n_n4778)) + ((!n_n4781) & (n_n4797) & (n_n4801) & (n_n4778)) + ((n_n4781) & (!n_n4797) & (!n_n4801) & (!n_n4778)) + ((n_n4781) & (!n_n4797) & (!n_n4801) & (n_n4778)) + ((n_n4781) & (!n_n4797) & (n_n4801) & (!n_n4778)) + ((n_n4781) & (!n_n4797) & (n_n4801) & (n_n4778)) + ((n_n4781) & (n_n4797) & (!n_n4801) & (!n_n4778)) + ((n_n4781) & (n_n4797) & (!n_n4801) & (n_n4778)) + ((n_n4781) & (n_n4797) & (n_n4801) & (!n_n4778)) + ((n_n4781) & (n_n4797) & (n_n4801) & (n_n4778)));
	assign x11676x = (((!n_n4817) & (!n_n4823) & (!n_n4742) & (!n_n4773) & (n_n4813)) + ((!n_n4817) & (!n_n4823) & (!n_n4742) & (n_n4773) & (!n_n4813)) + ((!n_n4817) & (!n_n4823) & (!n_n4742) & (n_n4773) & (n_n4813)) + ((!n_n4817) & (!n_n4823) & (n_n4742) & (!n_n4773) & (!n_n4813)) + ((!n_n4817) & (!n_n4823) & (n_n4742) & (!n_n4773) & (n_n4813)) + ((!n_n4817) & (!n_n4823) & (n_n4742) & (n_n4773) & (!n_n4813)) + ((!n_n4817) & (!n_n4823) & (n_n4742) & (n_n4773) & (n_n4813)) + ((!n_n4817) & (n_n4823) & (!n_n4742) & (!n_n4773) & (!n_n4813)) + ((!n_n4817) & (n_n4823) & (!n_n4742) & (!n_n4773) & (n_n4813)) + ((!n_n4817) & (n_n4823) & (!n_n4742) & (n_n4773) & (!n_n4813)) + ((!n_n4817) & (n_n4823) & (!n_n4742) & (n_n4773) & (n_n4813)) + ((!n_n4817) & (n_n4823) & (n_n4742) & (!n_n4773) & (!n_n4813)) + ((!n_n4817) & (n_n4823) & (n_n4742) & (!n_n4773) & (n_n4813)) + ((!n_n4817) & (n_n4823) & (n_n4742) & (n_n4773) & (!n_n4813)) + ((!n_n4817) & (n_n4823) & (n_n4742) & (n_n4773) & (n_n4813)) + ((n_n4817) & (!n_n4823) & (!n_n4742) & (!n_n4773) & (!n_n4813)) + ((n_n4817) & (!n_n4823) & (!n_n4742) & (!n_n4773) & (n_n4813)) + ((n_n4817) & (!n_n4823) & (!n_n4742) & (n_n4773) & (!n_n4813)) + ((n_n4817) & (!n_n4823) & (!n_n4742) & (n_n4773) & (n_n4813)) + ((n_n4817) & (!n_n4823) & (n_n4742) & (!n_n4773) & (!n_n4813)) + ((n_n4817) & (!n_n4823) & (n_n4742) & (!n_n4773) & (n_n4813)) + ((n_n4817) & (!n_n4823) & (n_n4742) & (n_n4773) & (!n_n4813)) + ((n_n4817) & (!n_n4823) & (n_n4742) & (n_n4773) & (n_n4813)) + ((n_n4817) & (n_n4823) & (!n_n4742) & (!n_n4773) & (!n_n4813)) + ((n_n4817) & (n_n4823) & (!n_n4742) & (!n_n4773) & (n_n4813)) + ((n_n4817) & (n_n4823) & (!n_n4742) & (n_n4773) & (!n_n4813)) + ((n_n4817) & (n_n4823) & (!n_n4742) & (n_n4773) & (n_n4813)) + ((n_n4817) & (n_n4823) & (n_n4742) & (!n_n4773) & (!n_n4813)) + ((n_n4817) & (n_n4823) & (n_n4742) & (!n_n4773) & (n_n4813)) + ((n_n4817) & (n_n4823) & (n_n4742) & (n_n4773) & (!n_n4813)) + ((n_n4817) & (n_n4823) & (n_n4742) & (n_n4773) & (n_n4813)));
	assign x12873x = (((!n_n5244) & (!n_n5241) & (!n_n5242) & (!n_n5243) & (n_n5234)) + ((!n_n5244) & (!n_n5241) & (!n_n5242) & (n_n5243) & (!n_n5234)) + ((!n_n5244) & (!n_n5241) & (!n_n5242) & (n_n5243) & (n_n5234)) + ((!n_n5244) & (!n_n5241) & (n_n5242) & (!n_n5243) & (!n_n5234)) + ((!n_n5244) & (!n_n5241) & (n_n5242) & (!n_n5243) & (n_n5234)) + ((!n_n5244) & (!n_n5241) & (n_n5242) & (n_n5243) & (!n_n5234)) + ((!n_n5244) & (!n_n5241) & (n_n5242) & (n_n5243) & (n_n5234)) + ((!n_n5244) & (n_n5241) & (!n_n5242) & (!n_n5243) & (!n_n5234)) + ((!n_n5244) & (n_n5241) & (!n_n5242) & (!n_n5243) & (n_n5234)) + ((!n_n5244) & (n_n5241) & (!n_n5242) & (n_n5243) & (!n_n5234)) + ((!n_n5244) & (n_n5241) & (!n_n5242) & (n_n5243) & (n_n5234)) + ((!n_n5244) & (n_n5241) & (n_n5242) & (!n_n5243) & (!n_n5234)) + ((!n_n5244) & (n_n5241) & (n_n5242) & (!n_n5243) & (n_n5234)) + ((!n_n5244) & (n_n5241) & (n_n5242) & (n_n5243) & (!n_n5234)) + ((!n_n5244) & (n_n5241) & (n_n5242) & (n_n5243) & (n_n5234)) + ((n_n5244) & (!n_n5241) & (!n_n5242) & (!n_n5243) & (!n_n5234)) + ((n_n5244) & (!n_n5241) & (!n_n5242) & (!n_n5243) & (n_n5234)) + ((n_n5244) & (!n_n5241) & (!n_n5242) & (n_n5243) & (!n_n5234)) + ((n_n5244) & (!n_n5241) & (!n_n5242) & (n_n5243) & (n_n5234)) + ((n_n5244) & (!n_n5241) & (n_n5242) & (!n_n5243) & (!n_n5234)) + ((n_n5244) & (!n_n5241) & (n_n5242) & (!n_n5243) & (n_n5234)) + ((n_n5244) & (!n_n5241) & (n_n5242) & (n_n5243) & (!n_n5234)) + ((n_n5244) & (!n_n5241) & (n_n5242) & (n_n5243) & (n_n5234)) + ((n_n5244) & (n_n5241) & (!n_n5242) & (!n_n5243) & (!n_n5234)) + ((n_n5244) & (n_n5241) & (!n_n5242) & (!n_n5243) & (n_n5234)) + ((n_n5244) & (n_n5241) & (!n_n5242) & (n_n5243) & (!n_n5234)) + ((n_n5244) & (n_n5241) & (!n_n5242) & (n_n5243) & (n_n5234)) + ((n_n5244) & (n_n5241) & (n_n5242) & (!n_n5243) & (!n_n5234)) + ((n_n5244) & (n_n5241) & (n_n5242) & (!n_n5243) & (n_n5234)) + ((n_n5244) & (n_n5241) & (n_n5242) & (n_n5243) & (!n_n5234)) + ((n_n5244) & (n_n5241) & (n_n5242) & (n_n5243) & (n_n5234)));
	assign n_n667 = (((!n_n5240) & (!n_n5238) & (!n_n5247) & (!n_n5246) & (x12873x)) + ((!n_n5240) & (!n_n5238) & (!n_n5247) & (n_n5246) & (!x12873x)) + ((!n_n5240) & (!n_n5238) & (!n_n5247) & (n_n5246) & (x12873x)) + ((!n_n5240) & (!n_n5238) & (n_n5247) & (!n_n5246) & (!x12873x)) + ((!n_n5240) & (!n_n5238) & (n_n5247) & (!n_n5246) & (x12873x)) + ((!n_n5240) & (!n_n5238) & (n_n5247) & (n_n5246) & (!x12873x)) + ((!n_n5240) & (!n_n5238) & (n_n5247) & (n_n5246) & (x12873x)) + ((!n_n5240) & (n_n5238) & (!n_n5247) & (!n_n5246) & (!x12873x)) + ((!n_n5240) & (n_n5238) & (!n_n5247) & (!n_n5246) & (x12873x)) + ((!n_n5240) & (n_n5238) & (!n_n5247) & (n_n5246) & (!x12873x)) + ((!n_n5240) & (n_n5238) & (!n_n5247) & (n_n5246) & (x12873x)) + ((!n_n5240) & (n_n5238) & (n_n5247) & (!n_n5246) & (!x12873x)) + ((!n_n5240) & (n_n5238) & (n_n5247) & (!n_n5246) & (x12873x)) + ((!n_n5240) & (n_n5238) & (n_n5247) & (n_n5246) & (!x12873x)) + ((!n_n5240) & (n_n5238) & (n_n5247) & (n_n5246) & (x12873x)) + ((n_n5240) & (!n_n5238) & (!n_n5247) & (!n_n5246) & (!x12873x)) + ((n_n5240) & (!n_n5238) & (!n_n5247) & (!n_n5246) & (x12873x)) + ((n_n5240) & (!n_n5238) & (!n_n5247) & (n_n5246) & (!x12873x)) + ((n_n5240) & (!n_n5238) & (!n_n5247) & (n_n5246) & (x12873x)) + ((n_n5240) & (!n_n5238) & (n_n5247) & (!n_n5246) & (!x12873x)) + ((n_n5240) & (!n_n5238) & (n_n5247) & (!n_n5246) & (x12873x)) + ((n_n5240) & (!n_n5238) & (n_n5247) & (n_n5246) & (!x12873x)) + ((n_n5240) & (!n_n5238) & (n_n5247) & (n_n5246) & (x12873x)) + ((n_n5240) & (n_n5238) & (!n_n5247) & (!n_n5246) & (!x12873x)) + ((n_n5240) & (n_n5238) & (!n_n5247) & (!n_n5246) & (x12873x)) + ((n_n5240) & (n_n5238) & (!n_n5247) & (n_n5246) & (!x12873x)) + ((n_n5240) & (n_n5238) & (!n_n5247) & (n_n5246) & (x12873x)) + ((n_n5240) & (n_n5238) & (n_n5247) & (!n_n5246) & (!x12873x)) + ((n_n5240) & (n_n5238) & (n_n5247) & (!n_n5246) & (x12873x)) + ((n_n5240) & (n_n5238) & (n_n5247) & (n_n5246) & (!x12873x)) + ((n_n5240) & (n_n5238) & (n_n5247) & (n_n5246) & (x12873x)));
	assign n_n761 = (((!x19x) & (!n_n535) & (!n_n520) & (!n_n5223) & (n_n5224)) + ((!x19x) & (!n_n535) & (!n_n520) & (n_n5223) & (!n_n5224)) + ((!x19x) & (!n_n535) & (!n_n520) & (n_n5223) & (n_n5224)) + ((!x19x) & (!n_n535) & (n_n520) & (!n_n5223) & (n_n5224)) + ((!x19x) & (!n_n535) & (n_n520) & (n_n5223) & (!n_n5224)) + ((!x19x) & (!n_n535) & (n_n520) & (n_n5223) & (n_n5224)) + ((!x19x) & (n_n535) & (!n_n520) & (!n_n5223) & (n_n5224)) + ((!x19x) & (n_n535) & (!n_n520) & (n_n5223) & (!n_n5224)) + ((!x19x) & (n_n535) & (!n_n520) & (n_n5223) & (n_n5224)) + ((!x19x) & (n_n535) & (n_n520) & (!n_n5223) & (n_n5224)) + ((!x19x) & (n_n535) & (n_n520) & (n_n5223) & (!n_n5224)) + ((!x19x) & (n_n535) & (n_n520) & (n_n5223) & (n_n5224)) + ((x19x) & (!n_n535) & (!n_n520) & (!n_n5223) & (n_n5224)) + ((x19x) & (!n_n535) & (!n_n520) & (n_n5223) & (!n_n5224)) + ((x19x) & (!n_n535) & (!n_n520) & (n_n5223) & (n_n5224)) + ((x19x) & (!n_n535) & (n_n520) & (!n_n5223) & (n_n5224)) + ((x19x) & (!n_n535) & (n_n520) & (n_n5223) & (!n_n5224)) + ((x19x) & (!n_n535) & (n_n520) & (n_n5223) & (n_n5224)) + ((x19x) & (n_n535) & (!n_n520) & (!n_n5223) & (n_n5224)) + ((x19x) & (n_n535) & (!n_n520) & (n_n5223) & (!n_n5224)) + ((x19x) & (n_n535) & (!n_n520) & (n_n5223) & (n_n5224)) + ((x19x) & (n_n535) & (n_n520) & (!n_n5223) & (!n_n5224)) + ((x19x) & (n_n535) & (n_n520) & (!n_n5223) & (n_n5224)) + ((x19x) & (n_n535) & (n_n520) & (n_n5223) & (!n_n5224)) + ((x19x) & (n_n535) & (n_n520) & (n_n5223) & (n_n5224)));
	assign x12878x = (((!n_n5229) & (!n_n5220) & (!x223x) & (n_n5208)) + ((!n_n5229) & (!n_n5220) & (x223x) & (!n_n5208)) + ((!n_n5229) & (!n_n5220) & (x223x) & (n_n5208)) + ((!n_n5229) & (n_n5220) & (!x223x) & (!n_n5208)) + ((!n_n5229) & (n_n5220) & (!x223x) & (n_n5208)) + ((!n_n5229) & (n_n5220) & (x223x) & (!n_n5208)) + ((!n_n5229) & (n_n5220) & (x223x) & (n_n5208)) + ((n_n5229) & (!n_n5220) & (!x223x) & (!n_n5208)) + ((n_n5229) & (!n_n5220) & (!x223x) & (n_n5208)) + ((n_n5229) & (!n_n5220) & (x223x) & (!n_n5208)) + ((n_n5229) & (!n_n5220) & (x223x) & (n_n5208)) + ((n_n5229) & (n_n5220) & (!x223x) & (!n_n5208)) + ((n_n5229) & (n_n5220) & (!x223x) & (n_n5208)) + ((n_n5229) & (n_n5220) & (x223x) & (!n_n5208)) + ((n_n5229) & (n_n5220) & (x223x) & (n_n5208)));
	assign x12879x = (((!n_n5217) & (!n_n5218) & (!n_n5215) & (n_n761)) + ((!n_n5217) & (!n_n5218) & (n_n5215) & (!n_n761)) + ((!n_n5217) & (!n_n5218) & (n_n5215) & (n_n761)) + ((!n_n5217) & (n_n5218) & (!n_n5215) & (!n_n761)) + ((!n_n5217) & (n_n5218) & (!n_n5215) & (n_n761)) + ((!n_n5217) & (n_n5218) & (n_n5215) & (!n_n761)) + ((!n_n5217) & (n_n5218) & (n_n5215) & (n_n761)) + ((n_n5217) & (!n_n5218) & (!n_n5215) & (!n_n761)) + ((n_n5217) & (!n_n5218) & (!n_n5215) & (n_n761)) + ((n_n5217) & (!n_n5218) & (n_n5215) & (!n_n761)) + ((n_n5217) & (!n_n5218) & (n_n5215) & (n_n761)) + ((n_n5217) & (n_n5218) & (!n_n5215) & (!n_n761)) + ((n_n5217) & (n_n5218) & (!n_n5215) & (n_n761)) + ((n_n5217) & (n_n5218) & (n_n5215) & (!n_n761)) + ((n_n5217) & (n_n5218) & (n_n5215) & (n_n761)));
	assign x12880x = (((!n_n5232) & (!n_n5233) & (!n_n5226) & (!x383x) & (x183x)) + ((!n_n5232) & (!n_n5233) & (!n_n5226) & (x383x) & (!x183x)) + ((!n_n5232) & (!n_n5233) & (!n_n5226) & (x383x) & (x183x)) + ((!n_n5232) & (!n_n5233) & (n_n5226) & (!x383x) & (!x183x)) + ((!n_n5232) & (!n_n5233) & (n_n5226) & (!x383x) & (x183x)) + ((!n_n5232) & (!n_n5233) & (n_n5226) & (x383x) & (!x183x)) + ((!n_n5232) & (!n_n5233) & (n_n5226) & (x383x) & (x183x)) + ((!n_n5232) & (n_n5233) & (!n_n5226) & (!x383x) & (!x183x)) + ((!n_n5232) & (n_n5233) & (!n_n5226) & (!x383x) & (x183x)) + ((!n_n5232) & (n_n5233) & (!n_n5226) & (x383x) & (!x183x)) + ((!n_n5232) & (n_n5233) & (!n_n5226) & (x383x) & (x183x)) + ((!n_n5232) & (n_n5233) & (n_n5226) & (!x383x) & (!x183x)) + ((!n_n5232) & (n_n5233) & (n_n5226) & (!x383x) & (x183x)) + ((!n_n5232) & (n_n5233) & (n_n5226) & (x383x) & (!x183x)) + ((!n_n5232) & (n_n5233) & (n_n5226) & (x383x) & (x183x)) + ((n_n5232) & (!n_n5233) & (!n_n5226) & (!x383x) & (!x183x)) + ((n_n5232) & (!n_n5233) & (!n_n5226) & (!x383x) & (x183x)) + ((n_n5232) & (!n_n5233) & (!n_n5226) & (x383x) & (!x183x)) + ((n_n5232) & (!n_n5233) & (!n_n5226) & (x383x) & (x183x)) + ((n_n5232) & (!n_n5233) & (n_n5226) & (!x383x) & (!x183x)) + ((n_n5232) & (!n_n5233) & (n_n5226) & (!x383x) & (x183x)) + ((n_n5232) & (!n_n5233) & (n_n5226) & (x383x) & (!x183x)) + ((n_n5232) & (!n_n5233) & (n_n5226) & (x383x) & (x183x)) + ((n_n5232) & (n_n5233) & (!n_n5226) & (!x383x) & (!x183x)) + ((n_n5232) & (n_n5233) & (!n_n5226) & (!x383x) & (x183x)) + ((n_n5232) & (n_n5233) & (!n_n5226) & (x383x) & (!x183x)) + ((n_n5232) & (n_n5233) & (!n_n5226) & (x383x) & (x183x)) + ((n_n5232) & (n_n5233) & (n_n5226) & (!x383x) & (!x183x)) + ((n_n5232) & (n_n5233) & (n_n5226) & (!x383x) & (x183x)) + ((n_n5232) & (n_n5233) & (n_n5226) & (x383x) & (!x183x)) + ((n_n5232) & (n_n5233) & (n_n5226) & (x383x) & (x183x)));
	assign n_n635 = (((!n_n667) & (!x12878x) & (!x12879x) & (x12880x)) + ((!n_n667) & (!x12878x) & (x12879x) & (!x12880x)) + ((!n_n667) & (!x12878x) & (x12879x) & (x12880x)) + ((!n_n667) & (x12878x) & (!x12879x) & (!x12880x)) + ((!n_n667) & (x12878x) & (!x12879x) & (x12880x)) + ((!n_n667) & (x12878x) & (x12879x) & (!x12880x)) + ((!n_n667) & (x12878x) & (x12879x) & (x12880x)) + ((n_n667) & (!x12878x) & (!x12879x) & (!x12880x)) + ((n_n667) & (!x12878x) & (!x12879x) & (x12880x)) + ((n_n667) & (!x12878x) & (x12879x) & (!x12880x)) + ((n_n667) & (!x12878x) & (x12879x) & (x12880x)) + ((n_n667) & (x12878x) & (!x12879x) & (!x12880x)) + ((n_n667) & (x12878x) & (!x12879x) & (x12880x)) + ((n_n667) & (x12878x) & (x12879x) & (!x12880x)) + ((n_n667) & (x12878x) & (x12879x) & (x12880x)));
	assign x12884x = (((!i_9_) & (n_n524) & (n_n130) & (n_n500)) + ((i_9_) & (n_n524) & (n_n130) & (n_n500)));
	assign n_n777 = (((!n_n522) & (!x12x) & (!n_n500) & (x12884x)) + ((!n_n522) & (!x12x) & (n_n500) & (x12884x)) + ((!n_n522) & (x12x) & (!n_n500) & (x12884x)) + ((!n_n522) & (x12x) & (n_n500) & (x12884x)) + ((n_n522) & (!x12x) & (!n_n500) & (x12884x)) + ((n_n522) & (!x12x) & (n_n500) & (x12884x)) + ((n_n522) & (x12x) & (!n_n500) & (x12884x)) + ((n_n522) & (x12x) & (n_n500) & (!x12884x)) + ((n_n522) & (x12x) & (n_n500) & (x12884x)));
	assign n_n3772 = (((!n_n532) & (!x12x) & (!n_n500) & (x155x)) + ((!n_n532) & (!x12x) & (n_n500) & (x155x)) + ((!n_n532) & (x12x) & (!n_n500) & (x155x)) + ((!n_n532) & (x12x) & (n_n500) & (x155x)) + ((n_n532) & (!x12x) & (!n_n500) & (x155x)) + ((n_n532) & (!x12x) & (n_n500) & (x155x)) + ((n_n532) & (x12x) & (!n_n500) & (x155x)) + ((n_n532) & (x12x) & (n_n500) & (!x155x)) + ((n_n532) & (x12x) & (n_n500) & (x155x)));
	assign x12889x = (((!n_n5156) & (!n_n5163) & (!n_n5157) & (!n_n5159) & (n_n5169)) + ((!n_n5156) & (!n_n5163) & (!n_n5157) & (n_n5159) & (!n_n5169)) + ((!n_n5156) & (!n_n5163) & (!n_n5157) & (n_n5159) & (n_n5169)) + ((!n_n5156) & (!n_n5163) & (n_n5157) & (!n_n5159) & (!n_n5169)) + ((!n_n5156) & (!n_n5163) & (n_n5157) & (!n_n5159) & (n_n5169)) + ((!n_n5156) & (!n_n5163) & (n_n5157) & (n_n5159) & (!n_n5169)) + ((!n_n5156) & (!n_n5163) & (n_n5157) & (n_n5159) & (n_n5169)) + ((!n_n5156) & (n_n5163) & (!n_n5157) & (!n_n5159) & (!n_n5169)) + ((!n_n5156) & (n_n5163) & (!n_n5157) & (!n_n5159) & (n_n5169)) + ((!n_n5156) & (n_n5163) & (!n_n5157) & (n_n5159) & (!n_n5169)) + ((!n_n5156) & (n_n5163) & (!n_n5157) & (n_n5159) & (n_n5169)) + ((!n_n5156) & (n_n5163) & (n_n5157) & (!n_n5159) & (!n_n5169)) + ((!n_n5156) & (n_n5163) & (n_n5157) & (!n_n5159) & (n_n5169)) + ((!n_n5156) & (n_n5163) & (n_n5157) & (n_n5159) & (!n_n5169)) + ((!n_n5156) & (n_n5163) & (n_n5157) & (n_n5159) & (n_n5169)) + ((n_n5156) & (!n_n5163) & (!n_n5157) & (!n_n5159) & (!n_n5169)) + ((n_n5156) & (!n_n5163) & (!n_n5157) & (!n_n5159) & (n_n5169)) + ((n_n5156) & (!n_n5163) & (!n_n5157) & (n_n5159) & (!n_n5169)) + ((n_n5156) & (!n_n5163) & (!n_n5157) & (n_n5159) & (n_n5169)) + ((n_n5156) & (!n_n5163) & (n_n5157) & (!n_n5159) & (!n_n5169)) + ((n_n5156) & (!n_n5163) & (n_n5157) & (!n_n5159) & (n_n5169)) + ((n_n5156) & (!n_n5163) & (n_n5157) & (n_n5159) & (!n_n5169)) + ((n_n5156) & (!n_n5163) & (n_n5157) & (n_n5159) & (n_n5169)) + ((n_n5156) & (n_n5163) & (!n_n5157) & (!n_n5159) & (!n_n5169)) + ((n_n5156) & (n_n5163) & (!n_n5157) & (!n_n5159) & (n_n5169)) + ((n_n5156) & (n_n5163) & (!n_n5157) & (n_n5159) & (!n_n5169)) + ((n_n5156) & (n_n5163) & (!n_n5157) & (n_n5159) & (n_n5169)) + ((n_n5156) & (n_n5163) & (n_n5157) & (!n_n5159) & (!n_n5169)) + ((n_n5156) & (n_n5163) & (n_n5157) & (!n_n5159) & (n_n5169)) + ((n_n5156) & (n_n5163) & (n_n5157) & (n_n5159) & (!n_n5169)) + ((n_n5156) & (n_n5163) & (n_n5157) & (n_n5159) & (n_n5169)));
	assign x12897x = (((!n_n5148) & (!n_n5153) & (!n_n3771) & (!n_n777) & (n_n3772)) + ((!n_n5148) & (!n_n5153) & (!n_n3771) & (n_n777) & (!n_n3772)) + ((!n_n5148) & (!n_n5153) & (!n_n3771) & (n_n777) & (n_n3772)) + ((!n_n5148) & (!n_n5153) & (n_n3771) & (!n_n777) & (!n_n3772)) + ((!n_n5148) & (!n_n5153) & (n_n3771) & (!n_n777) & (n_n3772)) + ((!n_n5148) & (!n_n5153) & (n_n3771) & (n_n777) & (!n_n3772)) + ((!n_n5148) & (!n_n5153) & (n_n3771) & (n_n777) & (n_n3772)) + ((!n_n5148) & (n_n5153) & (!n_n3771) & (!n_n777) & (!n_n3772)) + ((!n_n5148) & (n_n5153) & (!n_n3771) & (!n_n777) & (n_n3772)) + ((!n_n5148) & (n_n5153) & (!n_n3771) & (n_n777) & (!n_n3772)) + ((!n_n5148) & (n_n5153) & (!n_n3771) & (n_n777) & (n_n3772)) + ((!n_n5148) & (n_n5153) & (n_n3771) & (!n_n777) & (!n_n3772)) + ((!n_n5148) & (n_n5153) & (n_n3771) & (!n_n777) & (n_n3772)) + ((!n_n5148) & (n_n5153) & (n_n3771) & (n_n777) & (!n_n3772)) + ((!n_n5148) & (n_n5153) & (n_n3771) & (n_n777) & (n_n3772)) + ((n_n5148) & (!n_n5153) & (!n_n3771) & (!n_n777) & (!n_n3772)) + ((n_n5148) & (!n_n5153) & (!n_n3771) & (!n_n777) & (n_n3772)) + ((n_n5148) & (!n_n5153) & (!n_n3771) & (n_n777) & (!n_n3772)) + ((n_n5148) & (!n_n5153) & (!n_n3771) & (n_n777) & (n_n3772)) + ((n_n5148) & (!n_n5153) & (n_n3771) & (!n_n777) & (!n_n3772)) + ((n_n5148) & (!n_n5153) & (n_n3771) & (!n_n777) & (n_n3772)) + ((n_n5148) & (!n_n5153) & (n_n3771) & (n_n777) & (!n_n3772)) + ((n_n5148) & (!n_n5153) & (n_n3771) & (n_n777) & (n_n3772)) + ((n_n5148) & (n_n5153) & (!n_n3771) & (!n_n777) & (!n_n3772)) + ((n_n5148) & (n_n5153) & (!n_n3771) & (!n_n777) & (n_n3772)) + ((n_n5148) & (n_n5153) & (!n_n3771) & (n_n777) & (!n_n3772)) + ((n_n5148) & (n_n5153) & (!n_n3771) & (n_n777) & (n_n3772)) + ((n_n5148) & (n_n5153) & (n_n3771) & (!n_n777) & (!n_n3772)) + ((n_n5148) & (n_n5153) & (n_n3771) & (!n_n777) & (n_n3772)) + ((n_n5148) & (n_n5153) & (n_n3771) & (n_n777) & (!n_n3772)) + ((n_n5148) & (n_n5153) & (n_n3771) & (n_n777) & (n_n3772)));
	assign x12896x = (((!n_n5150) & (!n_n5149) & (!x126x) & (!n_n5144) & (x407x)) + ((!n_n5150) & (!n_n5149) & (!x126x) & (n_n5144) & (!x407x)) + ((!n_n5150) & (!n_n5149) & (!x126x) & (n_n5144) & (x407x)) + ((!n_n5150) & (!n_n5149) & (x126x) & (!n_n5144) & (!x407x)) + ((!n_n5150) & (!n_n5149) & (x126x) & (!n_n5144) & (x407x)) + ((!n_n5150) & (!n_n5149) & (x126x) & (n_n5144) & (!x407x)) + ((!n_n5150) & (!n_n5149) & (x126x) & (n_n5144) & (x407x)) + ((!n_n5150) & (n_n5149) & (!x126x) & (!n_n5144) & (!x407x)) + ((!n_n5150) & (n_n5149) & (!x126x) & (!n_n5144) & (x407x)) + ((!n_n5150) & (n_n5149) & (!x126x) & (n_n5144) & (!x407x)) + ((!n_n5150) & (n_n5149) & (!x126x) & (n_n5144) & (x407x)) + ((!n_n5150) & (n_n5149) & (x126x) & (!n_n5144) & (!x407x)) + ((!n_n5150) & (n_n5149) & (x126x) & (!n_n5144) & (x407x)) + ((!n_n5150) & (n_n5149) & (x126x) & (n_n5144) & (!x407x)) + ((!n_n5150) & (n_n5149) & (x126x) & (n_n5144) & (x407x)) + ((n_n5150) & (!n_n5149) & (!x126x) & (!n_n5144) & (!x407x)) + ((n_n5150) & (!n_n5149) & (!x126x) & (!n_n5144) & (x407x)) + ((n_n5150) & (!n_n5149) & (!x126x) & (n_n5144) & (!x407x)) + ((n_n5150) & (!n_n5149) & (!x126x) & (n_n5144) & (x407x)) + ((n_n5150) & (!n_n5149) & (x126x) & (!n_n5144) & (!x407x)) + ((n_n5150) & (!n_n5149) & (x126x) & (!n_n5144) & (x407x)) + ((n_n5150) & (!n_n5149) & (x126x) & (n_n5144) & (!x407x)) + ((n_n5150) & (!n_n5149) & (x126x) & (n_n5144) & (x407x)) + ((n_n5150) & (n_n5149) & (!x126x) & (!n_n5144) & (!x407x)) + ((n_n5150) & (n_n5149) & (!x126x) & (!n_n5144) & (x407x)) + ((n_n5150) & (n_n5149) & (!x126x) & (n_n5144) & (!x407x)) + ((n_n5150) & (n_n5149) & (!x126x) & (n_n5144) & (x407x)) + ((n_n5150) & (n_n5149) & (x126x) & (!n_n5144) & (!x407x)) + ((n_n5150) & (n_n5149) & (x126x) & (!n_n5144) & (x407x)) + ((n_n5150) & (n_n5149) & (x126x) & (n_n5144) & (!x407x)) + ((n_n5150) & (n_n5149) & (x126x) & (n_n5144) & (x407x)));
	assign x22203x = (((!n_n5167) & (!n_n5161) & (!n_n5162) & (!n_n5160)));
	assign n_n637 = (((!x12889x) & (!x12897x) & (!x12896x) & (!x22203x)) + ((!x12889x) & (!x12897x) & (x12896x) & (!x22203x)) + ((!x12889x) & (!x12897x) & (x12896x) & (x22203x)) + ((!x12889x) & (x12897x) & (!x12896x) & (!x22203x)) + ((!x12889x) & (x12897x) & (!x12896x) & (x22203x)) + ((!x12889x) & (x12897x) & (x12896x) & (!x22203x)) + ((!x12889x) & (x12897x) & (x12896x) & (x22203x)) + ((x12889x) & (!x12897x) & (!x12896x) & (!x22203x)) + ((x12889x) & (!x12897x) & (!x12896x) & (x22203x)) + ((x12889x) & (!x12897x) & (x12896x) & (!x22203x)) + ((x12889x) & (!x12897x) & (x12896x) & (x22203x)) + ((x12889x) & (x12897x) & (!x12896x) & (!x22203x)) + ((x12889x) & (x12897x) & (!x12896x) & (x22203x)) + ((x12889x) & (x12897x) & (x12896x) & (!x22203x)) + ((x12889x) & (x12897x) & (x12896x) & (x22203x)));
	assign x12647x = (((!n_n5165) & (!n_n5117) & (!n_n5135) & (n_n5158)) + ((!n_n5165) & (!n_n5117) & (n_n5135) & (!n_n5158)) + ((!n_n5165) & (!n_n5117) & (n_n5135) & (n_n5158)) + ((!n_n5165) & (n_n5117) & (!n_n5135) & (!n_n5158)) + ((!n_n5165) & (n_n5117) & (!n_n5135) & (n_n5158)) + ((!n_n5165) & (n_n5117) & (n_n5135) & (!n_n5158)) + ((!n_n5165) & (n_n5117) & (n_n5135) & (n_n5158)) + ((n_n5165) & (!n_n5117) & (!n_n5135) & (!n_n5158)) + ((n_n5165) & (!n_n5117) & (!n_n5135) & (n_n5158)) + ((n_n5165) & (!n_n5117) & (n_n5135) & (!n_n5158)) + ((n_n5165) & (!n_n5117) & (n_n5135) & (n_n5158)) + ((n_n5165) & (n_n5117) & (!n_n5135) & (!n_n5158)) + ((n_n5165) & (n_n5117) & (!n_n5135) & (n_n5158)) + ((n_n5165) & (n_n5117) & (n_n5135) & (!n_n5158)) + ((n_n5165) & (n_n5117) & (n_n5135) & (n_n5158)));
	assign x12648x = (((!n_n5123) & (!n_n5155) & (!n_n5121) & (!n_n5151) & (n_n5134)) + ((!n_n5123) & (!n_n5155) & (!n_n5121) & (n_n5151) & (!n_n5134)) + ((!n_n5123) & (!n_n5155) & (!n_n5121) & (n_n5151) & (n_n5134)) + ((!n_n5123) & (!n_n5155) & (n_n5121) & (!n_n5151) & (!n_n5134)) + ((!n_n5123) & (!n_n5155) & (n_n5121) & (!n_n5151) & (n_n5134)) + ((!n_n5123) & (!n_n5155) & (n_n5121) & (n_n5151) & (!n_n5134)) + ((!n_n5123) & (!n_n5155) & (n_n5121) & (n_n5151) & (n_n5134)) + ((!n_n5123) & (n_n5155) & (!n_n5121) & (!n_n5151) & (!n_n5134)) + ((!n_n5123) & (n_n5155) & (!n_n5121) & (!n_n5151) & (n_n5134)) + ((!n_n5123) & (n_n5155) & (!n_n5121) & (n_n5151) & (!n_n5134)) + ((!n_n5123) & (n_n5155) & (!n_n5121) & (n_n5151) & (n_n5134)) + ((!n_n5123) & (n_n5155) & (n_n5121) & (!n_n5151) & (!n_n5134)) + ((!n_n5123) & (n_n5155) & (n_n5121) & (!n_n5151) & (n_n5134)) + ((!n_n5123) & (n_n5155) & (n_n5121) & (n_n5151) & (!n_n5134)) + ((!n_n5123) & (n_n5155) & (n_n5121) & (n_n5151) & (n_n5134)) + ((n_n5123) & (!n_n5155) & (!n_n5121) & (!n_n5151) & (!n_n5134)) + ((n_n5123) & (!n_n5155) & (!n_n5121) & (!n_n5151) & (n_n5134)) + ((n_n5123) & (!n_n5155) & (!n_n5121) & (n_n5151) & (!n_n5134)) + ((n_n5123) & (!n_n5155) & (!n_n5121) & (n_n5151) & (n_n5134)) + ((n_n5123) & (!n_n5155) & (n_n5121) & (!n_n5151) & (!n_n5134)) + ((n_n5123) & (!n_n5155) & (n_n5121) & (!n_n5151) & (n_n5134)) + ((n_n5123) & (!n_n5155) & (n_n5121) & (n_n5151) & (!n_n5134)) + ((n_n5123) & (!n_n5155) & (n_n5121) & (n_n5151) & (n_n5134)) + ((n_n5123) & (n_n5155) & (!n_n5121) & (!n_n5151) & (!n_n5134)) + ((n_n5123) & (n_n5155) & (!n_n5121) & (!n_n5151) & (n_n5134)) + ((n_n5123) & (n_n5155) & (!n_n5121) & (n_n5151) & (!n_n5134)) + ((n_n5123) & (n_n5155) & (!n_n5121) & (n_n5151) & (n_n5134)) + ((n_n5123) & (n_n5155) & (n_n5121) & (!n_n5151) & (!n_n5134)) + ((n_n5123) & (n_n5155) & (n_n5121) & (!n_n5151) & (n_n5134)) + ((n_n5123) & (n_n5155) & (n_n5121) & (n_n5151) & (!n_n5134)) + ((n_n5123) & (n_n5155) & (n_n5121) & (n_n5151) & (n_n5134)));
	assign x22211x = (((!n_n4416) & (!n_n4415) & (!n_n4409) & (!n_n4417)));
	assign n_n4097 = (((!n_n4414) & (!n_n4411) & (!n_n4412) & (!x79x) & (!x22211x)) + ((!n_n4414) & (!n_n4411) & (!n_n4412) & (x79x) & (!x22211x)) + ((!n_n4414) & (!n_n4411) & (!n_n4412) & (x79x) & (x22211x)) + ((!n_n4414) & (!n_n4411) & (n_n4412) & (!x79x) & (!x22211x)) + ((!n_n4414) & (!n_n4411) & (n_n4412) & (!x79x) & (x22211x)) + ((!n_n4414) & (!n_n4411) & (n_n4412) & (x79x) & (!x22211x)) + ((!n_n4414) & (!n_n4411) & (n_n4412) & (x79x) & (x22211x)) + ((!n_n4414) & (n_n4411) & (!n_n4412) & (!x79x) & (!x22211x)) + ((!n_n4414) & (n_n4411) & (!n_n4412) & (!x79x) & (x22211x)) + ((!n_n4414) & (n_n4411) & (!n_n4412) & (x79x) & (!x22211x)) + ((!n_n4414) & (n_n4411) & (!n_n4412) & (x79x) & (x22211x)) + ((!n_n4414) & (n_n4411) & (n_n4412) & (!x79x) & (!x22211x)) + ((!n_n4414) & (n_n4411) & (n_n4412) & (!x79x) & (x22211x)) + ((!n_n4414) & (n_n4411) & (n_n4412) & (x79x) & (!x22211x)) + ((!n_n4414) & (n_n4411) & (n_n4412) & (x79x) & (x22211x)) + ((n_n4414) & (!n_n4411) & (!n_n4412) & (!x79x) & (!x22211x)) + ((n_n4414) & (!n_n4411) & (!n_n4412) & (!x79x) & (x22211x)) + ((n_n4414) & (!n_n4411) & (!n_n4412) & (x79x) & (!x22211x)) + ((n_n4414) & (!n_n4411) & (!n_n4412) & (x79x) & (x22211x)) + ((n_n4414) & (!n_n4411) & (n_n4412) & (!x79x) & (!x22211x)) + ((n_n4414) & (!n_n4411) & (n_n4412) & (!x79x) & (x22211x)) + ((n_n4414) & (!n_n4411) & (n_n4412) & (x79x) & (!x22211x)) + ((n_n4414) & (!n_n4411) & (n_n4412) & (x79x) & (x22211x)) + ((n_n4414) & (n_n4411) & (!n_n4412) & (!x79x) & (!x22211x)) + ((n_n4414) & (n_n4411) & (!n_n4412) & (!x79x) & (x22211x)) + ((n_n4414) & (n_n4411) & (!n_n4412) & (x79x) & (!x22211x)) + ((n_n4414) & (n_n4411) & (!n_n4412) & (x79x) & (x22211x)) + ((n_n4414) & (n_n4411) & (n_n4412) & (!x79x) & (!x22211x)) + ((n_n4414) & (n_n4411) & (n_n4412) & (!x79x) & (x22211x)) + ((n_n4414) & (n_n4411) & (n_n4412) & (x79x) & (!x22211x)) + ((n_n4414) & (n_n4411) & (n_n4412) & (x79x) & (x22211x)));
	assign x398x = (((!i_9_) & (n_n536) & (!n_n526) & (n_n528) & (n_n509)) + ((!i_9_) & (n_n536) & (n_n526) & (n_n528) & (n_n509)) + ((i_9_) & (n_n536) & (n_n526) & (!n_n528) & (n_n509)) + ((i_9_) & (n_n536) & (n_n526) & (n_n528) & (n_n509)));
	assign n_n4694 = (((i_9_) & (n_n390) & (n_n520) & (n_n464)));
	assign n_n4219 = (((!i_9_) & (!n_n526) & (n_n528) & (n_n325) & (n_n535)) + ((!i_9_) & (n_n526) & (n_n528) & (n_n325) & (n_n535)) + ((i_9_) & (!n_n526) & (n_n528) & (n_n325) & (n_n535)) + ((i_9_) & (n_n526) & (!n_n528) & (n_n325) & (n_n535)) + ((i_9_) & (n_n526) & (n_n528) & (n_n325) & (n_n535)));
	assign x30x = (((!i_9_) & (n_n325) & (n_n535) & (!n_n520) & (x20x)) + ((!i_9_) & (n_n325) & (n_n535) & (n_n520) & (x20x)) + ((i_9_) & (n_n325) & (n_n535) & (!n_n520) & (x20x)) + ((i_9_) & (n_n325) & (n_n535) & (n_n520) & (!x20x)) + ((i_9_) & (n_n325) & (n_n535) & (n_n520) & (x20x)));
	assign n_n4721 = (((!i_9_) & (n_n518) & (n_n526) & (n_n325)));
	assign x13293x = (((!n_n473) & (!n_n532) & (!n_n534) & (!x12x) & (n_n4129)) + ((!n_n473) & (!n_n532) & (!n_n534) & (x12x) & (n_n4129)) + ((!n_n473) & (!n_n532) & (n_n534) & (!x12x) & (n_n4129)) + ((!n_n473) & (!n_n532) & (n_n534) & (x12x) & (n_n4129)) + ((!n_n473) & (n_n532) & (!n_n534) & (!x12x) & (n_n4129)) + ((!n_n473) & (n_n532) & (!n_n534) & (x12x) & (n_n4129)) + ((!n_n473) & (n_n532) & (n_n534) & (!x12x) & (n_n4129)) + ((!n_n473) & (n_n532) & (n_n534) & (x12x) & (n_n4129)) + ((n_n473) & (!n_n532) & (!n_n534) & (!x12x) & (n_n4129)) + ((n_n473) & (!n_n532) & (!n_n534) & (x12x) & (n_n4129)) + ((n_n473) & (!n_n532) & (n_n534) & (!x12x) & (n_n4129)) + ((n_n473) & (!n_n532) & (n_n534) & (x12x) & (!n_n4129)) + ((n_n473) & (!n_n532) & (n_n534) & (x12x) & (n_n4129)) + ((n_n473) & (n_n532) & (!n_n534) & (!x12x) & (n_n4129)) + ((n_n473) & (n_n532) & (!n_n534) & (x12x) & (!n_n4129)) + ((n_n473) & (n_n532) & (!n_n534) & (x12x) & (n_n4129)) + ((n_n473) & (n_n532) & (n_n534) & (!x12x) & (n_n4129)) + ((n_n473) & (n_n532) & (n_n534) & (x12x) & (!n_n4129)) + ((n_n473) & (n_n532) & (n_n534) & (x12x) & (n_n4129)));
	assign x13296x = (((!n_n5167) & (!n_n5173) & (!n_n5166) & (n_n5172)) + ((!n_n5167) & (!n_n5173) & (n_n5166) & (!n_n5172)) + ((!n_n5167) & (!n_n5173) & (n_n5166) & (n_n5172)) + ((!n_n5167) & (n_n5173) & (!n_n5166) & (!n_n5172)) + ((!n_n5167) & (n_n5173) & (!n_n5166) & (n_n5172)) + ((!n_n5167) & (n_n5173) & (n_n5166) & (!n_n5172)) + ((!n_n5167) & (n_n5173) & (n_n5166) & (n_n5172)) + ((n_n5167) & (!n_n5173) & (!n_n5166) & (!n_n5172)) + ((n_n5167) & (!n_n5173) & (!n_n5166) & (n_n5172)) + ((n_n5167) & (!n_n5173) & (n_n5166) & (!n_n5172)) + ((n_n5167) & (!n_n5173) & (n_n5166) & (n_n5172)) + ((n_n5167) & (n_n5173) & (!n_n5166) & (!n_n5172)) + ((n_n5167) & (n_n5173) & (!n_n5166) & (n_n5172)) + ((n_n5167) & (n_n5173) & (n_n5166) & (!n_n5172)) + ((n_n5167) & (n_n5173) & (n_n5166) & (n_n5172)));
	assign x303x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n260) & (n_n535)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n260) & (n_n535)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n260) & (n_n535)) + ((i_9_) & (n_n524) & (n_n526) & (n_n260) & (n_n535)));
	assign x422x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n130) & (n_n500)) + ((!i_9_) & (n_n524) & (!n_n526) & (n_n130) & (n_n500)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n130) & (n_n500)));
	assign x13580x = (((!n_n5117) & (!n_n5119) & (!n_n5144) & (x422x)) + ((!n_n5117) & (!n_n5119) & (n_n5144) & (!x422x)) + ((!n_n5117) & (!n_n5119) & (n_n5144) & (x422x)) + ((!n_n5117) & (n_n5119) & (!n_n5144) & (!x422x)) + ((!n_n5117) & (n_n5119) & (!n_n5144) & (x422x)) + ((!n_n5117) & (n_n5119) & (n_n5144) & (!x422x)) + ((!n_n5117) & (n_n5119) & (n_n5144) & (x422x)) + ((n_n5117) & (!n_n5119) & (!n_n5144) & (!x422x)) + ((n_n5117) & (!n_n5119) & (!n_n5144) & (x422x)) + ((n_n5117) & (!n_n5119) & (n_n5144) & (!x422x)) + ((n_n5117) & (!n_n5119) & (n_n5144) & (x422x)) + ((n_n5117) & (n_n5119) & (!n_n5144) & (!x422x)) + ((n_n5117) & (n_n5119) & (!n_n5144) & (x422x)) + ((n_n5117) & (n_n5119) & (n_n5144) & (!x422x)) + ((n_n5117) & (n_n5119) & (n_n5144) & (x422x)));
	assign n_n3926 = (((!n_n5112) & (!n_n5123) & (!n_n5136) & (!n_n5104) & (x13580x)) + ((!n_n5112) & (!n_n5123) & (!n_n5136) & (n_n5104) & (!x13580x)) + ((!n_n5112) & (!n_n5123) & (!n_n5136) & (n_n5104) & (x13580x)) + ((!n_n5112) & (!n_n5123) & (n_n5136) & (!n_n5104) & (!x13580x)) + ((!n_n5112) & (!n_n5123) & (n_n5136) & (!n_n5104) & (x13580x)) + ((!n_n5112) & (!n_n5123) & (n_n5136) & (n_n5104) & (!x13580x)) + ((!n_n5112) & (!n_n5123) & (n_n5136) & (n_n5104) & (x13580x)) + ((!n_n5112) & (n_n5123) & (!n_n5136) & (!n_n5104) & (!x13580x)) + ((!n_n5112) & (n_n5123) & (!n_n5136) & (!n_n5104) & (x13580x)) + ((!n_n5112) & (n_n5123) & (!n_n5136) & (n_n5104) & (!x13580x)) + ((!n_n5112) & (n_n5123) & (!n_n5136) & (n_n5104) & (x13580x)) + ((!n_n5112) & (n_n5123) & (n_n5136) & (!n_n5104) & (!x13580x)) + ((!n_n5112) & (n_n5123) & (n_n5136) & (!n_n5104) & (x13580x)) + ((!n_n5112) & (n_n5123) & (n_n5136) & (n_n5104) & (!x13580x)) + ((!n_n5112) & (n_n5123) & (n_n5136) & (n_n5104) & (x13580x)) + ((n_n5112) & (!n_n5123) & (!n_n5136) & (!n_n5104) & (!x13580x)) + ((n_n5112) & (!n_n5123) & (!n_n5136) & (!n_n5104) & (x13580x)) + ((n_n5112) & (!n_n5123) & (!n_n5136) & (n_n5104) & (!x13580x)) + ((n_n5112) & (!n_n5123) & (!n_n5136) & (n_n5104) & (x13580x)) + ((n_n5112) & (!n_n5123) & (n_n5136) & (!n_n5104) & (!x13580x)) + ((n_n5112) & (!n_n5123) & (n_n5136) & (!n_n5104) & (x13580x)) + ((n_n5112) & (!n_n5123) & (n_n5136) & (n_n5104) & (!x13580x)) + ((n_n5112) & (!n_n5123) & (n_n5136) & (n_n5104) & (x13580x)) + ((n_n5112) & (n_n5123) & (!n_n5136) & (!n_n5104) & (!x13580x)) + ((n_n5112) & (n_n5123) & (!n_n5136) & (!n_n5104) & (x13580x)) + ((n_n5112) & (n_n5123) & (!n_n5136) & (n_n5104) & (!x13580x)) + ((n_n5112) & (n_n5123) & (!n_n5136) & (n_n5104) & (x13580x)) + ((n_n5112) & (n_n5123) & (n_n5136) & (!n_n5104) & (!x13580x)) + ((n_n5112) & (n_n5123) & (n_n5136) & (!n_n5104) & (x13580x)) + ((n_n5112) & (n_n5123) & (n_n5136) & (n_n5104) & (!x13580x)) + ((n_n5112) & (n_n5123) & (n_n5136) & (n_n5104) & (x13580x)));
	assign x13587x = (((!n_n5240) & (!n_n5222) & (!n_n5250) & (!n_n5227) & (n_n5219)) + ((!n_n5240) & (!n_n5222) & (!n_n5250) & (n_n5227) & (!n_n5219)) + ((!n_n5240) & (!n_n5222) & (!n_n5250) & (n_n5227) & (n_n5219)) + ((!n_n5240) & (!n_n5222) & (n_n5250) & (!n_n5227) & (!n_n5219)) + ((!n_n5240) & (!n_n5222) & (n_n5250) & (!n_n5227) & (n_n5219)) + ((!n_n5240) & (!n_n5222) & (n_n5250) & (n_n5227) & (!n_n5219)) + ((!n_n5240) & (!n_n5222) & (n_n5250) & (n_n5227) & (n_n5219)) + ((!n_n5240) & (n_n5222) & (!n_n5250) & (!n_n5227) & (!n_n5219)) + ((!n_n5240) & (n_n5222) & (!n_n5250) & (!n_n5227) & (n_n5219)) + ((!n_n5240) & (n_n5222) & (!n_n5250) & (n_n5227) & (!n_n5219)) + ((!n_n5240) & (n_n5222) & (!n_n5250) & (n_n5227) & (n_n5219)) + ((!n_n5240) & (n_n5222) & (n_n5250) & (!n_n5227) & (!n_n5219)) + ((!n_n5240) & (n_n5222) & (n_n5250) & (!n_n5227) & (n_n5219)) + ((!n_n5240) & (n_n5222) & (n_n5250) & (n_n5227) & (!n_n5219)) + ((!n_n5240) & (n_n5222) & (n_n5250) & (n_n5227) & (n_n5219)) + ((n_n5240) & (!n_n5222) & (!n_n5250) & (!n_n5227) & (!n_n5219)) + ((n_n5240) & (!n_n5222) & (!n_n5250) & (!n_n5227) & (n_n5219)) + ((n_n5240) & (!n_n5222) & (!n_n5250) & (n_n5227) & (!n_n5219)) + ((n_n5240) & (!n_n5222) & (!n_n5250) & (n_n5227) & (n_n5219)) + ((n_n5240) & (!n_n5222) & (n_n5250) & (!n_n5227) & (!n_n5219)) + ((n_n5240) & (!n_n5222) & (n_n5250) & (!n_n5227) & (n_n5219)) + ((n_n5240) & (!n_n5222) & (n_n5250) & (n_n5227) & (!n_n5219)) + ((n_n5240) & (!n_n5222) & (n_n5250) & (n_n5227) & (n_n5219)) + ((n_n5240) & (n_n5222) & (!n_n5250) & (!n_n5227) & (!n_n5219)) + ((n_n5240) & (n_n5222) & (!n_n5250) & (!n_n5227) & (n_n5219)) + ((n_n5240) & (n_n5222) & (!n_n5250) & (n_n5227) & (!n_n5219)) + ((n_n5240) & (n_n5222) & (!n_n5250) & (n_n5227) & (n_n5219)) + ((n_n5240) & (n_n5222) & (n_n5250) & (!n_n5227) & (!n_n5219)) + ((n_n5240) & (n_n5222) & (n_n5250) & (!n_n5227) & (n_n5219)) + ((n_n5240) & (n_n5222) & (n_n5250) & (n_n5227) & (!n_n5219)) + ((n_n5240) & (n_n5222) & (n_n5250) & (n_n5227) & (n_n5219)));
	assign n_n3924 = (((!n_n5236) & (!n_n5278) & (!n_n5260) & (!n_n5286) & (x13587x)) + ((!n_n5236) & (!n_n5278) & (!n_n5260) & (n_n5286) & (!x13587x)) + ((!n_n5236) & (!n_n5278) & (!n_n5260) & (n_n5286) & (x13587x)) + ((!n_n5236) & (!n_n5278) & (n_n5260) & (!n_n5286) & (!x13587x)) + ((!n_n5236) & (!n_n5278) & (n_n5260) & (!n_n5286) & (x13587x)) + ((!n_n5236) & (!n_n5278) & (n_n5260) & (n_n5286) & (!x13587x)) + ((!n_n5236) & (!n_n5278) & (n_n5260) & (n_n5286) & (x13587x)) + ((!n_n5236) & (n_n5278) & (!n_n5260) & (!n_n5286) & (!x13587x)) + ((!n_n5236) & (n_n5278) & (!n_n5260) & (!n_n5286) & (x13587x)) + ((!n_n5236) & (n_n5278) & (!n_n5260) & (n_n5286) & (!x13587x)) + ((!n_n5236) & (n_n5278) & (!n_n5260) & (n_n5286) & (x13587x)) + ((!n_n5236) & (n_n5278) & (n_n5260) & (!n_n5286) & (!x13587x)) + ((!n_n5236) & (n_n5278) & (n_n5260) & (!n_n5286) & (x13587x)) + ((!n_n5236) & (n_n5278) & (n_n5260) & (n_n5286) & (!x13587x)) + ((!n_n5236) & (n_n5278) & (n_n5260) & (n_n5286) & (x13587x)) + ((n_n5236) & (!n_n5278) & (!n_n5260) & (!n_n5286) & (!x13587x)) + ((n_n5236) & (!n_n5278) & (!n_n5260) & (!n_n5286) & (x13587x)) + ((n_n5236) & (!n_n5278) & (!n_n5260) & (n_n5286) & (!x13587x)) + ((n_n5236) & (!n_n5278) & (!n_n5260) & (n_n5286) & (x13587x)) + ((n_n5236) & (!n_n5278) & (n_n5260) & (!n_n5286) & (!x13587x)) + ((n_n5236) & (!n_n5278) & (n_n5260) & (!n_n5286) & (x13587x)) + ((n_n5236) & (!n_n5278) & (n_n5260) & (n_n5286) & (!x13587x)) + ((n_n5236) & (!n_n5278) & (n_n5260) & (n_n5286) & (x13587x)) + ((n_n5236) & (n_n5278) & (!n_n5260) & (!n_n5286) & (!x13587x)) + ((n_n5236) & (n_n5278) & (!n_n5260) & (!n_n5286) & (x13587x)) + ((n_n5236) & (n_n5278) & (!n_n5260) & (n_n5286) & (!x13587x)) + ((n_n5236) & (n_n5278) & (!n_n5260) & (n_n5286) & (x13587x)) + ((n_n5236) & (n_n5278) & (n_n5260) & (!n_n5286) & (!x13587x)) + ((n_n5236) & (n_n5278) & (n_n5260) & (!n_n5286) & (x13587x)) + ((n_n5236) & (n_n5278) & (n_n5260) & (n_n5286) & (!x13587x)) + ((n_n5236) & (n_n5278) & (n_n5260) & (n_n5286) & (x13587x)));
	assign x13592x = (((!n_n5293) & (!n_n5296) & (!n_n5311) & (n_n5323)) + ((!n_n5293) & (!n_n5296) & (n_n5311) & (!n_n5323)) + ((!n_n5293) & (!n_n5296) & (n_n5311) & (n_n5323)) + ((!n_n5293) & (n_n5296) & (!n_n5311) & (!n_n5323)) + ((!n_n5293) & (n_n5296) & (!n_n5311) & (n_n5323)) + ((!n_n5293) & (n_n5296) & (n_n5311) & (!n_n5323)) + ((!n_n5293) & (n_n5296) & (n_n5311) & (n_n5323)) + ((n_n5293) & (!n_n5296) & (!n_n5311) & (!n_n5323)) + ((n_n5293) & (!n_n5296) & (!n_n5311) & (n_n5323)) + ((n_n5293) & (!n_n5296) & (n_n5311) & (!n_n5323)) + ((n_n5293) & (!n_n5296) & (n_n5311) & (n_n5323)) + ((n_n5293) & (n_n5296) & (!n_n5311) & (!n_n5323)) + ((n_n5293) & (n_n5296) & (!n_n5311) & (n_n5323)) + ((n_n5293) & (n_n5296) & (n_n5311) & (!n_n5323)) + ((n_n5293) & (n_n5296) & (n_n5311) & (n_n5323)));
	assign x13593x = (((!n_n5297) & (!n_n5312) & (!n_n5289) & (!n_n5298) & (n_n5333)) + ((!n_n5297) & (!n_n5312) & (!n_n5289) & (n_n5298) & (!n_n5333)) + ((!n_n5297) & (!n_n5312) & (!n_n5289) & (n_n5298) & (n_n5333)) + ((!n_n5297) & (!n_n5312) & (n_n5289) & (!n_n5298) & (!n_n5333)) + ((!n_n5297) & (!n_n5312) & (n_n5289) & (!n_n5298) & (n_n5333)) + ((!n_n5297) & (!n_n5312) & (n_n5289) & (n_n5298) & (!n_n5333)) + ((!n_n5297) & (!n_n5312) & (n_n5289) & (n_n5298) & (n_n5333)) + ((!n_n5297) & (n_n5312) & (!n_n5289) & (!n_n5298) & (!n_n5333)) + ((!n_n5297) & (n_n5312) & (!n_n5289) & (!n_n5298) & (n_n5333)) + ((!n_n5297) & (n_n5312) & (!n_n5289) & (n_n5298) & (!n_n5333)) + ((!n_n5297) & (n_n5312) & (!n_n5289) & (n_n5298) & (n_n5333)) + ((!n_n5297) & (n_n5312) & (n_n5289) & (!n_n5298) & (!n_n5333)) + ((!n_n5297) & (n_n5312) & (n_n5289) & (!n_n5298) & (n_n5333)) + ((!n_n5297) & (n_n5312) & (n_n5289) & (n_n5298) & (!n_n5333)) + ((!n_n5297) & (n_n5312) & (n_n5289) & (n_n5298) & (n_n5333)) + ((n_n5297) & (!n_n5312) & (!n_n5289) & (!n_n5298) & (!n_n5333)) + ((n_n5297) & (!n_n5312) & (!n_n5289) & (!n_n5298) & (n_n5333)) + ((n_n5297) & (!n_n5312) & (!n_n5289) & (n_n5298) & (!n_n5333)) + ((n_n5297) & (!n_n5312) & (!n_n5289) & (n_n5298) & (n_n5333)) + ((n_n5297) & (!n_n5312) & (n_n5289) & (!n_n5298) & (!n_n5333)) + ((n_n5297) & (!n_n5312) & (n_n5289) & (!n_n5298) & (n_n5333)) + ((n_n5297) & (!n_n5312) & (n_n5289) & (n_n5298) & (!n_n5333)) + ((n_n5297) & (!n_n5312) & (n_n5289) & (n_n5298) & (n_n5333)) + ((n_n5297) & (n_n5312) & (!n_n5289) & (!n_n5298) & (!n_n5333)) + ((n_n5297) & (n_n5312) & (!n_n5289) & (!n_n5298) & (n_n5333)) + ((n_n5297) & (n_n5312) & (!n_n5289) & (n_n5298) & (!n_n5333)) + ((n_n5297) & (n_n5312) & (!n_n5289) & (n_n5298) & (n_n5333)) + ((n_n5297) & (n_n5312) & (n_n5289) & (!n_n5298) & (!n_n5333)) + ((n_n5297) & (n_n5312) & (n_n5289) & (!n_n5298) & (n_n5333)) + ((n_n5297) & (n_n5312) & (n_n5289) & (n_n5298) & (!n_n5333)) + ((n_n5297) & (n_n5312) & (n_n5289) & (n_n5298) & (n_n5333)));
	assign x13599x = (((!n_n4920) & (!n_n4987) & (!n_n4963) & (n_n4974)) + ((!n_n4920) & (!n_n4987) & (n_n4963) & (!n_n4974)) + ((!n_n4920) & (!n_n4987) & (n_n4963) & (n_n4974)) + ((!n_n4920) & (n_n4987) & (!n_n4963) & (!n_n4974)) + ((!n_n4920) & (n_n4987) & (!n_n4963) & (n_n4974)) + ((!n_n4920) & (n_n4987) & (n_n4963) & (!n_n4974)) + ((!n_n4920) & (n_n4987) & (n_n4963) & (n_n4974)) + ((n_n4920) & (!n_n4987) & (!n_n4963) & (!n_n4974)) + ((n_n4920) & (!n_n4987) & (!n_n4963) & (n_n4974)) + ((n_n4920) & (!n_n4987) & (n_n4963) & (!n_n4974)) + ((n_n4920) & (!n_n4987) & (n_n4963) & (n_n4974)) + ((n_n4920) & (n_n4987) & (!n_n4963) & (!n_n4974)) + ((n_n4920) & (n_n4987) & (!n_n4963) & (n_n4974)) + ((n_n4920) & (n_n4987) & (n_n4963) & (!n_n4974)) + ((n_n4920) & (n_n4987) & (n_n4963) & (n_n4974)));
	assign x13600x = (((!n_n4927) & (!n_n4958) & (!n_n4994) & (!n_n5009) & (n_n4961)) + ((!n_n4927) & (!n_n4958) & (!n_n4994) & (n_n5009) & (!n_n4961)) + ((!n_n4927) & (!n_n4958) & (!n_n4994) & (n_n5009) & (n_n4961)) + ((!n_n4927) & (!n_n4958) & (n_n4994) & (!n_n5009) & (!n_n4961)) + ((!n_n4927) & (!n_n4958) & (n_n4994) & (!n_n5009) & (n_n4961)) + ((!n_n4927) & (!n_n4958) & (n_n4994) & (n_n5009) & (!n_n4961)) + ((!n_n4927) & (!n_n4958) & (n_n4994) & (n_n5009) & (n_n4961)) + ((!n_n4927) & (n_n4958) & (!n_n4994) & (!n_n5009) & (!n_n4961)) + ((!n_n4927) & (n_n4958) & (!n_n4994) & (!n_n5009) & (n_n4961)) + ((!n_n4927) & (n_n4958) & (!n_n4994) & (n_n5009) & (!n_n4961)) + ((!n_n4927) & (n_n4958) & (!n_n4994) & (n_n5009) & (n_n4961)) + ((!n_n4927) & (n_n4958) & (n_n4994) & (!n_n5009) & (!n_n4961)) + ((!n_n4927) & (n_n4958) & (n_n4994) & (!n_n5009) & (n_n4961)) + ((!n_n4927) & (n_n4958) & (n_n4994) & (n_n5009) & (!n_n4961)) + ((!n_n4927) & (n_n4958) & (n_n4994) & (n_n5009) & (n_n4961)) + ((n_n4927) & (!n_n4958) & (!n_n4994) & (!n_n5009) & (!n_n4961)) + ((n_n4927) & (!n_n4958) & (!n_n4994) & (!n_n5009) & (n_n4961)) + ((n_n4927) & (!n_n4958) & (!n_n4994) & (n_n5009) & (!n_n4961)) + ((n_n4927) & (!n_n4958) & (!n_n4994) & (n_n5009) & (n_n4961)) + ((n_n4927) & (!n_n4958) & (n_n4994) & (!n_n5009) & (!n_n4961)) + ((n_n4927) & (!n_n4958) & (n_n4994) & (!n_n5009) & (n_n4961)) + ((n_n4927) & (!n_n4958) & (n_n4994) & (n_n5009) & (!n_n4961)) + ((n_n4927) & (!n_n4958) & (n_n4994) & (n_n5009) & (n_n4961)) + ((n_n4927) & (n_n4958) & (!n_n4994) & (!n_n5009) & (!n_n4961)) + ((n_n4927) & (n_n4958) & (!n_n4994) & (!n_n5009) & (n_n4961)) + ((n_n4927) & (n_n4958) & (!n_n4994) & (n_n5009) & (!n_n4961)) + ((n_n4927) & (n_n4958) & (!n_n4994) & (n_n5009) & (n_n4961)) + ((n_n4927) & (n_n4958) & (n_n4994) & (!n_n5009) & (!n_n4961)) + ((n_n4927) & (n_n4958) & (n_n4994) & (!n_n5009) & (n_n4961)) + ((n_n4927) & (n_n4958) & (n_n4994) & (n_n5009) & (!n_n4961)) + ((n_n4927) & (n_n4958) & (n_n4994) & (n_n5009) & (n_n4961)));
	assign x13950x = (((!n_n518) & (!x11x) & (!x24x) & (!n_n65) & (n_n5226)) + ((!n_n518) & (!x11x) & (!x24x) & (n_n65) & (n_n5226)) + ((!n_n518) & (!x11x) & (x24x) & (!n_n65) & (n_n5226)) + ((!n_n518) & (!x11x) & (x24x) & (n_n65) & (n_n5226)) + ((!n_n518) & (x11x) & (!x24x) & (!n_n65) & (n_n5226)) + ((!n_n518) & (x11x) & (!x24x) & (n_n65) & (n_n5226)) + ((!n_n518) & (x11x) & (x24x) & (!n_n65) & (n_n5226)) + ((!n_n518) & (x11x) & (x24x) & (n_n65) & (n_n5226)) + ((n_n518) & (!x11x) & (!x24x) & (!n_n65) & (n_n5226)) + ((n_n518) & (!x11x) & (!x24x) & (n_n65) & (n_n5226)) + ((n_n518) & (!x11x) & (x24x) & (!n_n65) & (n_n5226)) + ((n_n518) & (!x11x) & (x24x) & (n_n65) & (!n_n5226)) + ((n_n518) & (!x11x) & (x24x) & (n_n65) & (n_n5226)) + ((n_n518) & (x11x) & (!x24x) & (!n_n65) & (n_n5226)) + ((n_n518) & (x11x) & (!x24x) & (n_n65) & (!n_n5226)) + ((n_n518) & (x11x) & (!x24x) & (n_n65) & (n_n5226)) + ((n_n518) & (x11x) & (x24x) & (!n_n65) & (n_n5226)) + ((n_n518) & (x11x) & (x24x) & (n_n65) & (!n_n5226)) + ((n_n518) & (x11x) & (x24x) & (n_n65) & (n_n5226)));
	assign x14047x = (((!i_7_) & (!i_8_) & (!i_6_) & (x12x) & (n_n464)) + ((i_7_) & (i_8_) & (!i_6_) & (x12x) & (n_n464)));
	assign n_n3051 = (((!x25x) & (!n_n130) & (!n_n500) & (!n_n5127) & (n_n5126)) + ((!x25x) & (!n_n130) & (!n_n500) & (n_n5127) & (!n_n5126)) + ((!x25x) & (!n_n130) & (!n_n500) & (n_n5127) & (n_n5126)) + ((!x25x) & (!n_n130) & (n_n500) & (!n_n5127) & (n_n5126)) + ((!x25x) & (!n_n130) & (n_n500) & (n_n5127) & (!n_n5126)) + ((!x25x) & (!n_n130) & (n_n500) & (n_n5127) & (n_n5126)) + ((!x25x) & (n_n130) & (!n_n500) & (!n_n5127) & (n_n5126)) + ((!x25x) & (n_n130) & (!n_n500) & (n_n5127) & (!n_n5126)) + ((!x25x) & (n_n130) & (!n_n500) & (n_n5127) & (n_n5126)) + ((!x25x) & (n_n130) & (n_n500) & (!n_n5127) & (n_n5126)) + ((!x25x) & (n_n130) & (n_n500) & (n_n5127) & (!n_n5126)) + ((!x25x) & (n_n130) & (n_n500) & (n_n5127) & (n_n5126)) + ((x25x) & (!n_n130) & (!n_n500) & (!n_n5127) & (n_n5126)) + ((x25x) & (!n_n130) & (!n_n500) & (n_n5127) & (!n_n5126)) + ((x25x) & (!n_n130) & (!n_n500) & (n_n5127) & (n_n5126)) + ((x25x) & (!n_n130) & (n_n500) & (!n_n5127) & (n_n5126)) + ((x25x) & (!n_n130) & (n_n500) & (n_n5127) & (!n_n5126)) + ((x25x) & (!n_n130) & (n_n500) & (n_n5127) & (n_n5126)) + ((x25x) & (n_n130) & (!n_n500) & (!n_n5127) & (n_n5126)) + ((x25x) & (n_n130) & (!n_n500) & (n_n5127) & (!n_n5126)) + ((x25x) & (n_n130) & (!n_n500) & (n_n5127) & (n_n5126)) + ((x25x) & (n_n130) & (n_n500) & (!n_n5127) & (!n_n5126)) + ((x25x) & (n_n130) & (n_n500) & (!n_n5127) & (n_n5126)) + ((x25x) & (n_n130) & (n_n500) & (n_n5127) & (!n_n5126)) + ((x25x) & (n_n130) & (n_n500) & (n_n5127) & (n_n5126)));
	assign x15508x = (((!n_n4388) & (!n_n4392) & (!n_n4393) & (!n_n4396) & (n_n4399)) + ((!n_n4388) & (!n_n4392) & (!n_n4393) & (n_n4396) & (!n_n4399)) + ((!n_n4388) & (!n_n4392) & (!n_n4393) & (n_n4396) & (n_n4399)) + ((!n_n4388) & (!n_n4392) & (n_n4393) & (!n_n4396) & (!n_n4399)) + ((!n_n4388) & (!n_n4392) & (n_n4393) & (!n_n4396) & (n_n4399)) + ((!n_n4388) & (!n_n4392) & (n_n4393) & (n_n4396) & (!n_n4399)) + ((!n_n4388) & (!n_n4392) & (n_n4393) & (n_n4396) & (n_n4399)) + ((!n_n4388) & (n_n4392) & (!n_n4393) & (!n_n4396) & (!n_n4399)) + ((!n_n4388) & (n_n4392) & (!n_n4393) & (!n_n4396) & (n_n4399)) + ((!n_n4388) & (n_n4392) & (!n_n4393) & (n_n4396) & (!n_n4399)) + ((!n_n4388) & (n_n4392) & (!n_n4393) & (n_n4396) & (n_n4399)) + ((!n_n4388) & (n_n4392) & (n_n4393) & (!n_n4396) & (!n_n4399)) + ((!n_n4388) & (n_n4392) & (n_n4393) & (!n_n4396) & (n_n4399)) + ((!n_n4388) & (n_n4392) & (n_n4393) & (n_n4396) & (!n_n4399)) + ((!n_n4388) & (n_n4392) & (n_n4393) & (n_n4396) & (n_n4399)) + ((n_n4388) & (!n_n4392) & (!n_n4393) & (!n_n4396) & (!n_n4399)) + ((n_n4388) & (!n_n4392) & (!n_n4393) & (!n_n4396) & (n_n4399)) + ((n_n4388) & (!n_n4392) & (!n_n4393) & (n_n4396) & (!n_n4399)) + ((n_n4388) & (!n_n4392) & (!n_n4393) & (n_n4396) & (n_n4399)) + ((n_n4388) & (!n_n4392) & (n_n4393) & (!n_n4396) & (!n_n4399)) + ((n_n4388) & (!n_n4392) & (n_n4393) & (!n_n4396) & (n_n4399)) + ((n_n4388) & (!n_n4392) & (n_n4393) & (n_n4396) & (!n_n4399)) + ((n_n4388) & (!n_n4392) & (n_n4393) & (n_n4396) & (n_n4399)) + ((n_n4388) & (n_n4392) & (!n_n4393) & (!n_n4396) & (!n_n4399)) + ((n_n4388) & (n_n4392) & (!n_n4393) & (!n_n4396) & (n_n4399)) + ((n_n4388) & (n_n4392) & (!n_n4393) & (n_n4396) & (!n_n4399)) + ((n_n4388) & (n_n4392) & (!n_n4393) & (n_n4396) & (n_n4399)) + ((n_n4388) & (n_n4392) & (n_n4393) & (!n_n4396) & (!n_n4399)) + ((n_n4388) & (n_n4392) & (n_n4393) & (!n_n4396) & (n_n4399)) + ((n_n4388) & (n_n4392) & (n_n4393) & (n_n4396) & (!n_n4399)) + ((n_n4388) & (n_n4392) & (n_n4393) & (n_n4396) & (n_n4399)));
	assign x440x = (((!n_n473) & (!n_n325) & (!x23x) & (n_n4808)) + ((!n_n473) & (!n_n325) & (x23x) & (n_n4808)) + ((!n_n473) & (n_n325) & (!x23x) & (n_n4808)) + ((!n_n473) & (n_n325) & (x23x) & (n_n4808)) + ((n_n473) & (!n_n325) & (!x23x) & (n_n4808)) + ((n_n473) & (!n_n325) & (x23x) & (n_n4808)) + ((n_n473) & (n_n325) & (!x23x) & (n_n4808)) + ((n_n473) & (n_n325) & (x23x) & (!n_n4808)) + ((n_n473) & (n_n325) & (x23x) & (n_n4808)));
	assign x12460x = (((!n_n4403) & (!n_n4415) & (!n_n4405) & (!n_n4406) & (n_n4408)) + ((!n_n4403) & (!n_n4415) & (!n_n4405) & (n_n4406) & (!n_n4408)) + ((!n_n4403) & (!n_n4415) & (!n_n4405) & (n_n4406) & (n_n4408)) + ((!n_n4403) & (!n_n4415) & (n_n4405) & (!n_n4406) & (!n_n4408)) + ((!n_n4403) & (!n_n4415) & (n_n4405) & (!n_n4406) & (n_n4408)) + ((!n_n4403) & (!n_n4415) & (n_n4405) & (n_n4406) & (!n_n4408)) + ((!n_n4403) & (!n_n4415) & (n_n4405) & (n_n4406) & (n_n4408)) + ((!n_n4403) & (n_n4415) & (!n_n4405) & (!n_n4406) & (!n_n4408)) + ((!n_n4403) & (n_n4415) & (!n_n4405) & (!n_n4406) & (n_n4408)) + ((!n_n4403) & (n_n4415) & (!n_n4405) & (n_n4406) & (!n_n4408)) + ((!n_n4403) & (n_n4415) & (!n_n4405) & (n_n4406) & (n_n4408)) + ((!n_n4403) & (n_n4415) & (n_n4405) & (!n_n4406) & (!n_n4408)) + ((!n_n4403) & (n_n4415) & (n_n4405) & (!n_n4406) & (n_n4408)) + ((!n_n4403) & (n_n4415) & (n_n4405) & (n_n4406) & (!n_n4408)) + ((!n_n4403) & (n_n4415) & (n_n4405) & (n_n4406) & (n_n4408)) + ((n_n4403) & (!n_n4415) & (!n_n4405) & (!n_n4406) & (!n_n4408)) + ((n_n4403) & (!n_n4415) & (!n_n4405) & (!n_n4406) & (n_n4408)) + ((n_n4403) & (!n_n4415) & (!n_n4405) & (n_n4406) & (!n_n4408)) + ((n_n4403) & (!n_n4415) & (!n_n4405) & (n_n4406) & (n_n4408)) + ((n_n4403) & (!n_n4415) & (n_n4405) & (!n_n4406) & (!n_n4408)) + ((n_n4403) & (!n_n4415) & (n_n4405) & (!n_n4406) & (n_n4408)) + ((n_n4403) & (!n_n4415) & (n_n4405) & (n_n4406) & (!n_n4408)) + ((n_n4403) & (!n_n4415) & (n_n4405) & (n_n4406) & (n_n4408)) + ((n_n4403) & (n_n4415) & (!n_n4405) & (!n_n4406) & (!n_n4408)) + ((n_n4403) & (n_n4415) & (!n_n4405) & (!n_n4406) & (n_n4408)) + ((n_n4403) & (n_n4415) & (!n_n4405) & (n_n4406) & (!n_n4408)) + ((n_n4403) & (n_n4415) & (!n_n4405) & (n_n4406) & (n_n4408)) + ((n_n4403) & (n_n4415) & (n_n4405) & (!n_n4406) & (!n_n4408)) + ((n_n4403) & (n_n4415) & (n_n4405) & (!n_n4406) & (n_n4408)) + ((n_n4403) & (n_n4415) & (n_n4405) & (n_n4406) & (!n_n4408)) + ((n_n4403) & (n_n4415) & (n_n4405) & (n_n4406) & (n_n4408)));
	assign x360x = (((!i_9_) & (n_n536) & (n_n482) & (n_n532) & (!n_n530)) + ((!i_9_) & (n_n536) & (n_n482) & (n_n532) & (n_n530)) + ((i_9_) & (n_n536) & (n_n482) & (!n_n532) & (n_n530)) + ((i_9_) & (n_n536) & (n_n482) & (n_n532) & (n_n530)));
	assign x22142x = (((!n_n4431) & (!n_n4433) & (!n_n4392) & (!n_n4398) & (!n_n4429)));
	assign x12469x = (((!n_n4399) & (!n_n4421) & (!n_n4428) & (!x215x) & (!x22142x)) + ((!n_n4399) & (!n_n4421) & (!n_n4428) & (x215x) & (!x22142x)) + ((!n_n4399) & (!n_n4421) & (!n_n4428) & (x215x) & (x22142x)) + ((!n_n4399) & (!n_n4421) & (n_n4428) & (!x215x) & (!x22142x)) + ((!n_n4399) & (!n_n4421) & (n_n4428) & (!x215x) & (x22142x)) + ((!n_n4399) & (!n_n4421) & (n_n4428) & (x215x) & (!x22142x)) + ((!n_n4399) & (!n_n4421) & (n_n4428) & (x215x) & (x22142x)) + ((!n_n4399) & (n_n4421) & (!n_n4428) & (!x215x) & (!x22142x)) + ((!n_n4399) & (n_n4421) & (!n_n4428) & (!x215x) & (x22142x)) + ((!n_n4399) & (n_n4421) & (!n_n4428) & (x215x) & (!x22142x)) + ((!n_n4399) & (n_n4421) & (!n_n4428) & (x215x) & (x22142x)) + ((!n_n4399) & (n_n4421) & (n_n4428) & (!x215x) & (!x22142x)) + ((!n_n4399) & (n_n4421) & (n_n4428) & (!x215x) & (x22142x)) + ((!n_n4399) & (n_n4421) & (n_n4428) & (x215x) & (!x22142x)) + ((!n_n4399) & (n_n4421) & (n_n4428) & (x215x) & (x22142x)) + ((n_n4399) & (!n_n4421) & (!n_n4428) & (!x215x) & (!x22142x)) + ((n_n4399) & (!n_n4421) & (!n_n4428) & (!x215x) & (x22142x)) + ((n_n4399) & (!n_n4421) & (!n_n4428) & (x215x) & (!x22142x)) + ((n_n4399) & (!n_n4421) & (!n_n4428) & (x215x) & (x22142x)) + ((n_n4399) & (!n_n4421) & (n_n4428) & (!x215x) & (!x22142x)) + ((n_n4399) & (!n_n4421) & (n_n4428) & (!x215x) & (x22142x)) + ((n_n4399) & (!n_n4421) & (n_n4428) & (x215x) & (!x22142x)) + ((n_n4399) & (!n_n4421) & (n_n4428) & (x215x) & (x22142x)) + ((n_n4399) & (n_n4421) & (!n_n4428) & (!x215x) & (!x22142x)) + ((n_n4399) & (n_n4421) & (!n_n4428) & (!x215x) & (x22142x)) + ((n_n4399) & (n_n4421) & (!n_n4428) & (x215x) & (!x22142x)) + ((n_n4399) & (n_n4421) & (!n_n4428) & (x215x) & (x22142x)) + ((n_n4399) & (n_n4421) & (n_n4428) & (!x215x) & (!x22142x)) + ((n_n4399) & (n_n4421) & (n_n4428) & (!x215x) & (x22142x)) + ((n_n4399) & (n_n4421) & (n_n4428) & (x215x) & (!x22142x)) + ((n_n4399) & (n_n4421) & (n_n4428) & (x215x) & (x22142x)));
	assign x12468x = (((!n_n4401) & (!x216x) & (!x37x) & (!n_n4402) & (x360x)) + ((!n_n4401) & (!x216x) & (!x37x) & (n_n4402) & (!x360x)) + ((!n_n4401) & (!x216x) & (!x37x) & (n_n4402) & (x360x)) + ((!n_n4401) & (!x216x) & (x37x) & (!n_n4402) & (!x360x)) + ((!n_n4401) & (!x216x) & (x37x) & (!n_n4402) & (x360x)) + ((!n_n4401) & (!x216x) & (x37x) & (n_n4402) & (!x360x)) + ((!n_n4401) & (!x216x) & (x37x) & (n_n4402) & (x360x)) + ((!n_n4401) & (x216x) & (!x37x) & (!n_n4402) & (!x360x)) + ((!n_n4401) & (x216x) & (!x37x) & (!n_n4402) & (x360x)) + ((!n_n4401) & (x216x) & (!x37x) & (n_n4402) & (!x360x)) + ((!n_n4401) & (x216x) & (!x37x) & (n_n4402) & (x360x)) + ((!n_n4401) & (x216x) & (x37x) & (!n_n4402) & (!x360x)) + ((!n_n4401) & (x216x) & (x37x) & (!n_n4402) & (x360x)) + ((!n_n4401) & (x216x) & (x37x) & (n_n4402) & (!x360x)) + ((!n_n4401) & (x216x) & (x37x) & (n_n4402) & (x360x)) + ((n_n4401) & (!x216x) & (!x37x) & (!n_n4402) & (!x360x)) + ((n_n4401) & (!x216x) & (!x37x) & (!n_n4402) & (x360x)) + ((n_n4401) & (!x216x) & (!x37x) & (n_n4402) & (!x360x)) + ((n_n4401) & (!x216x) & (!x37x) & (n_n4402) & (x360x)) + ((n_n4401) & (!x216x) & (x37x) & (!n_n4402) & (!x360x)) + ((n_n4401) & (!x216x) & (x37x) & (!n_n4402) & (x360x)) + ((n_n4401) & (!x216x) & (x37x) & (n_n4402) & (!x360x)) + ((n_n4401) & (!x216x) & (x37x) & (n_n4402) & (x360x)) + ((n_n4401) & (x216x) & (!x37x) & (!n_n4402) & (!x360x)) + ((n_n4401) & (x216x) & (!x37x) & (!n_n4402) & (x360x)) + ((n_n4401) & (x216x) & (!x37x) & (n_n4402) & (!x360x)) + ((n_n4401) & (x216x) & (!x37x) & (n_n4402) & (x360x)) + ((n_n4401) & (x216x) & (x37x) & (!n_n4402) & (!x360x)) + ((n_n4401) & (x216x) & (x37x) & (!n_n4402) & (x360x)) + ((n_n4401) & (x216x) & (x37x) & (n_n4402) & (!x360x)) + ((n_n4401) & (x216x) & (x37x) & (n_n4402) & (x360x)));
	assign x22143x = (((!x21x) & (!x483x) & (!n_n4738) & (!n_n4744) & (!n_n4745)) + ((!x21x) & (x483x) & (!n_n4738) & (!n_n4744) & (!n_n4745)) + ((x21x) & (!x483x) & (!n_n4738) & (!n_n4744) & (!n_n4745)));
	assign x12357x = (((!x19x) & (!n_n528) & (!n_n500) & (!n_n530) & (x77x)) + ((!x19x) & (!n_n528) & (!n_n500) & (n_n530) & (x77x)) + ((!x19x) & (!n_n528) & (n_n500) & (!n_n530) & (x77x)) + ((!x19x) & (!n_n528) & (n_n500) & (n_n530) & (x77x)) + ((!x19x) & (n_n528) & (!n_n500) & (!n_n530) & (x77x)) + ((!x19x) & (n_n528) & (!n_n500) & (n_n530) & (x77x)) + ((!x19x) & (n_n528) & (n_n500) & (!n_n530) & (x77x)) + ((!x19x) & (n_n528) & (n_n500) & (n_n530) & (x77x)) + ((x19x) & (!n_n528) & (!n_n500) & (!n_n530) & (x77x)) + ((x19x) & (!n_n528) & (!n_n500) & (n_n530) & (x77x)) + ((x19x) & (!n_n528) & (n_n500) & (!n_n530) & (x77x)) + ((x19x) & (!n_n528) & (n_n500) & (n_n530) & (!x77x)) + ((x19x) & (!n_n528) & (n_n500) & (n_n530) & (x77x)) + ((x19x) & (n_n528) & (!n_n500) & (!n_n530) & (x77x)) + ((x19x) & (n_n528) & (!n_n500) & (n_n530) & (x77x)) + ((x19x) & (n_n528) & (n_n500) & (!n_n530) & (!x77x)) + ((x19x) & (n_n528) & (n_n500) & (!n_n530) & (x77x)) + ((x19x) & (n_n528) & (n_n500) & (n_n530) & (!x77x)) + ((x19x) & (n_n528) & (n_n500) & (n_n530) & (x77x)));
	assign x12358x = (((!x19x) & (!n_n526) & (!n_n500) & (!n_n5265) & (n_n1521)) + ((!x19x) & (!n_n526) & (!n_n500) & (n_n5265) & (!n_n1521)) + ((!x19x) & (!n_n526) & (!n_n500) & (n_n5265) & (n_n1521)) + ((!x19x) & (!n_n526) & (n_n500) & (!n_n5265) & (n_n1521)) + ((!x19x) & (!n_n526) & (n_n500) & (n_n5265) & (!n_n1521)) + ((!x19x) & (!n_n526) & (n_n500) & (n_n5265) & (n_n1521)) + ((!x19x) & (n_n526) & (!n_n500) & (!n_n5265) & (n_n1521)) + ((!x19x) & (n_n526) & (!n_n500) & (n_n5265) & (!n_n1521)) + ((!x19x) & (n_n526) & (!n_n500) & (n_n5265) & (n_n1521)) + ((!x19x) & (n_n526) & (n_n500) & (!n_n5265) & (n_n1521)) + ((!x19x) & (n_n526) & (n_n500) & (n_n5265) & (!n_n1521)) + ((!x19x) & (n_n526) & (n_n500) & (n_n5265) & (n_n1521)) + ((x19x) & (!n_n526) & (!n_n500) & (!n_n5265) & (n_n1521)) + ((x19x) & (!n_n526) & (!n_n500) & (n_n5265) & (!n_n1521)) + ((x19x) & (!n_n526) & (!n_n500) & (n_n5265) & (n_n1521)) + ((x19x) & (!n_n526) & (n_n500) & (!n_n5265) & (n_n1521)) + ((x19x) & (!n_n526) & (n_n500) & (n_n5265) & (!n_n1521)) + ((x19x) & (!n_n526) & (n_n500) & (n_n5265) & (n_n1521)) + ((x19x) & (n_n526) & (!n_n500) & (!n_n5265) & (n_n1521)) + ((x19x) & (n_n526) & (!n_n500) & (n_n5265) & (!n_n1521)) + ((x19x) & (n_n526) & (!n_n500) & (n_n5265) & (n_n1521)) + ((x19x) & (n_n526) & (n_n500) & (!n_n5265) & (!n_n1521)) + ((x19x) & (n_n526) & (n_n500) & (!n_n5265) & (n_n1521)) + ((x19x) & (n_n526) & (n_n500) & (n_n5265) & (!n_n1521)) + ((x19x) & (n_n526) & (n_n500) & (n_n5265) & (n_n1521)));
	assign n_n1404 = (((!n_n1435) & (!n_n1436) & (!x12357x) & (x12358x)) + ((!n_n1435) & (!n_n1436) & (x12357x) & (!x12358x)) + ((!n_n1435) & (!n_n1436) & (x12357x) & (x12358x)) + ((!n_n1435) & (n_n1436) & (!x12357x) & (!x12358x)) + ((!n_n1435) & (n_n1436) & (!x12357x) & (x12358x)) + ((!n_n1435) & (n_n1436) & (x12357x) & (!x12358x)) + ((!n_n1435) & (n_n1436) & (x12357x) & (x12358x)) + ((n_n1435) & (!n_n1436) & (!x12357x) & (!x12358x)) + ((n_n1435) & (!n_n1436) & (!x12357x) & (x12358x)) + ((n_n1435) & (!n_n1436) & (x12357x) & (!x12358x)) + ((n_n1435) & (!n_n1436) & (x12357x) & (x12358x)) + ((n_n1435) & (n_n1436) & (!x12357x) & (!x12358x)) + ((n_n1435) & (n_n1436) & (!x12357x) & (x12358x)) + ((n_n1435) & (n_n1436) & (x12357x) & (!x12358x)) + ((n_n1435) & (n_n1436) & (x12357x) & (x12358x)));
	assign x12321x = (((!x15x) & (!x11x) & (!n_n195) & (!n_n464) & (n_n5073)) + ((!x15x) & (!x11x) & (!n_n195) & (n_n464) & (n_n5073)) + ((!x15x) & (!x11x) & (n_n195) & (!n_n464) & (n_n5073)) + ((!x15x) & (!x11x) & (n_n195) & (n_n464) & (n_n5073)) + ((!x15x) & (x11x) & (!n_n195) & (!n_n464) & (n_n5073)) + ((!x15x) & (x11x) & (!n_n195) & (n_n464) & (n_n5073)) + ((!x15x) & (x11x) & (n_n195) & (!n_n464) & (n_n5073)) + ((!x15x) & (x11x) & (n_n195) & (n_n464) & (!n_n5073)) + ((!x15x) & (x11x) & (n_n195) & (n_n464) & (n_n5073)) + ((x15x) & (!x11x) & (!n_n195) & (!n_n464) & (n_n5073)) + ((x15x) & (!x11x) & (!n_n195) & (n_n464) & (n_n5073)) + ((x15x) & (!x11x) & (n_n195) & (!n_n464) & (n_n5073)) + ((x15x) & (!x11x) & (n_n195) & (n_n464) & (!n_n5073)) + ((x15x) & (!x11x) & (n_n195) & (n_n464) & (n_n5073)) + ((x15x) & (x11x) & (!n_n195) & (!n_n464) & (n_n5073)) + ((x15x) & (x11x) & (!n_n195) & (n_n464) & (n_n5073)) + ((x15x) & (x11x) & (n_n195) & (!n_n464) & (n_n5073)) + ((x15x) & (x11x) & (n_n195) & (n_n464) & (!n_n5073)) + ((x15x) & (x11x) & (n_n195) & (n_n464) & (n_n5073)));
	assign x12322x = (((!i_7_) & (!i_8_) & (i_6_) & (x18x) & (n_n464)) + ((!i_7_) & (i_8_) & (!i_6_) & (x18x) & (n_n464)) + ((i_7_) & (!i_8_) & (!i_6_) & (x18x) & (n_n464)) + ((i_7_) & (i_8_) & (!i_6_) & (x18x) & (n_n464)));
	assign x12333x = (((!n_n5085) & (!n_n5082) & (!n_n5084) & (n_n5079)) + ((!n_n5085) & (!n_n5082) & (n_n5084) & (!n_n5079)) + ((!n_n5085) & (!n_n5082) & (n_n5084) & (n_n5079)) + ((!n_n5085) & (n_n5082) & (!n_n5084) & (!n_n5079)) + ((!n_n5085) & (n_n5082) & (!n_n5084) & (n_n5079)) + ((!n_n5085) & (n_n5082) & (n_n5084) & (!n_n5079)) + ((!n_n5085) & (n_n5082) & (n_n5084) & (n_n5079)) + ((n_n5085) & (!n_n5082) & (!n_n5084) & (!n_n5079)) + ((n_n5085) & (!n_n5082) & (!n_n5084) & (n_n5079)) + ((n_n5085) & (!n_n5082) & (n_n5084) & (!n_n5079)) + ((n_n5085) & (!n_n5082) & (n_n5084) & (n_n5079)) + ((n_n5085) & (n_n5082) & (!n_n5084) & (!n_n5079)) + ((n_n5085) & (n_n5082) & (!n_n5084) & (n_n5079)) + ((n_n5085) & (n_n5082) & (n_n5084) & (!n_n5079)) + ((n_n5085) & (n_n5082) & (n_n5084) & (n_n5079)));
	assign x12334x = (((!n_n5087) & (!n_n5088) & (!n_n5078) & (!n_n5083) & (n_n5077)) + ((!n_n5087) & (!n_n5088) & (!n_n5078) & (n_n5083) & (!n_n5077)) + ((!n_n5087) & (!n_n5088) & (!n_n5078) & (n_n5083) & (n_n5077)) + ((!n_n5087) & (!n_n5088) & (n_n5078) & (!n_n5083) & (!n_n5077)) + ((!n_n5087) & (!n_n5088) & (n_n5078) & (!n_n5083) & (n_n5077)) + ((!n_n5087) & (!n_n5088) & (n_n5078) & (n_n5083) & (!n_n5077)) + ((!n_n5087) & (!n_n5088) & (n_n5078) & (n_n5083) & (n_n5077)) + ((!n_n5087) & (n_n5088) & (!n_n5078) & (!n_n5083) & (!n_n5077)) + ((!n_n5087) & (n_n5088) & (!n_n5078) & (!n_n5083) & (n_n5077)) + ((!n_n5087) & (n_n5088) & (!n_n5078) & (n_n5083) & (!n_n5077)) + ((!n_n5087) & (n_n5088) & (!n_n5078) & (n_n5083) & (n_n5077)) + ((!n_n5087) & (n_n5088) & (n_n5078) & (!n_n5083) & (!n_n5077)) + ((!n_n5087) & (n_n5088) & (n_n5078) & (!n_n5083) & (n_n5077)) + ((!n_n5087) & (n_n5088) & (n_n5078) & (n_n5083) & (!n_n5077)) + ((!n_n5087) & (n_n5088) & (n_n5078) & (n_n5083) & (n_n5077)) + ((n_n5087) & (!n_n5088) & (!n_n5078) & (!n_n5083) & (!n_n5077)) + ((n_n5087) & (!n_n5088) & (!n_n5078) & (!n_n5083) & (n_n5077)) + ((n_n5087) & (!n_n5088) & (!n_n5078) & (n_n5083) & (!n_n5077)) + ((n_n5087) & (!n_n5088) & (!n_n5078) & (n_n5083) & (n_n5077)) + ((n_n5087) & (!n_n5088) & (n_n5078) & (!n_n5083) & (!n_n5077)) + ((n_n5087) & (!n_n5088) & (n_n5078) & (!n_n5083) & (n_n5077)) + ((n_n5087) & (!n_n5088) & (n_n5078) & (n_n5083) & (!n_n5077)) + ((n_n5087) & (!n_n5088) & (n_n5078) & (n_n5083) & (n_n5077)) + ((n_n5087) & (n_n5088) & (!n_n5078) & (!n_n5083) & (!n_n5077)) + ((n_n5087) & (n_n5088) & (!n_n5078) & (!n_n5083) & (n_n5077)) + ((n_n5087) & (n_n5088) & (!n_n5078) & (n_n5083) & (!n_n5077)) + ((n_n5087) & (n_n5088) & (!n_n5078) & (n_n5083) & (n_n5077)) + ((n_n5087) & (n_n5088) & (n_n5078) & (!n_n5083) & (!n_n5077)) + ((n_n5087) & (n_n5088) & (n_n5078) & (!n_n5083) & (n_n5077)) + ((n_n5087) & (n_n5088) & (n_n5078) & (n_n5083) & (!n_n5077)) + ((n_n5087) & (n_n5088) & (n_n5078) & (n_n5083) & (n_n5077)));
	assign x12338x = (((!n_n5093) & (!n_n5091) & (!n_n5101) & (n_n5105)) + ((!n_n5093) & (!n_n5091) & (n_n5101) & (!n_n5105)) + ((!n_n5093) & (!n_n5091) & (n_n5101) & (n_n5105)) + ((!n_n5093) & (n_n5091) & (!n_n5101) & (!n_n5105)) + ((!n_n5093) & (n_n5091) & (!n_n5101) & (n_n5105)) + ((!n_n5093) & (n_n5091) & (n_n5101) & (!n_n5105)) + ((!n_n5093) & (n_n5091) & (n_n5101) & (n_n5105)) + ((n_n5093) & (!n_n5091) & (!n_n5101) & (!n_n5105)) + ((n_n5093) & (!n_n5091) & (!n_n5101) & (n_n5105)) + ((n_n5093) & (!n_n5091) & (n_n5101) & (!n_n5105)) + ((n_n5093) & (!n_n5091) & (n_n5101) & (n_n5105)) + ((n_n5093) & (n_n5091) & (!n_n5101) & (!n_n5105)) + ((n_n5093) & (n_n5091) & (!n_n5101) & (n_n5105)) + ((n_n5093) & (n_n5091) & (n_n5101) & (!n_n5105)) + ((n_n5093) & (n_n5091) & (n_n5101) & (n_n5105)));
	assign x12339x = (((!n_n5100) & (!n_n5098) & (!n_n5103) & (!n_n5095) & (x88x)) + ((!n_n5100) & (!n_n5098) & (!n_n5103) & (n_n5095) & (!x88x)) + ((!n_n5100) & (!n_n5098) & (!n_n5103) & (n_n5095) & (x88x)) + ((!n_n5100) & (!n_n5098) & (n_n5103) & (!n_n5095) & (!x88x)) + ((!n_n5100) & (!n_n5098) & (n_n5103) & (!n_n5095) & (x88x)) + ((!n_n5100) & (!n_n5098) & (n_n5103) & (n_n5095) & (!x88x)) + ((!n_n5100) & (!n_n5098) & (n_n5103) & (n_n5095) & (x88x)) + ((!n_n5100) & (n_n5098) & (!n_n5103) & (!n_n5095) & (!x88x)) + ((!n_n5100) & (n_n5098) & (!n_n5103) & (!n_n5095) & (x88x)) + ((!n_n5100) & (n_n5098) & (!n_n5103) & (n_n5095) & (!x88x)) + ((!n_n5100) & (n_n5098) & (!n_n5103) & (n_n5095) & (x88x)) + ((!n_n5100) & (n_n5098) & (n_n5103) & (!n_n5095) & (!x88x)) + ((!n_n5100) & (n_n5098) & (n_n5103) & (!n_n5095) & (x88x)) + ((!n_n5100) & (n_n5098) & (n_n5103) & (n_n5095) & (!x88x)) + ((!n_n5100) & (n_n5098) & (n_n5103) & (n_n5095) & (x88x)) + ((n_n5100) & (!n_n5098) & (!n_n5103) & (!n_n5095) & (!x88x)) + ((n_n5100) & (!n_n5098) & (!n_n5103) & (!n_n5095) & (x88x)) + ((n_n5100) & (!n_n5098) & (!n_n5103) & (n_n5095) & (!x88x)) + ((n_n5100) & (!n_n5098) & (!n_n5103) & (n_n5095) & (x88x)) + ((n_n5100) & (!n_n5098) & (n_n5103) & (!n_n5095) & (!x88x)) + ((n_n5100) & (!n_n5098) & (n_n5103) & (!n_n5095) & (x88x)) + ((n_n5100) & (!n_n5098) & (n_n5103) & (n_n5095) & (!x88x)) + ((n_n5100) & (!n_n5098) & (n_n5103) & (n_n5095) & (x88x)) + ((n_n5100) & (n_n5098) & (!n_n5103) & (!n_n5095) & (!x88x)) + ((n_n5100) & (n_n5098) & (!n_n5103) & (!n_n5095) & (x88x)) + ((n_n5100) & (n_n5098) & (!n_n5103) & (n_n5095) & (!x88x)) + ((n_n5100) & (n_n5098) & (!n_n5103) & (n_n5095) & (x88x)) + ((n_n5100) & (n_n5098) & (n_n5103) & (!n_n5095) & (!x88x)) + ((n_n5100) & (n_n5098) & (n_n5103) & (!n_n5095) & (x88x)) + ((n_n5100) & (n_n5098) & (n_n5103) & (n_n5095) & (!x88x)) + ((n_n5100) & (n_n5098) & (n_n5103) & (n_n5095) & (x88x)));
	assign x347x = (((!i_9_) & (n_n455) & (!n_n528) & (n_n500) & (n_n530)) + ((!i_9_) & (n_n455) & (n_n528) & (n_n500) & (!n_n530)) + ((!i_9_) & (n_n455) & (n_n528) & (n_n500) & (n_n530)));
	assign x12952x = (((!x21x) & (!n_n491) & (!n_n65) & (!n_n3382) & (n_n5280)) + ((!x21x) & (!n_n491) & (!n_n65) & (n_n3382) & (!n_n5280)) + ((!x21x) & (!n_n491) & (!n_n65) & (n_n3382) & (n_n5280)) + ((!x21x) & (!n_n491) & (n_n65) & (!n_n3382) & (n_n5280)) + ((!x21x) & (!n_n491) & (n_n65) & (n_n3382) & (!n_n5280)) + ((!x21x) & (!n_n491) & (n_n65) & (n_n3382) & (n_n5280)) + ((!x21x) & (n_n491) & (!n_n65) & (!n_n3382) & (n_n5280)) + ((!x21x) & (n_n491) & (!n_n65) & (n_n3382) & (!n_n5280)) + ((!x21x) & (n_n491) & (!n_n65) & (n_n3382) & (n_n5280)) + ((!x21x) & (n_n491) & (n_n65) & (!n_n3382) & (n_n5280)) + ((!x21x) & (n_n491) & (n_n65) & (n_n3382) & (!n_n5280)) + ((!x21x) & (n_n491) & (n_n65) & (n_n3382) & (n_n5280)) + ((x21x) & (!n_n491) & (!n_n65) & (!n_n3382) & (n_n5280)) + ((x21x) & (!n_n491) & (!n_n65) & (n_n3382) & (!n_n5280)) + ((x21x) & (!n_n491) & (!n_n65) & (n_n3382) & (n_n5280)) + ((x21x) & (!n_n491) & (n_n65) & (!n_n3382) & (n_n5280)) + ((x21x) & (!n_n491) & (n_n65) & (n_n3382) & (!n_n5280)) + ((x21x) & (!n_n491) & (n_n65) & (n_n3382) & (n_n5280)) + ((x21x) & (n_n491) & (!n_n65) & (!n_n3382) & (n_n5280)) + ((x21x) & (n_n491) & (!n_n65) & (n_n3382) & (!n_n5280)) + ((x21x) & (n_n491) & (!n_n65) & (n_n3382) & (n_n5280)) + ((x21x) & (n_n491) & (n_n65) & (!n_n3382) & (!n_n5280)) + ((x21x) & (n_n491) & (n_n65) & (!n_n3382) & (n_n5280)) + ((x21x) & (n_n491) & (n_n65) & (n_n3382) & (!n_n5280)) + ((x21x) & (n_n491) & (n_n65) & (n_n3382) & (n_n5280)));
	assign n_n664 = (((!n_n5274) & (!n_n5273) & (!n_n5275) & (!n_n5285) & (x12952x)) + ((!n_n5274) & (!n_n5273) & (!n_n5275) & (n_n5285) & (!x12952x)) + ((!n_n5274) & (!n_n5273) & (!n_n5275) & (n_n5285) & (x12952x)) + ((!n_n5274) & (!n_n5273) & (n_n5275) & (!n_n5285) & (!x12952x)) + ((!n_n5274) & (!n_n5273) & (n_n5275) & (!n_n5285) & (x12952x)) + ((!n_n5274) & (!n_n5273) & (n_n5275) & (n_n5285) & (!x12952x)) + ((!n_n5274) & (!n_n5273) & (n_n5275) & (n_n5285) & (x12952x)) + ((!n_n5274) & (n_n5273) & (!n_n5275) & (!n_n5285) & (!x12952x)) + ((!n_n5274) & (n_n5273) & (!n_n5275) & (!n_n5285) & (x12952x)) + ((!n_n5274) & (n_n5273) & (!n_n5275) & (n_n5285) & (!x12952x)) + ((!n_n5274) & (n_n5273) & (!n_n5275) & (n_n5285) & (x12952x)) + ((!n_n5274) & (n_n5273) & (n_n5275) & (!n_n5285) & (!x12952x)) + ((!n_n5274) & (n_n5273) & (n_n5275) & (!n_n5285) & (x12952x)) + ((!n_n5274) & (n_n5273) & (n_n5275) & (n_n5285) & (!x12952x)) + ((!n_n5274) & (n_n5273) & (n_n5275) & (n_n5285) & (x12952x)) + ((n_n5274) & (!n_n5273) & (!n_n5275) & (!n_n5285) & (!x12952x)) + ((n_n5274) & (!n_n5273) & (!n_n5275) & (!n_n5285) & (x12952x)) + ((n_n5274) & (!n_n5273) & (!n_n5275) & (n_n5285) & (!x12952x)) + ((n_n5274) & (!n_n5273) & (!n_n5275) & (n_n5285) & (x12952x)) + ((n_n5274) & (!n_n5273) & (n_n5275) & (!n_n5285) & (!x12952x)) + ((n_n5274) & (!n_n5273) & (n_n5275) & (!n_n5285) & (x12952x)) + ((n_n5274) & (!n_n5273) & (n_n5275) & (n_n5285) & (!x12952x)) + ((n_n5274) & (!n_n5273) & (n_n5275) & (n_n5285) & (x12952x)) + ((n_n5274) & (n_n5273) & (!n_n5275) & (!n_n5285) & (!x12952x)) + ((n_n5274) & (n_n5273) & (!n_n5275) & (!n_n5285) & (x12952x)) + ((n_n5274) & (n_n5273) & (!n_n5275) & (n_n5285) & (!x12952x)) + ((n_n5274) & (n_n5273) & (!n_n5275) & (n_n5285) & (x12952x)) + ((n_n5274) & (n_n5273) & (n_n5275) & (!n_n5285) & (!x12952x)) + ((n_n5274) & (n_n5273) & (n_n5275) & (!n_n5285) & (x12952x)) + ((n_n5274) & (n_n5273) & (n_n5275) & (n_n5285) & (!x12952x)) + ((n_n5274) & (n_n5273) & (n_n5275) & (n_n5285) & (x12952x)));
	assign x12958x = (((!n_n5254) & (!n_n5252) & (!n_n5260) & (n_n5253)) + ((!n_n5254) & (!n_n5252) & (n_n5260) & (!n_n5253)) + ((!n_n5254) & (!n_n5252) & (n_n5260) & (n_n5253)) + ((!n_n5254) & (n_n5252) & (!n_n5260) & (!n_n5253)) + ((!n_n5254) & (n_n5252) & (!n_n5260) & (n_n5253)) + ((!n_n5254) & (n_n5252) & (n_n5260) & (!n_n5253)) + ((!n_n5254) & (n_n5252) & (n_n5260) & (n_n5253)) + ((n_n5254) & (!n_n5252) & (!n_n5260) & (!n_n5253)) + ((n_n5254) & (!n_n5252) & (!n_n5260) & (n_n5253)) + ((n_n5254) & (!n_n5252) & (n_n5260) & (!n_n5253)) + ((n_n5254) & (!n_n5252) & (n_n5260) & (n_n5253)) + ((n_n5254) & (n_n5252) & (!n_n5260) & (!n_n5253)) + ((n_n5254) & (n_n5252) & (!n_n5260) & (n_n5253)) + ((n_n5254) & (n_n5252) & (n_n5260) & (!n_n5253)) + ((n_n5254) & (n_n5252) & (n_n5260) & (n_n5253)));
	assign x12960x = (((!n_n5267) & (!n_n5251) & (!x77x) & (!x446x) & (x205x)) + ((!n_n5267) & (!n_n5251) & (!x77x) & (x446x) & (!x205x)) + ((!n_n5267) & (!n_n5251) & (!x77x) & (x446x) & (x205x)) + ((!n_n5267) & (!n_n5251) & (x77x) & (!x446x) & (!x205x)) + ((!n_n5267) & (!n_n5251) & (x77x) & (!x446x) & (x205x)) + ((!n_n5267) & (!n_n5251) & (x77x) & (x446x) & (!x205x)) + ((!n_n5267) & (!n_n5251) & (x77x) & (x446x) & (x205x)) + ((!n_n5267) & (n_n5251) & (!x77x) & (!x446x) & (!x205x)) + ((!n_n5267) & (n_n5251) & (!x77x) & (!x446x) & (x205x)) + ((!n_n5267) & (n_n5251) & (!x77x) & (x446x) & (!x205x)) + ((!n_n5267) & (n_n5251) & (!x77x) & (x446x) & (x205x)) + ((!n_n5267) & (n_n5251) & (x77x) & (!x446x) & (!x205x)) + ((!n_n5267) & (n_n5251) & (x77x) & (!x446x) & (x205x)) + ((!n_n5267) & (n_n5251) & (x77x) & (x446x) & (!x205x)) + ((!n_n5267) & (n_n5251) & (x77x) & (x446x) & (x205x)) + ((n_n5267) & (!n_n5251) & (!x77x) & (!x446x) & (!x205x)) + ((n_n5267) & (!n_n5251) & (!x77x) & (!x446x) & (x205x)) + ((n_n5267) & (!n_n5251) & (!x77x) & (x446x) & (!x205x)) + ((n_n5267) & (!n_n5251) & (!x77x) & (x446x) & (x205x)) + ((n_n5267) & (!n_n5251) & (x77x) & (!x446x) & (!x205x)) + ((n_n5267) & (!n_n5251) & (x77x) & (!x446x) & (x205x)) + ((n_n5267) & (!n_n5251) & (x77x) & (x446x) & (!x205x)) + ((n_n5267) & (!n_n5251) & (x77x) & (x446x) & (x205x)) + ((n_n5267) & (n_n5251) & (!x77x) & (!x446x) & (!x205x)) + ((n_n5267) & (n_n5251) & (!x77x) & (!x446x) & (x205x)) + ((n_n5267) & (n_n5251) & (!x77x) & (x446x) & (!x205x)) + ((n_n5267) & (n_n5251) & (!x77x) & (x446x) & (x205x)) + ((n_n5267) & (n_n5251) & (x77x) & (!x446x) & (!x205x)) + ((n_n5267) & (n_n5251) & (x77x) & (!x446x) & (x205x)) + ((n_n5267) & (n_n5251) & (x77x) & (x446x) & (!x205x)) + ((n_n5267) & (n_n5251) & (x77x) & (x446x) & (x205x)));
	assign n_n634 = (((!n_n1521) & (!n_n3385) & (!n_n664) & (!x12958x) & (x12960x)) + ((!n_n1521) & (!n_n3385) & (!n_n664) & (x12958x) & (!x12960x)) + ((!n_n1521) & (!n_n3385) & (!n_n664) & (x12958x) & (x12960x)) + ((!n_n1521) & (!n_n3385) & (n_n664) & (!x12958x) & (!x12960x)) + ((!n_n1521) & (!n_n3385) & (n_n664) & (!x12958x) & (x12960x)) + ((!n_n1521) & (!n_n3385) & (n_n664) & (x12958x) & (!x12960x)) + ((!n_n1521) & (!n_n3385) & (n_n664) & (x12958x) & (x12960x)) + ((!n_n1521) & (n_n3385) & (!n_n664) & (!x12958x) & (!x12960x)) + ((!n_n1521) & (n_n3385) & (!n_n664) & (!x12958x) & (x12960x)) + ((!n_n1521) & (n_n3385) & (!n_n664) & (x12958x) & (!x12960x)) + ((!n_n1521) & (n_n3385) & (!n_n664) & (x12958x) & (x12960x)) + ((!n_n1521) & (n_n3385) & (n_n664) & (!x12958x) & (!x12960x)) + ((!n_n1521) & (n_n3385) & (n_n664) & (!x12958x) & (x12960x)) + ((!n_n1521) & (n_n3385) & (n_n664) & (x12958x) & (!x12960x)) + ((!n_n1521) & (n_n3385) & (n_n664) & (x12958x) & (x12960x)) + ((n_n1521) & (!n_n3385) & (!n_n664) & (!x12958x) & (!x12960x)) + ((n_n1521) & (!n_n3385) & (!n_n664) & (!x12958x) & (x12960x)) + ((n_n1521) & (!n_n3385) & (!n_n664) & (x12958x) & (!x12960x)) + ((n_n1521) & (!n_n3385) & (!n_n664) & (x12958x) & (x12960x)) + ((n_n1521) & (!n_n3385) & (n_n664) & (!x12958x) & (!x12960x)) + ((n_n1521) & (!n_n3385) & (n_n664) & (!x12958x) & (x12960x)) + ((n_n1521) & (!n_n3385) & (n_n664) & (x12958x) & (!x12960x)) + ((n_n1521) & (!n_n3385) & (n_n664) & (x12958x) & (x12960x)) + ((n_n1521) & (n_n3385) & (!n_n664) & (!x12958x) & (!x12960x)) + ((n_n1521) & (n_n3385) & (!n_n664) & (!x12958x) & (x12960x)) + ((n_n1521) & (n_n3385) & (!n_n664) & (x12958x) & (!x12960x)) + ((n_n1521) & (n_n3385) & (!n_n664) & (x12958x) & (x12960x)) + ((n_n1521) & (n_n3385) & (n_n664) & (!x12958x) & (!x12960x)) + ((n_n1521) & (n_n3385) & (n_n664) & (!x12958x) & (x12960x)) + ((n_n1521) & (n_n3385) & (n_n664) & (x12958x) & (!x12960x)) + ((n_n1521) & (n_n3385) & (n_n664) & (x12958x) & (x12960x)));
	assign x12902x = (((!x21x) & (!n_n473) & (!n_n195) & (!n_n5073) & (x160x)) + ((!x21x) & (!n_n473) & (!n_n195) & (n_n5073) & (!x160x)) + ((!x21x) & (!n_n473) & (!n_n195) & (n_n5073) & (x160x)) + ((!x21x) & (!n_n473) & (n_n195) & (!n_n5073) & (x160x)) + ((!x21x) & (!n_n473) & (n_n195) & (n_n5073) & (!x160x)) + ((!x21x) & (!n_n473) & (n_n195) & (n_n5073) & (x160x)) + ((!x21x) & (n_n473) & (!n_n195) & (!n_n5073) & (x160x)) + ((!x21x) & (n_n473) & (!n_n195) & (n_n5073) & (!x160x)) + ((!x21x) & (n_n473) & (!n_n195) & (n_n5073) & (x160x)) + ((!x21x) & (n_n473) & (n_n195) & (!n_n5073) & (x160x)) + ((!x21x) & (n_n473) & (n_n195) & (n_n5073) & (!x160x)) + ((!x21x) & (n_n473) & (n_n195) & (n_n5073) & (x160x)) + ((x21x) & (!n_n473) & (!n_n195) & (!n_n5073) & (x160x)) + ((x21x) & (!n_n473) & (!n_n195) & (n_n5073) & (!x160x)) + ((x21x) & (!n_n473) & (!n_n195) & (n_n5073) & (x160x)) + ((x21x) & (!n_n473) & (n_n195) & (!n_n5073) & (x160x)) + ((x21x) & (!n_n473) & (n_n195) & (n_n5073) & (!x160x)) + ((x21x) & (!n_n473) & (n_n195) & (n_n5073) & (x160x)) + ((x21x) & (n_n473) & (!n_n195) & (!n_n5073) & (x160x)) + ((x21x) & (n_n473) & (!n_n195) & (n_n5073) & (!x160x)) + ((x21x) & (n_n473) & (!n_n195) & (n_n5073) & (x160x)) + ((x21x) & (n_n473) & (n_n195) & (!n_n5073) & (!x160x)) + ((x21x) & (n_n473) & (n_n195) & (!n_n5073) & (x160x)) + ((x21x) & (n_n473) & (n_n195) & (n_n5073) & (!x160x)) + ((x21x) & (n_n473) & (n_n195) & (n_n5073) & (x160x)));
	assign x12903x = (((!n_n524) & (!n_n473) & (!x18x) & (!n_n5061) & (n_n789)) + ((!n_n524) & (!n_n473) & (!x18x) & (n_n5061) & (!n_n789)) + ((!n_n524) & (!n_n473) & (!x18x) & (n_n5061) & (n_n789)) + ((!n_n524) & (!n_n473) & (x18x) & (!n_n5061) & (n_n789)) + ((!n_n524) & (!n_n473) & (x18x) & (n_n5061) & (!n_n789)) + ((!n_n524) & (!n_n473) & (x18x) & (n_n5061) & (n_n789)) + ((!n_n524) & (n_n473) & (!x18x) & (!n_n5061) & (n_n789)) + ((!n_n524) & (n_n473) & (!x18x) & (n_n5061) & (!n_n789)) + ((!n_n524) & (n_n473) & (!x18x) & (n_n5061) & (n_n789)) + ((!n_n524) & (n_n473) & (x18x) & (!n_n5061) & (n_n789)) + ((!n_n524) & (n_n473) & (x18x) & (n_n5061) & (!n_n789)) + ((!n_n524) & (n_n473) & (x18x) & (n_n5061) & (n_n789)) + ((n_n524) & (!n_n473) & (!x18x) & (!n_n5061) & (n_n789)) + ((n_n524) & (!n_n473) & (!x18x) & (n_n5061) & (!n_n789)) + ((n_n524) & (!n_n473) & (!x18x) & (n_n5061) & (n_n789)) + ((n_n524) & (!n_n473) & (x18x) & (!n_n5061) & (n_n789)) + ((n_n524) & (!n_n473) & (x18x) & (n_n5061) & (!n_n789)) + ((n_n524) & (!n_n473) & (x18x) & (n_n5061) & (n_n789)) + ((n_n524) & (n_n473) & (!x18x) & (!n_n5061) & (n_n789)) + ((n_n524) & (n_n473) & (!x18x) & (n_n5061) & (!n_n789)) + ((n_n524) & (n_n473) & (!x18x) & (n_n5061) & (n_n789)) + ((n_n524) & (n_n473) & (x18x) & (!n_n5061) & (!n_n789)) + ((n_n524) & (n_n473) & (x18x) & (!n_n5061) & (n_n789)) + ((n_n524) & (n_n473) & (x18x) & (n_n5061) & (!n_n789)) + ((n_n524) & (n_n473) & (x18x) & (n_n5061) & (n_n789)));
	assign x22130x = (((!n_n5055) & (!n_n5054) & (!n_n5057) & (!n_n5047)));
	assign n_n681 = (((!n_n5050) & (!n_n5049) & (!x166x) & (!n_n5051) & (!x22130x)) + ((!n_n5050) & (!n_n5049) & (!x166x) & (n_n5051) & (!x22130x)) + ((!n_n5050) & (!n_n5049) & (!x166x) & (n_n5051) & (x22130x)) + ((!n_n5050) & (!n_n5049) & (x166x) & (!n_n5051) & (!x22130x)) + ((!n_n5050) & (!n_n5049) & (x166x) & (!n_n5051) & (x22130x)) + ((!n_n5050) & (!n_n5049) & (x166x) & (n_n5051) & (!x22130x)) + ((!n_n5050) & (!n_n5049) & (x166x) & (n_n5051) & (x22130x)) + ((!n_n5050) & (n_n5049) & (!x166x) & (!n_n5051) & (!x22130x)) + ((!n_n5050) & (n_n5049) & (!x166x) & (!n_n5051) & (x22130x)) + ((!n_n5050) & (n_n5049) & (!x166x) & (n_n5051) & (!x22130x)) + ((!n_n5050) & (n_n5049) & (!x166x) & (n_n5051) & (x22130x)) + ((!n_n5050) & (n_n5049) & (x166x) & (!n_n5051) & (!x22130x)) + ((!n_n5050) & (n_n5049) & (x166x) & (!n_n5051) & (x22130x)) + ((!n_n5050) & (n_n5049) & (x166x) & (n_n5051) & (!x22130x)) + ((!n_n5050) & (n_n5049) & (x166x) & (n_n5051) & (x22130x)) + ((n_n5050) & (!n_n5049) & (!x166x) & (!n_n5051) & (!x22130x)) + ((n_n5050) & (!n_n5049) & (!x166x) & (!n_n5051) & (x22130x)) + ((n_n5050) & (!n_n5049) & (!x166x) & (n_n5051) & (!x22130x)) + ((n_n5050) & (!n_n5049) & (!x166x) & (n_n5051) & (x22130x)) + ((n_n5050) & (!n_n5049) & (x166x) & (!n_n5051) & (!x22130x)) + ((n_n5050) & (!n_n5049) & (x166x) & (!n_n5051) & (x22130x)) + ((n_n5050) & (!n_n5049) & (x166x) & (n_n5051) & (!x22130x)) + ((n_n5050) & (!n_n5049) & (x166x) & (n_n5051) & (x22130x)) + ((n_n5050) & (n_n5049) & (!x166x) & (!n_n5051) & (!x22130x)) + ((n_n5050) & (n_n5049) & (!x166x) & (!n_n5051) & (x22130x)) + ((n_n5050) & (n_n5049) & (!x166x) & (n_n5051) & (!x22130x)) + ((n_n5050) & (n_n5049) & (!x166x) & (n_n5051) & (x22130x)) + ((n_n5050) & (n_n5049) & (x166x) & (!n_n5051) & (!x22130x)) + ((n_n5050) & (n_n5049) & (x166x) & (!n_n5051) & (x22130x)) + ((n_n5050) & (n_n5049) & (x166x) & (n_n5051) & (!x22130x)) + ((n_n5050) & (n_n5049) & (x166x) & (n_n5051) & (x22130x)));
	assign x209x = (((!i_9_) & (!n_n522) & (n_n195) & (x20x) & (n_n464)) + ((!i_9_) & (n_n522) & (n_n195) & (x20x) & (n_n464)) + ((i_9_) & (!n_n522) & (n_n195) & (x20x) & (n_n464)) + ((i_9_) & (n_n522) & (n_n195) & (!x20x) & (n_n464)) + ((i_9_) & (n_n522) & (n_n195) & (x20x) & (n_n464)));
	assign x12913x = (((!x18x) & (!x516x) & (!n_n5085) & (!n_n5081) & (n_n5082)) + ((!x18x) & (!x516x) & (!n_n5085) & (n_n5081) & (!n_n5082)) + ((!x18x) & (!x516x) & (!n_n5085) & (n_n5081) & (n_n5082)) + ((!x18x) & (!x516x) & (n_n5085) & (!n_n5081) & (!n_n5082)) + ((!x18x) & (!x516x) & (n_n5085) & (!n_n5081) & (n_n5082)) + ((!x18x) & (!x516x) & (n_n5085) & (n_n5081) & (!n_n5082)) + ((!x18x) & (!x516x) & (n_n5085) & (n_n5081) & (n_n5082)) + ((!x18x) & (x516x) & (!n_n5085) & (!n_n5081) & (n_n5082)) + ((!x18x) & (x516x) & (!n_n5085) & (n_n5081) & (!n_n5082)) + ((!x18x) & (x516x) & (!n_n5085) & (n_n5081) & (n_n5082)) + ((!x18x) & (x516x) & (n_n5085) & (!n_n5081) & (!n_n5082)) + ((!x18x) & (x516x) & (n_n5085) & (!n_n5081) & (n_n5082)) + ((!x18x) & (x516x) & (n_n5085) & (n_n5081) & (!n_n5082)) + ((!x18x) & (x516x) & (n_n5085) & (n_n5081) & (n_n5082)) + ((x18x) & (!x516x) & (!n_n5085) & (!n_n5081) & (n_n5082)) + ((x18x) & (!x516x) & (!n_n5085) & (n_n5081) & (!n_n5082)) + ((x18x) & (!x516x) & (!n_n5085) & (n_n5081) & (n_n5082)) + ((x18x) & (!x516x) & (n_n5085) & (!n_n5081) & (!n_n5082)) + ((x18x) & (!x516x) & (n_n5085) & (!n_n5081) & (n_n5082)) + ((x18x) & (!x516x) & (n_n5085) & (n_n5081) & (!n_n5082)) + ((x18x) & (!x516x) & (n_n5085) & (n_n5081) & (n_n5082)) + ((x18x) & (x516x) & (!n_n5085) & (!n_n5081) & (!n_n5082)) + ((x18x) & (x516x) & (!n_n5085) & (!n_n5081) & (n_n5082)) + ((x18x) & (x516x) & (!n_n5085) & (n_n5081) & (!n_n5082)) + ((x18x) & (x516x) & (!n_n5085) & (n_n5081) & (n_n5082)) + ((x18x) & (x516x) & (n_n5085) & (!n_n5081) & (!n_n5082)) + ((x18x) & (x516x) & (n_n5085) & (!n_n5081) & (n_n5082)) + ((x18x) & (x516x) & (n_n5085) & (n_n5081) & (!n_n5082)) + ((x18x) & (x516x) & (n_n5085) & (n_n5081) & (n_n5082)));
	assign x12914x = (((!n_n5076) & (!n_n5079) & (!n_n5083) & (!n_n5077) & (n_n5080)) + ((!n_n5076) & (!n_n5079) & (!n_n5083) & (n_n5077) & (!n_n5080)) + ((!n_n5076) & (!n_n5079) & (!n_n5083) & (n_n5077) & (n_n5080)) + ((!n_n5076) & (!n_n5079) & (n_n5083) & (!n_n5077) & (!n_n5080)) + ((!n_n5076) & (!n_n5079) & (n_n5083) & (!n_n5077) & (n_n5080)) + ((!n_n5076) & (!n_n5079) & (n_n5083) & (n_n5077) & (!n_n5080)) + ((!n_n5076) & (!n_n5079) & (n_n5083) & (n_n5077) & (n_n5080)) + ((!n_n5076) & (n_n5079) & (!n_n5083) & (!n_n5077) & (!n_n5080)) + ((!n_n5076) & (n_n5079) & (!n_n5083) & (!n_n5077) & (n_n5080)) + ((!n_n5076) & (n_n5079) & (!n_n5083) & (n_n5077) & (!n_n5080)) + ((!n_n5076) & (n_n5079) & (!n_n5083) & (n_n5077) & (n_n5080)) + ((!n_n5076) & (n_n5079) & (n_n5083) & (!n_n5077) & (!n_n5080)) + ((!n_n5076) & (n_n5079) & (n_n5083) & (!n_n5077) & (n_n5080)) + ((!n_n5076) & (n_n5079) & (n_n5083) & (n_n5077) & (!n_n5080)) + ((!n_n5076) & (n_n5079) & (n_n5083) & (n_n5077) & (n_n5080)) + ((n_n5076) & (!n_n5079) & (!n_n5083) & (!n_n5077) & (!n_n5080)) + ((n_n5076) & (!n_n5079) & (!n_n5083) & (!n_n5077) & (n_n5080)) + ((n_n5076) & (!n_n5079) & (!n_n5083) & (n_n5077) & (!n_n5080)) + ((n_n5076) & (!n_n5079) & (!n_n5083) & (n_n5077) & (n_n5080)) + ((n_n5076) & (!n_n5079) & (n_n5083) & (!n_n5077) & (!n_n5080)) + ((n_n5076) & (!n_n5079) & (n_n5083) & (!n_n5077) & (n_n5080)) + ((n_n5076) & (!n_n5079) & (n_n5083) & (n_n5077) & (!n_n5080)) + ((n_n5076) & (!n_n5079) & (n_n5083) & (n_n5077) & (n_n5080)) + ((n_n5076) & (n_n5079) & (!n_n5083) & (!n_n5077) & (!n_n5080)) + ((n_n5076) & (n_n5079) & (!n_n5083) & (!n_n5077) & (n_n5080)) + ((n_n5076) & (n_n5079) & (!n_n5083) & (n_n5077) & (!n_n5080)) + ((n_n5076) & (n_n5079) & (!n_n5083) & (n_n5077) & (n_n5080)) + ((n_n5076) & (n_n5079) & (n_n5083) & (!n_n5077) & (!n_n5080)) + ((n_n5076) & (n_n5079) & (n_n5083) & (!n_n5077) & (n_n5080)) + ((n_n5076) & (n_n5079) & (n_n5083) & (n_n5077) & (!n_n5080)) + ((n_n5076) & (n_n5079) & (n_n5083) & (n_n5077) & (n_n5080)));
	assign n_n639 = (((!x12902x) & (!x12903x) & (!n_n681) & (!x12913x) & (x12914x)) + ((!x12902x) & (!x12903x) & (!n_n681) & (x12913x) & (!x12914x)) + ((!x12902x) & (!x12903x) & (!n_n681) & (x12913x) & (x12914x)) + ((!x12902x) & (!x12903x) & (n_n681) & (!x12913x) & (!x12914x)) + ((!x12902x) & (!x12903x) & (n_n681) & (!x12913x) & (x12914x)) + ((!x12902x) & (!x12903x) & (n_n681) & (x12913x) & (!x12914x)) + ((!x12902x) & (!x12903x) & (n_n681) & (x12913x) & (x12914x)) + ((!x12902x) & (x12903x) & (!n_n681) & (!x12913x) & (!x12914x)) + ((!x12902x) & (x12903x) & (!n_n681) & (!x12913x) & (x12914x)) + ((!x12902x) & (x12903x) & (!n_n681) & (x12913x) & (!x12914x)) + ((!x12902x) & (x12903x) & (!n_n681) & (x12913x) & (x12914x)) + ((!x12902x) & (x12903x) & (n_n681) & (!x12913x) & (!x12914x)) + ((!x12902x) & (x12903x) & (n_n681) & (!x12913x) & (x12914x)) + ((!x12902x) & (x12903x) & (n_n681) & (x12913x) & (!x12914x)) + ((!x12902x) & (x12903x) & (n_n681) & (x12913x) & (x12914x)) + ((x12902x) & (!x12903x) & (!n_n681) & (!x12913x) & (!x12914x)) + ((x12902x) & (!x12903x) & (!n_n681) & (!x12913x) & (x12914x)) + ((x12902x) & (!x12903x) & (!n_n681) & (x12913x) & (!x12914x)) + ((x12902x) & (!x12903x) & (!n_n681) & (x12913x) & (x12914x)) + ((x12902x) & (!x12903x) & (n_n681) & (!x12913x) & (!x12914x)) + ((x12902x) & (!x12903x) & (n_n681) & (!x12913x) & (x12914x)) + ((x12902x) & (!x12903x) & (n_n681) & (x12913x) & (!x12914x)) + ((x12902x) & (!x12903x) & (n_n681) & (x12913x) & (x12914x)) + ((x12902x) & (x12903x) & (!n_n681) & (!x12913x) & (!x12914x)) + ((x12902x) & (x12903x) & (!n_n681) & (!x12913x) & (x12914x)) + ((x12902x) & (x12903x) & (!n_n681) & (x12913x) & (!x12914x)) + ((x12902x) & (x12903x) & (!n_n681) & (x12913x) & (x12914x)) + ((x12902x) & (x12903x) & (n_n681) & (!x12913x) & (!x12914x)) + ((x12902x) & (x12903x) & (n_n681) & (!x12913x) & (x12914x)) + ((x12902x) & (x12903x) & (n_n681) & (x12913x) & (!x12914x)) + ((x12902x) & (x12903x) & (n_n681) & (x12913x) & (x12914x)));
	assign x12921x = (((!n_n5129) & (!n_n5124) & (!n_n5120) & (n_n5126)) + ((!n_n5129) & (!n_n5124) & (n_n5120) & (!n_n5126)) + ((!n_n5129) & (!n_n5124) & (n_n5120) & (n_n5126)) + ((!n_n5129) & (n_n5124) & (!n_n5120) & (!n_n5126)) + ((!n_n5129) & (n_n5124) & (!n_n5120) & (n_n5126)) + ((!n_n5129) & (n_n5124) & (n_n5120) & (!n_n5126)) + ((!n_n5129) & (n_n5124) & (n_n5120) & (n_n5126)) + ((n_n5129) & (!n_n5124) & (!n_n5120) & (!n_n5126)) + ((n_n5129) & (!n_n5124) & (!n_n5120) & (n_n5126)) + ((n_n5129) & (!n_n5124) & (n_n5120) & (!n_n5126)) + ((n_n5129) & (!n_n5124) & (n_n5120) & (n_n5126)) + ((n_n5129) & (n_n5124) & (!n_n5120) & (!n_n5126)) + ((n_n5129) & (n_n5124) & (!n_n5120) & (n_n5126)) + ((n_n5129) & (n_n5124) & (n_n5120) & (!n_n5126)) + ((n_n5129) & (n_n5124) & (n_n5120) & (n_n5126)));
	assign x12920x = (((!n_n524) & (!n_n528) & (!n_n509) & (!x12x) & (n_n5119)) + ((!n_n524) & (!n_n528) & (!n_n509) & (x12x) & (n_n5119)) + ((!n_n524) & (!n_n528) & (n_n509) & (!x12x) & (n_n5119)) + ((!n_n524) & (!n_n528) & (n_n509) & (x12x) & (n_n5119)) + ((!n_n524) & (n_n528) & (!n_n509) & (!x12x) & (n_n5119)) + ((!n_n524) & (n_n528) & (!n_n509) & (x12x) & (n_n5119)) + ((!n_n524) & (n_n528) & (n_n509) & (!x12x) & (n_n5119)) + ((!n_n524) & (n_n528) & (n_n509) & (x12x) & (!n_n5119)) + ((!n_n524) & (n_n528) & (n_n509) & (x12x) & (n_n5119)) + ((n_n524) & (!n_n528) & (!n_n509) & (!x12x) & (n_n5119)) + ((n_n524) & (!n_n528) & (!n_n509) & (x12x) & (n_n5119)) + ((n_n524) & (!n_n528) & (n_n509) & (!x12x) & (n_n5119)) + ((n_n524) & (!n_n528) & (n_n509) & (x12x) & (!n_n5119)) + ((n_n524) & (!n_n528) & (n_n509) & (x12x) & (n_n5119)) + ((n_n524) & (n_n528) & (!n_n509) & (!x12x) & (n_n5119)) + ((n_n524) & (n_n528) & (!n_n509) & (x12x) & (n_n5119)) + ((n_n524) & (n_n528) & (n_n509) & (!x12x) & (n_n5119)) + ((n_n524) & (n_n528) & (n_n509) & (x12x) & (!n_n5119)) + ((n_n524) & (n_n528) & (n_n509) & (x12x) & (n_n5119)));
	assign x12922x = (((!n_n509) & (!n_n130) & (!x23x) & (!n_n5128) & (x12920x)) + ((!n_n509) & (!n_n130) & (!x23x) & (n_n5128) & (!x12920x)) + ((!n_n509) & (!n_n130) & (!x23x) & (n_n5128) & (x12920x)) + ((!n_n509) & (!n_n130) & (x23x) & (!n_n5128) & (x12920x)) + ((!n_n509) & (!n_n130) & (x23x) & (n_n5128) & (!x12920x)) + ((!n_n509) & (!n_n130) & (x23x) & (n_n5128) & (x12920x)) + ((!n_n509) & (n_n130) & (!x23x) & (!n_n5128) & (x12920x)) + ((!n_n509) & (n_n130) & (!x23x) & (n_n5128) & (!x12920x)) + ((!n_n509) & (n_n130) & (!x23x) & (n_n5128) & (x12920x)) + ((!n_n509) & (n_n130) & (x23x) & (!n_n5128) & (x12920x)) + ((!n_n509) & (n_n130) & (x23x) & (n_n5128) & (!x12920x)) + ((!n_n509) & (n_n130) & (x23x) & (n_n5128) & (x12920x)) + ((n_n509) & (!n_n130) & (!x23x) & (!n_n5128) & (x12920x)) + ((n_n509) & (!n_n130) & (!x23x) & (n_n5128) & (!x12920x)) + ((n_n509) & (!n_n130) & (!x23x) & (n_n5128) & (x12920x)) + ((n_n509) & (!n_n130) & (x23x) & (!n_n5128) & (x12920x)) + ((n_n509) & (!n_n130) & (x23x) & (n_n5128) & (!x12920x)) + ((n_n509) & (!n_n130) & (x23x) & (n_n5128) & (x12920x)) + ((n_n509) & (n_n130) & (!x23x) & (!n_n5128) & (x12920x)) + ((n_n509) & (n_n130) & (!x23x) & (n_n5128) & (!x12920x)) + ((n_n509) & (n_n130) & (!x23x) & (n_n5128) & (x12920x)) + ((n_n509) & (n_n130) & (x23x) & (!n_n5128) & (!x12920x)) + ((n_n509) & (n_n130) & (x23x) & (!n_n5128) & (x12920x)) + ((n_n509) & (n_n130) & (x23x) & (n_n5128) & (!x12920x)) + ((n_n509) & (n_n130) & (x23x) & (n_n5128) & (x12920x)));
	assign x12929x = (((!n_n5102) & (!n_n5106) & (!x28x) & (n_n783)) + ((!n_n5102) & (!n_n5106) & (x28x) & (!n_n783)) + ((!n_n5102) & (!n_n5106) & (x28x) & (n_n783)) + ((!n_n5102) & (n_n5106) & (!x28x) & (!n_n783)) + ((!n_n5102) & (n_n5106) & (!x28x) & (n_n783)) + ((!n_n5102) & (n_n5106) & (x28x) & (!n_n783)) + ((!n_n5102) & (n_n5106) & (x28x) & (n_n783)) + ((n_n5102) & (!n_n5106) & (!x28x) & (!n_n783)) + ((n_n5102) & (!n_n5106) & (!x28x) & (n_n783)) + ((n_n5102) & (!n_n5106) & (x28x) & (!n_n783)) + ((n_n5102) & (!n_n5106) & (x28x) & (n_n783)) + ((n_n5102) & (n_n5106) & (!x28x) & (!n_n783)) + ((n_n5102) & (n_n5106) & (!x28x) & (n_n783)) + ((n_n5102) & (n_n5106) & (x28x) & (!n_n783)) + ((n_n5102) & (n_n5106) & (x28x) & (n_n783)));
	assign x12928x = (((!n_n5112) & (!n_n5086) & (!x290x) & (!x122x) & (x143x)) + ((!n_n5112) & (!n_n5086) & (!x290x) & (x122x) & (!x143x)) + ((!n_n5112) & (!n_n5086) & (!x290x) & (x122x) & (x143x)) + ((!n_n5112) & (!n_n5086) & (x290x) & (!x122x) & (!x143x)) + ((!n_n5112) & (!n_n5086) & (x290x) & (!x122x) & (x143x)) + ((!n_n5112) & (!n_n5086) & (x290x) & (x122x) & (!x143x)) + ((!n_n5112) & (!n_n5086) & (x290x) & (x122x) & (x143x)) + ((!n_n5112) & (n_n5086) & (!x290x) & (!x122x) & (!x143x)) + ((!n_n5112) & (n_n5086) & (!x290x) & (!x122x) & (x143x)) + ((!n_n5112) & (n_n5086) & (!x290x) & (x122x) & (!x143x)) + ((!n_n5112) & (n_n5086) & (!x290x) & (x122x) & (x143x)) + ((!n_n5112) & (n_n5086) & (x290x) & (!x122x) & (!x143x)) + ((!n_n5112) & (n_n5086) & (x290x) & (!x122x) & (x143x)) + ((!n_n5112) & (n_n5086) & (x290x) & (x122x) & (!x143x)) + ((!n_n5112) & (n_n5086) & (x290x) & (x122x) & (x143x)) + ((n_n5112) & (!n_n5086) & (!x290x) & (!x122x) & (!x143x)) + ((n_n5112) & (!n_n5086) & (!x290x) & (!x122x) & (x143x)) + ((n_n5112) & (!n_n5086) & (!x290x) & (x122x) & (!x143x)) + ((n_n5112) & (!n_n5086) & (!x290x) & (x122x) & (x143x)) + ((n_n5112) & (!n_n5086) & (x290x) & (!x122x) & (!x143x)) + ((n_n5112) & (!n_n5086) & (x290x) & (!x122x) & (x143x)) + ((n_n5112) & (!n_n5086) & (x290x) & (x122x) & (!x143x)) + ((n_n5112) & (!n_n5086) & (x290x) & (x122x) & (x143x)) + ((n_n5112) & (n_n5086) & (!x290x) & (!x122x) & (!x143x)) + ((n_n5112) & (n_n5086) & (!x290x) & (!x122x) & (x143x)) + ((n_n5112) & (n_n5086) & (!x290x) & (x122x) & (!x143x)) + ((n_n5112) & (n_n5086) & (!x290x) & (x122x) & (x143x)) + ((n_n5112) & (n_n5086) & (x290x) & (!x122x) & (!x143x)) + ((n_n5112) & (n_n5086) & (x290x) & (!x122x) & (x143x)) + ((n_n5112) & (n_n5086) & (x290x) & (x122x) & (!x143x)) + ((n_n5112) & (n_n5086) & (x290x) & (x122x) & (x143x)));
	assign n_n638 = (((!x12921x) & (!x12922x) & (!x12929x) & (x12928x)) + ((!x12921x) & (!x12922x) & (x12929x) & (!x12928x)) + ((!x12921x) & (!x12922x) & (x12929x) & (x12928x)) + ((!x12921x) & (x12922x) & (!x12929x) & (!x12928x)) + ((!x12921x) & (x12922x) & (!x12929x) & (x12928x)) + ((!x12921x) & (x12922x) & (x12929x) & (!x12928x)) + ((!x12921x) & (x12922x) & (x12929x) & (x12928x)) + ((x12921x) & (!x12922x) & (!x12929x) & (!x12928x)) + ((x12921x) & (!x12922x) & (!x12929x) & (x12928x)) + ((x12921x) & (!x12922x) & (x12929x) & (!x12928x)) + ((x12921x) & (!x12922x) & (x12929x) & (x12928x)) + ((x12921x) & (x12922x) & (!x12929x) & (!x12928x)) + ((x12921x) & (x12922x) & (!x12929x) & (x12928x)) + ((x12921x) & (x12922x) & (x12929x) & (!x12928x)) + ((x12921x) & (x12922x) & (x12929x) & (x12928x)));
	assign n_n684 = (((!n_n5007) & (!n_n5016) & (!n_n3427) & (!x297x) & (x394x)) + ((!n_n5007) & (!n_n5016) & (!n_n3427) & (x297x) & (!x394x)) + ((!n_n5007) & (!n_n5016) & (!n_n3427) & (x297x) & (x394x)) + ((!n_n5007) & (!n_n5016) & (n_n3427) & (!x297x) & (!x394x)) + ((!n_n5007) & (!n_n5016) & (n_n3427) & (!x297x) & (x394x)) + ((!n_n5007) & (!n_n5016) & (n_n3427) & (x297x) & (!x394x)) + ((!n_n5007) & (!n_n5016) & (n_n3427) & (x297x) & (x394x)) + ((!n_n5007) & (n_n5016) & (!n_n3427) & (!x297x) & (!x394x)) + ((!n_n5007) & (n_n5016) & (!n_n3427) & (!x297x) & (x394x)) + ((!n_n5007) & (n_n5016) & (!n_n3427) & (x297x) & (!x394x)) + ((!n_n5007) & (n_n5016) & (!n_n3427) & (x297x) & (x394x)) + ((!n_n5007) & (n_n5016) & (n_n3427) & (!x297x) & (!x394x)) + ((!n_n5007) & (n_n5016) & (n_n3427) & (!x297x) & (x394x)) + ((!n_n5007) & (n_n5016) & (n_n3427) & (x297x) & (!x394x)) + ((!n_n5007) & (n_n5016) & (n_n3427) & (x297x) & (x394x)) + ((n_n5007) & (!n_n5016) & (!n_n3427) & (!x297x) & (!x394x)) + ((n_n5007) & (!n_n5016) & (!n_n3427) & (!x297x) & (x394x)) + ((n_n5007) & (!n_n5016) & (!n_n3427) & (x297x) & (!x394x)) + ((n_n5007) & (!n_n5016) & (!n_n3427) & (x297x) & (x394x)) + ((n_n5007) & (!n_n5016) & (n_n3427) & (!x297x) & (!x394x)) + ((n_n5007) & (!n_n5016) & (n_n3427) & (!x297x) & (x394x)) + ((n_n5007) & (!n_n5016) & (n_n3427) & (x297x) & (!x394x)) + ((n_n5007) & (!n_n5016) & (n_n3427) & (x297x) & (x394x)) + ((n_n5007) & (n_n5016) & (!n_n3427) & (!x297x) & (!x394x)) + ((n_n5007) & (n_n5016) & (!n_n3427) & (!x297x) & (x394x)) + ((n_n5007) & (n_n5016) & (!n_n3427) & (x297x) & (!x394x)) + ((n_n5007) & (n_n5016) & (!n_n3427) & (x297x) & (x394x)) + ((n_n5007) & (n_n5016) & (n_n3427) & (!x297x) & (!x394x)) + ((n_n5007) & (n_n5016) & (n_n3427) & (!x297x) & (x394x)) + ((n_n5007) & (n_n5016) & (n_n3427) & (x297x) & (!x394x)) + ((n_n5007) & (n_n5016) & (n_n3427) & (x297x) & (x394x)));
	assign x12939x = (((!n_n5031) & (!n_n5023) & (!n_n5029) & (x253x)) + ((!n_n5031) & (!n_n5023) & (n_n5029) & (!x253x)) + ((!n_n5031) & (!n_n5023) & (n_n5029) & (x253x)) + ((!n_n5031) & (n_n5023) & (!n_n5029) & (!x253x)) + ((!n_n5031) & (n_n5023) & (!n_n5029) & (x253x)) + ((!n_n5031) & (n_n5023) & (n_n5029) & (!x253x)) + ((!n_n5031) & (n_n5023) & (n_n5029) & (x253x)) + ((n_n5031) & (!n_n5023) & (!n_n5029) & (!x253x)) + ((n_n5031) & (!n_n5023) & (!n_n5029) & (x253x)) + ((n_n5031) & (!n_n5023) & (n_n5029) & (!x253x)) + ((n_n5031) & (!n_n5023) & (n_n5029) & (x253x)) + ((n_n5031) & (n_n5023) & (!n_n5029) & (!x253x)) + ((n_n5031) & (n_n5023) & (!n_n5029) & (x253x)) + ((n_n5031) & (n_n5023) & (n_n5029) & (!x253x)) + ((n_n5031) & (n_n5023) & (n_n5029) & (x253x)));
	assign n_n683 = (((!x492x) & (!x18x) & (!n_n5026) & (!x12939x) & (x265x)) + ((!x492x) & (!x18x) & (!n_n5026) & (x12939x) & (!x265x)) + ((!x492x) & (!x18x) & (!n_n5026) & (x12939x) & (x265x)) + ((!x492x) & (!x18x) & (n_n5026) & (!x12939x) & (!x265x)) + ((!x492x) & (!x18x) & (n_n5026) & (!x12939x) & (x265x)) + ((!x492x) & (!x18x) & (n_n5026) & (x12939x) & (!x265x)) + ((!x492x) & (!x18x) & (n_n5026) & (x12939x) & (x265x)) + ((!x492x) & (x18x) & (!n_n5026) & (!x12939x) & (x265x)) + ((!x492x) & (x18x) & (!n_n5026) & (x12939x) & (!x265x)) + ((!x492x) & (x18x) & (!n_n5026) & (x12939x) & (x265x)) + ((!x492x) & (x18x) & (n_n5026) & (!x12939x) & (!x265x)) + ((!x492x) & (x18x) & (n_n5026) & (!x12939x) & (x265x)) + ((!x492x) & (x18x) & (n_n5026) & (x12939x) & (!x265x)) + ((!x492x) & (x18x) & (n_n5026) & (x12939x) & (x265x)) + ((x492x) & (!x18x) & (!n_n5026) & (!x12939x) & (x265x)) + ((x492x) & (!x18x) & (!n_n5026) & (x12939x) & (!x265x)) + ((x492x) & (!x18x) & (!n_n5026) & (x12939x) & (x265x)) + ((x492x) & (!x18x) & (n_n5026) & (!x12939x) & (!x265x)) + ((x492x) & (!x18x) & (n_n5026) & (!x12939x) & (x265x)) + ((x492x) & (!x18x) & (n_n5026) & (x12939x) & (!x265x)) + ((x492x) & (!x18x) & (n_n5026) & (x12939x) & (x265x)) + ((x492x) & (x18x) & (!n_n5026) & (!x12939x) & (!x265x)) + ((x492x) & (x18x) & (!n_n5026) & (!x12939x) & (x265x)) + ((x492x) & (x18x) & (!n_n5026) & (x12939x) & (!x265x)) + ((x492x) & (x18x) & (!n_n5026) & (x12939x) & (x265x)) + ((x492x) & (x18x) & (n_n5026) & (!x12939x) & (!x265x)) + ((x492x) & (x18x) & (n_n5026) & (!x12939x) & (x265x)) + ((x492x) & (x18x) & (n_n5026) & (x12939x) & (!x265x)) + ((x492x) & (x18x) & (n_n5026) & (x12939x) & (x265x)));
	assign x12945x = (((!n_n5034) & (!n_n5035) & (!n_n5039) & (!x153x) & (!x22129x)) + ((!n_n5034) & (!n_n5035) & (!n_n5039) & (x153x) & (!x22129x)) + ((!n_n5034) & (!n_n5035) & (!n_n5039) & (x153x) & (x22129x)) + ((!n_n5034) & (!n_n5035) & (n_n5039) & (!x153x) & (!x22129x)) + ((!n_n5034) & (!n_n5035) & (n_n5039) & (!x153x) & (x22129x)) + ((!n_n5034) & (!n_n5035) & (n_n5039) & (x153x) & (!x22129x)) + ((!n_n5034) & (!n_n5035) & (n_n5039) & (x153x) & (x22129x)) + ((!n_n5034) & (n_n5035) & (!n_n5039) & (!x153x) & (!x22129x)) + ((!n_n5034) & (n_n5035) & (!n_n5039) & (!x153x) & (x22129x)) + ((!n_n5034) & (n_n5035) & (!n_n5039) & (x153x) & (!x22129x)) + ((!n_n5034) & (n_n5035) & (!n_n5039) & (x153x) & (x22129x)) + ((!n_n5034) & (n_n5035) & (n_n5039) & (!x153x) & (!x22129x)) + ((!n_n5034) & (n_n5035) & (n_n5039) & (!x153x) & (x22129x)) + ((!n_n5034) & (n_n5035) & (n_n5039) & (x153x) & (!x22129x)) + ((!n_n5034) & (n_n5035) & (n_n5039) & (x153x) & (x22129x)) + ((n_n5034) & (!n_n5035) & (!n_n5039) & (!x153x) & (!x22129x)) + ((n_n5034) & (!n_n5035) & (!n_n5039) & (!x153x) & (x22129x)) + ((n_n5034) & (!n_n5035) & (!n_n5039) & (x153x) & (!x22129x)) + ((n_n5034) & (!n_n5035) & (!n_n5039) & (x153x) & (x22129x)) + ((n_n5034) & (!n_n5035) & (n_n5039) & (!x153x) & (!x22129x)) + ((n_n5034) & (!n_n5035) & (n_n5039) & (!x153x) & (x22129x)) + ((n_n5034) & (!n_n5035) & (n_n5039) & (x153x) & (!x22129x)) + ((n_n5034) & (!n_n5035) & (n_n5039) & (x153x) & (x22129x)) + ((n_n5034) & (n_n5035) & (!n_n5039) & (!x153x) & (!x22129x)) + ((n_n5034) & (n_n5035) & (!n_n5039) & (!x153x) & (x22129x)) + ((n_n5034) & (n_n5035) & (!n_n5039) & (x153x) & (!x22129x)) + ((n_n5034) & (n_n5035) & (!n_n5039) & (x153x) & (x22129x)) + ((n_n5034) & (n_n5035) & (n_n5039) & (!x153x) & (!x22129x)) + ((n_n5034) & (n_n5035) & (n_n5039) & (!x153x) & (x22129x)) + ((n_n5034) & (n_n5035) & (n_n5039) & (x153x) & (!x22129x)) + ((n_n5034) & (n_n5035) & (n_n5039) & (x153x) & (x22129x)));
	assign x12947x = (((!n_n684) & (!n_n683) & (x12945x)) + ((!n_n684) & (n_n683) & (!x12945x)) + ((!n_n684) & (n_n683) & (x12945x)) + ((n_n684) & (!n_n683) & (!x12945x)) + ((n_n684) & (!n_n683) & (x12945x)) + ((n_n684) & (n_n683) & (!x12945x)) + ((n_n684) & (n_n683) & (x12945x)));
	assign x13533x = (((!n_n4389) & (!n_n4393) & (!n_n4384) & (!n_n4390) & (n_n4394)) + ((!n_n4389) & (!n_n4393) & (!n_n4384) & (n_n4390) & (!n_n4394)) + ((!n_n4389) & (!n_n4393) & (!n_n4384) & (n_n4390) & (n_n4394)) + ((!n_n4389) & (!n_n4393) & (n_n4384) & (!n_n4390) & (!n_n4394)) + ((!n_n4389) & (!n_n4393) & (n_n4384) & (!n_n4390) & (n_n4394)) + ((!n_n4389) & (!n_n4393) & (n_n4384) & (n_n4390) & (!n_n4394)) + ((!n_n4389) & (!n_n4393) & (n_n4384) & (n_n4390) & (n_n4394)) + ((!n_n4389) & (n_n4393) & (!n_n4384) & (!n_n4390) & (!n_n4394)) + ((!n_n4389) & (n_n4393) & (!n_n4384) & (!n_n4390) & (n_n4394)) + ((!n_n4389) & (n_n4393) & (!n_n4384) & (n_n4390) & (!n_n4394)) + ((!n_n4389) & (n_n4393) & (!n_n4384) & (n_n4390) & (n_n4394)) + ((!n_n4389) & (n_n4393) & (n_n4384) & (!n_n4390) & (!n_n4394)) + ((!n_n4389) & (n_n4393) & (n_n4384) & (!n_n4390) & (n_n4394)) + ((!n_n4389) & (n_n4393) & (n_n4384) & (n_n4390) & (!n_n4394)) + ((!n_n4389) & (n_n4393) & (n_n4384) & (n_n4390) & (n_n4394)) + ((n_n4389) & (!n_n4393) & (!n_n4384) & (!n_n4390) & (!n_n4394)) + ((n_n4389) & (!n_n4393) & (!n_n4384) & (!n_n4390) & (n_n4394)) + ((n_n4389) & (!n_n4393) & (!n_n4384) & (n_n4390) & (!n_n4394)) + ((n_n4389) & (!n_n4393) & (!n_n4384) & (n_n4390) & (n_n4394)) + ((n_n4389) & (!n_n4393) & (n_n4384) & (!n_n4390) & (!n_n4394)) + ((n_n4389) & (!n_n4393) & (n_n4384) & (!n_n4390) & (n_n4394)) + ((n_n4389) & (!n_n4393) & (n_n4384) & (n_n4390) & (!n_n4394)) + ((n_n4389) & (!n_n4393) & (n_n4384) & (n_n4390) & (n_n4394)) + ((n_n4389) & (n_n4393) & (!n_n4384) & (!n_n4390) & (!n_n4394)) + ((n_n4389) & (n_n4393) & (!n_n4384) & (!n_n4390) & (n_n4394)) + ((n_n4389) & (n_n4393) & (!n_n4384) & (n_n4390) & (!n_n4394)) + ((n_n4389) & (n_n4393) & (!n_n4384) & (n_n4390) & (n_n4394)) + ((n_n4389) & (n_n4393) & (n_n4384) & (!n_n4390) & (!n_n4394)) + ((n_n4389) & (n_n4393) & (n_n4384) & (!n_n4390) & (n_n4394)) + ((n_n4389) & (n_n4393) & (n_n4384) & (n_n4390) & (!n_n4394)) + ((n_n4389) & (n_n4393) & (n_n4384) & (n_n4390) & (n_n4394)));
	assign x13538x = (((!n_n4400) & (!n_n4404) & (!n_n4405) & (!n_n4406) & (n_n4396)) + ((!n_n4400) & (!n_n4404) & (!n_n4405) & (n_n4406) & (!n_n4396)) + ((!n_n4400) & (!n_n4404) & (!n_n4405) & (n_n4406) & (n_n4396)) + ((!n_n4400) & (!n_n4404) & (n_n4405) & (!n_n4406) & (!n_n4396)) + ((!n_n4400) & (!n_n4404) & (n_n4405) & (!n_n4406) & (n_n4396)) + ((!n_n4400) & (!n_n4404) & (n_n4405) & (n_n4406) & (!n_n4396)) + ((!n_n4400) & (!n_n4404) & (n_n4405) & (n_n4406) & (n_n4396)) + ((!n_n4400) & (n_n4404) & (!n_n4405) & (!n_n4406) & (!n_n4396)) + ((!n_n4400) & (n_n4404) & (!n_n4405) & (!n_n4406) & (n_n4396)) + ((!n_n4400) & (n_n4404) & (!n_n4405) & (n_n4406) & (!n_n4396)) + ((!n_n4400) & (n_n4404) & (!n_n4405) & (n_n4406) & (n_n4396)) + ((!n_n4400) & (n_n4404) & (n_n4405) & (!n_n4406) & (!n_n4396)) + ((!n_n4400) & (n_n4404) & (n_n4405) & (!n_n4406) & (n_n4396)) + ((!n_n4400) & (n_n4404) & (n_n4405) & (n_n4406) & (!n_n4396)) + ((!n_n4400) & (n_n4404) & (n_n4405) & (n_n4406) & (n_n4396)) + ((n_n4400) & (!n_n4404) & (!n_n4405) & (!n_n4406) & (!n_n4396)) + ((n_n4400) & (!n_n4404) & (!n_n4405) & (!n_n4406) & (n_n4396)) + ((n_n4400) & (!n_n4404) & (!n_n4405) & (n_n4406) & (!n_n4396)) + ((n_n4400) & (!n_n4404) & (!n_n4405) & (n_n4406) & (n_n4396)) + ((n_n4400) & (!n_n4404) & (n_n4405) & (!n_n4406) & (!n_n4396)) + ((n_n4400) & (!n_n4404) & (n_n4405) & (!n_n4406) & (n_n4396)) + ((n_n4400) & (!n_n4404) & (n_n4405) & (n_n4406) & (!n_n4396)) + ((n_n4400) & (!n_n4404) & (n_n4405) & (n_n4406) & (n_n4396)) + ((n_n4400) & (n_n4404) & (!n_n4405) & (!n_n4406) & (!n_n4396)) + ((n_n4400) & (n_n4404) & (!n_n4405) & (!n_n4406) & (n_n4396)) + ((n_n4400) & (n_n4404) & (!n_n4405) & (n_n4406) & (!n_n4396)) + ((n_n4400) & (n_n4404) & (!n_n4405) & (n_n4406) & (n_n4396)) + ((n_n4400) & (n_n4404) & (n_n4405) & (!n_n4406) & (!n_n4396)) + ((n_n4400) & (n_n4404) & (n_n4405) & (!n_n4406) & (n_n4396)) + ((n_n4400) & (n_n4404) & (n_n4405) & (n_n4406) & (!n_n4396)) + ((n_n4400) & (n_n4404) & (n_n4405) & (n_n4406) & (n_n4396)));
	assign x13539x = (((!n_n4401) & (!n_n4403) & (!n_n4397) & (!n_n4398) & (x13538x)) + ((!n_n4401) & (!n_n4403) & (!n_n4397) & (n_n4398) & (!x13538x)) + ((!n_n4401) & (!n_n4403) & (!n_n4397) & (n_n4398) & (x13538x)) + ((!n_n4401) & (!n_n4403) & (n_n4397) & (!n_n4398) & (!x13538x)) + ((!n_n4401) & (!n_n4403) & (n_n4397) & (!n_n4398) & (x13538x)) + ((!n_n4401) & (!n_n4403) & (n_n4397) & (n_n4398) & (!x13538x)) + ((!n_n4401) & (!n_n4403) & (n_n4397) & (n_n4398) & (x13538x)) + ((!n_n4401) & (n_n4403) & (!n_n4397) & (!n_n4398) & (!x13538x)) + ((!n_n4401) & (n_n4403) & (!n_n4397) & (!n_n4398) & (x13538x)) + ((!n_n4401) & (n_n4403) & (!n_n4397) & (n_n4398) & (!x13538x)) + ((!n_n4401) & (n_n4403) & (!n_n4397) & (n_n4398) & (x13538x)) + ((!n_n4401) & (n_n4403) & (n_n4397) & (!n_n4398) & (!x13538x)) + ((!n_n4401) & (n_n4403) & (n_n4397) & (!n_n4398) & (x13538x)) + ((!n_n4401) & (n_n4403) & (n_n4397) & (n_n4398) & (!x13538x)) + ((!n_n4401) & (n_n4403) & (n_n4397) & (n_n4398) & (x13538x)) + ((n_n4401) & (!n_n4403) & (!n_n4397) & (!n_n4398) & (!x13538x)) + ((n_n4401) & (!n_n4403) & (!n_n4397) & (!n_n4398) & (x13538x)) + ((n_n4401) & (!n_n4403) & (!n_n4397) & (n_n4398) & (!x13538x)) + ((n_n4401) & (!n_n4403) & (!n_n4397) & (n_n4398) & (x13538x)) + ((n_n4401) & (!n_n4403) & (n_n4397) & (!n_n4398) & (!x13538x)) + ((n_n4401) & (!n_n4403) & (n_n4397) & (!n_n4398) & (x13538x)) + ((n_n4401) & (!n_n4403) & (n_n4397) & (n_n4398) & (!x13538x)) + ((n_n4401) & (!n_n4403) & (n_n4397) & (n_n4398) & (x13538x)) + ((n_n4401) & (n_n4403) & (!n_n4397) & (!n_n4398) & (!x13538x)) + ((n_n4401) & (n_n4403) & (!n_n4397) & (!n_n4398) & (x13538x)) + ((n_n4401) & (n_n4403) & (!n_n4397) & (n_n4398) & (!x13538x)) + ((n_n4401) & (n_n4403) & (!n_n4397) & (n_n4398) & (x13538x)) + ((n_n4401) & (n_n4403) & (n_n4397) & (!n_n4398) & (!x13538x)) + ((n_n4401) & (n_n4403) & (n_n4397) & (!n_n4398) & (x13538x)) + ((n_n4401) & (n_n4403) & (n_n4397) & (n_n4398) & (!x13538x)) + ((n_n4401) & (n_n4403) & (n_n4397) & (n_n4398) & (x13538x)));
	assign x13943x = (((!x592x) & (!x20x) & (!n_n5308) & (!x200x) & (n_n5304)) + ((!x592x) & (!x20x) & (!n_n5308) & (x200x) & (!n_n5304)) + ((!x592x) & (!x20x) & (!n_n5308) & (x200x) & (n_n5304)) + ((!x592x) & (!x20x) & (n_n5308) & (!x200x) & (!n_n5304)) + ((!x592x) & (!x20x) & (n_n5308) & (!x200x) & (n_n5304)) + ((!x592x) & (!x20x) & (n_n5308) & (x200x) & (!n_n5304)) + ((!x592x) & (!x20x) & (n_n5308) & (x200x) & (n_n5304)) + ((!x592x) & (x20x) & (!n_n5308) & (!x200x) & (n_n5304)) + ((!x592x) & (x20x) & (!n_n5308) & (x200x) & (!n_n5304)) + ((!x592x) & (x20x) & (!n_n5308) & (x200x) & (n_n5304)) + ((!x592x) & (x20x) & (n_n5308) & (!x200x) & (!n_n5304)) + ((!x592x) & (x20x) & (n_n5308) & (!x200x) & (n_n5304)) + ((!x592x) & (x20x) & (n_n5308) & (x200x) & (!n_n5304)) + ((!x592x) & (x20x) & (n_n5308) & (x200x) & (n_n5304)) + ((x592x) & (!x20x) & (!n_n5308) & (!x200x) & (n_n5304)) + ((x592x) & (!x20x) & (!n_n5308) & (x200x) & (!n_n5304)) + ((x592x) & (!x20x) & (!n_n5308) & (x200x) & (n_n5304)) + ((x592x) & (!x20x) & (n_n5308) & (!x200x) & (!n_n5304)) + ((x592x) & (!x20x) & (n_n5308) & (!x200x) & (n_n5304)) + ((x592x) & (!x20x) & (n_n5308) & (x200x) & (!n_n5304)) + ((x592x) & (!x20x) & (n_n5308) & (x200x) & (n_n5304)) + ((x592x) & (x20x) & (!n_n5308) & (!x200x) & (!n_n5304)) + ((x592x) & (x20x) & (!n_n5308) & (!x200x) & (n_n5304)) + ((x592x) & (x20x) & (!n_n5308) & (x200x) & (!n_n5304)) + ((x592x) & (x20x) & (!n_n5308) & (x200x) & (n_n5304)) + ((x592x) & (x20x) & (n_n5308) & (!x200x) & (!n_n5304)) + ((x592x) & (x20x) & (n_n5308) & (!x200x) & (n_n5304)) + ((x592x) & (x20x) & (n_n5308) & (x200x) & (!n_n5304)) + ((x592x) & (x20x) & (n_n5308) & (x200x) & (n_n5304)));
	assign x434x = (((!i_9_) & (!n_n524) & (n_n509) & (x20x) & (n_n65)) + ((!i_9_) & (n_n524) & (n_n509) & (!x20x) & (n_n65)) + ((!i_9_) & (n_n524) & (n_n509) & (x20x) & (n_n65)) + ((i_9_) & (!n_n524) & (n_n509) & (x20x) & (n_n65)) + ((i_9_) & (n_n524) & (n_n509) & (x20x) & (n_n65)));
	assign x12476x = (((!x20x) & (!n_n4447) & (!x496x) & (!n_n4435) & (x421x)) + ((!x20x) & (!n_n4447) & (!x496x) & (n_n4435) & (!x421x)) + ((!x20x) & (!n_n4447) & (!x496x) & (n_n4435) & (x421x)) + ((!x20x) & (!n_n4447) & (x496x) & (!n_n4435) & (x421x)) + ((!x20x) & (!n_n4447) & (x496x) & (n_n4435) & (!x421x)) + ((!x20x) & (!n_n4447) & (x496x) & (n_n4435) & (x421x)) + ((!x20x) & (n_n4447) & (!x496x) & (!n_n4435) & (!x421x)) + ((!x20x) & (n_n4447) & (!x496x) & (!n_n4435) & (x421x)) + ((!x20x) & (n_n4447) & (!x496x) & (n_n4435) & (!x421x)) + ((!x20x) & (n_n4447) & (!x496x) & (n_n4435) & (x421x)) + ((!x20x) & (n_n4447) & (x496x) & (!n_n4435) & (!x421x)) + ((!x20x) & (n_n4447) & (x496x) & (!n_n4435) & (x421x)) + ((!x20x) & (n_n4447) & (x496x) & (n_n4435) & (!x421x)) + ((!x20x) & (n_n4447) & (x496x) & (n_n4435) & (x421x)) + ((x20x) & (!n_n4447) & (!x496x) & (!n_n4435) & (x421x)) + ((x20x) & (!n_n4447) & (!x496x) & (n_n4435) & (!x421x)) + ((x20x) & (!n_n4447) & (!x496x) & (n_n4435) & (x421x)) + ((x20x) & (!n_n4447) & (x496x) & (!n_n4435) & (!x421x)) + ((x20x) & (!n_n4447) & (x496x) & (!n_n4435) & (x421x)) + ((x20x) & (!n_n4447) & (x496x) & (n_n4435) & (!x421x)) + ((x20x) & (!n_n4447) & (x496x) & (n_n4435) & (x421x)) + ((x20x) & (n_n4447) & (!x496x) & (!n_n4435) & (!x421x)) + ((x20x) & (n_n4447) & (!x496x) & (!n_n4435) & (x421x)) + ((x20x) & (n_n4447) & (!x496x) & (n_n4435) & (!x421x)) + ((x20x) & (n_n4447) & (!x496x) & (n_n4435) & (x421x)) + ((x20x) & (n_n4447) & (x496x) & (!n_n4435) & (!x421x)) + ((x20x) & (n_n4447) & (x496x) & (!n_n4435) & (x421x)) + ((x20x) & (n_n4447) & (x496x) & (n_n4435) & (!x421x)) + ((x20x) & (n_n4447) & (x496x) & (n_n4435) & (x421x)));
	assign n_n2058 = (((!i_9_) & (n_n518) & (n_n455) & (!n_n532) & (n_n534)) + ((!i_9_) & (n_n518) & (n_n455) & (n_n532) & (!n_n534)) + ((!i_9_) & (n_n518) & (n_n455) & (n_n532) & (n_n534)) + ((i_9_) & (n_n518) & (n_n455) & (!n_n532) & (n_n534)) + ((i_9_) & (n_n518) & (n_n455) & (n_n532) & (n_n534)));
	assign x12485x = (((!n_n4448) & (!n_n4451) & (!n_n3162) & (!x55x) & (n_n2058)) + ((!n_n4448) & (!n_n4451) & (!n_n3162) & (x55x) & (!n_n2058)) + ((!n_n4448) & (!n_n4451) & (!n_n3162) & (x55x) & (n_n2058)) + ((!n_n4448) & (!n_n4451) & (n_n3162) & (!x55x) & (!n_n2058)) + ((!n_n4448) & (!n_n4451) & (n_n3162) & (!x55x) & (n_n2058)) + ((!n_n4448) & (!n_n4451) & (n_n3162) & (x55x) & (!n_n2058)) + ((!n_n4448) & (!n_n4451) & (n_n3162) & (x55x) & (n_n2058)) + ((!n_n4448) & (n_n4451) & (!n_n3162) & (!x55x) & (!n_n2058)) + ((!n_n4448) & (n_n4451) & (!n_n3162) & (!x55x) & (n_n2058)) + ((!n_n4448) & (n_n4451) & (!n_n3162) & (x55x) & (!n_n2058)) + ((!n_n4448) & (n_n4451) & (!n_n3162) & (x55x) & (n_n2058)) + ((!n_n4448) & (n_n4451) & (n_n3162) & (!x55x) & (!n_n2058)) + ((!n_n4448) & (n_n4451) & (n_n3162) & (!x55x) & (n_n2058)) + ((!n_n4448) & (n_n4451) & (n_n3162) & (x55x) & (!n_n2058)) + ((!n_n4448) & (n_n4451) & (n_n3162) & (x55x) & (n_n2058)) + ((n_n4448) & (!n_n4451) & (!n_n3162) & (!x55x) & (!n_n2058)) + ((n_n4448) & (!n_n4451) & (!n_n3162) & (!x55x) & (n_n2058)) + ((n_n4448) & (!n_n4451) & (!n_n3162) & (x55x) & (!n_n2058)) + ((n_n4448) & (!n_n4451) & (!n_n3162) & (x55x) & (n_n2058)) + ((n_n4448) & (!n_n4451) & (n_n3162) & (!x55x) & (!n_n2058)) + ((n_n4448) & (!n_n4451) & (n_n3162) & (!x55x) & (n_n2058)) + ((n_n4448) & (!n_n4451) & (n_n3162) & (x55x) & (!n_n2058)) + ((n_n4448) & (!n_n4451) & (n_n3162) & (x55x) & (n_n2058)) + ((n_n4448) & (n_n4451) & (!n_n3162) & (!x55x) & (!n_n2058)) + ((n_n4448) & (n_n4451) & (!n_n3162) & (!x55x) & (n_n2058)) + ((n_n4448) & (n_n4451) & (!n_n3162) & (x55x) & (!n_n2058)) + ((n_n4448) & (n_n4451) & (!n_n3162) & (x55x) & (n_n2058)) + ((n_n4448) & (n_n4451) & (n_n3162) & (!x55x) & (!n_n2058)) + ((n_n4448) & (n_n4451) & (n_n3162) & (!x55x) & (n_n2058)) + ((n_n4448) & (n_n4451) & (n_n3162) & (x55x) & (!n_n2058)) + ((n_n4448) & (n_n4451) & (n_n3162) & (x55x) & (n_n2058)));
	assign x12481x = (((!i_9_) & (!n_n455) & (!n_n535) & (!n_n522) & (x128x)) + ((!i_9_) & (!n_n455) & (!n_n535) & (n_n522) & (x128x)) + ((!i_9_) & (!n_n455) & (n_n535) & (!n_n522) & (x128x)) + ((!i_9_) & (!n_n455) & (n_n535) & (n_n522) & (x128x)) + ((!i_9_) & (n_n455) & (!n_n535) & (!n_n522) & (x128x)) + ((!i_9_) & (n_n455) & (!n_n535) & (n_n522) & (x128x)) + ((!i_9_) & (n_n455) & (n_n535) & (!n_n522) & (x128x)) + ((!i_9_) & (n_n455) & (n_n535) & (n_n522) & (!x128x)) + ((!i_9_) & (n_n455) & (n_n535) & (n_n522) & (x128x)) + ((i_9_) & (!n_n455) & (!n_n535) & (!n_n522) & (x128x)) + ((i_9_) & (!n_n455) & (!n_n535) & (n_n522) & (x128x)) + ((i_9_) & (!n_n455) & (n_n535) & (!n_n522) & (x128x)) + ((i_9_) & (!n_n455) & (n_n535) & (n_n522) & (x128x)) + ((i_9_) & (n_n455) & (!n_n535) & (!n_n522) & (x128x)) + ((i_9_) & (n_n455) & (!n_n535) & (n_n522) & (x128x)) + ((i_9_) & (n_n455) & (n_n535) & (!n_n522) & (x128x)) + ((i_9_) & (n_n455) & (n_n535) & (n_n522) & (!x128x)) + ((i_9_) & (n_n455) & (n_n535) & (n_n522) & (x128x)));
	assign x22141x = (((!n_n4440) & (!n_n4444) & (!x147x) & (!x32x) & (!n_n4465)));
	assign x22146x = (((!n_n4856) & (!n_n4854) & (!n_n4860) & (!n_n4864)));
	assign x263x = (((!i_9_) & (!n_n524) & (n_n526) & (n_n260) & (n_n500)) + ((!i_9_) & (n_n524) & (n_n526) & (n_n260) & (n_n500)) + ((i_9_) & (n_n524) & (!n_n526) & (n_n260) & (n_n500)) + ((i_9_) & (n_n524) & (n_n526) & (n_n260) & (n_n500)));
	assign x324x = (((!i_9_) & (n_n534) & (n_n260) & (n_n500)) + ((i_9_) & (n_n534) & (n_n260) & (n_n500)));
	assign x12217x = (((!i_9_) & (!n_n524) & (n_n509) & (n_n260) & (x23x)) + ((!i_9_) & (n_n524) & (n_n509) & (n_n260) & (!x23x)) + ((!i_9_) & (n_n524) & (n_n509) & (n_n260) & (x23x)) + ((i_9_) & (!n_n524) & (n_n509) & (n_n260) & (x23x)) + ((i_9_) & (n_n524) & (n_n509) & (n_n260) & (x23x)));
	assign x12164x = (((!n_n260) & (!x23x) & (!n_n464) & (!n_n4952) & (x210x)) + ((!n_n260) & (!x23x) & (!n_n464) & (n_n4952) & (!x210x)) + ((!n_n260) & (!x23x) & (!n_n464) & (n_n4952) & (x210x)) + ((!n_n260) & (!x23x) & (n_n464) & (!n_n4952) & (x210x)) + ((!n_n260) & (!x23x) & (n_n464) & (n_n4952) & (!x210x)) + ((!n_n260) & (!x23x) & (n_n464) & (n_n4952) & (x210x)) + ((!n_n260) & (x23x) & (!n_n464) & (!n_n4952) & (x210x)) + ((!n_n260) & (x23x) & (!n_n464) & (n_n4952) & (!x210x)) + ((!n_n260) & (x23x) & (!n_n464) & (n_n4952) & (x210x)) + ((!n_n260) & (x23x) & (n_n464) & (!n_n4952) & (x210x)) + ((!n_n260) & (x23x) & (n_n464) & (n_n4952) & (!x210x)) + ((!n_n260) & (x23x) & (n_n464) & (n_n4952) & (x210x)) + ((n_n260) & (!x23x) & (!n_n464) & (!n_n4952) & (x210x)) + ((n_n260) & (!x23x) & (!n_n464) & (n_n4952) & (!x210x)) + ((n_n260) & (!x23x) & (!n_n464) & (n_n4952) & (x210x)) + ((n_n260) & (!x23x) & (n_n464) & (!n_n4952) & (x210x)) + ((n_n260) & (!x23x) & (n_n464) & (n_n4952) & (!x210x)) + ((n_n260) & (!x23x) & (n_n464) & (n_n4952) & (x210x)) + ((n_n260) & (x23x) & (!n_n464) & (!n_n4952) & (x210x)) + ((n_n260) & (x23x) & (!n_n464) & (n_n4952) & (!x210x)) + ((n_n260) & (x23x) & (!n_n464) & (n_n4952) & (x210x)) + ((n_n260) & (x23x) & (n_n464) & (!n_n4952) & (!x210x)) + ((n_n260) & (x23x) & (n_n464) & (!n_n4952) & (x210x)) + ((n_n260) & (x23x) & (n_n464) & (n_n4952) & (!x210x)) + ((n_n260) & (x23x) & (n_n464) & (n_n4952) & (x210x)));
	assign x12165x = (((!n_n4958) & (!n_n4953) & (!n_n4956) & (!n_n4957) & (n_n4961)) + ((!n_n4958) & (!n_n4953) & (!n_n4956) & (n_n4957) & (!n_n4961)) + ((!n_n4958) & (!n_n4953) & (!n_n4956) & (n_n4957) & (n_n4961)) + ((!n_n4958) & (!n_n4953) & (n_n4956) & (!n_n4957) & (!n_n4961)) + ((!n_n4958) & (!n_n4953) & (n_n4956) & (!n_n4957) & (n_n4961)) + ((!n_n4958) & (!n_n4953) & (n_n4956) & (n_n4957) & (!n_n4961)) + ((!n_n4958) & (!n_n4953) & (n_n4956) & (n_n4957) & (n_n4961)) + ((!n_n4958) & (n_n4953) & (!n_n4956) & (!n_n4957) & (!n_n4961)) + ((!n_n4958) & (n_n4953) & (!n_n4956) & (!n_n4957) & (n_n4961)) + ((!n_n4958) & (n_n4953) & (!n_n4956) & (n_n4957) & (!n_n4961)) + ((!n_n4958) & (n_n4953) & (!n_n4956) & (n_n4957) & (n_n4961)) + ((!n_n4958) & (n_n4953) & (n_n4956) & (!n_n4957) & (!n_n4961)) + ((!n_n4958) & (n_n4953) & (n_n4956) & (!n_n4957) & (n_n4961)) + ((!n_n4958) & (n_n4953) & (n_n4956) & (n_n4957) & (!n_n4961)) + ((!n_n4958) & (n_n4953) & (n_n4956) & (n_n4957) & (n_n4961)) + ((n_n4958) & (!n_n4953) & (!n_n4956) & (!n_n4957) & (!n_n4961)) + ((n_n4958) & (!n_n4953) & (!n_n4956) & (!n_n4957) & (n_n4961)) + ((n_n4958) & (!n_n4953) & (!n_n4956) & (n_n4957) & (!n_n4961)) + ((n_n4958) & (!n_n4953) & (!n_n4956) & (n_n4957) & (n_n4961)) + ((n_n4958) & (!n_n4953) & (n_n4956) & (!n_n4957) & (!n_n4961)) + ((n_n4958) & (!n_n4953) & (n_n4956) & (!n_n4957) & (n_n4961)) + ((n_n4958) & (!n_n4953) & (n_n4956) & (n_n4957) & (!n_n4961)) + ((n_n4958) & (!n_n4953) & (n_n4956) & (n_n4957) & (n_n4961)) + ((n_n4958) & (n_n4953) & (!n_n4956) & (!n_n4957) & (!n_n4961)) + ((n_n4958) & (n_n4953) & (!n_n4956) & (!n_n4957) & (n_n4961)) + ((n_n4958) & (n_n4953) & (!n_n4956) & (n_n4957) & (!n_n4961)) + ((n_n4958) & (n_n4953) & (!n_n4956) & (n_n4957) & (n_n4961)) + ((n_n4958) & (n_n4953) & (n_n4956) & (!n_n4957) & (!n_n4961)) + ((n_n4958) & (n_n4953) & (n_n4956) & (!n_n4957) & (n_n4961)) + ((n_n4958) & (n_n4953) & (n_n4956) & (n_n4957) & (!n_n4961)) + ((n_n4958) & (n_n4953) & (n_n4956) & (n_n4957) & (n_n4961)));
	assign x142x = (((!n_n3805) & (!n_n4949) & (!n_n4939) & (!n_n4944) & (x331x)) + ((!n_n3805) & (!n_n4949) & (!n_n4939) & (n_n4944) & (!x331x)) + ((!n_n3805) & (!n_n4949) & (!n_n4939) & (n_n4944) & (x331x)) + ((!n_n3805) & (!n_n4949) & (n_n4939) & (!n_n4944) & (!x331x)) + ((!n_n3805) & (!n_n4949) & (n_n4939) & (!n_n4944) & (x331x)) + ((!n_n3805) & (!n_n4949) & (n_n4939) & (n_n4944) & (!x331x)) + ((!n_n3805) & (!n_n4949) & (n_n4939) & (n_n4944) & (x331x)) + ((!n_n3805) & (n_n4949) & (!n_n4939) & (!n_n4944) & (!x331x)) + ((!n_n3805) & (n_n4949) & (!n_n4939) & (!n_n4944) & (x331x)) + ((!n_n3805) & (n_n4949) & (!n_n4939) & (n_n4944) & (!x331x)) + ((!n_n3805) & (n_n4949) & (!n_n4939) & (n_n4944) & (x331x)) + ((!n_n3805) & (n_n4949) & (n_n4939) & (!n_n4944) & (!x331x)) + ((!n_n3805) & (n_n4949) & (n_n4939) & (!n_n4944) & (x331x)) + ((!n_n3805) & (n_n4949) & (n_n4939) & (n_n4944) & (!x331x)) + ((!n_n3805) & (n_n4949) & (n_n4939) & (n_n4944) & (x331x)) + ((n_n3805) & (!n_n4949) & (!n_n4939) & (!n_n4944) & (!x331x)) + ((n_n3805) & (!n_n4949) & (!n_n4939) & (!n_n4944) & (x331x)) + ((n_n3805) & (!n_n4949) & (!n_n4939) & (n_n4944) & (!x331x)) + ((n_n3805) & (!n_n4949) & (!n_n4939) & (n_n4944) & (x331x)) + ((n_n3805) & (!n_n4949) & (n_n4939) & (!n_n4944) & (!x331x)) + ((n_n3805) & (!n_n4949) & (n_n4939) & (!n_n4944) & (x331x)) + ((n_n3805) & (!n_n4949) & (n_n4939) & (n_n4944) & (!x331x)) + ((n_n3805) & (!n_n4949) & (n_n4939) & (n_n4944) & (x331x)) + ((n_n3805) & (n_n4949) & (!n_n4939) & (!n_n4944) & (!x331x)) + ((n_n3805) & (n_n4949) & (!n_n4939) & (!n_n4944) & (x331x)) + ((n_n3805) & (n_n4949) & (!n_n4939) & (n_n4944) & (!x331x)) + ((n_n3805) & (n_n4949) & (!n_n4939) & (n_n4944) & (x331x)) + ((n_n3805) & (n_n4949) & (n_n4939) & (!n_n4944) & (!x331x)) + ((n_n3805) & (n_n4949) & (n_n4939) & (!n_n4944) & (x331x)) + ((n_n3805) & (n_n4949) & (n_n4939) & (n_n4944) & (!x331x)) + ((n_n3805) & (n_n4949) & (n_n4939) & (n_n4944) & (x331x)));
	assign x22148x = (((!x17x) & (!x516x) & (!n_n4926) & (!n_n4934) & (!n_n4936)) + ((!x17x) & (x516x) & (!n_n4926) & (!n_n4934) & (!n_n4936)) + ((x17x) & (!x516x) & (!n_n4926) & (!n_n4934) & (!n_n4936)));
	assign x12176x = (((!x31x) & (!n_n4933) & (!n_n4931) & (!x42x) & (!x22148x)) + ((!x31x) & (!n_n4933) & (!n_n4931) & (x42x) & (!x22148x)) + ((!x31x) & (!n_n4933) & (!n_n4931) & (x42x) & (x22148x)) + ((!x31x) & (!n_n4933) & (n_n4931) & (!x42x) & (!x22148x)) + ((!x31x) & (!n_n4933) & (n_n4931) & (!x42x) & (x22148x)) + ((!x31x) & (!n_n4933) & (n_n4931) & (x42x) & (!x22148x)) + ((!x31x) & (!n_n4933) & (n_n4931) & (x42x) & (x22148x)) + ((!x31x) & (n_n4933) & (!n_n4931) & (!x42x) & (!x22148x)) + ((!x31x) & (n_n4933) & (!n_n4931) & (!x42x) & (x22148x)) + ((!x31x) & (n_n4933) & (!n_n4931) & (x42x) & (!x22148x)) + ((!x31x) & (n_n4933) & (!n_n4931) & (x42x) & (x22148x)) + ((!x31x) & (n_n4933) & (n_n4931) & (!x42x) & (!x22148x)) + ((!x31x) & (n_n4933) & (n_n4931) & (!x42x) & (x22148x)) + ((!x31x) & (n_n4933) & (n_n4931) & (x42x) & (!x22148x)) + ((!x31x) & (n_n4933) & (n_n4931) & (x42x) & (x22148x)) + ((x31x) & (!n_n4933) & (!n_n4931) & (!x42x) & (!x22148x)) + ((x31x) & (!n_n4933) & (!n_n4931) & (!x42x) & (x22148x)) + ((x31x) & (!n_n4933) & (!n_n4931) & (x42x) & (!x22148x)) + ((x31x) & (!n_n4933) & (!n_n4931) & (x42x) & (x22148x)) + ((x31x) & (!n_n4933) & (n_n4931) & (!x42x) & (!x22148x)) + ((x31x) & (!n_n4933) & (n_n4931) & (!x42x) & (x22148x)) + ((x31x) & (!n_n4933) & (n_n4931) & (x42x) & (!x22148x)) + ((x31x) & (!n_n4933) & (n_n4931) & (x42x) & (x22148x)) + ((x31x) & (n_n4933) & (!n_n4931) & (!x42x) & (!x22148x)) + ((x31x) & (n_n4933) & (!n_n4931) & (!x42x) & (x22148x)) + ((x31x) & (n_n4933) & (!n_n4931) & (x42x) & (!x22148x)) + ((x31x) & (n_n4933) & (!n_n4931) & (x42x) & (x22148x)) + ((x31x) & (n_n4933) & (n_n4931) & (!x42x) & (!x22148x)) + ((x31x) & (n_n4933) & (n_n4931) & (!x42x) & (x22148x)) + ((x31x) & (n_n4933) & (n_n4931) & (x42x) & (!x22148x)) + ((x31x) & (n_n4933) & (n_n4931) & (x42x) & (x22148x)));
	assign n_n1463 = (((!n_n4888) & (!n_n4895) & (!x260x) & (!x48x) & (x49x)) + ((!n_n4888) & (!n_n4895) & (!x260x) & (x48x) & (!x49x)) + ((!n_n4888) & (!n_n4895) & (!x260x) & (x48x) & (x49x)) + ((!n_n4888) & (!n_n4895) & (x260x) & (!x48x) & (!x49x)) + ((!n_n4888) & (!n_n4895) & (x260x) & (!x48x) & (x49x)) + ((!n_n4888) & (!n_n4895) & (x260x) & (x48x) & (!x49x)) + ((!n_n4888) & (!n_n4895) & (x260x) & (x48x) & (x49x)) + ((!n_n4888) & (n_n4895) & (!x260x) & (!x48x) & (!x49x)) + ((!n_n4888) & (n_n4895) & (!x260x) & (!x48x) & (x49x)) + ((!n_n4888) & (n_n4895) & (!x260x) & (x48x) & (!x49x)) + ((!n_n4888) & (n_n4895) & (!x260x) & (x48x) & (x49x)) + ((!n_n4888) & (n_n4895) & (x260x) & (!x48x) & (!x49x)) + ((!n_n4888) & (n_n4895) & (x260x) & (!x48x) & (x49x)) + ((!n_n4888) & (n_n4895) & (x260x) & (x48x) & (!x49x)) + ((!n_n4888) & (n_n4895) & (x260x) & (x48x) & (x49x)) + ((n_n4888) & (!n_n4895) & (!x260x) & (!x48x) & (!x49x)) + ((n_n4888) & (!n_n4895) & (!x260x) & (!x48x) & (x49x)) + ((n_n4888) & (!n_n4895) & (!x260x) & (x48x) & (!x49x)) + ((n_n4888) & (!n_n4895) & (!x260x) & (x48x) & (x49x)) + ((n_n4888) & (!n_n4895) & (x260x) & (!x48x) & (!x49x)) + ((n_n4888) & (!n_n4895) & (x260x) & (!x48x) & (x49x)) + ((n_n4888) & (!n_n4895) & (x260x) & (x48x) & (!x49x)) + ((n_n4888) & (!n_n4895) & (x260x) & (x48x) & (x49x)) + ((n_n4888) & (n_n4895) & (!x260x) & (!x48x) & (!x49x)) + ((n_n4888) & (n_n4895) & (!x260x) & (!x48x) & (x49x)) + ((n_n4888) & (n_n4895) & (!x260x) & (x48x) & (!x49x)) + ((n_n4888) & (n_n4895) & (!x260x) & (x48x) & (x49x)) + ((n_n4888) & (n_n4895) & (x260x) & (!x48x) & (!x49x)) + ((n_n4888) & (n_n4895) & (x260x) & (!x48x) & (x49x)) + ((n_n4888) & (n_n4895) & (x260x) & (x48x) & (!x49x)) + ((n_n4888) & (n_n4895) & (x260x) & (x48x) & (x49x)));
	assign x305x = (((!i_9_) & (n_n482) & (n_n260) & (n_n530)) + ((i_9_) & (n_n482) & (n_n260) & (n_n530)));
	assign x12188x = (((!n_n4914) & (!n_n4917) & (!n_n4915) & (n_n4910)) + ((!n_n4914) & (!n_n4917) & (n_n4915) & (!n_n4910)) + ((!n_n4914) & (!n_n4917) & (n_n4915) & (n_n4910)) + ((!n_n4914) & (n_n4917) & (!n_n4915) & (!n_n4910)) + ((!n_n4914) & (n_n4917) & (!n_n4915) & (n_n4910)) + ((!n_n4914) & (n_n4917) & (n_n4915) & (!n_n4910)) + ((!n_n4914) & (n_n4917) & (n_n4915) & (n_n4910)) + ((n_n4914) & (!n_n4917) & (!n_n4915) & (!n_n4910)) + ((n_n4914) & (!n_n4917) & (!n_n4915) & (n_n4910)) + ((n_n4914) & (!n_n4917) & (n_n4915) & (!n_n4910)) + ((n_n4914) & (!n_n4917) & (n_n4915) & (n_n4910)) + ((n_n4914) & (n_n4917) & (!n_n4915) & (!n_n4910)) + ((n_n4914) & (n_n4917) & (!n_n4915) & (n_n4910)) + ((n_n4914) & (n_n4917) & (n_n4915) & (!n_n4910)) + ((n_n4914) & (n_n4917) & (n_n4915) & (n_n4910)));
	assign x12190x = (((!n_n4913) & (!x353x) & (!n_n4905) & (!x306x) & (x305x)) + ((!n_n4913) & (!x353x) & (!n_n4905) & (x306x) & (!x305x)) + ((!n_n4913) & (!x353x) & (!n_n4905) & (x306x) & (x305x)) + ((!n_n4913) & (!x353x) & (n_n4905) & (!x306x) & (!x305x)) + ((!n_n4913) & (!x353x) & (n_n4905) & (!x306x) & (x305x)) + ((!n_n4913) & (!x353x) & (n_n4905) & (x306x) & (!x305x)) + ((!n_n4913) & (!x353x) & (n_n4905) & (x306x) & (x305x)) + ((!n_n4913) & (x353x) & (!n_n4905) & (!x306x) & (!x305x)) + ((!n_n4913) & (x353x) & (!n_n4905) & (!x306x) & (x305x)) + ((!n_n4913) & (x353x) & (!n_n4905) & (x306x) & (!x305x)) + ((!n_n4913) & (x353x) & (!n_n4905) & (x306x) & (x305x)) + ((!n_n4913) & (x353x) & (n_n4905) & (!x306x) & (!x305x)) + ((!n_n4913) & (x353x) & (n_n4905) & (!x306x) & (x305x)) + ((!n_n4913) & (x353x) & (n_n4905) & (x306x) & (!x305x)) + ((!n_n4913) & (x353x) & (n_n4905) & (x306x) & (x305x)) + ((n_n4913) & (!x353x) & (!n_n4905) & (!x306x) & (!x305x)) + ((n_n4913) & (!x353x) & (!n_n4905) & (!x306x) & (x305x)) + ((n_n4913) & (!x353x) & (!n_n4905) & (x306x) & (!x305x)) + ((n_n4913) & (!x353x) & (!n_n4905) & (x306x) & (x305x)) + ((n_n4913) & (!x353x) & (n_n4905) & (!x306x) & (!x305x)) + ((n_n4913) & (!x353x) & (n_n4905) & (!x306x) & (x305x)) + ((n_n4913) & (!x353x) & (n_n4905) & (x306x) & (!x305x)) + ((n_n4913) & (!x353x) & (n_n4905) & (x306x) & (x305x)) + ((n_n4913) & (x353x) & (!n_n4905) & (!x306x) & (!x305x)) + ((n_n4913) & (x353x) & (!n_n4905) & (!x306x) & (x305x)) + ((n_n4913) & (x353x) & (!n_n4905) & (x306x) & (!x305x)) + ((n_n4913) & (x353x) & (!n_n4905) & (x306x) & (x305x)) + ((n_n4913) & (x353x) & (n_n4905) & (!x306x) & (!x305x)) + ((n_n4913) & (x353x) & (n_n4905) & (!x306x) & (x305x)) + ((n_n4913) & (x353x) & (n_n4905) & (x306x) & (!x305x)) + ((n_n4913) & (x353x) & (n_n4905) & (x306x) & (x305x)));
	assign x22166x = (((!n_n4460) & (!n_n4456) & (!n_n4458) & (!n_n4457)));
	assign x12662x = (((!n_n518) & (n_n526) & (!n_n532) & (n_n509) & (x18x)) + ((!n_n518) & (n_n526) & (n_n532) & (n_n509) & (x18x)) + ((n_n518) & (!n_n526) & (n_n532) & (!n_n509) & (x18x)) + ((n_n518) & (!n_n526) & (n_n532) & (n_n509) & (x18x)) + ((n_n518) & (n_n526) & (!n_n532) & (!n_n509) & (x18x)) + ((n_n518) & (n_n526) & (!n_n532) & (n_n509) & (x18x)) + ((n_n518) & (n_n526) & (n_n532) & (!n_n509) & (x18x)) + ((n_n518) & (n_n526) & (n_n532) & (n_n509) & (x18x)));
	assign x22135x = (((!n_n4987) & (!n_n5019) & (!n_n5010) & (!n_n4966)));
	assign n_n551 = (((!n_n5011) & (!n_n4961) & (!x12662x) & (!x22135x)) + ((!n_n5011) & (!n_n4961) & (x12662x) & (!x22135x)) + ((!n_n5011) & (!n_n4961) & (x12662x) & (x22135x)) + ((!n_n5011) & (n_n4961) & (!x12662x) & (!x22135x)) + ((!n_n5011) & (n_n4961) & (!x12662x) & (x22135x)) + ((!n_n5011) & (n_n4961) & (x12662x) & (!x22135x)) + ((!n_n5011) & (n_n4961) & (x12662x) & (x22135x)) + ((n_n5011) & (!n_n4961) & (!x12662x) & (!x22135x)) + ((n_n5011) & (!n_n4961) & (!x12662x) & (x22135x)) + ((n_n5011) & (!n_n4961) & (x12662x) & (!x22135x)) + ((n_n5011) & (!n_n4961) & (x12662x) & (x22135x)) + ((n_n5011) & (n_n4961) & (!x12662x) & (!x22135x)) + ((n_n5011) & (n_n4961) & (!x12662x) & (x22135x)) + ((n_n5011) & (n_n4961) & (x12662x) & (!x22135x)) + ((n_n5011) & (n_n4961) & (x12662x) & (x22135x)));
	assign x12670x = (((!x18x) & (!x572x) & (!n_n5042) & (!n_n5022) & (n_n5067)) + ((!x18x) & (!x572x) & (!n_n5042) & (n_n5022) & (!n_n5067)) + ((!x18x) & (!x572x) & (!n_n5042) & (n_n5022) & (n_n5067)) + ((!x18x) & (!x572x) & (n_n5042) & (!n_n5022) & (!n_n5067)) + ((!x18x) & (!x572x) & (n_n5042) & (!n_n5022) & (n_n5067)) + ((!x18x) & (!x572x) & (n_n5042) & (n_n5022) & (!n_n5067)) + ((!x18x) & (!x572x) & (n_n5042) & (n_n5022) & (n_n5067)) + ((!x18x) & (x572x) & (!n_n5042) & (!n_n5022) & (n_n5067)) + ((!x18x) & (x572x) & (!n_n5042) & (n_n5022) & (!n_n5067)) + ((!x18x) & (x572x) & (!n_n5042) & (n_n5022) & (n_n5067)) + ((!x18x) & (x572x) & (n_n5042) & (!n_n5022) & (!n_n5067)) + ((!x18x) & (x572x) & (n_n5042) & (!n_n5022) & (n_n5067)) + ((!x18x) & (x572x) & (n_n5042) & (n_n5022) & (!n_n5067)) + ((!x18x) & (x572x) & (n_n5042) & (n_n5022) & (n_n5067)) + ((x18x) & (!x572x) & (!n_n5042) & (!n_n5022) & (n_n5067)) + ((x18x) & (!x572x) & (!n_n5042) & (n_n5022) & (!n_n5067)) + ((x18x) & (!x572x) & (!n_n5042) & (n_n5022) & (n_n5067)) + ((x18x) & (!x572x) & (n_n5042) & (!n_n5022) & (!n_n5067)) + ((x18x) & (!x572x) & (n_n5042) & (!n_n5022) & (n_n5067)) + ((x18x) & (!x572x) & (n_n5042) & (n_n5022) & (!n_n5067)) + ((x18x) & (!x572x) & (n_n5042) & (n_n5022) & (n_n5067)) + ((x18x) & (x572x) & (!n_n5042) & (!n_n5022) & (!n_n5067)) + ((x18x) & (x572x) & (!n_n5042) & (!n_n5022) & (n_n5067)) + ((x18x) & (x572x) & (!n_n5042) & (n_n5022) & (!n_n5067)) + ((x18x) & (x572x) & (!n_n5042) & (n_n5022) & (n_n5067)) + ((x18x) & (x572x) & (n_n5042) & (!n_n5022) & (!n_n5067)) + ((x18x) & (x572x) & (n_n5042) & (!n_n5022) & (n_n5067)) + ((x18x) & (x572x) & (n_n5042) & (n_n5022) & (!n_n5067)) + ((x18x) & (x572x) & (n_n5042) & (n_n5022) & (n_n5067)));
	assign x12671x = (((!n_n526) & (!x18x) & (!n_n464) & (!n_n5075) & (x12669x)) + ((!n_n526) & (!x18x) & (!n_n464) & (n_n5075) & (!x12669x)) + ((!n_n526) & (!x18x) & (!n_n464) & (n_n5075) & (x12669x)) + ((!n_n526) & (!x18x) & (n_n464) & (!n_n5075) & (x12669x)) + ((!n_n526) & (!x18x) & (n_n464) & (n_n5075) & (!x12669x)) + ((!n_n526) & (!x18x) & (n_n464) & (n_n5075) & (x12669x)) + ((!n_n526) & (x18x) & (!n_n464) & (!n_n5075) & (x12669x)) + ((!n_n526) & (x18x) & (!n_n464) & (n_n5075) & (!x12669x)) + ((!n_n526) & (x18x) & (!n_n464) & (n_n5075) & (x12669x)) + ((!n_n526) & (x18x) & (n_n464) & (!n_n5075) & (x12669x)) + ((!n_n526) & (x18x) & (n_n464) & (n_n5075) & (!x12669x)) + ((!n_n526) & (x18x) & (n_n464) & (n_n5075) & (x12669x)) + ((n_n526) & (!x18x) & (!n_n464) & (!n_n5075) & (x12669x)) + ((n_n526) & (!x18x) & (!n_n464) & (n_n5075) & (!x12669x)) + ((n_n526) & (!x18x) & (!n_n464) & (n_n5075) & (x12669x)) + ((n_n526) & (!x18x) & (n_n464) & (!n_n5075) & (x12669x)) + ((n_n526) & (!x18x) & (n_n464) & (n_n5075) & (!x12669x)) + ((n_n526) & (!x18x) & (n_n464) & (n_n5075) & (x12669x)) + ((n_n526) & (x18x) & (!n_n464) & (!n_n5075) & (x12669x)) + ((n_n526) & (x18x) & (!n_n464) & (n_n5075) & (!x12669x)) + ((n_n526) & (x18x) & (!n_n464) & (n_n5075) & (x12669x)) + ((n_n526) & (x18x) & (n_n464) & (!n_n5075) & (!x12669x)) + ((n_n526) & (x18x) & (n_n464) & (!n_n5075) & (x12669x)) + ((n_n526) & (x18x) & (n_n464) & (n_n5075) & (!x12669x)) + ((n_n526) & (x18x) & (n_n464) & (n_n5075) & (x12669x)));
	assign x12679x = (((!n_n4890) & (!n_n4886) & (!n_n4872) & (!n_n4873) & (n_n4892)) + ((!n_n4890) & (!n_n4886) & (!n_n4872) & (n_n4873) & (!n_n4892)) + ((!n_n4890) & (!n_n4886) & (!n_n4872) & (n_n4873) & (n_n4892)) + ((!n_n4890) & (!n_n4886) & (n_n4872) & (!n_n4873) & (!n_n4892)) + ((!n_n4890) & (!n_n4886) & (n_n4872) & (!n_n4873) & (n_n4892)) + ((!n_n4890) & (!n_n4886) & (n_n4872) & (n_n4873) & (!n_n4892)) + ((!n_n4890) & (!n_n4886) & (n_n4872) & (n_n4873) & (n_n4892)) + ((!n_n4890) & (n_n4886) & (!n_n4872) & (!n_n4873) & (!n_n4892)) + ((!n_n4890) & (n_n4886) & (!n_n4872) & (!n_n4873) & (n_n4892)) + ((!n_n4890) & (n_n4886) & (!n_n4872) & (n_n4873) & (!n_n4892)) + ((!n_n4890) & (n_n4886) & (!n_n4872) & (n_n4873) & (n_n4892)) + ((!n_n4890) & (n_n4886) & (n_n4872) & (!n_n4873) & (!n_n4892)) + ((!n_n4890) & (n_n4886) & (n_n4872) & (!n_n4873) & (n_n4892)) + ((!n_n4890) & (n_n4886) & (n_n4872) & (n_n4873) & (!n_n4892)) + ((!n_n4890) & (n_n4886) & (n_n4872) & (n_n4873) & (n_n4892)) + ((n_n4890) & (!n_n4886) & (!n_n4872) & (!n_n4873) & (!n_n4892)) + ((n_n4890) & (!n_n4886) & (!n_n4872) & (!n_n4873) & (n_n4892)) + ((n_n4890) & (!n_n4886) & (!n_n4872) & (n_n4873) & (!n_n4892)) + ((n_n4890) & (!n_n4886) & (!n_n4872) & (n_n4873) & (n_n4892)) + ((n_n4890) & (!n_n4886) & (n_n4872) & (!n_n4873) & (!n_n4892)) + ((n_n4890) & (!n_n4886) & (n_n4872) & (!n_n4873) & (n_n4892)) + ((n_n4890) & (!n_n4886) & (n_n4872) & (n_n4873) & (!n_n4892)) + ((n_n4890) & (!n_n4886) & (n_n4872) & (n_n4873) & (n_n4892)) + ((n_n4890) & (n_n4886) & (!n_n4872) & (!n_n4873) & (!n_n4892)) + ((n_n4890) & (n_n4886) & (!n_n4872) & (!n_n4873) & (n_n4892)) + ((n_n4890) & (n_n4886) & (!n_n4872) & (n_n4873) & (!n_n4892)) + ((n_n4890) & (n_n4886) & (!n_n4872) & (n_n4873) & (n_n4892)) + ((n_n4890) & (n_n4886) & (n_n4872) & (!n_n4873) & (!n_n4892)) + ((n_n4890) & (n_n4886) & (n_n4872) & (!n_n4873) & (n_n4892)) + ((n_n4890) & (n_n4886) & (n_n4872) & (n_n4873) & (!n_n4892)) + ((n_n4890) & (n_n4886) & (n_n4872) & (n_n4873) & (n_n4892)));
	assign x22122x = (((!n_n4497) & (!n_n4499) & (!n_n4500) & (!n_n4496)));
	assign x13450x = (((!n_n4575) & (!n_n4584) & (!n_n4586) & (n_n4583)) + ((!n_n4575) & (!n_n4584) & (n_n4586) & (!n_n4583)) + ((!n_n4575) & (!n_n4584) & (n_n4586) & (n_n4583)) + ((!n_n4575) & (n_n4584) & (!n_n4586) & (!n_n4583)) + ((!n_n4575) & (n_n4584) & (!n_n4586) & (n_n4583)) + ((!n_n4575) & (n_n4584) & (n_n4586) & (!n_n4583)) + ((!n_n4575) & (n_n4584) & (n_n4586) & (n_n4583)) + ((n_n4575) & (!n_n4584) & (!n_n4586) & (!n_n4583)) + ((n_n4575) & (!n_n4584) & (!n_n4586) & (n_n4583)) + ((n_n4575) & (!n_n4584) & (n_n4586) & (!n_n4583)) + ((n_n4575) & (!n_n4584) & (n_n4586) & (n_n4583)) + ((n_n4575) & (n_n4584) & (!n_n4586) & (!n_n4583)) + ((n_n4575) & (n_n4584) & (!n_n4586) & (n_n4583)) + ((n_n4575) & (n_n4584) & (n_n4586) & (!n_n4583)) + ((n_n4575) & (n_n4584) & (n_n4586) & (n_n4583)));
	assign x13451x = (((!n_n390) & (!n_n535) & (!x20x) & (!n_n4577) & (x13449x)) + ((!n_n390) & (!n_n535) & (!x20x) & (n_n4577) & (!x13449x)) + ((!n_n390) & (!n_n535) & (!x20x) & (n_n4577) & (x13449x)) + ((!n_n390) & (!n_n535) & (x20x) & (!n_n4577) & (x13449x)) + ((!n_n390) & (!n_n535) & (x20x) & (n_n4577) & (!x13449x)) + ((!n_n390) & (!n_n535) & (x20x) & (n_n4577) & (x13449x)) + ((!n_n390) & (n_n535) & (!x20x) & (!n_n4577) & (x13449x)) + ((!n_n390) & (n_n535) & (!x20x) & (n_n4577) & (!x13449x)) + ((!n_n390) & (n_n535) & (!x20x) & (n_n4577) & (x13449x)) + ((!n_n390) & (n_n535) & (x20x) & (!n_n4577) & (x13449x)) + ((!n_n390) & (n_n535) & (x20x) & (n_n4577) & (!x13449x)) + ((!n_n390) & (n_n535) & (x20x) & (n_n4577) & (x13449x)) + ((n_n390) & (!n_n535) & (!x20x) & (!n_n4577) & (x13449x)) + ((n_n390) & (!n_n535) & (!x20x) & (n_n4577) & (!x13449x)) + ((n_n390) & (!n_n535) & (!x20x) & (n_n4577) & (x13449x)) + ((n_n390) & (!n_n535) & (x20x) & (!n_n4577) & (x13449x)) + ((n_n390) & (!n_n535) & (x20x) & (n_n4577) & (!x13449x)) + ((n_n390) & (!n_n535) & (x20x) & (n_n4577) & (x13449x)) + ((n_n390) & (n_n535) & (!x20x) & (!n_n4577) & (x13449x)) + ((n_n390) & (n_n535) & (!x20x) & (n_n4577) & (!x13449x)) + ((n_n390) & (n_n535) & (!x20x) & (n_n4577) & (x13449x)) + ((n_n390) & (n_n535) & (x20x) & (!n_n4577) & (!x13449x)) + ((n_n390) & (n_n535) & (x20x) & (!n_n4577) & (x13449x)) + ((n_n390) & (n_n535) & (x20x) & (n_n4577) & (!x13449x)) + ((n_n390) & (n_n535) & (x20x) & (n_n4577) & (x13449x)));
	assign x401x = (((!i_9_) & (n_n528) & (n_n390) & (n_n500)) + ((i_9_) & (n_n528) & (n_n390) & (n_n500)));
	assign x13464x = (((!n_n4625) & (!n_n4631) & (!n_n4635) & (n_n4620)) + ((!n_n4625) & (!n_n4631) & (n_n4635) & (!n_n4620)) + ((!n_n4625) & (!n_n4631) & (n_n4635) & (n_n4620)) + ((!n_n4625) & (n_n4631) & (!n_n4635) & (!n_n4620)) + ((!n_n4625) & (n_n4631) & (!n_n4635) & (n_n4620)) + ((!n_n4625) & (n_n4631) & (n_n4635) & (!n_n4620)) + ((!n_n4625) & (n_n4631) & (n_n4635) & (n_n4620)) + ((n_n4625) & (!n_n4631) & (!n_n4635) & (!n_n4620)) + ((n_n4625) & (!n_n4631) & (!n_n4635) & (n_n4620)) + ((n_n4625) & (!n_n4631) & (n_n4635) & (!n_n4620)) + ((n_n4625) & (!n_n4631) & (n_n4635) & (n_n4620)) + ((n_n4625) & (n_n4631) & (!n_n4635) & (!n_n4620)) + ((n_n4625) & (n_n4631) & (!n_n4635) & (n_n4620)) + ((n_n4625) & (n_n4631) & (n_n4635) & (!n_n4620)) + ((n_n4625) & (n_n4631) & (n_n4635) & (n_n4620)));
	assign x13466x = (((!n_n4634) & (!x118x) & (!n_n4638) & (!x357x) & (x401x)) + ((!n_n4634) & (!x118x) & (!n_n4638) & (x357x) & (!x401x)) + ((!n_n4634) & (!x118x) & (!n_n4638) & (x357x) & (x401x)) + ((!n_n4634) & (!x118x) & (n_n4638) & (!x357x) & (!x401x)) + ((!n_n4634) & (!x118x) & (n_n4638) & (!x357x) & (x401x)) + ((!n_n4634) & (!x118x) & (n_n4638) & (x357x) & (!x401x)) + ((!n_n4634) & (!x118x) & (n_n4638) & (x357x) & (x401x)) + ((!n_n4634) & (x118x) & (!n_n4638) & (!x357x) & (!x401x)) + ((!n_n4634) & (x118x) & (!n_n4638) & (!x357x) & (x401x)) + ((!n_n4634) & (x118x) & (!n_n4638) & (x357x) & (!x401x)) + ((!n_n4634) & (x118x) & (!n_n4638) & (x357x) & (x401x)) + ((!n_n4634) & (x118x) & (n_n4638) & (!x357x) & (!x401x)) + ((!n_n4634) & (x118x) & (n_n4638) & (!x357x) & (x401x)) + ((!n_n4634) & (x118x) & (n_n4638) & (x357x) & (!x401x)) + ((!n_n4634) & (x118x) & (n_n4638) & (x357x) & (x401x)) + ((n_n4634) & (!x118x) & (!n_n4638) & (!x357x) & (!x401x)) + ((n_n4634) & (!x118x) & (!n_n4638) & (!x357x) & (x401x)) + ((n_n4634) & (!x118x) & (!n_n4638) & (x357x) & (!x401x)) + ((n_n4634) & (!x118x) & (!n_n4638) & (x357x) & (x401x)) + ((n_n4634) & (!x118x) & (n_n4638) & (!x357x) & (!x401x)) + ((n_n4634) & (!x118x) & (n_n4638) & (!x357x) & (x401x)) + ((n_n4634) & (!x118x) & (n_n4638) & (x357x) & (!x401x)) + ((n_n4634) & (!x118x) & (n_n4638) & (x357x) & (x401x)) + ((n_n4634) & (x118x) & (!n_n4638) & (!x357x) & (!x401x)) + ((n_n4634) & (x118x) & (!n_n4638) & (!x357x) & (x401x)) + ((n_n4634) & (x118x) & (!n_n4638) & (x357x) & (!x401x)) + ((n_n4634) & (x118x) & (!n_n4638) & (x357x) & (x401x)) + ((n_n4634) & (x118x) & (n_n4638) & (!x357x) & (!x401x)) + ((n_n4634) & (x118x) & (n_n4638) & (!x357x) & (x401x)) + ((n_n4634) & (x118x) & (n_n4638) & (x357x) & (!x401x)) + ((n_n4634) & (x118x) & (n_n4638) & (x357x) & (x401x)));
	assign x22207x = (((!x13x) & (!x506x) & (!n_n4542) & (!n_n4548) & (!n_n4543)) + ((!x13x) & (x506x) & (!n_n4542) & (!n_n4548) & (!n_n4543)) + ((x13x) & (!x506x) & (!n_n4542) & (!n_n4548) & (!n_n4543)));
	assign x16390x = (((!x25x) & (!x483x) & (!n_n4724) & (!n_n4727) & (x101x)) + ((!x25x) & (!x483x) & (!n_n4724) & (n_n4727) & (!x101x)) + ((!x25x) & (!x483x) & (!n_n4724) & (n_n4727) & (x101x)) + ((!x25x) & (!x483x) & (n_n4724) & (!n_n4727) & (!x101x)) + ((!x25x) & (!x483x) & (n_n4724) & (!n_n4727) & (x101x)) + ((!x25x) & (!x483x) & (n_n4724) & (n_n4727) & (!x101x)) + ((!x25x) & (!x483x) & (n_n4724) & (n_n4727) & (x101x)) + ((!x25x) & (x483x) & (!n_n4724) & (!n_n4727) & (x101x)) + ((!x25x) & (x483x) & (!n_n4724) & (n_n4727) & (!x101x)) + ((!x25x) & (x483x) & (!n_n4724) & (n_n4727) & (x101x)) + ((!x25x) & (x483x) & (n_n4724) & (!n_n4727) & (!x101x)) + ((!x25x) & (x483x) & (n_n4724) & (!n_n4727) & (x101x)) + ((!x25x) & (x483x) & (n_n4724) & (n_n4727) & (!x101x)) + ((!x25x) & (x483x) & (n_n4724) & (n_n4727) & (x101x)) + ((x25x) & (!x483x) & (!n_n4724) & (!n_n4727) & (x101x)) + ((x25x) & (!x483x) & (!n_n4724) & (n_n4727) & (!x101x)) + ((x25x) & (!x483x) & (!n_n4724) & (n_n4727) & (x101x)) + ((x25x) & (!x483x) & (n_n4724) & (!n_n4727) & (!x101x)) + ((x25x) & (!x483x) & (n_n4724) & (!n_n4727) & (x101x)) + ((x25x) & (!x483x) & (n_n4724) & (n_n4727) & (!x101x)) + ((x25x) & (!x483x) & (n_n4724) & (n_n4727) & (x101x)) + ((x25x) & (x483x) & (!n_n4724) & (!n_n4727) & (!x101x)) + ((x25x) & (x483x) & (!n_n4724) & (!n_n4727) & (x101x)) + ((x25x) & (x483x) & (!n_n4724) & (n_n4727) & (!x101x)) + ((x25x) & (x483x) & (!n_n4724) & (n_n4727) & (x101x)) + ((x25x) & (x483x) & (n_n4724) & (!n_n4727) & (!x101x)) + ((x25x) & (x483x) & (n_n4724) & (!n_n4727) & (x101x)) + ((x25x) & (x483x) & (n_n4724) & (n_n4727) & (!x101x)) + ((x25x) & (x483x) & (n_n4724) & (n_n4727) & (x101x)));
	assign x12492x = (((!i_9_) & (n_n455) & (!n_n532) & (n_n509) & (n_n530)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n509) & (!n_n530)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n509) & (n_n530)) + ((i_9_) & (n_n455) & (!n_n532) & (n_n509) & (n_n530)) + ((i_9_) & (n_n455) & (n_n532) & (n_n509) & (n_n530)));
	assign n_n1496 = (((!n_n4471) & (!n_n4472) & (!x194x) & (!x199x) & (x12492x)) + ((!n_n4471) & (!n_n4472) & (!x194x) & (x199x) & (!x12492x)) + ((!n_n4471) & (!n_n4472) & (!x194x) & (x199x) & (x12492x)) + ((!n_n4471) & (!n_n4472) & (x194x) & (!x199x) & (!x12492x)) + ((!n_n4471) & (!n_n4472) & (x194x) & (!x199x) & (x12492x)) + ((!n_n4471) & (!n_n4472) & (x194x) & (x199x) & (!x12492x)) + ((!n_n4471) & (!n_n4472) & (x194x) & (x199x) & (x12492x)) + ((!n_n4471) & (n_n4472) & (!x194x) & (!x199x) & (!x12492x)) + ((!n_n4471) & (n_n4472) & (!x194x) & (!x199x) & (x12492x)) + ((!n_n4471) & (n_n4472) & (!x194x) & (x199x) & (!x12492x)) + ((!n_n4471) & (n_n4472) & (!x194x) & (x199x) & (x12492x)) + ((!n_n4471) & (n_n4472) & (x194x) & (!x199x) & (!x12492x)) + ((!n_n4471) & (n_n4472) & (x194x) & (!x199x) & (x12492x)) + ((!n_n4471) & (n_n4472) & (x194x) & (x199x) & (!x12492x)) + ((!n_n4471) & (n_n4472) & (x194x) & (x199x) & (x12492x)) + ((n_n4471) & (!n_n4472) & (!x194x) & (!x199x) & (!x12492x)) + ((n_n4471) & (!n_n4472) & (!x194x) & (!x199x) & (x12492x)) + ((n_n4471) & (!n_n4472) & (!x194x) & (x199x) & (!x12492x)) + ((n_n4471) & (!n_n4472) & (!x194x) & (x199x) & (x12492x)) + ((n_n4471) & (!n_n4472) & (x194x) & (!x199x) & (!x12492x)) + ((n_n4471) & (!n_n4472) & (x194x) & (!x199x) & (x12492x)) + ((n_n4471) & (!n_n4472) & (x194x) & (x199x) & (!x12492x)) + ((n_n4471) & (!n_n4472) & (x194x) & (x199x) & (x12492x)) + ((n_n4471) & (n_n4472) & (!x194x) & (!x199x) & (!x12492x)) + ((n_n4471) & (n_n4472) & (!x194x) & (!x199x) & (x12492x)) + ((n_n4471) & (n_n4472) & (!x194x) & (x199x) & (!x12492x)) + ((n_n4471) & (n_n4472) & (!x194x) & (x199x) & (x12492x)) + ((n_n4471) & (n_n4472) & (x194x) & (!x199x) & (!x12492x)) + ((n_n4471) & (n_n4472) & (x194x) & (!x199x) & (x12492x)) + ((n_n4471) & (n_n4472) & (x194x) & (x199x) & (!x12492x)) + ((n_n4471) & (n_n4472) & (x194x) & (x199x) & (x12492x)));
	assign x12231x = (((!x15x) & (!x552x) & (!n_n4838) & (!n_n4833) & (x304x)) + ((!x15x) & (!x552x) & (!n_n4838) & (n_n4833) & (!x304x)) + ((!x15x) & (!x552x) & (!n_n4838) & (n_n4833) & (x304x)) + ((!x15x) & (!x552x) & (n_n4838) & (!n_n4833) & (!x304x)) + ((!x15x) & (!x552x) & (n_n4838) & (!n_n4833) & (x304x)) + ((!x15x) & (!x552x) & (n_n4838) & (n_n4833) & (!x304x)) + ((!x15x) & (!x552x) & (n_n4838) & (n_n4833) & (x304x)) + ((!x15x) & (x552x) & (!n_n4838) & (!n_n4833) & (x304x)) + ((!x15x) & (x552x) & (!n_n4838) & (n_n4833) & (!x304x)) + ((!x15x) & (x552x) & (!n_n4838) & (n_n4833) & (x304x)) + ((!x15x) & (x552x) & (n_n4838) & (!n_n4833) & (!x304x)) + ((!x15x) & (x552x) & (n_n4838) & (!n_n4833) & (x304x)) + ((!x15x) & (x552x) & (n_n4838) & (n_n4833) & (!x304x)) + ((!x15x) & (x552x) & (n_n4838) & (n_n4833) & (x304x)) + ((x15x) & (!x552x) & (!n_n4838) & (!n_n4833) & (x304x)) + ((x15x) & (!x552x) & (!n_n4838) & (n_n4833) & (!x304x)) + ((x15x) & (!x552x) & (!n_n4838) & (n_n4833) & (x304x)) + ((x15x) & (!x552x) & (n_n4838) & (!n_n4833) & (!x304x)) + ((x15x) & (!x552x) & (n_n4838) & (!n_n4833) & (x304x)) + ((x15x) & (!x552x) & (n_n4838) & (n_n4833) & (!x304x)) + ((x15x) & (!x552x) & (n_n4838) & (n_n4833) & (x304x)) + ((x15x) & (x552x) & (!n_n4838) & (!n_n4833) & (!x304x)) + ((x15x) & (x552x) & (!n_n4838) & (!n_n4833) & (x304x)) + ((x15x) & (x552x) & (!n_n4838) & (n_n4833) & (!x304x)) + ((x15x) & (x552x) & (!n_n4838) & (n_n4833) & (x304x)) + ((x15x) & (x552x) & (n_n4838) & (!n_n4833) & (!x304x)) + ((x15x) & (x552x) & (n_n4838) & (!n_n4833) & (x304x)) + ((x15x) & (x552x) & (n_n4838) & (n_n4833) & (!x304x)) + ((x15x) & (x552x) & (n_n4838) & (n_n4833) & (x304x)));
	assign n_n1468 = (((!n_n4830) & (!n_n4831) & (!n_n4827) & (!n_n4828) & (x12231x)) + ((!n_n4830) & (!n_n4831) & (!n_n4827) & (n_n4828) & (!x12231x)) + ((!n_n4830) & (!n_n4831) & (!n_n4827) & (n_n4828) & (x12231x)) + ((!n_n4830) & (!n_n4831) & (n_n4827) & (!n_n4828) & (!x12231x)) + ((!n_n4830) & (!n_n4831) & (n_n4827) & (!n_n4828) & (x12231x)) + ((!n_n4830) & (!n_n4831) & (n_n4827) & (n_n4828) & (!x12231x)) + ((!n_n4830) & (!n_n4831) & (n_n4827) & (n_n4828) & (x12231x)) + ((!n_n4830) & (n_n4831) & (!n_n4827) & (!n_n4828) & (!x12231x)) + ((!n_n4830) & (n_n4831) & (!n_n4827) & (!n_n4828) & (x12231x)) + ((!n_n4830) & (n_n4831) & (!n_n4827) & (n_n4828) & (!x12231x)) + ((!n_n4830) & (n_n4831) & (!n_n4827) & (n_n4828) & (x12231x)) + ((!n_n4830) & (n_n4831) & (n_n4827) & (!n_n4828) & (!x12231x)) + ((!n_n4830) & (n_n4831) & (n_n4827) & (!n_n4828) & (x12231x)) + ((!n_n4830) & (n_n4831) & (n_n4827) & (n_n4828) & (!x12231x)) + ((!n_n4830) & (n_n4831) & (n_n4827) & (n_n4828) & (x12231x)) + ((n_n4830) & (!n_n4831) & (!n_n4827) & (!n_n4828) & (!x12231x)) + ((n_n4830) & (!n_n4831) & (!n_n4827) & (!n_n4828) & (x12231x)) + ((n_n4830) & (!n_n4831) & (!n_n4827) & (n_n4828) & (!x12231x)) + ((n_n4830) & (!n_n4831) & (!n_n4827) & (n_n4828) & (x12231x)) + ((n_n4830) & (!n_n4831) & (n_n4827) & (!n_n4828) & (!x12231x)) + ((n_n4830) & (!n_n4831) & (n_n4827) & (!n_n4828) & (x12231x)) + ((n_n4830) & (!n_n4831) & (n_n4827) & (n_n4828) & (!x12231x)) + ((n_n4830) & (!n_n4831) & (n_n4827) & (n_n4828) & (x12231x)) + ((n_n4830) & (n_n4831) & (!n_n4827) & (!n_n4828) & (!x12231x)) + ((n_n4830) & (n_n4831) & (!n_n4827) & (!n_n4828) & (x12231x)) + ((n_n4830) & (n_n4831) & (!n_n4827) & (n_n4828) & (!x12231x)) + ((n_n4830) & (n_n4831) & (!n_n4827) & (n_n4828) & (x12231x)) + ((n_n4830) & (n_n4831) & (n_n4827) & (!n_n4828) & (!x12231x)) + ((n_n4830) & (n_n4831) & (n_n4827) & (!n_n4828) & (x12231x)) + ((n_n4830) & (n_n4831) & (n_n4827) & (n_n4828) & (!x12231x)) + ((n_n4830) & (n_n4831) & (n_n4827) & (n_n4828) & (x12231x)));
	assign x12235x = (((!n_n4849) & (!n_n4847) & (!n_n4843) & (n_n4846)) + ((!n_n4849) & (!n_n4847) & (n_n4843) & (!n_n4846)) + ((!n_n4849) & (!n_n4847) & (n_n4843) & (n_n4846)) + ((!n_n4849) & (n_n4847) & (!n_n4843) & (!n_n4846)) + ((!n_n4849) & (n_n4847) & (!n_n4843) & (n_n4846)) + ((!n_n4849) & (n_n4847) & (n_n4843) & (!n_n4846)) + ((!n_n4849) & (n_n4847) & (n_n4843) & (n_n4846)) + ((n_n4849) & (!n_n4847) & (!n_n4843) & (!n_n4846)) + ((n_n4849) & (!n_n4847) & (!n_n4843) & (n_n4846)) + ((n_n4849) & (!n_n4847) & (n_n4843) & (!n_n4846)) + ((n_n4849) & (!n_n4847) & (n_n4843) & (n_n4846)) + ((n_n4849) & (n_n4847) & (!n_n4843) & (!n_n4846)) + ((n_n4849) & (n_n4847) & (!n_n4843) & (n_n4846)) + ((n_n4849) & (n_n4847) & (n_n4843) & (!n_n4846)) + ((n_n4849) & (n_n4847) & (n_n4843) & (n_n4846)));
	assign x12236x = (((!x552x) & (!x23x) & (!n_n4848) & (!x372x) & (n_n4851)) + ((!x552x) & (!x23x) & (!n_n4848) & (x372x) & (!n_n4851)) + ((!x552x) & (!x23x) & (!n_n4848) & (x372x) & (n_n4851)) + ((!x552x) & (!x23x) & (n_n4848) & (!x372x) & (!n_n4851)) + ((!x552x) & (!x23x) & (n_n4848) & (!x372x) & (n_n4851)) + ((!x552x) & (!x23x) & (n_n4848) & (x372x) & (!n_n4851)) + ((!x552x) & (!x23x) & (n_n4848) & (x372x) & (n_n4851)) + ((!x552x) & (x23x) & (!n_n4848) & (!x372x) & (n_n4851)) + ((!x552x) & (x23x) & (!n_n4848) & (x372x) & (!n_n4851)) + ((!x552x) & (x23x) & (!n_n4848) & (x372x) & (n_n4851)) + ((!x552x) & (x23x) & (n_n4848) & (!x372x) & (!n_n4851)) + ((!x552x) & (x23x) & (n_n4848) & (!x372x) & (n_n4851)) + ((!x552x) & (x23x) & (n_n4848) & (x372x) & (!n_n4851)) + ((!x552x) & (x23x) & (n_n4848) & (x372x) & (n_n4851)) + ((x552x) & (!x23x) & (!n_n4848) & (!x372x) & (n_n4851)) + ((x552x) & (!x23x) & (!n_n4848) & (x372x) & (!n_n4851)) + ((x552x) & (!x23x) & (!n_n4848) & (x372x) & (n_n4851)) + ((x552x) & (!x23x) & (n_n4848) & (!x372x) & (!n_n4851)) + ((x552x) & (!x23x) & (n_n4848) & (!x372x) & (n_n4851)) + ((x552x) & (!x23x) & (n_n4848) & (x372x) & (!n_n4851)) + ((x552x) & (!x23x) & (n_n4848) & (x372x) & (n_n4851)) + ((x552x) & (x23x) & (!n_n4848) & (!x372x) & (!n_n4851)) + ((x552x) & (x23x) & (!n_n4848) & (!x372x) & (n_n4851)) + ((x552x) & (x23x) & (!n_n4848) & (x372x) & (!n_n4851)) + ((x552x) & (x23x) & (!n_n4848) & (x372x) & (n_n4851)) + ((x552x) & (x23x) & (n_n4848) & (!x372x) & (!n_n4851)) + ((x552x) & (x23x) & (n_n4848) & (!x372x) & (n_n4851)) + ((x552x) & (x23x) & (n_n4848) & (x372x) & (!n_n4851)) + ((x552x) & (x23x) & (n_n4848) & (x372x) & (n_n4851)));
	assign x12240x = (((!n_n4817) & (!n_n4824) & (!x185x) & (!x186x) & (n_n4196)) + ((!n_n4817) & (!n_n4824) & (!x185x) & (x186x) & (!n_n4196)) + ((!n_n4817) & (!n_n4824) & (!x185x) & (x186x) & (n_n4196)) + ((!n_n4817) & (!n_n4824) & (x185x) & (!x186x) & (!n_n4196)) + ((!n_n4817) & (!n_n4824) & (x185x) & (!x186x) & (n_n4196)) + ((!n_n4817) & (!n_n4824) & (x185x) & (x186x) & (!n_n4196)) + ((!n_n4817) & (!n_n4824) & (x185x) & (x186x) & (n_n4196)) + ((!n_n4817) & (n_n4824) & (!x185x) & (!x186x) & (!n_n4196)) + ((!n_n4817) & (n_n4824) & (!x185x) & (!x186x) & (n_n4196)) + ((!n_n4817) & (n_n4824) & (!x185x) & (x186x) & (!n_n4196)) + ((!n_n4817) & (n_n4824) & (!x185x) & (x186x) & (n_n4196)) + ((!n_n4817) & (n_n4824) & (x185x) & (!x186x) & (!n_n4196)) + ((!n_n4817) & (n_n4824) & (x185x) & (!x186x) & (n_n4196)) + ((!n_n4817) & (n_n4824) & (x185x) & (x186x) & (!n_n4196)) + ((!n_n4817) & (n_n4824) & (x185x) & (x186x) & (n_n4196)) + ((n_n4817) & (!n_n4824) & (!x185x) & (!x186x) & (!n_n4196)) + ((n_n4817) & (!n_n4824) & (!x185x) & (!x186x) & (n_n4196)) + ((n_n4817) & (!n_n4824) & (!x185x) & (x186x) & (!n_n4196)) + ((n_n4817) & (!n_n4824) & (!x185x) & (x186x) & (n_n4196)) + ((n_n4817) & (!n_n4824) & (x185x) & (!x186x) & (!n_n4196)) + ((n_n4817) & (!n_n4824) & (x185x) & (!x186x) & (n_n4196)) + ((n_n4817) & (!n_n4824) & (x185x) & (x186x) & (!n_n4196)) + ((n_n4817) & (!n_n4824) & (x185x) & (x186x) & (n_n4196)) + ((n_n4817) & (n_n4824) & (!x185x) & (!x186x) & (!n_n4196)) + ((n_n4817) & (n_n4824) & (!x185x) & (!x186x) & (n_n4196)) + ((n_n4817) & (n_n4824) & (!x185x) & (x186x) & (!n_n4196)) + ((n_n4817) & (n_n4824) & (!x185x) & (x186x) & (n_n4196)) + ((n_n4817) & (n_n4824) & (x185x) & (!x186x) & (!n_n4196)) + ((n_n4817) & (n_n4824) & (x185x) & (!x186x) & (n_n4196)) + ((n_n4817) & (n_n4824) & (x185x) & (x186x) & (!n_n4196)) + ((n_n4817) & (n_n4824) & (x185x) & (x186x) & (n_n4196)));
	assign x11867x = (((!n_n4711) & (!n_n4712) & (!n_n4715) & (n_n4714)) + ((!n_n4711) & (!n_n4712) & (n_n4715) & (!n_n4714)) + ((!n_n4711) & (!n_n4712) & (n_n4715) & (n_n4714)) + ((!n_n4711) & (n_n4712) & (!n_n4715) & (!n_n4714)) + ((!n_n4711) & (n_n4712) & (!n_n4715) & (n_n4714)) + ((!n_n4711) & (n_n4712) & (n_n4715) & (!n_n4714)) + ((!n_n4711) & (n_n4712) & (n_n4715) & (n_n4714)) + ((n_n4711) & (!n_n4712) & (!n_n4715) & (!n_n4714)) + ((n_n4711) & (!n_n4712) & (!n_n4715) & (n_n4714)) + ((n_n4711) & (!n_n4712) & (n_n4715) & (!n_n4714)) + ((n_n4711) & (!n_n4712) & (n_n4715) & (n_n4714)) + ((n_n4711) & (n_n4712) & (!n_n4715) & (!n_n4714)) + ((n_n4711) & (n_n4712) & (!n_n4715) & (n_n4714)) + ((n_n4711) & (n_n4712) & (n_n4715) & (!n_n4714)) + ((n_n4711) & (n_n4712) & (n_n4715) & (n_n4714)));
	assign x11868x = (((!x241x) & (!n_n4710) & (!n_n4719) & (n_n4716)) + ((!x241x) & (!n_n4710) & (n_n4719) & (!n_n4716)) + ((!x241x) & (!n_n4710) & (n_n4719) & (n_n4716)) + ((!x241x) & (n_n4710) & (!n_n4719) & (!n_n4716)) + ((!x241x) & (n_n4710) & (!n_n4719) & (n_n4716)) + ((!x241x) & (n_n4710) & (n_n4719) & (!n_n4716)) + ((!x241x) & (n_n4710) & (n_n4719) & (n_n4716)) + ((x241x) & (!n_n4710) & (!n_n4719) & (!n_n4716)) + ((x241x) & (!n_n4710) & (!n_n4719) & (n_n4716)) + ((x241x) & (!n_n4710) & (n_n4719) & (!n_n4716)) + ((x241x) & (!n_n4710) & (n_n4719) & (n_n4716)) + ((x241x) & (n_n4710) & (!n_n4719) & (!n_n4716)) + ((x241x) & (n_n4710) & (!n_n4719) & (n_n4716)) + ((x241x) & (n_n4710) & (n_n4719) & (!n_n4716)) + ((x241x) & (n_n4710) & (n_n4719) & (n_n4716)));
	assign x124x = (((!i_9_) & (n_n536) & (n_n518) & (!n_n522) & (x20x)) + ((!i_9_) & (n_n536) & (n_n518) & (n_n522) & (x20x)) + ((i_9_) & (n_n536) & (n_n518) & (!n_n522) & (x20x)) + ((i_9_) & (n_n536) & (n_n518) & (n_n522) & (!x20x)) + ((i_9_) & (n_n536) & (n_n518) & (n_n522) & (x20x)));
	assign x22089x = (((!n_n4344) & (!n_n4342) & (!n_n4352) & (!n_n4349)));
	assign n_n3010 = (((!n_n4340) & (!n_n4341) & (!x67x) & (!n_n4350) & (!x22089x)) + ((!n_n4340) & (!n_n4341) & (!x67x) & (n_n4350) & (!x22089x)) + ((!n_n4340) & (!n_n4341) & (!x67x) & (n_n4350) & (x22089x)) + ((!n_n4340) & (!n_n4341) & (x67x) & (!n_n4350) & (!x22089x)) + ((!n_n4340) & (!n_n4341) & (x67x) & (!n_n4350) & (x22089x)) + ((!n_n4340) & (!n_n4341) & (x67x) & (n_n4350) & (!x22089x)) + ((!n_n4340) & (!n_n4341) & (x67x) & (n_n4350) & (x22089x)) + ((!n_n4340) & (n_n4341) & (!x67x) & (!n_n4350) & (!x22089x)) + ((!n_n4340) & (n_n4341) & (!x67x) & (!n_n4350) & (x22089x)) + ((!n_n4340) & (n_n4341) & (!x67x) & (n_n4350) & (!x22089x)) + ((!n_n4340) & (n_n4341) & (!x67x) & (n_n4350) & (x22089x)) + ((!n_n4340) & (n_n4341) & (x67x) & (!n_n4350) & (!x22089x)) + ((!n_n4340) & (n_n4341) & (x67x) & (!n_n4350) & (x22089x)) + ((!n_n4340) & (n_n4341) & (x67x) & (n_n4350) & (!x22089x)) + ((!n_n4340) & (n_n4341) & (x67x) & (n_n4350) & (x22089x)) + ((n_n4340) & (!n_n4341) & (!x67x) & (!n_n4350) & (!x22089x)) + ((n_n4340) & (!n_n4341) & (!x67x) & (!n_n4350) & (x22089x)) + ((n_n4340) & (!n_n4341) & (!x67x) & (n_n4350) & (!x22089x)) + ((n_n4340) & (!n_n4341) & (!x67x) & (n_n4350) & (x22089x)) + ((n_n4340) & (!n_n4341) & (x67x) & (!n_n4350) & (!x22089x)) + ((n_n4340) & (!n_n4341) & (x67x) & (!n_n4350) & (x22089x)) + ((n_n4340) & (!n_n4341) & (x67x) & (n_n4350) & (!x22089x)) + ((n_n4340) & (!n_n4341) & (x67x) & (n_n4350) & (x22089x)) + ((n_n4340) & (n_n4341) & (!x67x) & (!n_n4350) & (!x22089x)) + ((n_n4340) & (n_n4341) & (!x67x) & (!n_n4350) & (x22089x)) + ((n_n4340) & (n_n4341) & (!x67x) & (n_n4350) & (!x22089x)) + ((n_n4340) & (n_n4341) & (!x67x) & (n_n4350) & (x22089x)) + ((n_n4340) & (n_n4341) & (x67x) & (!n_n4350) & (!x22089x)) + ((n_n4340) & (n_n4341) & (x67x) & (!n_n4350) & (x22089x)) + ((n_n4340) & (n_n4341) & (x67x) & (n_n4350) & (!x22089x)) + ((n_n4340) & (n_n4341) & (x67x) & (n_n4350) & (x22089x)));
	assign x22097x = (((!n_n4602) & (!n_n4601) & (!n_n4607) & (!n_n4600)));
	assign x51x = (((!n_n390) & (!n_n509) & (!x20x) & (!x23x) & (n_n4614)) + ((!n_n390) & (!n_n509) & (!x20x) & (x23x) & (n_n4614)) + ((!n_n390) & (!n_n509) & (x20x) & (!x23x) & (n_n4614)) + ((!n_n390) & (!n_n509) & (x20x) & (x23x) & (n_n4614)) + ((!n_n390) & (n_n509) & (!x20x) & (!x23x) & (n_n4614)) + ((!n_n390) & (n_n509) & (!x20x) & (x23x) & (n_n4614)) + ((!n_n390) & (n_n509) & (x20x) & (!x23x) & (n_n4614)) + ((!n_n390) & (n_n509) & (x20x) & (x23x) & (n_n4614)) + ((n_n390) & (!n_n509) & (!x20x) & (!x23x) & (n_n4614)) + ((n_n390) & (!n_n509) & (!x20x) & (x23x) & (n_n4614)) + ((n_n390) & (!n_n509) & (x20x) & (!x23x) & (n_n4614)) + ((n_n390) & (!n_n509) & (x20x) & (x23x) & (n_n4614)) + ((n_n390) & (n_n509) & (!x20x) & (!x23x) & (n_n4614)) + ((n_n390) & (n_n509) & (!x20x) & (x23x) & (!n_n4614)) + ((n_n390) & (n_n509) & (!x20x) & (x23x) & (n_n4614)) + ((n_n390) & (n_n509) & (x20x) & (!x23x) & (!n_n4614)) + ((n_n390) & (n_n509) & (x20x) & (!x23x) & (n_n4614)) + ((n_n390) & (n_n509) & (x20x) & (x23x) & (!n_n4614)) + ((n_n390) & (n_n509) & (x20x) & (x23x) & (n_n4614)));
	assign x22167x = (((!n_n4612) & (!n_n4611) & (!n_n4622) & (!n_n4620)));
	assign x12504x = (((!n_n4536) & (!n_n4537) & (!n_n4528) & (n_n4534)) + ((!n_n4536) & (!n_n4537) & (n_n4528) & (!n_n4534)) + ((!n_n4536) & (!n_n4537) & (n_n4528) & (n_n4534)) + ((!n_n4536) & (n_n4537) & (!n_n4528) & (!n_n4534)) + ((!n_n4536) & (n_n4537) & (!n_n4528) & (n_n4534)) + ((!n_n4536) & (n_n4537) & (n_n4528) & (!n_n4534)) + ((!n_n4536) & (n_n4537) & (n_n4528) & (n_n4534)) + ((n_n4536) & (!n_n4537) & (!n_n4528) & (!n_n4534)) + ((n_n4536) & (!n_n4537) & (!n_n4528) & (n_n4534)) + ((n_n4536) & (!n_n4537) & (n_n4528) & (!n_n4534)) + ((n_n4536) & (!n_n4537) & (n_n4528) & (n_n4534)) + ((n_n4536) & (n_n4537) & (!n_n4528) & (!n_n4534)) + ((n_n4536) & (n_n4537) & (!n_n4528) & (n_n4534)) + ((n_n4536) & (n_n4537) & (n_n4528) & (!n_n4534)) + ((n_n4536) & (n_n4537) & (n_n4528) & (n_n4534)));
	assign x12505x = (((!x13x) & (!n_n491) & (!n_n520) & (!n_n4247) & (x307x)) + ((!x13x) & (!n_n491) & (!n_n520) & (n_n4247) & (!x307x)) + ((!x13x) & (!n_n491) & (!n_n520) & (n_n4247) & (x307x)) + ((!x13x) & (!n_n491) & (n_n520) & (!n_n4247) & (x307x)) + ((!x13x) & (!n_n491) & (n_n520) & (n_n4247) & (!x307x)) + ((!x13x) & (!n_n491) & (n_n520) & (n_n4247) & (x307x)) + ((!x13x) & (n_n491) & (!n_n520) & (!n_n4247) & (x307x)) + ((!x13x) & (n_n491) & (!n_n520) & (n_n4247) & (!x307x)) + ((!x13x) & (n_n491) & (!n_n520) & (n_n4247) & (x307x)) + ((!x13x) & (n_n491) & (n_n520) & (!n_n4247) & (x307x)) + ((!x13x) & (n_n491) & (n_n520) & (n_n4247) & (!x307x)) + ((!x13x) & (n_n491) & (n_n520) & (n_n4247) & (x307x)) + ((x13x) & (!n_n491) & (!n_n520) & (!n_n4247) & (x307x)) + ((x13x) & (!n_n491) & (!n_n520) & (n_n4247) & (!x307x)) + ((x13x) & (!n_n491) & (!n_n520) & (n_n4247) & (x307x)) + ((x13x) & (!n_n491) & (n_n520) & (!n_n4247) & (x307x)) + ((x13x) & (!n_n491) & (n_n520) & (n_n4247) & (!x307x)) + ((x13x) & (!n_n491) & (n_n520) & (n_n4247) & (x307x)) + ((x13x) & (n_n491) & (!n_n520) & (!n_n4247) & (x307x)) + ((x13x) & (n_n491) & (!n_n520) & (n_n4247) & (!x307x)) + ((x13x) & (n_n491) & (!n_n520) & (n_n4247) & (x307x)) + ((x13x) & (n_n491) & (n_n520) & (!n_n4247) & (!x307x)) + ((x13x) & (n_n491) & (n_n520) & (!n_n4247) & (x307x)) + ((x13x) & (n_n491) & (n_n520) & (n_n4247) & (!x307x)) + ((x13x) & (n_n491) & (n_n520) & (n_n4247) & (x307x)));
	assign x12506x = (((!n_n4521) & (!x170x) & (!n_n4531) & (!x178x) & (x361x)) + ((!n_n4521) & (!x170x) & (!n_n4531) & (x178x) & (!x361x)) + ((!n_n4521) & (!x170x) & (!n_n4531) & (x178x) & (x361x)) + ((!n_n4521) & (!x170x) & (n_n4531) & (!x178x) & (!x361x)) + ((!n_n4521) & (!x170x) & (n_n4531) & (!x178x) & (x361x)) + ((!n_n4521) & (!x170x) & (n_n4531) & (x178x) & (!x361x)) + ((!n_n4521) & (!x170x) & (n_n4531) & (x178x) & (x361x)) + ((!n_n4521) & (x170x) & (!n_n4531) & (!x178x) & (!x361x)) + ((!n_n4521) & (x170x) & (!n_n4531) & (!x178x) & (x361x)) + ((!n_n4521) & (x170x) & (!n_n4531) & (x178x) & (!x361x)) + ((!n_n4521) & (x170x) & (!n_n4531) & (x178x) & (x361x)) + ((!n_n4521) & (x170x) & (n_n4531) & (!x178x) & (!x361x)) + ((!n_n4521) & (x170x) & (n_n4531) & (!x178x) & (x361x)) + ((!n_n4521) & (x170x) & (n_n4531) & (x178x) & (!x361x)) + ((!n_n4521) & (x170x) & (n_n4531) & (x178x) & (x361x)) + ((n_n4521) & (!x170x) & (!n_n4531) & (!x178x) & (!x361x)) + ((n_n4521) & (!x170x) & (!n_n4531) & (!x178x) & (x361x)) + ((n_n4521) & (!x170x) & (!n_n4531) & (x178x) & (!x361x)) + ((n_n4521) & (!x170x) & (!n_n4531) & (x178x) & (x361x)) + ((n_n4521) & (!x170x) & (n_n4531) & (!x178x) & (!x361x)) + ((n_n4521) & (!x170x) & (n_n4531) & (!x178x) & (x361x)) + ((n_n4521) & (!x170x) & (n_n4531) & (x178x) & (!x361x)) + ((n_n4521) & (!x170x) & (n_n4531) & (x178x) & (x361x)) + ((n_n4521) & (x170x) & (!n_n4531) & (!x178x) & (!x361x)) + ((n_n4521) & (x170x) & (!n_n4531) & (!x178x) & (x361x)) + ((n_n4521) & (x170x) & (!n_n4531) & (x178x) & (!x361x)) + ((n_n4521) & (x170x) & (!n_n4531) & (x178x) & (x361x)) + ((n_n4521) & (x170x) & (n_n4531) & (!x178x) & (!x361x)) + ((n_n4521) & (x170x) & (n_n4531) & (!x178x) & (x361x)) + ((n_n4521) & (x170x) & (n_n4531) & (x178x) & (!x361x)) + ((n_n4521) & (x170x) & (n_n4531) & (x178x) & (x361x)));
	assign x12369x = (((!n_n5318) & (!n_n5320) & (!n_n5312) & (!n_n5311) & (n_n5309)) + ((!n_n5318) & (!n_n5320) & (!n_n5312) & (n_n5311) & (!n_n5309)) + ((!n_n5318) & (!n_n5320) & (!n_n5312) & (n_n5311) & (n_n5309)) + ((!n_n5318) & (!n_n5320) & (n_n5312) & (!n_n5311) & (!n_n5309)) + ((!n_n5318) & (!n_n5320) & (n_n5312) & (!n_n5311) & (n_n5309)) + ((!n_n5318) & (!n_n5320) & (n_n5312) & (n_n5311) & (!n_n5309)) + ((!n_n5318) & (!n_n5320) & (n_n5312) & (n_n5311) & (n_n5309)) + ((!n_n5318) & (n_n5320) & (!n_n5312) & (!n_n5311) & (!n_n5309)) + ((!n_n5318) & (n_n5320) & (!n_n5312) & (!n_n5311) & (n_n5309)) + ((!n_n5318) & (n_n5320) & (!n_n5312) & (n_n5311) & (!n_n5309)) + ((!n_n5318) & (n_n5320) & (!n_n5312) & (n_n5311) & (n_n5309)) + ((!n_n5318) & (n_n5320) & (n_n5312) & (!n_n5311) & (!n_n5309)) + ((!n_n5318) & (n_n5320) & (n_n5312) & (!n_n5311) & (n_n5309)) + ((!n_n5318) & (n_n5320) & (n_n5312) & (n_n5311) & (!n_n5309)) + ((!n_n5318) & (n_n5320) & (n_n5312) & (n_n5311) & (n_n5309)) + ((n_n5318) & (!n_n5320) & (!n_n5312) & (!n_n5311) & (!n_n5309)) + ((n_n5318) & (!n_n5320) & (!n_n5312) & (!n_n5311) & (n_n5309)) + ((n_n5318) & (!n_n5320) & (!n_n5312) & (n_n5311) & (!n_n5309)) + ((n_n5318) & (!n_n5320) & (!n_n5312) & (n_n5311) & (n_n5309)) + ((n_n5318) & (!n_n5320) & (n_n5312) & (!n_n5311) & (!n_n5309)) + ((n_n5318) & (!n_n5320) & (n_n5312) & (!n_n5311) & (n_n5309)) + ((n_n5318) & (!n_n5320) & (n_n5312) & (n_n5311) & (!n_n5309)) + ((n_n5318) & (!n_n5320) & (n_n5312) & (n_n5311) & (n_n5309)) + ((n_n5318) & (n_n5320) & (!n_n5312) & (!n_n5311) & (!n_n5309)) + ((n_n5318) & (n_n5320) & (!n_n5312) & (!n_n5311) & (n_n5309)) + ((n_n5318) & (n_n5320) & (!n_n5312) & (n_n5311) & (!n_n5309)) + ((n_n5318) & (n_n5320) & (!n_n5312) & (n_n5311) & (n_n5309)) + ((n_n5318) & (n_n5320) & (n_n5312) & (!n_n5311) & (!n_n5309)) + ((n_n5318) & (n_n5320) & (n_n5312) & (!n_n5311) & (n_n5309)) + ((n_n5318) & (n_n5320) & (n_n5312) & (n_n5311) & (!n_n5309)) + ((n_n5318) & (n_n5320) & (n_n5312) & (n_n5311) & (n_n5309)));
	assign n_n1429 = (((!n_n5325) & (!n_n5332) & (!n_n5324) & (!n_n5334) & (x12364x)) + ((!n_n5325) & (!n_n5332) & (!n_n5324) & (n_n5334) & (!x12364x)) + ((!n_n5325) & (!n_n5332) & (!n_n5324) & (n_n5334) & (x12364x)) + ((!n_n5325) & (!n_n5332) & (n_n5324) & (!n_n5334) & (!x12364x)) + ((!n_n5325) & (!n_n5332) & (n_n5324) & (!n_n5334) & (x12364x)) + ((!n_n5325) & (!n_n5332) & (n_n5324) & (n_n5334) & (!x12364x)) + ((!n_n5325) & (!n_n5332) & (n_n5324) & (n_n5334) & (x12364x)) + ((!n_n5325) & (n_n5332) & (!n_n5324) & (!n_n5334) & (!x12364x)) + ((!n_n5325) & (n_n5332) & (!n_n5324) & (!n_n5334) & (x12364x)) + ((!n_n5325) & (n_n5332) & (!n_n5324) & (n_n5334) & (!x12364x)) + ((!n_n5325) & (n_n5332) & (!n_n5324) & (n_n5334) & (x12364x)) + ((!n_n5325) & (n_n5332) & (n_n5324) & (!n_n5334) & (!x12364x)) + ((!n_n5325) & (n_n5332) & (n_n5324) & (!n_n5334) & (x12364x)) + ((!n_n5325) & (n_n5332) & (n_n5324) & (n_n5334) & (!x12364x)) + ((!n_n5325) & (n_n5332) & (n_n5324) & (n_n5334) & (x12364x)) + ((n_n5325) & (!n_n5332) & (!n_n5324) & (!n_n5334) & (!x12364x)) + ((n_n5325) & (!n_n5332) & (!n_n5324) & (!n_n5334) & (x12364x)) + ((n_n5325) & (!n_n5332) & (!n_n5324) & (n_n5334) & (!x12364x)) + ((n_n5325) & (!n_n5332) & (!n_n5324) & (n_n5334) & (x12364x)) + ((n_n5325) & (!n_n5332) & (n_n5324) & (!n_n5334) & (!x12364x)) + ((n_n5325) & (!n_n5332) & (n_n5324) & (!n_n5334) & (x12364x)) + ((n_n5325) & (!n_n5332) & (n_n5324) & (n_n5334) & (!x12364x)) + ((n_n5325) & (!n_n5332) & (n_n5324) & (n_n5334) & (x12364x)) + ((n_n5325) & (n_n5332) & (!n_n5324) & (!n_n5334) & (!x12364x)) + ((n_n5325) & (n_n5332) & (!n_n5324) & (!n_n5334) & (x12364x)) + ((n_n5325) & (n_n5332) & (!n_n5324) & (n_n5334) & (!x12364x)) + ((n_n5325) & (n_n5332) & (!n_n5324) & (n_n5334) & (x12364x)) + ((n_n5325) & (n_n5332) & (n_n5324) & (!n_n5334) & (!x12364x)) + ((n_n5325) & (n_n5332) & (n_n5324) & (!n_n5334) & (x12364x)) + ((n_n5325) & (n_n5332) & (n_n5324) & (n_n5334) & (!x12364x)) + ((n_n5325) & (n_n5332) & (n_n5324) & (n_n5334) & (x12364x)));
	assign x12368x = (((!x19x) & (!n_n524) & (!n_n473) & (!n_n5322) & (x115x)) + ((!x19x) & (!n_n524) & (!n_n473) & (n_n5322) & (!x115x)) + ((!x19x) & (!n_n524) & (!n_n473) & (n_n5322) & (x115x)) + ((!x19x) & (!n_n524) & (n_n473) & (!n_n5322) & (x115x)) + ((!x19x) & (!n_n524) & (n_n473) & (n_n5322) & (!x115x)) + ((!x19x) & (!n_n524) & (n_n473) & (n_n5322) & (x115x)) + ((!x19x) & (n_n524) & (!n_n473) & (!n_n5322) & (x115x)) + ((!x19x) & (n_n524) & (!n_n473) & (n_n5322) & (!x115x)) + ((!x19x) & (n_n524) & (!n_n473) & (n_n5322) & (x115x)) + ((!x19x) & (n_n524) & (n_n473) & (!n_n5322) & (x115x)) + ((!x19x) & (n_n524) & (n_n473) & (n_n5322) & (!x115x)) + ((!x19x) & (n_n524) & (n_n473) & (n_n5322) & (x115x)) + ((x19x) & (!n_n524) & (!n_n473) & (!n_n5322) & (x115x)) + ((x19x) & (!n_n524) & (!n_n473) & (n_n5322) & (!x115x)) + ((x19x) & (!n_n524) & (!n_n473) & (n_n5322) & (x115x)) + ((x19x) & (!n_n524) & (n_n473) & (!n_n5322) & (x115x)) + ((x19x) & (!n_n524) & (n_n473) & (n_n5322) & (!x115x)) + ((x19x) & (!n_n524) & (n_n473) & (n_n5322) & (x115x)) + ((x19x) & (n_n524) & (!n_n473) & (!n_n5322) & (x115x)) + ((x19x) & (n_n524) & (!n_n473) & (n_n5322) & (!x115x)) + ((x19x) & (n_n524) & (!n_n473) & (n_n5322) & (x115x)) + ((x19x) & (n_n524) & (n_n473) & (!n_n5322) & (!x115x)) + ((x19x) & (n_n524) & (n_n473) & (!n_n5322) & (x115x)) + ((x19x) & (n_n524) & (n_n473) & (n_n5322) & (!x115x)) + ((x19x) & (n_n524) & (n_n473) & (n_n5322) & (x115x)));
	assign x12379x = (((!n_n5305) & (!x592x) & (!x21x) & (!n_n3019) & (x204x)) + ((!n_n5305) & (!x592x) & (!x21x) & (n_n3019) & (!x204x)) + ((!n_n5305) & (!x592x) & (!x21x) & (n_n3019) & (x204x)) + ((!n_n5305) & (!x592x) & (x21x) & (!n_n3019) & (x204x)) + ((!n_n5305) & (!x592x) & (x21x) & (n_n3019) & (!x204x)) + ((!n_n5305) & (!x592x) & (x21x) & (n_n3019) & (x204x)) + ((!n_n5305) & (x592x) & (!x21x) & (!n_n3019) & (x204x)) + ((!n_n5305) & (x592x) & (!x21x) & (n_n3019) & (!x204x)) + ((!n_n5305) & (x592x) & (!x21x) & (n_n3019) & (x204x)) + ((!n_n5305) & (x592x) & (x21x) & (!n_n3019) & (!x204x)) + ((!n_n5305) & (x592x) & (x21x) & (!n_n3019) & (x204x)) + ((!n_n5305) & (x592x) & (x21x) & (n_n3019) & (!x204x)) + ((!n_n5305) & (x592x) & (x21x) & (n_n3019) & (x204x)) + ((n_n5305) & (!x592x) & (!x21x) & (!n_n3019) & (!x204x)) + ((n_n5305) & (!x592x) & (!x21x) & (!n_n3019) & (x204x)) + ((n_n5305) & (!x592x) & (!x21x) & (n_n3019) & (!x204x)) + ((n_n5305) & (!x592x) & (!x21x) & (n_n3019) & (x204x)) + ((n_n5305) & (!x592x) & (x21x) & (!n_n3019) & (!x204x)) + ((n_n5305) & (!x592x) & (x21x) & (!n_n3019) & (x204x)) + ((n_n5305) & (!x592x) & (x21x) & (n_n3019) & (!x204x)) + ((n_n5305) & (!x592x) & (x21x) & (n_n3019) & (x204x)) + ((n_n5305) & (x592x) & (!x21x) & (!n_n3019) & (!x204x)) + ((n_n5305) & (x592x) & (!x21x) & (!n_n3019) & (x204x)) + ((n_n5305) & (x592x) & (!x21x) & (n_n3019) & (!x204x)) + ((n_n5305) & (x592x) & (!x21x) & (n_n3019) & (x204x)) + ((n_n5305) & (x592x) & (x21x) & (!n_n3019) & (!x204x)) + ((n_n5305) & (x592x) & (x21x) & (!n_n3019) & (x204x)) + ((n_n5305) & (x592x) & (x21x) & (n_n3019) & (!x204x)) + ((n_n5305) & (x592x) & (x21x) & (n_n3019) & (x204x)));
	assign x12381x = (((!x12369x) & (!n_n1429) & (!x12368x) & (x12379x)) + ((!x12369x) & (!n_n1429) & (x12368x) & (!x12379x)) + ((!x12369x) & (!n_n1429) & (x12368x) & (x12379x)) + ((!x12369x) & (n_n1429) & (!x12368x) & (!x12379x)) + ((!x12369x) & (n_n1429) & (!x12368x) & (x12379x)) + ((!x12369x) & (n_n1429) & (x12368x) & (!x12379x)) + ((!x12369x) & (n_n1429) & (x12368x) & (x12379x)) + ((x12369x) & (!n_n1429) & (!x12368x) & (!x12379x)) + ((x12369x) & (!n_n1429) & (!x12368x) & (x12379x)) + ((x12369x) & (!n_n1429) & (x12368x) & (!x12379x)) + ((x12369x) & (!n_n1429) & (x12368x) & (x12379x)) + ((x12369x) & (n_n1429) & (!x12368x) & (!x12379x)) + ((x12369x) & (n_n1429) & (!x12368x) & (x12379x)) + ((x12369x) & (n_n1429) & (x12368x) & (!x12379x)) + ((x12369x) & (n_n1429) & (x12368x) & (x12379x)));
	assign x12380x = (((!n_n1432) & (!n_n5286) & (!x218x) & (!x63x) & (x60x)) + ((!n_n1432) & (!n_n5286) & (!x218x) & (x63x) & (!x60x)) + ((!n_n1432) & (!n_n5286) & (!x218x) & (x63x) & (x60x)) + ((!n_n1432) & (!n_n5286) & (x218x) & (!x63x) & (!x60x)) + ((!n_n1432) & (!n_n5286) & (x218x) & (!x63x) & (x60x)) + ((!n_n1432) & (!n_n5286) & (x218x) & (x63x) & (!x60x)) + ((!n_n1432) & (!n_n5286) & (x218x) & (x63x) & (x60x)) + ((!n_n1432) & (n_n5286) & (!x218x) & (!x63x) & (!x60x)) + ((!n_n1432) & (n_n5286) & (!x218x) & (!x63x) & (x60x)) + ((!n_n1432) & (n_n5286) & (!x218x) & (x63x) & (!x60x)) + ((!n_n1432) & (n_n5286) & (!x218x) & (x63x) & (x60x)) + ((!n_n1432) & (n_n5286) & (x218x) & (!x63x) & (!x60x)) + ((!n_n1432) & (n_n5286) & (x218x) & (!x63x) & (x60x)) + ((!n_n1432) & (n_n5286) & (x218x) & (x63x) & (!x60x)) + ((!n_n1432) & (n_n5286) & (x218x) & (x63x) & (x60x)) + ((n_n1432) & (!n_n5286) & (!x218x) & (!x63x) & (!x60x)) + ((n_n1432) & (!n_n5286) & (!x218x) & (!x63x) & (x60x)) + ((n_n1432) & (!n_n5286) & (!x218x) & (x63x) & (!x60x)) + ((n_n1432) & (!n_n5286) & (!x218x) & (x63x) & (x60x)) + ((n_n1432) & (!n_n5286) & (x218x) & (!x63x) & (!x60x)) + ((n_n1432) & (!n_n5286) & (x218x) & (!x63x) & (x60x)) + ((n_n1432) & (!n_n5286) & (x218x) & (x63x) & (!x60x)) + ((n_n1432) & (!n_n5286) & (x218x) & (x63x) & (x60x)) + ((n_n1432) & (n_n5286) & (!x218x) & (!x63x) & (!x60x)) + ((n_n1432) & (n_n5286) & (!x218x) & (!x63x) & (x60x)) + ((n_n1432) & (n_n5286) & (!x218x) & (x63x) & (!x60x)) + ((n_n1432) & (n_n5286) & (!x218x) & (x63x) & (x60x)) + ((n_n1432) & (n_n5286) & (x218x) & (!x63x) & (!x60x)) + ((n_n1432) & (n_n5286) & (x218x) & (!x63x) & (x60x)) + ((n_n1432) & (n_n5286) & (x218x) & (x63x) & (!x60x)) + ((n_n1432) & (n_n5286) & (x218x) & (x63x) & (x60x)));
	assign x11660x = (((!n_n4455) & (!n_n4420) & (!n_n4430) & (n_n4429)) + ((!n_n4455) & (!n_n4420) & (n_n4430) & (!n_n4429)) + ((!n_n4455) & (!n_n4420) & (n_n4430) & (n_n4429)) + ((!n_n4455) & (n_n4420) & (!n_n4430) & (!n_n4429)) + ((!n_n4455) & (n_n4420) & (!n_n4430) & (n_n4429)) + ((!n_n4455) & (n_n4420) & (n_n4430) & (!n_n4429)) + ((!n_n4455) & (n_n4420) & (n_n4430) & (n_n4429)) + ((n_n4455) & (!n_n4420) & (!n_n4430) & (!n_n4429)) + ((n_n4455) & (!n_n4420) & (!n_n4430) & (n_n4429)) + ((n_n4455) & (!n_n4420) & (n_n4430) & (!n_n4429)) + ((n_n4455) & (!n_n4420) & (n_n4430) & (n_n4429)) + ((n_n4455) & (n_n4420) & (!n_n4430) & (!n_n4429)) + ((n_n4455) & (n_n4420) & (!n_n4430) & (n_n4429)) + ((n_n4455) & (n_n4420) & (n_n4430) & (!n_n4429)) + ((n_n4455) & (n_n4420) & (n_n4430) & (n_n4429)));
	assign x11661x = (((!n_n4433) & (!x23x) & (!x496x) & (!n_n4394) & (x427x)) + ((!n_n4433) & (!x23x) & (!x496x) & (n_n4394) & (!x427x)) + ((!n_n4433) & (!x23x) & (!x496x) & (n_n4394) & (x427x)) + ((!n_n4433) & (!x23x) & (x496x) & (!n_n4394) & (x427x)) + ((!n_n4433) & (!x23x) & (x496x) & (n_n4394) & (!x427x)) + ((!n_n4433) & (!x23x) & (x496x) & (n_n4394) & (x427x)) + ((!n_n4433) & (x23x) & (!x496x) & (!n_n4394) & (x427x)) + ((!n_n4433) & (x23x) & (!x496x) & (n_n4394) & (!x427x)) + ((!n_n4433) & (x23x) & (!x496x) & (n_n4394) & (x427x)) + ((!n_n4433) & (x23x) & (x496x) & (!n_n4394) & (!x427x)) + ((!n_n4433) & (x23x) & (x496x) & (!n_n4394) & (x427x)) + ((!n_n4433) & (x23x) & (x496x) & (n_n4394) & (!x427x)) + ((!n_n4433) & (x23x) & (x496x) & (n_n4394) & (x427x)) + ((n_n4433) & (!x23x) & (!x496x) & (!n_n4394) & (!x427x)) + ((n_n4433) & (!x23x) & (!x496x) & (!n_n4394) & (x427x)) + ((n_n4433) & (!x23x) & (!x496x) & (n_n4394) & (!x427x)) + ((n_n4433) & (!x23x) & (!x496x) & (n_n4394) & (x427x)) + ((n_n4433) & (!x23x) & (x496x) & (!n_n4394) & (!x427x)) + ((n_n4433) & (!x23x) & (x496x) & (!n_n4394) & (x427x)) + ((n_n4433) & (!x23x) & (x496x) & (n_n4394) & (!x427x)) + ((n_n4433) & (!x23x) & (x496x) & (n_n4394) & (x427x)) + ((n_n4433) & (x23x) & (!x496x) & (!n_n4394) & (!x427x)) + ((n_n4433) & (x23x) & (!x496x) & (!n_n4394) & (x427x)) + ((n_n4433) & (x23x) & (!x496x) & (n_n4394) & (!x427x)) + ((n_n4433) & (x23x) & (!x496x) & (n_n4394) & (x427x)) + ((n_n4433) & (x23x) & (x496x) & (!n_n4394) & (!x427x)) + ((n_n4433) & (x23x) & (x496x) & (!n_n4394) & (x427x)) + ((n_n4433) & (x23x) & (x496x) & (n_n4394) & (!x427x)) + ((n_n4433) & (x23x) & (x496x) & (n_n4394) & (x427x)));
	assign x11667x = (((!n_n4477) & (!n_n4505) & (!n_n4496) & (n_n4490)) + ((!n_n4477) & (!n_n4505) & (n_n4496) & (!n_n4490)) + ((!n_n4477) & (!n_n4505) & (n_n4496) & (n_n4490)) + ((!n_n4477) & (n_n4505) & (!n_n4496) & (!n_n4490)) + ((!n_n4477) & (n_n4505) & (!n_n4496) & (n_n4490)) + ((!n_n4477) & (n_n4505) & (n_n4496) & (!n_n4490)) + ((!n_n4477) & (n_n4505) & (n_n4496) & (n_n4490)) + ((n_n4477) & (!n_n4505) & (!n_n4496) & (!n_n4490)) + ((n_n4477) & (!n_n4505) & (!n_n4496) & (n_n4490)) + ((n_n4477) & (!n_n4505) & (n_n4496) & (!n_n4490)) + ((n_n4477) & (!n_n4505) & (n_n4496) & (n_n4490)) + ((n_n4477) & (n_n4505) & (!n_n4496) & (!n_n4490)) + ((n_n4477) & (n_n4505) & (!n_n4496) & (n_n4490)) + ((n_n4477) & (n_n4505) & (n_n4496) & (!n_n4490)) + ((n_n4477) & (n_n4505) & (n_n4496) & (n_n4490)));
	assign x11668x = (((!n_n4468) & (!n_n4518) & (!n_n4500) & (!n_n4479) & (n_n4476)) + ((!n_n4468) & (!n_n4518) & (!n_n4500) & (n_n4479) & (!n_n4476)) + ((!n_n4468) & (!n_n4518) & (!n_n4500) & (n_n4479) & (n_n4476)) + ((!n_n4468) & (!n_n4518) & (n_n4500) & (!n_n4479) & (!n_n4476)) + ((!n_n4468) & (!n_n4518) & (n_n4500) & (!n_n4479) & (n_n4476)) + ((!n_n4468) & (!n_n4518) & (n_n4500) & (n_n4479) & (!n_n4476)) + ((!n_n4468) & (!n_n4518) & (n_n4500) & (n_n4479) & (n_n4476)) + ((!n_n4468) & (n_n4518) & (!n_n4500) & (!n_n4479) & (!n_n4476)) + ((!n_n4468) & (n_n4518) & (!n_n4500) & (!n_n4479) & (n_n4476)) + ((!n_n4468) & (n_n4518) & (!n_n4500) & (n_n4479) & (!n_n4476)) + ((!n_n4468) & (n_n4518) & (!n_n4500) & (n_n4479) & (n_n4476)) + ((!n_n4468) & (n_n4518) & (n_n4500) & (!n_n4479) & (!n_n4476)) + ((!n_n4468) & (n_n4518) & (n_n4500) & (!n_n4479) & (n_n4476)) + ((!n_n4468) & (n_n4518) & (n_n4500) & (n_n4479) & (!n_n4476)) + ((!n_n4468) & (n_n4518) & (n_n4500) & (n_n4479) & (n_n4476)) + ((n_n4468) & (!n_n4518) & (!n_n4500) & (!n_n4479) & (!n_n4476)) + ((n_n4468) & (!n_n4518) & (!n_n4500) & (!n_n4479) & (n_n4476)) + ((n_n4468) & (!n_n4518) & (!n_n4500) & (n_n4479) & (!n_n4476)) + ((n_n4468) & (!n_n4518) & (!n_n4500) & (n_n4479) & (n_n4476)) + ((n_n4468) & (!n_n4518) & (n_n4500) & (!n_n4479) & (!n_n4476)) + ((n_n4468) & (!n_n4518) & (n_n4500) & (!n_n4479) & (n_n4476)) + ((n_n4468) & (!n_n4518) & (n_n4500) & (n_n4479) & (!n_n4476)) + ((n_n4468) & (!n_n4518) & (n_n4500) & (n_n4479) & (n_n4476)) + ((n_n4468) & (n_n4518) & (!n_n4500) & (!n_n4479) & (!n_n4476)) + ((n_n4468) & (n_n4518) & (!n_n4500) & (!n_n4479) & (n_n4476)) + ((n_n4468) & (n_n4518) & (!n_n4500) & (n_n4479) & (!n_n4476)) + ((n_n4468) & (n_n4518) & (!n_n4500) & (n_n4479) & (n_n4476)) + ((n_n4468) & (n_n4518) & (n_n4500) & (!n_n4479) & (!n_n4476)) + ((n_n4468) & (n_n4518) & (n_n4500) & (!n_n4479) & (n_n4476)) + ((n_n4468) & (n_n4518) & (n_n4500) & (n_n4479) & (!n_n4476)) + ((n_n4468) & (n_n4518) & (n_n4500) & (n_n4479) & (n_n4476)));
	assign n_n951 = (((!n_n4830) & (!n_n4831) & (!n_n4857) & (!n_n4847) & (x11682x)) + ((!n_n4830) & (!n_n4831) & (!n_n4857) & (n_n4847) & (!x11682x)) + ((!n_n4830) & (!n_n4831) & (!n_n4857) & (n_n4847) & (x11682x)) + ((!n_n4830) & (!n_n4831) & (n_n4857) & (!n_n4847) & (!x11682x)) + ((!n_n4830) & (!n_n4831) & (n_n4857) & (!n_n4847) & (x11682x)) + ((!n_n4830) & (!n_n4831) & (n_n4857) & (n_n4847) & (!x11682x)) + ((!n_n4830) & (!n_n4831) & (n_n4857) & (n_n4847) & (x11682x)) + ((!n_n4830) & (n_n4831) & (!n_n4857) & (!n_n4847) & (!x11682x)) + ((!n_n4830) & (n_n4831) & (!n_n4857) & (!n_n4847) & (x11682x)) + ((!n_n4830) & (n_n4831) & (!n_n4857) & (n_n4847) & (!x11682x)) + ((!n_n4830) & (n_n4831) & (!n_n4857) & (n_n4847) & (x11682x)) + ((!n_n4830) & (n_n4831) & (n_n4857) & (!n_n4847) & (!x11682x)) + ((!n_n4830) & (n_n4831) & (n_n4857) & (!n_n4847) & (x11682x)) + ((!n_n4830) & (n_n4831) & (n_n4857) & (n_n4847) & (!x11682x)) + ((!n_n4830) & (n_n4831) & (n_n4857) & (n_n4847) & (x11682x)) + ((n_n4830) & (!n_n4831) & (!n_n4857) & (!n_n4847) & (!x11682x)) + ((n_n4830) & (!n_n4831) & (!n_n4857) & (!n_n4847) & (x11682x)) + ((n_n4830) & (!n_n4831) & (!n_n4857) & (n_n4847) & (!x11682x)) + ((n_n4830) & (!n_n4831) & (!n_n4857) & (n_n4847) & (x11682x)) + ((n_n4830) & (!n_n4831) & (n_n4857) & (!n_n4847) & (!x11682x)) + ((n_n4830) & (!n_n4831) & (n_n4857) & (!n_n4847) & (x11682x)) + ((n_n4830) & (!n_n4831) & (n_n4857) & (n_n4847) & (!x11682x)) + ((n_n4830) & (!n_n4831) & (n_n4857) & (n_n4847) & (x11682x)) + ((n_n4830) & (n_n4831) & (!n_n4857) & (!n_n4847) & (!x11682x)) + ((n_n4830) & (n_n4831) & (!n_n4857) & (!n_n4847) & (x11682x)) + ((n_n4830) & (n_n4831) & (!n_n4857) & (n_n4847) & (!x11682x)) + ((n_n4830) & (n_n4831) & (!n_n4857) & (n_n4847) & (x11682x)) + ((n_n4830) & (n_n4831) & (n_n4857) & (!n_n4847) & (!x11682x)) + ((n_n4830) & (n_n4831) & (n_n4857) & (!n_n4847) & (x11682x)) + ((n_n4830) & (n_n4831) & (n_n4857) & (n_n4847) & (!x11682x)) + ((n_n4830) & (n_n4831) & (n_n4857) & (n_n4847) & (x11682x)));
	assign x11688x = (((!n_n4907) & (!n_n4879) & (!n_n4936) & (n_n4947)) + ((!n_n4907) & (!n_n4879) & (n_n4936) & (!n_n4947)) + ((!n_n4907) & (!n_n4879) & (n_n4936) & (n_n4947)) + ((!n_n4907) & (n_n4879) & (!n_n4936) & (!n_n4947)) + ((!n_n4907) & (n_n4879) & (!n_n4936) & (n_n4947)) + ((!n_n4907) & (n_n4879) & (n_n4936) & (!n_n4947)) + ((!n_n4907) & (n_n4879) & (n_n4936) & (n_n4947)) + ((n_n4907) & (!n_n4879) & (!n_n4936) & (!n_n4947)) + ((n_n4907) & (!n_n4879) & (!n_n4936) & (n_n4947)) + ((n_n4907) & (!n_n4879) & (n_n4936) & (!n_n4947)) + ((n_n4907) & (!n_n4879) & (n_n4936) & (n_n4947)) + ((n_n4907) & (n_n4879) & (!n_n4936) & (!n_n4947)) + ((n_n4907) & (n_n4879) & (!n_n4936) & (n_n4947)) + ((n_n4907) & (n_n4879) & (n_n4936) & (!n_n4947)) + ((n_n4907) & (n_n4879) & (n_n4936) & (n_n4947)));
	assign x11689x = (((!n_n4998) & (!n_n4887) & (!n_n4967) & (!n_n4986) & (n_n4915)) + ((!n_n4998) & (!n_n4887) & (!n_n4967) & (n_n4986) & (!n_n4915)) + ((!n_n4998) & (!n_n4887) & (!n_n4967) & (n_n4986) & (n_n4915)) + ((!n_n4998) & (!n_n4887) & (n_n4967) & (!n_n4986) & (!n_n4915)) + ((!n_n4998) & (!n_n4887) & (n_n4967) & (!n_n4986) & (n_n4915)) + ((!n_n4998) & (!n_n4887) & (n_n4967) & (n_n4986) & (!n_n4915)) + ((!n_n4998) & (!n_n4887) & (n_n4967) & (n_n4986) & (n_n4915)) + ((!n_n4998) & (n_n4887) & (!n_n4967) & (!n_n4986) & (!n_n4915)) + ((!n_n4998) & (n_n4887) & (!n_n4967) & (!n_n4986) & (n_n4915)) + ((!n_n4998) & (n_n4887) & (!n_n4967) & (n_n4986) & (!n_n4915)) + ((!n_n4998) & (n_n4887) & (!n_n4967) & (n_n4986) & (n_n4915)) + ((!n_n4998) & (n_n4887) & (n_n4967) & (!n_n4986) & (!n_n4915)) + ((!n_n4998) & (n_n4887) & (n_n4967) & (!n_n4986) & (n_n4915)) + ((!n_n4998) & (n_n4887) & (n_n4967) & (n_n4986) & (!n_n4915)) + ((!n_n4998) & (n_n4887) & (n_n4967) & (n_n4986) & (n_n4915)) + ((n_n4998) & (!n_n4887) & (!n_n4967) & (!n_n4986) & (!n_n4915)) + ((n_n4998) & (!n_n4887) & (!n_n4967) & (!n_n4986) & (n_n4915)) + ((n_n4998) & (!n_n4887) & (!n_n4967) & (n_n4986) & (!n_n4915)) + ((n_n4998) & (!n_n4887) & (!n_n4967) & (n_n4986) & (n_n4915)) + ((n_n4998) & (!n_n4887) & (n_n4967) & (!n_n4986) & (!n_n4915)) + ((n_n4998) & (!n_n4887) & (n_n4967) & (!n_n4986) & (n_n4915)) + ((n_n4998) & (!n_n4887) & (n_n4967) & (n_n4986) & (!n_n4915)) + ((n_n4998) & (!n_n4887) & (n_n4967) & (n_n4986) & (n_n4915)) + ((n_n4998) & (n_n4887) & (!n_n4967) & (!n_n4986) & (!n_n4915)) + ((n_n4998) & (n_n4887) & (!n_n4967) & (!n_n4986) & (n_n4915)) + ((n_n4998) & (n_n4887) & (!n_n4967) & (n_n4986) & (!n_n4915)) + ((n_n4998) & (n_n4887) & (!n_n4967) & (n_n4986) & (n_n4915)) + ((n_n4998) & (n_n4887) & (n_n4967) & (!n_n4986) & (!n_n4915)) + ((n_n4998) & (n_n4887) & (n_n4967) & (!n_n4986) & (n_n4915)) + ((n_n4998) & (n_n4887) & (n_n4967) & (n_n4986) & (!n_n4915)) + ((n_n4998) & (n_n4887) & (n_n4967) & (n_n4986) & (n_n4915)));
	assign n_n941 = (((!x11675x) & (!x11676x) & (!n_n951) & (!x11688x) & (x11689x)) + ((!x11675x) & (!x11676x) & (!n_n951) & (x11688x) & (!x11689x)) + ((!x11675x) & (!x11676x) & (!n_n951) & (x11688x) & (x11689x)) + ((!x11675x) & (!x11676x) & (n_n951) & (!x11688x) & (!x11689x)) + ((!x11675x) & (!x11676x) & (n_n951) & (!x11688x) & (x11689x)) + ((!x11675x) & (!x11676x) & (n_n951) & (x11688x) & (!x11689x)) + ((!x11675x) & (!x11676x) & (n_n951) & (x11688x) & (x11689x)) + ((!x11675x) & (x11676x) & (!n_n951) & (!x11688x) & (!x11689x)) + ((!x11675x) & (x11676x) & (!n_n951) & (!x11688x) & (x11689x)) + ((!x11675x) & (x11676x) & (!n_n951) & (x11688x) & (!x11689x)) + ((!x11675x) & (x11676x) & (!n_n951) & (x11688x) & (x11689x)) + ((!x11675x) & (x11676x) & (n_n951) & (!x11688x) & (!x11689x)) + ((!x11675x) & (x11676x) & (n_n951) & (!x11688x) & (x11689x)) + ((!x11675x) & (x11676x) & (n_n951) & (x11688x) & (!x11689x)) + ((!x11675x) & (x11676x) & (n_n951) & (x11688x) & (x11689x)) + ((x11675x) & (!x11676x) & (!n_n951) & (!x11688x) & (!x11689x)) + ((x11675x) & (!x11676x) & (!n_n951) & (!x11688x) & (x11689x)) + ((x11675x) & (!x11676x) & (!n_n951) & (x11688x) & (!x11689x)) + ((x11675x) & (!x11676x) & (!n_n951) & (x11688x) & (x11689x)) + ((x11675x) & (!x11676x) & (n_n951) & (!x11688x) & (!x11689x)) + ((x11675x) & (!x11676x) & (n_n951) & (!x11688x) & (x11689x)) + ((x11675x) & (!x11676x) & (n_n951) & (x11688x) & (!x11689x)) + ((x11675x) & (!x11676x) & (n_n951) & (x11688x) & (x11689x)) + ((x11675x) & (x11676x) & (!n_n951) & (!x11688x) & (!x11689x)) + ((x11675x) & (x11676x) & (!n_n951) & (!x11688x) & (x11689x)) + ((x11675x) & (x11676x) & (!n_n951) & (x11688x) & (!x11689x)) + ((x11675x) & (x11676x) & (!n_n951) & (x11688x) & (x11689x)) + ((x11675x) & (x11676x) & (n_n951) & (!x11688x) & (!x11689x)) + ((x11675x) & (x11676x) & (n_n951) & (!x11688x) & (x11689x)) + ((x11675x) & (x11676x) & (n_n951) & (x11688x) & (!x11689x)) + ((x11675x) & (x11676x) & (n_n951) & (x11688x) & (x11689x)));
	assign x11719x = (((!n_n5085) & (!n_n5087) & (!n_n5106) & (n_n5070)) + ((!n_n5085) & (!n_n5087) & (n_n5106) & (!n_n5070)) + ((!n_n5085) & (!n_n5087) & (n_n5106) & (n_n5070)) + ((!n_n5085) & (n_n5087) & (!n_n5106) & (!n_n5070)) + ((!n_n5085) & (n_n5087) & (!n_n5106) & (n_n5070)) + ((!n_n5085) & (n_n5087) & (n_n5106) & (!n_n5070)) + ((!n_n5085) & (n_n5087) & (n_n5106) & (n_n5070)) + ((n_n5085) & (!n_n5087) & (!n_n5106) & (!n_n5070)) + ((n_n5085) & (!n_n5087) & (!n_n5106) & (n_n5070)) + ((n_n5085) & (!n_n5087) & (n_n5106) & (!n_n5070)) + ((n_n5085) & (!n_n5087) & (n_n5106) & (n_n5070)) + ((n_n5085) & (n_n5087) & (!n_n5106) & (!n_n5070)) + ((n_n5085) & (n_n5087) & (!n_n5106) & (n_n5070)) + ((n_n5085) & (n_n5087) & (n_n5106) & (!n_n5070)) + ((n_n5085) & (n_n5087) & (n_n5106) & (n_n5070)));
	assign x11720x = (((!n_n5093) & (!n_n5054) & (!n_n5063) & (!n_n5075) & (n_n5068)) + ((!n_n5093) & (!n_n5054) & (!n_n5063) & (n_n5075) & (!n_n5068)) + ((!n_n5093) & (!n_n5054) & (!n_n5063) & (n_n5075) & (n_n5068)) + ((!n_n5093) & (!n_n5054) & (n_n5063) & (!n_n5075) & (!n_n5068)) + ((!n_n5093) & (!n_n5054) & (n_n5063) & (!n_n5075) & (n_n5068)) + ((!n_n5093) & (!n_n5054) & (n_n5063) & (n_n5075) & (!n_n5068)) + ((!n_n5093) & (!n_n5054) & (n_n5063) & (n_n5075) & (n_n5068)) + ((!n_n5093) & (n_n5054) & (!n_n5063) & (!n_n5075) & (!n_n5068)) + ((!n_n5093) & (n_n5054) & (!n_n5063) & (!n_n5075) & (n_n5068)) + ((!n_n5093) & (n_n5054) & (!n_n5063) & (n_n5075) & (!n_n5068)) + ((!n_n5093) & (n_n5054) & (!n_n5063) & (n_n5075) & (n_n5068)) + ((!n_n5093) & (n_n5054) & (n_n5063) & (!n_n5075) & (!n_n5068)) + ((!n_n5093) & (n_n5054) & (n_n5063) & (!n_n5075) & (n_n5068)) + ((!n_n5093) & (n_n5054) & (n_n5063) & (n_n5075) & (!n_n5068)) + ((!n_n5093) & (n_n5054) & (n_n5063) & (n_n5075) & (n_n5068)) + ((n_n5093) & (!n_n5054) & (!n_n5063) & (!n_n5075) & (!n_n5068)) + ((n_n5093) & (!n_n5054) & (!n_n5063) & (!n_n5075) & (n_n5068)) + ((n_n5093) & (!n_n5054) & (!n_n5063) & (n_n5075) & (!n_n5068)) + ((n_n5093) & (!n_n5054) & (!n_n5063) & (n_n5075) & (n_n5068)) + ((n_n5093) & (!n_n5054) & (n_n5063) & (!n_n5075) & (!n_n5068)) + ((n_n5093) & (!n_n5054) & (n_n5063) & (!n_n5075) & (n_n5068)) + ((n_n5093) & (!n_n5054) & (n_n5063) & (n_n5075) & (!n_n5068)) + ((n_n5093) & (!n_n5054) & (n_n5063) & (n_n5075) & (n_n5068)) + ((n_n5093) & (n_n5054) & (!n_n5063) & (!n_n5075) & (!n_n5068)) + ((n_n5093) & (n_n5054) & (!n_n5063) & (!n_n5075) & (n_n5068)) + ((n_n5093) & (n_n5054) & (!n_n5063) & (n_n5075) & (!n_n5068)) + ((n_n5093) & (n_n5054) & (!n_n5063) & (n_n5075) & (n_n5068)) + ((n_n5093) & (n_n5054) & (n_n5063) & (!n_n5075) & (!n_n5068)) + ((n_n5093) & (n_n5054) & (n_n5063) & (!n_n5075) & (n_n5068)) + ((n_n5093) & (n_n5054) & (n_n5063) & (n_n5075) & (!n_n5068)) + ((n_n5093) & (n_n5054) & (n_n5063) & (n_n5075) & (n_n5068)));
	assign x11726x = (((!n_n5025) & (!n_n5049) & (!n_n5047) & (n_n5051)) + ((!n_n5025) & (!n_n5049) & (n_n5047) & (!n_n5051)) + ((!n_n5025) & (!n_n5049) & (n_n5047) & (n_n5051)) + ((!n_n5025) & (n_n5049) & (!n_n5047) & (!n_n5051)) + ((!n_n5025) & (n_n5049) & (!n_n5047) & (n_n5051)) + ((!n_n5025) & (n_n5049) & (n_n5047) & (!n_n5051)) + ((!n_n5025) & (n_n5049) & (n_n5047) & (n_n5051)) + ((n_n5025) & (!n_n5049) & (!n_n5047) & (!n_n5051)) + ((n_n5025) & (!n_n5049) & (!n_n5047) & (n_n5051)) + ((n_n5025) & (!n_n5049) & (n_n5047) & (!n_n5051)) + ((n_n5025) & (!n_n5049) & (n_n5047) & (n_n5051)) + ((n_n5025) & (n_n5049) & (!n_n5047) & (!n_n5051)) + ((n_n5025) & (n_n5049) & (!n_n5047) & (n_n5051)) + ((n_n5025) & (n_n5049) & (n_n5047) & (!n_n5051)) + ((n_n5025) & (n_n5049) & (n_n5047) & (n_n5051)));
	assign x11727x = (((!n_n5040) & (!n_n4999) & (!n_n5044) & (!n_n5011) & (n_n5024)) + ((!n_n5040) & (!n_n4999) & (!n_n5044) & (n_n5011) & (!n_n5024)) + ((!n_n5040) & (!n_n4999) & (!n_n5044) & (n_n5011) & (n_n5024)) + ((!n_n5040) & (!n_n4999) & (n_n5044) & (!n_n5011) & (!n_n5024)) + ((!n_n5040) & (!n_n4999) & (n_n5044) & (!n_n5011) & (n_n5024)) + ((!n_n5040) & (!n_n4999) & (n_n5044) & (n_n5011) & (!n_n5024)) + ((!n_n5040) & (!n_n4999) & (n_n5044) & (n_n5011) & (n_n5024)) + ((!n_n5040) & (n_n4999) & (!n_n5044) & (!n_n5011) & (!n_n5024)) + ((!n_n5040) & (n_n4999) & (!n_n5044) & (!n_n5011) & (n_n5024)) + ((!n_n5040) & (n_n4999) & (!n_n5044) & (n_n5011) & (!n_n5024)) + ((!n_n5040) & (n_n4999) & (!n_n5044) & (n_n5011) & (n_n5024)) + ((!n_n5040) & (n_n4999) & (n_n5044) & (!n_n5011) & (!n_n5024)) + ((!n_n5040) & (n_n4999) & (n_n5044) & (!n_n5011) & (n_n5024)) + ((!n_n5040) & (n_n4999) & (n_n5044) & (n_n5011) & (!n_n5024)) + ((!n_n5040) & (n_n4999) & (n_n5044) & (n_n5011) & (n_n5024)) + ((n_n5040) & (!n_n4999) & (!n_n5044) & (!n_n5011) & (!n_n5024)) + ((n_n5040) & (!n_n4999) & (!n_n5044) & (!n_n5011) & (n_n5024)) + ((n_n5040) & (!n_n4999) & (!n_n5044) & (n_n5011) & (!n_n5024)) + ((n_n5040) & (!n_n4999) & (!n_n5044) & (n_n5011) & (n_n5024)) + ((n_n5040) & (!n_n4999) & (n_n5044) & (!n_n5011) & (!n_n5024)) + ((n_n5040) & (!n_n4999) & (n_n5044) & (!n_n5011) & (n_n5024)) + ((n_n5040) & (!n_n4999) & (n_n5044) & (n_n5011) & (!n_n5024)) + ((n_n5040) & (!n_n4999) & (n_n5044) & (n_n5011) & (n_n5024)) + ((n_n5040) & (n_n4999) & (!n_n5044) & (!n_n5011) & (!n_n5024)) + ((n_n5040) & (n_n4999) & (!n_n5044) & (!n_n5011) & (n_n5024)) + ((n_n5040) & (n_n4999) & (!n_n5044) & (n_n5011) & (!n_n5024)) + ((n_n5040) & (n_n4999) & (!n_n5044) & (n_n5011) & (n_n5024)) + ((n_n5040) & (n_n4999) & (n_n5044) & (!n_n5011) & (!n_n5024)) + ((n_n5040) & (n_n4999) & (n_n5044) & (!n_n5011) & (n_n5024)) + ((n_n5040) & (n_n4999) & (n_n5044) & (n_n5011) & (!n_n5024)) + ((n_n5040) & (n_n4999) & (n_n5044) & (n_n5011) & (n_n5024)));
	assign x13343x = (((!n_n5239) & (!n_n5245) & (!n_n5241) & (!n_n5242) & (n_n5249)) + ((!n_n5239) & (!n_n5245) & (!n_n5241) & (n_n5242) & (!n_n5249)) + ((!n_n5239) & (!n_n5245) & (!n_n5241) & (n_n5242) & (n_n5249)) + ((!n_n5239) & (!n_n5245) & (n_n5241) & (!n_n5242) & (!n_n5249)) + ((!n_n5239) & (!n_n5245) & (n_n5241) & (!n_n5242) & (n_n5249)) + ((!n_n5239) & (!n_n5245) & (n_n5241) & (n_n5242) & (!n_n5249)) + ((!n_n5239) & (!n_n5245) & (n_n5241) & (n_n5242) & (n_n5249)) + ((!n_n5239) & (n_n5245) & (!n_n5241) & (!n_n5242) & (!n_n5249)) + ((!n_n5239) & (n_n5245) & (!n_n5241) & (!n_n5242) & (n_n5249)) + ((!n_n5239) & (n_n5245) & (!n_n5241) & (n_n5242) & (!n_n5249)) + ((!n_n5239) & (n_n5245) & (!n_n5241) & (n_n5242) & (n_n5249)) + ((!n_n5239) & (n_n5245) & (n_n5241) & (!n_n5242) & (!n_n5249)) + ((!n_n5239) & (n_n5245) & (n_n5241) & (!n_n5242) & (n_n5249)) + ((!n_n5239) & (n_n5245) & (n_n5241) & (n_n5242) & (!n_n5249)) + ((!n_n5239) & (n_n5245) & (n_n5241) & (n_n5242) & (n_n5249)) + ((n_n5239) & (!n_n5245) & (!n_n5241) & (!n_n5242) & (!n_n5249)) + ((n_n5239) & (!n_n5245) & (!n_n5241) & (!n_n5242) & (n_n5249)) + ((n_n5239) & (!n_n5245) & (!n_n5241) & (n_n5242) & (!n_n5249)) + ((n_n5239) & (!n_n5245) & (!n_n5241) & (n_n5242) & (n_n5249)) + ((n_n5239) & (!n_n5245) & (n_n5241) & (!n_n5242) & (!n_n5249)) + ((n_n5239) & (!n_n5245) & (n_n5241) & (!n_n5242) & (n_n5249)) + ((n_n5239) & (!n_n5245) & (n_n5241) & (n_n5242) & (!n_n5249)) + ((n_n5239) & (!n_n5245) & (n_n5241) & (n_n5242) & (n_n5249)) + ((n_n5239) & (n_n5245) & (!n_n5241) & (!n_n5242) & (!n_n5249)) + ((n_n5239) & (n_n5245) & (!n_n5241) & (!n_n5242) & (n_n5249)) + ((n_n5239) & (n_n5245) & (!n_n5241) & (n_n5242) & (!n_n5249)) + ((n_n5239) & (n_n5245) & (!n_n5241) & (n_n5242) & (n_n5249)) + ((n_n5239) & (n_n5245) & (n_n5241) & (!n_n5242) & (!n_n5249)) + ((n_n5239) & (n_n5245) & (n_n5241) & (!n_n5242) & (n_n5249)) + ((n_n5239) & (n_n5245) & (n_n5241) & (n_n5242) & (!n_n5249)) + ((n_n5239) & (n_n5245) & (n_n5241) & (n_n5242) & (n_n5249)));
	assign x14296x = (((!n_n4613) & (!n_n4619) & (!n_n4632) & (!n_n4610) & (n_n4627)) + ((!n_n4613) & (!n_n4619) & (!n_n4632) & (n_n4610) & (!n_n4627)) + ((!n_n4613) & (!n_n4619) & (!n_n4632) & (n_n4610) & (n_n4627)) + ((!n_n4613) & (!n_n4619) & (n_n4632) & (!n_n4610) & (!n_n4627)) + ((!n_n4613) & (!n_n4619) & (n_n4632) & (!n_n4610) & (n_n4627)) + ((!n_n4613) & (!n_n4619) & (n_n4632) & (n_n4610) & (!n_n4627)) + ((!n_n4613) & (!n_n4619) & (n_n4632) & (n_n4610) & (n_n4627)) + ((!n_n4613) & (n_n4619) & (!n_n4632) & (!n_n4610) & (!n_n4627)) + ((!n_n4613) & (n_n4619) & (!n_n4632) & (!n_n4610) & (n_n4627)) + ((!n_n4613) & (n_n4619) & (!n_n4632) & (n_n4610) & (!n_n4627)) + ((!n_n4613) & (n_n4619) & (!n_n4632) & (n_n4610) & (n_n4627)) + ((!n_n4613) & (n_n4619) & (n_n4632) & (!n_n4610) & (!n_n4627)) + ((!n_n4613) & (n_n4619) & (n_n4632) & (!n_n4610) & (n_n4627)) + ((!n_n4613) & (n_n4619) & (n_n4632) & (n_n4610) & (!n_n4627)) + ((!n_n4613) & (n_n4619) & (n_n4632) & (n_n4610) & (n_n4627)) + ((n_n4613) & (!n_n4619) & (!n_n4632) & (!n_n4610) & (!n_n4627)) + ((n_n4613) & (!n_n4619) & (!n_n4632) & (!n_n4610) & (n_n4627)) + ((n_n4613) & (!n_n4619) & (!n_n4632) & (n_n4610) & (!n_n4627)) + ((n_n4613) & (!n_n4619) & (!n_n4632) & (n_n4610) & (n_n4627)) + ((n_n4613) & (!n_n4619) & (n_n4632) & (!n_n4610) & (!n_n4627)) + ((n_n4613) & (!n_n4619) & (n_n4632) & (!n_n4610) & (n_n4627)) + ((n_n4613) & (!n_n4619) & (n_n4632) & (n_n4610) & (!n_n4627)) + ((n_n4613) & (!n_n4619) & (n_n4632) & (n_n4610) & (n_n4627)) + ((n_n4613) & (n_n4619) & (!n_n4632) & (!n_n4610) & (!n_n4627)) + ((n_n4613) & (n_n4619) & (!n_n4632) & (!n_n4610) & (n_n4627)) + ((n_n4613) & (n_n4619) & (!n_n4632) & (n_n4610) & (!n_n4627)) + ((n_n4613) & (n_n4619) & (!n_n4632) & (n_n4610) & (n_n4627)) + ((n_n4613) & (n_n4619) & (n_n4632) & (!n_n4610) & (!n_n4627)) + ((n_n4613) & (n_n4619) & (n_n4632) & (!n_n4610) & (n_n4627)) + ((n_n4613) & (n_n4619) & (n_n4632) & (n_n4610) & (!n_n4627)) + ((n_n4613) & (n_n4619) & (n_n4632) & (n_n4610) & (n_n4627)));
	assign n_n2036 = (((!i_9_) & (!n_n528) & (n_n390) & (n_n509) & (n_n530)) + ((!i_9_) & (n_n528) & (n_n390) & (n_n509) & (!n_n530)) + ((!i_9_) & (n_n528) & (n_n390) & (n_n509) & (n_n530)) + ((i_9_) & (n_n528) & (n_n390) & (n_n509) & (!n_n530)) + ((i_9_) & (n_n528) & (n_n390) & (n_n509) & (n_n530)));
	assign x22139x = (((!x21x) & (!x20x) & (!n_n4571) & (!n_n4570) & (!x523x)) + ((!x21x) & (!x20x) & (!n_n4571) & (!n_n4570) & (x523x)) + ((!x21x) & (x20x) & (!n_n4571) & (!n_n4570) & (!x523x)) + ((x21x) & (!x20x) & (!n_n4571) & (!n_n4570) & (!x523x)) + ((x21x) & (x20x) & (!n_n4571) & (!n_n4570) & (!x523x)));
	assign n_n1489 = (((!n_n4561) & (!n_n4568) & (!n_n4572) & (!x238x) & (!x22139x)) + ((!n_n4561) & (!n_n4568) & (!n_n4572) & (x238x) & (!x22139x)) + ((!n_n4561) & (!n_n4568) & (!n_n4572) & (x238x) & (x22139x)) + ((!n_n4561) & (!n_n4568) & (n_n4572) & (!x238x) & (!x22139x)) + ((!n_n4561) & (!n_n4568) & (n_n4572) & (!x238x) & (x22139x)) + ((!n_n4561) & (!n_n4568) & (n_n4572) & (x238x) & (!x22139x)) + ((!n_n4561) & (!n_n4568) & (n_n4572) & (x238x) & (x22139x)) + ((!n_n4561) & (n_n4568) & (!n_n4572) & (!x238x) & (!x22139x)) + ((!n_n4561) & (n_n4568) & (!n_n4572) & (!x238x) & (x22139x)) + ((!n_n4561) & (n_n4568) & (!n_n4572) & (x238x) & (!x22139x)) + ((!n_n4561) & (n_n4568) & (!n_n4572) & (x238x) & (x22139x)) + ((!n_n4561) & (n_n4568) & (n_n4572) & (!x238x) & (!x22139x)) + ((!n_n4561) & (n_n4568) & (n_n4572) & (!x238x) & (x22139x)) + ((!n_n4561) & (n_n4568) & (n_n4572) & (x238x) & (!x22139x)) + ((!n_n4561) & (n_n4568) & (n_n4572) & (x238x) & (x22139x)) + ((n_n4561) & (!n_n4568) & (!n_n4572) & (!x238x) & (!x22139x)) + ((n_n4561) & (!n_n4568) & (!n_n4572) & (!x238x) & (x22139x)) + ((n_n4561) & (!n_n4568) & (!n_n4572) & (x238x) & (!x22139x)) + ((n_n4561) & (!n_n4568) & (!n_n4572) & (x238x) & (x22139x)) + ((n_n4561) & (!n_n4568) & (n_n4572) & (!x238x) & (!x22139x)) + ((n_n4561) & (!n_n4568) & (n_n4572) & (!x238x) & (x22139x)) + ((n_n4561) & (!n_n4568) & (n_n4572) & (x238x) & (!x22139x)) + ((n_n4561) & (!n_n4568) & (n_n4572) & (x238x) & (x22139x)) + ((n_n4561) & (n_n4568) & (!n_n4572) & (!x238x) & (!x22139x)) + ((n_n4561) & (n_n4568) & (!n_n4572) & (!x238x) & (x22139x)) + ((n_n4561) & (n_n4568) & (!n_n4572) & (x238x) & (!x22139x)) + ((n_n4561) & (n_n4568) & (!n_n4572) & (x238x) & (x22139x)) + ((n_n4561) & (n_n4568) & (n_n4572) & (!x238x) & (!x22139x)) + ((n_n4561) & (n_n4568) & (n_n4572) & (!x238x) & (x22139x)) + ((n_n4561) & (n_n4568) & (n_n4572) & (x238x) & (!x22139x)) + ((n_n4561) & (n_n4568) & (n_n4572) & (x238x) & (x22139x)));
	assign x12531x = (((!n_n4554) & (!n_n4584) & (!n_n4577) & (n_n4556)) + ((!n_n4554) & (!n_n4584) & (n_n4577) & (!n_n4556)) + ((!n_n4554) & (!n_n4584) & (n_n4577) & (n_n4556)) + ((!n_n4554) & (n_n4584) & (!n_n4577) & (!n_n4556)) + ((!n_n4554) & (n_n4584) & (!n_n4577) & (n_n4556)) + ((!n_n4554) & (n_n4584) & (n_n4577) & (!n_n4556)) + ((!n_n4554) & (n_n4584) & (n_n4577) & (n_n4556)) + ((n_n4554) & (!n_n4584) & (!n_n4577) & (!n_n4556)) + ((n_n4554) & (!n_n4584) & (!n_n4577) & (n_n4556)) + ((n_n4554) & (!n_n4584) & (n_n4577) & (!n_n4556)) + ((n_n4554) & (!n_n4584) & (n_n4577) & (n_n4556)) + ((n_n4554) & (n_n4584) & (!n_n4577) & (!n_n4556)) + ((n_n4554) & (n_n4584) & (!n_n4577) & (n_n4556)) + ((n_n4554) & (n_n4584) & (n_n4577) & (!n_n4556)) + ((n_n4554) & (n_n4584) & (n_n4577) & (n_n4556)));
	assign x12533x = (((!n_n4557) & (!n_n4560) & (!x213x) & (!x276x) & (x237x)) + ((!n_n4557) & (!n_n4560) & (!x213x) & (x276x) & (!x237x)) + ((!n_n4557) & (!n_n4560) & (!x213x) & (x276x) & (x237x)) + ((!n_n4557) & (!n_n4560) & (x213x) & (!x276x) & (!x237x)) + ((!n_n4557) & (!n_n4560) & (x213x) & (!x276x) & (x237x)) + ((!n_n4557) & (!n_n4560) & (x213x) & (x276x) & (!x237x)) + ((!n_n4557) & (!n_n4560) & (x213x) & (x276x) & (x237x)) + ((!n_n4557) & (n_n4560) & (!x213x) & (!x276x) & (!x237x)) + ((!n_n4557) & (n_n4560) & (!x213x) & (!x276x) & (x237x)) + ((!n_n4557) & (n_n4560) & (!x213x) & (x276x) & (!x237x)) + ((!n_n4557) & (n_n4560) & (!x213x) & (x276x) & (x237x)) + ((!n_n4557) & (n_n4560) & (x213x) & (!x276x) & (!x237x)) + ((!n_n4557) & (n_n4560) & (x213x) & (!x276x) & (x237x)) + ((!n_n4557) & (n_n4560) & (x213x) & (x276x) & (!x237x)) + ((!n_n4557) & (n_n4560) & (x213x) & (x276x) & (x237x)) + ((n_n4557) & (!n_n4560) & (!x213x) & (!x276x) & (!x237x)) + ((n_n4557) & (!n_n4560) & (!x213x) & (!x276x) & (x237x)) + ((n_n4557) & (!n_n4560) & (!x213x) & (x276x) & (!x237x)) + ((n_n4557) & (!n_n4560) & (!x213x) & (x276x) & (x237x)) + ((n_n4557) & (!n_n4560) & (x213x) & (!x276x) & (!x237x)) + ((n_n4557) & (!n_n4560) & (x213x) & (!x276x) & (x237x)) + ((n_n4557) & (!n_n4560) & (x213x) & (x276x) & (!x237x)) + ((n_n4557) & (!n_n4560) & (x213x) & (x276x) & (x237x)) + ((n_n4557) & (n_n4560) & (!x213x) & (!x276x) & (!x237x)) + ((n_n4557) & (n_n4560) & (!x213x) & (!x276x) & (x237x)) + ((n_n4557) & (n_n4560) & (!x213x) & (x276x) & (!x237x)) + ((n_n4557) & (n_n4560) & (!x213x) & (x276x) & (x237x)) + ((n_n4557) & (n_n4560) & (x213x) & (!x276x) & (!x237x)) + ((n_n4557) & (n_n4560) & (x213x) & (!x276x) & (x237x)) + ((n_n4557) & (n_n4560) & (x213x) & (x276x) & (!x237x)) + ((n_n4557) & (n_n4560) & (x213x) & (x276x) & (x237x)));
	assign n_n1422 = (((!n_n3871) & (!n_n2401) & (!n_n1489) & (!x12531x) & (x12533x)) + ((!n_n3871) & (!n_n2401) & (!n_n1489) & (x12531x) & (!x12533x)) + ((!n_n3871) & (!n_n2401) & (!n_n1489) & (x12531x) & (x12533x)) + ((!n_n3871) & (!n_n2401) & (n_n1489) & (!x12531x) & (!x12533x)) + ((!n_n3871) & (!n_n2401) & (n_n1489) & (!x12531x) & (x12533x)) + ((!n_n3871) & (!n_n2401) & (n_n1489) & (x12531x) & (!x12533x)) + ((!n_n3871) & (!n_n2401) & (n_n1489) & (x12531x) & (x12533x)) + ((!n_n3871) & (n_n2401) & (!n_n1489) & (!x12531x) & (!x12533x)) + ((!n_n3871) & (n_n2401) & (!n_n1489) & (!x12531x) & (x12533x)) + ((!n_n3871) & (n_n2401) & (!n_n1489) & (x12531x) & (!x12533x)) + ((!n_n3871) & (n_n2401) & (!n_n1489) & (x12531x) & (x12533x)) + ((!n_n3871) & (n_n2401) & (n_n1489) & (!x12531x) & (!x12533x)) + ((!n_n3871) & (n_n2401) & (n_n1489) & (!x12531x) & (x12533x)) + ((!n_n3871) & (n_n2401) & (n_n1489) & (x12531x) & (!x12533x)) + ((!n_n3871) & (n_n2401) & (n_n1489) & (x12531x) & (x12533x)) + ((n_n3871) & (!n_n2401) & (!n_n1489) & (!x12531x) & (!x12533x)) + ((n_n3871) & (!n_n2401) & (!n_n1489) & (!x12531x) & (x12533x)) + ((n_n3871) & (!n_n2401) & (!n_n1489) & (x12531x) & (!x12533x)) + ((n_n3871) & (!n_n2401) & (!n_n1489) & (x12531x) & (x12533x)) + ((n_n3871) & (!n_n2401) & (n_n1489) & (!x12531x) & (!x12533x)) + ((n_n3871) & (!n_n2401) & (n_n1489) & (!x12531x) & (x12533x)) + ((n_n3871) & (!n_n2401) & (n_n1489) & (x12531x) & (!x12533x)) + ((n_n3871) & (!n_n2401) & (n_n1489) & (x12531x) & (x12533x)) + ((n_n3871) & (n_n2401) & (!n_n1489) & (!x12531x) & (!x12533x)) + ((n_n3871) & (n_n2401) & (!n_n1489) & (!x12531x) & (x12533x)) + ((n_n3871) & (n_n2401) & (!n_n1489) & (x12531x) & (!x12533x)) + ((n_n3871) & (n_n2401) & (!n_n1489) & (x12531x) & (x12533x)) + ((n_n3871) & (n_n2401) & (n_n1489) & (!x12531x) & (!x12533x)) + ((n_n3871) & (n_n2401) & (n_n1489) & (!x12531x) & (x12533x)) + ((n_n3871) & (n_n2401) & (n_n1489) & (x12531x) & (!x12533x)) + ((n_n3871) & (n_n2401) & (n_n1489) & (x12531x) & (x12533x)));
	assign x12513x = (((!n_n4504) & (!n_n4503) & (!n_n4507) & (n_n4509)) + ((!n_n4504) & (!n_n4503) & (n_n4507) & (!n_n4509)) + ((!n_n4504) & (!n_n4503) & (n_n4507) & (n_n4509)) + ((!n_n4504) & (n_n4503) & (!n_n4507) & (!n_n4509)) + ((!n_n4504) & (n_n4503) & (!n_n4507) & (n_n4509)) + ((!n_n4504) & (n_n4503) & (n_n4507) & (!n_n4509)) + ((!n_n4504) & (n_n4503) & (n_n4507) & (n_n4509)) + ((n_n4504) & (!n_n4503) & (!n_n4507) & (!n_n4509)) + ((n_n4504) & (!n_n4503) & (!n_n4507) & (n_n4509)) + ((n_n4504) & (!n_n4503) & (n_n4507) & (!n_n4509)) + ((n_n4504) & (!n_n4503) & (n_n4507) & (n_n4509)) + ((n_n4504) & (n_n4503) & (!n_n4507) & (!n_n4509)) + ((n_n4504) & (n_n4503) & (!n_n4507) & (n_n4509)) + ((n_n4504) & (n_n4503) & (n_n4507) & (!n_n4509)) + ((n_n4504) & (n_n4503) & (n_n4507) & (n_n4509)));
	assign x12514x = (((!n_n4511) & (!n_n4499) & (!n_n4505) & (!n_n4510) & (n_n4501)) + ((!n_n4511) & (!n_n4499) & (!n_n4505) & (n_n4510) & (!n_n4501)) + ((!n_n4511) & (!n_n4499) & (!n_n4505) & (n_n4510) & (n_n4501)) + ((!n_n4511) & (!n_n4499) & (n_n4505) & (!n_n4510) & (!n_n4501)) + ((!n_n4511) & (!n_n4499) & (n_n4505) & (!n_n4510) & (n_n4501)) + ((!n_n4511) & (!n_n4499) & (n_n4505) & (n_n4510) & (!n_n4501)) + ((!n_n4511) & (!n_n4499) & (n_n4505) & (n_n4510) & (n_n4501)) + ((!n_n4511) & (n_n4499) & (!n_n4505) & (!n_n4510) & (!n_n4501)) + ((!n_n4511) & (n_n4499) & (!n_n4505) & (!n_n4510) & (n_n4501)) + ((!n_n4511) & (n_n4499) & (!n_n4505) & (n_n4510) & (!n_n4501)) + ((!n_n4511) & (n_n4499) & (!n_n4505) & (n_n4510) & (n_n4501)) + ((!n_n4511) & (n_n4499) & (n_n4505) & (!n_n4510) & (!n_n4501)) + ((!n_n4511) & (n_n4499) & (n_n4505) & (!n_n4510) & (n_n4501)) + ((!n_n4511) & (n_n4499) & (n_n4505) & (n_n4510) & (!n_n4501)) + ((!n_n4511) & (n_n4499) & (n_n4505) & (n_n4510) & (n_n4501)) + ((n_n4511) & (!n_n4499) & (!n_n4505) & (!n_n4510) & (!n_n4501)) + ((n_n4511) & (!n_n4499) & (!n_n4505) & (!n_n4510) & (n_n4501)) + ((n_n4511) & (!n_n4499) & (!n_n4505) & (n_n4510) & (!n_n4501)) + ((n_n4511) & (!n_n4499) & (!n_n4505) & (n_n4510) & (n_n4501)) + ((n_n4511) & (!n_n4499) & (n_n4505) & (!n_n4510) & (!n_n4501)) + ((n_n4511) & (!n_n4499) & (n_n4505) & (!n_n4510) & (n_n4501)) + ((n_n4511) & (!n_n4499) & (n_n4505) & (n_n4510) & (!n_n4501)) + ((n_n4511) & (!n_n4499) & (n_n4505) & (n_n4510) & (n_n4501)) + ((n_n4511) & (n_n4499) & (!n_n4505) & (!n_n4510) & (!n_n4501)) + ((n_n4511) & (n_n4499) & (!n_n4505) & (!n_n4510) & (n_n4501)) + ((n_n4511) & (n_n4499) & (!n_n4505) & (n_n4510) & (!n_n4501)) + ((n_n4511) & (n_n4499) & (!n_n4505) & (n_n4510) & (n_n4501)) + ((n_n4511) & (n_n4499) & (n_n4505) & (!n_n4510) & (!n_n4501)) + ((n_n4511) & (n_n4499) & (n_n4505) & (!n_n4510) & (n_n4501)) + ((n_n4511) & (n_n4499) & (n_n4505) & (n_n4510) & (!n_n4501)) + ((n_n4511) & (n_n4499) & (n_n4505) & (n_n4510) & (n_n4501)));
	assign x22140x = (((!n_n4497) & (!x428x) & (!x66x) & (!n_n4493) & (!n_n1677)));
	assign x12415x = (((!x241x) & (!n_n4715) & (!n_n4716) & (n_n4713)) + ((!x241x) & (!n_n4715) & (n_n4716) & (!n_n4713)) + ((!x241x) & (!n_n4715) & (n_n4716) & (n_n4713)) + ((!x241x) & (n_n4715) & (!n_n4716) & (!n_n4713)) + ((!x241x) & (n_n4715) & (!n_n4716) & (n_n4713)) + ((!x241x) & (n_n4715) & (n_n4716) & (!n_n4713)) + ((!x241x) & (n_n4715) & (n_n4716) & (n_n4713)) + ((x241x) & (!n_n4715) & (!n_n4716) & (!n_n4713)) + ((x241x) & (!n_n4715) & (!n_n4716) & (n_n4713)) + ((x241x) & (!n_n4715) & (n_n4716) & (!n_n4713)) + ((x241x) & (!n_n4715) & (n_n4716) & (n_n4713)) + ((x241x) & (n_n4715) & (!n_n4716) & (!n_n4713)) + ((x241x) & (n_n4715) & (!n_n4716) & (n_n4713)) + ((x241x) & (n_n4715) & (n_n4716) & (!n_n4713)) + ((x241x) & (n_n4715) & (n_n4716) & (n_n4713)));
	assign x12416x = (((!n_n4704) & (!n_n4711) & (!x30x) & (x12415x)) + ((!n_n4704) & (!n_n4711) & (x30x) & (!x12415x)) + ((!n_n4704) & (!n_n4711) & (x30x) & (x12415x)) + ((!n_n4704) & (n_n4711) & (!x30x) & (!x12415x)) + ((!n_n4704) & (n_n4711) & (!x30x) & (x12415x)) + ((!n_n4704) & (n_n4711) & (x30x) & (!x12415x)) + ((!n_n4704) & (n_n4711) & (x30x) & (x12415x)) + ((n_n4704) & (!n_n4711) & (!x30x) & (!x12415x)) + ((n_n4704) & (!n_n4711) & (!x30x) & (x12415x)) + ((n_n4704) & (!n_n4711) & (x30x) & (!x12415x)) + ((n_n4704) & (!n_n4711) & (x30x) & (x12415x)) + ((n_n4704) & (n_n4711) & (!x30x) & (!x12415x)) + ((n_n4704) & (n_n4711) & (!x30x) & (x12415x)) + ((n_n4704) & (n_n4711) & (x30x) & (!x12415x)) + ((n_n4704) & (n_n4711) & (x30x) & (x12415x)));
	assign x12404x = (((!x25x) & (!x11x) & (!n_n325) & (!n_n535) & (x221x)) + ((!x25x) & (!x11x) & (!n_n325) & (n_n535) & (x221x)) + ((!x25x) & (!x11x) & (n_n325) & (!n_n535) & (x221x)) + ((!x25x) & (!x11x) & (n_n325) & (n_n535) & (x221x)) + ((!x25x) & (x11x) & (!n_n325) & (!n_n535) & (x221x)) + ((!x25x) & (x11x) & (!n_n325) & (n_n535) & (x221x)) + ((!x25x) & (x11x) & (n_n325) & (!n_n535) & (x221x)) + ((!x25x) & (x11x) & (n_n325) & (n_n535) & (!x221x)) + ((!x25x) & (x11x) & (n_n325) & (n_n535) & (x221x)) + ((x25x) & (!x11x) & (!n_n325) & (!n_n535) & (x221x)) + ((x25x) & (!x11x) & (!n_n325) & (n_n535) & (x221x)) + ((x25x) & (!x11x) & (n_n325) & (!n_n535) & (x221x)) + ((x25x) & (!x11x) & (n_n325) & (n_n535) & (!x221x)) + ((x25x) & (!x11x) & (n_n325) & (n_n535) & (x221x)) + ((x25x) & (x11x) & (!n_n325) & (!n_n535) & (x221x)) + ((x25x) & (x11x) & (!n_n325) & (n_n535) & (x221x)) + ((x25x) & (x11x) & (n_n325) & (!n_n535) & (x221x)) + ((x25x) & (x11x) & (n_n325) & (n_n535) & (!x221x)) + ((x25x) & (x11x) & (n_n325) & (n_n535) & (x221x)));
	assign x12405x = (((!n_n4701) & (!n_n4696) & (!n_n4695) & (!n_n4702) & (n_n4700)) + ((!n_n4701) & (!n_n4696) & (!n_n4695) & (n_n4702) & (!n_n4700)) + ((!n_n4701) & (!n_n4696) & (!n_n4695) & (n_n4702) & (n_n4700)) + ((!n_n4701) & (!n_n4696) & (n_n4695) & (!n_n4702) & (!n_n4700)) + ((!n_n4701) & (!n_n4696) & (n_n4695) & (!n_n4702) & (n_n4700)) + ((!n_n4701) & (!n_n4696) & (n_n4695) & (n_n4702) & (!n_n4700)) + ((!n_n4701) & (!n_n4696) & (n_n4695) & (n_n4702) & (n_n4700)) + ((!n_n4701) & (n_n4696) & (!n_n4695) & (!n_n4702) & (!n_n4700)) + ((!n_n4701) & (n_n4696) & (!n_n4695) & (!n_n4702) & (n_n4700)) + ((!n_n4701) & (n_n4696) & (!n_n4695) & (n_n4702) & (!n_n4700)) + ((!n_n4701) & (n_n4696) & (!n_n4695) & (n_n4702) & (n_n4700)) + ((!n_n4701) & (n_n4696) & (n_n4695) & (!n_n4702) & (!n_n4700)) + ((!n_n4701) & (n_n4696) & (n_n4695) & (!n_n4702) & (n_n4700)) + ((!n_n4701) & (n_n4696) & (n_n4695) & (n_n4702) & (!n_n4700)) + ((!n_n4701) & (n_n4696) & (n_n4695) & (n_n4702) & (n_n4700)) + ((n_n4701) & (!n_n4696) & (!n_n4695) & (!n_n4702) & (!n_n4700)) + ((n_n4701) & (!n_n4696) & (!n_n4695) & (!n_n4702) & (n_n4700)) + ((n_n4701) & (!n_n4696) & (!n_n4695) & (n_n4702) & (!n_n4700)) + ((n_n4701) & (!n_n4696) & (!n_n4695) & (n_n4702) & (n_n4700)) + ((n_n4701) & (!n_n4696) & (n_n4695) & (!n_n4702) & (!n_n4700)) + ((n_n4701) & (!n_n4696) & (n_n4695) & (!n_n4702) & (n_n4700)) + ((n_n4701) & (!n_n4696) & (n_n4695) & (n_n4702) & (!n_n4700)) + ((n_n4701) & (!n_n4696) & (n_n4695) & (n_n4702) & (n_n4700)) + ((n_n4701) & (n_n4696) & (!n_n4695) & (!n_n4702) & (!n_n4700)) + ((n_n4701) & (n_n4696) & (!n_n4695) & (!n_n4702) & (n_n4700)) + ((n_n4701) & (n_n4696) & (!n_n4695) & (n_n4702) & (!n_n4700)) + ((n_n4701) & (n_n4696) & (!n_n4695) & (n_n4702) & (n_n4700)) + ((n_n4701) & (n_n4696) & (n_n4695) & (!n_n4702) & (!n_n4700)) + ((n_n4701) & (n_n4696) & (n_n4695) & (!n_n4702) & (n_n4700)) + ((n_n4701) & (n_n4696) & (n_n4695) & (n_n4702) & (!n_n4700)) + ((n_n4701) & (n_n4696) & (n_n4695) & (n_n4702) & (n_n4700)));
	assign n_n1476 = (((!x25x) & (!x483x) & (!n_n4727) & (!x242x) & (x12410x)) + ((!x25x) & (!x483x) & (!n_n4727) & (x242x) & (!x12410x)) + ((!x25x) & (!x483x) & (!n_n4727) & (x242x) & (x12410x)) + ((!x25x) & (!x483x) & (n_n4727) & (!x242x) & (!x12410x)) + ((!x25x) & (!x483x) & (n_n4727) & (!x242x) & (x12410x)) + ((!x25x) & (!x483x) & (n_n4727) & (x242x) & (!x12410x)) + ((!x25x) & (!x483x) & (n_n4727) & (x242x) & (x12410x)) + ((!x25x) & (x483x) & (!n_n4727) & (!x242x) & (x12410x)) + ((!x25x) & (x483x) & (!n_n4727) & (x242x) & (!x12410x)) + ((!x25x) & (x483x) & (!n_n4727) & (x242x) & (x12410x)) + ((!x25x) & (x483x) & (n_n4727) & (!x242x) & (!x12410x)) + ((!x25x) & (x483x) & (n_n4727) & (!x242x) & (x12410x)) + ((!x25x) & (x483x) & (n_n4727) & (x242x) & (!x12410x)) + ((!x25x) & (x483x) & (n_n4727) & (x242x) & (x12410x)) + ((x25x) & (!x483x) & (!n_n4727) & (!x242x) & (x12410x)) + ((x25x) & (!x483x) & (!n_n4727) & (x242x) & (!x12410x)) + ((x25x) & (!x483x) & (!n_n4727) & (x242x) & (x12410x)) + ((x25x) & (!x483x) & (n_n4727) & (!x242x) & (!x12410x)) + ((x25x) & (!x483x) & (n_n4727) & (!x242x) & (x12410x)) + ((x25x) & (!x483x) & (n_n4727) & (x242x) & (!x12410x)) + ((x25x) & (!x483x) & (n_n4727) & (x242x) & (x12410x)) + ((x25x) & (x483x) & (!n_n4727) & (!x242x) & (!x12410x)) + ((x25x) & (x483x) & (!n_n4727) & (!x242x) & (x12410x)) + ((x25x) & (x483x) & (!n_n4727) & (x242x) & (!x12410x)) + ((x25x) & (x483x) & (!n_n4727) & (x242x) & (x12410x)) + ((x25x) & (x483x) & (n_n4727) & (!x242x) & (!x12410x)) + ((x25x) & (x483x) & (n_n4727) & (!x242x) & (x12410x)) + ((x25x) & (x483x) & (n_n4727) & (x242x) & (!x12410x)) + ((x25x) & (x483x) & (n_n4727) & (x242x) & (x12410x)));
	assign x22206x = (((!n_n4690) & (!n_n4688) & (!n_n4685) & (!n_n4687) & (!n_n3848)));
	assign x13351x = (((!i_7_) & (!i_8_) & (!i_6_) & (x19x) & (n_n518)) + ((!i_7_) & (!i_8_) & (i_6_) & (x19x) & (n_n518)));
	assign x13353x = (((!n_n518) & (!x11x) & (!n_n65) & (!n_n5232) & (n_n5233)) + ((!n_n518) & (!x11x) & (!n_n65) & (n_n5232) & (!n_n5233)) + ((!n_n518) & (!x11x) & (!n_n65) & (n_n5232) & (n_n5233)) + ((!n_n518) & (!x11x) & (n_n65) & (!n_n5232) & (n_n5233)) + ((!n_n518) & (!x11x) & (n_n65) & (n_n5232) & (!n_n5233)) + ((!n_n518) & (!x11x) & (n_n65) & (n_n5232) & (n_n5233)) + ((!n_n518) & (x11x) & (!n_n65) & (!n_n5232) & (n_n5233)) + ((!n_n518) & (x11x) & (!n_n65) & (n_n5232) & (!n_n5233)) + ((!n_n518) & (x11x) & (!n_n65) & (n_n5232) & (n_n5233)) + ((!n_n518) & (x11x) & (n_n65) & (!n_n5232) & (n_n5233)) + ((!n_n518) & (x11x) & (n_n65) & (n_n5232) & (!n_n5233)) + ((!n_n518) & (x11x) & (n_n65) & (n_n5232) & (n_n5233)) + ((n_n518) & (!x11x) & (!n_n65) & (!n_n5232) & (n_n5233)) + ((n_n518) & (!x11x) & (!n_n65) & (n_n5232) & (!n_n5233)) + ((n_n518) & (!x11x) & (!n_n65) & (n_n5232) & (n_n5233)) + ((n_n518) & (!x11x) & (n_n65) & (!n_n5232) & (n_n5233)) + ((n_n518) & (!x11x) & (n_n65) & (n_n5232) & (!n_n5233)) + ((n_n518) & (!x11x) & (n_n65) & (n_n5232) & (n_n5233)) + ((n_n518) & (x11x) & (!n_n65) & (!n_n5232) & (n_n5233)) + ((n_n518) & (x11x) & (!n_n65) & (n_n5232) & (!n_n5233)) + ((n_n518) & (x11x) & (!n_n65) & (n_n5232) & (n_n5233)) + ((n_n518) & (x11x) & (n_n65) & (!n_n5232) & (!n_n5233)) + ((n_n518) & (x11x) & (n_n65) & (!n_n5232) & (n_n5233)) + ((n_n518) & (x11x) & (n_n65) & (n_n5232) & (!n_n5233)) + ((n_n518) & (x11x) & (n_n65) & (n_n5232) & (n_n5233)));
	assign x13027x = (((!i_9_) & (n_n526) & (n_n455) & (n_n500)) + ((i_9_) & (n_n526) & (n_n455) & (n_n500)));
	assign x22137x = (((!x492x) & (!x10x) & (!n_n4648) & (!n_n4646) & (!n_n4650)) + ((!x492x) & (x10x) & (!n_n4648) & (!n_n4646) & (!n_n4650)) + ((x492x) & (!x10x) & (!n_n4648) & (!n_n4646) & (!n_n4650)));
	assign n_n1482 = (((!x311x) & (!n_n4656) & (!n_n4654) & (!n_n4657) & (!x22137x)) + ((!x311x) & (!n_n4656) & (!n_n4654) & (n_n4657) & (!x22137x)) + ((!x311x) & (!n_n4656) & (!n_n4654) & (n_n4657) & (x22137x)) + ((!x311x) & (!n_n4656) & (n_n4654) & (!n_n4657) & (!x22137x)) + ((!x311x) & (!n_n4656) & (n_n4654) & (!n_n4657) & (x22137x)) + ((!x311x) & (!n_n4656) & (n_n4654) & (n_n4657) & (!x22137x)) + ((!x311x) & (!n_n4656) & (n_n4654) & (n_n4657) & (x22137x)) + ((!x311x) & (n_n4656) & (!n_n4654) & (!n_n4657) & (!x22137x)) + ((!x311x) & (n_n4656) & (!n_n4654) & (!n_n4657) & (x22137x)) + ((!x311x) & (n_n4656) & (!n_n4654) & (n_n4657) & (!x22137x)) + ((!x311x) & (n_n4656) & (!n_n4654) & (n_n4657) & (x22137x)) + ((!x311x) & (n_n4656) & (n_n4654) & (!n_n4657) & (!x22137x)) + ((!x311x) & (n_n4656) & (n_n4654) & (!n_n4657) & (x22137x)) + ((!x311x) & (n_n4656) & (n_n4654) & (n_n4657) & (!x22137x)) + ((!x311x) & (n_n4656) & (n_n4654) & (n_n4657) & (x22137x)) + ((x311x) & (!n_n4656) & (!n_n4654) & (!n_n4657) & (!x22137x)) + ((x311x) & (!n_n4656) & (!n_n4654) & (!n_n4657) & (x22137x)) + ((x311x) & (!n_n4656) & (!n_n4654) & (n_n4657) & (!x22137x)) + ((x311x) & (!n_n4656) & (!n_n4654) & (n_n4657) & (x22137x)) + ((x311x) & (!n_n4656) & (n_n4654) & (!n_n4657) & (!x22137x)) + ((x311x) & (!n_n4656) & (n_n4654) & (!n_n4657) & (x22137x)) + ((x311x) & (!n_n4656) & (n_n4654) & (n_n4657) & (!x22137x)) + ((x311x) & (!n_n4656) & (n_n4654) & (n_n4657) & (x22137x)) + ((x311x) & (n_n4656) & (!n_n4654) & (!n_n4657) & (!x22137x)) + ((x311x) & (n_n4656) & (!n_n4654) & (!n_n4657) & (x22137x)) + ((x311x) & (n_n4656) & (!n_n4654) & (n_n4657) & (!x22137x)) + ((x311x) & (n_n4656) & (!n_n4654) & (n_n4657) & (x22137x)) + ((x311x) & (n_n4656) & (n_n4654) & (!n_n4657) & (!x22137x)) + ((x311x) & (n_n4656) & (n_n4654) & (!n_n4657) & (x22137x)) + ((x311x) & (n_n4656) & (n_n4654) & (n_n4657) & (!x22137x)) + ((x311x) & (n_n4656) & (n_n4654) & (n_n4657) & (x22137x)));
	assign x270x = (((!i_9_) & (n_n390) & (n_n532) & (!n_n534) & (n_n500)) + ((!i_9_) & (n_n390) & (n_n532) & (n_n534) & (n_n500)) + ((i_9_) & (n_n390) & (!n_n532) & (n_n534) & (n_n500)) + ((i_9_) & (n_n390) & (n_n532) & (n_n534) & (n_n500)));
	assign x22138x = (((!n_n4612) & (!n_n4608) & (!n_n4611) & (!n_n4620)));
	assign n_n1485 = (((!n_n4615) & (!n_n4609) & (!n_n4614) & (!x270x) & (!x22138x)) + ((!n_n4615) & (!n_n4609) & (!n_n4614) & (x270x) & (!x22138x)) + ((!n_n4615) & (!n_n4609) & (!n_n4614) & (x270x) & (x22138x)) + ((!n_n4615) & (!n_n4609) & (n_n4614) & (!x270x) & (!x22138x)) + ((!n_n4615) & (!n_n4609) & (n_n4614) & (!x270x) & (x22138x)) + ((!n_n4615) & (!n_n4609) & (n_n4614) & (x270x) & (!x22138x)) + ((!n_n4615) & (!n_n4609) & (n_n4614) & (x270x) & (x22138x)) + ((!n_n4615) & (n_n4609) & (!n_n4614) & (!x270x) & (!x22138x)) + ((!n_n4615) & (n_n4609) & (!n_n4614) & (!x270x) & (x22138x)) + ((!n_n4615) & (n_n4609) & (!n_n4614) & (x270x) & (!x22138x)) + ((!n_n4615) & (n_n4609) & (!n_n4614) & (x270x) & (x22138x)) + ((!n_n4615) & (n_n4609) & (n_n4614) & (!x270x) & (!x22138x)) + ((!n_n4615) & (n_n4609) & (n_n4614) & (!x270x) & (x22138x)) + ((!n_n4615) & (n_n4609) & (n_n4614) & (x270x) & (!x22138x)) + ((!n_n4615) & (n_n4609) & (n_n4614) & (x270x) & (x22138x)) + ((n_n4615) & (!n_n4609) & (!n_n4614) & (!x270x) & (!x22138x)) + ((n_n4615) & (!n_n4609) & (!n_n4614) & (!x270x) & (x22138x)) + ((n_n4615) & (!n_n4609) & (!n_n4614) & (x270x) & (!x22138x)) + ((n_n4615) & (!n_n4609) & (!n_n4614) & (x270x) & (x22138x)) + ((n_n4615) & (!n_n4609) & (n_n4614) & (!x270x) & (!x22138x)) + ((n_n4615) & (!n_n4609) & (n_n4614) & (!x270x) & (x22138x)) + ((n_n4615) & (!n_n4609) & (n_n4614) & (x270x) & (!x22138x)) + ((n_n4615) & (!n_n4609) & (n_n4614) & (x270x) & (x22138x)) + ((n_n4615) & (n_n4609) & (!n_n4614) & (!x270x) & (!x22138x)) + ((n_n4615) & (n_n4609) & (!n_n4614) & (!x270x) & (x22138x)) + ((n_n4615) & (n_n4609) & (!n_n4614) & (x270x) & (!x22138x)) + ((n_n4615) & (n_n4609) & (!n_n4614) & (x270x) & (x22138x)) + ((n_n4615) & (n_n4609) & (n_n4614) & (!x270x) & (!x22138x)) + ((n_n4615) & (n_n4609) & (n_n4614) & (!x270x) & (x22138x)) + ((n_n4615) & (n_n4609) & (n_n4614) & (x270x) & (!x22138x)) + ((n_n4615) & (n_n4609) & (n_n4614) & (x270x) & (x22138x)));
	assign x22209x = (((!x20x) & (!x583x) & (!n_n4598) & (!n_n4596) & (!n_n4590)) + ((!x20x) & (x583x) & (!n_n4598) & (!n_n4596) & (!n_n4590)) + ((x20x) & (!x583x) & (!n_n4598) & (!n_n4596) & (!n_n4590)));
	assign n_n1487 = (((!n_n4593) & (!n_n4595) & (!n_n4594) & (!x365x) & (!x22209x)) + ((!n_n4593) & (!n_n4595) & (!n_n4594) & (x365x) & (!x22209x)) + ((!n_n4593) & (!n_n4595) & (!n_n4594) & (x365x) & (x22209x)) + ((!n_n4593) & (!n_n4595) & (n_n4594) & (!x365x) & (!x22209x)) + ((!n_n4593) & (!n_n4595) & (n_n4594) & (!x365x) & (x22209x)) + ((!n_n4593) & (!n_n4595) & (n_n4594) & (x365x) & (!x22209x)) + ((!n_n4593) & (!n_n4595) & (n_n4594) & (x365x) & (x22209x)) + ((!n_n4593) & (n_n4595) & (!n_n4594) & (!x365x) & (!x22209x)) + ((!n_n4593) & (n_n4595) & (!n_n4594) & (!x365x) & (x22209x)) + ((!n_n4593) & (n_n4595) & (!n_n4594) & (x365x) & (!x22209x)) + ((!n_n4593) & (n_n4595) & (!n_n4594) & (x365x) & (x22209x)) + ((!n_n4593) & (n_n4595) & (n_n4594) & (!x365x) & (!x22209x)) + ((!n_n4593) & (n_n4595) & (n_n4594) & (!x365x) & (x22209x)) + ((!n_n4593) & (n_n4595) & (n_n4594) & (x365x) & (!x22209x)) + ((!n_n4593) & (n_n4595) & (n_n4594) & (x365x) & (x22209x)) + ((n_n4593) & (!n_n4595) & (!n_n4594) & (!x365x) & (!x22209x)) + ((n_n4593) & (!n_n4595) & (!n_n4594) & (!x365x) & (x22209x)) + ((n_n4593) & (!n_n4595) & (!n_n4594) & (x365x) & (!x22209x)) + ((n_n4593) & (!n_n4595) & (!n_n4594) & (x365x) & (x22209x)) + ((n_n4593) & (!n_n4595) & (n_n4594) & (!x365x) & (!x22209x)) + ((n_n4593) & (!n_n4595) & (n_n4594) & (!x365x) & (x22209x)) + ((n_n4593) & (!n_n4595) & (n_n4594) & (x365x) & (!x22209x)) + ((n_n4593) & (!n_n4595) & (n_n4594) & (x365x) & (x22209x)) + ((n_n4593) & (n_n4595) & (!n_n4594) & (!x365x) & (!x22209x)) + ((n_n4593) & (n_n4595) & (!n_n4594) & (!x365x) & (x22209x)) + ((n_n4593) & (n_n4595) & (!n_n4594) & (x365x) & (!x22209x)) + ((n_n4593) & (n_n4595) & (!n_n4594) & (x365x) & (x22209x)) + ((n_n4593) & (n_n4595) & (n_n4594) & (!x365x) & (!x22209x)) + ((n_n4593) & (n_n4595) & (n_n4594) & (!x365x) & (x22209x)) + ((n_n4593) & (n_n4595) & (n_n4594) & (x365x) & (!x22209x)) + ((n_n4593) & (n_n4595) & (n_n4594) & (x365x) & (x22209x)));
	assign x12559x = (((!n_n1649) & (!n_n4621) & (!n_n4640) & (!n_n1648) & (n_n1646)) + ((!n_n1649) & (!n_n4621) & (!n_n4640) & (n_n1648) & (!n_n1646)) + ((!n_n1649) & (!n_n4621) & (!n_n4640) & (n_n1648) & (n_n1646)) + ((!n_n1649) & (!n_n4621) & (n_n4640) & (!n_n1648) & (!n_n1646)) + ((!n_n1649) & (!n_n4621) & (n_n4640) & (!n_n1648) & (n_n1646)) + ((!n_n1649) & (!n_n4621) & (n_n4640) & (n_n1648) & (!n_n1646)) + ((!n_n1649) & (!n_n4621) & (n_n4640) & (n_n1648) & (n_n1646)) + ((!n_n1649) & (n_n4621) & (!n_n4640) & (!n_n1648) & (!n_n1646)) + ((!n_n1649) & (n_n4621) & (!n_n4640) & (!n_n1648) & (n_n1646)) + ((!n_n1649) & (n_n4621) & (!n_n4640) & (n_n1648) & (!n_n1646)) + ((!n_n1649) & (n_n4621) & (!n_n4640) & (n_n1648) & (n_n1646)) + ((!n_n1649) & (n_n4621) & (n_n4640) & (!n_n1648) & (!n_n1646)) + ((!n_n1649) & (n_n4621) & (n_n4640) & (!n_n1648) & (n_n1646)) + ((!n_n1649) & (n_n4621) & (n_n4640) & (n_n1648) & (!n_n1646)) + ((!n_n1649) & (n_n4621) & (n_n4640) & (n_n1648) & (n_n1646)) + ((n_n1649) & (!n_n4621) & (!n_n4640) & (!n_n1648) & (!n_n1646)) + ((n_n1649) & (!n_n4621) & (!n_n4640) & (!n_n1648) & (n_n1646)) + ((n_n1649) & (!n_n4621) & (!n_n4640) & (n_n1648) & (!n_n1646)) + ((n_n1649) & (!n_n4621) & (!n_n4640) & (n_n1648) & (n_n1646)) + ((n_n1649) & (!n_n4621) & (n_n4640) & (!n_n1648) & (!n_n1646)) + ((n_n1649) & (!n_n4621) & (n_n4640) & (!n_n1648) & (n_n1646)) + ((n_n1649) & (!n_n4621) & (n_n4640) & (n_n1648) & (!n_n1646)) + ((n_n1649) & (!n_n4621) & (n_n4640) & (n_n1648) & (n_n1646)) + ((n_n1649) & (n_n4621) & (!n_n4640) & (!n_n1648) & (!n_n1646)) + ((n_n1649) & (n_n4621) & (!n_n4640) & (!n_n1648) & (n_n1646)) + ((n_n1649) & (n_n4621) & (!n_n4640) & (n_n1648) & (!n_n1646)) + ((n_n1649) & (n_n4621) & (!n_n4640) & (n_n1648) & (n_n1646)) + ((n_n1649) & (n_n4621) & (n_n4640) & (!n_n1648) & (!n_n1646)) + ((n_n1649) & (n_n4621) & (n_n4640) & (!n_n1648) & (n_n1646)) + ((n_n1649) & (n_n4621) & (n_n4640) & (n_n1648) & (!n_n1646)) + ((n_n1649) & (n_n4621) & (n_n4640) & (n_n1648) & (n_n1646)));
	assign x12558x = (((!n_n4641) & (!n_n4643) & (!x349x) & (!n_n4630) & (x401x)) + ((!n_n4641) & (!n_n4643) & (!x349x) & (n_n4630) & (!x401x)) + ((!n_n4641) & (!n_n4643) & (!x349x) & (n_n4630) & (x401x)) + ((!n_n4641) & (!n_n4643) & (x349x) & (!n_n4630) & (!x401x)) + ((!n_n4641) & (!n_n4643) & (x349x) & (!n_n4630) & (x401x)) + ((!n_n4641) & (!n_n4643) & (x349x) & (n_n4630) & (!x401x)) + ((!n_n4641) & (!n_n4643) & (x349x) & (n_n4630) & (x401x)) + ((!n_n4641) & (n_n4643) & (!x349x) & (!n_n4630) & (!x401x)) + ((!n_n4641) & (n_n4643) & (!x349x) & (!n_n4630) & (x401x)) + ((!n_n4641) & (n_n4643) & (!x349x) & (n_n4630) & (!x401x)) + ((!n_n4641) & (n_n4643) & (!x349x) & (n_n4630) & (x401x)) + ((!n_n4641) & (n_n4643) & (x349x) & (!n_n4630) & (!x401x)) + ((!n_n4641) & (n_n4643) & (x349x) & (!n_n4630) & (x401x)) + ((!n_n4641) & (n_n4643) & (x349x) & (n_n4630) & (!x401x)) + ((!n_n4641) & (n_n4643) & (x349x) & (n_n4630) & (x401x)) + ((n_n4641) & (!n_n4643) & (!x349x) & (!n_n4630) & (!x401x)) + ((n_n4641) & (!n_n4643) & (!x349x) & (!n_n4630) & (x401x)) + ((n_n4641) & (!n_n4643) & (!x349x) & (n_n4630) & (!x401x)) + ((n_n4641) & (!n_n4643) & (!x349x) & (n_n4630) & (x401x)) + ((n_n4641) & (!n_n4643) & (x349x) & (!n_n4630) & (!x401x)) + ((n_n4641) & (!n_n4643) & (x349x) & (!n_n4630) & (x401x)) + ((n_n4641) & (!n_n4643) & (x349x) & (n_n4630) & (!x401x)) + ((n_n4641) & (!n_n4643) & (x349x) & (n_n4630) & (x401x)) + ((n_n4641) & (n_n4643) & (!x349x) & (!n_n4630) & (!x401x)) + ((n_n4641) & (n_n4643) & (!x349x) & (!n_n4630) & (x401x)) + ((n_n4641) & (n_n4643) & (!x349x) & (n_n4630) & (!x401x)) + ((n_n4641) & (n_n4643) & (!x349x) & (n_n4630) & (x401x)) + ((n_n4641) & (n_n4643) & (x349x) & (!n_n4630) & (!x401x)) + ((n_n4641) & (n_n4643) & (x349x) & (!n_n4630) & (x401x)) + ((n_n4641) & (n_n4643) & (x349x) & (n_n4630) & (!x401x)) + ((n_n4641) & (n_n4643) & (x349x) & (n_n4630) & (x401x)));
	assign n_n1420 = (((!n_n1482) & (!x12559x) & (x12558x)) + ((!n_n1482) & (x12559x) & (!x12558x)) + ((!n_n1482) & (x12559x) & (x12558x)) + ((n_n1482) & (!x12559x) & (!x12558x)) + ((n_n1482) & (!x12559x) & (x12558x)) + ((n_n1482) & (x12559x) & (!x12558x)) + ((n_n1482) & (x12559x) & (x12558x)));
	assign x12565x = (((!n_n4603) & (!x256x) & (!n_n2036) & (!x22170x)) + ((!n_n4603) & (!x256x) & (n_n2036) & (!x22170x)) + ((!n_n4603) & (!x256x) & (n_n2036) & (x22170x)) + ((!n_n4603) & (x256x) & (!n_n2036) & (!x22170x)) + ((!n_n4603) & (x256x) & (!n_n2036) & (x22170x)) + ((!n_n4603) & (x256x) & (n_n2036) & (!x22170x)) + ((!n_n4603) & (x256x) & (n_n2036) & (x22170x)) + ((n_n4603) & (!x256x) & (!n_n2036) & (!x22170x)) + ((n_n4603) & (!x256x) & (!n_n2036) & (x22170x)) + ((n_n4603) & (!x256x) & (n_n2036) & (!x22170x)) + ((n_n4603) & (!x256x) & (n_n2036) & (x22170x)) + ((n_n4603) & (x256x) & (!n_n2036) & (!x22170x)) + ((n_n4603) & (x256x) & (!n_n2036) & (x22170x)) + ((n_n4603) & (x256x) & (n_n2036) & (!x22170x)) + ((n_n4603) & (x256x) & (n_n2036) & (x22170x)));
	assign n_n1703 = (((!i_9_) & (n_n536) & (n_n524) & (n_n535) & (!n_n522)) + ((!i_9_) & (n_n536) & (n_n524) & (n_n535) & (n_n522)) + ((i_9_) & (n_n536) & (!n_n524) & (n_n535) & (n_n522)) + ((i_9_) & (n_n536) & (n_n524) & (n_n535) & (!n_n522)) + ((i_9_) & (n_n536) & (n_n524) & (n_n535) & (n_n522)));
	assign x448x = (((!i_9_) & (n_n536) & (n_n518) & (!n_n526) & (n_n528)) + ((!i_9_) & (n_n536) & (n_n518) & (n_n526) & (!n_n528)) + ((!i_9_) & (n_n536) & (n_n518) & (n_n526) & (n_n528)) + ((i_9_) & (n_n536) & (n_n518) & (n_n526) & (!n_n528)) + ((i_9_) & (n_n536) & (n_n518) & (n_n526) & (n_n528)));
	assign x12575x = (((!x25x) & (!n_n536) & (!x11x) & (!n_n535) & (n_n4321)) + ((!x25x) & (!n_n536) & (!x11x) & (n_n535) & (n_n4321)) + ((!x25x) & (!n_n536) & (x11x) & (!n_n535) & (n_n4321)) + ((!x25x) & (!n_n536) & (x11x) & (n_n535) & (n_n4321)) + ((!x25x) & (n_n536) & (!x11x) & (!n_n535) & (n_n4321)) + ((!x25x) & (n_n536) & (!x11x) & (n_n535) & (n_n4321)) + ((!x25x) & (n_n536) & (x11x) & (!n_n535) & (n_n4321)) + ((!x25x) & (n_n536) & (x11x) & (n_n535) & (!n_n4321)) + ((!x25x) & (n_n536) & (x11x) & (n_n535) & (n_n4321)) + ((x25x) & (!n_n536) & (!x11x) & (!n_n535) & (n_n4321)) + ((x25x) & (!n_n536) & (!x11x) & (n_n535) & (n_n4321)) + ((x25x) & (!n_n536) & (x11x) & (!n_n535) & (n_n4321)) + ((x25x) & (!n_n536) & (x11x) & (n_n535) & (n_n4321)) + ((x25x) & (n_n536) & (!x11x) & (!n_n535) & (n_n4321)) + ((x25x) & (n_n536) & (!x11x) & (n_n535) & (!n_n4321)) + ((x25x) & (n_n536) & (!x11x) & (n_n535) & (n_n4321)) + ((x25x) & (n_n536) & (x11x) & (!n_n535) & (n_n4321)) + ((x25x) & (n_n536) & (x11x) & (n_n535) & (!n_n4321)) + ((x25x) & (n_n536) & (x11x) & (n_n535) & (n_n4321)));
	assign x15837x = (((!n_n4473) & (!n_n4497) & (!n_n4474) & (!n_n4486) & (x617x)) + ((!n_n4473) & (!n_n4497) & (!n_n4474) & (n_n4486) & (!x617x)) + ((!n_n4473) & (!n_n4497) & (!n_n4474) & (n_n4486) & (x617x)) + ((!n_n4473) & (!n_n4497) & (n_n4474) & (!n_n4486) & (!x617x)) + ((!n_n4473) & (!n_n4497) & (n_n4474) & (!n_n4486) & (x617x)) + ((!n_n4473) & (!n_n4497) & (n_n4474) & (n_n4486) & (!x617x)) + ((!n_n4473) & (!n_n4497) & (n_n4474) & (n_n4486) & (x617x)) + ((!n_n4473) & (n_n4497) & (!n_n4474) & (!n_n4486) & (!x617x)) + ((!n_n4473) & (n_n4497) & (!n_n4474) & (!n_n4486) & (x617x)) + ((!n_n4473) & (n_n4497) & (!n_n4474) & (n_n4486) & (!x617x)) + ((!n_n4473) & (n_n4497) & (!n_n4474) & (n_n4486) & (x617x)) + ((!n_n4473) & (n_n4497) & (n_n4474) & (!n_n4486) & (!x617x)) + ((!n_n4473) & (n_n4497) & (n_n4474) & (!n_n4486) & (x617x)) + ((!n_n4473) & (n_n4497) & (n_n4474) & (n_n4486) & (!x617x)) + ((!n_n4473) & (n_n4497) & (n_n4474) & (n_n4486) & (x617x)) + ((n_n4473) & (!n_n4497) & (!n_n4474) & (!n_n4486) & (!x617x)) + ((n_n4473) & (!n_n4497) & (!n_n4474) & (!n_n4486) & (x617x)) + ((n_n4473) & (!n_n4497) & (!n_n4474) & (n_n4486) & (!x617x)) + ((n_n4473) & (!n_n4497) & (!n_n4474) & (n_n4486) & (x617x)) + ((n_n4473) & (!n_n4497) & (n_n4474) & (!n_n4486) & (!x617x)) + ((n_n4473) & (!n_n4497) & (n_n4474) & (!n_n4486) & (x617x)) + ((n_n4473) & (!n_n4497) & (n_n4474) & (n_n4486) & (!x617x)) + ((n_n4473) & (!n_n4497) & (n_n4474) & (n_n4486) & (x617x)) + ((n_n4473) & (n_n4497) & (!n_n4474) & (!n_n4486) & (!x617x)) + ((n_n4473) & (n_n4497) & (!n_n4474) & (!n_n4486) & (x617x)) + ((n_n4473) & (n_n4497) & (!n_n4474) & (n_n4486) & (!x617x)) + ((n_n4473) & (n_n4497) & (!n_n4474) & (n_n4486) & (x617x)) + ((n_n4473) & (n_n4497) & (n_n4474) & (!n_n4486) & (!x617x)) + ((n_n4473) & (n_n4497) & (n_n4474) & (!n_n4486) & (x617x)) + ((n_n4473) & (n_n4497) & (n_n4474) & (n_n4486) & (!x617x)) + ((n_n4473) & (n_n4497) & (n_n4474) & (n_n4486) & (x617x)));
	assign x15838x = (((!n_n4471) & (!n_n4478) & (!n_n4502) & (!n_n4509) & (x15837x)) + ((!n_n4471) & (!n_n4478) & (!n_n4502) & (n_n4509) & (!x15837x)) + ((!n_n4471) & (!n_n4478) & (!n_n4502) & (n_n4509) & (x15837x)) + ((!n_n4471) & (!n_n4478) & (n_n4502) & (!n_n4509) & (!x15837x)) + ((!n_n4471) & (!n_n4478) & (n_n4502) & (!n_n4509) & (x15837x)) + ((!n_n4471) & (!n_n4478) & (n_n4502) & (n_n4509) & (!x15837x)) + ((!n_n4471) & (!n_n4478) & (n_n4502) & (n_n4509) & (x15837x)) + ((!n_n4471) & (n_n4478) & (!n_n4502) & (!n_n4509) & (!x15837x)) + ((!n_n4471) & (n_n4478) & (!n_n4502) & (!n_n4509) & (x15837x)) + ((!n_n4471) & (n_n4478) & (!n_n4502) & (n_n4509) & (!x15837x)) + ((!n_n4471) & (n_n4478) & (!n_n4502) & (n_n4509) & (x15837x)) + ((!n_n4471) & (n_n4478) & (n_n4502) & (!n_n4509) & (!x15837x)) + ((!n_n4471) & (n_n4478) & (n_n4502) & (!n_n4509) & (x15837x)) + ((!n_n4471) & (n_n4478) & (n_n4502) & (n_n4509) & (!x15837x)) + ((!n_n4471) & (n_n4478) & (n_n4502) & (n_n4509) & (x15837x)) + ((n_n4471) & (!n_n4478) & (!n_n4502) & (!n_n4509) & (!x15837x)) + ((n_n4471) & (!n_n4478) & (!n_n4502) & (!n_n4509) & (x15837x)) + ((n_n4471) & (!n_n4478) & (!n_n4502) & (n_n4509) & (!x15837x)) + ((n_n4471) & (!n_n4478) & (!n_n4502) & (n_n4509) & (x15837x)) + ((n_n4471) & (!n_n4478) & (n_n4502) & (!n_n4509) & (!x15837x)) + ((n_n4471) & (!n_n4478) & (n_n4502) & (!n_n4509) & (x15837x)) + ((n_n4471) & (!n_n4478) & (n_n4502) & (n_n4509) & (!x15837x)) + ((n_n4471) & (!n_n4478) & (n_n4502) & (n_n4509) & (x15837x)) + ((n_n4471) & (n_n4478) & (!n_n4502) & (!n_n4509) & (!x15837x)) + ((n_n4471) & (n_n4478) & (!n_n4502) & (!n_n4509) & (x15837x)) + ((n_n4471) & (n_n4478) & (!n_n4502) & (n_n4509) & (!x15837x)) + ((n_n4471) & (n_n4478) & (!n_n4502) & (n_n4509) & (x15837x)) + ((n_n4471) & (n_n4478) & (n_n4502) & (!n_n4509) & (!x15837x)) + ((n_n4471) & (n_n4478) & (n_n4502) & (!n_n4509) & (x15837x)) + ((n_n4471) & (n_n4478) & (n_n4502) & (n_n4509) & (!x15837x)) + ((n_n4471) & (n_n4478) & (n_n4502) & (n_n4509) & (x15837x)));
	assign x15823x = (((!n_n4513) & (!n_n4515) & (!n_n4511) & (n_n4590)) + ((!n_n4513) & (!n_n4515) & (n_n4511) & (!n_n4590)) + ((!n_n4513) & (!n_n4515) & (n_n4511) & (n_n4590)) + ((!n_n4513) & (n_n4515) & (!n_n4511) & (!n_n4590)) + ((!n_n4513) & (n_n4515) & (!n_n4511) & (n_n4590)) + ((!n_n4513) & (n_n4515) & (n_n4511) & (!n_n4590)) + ((!n_n4513) & (n_n4515) & (n_n4511) & (n_n4590)) + ((n_n4513) & (!n_n4515) & (!n_n4511) & (!n_n4590)) + ((n_n4513) & (!n_n4515) & (!n_n4511) & (n_n4590)) + ((n_n4513) & (!n_n4515) & (n_n4511) & (!n_n4590)) + ((n_n4513) & (!n_n4515) & (n_n4511) & (n_n4590)) + ((n_n4513) & (n_n4515) & (!n_n4511) & (!n_n4590)) + ((n_n4513) & (n_n4515) & (!n_n4511) & (n_n4590)) + ((n_n4513) & (n_n4515) & (n_n4511) & (!n_n4590)) + ((n_n4513) & (n_n4515) & (n_n4511) & (n_n4590)));
	assign x15824x = (((!n_n4593) & (!n_n4594) & (!n_n4572) & (!n_n4518) & (n_n4552)) + ((!n_n4593) & (!n_n4594) & (!n_n4572) & (n_n4518) & (!n_n4552)) + ((!n_n4593) & (!n_n4594) & (!n_n4572) & (n_n4518) & (n_n4552)) + ((!n_n4593) & (!n_n4594) & (n_n4572) & (!n_n4518) & (!n_n4552)) + ((!n_n4593) & (!n_n4594) & (n_n4572) & (!n_n4518) & (n_n4552)) + ((!n_n4593) & (!n_n4594) & (n_n4572) & (n_n4518) & (!n_n4552)) + ((!n_n4593) & (!n_n4594) & (n_n4572) & (n_n4518) & (n_n4552)) + ((!n_n4593) & (n_n4594) & (!n_n4572) & (!n_n4518) & (!n_n4552)) + ((!n_n4593) & (n_n4594) & (!n_n4572) & (!n_n4518) & (n_n4552)) + ((!n_n4593) & (n_n4594) & (!n_n4572) & (n_n4518) & (!n_n4552)) + ((!n_n4593) & (n_n4594) & (!n_n4572) & (n_n4518) & (n_n4552)) + ((!n_n4593) & (n_n4594) & (n_n4572) & (!n_n4518) & (!n_n4552)) + ((!n_n4593) & (n_n4594) & (n_n4572) & (!n_n4518) & (n_n4552)) + ((!n_n4593) & (n_n4594) & (n_n4572) & (n_n4518) & (!n_n4552)) + ((!n_n4593) & (n_n4594) & (n_n4572) & (n_n4518) & (n_n4552)) + ((n_n4593) & (!n_n4594) & (!n_n4572) & (!n_n4518) & (!n_n4552)) + ((n_n4593) & (!n_n4594) & (!n_n4572) & (!n_n4518) & (n_n4552)) + ((n_n4593) & (!n_n4594) & (!n_n4572) & (n_n4518) & (!n_n4552)) + ((n_n4593) & (!n_n4594) & (!n_n4572) & (n_n4518) & (n_n4552)) + ((n_n4593) & (!n_n4594) & (n_n4572) & (!n_n4518) & (!n_n4552)) + ((n_n4593) & (!n_n4594) & (n_n4572) & (!n_n4518) & (n_n4552)) + ((n_n4593) & (!n_n4594) & (n_n4572) & (n_n4518) & (!n_n4552)) + ((n_n4593) & (!n_n4594) & (n_n4572) & (n_n4518) & (n_n4552)) + ((n_n4593) & (n_n4594) & (!n_n4572) & (!n_n4518) & (!n_n4552)) + ((n_n4593) & (n_n4594) & (!n_n4572) & (!n_n4518) & (n_n4552)) + ((n_n4593) & (n_n4594) & (!n_n4572) & (n_n4518) & (!n_n4552)) + ((n_n4593) & (n_n4594) & (!n_n4572) & (n_n4518) & (n_n4552)) + ((n_n4593) & (n_n4594) & (n_n4572) & (!n_n4518) & (!n_n4552)) + ((n_n4593) & (n_n4594) & (n_n4572) & (!n_n4518) & (n_n4552)) + ((n_n4593) & (n_n4594) & (n_n4572) & (n_n4518) & (!n_n4552)) + ((n_n4593) & (n_n4594) & (n_n4572) & (n_n4518) & (n_n4552)));
	assign x15829x = (((!n_n4641) & (!n_n4648) & (!n_n4651) & (n_n4622)) + ((!n_n4641) & (!n_n4648) & (n_n4651) & (!n_n4622)) + ((!n_n4641) & (!n_n4648) & (n_n4651) & (n_n4622)) + ((!n_n4641) & (n_n4648) & (!n_n4651) & (!n_n4622)) + ((!n_n4641) & (n_n4648) & (!n_n4651) & (n_n4622)) + ((!n_n4641) & (n_n4648) & (n_n4651) & (!n_n4622)) + ((!n_n4641) & (n_n4648) & (n_n4651) & (n_n4622)) + ((n_n4641) & (!n_n4648) & (!n_n4651) & (!n_n4622)) + ((n_n4641) & (!n_n4648) & (!n_n4651) & (n_n4622)) + ((n_n4641) & (!n_n4648) & (n_n4651) & (!n_n4622)) + ((n_n4641) & (!n_n4648) & (n_n4651) & (n_n4622)) + ((n_n4641) & (n_n4648) & (!n_n4651) & (!n_n4622)) + ((n_n4641) & (n_n4648) & (!n_n4651) & (n_n4622)) + ((n_n4641) & (n_n4648) & (n_n4651) & (!n_n4622)) + ((n_n4641) & (n_n4648) & (n_n4651) & (n_n4622)));
	assign x15830x = (((!n_n4597) & (!n_n4596) & (!n_n4631) & (!n_n4620) & (n_n4627)) + ((!n_n4597) & (!n_n4596) & (!n_n4631) & (n_n4620) & (!n_n4627)) + ((!n_n4597) & (!n_n4596) & (!n_n4631) & (n_n4620) & (n_n4627)) + ((!n_n4597) & (!n_n4596) & (n_n4631) & (!n_n4620) & (!n_n4627)) + ((!n_n4597) & (!n_n4596) & (n_n4631) & (!n_n4620) & (n_n4627)) + ((!n_n4597) & (!n_n4596) & (n_n4631) & (n_n4620) & (!n_n4627)) + ((!n_n4597) & (!n_n4596) & (n_n4631) & (n_n4620) & (n_n4627)) + ((!n_n4597) & (n_n4596) & (!n_n4631) & (!n_n4620) & (!n_n4627)) + ((!n_n4597) & (n_n4596) & (!n_n4631) & (!n_n4620) & (n_n4627)) + ((!n_n4597) & (n_n4596) & (!n_n4631) & (n_n4620) & (!n_n4627)) + ((!n_n4597) & (n_n4596) & (!n_n4631) & (n_n4620) & (n_n4627)) + ((!n_n4597) & (n_n4596) & (n_n4631) & (!n_n4620) & (!n_n4627)) + ((!n_n4597) & (n_n4596) & (n_n4631) & (!n_n4620) & (n_n4627)) + ((!n_n4597) & (n_n4596) & (n_n4631) & (n_n4620) & (!n_n4627)) + ((!n_n4597) & (n_n4596) & (n_n4631) & (n_n4620) & (n_n4627)) + ((n_n4597) & (!n_n4596) & (!n_n4631) & (!n_n4620) & (!n_n4627)) + ((n_n4597) & (!n_n4596) & (!n_n4631) & (!n_n4620) & (n_n4627)) + ((n_n4597) & (!n_n4596) & (!n_n4631) & (n_n4620) & (!n_n4627)) + ((n_n4597) & (!n_n4596) & (!n_n4631) & (n_n4620) & (n_n4627)) + ((n_n4597) & (!n_n4596) & (n_n4631) & (!n_n4620) & (!n_n4627)) + ((n_n4597) & (!n_n4596) & (n_n4631) & (!n_n4620) & (n_n4627)) + ((n_n4597) & (!n_n4596) & (n_n4631) & (n_n4620) & (!n_n4627)) + ((n_n4597) & (!n_n4596) & (n_n4631) & (n_n4620) & (n_n4627)) + ((n_n4597) & (n_n4596) & (!n_n4631) & (!n_n4620) & (!n_n4627)) + ((n_n4597) & (n_n4596) & (!n_n4631) & (!n_n4620) & (n_n4627)) + ((n_n4597) & (n_n4596) & (!n_n4631) & (n_n4620) & (!n_n4627)) + ((n_n4597) & (n_n4596) & (!n_n4631) & (n_n4620) & (n_n4627)) + ((n_n4597) & (n_n4596) & (n_n4631) & (!n_n4620) & (!n_n4627)) + ((n_n4597) & (n_n4596) & (n_n4631) & (!n_n4620) & (n_n4627)) + ((n_n4597) & (n_n4596) & (n_n4631) & (n_n4620) & (!n_n4627)) + ((n_n4597) & (n_n4596) & (n_n4631) & (n_n4620) & (n_n4627)));
	assign x15909x = (((!n_n4373) & (!n_n4392) & (!n_n4426) & (n_n4419)) + ((!n_n4373) & (!n_n4392) & (n_n4426) & (!n_n4419)) + ((!n_n4373) & (!n_n4392) & (n_n4426) & (n_n4419)) + ((!n_n4373) & (n_n4392) & (!n_n4426) & (!n_n4419)) + ((!n_n4373) & (n_n4392) & (!n_n4426) & (n_n4419)) + ((!n_n4373) & (n_n4392) & (n_n4426) & (!n_n4419)) + ((!n_n4373) & (n_n4392) & (n_n4426) & (n_n4419)) + ((n_n4373) & (!n_n4392) & (!n_n4426) & (!n_n4419)) + ((n_n4373) & (!n_n4392) & (!n_n4426) & (n_n4419)) + ((n_n4373) & (!n_n4392) & (n_n4426) & (!n_n4419)) + ((n_n4373) & (!n_n4392) & (n_n4426) & (n_n4419)) + ((n_n4373) & (n_n4392) & (!n_n4426) & (!n_n4419)) + ((n_n4373) & (n_n4392) & (!n_n4426) & (n_n4419)) + ((n_n4373) & (n_n4392) & (n_n4426) & (!n_n4419)) + ((n_n4373) & (n_n4392) & (n_n4426) & (n_n4419)));
	assign x15910x = (((!n_n4420) & (!n_n4407) & (!n_n4394) & (!n_n4376) & (n_n4412)) + ((!n_n4420) & (!n_n4407) & (!n_n4394) & (n_n4376) & (!n_n4412)) + ((!n_n4420) & (!n_n4407) & (!n_n4394) & (n_n4376) & (n_n4412)) + ((!n_n4420) & (!n_n4407) & (n_n4394) & (!n_n4376) & (!n_n4412)) + ((!n_n4420) & (!n_n4407) & (n_n4394) & (!n_n4376) & (n_n4412)) + ((!n_n4420) & (!n_n4407) & (n_n4394) & (n_n4376) & (!n_n4412)) + ((!n_n4420) & (!n_n4407) & (n_n4394) & (n_n4376) & (n_n4412)) + ((!n_n4420) & (n_n4407) & (!n_n4394) & (!n_n4376) & (!n_n4412)) + ((!n_n4420) & (n_n4407) & (!n_n4394) & (!n_n4376) & (n_n4412)) + ((!n_n4420) & (n_n4407) & (!n_n4394) & (n_n4376) & (!n_n4412)) + ((!n_n4420) & (n_n4407) & (!n_n4394) & (n_n4376) & (n_n4412)) + ((!n_n4420) & (n_n4407) & (n_n4394) & (!n_n4376) & (!n_n4412)) + ((!n_n4420) & (n_n4407) & (n_n4394) & (!n_n4376) & (n_n4412)) + ((!n_n4420) & (n_n4407) & (n_n4394) & (n_n4376) & (!n_n4412)) + ((!n_n4420) & (n_n4407) & (n_n4394) & (n_n4376) & (n_n4412)) + ((n_n4420) & (!n_n4407) & (!n_n4394) & (!n_n4376) & (!n_n4412)) + ((n_n4420) & (!n_n4407) & (!n_n4394) & (!n_n4376) & (n_n4412)) + ((n_n4420) & (!n_n4407) & (!n_n4394) & (n_n4376) & (!n_n4412)) + ((n_n4420) & (!n_n4407) & (!n_n4394) & (n_n4376) & (n_n4412)) + ((n_n4420) & (!n_n4407) & (n_n4394) & (!n_n4376) & (!n_n4412)) + ((n_n4420) & (!n_n4407) & (n_n4394) & (!n_n4376) & (n_n4412)) + ((n_n4420) & (!n_n4407) & (n_n4394) & (n_n4376) & (!n_n4412)) + ((n_n4420) & (!n_n4407) & (n_n4394) & (n_n4376) & (n_n4412)) + ((n_n4420) & (n_n4407) & (!n_n4394) & (!n_n4376) & (!n_n4412)) + ((n_n4420) & (n_n4407) & (!n_n4394) & (!n_n4376) & (n_n4412)) + ((n_n4420) & (n_n4407) & (!n_n4394) & (n_n4376) & (!n_n4412)) + ((n_n4420) & (n_n4407) & (!n_n4394) & (n_n4376) & (n_n4412)) + ((n_n4420) & (n_n4407) & (n_n4394) & (!n_n4376) & (!n_n4412)) + ((n_n4420) & (n_n4407) & (n_n4394) & (!n_n4376) & (n_n4412)) + ((n_n4420) & (n_n4407) & (n_n4394) & (n_n4376) & (!n_n4412)) + ((n_n4420) & (n_n4407) & (n_n4394) & (n_n4376) & (n_n4412)));
	assign x15915x = (((!n_n4464) & (!n_n4433) & (!n_n4455) & (n_n4441)) + ((!n_n4464) & (!n_n4433) & (n_n4455) & (!n_n4441)) + ((!n_n4464) & (!n_n4433) & (n_n4455) & (n_n4441)) + ((!n_n4464) & (n_n4433) & (!n_n4455) & (!n_n4441)) + ((!n_n4464) & (n_n4433) & (!n_n4455) & (n_n4441)) + ((!n_n4464) & (n_n4433) & (n_n4455) & (!n_n4441)) + ((!n_n4464) & (n_n4433) & (n_n4455) & (n_n4441)) + ((n_n4464) & (!n_n4433) & (!n_n4455) & (!n_n4441)) + ((n_n4464) & (!n_n4433) & (!n_n4455) & (n_n4441)) + ((n_n4464) & (!n_n4433) & (n_n4455) & (!n_n4441)) + ((n_n4464) & (!n_n4433) & (n_n4455) & (n_n4441)) + ((n_n4464) & (n_n4433) & (!n_n4455) & (!n_n4441)) + ((n_n4464) & (n_n4433) & (!n_n4455) & (n_n4441)) + ((n_n4464) & (n_n4433) & (n_n4455) & (!n_n4441)) + ((n_n4464) & (n_n4433) & (n_n4455) & (n_n4441)));
	assign x15916x = (((!n_n4432) & (!n_n4451) & (!n_n4468) & (!n_n4458) & (n_n4435)) + ((!n_n4432) & (!n_n4451) & (!n_n4468) & (n_n4458) & (!n_n4435)) + ((!n_n4432) & (!n_n4451) & (!n_n4468) & (n_n4458) & (n_n4435)) + ((!n_n4432) & (!n_n4451) & (n_n4468) & (!n_n4458) & (!n_n4435)) + ((!n_n4432) & (!n_n4451) & (n_n4468) & (!n_n4458) & (n_n4435)) + ((!n_n4432) & (!n_n4451) & (n_n4468) & (n_n4458) & (!n_n4435)) + ((!n_n4432) & (!n_n4451) & (n_n4468) & (n_n4458) & (n_n4435)) + ((!n_n4432) & (n_n4451) & (!n_n4468) & (!n_n4458) & (!n_n4435)) + ((!n_n4432) & (n_n4451) & (!n_n4468) & (!n_n4458) & (n_n4435)) + ((!n_n4432) & (n_n4451) & (!n_n4468) & (n_n4458) & (!n_n4435)) + ((!n_n4432) & (n_n4451) & (!n_n4468) & (n_n4458) & (n_n4435)) + ((!n_n4432) & (n_n4451) & (n_n4468) & (!n_n4458) & (!n_n4435)) + ((!n_n4432) & (n_n4451) & (n_n4468) & (!n_n4458) & (n_n4435)) + ((!n_n4432) & (n_n4451) & (n_n4468) & (n_n4458) & (!n_n4435)) + ((!n_n4432) & (n_n4451) & (n_n4468) & (n_n4458) & (n_n4435)) + ((n_n4432) & (!n_n4451) & (!n_n4468) & (!n_n4458) & (!n_n4435)) + ((n_n4432) & (!n_n4451) & (!n_n4468) & (!n_n4458) & (n_n4435)) + ((n_n4432) & (!n_n4451) & (!n_n4468) & (n_n4458) & (!n_n4435)) + ((n_n4432) & (!n_n4451) & (!n_n4468) & (n_n4458) & (n_n4435)) + ((n_n4432) & (!n_n4451) & (n_n4468) & (!n_n4458) & (!n_n4435)) + ((n_n4432) & (!n_n4451) & (n_n4468) & (!n_n4458) & (n_n4435)) + ((n_n4432) & (!n_n4451) & (n_n4468) & (n_n4458) & (!n_n4435)) + ((n_n4432) & (!n_n4451) & (n_n4468) & (n_n4458) & (n_n4435)) + ((n_n4432) & (n_n4451) & (!n_n4468) & (!n_n4458) & (!n_n4435)) + ((n_n4432) & (n_n4451) & (!n_n4468) & (!n_n4458) & (n_n4435)) + ((n_n4432) & (n_n4451) & (!n_n4468) & (n_n4458) & (!n_n4435)) + ((n_n4432) & (n_n4451) & (!n_n4468) & (n_n4458) & (n_n4435)) + ((n_n4432) & (n_n4451) & (n_n4468) & (!n_n4458) & (!n_n4435)) + ((n_n4432) & (n_n4451) & (n_n4468) & (!n_n4458) & (n_n4435)) + ((n_n4432) & (n_n4451) & (n_n4468) & (n_n4458) & (!n_n4435)) + ((n_n4432) & (n_n4451) & (n_n4468) & (n_n4458) & (n_n4435)));
	assign x22074x = (((!n_n4784) & (!n_n4754) & (!n_n4787) & (!n_n4781)));
	assign x15932x = (((!n_n4748) & (!n_n4766) & (!n_n4772) & (!x164x) & (!x22074x)) + ((!n_n4748) & (!n_n4766) & (!n_n4772) & (x164x) & (!x22074x)) + ((!n_n4748) & (!n_n4766) & (!n_n4772) & (x164x) & (x22074x)) + ((!n_n4748) & (!n_n4766) & (n_n4772) & (!x164x) & (!x22074x)) + ((!n_n4748) & (!n_n4766) & (n_n4772) & (!x164x) & (x22074x)) + ((!n_n4748) & (!n_n4766) & (n_n4772) & (x164x) & (!x22074x)) + ((!n_n4748) & (!n_n4766) & (n_n4772) & (x164x) & (x22074x)) + ((!n_n4748) & (n_n4766) & (!n_n4772) & (!x164x) & (!x22074x)) + ((!n_n4748) & (n_n4766) & (!n_n4772) & (!x164x) & (x22074x)) + ((!n_n4748) & (n_n4766) & (!n_n4772) & (x164x) & (!x22074x)) + ((!n_n4748) & (n_n4766) & (!n_n4772) & (x164x) & (x22074x)) + ((!n_n4748) & (n_n4766) & (n_n4772) & (!x164x) & (!x22074x)) + ((!n_n4748) & (n_n4766) & (n_n4772) & (!x164x) & (x22074x)) + ((!n_n4748) & (n_n4766) & (n_n4772) & (x164x) & (!x22074x)) + ((!n_n4748) & (n_n4766) & (n_n4772) & (x164x) & (x22074x)) + ((n_n4748) & (!n_n4766) & (!n_n4772) & (!x164x) & (!x22074x)) + ((n_n4748) & (!n_n4766) & (!n_n4772) & (!x164x) & (x22074x)) + ((n_n4748) & (!n_n4766) & (!n_n4772) & (x164x) & (!x22074x)) + ((n_n4748) & (!n_n4766) & (!n_n4772) & (x164x) & (x22074x)) + ((n_n4748) & (!n_n4766) & (n_n4772) & (!x164x) & (!x22074x)) + ((n_n4748) & (!n_n4766) & (n_n4772) & (!x164x) & (x22074x)) + ((n_n4748) & (!n_n4766) & (n_n4772) & (x164x) & (!x22074x)) + ((n_n4748) & (!n_n4766) & (n_n4772) & (x164x) & (x22074x)) + ((n_n4748) & (n_n4766) & (!n_n4772) & (!x164x) & (!x22074x)) + ((n_n4748) & (n_n4766) & (!n_n4772) & (!x164x) & (x22074x)) + ((n_n4748) & (n_n4766) & (!n_n4772) & (x164x) & (!x22074x)) + ((n_n4748) & (n_n4766) & (!n_n4772) & (x164x) & (x22074x)) + ((n_n4748) & (n_n4766) & (n_n4772) & (!x164x) & (!x22074x)) + ((n_n4748) & (n_n4766) & (n_n4772) & (!x164x) & (x22074x)) + ((n_n4748) & (n_n4766) & (n_n4772) & (x164x) & (!x22074x)) + ((n_n4748) & (n_n4766) & (n_n4772) & (x164x) & (x22074x)));
	assign x15920x = (((!n_n4656) & (!n_n4676) & (!n_n4655) & (n_n4657)) + ((!n_n4656) & (!n_n4676) & (n_n4655) & (!n_n4657)) + ((!n_n4656) & (!n_n4676) & (n_n4655) & (n_n4657)) + ((!n_n4656) & (n_n4676) & (!n_n4655) & (!n_n4657)) + ((!n_n4656) & (n_n4676) & (!n_n4655) & (n_n4657)) + ((!n_n4656) & (n_n4676) & (n_n4655) & (!n_n4657)) + ((!n_n4656) & (n_n4676) & (n_n4655) & (n_n4657)) + ((n_n4656) & (!n_n4676) & (!n_n4655) & (!n_n4657)) + ((n_n4656) & (!n_n4676) & (!n_n4655) & (n_n4657)) + ((n_n4656) & (!n_n4676) & (n_n4655) & (!n_n4657)) + ((n_n4656) & (!n_n4676) & (n_n4655) & (n_n4657)) + ((n_n4656) & (n_n4676) & (!n_n4655) & (!n_n4657)) + ((n_n4656) & (n_n4676) & (!n_n4655) & (n_n4657)) + ((n_n4656) & (n_n4676) & (n_n4655) & (!n_n4657)) + ((n_n4656) & (n_n4676) & (n_n4655) & (n_n4657)));
	assign x15921x = (((!x10x) & (!n_n473) & (!n_n520) & (!n_n1764) & (n_n4687)) + ((!x10x) & (!n_n473) & (!n_n520) & (n_n1764) & (!n_n4687)) + ((!x10x) & (!n_n473) & (!n_n520) & (n_n1764) & (n_n4687)) + ((!x10x) & (!n_n473) & (n_n520) & (!n_n1764) & (n_n4687)) + ((!x10x) & (!n_n473) & (n_n520) & (n_n1764) & (!n_n4687)) + ((!x10x) & (!n_n473) & (n_n520) & (n_n1764) & (n_n4687)) + ((!x10x) & (n_n473) & (!n_n520) & (!n_n1764) & (n_n4687)) + ((!x10x) & (n_n473) & (!n_n520) & (n_n1764) & (!n_n4687)) + ((!x10x) & (n_n473) & (!n_n520) & (n_n1764) & (n_n4687)) + ((!x10x) & (n_n473) & (n_n520) & (!n_n1764) & (n_n4687)) + ((!x10x) & (n_n473) & (n_n520) & (n_n1764) & (!n_n4687)) + ((!x10x) & (n_n473) & (n_n520) & (n_n1764) & (n_n4687)) + ((x10x) & (!n_n473) & (!n_n520) & (!n_n1764) & (n_n4687)) + ((x10x) & (!n_n473) & (!n_n520) & (n_n1764) & (!n_n4687)) + ((x10x) & (!n_n473) & (!n_n520) & (n_n1764) & (n_n4687)) + ((x10x) & (!n_n473) & (n_n520) & (!n_n1764) & (n_n4687)) + ((x10x) & (!n_n473) & (n_n520) & (n_n1764) & (!n_n4687)) + ((x10x) & (!n_n473) & (n_n520) & (n_n1764) & (n_n4687)) + ((x10x) & (n_n473) & (!n_n520) & (!n_n1764) & (n_n4687)) + ((x10x) & (n_n473) & (!n_n520) & (n_n1764) & (!n_n4687)) + ((x10x) & (n_n473) & (!n_n520) & (n_n1764) & (n_n4687)) + ((x10x) & (n_n473) & (n_n520) & (!n_n1764) & (!n_n4687)) + ((x10x) & (n_n473) & (n_n520) & (!n_n1764) & (n_n4687)) + ((x10x) & (n_n473) & (n_n520) & (n_n1764) & (!n_n4687)) + ((x10x) & (n_n473) & (n_n520) & (n_n1764) & (n_n4687)));
	assign x15924x = (((!x10x) & (!x516x) & (!n_n4727) & (!n_n4711) & (n_n4688)) + ((!x10x) & (!x516x) & (!n_n4727) & (n_n4711) & (!n_n4688)) + ((!x10x) & (!x516x) & (!n_n4727) & (n_n4711) & (n_n4688)) + ((!x10x) & (!x516x) & (n_n4727) & (!n_n4711) & (!n_n4688)) + ((!x10x) & (!x516x) & (n_n4727) & (!n_n4711) & (n_n4688)) + ((!x10x) & (!x516x) & (n_n4727) & (n_n4711) & (!n_n4688)) + ((!x10x) & (!x516x) & (n_n4727) & (n_n4711) & (n_n4688)) + ((!x10x) & (x516x) & (!n_n4727) & (!n_n4711) & (n_n4688)) + ((!x10x) & (x516x) & (!n_n4727) & (n_n4711) & (!n_n4688)) + ((!x10x) & (x516x) & (!n_n4727) & (n_n4711) & (n_n4688)) + ((!x10x) & (x516x) & (n_n4727) & (!n_n4711) & (!n_n4688)) + ((!x10x) & (x516x) & (n_n4727) & (!n_n4711) & (n_n4688)) + ((!x10x) & (x516x) & (n_n4727) & (n_n4711) & (!n_n4688)) + ((!x10x) & (x516x) & (n_n4727) & (n_n4711) & (n_n4688)) + ((x10x) & (!x516x) & (!n_n4727) & (!n_n4711) & (n_n4688)) + ((x10x) & (!x516x) & (!n_n4727) & (n_n4711) & (!n_n4688)) + ((x10x) & (!x516x) & (!n_n4727) & (n_n4711) & (n_n4688)) + ((x10x) & (!x516x) & (n_n4727) & (!n_n4711) & (!n_n4688)) + ((x10x) & (!x516x) & (n_n4727) & (!n_n4711) & (n_n4688)) + ((x10x) & (!x516x) & (n_n4727) & (n_n4711) & (!n_n4688)) + ((x10x) & (!x516x) & (n_n4727) & (n_n4711) & (n_n4688)) + ((x10x) & (x516x) & (!n_n4727) & (!n_n4711) & (!n_n4688)) + ((x10x) & (x516x) & (!n_n4727) & (!n_n4711) & (n_n4688)) + ((x10x) & (x516x) & (!n_n4727) & (n_n4711) & (!n_n4688)) + ((x10x) & (x516x) & (!n_n4727) & (n_n4711) & (n_n4688)) + ((x10x) & (x516x) & (n_n4727) & (!n_n4711) & (!n_n4688)) + ((x10x) & (x516x) & (n_n4727) & (!n_n4711) & (n_n4688)) + ((x10x) & (x516x) & (n_n4727) & (n_n4711) & (!n_n4688)) + ((x10x) & (x516x) & (n_n4727) & (n_n4711) & (n_n4688)));
	assign x15925x = (((!n_n518) & (!n_n325) & (!x20x) & (!n_n4700) & (n_n1760)) + ((!n_n518) & (!n_n325) & (!x20x) & (n_n4700) & (!n_n1760)) + ((!n_n518) & (!n_n325) & (!x20x) & (n_n4700) & (n_n1760)) + ((!n_n518) & (!n_n325) & (x20x) & (!n_n4700) & (n_n1760)) + ((!n_n518) & (!n_n325) & (x20x) & (n_n4700) & (!n_n1760)) + ((!n_n518) & (!n_n325) & (x20x) & (n_n4700) & (n_n1760)) + ((!n_n518) & (n_n325) & (!x20x) & (!n_n4700) & (n_n1760)) + ((!n_n518) & (n_n325) & (!x20x) & (n_n4700) & (!n_n1760)) + ((!n_n518) & (n_n325) & (!x20x) & (n_n4700) & (n_n1760)) + ((!n_n518) & (n_n325) & (x20x) & (!n_n4700) & (n_n1760)) + ((!n_n518) & (n_n325) & (x20x) & (n_n4700) & (!n_n1760)) + ((!n_n518) & (n_n325) & (x20x) & (n_n4700) & (n_n1760)) + ((n_n518) & (!n_n325) & (!x20x) & (!n_n4700) & (n_n1760)) + ((n_n518) & (!n_n325) & (!x20x) & (n_n4700) & (!n_n1760)) + ((n_n518) & (!n_n325) & (!x20x) & (n_n4700) & (n_n1760)) + ((n_n518) & (!n_n325) & (x20x) & (!n_n4700) & (n_n1760)) + ((n_n518) & (!n_n325) & (x20x) & (n_n4700) & (!n_n1760)) + ((n_n518) & (!n_n325) & (x20x) & (n_n4700) & (n_n1760)) + ((n_n518) & (n_n325) & (!x20x) & (!n_n4700) & (n_n1760)) + ((n_n518) & (n_n325) & (!x20x) & (n_n4700) & (!n_n1760)) + ((n_n518) & (n_n325) & (!x20x) & (n_n4700) & (n_n1760)) + ((n_n518) & (n_n325) & (x20x) & (!n_n4700) & (!n_n1760)) + ((n_n518) & (n_n325) & (x20x) & (!n_n4700) & (n_n1760)) + ((n_n518) & (n_n325) & (x20x) & (n_n4700) & (!n_n1760)) + ((n_n518) & (n_n325) & (x20x) & (n_n4700) & (n_n1760)));
	assign x12425x = (((!i_9_) & (n_n390) & (n_n473) & (!n_n534) & (n_n530)) + ((!i_9_) & (n_n390) & (n_n473) & (n_n534) & (!n_n530)) + ((!i_9_) & (n_n390) & (n_n473) & (n_n534) & (n_n530)) + ((i_9_) & (n_n390) & (n_n473) & (!n_n534) & (n_n530)) + ((i_9_) & (n_n390) & (n_n473) & (n_n534) & (!n_n530)) + ((i_9_) & (n_n390) & (n_n473) & (n_n534) & (n_n530)));
	assign x12364x = (((!x19x) & (!x516x) & (!n_n5327) & (!n_n5323) & (n_n5333)) + ((!x19x) & (!x516x) & (!n_n5327) & (n_n5323) & (!n_n5333)) + ((!x19x) & (!x516x) & (!n_n5327) & (n_n5323) & (n_n5333)) + ((!x19x) & (!x516x) & (n_n5327) & (!n_n5323) & (!n_n5333)) + ((!x19x) & (!x516x) & (n_n5327) & (!n_n5323) & (n_n5333)) + ((!x19x) & (!x516x) & (n_n5327) & (n_n5323) & (!n_n5333)) + ((!x19x) & (!x516x) & (n_n5327) & (n_n5323) & (n_n5333)) + ((!x19x) & (x516x) & (!n_n5327) & (!n_n5323) & (n_n5333)) + ((!x19x) & (x516x) & (!n_n5327) & (n_n5323) & (!n_n5333)) + ((!x19x) & (x516x) & (!n_n5327) & (n_n5323) & (n_n5333)) + ((!x19x) & (x516x) & (n_n5327) & (!n_n5323) & (!n_n5333)) + ((!x19x) & (x516x) & (n_n5327) & (!n_n5323) & (n_n5333)) + ((!x19x) & (x516x) & (n_n5327) & (n_n5323) & (!n_n5333)) + ((!x19x) & (x516x) & (n_n5327) & (n_n5323) & (n_n5333)) + ((x19x) & (!x516x) & (!n_n5327) & (!n_n5323) & (n_n5333)) + ((x19x) & (!x516x) & (!n_n5327) & (n_n5323) & (!n_n5333)) + ((x19x) & (!x516x) & (!n_n5327) & (n_n5323) & (n_n5333)) + ((x19x) & (!x516x) & (n_n5327) & (!n_n5323) & (!n_n5333)) + ((x19x) & (!x516x) & (n_n5327) & (!n_n5323) & (n_n5333)) + ((x19x) & (!x516x) & (n_n5327) & (n_n5323) & (!n_n5333)) + ((x19x) & (!x516x) & (n_n5327) & (n_n5323) & (n_n5333)) + ((x19x) & (x516x) & (!n_n5327) & (!n_n5323) & (!n_n5333)) + ((x19x) & (x516x) & (!n_n5327) & (!n_n5323) & (n_n5333)) + ((x19x) & (x516x) & (!n_n5327) & (n_n5323) & (!n_n5333)) + ((x19x) & (x516x) & (!n_n5327) & (n_n5323) & (n_n5333)) + ((x19x) & (x516x) & (n_n5327) & (!n_n5323) & (!n_n5333)) + ((x19x) & (x516x) & (n_n5327) & (!n_n5323) & (n_n5333)) + ((x19x) & (x516x) & (n_n5327) & (n_n5323) & (!n_n5333)) + ((x19x) & (x516x) & (n_n5327) & (n_n5323) & (n_n5333)));
	assign x261x = (((!i_9_) & (n_n534) & (n_n260) & (n_n491)) + ((i_9_) & (n_n534) & (n_n260) & (n_n491)));
	assign x22106x = (((!x19x) & (!n_n5310) & (!x502x) & (!n_n5311) & (!n_n5317)) + ((!x19x) & (!n_n5310) & (x502x) & (!n_n5311) & (!n_n5317)) + ((x19x) & (!n_n5310) & (!x502x) & (!n_n5311) & (!n_n5317)));
	assign x22178x = (((!n_n4717) & (!n_n4719) & (!n_n4715) & (!n_n4714)));
	assign n_n2982 = (((!n_n4720) & (!x39x) & (!n_n4716) & (!n_n4713) & (!x22178x)) + ((!n_n4720) & (!x39x) & (!n_n4716) & (n_n4713) & (!x22178x)) + ((!n_n4720) & (!x39x) & (!n_n4716) & (n_n4713) & (x22178x)) + ((!n_n4720) & (!x39x) & (n_n4716) & (!n_n4713) & (!x22178x)) + ((!n_n4720) & (!x39x) & (n_n4716) & (!n_n4713) & (x22178x)) + ((!n_n4720) & (!x39x) & (n_n4716) & (n_n4713) & (!x22178x)) + ((!n_n4720) & (!x39x) & (n_n4716) & (n_n4713) & (x22178x)) + ((!n_n4720) & (x39x) & (!n_n4716) & (!n_n4713) & (!x22178x)) + ((!n_n4720) & (x39x) & (!n_n4716) & (!n_n4713) & (x22178x)) + ((!n_n4720) & (x39x) & (!n_n4716) & (n_n4713) & (!x22178x)) + ((!n_n4720) & (x39x) & (!n_n4716) & (n_n4713) & (x22178x)) + ((!n_n4720) & (x39x) & (n_n4716) & (!n_n4713) & (!x22178x)) + ((!n_n4720) & (x39x) & (n_n4716) & (!n_n4713) & (x22178x)) + ((!n_n4720) & (x39x) & (n_n4716) & (n_n4713) & (!x22178x)) + ((!n_n4720) & (x39x) & (n_n4716) & (n_n4713) & (x22178x)) + ((n_n4720) & (!x39x) & (!n_n4716) & (!n_n4713) & (!x22178x)) + ((n_n4720) & (!x39x) & (!n_n4716) & (!n_n4713) & (x22178x)) + ((n_n4720) & (!x39x) & (!n_n4716) & (n_n4713) & (!x22178x)) + ((n_n4720) & (!x39x) & (!n_n4716) & (n_n4713) & (x22178x)) + ((n_n4720) & (!x39x) & (n_n4716) & (!n_n4713) & (!x22178x)) + ((n_n4720) & (!x39x) & (n_n4716) & (!n_n4713) & (x22178x)) + ((n_n4720) & (!x39x) & (n_n4716) & (n_n4713) & (!x22178x)) + ((n_n4720) & (!x39x) & (n_n4716) & (n_n4713) & (x22178x)) + ((n_n4720) & (x39x) & (!n_n4716) & (!n_n4713) & (!x22178x)) + ((n_n4720) & (x39x) & (!n_n4716) & (!n_n4713) & (x22178x)) + ((n_n4720) & (x39x) & (!n_n4716) & (n_n4713) & (!x22178x)) + ((n_n4720) & (x39x) & (!n_n4716) & (n_n4713) & (x22178x)) + ((n_n4720) & (x39x) & (n_n4716) & (!n_n4713) & (!x22178x)) + ((n_n4720) & (x39x) & (n_n4716) & (!n_n4713) & (x22178x)) + ((n_n4720) & (x39x) & (n_n4716) & (n_n4713) & (!x22178x)) + ((n_n4720) & (x39x) & (n_n4716) & (n_n4713) & (x22178x)));
	assign x15607x = (((!n_n5091) & (!n_n5100) & (!n_n5089) & (!n_n5098) & (n_n5095)) + ((!n_n5091) & (!n_n5100) & (!n_n5089) & (n_n5098) & (!n_n5095)) + ((!n_n5091) & (!n_n5100) & (!n_n5089) & (n_n5098) & (n_n5095)) + ((!n_n5091) & (!n_n5100) & (n_n5089) & (!n_n5098) & (!n_n5095)) + ((!n_n5091) & (!n_n5100) & (n_n5089) & (!n_n5098) & (n_n5095)) + ((!n_n5091) & (!n_n5100) & (n_n5089) & (n_n5098) & (!n_n5095)) + ((!n_n5091) & (!n_n5100) & (n_n5089) & (n_n5098) & (n_n5095)) + ((!n_n5091) & (n_n5100) & (!n_n5089) & (!n_n5098) & (!n_n5095)) + ((!n_n5091) & (n_n5100) & (!n_n5089) & (!n_n5098) & (n_n5095)) + ((!n_n5091) & (n_n5100) & (!n_n5089) & (n_n5098) & (!n_n5095)) + ((!n_n5091) & (n_n5100) & (!n_n5089) & (n_n5098) & (n_n5095)) + ((!n_n5091) & (n_n5100) & (n_n5089) & (!n_n5098) & (!n_n5095)) + ((!n_n5091) & (n_n5100) & (n_n5089) & (!n_n5098) & (n_n5095)) + ((!n_n5091) & (n_n5100) & (n_n5089) & (n_n5098) & (!n_n5095)) + ((!n_n5091) & (n_n5100) & (n_n5089) & (n_n5098) & (n_n5095)) + ((n_n5091) & (!n_n5100) & (!n_n5089) & (!n_n5098) & (!n_n5095)) + ((n_n5091) & (!n_n5100) & (!n_n5089) & (!n_n5098) & (n_n5095)) + ((n_n5091) & (!n_n5100) & (!n_n5089) & (n_n5098) & (!n_n5095)) + ((n_n5091) & (!n_n5100) & (!n_n5089) & (n_n5098) & (n_n5095)) + ((n_n5091) & (!n_n5100) & (n_n5089) & (!n_n5098) & (!n_n5095)) + ((n_n5091) & (!n_n5100) & (n_n5089) & (!n_n5098) & (n_n5095)) + ((n_n5091) & (!n_n5100) & (n_n5089) & (n_n5098) & (!n_n5095)) + ((n_n5091) & (!n_n5100) & (n_n5089) & (n_n5098) & (n_n5095)) + ((n_n5091) & (n_n5100) & (!n_n5089) & (!n_n5098) & (!n_n5095)) + ((n_n5091) & (n_n5100) & (!n_n5089) & (!n_n5098) & (n_n5095)) + ((n_n5091) & (n_n5100) & (!n_n5089) & (n_n5098) & (!n_n5095)) + ((n_n5091) & (n_n5100) & (!n_n5089) & (n_n5098) & (n_n5095)) + ((n_n5091) & (n_n5100) & (n_n5089) & (!n_n5098) & (!n_n5095)) + ((n_n5091) & (n_n5100) & (n_n5089) & (!n_n5098) & (n_n5095)) + ((n_n5091) & (n_n5100) & (n_n5089) & (n_n5098) & (!n_n5095)) + ((n_n5091) & (n_n5100) & (n_n5089) & (n_n5098) & (n_n5095)));
	assign x15611x = (((!n_n5057) & (!n_n5058) & (!n_n5072) & (!n_n5061) & (n_n5065)) + ((!n_n5057) & (!n_n5058) & (!n_n5072) & (n_n5061) & (!n_n5065)) + ((!n_n5057) & (!n_n5058) & (!n_n5072) & (n_n5061) & (n_n5065)) + ((!n_n5057) & (!n_n5058) & (n_n5072) & (!n_n5061) & (!n_n5065)) + ((!n_n5057) & (!n_n5058) & (n_n5072) & (!n_n5061) & (n_n5065)) + ((!n_n5057) & (!n_n5058) & (n_n5072) & (n_n5061) & (!n_n5065)) + ((!n_n5057) & (!n_n5058) & (n_n5072) & (n_n5061) & (n_n5065)) + ((!n_n5057) & (n_n5058) & (!n_n5072) & (!n_n5061) & (!n_n5065)) + ((!n_n5057) & (n_n5058) & (!n_n5072) & (!n_n5061) & (n_n5065)) + ((!n_n5057) & (n_n5058) & (!n_n5072) & (n_n5061) & (!n_n5065)) + ((!n_n5057) & (n_n5058) & (!n_n5072) & (n_n5061) & (n_n5065)) + ((!n_n5057) & (n_n5058) & (n_n5072) & (!n_n5061) & (!n_n5065)) + ((!n_n5057) & (n_n5058) & (n_n5072) & (!n_n5061) & (n_n5065)) + ((!n_n5057) & (n_n5058) & (n_n5072) & (n_n5061) & (!n_n5065)) + ((!n_n5057) & (n_n5058) & (n_n5072) & (n_n5061) & (n_n5065)) + ((n_n5057) & (!n_n5058) & (!n_n5072) & (!n_n5061) & (!n_n5065)) + ((n_n5057) & (!n_n5058) & (!n_n5072) & (!n_n5061) & (n_n5065)) + ((n_n5057) & (!n_n5058) & (!n_n5072) & (n_n5061) & (!n_n5065)) + ((n_n5057) & (!n_n5058) & (!n_n5072) & (n_n5061) & (n_n5065)) + ((n_n5057) & (!n_n5058) & (n_n5072) & (!n_n5061) & (!n_n5065)) + ((n_n5057) & (!n_n5058) & (n_n5072) & (!n_n5061) & (n_n5065)) + ((n_n5057) & (!n_n5058) & (n_n5072) & (n_n5061) & (!n_n5065)) + ((n_n5057) & (!n_n5058) & (n_n5072) & (n_n5061) & (n_n5065)) + ((n_n5057) & (n_n5058) & (!n_n5072) & (!n_n5061) & (!n_n5065)) + ((n_n5057) & (n_n5058) & (!n_n5072) & (!n_n5061) & (n_n5065)) + ((n_n5057) & (n_n5058) & (!n_n5072) & (n_n5061) & (!n_n5065)) + ((n_n5057) & (n_n5058) & (!n_n5072) & (n_n5061) & (n_n5065)) + ((n_n5057) & (n_n5058) & (n_n5072) & (!n_n5061) & (!n_n5065)) + ((n_n5057) & (n_n5058) & (n_n5072) & (!n_n5061) & (n_n5065)) + ((n_n5057) & (n_n5058) & (n_n5072) & (n_n5061) & (!n_n5065)) + ((n_n5057) & (n_n5058) & (n_n5072) & (n_n5061) & (n_n5065)));
	assign x22088x = (((!x18x) & (!x516x) & (!n_n5085) & (!n_n5081) & (!n_n5075)) + ((!x18x) & (x516x) & (!n_n5085) & (!n_n5081) & (!n_n5075)) + ((x18x) & (!x516x) & (!n_n5085) & (!n_n5081) & (!n_n5075)));
	assign x15618x = (((!n_n5086) & (!n_n5073) & (!n_n5079) & (!x209x) & (!x22088x)) + ((!n_n5086) & (!n_n5073) & (!n_n5079) & (x209x) & (!x22088x)) + ((!n_n5086) & (!n_n5073) & (!n_n5079) & (x209x) & (x22088x)) + ((!n_n5086) & (!n_n5073) & (n_n5079) & (!x209x) & (!x22088x)) + ((!n_n5086) & (!n_n5073) & (n_n5079) & (!x209x) & (x22088x)) + ((!n_n5086) & (!n_n5073) & (n_n5079) & (x209x) & (!x22088x)) + ((!n_n5086) & (!n_n5073) & (n_n5079) & (x209x) & (x22088x)) + ((!n_n5086) & (n_n5073) & (!n_n5079) & (!x209x) & (!x22088x)) + ((!n_n5086) & (n_n5073) & (!n_n5079) & (!x209x) & (x22088x)) + ((!n_n5086) & (n_n5073) & (!n_n5079) & (x209x) & (!x22088x)) + ((!n_n5086) & (n_n5073) & (!n_n5079) & (x209x) & (x22088x)) + ((!n_n5086) & (n_n5073) & (n_n5079) & (!x209x) & (!x22088x)) + ((!n_n5086) & (n_n5073) & (n_n5079) & (!x209x) & (x22088x)) + ((!n_n5086) & (n_n5073) & (n_n5079) & (x209x) & (!x22088x)) + ((!n_n5086) & (n_n5073) & (n_n5079) & (x209x) & (x22088x)) + ((n_n5086) & (!n_n5073) & (!n_n5079) & (!x209x) & (!x22088x)) + ((n_n5086) & (!n_n5073) & (!n_n5079) & (!x209x) & (x22088x)) + ((n_n5086) & (!n_n5073) & (!n_n5079) & (x209x) & (!x22088x)) + ((n_n5086) & (!n_n5073) & (!n_n5079) & (x209x) & (x22088x)) + ((n_n5086) & (!n_n5073) & (n_n5079) & (!x209x) & (!x22088x)) + ((n_n5086) & (!n_n5073) & (n_n5079) & (!x209x) & (x22088x)) + ((n_n5086) & (!n_n5073) & (n_n5079) & (x209x) & (!x22088x)) + ((n_n5086) & (!n_n5073) & (n_n5079) & (x209x) & (x22088x)) + ((n_n5086) & (n_n5073) & (!n_n5079) & (!x209x) & (!x22088x)) + ((n_n5086) & (n_n5073) & (!n_n5079) & (!x209x) & (x22088x)) + ((n_n5086) & (n_n5073) & (!n_n5079) & (x209x) & (!x22088x)) + ((n_n5086) & (n_n5073) & (!n_n5079) & (x209x) & (x22088x)) + ((n_n5086) & (n_n5073) & (n_n5079) & (!x209x) & (!x22088x)) + ((n_n5086) & (n_n5073) & (n_n5079) & (!x209x) & (x22088x)) + ((n_n5086) & (n_n5073) & (n_n5079) & (x209x) & (!x22088x)) + ((n_n5086) & (n_n5073) & (n_n5079) & (x209x) & (x22088x)));
	assign x22087x = (((!n_n5099) & (!n_n5101) & (!x344x) & (!x159x) & (!x143x)));
	assign x22086x = (((!n_n5109) & (!n_n5103) & (!n_n5104) & (!n_n5102)));
	assign x15626x = (((!i_9_) & (!n_n528) & (n_n532) & (n_n509) & (n_n130)) + ((!i_9_) & (n_n528) & (!n_n532) & (n_n509) & (n_n130)) + ((!i_9_) & (n_n528) & (n_n532) & (n_n509) & (n_n130)));
	assign x15638x = (((!i_9_) & (!x492x) & (!n_n195) & (!n_n5032) & (x265x)) + ((!i_9_) & (!x492x) & (!n_n195) & (n_n5032) & (!x265x)) + ((!i_9_) & (!x492x) & (!n_n195) & (n_n5032) & (x265x)) + ((!i_9_) & (!x492x) & (n_n195) & (!n_n5032) & (x265x)) + ((!i_9_) & (!x492x) & (n_n195) & (n_n5032) & (!x265x)) + ((!i_9_) & (!x492x) & (n_n195) & (n_n5032) & (x265x)) + ((!i_9_) & (x492x) & (!n_n195) & (!n_n5032) & (x265x)) + ((!i_9_) & (x492x) & (!n_n195) & (n_n5032) & (!x265x)) + ((!i_9_) & (x492x) & (!n_n195) & (n_n5032) & (x265x)) + ((!i_9_) & (x492x) & (n_n195) & (!n_n5032) & (x265x)) + ((!i_9_) & (x492x) & (n_n195) & (n_n5032) & (!x265x)) + ((!i_9_) & (x492x) & (n_n195) & (n_n5032) & (x265x)) + ((i_9_) & (!x492x) & (!n_n195) & (!n_n5032) & (x265x)) + ((i_9_) & (!x492x) & (!n_n195) & (n_n5032) & (!x265x)) + ((i_9_) & (!x492x) & (!n_n195) & (n_n5032) & (x265x)) + ((i_9_) & (!x492x) & (n_n195) & (!n_n5032) & (x265x)) + ((i_9_) & (!x492x) & (n_n195) & (n_n5032) & (!x265x)) + ((i_9_) & (!x492x) & (n_n195) & (n_n5032) & (x265x)) + ((i_9_) & (x492x) & (!n_n195) & (!n_n5032) & (x265x)) + ((i_9_) & (x492x) & (!n_n195) & (n_n5032) & (!x265x)) + ((i_9_) & (x492x) & (!n_n195) & (n_n5032) & (x265x)) + ((i_9_) & (x492x) & (n_n195) & (!n_n5032) & (!x265x)) + ((i_9_) & (x492x) & (n_n195) & (!n_n5032) & (x265x)) + ((i_9_) & (x492x) & (n_n195) & (n_n5032) & (!x265x)) + ((i_9_) & (x492x) & (n_n195) & (n_n5032) & (x265x)));
	assign x15639x = (((!n_n5034) & (!n_n5035) & (!n_n5036) & (!n_n5031) & (n_n5029)) + ((!n_n5034) & (!n_n5035) & (!n_n5036) & (n_n5031) & (!n_n5029)) + ((!n_n5034) & (!n_n5035) & (!n_n5036) & (n_n5031) & (n_n5029)) + ((!n_n5034) & (!n_n5035) & (n_n5036) & (!n_n5031) & (!n_n5029)) + ((!n_n5034) & (!n_n5035) & (n_n5036) & (!n_n5031) & (n_n5029)) + ((!n_n5034) & (!n_n5035) & (n_n5036) & (n_n5031) & (!n_n5029)) + ((!n_n5034) & (!n_n5035) & (n_n5036) & (n_n5031) & (n_n5029)) + ((!n_n5034) & (n_n5035) & (!n_n5036) & (!n_n5031) & (!n_n5029)) + ((!n_n5034) & (n_n5035) & (!n_n5036) & (!n_n5031) & (n_n5029)) + ((!n_n5034) & (n_n5035) & (!n_n5036) & (n_n5031) & (!n_n5029)) + ((!n_n5034) & (n_n5035) & (!n_n5036) & (n_n5031) & (n_n5029)) + ((!n_n5034) & (n_n5035) & (n_n5036) & (!n_n5031) & (!n_n5029)) + ((!n_n5034) & (n_n5035) & (n_n5036) & (!n_n5031) & (n_n5029)) + ((!n_n5034) & (n_n5035) & (n_n5036) & (n_n5031) & (!n_n5029)) + ((!n_n5034) & (n_n5035) & (n_n5036) & (n_n5031) & (n_n5029)) + ((n_n5034) & (!n_n5035) & (!n_n5036) & (!n_n5031) & (!n_n5029)) + ((n_n5034) & (!n_n5035) & (!n_n5036) & (!n_n5031) & (n_n5029)) + ((n_n5034) & (!n_n5035) & (!n_n5036) & (n_n5031) & (!n_n5029)) + ((n_n5034) & (!n_n5035) & (!n_n5036) & (n_n5031) & (n_n5029)) + ((n_n5034) & (!n_n5035) & (n_n5036) & (!n_n5031) & (!n_n5029)) + ((n_n5034) & (!n_n5035) & (n_n5036) & (!n_n5031) & (n_n5029)) + ((n_n5034) & (!n_n5035) & (n_n5036) & (n_n5031) & (!n_n5029)) + ((n_n5034) & (!n_n5035) & (n_n5036) & (n_n5031) & (n_n5029)) + ((n_n5034) & (n_n5035) & (!n_n5036) & (!n_n5031) & (!n_n5029)) + ((n_n5034) & (n_n5035) & (!n_n5036) & (!n_n5031) & (n_n5029)) + ((n_n5034) & (n_n5035) & (!n_n5036) & (n_n5031) & (!n_n5029)) + ((n_n5034) & (n_n5035) & (!n_n5036) & (n_n5031) & (n_n5029)) + ((n_n5034) & (n_n5035) & (n_n5036) & (!n_n5031) & (!n_n5029)) + ((n_n5034) & (n_n5035) & (n_n5036) & (!n_n5031) & (n_n5029)) + ((n_n5034) & (n_n5035) & (n_n5036) & (n_n5031) & (!n_n5029)) + ((n_n5034) & (n_n5035) & (n_n5036) & (n_n5031) & (n_n5029)));
	assign x22224x = (((!n_n4464) & (!n_n4471) & (!n_n4472) & (!n_n4469)));
	assign x16182x = (((!i_9_) & (!n_n528) & (n_n260) & (n_n491) & (x23x)) + ((!i_9_) & (n_n528) & (n_n260) & (n_n491) & (!x23x)) + ((!i_9_) & (n_n528) & (n_n260) & (n_n491) & (x23x)) + ((i_9_) & (!n_n528) & (n_n260) & (n_n491) & (x23x)) + ((i_9_) & (n_n528) & (n_n260) & (n_n491) & (x23x)));
	assign n_n1854 = (((!n_n4901) & (!x96x) & (!x352x) & (!x227x) & (x16182x)) + ((!n_n4901) & (!x96x) & (!x352x) & (x227x) & (!x16182x)) + ((!n_n4901) & (!x96x) & (!x352x) & (x227x) & (x16182x)) + ((!n_n4901) & (!x96x) & (x352x) & (!x227x) & (!x16182x)) + ((!n_n4901) & (!x96x) & (x352x) & (!x227x) & (x16182x)) + ((!n_n4901) & (!x96x) & (x352x) & (x227x) & (!x16182x)) + ((!n_n4901) & (!x96x) & (x352x) & (x227x) & (x16182x)) + ((!n_n4901) & (x96x) & (!x352x) & (!x227x) & (!x16182x)) + ((!n_n4901) & (x96x) & (!x352x) & (!x227x) & (x16182x)) + ((!n_n4901) & (x96x) & (!x352x) & (x227x) & (!x16182x)) + ((!n_n4901) & (x96x) & (!x352x) & (x227x) & (x16182x)) + ((!n_n4901) & (x96x) & (x352x) & (!x227x) & (!x16182x)) + ((!n_n4901) & (x96x) & (x352x) & (!x227x) & (x16182x)) + ((!n_n4901) & (x96x) & (x352x) & (x227x) & (!x16182x)) + ((!n_n4901) & (x96x) & (x352x) & (x227x) & (x16182x)) + ((n_n4901) & (!x96x) & (!x352x) & (!x227x) & (!x16182x)) + ((n_n4901) & (!x96x) & (!x352x) & (!x227x) & (x16182x)) + ((n_n4901) & (!x96x) & (!x352x) & (x227x) & (!x16182x)) + ((n_n4901) & (!x96x) & (!x352x) & (x227x) & (x16182x)) + ((n_n4901) & (!x96x) & (x352x) & (!x227x) & (!x16182x)) + ((n_n4901) & (!x96x) & (x352x) & (!x227x) & (x16182x)) + ((n_n4901) & (!x96x) & (x352x) & (x227x) & (!x16182x)) + ((n_n4901) & (!x96x) & (x352x) & (x227x) & (x16182x)) + ((n_n4901) & (x96x) & (!x352x) & (!x227x) & (!x16182x)) + ((n_n4901) & (x96x) & (!x352x) & (!x227x) & (x16182x)) + ((n_n4901) & (x96x) & (!x352x) & (x227x) & (!x16182x)) + ((n_n4901) & (x96x) & (!x352x) & (x227x) & (x16182x)) + ((n_n4901) & (x96x) & (x352x) & (!x227x) & (!x16182x)) + ((n_n4901) & (x96x) & (x352x) & (!x227x) & (x16182x)) + ((n_n4901) & (x96x) & (x352x) & (x227x) & (!x16182x)) + ((n_n4901) & (x96x) & (x352x) & (x227x) & (x16182x)));
	assign x22076x = (((!n_n5181) & (!n_n5184) & (!n_n5185) & (!n_n5183)));
	assign x22072x = (((!n_n4749) & (!n_n4747) & (!n_n4755) & (!n_n4752)));
	assign x22177x = (((!n_n4718) & (!n_n4717) & (!n_n4715) & (!n_n4714)));
	assign x16248x = (((!n_n5173) & (!n_n5172) & (!n_n5168) & (n_n5169)) + ((!n_n5173) & (!n_n5172) & (n_n5168) & (!n_n5169)) + ((!n_n5173) & (!n_n5172) & (n_n5168) & (n_n5169)) + ((!n_n5173) & (n_n5172) & (!n_n5168) & (!n_n5169)) + ((!n_n5173) & (n_n5172) & (!n_n5168) & (n_n5169)) + ((!n_n5173) & (n_n5172) & (n_n5168) & (!n_n5169)) + ((!n_n5173) & (n_n5172) & (n_n5168) & (n_n5169)) + ((n_n5173) & (!n_n5172) & (!n_n5168) & (!n_n5169)) + ((n_n5173) & (!n_n5172) & (!n_n5168) & (n_n5169)) + ((n_n5173) & (!n_n5172) & (n_n5168) & (!n_n5169)) + ((n_n5173) & (!n_n5172) & (n_n5168) & (n_n5169)) + ((n_n5173) & (n_n5172) & (!n_n5168) & (!n_n5169)) + ((n_n5173) & (n_n5172) & (!n_n5168) & (n_n5169)) + ((n_n5173) & (n_n5172) & (n_n5168) & (!n_n5169)) + ((n_n5173) & (n_n5172) & (n_n5168) & (n_n5169)));
	assign n_n1840 = (((!n_n5082) & (!n_n5079) & (!x123x) & (!n_n1952) & (x209x)) + ((!n_n5082) & (!n_n5079) & (!x123x) & (n_n1952) & (!x209x)) + ((!n_n5082) & (!n_n5079) & (!x123x) & (n_n1952) & (x209x)) + ((!n_n5082) & (!n_n5079) & (x123x) & (!n_n1952) & (!x209x)) + ((!n_n5082) & (!n_n5079) & (x123x) & (!n_n1952) & (x209x)) + ((!n_n5082) & (!n_n5079) & (x123x) & (n_n1952) & (!x209x)) + ((!n_n5082) & (!n_n5079) & (x123x) & (n_n1952) & (x209x)) + ((!n_n5082) & (n_n5079) & (!x123x) & (!n_n1952) & (!x209x)) + ((!n_n5082) & (n_n5079) & (!x123x) & (!n_n1952) & (x209x)) + ((!n_n5082) & (n_n5079) & (!x123x) & (n_n1952) & (!x209x)) + ((!n_n5082) & (n_n5079) & (!x123x) & (n_n1952) & (x209x)) + ((!n_n5082) & (n_n5079) & (x123x) & (!n_n1952) & (!x209x)) + ((!n_n5082) & (n_n5079) & (x123x) & (!n_n1952) & (x209x)) + ((!n_n5082) & (n_n5079) & (x123x) & (n_n1952) & (!x209x)) + ((!n_n5082) & (n_n5079) & (x123x) & (n_n1952) & (x209x)) + ((n_n5082) & (!n_n5079) & (!x123x) & (!n_n1952) & (!x209x)) + ((n_n5082) & (!n_n5079) & (!x123x) & (!n_n1952) & (x209x)) + ((n_n5082) & (!n_n5079) & (!x123x) & (n_n1952) & (!x209x)) + ((n_n5082) & (!n_n5079) & (!x123x) & (n_n1952) & (x209x)) + ((n_n5082) & (!n_n5079) & (x123x) & (!n_n1952) & (!x209x)) + ((n_n5082) & (!n_n5079) & (x123x) & (!n_n1952) & (x209x)) + ((n_n5082) & (!n_n5079) & (x123x) & (n_n1952) & (!x209x)) + ((n_n5082) & (!n_n5079) & (x123x) & (n_n1952) & (x209x)) + ((n_n5082) & (n_n5079) & (!x123x) & (!n_n1952) & (!x209x)) + ((n_n5082) & (n_n5079) & (!x123x) & (!n_n1952) & (x209x)) + ((n_n5082) & (n_n5079) & (!x123x) & (n_n1952) & (!x209x)) + ((n_n5082) & (n_n5079) & (!x123x) & (n_n1952) & (x209x)) + ((n_n5082) & (n_n5079) & (x123x) & (!n_n1952) & (!x209x)) + ((n_n5082) & (n_n5079) & (x123x) & (!n_n1952) & (x209x)) + ((n_n5082) & (n_n5079) & (x123x) & (n_n1952) & (!x209x)) + ((n_n5082) & (n_n5079) & (x123x) & (n_n1952) & (x209x)));
	assign x22066x = (((!n_n5092) & (!n_n5093) & (!n_n5089) & (!n_n5086)));
	assign n_n1839 = (((!n_n5091) & (!n_n5088) & (!n_n5090) & (!x279x) & (!x22066x)) + ((!n_n5091) & (!n_n5088) & (!n_n5090) & (x279x) & (!x22066x)) + ((!n_n5091) & (!n_n5088) & (!n_n5090) & (x279x) & (x22066x)) + ((!n_n5091) & (!n_n5088) & (n_n5090) & (!x279x) & (!x22066x)) + ((!n_n5091) & (!n_n5088) & (n_n5090) & (!x279x) & (x22066x)) + ((!n_n5091) & (!n_n5088) & (n_n5090) & (x279x) & (!x22066x)) + ((!n_n5091) & (!n_n5088) & (n_n5090) & (x279x) & (x22066x)) + ((!n_n5091) & (n_n5088) & (!n_n5090) & (!x279x) & (!x22066x)) + ((!n_n5091) & (n_n5088) & (!n_n5090) & (!x279x) & (x22066x)) + ((!n_n5091) & (n_n5088) & (!n_n5090) & (x279x) & (!x22066x)) + ((!n_n5091) & (n_n5088) & (!n_n5090) & (x279x) & (x22066x)) + ((!n_n5091) & (n_n5088) & (n_n5090) & (!x279x) & (!x22066x)) + ((!n_n5091) & (n_n5088) & (n_n5090) & (!x279x) & (x22066x)) + ((!n_n5091) & (n_n5088) & (n_n5090) & (x279x) & (!x22066x)) + ((!n_n5091) & (n_n5088) & (n_n5090) & (x279x) & (x22066x)) + ((n_n5091) & (!n_n5088) & (!n_n5090) & (!x279x) & (!x22066x)) + ((n_n5091) & (!n_n5088) & (!n_n5090) & (!x279x) & (x22066x)) + ((n_n5091) & (!n_n5088) & (!n_n5090) & (x279x) & (!x22066x)) + ((n_n5091) & (!n_n5088) & (!n_n5090) & (x279x) & (x22066x)) + ((n_n5091) & (!n_n5088) & (n_n5090) & (!x279x) & (!x22066x)) + ((n_n5091) & (!n_n5088) & (n_n5090) & (!x279x) & (x22066x)) + ((n_n5091) & (!n_n5088) & (n_n5090) & (x279x) & (!x22066x)) + ((n_n5091) & (!n_n5088) & (n_n5090) & (x279x) & (x22066x)) + ((n_n5091) & (n_n5088) & (!n_n5090) & (!x279x) & (!x22066x)) + ((n_n5091) & (n_n5088) & (!n_n5090) & (!x279x) & (x22066x)) + ((n_n5091) & (n_n5088) & (!n_n5090) & (x279x) & (!x22066x)) + ((n_n5091) & (n_n5088) & (!n_n5090) & (x279x) & (x22066x)) + ((n_n5091) & (n_n5088) & (n_n5090) & (!x279x) & (!x22066x)) + ((n_n5091) & (n_n5088) & (n_n5090) & (!x279x) & (x22066x)) + ((n_n5091) & (n_n5088) & (n_n5090) & (x279x) & (!x22066x)) + ((n_n5091) & (n_n5088) & (n_n5090) & (x279x) & (x22066x)));
	assign x15956x = (((!n_n5064) & (!n_n5057) & (!n_n5058) & (!n_n5067) & (n_n5065)) + ((!n_n5064) & (!n_n5057) & (!n_n5058) & (n_n5067) & (!n_n5065)) + ((!n_n5064) & (!n_n5057) & (!n_n5058) & (n_n5067) & (n_n5065)) + ((!n_n5064) & (!n_n5057) & (n_n5058) & (!n_n5067) & (!n_n5065)) + ((!n_n5064) & (!n_n5057) & (n_n5058) & (!n_n5067) & (n_n5065)) + ((!n_n5064) & (!n_n5057) & (n_n5058) & (n_n5067) & (!n_n5065)) + ((!n_n5064) & (!n_n5057) & (n_n5058) & (n_n5067) & (n_n5065)) + ((!n_n5064) & (n_n5057) & (!n_n5058) & (!n_n5067) & (!n_n5065)) + ((!n_n5064) & (n_n5057) & (!n_n5058) & (!n_n5067) & (n_n5065)) + ((!n_n5064) & (n_n5057) & (!n_n5058) & (n_n5067) & (!n_n5065)) + ((!n_n5064) & (n_n5057) & (!n_n5058) & (n_n5067) & (n_n5065)) + ((!n_n5064) & (n_n5057) & (n_n5058) & (!n_n5067) & (!n_n5065)) + ((!n_n5064) & (n_n5057) & (n_n5058) & (!n_n5067) & (n_n5065)) + ((!n_n5064) & (n_n5057) & (n_n5058) & (n_n5067) & (!n_n5065)) + ((!n_n5064) & (n_n5057) & (n_n5058) & (n_n5067) & (n_n5065)) + ((n_n5064) & (!n_n5057) & (!n_n5058) & (!n_n5067) & (!n_n5065)) + ((n_n5064) & (!n_n5057) & (!n_n5058) & (!n_n5067) & (n_n5065)) + ((n_n5064) & (!n_n5057) & (!n_n5058) & (n_n5067) & (!n_n5065)) + ((n_n5064) & (!n_n5057) & (!n_n5058) & (n_n5067) & (n_n5065)) + ((n_n5064) & (!n_n5057) & (n_n5058) & (!n_n5067) & (!n_n5065)) + ((n_n5064) & (!n_n5057) & (n_n5058) & (!n_n5067) & (n_n5065)) + ((n_n5064) & (!n_n5057) & (n_n5058) & (n_n5067) & (!n_n5065)) + ((n_n5064) & (!n_n5057) & (n_n5058) & (n_n5067) & (n_n5065)) + ((n_n5064) & (n_n5057) & (!n_n5058) & (!n_n5067) & (!n_n5065)) + ((n_n5064) & (n_n5057) & (!n_n5058) & (!n_n5067) & (n_n5065)) + ((n_n5064) & (n_n5057) & (!n_n5058) & (n_n5067) & (!n_n5065)) + ((n_n5064) & (n_n5057) & (!n_n5058) & (n_n5067) & (n_n5065)) + ((n_n5064) & (n_n5057) & (n_n5058) & (!n_n5067) & (!n_n5065)) + ((n_n5064) & (n_n5057) & (n_n5058) & (!n_n5067) & (n_n5065)) + ((n_n5064) & (n_n5057) & (n_n5058) & (n_n5067) & (!n_n5065)) + ((n_n5064) & (n_n5057) & (n_n5058) & (n_n5067) & (n_n5065)));
	assign x15957x = (((!n_n5060) & (!n_n5054) & (!x160x) & (x15956x)) + ((!n_n5060) & (!n_n5054) & (x160x) & (!x15956x)) + ((!n_n5060) & (!n_n5054) & (x160x) & (x15956x)) + ((!n_n5060) & (n_n5054) & (!x160x) & (!x15956x)) + ((!n_n5060) & (n_n5054) & (!x160x) & (x15956x)) + ((!n_n5060) & (n_n5054) & (x160x) & (!x15956x)) + ((!n_n5060) & (n_n5054) & (x160x) & (x15956x)) + ((n_n5060) & (!n_n5054) & (!x160x) & (!x15956x)) + ((n_n5060) & (!n_n5054) & (!x160x) & (x15956x)) + ((n_n5060) & (!n_n5054) & (x160x) & (!x15956x)) + ((n_n5060) & (!n_n5054) & (x160x) & (x15956x)) + ((n_n5060) & (n_n5054) & (!x160x) & (!x15956x)) + ((n_n5060) & (n_n5054) & (!x160x) & (x15956x)) + ((n_n5060) & (n_n5054) & (x160x) & (!x15956x)) + ((n_n5060) & (n_n5054) & (x160x) & (x15956x)));
	assign n_n1801 = (((!n_n1840) & (!n_n1839) & (x15957x)) + ((!n_n1840) & (n_n1839) & (!x15957x)) + ((!n_n1840) & (n_n1839) & (x15957x)) + ((n_n1840) & (!n_n1839) & (!x15957x)) + ((n_n1840) & (!n_n1839) & (x15957x)) + ((n_n1840) & (n_n1839) & (!x15957x)) + ((n_n1840) & (n_n1839) & (x15957x)));
	assign x15962x = (((!n_n5123) & (!n_n5124) & (!n_n5114) & (n_n5126)) + ((!n_n5123) & (!n_n5124) & (n_n5114) & (!n_n5126)) + ((!n_n5123) & (!n_n5124) & (n_n5114) & (n_n5126)) + ((!n_n5123) & (n_n5124) & (!n_n5114) & (!n_n5126)) + ((!n_n5123) & (n_n5124) & (!n_n5114) & (n_n5126)) + ((!n_n5123) & (n_n5124) & (n_n5114) & (!n_n5126)) + ((!n_n5123) & (n_n5124) & (n_n5114) & (n_n5126)) + ((n_n5123) & (!n_n5124) & (!n_n5114) & (!n_n5126)) + ((n_n5123) & (!n_n5124) & (!n_n5114) & (n_n5126)) + ((n_n5123) & (!n_n5124) & (n_n5114) & (!n_n5126)) + ((n_n5123) & (!n_n5124) & (n_n5114) & (n_n5126)) + ((n_n5123) & (n_n5124) & (!n_n5114) & (!n_n5126)) + ((n_n5123) & (n_n5124) & (!n_n5114) & (n_n5126)) + ((n_n5123) & (n_n5124) & (n_n5114) & (!n_n5126)) + ((n_n5123) & (n_n5124) & (n_n5114) & (n_n5126)));
	assign x15963x = (((!n_n5115) & (!n_n5121) & (!n_n5122) & (!n_n5128) & (n_n5118)) + ((!n_n5115) & (!n_n5121) & (!n_n5122) & (n_n5128) & (!n_n5118)) + ((!n_n5115) & (!n_n5121) & (!n_n5122) & (n_n5128) & (n_n5118)) + ((!n_n5115) & (!n_n5121) & (n_n5122) & (!n_n5128) & (!n_n5118)) + ((!n_n5115) & (!n_n5121) & (n_n5122) & (!n_n5128) & (n_n5118)) + ((!n_n5115) & (!n_n5121) & (n_n5122) & (n_n5128) & (!n_n5118)) + ((!n_n5115) & (!n_n5121) & (n_n5122) & (n_n5128) & (n_n5118)) + ((!n_n5115) & (n_n5121) & (!n_n5122) & (!n_n5128) & (!n_n5118)) + ((!n_n5115) & (n_n5121) & (!n_n5122) & (!n_n5128) & (n_n5118)) + ((!n_n5115) & (n_n5121) & (!n_n5122) & (n_n5128) & (!n_n5118)) + ((!n_n5115) & (n_n5121) & (!n_n5122) & (n_n5128) & (n_n5118)) + ((!n_n5115) & (n_n5121) & (n_n5122) & (!n_n5128) & (!n_n5118)) + ((!n_n5115) & (n_n5121) & (n_n5122) & (!n_n5128) & (n_n5118)) + ((!n_n5115) & (n_n5121) & (n_n5122) & (n_n5128) & (!n_n5118)) + ((!n_n5115) & (n_n5121) & (n_n5122) & (n_n5128) & (n_n5118)) + ((n_n5115) & (!n_n5121) & (!n_n5122) & (!n_n5128) & (!n_n5118)) + ((n_n5115) & (!n_n5121) & (!n_n5122) & (!n_n5128) & (n_n5118)) + ((n_n5115) & (!n_n5121) & (!n_n5122) & (n_n5128) & (!n_n5118)) + ((n_n5115) & (!n_n5121) & (!n_n5122) & (n_n5128) & (n_n5118)) + ((n_n5115) & (!n_n5121) & (n_n5122) & (!n_n5128) & (!n_n5118)) + ((n_n5115) & (!n_n5121) & (n_n5122) & (!n_n5128) & (n_n5118)) + ((n_n5115) & (!n_n5121) & (n_n5122) & (n_n5128) & (!n_n5118)) + ((n_n5115) & (!n_n5121) & (n_n5122) & (n_n5128) & (n_n5118)) + ((n_n5115) & (n_n5121) & (!n_n5122) & (!n_n5128) & (!n_n5118)) + ((n_n5115) & (n_n5121) & (!n_n5122) & (!n_n5128) & (n_n5118)) + ((n_n5115) & (n_n5121) & (!n_n5122) & (n_n5128) & (!n_n5118)) + ((n_n5115) & (n_n5121) & (!n_n5122) & (n_n5128) & (n_n5118)) + ((n_n5115) & (n_n5121) & (n_n5122) & (!n_n5128) & (!n_n5118)) + ((n_n5115) & (n_n5121) & (n_n5122) & (!n_n5128) & (n_n5118)) + ((n_n5115) & (n_n5121) & (n_n5122) & (n_n5128) & (!n_n5118)) + ((n_n5115) & (n_n5121) & (n_n5122) & (n_n5128) & (n_n5118)));
	assign x15967x = (((!n_n5112) & (!n_n5109) & (!n_n5110) & (n_n5107)) + ((!n_n5112) & (!n_n5109) & (n_n5110) & (!n_n5107)) + ((!n_n5112) & (!n_n5109) & (n_n5110) & (n_n5107)) + ((!n_n5112) & (n_n5109) & (!n_n5110) & (!n_n5107)) + ((!n_n5112) & (n_n5109) & (!n_n5110) & (n_n5107)) + ((!n_n5112) & (n_n5109) & (n_n5110) & (!n_n5107)) + ((!n_n5112) & (n_n5109) & (n_n5110) & (n_n5107)) + ((n_n5112) & (!n_n5109) & (!n_n5110) & (!n_n5107)) + ((n_n5112) & (!n_n5109) & (!n_n5110) & (n_n5107)) + ((n_n5112) & (!n_n5109) & (n_n5110) & (!n_n5107)) + ((n_n5112) & (!n_n5109) & (n_n5110) & (n_n5107)) + ((n_n5112) & (n_n5109) & (!n_n5110) & (!n_n5107)) + ((n_n5112) & (n_n5109) & (!n_n5110) & (n_n5107)) + ((n_n5112) & (n_n5109) & (n_n5110) & (!n_n5107)) + ((n_n5112) & (n_n5109) & (n_n5110) & (n_n5107)));
	assign x15968x = (((!n_n5099) & (!n_n5101) & (!n_n5113) & (!n_n5104) & (n_n5106)) + ((!n_n5099) & (!n_n5101) & (!n_n5113) & (n_n5104) & (!n_n5106)) + ((!n_n5099) & (!n_n5101) & (!n_n5113) & (n_n5104) & (n_n5106)) + ((!n_n5099) & (!n_n5101) & (n_n5113) & (!n_n5104) & (!n_n5106)) + ((!n_n5099) & (!n_n5101) & (n_n5113) & (!n_n5104) & (n_n5106)) + ((!n_n5099) & (!n_n5101) & (n_n5113) & (n_n5104) & (!n_n5106)) + ((!n_n5099) & (!n_n5101) & (n_n5113) & (n_n5104) & (n_n5106)) + ((!n_n5099) & (n_n5101) & (!n_n5113) & (!n_n5104) & (!n_n5106)) + ((!n_n5099) & (n_n5101) & (!n_n5113) & (!n_n5104) & (n_n5106)) + ((!n_n5099) & (n_n5101) & (!n_n5113) & (n_n5104) & (!n_n5106)) + ((!n_n5099) & (n_n5101) & (!n_n5113) & (n_n5104) & (n_n5106)) + ((!n_n5099) & (n_n5101) & (n_n5113) & (!n_n5104) & (!n_n5106)) + ((!n_n5099) & (n_n5101) & (n_n5113) & (!n_n5104) & (n_n5106)) + ((!n_n5099) & (n_n5101) & (n_n5113) & (n_n5104) & (!n_n5106)) + ((!n_n5099) & (n_n5101) & (n_n5113) & (n_n5104) & (n_n5106)) + ((n_n5099) & (!n_n5101) & (!n_n5113) & (!n_n5104) & (!n_n5106)) + ((n_n5099) & (!n_n5101) & (!n_n5113) & (!n_n5104) & (n_n5106)) + ((n_n5099) & (!n_n5101) & (!n_n5113) & (n_n5104) & (!n_n5106)) + ((n_n5099) & (!n_n5101) & (!n_n5113) & (n_n5104) & (n_n5106)) + ((n_n5099) & (!n_n5101) & (n_n5113) & (!n_n5104) & (!n_n5106)) + ((n_n5099) & (!n_n5101) & (n_n5113) & (!n_n5104) & (n_n5106)) + ((n_n5099) & (!n_n5101) & (n_n5113) & (n_n5104) & (!n_n5106)) + ((n_n5099) & (!n_n5101) & (n_n5113) & (n_n5104) & (n_n5106)) + ((n_n5099) & (n_n5101) & (!n_n5113) & (!n_n5104) & (!n_n5106)) + ((n_n5099) & (n_n5101) & (!n_n5113) & (!n_n5104) & (n_n5106)) + ((n_n5099) & (n_n5101) & (!n_n5113) & (n_n5104) & (!n_n5106)) + ((n_n5099) & (n_n5101) & (!n_n5113) & (n_n5104) & (n_n5106)) + ((n_n5099) & (n_n5101) & (n_n5113) & (!n_n5104) & (!n_n5106)) + ((n_n5099) & (n_n5101) & (n_n5113) & (!n_n5104) & (n_n5106)) + ((n_n5099) & (n_n5101) & (n_n5113) & (n_n5104) & (!n_n5106)) + ((n_n5099) & (n_n5101) & (n_n5113) & (n_n5104) & (n_n5106)));
	assign x15972x = (((!n_n522) & (!x12x) & (!n_n500) & (!n_n530) & (n_n1162)) + ((!n_n522) & (!x12x) & (!n_n500) & (n_n530) & (n_n1162)) + ((!n_n522) & (!x12x) & (n_n500) & (!n_n530) & (n_n1162)) + ((!n_n522) & (!x12x) & (n_n500) & (n_n530) & (n_n1162)) + ((!n_n522) & (x12x) & (!n_n500) & (!n_n530) & (n_n1162)) + ((!n_n522) & (x12x) & (!n_n500) & (n_n530) & (n_n1162)) + ((!n_n522) & (x12x) & (n_n500) & (!n_n530) & (n_n1162)) + ((!n_n522) & (x12x) & (n_n500) & (n_n530) & (!n_n1162)) + ((!n_n522) & (x12x) & (n_n500) & (n_n530) & (n_n1162)) + ((n_n522) & (!x12x) & (!n_n500) & (!n_n530) & (n_n1162)) + ((n_n522) & (!x12x) & (!n_n500) & (n_n530) & (n_n1162)) + ((n_n522) & (!x12x) & (n_n500) & (!n_n530) & (n_n1162)) + ((n_n522) & (!x12x) & (n_n500) & (n_n530) & (n_n1162)) + ((n_n522) & (x12x) & (!n_n500) & (!n_n530) & (n_n1162)) + ((n_n522) & (x12x) & (!n_n500) & (n_n530) & (n_n1162)) + ((n_n522) & (x12x) & (n_n500) & (!n_n530) & (!n_n1162)) + ((n_n522) & (x12x) & (n_n500) & (!n_n530) & (n_n1162)) + ((n_n522) & (x12x) & (n_n500) & (n_n530) & (!n_n1162)) + ((n_n522) & (x12x) & (n_n500) & (n_n530) & (n_n1162)));
	assign x15973x = (((!n_n5130) & (!n_n5129) & (!x422x) & (x15972x)) + ((!n_n5130) & (!n_n5129) & (x422x) & (!x15972x)) + ((!n_n5130) & (!n_n5129) & (x422x) & (x15972x)) + ((!n_n5130) & (n_n5129) & (!x422x) & (!x15972x)) + ((!n_n5130) & (n_n5129) & (!x422x) & (x15972x)) + ((!n_n5130) & (n_n5129) & (x422x) & (!x15972x)) + ((!n_n5130) & (n_n5129) & (x422x) & (x15972x)) + ((n_n5130) & (!n_n5129) & (!x422x) & (!x15972x)) + ((n_n5130) & (!n_n5129) & (!x422x) & (x15972x)) + ((n_n5130) & (!n_n5129) & (x422x) & (!x15972x)) + ((n_n5130) & (!n_n5129) & (x422x) & (x15972x)) + ((n_n5130) & (n_n5129) & (!x422x) & (!x15972x)) + ((n_n5130) & (n_n5129) & (!x422x) & (x15972x)) + ((n_n5130) & (n_n5129) & (x422x) & (!x15972x)) + ((n_n5130) & (n_n5129) & (x422x) & (x15972x)));
	assign n_n1800 = (((!x15962x) & (!x15963x) & (!x15967x) & (!x15968x) & (x15973x)) + ((!x15962x) & (!x15963x) & (!x15967x) & (x15968x) & (!x15973x)) + ((!x15962x) & (!x15963x) & (!x15967x) & (x15968x) & (x15973x)) + ((!x15962x) & (!x15963x) & (x15967x) & (!x15968x) & (!x15973x)) + ((!x15962x) & (!x15963x) & (x15967x) & (!x15968x) & (x15973x)) + ((!x15962x) & (!x15963x) & (x15967x) & (x15968x) & (!x15973x)) + ((!x15962x) & (!x15963x) & (x15967x) & (x15968x) & (x15973x)) + ((!x15962x) & (x15963x) & (!x15967x) & (!x15968x) & (!x15973x)) + ((!x15962x) & (x15963x) & (!x15967x) & (!x15968x) & (x15973x)) + ((!x15962x) & (x15963x) & (!x15967x) & (x15968x) & (!x15973x)) + ((!x15962x) & (x15963x) & (!x15967x) & (x15968x) & (x15973x)) + ((!x15962x) & (x15963x) & (x15967x) & (!x15968x) & (!x15973x)) + ((!x15962x) & (x15963x) & (x15967x) & (!x15968x) & (x15973x)) + ((!x15962x) & (x15963x) & (x15967x) & (x15968x) & (!x15973x)) + ((!x15962x) & (x15963x) & (x15967x) & (x15968x) & (x15973x)) + ((x15962x) & (!x15963x) & (!x15967x) & (!x15968x) & (!x15973x)) + ((x15962x) & (!x15963x) & (!x15967x) & (!x15968x) & (x15973x)) + ((x15962x) & (!x15963x) & (!x15967x) & (x15968x) & (!x15973x)) + ((x15962x) & (!x15963x) & (!x15967x) & (x15968x) & (x15973x)) + ((x15962x) & (!x15963x) & (x15967x) & (!x15968x) & (!x15973x)) + ((x15962x) & (!x15963x) & (x15967x) & (!x15968x) & (x15973x)) + ((x15962x) & (!x15963x) & (x15967x) & (x15968x) & (!x15973x)) + ((x15962x) & (!x15963x) & (x15967x) & (x15968x) & (x15973x)) + ((x15962x) & (x15963x) & (!x15967x) & (!x15968x) & (!x15973x)) + ((x15962x) & (x15963x) & (!x15967x) & (!x15968x) & (x15973x)) + ((x15962x) & (x15963x) & (!x15967x) & (x15968x) & (!x15973x)) + ((x15962x) & (x15963x) & (!x15967x) & (x15968x) & (x15973x)) + ((x15962x) & (x15963x) & (x15967x) & (!x15968x) & (!x15973x)) + ((x15962x) & (x15963x) & (x15967x) & (!x15968x) & (x15973x)) + ((x15962x) & (x15963x) & (x15967x) & (x15968x) & (!x15973x)) + ((x15962x) & (x15963x) & (x15967x) & (x15968x) & (x15973x)));
	assign x15983x = (((!n_n5026) & (!n_n5014) & (!n_n5015) & (!n_n5020) & (n_n5016)) + ((!n_n5026) & (!n_n5014) & (!n_n5015) & (n_n5020) & (!n_n5016)) + ((!n_n5026) & (!n_n5014) & (!n_n5015) & (n_n5020) & (n_n5016)) + ((!n_n5026) & (!n_n5014) & (n_n5015) & (!n_n5020) & (!n_n5016)) + ((!n_n5026) & (!n_n5014) & (n_n5015) & (!n_n5020) & (n_n5016)) + ((!n_n5026) & (!n_n5014) & (n_n5015) & (n_n5020) & (!n_n5016)) + ((!n_n5026) & (!n_n5014) & (n_n5015) & (n_n5020) & (n_n5016)) + ((!n_n5026) & (n_n5014) & (!n_n5015) & (!n_n5020) & (!n_n5016)) + ((!n_n5026) & (n_n5014) & (!n_n5015) & (!n_n5020) & (n_n5016)) + ((!n_n5026) & (n_n5014) & (!n_n5015) & (n_n5020) & (!n_n5016)) + ((!n_n5026) & (n_n5014) & (!n_n5015) & (n_n5020) & (n_n5016)) + ((!n_n5026) & (n_n5014) & (n_n5015) & (!n_n5020) & (!n_n5016)) + ((!n_n5026) & (n_n5014) & (n_n5015) & (!n_n5020) & (n_n5016)) + ((!n_n5026) & (n_n5014) & (n_n5015) & (n_n5020) & (!n_n5016)) + ((!n_n5026) & (n_n5014) & (n_n5015) & (n_n5020) & (n_n5016)) + ((n_n5026) & (!n_n5014) & (!n_n5015) & (!n_n5020) & (!n_n5016)) + ((n_n5026) & (!n_n5014) & (!n_n5015) & (!n_n5020) & (n_n5016)) + ((n_n5026) & (!n_n5014) & (!n_n5015) & (n_n5020) & (!n_n5016)) + ((n_n5026) & (!n_n5014) & (!n_n5015) & (n_n5020) & (n_n5016)) + ((n_n5026) & (!n_n5014) & (n_n5015) & (!n_n5020) & (!n_n5016)) + ((n_n5026) & (!n_n5014) & (n_n5015) & (!n_n5020) & (n_n5016)) + ((n_n5026) & (!n_n5014) & (n_n5015) & (n_n5020) & (!n_n5016)) + ((n_n5026) & (!n_n5014) & (n_n5015) & (n_n5020) & (n_n5016)) + ((n_n5026) & (n_n5014) & (!n_n5015) & (!n_n5020) & (!n_n5016)) + ((n_n5026) & (n_n5014) & (!n_n5015) & (!n_n5020) & (n_n5016)) + ((n_n5026) & (n_n5014) & (!n_n5015) & (n_n5020) & (!n_n5016)) + ((n_n5026) & (n_n5014) & (!n_n5015) & (n_n5020) & (n_n5016)) + ((n_n5026) & (n_n5014) & (n_n5015) & (!n_n5020) & (!n_n5016)) + ((n_n5026) & (n_n5014) & (n_n5015) & (!n_n5020) & (n_n5016)) + ((n_n5026) & (n_n5014) & (n_n5015) & (n_n5020) & (!n_n5016)) + ((n_n5026) & (n_n5014) & (n_n5015) & (n_n5020) & (n_n5016)));
	assign x12784x = (((!n_n325) & (!n_n535) & (!x23x) & (!n_n4712) & (x30x)) + ((!n_n325) & (!n_n535) & (!x23x) & (n_n4712) & (!x30x)) + ((!n_n325) & (!n_n535) & (!x23x) & (n_n4712) & (x30x)) + ((!n_n325) & (!n_n535) & (x23x) & (!n_n4712) & (x30x)) + ((!n_n325) & (!n_n535) & (x23x) & (n_n4712) & (!x30x)) + ((!n_n325) & (!n_n535) & (x23x) & (n_n4712) & (x30x)) + ((!n_n325) & (n_n535) & (!x23x) & (!n_n4712) & (x30x)) + ((!n_n325) & (n_n535) & (!x23x) & (n_n4712) & (!x30x)) + ((!n_n325) & (n_n535) & (!x23x) & (n_n4712) & (x30x)) + ((!n_n325) & (n_n535) & (x23x) & (!n_n4712) & (x30x)) + ((!n_n325) & (n_n535) & (x23x) & (n_n4712) & (!x30x)) + ((!n_n325) & (n_n535) & (x23x) & (n_n4712) & (x30x)) + ((n_n325) & (!n_n535) & (!x23x) & (!n_n4712) & (x30x)) + ((n_n325) & (!n_n535) & (!x23x) & (n_n4712) & (!x30x)) + ((n_n325) & (!n_n535) & (!x23x) & (n_n4712) & (x30x)) + ((n_n325) & (!n_n535) & (x23x) & (!n_n4712) & (x30x)) + ((n_n325) & (!n_n535) & (x23x) & (n_n4712) & (!x30x)) + ((n_n325) & (!n_n535) & (x23x) & (n_n4712) & (x30x)) + ((n_n325) & (n_n535) & (!x23x) & (!n_n4712) & (x30x)) + ((n_n325) & (n_n535) & (!x23x) & (n_n4712) & (!x30x)) + ((n_n325) & (n_n535) & (!x23x) & (n_n4712) & (x30x)) + ((n_n325) & (n_n535) & (x23x) & (!n_n4712) & (!x30x)) + ((n_n325) & (n_n535) & (x23x) & (!n_n4712) & (x30x)) + ((n_n325) & (n_n535) & (x23x) & (n_n4712) & (!x30x)) + ((n_n325) & (n_n535) & (x23x) & (n_n4712) & (x30x)));
	assign x12785x = (((!n_n4705) & (!n_n4708) & (!n_n4706) & (!n_n4707) & (n_n4713)) + ((!n_n4705) & (!n_n4708) & (!n_n4706) & (n_n4707) & (!n_n4713)) + ((!n_n4705) & (!n_n4708) & (!n_n4706) & (n_n4707) & (n_n4713)) + ((!n_n4705) & (!n_n4708) & (n_n4706) & (!n_n4707) & (!n_n4713)) + ((!n_n4705) & (!n_n4708) & (n_n4706) & (!n_n4707) & (n_n4713)) + ((!n_n4705) & (!n_n4708) & (n_n4706) & (n_n4707) & (!n_n4713)) + ((!n_n4705) & (!n_n4708) & (n_n4706) & (n_n4707) & (n_n4713)) + ((!n_n4705) & (n_n4708) & (!n_n4706) & (!n_n4707) & (!n_n4713)) + ((!n_n4705) & (n_n4708) & (!n_n4706) & (!n_n4707) & (n_n4713)) + ((!n_n4705) & (n_n4708) & (!n_n4706) & (n_n4707) & (!n_n4713)) + ((!n_n4705) & (n_n4708) & (!n_n4706) & (n_n4707) & (n_n4713)) + ((!n_n4705) & (n_n4708) & (n_n4706) & (!n_n4707) & (!n_n4713)) + ((!n_n4705) & (n_n4708) & (n_n4706) & (!n_n4707) & (n_n4713)) + ((!n_n4705) & (n_n4708) & (n_n4706) & (n_n4707) & (!n_n4713)) + ((!n_n4705) & (n_n4708) & (n_n4706) & (n_n4707) & (n_n4713)) + ((n_n4705) & (!n_n4708) & (!n_n4706) & (!n_n4707) & (!n_n4713)) + ((n_n4705) & (!n_n4708) & (!n_n4706) & (!n_n4707) & (n_n4713)) + ((n_n4705) & (!n_n4708) & (!n_n4706) & (n_n4707) & (!n_n4713)) + ((n_n4705) & (!n_n4708) & (!n_n4706) & (n_n4707) & (n_n4713)) + ((n_n4705) & (!n_n4708) & (n_n4706) & (!n_n4707) & (!n_n4713)) + ((n_n4705) & (!n_n4708) & (n_n4706) & (!n_n4707) & (n_n4713)) + ((n_n4705) & (!n_n4708) & (n_n4706) & (n_n4707) & (!n_n4713)) + ((n_n4705) & (!n_n4708) & (n_n4706) & (n_n4707) & (n_n4713)) + ((n_n4705) & (n_n4708) & (!n_n4706) & (!n_n4707) & (!n_n4713)) + ((n_n4705) & (n_n4708) & (!n_n4706) & (!n_n4707) & (n_n4713)) + ((n_n4705) & (n_n4708) & (!n_n4706) & (n_n4707) & (!n_n4713)) + ((n_n4705) & (n_n4708) & (!n_n4706) & (n_n4707) & (n_n4713)) + ((n_n4705) & (n_n4708) & (n_n4706) & (!n_n4707) & (!n_n4713)) + ((n_n4705) & (n_n4708) & (n_n4706) & (!n_n4707) & (n_n4713)) + ((n_n4705) & (n_n4708) & (n_n4706) & (n_n4707) & (!n_n4713)) + ((n_n4705) & (n_n4708) & (n_n4706) & (n_n4707) & (n_n4713)));
	assign n_n691 = (((!n_n4921) & (!n_n4929) & (!x249x) & (!n_n4932) & (x42x)) + ((!n_n4921) & (!n_n4929) & (!x249x) & (n_n4932) & (!x42x)) + ((!n_n4921) & (!n_n4929) & (!x249x) & (n_n4932) & (x42x)) + ((!n_n4921) & (!n_n4929) & (x249x) & (!n_n4932) & (!x42x)) + ((!n_n4921) & (!n_n4929) & (x249x) & (!n_n4932) & (x42x)) + ((!n_n4921) & (!n_n4929) & (x249x) & (n_n4932) & (!x42x)) + ((!n_n4921) & (!n_n4929) & (x249x) & (n_n4932) & (x42x)) + ((!n_n4921) & (n_n4929) & (!x249x) & (!n_n4932) & (!x42x)) + ((!n_n4921) & (n_n4929) & (!x249x) & (!n_n4932) & (x42x)) + ((!n_n4921) & (n_n4929) & (!x249x) & (n_n4932) & (!x42x)) + ((!n_n4921) & (n_n4929) & (!x249x) & (n_n4932) & (x42x)) + ((!n_n4921) & (n_n4929) & (x249x) & (!n_n4932) & (!x42x)) + ((!n_n4921) & (n_n4929) & (x249x) & (!n_n4932) & (x42x)) + ((!n_n4921) & (n_n4929) & (x249x) & (n_n4932) & (!x42x)) + ((!n_n4921) & (n_n4929) & (x249x) & (n_n4932) & (x42x)) + ((n_n4921) & (!n_n4929) & (!x249x) & (!n_n4932) & (!x42x)) + ((n_n4921) & (!n_n4929) & (!x249x) & (!n_n4932) & (x42x)) + ((n_n4921) & (!n_n4929) & (!x249x) & (n_n4932) & (!x42x)) + ((n_n4921) & (!n_n4929) & (!x249x) & (n_n4932) & (x42x)) + ((n_n4921) & (!n_n4929) & (x249x) & (!n_n4932) & (!x42x)) + ((n_n4921) & (!n_n4929) & (x249x) & (!n_n4932) & (x42x)) + ((n_n4921) & (!n_n4929) & (x249x) & (n_n4932) & (!x42x)) + ((n_n4921) & (!n_n4929) & (x249x) & (n_n4932) & (x42x)) + ((n_n4921) & (n_n4929) & (!x249x) & (!n_n4932) & (!x42x)) + ((n_n4921) & (n_n4929) & (!x249x) & (!n_n4932) & (x42x)) + ((n_n4921) & (n_n4929) & (!x249x) & (n_n4932) & (!x42x)) + ((n_n4921) & (n_n4929) & (!x249x) & (n_n4932) & (x42x)) + ((n_n4921) & (n_n4929) & (x249x) & (!n_n4932) & (!x42x)) + ((n_n4921) & (n_n4929) & (x249x) & (!n_n4932) & (x42x)) + ((n_n4921) & (n_n4929) & (x249x) & (n_n4932) & (!x42x)) + ((n_n4921) & (n_n4929) & (x249x) & (n_n4932) & (x42x)));
	assign x12724x = (((!n_n4898) & (!n_n4901) & (!n_n4904) & (n_n4899)) + ((!n_n4898) & (!n_n4901) & (n_n4904) & (!n_n4899)) + ((!n_n4898) & (!n_n4901) & (n_n4904) & (n_n4899)) + ((!n_n4898) & (n_n4901) & (!n_n4904) & (!n_n4899)) + ((!n_n4898) & (n_n4901) & (!n_n4904) & (n_n4899)) + ((!n_n4898) & (n_n4901) & (n_n4904) & (!n_n4899)) + ((!n_n4898) & (n_n4901) & (n_n4904) & (n_n4899)) + ((n_n4898) & (!n_n4901) & (!n_n4904) & (!n_n4899)) + ((n_n4898) & (!n_n4901) & (!n_n4904) & (n_n4899)) + ((n_n4898) & (!n_n4901) & (n_n4904) & (!n_n4899)) + ((n_n4898) & (!n_n4901) & (n_n4904) & (n_n4899)) + ((n_n4898) & (n_n4901) & (!n_n4904) & (!n_n4899)) + ((n_n4898) & (n_n4901) & (!n_n4904) & (n_n4899)) + ((n_n4898) & (n_n4901) & (n_n4904) & (!n_n4899)) + ((n_n4898) & (n_n4901) & (n_n4904) & (n_n4899)));
	assign x12725x = (((!n_n4897) & (!n_n4893) & (!x154x) & (n_n4896)) + ((!n_n4897) & (!n_n4893) & (x154x) & (!n_n4896)) + ((!n_n4897) & (!n_n4893) & (x154x) & (n_n4896)) + ((!n_n4897) & (n_n4893) & (!x154x) & (!n_n4896)) + ((!n_n4897) & (n_n4893) & (!x154x) & (n_n4896)) + ((!n_n4897) & (n_n4893) & (x154x) & (!n_n4896)) + ((!n_n4897) & (n_n4893) & (x154x) & (n_n4896)) + ((n_n4897) & (!n_n4893) & (!x154x) & (!n_n4896)) + ((n_n4897) & (!n_n4893) & (!x154x) & (n_n4896)) + ((n_n4897) & (!n_n4893) & (x154x) & (!n_n4896)) + ((n_n4897) & (!n_n4893) & (x154x) & (n_n4896)) + ((n_n4897) & (n_n4893) & (!x154x) & (!n_n4896)) + ((n_n4897) & (n_n4893) & (!x154x) & (n_n4896)) + ((n_n4897) & (n_n4893) & (x154x) & (!n_n4896)) + ((n_n4897) & (n_n4893) & (x154x) & (n_n4896)));
	assign x22191x = (((!x19x) & (!n_n5331) & (!x516x) & (!n_n5327) & (!n_n5328)) + ((!x19x) & (!n_n5331) & (x516x) & (!n_n5327) & (!n_n5328)) + ((x19x) & (!n_n5331) & (!x516x) & (!n_n5327) & (!n_n5328)));
	assign n_n632 = (((!n_n659) & (!n_n5325) & (!n_n5324) & (!n_n1900) & (!x22191x)) + ((!n_n659) & (!n_n5325) & (!n_n5324) & (n_n1900) & (!x22191x)) + ((!n_n659) & (!n_n5325) & (!n_n5324) & (n_n1900) & (x22191x)) + ((!n_n659) & (!n_n5325) & (n_n5324) & (!n_n1900) & (!x22191x)) + ((!n_n659) & (!n_n5325) & (n_n5324) & (!n_n1900) & (x22191x)) + ((!n_n659) & (!n_n5325) & (n_n5324) & (n_n1900) & (!x22191x)) + ((!n_n659) & (!n_n5325) & (n_n5324) & (n_n1900) & (x22191x)) + ((!n_n659) & (n_n5325) & (!n_n5324) & (!n_n1900) & (!x22191x)) + ((!n_n659) & (n_n5325) & (!n_n5324) & (!n_n1900) & (x22191x)) + ((!n_n659) & (n_n5325) & (!n_n5324) & (n_n1900) & (!x22191x)) + ((!n_n659) & (n_n5325) & (!n_n5324) & (n_n1900) & (x22191x)) + ((!n_n659) & (n_n5325) & (n_n5324) & (!n_n1900) & (!x22191x)) + ((!n_n659) & (n_n5325) & (n_n5324) & (!n_n1900) & (x22191x)) + ((!n_n659) & (n_n5325) & (n_n5324) & (n_n1900) & (!x22191x)) + ((!n_n659) & (n_n5325) & (n_n5324) & (n_n1900) & (x22191x)) + ((n_n659) & (!n_n5325) & (!n_n5324) & (!n_n1900) & (!x22191x)) + ((n_n659) & (!n_n5325) & (!n_n5324) & (!n_n1900) & (x22191x)) + ((n_n659) & (!n_n5325) & (!n_n5324) & (n_n1900) & (!x22191x)) + ((n_n659) & (!n_n5325) & (!n_n5324) & (n_n1900) & (x22191x)) + ((n_n659) & (!n_n5325) & (n_n5324) & (!n_n1900) & (!x22191x)) + ((n_n659) & (!n_n5325) & (n_n5324) & (!n_n1900) & (x22191x)) + ((n_n659) & (!n_n5325) & (n_n5324) & (n_n1900) & (!x22191x)) + ((n_n659) & (!n_n5325) & (n_n5324) & (n_n1900) & (x22191x)) + ((n_n659) & (n_n5325) & (!n_n5324) & (!n_n1900) & (!x22191x)) + ((n_n659) & (n_n5325) & (!n_n5324) & (!n_n1900) & (x22191x)) + ((n_n659) & (n_n5325) & (!n_n5324) & (n_n1900) & (!x22191x)) + ((n_n659) & (n_n5325) & (!n_n5324) & (n_n1900) & (x22191x)) + ((n_n659) & (n_n5325) & (n_n5324) & (!n_n1900) & (!x22191x)) + ((n_n659) & (n_n5325) & (n_n5324) & (!n_n1900) & (x22191x)) + ((n_n659) & (n_n5325) & (n_n5324) & (n_n1900) & (!x22191x)) + ((n_n659) & (n_n5325) & (n_n5324) & (n_n1900) & (x22191x)));
	assign x12767x = (((!n_n4789) & (!n_n2003) & (!x292x) & (!n_n4797) & (x380x)) + ((!n_n4789) & (!n_n2003) & (!x292x) & (n_n4797) & (!x380x)) + ((!n_n4789) & (!n_n2003) & (!x292x) & (n_n4797) & (x380x)) + ((!n_n4789) & (!n_n2003) & (x292x) & (!n_n4797) & (!x380x)) + ((!n_n4789) & (!n_n2003) & (x292x) & (!n_n4797) & (x380x)) + ((!n_n4789) & (!n_n2003) & (x292x) & (n_n4797) & (!x380x)) + ((!n_n4789) & (!n_n2003) & (x292x) & (n_n4797) & (x380x)) + ((!n_n4789) & (n_n2003) & (!x292x) & (!n_n4797) & (!x380x)) + ((!n_n4789) & (n_n2003) & (!x292x) & (!n_n4797) & (x380x)) + ((!n_n4789) & (n_n2003) & (!x292x) & (n_n4797) & (!x380x)) + ((!n_n4789) & (n_n2003) & (!x292x) & (n_n4797) & (x380x)) + ((!n_n4789) & (n_n2003) & (x292x) & (!n_n4797) & (!x380x)) + ((!n_n4789) & (n_n2003) & (x292x) & (!n_n4797) & (x380x)) + ((!n_n4789) & (n_n2003) & (x292x) & (n_n4797) & (!x380x)) + ((!n_n4789) & (n_n2003) & (x292x) & (n_n4797) & (x380x)) + ((n_n4789) & (!n_n2003) & (!x292x) & (!n_n4797) & (!x380x)) + ((n_n4789) & (!n_n2003) & (!x292x) & (!n_n4797) & (x380x)) + ((n_n4789) & (!n_n2003) & (!x292x) & (n_n4797) & (!x380x)) + ((n_n4789) & (!n_n2003) & (!x292x) & (n_n4797) & (x380x)) + ((n_n4789) & (!n_n2003) & (x292x) & (!n_n4797) & (!x380x)) + ((n_n4789) & (!n_n2003) & (x292x) & (!n_n4797) & (x380x)) + ((n_n4789) & (!n_n2003) & (x292x) & (n_n4797) & (!x380x)) + ((n_n4789) & (!n_n2003) & (x292x) & (n_n4797) & (x380x)) + ((n_n4789) & (n_n2003) & (!x292x) & (!n_n4797) & (!x380x)) + ((n_n4789) & (n_n2003) & (!x292x) & (!n_n4797) & (x380x)) + ((n_n4789) & (n_n2003) & (!x292x) & (n_n4797) & (!x380x)) + ((n_n4789) & (n_n2003) & (!x292x) & (n_n4797) & (x380x)) + ((n_n4789) & (n_n2003) & (x292x) & (!n_n4797) & (!x380x)) + ((n_n4789) & (n_n2003) & (x292x) & (!n_n4797) & (x380x)) + ((n_n4789) & (n_n2003) & (x292x) & (n_n4797) & (!x380x)) + ((n_n4789) & (n_n2003) & (x292x) & (n_n4797) & (x380x)));
	assign x12757x = (((!i_9_) & (!n_n532) & (!x530x) & (!n_n4807) & (x381x)) + ((!i_9_) & (!n_n532) & (!x530x) & (n_n4807) & (!x381x)) + ((!i_9_) & (!n_n532) & (!x530x) & (n_n4807) & (x381x)) + ((!i_9_) & (!n_n532) & (x530x) & (!n_n4807) & (x381x)) + ((!i_9_) & (!n_n532) & (x530x) & (n_n4807) & (!x381x)) + ((!i_9_) & (!n_n532) & (x530x) & (n_n4807) & (x381x)) + ((!i_9_) & (n_n532) & (!x530x) & (!n_n4807) & (x381x)) + ((!i_9_) & (n_n532) & (!x530x) & (n_n4807) & (!x381x)) + ((!i_9_) & (n_n532) & (!x530x) & (n_n4807) & (x381x)) + ((!i_9_) & (n_n532) & (x530x) & (!n_n4807) & (!x381x)) + ((!i_9_) & (n_n532) & (x530x) & (!n_n4807) & (x381x)) + ((!i_9_) & (n_n532) & (x530x) & (n_n4807) & (!x381x)) + ((!i_9_) & (n_n532) & (x530x) & (n_n4807) & (x381x)) + ((i_9_) & (!n_n532) & (!x530x) & (!n_n4807) & (x381x)) + ((i_9_) & (!n_n532) & (!x530x) & (n_n4807) & (!x381x)) + ((i_9_) & (!n_n532) & (!x530x) & (n_n4807) & (x381x)) + ((i_9_) & (!n_n532) & (x530x) & (!n_n4807) & (x381x)) + ((i_9_) & (!n_n532) & (x530x) & (n_n4807) & (!x381x)) + ((i_9_) & (!n_n532) & (x530x) & (n_n4807) & (x381x)) + ((i_9_) & (n_n532) & (!x530x) & (!n_n4807) & (x381x)) + ((i_9_) & (n_n532) & (!x530x) & (n_n4807) & (!x381x)) + ((i_9_) & (n_n532) & (!x530x) & (n_n4807) & (x381x)) + ((i_9_) & (n_n532) & (x530x) & (!n_n4807) & (x381x)) + ((i_9_) & (n_n532) & (x530x) & (n_n4807) & (!x381x)) + ((i_9_) & (n_n532) & (x530x) & (n_n4807) & (x381x)));
	assign x12758x = (((!x25x) & (!x530x) & (!x71x) & (!n_n4808) & (n_n4799)) + ((!x25x) & (!x530x) & (!x71x) & (n_n4808) & (!n_n4799)) + ((!x25x) & (!x530x) & (!x71x) & (n_n4808) & (n_n4799)) + ((!x25x) & (!x530x) & (x71x) & (!n_n4808) & (!n_n4799)) + ((!x25x) & (!x530x) & (x71x) & (!n_n4808) & (n_n4799)) + ((!x25x) & (!x530x) & (x71x) & (n_n4808) & (!n_n4799)) + ((!x25x) & (!x530x) & (x71x) & (n_n4808) & (n_n4799)) + ((!x25x) & (x530x) & (!x71x) & (!n_n4808) & (n_n4799)) + ((!x25x) & (x530x) & (!x71x) & (n_n4808) & (!n_n4799)) + ((!x25x) & (x530x) & (!x71x) & (n_n4808) & (n_n4799)) + ((!x25x) & (x530x) & (x71x) & (!n_n4808) & (!n_n4799)) + ((!x25x) & (x530x) & (x71x) & (!n_n4808) & (n_n4799)) + ((!x25x) & (x530x) & (x71x) & (n_n4808) & (!n_n4799)) + ((!x25x) & (x530x) & (x71x) & (n_n4808) & (n_n4799)) + ((x25x) & (!x530x) & (!x71x) & (!n_n4808) & (n_n4799)) + ((x25x) & (!x530x) & (!x71x) & (n_n4808) & (!n_n4799)) + ((x25x) & (!x530x) & (!x71x) & (n_n4808) & (n_n4799)) + ((x25x) & (!x530x) & (x71x) & (!n_n4808) & (!n_n4799)) + ((x25x) & (!x530x) & (x71x) & (!n_n4808) & (n_n4799)) + ((x25x) & (!x530x) & (x71x) & (n_n4808) & (!n_n4799)) + ((x25x) & (!x530x) & (x71x) & (n_n4808) & (n_n4799)) + ((x25x) & (x530x) & (!x71x) & (!n_n4808) & (!n_n4799)) + ((x25x) & (x530x) & (!x71x) & (!n_n4808) & (n_n4799)) + ((x25x) & (x530x) & (!x71x) & (n_n4808) & (!n_n4799)) + ((x25x) & (x530x) & (!x71x) & (n_n4808) & (n_n4799)) + ((x25x) & (x530x) & (x71x) & (!n_n4808) & (!n_n4799)) + ((x25x) & (x530x) & (x71x) & (!n_n4808) & (n_n4799)) + ((x25x) & (x530x) & (x71x) & (n_n4808) & (!n_n4799)) + ((x25x) & (x530x) & (x71x) & (n_n4808) & (n_n4799)));
	assign n_n702 = (((!n_n4782) & (!n_n4779) & (!n_n4781) & (!n_n4777) & (x12763x)) + ((!n_n4782) & (!n_n4779) & (!n_n4781) & (n_n4777) & (!x12763x)) + ((!n_n4782) & (!n_n4779) & (!n_n4781) & (n_n4777) & (x12763x)) + ((!n_n4782) & (!n_n4779) & (n_n4781) & (!n_n4777) & (!x12763x)) + ((!n_n4782) & (!n_n4779) & (n_n4781) & (!n_n4777) & (x12763x)) + ((!n_n4782) & (!n_n4779) & (n_n4781) & (n_n4777) & (!x12763x)) + ((!n_n4782) & (!n_n4779) & (n_n4781) & (n_n4777) & (x12763x)) + ((!n_n4782) & (n_n4779) & (!n_n4781) & (!n_n4777) & (!x12763x)) + ((!n_n4782) & (n_n4779) & (!n_n4781) & (!n_n4777) & (x12763x)) + ((!n_n4782) & (n_n4779) & (!n_n4781) & (n_n4777) & (!x12763x)) + ((!n_n4782) & (n_n4779) & (!n_n4781) & (n_n4777) & (x12763x)) + ((!n_n4782) & (n_n4779) & (n_n4781) & (!n_n4777) & (!x12763x)) + ((!n_n4782) & (n_n4779) & (n_n4781) & (!n_n4777) & (x12763x)) + ((!n_n4782) & (n_n4779) & (n_n4781) & (n_n4777) & (!x12763x)) + ((!n_n4782) & (n_n4779) & (n_n4781) & (n_n4777) & (x12763x)) + ((n_n4782) & (!n_n4779) & (!n_n4781) & (!n_n4777) & (!x12763x)) + ((n_n4782) & (!n_n4779) & (!n_n4781) & (!n_n4777) & (x12763x)) + ((n_n4782) & (!n_n4779) & (!n_n4781) & (n_n4777) & (!x12763x)) + ((n_n4782) & (!n_n4779) & (!n_n4781) & (n_n4777) & (x12763x)) + ((n_n4782) & (!n_n4779) & (n_n4781) & (!n_n4777) & (!x12763x)) + ((n_n4782) & (!n_n4779) & (n_n4781) & (!n_n4777) & (x12763x)) + ((n_n4782) & (!n_n4779) & (n_n4781) & (n_n4777) & (!x12763x)) + ((n_n4782) & (!n_n4779) & (n_n4781) & (n_n4777) & (x12763x)) + ((n_n4782) & (n_n4779) & (!n_n4781) & (!n_n4777) & (!x12763x)) + ((n_n4782) & (n_n4779) & (!n_n4781) & (!n_n4777) & (x12763x)) + ((n_n4782) & (n_n4779) & (!n_n4781) & (n_n4777) & (!x12763x)) + ((n_n4782) & (n_n4779) & (!n_n4781) & (n_n4777) & (x12763x)) + ((n_n4782) & (n_n4779) & (n_n4781) & (!n_n4777) & (!x12763x)) + ((n_n4782) & (n_n4779) & (n_n4781) & (!n_n4777) & (x12763x)) + ((n_n4782) & (n_n4779) & (n_n4781) & (n_n4777) & (!x12763x)) + ((n_n4782) & (n_n4779) & (n_n4781) & (n_n4777) & (x12763x)));
	assign n_n646 = (((!x12767x) & (!x12757x) & (!x12758x) & (n_n702)) + ((!x12767x) & (!x12757x) & (x12758x) & (!n_n702)) + ((!x12767x) & (!x12757x) & (x12758x) & (n_n702)) + ((!x12767x) & (x12757x) & (!x12758x) & (!n_n702)) + ((!x12767x) & (x12757x) & (!x12758x) & (n_n702)) + ((!x12767x) & (x12757x) & (x12758x) & (!n_n702)) + ((!x12767x) & (x12757x) & (x12758x) & (n_n702)) + ((x12767x) & (!x12757x) & (!x12758x) & (!n_n702)) + ((x12767x) & (!x12757x) & (!x12758x) & (n_n702)) + ((x12767x) & (!x12757x) & (x12758x) & (!n_n702)) + ((x12767x) & (!x12757x) & (x12758x) & (n_n702)) + ((x12767x) & (x12757x) & (!x12758x) & (!n_n702)) + ((x12767x) & (x12757x) & (!x12758x) & (n_n702)) + ((x12767x) & (x12757x) & (x12758x) & (!n_n702)) + ((x12767x) & (x12757x) & (x12758x) & (n_n702)));
	assign x12773x = (((!n_n4888) & (!n_n4882) & (!n_n4881) & (!n_n4889) & (x12772x)) + ((!n_n4888) & (!n_n4882) & (!n_n4881) & (n_n4889) & (!x12772x)) + ((!n_n4888) & (!n_n4882) & (!n_n4881) & (n_n4889) & (x12772x)) + ((!n_n4888) & (!n_n4882) & (n_n4881) & (!n_n4889) & (!x12772x)) + ((!n_n4888) & (!n_n4882) & (n_n4881) & (!n_n4889) & (x12772x)) + ((!n_n4888) & (!n_n4882) & (n_n4881) & (n_n4889) & (!x12772x)) + ((!n_n4888) & (!n_n4882) & (n_n4881) & (n_n4889) & (x12772x)) + ((!n_n4888) & (n_n4882) & (!n_n4881) & (!n_n4889) & (!x12772x)) + ((!n_n4888) & (n_n4882) & (!n_n4881) & (!n_n4889) & (x12772x)) + ((!n_n4888) & (n_n4882) & (!n_n4881) & (n_n4889) & (!x12772x)) + ((!n_n4888) & (n_n4882) & (!n_n4881) & (n_n4889) & (x12772x)) + ((!n_n4888) & (n_n4882) & (n_n4881) & (!n_n4889) & (!x12772x)) + ((!n_n4888) & (n_n4882) & (n_n4881) & (!n_n4889) & (x12772x)) + ((!n_n4888) & (n_n4882) & (n_n4881) & (n_n4889) & (!x12772x)) + ((!n_n4888) & (n_n4882) & (n_n4881) & (n_n4889) & (x12772x)) + ((n_n4888) & (!n_n4882) & (!n_n4881) & (!n_n4889) & (!x12772x)) + ((n_n4888) & (!n_n4882) & (!n_n4881) & (!n_n4889) & (x12772x)) + ((n_n4888) & (!n_n4882) & (!n_n4881) & (n_n4889) & (!x12772x)) + ((n_n4888) & (!n_n4882) & (!n_n4881) & (n_n4889) & (x12772x)) + ((n_n4888) & (!n_n4882) & (n_n4881) & (!n_n4889) & (!x12772x)) + ((n_n4888) & (!n_n4882) & (n_n4881) & (!n_n4889) & (x12772x)) + ((n_n4888) & (!n_n4882) & (n_n4881) & (n_n4889) & (!x12772x)) + ((n_n4888) & (!n_n4882) & (n_n4881) & (n_n4889) & (x12772x)) + ((n_n4888) & (n_n4882) & (!n_n4881) & (!n_n4889) & (!x12772x)) + ((n_n4888) & (n_n4882) & (!n_n4881) & (!n_n4889) & (x12772x)) + ((n_n4888) & (n_n4882) & (!n_n4881) & (n_n4889) & (!x12772x)) + ((n_n4888) & (n_n4882) & (!n_n4881) & (n_n4889) & (x12772x)) + ((n_n4888) & (n_n4882) & (n_n4881) & (!n_n4889) & (!x12772x)) + ((n_n4888) & (n_n4882) & (n_n4881) & (!n_n4889) & (x12772x)) + ((n_n4888) & (n_n4882) & (n_n4881) & (n_n4889) & (!x12772x)) + ((n_n4888) & (n_n4882) & (n_n4881) & (n_n4889) & (x12772x)));
	assign x12775x = (((!x12729x) & (!x12730x) & (!n_n696) & (x12773x)) + ((!x12729x) & (!x12730x) & (n_n696) & (!x12773x)) + ((!x12729x) & (!x12730x) & (n_n696) & (x12773x)) + ((!x12729x) & (x12730x) & (!n_n696) & (!x12773x)) + ((!x12729x) & (x12730x) & (!n_n696) & (x12773x)) + ((!x12729x) & (x12730x) & (n_n696) & (!x12773x)) + ((!x12729x) & (x12730x) & (n_n696) & (x12773x)) + ((x12729x) & (!x12730x) & (!n_n696) & (!x12773x)) + ((x12729x) & (!x12730x) & (!n_n696) & (x12773x)) + ((x12729x) & (!x12730x) & (n_n696) & (!x12773x)) + ((x12729x) & (!x12730x) & (n_n696) & (x12773x)) + ((x12729x) & (x12730x) & (!n_n696) & (!x12773x)) + ((x12729x) & (x12730x) & (!n_n696) & (x12773x)) + ((x12729x) & (x12730x) & (n_n696) & (!x12773x)) + ((x12729x) & (x12730x) & (n_n696) & (x12773x)));
	assign x12751x = (((!n_n4843) & (!n_n4845) & (!x52x) & (!x150x) & (x326x)) + ((!n_n4843) & (!n_n4845) & (!x52x) & (x150x) & (!x326x)) + ((!n_n4843) & (!n_n4845) & (!x52x) & (x150x) & (x326x)) + ((!n_n4843) & (!n_n4845) & (x52x) & (!x150x) & (!x326x)) + ((!n_n4843) & (!n_n4845) & (x52x) & (!x150x) & (x326x)) + ((!n_n4843) & (!n_n4845) & (x52x) & (x150x) & (!x326x)) + ((!n_n4843) & (!n_n4845) & (x52x) & (x150x) & (x326x)) + ((!n_n4843) & (n_n4845) & (!x52x) & (!x150x) & (!x326x)) + ((!n_n4843) & (n_n4845) & (!x52x) & (!x150x) & (x326x)) + ((!n_n4843) & (n_n4845) & (!x52x) & (x150x) & (!x326x)) + ((!n_n4843) & (n_n4845) & (!x52x) & (x150x) & (x326x)) + ((!n_n4843) & (n_n4845) & (x52x) & (!x150x) & (!x326x)) + ((!n_n4843) & (n_n4845) & (x52x) & (!x150x) & (x326x)) + ((!n_n4843) & (n_n4845) & (x52x) & (x150x) & (!x326x)) + ((!n_n4843) & (n_n4845) & (x52x) & (x150x) & (x326x)) + ((n_n4843) & (!n_n4845) & (!x52x) & (!x150x) & (!x326x)) + ((n_n4843) & (!n_n4845) & (!x52x) & (!x150x) & (x326x)) + ((n_n4843) & (!n_n4845) & (!x52x) & (x150x) & (!x326x)) + ((n_n4843) & (!n_n4845) & (!x52x) & (x150x) & (x326x)) + ((n_n4843) & (!n_n4845) & (x52x) & (!x150x) & (!x326x)) + ((n_n4843) & (!n_n4845) & (x52x) & (!x150x) & (x326x)) + ((n_n4843) & (!n_n4845) & (x52x) & (x150x) & (!x326x)) + ((n_n4843) & (!n_n4845) & (x52x) & (x150x) & (x326x)) + ((n_n4843) & (n_n4845) & (!x52x) & (!x150x) & (!x326x)) + ((n_n4843) & (n_n4845) & (!x52x) & (!x150x) & (x326x)) + ((n_n4843) & (n_n4845) & (!x52x) & (x150x) & (!x326x)) + ((n_n4843) & (n_n4845) & (!x52x) & (x150x) & (x326x)) + ((n_n4843) & (n_n4845) & (x52x) & (!x150x) & (!x326x)) + ((n_n4843) & (n_n4845) & (x52x) & (!x150x) & (x326x)) + ((n_n4843) & (n_n4845) & (x52x) & (x150x) & (!x326x)) + ((n_n4843) & (n_n4845) & (x52x) & (x150x) & (x326x)));
	assign n_n856 = (((!i_9_) & (!n_n532) & (!n_n534) & (!x483x) & (n_n4734)) + ((!i_9_) & (!n_n532) & (!n_n534) & (x483x) & (n_n4734)) + ((!i_9_) & (!n_n532) & (n_n534) & (!x483x) & (n_n4734)) + ((!i_9_) & (!n_n532) & (n_n534) & (x483x) & (!n_n4734)) + ((!i_9_) & (!n_n532) & (n_n534) & (x483x) & (n_n4734)) + ((!i_9_) & (n_n532) & (!n_n534) & (!x483x) & (n_n4734)) + ((!i_9_) & (n_n532) & (!n_n534) & (x483x) & (!n_n4734)) + ((!i_9_) & (n_n532) & (!n_n534) & (x483x) & (n_n4734)) + ((!i_9_) & (n_n532) & (n_n534) & (!x483x) & (n_n4734)) + ((!i_9_) & (n_n532) & (n_n534) & (x483x) & (!n_n4734)) + ((!i_9_) & (n_n532) & (n_n534) & (x483x) & (n_n4734)) + ((i_9_) & (!n_n532) & (!n_n534) & (!x483x) & (n_n4734)) + ((i_9_) & (!n_n532) & (!n_n534) & (x483x) & (n_n4734)) + ((i_9_) & (!n_n532) & (n_n534) & (!x483x) & (n_n4734)) + ((i_9_) & (!n_n532) & (n_n534) & (x483x) & (n_n4734)) + ((i_9_) & (n_n532) & (!n_n534) & (!x483x) & (n_n4734)) + ((i_9_) & (n_n532) & (!n_n534) & (x483x) & (n_n4734)) + ((i_9_) & (n_n532) & (n_n534) & (!x483x) & (n_n4734)) + ((i_9_) & (n_n532) & (n_n534) & (x483x) & (n_n4734)));
	assign n_n706 = (((!n_n4720) & (!n_n4717) & (!n_n4728) & (!n_n4719) & (x12791x)) + ((!n_n4720) & (!n_n4717) & (!n_n4728) & (n_n4719) & (!x12791x)) + ((!n_n4720) & (!n_n4717) & (!n_n4728) & (n_n4719) & (x12791x)) + ((!n_n4720) & (!n_n4717) & (n_n4728) & (!n_n4719) & (!x12791x)) + ((!n_n4720) & (!n_n4717) & (n_n4728) & (!n_n4719) & (x12791x)) + ((!n_n4720) & (!n_n4717) & (n_n4728) & (n_n4719) & (!x12791x)) + ((!n_n4720) & (!n_n4717) & (n_n4728) & (n_n4719) & (x12791x)) + ((!n_n4720) & (n_n4717) & (!n_n4728) & (!n_n4719) & (!x12791x)) + ((!n_n4720) & (n_n4717) & (!n_n4728) & (!n_n4719) & (x12791x)) + ((!n_n4720) & (n_n4717) & (!n_n4728) & (n_n4719) & (!x12791x)) + ((!n_n4720) & (n_n4717) & (!n_n4728) & (n_n4719) & (x12791x)) + ((!n_n4720) & (n_n4717) & (n_n4728) & (!n_n4719) & (!x12791x)) + ((!n_n4720) & (n_n4717) & (n_n4728) & (!n_n4719) & (x12791x)) + ((!n_n4720) & (n_n4717) & (n_n4728) & (n_n4719) & (!x12791x)) + ((!n_n4720) & (n_n4717) & (n_n4728) & (n_n4719) & (x12791x)) + ((n_n4720) & (!n_n4717) & (!n_n4728) & (!n_n4719) & (!x12791x)) + ((n_n4720) & (!n_n4717) & (!n_n4728) & (!n_n4719) & (x12791x)) + ((n_n4720) & (!n_n4717) & (!n_n4728) & (n_n4719) & (!x12791x)) + ((n_n4720) & (!n_n4717) & (!n_n4728) & (n_n4719) & (x12791x)) + ((n_n4720) & (!n_n4717) & (n_n4728) & (!n_n4719) & (!x12791x)) + ((n_n4720) & (!n_n4717) & (n_n4728) & (!n_n4719) & (x12791x)) + ((n_n4720) & (!n_n4717) & (n_n4728) & (n_n4719) & (!x12791x)) + ((n_n4720) & (!n_n4717) & (n_n4728) & (n_n4719) & (x12791x)) + ((n_n4720) & (n_n4717) & (!n_n4728) & (!n_n4719) & (!x12791x)) + ((n_n4720) & (n_n4717) & (!n_n4728) & (!n_n4719) & (x12791x)) + ((n_n4720) & (n_n4717) & (!n_n4728) & (n_n4719) & (!x12791x)) + ((n_n4720) & (n_n4717) & (!n_n4728) & (n_n4719) & (x12791x)) + ((n_n4720) & (n_n4717) & (n_n4728) & (!n_n4719) & (!x12791x)) + ((n_n4720) & (n_n4717) & (n_n4728) & (!n_n4719) & (x12791x)) + ((n_n4720) & (n_n4717) & (n_n4728) & (n_n4719) & (!x12791x)) + ((n_n4720) & (n_n4717) & (n_n4728) & (n_n4719) & (x12791x)));
	assign x12794x = (((!n_n4697) & (!n_n4696) & (!n_n4695) & (n_n4699)) + ((!n_n4697) & (!n_n4696) & (n_n4695) & (!n_n4699)) + ((!n_n4697) & (!n_n4696) & (n_n4695) & (n_n4699)) + ((!n_n4697) & (n_n4696) & (!n_n4695) & (!n_n4699)) + ((!n_n4697) & (n_n4696) & (!n_n4695) & (n_n4699)) + ((!n_n4697) & (n_n4696) & (n_n4695) & (!n_n4699)) + ((!n_n4697) & (n_n4696) & (n_n4695) & (n_n4699)) + ((n_n4697) & (!n_n4696) & (!n_n4695) & (!n_n4699)) + ((n_n4697) & (!n_n4696) & (!n_n4695) & (n_n4699)) + ((n_n4697) & (!n_n4696) & (n_n4695) & (!n_n4699)) + ((n_n4697) & (!n_n4696) & (n_n4695) & (n_n4699)) + ((n_n4697) & (n_n4696) & (!n_n4695) & (!n_n4699)) + ((n_n4697) & (n_n4696) & (!n_n4695) & (n_n4699)) + ((n_n4697) & (n_n4696) & (n_n4695) & (!n_n4699)) + ((n_n4697) & (n_n4696) & (n_n4695) & (n_n4699)));
	assign x12795x = (((!n_n528) & (!x14x) & (!n_n535) & (!n_n3849) & (n_n4694)) + ((!n_n528) & (!x14x) & (!n_n535) & (n_n3849) & (!n_n4694)) + ((!n_n528) & (!x14x) & (!n_n535) & (n_n3849) & (n_n4694)) + ((!n_n528) & (!x14x) & (n_n535) & (!n_n3849) & (n_n4694)) + ((!n_n528) & (!x14x) & (n_n535) & (n_n3849) & (!n_n4694)) + ((!n_n528) & (!x14x) & (n_n535) & (n_n3849) & (n_n4694)) + ((!n_n528) & (x14x) & (!n_n535) & (!n_n3849) & (n_n4694)) + ((!n_n528) & (x14x) & (!n_n535) & (n_n3849) & (!n_n4694)) + ((!n_n528) & (x14x) & (!n_n535) & (n_n3849) & (n_n4694)) + ((!n_n528) & (x14x) & (n_n535) & (!n_n3849) & (n_n4694)) + ((!n_n528) & (x14x) & (n_n535) & (n_n3849) & (!n_n4694)) + ((!n_n528) & (x14x) & (n_n535) & (n_n3849) & (n_n4694)) + ((n_n528) & (!x14x) & (!n_n535) & (!n_n3849) & (n_n4694)) + ((n_n528) & (!x14x) & (!n_n535) & (n_n3849) & (!n_n4694)) + ((n_n528) & (!x14x) & (!n_n535) & (n_n3849) & (n_n4694)) + ((n_n528) & (!x14x) & (n_n535) & (!n_n3849) & (n_n4694)) + ((n_n528) & (!x14x) & (n_n535) & (n_n3849) & (!n_n4694)) + ((n_n528) & (!x14x) & (n_n535) & (n_n3849) & (n_n4694)) + ((n_n528) & (x14x) & (!n_n535) & (!n_n3849) & (n_n4694)) + ((n_n528) & (x14x) & (!n_n535) & (n_n3849) & (!n_n4694)) + ((n_n528) & (x14x) & (!n_n535) & (n_n3849) & (n_n4694)) + ((n_n528) & (x14x) & (n_n535) & (!n_n3849) & (!n_n4694)) + ((n_n528) & (x14x) & (n_n535) & (!n_n3849) & (n_n4694)) + ((n_n528) & (x14x) & (n_n535) & (n_n3849) & (!n_n4694)) + ((n_n528) & (x14x) & (n_n535) & (n_n3849) & (n_n4694)));
	assign n_n648 = (((!x12784x) & (!x12785x) & (!n_n706) & (!x12794x) & (x12795x)) + ((!x12784x) & (!x12785x) & (!n_n706) & (x12794x) & (!x12795x)) + ((!x12784x) & (!x12785x) & (!n_n706) & (x12794x) & (x12795x)) + ((!x12784x) & (!x12785x) & (n_n706) & (!x12794x) & (!x12795x)) + ((!x12784x) & (!x12785x) & (n_n706) & (!x12794x) & (x12795x)) + ((!x12784x) & (!x12785x) & (n_n706) & (x12794x) & (!x12795x)) + ((!x12784x) & (!x12785x) & (n_n706) & (x12794x) & (x12795x)) + ((!x12784x) & (x12785x) & (!n_n706) & (!x12794x) & (!x12795x)) + ((!x12784x) & (x12785x) & (!n_n706) & (!x12794x) & (x12795x)) + ((!x12784x) & (x12785x) & (!n_n706) & (x12794x) & (!x12795x)) + ((!x12784x) & (x12785x) & (!n_n706) & (x12794x) & (x12795x)) + ((!x12784x) & (x12785x) & (n_n706) & (!x12794x) & (!x12795x)) + ((!x12784x) & (x12785x) & (n_n706) & (!x12794x) & (x12795x)) + ((!x12784x) & (x12785x) & (n_n706) & (x12794x) & (!x12795x)) + ((!x12784x) & (x12785x) & (n_n706) & (x12794x) & (x12795x)) + ((x12784x) & (!x12785x) & (!n_n706) & (!x12794x) & (!x12795x)) + ((x12784x) & (!x12785x) & (!n_n706) & (!x12794x) & (x12795x)) + ((x12784x) & (!x12785x) & (!n_n706) & (x12794x) & (!x12795x)) + ((x12784x) & (!x12785x) & (!n_n706) & (x12794x) & (x12795x)) + ((x12784x) & (!x12785x) & (n_n706) & (!x12794x) & (!x12795x)) + ((x12784x) & (!x12785x) & (n_n706) & (!x12794x) & (x12795x)) + ((x12784x) & (!x12785x) & (n_n706) & (x12794x) & (!x12795x)) + ((x12784x) & (!x12785x) & (n_n706) & (x12794x) & (x12795x)) + ((x12784x) & (x12785x) & (!n_n706) & (!x12794x) & (!x12795x)) + ((x12784x) & (x12785x) & (!n_n706) & (!x12794x) & (x12795x)) + ((x12784x) & (x12785x) & (!n_n706) & (x12794x) & (!x12795x)) + ((x12784x) & (x12785x) & (!n_n706) & (x12794x) & (x12795x)) + ((x12784x) & (x12785x) & (n_n706) & (!x12794x) & (!x12795x)) + ((x12784x) & (x12785x) & (n_n706) & (!x12794x) & (x12795x)) + ((x12784x) & (x12785x) & (n_n706) & (x12794x) & (!x12795x)) + ((x12784x) & (x12785x) & (n_n706) & (x12794x) & (x12795x)));
	assign n_n709 = (((!n_n4677) & (!x426x) & (!n_n4685) & (!n_n1636) & (x417x)) + ((!n_n4677) & (!x426x) & (!n_n4685) & (n_n1636) & (!x417x)) + ((!n_n4677) & (!x426x) & (!n_n4685) & (n_n1636) & (x417x)) + ((!n_n4677) & (!x426x) & (n_n4685) & (!n_n1636) & (!x417x)) + ((!n_n4677) & (!x426x) & (n_n4685) & (!n_n1636) & (x417x)) + ((!n_n4677) & (!x426x) & (n_n4685) & (n_n1636) & (!x417x)) + ((!n_n4677) & (!x426x) & (n_n4685) & (n_n1636) & (x417x)) + ((!n_n4677) & (x426x) & (!n_n4685) & (!n_n1636) & (!x417x)) + ((!n_n4677) & (x426x) & (!n_n4685) & (!n_n1636) & (x417x)) + ((!n_n4677) & (x426x) & (!n_n4685) & (n_n1636) & (!x417x)) + ((!n_n4677) & (x426x) & (!n_n4685) & (n_n1636) & (x417x)) + ((!n_n4677) & (x426x) & (n_n4685) & (!n_n1636) & (!x417x)) + ((!n_n4677) & (x426x) & (n_n4685) & (!n_n1636) & (x417x)) + ((!n_n4677) & (x426x) & (n_n4685) & (n_n1636) & (!x417x)) + ((!n_n4677) & (x426x) & (n_n4685) & (n_n1636) & (x417x)) + ((n_n4677) & (!x426x) & (!n_n4685) & (!n_n1636) & (!x417x)) + ((n_n4677) & (!x426x) & (!n_n4685) & (!n_n1636) & (x417x)) + ((n_n4677) & (!x426x) & (!n_n4685) & (n_n1636) & (!x417x)) + ((n_n4677) & (!x426x) & (!n_n4685) & (n_n1636) & (x417x)) + ((n_n4677) & (!x426x) & (n_n4685) & (!n_n1636) & (!x417x)) + ((n_n4677) & (!x426x) & (n_n4685) & (!n_n1636) & (x417x)) + ((n_n4677) & (!x426x) & (n_n4685) & (n_n1636) & (!x417x)) + ((n_n4677) & (!x426x) & (n_n4685) & (n_n1636) & (x417x)) + ((n_n4677) & (x426x) & (!n_n4685) & (!n_n1636) & (!x417x)) + ((n_n4677) & (x426x) & (!n_n4685) & (!n_n1636) & (x417x)) + ((n_n4677) & (x426x) & (!n_n4685) & (n_n1636) & (!x417x)) + ((n_n4677) & (x426x) & (!n_n4685) & (n_n1636) & (x417x)) + ((n_n4677) & (x426x) & (n_n4685) & (!n_n1636) & (!x417x)) + ((n_n4677) & (x426x) & (n_n4685) & (!n_n1636) & (x417x)) + ((n_n4677) & (x426x) & (n_n4685) & (n_n1636) & (!x417x)) + ((n_n4677) & (x426x) & (n_n4685) & (n_n1636) & (x417x)));
	assign n_n710 = (((!n_n4669) & (!n_n4675) & (!n_n4671) & (!x339x) & (x12804x)) + ((!n_n4669) & (!n_n4675) & (!n_n4671) & (x339x) & (!x12804x)) + ((!n_n4669) & (!n_n4675) & (!n_n4671) & (x339x) & (x12804x)) + ((!n_n4669) & (!n_n4675) & (n_n4671) & (!x339x) & (!x12804x)) + ((!n_n4669) & (!n_n4675) & (n_n4671) & (!x339x) & (x12804x)) + ((!n_n4669) & (!n_n4675) & (n_n4671) & (x339x) & (!x12804x)) + ((!n_n4669) & (!n_n4675) & (n_n4671) & (x339x) & (x12804x)) + ((!n_n4669) & (n_n4675) & (!n_n4671) & (!x339x) & (!x12804x)) + ((!n_n4669) & (n_n4675) & (!n_n4671) & (!x339x) & (x12804x)) + ((!n_n4669) & (n_n4675) & (!n_n4671) & (x339x) & (!x12804x)) + ((!n_n4669) & (n_n4675) & (!n_n4671) & (x339x) & (x12804x)) + ((!n_n4669) & (n_n4675) & (n_n4671) & (!x339x) & (!x12804x)) + ((!n_n4669) & (n_n4675) & (n_n4671) & (!x339x) & (x12804x)) + ((!n_n4669) & (n_n4675) & (n_n4671) & (x339x) & (!x12804x)) + ((!n_n4669) & (n_n4675) & (n_n4671) & (x339x) & (x12804x)) + ((n_n4669) & (!n_n4675) & (!n_n4671) & (!x339x) & (!x12804x)) + ((n_n4669) & (!n_n4675) & (!n_n4671) & (!x339x) & (x12804x)) + ((n_n4669) & (!n_n4675) & (!n_n4671) & (x339x) & (!x12804x)) + ((n_n4669) & (!n_n4675) & (!n_n4671) & (x339x) & (x12804x)) + ((n_n4669) & (!n_n4675) & (n_n4671) & (!x339x) & (!x12804x)) + ((n_n4669) & (!n_n4675) & (n_n4671) & (!x339x) & (x12804x)) + ((n_n4669) & (!n_n4675) & (n_n4671) & (x339x) & (!x12804x)) + ((n_n4669) & (!n_n4675) & (n_n4671) & (x339x) & (x12804x)) + ((n_n4669) & (n_n4675) & (!n_n4671) & (!x339x) & (!x12804x)) + ((n_n4669) & (n_n4675) & (!n_n4671) & (!x339x) & (x12804x)) + ((n_n4669) & (n_n4675) & (!n_n4671) & (x339x) & (!x12804x)) + ((n_n4669) & (n_n4675) & (!n_n4671) & (x339x) & (x12804x)) + ((n_n4669) & (n_n4675) & (n_n4671) & (!x339x) & (!x12804x)) + ((n_n4669) & (n_n4675) & (n_n4671) & (!x339x) & (x12804x)) + ((n_n4669) & (n_n4675) & (n_n4671) & (x339x) & (!x12804x)) + ((n_n4669) & (n_n4675) & (n_n4671) & (x339x) & (x12804x)));
	assign x12811x = (((!n_n4662) & (!n_n4659) & (!n_n4655) & (n_n4658)) + ((!n_n4662) & (!n_n4659) & (n_n4655) & (!n_n4658)) + ((!n_n4662) & (!n_n4659) & (n_n4655) & (n_n4658)) + ((!n_n4662) & (n_n4659) & (!n_n4655) & (!n_n4658)) + ((!n_n4662) & (n_n4659) & (!n_n4655) & (n_n4658)) + ((!n_n4662) & (n_n4659) & (n_n4655) & (!n_n4658)) + ((!n_n4662) & (n_n4659) & (n_n4655) & (n_n4658)) + ((n_n4662) & (!n_n4659) & (!n_n4655) & (!n_n4658)) + ((n_n4662) & (!n_n4659) & (!n_n4655) & (n_n4658)) + ((n_n4662) & (!n_n4659) & (n_n4655) & (!n_n4658)) + ((n_n4662) & (!n_n4659) & (n_n4655) & (n_n4658)) + ((n_n4662) & (n_n4659) & (!n_n4655) & (!n_n4658)) + ((n_n4662) & (n_n4659) & (!n_n4655) & (n_n4658)) + ((n_n4662) & (n_n4659) & (n_n4655) & (!n_n4658)) + ((n_n4662) & (n_n4659) & (n_n4655) & (n_n4658)));
	assign x12812x = (((!n_n4644) & (!n_n4649) & (!n_n4652) & (!n_n4663) & (n_n4657)) + ((!n_n4644) & (!n_n4649) & (!n_n4652) & (n_n4663) & (!n_n4657)) + ((!n_n4644) & (!n_n4649) & (!n_n4652) & (n_n4663) & (n_n4657)) + ((!n_n4644) & (!n_n4649) & (n_n4652) & (!n_n4663) & (!n_n4657)) + ((!n_n4644) & (!n_n4649) & (n_n4652) & (!n_n4663) & (n_n4657)) + ((!n_n4644) & (!n_n4649) & (n_n4652) & (n_n4663) & (!n_n4657)) + ((!n_n4644) & (!n_n4649) & (n_n4652) & (n_n4663) & (n_n4657)) + ((!n_n4644) & (n_n4649) & (!n_n4652) & (!n_n4663) & (!n_n4657)) + ((!n_n4644) & (n_n4649) & (!n_n4652) & (!n_n4663) & (n_n4657)) + ((!n_n4644) & (n_n4649) & (!n_n4652) & (n_n4663) & (!n_n4657)) + ((!n_n4644) & (n_n4649) & (!n_n4652) & (n_n4663) & (n_n4657)) + ((!n_n4644) & (n_n4649) & (n_n4652) & (!n_n4663) & (!n_n4657)) + ((!n_n4644) & (n_n4649) & (n_n4652) & (!n_n4663) & (n_n4657)) + ((!n_n4644) & (n_n4649) & (n_n4652) & (n_n4663) & (!n_n4657)) + ((!n_n4644) & (n_n4649) & (n_n4652) & (n_n4663) & (n_n4657)) + ((n_n4644) & (!n_n4649) & (!n_n4652) & (!n_n4663) & (!n_n4657)) + ((n_n4644) & (!n_n4649) & (!n_n4652) & (!n_n4663) & (n_n4657)) + ((n_n4644) & (!n_n4649) & (!n_n4652) & (n_n4663) & (!n_n4657)) + ((n_n4644) & (!n_n4649) & (!n_n4652) & (n_n4663) & (n_n4657)) + ((n_n4644) & (!n_n4649) & (n_n4652) & (!n_n4663) & (!n_n4657)) + ((n_n4644) & (!n_n4649) & (n_n4652) & (!n_n4663) & (n_n4657)) + ((n_n4644) & (!n_n4649) & (n_n4652) & (n_n4663) & (!n_n4657)) + ((n_n4644) & (!n_n4649) & (n_n4652) & (n_n4663) & (n_n4657)) + ((n_n4644) & (n_n4649) & (!n_n4652) & (!n_n4663) & (!n_n4657)) + ((n_n4644) & (n_n4649) & (!n_n4652) & (!n_n4663) & (n_n4657)) + ((n_n4644) & (n_n4649) & (!n_n4652) & (n_n4663) & (!n_n4657)) + ((n_n4644) & (n_n4649) & (!n_n4652) & (n_n4663) & (n_n4657)) + ((n_n4644) & (n_n4649) & (n_n4652) & (!n_n4663) & (!n_n4657)) + ((n_n4644) & (n_n4649) & (n_n4652) & (!n_n4663) & (n_n4657)) + ((n_n4644) & (n_n4649) & (n_n4652) & (n_n4663) & (!n_n4657)) + ((n_n4644) & (n_n4649) & (n_n4652) & (n_n4663) & (n_n4657)));
	assign n_n649 = (((!n_n709) & (!n_n710) & (!x12811x) & (x12812x)) + ((!n_n709) & (!n_n710) & (x12811x) & (!x12812x)) + ((!n_n709) & (!n_n710) & (x12811x) & (x12812x)) + ((!n_n709) & (n_n710) & (!x12811x) & (!x12812x)) + ((!n_n709) & (n_n710) & (!x12811x) & (x12812x)) + ((!n_n709) & (n_n710) & (x12811x) & (!x12812x)) + ((!n_n709) & (n_n710) & (x12811x) & (x12812x)) + ((n_n709) & (!n_n710) & (!x12811x) & (!x12812x)) + ((n_n709) & (!n_n710) & (!x12811x) & (x12812x)) + ((n_n709) & (!n_n710) & (x12811x) & (!x12812x)) + ((n_n709) & (!n_n710) & (x12811x) & (x12812x)) + ((n_n709) & (n_n710) & (!x12811x) & (!x12812x)) + ((n_n709) & (n_n710) & (!x12811x) & (x12812x)) + ((n_n709) & (n_n710) & (x12811x) & (!x12812x)) + ((n_n709) & (n_n710) & (x12811x) & (x12812x)));
	assign x22132x = (((!n_n4757) & (!n_n4747) & (!n_n4755) & (!n_n4758)));
	assign n_n704 = (((!n_n4751) & (!n_n4752) & (!x47x) & (!n_n4745) & (!x22132x)) + ((!n_n4751) & (!n_n4752) & (!x47x) & (n_n4745) & (!x22132x)) + ((!n_n4751) & (!n_n4752) & (!x47x) & (n_n4745) & (x22132x)) + ((!n_n4751) & (!n_n4752) & (x47x) & (!n_n4745) & (!x22132x)) + ((!n_n4751) & (!n_n4752) & (x47x) & (!n_n4745) & (x22132x)) + ((!n_n4751) & (!n_n4752) & (x47x) & (n_n4745) & (!x22132x)) + ((!n_n4751) & (!n_n4752) & (x47x) & (n_n4745) & (x22132x)) + ((!n_n4751) & (n_n4752) & (!x47x) & (!n_n4745) & (!x22132x)) + ((!n_n4751) & (n_n4752) & (!x47x) & (!n_n4745) & (x22132x)) + ((!n_n4751) & (n_n4752) & (!x47x) & (n_n4745) & (!x22132x)) + ((!n_n4751) & (n_n4752) & (!x47x) & (n_n4745) & (x22132x)) + ((!n_n4751) & (n_n4752) & (x47x) & (!n_n4745) & (!x22132x)) + ((!n_n4751) & (n_n4752) & (x47x) & (!n_n4745) & (x22132x)) + ((!n_n4751) & (n_n4752) & (x47x) & (n_n4745) & (!x22132x)) + ((!n_n4751) & (n_n4752) & (x47x) & (n_n4745) & (x22132x)) + ((n_n4751) & (!n_n4752) & (!x47x) & (!n_n4745) & (!x22132x)) + ((n_n4751) & (!n_n4752) & (!x47x) & (!n_n4745) & (x22132x)) + ((n_n4751) & (!n_n4752) & (!x47x) & (n_n4745) & (!x22132x)) + ((n_n4751) & (!n_n4752) & (!x47x) & (n_n4745) & (x22132x)) + ((n_n4751) & (!n_n4752) & (x47x) & (!n_n4745) & (!x22132x)) + ((n_n4751) & (!n_n4752) & (x47x) & (!n_n4745) & (x22132x)) + ((n_n4751) & (!n_n4752) & (x47x) & (n_n4745) & (!x22132x)) + ((n_n4751) & (!n_n4752) & (x47x) & (n_n4745) & (x22132x)) + ((n_n4751) & (n_n4752) & (!x47x) & (!n_n4745) & (!x22132x)) + ((n_n4751) & (n_n4752) & (!x47x) & (!n_n4745) & (x22132x)) + ((n_n4751) & (n_n4752) & (!x47x) & (n_n4745) & (!x22132x)) + ((n_n4751) & (n_n4752) & (!x47x) & (n_n4745) & (x22132x)) + ((n_n4751) & (n_n4752) & (x47x) & (!n_n4745) & (!x22132x)) + ((n_n4751) & (n_n4752) & (x47x) & (!n_n4745) & (x22132x)) + ((n_n4751) & (n_n4752) & (x47x) & (n_n4745) & (!x22132x)) + ((n_n4751) & (n_n4752) & (x47x) & (n_n4745) & (x22132x)));
	assign x12824x = (((!n_n4760) & (!n_n4762) & (!n_n4769) & (n_n856)) + ((!n_n4760) & (!n_n4762) & (n_n4769) & (!n_n856)) + ((!n_n4760) & (!n_n4762) & (n_n4769) & (n_n856)) + ((!n_n4760) & (n_n4762) & (!n_n4769) & (!n_n856)) + ((!n_n4760) & (n_n4762) & (!n_n4769) & (n_n856)) + ((!n_n4760) & (n_n4762) & (n_n4769) & (!n_n856)) + ((!n_n4760) & (n_n4762) & (n_n4769) & (n_n856)) + ((n_n4760) & (!n_n4762) & (!n_n4769) & (!n_n856)) + ((n_n4760) & (!n_n4762) & (!n_n4769) & (n_n856)) + ((n_n4760) & (!n_n4762) & (n_n4769) & (!n_n856)) + ((n_n4760) & (!n_n4762) & (n_n4769) & (n_n856)) + ((n_n4760) & (n_n4762) & (!n_n4769) & (!n_n856)) + ((n_n4760) & (n_n4762) & (!n_n4769) & (n_n856)) + ((n_n4760) & (n_n4762) & (n_n4769) & (!n_n856)) + ((n_n4760) & (n_n4762) & (n_n4769) & (n_n856)));
	assign x12827x = (((!n_n4205) & (!n_n4204) & (!x456x) & (!n_n704) & (x12824x)) + ((!n_n4205) & (!n_n4204) & (!x456x) & (n_n704) & (!x12824x)) + ((!n_n4205) & (!n_n4204) & (!x456x) & (n_n704) & (x12824x)) + ((!n_n4205) & (!n_n4204) & (x456x) & (!n_n704) & (!x12824x)) + ((!n_n4205) & (!n_n4204) & (x456x) & (!n_n704) & (x12824x)) + ((!n_n4205) & (!n_n4204) & (x456x) & (n_n704) & (!x12824x)) + ((!n_n4205) & (!n_n4204) & (x456x) & (n_n704) & (x12824x)) + ((!n_n4205) & (n_n4204) & (!x456x) & (!n_n704) & (!x12824x)) + ((!n_n4205) & (n_n4204) & (!x456x) & (!n_n704) & (x12824x)) + ((!n_n4205) & (n_n4204) & (!x456x) & (n_n704) & (!x12824x)) + ((!n_n4205) & (n_n4204) & (!x456x) & (n_n704) & (x12824x)) + ((!n_n4205) & (n_n4204) & (x456x) & (!n_n704) & (!x12824x)) + ((!n_n4205) & (n_n4204) & (x456x) & (!n_n704) & (x12824x)) + ((!n_n4205) & (n_n4204) & (x456x) & (n_n704) & (!x12824x)) + ((!n_n4205) & (n_n4204) & (x456x) & (n_n704) & (x12824x)) + ((n_n4205) & (!n_n4204) & (!x456x) & (!n_n704) & (!x12824x)) + ((n_n4205) & (!n_n4204) & (!x456x) & (!n_n704) & (x12824x)) + ((n_n4205) & (!n_n4204) & (!x456x) & (n_n704) & (!x12824x)) + ((n_n4205) & (!n_n4204) & (!x456x) & (n_n704) & (x12824x)) + ((n_n4205) & (!n_n4204) & (x456x) & (!n_n704) & (!x12824x)) + ((n_n4205) & (!n_n4204) & (x456x) & (!n_n704) & (x12824x)) + ((n_n4205) & (!n_n4204) & (x456x) & (n_n704) & (!x12824x)) + ((n_n4205) & (!n_n4204) & (x456x) & (n_n704) & (x12824x)) + ((n_n4205) & (n_n4204) & (!x456x) & (!n_n704) & (!x12824x)) + ((n_n4205) & (n_n4204) & (!x456x) & (!n_n704) & (x12824x)) + ((n_n4205) & (n_n4204) & (!x456x) & (n_n704) & (!x12824x)) + ((n_n4205) & (n_n4204) & (!x456x) & (n_n704) & (x12824x)) + ((n_n4205) & (n_n4204) & (x456x) & (!n_n704) & (!x12824x)) + ((n_n4205) & (n_n4204) & (x456x) & (!n_n704) & (x12824x)) + ((n_n4205) & (n_n4204) & (x456x) & (n_n704) & (!x12824x)) + ((n_n4205) & (n_n4204) & (x456x) & (n_n704) & (x12824x)));
	assign n_n689 = (((!n_n4952) & (!n_n4949) & (!n_n4959) & (!n_n4957) & (x12834x)) + ((!n_n4952) & (!n_n4949) & (!n_n4959) & (n_n4957) & (!x12834x)) + ((!n_n4952) & (!n_n4949) & (!n_n4959) & (n_n4957) & (x12834x)) + ((!n_n4952) & (!n_n4949) & (n_n4959) & (!n_n4957) & (!x12834x)) + ((!n_n4952) & (!n_n4949) & (n_n4959) & (!n_n4957) & (x12834x)) + ((!n_n4952) & (!n_n4949) & (n_n4959) & (n_n4957) & (!x12834x)) + ((!n_n4952) & (!n_n4949) & (n_n4959) & (n_n4957) & (x12834x)) + ((!n_n4952) & (n_n4949) & (!n_n4959) & (!n_n4957) & (!x12834x)) + ((!n_n4952) & (n_n4949) & (!n_n4959) & (!n_n4957) & (x12834x)) + ((!n_n4952) & (n_n4949) & (!n_n4959) & (n_n4957) & (!x12834x)) + ((!n_n4952) & (n_n4949) & (!n_n4959) & (n_n4957) & (x12834x)) + ((!n_n4952) & (n_n4949) & (n_n4959) & (!n_n4957) & (!x12834x)) + ((!n_n4952) & (n_n4949) & (n_n4959) & (!n_n4957) & (x12834x)) + ((!n_n4952) & (n_n4949) & (n_n4959) & (n_n4957) & (!x12834x)) + ((!n_n4952) & (n_n4949) & (n_n4959) & (n_n4957) & (x12834x)) + ((n_n4952) & (!n_n4949) & (!n_n4959) & (!n_n4957) & (!x12834x)) + ((n_n4952) & (!n_n4949) & (!n_n4959) & (!n_n4957) & (x12834x)) + ((n_n4952) & (!n_n4949) & (!n_n4959) & (n_n4957) & (!x12834x)) + ((n_n4952) & (!n_n4949) & (!n_n4959) & (n_n4957) & (x12834x)) + ((n_n4952) & (!n_n4949) & (n_n4959) & (!n_n4957) & (!x12834x)) + ((n_n4952) & (!n_n4949) & (n_n4959) & (!n_n4957) & (x12834x)) + ((n_n4952) & (!n_n4949) & (n_n4959) & (n_n4957) & (!x12834x)) + ((n_n4952) & (!n_n4949) & (n_n4959) & (n_n4957) & (x12834x)) + ((n_n4952) & (n_n4949) & (!n_n4959) & (!n_n4957) & (!x12834x)) + ((n_n4952) & (n_n4949) & (!n_n4959) & (!n_n4957) & (x12834x)) + ((n_n4952) & (n_n4949) & (!n_n4959) & (n_n4957) & (!x12834x)) + ((n_n4952) & (n_n4949) & (!n_n4959) & (n_n4957) & (x12834x)) + ((n_n4952) & (n_n4949) & (n_n4959) & (!n_n4957) & (!x12834x)) + ((n_n4952) & (n_n4949) & (n_n4959) & (!n_n4957) & (x12834x)) + ((n_n4952) & (n_n4949) & (n_n4959) & (n_n4957) & (!x12834x)) + ((n_n4952) & (n_n4949) & (n_n4959) & (n_n4957) & (x12834x)));
	assign x12840x = (((!n_n4960) & (!n_n4964) & (!n_n4938) & (n_n4933)) + ((!n_n4960) & (!n_n4964) & (n_n4938) & (!n_n4933)) + ((!n_n4960) & (!n_n4964) & (n_n4938) & (n_n4933)) + ((!n_n4960) & (n_n4964) & (!n_n4938) & (!n_n4933)) + ((!n_n4960) & (n_n4964) & (!n_n4938) & (n_n4933)) + ((!n_n4960) & (n_n4964) & (n_n4938) & (!n_n4933)) + ((!n_n4960) & (n_n4964) & (n_n4938) & (n_n4933)) + ((n_n4960) & (!n_n4964) & (!n_n4938) & (!n_n4933)) + ((n_n4960) & (!n_n4964) & (!n_n4938) & (n_n4933)) + ((n_n4960) & (!n_n4964) & (n_n4938) & (!n_n4933)) + ((n_n4960) & (!n_n4964) & (n_n4938) & (n_n4933)) + ((n_n4960) & (n_n4964) & (!n_n4938) & (!n_n4933)) + ((n_n4960) & (n_n4964) & (!n_n4938) & (n_n4933)) + ((n_n4960) & (n_n4964) & (n_n4938) & (!n_n4933)) + ((n_n4960) & (n_n4964) & (n_n4938) & (n_n4933)));
	assign x12841x = (((!n_n4934) & (!n_n3805) & (!n_n4935) & (n_n4971)) + ((!n_n4934) & (!n_n3805) & (n_n4935) & (!n_n4971)) + ((!n_n4934) & (!n_n3805) & (n_n4935) & (n_n4971)) + ((!n_n4934) & (n_n3805) & (!n_n4935) & (!n_n4971)) + ((!n_n4934) & (n_n3805) & (!n_n4935) & (n_n4971)) + ((!n_n4934) & (n_n3805) & (n_n4935) & (!n_n4971)) + ((!n_n4934) & (n_n3805) & (n_n4935) & (n_n4971)) + ((n_n4934) & (!n_n3805) & (!n_n4935) & (!n_n4971)) + ((n_n4934) & (!n_n3805) & (!n_n4935) & (n_n4971)) + ((n_n4934) & (!n_n3805) & (n_n4935) & (!n_n4971)) + ((n_n4934) & (!n_n3805) & (n_n4935) & (n_n4971)) + ((n_n4934) & (n_n3805) & (!n_n4935) & (!n_n4971)) + ((n_n4934) & (n_n3805) & (!n_n4935) & (n_n4971)) + ((n_n4934) & (n_n3805) & (n_n4935) & (!n_n4971)) + ((n_n4934) & (n_n3805) & (n_n4935) & (n_n4971)));
	assign x12842x = (((!n_n4963) & (!n_n4962) & (!x411x) & (!x341x) & (x362x)) + ((!n_n4963) & (!n_n4962) & (!x411x) & (x341x) & (!x362x)) + ((!n_n4963) & (!n_n4962) & (!x411x) & (x341x) & (x362x)) + ((!n_n4963) & (!n_n4962) & (x411x) & (!x341x) & (!x362x)) + ((!n_n4963) & (!n_n4962) & (x411x) & (!x341x) & (x362x)) + ((!n_n4963) & (!n_n4962) & (x411x) & (x341x) & (!x362x)) + ((!n_n4963) & (!n_n4962) & (x411x) & (x341x) & (x362x)) + ((!n_n4963) & (n_n4962) & (!x411x) & (!x341x) & (!x362x)) + ((!n_n4963) & (n_n4962) & (!x411x) & (!x341x) & (x362x)) + ((!n_n4963) & (n_n4962) & (!x411x) & (x341x) & (!x362x)) + ((!n_n4963) & (n_n4962) & (!x411x) & (x341x) & (x362x)) + ((!n_n4963) & (n_n4962) & (x411x) & (!x341x) & (!x362x)) + ((!n_n4963) & (n_n4962) & (x411x) & (!x341x) & (x362x)) + ((!n_n4963) & (n_n4962) & (x411x) & (x341x) & (!x362x)) + ((!n_n4963) & (n_n4962) & (x411x) & (x341x) & (x362x)) + ((n_n4963) & (!n_n4962) & (!x411x) & (!x341x) & (!x362x)) + ((n_n4963) & (!n_n4962) & (!x411x) & (!x341x) & (x362x)) + ((n_n4963) & (!n_n4962) & (!x411x) & (x341x) & (!x362x)) + ((n_n4963) & (!n_n4962) & (!x411x) & (x341x) & (x362x)) + ((n_n4963) & (!n_n4962) & (x411x) & (!x341x) & (!x362x)) + ((n_n4963) & (!n_n4962) & (x411x) & (!x341x) & (x362x)) + ((n_n4963) & (!n_n4962) & (x411x) & (x341x) & (!x362x)) + ((n_n4963) & (!n_n4962) & (x411x) & (x341x) & (x362x)) + ((n_n4963) & (n_n4962) & (!x411x) & (!x341x) & (!x362x)) + ((n_n4963) & (n_n4962) & (!x411x) & (!x341x) & (x362x)) + ((n_n4963) & (n_n4962) & (!x411x) & (x341x) & (!x362x)) + ((n_n4963) & (n_n4962) & (!x411x) & (x341x) & (x362x)) + ((n_n4963) & (n_n4962) & (x411x) & (!x341x) & (!x362x)) + ((n_n4963) & (n_n4962) & (x411x) & (!x341x) & (x362x)) + ((n_n4963) & (n_n4962) & (x411x) & (x341x) & (!x362x)) + ((n_n4963) & (n_n4962) & (x411x) & (x341x) & (x362x)));
	assign n_n642 = (((!n_n689) & (!x12840x) & (!x12841x) & (x12842x)) + ((!n_n689) & (!x12840x) & (x12841x) & (!x12842x)) + ((!n_n689) & (!x12840x) & (x12841x) & (x12842x)) + ((!n_n689) & (x12840x) & (!x12841x) & (!x12842x)) + ((!n_n689) & (x12840x) & (!x12841x) & (x12842x)) + ((!n_n689) & (x12840x) & (x12841x) & (!x12842x)) + ((!n_n689) & (x12840x) & (x12841x) & (x12842x)) + ((n_n689) & (!x12840x) & (!x12841x) & (!x12842x)) + ((n_n689) & (!x12840x) & (!x12841x) & (x12842x)) + ((n_n689) & (!x12840x) & (x12841x) & (!x12842x)) + ((n_n689) & (!x12840x) & (x12841x) & (x12842x)) + ((n_n689) & (x12840x) & (!x12841x) & (!x12842x)) + ((n_n689) & (x12840x) & (!x12841x) & (x12842x)) + ((n_n689) & (x12840x) & (x12841x) & (!x12842x)) + ((n_n689) & (x12840x) & (x12841x) & (x12842x)));
	assign n_n686 = (((!n_n4983) & (!x134x) & (!n_n4984) & (!n_n4986) & (!x22131x)) + ((!n_n4983) & (!x134x) & (!n_n4984) & (n_n4986) & (!x22131x)) + ((!n_n4983) & (!x134x) & (!n_n4984) & (n_n4986) & (x22131x)) + ((!n_n4983) & (!x134x) & (n_n4984) & (!n_n4986) & (!x22131x)) + ((!n_n4983) & (!x134x) & (n_n4984) & (!n_n4986) & (x22131x)) + ((!n_n4983) & (!x134x) & (n_n4984) & (n_n4986) & (!x22131x)) + ((!n_n4983) & (!x134x) & (n_n4984) & (n_n4986) & (x22131x)) + ((!n_n4983) & (x134x) & (!n_n4984) & (!n_n4986) & (!x22131x)) + ((!n_n4983) & (x134x) & (!n_n4984) & (!n_n4986) & (x22131x)) + ((!n_n4983) & (x134x) & (!n_n4984) & (n_n4986) & (!x22131x)) + ((!n_n4983) & (x134x) & (!n_n4984) & (n_n4986) & (x22131x)) + ((!n_n4983) & (x134x) & (n_n4984) & (!n_n4986) & (!x22131x)) + ((!n_n4983) & (x134x) & (n_n4984) & (!n_n4986) & (x22131x)) + ((!n_n4983) & (x134x) & (n_n4984) & (n_n4986) & (!x22131x)) + ((!n_n4983) & (x134x) & (n_n4984) & (n_n4986) & (x22131x)) + ((n_n4983) & (!x134x) & (!n_n4984) & (!n_n4986) & (!x22131x)) + ((n_n4983) & (!x134x) & (!n_n4984) & (!n_n4986) & (x22131x)) + ((n_n4983) & (!x134x) & (!n_n4984) & (n_n4986) & (!x22131x)) + ((n_n4983) & (!x134x) & (!n_n4984) & (n_n4986) & (x22131x)) + ((n_n4983) & (!x134x) & (n_n4984) & (!n_n4986) & (!x22131x)) + ((n_n4983) & (!x134x) & (n_n4984) & (!n_n4986) & (x22131x)) + ((n_n4983) & (!x134x) & (n_n4984) & (n_n4986) & (!x22131x)) + ((n_n4983) & (!x134x) & (n_n4984) & (n_n4986) & (x22131x)) + ((n_n4983) & (x134x) & (!n_n4984) & (!n_n4986) & (!x22131x)) + ((n_n4983) & (x134x) & (!n_n4984) & (!n_n4986) & (x22131x)) + ((n_n4983) & (x134x) & (!n_n4984) & (n_n4986) & (!x22131x)) + ((n_n4983) & (x134x) & (!n_n4984) & (n_n4986) & (x22131x)) + ((n_n4983) & (x134x) & (n_n4984) & (!n_n4986) & (!x22131x)) + ((n_n4983) & (x134x) & (n_n4984) & (!n_n4986) & (x22131x)) + ((n_n4983) & (x134x) & (n_n4984) & (n_n4986) & (!x22131x)) + ((n_n4983) & (x134x) & (n_n4984) & (n_n4986) & (x22131x)));
	assign x12854x = (((!n_n4975) & (!n_n4999) & (!n_n4981) & (n_n5002)) + ((!n_n4975) & (!n_n4999) & (n_n4981) & (!n_n5002)) + ((!n_n4975) & (!n_n4999) & (n_n4981) & (n_n5002)) + ((!n_n4975) & (n_n4999) & (!n_n4981) & (!n_n5002)) + ((!n_n4975) & (n_n4999) & (!n_n4981) & (n_n5002)) + ((!n_n4975) & (n_n4999) & (n_n4981) & (!n_n5002)) + ((!n_n4975) & (n_n4999) & (n_n4981) & (n_n5002)) + ((n_n4975) & (!n_n4999) & (!n_n4981) & (!n_n5002)) + ((n_n4975) & (!n_n4999) & (!n_n4981) & (n_n5002)) + ((n_n4975) & (!n_n4999) & (n_n4981) & (!n_n5002)) + ((n_n4975) & (!n_n4999) & (n_n4981) & (n_n5002)) + ((n_n4975) & (n_n4999) & (!n_n4981) & (!n_n5002)) + ((n_n4975) & (n_n4999) & (!n_n4981) & (n_n5002)) + ((n_n4975) & (n_n4999) & (n_n4981) & (!n_n5002)) + ((n_n4975) & (n_n4999) & (n_n4981) & (n_n5002)));
	assign x12856x = (((!x103x) & (!x252x) & (!x247x) & (!n_n4979) & (n_n4978)) + ((!x103x) & (!x252x) & (!x247x) & (n_n4979) & (!n_n4978)) + ((!x103x) & (!x252x) & (!x247x) & (n_n4979) & (n_n4978)) + ((!x103x) & (!x252x) & (x247x) & (!n_n4979) & (!n_n4978)) + ((!x103x) & (!x252x) & (x247x) & (!n_n4979) & (n_n4978)) + ((!x103x) & (!x252x) & (x247x) & (n_n4979) & (!n_n4978)) + ((!x103x) & (!x252x) & (x247x) & (n_n4979) & (n_n4978)) + ((!x103x) & (x252x) & (!x247x) & (!n_n4979) & (!n_n4978)) + ((!x103x) & (x252x) & (!x247x) & (!n_n4979) & (n_n4978)) + ((!x103x) & (x252x) & (!x247x) & (n_n4979) & (!n_n4978)) + ((!x103x) & (x252x) & (!x247x) & (n_n4979) & (n_n4978)) + ((!x103x) & (x252x) & (x247x) & (!n_n4979) & (!n_n4978)) + ((!x103x) & (x252x) & (x247x) & (!n_n4979) & (n_n4978)) + ((!x103x) & (x252x) & (x247x) & (n_n4979) & (!n_n4978)) + ((!x103x) & (x252x) & (x247x) & (n_n4979) & (n_n4978)) + ((x103x) & (!x252x) & (!x247x) & (!n_n4979) & (!n_n4978)) + ((x103x) & (!x252x) & (!x247x) & (!n_n4979) & (n_n4978)) + ((x103x) & (!x252x) & (!x247x) & (n_n4979) & (!n_n4978)) + ((x103x) & (!x252x) & (!x247x) & (n_n4979) & (n_n4978)) + ((x103x) & (!x252x) & (x247x) & (!n_n4979) & (!n_n4978)) + ((x103x) & (!x252x) & (x247x) & (!n_n4979) & (n_n4978)) + ((x103x) & (!x252x) & (x247x) & (n_n4979) & (!n_n4978)) + ((x103x) & (!x252x) & (x247x) & (n_n4979) & (n_n4978)) + ((x103x) & (x252x) & (!x247x) & (!n_n4979) & (!n_n4978)) + ((x103x) & (x252x) & (!x247x) & (!n_n4979) & (n_n4978)) + ((x103x) & (x252x) & (!x247x) & (n_n4979) & (!n_n4978)) + ((x103x) & (x252x) & (!x247x) & (n_n4979) & (n_n4978)) + ((x103x) & (x252x) & (x247x) & (!n_n4979) & (!n_n4978)) + ((x103x) & (x252x) & (x247x) & (!n_n4979) & (n_n4978)) + ((x103x) & (x252x) & (x247x) & (n_n4979) & (!n_n4978)) + ((x103x) & (x252x) & (x247x) & (n_n4979) & (n_n4978)));
	assign n_n641 = (((!x29x) & (!n_n801) & (!n_n686) & (!x12854x) & (x12856x)) + ((!x29x) & (!n_n801) & (!n_n686) & (x12854x) & (!x12856x)) + ((!x29x) & (!n_n801) & (!n_n686) & (x12854x) & (x12856x)) + ((!x29x) & (!n_n801) & (n_n686) & (!x12854x) & (!x12856x)) + ((!x29x) & (!n_n801) & (n_n686) & (!x12854x) & (x12856x)) + ((!x29x) & (!n_n801) & (n_n686) & (x12854x) & (!x12856x)) + ((!x29x) & (!n_n801) & (n_n686) & (x12854x) & (x12856x)) + ((!x29x) & (n_n801) & (!n_n686) & (!x12854x) & (!x12856x)) + ((!x29x) & (n_n801) & (!n_n686) & (!x12854x) & (x12856x)) + ((!x29x) & (n_n801) & (!n_n686) & (x12854x) & (!x12856x)) + ((!x29x) & (n_n801) & (!n_n686) & (x12854x) & (x12856x)) + ((!x29x) & (n_n801) & (n_n686) & (!x12854x) & (!x12856x)) + ((!x29x) & (n_n801) & (n_n686) & (!x12854x) & (x12856x)) + ((!x29x) & (n_n801) & (n_n686) & (x12854x) & (!x12856x)) + ((!x29x) & (n_n801) & (n_n686) & (x12854x) & (x12856x)) + ((x29x) & (!n_n801) & (!n_n686) & (!x12854x) & (!x12856x)) + ((x29x) & (!n_n801) & (!n_n686) & (!x12854x) & (x12856x)) + ((x29x) & (!n_n801) & (!n_n686) & (x12854x) & (!x12856x)) + ((x29x) & (!n_n801) & (!n_n686) & (x12854x) & (x12856x)) + ((x29x) & (!n_n801) & (n_n686) & (!x12854x) & (!x12856x)) + ((x29x) & (!n_n801) & (n_n686) & (!x12854x) & (x12856x)) + ((x29x) & (!n_n801) & (n_n686) & (x12854x) & (!x12856x)) + ((x29x) & (!n_n801) & (n_n686) & (x12854x) & (x12856x)) + ((x29x) & (n_n801) & (!n_n686) & (!x12854x) & (!x12856x)) + ((x29x) & (n_n801) & (!n_n686) & (!x12854x) & (x12856x)) + ((x29x) & (n_n801) & (!n_n686) & (x12854x) & (!x12856x)) + ((x29x) & (n_n801) & (!n_n686) & (x12854x) & (x12856x)) + ((x29x) & (n_n801) & (n_n686) & (!x12854x) & (!x12856x)) + ((x29x) & (n_n801) & (n_n686) & (!x12854x) & (x12856x)) + ((x29x) & (n_n801) & (n_n686) & (x12854x) & (!x12856x)) + ((x29x) & (n_n801) & (n_n686) & (x12854x) & (x12856x)));
	assign x12865x = (((!n_n691) & (!x12724x) & (!x12725x) & (x12863x)) + ((!n_n691) & (!x12724x) & (x12725x) & (!x12863x)) + ((!n_n691) & (!x12724x) & (x12725x) & (x12863x)) + ((!n_n691) & (x12724x) & (!x12725x) & (!x12863x)) + ((!n_n691) & (x12724x) & (!x12725x) & (x12863x)) + ((!n_n691) & (x12724x) & (x12725x) & (!x12863x)) + ((!n_n691) & (x12724x) & (x12725x) & (x12863x)) + ((n_n691) & (!x12724x) & (!x12725x) & (!x12863x)) + ((n_n691) & (!x12724x) & (!x12725x) & (x12863x)) + ((n_n691) & (!x12724x) & (x12725x) & (!x12863x)) + ((n_n691) & (!x12724x) & (x12725x) & (x12863x)) + ((n_n691) & (x12724x) & (!x12725x) & (!x12863x)) + ((n_n691) & (x12724x) & (!x12725x) & (x12863x)) + ((n_n691) & (x12724x) & (x12725x) & (!x12863x)) + ((n_n691) & (x12724x) & (x12725x) & (x12863x)));
	assign x13657x = (((!n_n4608) & (!n_n4639) & (!n_n4646) & (!n_n4611) & (n_n4647)) + ((!n_n4608) & (!n_n4639) & (!n_n4646) & (n_n4611) & (!n_n4647)) + ((!n_n4608) & (!n_n4639) & (!n_n4646) & (n_n4611) & (n_n4647)) + ((!n_n4608) & (!n_n4639) & (n_n4646) & (!n_n4611) & (!n_n4647)) + ((!n_n4608) & (!n_n4639) & (n_n4646) & (!n_n4611) & (n_n4647)) + ((!n_n4608) & (!n_n4639) & (n_n4646) & (n_n4611) & (!n_n4647)) + ((!n_n4608) & (!n_n4639) & (n_n4646) & (n_n4611) & (n_n4647)) + ((!n_n4608) & (n_n4639) & (!n_n4646) & (!n_n4611) & (!n_n4647)) + ((!n_n4608) & (n_n4639) & (!n_n4646) & (!n_n4611) & (n_n4647)) + ((!n_n4608) & (n_n4639) & (!n_n4646) & (n_n4611) & (!n_n4647)) + ((!n_n4608) & (n_n4639) & (!n_n4646) & (n_n4611) & (n_n4647)) + ((!n_n4608) & (n_n4639) & (n_n4646) & (!n_n4611) & (!n_n4647)) + ((!n_n4608) & (n_n4639) & (n_n4646) & (!n_n4611) & (n_n4647)) + ((!n_n4608) & (n_n4639) & (n_n4646) & (n_n4611) & (!n_n4647)) + ((!n_n4608) & (n_n4639) & (n_n4646) & (n_n4611) & (n_n4647)) + ((n_n4608) & (!n_n4639) & (!n_n4646) & (!n_n4611) & (!n_n4647)) + ((n_n4608) & (!n_n4639) & (!n_n4646) & (!n_n4611) & (n_n4647)) + ((n_n4608) & (!n_n4639) & (!n_n4646) & (n_n4611) & (!n_n4647)) + ((n_n4608) & (!n_n4639) & (!n_n4646) & (n_n4611) & (n_n4647)) + ((n_n4608) & (!n_n4639) & (n_n4646) & (!n_n4611) & (!n_n4647)) + ((n_n4608) & (!n_n4639) & (n_n4646) & (!n_n4611) & (n_n4647)) + ((n_n4608) & (!n_n4639) & (n_n4646) & (n_n4611) & (!n_n4647)) + ((n_n4608) & (!n_n4639) & (n_n4646) & (n_n4611) & (n_n4647)) + ((n_n4608) & (n_n4639) & (!n_n4646) & (!n_n4611) & (!n_n4647)) + ((n_n4608) & (n_n4639) & (!n_n4646) & (!n_n4611) & (n_n4647)) + ((n_n4608) & (n_n4639) & (!n_n4646) & (n_n4611) & (!n_n4647)) + ((n_n4608) & (n_n4639) & (!n_n4646) & (n_n4611) & (n_n4647)) + ((n_n4608) & (n_n4639) & (n_n4646) & (!n_n4611) & (!n_n4647)) + ((n_n4608) & (n_n4639) & (n_n4646) & (!n_n4611) & (n_n4647)) + ((n_n4608) & (n_n4639) & (n_n4646) & (n_n4611) & (!n_n4647)) + ((n_n4608) & (n_n4639) & (n_n4646) & (n_n4611) & (n_n4647)));
	assign x14467x = (((!n_n4361) & (!n_n4363) & (!n_n4358) & (!n_n4356) & (n_n4354)) + ((!n_n4361) & (!n_n4363) & (!n_n4358) & (n_n4356) & (!n_n4354)) + ((!n_n4361) & (!n_n4363) & (!n_n4358) & (n_n4356) & (n_n4354)) + ((!n_n4361) & (!n_n4363) & (n_n4358) & (!n_n4356) & (!n_n4354)) + ((!n_n4361) & (!n_n4363) & (n_n4358) & (!n_n4356) & (n_n4354)) + ((!n_n4361) & (!n_n4363) & (n_n4358) & (n_n4356) & (!n_n4354)) + ((!n_n4361) & (!n_n4363) & (n_n4358) & (n_n4356) & (n_n4354)) + ((!n_n4361) & (n_n4363) & (!n_n4358) & (!n_n4356) & (!n_n4354)) + ((!n_n4361) & (n_n4363) & (!n_n4358) & (!n_n4356) & (n_n4354)) + ((!n_n4361) & (n_n4363) & (!n_n4358) & (n_n4356) & (!n_n4354)) + ((!n_n4361) & (n_n4363) & (!n_n4358) & (n_n4356) & (n_n4354)) + ((!n_n4361) & (n_n4363) & (n_n4358) & (!n_n4356) & (!n_n4354)) + ((!n_n4361) & (n_n4363) & (n_n4358) & (!n_n4356) & (n_n4354)) + ((!n_n4361) & (n_n4363) & (n_n4358) & (n_n4356) & (!n_n4354)) + ((!n_n4361) & (n_n4363) & (n_n4358) & (n_n4356) & (n_n4354)) + ((n_n4361) & (!n_n4363) & (!n_n4358) & (!n_n4356) & (!n_n4354)) + ((n_n4361) & (!n_n4363) & (!n_n4358) & (!n_n4356) & (n_n4354)) + ((n_n4361) & (!n_n4363) & (!n_n4358) & (n_n4356) & (!n_n4354)) + ((n_n4361) & (!n_n4363) & (!n_n4358) & (n_n4356) & (n_n4354)) + ((n_n4361) & (!n_n4363) & (n_n4358) & (!n_n4356) & (!n_n4354)) + ((n_n4361) & (!n_n4363) & (n_n4358) & (!n_n4356) & (n_n4354)) + ((n_n4361) & (!n_n4363) & (n_n4358) & (n_n4356) & (!n_n4354)) + ((n_n4361) & (!n_n4363) & (n_n4358) & (n_n4356) & (n_n4354)) + ((n_n4361) & (n_n4363) & (!n_n4358) & (!n_n4356) & (!n_n4354)) + ((n_n4361) & (n_n4363) & (!n_n4358) & (!n_n4356) & (n_n4354)) + ((n_n4361) & (n_n4363) & (!n_n4358) & (n_n4356) & (!n_n4354)) + ((n_n4361) & (n_n4363) & (!n_n4358) & (n_n4356) & (n_n4354)) + ((n_n4361) & (n_n4363) & (n_n4358) & (!n_n4356) & (!n_n4354)) + ((n_n4361) & (n_n4363) & (n_n4358) & (!n_n4356) & (n_n4354)) + ((n_n4361) & (n_n4363) & (n_n4358) & (n_n4356) & (!n_n4354)) + ((n_n4361) & (n_n4363) & (n_n4358) & (n_n4356) & (n_n4354)));
	assign x14739x = (((!n_n260) & (!n_n491) & (!x20x) & (!n_n4905) & (n_n2718)) + ((!n_n260) & (!n_n491) & (!x20x) & (n_n4905) & (!n_n2718)) + ((!n_n260) & (!n_n491) & (!x20x) & (n_n4905) & (n_n2718)) + ((!n_n260) & (!n_n491) & (x20x) & (!n_n4905) & (n_n2718)) + ((!n_n260) & (!n_n491) & (x20x) & (n_n4905) & (!n_n2718)) + ((!n_n260) & (!n_n491) & (x20x) & (n_n4905) & (n_n2718)) + ((!n_n260) & (n_n491) & (!x20x) & (!n_n4905) & (n_n2718)) + ((!n_n260) & (n_n491) & (!x20x) & (n_n4905) & (!n_n2718)) + ((!n_n260) & (n_n491) & (!x20x) & (n_n4905) & (n_n2718)) + ((!n_n260) & (n_n491) & (x20x) & (!n_n4905) & (n_n2718)) + ((!n_n260) & (n_n491) & (x20x) & (n_n4905) & (!n_n2718)) + ((!n_n260) & (n_n491) & (x20x) & (n_n4905) & (n_n2718)) + ((n_n260) & (!n_n491) & (!x20x) & (!n_n4905) & (n_n2718)) + ((n_n260) & (!n_n491) & (!x20x) & (n_n4905) & (!n_n2718)) + ((n_n260) & (!n_n491) & (!x20x) & (n_n4905) & (n_n2718)) + ((n_n260) & (!n_n491) & (x20x) & (!n_n4905) & (n_n2718)) + ((n_n260) & (!n_n491) & (x20x) & (n_n4905) & (!n_n2718)) + ((n_n260) & (!n_n491) & (x20x) & (n_n4905) & (n_n2718)) + ((n_n260) & (n_n491) & (!x20x) & (!n_n4905) & (n_n2718)) + ((n_n260) & (n_n491) & (!x20x) & (n_n4905) & (!n_n2718)) + ((n_n260) & (n_n491) & (!x20x) & (n_n4905) & (n_n2718)) + ((n_n260) & (n_n491) & (x20x) & (!n_n4905) & (!n_n2718)) + ((n_n260) & (n_n491) & (x20x) & (!n_n4905) & (n_n2718)) + ((n_n260) & (n_n491) & (x20x) & (n_n4905) & (!n_n2718)) + ((n_n260) & (n_n491) & (x20x) & (n_n4905) & (n_n2718)));
	assign x15649x = (((!n_n5321) & (!n_n5326) & (!n_n5323) & (n_n5324)) + ((!n_n5321) & (!n_n5326) & (n_n5323) & (!n_n5324)) + ((!n_n5321) & (!n_n5326) & (n_n5323) & (n_n5324)) + ((!n_n5321) & (n_n5326) & (!n_n5323) & (!n_n5324)) + ((!n_n5321) & (n_n5326) & (!n_n5323) & (n_n5324)) + ((!n_n5321) & (n_n5326) & (n_n5323) & (!n_n5324)) + ((!n_n5321) & (n_n5326) & (n_n5323) & (n_n5324)) + ((n_n5321) & (!n_n5326) & (!n_n5323) & (!n_n5324)) + ((n_n5321) & (!n_n5326) & (!n_n5323) & (n_n5324)) + ((n_n5321) & (!n_n5326) & (n_n5323) & (!n_n5324)) + ((n_n5321) & (!n_n5326) & (n_n5323) & (n_n5324)) + ((n_n5321) & (n_n5326) & (!n_n5323) & (!n_n5324)) + ((n_n5321) & (n_n5326) & (!n_n5323) & (n_n5324)) + ((n_n5321) & (n_n5326) & (n_n5323) & (!n_n5324)) + ((n_n5321) & (n_n5326) & (n_n5323) & (n_n5324)));
	assign x15650x = (((!n_n5318) & (!n_n5320) & (!n_n5322) & (!n_n5317) & (n_n5315)) + ((!n_n5318) & (!n_n5320) & (!n_n5322) & (n_n5317) & (!n_n5315)) + ((!n_n5318) & (!n_n5320) & (!n_n5322) & (n_n5317) & (n_n5315)) + ((!n_n5318) & (!n_n5320) & (n_n5322) & (!n_n5317) & (!n_n5315)) + ((!n_n5318) & (!n_n5320) & (n_n5322) & (!n_n5317) & (n_n5315)) + ((!n_n5318) & (!n_n5320) & (n_n5322) & (n_n5317) & (!n_n5315)) + ((!n_n5318) & (!n_n5320) & (n_n5322) & (n_n5317) & (n_n5315)) + ((!n_n5318) & (n_n5320) & (!n_n5322) & (!n_n5317) & (!n_n5315)) + ((!n_n5318) & (n_n5320) & (!n_n5322) & (!n_n5317) & (n_n5315)) + ((!n_n5318) & (n_n5320) & (!n_n5322) & (n_n5317) & (!n_n5315)) + ((!n_n5318) & (n_n5320) & (!n_n5322) & (n_n5317) & (n_n5315)) + ((!n_n5318) & (n_n5320) & (n_n5322) & (!n_n5317) & (!n_n5315)) + ((!n_n5318) & (n_n5320) & (n_n5322) & (!n_n5317) & (n_n5315)) + ((!n_n5318) & (n_n5320) & (n_n5322) & (n_n5317) & (!n_n5315)) + ((!n_n5318) & (n_n5320) & (n_n5322) & (n_n5317) & (n_n5315)) + ((n_n5318) & (!n_n5320) & (!n_n5322) & (!n_n5317) & (!n_n5315)) + ((n_n5318) & (!n_n5320) & (!n_n5322) & (!n_n5317) & (n_n5315)) + ((n_n5318) & (!n_n5320) & (!n_n5322) & (n_n5317) & (!n_n5315)) + ((n_n5318) & (!n_n5320) & (!n_n5322) & (n_n5317) & (n_n5315)) + ((n_n5318) & (!n_n5320) & (n_n5322) & (!n_n5317) & (!n_n5315)) + ((n_n5318) & (!n_n5320) & (n_n5322) & (!n_n5317) & (n_n5315)) + ((n_n5318) & (!n_n5320) & (n_n5322) & (n_n5317) & (!n_n5315)) + ((n_n5318) & (!n_n5320) & (n_n5322) & (n_n5317) & (n_n5315)) + ((n_n5318) & (n_n5320) & (!n_n5322) & (!n_n5317) & (!n_n5315)) + ((n_n5318) & (n_n5320) & (!n_n5322) & (!n_n5317) & (n_n5315)) + ((n_n5318) & (n_n5320) & (!n_n5322) & (n_n5317) & (!n_n5315)) + ((n_n5318) & (n_n5320) & (!n_n5322) & (n_n5317) & (n_n5315)) + ((n_n5318) & (n_n5320) & (n_n5322) & (!n_n5317) & (!n_n5315)) + ((n_n5318) & (n_n5320) & (n_n5322) & (!n_n5317) & (n_n5315)) + ((n_n5318) & (n_n5320) & (n_n5322) & (n_n5317) & (!n_n5315)) + ((n_n5318) & (n_n5320) & (n_n5322) & (n_n5317) & (n_n5315)));
	assign x15763x = (((!i_7_) & (!i_8_) & (i_6_) & (x14x) & (n_n491)) + ((i_7_) & (i_8_) & (!i_6_) & (x14x) & (n_n491)));
	assign x15766x = (((!n_n4770) & (!n_n4765) & (!x316x) & (!x350x) & (x15763x)) + ((!n_n4770) & (!n_n4765) & (!x316x) & (x350x) & (!x15763x)) + ((!n_n4770) & (!n_n4765) & (!x316x) & (x350x) & (x15763x)) + ((!n_n4770) & (!n_n4765) & (x316x) & (!x350x) & (!x15763x)) + ((!n_n4770) & (!n_n4765) & (x316x) & (!x350x) & (x15763x)) + ((!n_n4770) & (!n_n4765) & (x316x) & (x350x) & (!x15763x)) + ((!n_n4770) & (!n_n4765) & (x316x) & (x350x) & (x15763x)) + ((!n_n4770) & (n_n4765) & (!x316x) & (!x350x) & (!x15763x)) + ((!n_n4770) & (n_n4765) & (!x316x) & (!x350x) & (x15763x)) + ((!n_n4770) & (n_n4765) & (!x316x) & (x350x) & (!x15763x)) + ((!n_n4770) & (n_n4765) & (!x316x) & (x350x) & (x15763x)) + ((!n_n4770) & (n_n4765) & (x316x) & (!x350x) & (!x15763x)) + ((!n_n4770) & (n_n4765) & (x316x) & (!x350x) & (x15763x)) + ((!n_n4770) & (n_n4765) & (x316x) & (x350x) & (!x15763x)) + ((!n_n4770) & (n_n4765) & (x316x) & (x350x) & (x15763x)) + ((n_n4770) & (!n_n4765) & (!x316x) & (!x350x) & (!x15763x)) + ((n_n4770) & (!n_n4765) & (!x316x) & (!x350x) & (x15763x)) + ((n_n4770) & (!n_n4765) & (!x316x) & (x350x) & (!x15763x)) + ((n_n4770) & (!n_n4765) & (!x316x) & (x350x) & (x15763x)) + ((n_n4770) & (!n_n4765) & (x316x) & (!x350x) & (!x15763x)) + ((n_n4770) & (!n_n4765) & (x316x) & (!x350x) & (x15763x)) + ((n_n4770) & (!n_n4765) & (x316x) & (x350x) & (!x15763x)) + ((n_n4770) & (!n_n4765) & (x316x) & (x350x) & (x15763x)) + ((n_n4770) & (n_n4765) & (!x316x) & (!x350x) & (!x15763x)) + ((n_n4770) & (n_n4765) & (!x316x) & (!x350x) & (x15763x)) + ((n_n4770) & (n_n4765) & (!x316x) & (x350x) & (!x15763x)) + ((n_n4770) & (n_n4765) & (!x316x) & (x350x) & (x15763x)) + ((n_n4770) & (n_n4765) & (x316x) & (!x350x) & (!x15763x)) + ((n_n4770) & (n_n4765) & (x316x) & (!x350x) & (x15763x)) + ((n_n4770) & (n_n4765) & (x316x) & (x350x) & (!x15763x)) + ((n_n4770) & (n_n4765) & (x316x) & (x350x) & (x15763x)));
	assign x15329x = (((!n_n4609) & (!n_n4606) & (!n_n4622) & (!n_n4600) & (n_n4623)) + ((!n_n4609) & (!n_n4606) & (!n_n4622) & (n_n4600) & (!n_n4623)) + ((!n_n4609) & (!n_n4606) & (!n_n4622) & (n_n4600) & (n_n4623)) + ((!n_n4609) & (!n_n4606) & (n_n4622) & (!n_n4600) & (!n_n4623)) + ((!n_n4609) & (!n_n4606) & (n_n4622) & (!n_n4600) & (n_n4623)) + ((!n_n4609) & (!n_n4606) & (n_n4622) & (n_n4600) & (!n_n4623)) + ((!n_n4609) & (!n_n4606) & (n_n4622) & (n_n4600) & (n_n4623)) + ((!n_n4609) & (n_n4606) & (!n_n4622) & (!n_n4600) & (!n_n4623)) + ((!n_n4609) & (n_n4606) & (!n_n4622) & (!n_n4600) & (n_n4623)) + ((!n_n4609) & (n_n4606) & (!n_n4622) & (n_n4600) & (!n_n4623)) + ((!n_n4609) & (n_n4606) & (!n_n4622) & (n_n4600) & (n_n4623)) + ((!n_n4609) & (n_n4606) & (n_n4622) & (!n_n4600) & (!n_n4623)) + ((!n_n4609) & (n_n4606) & (n_n4622) & (!n_n4600) & (n_n4623)) + ((!n_n4609) & (n_n4606) & (n_n4622) & (n_n4600) & (!n_n4623)) + ((!n_n4609) & (n_n4606) & (n_n4622) & (n_n4600) & (n_n4623)) + ((n_n4609) & (!n_n4606) & (!n_n4622) & (!n_n4600) & (!n_n4623)) + ((n_n4609) & (!n_n4606) & (!n_n4622) & (!n_n4600) & (n_n4623)) + ((n_n4609) & (!n_n4606) & (!n_n4622) & (n_n4600) & (!n_n4623)) + ((n_n4609) & (!n_n4606) & (!n_n4622) & (n_n4600) & (n_n4623)) + ((n_n4609) & (!n_n4606) & (n_n4622) & (!n_n4600) & (!n_n4623)) + ((n_n4609) & (!n_n4606) & (n_n4622) & (!n_n4600) & (n_n4623)) + ((n_n4609) & (!n_n4606) & (n_n4622) & (n_n4600) & (!n_n4623)) + ((n_n4609) & (!n_n4606) & (n_n4622) & (n_n4600) & (n_n4623)) + ((n_n4609) & (n_n4606) & (!n_n4622) & (!n_n4600) & (!n_n4623)) + ((n_n4609) & (n_n4606) & (!n_n4622) & (!n_n4600) & (n_n4623)) + ((n_n4609) & (n_n4606) & (!n_n4622) & (n_n4600) & (!n_n4623)) + ((n_n4609) & (n_n4606) & (!n_n4622) & (n_n4600) & (n_n4623)) + ((n_n4609) & (n_n4606) & (n_n4622) & (!n_n4600) & (!n_n4623)) + ((n_n4609) & (n_n4606) & (n_n4622) & (!n_n4600) & (n_n4623)) + ((n_n4609) & (n_n4606) & (n_n4622) & (n_n4600) & (!n_n4623)) + ((n_n4609) & (n_n4606) & (n_n4622) & (n_n4600) & (n_n4623)));
	assign x22078x = (((!n_n4344) & (!n_n4347) & (!n_n4349) & (!n_n4348)));
	assign x16080x = (((!i_9_) & (n_n536) & (n_n534) & (n_n535) & (!n_n520)) + ((!i_9_) & (n_n536) & (n_n534) & (n_n535) & (n_n520)) + ((i_9_) & (n_n536) & (!n_n534) & (n_n535) & (n_n520)) + ((i_9_) & (n_n536) & (n_n534) & (n_n535) & (n_n520)));
	assign x16135x = (((!n_n4697) & (!n_n4701) & (!n_n4696) & (!n_n4692) & (n_n4695)) + ((!n_n4697) & (!n_n4701) & (!n_n4696) & (n_n4692) & (!n_n4695)) + ((!n_n4697) & (!n_n4701) & (!n_n4696) & (n_n4692) & (n_n4695)) + ((!n_n4697) & (!n_n4701) & (n_n4696) & (!n_n4692) & (!n_n4695)) + ((!n_n4697) & (!n_n4701) & (n_n4696) & (!n_n4692) & (n_n4695)) + ((!n_n4697) & (!n_n4701) & (n_n4696) & (n_n4692) & (!n_n4695)) + ((!n_n4697) & (!n_n4701) & (n_n4696) & (n_n4692) & (n_n4695)) + ((!n_n4697) & (n_n4701) & (!n_n4696) & (!n_n4692) & (!n_n4695)) + ((!n_n4697) & (n_n4701) & (!n_n4696) & (!n_n4692) & (n_n4695)) + ((!n_n4697) & (n_n4701) & (!n_n4696) & (n_n4692) & (!n_n4695)) + ((!n_n4697) & (n_n4701) & (!n_n4696) & (n_n4692) & (n_n4695)) + ((!n_n4697) & (n_n4701) & (n_n4696) & (!n_n4692) & (!n_n4695)) + ((!n_n4697) & (n_n4701) & (n_n4696) & (!n_n4692) & (n_n4695)) + ((!n_n4697) & (n_n4701) & (n_n4696) & (n_n4692) & (!n_n4695)) + ((!n_n4697) & (n_n4701) & (n_n4696) & (n_n4692) & (n_n4695)) + ((n_n4697) & (!n_n4701) & (!n_n4696) & (!n_n4692) & (!n_n4695)) + ((n_n4697) & (!n_n4701) & (!n_n4696) & (!n_n4692) & (n_n4695)) + ((n_n4697) & (!n_n4701) & (!n_n4696) & (n_n4692) & (!n_n4695)) + ((n_n4697) & (!n_n4701) & (!n_n4696) & (n_n4692) & (n_n4695)) + ((n_n4697) & (!n_n4701) & (n_n4696) & (!n_n4692) & (!n_n4695)) + ((n_n4697) & (!n_n4701) & (n_n4696) & (!n_n4692) & (n_n4695)) + ((n_n4697) & (!n_n4701) & (n_n4696) & (n_n4692) & (!n_n4695)) + ((n_n4697) & (!n_n4701) & (n_n4696) & (n_n4692) & (n_n4695)) + ((n_n4697) & (n_n4701) & (!n_n4696) & (!n_n4692) & (!n_n4695)) + ((n_n4697) & (n_n4701) & (!n_n4696) & (!n_n4692) & (n_n4695)) + ((n_n4697) & (n_n4701) & (!n_n4696) & (n_n4692) & (!n_n4695)) + ((n_n4697) & (n_n4701) & (!n_n4696) & (n_n4692) & (n_n4695)) + ((n_n4697) & (n_n4701) & (n_n4696) & (!n_n4692) & (!n_n4695)) + ((n_n4697) & (n_n4701) & (n_n4696) & (!n_n4692) & (n_n4695)) + ((n_n4697) & (n_n4701) & (n_n4696) & (n_n4692) & (!n_n4695)) + ((n_n4697) & (n_n4701) & (n_n4696) & (n_n4692) & (n_n4695)));
	assign x464x = (((!n_n325) & (!n_n535) & (!x20x) & (!n_n4710) & (n_n4219)) + ((!n_n325) & (!n_n535) & (!x20x) & (n_n4710) & (!n_n4219)) + ((!n_n325) & (!n_n535) & (!x20x) & (n_n4710) & (n_n4219)) + ((!n_n325) & (!n_n535) & (x20x) & (!n_n4710) & (n_n4219)) + ((!n_n325) & (!n_n535) & (x20x) & (n_n4710) & (!n_n4219)) + ((!n_n325) & (!n_n535) & (x20x) & (n_n4710) & (n_n4219)) + ((!n_n325) & (n_n535) & (!x20x) & (!n_n4710) & (n_n4219)) + ((!n_n325) & (n_n535) & (!x20x) & (n_n4710) & (!n_n4219)) + ((!n_n325) & (n_n535) & (!x20x) & (n_n4710) & (n_n4219)) + ((!n_n325) & (n_n535) & (x20x) & (!n_n4710) & (n_n4219)) + ((!n_n325) & (n_n535) & (x20x) & (n_n4710) & (!n_n4219)) + ((!n_n325) & (n_n535) & (x20x) & (n_n4710) & (n_n4219)) + ((n_n325) & (!n_n535) & (!x20x) & (!n_n4710) & (n_n4219)) + ((n_n325) & (!n_n535) & (!x20x) & (n_n4710) & (!n_n4219)) + ((n_n325) & (!n_n535) & (!x20x) & (n_n4710) & (n_n4219)) + ((n_n325) & (!n_n535) & (x20x) & (!n_n4710) & (n_n4219)) + ((n_n325) & (!n_n535) & (x20x) & (n_n4710) & (!n_n4219)) + ((n_n325) & (!n_n535) & (x20x) & (n_n4710) & (n_n4219)) + ((n_n325) & (n_n535) & (!x20x) & (!n_n4710) & (n_n4219)) + ((n_n325) & (n_n535) & (!x20x) & (n_n4710) & (!n_n4219)) + ((n_n325) & (n_n535) & (!x20x) & (n_n4710) & (n_n4219)) + ((n_n325) & (n_n535) & (x20x) & (!n_n4710) & (!n_n4219)) + ((n_n325) & (n_n535) & (x20x) & (!n_n4710) & (n_n4219)) + ((n_n325) & (n_n535) & (x20x) & (n_n4710) & (!n_n4219)) + ((n_n325) & (n_n535) & (x20x) & (n_n4710) & (n_n4219)));
	assign x16144x = (((!x426x) & (!n_n4680) & (!n_n4708) & (!n_n4707) & (x464x)) + ((!x426x) & (!n_n4680) & (!n_n4708) & (n_n4707) & (!x464x)) + ((!x426x) & (!n_n4680) & (!n_n4708) & (n_n4707) & (x464x)) + ((!x426x) & (!n_n4680) & (n_n4708) & (!n_n4707) & (!x464x)) + ((!x426x) & (!n_n4680) & (n_n4708) & (!n_n4707) & (x464x)) + ((!x426x) & (!n_n4680) & (n_n4708) & (n_n4707) & (!x464x)) + ((!x426x) & (!n_n4680) & (n_n4708) & (n_n4707) & (x464x)) + ((!x426x) & (n_n4680) & (!n_n4708) & (!n_n4707) & (!x464x)) + ((!x426x) & (n_n4680) & (!n_n4708) & (!n_n4707) & (x464x)) + ((!x426x) & (n_n4680) & (!n_n4708) & (n_n4707) & (!x464x)) + ((!x426x) & (n_n4680) & (!n_n4708) & (n_n4707) & (x464x)) + ((!x426x) & (n_n4680) & (n_n4708) & (!n_n4707) & (!x464x)) + ((!x426x) & (n_n4680) & (n_n4708) & (!n_n4707) & (x464x)) + ((!x426x) & (n_n4680) & (n_n4708) & (n_n4707) & (!x464x)) + ((!x426x) & (n_n4680) & (n_n4708) & (n_n4707) & (x464x)) + ((x426x) & (!n_n4680) & (!n_n4708) & (!n_n4707) & (!x464x)) + ((x426x) & (!n_n4680) & (!n_n4708) & (!n_n4707) & (x464x)) + ((x426x) & (!n_n4680) & (!n_n4708) & (n_n4707) & (!x464x)) + ((x426x) & (!n_n4680) & (!n_n4708) & (n_n4707) & (x464x)) + ((x426x) & (!n_n4680) & (n_n4708) & (!n_n4707) & (!x464x)) + ((x426x) & (!n_n4680) & (n_n4708) & (!n_n4707) & (x464x)) + ((x426x) & (!n_n4680) & (n_n4708) & (n_n4707) & (!x464x)) + ((x426x) & (!n_n4680) & (n_n4708) & (n_n4707) & (x464x)) + ((x426x) & (n_n4680) & (!n_n4708) & (!n_n4707) & (!x464x)) + ((x426x) & (n_n4680) & (!n_n4708) & (!n_n4707) & (x464x)) + ((x426x) & (n_n4680) & (!n_n4708) & (n_n4707) & (!x464x)) + ((x426x) & (n_n4680) & (!n_n4708) & (n_n4707) & (x464x)) + ((x426x) & (n_n4680) & (n_n4708) & (!n_n4707) & (!x464x)) + ((x426x) & (n_n4680) & (n_n4708) & (!n_n4707) & (x464x)) + ((x426x) & (n_n4680) & (n_n4708) & (n_n4707) & (!x464x)) + ((x426x) & (n_n4680) & (n_n4708) & (n_n4707) & (x464x)));
	assign x16141x = (((!n_n4689) & (!n_n4712) & (!n_n4681) & (n_n4705)) + ((!n_n4689) & (!n_n4712) & (n_n4681) & (!n_n4705)) + ((!n_n4689) & (!n_n4712) & (n_n4681) & (n_n4705)) + ((!n_n4689) & (n_n4712) & (!n_n4681) & (!n_n4705)) + ((!n_n4689) & (n_n4712) & (!n_n4681) & (n_n4705)) + ((!n_n4689) & (n_n4712) & (n_n4681) & (!n_n4705)) + ((!n_n4689) & (n_n4712) & (n_n4681) & (n_n4705)) + ((n_n4689) & (!n_n4712) & (!n_n4681) & (!n_n4705)) + ((n_n4689) & (!n_n4712) & (!n_n4681) & (n_n4705)) + ((n_n4689) & (!n_n4712) & (n_n4681) & (!n_n4705)) + ((n_n4689) & (!n_n4712) & (n_n4681) & (n_n4705)) + ((n_n4689) & (n_n4712) & (!n_n4681) & (!n_n4705)) + ((n_n4689) & (n_n4712) & (!n_n4681) & (n_n4705)) + ((n_n4689) & (n_n4712) & (n_n4681) & (!n_n4705)) + ((n_n4689) & (n_n4712) & (n_n4681) & (n_n4705)));
	assign x22071x = (((!n_n4691) & (!x219x) & (!x80x) & (!x221x) & (!n_n4693)));
	assign x22218x = (((!n_n5201) & (!n_n5199) & (!x223x) & (!n_n5208)));
	assign x16146x = (((!i_7_) & (i_8_) & (!i_6_) & (n_n509) & (x18x)) + ((i_7_) & (i_8_) & (!i_6_) & (n_n509) & (x18x)));
	assign n_n1846 = (((!n_n4999) & (!n_n4986) & (!x41x) & (!x133x) & (x16146x)) + ((!n_n4999) & (!n_n4986) & (!x41x) & (x133x) & (!x16146x)) + ((!n_n4999) & (!n_n4986) & (!x41x) & (x133x) & (x16146x)) + ((!n_n4999) & (!n_n4986) & (x41x) & (!x133x) & (!x16146x)) + ((!n_n4999) & (!n_n4986) & (x41x) & (!x133x) & (x16146x)) + ((!n_n4999) & (!n_n4986) & (x41x) & (x133x) & (!x16146x)) + ((!n_n4999) & (!n_n4986) & (x41x) & (x133x) & (x16146x)) + ((!n_n4999) & (n_n4986) & (!x41x) & (!x133x) & (!x16146x)) + ((!n_n4999) & (n_n4986) & (!x41x) & (!x133x) & (x16146x)) + ((!n_n4999) & (n_n4986) & (!x41x) & (x133x) & (!x16146x)) + ((!n_n4999) & (n_n4986) & (!x41x) & (x133x) & (x16146x)) + ((!n_n4999) & (n_n4986) & (x41x) & (!x133x) & (!x16146x)) + ((!n_n4999) & (n_n4986) & (x41x) & (!x133x) & (x16146x)) + ((!n_n4999) & (n_n4986) & (x41x) & (x133x) & (!x16146x)) + ((!n_n4999) & (n_n4986) & (x41x) & (x133x) & (x16146x)) + ((n_n4999) & (!n_n4986) & (!x41x) & (!x133x) & (!x16146x)) + ((n_n4999) & (!n_n4986) & (!x41x) & (!x133x) & (x16146x)) + ((n_n4999) & (!n_n4986) & (!x41x) & (x133x) & (!x16146x)) + ((n_n4999) & (!n_n4986) & (!x41x) & (x133x) & (x16146x)) + ((n_n4999) & (!n_n4986) & (x41x) & (!x133x) & (!x16146x)) + ((n_n4999) & (!n_n4986) & (x41x) & (!x133x) & (x16146x)) + ((n_n4999) & (!n_n4986) & (x41x) & (x133x) & (!x16146x)) + ((n_n4999) & (!n_n4986) & (x41x) & (x133x) & (x16146x)) + ((n_n4999) & (n_n4986) & (!x41x) & (!x133x) & (!x16146x)) + ((n_n4999) & (n_n4986) & (!x41x) & (!x133x) & (x16146x)) + ((n_n4999) & (n_n4986) & (!x41x) & (x133x) & (!x16146x)) + ((n_n4999) & (n_n4986) & (!x41x) & (x133x) & (x16146x)) + ((n_n4999) & (n_n4986) & (x41x) & (!x133x) & (!x16146x)) + ((n_n4999) & (n_n4986) & (x41x) & (!x133x) & (x16146x)) + ((n_n4999) & (n_n4986) & (x41x) & (x133x) & (!x16146x)) + ((n_n4999) & (n_n4986) & (x41x) & (x133x) & (x16146x)));
	assign x16155x = (((!n_n518) & (!x21x) & (!n_n195) & (!n_n4985) & (x405x)) + ((!n_n518) & (!x21x) & (!n_n195) & (n_n4985) & (!x405x)) + ((!n_n518) & (!x21x) & (!n_n195) & (n_n4985) & (x405x)) + ((!n_n518) & (!x21x) & (n_n195) & (!n_n4985) & (x405x)) + ((!n_n518) & (!x21x) & (n_n195) & (n_n4985) & (!x405x)) + ((!n_n518) & (!x21x) & (n_n195) & (n_n4985) & (x405x)) + ((!n_n518) & (x21x) & (!n_n195) & (!n_n4985) & (x405x)) + ((!n_n518) & (x21x) & (!n_n195) & (n_n4985) & (!x405x)) + ((!n_n518) & (x21x) & (!n_n195) & (n_n4985) & (x405x)) + ((!n_n518) & (x21x) & (n_n195) & (!n_n4985) & (x405x)) + ((!n_n518) & (x21x) & (n_n195) & (n_n4985) & (!x405x)) + ((!n_n518) & (x21x) & (n_n195) & (n_n4985) & (x405x)) + ((n_n518) & (!x21x) & (!n_n195) & (!n_n4985) & (x405x)) + ((n_n518) & (!x21x) & (!n_n195) & (n_n4985) & (!x405x)) + ((n_n518) & (!x21x) & (!n_n195) & (n_n4985) & (x405x)) + ((n_n518) & (!x21x) & (n_n195) & (!n_n4985) & (x405x)) + ((n_n518) & (!x21x) & (n_n195) & (n_n4985) & (!x405x)) + ((n_n518) & (!x21x) & (n_n195) & (n_n4985) & (x405x)) + ((n_n518) & (x21x) & (!n_n195) & (!n_n4985) & (x405x)) + ((n_n518) & (x21x) & (!n_n195) & (n_n4985) & (!x405x)) + ((n_n518) & (x21x) & (!n_n195) & (n_n4985) & (x405x)) + ((n_n518) & (x21x) & (n_n195) & (!n_n4985) & (!x405x)) + ((n_n518) & (x21x) & (n_n195) & (!n_n4985) & (x405x)) + ((n_n518) & (x21x) & (n_n195) & (n_n4985) & (!x405x)) + ((n_n518) & (x21x) & (n_n195) & (n_n4985) & (x405x)));
	assign x16157x = (((!n_n4975) & (!n_n5000) & (!x299x) & (x16155x)) + ((!n_n4975) & (!n_n5000) & (x299x) & (!x16155x)) + ((!n_n4975) & (!n_n5000) & (x299x) & (x16155x)) + ((!n_n4975) & (n_n5000) & (!x299x) & (!x16155x)) + ((!n_n4975) & (n_n5000) & (!x299x) & (x16155x)) + ((!n_n4975) & (n_n5000) & (x299x) & (!x16155x)) + ((!n_n4975) & (n_n5000) & (x299x) & (x16155x)) + ((n_n4975) & (!n_n5000) & (!x299x) & (!x16155x)) + ((n_n4975) & (!n_n5000) & (!x299x) & (x16155x)) + ((n_n4975) & (!n_n5000) & (x299x) & (!x16155x)) + ((n_n4975) & (!n_n5000) & (x299x) & (x16155x)) + ((n_n4975) & (n_n5000) & (!x299x) & (!x16155x)) + ((n_n4975) & (n_n5000) & (!x299x) & (x16155x)) + ((n_n4975) & (n_n5000) & (x299x) & (!x16155x)) + ((n_n4975) & (n_n5000) & (x299x) & (x16155x)));
	assign n_n1852 = (((!n_n4920) & (!n_n4928) & (!x249x) & (!n_n4932) & (x42x)) + ((!n_n4920) & (!n_n4928) & (!x249x) & (n_n4932) & (!x42x)) + ((!n_n4920) & (!n_n4928) & (!x249x) & (n_n4932) & (x42x)) + ((!n_n4920) & (!n_n4928) & (x249x) & (!n_n4932) & (!x42x)) + ((!n_n4920) & (!n_n4928) & (x249x) & (!n_n4932) & (x42x)) + ((!n_n4920) & (!n_n4928) & (x249x) & (n_n4932) & (!x42x)) + ((!n_n4920) & (!n_n4928) & (x249x) & (n_n4932) & (x42x)) + ((!n_n4920) & (n_n4928) & (!x249x) & (!n_n4932) & (!x42x)) + ((!n_n4920) & (n_n4928) & (!x249x) & (!n_n4932) & (x42x)) + ((!n_n4920) & (n_n4928) & (!x249x) & (n_n4932) & (!x42x)) + ((!n_n4920) & (n_n4928) & (!x249x) & (n_n4932) & (x42x)) + ((!n_n4920) & (n_n4928) & (x249x) & (!n_n4932) & (!x42x)) + ((!n_n4920) & (n_n4928) & (x249x) & (!n_n4932) & (x42x)) + ((!n_n4920) & (n_n4928) & (x249x) & (n_n4932) & (!x42x)) + ((!n_n4920) & (n_n4928) & (x249x) & (n_n4932) & (x42x)) + ((n_n4920) & (!n_n4928) & (!x249x) & (!n_n4932) & (!x42x)) + ((n_n4920) & (!n_n4928) & (!x249x) & (!n_n4932) & (x42x)) + ((n_n4920) & (!n_n4928) & (!x249x) & (n_n4932) & (!x42x)) + ((n_n4920) & (!n_n4928) & (!x249x) & (n_n4932) & (x42x)) + ((n_n4920) & (!n_n4928) & (x249x) & (!n_n4932) & (!x42x)) + ((n_n4920) & (!n_n4928) & (x249x) & (!n_n4932) & (x42x)) + ((n_n4920) & (!n_n4928) & (x249x) & (n_n4932) & (!x42x)) + ((n_n4920) & (!n_n4928) & (x249x) & (n_n4932) & (x42x)) + ((n_n4920) & (n_n4928) & (!x249x) & (!n_n4932) & (!x42x)) + ((n_n4920) & (n_n4928) & (!x249x) & (!n_n4932) & (x42x)) + ((n_n4920) & (n_n4928) & (!x249x) & (n_n4932) & (!x42x)) + ((n_n4920) & (n_n4928) & (!x249x) & (n_n4932) & (x42x)) + ((n_n4920) & (n_n4928) & (x249x) & (!n_n4932) & (!x42x)) + ((n_n4920) & (n_n4928) & (x249x) & (!n_n4932) & (x42x)) + ((n_n4920) & (n_n4928) & (x249x) & (n_n4932) & (!x42x)) + ((n_n4920) & (n_n4928) & (x249x) & (n_n4932) & (x42x)));
	assign x16166x = (((!n_n4907) & (!n_n4942) & (!n_n4936) & (n_n4933)) + ((!n_n4907) & (!n_n4942) & (n_n4936) & (!n_n4933)) + ((!n_n4907) & (!n_n4942) & (n_n4936) & (n_n4933)) + ((!n_n4907) & (n_n4942) & (!n_n4936) & (!n_n4933)) + ((!n_n4907) & (n_n4942) & (!n_n4936) & (n_n4933)) + ((!n_n4907) & (n_n4942) & (n_n4936) & (!n_n4933)) + ((!n_n4907) & (n_n4942) & (n_n4936) & (n_n4933)) + ((n_n4907) & (!n_n4942) & (!n_n4936) & (!n_n4933)) + ((n_n4907) & (!n_n4942) & (!n_n4936) & (n_n4933)) + ((n_n4907) & (!n_n4942) & (n_n4936) & (!n_n4933)) + ((n_n4907) & (!n_n4942) & (n_n4936) & (n_n4933)) + ((n_n4907) & (n_n4942) & (!n_n4936) & (!n_n4933)) + ((n_n4907) & (n_n4942) & (!n_n4936) & (n_n4933)) + ((n_n4907) & (n_n4942) & (n_n4936) & (!n_n4933)) + ((n_n4907) & (n_n4942) & (n_n4936) & (n_n4933)));
	assign x16167x = (((!n_n4934) & (!n_n4935) & (!x411x) & (!x331x) & (x305x)) + ((!n_n4934) & (!n_n4935) & (!x411x) & (x331x) & (!x305x)) + ((!n_n4934) & (!n_n4935) & (!x411x) & (x331x) & (x305x)) + ((!n_n4934) & (!n_n4935) & (x411x) & (!x331x) & (!x305x)) + ((!n_n4934) & (!n_n4935) & (x411x) & (!x331x) & (x305x)) + ((!n_n4934) & (!n_n4935) & (x411x) & (x331x) & (!x305x)) + ((!n_n4934) & (!n_n4935) & (x411x) & (x331x) & (x305x)) + ((!n_n4934) & (n_n4935) & (!x411x) & (!x331x) & (!x305x)) + ((!n_n4934) & (n_n4935) & (!x411x) & (!x331x) & (x305x)) + ((!n_n4934) & (n_n4935) & (!x411x) & (x331x) & (!x305x)) + ((!n_n4934) & (n_n4935) & (!x411x) & (x331x) & (x305x)) + ((!n_n4934) & (n_n4935) & (x411x) & (!x331x) & (!x305x)) + ((!n_n4934) & (n_n4935) & (x411x) & (!x331x) & (x305x)) + ((!n_n4934) & (n_n4935) & (x411x) & (x331x) & (!x305x)) + ((!n_n4934) & (n_n4935) & (x411x) & (x331x) & (x305x)) + ((n_n4934) & (!n_n4935) & (!x411x) & (!x331x) & (!x305x)) + ((n_n4934) & (!n_n4935) & (!x411x) & (!x331x) & (x305x)) + ((n_n4934) & (!n_n4935) & (!x411x) & (x331x) & (!x305x)) + ((n_n4934) & (!n_n4935) & (!x411x) & (x331x) & (x305x)) + ((n_n4934) & (!n_n4935) & (x411x) & (!x331x) & (!x305x)) + ((n_n4934) & (!n_n4935) & (x411x) & (!x331x) & (x305x)) + ((n_n4934) & (!n_n4935) & (x411x) & (x331x) & (!x305x)) + ((n_n4934) & (!n_n4935) & (x411x) & (x331x) & (x305x)) + ((n_n4934) & (n_n4935) & (!x411x) & (!x331x) & (!x305x)) + ((n_n4934) & (n_n4935) & (!x411x) & (!x331x) & (x305x)) + ((n_n4934) & (n_n4935) & (!x411x) & (x331x) & (!x305x)) + ((n_n4934) & (n_n4935) & (!x411x) & (x331x) & (x305x)) + ((n_n4934) & (n_n4935) & (x411x) & (!x331x) & (!x305x)) + ((n_n4934) & (n_n4935) & (x411x) & (!x331x) & (x305x)) + ((n_n4934) & (n_n4935) & (x411x) & (x331x) & (!x305x)) + ((n_n4934) & (n_n4935) & (x411x) & (x331x) & (x305x)));
	assign n_n1805 = (((!x138x) & (!n_n1852) & (!x16166x) & (x16167x)) + ((!x138x) & (!n_n1852) & (x16166x) & (!x16167x)) + ((!x138x) & (!n_n1852) & (x16166x) & (x16167x)) + ((!x138x) & (n_n1852) & (!x16166x) & (!x16167x)) + ((!x138x) & (n_n1852) & (!x16166x) & (x16167x)) + ((!x138x) & (n_n1852) & (x16166x) & (!x16167x)) + ((!x138x) & (n_n1852) & (x16166x) & (x16167x)) + ((x138x) & (!n_n1852) & (!x16166x) & (!x16167x)) + ((x138x) & (!n_n1852) & (!x16166x) & (x16167x)) + ((x138x) & (!n_n1852) & (x16166x) & (!x16167x)) + ((x138x) & (!n_n1852) & (x16166x) & (x16167x)) + ((x138x) & (n_n1852) & (!x16166x) & (!x16167x)) + ((x138x) & (n_n1852) & (!x16166x) & (x16167x)) + ((x138x) & (n_n1852) & (x16166x) & (!x16167x)) + ((x138x) & (n_n1852) & (x16166x) & (x16167x)));
	assign n_n1850 = (((!n_n4950) & (!n_n4948) & (!x14962x) & (!x58x) & (x317x)) + ((!n_n4950) & (!n_n4948) & (!x14962x) & (x58x) & (!x317x)) + ((!n_n4950) & (!n_n4948) & (!x14962x) & (x58x) & (x317x)) + ((!n_n4950) & (!n_n4948) & (x14962x) & (!x58x) & (!x317x)) + ((!n_n4950) & (!n_n4948) & (x14962x) & (!x58x) & (x317x)) + ((!n_n4950) & (!n_n4948) & (x14962x) & (x58x) & (!x317x)) + ((!n_n4950) & (!n_n4948) & (x14962x) & (x58x) & (x317x)) + ((!n_n4950) & (n_n4948) & (!x14962x) & (!x58x) & (!x317x)) + ((!n_n4950) & (n_n4948) & (!x14962x) & (!x58x) & (x317x)) + ((!n_n4950) & (n_n4948) & (!x14962x) & (x58x) & (!x317x)) + ((!n_n4950) & (n_n4948) & (!x14962x) & (x58x) & (x317x)) + ((!n_n4950) & (n_n4948) & (x14962x) & (!x58x) & (!x317x)) + ((!n_n4950) & (n_n4948) & (x14962x) & (!x58x) & (x317x)) + ((!n_n4950) & (n_n4948) & (x14962x) & (x58x) & (!x317x)) + ((!n_n4950) & (n_n4948) & (x14962x) & (x58x) & (x317x)) + ((n_n4950) & (!n_n4948) & (!x14962x) & (!x58x) & (!x317x)) + ((n_n4950) & (!n_n4948) & (!x14962x) & (!x58x) & (x317x)) + ((n_n4950) & (!n_n4948) & (!x14962x) & (x58x) & (!x317x)) + ((n_n4950) & (!n_n4948) & (!x14962x) & (x58x) & (x317x)) + ((n_n4950) & (!n_n4948) & (x14962x) & (!x58x) & (!x317x)) + ((n_n4950) & (!n_n4948) & (x14962x) & (!x58x) & (x317x)) + ((n_n4950) & (!n_n4948) & (x14962x) & (x58x) & (!x317x)) + ((n_n4950) & (!n_n4948) & (x14962x) & (x58x) & (x317x)) + ((n_n4950) & (n_n4948) & (!x14962x) & (!x58x) & (!x317x)) + ((n_n4950) & (n_n4948) & (!x14962x) & (!x58x) & (x317x)) + ((n_n4950) & (n_n4948) & (!x14962x) & (x58x) & (!x317x)) + ((n_n4950) & (n_n4948) & (!x14962x) & (x58x) & (x317x)) + ((n_n4950) & (n_n4948) & (x14962x) & (!x58x) & (!x317x)) + ((n_n4950) & (n_n4948) & (x14962x) & (!x58x) & (x317x)) + ((n_n4950) & (n_n4948) & (x14962x) & (x58x) & (!x317x)) + ((n_n4950) & (n_n4948) & (x14962x) & (x58x) & (x317x)));
	assign x16177x = (((!n_n4952) & (!n_n4953) & (!x68x) & (!n_n4954) & (x210x)) + ((!n_n4952) & (!n_n4953) & (!x68x) & (n_n4954) & (!x210x)) + ((!n_n4952) & (!n_n4953) & (!x68x) & (n_n4954) & (x210x)) + ((!n_n4952) & (!n_n4953) & (x68x) & (!n_n4954) & (!x210x)) + ((!n_n4952) & (!n_n4953) & (x68x) & (!n_n4954) & (x210x)) + ((!n_n4952) & (!n_n4953) & (x68x) & (n_n4954) & (!x210x)) + ((!n_n4952) & (!n_n4953) & (x68x) & (n_n4954) & (x210x)) + ((!n_n4952) & (n_n4953) & (!x68x) & (!n_n4954) & (!x210x)) + ((!n_n4952) & (n_n4953) & (!x68x) & (!n_n4954) & (x210x)) + ((!n_n4952) & (n_n4953) & (!x68x) & (n_n4954) & (!x210x)) + ((!n_n4952) & (n_n4953) & (!x68x) & (n_n4954) & (x210x)) + ((!n_n4952) & (n_n4953) & (x68x) & (!n_n4954) & (!x210x)) + ((!n_n4952) & (n_n4953) & (x68x) & (!n_n4954) & (x210x)) + ((!n_n4952) & (n_n4953) & (x68x) & (n_n4954) & (!x210x)) + ((!n_n4952) & (n_n4953) & (x68x) & (n_n4954) & (x210x)) + ((n_n4952) & (!n_n4953) & (!x68x) & (!n_n4954) & (!x210x)) + ((n_n4952) & (!n_n4953) & (!x68x) & (!n_n4954) & (x210x)) + ((n_n4952) & (!n_n4953) & (!x68x) & (n_n4954) & (!x210x)) + ((n_n4952) & (!n_n4953) & (!x68x) & (n_n4954) & (x210x)) + ((n_n4952) & (!n_n4953) & (x68x) & (!n_n4954) & (!x210x)) + ((n_n4952) & (!n_n4953) & (x68x) & (!n_n4954) & (x210x)) + ((n_n4952) & (!n_n4953) & (x68x) & (n_n4954) & (!x210x)) + ((n_n4952) & (!n_n4953) & (x68x) & (n_n4954) & (x210x)) + ((n_n4952) & (n_n4953) & (!x68x) & (!n_n4954) & (!x210x)) + ((n_n4952) & (n_n4953) & (!x68x) & (!n_n4954) & (x210x)) + ((n_n4952) & (n_n4953) & (!x68x) & (n_n4954) & (!x210x)) + ((n_n4952) & (n_n4953) & (!x68x) & (n_n4954) & (x210x)) + ((n_n4952) & (n_n4953) & (x68x) & (!n_n4954) & (!x210x)) + ((n_n4952) & (n_n4953) & (x68x) & (!n_n4954) & (x210x)) + ((n_n4952) & (n_n4953) & (x68x) & (n_n4954) & (!x210x)) + ((n_n4952) & (n_n4953) & (x68x) & (n_n4954) & (x210x)));
	assign x16178x = (((!n_n4962) & (!x29x) & (!n_n4971) & (!n_n4172) & (n_n1970)) + ((!n_n4962) & (!x29x) & (!n_n4971) & (n_n4172) & (!n_n1970)) + ((!n_n4962) & (!x29x) & (!n_n4971) & (n_n4172) & (n_n1970)) + ((!n_n4962) & (!x29x) & (n_n4971) & (!n_n4172) & (!n_n1970)) + ((!n_n4962) & (!x29x) & (n_n4971) & (!n_n4172) & (n_n1970)) + ((!n_n4962) & (!x29x) & (n_n4971) & (n_n4172) & (!n_n1970)) + ((!n_n4962) & (!x29x) & (n_n4971) & (n_n4172) & (n_n1970)) + ((!n_n4962) & (x29x) & (!n_n4971) & (!n_n4172) & (!n_n1970)) + ((!n_n4962) & (x29x) & (!n_n4971) & (!n_n4172) & (n_n1970)) + ((!n_n4962) & (x29x) & (!n_n4971) & (n_n4172) & (!n_n1970)) + ((!n_n4962) & (x29x) & (!n_n4971) & (n_n4172) & (n_n1970)) + ((!n_n4962) & (x29x) & (n_n4971) & (!n_n4172) & (!n_n1970)) + ((!n_n4962) & (x29x) & (n_n4971) & (!n_n4172) & (n_n1970)) + ((!n_n4962) & (x29x) & (n_n4971) & (n_n4172) & (!n_n1970)) + ((!n_n4962) & (x29x) & (n_n4971) & (n_n4172) & (n_n1970)) + ((n_n4962) & (!x29x) & (!n_n4971) & (!n_n4172) & (!n_n1970)) + ((n_n4962) & (!x29x) & (!n_n4971) & (!n_n4172) & (n_n1970)) + ((n_n4962) & (!x29x) & (!n_n4971) & (n_n4172) & (!n_n1970)) + ((n_n4962) & (!x29x) & (!n_n4971) & (n_n4172) & (n_n1970)) + ((n_n4962) & (!x29x) & (n_n4971) & (!n_n4172) & (!n_n1970)) + ((n_n4962) & (!x29x) & (n_n4971) & (!n_n4172) & (n_n1970)) + ((n_n4962) & (!x29x) & (n_n4971) & (n_n4172) & (!n_n1970)) + ((n_n4962) & (!x29x) & (n_n4971) & (n_n4172) & (n_n1970)) + ((n_n4962) & (x29x) & (!n_n4971) & (!n_n4172) & (!n_n1970)) + ((n_n4962) & (x29x) & (!n_n4971) & (!n_n4172) & (n_n1970)) + ((n_n4962) & (x29x) & (!n_n4971) & (n_n4172) & (!n_n1970)) + ((n_n4962) & (x29x) & (!n_n4971) & (n_n4172) & (n_n1970)) + ((n_n4962) & (x29x) & (n_n4971) & (!n_n4172) & (!n_n1970)) + ((n_n4962) & (x29x) & (n_n4971) & (!n_n4172) & (n_n1970)) + ((n_n4962) & (x29x) & (n_n4971) & (n_n4172) & (!n_n1970)) + ((n_n4962) & (x29x) & (n_n4971) & (n_n4172) & (n_n1970)));
	assign x16180x = (((!n_n1850) & (!x16177x) & (x16178x)) + ((!n_n1850) & (x16177x) & (!x16178x)) + ((!n_n1850) & (x16177x) & (x16178x)) + ((n_n1850) & (!x16177x) & (!x16178x)) + ((n_n1850) & (!x16177x) & (x16178x)) + ((n_n1850) & (x16177x) & (!x16178x)) + ((n_n1850) & (x16177x) & (x16178x)));
	assign x16156x = (((!n_n4983) & (!x252x) & (!x393x) & (!n_n4984) & (x228x)) + ((!n_n4983) & (!x252x) & (!x393x) & (n_n4984) & (!x228x)) + ((!n_n4983) & (!x252x) & (!x393x) & (n_n4984) & (x228x)) + ((!n_n4983) & (!x252x) & (x393x) & (!n_n4984) & (!x228x)) + ((!n_n4983) & (!x252x) & (x393x) & (!n_n4984) & (x228x)) + ((!n_n4983) & (!x252x) & (x393x) & (n_n4984) & (!x228x)) + ((!n_n4983) & (!x252x) & (x393x) & (n_n4984) & (x228x)) + ((!n_n4983) & (x252x) & (!x393x) & (!n_n4984) & (!x228x)) + ((!n_n4983) & (x252x) & (!x393x) & (!n_n4984) & (x228x)) + ((!n_n4983) & (x252x) & (!x393x) & (n_n4984) & (!x228x)) + ((!n_n4983) & (x252x) & (!x393x) & (n_n4984) & (x228x)) + ((!n_n4983) & (x252x) & (x393x) & (!n_n4984) & (!x228x)) + ((!n_n4983) & (x252x) & (x393x) & (!n_n4984) & (x228x)) + ((!n_n4983) & (x252x) & (x393x) & (n_n4984) & (!x228x)) + ((!n_n4983) & (x252x) & (x393x) & (n_n4984) & (x228x)) + ((n_n4983) & (!x252x) & (!x393x) & (!n_n4984) & (!x228x)) + ((n_n4983) & (!x252x) & (!x393x) & (!n_n4984) & (x228x)) + ((n_n4983) & (!x252x) & (!x393x) & (n_n4984) & (!x228x)) + ((n_n4983) & (!x252x) & (!x393x) & (n_n4984) & (x228x)) + ((n_n4983) & (!x252x) & (x393x) & (!n_n4984) & (!x228x)) + ((n_n4983) & (!x252x) & (x393x) & (!n_n4984) & (x228x)) + ((n_n4983) & (!x252x) & (x393x) & (n_n4984) & (!x228x)) + ((n_n4983) & (!x252x) & (x393x) & (n_n4984) & (x228x)) + ((n_n4983) & (x252x) & (!x393x) & (!n_n4984) & (!x228x)) + ((n_n4983) & (x252x) & (!x393x) & (!n_n4984) & (x228x)) + ((n_n4983) & (x252x) & (!x393x) & (n_n4984) & (!x228x)) + ((n_n4983) & (x252x) & (!x393x) & (n_n4984) & (x228x)) + ((n_n4983) & (x252x) & (x393x) & (!n_n4984) & (!x228x)) + ((n_n4983) & (x252x) & (x393x) & (!n_n4984) & (x228x)) + ((n_n4983) & (x252x) & (x393x) & (n_n4984) & (!x228x)) + ((n_n4983) & (x252x) & (x393x) & (n_n4984) & (x228x)));
	assign x15845x = (((!x592x) & (!x11x) & (!x24x) & (!n_n5302) & (n_n5254)) + ((!x592x) & (!x11x) & (!x24x) & (n_n5302) & (!n_n5254)) + ((!x592x) & (!x11x) & (!x24x) & (n_n5302) & (n_n5254)) + ((!x592x) & (!x11x) & (x24x) & (!n_n5302) & (n_n5254)) + ((!x592x) & (!x11x) & (x24x) & (n_n5302) & (!n_n5254)) + ((!x592x) & (!x11x) & (x24x) & (n_n5302) & (n_n5254)) + ((!x592x) & (x11x) & (!x24x) & (!n_n5302) & (n_n5254)) + ((!x592x) & (x11x) & (!x24x) & (n_n5302) & (!n_n5254)) + ((!x592x) & (x11x) & (!x24x) & (n_n5302) & (n_n5254)) + ((!x592x) & (x11x) & (x24x) & (!n_n5302) & (n_n5254)) + ((!x592x) & (x11x) & (x24x) & (n_n5302) & (!n_n5254)) + ((!x592x) & (x11x) & (x24x) & (n_n5302) & (n_n5254)) + ((x592x) & (!x11x) & (!x24x) & (!n_n5302) & (n_n5254)) + ((x592x) & (!x11x) & (!x24x) & (n_n5302) & (!n_n5254)) + ((x592x) & (!x11x) & (!x24x) & (n_n5302) & (n_n5254)) + ((x592x) & (!x11x) & (x24x) & (!n_n5302) & (!n_n5254)) + ((x592x) & (!x11x) & (x24x) & (!n_n5302) & (n_n5254)) + ((x592x) & (!x11x) & (x24x) & (n_n5302) & (!n_n5254)) + ((x592x) & (!x11x) & (x24x) & (n_n5302) & (n_n5254)) + ((x592x) & (x11x) & (!x24x) & (!n_n5302) & (!n_n5254)) + ((x592x) & (x11x) & (!x24x) & (!n_n5302) & (n_n5254)) + ((x592x) & (x11x) & (!x24x) & (n_n5302) & (!n_n5254)) + ((x592x) & (x11x) & (!x24x) & (n_n5302) & (n_n5254)) + ((x592x) & (x11x) & (x24x) & (!n_n5302) & (!n_n5254)) + ((x592x) & (x11x) & (x24x) & (!n_n5302) & (n_n5254)) + ((x592x) & (x11x) & (x24x) & (n_n5302) & (!n_n5254)) + ((x592x) & (x11x) & (x24x) & (n_n5302) & (n_n5254)));
	assign x15846x = (((!n_n5238) & (!n_n5245) & (!n_n5253) & (!n_n5257) & (n_n5280)) + ((!n_n5238) & (!n_n5245) & (!n_n5253) & (n_n5257) & (!n_n5280)) + ((!n_n5238) & (!n_n5245) & (!n_n5253) & (n_n5257) & (n_n5280)) + ((!n_n5238) & (!n_n5245) & (n_n5253) & (!n_n5257) & (!n_n5280)) + ((!n_n5238) & (!n_n5245) & (n_n5253) & (!n_n5257) & (n_n5280)) + ((!n_n5238) & (!n_n5245) & (n_n5253) & (n_n5257) & (!n_n5280)) + ((!n_n5238) & (!n_n5245) & (n_n5253) & (n_n5257) & (n_n5280)) + ((!n_n5238) & (n_n5245) & (!n_n5253) & (!n_n5257) & (!n_n5280)) + ((!n_n5238) & (n_n5245) & (!n_n5253) & (!n_n5257) & (n_n5280)) + ((!n_n5238) & (n_n5245) & (!n_n5253) & (n_n5257) & (!n_n5280)) + ((!n_n5238) & (n_n5245) & (!n_n5253) & (n_n5257) & (n_n5280)) + ((!n_n5238) & (n_n5245) & (n_n5253) & (!n_n5257) & (!n_n5280)) + ((!n_n5238) & (n_n5245) & (n_n5253) & (!n_n5257) & (n_n5280)) + ((!n_n5238) & (n_n5245) & (n_n5253) & (n_n5257) & (!n_n5280)) + ((!n_n5238) & (n_n5245) & (n_n5253) & (n_n5257) & (n_n5280)) + ((n_n5238) & (!n_n5245) & (!n_n5253) & (!n_n5257) & (!n_n5280)) + ((n_n5238) & (!n_n5245) & (!n_n5253) & (!n_n5257) & (n_n5280)) + ((n_n5238) & (!n_n5245) & (!n_n5253) & (n_n5257) & (!n_n5280)) + ((n_n5238) & (!n_n5245) & (!n_n5253) & (n_n5257) & (n_n5280)) + ((n_n5238) & (!n_n5245) & (n_n5253) & (!n_n5257) & (!n_n5280)) + ((n_n5238) & (!n_n5245) & (n_n5253) & (!n_n5257) & (n_n5280)) + ((n_n5238) & (!n_n5245) & (n_n5253) & (n_n5257) & (!n_n5280)) + ((n_n5238) & (!n_n5245) & (n_n5253) & (n_n5257) & (n_n5280)) + ((n_n5238) & (n_n5245) & (!n_n5253) & (!n_n5257) & (!n_n5280)) + ((n_n5238) & (n_n5245) & (!n_n5253) & (!n_n5257) & (n_n5280)) + ((n_n5238) & (n_n5245) & (!n_n5253) & (n_n5257) & (!n_n5280)) + ((n_n5238) & (n_n5245) & (!n_n5253) & (n_n5257) & (n_n5280)) + ((n_n5238) & (n_n5245) & (n_n5253) & (!n_n5257) & (!n_n5280)) + ((n_n5238) & (n_n5245) & (n_n5253) & (!n_n5257) & (n_n5280)) + ((n_n5238) & (n_n5245) & (n_n5253) & (n_n5257) & (!n_n5280)) + ((n_n5238) & (n_n5245) & (n_n5253) & (n_n5257) & (n_n5280)));
	assign x11698x = (((!n_n5222) & (!n_n5214) & (!n_n5254) & (n_n5218)) + ((!n_n5222) & (!n_n5214) & (n_n5254) & (!n_n5218)) + ((!n_n5222) & (!n_n5214) & (n_n5254) & (n_n5218)) + ((!n_n5222) & (n_n5214) & (!n_n5254) & (!n_n5218)) + ((!n_n5222) & (n_n5214) & (!n_n5254) & (n_n5218)) + ((!n_n5222) & (n_n5214) & (n_n5254) & (!n_n5218)) + ((!n_n5222) & (n_n5214) & (n_n5254) & (n_n5218)) + ((n_n5222) & (!n_n5214) & (!n_n5254) & (!n_n5218)) + ((n_n5222) & (!n_n5214) & (!n_n5254) & (n_n5218)) + ((n_n5222) & (!n_n5214) & (n_n5254) & (!n_n5218)) + ((n_n5222) & (!n_n5214) & (n_n5254) & (n_n5218)) + ((n_n5222) & (n_n5214) & (!n_n5254) & (!n_n5218)) + ((n_n5222) & (n_n5214) & (!n_n5254) & (n_n5218)) + ((n_n5222) & (n_n5214) & (n_n5254) & (!n_n5218)) + ((n_n5222) & (n_n5214) & (n_n5254) & (n_n5218)));
	assign x11699x = (((!n_n5232) & (!n_n5216) & (!n_n5227) & (!n_n5213) & (n_n5248)) + ((!n_n5232) & (!n_n5216) & (!n_n5227) & (n_n5213) & (!n_n5248)) + ((!n_n5232) & (!n_n5216) & (!n_n5227) & (n_n5213) & (n_n5248)) + ((!n_n5232) & (!n_n5216) & (n_n5227) & (!n_n5213) & (!n_n5248)) + ((!n_n5232) & (!n_n5216) & (n_n5227) & (!n_n5213) & (n_n5248)) + ((!n_n5232) & (!n_n5216) & (n_n5227) & (n_n5213) & (!n_n5248)) + ((!n_n5232) & (!n_n5216) & (n_n5227) & (n_n5213) & (n_n5248)) + ((!n_n5232) & (n_n5216) & (!n_n5227) & (!n_n5213) & (!n_n5248)) + ((!n_n5232) & (n_n5216) & (!n_n5227) & (!n_n5213) & (n_n5248)) + ((!n_n5232) & (n_n5216) & (!n_n5227) & (n_n5213) & (!n_n5248)) + ((!n_n5232) & (n_n5216) & (!n_n5227) & (n_n5213) & (n_n5248)) + ((!n_n5232) & (n_n5216) & (n_n5227) & (!n_n5213) & (!n_n5248)) + ((!n_n5232) & (n_n5216) & (n_n5227) & (!n_n5213) & (n_n5248)) + ((!n_n5232) & (n_n5216) & (n_n5227) & (n_n5213) & (!n_n5248)) + ((!n_n5232) & (n_n5216) & (n_n5227) & (n_n5213) & (n_n5248)) + ((n_n5232) & (!n_n5216) & (!n_n5227) & (!n_n5213) & (!n_n5248)) + ((n_n5232) & (!n_n5216) & (!n_n5227) & (!n_n5213) & (n_n5248)) + ((n_n5232) & (!n_n5216) & (!n_n5227) & (n_n5213) & (!n_n5248)) + ((n_n5232) & (!n_n5216) & (!n_n5227) & (n_n5213) & (n_n5248)) + ((n_n5232) & (!n_n5216) & (n_n5227) & (!n_n5213) & (!n_n5248)) + ((n_n5232) & (!n_n5216) & (n_n5227) & (!n_n5213) & (n_n5248)) + ((n_n5232) & (!n_n5216) & (n_n5227) & (n_n5213) & (!n_n5248)) + ((n_n5232) & (!n_n5216) & (n_n5227) & (n_n5213) & (n_n5248)) + ((n_n5232) & (n_n5216) & (!n_n5227) & (!n_n5213) & (!n_n5248)) + ((n_n5232) & (n_n5216) & (!n_n5227) & (!n_n5213) & (n_n5248)) + ((n_n5232) & (n_n5216) & (!n_n5227) & (n_n5213) & (!n_n5248)) + ((n_n5232) & (n_n5216) & (!n_n5227) & (n_n5213) & (n_n5248)) + ((n_n5232) & (n_n5216) & (n_n5227) & (!n_n5213) & (!n_n5248)) + ((n_n5232) & (n_n5216) & (n_n5227) & (!n_n5213) & (n_n5248)) + ((n_n5232) & (n_n5216) & (n_n5227) & (n_n5213) & (!n_n5248)) + ((n_n5232) & (n_n5216) & (n_n5227) & (n_n5213) & (n_n5248)));
	assign x22212x = (((!n_n4416) & (!n_n4415) & (!n_n4413) & (!n_n4412) & (!x79x)));
	assign n_n730 = (((!n_n4420) & (!n_n4410) & (!n_n4414) & (!x22212x)) + ((!n_n4420) & (!n_n4410) & (n_n4414) & (!x22212x)) + ((!n_n4420) & (!n_n4410) & (n_n4414) & (x22212x)) + ((!n_n4420) & (n_n4410) & (!n_n4414) & (!x22212x)) + ((!n_n4420) & (n_n4410) & (!n_n4414) & (x22212x)) + ((!n_n4420) & (n_n4410) & (n_n4414) & (!x22212x)) + ((!n_n4420) & (n_n4410) & (n_n4414) & (x22212x)) + ((n_n4420) & (!n_n4410) & (!n_n4414) & (!x22212x)) + ((n_n4420) & (!n_n4410) & (!n_n4414) & (x22212x)) + ((n_n4420) & (!n_n4410) & (n_n4414) & (!x22212x)) + ((n_n4420) & (!n_n4410) & (n_n4414) & (x22212x)) + ((n_n4420) & (n_n4410) & (!n_n4414) & (!x22212x)) + ((n_n4420) & (n_n4410) & (!n_n4414) & (x22212x)) + ((n_n4420) & (n_n4410) & (n_n4414) & (!x22212x)) + ((n_n4420) & (n_n4410) & (n_n4414) & (x22212x)));
	assign x22131x = (((!n_n4991) & (!n_n4995) & (!n_n4993) & (!n_n4994)));
	assign x12834x = (((!x25x) & (!x24x) & (!n_n535) & (!n_n195) & (n_n814)) + ((!x25x) & (!x24x) & (!n_n535) & (n_n195) & (n_n814)) + ((!x25x) & (!x24x) & (n_n535) & (!n_n195) & (n_n814)) + ((!x25x) & (!x24x) & (n_n535) & (n_n195) & (n_n814)) + ((!x25x) & (x24x) & (!n_n535) & (!n_n195) & (n_n814)) + ((!x25x) & (x24x) & (!n_n535) & (n_n195) & (n_n814)) + ((!x25x) & (x24x) & (n_n535) & (!n_n195) & (n_n814)) + ((!x25x) & (x24x) & (n_n535) & (n_n195) & (!n_n814)) + ((!x25x) & (x24x) & (n_n535) & (n_n195) & (n_n814)) + ((x25x) & (!x24x) & (!n_n535) & (!n_n195) & (n_n814)) + ((x25x) & (!x24x) & (!n_n535) & (n_n195) & (n_n814)) + ((x25x) & (!x24x) & (n_n535) & (!n_n195) & (n_n814)) + ((x25x) & (!x24x) & (n_n535) & (n_n195) & (!n_n814)) + ((x25x) & (!x24x) & (n_n535) & (n_n195) & (n_n814)) + ((x25x) & (x24x) & (!n_n535) & (!n_n195) & (n_n814)) + ((x25x) & (x24x) & (!n_n535) & (n_n195) & (n_n814)) + ((x25x) & (x24x) & (n_n535) & (!n_n195) & (n_n814)) + ((x25x) & (x24x) & (n_n535) & (n_n195) & (!n_n814)) + ((x25x) & (x24x) & (n_n535) & (n_n195) & (n_n814)));
	assign n_n662 = (((!n_n5307) & (!x462x) & (!n_n5308) & (n_n5309)) + ((!n_n5307) & (!x462x) & (n_n5308) & (!n_n5309)) + ((!n_n5307) & (!x462x) & (n_n5308) & (n_n5309)) + ((!n_n5307) & (x462x) & (!n_n5308) & (!n_n5309)) + ((!n_n5307) & (x462x) & (!n_n5308) & (n_n5309)) + ((!n_n5307) & (x462x) & (n_n5308) & (!n_n5309)) + ((!n_n5307) & (x462x) & (n_n5308) & (n_n5309)) + ((n_n5307) & (!x462x) & (!n_n5308) & (!n_n5309)) + ((n_n5307) & (!x462x) & (!n_n5308) & (n_n5309)) + ((n_n5307) & (!x462x) & (n_n5308) & (!n_n5309)) + ((n_n5307) & (!x462x) & (n_n5308) & (n_n5309)) + ((n_n5307) & (x462x) & (!n_n5308) & (!n_n5309)) + ((n_n5307) & (x462x) & (!n_n5308) & (n_n5309)) + ((n_n5307) & (x462x) & (n_n5308) & (!n_n5309)) + ((n_n5307) & (x462x) & (n_n5308) & (n_n5309)));
	assign x12975x = (((!n_n5318) & (!n_n5320) & (!n_n5319) & (!n_n5313) & (n_n5315)) + ((!n_n5318) & (!n_n5320) & (!n_n5319) & (n_n5313) & (!n_n5315)) + ((!n_n5318) & (!n_n5320) & (!n_n5319) & (n_n5313) & (n_n5315)) + ((!n_n5318) & (!n_n5320) & (n_n5319) & (!n_n5313) & (!n_n5315)) + ((!n_n5318) & (!n_n5320) & (n_n5319) & (!n_n5313) & (n_n5315)) + ((!n_n5318) & (!n_n5320) & (n_n5319) & (n_n5313) & (!n_n5315)) + ((!n_n5318) & (!n_n5320) & (n_n5319) & (n_n5313) & (n_n5315)) + ((!n_n5318) & (n_n5320) & (!n_n5319) & (!n_n5313) & (!n_n5315)) + ((!n_n5318) & (n_n5320) & (!n_n5319) & (!n_n5313) & (n_n5315)) + ((!n_n5318) & (n_n5320) & (!n_n5319) & (n_n5313) & (!n_n5315)) + ((!n_n5318) & (n_n5320) & (!n_n5319) & (n_n5313) & (n_n5315)) + ((!n_n5318) & (n_n5320) & (n_n5319) & (!n_n5313) & (!n_n5315)) + ((!n_n5318) & (n_n5320) & (n_n5319) & (!n_n5313) & (n_n5315)) + ((!n_n5318) & (n_n5320) & (n_n5319) & (n_n5313) & (!n_n5315)) + ((!n_n5318) & (n_n5320) & (n_n5319) & (n_n5313) & (n_n5315)) + ((n_n5318) & (!n_n5320) & (!n_n5319) & (!n_n5313) & (!n_n5315)) + ((n_n5318) & (!n_n5320) & (!n_n5319) & (!n_n5313) & (n_n5315)) + ((n_n5318) & (!n_n5320) & (!n_n5319) & (n_n5313) & (!n_n5315)) + ((n_n5318) & (!n_n5320) & (!n_n5319) & (n_n5313) & (n_n5315)) + ((n_n5318) & (!n_n5320) & (n_n5319) & (!n_n5313) & (!n_n5315)) + ((n_n5318) & (!n_n5320) & (n_n5319) & (!n_n5313) & (n_n5315)) + ((n_n5318) & (!n_n5320) & (n_n5319) & (n_n5313) & (!n_n5315)) + ((n_n5318) & (!n_n5320) & (n_n5319) & (n_n5313) & (n_n5315)) + ((n_n5318) & (n_n5320) & (!n_n5319) & (!n_n5313) & (!n_n5315)) + ((n_n5318) & (n_n5320) & (!n_n5319) & (!n_n5313) & (n_n5315)) + ((n_n5318) & (n_n5320) & (!n_n5319) & (n_n5313) & (!n_n5315)) + ((n_n5318) & (n_n5320) & (!n_n5319) & (n_n5313) & (n_n5315)) + ((n_n5318) & (n_n5320) & (n_n5319) & (!n_n5313) & (!n_n5315)) + ((n_n5318) & (n_n5320) & (n_n5319) & (!n_n5313) & (n_n5315)) + ((n_n5318) & (n_n5320) & (n_n5319) & (n_n5313) & (!n_n5315)) + ((n_n5318) & (n_n5320) & (n_n5319) & (n_n5313) & (n_n5315)));
	assign n_n661 = (((!n_n5310) & (!n_n5316) & (!n_n5312) & (!n_n5311) & (x12975x)) + ((!n_n5310) & (!n_n5316) & (!n_n5312) & (n_n5311) & (!x12975x)) + ((!n_n5310) & (!n_n5316) & (!n_n5312) & (n_n5311) & (x12975x)) + ((!n_n5310) & (!n_n5316) & (n_n5312) & (!n_n5311) & (!x12975x)) + ((!n_n5310) & (!n_n5316) & (n_n5312) & (!n_n5311) & (x12975x)) + ((!n_n5310) & (!n_n5316) & (n_n5312) & (n_n5311) & (!x12975x)) + ((!n_n5310) & (!n_n5316) & (n_n5312) & (n_n5311) & (x12975x)) + ((!n_n5310) & (n_n5316) & (!n_n5312) & (!n_n5311) & (!x12975x)) + ((!n_n5310) & (n_n5316) & (!n_n5312) & (!n_n5311) & (x12975x)) + ((!n_n5310) & (n_n5316) & (!n_n5312) & (n_n5311) & (!x12975x)) + ((!n_n5310) & (n_n5316) & (!n_n5312) & (n_n5311) & (x12975x)) + ((!n_n5310) & (n_n5316) & (n_n5312) & (!n_n5311) & (!x12975x)) + ((!n_n5310) & (n_n5316) & (n_n5312) & (!n_n5311) & (x12975x)) + ((!n_n5310) & (n_n5316) & (n_n5312) & (n_n5311) & (!x12975x)) + ((!n_n5310) & (n_n5316) & (n_n5312) & (n_n5311) & (x12975x)) + ((n_n5310) & (!n_n5316) & (!n_n5312) & (!n_n5311) & (!x12975x)) + ((n_n5310) & (!n_n5316) & (!n_n5312) & (!n_n5311) & (x12975x)) + ((n_n5310) & (!n_n5316) & (!n_n5312) & (n_n5311) & (!x12975x)) + ((n_n5310) & (!n_n5316) & (!n_n5312) & (n_n5311) & (x12975x)) + ((n_n5310) & (!n_n5316) & (n_n5312) & (!n_n5311) & (!x12975x)) + ((n_n5310) & (!n_n5316) & (n_n5312) & (!n_n5311) & (x12975x)) + ((n_n5310) & (!n_n5316) & (n_n5312) & (n_n5311) & (!x12975x)) + ((n_n5310) & (!n_n5316) & (n_n5312) & (n_n5311) & (x12975x)) + ((n_n5310) & (n_n5316) & (!n_n5312) & (!n_n5311) & (!x12975x)) + ((n_n5310) & (n_n5316) & (!n_n5312) & (!n_n5311) & (x12975x)) + ((n_n5310) & (n_n5316) & (!n_n5312) & (n_n5311) & (!x12975x)) + ((n_n5310) & (n_n5316) & (!n_n5312) & (n_n5311) & (x12975x)) + ((n_n5310) & (n_n5316) & (n_n5312) & (!n_n5311) & (!x12975x)) + ((n_n5310) & (n_n5316) & (n_n5312) & (!n_n5311) & (x12975x)) + ((n_n5310) & (n_n5316) & (n_n5312) & (n_n5311) & (!x12975x)) + ((n_n5310) & (n_n5316) & (n_n5312) & (n_n5311) & (x12975x)));
	assign x12981x = (((!x592x) & (!x21x) & (!x11x) & (!x207x) & (x12980x)) + ((!x592x) & (!x21x) & (!x11x) & (x207x) & (!x12980x)) + ((!x592x) & (!x21x) & (!x11x) & (x207x) & (x12980x)) + ((!x592x) & (!x21x) & (x11x) & (!x207x) & (x12980x)) + ((!x592x) & (!x21x) & (x11x) & (x207x) & (!x12980x)) + ((!x592x) & (!x21x) & (x11x) & (x207x) & (x12980x)) + ((!x592x) & (x21x) & (!x11x) & (!x207x) & (x12980x)) + ((!x592x) & (x21x) & (!x11x) & (x207x) & (!x12980x)) + ((!x592x) & (x21x) & (!x11x) & (x207x) & (x12980x)) + ((!x592x) & (x21x) & (x11x) & (!x207x) & (x12980x)) + ((!x592x) & (x21x) & (x11x) & (x207x) & (!x12980x)) + ((!x592x) & (x21x) & (x11x) & (x207x) & (x12980x)) + ((x592x) & (!x21x) & (!x11x) & (!x207x) & (x12980x)) + ((x592x) & (!x21x) & (!x11x) & (x207x) & (!x12980x)) + ((x592x) & (!x21x) & (!x11x) & (x207x) & (x12980x)) + ((x592x) & (!x21x) & (x11x) & (!x207x) & (!x12980x)) + ((x592x) & (!x21x) & (x11x) & (!x207x) & (x12980x)) + ((x592x) & (!x21x) & (x11x) & (x207x) & (!x12980x)) + ((x592x) & (!x21x) & (x11x) & (x207x) & (x12980x)) + ((x592x) & (x21x) & (!x11x) & (!x207x) & (!x12980x)) + ((x592x) & (x21x) & (!x11x) & (!x207x) & (x12980x)) + ((x592x) & (x21x) & (!x11x) & (x207x) & (!x12980x)) + ((x592x) & (x21x) & (!x11x) & (x207x) & (x12980x)) + ((x592x) & (x21x) & (x11x) & (!x207x) & (!x12980x)) + ((x592x) & (x21x) & (x11x) & (!x207x) & (x12980x)) + ((x592x) & (x21x) & (x11x) & (x207x) & (!x12980x)) + ((x592x) & (x21x) & (x11x) & (x207x) & (x12980x)));
	assign x12984x = (((!n_n632) & (!n_n662) & (!n_n661) & (x12981x)) + ((!n_n632) & (!n_n662) & (n_n661) & (!x12981x)) + ((!n_n632) & (!n_n662) & (n_n661) & (x12981x)) + ((!n_n632) & (n_n662) & (!n_n661) & (!x12981x)) + ((!n_n632) & (n_n662) & (!n_n661) & (x12981x)) + ((!n_n632) & (n_n662) & (n_n661) & (!x12981x)) + ((!n_n632) & (n_n662) & (n_n661) & (x12981x)) + ((n_n632) & (!n_n662) & (!n_n661) & (!x12981x)) + ((n_n632) & (!n_n662) & (!n_n661) & (x12981x)) + ((n_n632) & (!n_n662) & (n_n661) & (!x12981x)) + ((n_n632) & (!n_n662) & (n_n661) & (x12981x)) + ((n_n632) & (n_n662) & (!n_n661) & (!x12981x)) + ((n_n632) & (n_n662) & (!n_n661) & (x12981x)) + ((n_n632) & (n_n662) & (n_n661) & (!x12981x)) + ((n_n632) & (n_n662) & (n_n661) & (x12981x)));
	assign x12989x = (((!n_n5203) & (!n_n5205) & (!n_n5197) & (x36x)) + ((!n_n5203) & (!n_n5205) & (n_n5197) & (!x36x)) + ((!n_n5203) & (!n_n5205) & (n_n5197) & (x36x)) + ((!n_n5203) & (n_n5205) & (!n_n5197) & (!x36x)) + ((!n_n5203) & (n_n5205) & (!n_n5197) & (x36x)) + ((!n_n5203) & (n_n5205) & (n_n5197) & (!x36x)) + ((!n_n5203) & (n_n5205) & (n_n5197) & (x36x)) + ((n_n5203) & (!n_n5205) & (!n_n5197) & (!x36x)) + ((n_n5203) & (!n_n5205) & (!n_n5197) & (x36x)) + ((n_n5203) & (!n_n5205) & (n_n5197) & (!x36x)) + ((n_n5203) & (!n_n5205) & (n_n5197) & (x36x)) + ((n_n5203) & (n_n5205) & (!n_n5197) & (!x36x)) + ((n_n5203) & (n_n5205) & (!n_n5197) & (x36x)) + ((n_n5203) & (n_n5205) & (n_n5197) & (!x36x)) + ((n_n5203) & (n_n5205) & (n_n5197) & (x36x)));
	assign n_n670 = (((!n_n5207) & (!n_n5199) & (!x452x) & (x12989x)) + ((!n_n5207) & (!n_n5199) & (x452x) & (!x12989x)) + ((!n_n5207) & (!n_n5199) & (x452x) & (x12989x)) + ((!n_n5207) & (n_n5199) & (!x452x) & (!x12989x)) + ((!n_n5207) & (n_n5199) & (!x452x) & (x12989x)) + ((!n_n5207) & (n_n5199) & (x452x) & (!x12989x)) + ((!n_n5207) & (n_n5199) & (x452x) & (x12989x)) + ((n_n5207) & (!n_n5199) & (!x452x) & (!x12989x)) + ((n_n5207) & (!n_n5199) & (!x452x) & (x12989x)) + ((n_n5207) & (!n_n5199) & (x452x) & (!x12989x)) + ((n_n5207) & (!n_n5199) & (x452x) & (x12989x)) + ((n_n5207) & (n_n5199) & (!x452x) & (!x12989x)) + ((n_n5207) & (n_n5199) & (!x452x) & (x12989x)) + ((n_n5207) & (n_n5199) & (x452x) & (!x12989x)) + ((n_n5207) & (n_n5199) & (x452x) & (x12989x)));
	assign n_n671 = (((!x112x) & (!n_n5188) & (!n_n5192) & (!n_n1927) & (x188x)) + ((!x112x) & (!n_n5188) & (!n_n5192) & (n_n1927) & (!x188x)) + ((!x112x) & (!n_n5188) & (!n_n5192) & (n_n1927) & (x188x)) + ((!x112x) & (!n_n5188) & (n_n5192) & (!n_n1927) & (!x188x)) + ((!x112x) & (!n_n5188) & (n_n5192) & (!n_n1927) & (x188x)) + ((!x112x) & (!n_n5188) & (n_n5192) & (n_n1927) & (!x188x)) + ((!x112x) & (!n_n5188) & (n_n5192) & (n_n1927) & (x188x)) + ((!x112x) & (n_n5188) & (!n_n5192) & (!n_n1927) & (!x188x)) + ((!x112x) & (n_n5188) & (!n_n5192) & (!n_n1927) & (x188x)) + ((!x112x) & (n_n5188) & (!n_n5192) & (n_n1927) & (!x188x)) + ((!x112x) & (n_n5188) & (!n_n5192) & (n_n1927) & (x188x)) + ((!x112x) & (n_n5188) & (n_n5192) & (!n_n1927) & (!x188x)) + ((!x112x) & (n_n5188) & (n_n5192) & (!n_n1927) & (x188x)) + ((!x112x) & (n_n5188) & (n_n5192) & (n_n1927) & (!x188x)) + ((!x112x) & (n_n5188) & (n_n5192) & (n_n1927) & (x188x)) + ((x112x) & (!n_n5188) & (!n_n5192) & (!n_n1927) & (!x188x)) + ((x112x) & (!n_n5188) & (!n_n5192) & (!n_n1927) & (x188x)) + ((x112x) & (!n_n5188) & (!n_n5192) & (n_n1927) & (!x188x)) + ((x112x) & (!n_n5188) & (!n_n5192) & (n_n1927) & (x188x)) + ((x112x) & (!n_n5188) & (n_n5192) & (!n_n1927) & (!x188x)) + ((x112x) & (!n_n5188) & (n_n5192) & (!n_n1927) & (x188x)) + ((x112x) & (!n_n5188) & (n_n5192) & (n_n1927) & (!x188x)) + ((x112x) & (!n_n5188) & (n_n5192) & (n_n1927) & (x188x)) + ((x112x) & (n_n5188) & (!n_n5192) & (!n_n1927) & (!x188x)) + ((x112x) & (n_n5188) & (!n_n5192) & (!n_n1927) & (x188x)) + ((x112x) & (n_n5188) & (!n_n5192) & (n_n1927) & (!x188x)) + ((x112x) & (n_n5188) & (!n_n5192) & (n_n1927) & (x188x)) + ((x112x) & (n_n5188) & (n_n5192) & (!n_n1927) & (!x188x)) + ((x112x) & (n_n5188) & (n_n5192) & (!n_n1927) & (x188x)) + ((x112x) & (n_n5188) & (n_n5192) & (n_n1927) & (!x188x)) + ((x112x) & (n_n5188) & (n_n5192) & (n_n1927) & (x188x)));
	assign x12999x = (((!n_n670) & (!n_n671) & (!x12995x) & (x12996x)) + ((!n_n670) & (!n_n671) & (x12995x) & (!x12996x)) + ((!n_n670) & (!n_n671) & (x12995x) & (x12996x)) + ((!n_n670) & (n_n671) & (!x12995x) & (!x12996x)) + ((!n_n670) & (n_n671) & (!x12995x) & (x12996x)) + ((!n_n670) & (n_n671) & (x12995x) & (!x12996x)) + ((!n_n670) & (n_n671) & (x12995x) & (x12996x)) + ((n_n670) & (!n_n671) & (!x12995x) & (!x12996x)) + ((n_n670) & (!n_n671) & (!x12995x) & (x12996x)) + ((n_n670) & (!n_n671) & (x12995x) & (!x12996x)) + ((n_n670) & (!n_n671) & (x12995x) & (x12996x)) + ((n_n670) & (n_n671) & (!x12995x) & (!x12996x)) + ((n_n670) & (n_n671) & (!x12995x) & (x12996x)) + ((n_n670) & (n_n671) & (x12995x) & (!x12996x)) + ((n_n670) & (n_n671) & (x12995x) & (x12996x)));
	assign x14472x = (((!n_n4372) & (!n_n4371) & (!n_n4366) & (!n_n4376) & (n_n4375)) + ((!n_n4372) & (!n_n4371) & (!n_n4366) & (n_n4376) & (!n_n4375)) + ((!n_n4372) & (!n_n4371) & (!n_n4366) & (n_n4376) & (n_n4375)) + ((!n_n4372) & (!n_n4371) & (n_n4366) & (!n_n4376) & (!n_n4375)) + ((!n_n4372) & (!n_n4371) & (n_n4366) & (!n_n4376) & (n_n4375)) + ((!n_n4372) & (!n_n4371) & (n_n4366) & (n_n4376) & (!n_n4375)) + ((!n_n4372) & (!n_n4371) & (n_n4366) & (n_n4376) & (n_n4375)) + ((!n_n4372) & (n_n4371) & (!n_n4366) & (!n_n4376) & (!n_n4375)) + ((!n_n4372) & (n_n4371) & (!n_n4366) & (!n_n4376) & (n_n4375)) + ((!n_n4372) & (n_n4371) & (!n_n4366) & (n_n4376) & (!n_n4375)) + ((!n_n4372) & (n_n4371) & (!n_n4366) & (n_n4376) & (n_n4375)) + ((!n_n4372) & (n_n4371) & (n_n4366) & (!n_n4376) & (!n_n4375)) + ((!n_n4372) & (n_n4371) & (n_n4366) & (!n_n4376) & (n_n4375)) + ((!n_n4372) & (n_n4371) & (n_n4366) & (n_n4376) & (!n_n4375)) + ((!n_n4372) & (n_n4371) & (n_n4366) & (n_n4376) & (n_n4375)) + ((n_n4372) & (!n_n4371) & (!n_n4366) & (!n_n4376) & (!n_n4375)) + ((n_n4372) & (!n_n4371) & (!n_n4366) & (!n_n4376) & (n_n4375)) + ((n_n4372) & (!n_n4371) & (!n_n4366) & (n_n4376) & (!n_n4375)) + ((n_n4372) & (!n_n4371) & (!n_n4366) & (n_n4376) & (n_n4375)) + ((n_n4372) & (!n_n4371) & (n_n4366) & (!n_n4376) & (!n_n4375)) + ((n_n4372) & (!n_n4371) & (n_n4366) & (!n_n4376) & (n_n4375)) + ((n_n4372) & (!n_n4371) & (n_n4366) & (n_n4376) & (!n_n4375)) + ((n_n4372) & (!n_n4371) & (n_n4366) & (n_n4376) & (n_n4375)) + ((n_n4372) & (n_n4371) & (!n_n4366) & (!n_n4376) & (!n_n4375)) + ((n_n4372) & (n_n4371) & (!n_n4366) & (!n_n4376) & (n_n4375)) + ((n_n4372) & (n_n4371) & (!n_n4366) & (n_n4376) & (!n_n4375)) + ((n_n4372) & (n_n4371) & (!n_n4366) & (n_n4376) & (n_n4375)) + ((n_n4372) & (n_n4371) & (n_n4366) & (!n_n4376) & (!n_n4375)) + ((n_n4372) & (n_n4371) & (n_n4366) & (!n_n4376) & (n_n4375)) + ((n_n4372) & (n_n4371) & (n_n4366) & (n_n4376) & (!n_n4375)) + ((n_n4372) & (n_n4371) & (n_n4366) & (n_n4376) & (n_n4375)));
	assign x15471x = (((!n_n4642) & (!n_n4644) & (!n_n4658) & (!x13454x) & (x432x)) + ((!n_n4642) & (!n_n4644) & (!n_n4658) & (x13454x) & (!x432x)) + ((!n_n4642) & (!n_n4644) & (!n_n4658) & (x13454x) & (x432x)) + ((!n_n4642) & (!n_n4644) & (n_n4658) & (!x13454x) & (!x432x)) + ((!n_n4642) & (!n_n4644) & (n_n4658) & (!x13454x) & (x432x)) + ((!n_n4642) & (!n_n4644) & (n_n4658) & (x13454x) & (!x432x)) + ((!n_n4642) & (!n_n4644) & (n_n4658) & (x13454x) & (x432x)) + ((!n_n4642) & (n_n4644) & (!n_n4658) & (!x13454x) & (!x432x)) + ((!n_n4642) & (n_n4644) & (!n_n4658) & (!x13454x) & (x432x)) + ((!n_n4642) & (n_n4644) & (!n_n4658) & (x13454x) & (!x432x)) + ((!n_n4642) & (n_n4644) & (!n_n4658) & (x13454x) & (x432x)) + ((!n_n4642) & (n_n4644) & (n_n4658) & (!x13454x) & (!x432x)) + ((!n_n4642) & (n_n4644) & (n_n4658) & (!x13454x) & (x432x)) + ((!n_n4642) & (n_n4644) & (n_n4658) & (x13454x) & (!x432x)) + ((!n_n4642) & (n_n4644) & (n_n4658) & (x13454x) & (x432x)) + ((n_n4642) & (!n_n4644) & (!n_n4658) & (!x13454x) & (!x432x)) + ((n_n4642) & (!n_n4644) & (!n_n4658) & (!x13454x) & (x432x)) + ((n_n4642) & (!n_n4644) & (!n_n4658) & (x13454x) & (!x432x)) + ((n_n4642) & (!n_n4644) & (!n_n4658) & (x13454x) & (x432x)) + ((n_n4642) & (!n_n4644) & (n_n4658) & (!x13454x) & (!x432x)) + ((n_n4642) & (!n_n4644) & (n_n4658) & (!x13454x) & (x432x)) + ((n_n4642) & (!n_n4644) & (n_n4658) & (x13454x) & (!x432x)) + ((n_n4642) & (!n_n4644) & (n_n4658) & (x13454x) & (x432x)) + ((n_n4642) & (n_n4644) & (!n_n4658) & (!x13454x) & (!x432x)) + ((n_n4642) & (n_n4644) & (!n_n4658) & (!x13454x) & (x432x)) + ((n_n4642) & (n_n4644) & (!n_n4658) & (x13454x) & (!x432x)) + ((n_n4642) & (n_n4644) & (!n_n4658) & (x13454x) & (x432x)) + ((n_n4642) & (n_n4644) & (n_n4658) & (!x13454x) & (!x432x)) + ((n_n4642) & (n_n4644) & (n_n4658) & (!x13454x) & (x432x)) + ((n_n4642) & (n_n4644) & (n_n4658) & (x13454x) & (!x432x)) + ((n_n4642) & (n_n4644) & (n_n4658) & (x13454x) & (x432x)));
	assign x15470x = (((!n_n4666) & (!n_n4648) & (!x309x) & (!x157x) & (x139x)) + ((!n_n4666) & (!n_n4648) & (!x309x) & (x157x) & (!x139x)) + ((!n_n4666) & (!n_n4648) & (!x309x) & (x157x) & (x139x)) + ((!n_n4666) & (!n_n4648) & (x309x) & (!x157x) & (!x139x)) + ((!n_n4666) & (!n_n4648) & (x309x) & (!x157x) & (x139x)) + ((!n_n4666) & (!n_n4648) & (x309x) & (x157x) & (!x139x)) + ((!n_n4666) & (!n_n4648) & (x309x) & (x157x) & (x139x)) + ((!n_n4666) & (n_n4648) & (!x309x) & (!x157x) & (!x139x)) + ((!n_n4666) & (n_n4648) & (!x309x) & (!x157x) & (x139x)) + ((!n_n4666) & (n_n4648) & (!x309x) & (x157x) & (!x139x)) + ((!n_n4666) & (n_n4648) & (!x309x) & (x157x) & (x139x)) + ((!n_n4666) & (n_n4648) & (x309x) & (!x157x) & (!x139x)) + ((!n_n4666) & (n_n4648) & (x309x) & (!x157x) & (x139x)) + ((!n_n4666) & (n_n4648) & (x309x) & (x157x) & (!x139x)) + ((!n_n4666) & (n_n4648) & (x309x) & (x157x) & (x139x)) + ((n_n4666) & (!n_n4648) & (!x309x) & (!x157x) & (!x139x)) + ((n_n4666) & (!n_n4648) & (!x309x) & (!x157x) & (x139x)) + ((n_n4666) & (!n_n4648) & (!x309x) & (x157x) & (!x139x)) + ((n_n4666) & (!n_n4648) & (!x309x) & (x157x) & (x139x)) + ((n_n4666) & (!n_n4648) & (x309x) & (!x157x) & (!x139x)) + ((n_n4666) & (!n_n4648) & (x309x) & (!x157x) & (x139x)) + ((n_n4666) & (!n_n4648) & (x309x) & (x157x) & (!x139x)) + ((n_n4666) & (!n_n4648) & (x309x) & (x157x) & (x139x)) + ((n_n4666) & (n_n4648) & (!x309x) & (!x157x) & (!x139x)) + ((n_n4666) & (n_n4648) & (!x309x) & (!x157x) & (x139x)) + ((n_n4666) & (n_n4648) & (!x309x) & (x157x) & (!x139x)) + ((n_n4666) & (n_n4648) & (!x309x) & (x157x) & (x139x)) + ((n_n4666) & (n_n4648) & (x309x) & (!x157x) & (!x139x)) + ((n_n4666) & (n_n4648) & (x309x) & (!x157x) & (x139x)) + ((n_n4666) & (n_n4648) & (x309x) & (x157x) & (!x139x)) + ((n_n4666) & (n_n4648) & (x309x) & (x157x) & (x139x)));
	assign x15348x = (((!n_n4898) & (!n_n4877) & (!n_n4876) & (n_n4899)) + ((!n_n4898) & (!n_n4877) & (n_n4876) & (!n_n4899)) + ((!n_n4898) & (!n_n4877) & (n_n4876) & (n_n4899)) + ((!n_n4898) & (n_n4877) & (!n_n4876) & (!n_n4899)) + ((!n_n4898) & (n_n4877) & (!n_n4876) & (n_n4899)) + ((!n_n4898) & (n_n4877) & (n_n4876) & (!n_n4899)) + ((!n_n4898) & (n_n4877) & (n_n4876) & (n_n4899)) + ((n_n4898) & (!n_n4877) & (!n_n4876) & (!n_n4899)) + ((n_n4898) & (!n_n4877) & (!n_n4876) & (n_n4899)) + ((n_n4898) & (!n_n4877) & (n_n4876) & (!n_n4899)) + ((n_n4898) & (!n_n4877) & (n_n4876) & (n_n4899)) + ((n_n4898) & (n_n4877) & (!n_n4876) & (!n_n4899)) + ((n_n4898) & (n_n4877) & (!n_n4876) & (n_n4899)) + ((n_n4898) & (n_n4877) & (n_n4876) & (!n_n4899)) + ((n_n4898) & (n_n4877) & (n_n4876) & (n_n4899)));
	assign x15349x = (((!n_n4886) & (!n_n4915) & (!x154x) & (n_n4874)) + ((!n_n4886) & (!n_n4915) & (x154x) & (!n_n4874)) + ((!n_n4886) & (!n_n4915) & (x154x) & (n_n4874)) + ((!n_n4886) & (n_n4915) & (!x154x) & (!n_n4874)) + ((!n_n4886) & (n_n4915) & (!x154x) & (n_n4874)) + ((!n_n4886) & (n_n4915) & (x154x) & (!n_n4874)) + ((!n_n4886) & (n_n4915) & (x154x) & (n_n4874)) + ((n_n4886) & (!n_n4915) & (!x154x) & (!n_n4874)) + ((n_n4886) & (!n_n4915) & (!x154x) & (n_n4874)) + ((n_n4886) & (!n_n4915) & (x154x) & (!n_n4874)) + ((n_n4886) & (!n_n4915) & (x154x) & (n_n4874)) + ((n_n4886) & (n_n4915) & (!x154x) & (!n_n4874)) + ((n_n4886) & (n_n4915) & (!x154x) & (n_n4874)) + ((n_n4886) & (n_n4915) & (x154x) & (!n_n4874)) + ((n_n4886) & (n_n4915) & (x154x) & (n_n4874)));
	assign x13056x = (((!i_9_) & (n_n536) & (!n_n526) & (n_n528) & (n_n500)) + ((!i_9_) & (n_n536) & (n_n526) & (!n_n528) & (n_n500)) + ((!i_9_) & (n_n536) & (n_n526) & (n_n528) & (n_n500)) + ((i_9_) & (n_n536) & (n_n526) & (!n_n528) & (n_n500)) + ((i_9_) & (n_n536) & (n_n526) & (n_n528) & (n_n500)));
	assign x16089x = (((!i_9_) & (n_n536) & (!n_n522) & (n_n520) & (n_n500)) + ((!i_9_) & (n_n536) & (n_n522) & (n_n520) & (n_n500)) + ((i_9_) & (n_n536) & (!n_n522) & (n_n520) & (n_n500)) + ((i_9_) & (n_n536) & (n_n522) & (!n_n520) & (n_n500)) + ((i_9_) & (n_n536) & (n_n522) & (n_n520) & (n_n500)));
	assign x16189x = (((!n_n4800) & (!n_n4806) & (!n_n4807) & (n_n4808)) + ((!n_n4800) & (!n_n4806) & (n_n4807) & (!n_n4808)) + ((!n_n4800) & (!n_n4806) & (n_n4807) & (n_n4808)) + ((!n_n4800) & (n_n4806) & (!n_n4807) & (!n_n4808)) + ((!n_n4800) & (n_n4806) & (!n_n4807) & (n_n4808)) + ((!n_n4800) & (n_n4806) & (n_n4807) & (!n_n4808)) + ((!n_n4800) & (n_n4806) & (n_n4807) & (n_n4808)) + ((n_n4800) & (!n_n4806) & (!n_n4807) & (!n_n4808)) + ((n_n4800) & (!n_n4806) & (!n_n4807) & (n_n4808)) + ((n_n4800) & (!n_n4806) & (n_n4807) & (!n_n4808)) + ((n_n4800) & (!n_n4806) & (n_n4807) & (n_n4808)) + ((n_n4800) & (n_n4806) & (!n_n4807) & (!n_n4808)) + ((n_n4800) & (n_n4806) & (!n_n4807) & (n_n4808)) + ((n_n4800) & (n_n4806) & (n_n4807) & (!n_n4808)) + ((n_n4800) & (n_n4806) & (n_n4807) & (n_n4808)));
	assign x16190x = (((!n_n4803) & (!n_n4804) & (!n_n4802) & (!n_n4805) & (n_n4799)) + ((!n_n4803) & (!n_n4804) & (!n_n4802) & (n_n4805) & (!n_n4799)) + ((!n_n4803) & (!n_n4804) & (!n_n4802) & (n_n4805) & (n_n4799)) + ((!n_n4803) & (!n_n4804) & (n_n4802) & (!n_n4805) & (!n_n4799)) + ((!n_n4803) & (!n_n4804) & (n_n4802) & (!n_n4805) & (n_n4799)) + ((!n_n4803) & (!n_n4804) & (n_n4802) & (n_n4805) & (!n_n4799)) + ((!n_n4803) & (!n_n4804) & (n_n4802) & (n_n4805) & (n_n4799)) + ((!n_n4803) & (n_n4804) & (!n_n4802) & (!n_n4805) & (!n_n4799)) + ((!n_n4803) & (n_n4804) & (!n_n4802) & (!n_n4805) & (n_n4799)) + ((!n_n4803) & (n_n4804) & (!n_n4802) & (n_n4805) & (!n_n4799)) + ((!n_n4803) & (n_n4804) & (!n_n4802) & (n_n4805) & (n_n4799)) + ((!n_n4803) & (n_n4804) & (n_n4802) & (!n_n4805) & (!n_n4799)) + ((!n_n4803) & (n_n4804) & (n_n4802) & (!n_n4805) & (n_n4799)) + ((!n_n4803) & (n_n4804) & (n_n4802) & (n_n4805) & (!n_n4799)) + ((!n_n4803) & (n_n4804) & (n_n4802) & (n_n4805) & (n_n4799)) + ((n_n4803) & (!n_n4804) & (!n_n4802) & (!n_n4805) & (!n_n4799)) + ((n_n4803) & (!n_n4804) & (!n_n4802) & (!n_n4805) & (n_n4799)) + ((n_n4803) & (!n_n4804) & (!n_n4802) & (n_n4805) & (!n_n4799)) + ((n_n4803) & (!n_n4804) & (!n_n4802) & (n_n4805) & (n_n4799)) + ((n_n4803) & (!n_n4804) & (n_n4802) & (!n_n4805) & (!n_n4799)) + ((n_n4803) & (!n_n4804) & (n_n4802) & (!n_n4805) & (n_n4799)) + ((n_n4803) & (!n_n4804) & (n_n4802) & (n_n4805) & (!n_n4799)) + ((n_n4803) & (!n_n4804) & (n_n4802) & (n_n4805) & (n_n4799)) + ((n_n4803) & (n_n4804) & (!n_n4802) & (!n_n4805) & (!n_n4799)) + ((n_n4803) & (n_n4804) & (!n_n4802) & (!n_n4805) & (n_n4799)) + ((n_n4803) & (n_n4804) & (!n_n4802) & (n_n4805) & (!n_n4799)) + ((n_n4803) & (n_n4804) & (!n_n4802) & (n_n4805) & (n_n4799)) + ((n_n4803) & (n_n4804) & (n_n4802) & (!n_n4805) & (!n_n4799)) + ((n_n4803) & (n_n4804) & (n_n4802) & (!n_n4805) & (n_n4799)) + ((n_n4803) & (n_n4804) & (n_n4802) & (n_n4805) & (!n_n4799)) + ((n_n4803) & (n_n4804) & (n_n4802) & (n_n4805) & (n_n4799)));
	assign x16192x = (((!i_9_) & (n_n534) & (n_n260) & (n_n535)) + ((i_9_) & (n_n534) & (n_n260) & (n_n535)));
	assign x16198x = (((!n_n4832) & (!n_n4812) & (!x388x) & (!n_n4197) & (x16192x)) + ((!n_n4832) & (!n_n4812) & (!x388x) & (n_n4197) & (!x16192x)) + ((!n_n4832) & (!n_n4812) & (!x388x) & (n_n4197) & (x16192x)) + ((!n_n4832) & (!n_n4812) & (x388x) & (!n_n4197) & (!x16192x)) + ((!n_n4832) & (!n_n4812) & (x388x) & (!n_n4197) & (x16192x)) + ((!n_n4832) & (!n_n4812) & (x388x) & (n_n4197) & (!x16192x)) + ((!n_n4832) & (!n_n4812) & (x388x) & (n_n4197) & (x16192x)) + ((!n_n4832) & (n_n4812) & (!x388x) & (!n_n4197) & (!x16192x)) + ((!n_n4832) & (n_n4812) & (!x388x) & (!n_n4197) & (x16192x)) + ((!n_n4832) & (n_n4812) & (!x388x) & (n_n4197) & (!x16192x)) + ((!n_n4832) & (n_n4812) & (!x388x) & (n_n4197) & (x16192x)) + ((!n_n4832) & (n_n4812) & (x388x) & (!n_n4197) & (!x16192x)) + ((!n_n4832) & (n_n4812) & (x388x) & (!n_n4197) & (x16192x)) + ((!n_n4832) & (n_n4812) & (x388x) & (n_n4197) & (!x16192x)) + ((!n_n4832) & (n_n4812) & (x388x) & (n_n4197) & (x16192x)) + ((n_n4832) & (!n_n4812) & (!x388x) & (!n_n4197) & (!x16192x)) + ((n_n4832) & (!n_n4812) & (!x388x) & (!n_n4197) & (x16192x)) + ((n_n4832) & (!n_n4812) & (!x388x) & (n_n4197) & (!x16192x)) + ((n_n4832) & (!n_n4812) & (!x388x) & (n_n4197) & (x16192x)) + ((n_n4832) & (!n_n4812) & (x388x) & (!n_n4197) & (!x16192x)) + ((n_n4832) & (!n_n4812) & (x388x) & (!n_n4197) & (x16192x)) + ((n_n4832) & (!n_n4812) & (x388x) & (n_n4197) & (!x16192x)) + ((n_n4832) & (!n_n4812) & (x388x) & (n_n4197) & (x16192x)) + ((n_n4832) & (n_n4812) & (!x388x) & (!n_n4197) & (!x16192x)) + ((n_n4832) & (n_n4812) & (!x388x) & (!n_n4197) & (x16192x)) + ((n_n4832) & (n_n4812) & (!x388x) & (n_n4197) & (!x16192x)) + ((n_n4832) & (n_n4812) & (!x388x) & (n_n4197) & (x16192x)) + ((n_n4832) & (n_n4812) & (x388x) & (!n_n4197) & (!x16192x)) + ((n_n4832) & (n_n4812) & (x388x) & (!n_n4197) & (x16192x)) + ((n_n4832) & (n_n4812) & (x388x) & (n_n4197) & (!x16192x)) + ((n_n4832) & (n_n4812) & (x388x) & (n_n4197) & (x16192x)));
	assign x16197x = (((!n_n4816) & (!n_n4818) & (!n_n4815) & (!x150x) & (x303x)) + ((!n_n4816) & (!n_n4818) & (!n_n4815) & (x150x) & (!x303x)) + ((!n_n4816) & (!n_n4818) & (!n_n4815) & (x150x) & (x303x)) + ((!n_n4816) & (!n_n4818) & (n_n4815) & (!x150x) & (!x303x)) + ((!n_n4816) & (!n_n4818) & (n_n4815) & (!x150x) & (x303x)) + ((!n_n4816) & (!n_n4818) & (n_n4815) & (x150x) & (!x303x)) + ((!n_n4816) & (!n_n4818) & (n_n4815) & (x150x) & (x303x)) + ((!n_n4816) & (n_n4818) & (!n_n4815) & (!x150x) & (!x303x)) + ((!n_n4816) & (n_n4818) & (!n_n4815) & (!x150x) & (x303x)) + ((!n_n4816) & (n_n4818) & (!n_n4815) & (x150x) & (!x303x)) + ((!n_n4816) & (n_n4818) & (!n_n4815) & (x150x) & (x303x)) + ((!n_n4816) & (n_n4818) & (n_n4815) & (!x150x) & (!x303x)) + ((!n_n4816) & (n_n4818) & (n_n4815) & (!x150x) & (x303x)) + ((!n_n4816) & (n_n4818) & (n_n4815) & (x150x) & (!x303x)) + ((!n_n4816) & (n_n4818) & (n_n4815) & (x150x) & (x303x)) + ((n_n4816) & (!n_n4818) & (!n_n4815) & (!x150x) & (!x303x)) + ((n_n4816) & (!n_n4818) & (!n_n4815) & (!x150x) & (x303x)) + ((n_n4816) & (!n_n4818) & (!n_n4815) & (x150x) & (!x303x)) + ((n_n4816) & (!n_n4818) & (!n_n4815) & (x150x) & (x303x)) + ((n_n4816) & (!n_n4818) & (n_n4815) & (!x150x) & (!x303x)) + ((n_n4816) & (!n_n4818) & (n_n4815) & (!x150x) & (x303x)) + ((n_n4816) & (!n_n4818) & (n_n4815) & (x150x) & (!x303x)) + ((n_n4816) & (!n_n4818) & (n_n4815) & (x150x) & (x303x)) + ((n_n4816) & (n_n4818) & (!n_n4815) & (!x150x) & (!x303x)) + ((n_n4816) & (n_n4818) & (!n_n4815) & (!x150x) & (x303x)) + ((n_n4816) & (n_n4818) & (!n_n4815) & (x150x) & (!x303x)) + ((n_n4816) & (n_n4818) & (!n_n4815) & (x150x) & (x303x)) + ((n_n4816) & (n_n4818) & (n_n4815) & (!x150x) & (!x303x)) + ((n_n4816) & (n_n4818) & (n_n4815) & (!x150x) & (x303x)) + ((n_n4816) & (n_n4818) & (n_n4815) & (x150x) & (!x303x)) + ((n_n4816) & (n_n4818) & (n_n4815) & (x150x) & (x303x)));
	assign n_n1808 = (((!x16189x) & (!x16190x) & (!x16198x) & (x16197x)) + ((!x16189x) & (!x16190x) & (x16198x) & (!x16197x)) + ((!x16189x) & (!x16190x) & (x16198x) & (x16197x)) + ((!x16189x) & (x16190x) & (!x16198x) & (!x16197x)) + ((!x16189x) & (x16190x) & (!x16198x) & (x16197x)) + ((!x16189x) & (x16190x) & (x16198x) & (!x16197x)) + ((!x16189x) & (x16190x) & (x16198x) & (x16197x)) + ((x16189x) & (!x16190x) & (!x16198x) & (!x16197x)) + ((x16189x) & (!x16190x) & (!x16198x) & (x16197x)) + ((x16189x) & (!x16190x) & (x16198x) & (!x16197x)) + ((x16189x) & (!x16190x) & (x16198x) & (x16197x)) + ((x16189x) & (x16190x) & (!x16198x) & (!x16197x)) + ((x16189x) & (x16190x) & (!x16198x) & (x16197x)) + ((x16189x) & (x16190x) & (x16198x) & (!x16197x)) + ((x16189x) & (x16190x) & (x16198x) & (x16197x)));
	assign x22070x = (((!n_n4857) & (!n_n4854) & (!n_n4855) & (!n_n4858)));
	assign n_n1858 = (((!n_n4847) & (!n_n4846) & (!n_n4848) & (!x375x) & (!x22070x)) + ((!n_n4847) & (!n_n4846) & (!n_n4848) & (x375x) & (!x22070x)) + ((!n_n4847) & (!n_n4846) & (!n_n4848) & (x375x) & (x22070x)) + ((!n_n4847) & (!n_n4846) & (n_n4848) & (!x375x) & (!x22070x)) + ((!n_n4847) & (!n_n4846) & (n_n4848) & (!x375x) & (x22070x)) + ((!n_n4847) & (!n_n4846) & (n_n4848) & (x375x) & (!x22070x)) + ((!n_n4847) & (!n_n4846) & (n_n4848) & (x375x) & (x22070x)) + ((!n_n4847) & (n_n4846) & (!n_n4848) & (!x375x) & (!x22070x)) + ((!n_n4847) & (n_n4846) & (!n_n4848) & (!x375x) & (x22070x)) + ((!n_n4847) & (n_n4846) & (!n_n4848) & (x375x) & (!x22070x)) + ((!n_n4847) & (n_n4846) & (!n_n4848) & (x375x) & (x22070x)) + ((!n_n4847) & (n_n4846) & (n_n4848) & (!x375x) & (!x22070x)) + ((!n_n4847) & (n_n4846) & (n_n4848) & (!x375x) & (x22070x)) + ((!n_n4847) & (n_n4846) & (n_n4848) & (x375x) & (!x22070x)) + ((!n_n4847) & (n_n4846) & (n_n4848) & (x375x) & (x22070x)) + ((n_n4847) & (!n_n4846) & (!n_n4848) & (!x375x) & (!x22070x)) + ((n_n4847) & (!n_n4846) & (!n_n4848) & (!x375x) & (x22070x)) + ((n_n4847) & (!n_n4846) & (!n_n4848) & (x375x) & (!x22070x)) + ((n_n4847) & (!n_n4846) & (!n_n4848) & (x375x) & (x22070x)) + ((n_n4847) & (!n_n4846) & (n_n4848) & (!x375x) & (!x22070x)) + ((n_n4847) & (!n_n4846) & (n_n4848) & (!x375x) & (x22070x)) + ((n_n4847) & (!n_n4846) & (n_n4848) & (x375x) & (!x22070x)) + ((n_n4847) & (!n_n4846) & (n_n4848) & (x375x) & (x22070x)) + ((n_n4847) & (n_n4846) & (!n_n4848) & (!x375x) & (!x22070x)) + ((n_n4847) & (n_n4846) & (!n_n4848) & (!x375x) & (x22070x)) + ((n_n4847) & (n_n4846) & (!n_n4848) & (x375x) & (!x22070x)) + ((n_n4847) & (n_n4846) & (!n_n4848) & (x375x) & (x22070x)) + ((n_n4847) & (n_n4846) & (n_n4848) & (!x375x) & (!x22070x)) + ((n_n4847) & (n_n4846) & (n_n4848) & (!x375x) & (x22070x)) + ((n_n4847) & (n_n4846) & (n_n4848) & (x375x) & (!x22070x)) + ((n_n4847) & (n_n4846) & (n_n4848) & (x375x) & (x22070x)));
	assign n_n1857 = (((!x40x) & (!n_n4859) & (!n_n4864) & (!x246x) & (n_n1988)) + ((!x40x) & (!n_n4859) & (!n_n4864) & (x246x) & (!n_n1988)) + ((!x40x) & (!n_n4859) & (!n_n4864) & (x246x) & (n_n1988)) + ((!x40x) & (!n_n4859) & (n_n4864) & (!x246x) & (!n_n1988)) + ((!x40x) & (!n_n4859) & (n_n4864) & (!x246x) & (n_n1988)) + ((!x40x) & (!n_n4859) & (n_n4864) & (x246x) & (!n_n1988)) + ((!x40x) & (!n_n4859) & (n_n4864) & (x246x) & (n_n1988)) + ((!x40x) & (n_n4859) & (!n_n4864) & (!x246x) & (!n_n1988)) + ((!x40x) & (n_n4859) & (!n_n4864) & (!x246x) & (n_n1988)) + ((!x40x) & (n_n4859) & (!n_n4864) & (x246x) & (!n_n1988)) + ((!x40x) & (n_n4859) & (!n_n4864) & (x246x) & (n_n1988)) + ((!x40x) & (n_n4859) & (n_n4864) & (!x246x) & (!n_n1988)) + ((!x40x) & (n_n4859) & (n_n4864) & (!x246x) & (n_n1988)) + ((!x40x) & (n_n4859) & (n_n4864) & (x246x) & (!n_n1988)) + ((!x40x) & (n_n4859) & (n_n4864) & (x246x) & (n_n1988)) + ((x40x) & (!n_n4859) & (!n_n4864) & (!x246x) & (!n_n1988)) + ((x40x) & (!n_n4859) & (!n_n4864) & (!x246x) & (n_n1988)) + ((x40x) & (!n_n4859) & (!n_n4864) & (x246x) & (!n_n1988)) + ((x40x) & (!n_n4859) & (!n_n4864) & (x246x) & (n_n1988)) + ((x40x) & (!n_n4859) & (n_n4864) & (!x246x) & (!n_n1988)) + ((x40x) & (!n_n4859) & (n_n4864) & (!x246x) & (n_n1988)) + ((x40x) & (!n_n4859) & (n_n4864) & (x246x) & (!n_n1988)) + ((x40x) & (!n_n4859) & (n_n4864) & (x246x) & (n_n1988)) + ((x40x) & (n_n4859) & (!n_n4864) & (!x246x) & (!n_n1988)) + ((x40x) & (n_n4859) & (!n_n4864) & (!x246x) & (n_n1988)) + ((x40x) & (n_n4859) & (!n_n4864) & (x246x) & (!n_n1988)) + ((x40x) & (n_n4859) & (!n_n4864) & (x246x) & (n_n1988)) + ((x40x) & (n_n4859) & (n_n4864) & (!x246x) & (!n_n1988)) + ((x40x) & (n_n4859) & (n_n4864) & (!x246x) & (n_n1988)) + ((x40x) & (n_n4859) & (n_n4864) & (x246x) & (!n_n1988)) + ((x40x) & (n_n4859) & (n_n4864) & (x246x) & (n_n1988)));
	assign x16211x = (((!i_9_) & (!n_n524) & (!x552x) & (!n_n4843) & (x177x)) + ((!i_9_) & (!n_n524) & (!x552x) & (n_n4843) & (!x177x)) + ((!i_9_) & (!n_n524) & (!x552x) & (n_n4843) & (x177x)) + ((!i_9_) & (!n_n524) & (x552x) & (!n_n4843) & (x177x)) + ((!i_9_) & (!n_n524) & (x552x) & (n_n4843) & (!x177x)) + ((!i_9_) & (!n_n524) & (x552x) & (n_n4843) & (x177x)) + ((!i_9_) & (n_n524) & (!x552x) & (!n_n4843) & (x177x)) + ((!i_9_) & (n_n524) & (!x552x) & (n_n4843) & (!x177x)) + ((!i_9_) & (n_n524) & (!x552x) & (n_n4843) & (x177x)) + ((!i_9_) & (n_n524) & (x552x) & (!n_n4843) & (!x177x)) + ((!i_9_) & (n_n524) & (x552x) & (!n_n4843) & (x177x)) + ((!i_9_) & (n_n524) & (x552x) & (n_n4843) & (!x177x)) + ((!i_9_) & (n_n524) & (x552x) & (n_n4843) & (x177x)) + ((i_9_) & (!n_n524) & (!x552x) & (!n_n4843) & (x177x)) + ((i_9_) & (!n_n524) & (!x552x) & (n_n4843) & (!x177x)) + ((i_9_) & (!n_n524) & (!x552x) & (n_n4843) & (x177x)) + ((i_9_) & (!n_n524) & (x552x) & (!n_n4843) & (x177x)) + ((i_9_) & (!n_n524) & (x552x) & (n_n4843) & (!x177x)) + ((i_9_) & (!n_n524) & (x552x) & (n_n4843) & (x177x)) + ((i_9_) & (n_n524) & (!x552x) & (!n_n4843) & (x177x)) + ((i_9_) & (n_n524) & (!x552x) & (n_n4843) & (!x177x)) + ((i_9_) & (n_n524) & (!x552x) & (n_n4843) & (x177x)) + ((i_9_) & (n_n524) & (x552x) & (!n_n4843) & (x177x)) + ((i_9_) & (n_n524) & (x552x) & (n_n4843) & (!x177x)) + ((i_9_) & (n_n524) & (x552x) & (n_n4843) & (x177x)));
	assign x16212x = (((!n_n4845) & (!n_n4836) & (!n_n4838) & (!n_n4841) & (n_n4844)) + ((!n_n4845) & (!n_n4836) & (!n_n4838) & (n_n4841) & (!n_n4844)) + ((!n_n4845) & (!n_n4836) & (!n_n4838) & (n_n4841) & (n_n4844)) + ((!n_n4845) & (!n_n4836) & (n_n4838) & (!n_n4841) & (!n_n4844)) + ((!n_n4845) & (!n_n4836) & (n_n4838) & (!n_n4841) & (n_n4844)) + ((!n_n4845) & (!n_n4836) & (n_n4838) & (n_n4841) & (!n_n4844)) + ((!n_n4845) & (!n_n4836) & (n_n4838) & (n_n4841) & (n_n4844)) + ((!n_n4845) & (n_n4836) & (!n_n4838) & (!n_n4841) & (!n_n4844)) + ((!n_n4845) & (n_n4836) & (!n_n4838) & (!n_n4841) & (n_n4844)) + ((!n_n4845) & (n_n4836) & (!n_n4838) & (n_n4841) & (!n_n4844)) + ((!n_n4845) & (n_n4836) & (!n_n4838) & (n_n4841) & (n_n4844)) + ((!n_n4845) & (n_n4836) & (n_n4838) & (!n_n4841) & (!n_n4844)) + ((!n_n4845) & (n_n4836) & (n_n4838) & (!n_n4841) & (n_n4844)) + ((!n_n4845) & (n_n4836) & (n_n4838) & (n_n4841) & (!n_n4844)) + ((!n_n4845) & (n_n4836) & (n_n4838) & (n_n4841) & (n_n4844)) + ((n_n4845) & (!n_n4836) & (!n_n4838) & (!n_n4841) & (!n_n4844)) + ((n_n4845) & (!n_n4836) & (!n_n4838) & (!n_n4841) & (n_n4844)) + ((n_n4845) & (!n_n4836) & (!n_n4838) & (n_n4841) & (!n_n4844)) + ((n_n4845) & (!n_n4836) & (!n_n4838) & (n_n4841) & (n_n4844)) + ((n_n4845) & (!n_n4836) & (n_n4838) & (!n_n4841) & (!n_n4844)) + ((n_n4845) & (!n_n4836) & (n_n4838) & (!n_n4841) & (n_n4844)) + ((n_n4845) & (!n_n4836) & (n_n4838) & (n_n4841) & (!n_n4844)) + ((n_n4845) & (!n_n4836) & (n_n4838) & (n_n4841) & (n_n4844)) + ((n_n4845) & (n_n4836) & (!n_n4838) & (!n_n4841) & (!n_n4844)) + ((n_n4845) & (n_n4836) & (!n_n4838) & (!n_n4841) & (n_n4844)) + ((n_n4845) & (n_n4836) & (!n_n4838) & (n_n4841) & (!n_n4844)) + ((n_n4845) & (n_n4836) & (!n_n4838) & (n_n4841) & (n_n4844)) + ((n_n4845) & (n_n4836) & (n_n4838) & (!n_n4841) & (!n_n4844)) + ((n_n4845) & (n_n4836) & (n_n4838) & (!n_n4841) & (n_n4844)) + ((n_n4845) & (n_n4836) & (n_n4838) & (n_n4841) & (!n_n4844)) + ((n_n4845) & (n_n4836) & (n_n4838) & (n_n4841) & (n_n4844)));
	assign n_n1807 = (((!n_n1858) & (!n_n1857) & (!x16211x) & (x16212x)) + ((!n_n1858) & (!n_n1857) & (x16211x) & (!x16212x)) + ((!n_n1858) & (!n_n1857) & (x16211x) & (x16212x)) + ((!n_n1858) & (n_n1857) & (!x16211x) & (!x16212x)) + ((!n_n1858) & (n_n1857) & (!x16211x) & (x16212x)) + ((!n_n1858) & (n_n1857) & (x16211x) & (!x16212x)) + ((!n_n1858) & (n_n1857) & (x16211x) & (x16212x)) + ((n_n1858) & (!n_n1857) & (!x16211x) & (!x16212x)) + ((n_n1858) & (!n_n1857) & (!x16211x) & (x16212x)) + ((n_n1858) & (!n_n1857) & (x16211x) & (!x16212x)) + ((n_n1858) & (!n_n1857) & (x16211x) & (x16212x)) + ((n_n1858) & (n_n1857) & (!x16211x) & (!x16212x)) + ((n_n1858) & (n_n1857) & (!x16211x) & (x16212x)) + ((n_n1858) & (n_n1857) & (x16211x) & (!x16212x)) + ((n_n1858) & (n_n1857) & (x16211x) & (x16212x)));
	assign x16215x = (((!i_9_) & (n_n528) & (n_n260) & (n_n500)) + ((i_9_) & (n_n528) & (n_n260) & (n_n500)));
	assign n_n1856 = (((!n_n4875) & (!n_n4876) & (!x461x) & (!x263x) & (x16215x)) + ((!n_n4875) & (!n_n4876) & (!x461x) & (x263x) & (!x16215x)) + ((!n_n4875) & (!n_n4876) & (!x461x) & (x263x) & (x16215x)) + ((!n_n4875) & (!n_n4876) & (x461x) & (!x263x) & (!x16215x)) + ((!n_n4875) & (!n_n4876) & (x461x) & (!x263x) & (x16215x)) + ((!n_n4875) & (!n_n4876) & (x461x) & (x263x) & (!x16215x)) + ((!n_n4875) & (!n_n4876) & (x461x) & (x263x) & (x16215x)) + ((!n_n4875) & (n_n4876) & (!x461x) & (!x263x) & (!x16215x)) + ((!n_n4875) & (n_n4876) & (!x461x) & (!x263x) & (x16215x)) + ((!n_n4875) & (n_n4876) & (!x461x) & (x263x) & (!x16215x)) + ((!n_n4875) & (n_n4876) & (!x461x) & (x263x) & (x16215x)) + ((!n_n4875) & (n_n4876) & (x461x) & (!x263x) & (!x16215x)) + ((!n_n4875) & (n_n4876) & (x461x) & (!x263x) & (x16215x)) + ((!n_n4875) & (n_n4876) & (x461x) & (x263x) & (!x16215x)) + ((!n_n4875) & (n_n4876) & (x461x) & (x263x) & (x16215x)) + ((n_n4875) & (!n_n4876) & (!x461x) & (!x263x) & (!x16215x)) + ((n_n4875) & (!n_n4876) & (!x461x) & (!x263x) & (x16215x)) + ((n_n4875) & (!n_n4876) & (!x461x) & (x263x) & (!x16215x)) + ((n_n4875) & (!n_n4876) & (!x461x) & (x263x) & (x16215x)) + ((n_n4875) & (!n_n4876) & (x461x) & (!x263x) & (!x16215x)) + ((n_n4875) & (!n_n4876) & (x461x) & (!x263x) & (x16215x)) + ((n_n4875) & (!n_n4876) & (x461x) & (x263x) & (!x16215x)) + ((n_n4875) & (!n_n4876) & (x461x) & (x263x) & (x16215x)) + ((n_n4875) & (n_n4876) & (!x461x) & (!x263x) & (!x16215x)) + ((n_n4875) & (n_n4876) & (!x461x) & (!x263x) & (x16215x)) + ((n_n4875) & (n_n4876) & (!x461x) & (x263x) & (!x16215x)) + ((n_n4875) & (n_n4876) & (!x461x) & (x263x) & (x16215x)) + ((n_n4875) & (n_n4876) & (x461x) & (!x263x) & (!x16215x)) + ((n_n4875) & (n_n4876) & (x461x) & (!x263x) & (x16215x)) + ((n_n4875) & (n_n4876) & (x461x) & (x263x) & (!x16215x)) + ((n_n4875) & (n_n4876) & (x461x) & (x263x) & (x16215x)));
	assign x16222x = (((!n_n4886) & (!x264x) & (!n_n4891) & (!n_n1985) & (x261x)) + ((!n_n4886) & (!x264x) & (!n_n4891) & (n_n1985) & (!x261x)) + ((!n_n4886) & (!x264x) & (!n_n4891) & (n_n1985) & (x261x)) + ((!n_n4886) & (!x264x) & (n_n4891) & (!n_n1985) & (!x261x)) + ((!n_n4886) & (!x264x) & (n_n4891) & (!n_n1985) & (x261x)) + ((!n_n4886) & (!x264x) & (n_n4891) & (n_n1985) & (!x261x)) + ((!n_n4886) & (!x264x) & (n_n4891) & (n_n1985) & (x261x)) + ((!n_n4886) & (x264x) & (!n_n4891) & (!n_n1985) & (!x261x)) + ((!n_n4886) & (x264x) & (!n_n4891) & (!n_n1985) & (x261x)) + ((!n_n4886) & (x264x) & (!n_n4891) & (n_n1985) & (!x261x)) + ((!n_n4886) & (x264x) & (!n_n4891) & (n_n1985) & (x261x)) + ((!n_n4886) & (x264x) & (n_n4891) & (!n_n1985) & (!x261x)) + ((!n_n4886) & (x264x) & (n_n4891) & (!n_n1985) & (x261x)) + ((!n_n4886) & (x264x) & (n_n4891) & (n_n1985) & (!x261x)) + ((!n_n4886) & (x264x) & (n_n4891) & (n_n1985) & (x261x)) + ((n_n4886) & (!x264x) & (!n_n4891) & (!n_n1985) & (!x261x)) + ((n_n4886) & (!x264x) & (!n_n4891) & (!n_n1985) & (x261x)) + ((n_n4886) & (!x264x) & (!n_n4891) & (n_n1985) & (!x261x)) + ((n_n4886) & (!x264x) & (!n_n4891) & (n_n1985) & (x261x)) + ((n_n4886) & (!x264x) & (n_n4891) & (!n_n1985) & (!x261x)) + ((n_n4886) & (!x264x) & (n_n4891) & (!n_n1985) & (x261x)) + ((n_n4886) & (!x264x) & (n_n4891) & (n_n1985) & (!x261x)) + ((n_n4886) & (!x264x) & (n_n4891) & (n_n1985) & (x261x)) + ((n_n4886) & (x264x) & (!n_n4891) & (!n_n1985) & (!x261x)) + ((n_n4886) & (x264x) & (!n_n4891) & (!n_n1985) & (x261x)) + ((n_n4886) & (x264x) & (!n_n4891) & (n_n1985) & (!x261x)) + ((n_n4886) & (x264x) & (!n_n4891) & (n_n1985) & (x261x)) + ((n_n4886) & (x264x) & (n_n4891) & (!n_n1985) & (!x261x)) + ((n_n4886) & (x264x) & (n_n4891) & (!n_n1985) & (x261x)) + ((n_n4886) & (x264x) & (n_n4891) & (n_n1985) & (!x261x)) + ((n_n4886) & (x264x) & (n_n4891) & (n_n1985) & (x261x)));
	assign x15852x = (((!x20x) & (!n_n4860) & (!n_n4868) & (!x530x) & (n_n4842)) + ((!x20x) & (!n_n4860) & (!n_n4868) & (x530x) & (n_n4842)) + ((!x20x) & (!n_n4860) & (n_n4868) & (!x530x) & (!n_n4842)) + ((!x20x) & (!n_n4860) & (n_n4868) & (!x530x) & (n_n4842)) + ((!x20x) & (!n_n4860) & (n_n4868) & (x530x) & (!n_n4842)) + ((!x20x) & (!n_n4860) & (n_n4868) & (x530x) & (n_n4842)) + ((!x20x) & (n_n4860) & (!n_n4868) & (!x530x) & (!n_n4842)) + ((!x20x) & (n_n4860) & (!n_n4868) & (!x530x) & (n_n4842)) + ((!x20x) & (n_n4860) & (!n_n4868) & (x530x) & (!n_n4842)) + ((!x20x) & (n_n4860) & (!n_n4868) & (x530x) & (n_n4842)) + ((!x20x) & (n_n4860) & (n_n4868) & (!x530x) & (!n_n4842)) + ((!x20x) & (n_n4860) & (n_n4868) & (!x530x) & (n_n4842)) + ((!x20x) & (n_n4860) & (n_n4868) & (x530x) & (!n_n4842)) + ((!x20x) & (n_n4860) & (n_n4868) & (x530x) & (n_n4842)) + ((x20x) & (!n_n4860) & (!n_n4868) & (!x530x) & (n_n4842)) + ((x20x) & (!n_n4860) & (!n_n4868) & (x530x) & (!n_n4842)) + ((x20x) & (!n_n4860) & (!n_n4868) & (x530x) & (n_n4842)) + ((x20x) & (!n_n4860) & (n_n4868) & (!x530x) & (!n_n4842)) + ((x20x) & (!n_n4860) & (n_n4868) & (!x530x) & (n_n4842)) + ((x20x) & (!n_n4860) & (n_n4868) & (x530x) & (!n_n4842)) + ((x20x) & (!n_n4860) & (n_n4868) & (x530x) & (n_n4842)) + ((x20x) & (n_n4860) & (!n_n4868) & (!x530x) & (!n_n4842)) + ((x20x) & (n_n4860) & (!n_n4868) & (!x530x) & (n_n4842)) + ((x20x) & (n_n4860) & (!n_n4868) & (x530x) & (!n_n4842)) + ((x20x) & (n_n4860) & (!n_n4868) & (x530x) & (n_n4842)) + ((x20x) & (n_n4860) & (n_n4868) & (!x530x) & (!n_n4842)) + ((x20x) & (n_n4860) & (n_n4868) & (!x530x) & (n_n4842)) + ((x20x) & (n_n4860) & (n_n4868) & (x530x) & (!n_n4842)) + ((x20x) & (n_n4860) & (n_n4868) & (x530x) & (n_n4842)));
	assign x15853x = (((!n_n4849) & (!n_n4790) & (!n_n4801) & (!n_n4820) & (n_n4813)) + ((!n_n4849) & (!n_n4790) & (!n_n4801) & (n_n4820) & (!n_n4813)) + ((!n_n4849) & (!n_n4790) & (!n_n4801) & (n_n4820) & (n_n4813)) + ((!n_n4849) & (!n_n4790) & (n_n4801) & (!n_n4820) & (!n_n4813)) + ((!n_n4849) & (!n_n4790) & (n_n4801) & (!n_n4820) & (n_n4813)) + ((!n_n4849) & (!n_n4790) & (n_n4801) & (n_n4820) & (!n_n4813)) + ((!n_n4849) & (!n_n4790) & (n_n4801) & (n_n4820) & (n_n4813)) + ((!n_n4849) & (n_n4790) & (!n_n4801) & (!n_n4820) & (!n_n4813)) + ((!n_n4849) & (n_n4790) & (!n_n4801) & (!n_n4820) & (n_n4813)) + ((!n_n4849) & (n_n4790) & (!n_n4801) & (n_n4820) & (!n_n4813)) + ((!n_n4849) & (n_n4790) & (!n_n4801) & (n_n4820) & (n_n4813)) + ((!n_n4849) & (n_n4790) & (n_n4801) & (!n_n4820) & (!n_n4813)) + ((!n_n4849) & (n_n4790) & (n_n4801) & (!n_n4820) & (n_n4813)) + ((!n_n4849) & (n_n4790) & (n_n4801) & (n_n4820) & (!n_n4813)) + ((!n_n4849) & (n_n4790) & (n_n4801) & (n_n4820) & (n_n4813)) + ((n_n4849) & (!n_n4790) & (!n_n4801) & (!n_n4820) & (!n_n4813)) + ((n_n4849) & (!n_n4790) & (!n_n4801) & (!n_n4820) & (n_n4813)) + ((n_n4849) & (!n_n4790) & (!n_n4801) & (n_n4820) & (!n_n4813)) + ((n_n4849) & (!n_n4790) & (!n_n4801) & (n_n4820) & (n_n4813)) + ((n_n4849) & (!n_n4790) & (n_n4801) & (!n_n4820) & (!n_n4813)) + ((n_n4849) & (!n_n4790) & (n_n4801) & (!n_n4820) & (n_n4813)) + ((n_n4849) & (!n_n4790) & (n_n4801) & (n_n4820) & (!n_n4813)) + ((n_n4849) & (!n_n4790) & (n_n4801) & (n_n4820) & (n_n4813)) + ((n_n4849) & (n_n4790) & (!n_n4801) & (!n_n4820) & (!n_n4813)) + ((n_n4849) & (n_n4790) & (!n_n4801) & (!n_n4820) & (n_n4813)) + ((n_n4849) & (n_n4790) & (!n_n4801) & (n_n4820) & (!n_n4813)) + ((n_n4849) & (n_n4790) & (!n_n4801) & (n_n4820) & (n_n4813)) + ((n_n4849) & (n_n4790) & (n_n4801) & (!n_n4820) & (!n_n4813)) + ((n_n4849) & (n_n4790) & (n_n4801) & (!n_n4820) & (n_n4813)) + ((n_n4849) & (n_n4790) & (n_n4801) & (n_n4820) & (!n_n4813)) + ((n_n4849) & (n_n4790) & (n_n4801) & (n_n4820) & (n_n4813)));
	assign x15859x = (((!n_n4912) & (!n_n4968) & (!n_n4967) & (n_n4899)) + ((!n_n4912) & (!n_n4968) & (n_n4967) & (!n_n4899)) + ((!n_n4912) & (!n_n4968) & (n_n4967) & (n_n4899)) + ((!n_n4912) & (n_n4968) & (!n_n4967) & (!n_n4899)) + ((!n_n4912) & (n_n4968) & (!n_n4967) & (n_n4899)) + ((!n_n4912) & (n_n4968) & (n_n4967) & (!n_n4899)) + ((!n_n4912) & (n_n4968) & (n_n4967) & (n_n4899)) + ((n_n4912) & (!n_n4968) & (!n_n4967) & (!n_n4899)) + ((n_n4912) & (!n_n4968) & (!n_n4967) & (n_n4899)) + ((n_n4912) & (!n_n4968) & (n_n4967) & (!n_n4899)) + ((n_n4912) & (!n_n4968) & (n_n4967) & (n_n4899)) + ((n_n4912) & (n_n4968) & (!n_n4967) & (!n_n4899)) + ((n_n4912) & (n_n4968) & (!n_n4967) & (n_n4899)) + ((n_n4912) & (n_n4968) & (n_n4967) & (!n_n4899)) + ((n_n4912) & (n_n4968) & (n_n4967) & (n_n4899)));
	assign x15860x = (((!n_n4887) & (!n_n4929) & (!n_n4930) & (!n_n4915) & (n_n4961)) + ((!n_n4887) & (!n_n4929) & (!n_n4930) & (n_n4915) & (!n_n4961)) + ((!n_n4887) & (!n_n4929) & (!n_n4930) & (n_n4915) & (n_n4961)) + ((!n_n4887) & (!n_n4929) & (n_n4930) & (!n_n4915) & (!n_n4961)) + ((!n_n4887) & (!n_n4929) & (n_n4930) & (!n_n4915) & (n_n4961)) + ((!n_n4887) & (!n_n4929) & (n_n4930) & (n_n4915) & (!n_n4961)) + ((!n_n4887) & (!n_n4929) & (n_n4930) & (n_n4915) & (n_n4961)) + ((!n_n4887) & (n_n4929) & (!n_n4930) & (!n_n4915) & (!n_n4961)) + ((!n_n4887) & (n_n4929) & (!n_n4930) & (!n_n4915) & (n_n4961)) + ((!n_n4887) & (n_n4929) & (!n_n4930) & (n_n4915) & (!n_n4961)) + ((!n_n4887) & (n_n4929) & (!n_n4930) & (n_n4915) & (n_n4961)) + ((!n_n4887) & (n_n4929) & (n_n4930) & (!n_n4915) & (!n_n4961)) + ((!n_n4887) & (n_n4929) & (n_n4930) & (!n_n4915) & (n_n4961)) + ((!n_n4887) & (n_n4929) & (n_n4930) & (n_n4915) & (!n_n4961)) + ((!n_n4887) & (n_n4929) & (n_n4930) & (n_n4915) & (n_n4961)) + ((n_n4887) & (!n_n4929) & (!n_n4930) & (!n_n4915) & (!n_n4961)) + ((n_n4887) & (!n_n4929) & (!n_n4930) & (!n_n4915) & (n_n4961)) + ((n_n4887) & (!n_n4929) & (!n_n4930) & (n_n4915) & (!n_n4961)) + ((n_n4887) & (!n_n4929) & (!n_n4930) & (n_n4915) & (n_n4961)) + ((n_n4887) & (!n_n4929) & (n_n4930) & (!n_n4915) & (!n_n4961)) + ((n_n4887) & (!n_n4929) & (n_n4930) & (!n_n4915) & (n_n4961)) + ((n_n4887) & (!n_n4929) & (n_n4930) & (n_n4915) & (!n_n4961)) + ((n_n4887) & (!n_n4929) & (n_n4930) & (n_n4915) & (n_n4961)) + ((n_n4887) & (n_n4929) & (!n_n4930) & (!n_n4915) & (!n_n4961)) + ((n_n4887) & (n_n4929) & (!n_n4930) & (!n_n4915) & (n_n4961)) + ((n_n4887) & (n_n4929) & (!n_n4930) & (n_n4915) & (!n_n4961)) + ((n_n4887) & (n_n4929) & (!n_n4930) & (n_n4915) & (n_n4961)) + ((n_n4887) & (n_n4929) & (n_n4930) & (!n_n4915) & (!n_n4961)) + ((n_n4887) & (n_n4929) & (n_n4930) & (!n_n4915) & (n_n4961)) + ((n_n4887) & (n_n4929) & (n_n4930) & (n_n4915) & (!n_n4961)) + ((n_n4887) & (n_n4929) & (n_n4930) & (n_n4915) & (n_n4961)));
	assign x22075x = (((!n_n5001) & (!n_n4993) & (!n_n4994) & (!n_n5006) & (!n_n5007)));
	assign n_n1720 = (((!n_n5009) & (!n_n4978) & (!x248x) & (!x22075x)) + ((!n_n5009) & (!n_n4978) & (x248x) & (!x22075x)) + ((!n_n5009) & (!n_n4978) & (x248x) & (x22075x)) + ((!n_n5009) & (n_n4978) & (!x248x) & (!x22075x)) + ((!n_n5009) & (n_n4978) & (!x248x) & (x22075x)) + ((!n_n5009) & (n_n4978) & (x248x) & (!x22075x)) + ((!n_n5009) & (n_n4978) & (x248x) & (x22075x)) + ((n_n5009) & (!n_n4978) & (!x248x) & (!x22075x)) + ((n_n5009) & (!n_n4978) & (!x248x) & (x22075x)) + ((n_n5009) & (!n_n4978) & (x248x) & (!x22075x)) + ((n_n5009) & (!n_n4978) & (x248x) & (x22075x)) + ((n_n5009) & (n_n4978) & (!x248x) & (!x22075x)) + ((n_n5009) & (n_n4978) & (!x248x) & (x22075x)) + ((n_n5009) & (n_n4978) & (x248x) & (!x22075x)) + ((n_n5009) & (n_n4978) & (x248x) & (x22075x)));
	assign x15886x = (((!n_n5034) & (!n_n5050) & (!n_n5063) & (!n_n5052) & (n_n5033)) + ((!n_n5034) & (!n_n5050) & (!n_n5063) & (n_n5052) & (!n_n5033)) + ((!n_n5034) & (!n_n5050) & (!n_n5063) & (n_n5052) & (n_n5033)) + ((!n_n5034) & (!n_n5050) & (n_n5063) & (!n_n5052) & (!n_n5033)) + ((!n_n5034) & (!n_n5050) & (n_n5063) & (!n_n5052) & (n_n5033)) + ((!n_n5034) & (!n_n5050) & (n_n5063) & (n_n5052) & (!n_n5033)) + ((!n_n5034) & (!n_n5050) & (n_n5063) & (n_n5052) & (n_n5033)) + ((!n_n5034) & (n_n5050) & (!n_n5063) & (!n_n5052) & (!n_n5033)) + ((!n_n5034) & (n_n5050) & (!n_n5063) & (!n_n5052) & (n_n5033)) + ((!n_n5034) & (n_n5050) & (!n_n5063) & (n_n5052) & (!n_n5033)) + ((!n_n5034) & (n_n5050) & (!n_n5063) & (n_n5052) & (n_n5033)) + ((!n_n5034) & (n_n5050) & (n_n5063) & (!n_n5052) & (!n_n5033)) + ((!n_n5034) & (n_n5050) & (n_n5063) & (!n_n5052) & (n_n5033)) + ((!n_n5034) & (n_n5050) & (n_n5063) & (n_n5052) & (!n_n5033)) + ((!n_n5034) & (n_n5050) & (n_n5063) & (n_n5052) & (n_n5033)) + ((n_n5034) & (!n_n5050) & (!n_n5063) & (!n_n5052) & (!n_n5033)) + ((n_n5034) & (!n_n5050) & (!n_n5063) & (!n_n5052) & (n_n5033)) + ((n_n5034) & (!n_n5050) & (!n_n5063) & (n_n5052) & (!n_n5033)) + ((n_n5034) & (!n_n5050) & (!n_n5063) & (n_n5052) & (n_n5033)) + ((n_n5034) & (!n_n5050) & (n_n5063) & (!n_n5052) & (!n_n5033)) + ((n_n5034) & (!n_n5050) & (n_n5063) & (!n_n5052) & (n_n5033)) + ((n_n5034) & (!n_n5050) & (n_n5063) & (n_n5052) & (!n_n5033)) + ((n_n5034) & (!n_n5050) & (n_n5063) & (n_n5052) & (n_n5033)) + ((n_n5034) & (n_n5050) & (!n_n5063) & (!n_n5052) & (!n_n5033)) + ((n_n5034) & (n_n5050) & (!n_n5063) & (!n_n5052) & (n_n5033)) + ((n_n5034) & (n_n5050) & (!n_n5063) & (n_n5052) & (!n_n5033)) + ((n_n5034) & (n_n5050) & (!n_n5063) & (n_n5052) & (n_n5033)) + ((n_n5034) & (n_n5050) & (n_n5063) & (!n_n5052) & (!n_n5033)) + ((n_n5034) & (n_n5050) & (n_n5063) & (!n_n5052) & (n_n5033)) + ((n_n5034) & (n_n5050) & (n_n5063) & (n_n5052) & (!n_n5033)) + ((n_n5034) & (n_n5050) & (n_n5063) & (n_n5052) & (n_n5033)));
	assign x15887x = (((!n_n5059) & (!n_n5046) & (!n_n5018) & (!n_n5022) & (x15886x)) + ((!n_n5059) & (!n_n5046) & (!n_n5018) & (n_n5022) & (!x15886x)) + ((!n_n5059) & (!n_n5046) & (!n_n5018) & (n_n5022) & (x15886x)) + ((!n_n5059) & (!n_n5046) & (n_n5018) & (!n_n5022) & (!x15886x)) + ((!n_n5059) & (!n_n5046) & (n_n5018) & (!n_n5022) & (x15886x)) + ((!n_n5059) & (!n_n5046) & (n_n5018) & (n_n5022) & (!x15886x)) + ((!n_n5059) & (!n_n5046) & (n_n5018) & (n_n5022) & (x15886x)) + ((!n_n5059) & (n_n5046) & (!n_n5018) & (!n_n5022) & (!x15886x)) + ((!n_n5059) & (n_n5046) & (!n_n5018) & (!n_n5022) & (x15886x)) + ((!n_n5059) & (n_n5046) & (!n_n5018) & (n_n5022) & (!x15886x)) + ((!n_n5059) & (n_n5046) & (!n_n5018) & (n_n5022) & (x15886x)) + ((!n_n5059) & (n_n5046) & (n_n5018) & (!n_n5022) & (!x15886x)) + ((!n_n5059) & (n_n5046) & (n_n5018) & (!n_n5022) & (x15886x)) + ((!n_n5059) & (n_n5046) & (n_n5018) & (n_n5022) & (!x15886x)) + ((!n_n5059) & (n_n5046) & (n_n5018) & (n_n5022) & (x15886x)) + ((n_n5059) & (!n_n5046) & (!n_n5018) & (!n_n5022) & (!x15886x)) + ((n_n5059) & (!n_n5046) & (!n_n5018) & (!n_n5022) & (x15886x)) + ((n_n5059) & (!n_n5046) & (!n_n5018) & (n_n5022) & (!x15886x)) + ((n_n5059) & (!n_n5046) & (!n_n5018) & (n_n5022) & (x15886x)) + ((n_n5059) & (!n_n5046) & (n_n5018) & (!n_n5022) & (!x15886x)) + ((n_n5059) & (!n_n5046) & (n_n5018) & (!n_n5022) & (x15886x)) + ((n_n5059) & (!n_n5046) & (n_n5018) & (n_n5022) & (!x15886x)) + ((n_n5059) & (!n_n5046) & (n_n5018) & (n_n5022) & (x15886x)) + ((n_n5059) & (n_n5046) & (!n_n5018) & (!n_n5022) & (!x15886x)) + ((n_n5059) & (n_n5046) & (!n_n5018) & (!n_n5022) & (x15886x)) + ((n_n5059) & (n_n5046) & (!n_n5018) & (n_n5022) & (!x15886x)) + ((n_n5059) & (n_n5046) & (!n_n5018) & (n_n5022) & (x15886x)) + ((n_n5059) & (n_n5046) & (n_n5018) & (!n_n5022) & (!x15886x)) + ((n_n5059) & (n_n5046) & (n_n5018) & (!n_n5022) & (x15886x)) + ((n_n5059) & (n_n5046) & (n_n5018) & (n_n5022) & (!x15886x)) + ((n_n5059) & (n_n5046) & (n_n5018) & (n_n5022) & (x15886x)));
	assign x15871x = (((!n_n5116) & (!n_n5098) & (!n_n5087) & (n_n5102)) + ((!n_n5116) & (!n_n5098) & (n_n5087) & (!n_n5102)) + ((!n_n5116) & (!n_n5098) & (n_n5087) & (n_n5102)) + ((!n_n5116) & (n_n5098) & (!n_n5087) & (!n_n5102)) + ((!n_n5116) & (n_n5098) & (!n_n5087) & (n_n5102)) + ((!n_n5116) & (n_n5098) & (n_n5087) & (!n_n5102)) + ((!n_n5116) & (n_n5098) & (n_n5087) & (n_n5102)) + ((n_n5116) & (!n_n5098) & (!n_n5087) & (!n_n5102)) + ((n_n5116) & (!n_n5098) & (!n_n5087) & (n_n5102)) + ((n_n5116) & (!n_n5098) & (n_n5087) & (!n_n5102)) + ((n_n5116) & (!n_n5098) & (n_n5087) & (n_n5102)) + ((n_n5116) & (n_n5098) & (!n_n5087) & (!n_n5102)) + ((n_n5116) & (n_n5098) & (!n_n5087) & (n_n5102)) + ((n_n5116) & (n_n5098) & (n_n5087) & (!n_n5102)) + ((n_n5116) & (n_n5098) & (n_n5087) & (n_n5102)));
	assign x15872x = (((!n_n5111) & (!n_n5081) & (!n_n5108) & (!n_n5078) & (n_n5080)) + ((!n_n5111) & (!n_n5081) & (!n_n5108) & (n_n5078) & (!n_n5080)) + ((!n_n5111) & (!n_n5081) & (!n_n5108) & (n_n5078) & (n_n5080)) + ((!n_n5111) & (!n_n5081) & (n_n5108) & (!n_n5078) & (!n_n5080)) + ((!n_n5111) & (!n_n5081) & (n_n5108) & (!n_n5078) & (n_n5080)) + ((!n_n5111) & (!n_n5081) & (n_n5108) & (n_n5078) & (!n_n5080)) + ((!n_n5111) & (!n_n5081) & (n_n5108) & (n_n5078) & (n_n5080)) + ((!n_n5111) & (n_n5081) & (!n_n5108) & (!n_n5078) & (!n_n5080)) + ((!n_n5111) & (n_n5081) & (!n_n5108) & (!n_n5078) & (n_n5080)) + ((!n_n5111) & (n_n5081) & (!n_n5108) & (n_n5078) & (!n_n5080)) + ((!n_n5111) & (n_n5081) & (!n_n5108) & (n_n5078) & (n_n5080)) + ((!n_n5111) & (n_n5081) & (n_n5108) & (!n_n5078) & (!n_n5080)) + ((!n_n5111) & (n_n5081) & (n_n5108) & (!n_n5078) & (n_n5080)) + ((!n_n5111) & (n_n5081) & (n_n5108) & (n_n5078) & (!n_n5080)) + ((!n_n5111) & (n_n5081) & (n_n5108) & (n_n5078) & (n_n5080)) + ((n_n5111) & (!n_n5081) & (!n_n5108) & (!n_n5078) & (!n_n5080)) + ((n_n5111) & (!n_n5081) & (!n_n5108) & (!n_n5078) & (n_n5080)) + ((n_n5111) & (!n_n5081) & (!n_n5108) & (n_n5078) & (!n_n5080)) + ((n_n5111) & (!n_n5081) & (!n_n5108) & (n_n5078) & (n_n5080)) + ((n_n5111) & (!n_n5081) & (n_n5108) & (!n_n5078) & (!n_n5080)) + ((n_n5111) & (!n_n5081) & (n_n5108) & (!n_n5078) & (n_n5080)) + ((n_n5111) & (!n_n5081) & (n_n5108) & (n_n5078) & (!n_n5080)) + ((n_n5111) & (!n_n5081) & (n_n5108) & (n_n5078) & (n_n5080)) + ((n_n5111) & (n_n5081) & (!n_n5108) & (!n_n5078) & (!n_n5080)) + ((n_n5111) & (n_n5081) & (!n_n5108) & (!n_n5078) & (n_n5080)) + ((n_n5111) & (n_n5081) & (!n_n5108) & (n_n5078) & (!n_n5080)) + ((n_n5111) & (n_n5081) & (!n_n5108) & (n_n5078) & (n_n5080)) + ((n_n5111) & (n_n5081) & (n_n5108) & (!n_n5078) & (!n_n5080)) + ((n_n5111) & (n_n5081) & (n_n5108) & (!n_n5078) & (n_n5080)) + ((n_n5111) & (n_n5081) & (n_n5108) & (n_n5078) & (!n_n5080)) + ((n_n5111) & (n_n5081) & (n_n5108) & (n_n5078) & (n_n5080)));
	assign n_n1717 = (((!n_n5131) & (!n_n5127) & (!n_n5190) & (!n_n5188) & (x15879x)) + ((!n_n5131) & (!n_n5127) & (!n_n5190) & (n_n5188) & (!x15879x)) + ((!n_n5131) & (!n_n5127) & (!n_n5190) & (n_n5188) & (x15879x)) + ((!n_n5131) & (!n_n5127) & (n_n5190) & (!n_n5188) & (!x15879x)) + ((!n_n5131) & (!n_n5127) & (n_n5190) & (!n_n5188) & (x15879x)) + ((!n_n5131) & (!n_n5127) & (n_n5190) & (n_n5188) & (!x15879x)) + ((!n_n5131) & (!n_n5127) & (n_n5190) & (n_n5188) & (x15879x)) + ((!n_n5131) & (n_n5127) & (!n_n5190) & (!n_n5188) & (!x15879x)) + ((!n_n5131) & (n_n5127) & (!n_n5190) & (!n_n5188) & (x15879x)) + ((!n_n5131) & (n_n5127) & (!n_n5190) & (n_n5188) & (!x15879x)) + ((!n_n5131) & (n_n5127) & (!n_n5190) & (n_n5188) & (x15879x)) + ((!n_n5131) & (n_n5127) & (n_n5190) & (!n_n5188) & (!x15879x)) + ((!n_n5131) & (n_n5127) & (n_n5190) & (!n_n5188) & (x15879x)) + ((!n_n5131) & (n_n5127) & (n_n5190) & (n_n5188) & (!x15879x)) + ((!n_n5131) & (n_n5127) & (n_n5190) & (n_n5188) & (x15879x)) + ((n_n5131) & (!n_n5127) & (!n_n5190) & (!n_n5188) & (!x15879x)) + ((n_n5131) & (!n_n5127) & (!n_n5190) & (!n_n5188) & (x15879x)) + ((n_n5131) & (!n_n5127) & (!n_n5190) & (n_n5188) & (!x15879x)) + ((n_n5131) & (!n_n5127) & (!n_n5190) & (n_n5188) & (x15879x)) + ((n_n5131) & (!n_n5127) & (n_n5190) & (!n_n5188) & (!x15879x)) + ((n_n5131) & (!n_n5127) & (n_n5190) & (!n_n5188) & (x15879x)) + ((n_n5131) & (!n_n5127) & (n_n5190) & (n_n5188) & (!x15879x)) + ((n_n5131) & (!n_n5127) & (n_n5190) & (n_n5188) & (x15879x)) + ((n_n5131) & (n_n5127) & (!n_n5190) & (!n_n5188) & (!x15879x)) + ((n_n5131) & (n_n5127) & (!n_n5190) & (!n_n5188) & (x15879x)) + ((n_n5131) & (n_n5127) & (!n_n5190) & (n_n5188) & (!x15879x)) + ((n_n5131) & (n_n5127) & (!n_n5190) & (n_n5188) & (x15879x)) + ((n_n5131) & (n_n5127) & (n_n5190) & (!n_n5188) & (!x15879x)) + ((n_n5131) & (n_n5127) & (n_n5190) & (!n_n5188) & (x15879x)) + ((n_n5131) & (n_n5127) & (n_n5190) & (n_n5188) & (!x15879x)) + ((n_n5131) & (n_n5127) & (n_n5190) & (n_n5188) & (x15879x)));
	assign x15894x = (((!n_n5214) & (!n_n5207) & (!n_n5229) & (n_n5221)) + ((!n_n5214) & (!n_n5207) & (n_n5229) & (!n_n5221)) + ((!n_n5214) & (!n_n5207) & (n_n5229) & (n_n5221)) + ((!n_n5214) & (n_n5207) & (!n_n5229) & (!n_n5221)) + ((!n_n5214) & (n_n5207) & (!n_n5229) & (n_n5221)) + ((!n_n5214) & (n_n5207) & (n_n5229) & (!n_n5221)) + ((!n_n5214) & (n_n5207) & (n_n5229) & (n_n5221)) + ((n_n5214) & (!n_n5207) & (!n_n5229) & (!n_n5221)) + ((n_n5214) & (!n_n5207) & (!n_n5229) & (n_n5221)) + ((n_n5214) & (!n_n5207) & (n_n5229) & (!n_n5221)) + ((n_n5214) & (!n_n5207) & (n_n5229) & (n_n5221)) + ((n_n5214) & (n_n5207) & (!n_n5229) & (!n_n5221)) + ((n_n5214) & (n_n5207) & (!n_n5229) & (n_n5221)) + ((n_n5214) & (n_n5207) & (n_n5229) & (!n_n5221)) + ((n_n5214) & (n_n5207) & (n_n5229) & (n_n5221)));
	assign x15895x = (((!n_n5200) & (!n_n5222) & (!n_n5218) & (!n_n5219) & (n_n5203)) + ((!n_n5200) & (!n_n5222) & (!n_n5218) & (n_n5219) & (!n_n5203)) + ((!n_n5200) & (!n_n5222) & (!n_n5218) & (n_n5219) & (n_n5203)) + ((!n_n5200) & (!n_n5222) & (n_n5218) & (!n_n5219) & (!n_n5203)) + ((!n_n5200) & (!n_n5222) & (n_n5218) & (!n_n5219) & (n_n5203)) + ((!n_n5200) & (!n_n5222) & (n_n5218) & (n_n5219) & (!n_n5203)) + ((!n_n5200) & (!n_n5222) & (n_n5218) & (n_n5219) & (n_n5203)) + ((!n_n5200) & (n_n5222) & (!n_n5218) & (!n_n5219) & (!n_n5203)) + ((!n_n5200) & (n_n5222) & (!n_n5218) & (!n_n5219) & (n_n5203)) + ((!n_n5200) & (n_n5222) & (!n_n5218) & (n_n5219) & (!n_n5203)) + ((!n_n5200) & (n_n5222) & (!n_n5218) & (n_n5219) & (n_n5203)) + ((!n_n5200) & (n_n5222) & (n_n5218) & (!n_n5219) & (!n_n5203)) + ((!n_n5200) & (n_n5222) & (n_n5218) & (!n_n5219) & (n_n5203)) + ((!n_n5200) & (n_n5222) & (n_n5218) & (n_n5219) & (!n_n5203)) + ((!n_n5200) & (n_n5222) & (n_n5218) & (n_n5219) & (n_n5203)) + ((n_n5200) & (!n_n5222) & (!n_n5218) & (!n_n5219) & (!n_n5203)) + ((n_n5200) & (!n_n5222) & (!n_n5218) & (!n_n5219) & (n_n5203)) + ((n_n5200) & (!n_n5222) & (!n_n5218) & (n_n5219) & (!n_n5203)) + ((n_n5200) & (!n_n5222) & (!n_n5218) & (n_n5219) & (n_n5203)) + ((n_n5200) & (!n_n5222) & (n_n5218) & (!n_n5219) & (!n_n5203)) + ((n_n5200) & (!n_n5222) & (n_n5218) & (!n_n5219) & (n_n5203)) + ((n_n5200) & (!n_n5222) & (n_n5218) & (n_n5219) & (!n_n5203)) + ((n_n5200) & (!n_n5222) & (n_n5218) & (n_n5219) & (n_n5203)) + ((n_n5200) & (n_n5222) & (!n_n5218) & (!n_n5219) & (!n_n5203)) + ((n_n5200) & (n_n5222) & (!n_n5218) & (!n_n5219) & (n_n5203)) + ((n_n5200) & (n_n5222) & (!n_n5218) & (n_n5219) & (!n_n5203)) + ((n_n5200) & (n_n5222) & (!n_n5218) & (n_n5219) & (n_n5203)) + ((n_n5200) & (n_n5222) & (n_n5218) & (!n_n5219) & (!n_n5203)) + ((n_n5200) & (n_n5222) & (n_n5218) & (!n_n5219) & (n_n5203)) + ((n_n5200) & (n_n5222) & (n_n5218) & (n_n5219) & (!n_n5203)) + ((n_n5200) & (n_n5222) & (n_n5218) & (n_n5219) & (n_n5203)));
	assign x11705x = (((!x12x) & (!x502x) & (!n_n5206) & (!n_n5182) & (n_n5172)) + ((!x12x) & (!x502x) & (!n_n5206) & (n_n5182) & (!n_n5172)) + ((!x12x) & (!x502x) & (!n_n5206) & (n_n5182) & (n_n5172)) + ((!x12x) & (!x502x) & (n_n5206) & (!n_n5182) & (!n_n5172)) + ((!x12x) & (!x502x) & (n_n5206) & (!n_n5182) & (n_n5172)) + ((!x12x) & (!x502x) & (n_n5206) & (n_n5182) & (!n_n5172)) + ((!x12x) & (!x502x) & (n_n5206) & (n_n5182) & (n_n5172)) + ((!x12x) & (x502x) & (!n_n5206) & (!n_n5182) & (n_n5172)) + ((!x12x) & (x502x) & (!n_n5206) & (n_n5182) & (!n_n5172)) + ((!x12x) & (x502x) & (!n_n5206) & (n_n5182) & (n_n5172)) + ((!x12x) & (x502x) & (n_n5206) & (!n_n5182) & (!n_n5172)) + ((!x12x) & (x502x) & (n_n5206) & (!n_n5182) & (n_n5172)) + ((!x12x) & (x502x) & (n_n5206) & (n_n5182) & (!n_n5172)) + ((!x12x) & (x502x) & (n_n5206) & (n_n5182) & (n_n5172)) + ((x12x) & (!x502x) & (!n_n5206) & (!n_n5182) & (n_n5172)) + ((x12x) & (!x502x) & (!n_n5206) & (n_n5182) & (!n_n5172)) + ((x12x) & (!x502x) & (!n_n5206) & (n_n5182) & (n_n5172)) + ((x12x) & (!x502x) & (n_n5206) & (!n_n5182) & (!n_n5172)) + ((x12x) & (!x502x) & (n_n5206) & (!n_n5182) & (n_n5172)) + ((x12x) & (!x502x) & (n_n5206) & (n_n5182) & (!n_n5172)) + ((x12x) & (!x502x) & (n_n5206) & (n_n5182) & (n_n5172)) + ((x12x) & (x502x) & (!n_n5206) & (!n_n5182) & (!n_n5172)) + ((x12x) & (x502x) & (!n_n5206) & (!n_n5182) & (n_n5172)) + ((x12x) & (x502x) & (!n_n5206) & (n_n5182) & (!n_n5172)) + ((x12x) & (x502x) & (!n_n5206) & (n_n5182) & (n_n5172)) + ((x12x) & (x502x) & (n_n5206) & (!n_n5182) & (!n_n5172)) + ((x12x) & (x502x) & (n_n5206) & (!n_n5182) & (n_n5172)) + ((x12x) & (x502x) & (n_n5206) & (n_n5182) & (!n_n5172)) + ((x12x) & (x502x) & (n_n5206) & (n_n5182) & (n_n5172)));
	assign x11706x = (((!n_n5191) & (!n_n5199) & (!n_n5209) & (!n_n5192) & (n_n5197)) + ((!n_n5191) & (!n_n5199) & (!n_n5209) & (n_n5192) & (!n_n5197)) + ((!n_n5191) & (!n_n5199) & (!n_n5209) & (n_n5192) & (n_n5197)) + ((!n_n5191) & (!n_n5199) & (n_n5209) & (!n_n5192) & (!n_n5197)) + ((!n_n5191) & (!n_n5199) & (n_n5209) & (!n_n5192) & (n_n5197)) + ((!n_n5191) & (!n_n5199) & (n_n5209) & (n_n5192) & (!n_n5197)) + ((!n_n5191) & (!n_n5199) & (n_n5209) & (n_n5192) & (n_n5197)) + ((!n_n5191) & (n_n5199) & (!n_n5209) & (!n_n5192) & (!n_n5197)) + ((!n_n5191) & (n_n5199) & (!n_n5209) & (!n_n5192) & (n_n5197)) + ((!n_n5191) & (n_n5199) & (!n_n5209) & (n_n5192) & (!n_n5197)) + ((!n_n5191) & (n_n5199) & (!n_n5209) & (n_n5192) & (n_n5197)) + ((!n_n5191) & (n_n5199) & (n_n5209) & (!n_n5192) & (!n_n5197)) + ((!n_n5191) & (n_n5199) & (n_n5209) & (!n_n5192) & (n_n5197)) + ((!n_n5191) & (n_n5199) & (n_n5209) & (n_n5192) & (!n_n5197)) + ((!n_n5191) & (n_n5199) & (n_n5209) & (n_n5192) & (n_n5197)) + ((n_n5191) & (!n_n5199) & (!n_n5209) & (!n_n5192) & (!n_n5197)) + ((n_n5191) & (!n_n5199) & (!n_n5209) & (!n_n5192) & (n_n5197)) + ((n_n5191) & (!n_n5199) & (!n_n5209) & (n_n5192) & (!n_n5197)) + ((n_n5191) & (!n_n5199) & (!n_n5209) & (n_n5192) & (n_n5197)) + ((n_n5191) & (!n_n5199) & (n_n5209) & (!n_n5192) & (!n_n5197)) + ((n_n5191) & (!n_n5199) & (n_n5209) & (!n_n5192) & (n_n5197)) + ((n_n5191) & (!n_n5199) & (n_n5209) & (n_n5192) & (!n_n5197)) + ((n_n5191) & (!n_n5199) & (n_n5209) & (n_n5192) & (n_n5197)) + ((n_n5191) & (n_n5199) & (!n_n5209) & (!n_n5192) & (!n_n5197)) + ((n_n5191) & (n_n5199) & (!n_n5209) & (!n_n5192) & (n_n5197)) + ((n_n5191) & (n_n5199) & (!n_n5209) & (n_n5192) & (!n_n5197)) + ((n_n5191) & (n_n5199) & (!n_n5209) & (n_n5192) & (n_n5197)) + ((n_n5191) & (n_n5199) & (n_n5209) & (!n_n5192) & (!n_n5197)) + ((n_n5191) & (n_n5199) & (n_n5209) & (!n_n5192) & (n_n5197)) + ((n_n5191) & (n_n5199) & (n_n5209) & (n_n5192) & (!n_n5197)) + ((n_n5191) & (n_n5199) & (n_n5209) & (n_n5192) & (n_n5197)));
	assign n_n738 = (((!n_n4318) & (!x171x) & (!n_n4322) & (!x284x) & (x364x)) + ((!n_n4318) & (!x171x) & (!n_n4322) & (x284x) & (!x364x)) + ((!n_n4318) & (!x171x) & (!n_n4322) & (x284x) & (x364x)) + ((!n_n4318) & (!x171x) & (n_n4322) & (!x284x) & (!x364x)) + ((!n_n4318) & (!x171x) & (n_n4322) & (!x284x) & (x364x)) + ((!n_n4318) & (!x171x) & (n_n4322) & (x284x) & (!x364x)) + ((!n_n4318) & (!x171x) & (n_n4322) & (x284x) & (x364x)) + ((!n_n4318) & (x171x) & (!n_n4322) & (!x284x) & (!x364x)) + ((!n_n4318) & (x171x) & (!n_n4322) & (!x284x) & (x364x)) + ((!n_n4318) & (x171x) & (!n_n4322) & (x284x) & (!x364x)) + ((!n_n4318) & (x171x) & (!n_n4322) & (x284x) & (x364x)) + ((!n_n4318) & (x171x) & (n_n4322) & (!x284x) & (!x364x)) + ((!n_n4318) & (x171x) & (n_n4322) & (!x284x) & (x364x)) + ((!n_n4318) & (x171x) & (n_n4322) & (x284x) & (!x364x)) + ((!n_n4318) & (x171x) & (n_n4322) & (x284x) & (x364x)) + ((n_n4318) & (!x171x) & (!n_n4322) & (!x284x) & (!x364x)) + ((n_n4318) & (!x171x) & (!n_n4322) & (!x284x) & (x364x)) + ((n_n4318) & (!x171x) & (!n_n4322) & (x284x) & (!x364x)) + ((n_n4318) & (!x171x) & (!n_n4322) & (x284x) & (x364x)) + ((n_n4318) & (!x171x) & (n_n4322) & (!x284x) & (!x364x)) + ((n_n4318) & (!x171x) & (n_n4322) & (!x284x) & (x364x)) + ((n_n4318) & (!x171x) & (n_n4322) & (x284x) & (!x364x)) + ((n_n4318) & (!x171x) & (n_n4322) & (x284x) & (x364x)) + ((n_n4318) & (x171x) & (!n_n4322) & (!x284x) & (!x364x)) + ((n_n4318) & (x171x) & (!n_n4322) & (!x284x) & (x364x)) + ((n_n4318) & (x171x) & (!n_n4322) & (x284x) & (!x364x)) + ((n_n4318) & (x171x) & (!n_n4322) & (x284x) & (x364x)) + ((n_n4318) & (x171x) & (n_n4322) & (!x284x) & (!x364x)) + ((n_n4318) & (x171x) & (n_n4322) & (!x284x) & (x364x)) + ((n_n4318) & (x171x) & (n_n4322) & (x284x) & (!x364x)) + ((n_n4318) & (x171x) & (n_n4322) & (x284x) & (x364x)));
	assign x13029x = (((!i_9_) & (!n_n526) & (n_n455) & (n_n528) & (n_n491)) + ((!i_9_) & (n_n526) & (n_n455) & (!n_n528) & (n_n491)) + ((!i_9_) & (n_n526) & (n_n455) & (n_n528) & (n_n491)) + ((i_9_) & (!n_n526) & (n_n455) & (n_n528) & (n_n491)) + ((i_9_) & (n_n526) & (n_n455) & (n_n528) & (n_n491)));
	assign n_n722 = (((!n_n4247) & (!x387x) & (x13029x)) + ((!n_n4247) & (x387x) & (!x13029x)) + ((!n_n4247) & (x387x) & (x13029x)) + ((n_n4247) & (!x387x) & (!x13029x)) + ((n_n4247) & (!x387x) & (x13029x)) + ((n_n4247) & (x387x) & (!x13029x)) + ((n_n4247) & (x387x) & (x13029x)));
	assign x346x = (((!i_9_) & (!n_n455) & (!n_n534) & (!n_n491) & (n_n4503)) + ((!i_9_) & (!n_n455) & (!n_n534) & (n_n491) & (n_n4503)) + ((!i_9_) & (!n_n455) & (n_n534) & (!n_n491) & (n_n4503)) + ((!i_9_) & (!n_n455) & (n_n534) & (n_n491) & (n_n4503)) + ((!i_9_) & (n_n455) & (!n_n534) & (!n_n491) & (n_n4503)) + ((!i_9_) & (n_n455) & (!n_n534) & (n_n491) & (n_n4503)) + ((!i_9_) & (n_n455) & (n_n534) & (!n_n491) & (n_n4503)) + ((!i_9_) & (n_n455) & (n_n534) & (n_n491) & (n_n4503)) + ((i_9_) & (!n_n455) & (!n_n534) & (!n_n491) & (n_n4503)) + ((i_9_) & (!n_n455) & (!n_n534) & (n_n491) & (n_n4503)) + ((i_9_) & (!n_n455) & (n_n534) & (!n_n491) & (n_n4503)) + ((i_9_) & (!n_n455) & (n_n534) & (n_n491) & (n_n4503)) + ((i_9_) & (n_n455) & (!n_n534) & (!n_n491) & (n_n4503)) + ((i_9_) & (n_n455) & (!n_n534) & (n_n491) & (n_n4503)) + ((i_9_) & (n_n455) & (n_n534) & (!n_n491) & (n_n4503)) + ((i_9_) & (n_n455) & (n_n534) & (n_n491) & (!n_n4503)) + ((i_9_) & (n_n455) & (n_n534) & (n_n491) & (n_n4503)));
	assign x13036x = (((!n_n4522) & (!n_n4525) & (!n_n4499) & (n_n4505)) + ((!n_n4522) & (!n_n4525) & (n_n4499) & (!n_n4505)) + ((!n_n4522) & (!n_n4525) & (n_n4499) & (n_n4505)) + ((!n_n4522) & (n_n4525) & (!n_n4499) & (!n_n4505)) + ((!n_n4522) & (n_n4525) & (!n_n4499) & (n_n4505)) + ((!n_n4522) & (n_n4525) & (n_n4499) & (!n_n4505)) + ((!n_n4522) & (n_n4525) & (n_n4499) & (n_n4505)) + ((n_n4522) & (!n_n4525) & (!n_n4499) & (!n_n4505)) + ((n_n4522) & (!n_n4525) & (!n_n4499) & (n_n4505)) + ((n_n4522) & (!n_n4525) & (n_n4499) & (!n_n4505)) + ((n_n4522) & (!n_n4525) & (n_n4499) & (n_n4505)) + ((n_n4522) & (n_n4525) & (!n_n4499) & (!n_n4505)) + ((n_n4522) & (n_n4525) & (!n_n4499) & (n_n4505)) + ((n_n4522) & (n_n4525) & (n_n4499) & (!n_n4505)) + ((n_n4522) & (n_n4525) & (n_n4499) & (n_n4505)));
	assign x13037x = (((!n_n4518) & (!n_n4498) & (!x307x) & (x13027x)) + ((!n_n4518) & (!n_n4498) & (x307x) & (!x13027x)) + ((!n_n4518) & (!n_n4498) & (x307x) & (x13027x)) + ((!n_n4518) & (n_n4498) & (!x307x) & (!x13027x)) + ((!n_n4518) & (n_n4498) & (!x307x) & (x13027x)) + ((!n_n4518) & (n_n4498) & (x307x) & (!x13027x)) + ((!n_n4518) & (n_n4498) & (x307x) & (x13027x)) + ((n_n4518) & (!n_n4498) & (!x307x) & (!x13027x)) + ((n_n4518) & (!n_n4498) & (!x307x) & (x13027x)) + ((n_n4518) & (!n_n4498) & (x307x) & (!x13027x)) + ((n_n4518) & (!n_n4498) & (x307x) & (x13027x)) + ((n_n4518) & (n_n4498) & (!x307x) & (!x13027x)) + ((n_n4518) & (n_n4498) & (!x307x) & (x13027x)) + ((n_n4518) & (n_n4498) & (x307x) & (!x13027x)) + ((n_n4518) & (n_n4498) & (x307x) & (x13027x)));
	assign x13038x = (((!n_n4521) & (!n_n4524) & (!x378x) & (!x162x) & (x346x)) + ((!n_n4521) & (!n_n4524) & (!x378x) & (x162x) & (!x346x)) + ((!n_n4521) & (!n_n4524) & (!x378x) & (x162x) & (x346x)) + ((!n_n4521) & (!n_n4524) & (x378x) & (!x162x) & (!x346x)) + ((!n_n4521) & (!n_n4524) & (x378x) & (!x162x) & (x346x)) + ((!n_n4521) & (!n_n4524) & (x378x) & (x162x) & (!x346x)) + ((!n_n4521) & (!n_n4524) & (x378x) & (x162x) & (x346x)) + ((!n_n4521) & (n_n4524) & (!x378x) & (!x162x) & (!x346x)) + ((!n_n4521) & (n_n4524) & (!x378x) & (!x162x) & (x346x)) + ((!n_n4521) & (n_n4524) & (!x378x) & (x162x) & (!x346x)) + ((!n_n4521) & (n_n4524) & (!x378x) & (x162x) & (x346x)) + ((!n_n4521) & (n_n4524) & (x378x) & (!x162x) & (!x346x)) + ((!n_n4521) & (n_n4524) & (x378x) & (!x162x) & (x346x)) + ((!n_n4521) & (n_n4524) & (x378x) & (x162x) & (!x346x)) + ((!n_n4521) & (n_n4524) & (x378x) & (x162x) & (x346x)) + ((n_n4521) & (!n_n4524) & (!x378x) & (!x162x) & (!x346x)) + ((n_n4521) & (!n_n4524) & (!x378x) & (!x162x) & (x346x)) + ((n_n4521) & (!n_n4524) & (!x378x) & (x162x) & (!x346x)) + ((n_n4521) & (!n_n4524) & (!x378x) & (x162x) & (x346x)) + ((n_n4521) & (!n_n4524) & (x378x) & (!x162x) & (!x346x)) + ((n_n4521) & (!n_n4524) & (x378x) & (!x162x) & (x346x)) + ((n_n4521) & (!n_n4524) & (x378x) & (x162x) & (!x346x)) + ((n_n4521) & (!n_n4524) & (x378x) & (x162x) & (x346x)) + ((n_n4521) & (n_n4524) & (!x378x) & (!x162x) & (!x346x)) + ((n_n4521) & (n_n4524) & (!x378x) & (!x162x) & (x346x)) + ((n_n4521) & (n_n4524) & (!x378x) & (x162x) & (!x346x)) + ((n_n4521) & (n_n4524) & (!x378x) & (x162x) & (x346x)) + ((n_n4521) & (n_n4524) & (x378x) & (!x162x) & (!x346x)) + ((n_n4521) & (n_n4524) & (x378x) & (!x162x) & (x346x)) + ((n_n4521) & (n_n4524) & (x378x) & (x162x) & (!x346x)) + ((n_n4521) & (n_n4524) & (x378x) & (x162x) & (x346x)));
	assign n_n653 = (((!n_n722) & (!x13036x) & (!x13037x) & (x13038x)) + ((!n_n722) & (!x13036x) & (x13037x) & (!x13038x)) + ((!n_n722) & (!x13036x) & (x13037x) & (x13038x)) + ((!n_n722) & (x13036x) & (!x13037x) & (!x13038x)) + ((!n_n722) & (x13036x) & (!x13037x) & (x13038x)) + ((!n_n722) & (x13036x) & (x13037x) & (!x13038x)) + ((!n_n722) & (x13036x) & (x13037x) & (x13038x)) + ((n_n722) & (!x13036x) & (!x13037x) & (!x13038x)) + ((n_n722) & (!x13036x) & (!x13037x) & (x13038x)) + ((n_n722) & (!x13036x) & (x13037x) & (!x13038x)) + ((n_n722) & (!x13036x) & (x13037x) & (x13038x)) + ((n_n722) & (x13036x) & (!x13037x) & (!x13038x)) + ((n_n722) & (x13036x) & (!x13037x) & (x13038x)) + ((n_n722) & (x13036x) & (x13037x) & (!x13038x)) + ((n_n722) & (x13036x) & (x13037x) & (x13038x)));
	assign x13044x = (((!x412x) & (!n_n4469) & (!n_n4462) & (!x322x) & (n_n2058)) + ((!x412x) & (!n_n4469) & (!n_n4462) & (x322x) & (!n_n2058)) + ((!x412x) & (!n_n4469) & (!n_n4462) & (x322x) & (n_n2058)) + ((!x412x) & (!n_n4469) & (n_n4462) & (!x322x) & (!n_n2058)) + ((!x412x) & (!n_n4469) & (n_n4462) & (!x322x) & (n_n2058)) + ((!x412x) & (!n_n4469) & (n_n4462) & (x322x) & (!n_n2058)) + ((!x412x) & (!n_n4469) & (n_n4462) & (x322x) & (n_n2058)) + ((!x412x) & (n_n4469) & (!n_n4462) & (!x322x) & (!n_n2058)) + ((!x412x) & (n_n4469) & (!n_n4462) & (!x322x) & (n_n2058)) + ((!x412x) & (n_n4469) & (!n_n4462) & (x322x) & (!n_n2058)) + ((!x412x) & (n_n4469) & (!n_n4462) & (x322x) & (n_n2058)) + ((!x412x) & (n_n4469) & (n_n4462) & (!x322x) & (!n_n2058)) + ((!x412x) & (n_n4469) & (n_n4462) & (!x322x) & (n_n2058)) + ((!x412x) & (n_n4469) & (n_n4462) & (x322x) & (!n_n2058)) + ((!x412x) & (n_n4469) & (n_n4462) & (x322x) & (n_n2058)) + ((x412x) & (!n_n4469) & (!n_n4462) & (!x322x) & (!n_n2058)) + ((x412x) & (!n_n4469) & (!n_n4462) & (!x322x) & (n_n2058)) + ((x412x) & (!n_n4469) & (!n_n4462) & (x322x) & (!n_n2058)) + ((x412x) & (!n_n4469) & (!n_n4462) & (x322x) & (n_n2058)) + ((x412x) & (!n_n4469) & (n_n4462) & (!x322x) & (!n_n2058)) + ((x412x) & (!n_n4469) & (n_n4462) & (!x322x) & (n_n2058)) + ((x412x) & (!n_n4469) & (n_n4462) & (x322x) & (!n_n2058)) + ((x412x) & (!n_n4469) & (n_n4462) & (x322x) & (n_n2058)) + ((x412x) & (n_n4469) & (!n_n4462) & (!x322x) & (!n_n2058)) + ((x412x) & (n_n4469) & (!n_n4462) & (!x322x) & (n_n2058)) + ((x412x) & (n_n4469) & (!n_n4462) & (x322x) & (!n_n2058)) + ((x412x) & (n_n4469) & (!n_n4462) & (x322x) & (n_n2058)) + ((x412x) & (n_n4469) & (n_n4462) & (!x322x) & (!n_n2058)) + ((x412x) & (n_n4469) & (n_n4462) & (!x322x) & (n_n2058)) + ((x412x) & (n_n4469) & (n_n4462) & (x322x) & (!n_n2058)) + ((x412x) & (n_n4469) & (n_n4462) & (x322x) & (n_n2058)));
	assign x13046x = (((!n_n725) & (!x13025x) & (!x13026x) & (x13044x)) + ((!n_n725) & (!x13025x) & (x13026x) & (!x13044x)) + ((!n_n725) & (!x13025x) & (x13026x) & (x13044x)) + ((!n_n725) & (x13025x) & (!x13026x) & (!x13044x)) + ((!n_n725) & (x13025x) & (!x13026x) & (x13044x)) + ((!n_n725) & (x13025x) & (x13026x) & (!x13044x)) + ((!n_n725) & (x13025x) & (x13026x) & (x13044x)) + ((n_n725) & (!x13025x) & (!x13026x) & (!x13044x)) + ((n_n725) & (!x13025x) & (!x13026x) & (x13044x)) + ((n_n725) & (!x13025x) & (x13026x) & (!x13044x)) + ((n_n725) & (!x13025x) & (x13026x) & (x13044x)) + ((n_n725) & (x13025x) & (!x13026x) & (!x13044x)) + ((n_n725) & (x13025x) & (!x13026x) & (x13044x)) + ((n_n725) & (x13025x) & (x13026x) & (!x13044x)) + ((n_n725) & (x13025x) & (x13026x) & (x13044x)));
	assign x13015x = (((!x233x) & (!x234x) & (!n_n4430) & (!n_n4426) & (x37x)) + ((!x233x) & (!x234x) & (!n_n4430) & (n_n4426) & (!x37x)) + ((!x233x) & (!x234x) & (!n_n4430) & (n_n4426) & (x37x)) + ((!x233x) & (!x234x) & (n_n4430) & (!n_n4426) & (!x37x)) + ((!x233x) & (!x234x) & (n_n4430) & (!n_n4426) & (x37x)) + ((!x233x) & (!x234x) & (n_n4430) & (n_n4426) & (!x37x)) + ((!x233x) & (!x234x) & (n_n4430) & (n_n4426) & (x37x)) + ((!x233x) & (x234x) & (!n_n4430) & (!n_n4426) & (!x37x)) + ((!x233x) & (x234x) & (!n_n4430) & (!n_n4426) & (x37x)) + ((!x233x) & (x234x) & (!n_n4430) & (n_n4426) & (!x37x)) + ((!x233x) & (x234x) & (!n_n4430) & (n_n4426) & (x37x)) + ((!x233x) & (x234x) & (n_n4430) & (!n_n4426) & (!x37x)) + ((!x233x) & (x234x) & (n_n4430) & (!n_n4426) & (x37x)) + ((!x233x) & (x234x) & (n_n4430) & (n_n4426) & (!x37x)) + ((!x233x) & (x234x) & (n_n4430) & (n_n4426) & (x37x)) + ((x233x) & (!x234x) & (!n_n4430) & (!n_n4426) & (!x37x)) + ((x233x) & (!x234x) & (!n_n4430) & (!n_n4426) & (x37x)) + ((x233x) & (!x234x) & (!n_n4430) & (n_n4426) & (!x37x)) + ((x233x) & (!x234x) & (!n_n4430) & (n_n4426) & (x37x)) + ((x233x) & (!x234x) & (n_n4430) & (!n_n4426) & (!x37x)) + ((x233x) & (!x234x) & (n_n4430) & (!n_n4426) & (x37x)) + ((x233x) & (!x234x) & (n_n4430) & (n_n4426) & (!x37x)) + ((x233x) & (!x234x) & (n_n4430) & (n_n4426) & (x37x)) + ((x233x) & (x234x) & (!n_n4430) & (!n_n4426) & (!x37x)) + ((x233x) & (x234x) & (!n_n4430) & (!n_n4426) & (x37x)) + ((x233x) & (x234x) & (!n_n4430) & (n_n4426) & (!x37x)) + ((x233x) & (x234x) & (!n_n4430) & (n_n4426) & (x37x)) + ((x233x) & (x234x) & (n_n4430) & (!n_n4426) & (!x37x)) + ((x233x) & (x234x) & (n_n4430) & (!n_n4426) & (x37x)) + ((x233x) & (x234x) & (n_n4430) & (n_n4426) & (!x37x)) + ((x233x) & (x234x) & (n_n4430) & (n_n4426) & (x37x)));
	assign x22173x = (((!n_n4927) & (!n_n4926) & (!n_n4925) & (!n_n4931)));
	assign n_n3691 = (((!n_n4934) & (!x31x) & (!n_n4935) & (!n_n4932) & (!x22173x)) + ((!n_n4934) & (!x31x) & (!n_n4935) & (n_n4932) & (!x22173x)) + ((!n_n4934) & (!x31x) & (!n_n4935) & (n_n4932) & (x22173x)) + ((!n_n4934) & (!x31x) & (n_n4935) & (!n_n4932) & (!x22173x)) + ((!n_n4934) & (!x31x) & (n_n4935) & (!n_n4932) & (x22173x)) + ((!n_n4934) & (!x31x) & (n_n4935) & (n_n4932) & (!x22173x)) + ((!n_n4934) & (!x31x) & (n_n4935) & (n_n4932) & (x22173x)) + ((!n_n4934) & (x31x) & (!n_n4935) & (!n_n4932) & (!x22173x)) + ((!n_n4934) & (x31x) & (!n_n4935) & (!n_n4932) & (x22173x)) + ((!n_n4934) & (x31x) & (!n_n4935) & (n_n4932) & (!x22173x)) + ((!n_n4934) & (x31x) & (!n_n4935) & (n_n4932) & (x22173x)) + ((!n_n4934) & (x31x) & (n_n4935) & (!n_n4932) & (!x22173x)) + ((!n_n4934) & (x31x) & (n_n4935) & (!n_n4932) & (x22173x)) + ((!n_n4934) & (x31x) & (n_n4935) & (n_n4932) & (!x22173x)) + ((!n_n4934) & (x31x) & (n_n4935) & (n_n4932) & (x22173x)) + ((n_n4934) & (!x31x) & (!n_n4935) & (!n_n4932) & (!x22173x)) + ((n_n4934) & (!x31x) & (!n_n4935) & (!n_n4932) & (x22173x)) + ((n_n4934) & (!x31x) & (!n_n4935) & (n_n4932) & (!x22173x)) + ((n_n4934) & (!x31x) & (!n_n4935) & (n_n4932) & (x22173x)) + ((n_n4934) & (!x31x) & (n_n4935) & (!n_n4932) & (!x22173x)) + ((n_n4934) & (!x31x) & (n_n4935) & (!n_n4932) & (x22173x)) + ((n_n4934) & (!x31x) & (n_n4935) & (n_n4932) & (!x22173x)) + ((n_n4934) & (!x31x) & (n_n4935) & (n_n4932) & (x22173x)) + ((n_n4934) & (x31x) & (!n_n4935) & (!n_n4932) & (!x22173x)) + ((n_n4934) & (x31x) & (!n_n4935) & (!n_n4932) & (x22173x)) + ((n_n4934) & (x31x) & (!n_n4935) & (n_n4932) & (!x22173x)) + ((n_n4934) & (x31x) & (!n_n4935) & (n_n4932) & (x22173x)) + ((n_n4934) & (x31x) & (n_n4935) & (!n_n4932) & (!x22173x)) + ((n_n4934) & (x31x) & (n_n4935) & (!n_n4932) & (x22173x)) + ((n_n4934) & (x31x) & (n_n4935) & (n_n4932) & (!x22173x)) + ((n_n4934) & (x31x) & (n_n4935) & (n_n4932) & (x22173x)));
	assign x14598x = (((!n_n522) & (!n_n491) & (!x12x) & (!n_n5157) & (x406x)) + ((!n_n522) & (!n_n491) & (!x12x) & (n_n5157) & (!x406x)) + ((!n_n522) & (!n_n491) & (!x12x) & (n_n5157) & (x406x)) + ((!n_n522) & (!n_n491) & (x12x) & (!n_n5157) & (x406x)) + ((!n_n522) & (!n_n491) & (x12x) & (n_n5157) & (!x406x)) + ((!n_n522) & (!n_n491) & (x12x) & (n_n5157) & (x406x)) + ((!n_n522) & (n_n491) & (!x12x) & (!n_n5157) & (x406x)) + ((!n_n522) & (n_n491) & (!x12x) & (n_n5157) & (!x406x)) + ((!n_n522) & (n_n491) & (!x12x) & (n_n5157) & (x406x)) + ((!n_n522) & (n_n491) & (x12x) & (!n_n5157) & (x406x)) + ((!n_n522) & (n_n491) & (x12x) & (n_n5157) & (!x406x)) + ((!n_n522) & (n_n491) & (x12x) & (n_n5157) & (x406x)) + ((n_n522) & (!n_n491) & (!x12x) & (!n_n5157) & (x406x)) + ((n_n522) & (!n_n491) & (!x12x) & (n_n5157) & (!x406x)) + ((n_n522) & (!n_n491) & (!x12x) & (n_n5157) & (x406x)) + ((n_n522) & (!n_n491) & (x12x) & (!n_n5157) & (x406x)) + ((n_n522) & (!n_n491) & (x12x) & (n_n5157) & (!x406x)) + ((n_n522) & (!n_n491) & (x12x) & (n_n5157) & (x406x)) + ((n_n522) & (n_n491) & (!x12x) & (!n_n5157) & (x406x)) + ((n_n522) & (n_n491) & (!x12x) & (n_n5157) & (!x406x)) + ((n_n522) & (n_n491) & (!x12x) & (n_n5157) & (x406x)) + ((n_n522) & (n_n491) & (x12x) & (!n_n5157) & (!x406x)) + ((n_n522) & (n_n491) & (x12x) & (!n_n5157) & (x406x)) + ((n_n522) & (n_n491) & (x12x) & (n_n5157) & (!x406x)) + ((n_n522) & (n_n491) & (x12x) & (n_n5157) & (x406x)));
	assign x22186x = (((!x19x) & (!n_n520) & (!n_n500) & (!x203x) & (!x438x)) + ((!x19x) & (!n_n520) & (n_n500) & (!x203x) & (!x438x)) + ((!x19x) & (n_n520) & (!n_n500) & (!x203x) & (!x438x)) + ((!x19x) & (n_n520) & (n_n500) & (!x203x) & (!x438x)) + ((x19x) & (!n_n520) & (!n_n500) & (!x203x) & (!x438x)) + ((x19x) & (!n_n520) & (n_n500) & (!x203x) & (!x438x)) + ((x19x) & (n_n520) & (!n_n500) & (!x203x) & (!x438x)));
	assign x15519x = (((!i_9_) & (n_n536) & (!n_n532) & (n_n535) & (x20x)) + ((!i_9_) & (n_n536) & (n_n532) & (n_n535) & (x20x)) + ((i_9_) & (n_n536) & (!n_n532) & (n_n535) & (x20x)) + ((i_9_) & (n_n536) & (n_n532) & (n_n535) & (!x20x)) + ((i_9_) & (n_n536) & (n_n532) & (n_n535) & (x20x)));
	assign n_n3012 = (((!n_n4317) & (!n_n4326) & (!n_n4328) & (!x363x) & (x15519x)) + ((!n_n4317) & (!n_n4326) & (!n_n4328) & (x363x) & (!x15519x)) + ((!n_n4317) & (!n_n4326) & (!n_n4328) & (x363x) & (x15519x)) + ((!n_n4317) & (!n_n4326) & (n_n4328) & (!x363x) & (!x15519x)) + ((!n_n4317) & (!n_n4326) & (n_n4328) & (!x363x) & (x15519x)) + ((!n_n4317) & (!n_n4326) & (n_n4328) & (x363x) & (!x15519x)) + ((!n_n4317) & (!n_n4326) & (n_n4328) & (x363x) & (x15519x)) + ((!n_n4317) & (n_n4326) & (!n_n4328) & (!x363x) & (!x15519x)) + ((!n_n4317) & (n_n4326) & (!n_n4328) & (!x363x) & (x15519x)) + ((!n_n4317) & (n_n4326) & (!n_n4328) & (x363x) & (!x15519x)) + ((!n_n4317) & (n_n4326) & (!n_n4328) & (x363x) & (x15519x)) + ((!n_n4317) & (n_n4326) & (n_n4328) & (!x363x) & (!x15519x)) + ((!n_n4317) & (n_n4326) & (n_n4328) & (!x363x) & (x15519x)) + ((!n_n4317) & (n_n4326) & (n_n4328) & (x363x) & (!x15519x)) + ((!n_n4317) & (n_n4326) & (n_n4328) & (x363x) & (x15519x)) + ((n_n4317) & (!n_n4326) & (!n_n4328) & (!x363x) & (!x15519x)) + ((n_n4317) & (!n_n4326) & (!n_n4328) & (!x363x) & (x15519x)) + ((n_n4317) & (!n_n4326) & (!n_n4328) & (x363x) & (!x15519x)) + ((n_n4317) & (!n_n4326) & (!n_n4328) & (x363x) & (x15519x)) + ((n_n4317) & (!n_n4326) & (n_n4328) & (!x363x) & (!x15519x)) + ((n_n4317) & (!n_n4326) & (n_n4328) & (!x363x) & (x15519x)) + ((n_n4317) & (!n_n4326) & (n_n4328) & (x363x) & (!x15519x)) + ((n_n4317) & (!n_n4326) & (n_n4328) & (x363x) & (x15519x)) + ((n_n4317) & (n_n4326) & (!n_n4328) & (!x363x) & (!x15519x)) + ((n_n4317) & (n_n4326) & (!n_n4328) & (!x363x) & (x15519x)) + ((n_n4317) & (n_n4326) & (!n_n4328) & (x363x) & (!x15519x)) + ((n_n4317) & (n_n4326) & (!n_n4328) & (x363x) & (x15519x)) + ((n_n4317) & (n_n4326) & (n_n4328) & (!x363x) & (!x15519x)) + ((n_n4317) & (n_n4326) & (n_n4328) & (!x363x) & (x15519x)) + ((n_n4317) & (n_n4326) & (n_n4328) & (x363x) & (!x15519x)) + ((n_n4317) & (n_n4326) & (n_n4328) & (x363x) & (x15519x)));
	assign x22213x = (((!x25x) & (!n_n536) & (!n_n518) & (!x24x) & (!n_n4336)) + ((!x25x) & (!n_n536) & (!n_n518) & (x24x) & (!n_n4336)) + ((!x25x) & (!n_n536) & (n_n518) & (!x24x) & (!n_n4336)) + ((!x25x) & (!n_n536) & (n_n518) & (x24x) & (!n_n4336)) + ((!x25x) & (n_n536) & (!n_n518) & (!x24x) & (!n_n4336)) + ((!x25x) & (n_n536) & (!n_n518) & (x24x) & (!n_n4336)) + ((!x25x) & (n_n536) & (n_n518) & (!x24x) & (!n_n4336)) + ((x25x) & (!n_n536) & (!n_n518) & (!x24x) & (!n_n4336)) + ((x25x) & (!n_n536) & (!n_n518) & (x24x) & (!n_n4336)) + ((x25x) & (!n_n536) & (n_n518) & (!x24x) & (!n_n4336)) + ((x25x) & (!n_n536) & (n_n518) & (x24x) & (!n_n4336)) + ((x25x) & (n_n536) & (!n_n518) & (!x24x) & (!n_n4336)) + ((x25x) & (n_n536) & (!n_n518) & (x24x) & (!n_n4336)));
	assign x15527x = (((!n_n4337) & (!n_n4332) & (!x53x) & (!x443x) & (!x22213x)) + ((!n_n4337) & (!n_n4332) & (!x53x) & (x443x) & (!x22213x)) + ((!n_n4337) & (!n_n4332) & (!x53x) & (x443x) & (x22213x)) + ((!n_n4337) & (!n_n4332) & (x53x) & (!x443x) & (!x22213x)) + ((!n_n4337) & (!n_n4332) & (x53x) & (!x443x) & (x22213x)) + ((!n_n4337) & (!n_n4332) & (x53x) & (x443x) & (!x22213x)) + ((!n_n4337) & (!n_n4332) & (x53x) & (x443x) & (x22213x)) + ((!n_n4337) & (n_n4332) & (!x53x) & (!x443x) & (!x22213x)) + ((!n_n4337) & (n_n4332) & (!x53x) & (!x443x) & (x22213x)) + ((!n_n4337) & (n_n4332) & (!x53x) & (x443x) & (!x22213x)) + ((!n_n4337) & (n_n4332) & (!x53x) & (x443x) & (x22213x)) + ((!n_n4337) & (n_n4332) & (x53x) & (!x443x) & (!x22213x)) + ((!n_n4337) & (n_n4332) & (x53x) & (!x443x) & (x22213x)) + ((!n_n4337) & (n_n4332) & (x53x) & (x443x) & (!x22213x)) + ((!n_n4337) & (n_n4332) & (x53x) & (x443x) & (x22213x)) + ((n_n4337) & (!n_n4332) & (!x53x) & (!x443x) & (!x22213x)) + ((n_n4337) & (!n_n4332) & (!x53x) & (!x443x) & (x22213x)) + ((n_n4337) & (!n_n4332) & (!x53x) & (x443x) & (!x22213x)) + ((n_n4337) & (!n_n4332) & (!x53x) & (x443x) & (x22213x)) + ((n_n4337) & (!n_n4332) & (x53x) & (!x443x) & (!x22213x)) + ((n_n4337) & (!n_n4332) & (x53x) & (!x443x) & (x22213x)) + ((n_n4337) & (!n_n4332) & (x53x) & (x443x) & (!x22213x)) + ((n_n4337) & (!n_n4332) & (x53x) & (x443x) & (x22213x)) + ((n_n4337) & (n_n4332) & (!x53x) & (!x443x) & (!x22213x)) + ((n_n4337) & (n_n4332) & (!x53x) & (!x443x) & (x22213x)) + ((n_n4337) & (n_n4332) & (!x53x) & (x443x) & (!x22213x)) + ((n_n4337) & (n_n4332) & (!x53x) & (x443x) & (x22213x)) + ((n_n4337) & (n_n4332) & (x53x) & (!x443x) & (!x22213x)) + ((n_n4337) & (n_n4332) & (x53x) & (!x443x) & (x22213x)) + ((n_n4337) & (n_n4332) & (x53x) & (x443x) & (!x22213x)) + ((n_n4337) & (n_n4332) & (x53x) & (x443x) & (x22213x)));
	assign x15771x = (((!n_n4674) & (!n_n4683) & (!n_n4681) & (!n_n4678) & (n_n4684)) + ((!n_n4674) & (!n_n4683) & (!n_n4681) & (n_n4678) & (!n_n4684)) + ((!n_n4674) & (!n_n4683) & (!n_n4681) & (n_n4678) & (n_n4684)) + ((!n_n4674) & (!n_n4683) & (n_n4681) & (!n_n4678) & (!n_n4684)) + ((!n_n4674) & (!n_n4683) & (n_n4681) & (!n_n4678) & (n_n4684)) + ((!n_n4674) & (!n_n4683) & (n_n4681) & (n_n4678) & (!n_n4684)) + ((!n_n4674) & (!n_n4683) & (n_n4681) & (n_n4678) & (n_n4684)) + ((!n_n4674) & (n_n4683) & (!n_n4681) & (!n_n4678) & (!n_n4684)) + ((!n_n4674) & (n_n4683) & (!n_n4681) & (!n_n4678) & (n_n4684)) + ((!n_n4674) & (n_n4683) & (!n_n4681) & (n_n4678) & (!n_n4684)) + ((!n_n4674) & (n_n4683) & (!n_n4681) & (n_n4678) & (n_n4684)) + ((!n_n4674) & (n_n4683) & (n_n4681) & (!n_n4678) & (!n_n4684)) + ((!n_n4674) & (n_n4683) & (n_n4681) & (!n_n4678) & (n_n4684)) + ((!n_n4674) & (n_n4683) & (n_n4681) & (n_n4678) & (!n_n4684)) + ((!n_n4674) & (n_n4683) & (n_n4681) & (n_n4678) & (n_n4684)) + ((n_n4674) & (!n_n4683) & (!n_n4681) & (!n_n4678) & (!n_n4684)) + ((n_n4674) & (!n_n4683) & (!n_n4681) & (!n_n4678) & (n_n4684)) + ((n_n4674) & (!n_n4683) & (!n_n4681) & (n_n4678) & (!n_n4684)) + ((n_n4674) & (!n_n4683) & (!n_n4681) & (n_n4678) & (n_n4684)) + ((n_n4674) & (!n_n4683) & (n_n4681) & (!n_n4678) & (!n_n4684)) + ((n_n4674) & (!n_n4683) & (n_n4681) & (!n_n4678) & (n_n4684)) + ((n_n4674) & (!n_n4683) & (n_n4681) & (n_n4678) & (!n_n4684)) + ((n_n4674) & (!n_n4683) & (n_n4681) & (n_n4678) & (n_n4684)) + ((n_n4674) & (n_n4683) & (!n_n4681) & (!n_n4678) & (!n_n4684)) + ((n_n4674) & (n_n4683) & (!n_n4681) & (!n_n4678) & (n_n4684)) + ((n_n4674) & (n_n4683) & (!n_n4681) & (n_n4678) & (!n_n4684)) + ((n_n4674) & (n_n4683) & (!n_n4681) & (n_n4678) & (n_n4684)) + ((n_n4674) & (n_n4683) & (n_n4681) & (!n_n4678) & (!n_n4684)) + ((n_n4674) & (n_n4683) & (n_n4681) & (!n_n4678) & (n_n4684)) + ((n_n4674) & (n_n4683) & (n_n4681) & (n_n4678) & (!n_n4684)) + ((n_n4674) & (n_n4683) & (n_n4681) & (n_n4678) & (n_n4684)));
	assign x15778x = (((!n_n3125) & (!n_n4219) & (!x30x) & (n_n3124)) + ((!n_n3125) & (!n_n4219) & (x30x) & (!n_n3124)) + ((!n_n3125) & (!n_n4219) & (x30x) & (n_n3124)) + ((!n_n3125) & (n_n4219) & (!x30x) & (!n_n3124)) + ((!n_n3125) & (n_n4219) & (!x30x) & (n_n3124)) + ((!n_n3125) & (n_n4219) & (x30x) & (!n_n3124)) + ((!n_n3125) & (n_n4219) & (x30x) & (n_n3124)) + ((n_n3125) & (!n_n4219) & (!x30x) & (!n_n3124)) + ((n_n3125) & (!n_n4219) & (!x30x) & (n_n3124)) + ((n_n3125) & (!n_n4219) & (x30x) & (!n_n3124)) + ((n_n3125) & (!n_n4219) & (x30x) & (n_n3124)) + ((n_n3125) & (n_n4219) & (!x30x) & (!n_n3124)) + ((n_n3125) & (n_n4219) & (!x30x) & (n_n3124)) + ((n_n3125) & (n_n4219) & (x30x) & (!n_n3124)) + ((n_n3125) & (n_n4219) & (x30x) & (n_n3124)));
	assign x15777x = (((!x10x) & (!x516x) & (!n_n4688) & (!n_n4693) & (x15775x)) + ((!x10x) & (!x516x) & (!n_n4688) & (n_n4693) & (!x15775x)) + ((!x10x) & (!x516x) & (!n_n4688) & (n_n4693) & (x15775x)) + ((!x10x) & (!x516x) & (n_n4688) & (!n_n4693) & (!x15775x)) + ((!x10x) & (!x516x) & (n_n4688) & (!n_n4693) & (x15775x)) + ((!x10x) & (!x516x) & (n_n4688) & (n_n4693) & (!x15775x)) + ((!x10x) & (!x516x) & (n_n4688) & (n_n4693) & (x15775x)) + ((!x10x) & (x516x) & (!n_n4688) & (!n_n4693) & (x15775x)) + ((!x10x) & (x516x) & (!n_n4688) & (n_n4693) & (!x15775x)) + ((!x10x) & (x516x) & (!n_n4688) & (n_n4693) & (x15775x)) + ((!x10x) & (x516x) & (n_n4688) & (!n_n4693) & (!x15775x)) + ((!x10x) & (x516x) & (n_n4688) & (!n_n4693) & (x15775x)) + ((!x10x) & (x516x) & (n_n4688) & (n_n4693) & (!x15775x)) + ((!x10x) & (x516x) & (n_n4688) & (n_n4693) & (x15775x)) + ((x10x) & (!x516x) & (!n_n4688) & (!n_n4693) & (x15775x)) + ((x10x) & (!x516x) & (!n_n4688) & (n_n4693) & (!x15775x)) + ((x10x) & (!x516x) & (!n_n4688) & (n_n4693) & (x15775x)) + ((x10x) & (!x516x) & (n_n4688) & (!n_n4693) & (!x15775x)) + ((x10x) & (!x516x) & (n_n4688) & (!n_n4693) & (x15775x)) + ((x10x) & (!x516x) & (n_n4688) & (n_n4693) & (!x15775x)) + ((x10x) & (!x516x) & (n_n4688) & (n_n4693) & (x15775x)) + ((x10x) & (x516x) & (!n_n4688) & (!n_n4693) & (!x15775x)) + ((x10x) & (x516x) & (!n_n4688) & (!n_n4693) & (x15775x)) + ((x10x) & (x516x) & (!n_n4688) & (n_n4693) & (!x15775x)) + ((x10x) & (x516x) & (!n_n4688) & (n_n4693) & (x15775x)) + ((x10x) & (x516x) & (n_n4688) & (!n_n4693) & (!x15775x)) + ((x10x) & (x516x) & (n_n4688) & (!n_n4693) & (x15775x)) + ((x10x) & (x516x) & (n_n4688) & (n_n4693) & (!x15775x)) + ((x10x) & (x516x) & (n_n4688) & (n_n4693) & (x15775x)));
	assign n_n2925 = (((!x193x) & (!x80x) & (!x15771x) & (!x15778x) & (x15777x)) + ((!x193x) & (!x80x) & (!x15771x) & (x15778x) & (!x15777x)) + ((!x193x) & (!x80x) & (!x15771x) & (x15778x) & (x15777x)) + ((!x193x) & (!x80x) & (x15771x) & (!x15778x) & (!x15777x)) + ((!x193x) & (!x80x) & (x15771x) & (!x15778x) & (x15777x)) + ((!x193x) & (!x80x) & (x15771x) & (x15778x) & (!x15777x)) + ((!x193x) & (!x80x) & (x15771x) & (x15778x) & (x15777x)) + ((!x193x) & (x80x) & (!x15771x) & (!x15778x) & (!x15777x)) + ((!x193x) & (x80x) & (!x15771x) & (!x15778x) & (x15777x)) + ((!x193x) & (x80x) & (!x15771x) & (x15778x) & (!x15777x)) + ((!x193x) & (x80x) & (!x15771x) & (x15778x) & (x15777x)) + ((!x193x) & (x80x) & (x15771x) & (!x15778x) & (!x15777x)) + ((!x193x) & (x80x) & (x15771x) & (!x15778x) & (x15777x)) + ((!x193x) & (x80x) & (x15771x) & (x15778x) & (!x15777x)) + ((!x193x) & (x80x) & (x15771x) & (x15778x) & (x15777x)) + ((x193x) & (!x80x) & (!x15771x) & (!x15778x) & (!x15777x)) + ((x193x) & (!x80x) & (!x15771x) & (!x15778x) & (x15777x)) + ((x193x) & (!x80x) & (!x15771x) & (x15778x) & (!x15777x)) + ((x193x) & (!x80x) & (!x15771x) & (x15778x) & (x15777x)) + ((x193x) & (!x80x) & (x15771x) & (!x15778x) & (!x15777x)) + ((x193x) & (!x80x) & (x15771x) & (!x15778x) & (x15777x)) + ((x193x) & (!x80x) & (x15771x) & (x15778x) & (!x15777x)) + ((x193x) & (!x80x) & (x15771x) & (x15778x) & (x15777x)) + ((x193x) & (x80x) & (!x15771x) & (!x15778x) & (!x15777x)) + ((x193x) & (x80x) & (!x15771x) & (!x15778x) & (x15777x)) + ((x193x) & (x80x) & (!x15771x) & (x15778x) & (!x15777x)) + ((x193x) & (x80x) & (!x15771x) & (x15778x) & (x15777x)) + ((x193x) & (x80x) & (x15771x) & (!x15778x) & (!x15777x)) + ((x193x) & (x80x) & (x15771x) & (!x15778x) & (x15777x)) + ((x193x) & (x80x) & (x15771x) & (x15778x) & (!x15777x)) + ((x193x) & (x80x) & (x15771x) & (x15778x) & (x15777x)));
	assign x15413x = (((!n_n4863) & (!n_n4865) & (!n_n4852) & (!n_n4872) & (n_n4826)) + ((!n_n4863) & (!n_n4865) & (!n_n4852) & (n_n4872) & (!n_n4826)) + ((!n_n4863) & (!n_n4865) & (!n_n4852) & (n_n4872) & (n_n4826)) + ((!n_n4863) & (!n_n4865) & (n_n4852) & (!n_n4872) & (!n_n4826)) + ((!n_n4863) & (!n_n4865) & (n_n4852) & (!n_n4872) & (n_n4826)) + ((!n_n4863) & (!n_n4865) & (n_n4852) & (n_n4872) & (!n_n4826)) + ((!n_n4863) & (!n_n4865) & (n_n4852) & (n_n4872) & (n_n4826)) + ((!n_n4863) & (n_n4865) & (!n_n4852) & (!n_n4872) & (!n_n4826)) + ((!n_n4863) & (n_n4865) & (!n_n4852) & (!n_n4872) & (n_n4826)) + ((!n_n4863) & (n_n4865) & (!n_n4852) & (n_n4872) & (!n_n4826)) + ((!n_n4863) & (n_n4865) & (!n_n4852) & (n_n4872) & (n_n4826)) + ((!n_n4863) & (n_n4865) & (n_n4852) & (!n_n4872) & (!n_n4826)) + ((!n_n4863) & (n_n4865) & (n_n4852) & (!n_n4872) & (n_n4826)) + ((!n_n4863) & (n_n4865) & (n_n4852) & (n_n4872) & (!n_n4826)) + ((!n_n4863) & (n_n4865) & (n_n4852) & (n_n4872) & (n_n4826)) + ((n_n4863) & (!n_n4865) & (!n_n4852) & (!n_n4872) & (!n_n4826)) + ((n_n4863) & (!n_n4865) & (!n_n4852) & (!n_n4872) & (n_n4826)) + ((n_n4863) & (!n_n4865) & (!n_n4852) & (n_n4872) & (!n_n4826)) + ((n_n4863) & (!n_n4865) & (!n_n4852) & (n_n4872) & (n_n4826)) + ((n_n4863) & (!n_n4865) & (n_n4852) & (!n_n4872) & (!n_n4826)) + ((n_n4863) & (!n_n4865) & (n_n4852) & (!n_n4872) & (n_n4826)) + ((n_n4863) & (!n_n4865) & (n_n4852) & (n_n4872) & (!n_n4826)) + ((n_n4863) & (!n_n4865) & (n_n4852) & (n_n4872) & (n_n4826)) + ((n_n4863) & (n_n4865) & (!n_n4852) & (!n_n4872) & (!n_n4826)) + ((n_n4863) & (n_n4865) & (!n_n4852) & (!n_n4872) & (n_n4826)) + ((n_n4863) & (n_n4865) & (!n_n4852) & (n_n4872) & (!n_n4826)) + ((n_n4863) & (n_n4865) & (!n_n4852) & (n_n4872) & (n_n4826)) + ((n_n4863) & (n_n4865) & (n_n4852) & (!n_n4872) & (!n_n4826)) + ((n_n4863) & (n_n4865) & (n_n4852) & (!n_n4872) & (n_n4826)) + ((n_n4863) & (n_n4865) & (n_n4852) & (n_n4872) & (!n_n4826)) + ((n_n4863) & (n_n4865) & (n_n4852) & (n_n4872) & (n_n4826)));
	assign x15367x = (((!n_n5092) & (!n_n5069) & (!n_n5084) & (n_n5078)) + ((!n_n5092) & (!n_n5069) & (n_n5084) & (!n_n5078)) + ((!n_n5092) & (!n_n5069) & (n_n5084) & (n_n5078)) + ((!n_n5092) & (n_n5069) & (!n_n5084) & (!n_n5078)) + ((!n_n5092) & (n_n5069) & (!n_n5084) & (n_n5078)) + ((!n_n5092) & (n_n5069) & (n_n5084) & (!n_n5078)) + ((!n_n5092) & (n_n5069) & (n_n5084) & (n_n5078)) + ((n_n5092) & (!n_n5069) & (!n_n5084) & (!n_n5078)) + ((n_n5092) & (!n_n5069) & (!n_n5084) & (n_n5078)) + ((n_n5092) & (!n_n5069) & (n_n5084) & (!n_n5078)) + ((n_n5092) & (!n_n5069) & (n_n5084) & (n_n5078)) + ((n_n5092) & (n_n5069) & (!n_n5084) & (!n_n5078)) + ((n_n5092) & (n_n5069) & (!n_n5084) & (n_n5078)) + ((n_n5092) & (n_n5069) & (n_n5084) & (!n_n5078)) + ((n_n5092) & (n_n5069) & (n_n5084) & (n_n5078)));
	assign x15355x = (((!n_n5161) & (!n_n5120) & (!n_n5135) & (n_n5147)) + ((!n_n5161) & (!n_n5120) & (n_n5135) & (!n_n5147)) + ((!n_n5161) & (!n_n5120) & (n_n5135) & (n_n5147)) + ((!n_n5161) & (n_n5120) & (!n_n5135) & (!n_n5147)) + ((!n_n5161) & (n_n5120) & (!n_n5135) & (n_n5147)) + ((!n_n5161) & (n_n5120) & (n_n5135) & (!n_n5147)) + ((!n_n5161) & (n_n5120) & (n_n5135) & (n_n5147)) + ((n_n5161) & (!n_n5120) & (!n_n5135) & (!n_n5147)) + ((n_n5161) & (!n_n5120) & (!n_n5135) & (n_n5147)) + ((n_n5161) & (!n_n5120) & (n_n5135) & (!n_n5147)) + ((n_n5161) & (!n_n5120) & (n_n5135) & (n_n5147)) + ((n_n5161) & (n_n5120) & (!n_n5135) & (!n_n5147)) + ((n_n5161) & (n_n5120) & (!n_n5135) & (n_n5147)) + ((n_n5161) & (n_n5120) & (n_n5135) & (!n_n5147)) + ((n_n5161) & (n_n5120) & (n_n5135) & (n_n5147)));
	assign x15356x = (((!n_n5111) & (!n_n5113) & (!n_n5140) & (!n_n5144) & (n_n5143)) + ((!n_n5111) & (!n_n5113) & (!n_n5140) & (n_n5144) & (!n_n5143)) + ((!n_n5111) & (!n_n5113) & (!n_n5140) & (n_n5144) & (n_n5143)) + ((!n_n5111) & (!n_n5113) & (n_n5140) & (!n_n5144) & (!n_n5143)) + ((!n_n5111) & (!n_n5113) & (n_n5140) & (!n_n5144) & (n_n5143)) + ((!n_n5111) & (!n_n5113) & (n_n5140) & (n_n5144) & (!n_n5143)) + ((!n_n5111) & (!n_n5113) & (n_n5140) & (n_n5144) & (n_n5143)) + ((!n_n5111) & (n_n5113) & (!n_n5140) & (!n_n5144) & (!n_n5143)) + ((!n_n5111) & (n_n5113) & (!n_n5140) & (!n_n5144) & (n_n5143)) + ((!n_n5111) & (n_n5113) & (!n_n5140) & (n_n5144) & (!n_n5143)) + ((!n_n5111) & (n_n5113) & (!n_n5140) & (n_n5144) & (n_n5143)) + ((!n_n5111) & (n_n5113) & (n_n5140) & (!n_n5144) & (!n_n5143)) + ((!n_n5111) & (n_n5113) & (n_n5140) & (!n_n5144) & (n_n5143)) + ((!n_n5111) & (n_n5113) & (n_n5140) & (n_n5144) & (!n_n5143)) + ((!n_n5111) & (n_n5113) & (n_n5140) & (n_n5144) & (n_n5143)) + ((n_n5111) & (!n_n5113) & (!n_n5140) & (!n_n5144) & (!n_n5143)) + ((n_n5111) & (!n_n5113) & (!n_n5140) & (!n_n5144) & (n_n5143)) + ((n_n5111) & (!n_n5113) & (!n_n5140) & (n_n5144) & (!n_n5143)) + ((n_n5111) & (!n_n5113) & (!n_n5140) & (n_n5144) & (n_n5143)) + ((n_n5111) & (!n_n5113) & (n_n5140) & (!n_n5144) & (!n_n5143)) + ((n_n5111) & (!n_n5113) & (n_n5140) & (!n_n5144) & (n_n5143)) + ((n_n5111) & (!n_n5113) & (n_n5140) & (n_n5144) & (!n_n5143)) + ((n_n5111) & (!n_n5113) & (n_n5140) & (n_n5144) & (n_n5143)) + ((n_n5111) & (n_n5113) & (!n_n5140) & (!n_n5144) & (!n_n5143)) + ((n_n5111) & (n_n5113) & (!n_n5140) & (!n_n5144) & (n_n5143)) + ((n_n5111) & (n_n5113) & (!n_n5140) & (n_n5144) & (!n_n5143)) + ((n_n5111) & (n_n5113) & (!n_n5140) & (n_n5144) & (n_n5143)) + ((n_n5111) & (n_n5113) & (n_n5140) & (!n_n5144) & (!n_n5143)) + ((n_n5111) & (n_n5113) & (n_n5140) & (!n_n5144) & (n_n5143)) + ((n_n5111) & (n_n5113) & (n_n5140) & (n_n5144) & (!n_n5143)) + ((n_n5111) & (n_n5113) & (n_n5140) & (n_n5144) & (n_n5143)));
	assign x15361x = (((!n_n4990) & (!n_n5027) & (!n_n5048) & (n_n5053)) + ((!n_n4990) & (!n_n5027) & (n_n5048) & (!n_n5053)) + ((!n_n4990) & (!n_n5027) & (n_n5048) & (n_n5053)) + ((!n_n4990) & (n_n5027) & (!n_n5048) & (!n_n5053)) + ((!n_n4990) & (n_n5027) & (!n_n5048) & (n_n5053)) + ((!n_n4990) & (n_n5027) & (n_n5048) & (!n_n5053)) + ((!n_n4990) & (n_n5027) & (n_n5048) & (n_n5053)) + ((n_n4990) & (!n_n5027) & (!n_n5048) & (!n_n5053)) + ((n_n4990) & (!n_n5027) & (!n_n5048) & (n_n5053)) + ((n_n4990) & (!n_n5027) & (n_n5048) & (!n_n5053)) + ((n_n4990) & (!n_n5027) & (n_n5048) & (n_n5053)) + ((n_n4990) & (n_n5027) & (!n_n5048) & (!n_n5053)) + ((n_n4990) & (n_n5027) & (!n_n5048) & (n_n5053)) + ((n_n4990) & (n_n5027) & (n_n5048) & (!n_n5053)) + ((n_n4990) & (n_n5027) & (n_n5048) & (n_n5053)));
	assign x15362x = (((!n_n5001) & (!x120x) & (!n_n4989) & (n_n5033)) + ((!n_n5001) & (!x120x) & (n_n4989) & (!n_n5033)) + ((!n_n5001) & (!x120x) & (n_n4989) & (n_n5033)) + ((!n_n5001) & (x120x) & (!n_n4989) & (!n_n5033)) + ((!n_n5001) & (x120x) & (!n_n4989) & (n_n5033)) + ((!n_n5001) & (x120x) & (n_n4989) & (!n_n5033)) + ((!n_n5001) & (x120x) & (n_n4989) & (n_n5033)) + ((n_n5001) & (!x120x) & (!n_n4989) & (!n_n5033)) + ((n_n5001) & (!x120x) & (!n_n4989) & (n_n5033)) + ((n_n5001) & (!x120x) & (n_n4989) & (!n_n5033)) + ((n_n5001) & (!x120x) & (n_n4989) & (n_n5033)) + ((n_n5001) & (x120x) & (!n_n4989) & (!n_n5033)) + ((n_n5001) & (x120x) & (!n_n4989) & (n_n5033)) + ((n_n5001) & (x120x) & (n_n4989) & (!n_n5033)) + ((n_n5001) & (x120x) & (n_n4989) & (n_n5033)));
	assign x15374x = (((!n_n5171) & (!n_n5230) & (!n_n5168) & (n_n5170)) + ((!n_n5171) & (!n_n5230) & (n_n5168) & (!n_n5170)) + ((!n_n5171) & (!n_n5230) & (n_n5168) & (n_n5170)) + ((!n_n5171) & (n_n5230) & (!n_n5168) & (!n_n5170)) + ((!n_n5171) & (n_n5230) & (!n_n5168) & (n_n5170)) + ((!n_n5171) & (n_n5230) & (n_n5168) & (!n_n5170)) + ((!n_n5171) & (n_n5230) & (n_n5168) & (n_n5170)) + ((n_n5171) & (!n_n5230) & (!n_n5168) & (!n_n5170)) + ((n_n5171) & (!n_n5230) & (!n_n5168) & (n_n5170)) + ((n_n5171) & (!n_n5230) & (n_n5168) & (!n_n5170)) + ((n_n5171) & (!n_n5230) & (n_n5168) & (n_n5170)) + ((n_n5171) & (n_n5230) & (!n_n5168) & (!n_n5170)) + ((n_n5171) & (n_n5230) & (!n_n5168) & (n_n5170)) + ((n_n5171) & (n_n5230) & (n_n5168) & (!n_n5170)) + ((n_n5171) & (n_n5230) & (n_n5168) & (n_n5170)));
	assign x15375x = (((!n_n5217) & (!n_n5169) & (!x33x) & (n_n5235)) + ((!n_n5217) & (!n_n5169) & (x33x) & (!n_n5235)) + ((!n_n5217) & (!n_n5169) & (x33x) & (n_n5235)) + ((!n_n5217) & (n_n5169) & (!x33x) & (!n_n5235)) + ((!n_n5217) & (n_n5169) & (!x33x) & (n_n5235)) + ((!n_n5217) & (n_n5169) & (x33x) & (!n_n5235)) + ((!n_n5217) & (n_n5169) & (x33x) & (n_n5235)) + ((n_n5217) & (!n_n5169) & (!x33x) & (!n_n5235)) + ((n_n5217) & (!n_n5169) & (!x33x) & (n_n5235)) + ((n_n5217) & (!n_n5169) & (x33x) & (!n_n5235)) + ((n_n5217) & (!n_n5169) & (x33x) & (n_n5235)) + ((n_n5217) & (n_n5169) & (!x33x) & (!n_n5235)) + ((n_n5217) & (n_n5169) & (!x33x) & (n_n5235)) + ((n_n5217) & (n_n5169) & (x33x) & (!n_n5235)) + ((n_n5217) & (n_n5169) & (x33x) & (n_n5235)));
	assign x15381x = (((!n_n5325) & (!n_n5329) & (!n_n5236) & (n_n5237)) + ((!n_n5325) & (!n_n5329) & (n_n5236) & (!n_n5237)) + ((!n_n5325) & (!n_n5329) & (n_n5236) & (n_n5237)) + ((!n_n5325) & (n_n5329) & (!n_n5236) & (!n_n5237)) + ((!n_n5325) & (n_n5329) & (!n_n5236) & (n_n5237)) + ((!n_n5325) & (n_n5329) & (n_n5236) & (!n_n5237)) + ((!n_n5325) & (n_n5329) & (n_n5236) & (n_n5237)) + ((n_n5325) & (!n_n5329) & (!n_n5236) & (!n_n5237)) + ((n_n5325) & (!n_n5329) & (!n_n5236) & (n_n5237)) + ((n_n5325) & (!n_n5329) & (n_n5236) & (!n_n5237)) + ((n_n5325) & (!n_n5329) & (n_n5236) & (n_n5237)) + ((n_n5325) & (n_n5329) & (!n_n5236) & (!n_n5237)) + ((n_n5325) & (n_n5329) & (!n_n5236) & (n_n5237)) + ((n_n5325) & (n_n5329) & (n_n5236) & (!n_n5237)) + ((n_n5325) & (n_n5329) & (n_n5236) & (n_n5237)));
	assign x15382x = (((!n_n5302) & (!n_n5273) & (!n_n5327) & (n_n5254)) + ((!n_n5302) & (!n_n5273) & (n_n5327) & (!n_n5254)) + ((!n_n5302) & (!n_n5273) & (n_n5327) & (n_n5254)) + ((!n_n5302) & (n_n5273) & (!n_n5327) & (!n_n5254)) + ((!n_n5302) & (n_n5273) & (!n_n5327) & (n_n5254)) + ((!n_n5302) & (n_n5273) & (n_n5327) & (!n_n5254)) + ((!n_n5302) & (n_n5273) & (n_n5327) & (n_n5254)) + ((n_n5302) & (!n_n5273) & (!n_n5327) & (!n_n5254)) + ((n_n5302) & (!n_n5273) & (!n_n5327) & (n_n5254)) + ((n_n5302) & (!n_n5273) & (n_n5327) & (!n_n5254)) + ((n_n5302) & (!n_n5273) & (n_n5327) & (n_n5254)) + ((n_n5302) & (n_n5273) & (!n_n5327) & (!n_n5254)) + ((n_n5302) & (n_n5273) & (!n_n5327) & (n_n5254)) + ((n_n5302) & (n_n5273) & (n_n5327) & (!n_n5254)) + ((n_n5302) & (n_n5273) & (n_n5327) & (n_n5254)));
	assign x15383x = (((!n_n5296) & (!n_n5319) & (!n_n5278) & (!n_n5298) & (n_n5282)) + ((!n_n5296) & (!n_n5319) & (!n_n5278) & (n_n5298) & (!n_n5282)) + ((!n_n5296) & (!n_n5319) & (!n_n5278) & (n_n5298) & (n_n5282)) + ((!n_n5296) & (!n_n5319) & (n_n5278) & (!n_n5298) & (!n_n5282)) + ((!n_n5296) & (!n_n5319) & (n_n5278) & (!n_n5298) & (n_n5282)) + ((!n_n5296) & (!n_n5319) & (n_n5278) & (n_n5298) & (!n_n5282)) + ((!n_n5296) & (!n_n5319) & (n_n5278) & (n_n5298) & (n_n5282)) + ((!n_n5296) & (n_n5319) & (!n_n5278) & (!n_n5298) & (!n_n5282)) + ((!n_n5296) & (n_n5319) & (!n_n5278) & (!n_n5298) & (n_n5282)) + ((!n_n5296) & (n_n5319) & (!n_n5278) & (n_n5298) & (!n_n5282)) + ((!n_n5296) & (n_n5319) & (!n_n5278) & (n_n5298) & (n_n5282)) + ((!n_n5296) & (n_n5319) & (n_n5278) & (!n_n5298) & (!n_n5282)) + ((!n_n5296) & (n_n5319) & (n_n5278) & (!n_n5298) & (n_n5282)) + ((!n_n5296) & (n_n5319) & (n_n5278) & (n_n5298) & (!n_n5282)) + ((!n_n5296) & (n_n5319) & (n_n5278) & (n_n5298) & (n_n5282)) + ((n_n5296) & (!n_n5319) & (!n_n5278) & (!n_n5298) & (!n_n5282)) + ((n_n5296) & (!n_n5319) & (!n_n5278) & (!n_n5298) & (n_n5282)) + ((n_n5296) & (!n_n5319) & (!n_n5278) & (n_n5298) & (!n_n5282)) + ((n_n5296) & (!n_n5319) & (!n_n5278) & (n_n5298) & (n_n5282)) + ((n_n5296) & (!n_n5319) & (n_n5278) & (!n_n5298) & (!n_n5282)) + ((n_n5296) & (!n_n5319) & (n_n5278) & (!n_n5298) & (n_n5282)) + ((n_n5296) & (!n_n5319) & (n_n5278) & (n_n5298) & (!n_n5282)) + ((n_n5296) & (!n_n5319) & (n_n5278) & (n_n5298) & (n_n5282)) + ((n_n5296) & (n_n5319) & (!n_n5278) & (!n_n5298) & (!n_n5282)) + ((n_n5296) & (n_n5319) & (!n_n5278) & (!n_n5298) & (n_n5282)) + ((n_n5296) & (n_n5319) & (!n_n5278) & (n_n5298) & (!n_n5282)) + ((n_n5296) & (n_n5319) & (!n_n5278) & (n_n5298) & (n_n5282)) + ((n_n5296) & (n_n5319) & (n_n5278) & (!n_n5298) & (!n_n5282)) + ((n_n5296) & (n_n5319) & (n_n5278) & (!n_n5298) & (n_n5282)) + ((n_n5296) & (n_n5319) & (n_n5278) & (n_n5298) & (!n_n5282)) + ((n_n5296) & (n_n5319) & (n_n5278) & (n_n5298) & (n_n5282)));
	assign x22083x = (((!n_n4980) & (!n_n4963) & (!n_n4964) & (!n_n4986)));
	assign n_n2835 = (((!n_n4974) & (!n_n4967) & (!n_n4961) & (!x210x) & (!x22083x)) + ((!n_n4974) & (!n_n4967) & (!n_n4961) & (x210x) & (!x22083x)) + ((!n_n4974) & (!n_n4967) & (!n_n4961) & (x210x) & (x22083x)) + ((!n_n4974) & (!n_n4967) & (n_n4961) & (!x210x) & (!x22083x)) + ((!n_n4974) & (!n_n4967) & (n_n4961) & (!x210x) & (x22083x)) + ((!n_n4974) & (!n_n4967) & (n_n4961) & (x210x) & (!x22083x)) + ((!n_n4974) & (!n_n4967) & (n_n4961) & (x210x) & (x22083x)) + ((!n_n4974) & (n_n4967) & (!n_n4961) & (!x210x) & (!x22083x)) + ((!n_n4974) & (n_n4967) & (!n_n4961) & (!x210x) & (x22083x)) + ((!n_n4974) & (n_n4967) & (!n_n4961) & (x210x) & (!x22083x)) + ((!n_n4974) & (n_n4967) & (!n_n4961) & (x210x) & (x22083x)) + ((!n_n4974) & (n_n4967) & (n_n4961) & (!x210x) & (!x22083x)) + ((!n_n4974) & (n_n4967) & (n_n4961) & (!x210x) & (x22083x)) + ((!n_n4974) & (n_n4967) & (n_n4961) & (x210x) & (!x22083x)) + ((!n_n4974) & (n_n4967) & (n_n4961) & (x210x) & (x22083x)) + ((n_n4974) & (!n_n4967) & (!n_n4961) & (!x210x) & (!x22083x)) + ((n_n4974) & (!n_n4967) & (!n_n4961) & (!x210x) & (x22083x)) + ((n_n4974) & (!n_n4967) & (!n_n4961) & (x210x) & (!x22083x)) + ((n_n4974) & (!n_n4967) & (!n_n4961) & (x210x) & (x22083x)) + ((n_n4974) & (!n_n4967) & (n_n4961) & (!x210x) & (!x22083x)) + ((n_n4974) & (!n_n4967) & (n_n4961) & (!x210x) & (x22083x)) + ((n_n4974) & (!n_n4967) & (n_n4961) & (x210x) & (!x22083x)) + ((n_n4974) & (!n_n4967) & (n_n4961) & (x210x) & (x22083x)) + ((n_n4974) & (n_n4967) & (!n_n4961) & (!x210x) & (!x22083x)) + ((n_n4974) & (n_n4967) & (!n_n4961) & (!x210x) & (x22083x)) + ((n_n4974) & (n_n4967) & (!n_n4961) & (x210x) & (!x22083x)) + ((n_n4974) & (n_n4967) & (!n_n4961) & (x210x) & (x22083x)) + ((n_n4974) & (n_n4967) & (n_n4961) & (!x210x) & (!x22083x)) + ((n_n4974) & (n_n4967) & (n_n4961) & (!x210x) & (x22083x)) + ((n_n4974) & (n_n4967) & (n_n4961) & (x210x) & (!x22083x)) + ((n_n4974) & (n_n4967) & (n_n4961) & (x210x) & (x22083x)));
	assign x15082x = (((!i_9_) & (n_n455) & (!n_n534) & (n_n509) & (n_n530)) + ((!i_9_) & (n_n455) & (n_n534) & (n_n509) & (!n_n530)) + ((!i_9_) & (n_n455) & (n_n534) & (n_n509) & (n_n530)));
	assign x16095x = (((!i_9_) & (!n_n536) & (!x502x) & (!n_n4414) & (n_n2803)) + ((!i_9_) & (!n_n536) & (!x502x) & (n_n4414) & (!n_n2803)) + ((!i_9_) & (!n_n536) & (!x502x) & (n_n4414) & (n_n2803)) + ((!i_9_) & (!n_n536) & (x502x) & (!n_n4414) & (n_n2803)) + ((!i_9_) & (!n_n536) & (x502x) & (n_n4414) & (!n_n2803)) + ((!i_9_) & (!n_n536) & (x502x) & (n_n4414) & (n_n2803)) + ((!i_9_) & (n_n536) & (!x502x) & (!n_n4414) & (n_n2803)) + ((!i_9_) & (n_n536) & (!x502x) & (n_n4414) & (!n_n2803)) + ((!i_9_) & (n_n536) & (!x502x) & (n_n4414) & (n_n2803)) + ((!i_9_) & (n_n536) & (x502x) & (!n_n4414) & (n_n2803)) + ((!i_9_) & (n_n536) & (x502x) & (n_n4414) & (!n_n2803)) + ((!i_9_) & (n_n536) & (x502x) & (n_n4414) & (n_n2803)) + ((i_9_) & (!n_n536) & (!x502x) & (!n_n4414) & (n_n2803)) + ((i_9_) & (!n_n536) & (!x502x) & (n_n4414) & (!n_n2803)) + ((i_9_) & (!n_n536) & (!x502x) & (n_n4414) & (n_n2803)) + ((i_9_) & (!n_n536) & (x502x) & (!n_n4414) & (n_n2803)) + ((i_9_) & (!n_n536) & (x502x) & (n_n4414) & (!n_n2803)) + ((i_9_) & (!n_n536) & (x502x) & (n_n4414) & (n_n2803)) + ((i_9_) & (n_n536) & (!x502x) & (!n_n4414) & (n_n2803)) + ((i_9_) & (n_n536) & (!x502x) & (n_n4414) & (!n_n2803)) + ((i_9_) & (n_n536) & (!x502x) & (n_n4414) & (n_n2803)) + ((i_9_) & (n_n536) & (x502x) & (!n_n4414) & (!n_n2803)) + ((i_9_) & (n_n536) & (x502x) & (!n_n4414) & (n_n2803)) + ((i_9_) & (n_n536) & (x502x) & (n_n4414) & (!n_n2803)) + ((i_9_) & (n_n536) & (x502x) & (n_n4414) & (n_n2803)));
	assign n_n1890 = (((!n_n4416) & (!n_n4430) & (!x37x) & (x16095x)) + ((!n_n4416) & (!n_n4430) & (x37x) & (!x16095x)) + ((!n_n4416) & (!n_n4430) & (x37x) & (x16095x)) + ((!n_n4416) & (n_n4430) & (!x37x) & (!x16095x)) + ((!n_n4416) & (n_n4430) & (!x37x) & (x16095x)) + ((!n_n4416) & (n_n4430) & (x37x) & (!x16095x)) + ((!n_n4416) & (n_n4430) & (x37x) & (x16095x)) + ((n_n4416) & (!n_n4430) & (!x37x) & (!x16095x)) + ((n_n4416) & (!n_n4430) & (!x37x) & (x16095x)) + ((n_n4416) & (!n_n4430) & (x37x) & (!x16095x)) + ((n_n4416) & (!n_n4430) & (x37x) & (x16095x)) + ((n_n4416) & (n_n4430) & (!x37x) & (!x16095x)) + ((n_n4416) & (n_n4430) & (!x37x) & (x16095x)) + ((n_n4416) & (n_n4430) & (x37x) & (!x16095x)) + ((n_n4416) & (n_n4430) & (x37x) & (x16095x)));
	assign x16099x = (((!n_n4389) & (!n_n4388) & (!n_n4393) & (n_n4390)) + ((!n_n4389) & (!n_n4388) & (n_n4393) & (!n_n4390)) + ((!n_n4389) & (!n_n4388) & (n_n4393) & (n_n4390)) + ((!n_n4389) & (n_n4388) & (!n_n4393) & (!n_n4390)) + ((!n_n4389) & (n_n4388) & (!n_n4393) & (n_n4390)) + ((!n_n4389) & (n_n4388) & (n_n4393) & (!n_n4390)) + ((!n_n4389) & (n_n4388) & (n_n4393) & (n_n4390)) + ((n_n4389) & (!n_n4388) & (!n_n4393) & (!n_n4390)) + ((n_n4389) & (!n_n4388) & (!n_n4393) & (n_n4390)) + ((n_n4389) & (!n_n4388) & (n_n4393) & (!n_n4390)) + ((n_n4389) & (!n_n4388) & (n_n4393) & (n_n4390)) + ((n_n4389) & (n_n4388) & (!n_n4393) & (!n_n4390)) + ((n_n4389) & (n_n4388) & (!n_n4393) & (n_n4390)) + ((n_n4389) & (n_n4388) & (n_n4393) & (!n_n4390)) + ((n_n4389) & (n_n4388) & (n_n4393) & (n_n4390)));
	assign x16100x = (((!n_n4391) & (!n_n4397) & (!n_n4398) & (!n_n4396) & (n_n4399)) + ((!n_n4391) & (!n_n4397) & (!n_n4398) & (n_n4396) & (!n_n4399)) + ((!n_n4391) & (!n_n4397) & (!n_n4398) & (n_n4396) & (n_n4399)) + ((!n_n4391) & (!n_n4397) & (n_n4398) & (!n_n4396) & (!n_n4399)) + ((!n_n4391) & (!n_n4397) & (n_n4398) & (!n_n4396) & (n_n4399)) + ((!n_n4391) & (!n_n4397) & (n_n4398) & (n_n4396) & (!n_n4399)) + ((!n_n4391) & (!n_n4397) & (n_n4398) & (n_n4396) & (n_n4399)) + ((!n_n4391) & (n_n4397) & (!n_n4398) & (!n_n4396) & (!n_n4399)) + ((!n_n4391) & (n_n4397) & (!n_n4398) & (!n_n4396) & (n_n4399)) + ((!n_n4391) & (n_n4397) & (!n_n4398) & (n_n4396) & (!n_n4399)) + ((!n_n4391) & (n_n4397) & (!n_n4398) & (n_n4396) & (n_n4399)) + ((!n_n4391) & (n_n4397) & (n_n4398) & (!n_n4396) & (!n_n4399)) + ((!n_n4391) & (n_n4397) & (n_n4398) & (!n_n4396) & (n_n4399)) + ((!n_n4391) & (n_n4397) & (n_n4398) & (n_n4396) & (!n_n4399)) + ((!n_n4391) & (n_n4397) & (n_n4398) & (n_n4396) & (n_n4399)) + ((n_n4391) & (!n_n4397) & (!n_n4398) & (!n_n4396) & (!n_n4399)) + ((n_n4391) & (!n_n4397) & (!n_n4398) & (!n_n4396) & (n_n4399)) + ((n_n4391) & (!n_n4397) & (!n_n4398) & (n_n4396) & (!n_n4399)) + ((n_n4391) & (!n_n4397) & (!n_n4398) & (n_n4396) & (n_n4399)) + ((n_n4391) & (!n_n4397) & (n_n4398) & (!n_n4396) & (!n_n4399)) + ((n_n4391) & (!n_n4397) & (n_n4398) & (!n_n4396) & (n_n4399)) + ((n_n4391) & (!n_n4397) & (n_n4398) & (n_n4396) & (!n_n4399)) + ((n_n4391) & (!n_n4397) & (n_n4398) & (n_n4396) & (n_n4399)) + ((n_n4391) & (n_n4397) & (!n_n4398) & (!n_n4396) & (!n_n4399)) + ((n_n4391) & (n_n4397) & (!n_n4398) & (!n_n4396) & (n_n4399)) + ((n_n4391) & (n_n4397) & (!n_n4398) & (n_n4396) & (!n_n4399)) + ((n_n4391) & (n_n4397) & (!n_n4398) & (n_n4396) & (n_n4399)) + ((n_n4391) & (n_n4397) & (n_n4398) & (!n_n4396) & (!n_n4399)) + ((n_n4391) & (n_n4397) & (n_n4398) & (!n_n4396) & (n_n4399)) + ((n_n4391) & (n_n4397) & (n_n4398) & (n_n4396) & (!n_n4399)) + ((n_n4391) & (n_n4397) & (n_n4398) & (n_n4396) & (n_n4399)));
	assign x16104x = (((!n_n4403) & (!n_n4400) & (!n_n4405) & (!n_n4406) & (n_n4411)) + ((!n_n4403) & (!n_n4400) & (!n_n4405) & (n_n4406) & (!n_n4411)) + ((!n_n4403) & (!n_n4400) & (!n_n4405) & (n_n4406) & (n_n4411)) + ((!n_n4403) & (!n_n4400) & (n_n4405) & (!n_n4406) & (!n_n4411)) + ((!n_n4403) & (!n_n4400) & (n_n4405) & (!n_n4406) & (n_n4411)) + ((!n_n4403) & (!n_n4400) & (n_n4405) & (n_n4406) & (!n_n4411)) + ((!n_n4403) & (!n_n4400) & (n_n4405) & (n_n4406) & (n_n4411)) + ((!n_n4403) & (n_n4400) & (!n_n4405) & (!n_n4406) & (!n_n4411)) + ((!n_n4403) & (n_n4400) & (!n_n4405) & (!n_n4406) & (n_n4411)) + ((!n_n4403) & (n_n4400) & (!n_n4405) & (n_n4406) & (!n_n4411)) + ((!n_n4403) & (n_n4400) & (!n_n4405) & (n_n4406) & (n_n4411)) + ((!n_n4403) & (n_n4400) & (n_n4405) & (!n_n4406) & (!n_n4411)) + ((!n_n4403) & (n_n4400) & (n_n4405) & (!n_n4406) & (n_n4411)) + ((!n_n4403) & (n_n4400) & (n_n4405) & (n_n4406) & (!n_n4411)) + ((!n_n4403) & (n_n4400) & (n_n4405) & (n_n4406) & (n_n4411)) + ((n_n4403) & (!n_n4400) & (!n_n4405) & (!n_n4406) & (!n_n4411)) + ((n_n4403) & (!n_n4400) & (!n_n4405) & (!n_n4406) & (n_n4411)) + ((n_n4403) & (!n_n4400) & (!n_n4405) & (n_n4406) & (!n_n4411)) + ((n_n4403) & (!n_n4400) & (!n_n4405) & (n_n4406) & (n_n4411)) + ((n_n4403) & (!n_n4400) & (n_n4405) & (!n_n4406) & (!n_n4411)) + ((n_n4403) & (!n_n4400) & (n_n4405) & (!n_n4406) & (n_n4411)) + ((n_n4403) & (!n_n4400) & (n_n4405) & (n_n4406) & (!n_n4411)) + ((n_n4403) & (!n_n4400) & (n_n4405) & (n_n4406) & (n_n4411)) + ((n_n4403) & (n_n4400) & (!n_n4405) & (!n_n4406) & (!n_n4411)) + ((n_n4403) & (n_n4400) & (!n_n4405) & (!n_n4406) & (n_n4411)) + ((n_n4403) & (n_n4400) & (!n_n4405) & (n_n4406) & (!n_n4411)) + ((n_n4403) & (n_n4400) & (!n_n4405) & (n_n4406) & (n_n4411)) + ((n_n4403) & (n_n4400) & (n_n4405) & (!n_n4406) & (!n_n4411)) + ((n_n4403) & (n_n4400) & (n_n4405) & (!n_n4406) & (n_n4411)) + ((n_n4403) & (n_n4400) & (n_n4405) & (n_n4406) & (!n_n4411)) + ((n_n4403) & (n_n4400) & (n_n4405) & (n_n4406) & (n_n4411)));
	assign x16105x = (((!n_n4401) & (!n_n4402) & (!n_n4409) & (!n_n4410) & (x16104x)) + ((!n_n4401) & (!n_n4402) & (!n_n4409) & (n_n4410) & (!x16104x)) + ((!n_n4401) & (!n_n4402) & (!n_n4409) & (n_n4410) & (x16104x)) + ((!n_n4401) & (!n_n4402) & (n_n4409) & (!n_n4410) & (!x16104x)) + ((!n_n4401) & (!n_n4402) & (n_n4409) & (!n_n4410) & (x16104x)) + ((!n_n4401) & (!n_n4402) & (n_n4409) & (n_n4410) & (!x16104x)) + ((!n_n4401) & (!n_n4402) & (n_n4409) & (n_n4410) & (x16104x)) + ((!n_n4401) & (n_n4402) & (!n_n4409) & (!n_n4410) & (!x16104x)) + ((!n_n4401) & (n_n4402) & (!n_n4409) & (!n_n4410) & (x16104x)) + ((!n_n4401) & (n_n4402) & (!n_n4409) & (n_n4410) & (!x16104x)) + ((!n_n4401) & (n_n4402) & (!n_n4409) & (n_n4410) & (x16104x)) + ((!n_n4401) & (n_n4402) & (n_n4409) & (!n_n4410) & (!x16104x)) + ((!n_n4401) & (n_n4402) & (n_n4409) & (!n_n4410) & (x16104x)) + ((!n_n4401) & (n_n4402) & (n_n4409) & (n_n4410) & (!x16104x)) + ((!n_n4401) & (n_n4402) & (n_n4409) & (n_n4410) & (x16104x)) + ((n_n4401) & (!n_n4402) & (!n_n4409) & (!n_n4410) & (!x16104x)) + ((n_n4401) & (!n_n4402) & (!n_n4409) & (!n_n4410) & (x16104x)) + ((n_n4401) & (!n_n4402) & (!n_n4409) & (n_n4410) & (!x16104x)) + ((n_n4401) & (!n_n4402) & (!n_n4409) & (n_n4410) & (x16104x)) + ((n_n4401) & (!n_n4402) & (n_n4409) & (!n_n4410) & (!x16104x)) + ((n_n4401) & (!n_n4402) & (n_n4409) & (!n_n4410) & (x16104x)) + ((n_n4401) & (!n_n4402) & (n_n4409) & (n_n4410) & (!x16104x)) + ((n_n4401) & (!n_n4402) & (n_n4409) & (n_n4410) & (x16104x)) + ((n_n4401) & (n_n4402) & (!n_n4409) & (!n_n4410) & (!x16104x)) + ((n_n4401) & (n_n4402) & (!n_n4409) & (!n_n4410) & (x16104x)) + ((n_n4401) & (n_n4402) & (!n_n4409) & (n_n4410) & (!x16104x)) + ((n_n4401) & (n_n4402) & (!n_n4409) & (n_n4410) & (x16104x)) + ((n_n4401) & (n_n4402) & (n_n4409) & (!n_n4410) & (!x16104x)) + ((n_n4401) & (n_n4402) & (n_n4409) & (!n_n4410) & (x16104x)) + ((n_n4401) & (n_n4402) & (n_n4409) & (n_n4410) & (!x16104x)) + ((n_n4401) & (n_n4402) & (n_n4409) & (n_n4410) & (x16104x)));
	assign x16227x = (((!x15x) & (n_n482) & (!n_n473) & (n_n325) & (x20x)) + ((!x15x) & (n_n482) & (n_n473) & (n_n325) & (x20x)) + ((x15x) & (!n_n482) & (n_n473) & (n_n325) & (!x20x)) + ((x15x) & (!n_n482) & (n_n473) & (n_n325) & (x20x)) + ((x15x) & (n_n482) & (!n_n473) & (n_n325) & (x20x)) + ((x15x) & (n_n482) & (n_n473) & (n_n325) & (!x20x)) + ((x15x) & (n_n482) & (n_n473) & (n_n325) & (x20x)));
	assign n_n1863 = (((!n_n4791) & (!n_n4792) & (!n_n2003) & (!x380x) & (x16227x)) + ((!n_n4791) & (!n_n4792) & (!n_n2003) & (x380x) & (!x16227x)) + ((!n_n4791) & (!n_n4792) & (!n_n2003) & (x380x) & (x16227x)) + ((!n_n4791) & (!n_n4792) & (n_n2003) & (!x380x) & (!x16227x)) + ((!n_n4791) & (!n_n4792) & (n_n2003) & (!x380x) & (x16227x)) + ((!n_n4791) & (!n_n4792) & (n_n2003) & (x380x) & (!x16227x)) + ((!n_n4791) & (!n_n4792) & (n_n2003) & (x380x) & (x16227x)) + ((!n_n4791) & (n_n4792) & (!n_n2003) & (!x380x) & (!x16227x)) + ((!n_n4791) & (n_n4792) & (!n_n2003) & (!x380x) & (x16227x)) + ((!n_n4791) & (n_n4792) & (!n_n2003) & (x380x) & (!x16227x)) + ((!n_n4791) & (n_n4792) & (!n_n2003) & (x380x) & (x16227x)) + ((!n_n4791) & (n_n4792) & (n_n2003) & (!x380x) & (!x16227x)) + ((!n_n4791) & (n_n4792) & (n_n2003) & (!x380x) & (x16227x)) + ((!n_n4791) & (n_n4792) & (n_n2003) & (x380x) & (!x16227x)) + ((!n_n4791) & (n_n4792) & (n_n2003) & (x380x) & (x16227x)) + ((n_n4791) & (!n_n4792) & (!n_n2003) & (!x380x) & (!x16227x)) + ((n_n4791) & (!n_n4792) & (!n_n2003) & (!x380x) & (x16227x)) + ((n_n4791) & (!n_n4792) & (!n_n2003) & (x380x) & (!x16227x)) + ((n_n4791) & (!n_n4792) & (!n_n2003) & (x380x) & (x16227x)) + ((n_n4791) & (!n_n4792) & (n_n2003) & (!x380x) & (!x16227x)) + ((n_n4791) & (!n_n4792) & (n_n2003) & (!x380x) & (x16227x)) + ((n_n4791) & (!n_n4792) & (n_n2003) & (x380x) & (!x16227x)) + ((n_n4791) & (!n_n4792) & (n_n2003) & (x380x) & (x16227x)) + ((n_n4791) & (n_n4792) & (!n_n2003) & (!x380x) & (!x16227x)) + ((n_n4791) & (n_n4792) & (!n_n2003) & (!x380x) & (x16227x)) + ((n_n4791) & (n_n4792) & (!n_n2003) & (x380x) & (!x16227x)) + ((n_n4791) & (n_n4792) & (!n_n2003) & (x380x) & (x16227x)) + ((n_n4791) & (n_n4792) & (n_n2003) & (!x380x) & (!x16227x)) + ((n_n4791) & (n_n4792) & (n_n2003) & (!x380x) & (x16227x)) + ((n_n4791) & (n_n4792) & (n_n2003) & (x380x) & (!x16227x)) + ((n_n4791) & (n_n4792) & (n_n2003) & (x380x) & (x16227x)));
	assign x16233x = (((!n_n4757) & (!n_n4759) & (!n_n4760) & (n_n4767)) + ((!n_n4757) & (!n_n4759) & (n_n4760) & (!n_n4767)) + ((!n_n4757) & (!n_n4759) & (n_n4760) & (n_n4767)) + ((!n_n4757) & (n_n4759) & (!n_n4760) & (!n_n4767)) + ((!n_n4757) & (n_n4759) & (!n_n4760) & (n_n4767)) + ((!n_n4757) & (n_n4759) & (n_n4760) & (!n_n4767)) + ((!n_n4757) & (n_n4759) & (n_n4760) & (n_n4767)) + ((n_n4757) & (!n_n4759) & (!n_n4760) & (!n_n4767)) + ((n_n4757) & (!n_n4759) & (!n_n4760) & (n_n4767)) + ((n_n4757) & (!n_n4759) & (n_n4760) & (!n_n4767)) + ((n_n4757) & (!n_n4759) & (n_n4760) & (n_n4767)) + ((n_n4757) & (n_n4759) & (!n_n4760) & (!n_n4767)) + ((n_n4757) & (n_n4759) & (!n_n4760) & (n_n4767)) + ((n_n4757) & (n_n4759) & (n_n4760) & (!n_n4767)) + ((n_n4757) & (n_n4759) & (n_n4760) & (n_n4767)));
	assign x16234x = (((!n_n4761) & (!n_n4762) & (!n_n4764) & (!n_n4765) & (n_n4763)) + ((!n_n4761) & (!n_n4762) & (!n_n4764) & (n_n4765) & (!n_n4763)) + ((!n_n4761) & (!n_n4762) & (!n_n4764) & (n_n4765) & (n_n4763)) + ((!n_n4761) & (!n_n4762) & (n_n4764) & (!n_n4765) & (!n_n4763)) + ((!n_n4761) & (!n_n4762) & (n_n4764) & (!n_n4765) & (n_n4763)) + ((!n_n4761) & (!n_n4762) & (n_n4764) & (n_n4765) & (!n_n4763)) + ((!n_n4761) & (!n_n4762) & (n_n4764) & (n_n4765) & (n_n4763)) + ((!n_n4761) & (n_n4762) & (!n_n4764) & (!n_n4765) & (!n_n4763)) + ((!n_n4761) & (n_n4762) & (!n_n4764) & (!n_n4765) & (n_n4763)) + ((!n_n4761) & (n_n4762) & (!n_n4764) & (n_n4765) & (!n_n4763)) + ((!n_n4761) & (n_n4762) & (!n_n4764) & (n_n4765) & (n_n4763)) + ((!n_n4761) & (n_n4762) & (n_n4764) & (!n_n4765) & (!n_n4763)) + ((!n_n4761) & (n_n4762) & (n_n4764) & (!n_n4765) & (n_n4763)) + ((!n_n4761) & (n_n4762) & (n_n4764) & (n_n4765) & (!n_n4763)) + ((!n_n4761) & (n_n4762) & (n_n4764) & (n_n4765) & (n_n4763)) + ((n_n4761) & (!n_n4762) & (!n_n4764) & (!n_n4765) & (!n_n4763)) + ((n_n4761) & (!n_n4762) & (!n_n4764) & (!n_n4765) & (n_n4763)) + ((n_n4761) & (!n_n4762) & (!n_n4764) & (n_n4765) & (!n_n4763)) + ((n_n4761) & (!n_n4762) & (!n_n4764) & (n_n4765) & (n_n4763)) + ((n_n4761) & (!n_n4762) & (n_n4764) & (!n_n4765) & (!n_n4763)) + ((n_n4761) & (!n_n4762) & (n_n4764) & (!n_n4765) & (n_n4763)) + ((n_n4761) & (!n_n4762) & (n_n4764) & (n_n4765) & (!n_n4763)) + ((n_n4761) & (!n_n4762) & (n_n4764) & (n_n4765) & (n_n4763)) + ((n_n4761) & (n_n4762) & (!n_n4764) & (!n_n4765) & (!n_n4763)) + ((n_n4761) & (n_n4762) & (!n_n4764) & (!n_n4765) & (n_n4763)) + ((n_n4761) & (n_n4762) & (!n_n4764) & (n_n4765) & (!n_n4763)) + ((n_n4761) & (n_n4762) & (!n_n4764) & (n_n4765) & (n_n4763)) + ((n_n4761) & (n_n4762) & (n_n4764) & (!n_n4765) & (!n_n4763)) + ((n_n4761) & (n_n4762) & (n_n4764) & (!n_n4765) & (n_n4763)) + ((n_n4761) & (n_n4762) & (n_n4764) & (n_n4765) & (!n_n4763)) + ((n_n4761) & (n_n4762) & (n_n4764) & (n_n4765) & (n_n4763)));
	assign x12410x = (((!n_n4725) & (!n_n4726) & (!n_n4730) & (!n_n4722) & (n_n4721)) + ((!n_n4725) & (!n_n4726) & (!n_n4730) & (n_n4722) & (!n_n4721)) + ((!n_n4725) & (!n_n4726) & (!n_n4730) & (n_n4722) & (n_n4721)) + ((!n_n4725) & (!n_n4726) & (n_n4730) & (!n_n4722) & (!n_n4721)) + ((!n_n4725) & (!n_n4726) & (n_n4730) & (!n_n4722) & (n_n4721)) + ((!n_n4725) & (!n_n4726) & (n_n4730) & (n_n4722) & (!n_n4721)) + ((!n_n4725) & (!n_n4726) & (n_n4730) & (n_n4722) & (n_n4721)) + ((!n_n4725) & (n_n4726) & (!n_n4730) & (!n_n4722) & (!n_n4721)) + ((!n_n4725) & (n_n4726) & (!n_n4730) & (!n_n4722) & (n_n4721)) + ((!n_n4725) & (n_n4726) & (!n_n4730) & (n_n4722) & (!n_n4721)) + ((!n_n4725) & (n_n4726) & (!n_n4730) & (n_n4722) & (n_n4721)) + ((!n_n4725) & (n_n4726) & (n_n4730) & (!n_n4722) & (!n_n4721)) + ((!n_n4725) & (n_n4726) & (n_n4730) & (!n_n4722) & (n_n4721)) + ((!n_n4725) & (n_n4726) & (n_n4730) & (n_n4722) & (!n_n4721)) + ((!n_n4725) & (n_n4726) & (n_n4730) & (n_n4722) & (n_n4721)) + ((n_n4725) & (!n_n4726) & (!n_n4730) & (!n_n4722) & (!n_n4721)) + ((n_n4725) & (!n_n4726) & (!n_n4730) & (!n_n4722) & (n_n4721)) + ((n_n4725) & (!n_n4726) & (!n_n4730) & (n_n4722) & (!n_n4721)) + ((n_n4725) & (!n_n4726) & (!n_n4730) & (n_n4722) & (n_n4721)) + ((n_n4725) & (!n_n4726) & (n_n4730) & (!n_n4722) & (!n_n4721)) + ((n_n4725) & (!n_n4726) & (n_n4730) & (!n_n4722) & (n_n4721)) + ((n_n4725) & (!n_n4726) & (n_n4730) & (n_n4722) & (!n_n4721)) + ((n_n4725) & (!n_n4726) & (n_n4730) & (n_n4722) & (n_n4721)) + ((n_n4725) & (n_n4726) & (!n_n4730) & (!n_n4722) & (!n_n4721)) + ((n_n4725) & (n_n4726) & (!n_n4730) & (!n_n4722) & (n_n4721)) + ((n_n4725) & (n_n4726) & (!n_n4730) & (n_n4722) & (!n_n4721)) + ((n_n4725) & (n_n4726) & (!n_n4730) & (n_n4722) & (n_n4721)) + ((n_n4725) & (n_n4726) & (n_n4730) & (!n_n4722) & (!n_n4721)) + ((n_n4725) & (n_n4726) & (n_n4730) & (!n_n4722) & (n_n4721)) + ((n_n4725) & (n_n4726) & (n_n4730) & (n_n4722) & (!n_n4721)) + ((n_n4725) & (n_n4726) & (n_n4730) & (n_n4722) & (n_n4721)));
	assign x11713x = (((!n_n5142) & (!n_n5130) & (!n_n5108) & (!n_n5118) & (n_n5119)) + ((!n_n5142) & (!n_n5130) & (!n_n5108) & (n_n5118) & (!n_n5119)) + ((!n_n5142) & (!n_n5130) & (!n_n5108) & (n_n5118) & (n_n5119)) + ((!n_n5142) & (!n_n5130) & (n_n5108) & (!n_n5118) & (!n_n5119)) + ((!n_n5142) & (!n_n5130) & (n_n5108) & (!n_n5118) & (n_n5119)) + ((!n_n5142) & (!n_n5130) & (n_n5108) & (n_n5118) & (!n_n5119)) + ((!n_n5142) & (!n_n5130) & (n_n5108) & (n_n5118) & (n_n5119)) + ((!n_n5142) & (n_n5130) & (!n_n5108) & (!n_n5118) & (!n_n5119)) + ((!n_n5142) & (n_n5130) & (!n_n5108) & (!n_n5118) & (n_n5119)) + ((!n_n5142) & (n_n5130) & (!n_n5108) & (n_n5118) & (!n_n5119)) + ((!n_n5142) & (n_n5130) & (!n_n5108) & (n_n5118) & (n_n5119)) + ((!n_n5142) & (n_n5130) & (n_n5108) & (!n_n5118) & (!n_n5119)) + ((!n_n5142) & (n_n5130) & (n_n5108) & (!n_n5118) & (n_n5119)) + ((!n_n5142) & (n_n5130) & (n_n5108) & (n_n5118) & (!n_n5119)) + ((!n_n5142) & (n_n5130) & (n_n5108) & (n_n5118) & (n_n5119)) + ((n_n5142) & (!n_n5130) & (!n_n5108) & (!n_n5118) & (!n_n5119)) + ((n_n5142) & (!n_n5130) & (!n_n5108) & (!n_n5118) & (n_n5119)) + ((n_n5142) & (!n_n5130) & (!n_n5108) & (n_n5118) & (!n_n5119)) + ((n_n5142) & (!n_n5130) & (!n_n5108) & (n_n5118) & (n_n5119)) + ((n_n5142) & (!n_n5130) & (n_n5108) & (!n_n5118) & (!n_n5119)) + ((n_n5142) & (!n_n5130) & (n_n5108) & (!n_n5118) & (n_n5119)) + ((n_n5142) & (!n_n5130) & (n_n5108) & (n_n5118) & (!n_n5119)) + ((n_n5142) & (!n_n5130) & (n_n5108) & (n_n5118) & (n_n5119)) + ((n_n5142) & (n_n5130) & (!n_n5108) & (!n_n5118) & (!n_n5119)) + ((n_n5142) & (n_n5130) & (!n_n5108) & (!n_n5118) & (n_n5119)) + ((n_n5142) & (n_n5130) & (!n_n5108) & (n_n5118) & (!n_n5119)) + ((n_n5142) & (n_n5130) & (!n_n5108) & (n_n5118) & (n_n5119)) + ((n_n5142) & (n_n5130) & (n_n5108) & (!n_n5118) & (!n_n5119)) + ((n_n5142) & (n_n5130) & (n_n5108) & (!n_n5118) & (n_n5119)) + ((n_n5142) & (n_n5130) & (n_n5108) & (n_n5118) & (!n_n5119)) + ((n_n5142) & (n_n5130) & (n_n5108) & (n_n5118) & (n_n5119)));
	assign n_n947 = (((!n_n5113) & (!n_n5155) & (!n_n5161) & (!n_n5127) & (x11713x)) + ((!n_n5113) & (!n_n5155) & (!n_n5161) & (n_n5127) & (!x11713x)) + ((!n_n5113) & (!n_n5155) & (!n_n5161) & (n_n5127) & (x11713x)) + ((!n_n5113) & (!n_n5155) & (n_n5161) & (!n_n5127) & (!x11713x)) + ((!n_n5113) & (!n_n5155) & (n_n5161) & (!n_n5127) & (x11713x)) + ((!n_n5113) & (!n_n5155) & (n_n5161) & (n_n5127) & (!x11713x)) + ((!n_n5113) & (!n_n5155) & (n_n5161) & (n_n5127) & (x11713x)) + ((!n_n5113) & (n_n5155) & (!n_n5161) & (!n_n5127) & (!x11713x)) + ((!n_n5113) & (n_n5155) & (!n_n5161) & (!n_n5127) & (x11713x)) + ((!n_n5113) & (n_n5155) & (!n_n5161) & (n_n5127) & (!x11713x)) + ((!n_n5113) & (n_n5155) & (!n_n5161) & (n_n5127) & (x11713x)) + ((!n_n5113) & (n_n5155) & (n_n5161) & (!n_n5127) & (!x11713x)) + ((!n_n5113) & (n_n5155) & (n_n5161) & (!n_n5127) & (x11713x)) + ((!n_n5113) & (n_n5155) & (n_n5161) & (n_n5127) & (!x11713x)) + ((!n_n5113) & (n_n5155) & (n_n5161) & (n_n5127) & (x11713x)) + ((n_n5113) & (!n_n5155) & (!n_n5161) & (!n_n5127) & (!x11713x)) + ((n_n5113) & (!n_n5155) & (!n_n5161) & (!n_n5127) & (x11713x)) + ((n_n5113) & (!n_n5155) & (!n_n5161) & (n_n5127) & (!x11713x)) + ((n_n5113) & (!n_n5155) & (!n_n5161) & (n_n5127) & (x11713x)) + ((n_n5113) & (!n_n5155) & (n_n5161) & (!n_n5127) & (!x11713x)) + ((n_n5113) & (!n_n5155) & (n_n5161) & (!n_n5127) & (x11713x)) + ((n_n5113) & (!n_n5155) & (n_n5161) & (n_n5127) & (!x11713x)) + ((n_n5113) & (!n_n5155) & (n_n5161) & (n_n5127) & (x11713x)) + ((n_n5113) & (n_n5155) & (!n_n5161) & (!n_n5127) & (!x11713x)) + ((n_n5113) & (n_n5155) & (!n_n5161) & (!n_n5127) & (x11713x)) + ((n_n5113) & (n_n5155) & (!n_n5161) & (n_n5127) & (!x11713x)) + ((n_n5113) & (n_n5155) & (!n_n5161) & (n_n5127) & (x11713x)) + ((n_n5113) & (n_n5155) & (n_n5161) & (!n_n5127) & (!x11713x)) + ((n_n5113) & (n_n5155) & (n_n5161) & (!n_n5127) & (x11713x)) + ((n_n5113) & (n_n5155) & (n_n5161) & (n_n5127) & (!x11713x)) + ((n_n5113) & (n_n5155) & (n_n5161) & (n_n5127) & (x11713x)));
	assign x13051x = (((!i_9_) & (!n_n536) & (!n_n518) & (!n_n534) & (n_n4325)) + ((!i_9_) & (!n_n536) & (!n_n518) & (n_n534) & (n_n4325)) + ((!i_9_) & (!n_n536) & (n_n518) & (!n_n534) & (n_n4325)) + ((!i_9_) & (!n_n536) & (n_n518) & (n_n534) & (n_n4325)) + ((!i_9_) & (n_n536) & (!n_n518) & (!n_n534) & (n_n4325)) + ((!i_9_) & (n_n536) & (!n_n518) & (n_n534) & (n_n4325)) + ((!i_9_) & (n_n536) & (n_n518) & (!n_n534) & (n_n4325)) + ((!i_9_) & (n_n536) & (n_n518) & (n_n534) & (!n_n4325)) + ((!i_9_) & (n_n536) & (n_n518) & (n_n534) & (n_n4325)) + ((i_9_) & (!n_n536) & (!n_n518) & (!n_n534) & (n_n4325)) + ((i_9_) & (!n_n536) & (!n_n518) & (n_n534) & (n_n4325)) + ((i_9_) & (!n_n536) & (n_n518) & (!n_n534) & (n_n4325)) + ((i_9_) & (!n_n536) & (n_n518) & (n_n534) & (n_n4325)) + ((i_9_) & (n_n536) & (!n_n518) & (!n_n534) & (n_n4325)) + ((i_9_) & (n_n536) & (!n_n518) & (n_n534) & (n_n4325)) + ((i_9_) & (n_n536) & (n_n518) & (!n_n534) & (n_n4325)) + ((i_9_) & (n_n536) & (n_n518) & (n_n534) & (n_n4325)));
	assign n_n737 = (((!n_n4330) & (!n_n4323) & (!x443x) & (!x448x) & (x13051x)) + ((!n_n4330) & (!n_n4323) & (!x443x) & (x448x) & (!x13051x)) + ((!n_n4330) & (!n_n4323) & (!x443x) & (x448x) & (x13051x)) + ((!n_n4330) & (!n_n4323) & (x443x) & (!x448x) & (!x13051x)) + ((!n_n4330) & (!n_n4323) & (x443x) & (!x448x) & (x13051x)) + ((!n_n4330) & (!n_n4323) & (x443x) & (x448x) & (!x13051x)) + ((!n_n4330) & (!n_n4323) & (x443x) & (x448x) & (x13051x)) + ((!n_n4330) & (n_n4323) & (!x443x) & (!x448x) & (!x13051x)) + ((!n_n4330) & (n_n4323) & (!x443x) & (!x448x) & (x13051x)) + ((!n_n4330) & (n_n4323) & (!x443x) & (x448x) & (!x13051x)) + ((!n_n4330) & (n_n4323) & (!x443x) & (x448x) & (x13051x)) + ((!n_n4330) & (n_n4323) & (x443x) & (!x448x) & (!x13051x)) + ((!n_n4330) & (n_n4323) & (x443x) & (!x448x) & (x13051x)) + ((!n_n4330) & (n_n4323) & (x443x) & (x448x) & (!x13051x)) + ((!n_n4330) & (n_n4323) & (x443x) & (x448x) & (x13051x)) + ((n_n4330) & (!n_n4323) & (!x443x) & (!x448x) & (!x13051x)) + ((n_n4330) & (!n_n4323) & (!x443x) & (!x448x) & (x13051x)) + ((n_n4330) & (!n_n4323) & (!x443x) & (x448x) & (!x13051x)) + ((n_n4330) & (!n_n4323) & (!x443x) & (x448x) & (x13051x)) + ((n_n4330) & (!n_n4323) & (x443x) & (!x448x) & (!x13051x)) + ((n_n4330) & (!n_n4323) & (x443x) & (!x448x) & (x13051x)) + ((n_n4330) & (!n_n4323) & (x443x) & (x448x) & (!x13051x)) + ((n_n4330) & (!n_n4323) & (x443x) & (x448x) & (x13051x)) + ((n_n4330) & (n_n4323) & (!x443x) & (!x448x) & (!x13051x)) + ((n_n4330) & (n_n4323) & (!x443x) & (!x448x) & (x13051x)) + ((n_n4330) & (n_n4323) & (!x443x) & (x448x) & (!x13051x)) + ((n_n4330) & (n_n4323) & (!x443x) & (x448x) & (x13051x)) + ((n_n4330) & (n_n4323) & (x443x) & (!x448x) & (!x13051x)) + ((n_n4330) & (n_n4323) & (x443x) & (!x448x) & (x13051x)) + ((n_n4330) & (n_n4323) & (x443x) & (x448x) & (!x13051x)) + ((n_n4330) & (n_n4323) & (x443x) & (x448x) & (x13051x)));
	assign x22134x = (((!x13x) & (!x506x) & (!n_n4544) & (!n_n4542) & (!n_n4541)) + ((!x13x) & (x506x) & (!n_n4544) & (!n_n4542) & (!n_n4541)) + ((x13x) & (!x506x) & (!n_n4544) & (!n_n4542) & (!n_n4541)));
	assign n_n719 = (((!n_n4548) & (!n_n4551) & (!n_n4545) & (!x13091x) & (!x22134x)) + ((!n_n4548) & (!n_n4551) & (!n_n4545) & (x13091x) & (!x22134x)) + ((!n_n4548) & (!n_n4551) & (!n_n4545) & (x13091x) & (x22134x)) + ((!n_n4548) & (!n_n4551) & (n_n4545) & (!x13091x) & (!x22134x)) + ((!n_n4548) & (!n_n4551) & (n_n4545) & (!x13091x) & (x22134x)) + ((!n_n4548) & (!n_n4551) & (n_n4545) & (x13091x) & (!x22134x)) + ((!n_n4548) & (!n_n4551) & (n_n4545) & (x13091x) & (x22134x)) + ((!n_n4548) & (n_n4551) & (!n_n4545) & (!x13091x) & (!x22134x)) + ((!n_n4548) & (n_n4551) & (!n_n4545) & (!x13091x) & (x22134x)) + ((!n_n4548) & (n_n4551) & (!n_n4545) & (x13091x) & (!x22134x)) + ((!n_n4548) & (n_n4551) & (!n_n4545) & (x13091x) & (x22134x)) + ((!n_n4548) & (n_n4551) & (n_n4545) & (!x13091x) & (!x22134x)) + ((!n_n4548) & (n_n4551) & (n_n4545) & (!x13091x) & (x22134x)) + ((!n_n4548) & (n_n4551) & (n_n4545) & (x13091x) & (!x22134x)) + ((!n_n4548) & (n_n4551) & (n_n4545) & (x13091x) & (x22134x)) + ((n_n4548) & (!n_n4551) & (!n_n4545) & (!x13091x) & (!x22134x)) + ((n_n4548) & (!n_n4551) & (!n_n4545) & (!x13091x) & (x22134x)) + ((n_n4548) & (!n_n4551) & (!n_n4545) & (x13091x) & (!x22134x)) + ((n_n4548) & (!n_n4551) & (!n_n4545) & (x13091x) & (x22134x)) + ((n_n4548) & (!n_n4551) & (n_n4545) & (!x13091x) & (!x22134x)) + ((n_n4548) & (!n_n4551) & (n_n4545) & (!x13091x) & (x22134x)) + ((n_n4548) & (!n_n4551) & (n_n4545) & (x13091x) & (!x22134x)) + ((n_n4548) & (!n_n4551) & (n_n4545) & (x13091x) & (x22134x)) + ((n_n4548) & (n_n4551) & (!n_n4545) & (!x13091x) & (!x22134x)) + ((n_n4548) & (n_n4551) & (!n_n4545) & (!x13091x) & (x22134x)) + ((n_n4548) & (n_n4551) & (!n_n4545) & (x13091x) & (!x22134x)) + ((n_n4548) & (n_n4551) & (!n_n4545) & (x13091x) & (x22134x)) + ((n_n4548) & (n_n4551) & (n_n4545) & (!x13091x) & (!x22134x)) + ((n_n4548) & (n_n4551) & (n_n4545) & (!x13091x) & (x22134x)) + ((n_n4548) & (n_n4551) & (n_n4545) & (x13091x) & (!x22134x)) + ((n_n4548) & (n_n4551) & (n_n4545) & (x13091x) & (x22134x)));
	assign x12804x = (((!i_9_) & (n_n390) & (n_n473) & (!n_n532) & (n_n534)) + ((!i_9_) & (n_n390) & (n_n473) & (n_n532) & (!n_n534)) + ((!i_9_) & (n_n390) & (n_n473) & (n_n532) & (n_n534)) + ((i_9_) & (n_n390) & (n_n473) & (!n_n532) & (n_n534)) + ((i_9_) & (n_n390) & (n_n473) & (n_n532) & (!n_n534)) + ((i_9_) & (n_n390) & (n_n473) & (n_n532) & (n_n534)));
	assign x13060x = (((!n_n4359) & (!n_n4357) & (!n_n4358) & (!n_n4354) & (n_n4349)) + ((!n_n4359) & (!n_n4357) & (!n_n4358) & (n_n4354) & (!n_n4349)) + ((!n_n4359) & (!n_n4357) & (!n_n4358) & (n_n4354) & (n_n4349)) + ((!n_n4359) & (!n_n4357) & (n_n4358) & (!n_n4354) & (!n_n4349)) + ((!n_n4359) & (!n_n4357) & (n_n4358) & (!n_n4354) & (n_n4349)) + ((!n_n4359) & (!n_n4357) & (n_n4358) & (n_n4354) & (!n_n4349)) + ((!n_n4359) & (!n_n4357) & (n_n4358) & (n_n4354) & (n_n4349)) + ((!n_n4359) & (n_n4357) & (!n_n4358) & (!n_n4354) & (!n_n4349)) + ((!n_n4359) & (n_n4357) & (!n_n4358) & (!n_n4354) & (n_n4349)) + ((!n_n4359) & (n_n4357) & (!n_n4358) & (n_n4354) & (!n_n4349)) + ((!n_n4359) & (n_n4357) & (!n_n4358) & (n_n4354) & (n_n4349)) + ((!n_n4359) & (n_n4357) & (n_n4358) & (!n_n4354) & (!n_n4349)) + ((!n_n4359) & (n_n4357) & (n_n4358) & (!n_n4354) & (n_n4349)) + ((!n_n4359) & (n_n4357) & (n_n4358) & (n_n4354) & (!n_n4349)) + ((!n_n4359) & (n_n4357) & (n_n4358) & (n_n4354) & (n_n4349)) + ((n_n4359) & (!n_n4357) & (!n_n4358) & (!n_n4354) & (!n_n4349)) + ((n_n4359) & (!n_n4357) & (!n_n4358) & (!n_n4354) & (n_n4349)) + ((n_n4359) & (!n_n4357) & (!n_n4358) & (n_n4354) & (!n_n4349)) + ((n_n4359) & (!n_n4357) & (!n_n4358) & (n_n4354) & (n_n4349)) + ((n_n4359) & (!n_n4357) & (n_n4358) & (!n_n4354) & (!n_n4349)) + ((n_n4359) & (!n_n4357) & (n_n4358) & (!n_n4354) & (n_n4349)) + ((n_n4359) & (!n_n4357) & (n_n4358) & (n_n4354) & (!n_n4349)) + ((n_n4359) & (!n_n4357) & (n_n4358) & (n_n4354) & (n_n4349)) + ((n_n4359) & (n_n4357) & (!n_n4358) & (!n_n4354) & (!n_n4349)) + ((n_n4359) & (n_n4357) & (!n_n4358) & (!n_n4354) & (n_n4349)) + ((n_n4359) & (n_n4357) & (!n_n4358) & (n_n4354) & (!n_n4349)) + ((n_n4359) & (n_n4357) & (!n_n4358) & (n_n4354) & (n_n4349)) + ((n_n4359) & (n_n4357) & (n_n4358) & (!n_n4354) & (!n_n4349)) + ((n_n4359) & (n_n4357) & (n_n4358) & (!n_n4354) & (n_n4349)) + ((n_n4359) & (n_n4357) & (n_n4358) & (n_n4354) & (!n_n4349)) + ((n_n4359) & (n_n4357) & (n_n4358) & (n_n4354) & (n_n4349)));
	assign x13065x = (((!n_n4361) & (!n_n4370) & (!n_n4275) & (!n_n3176) & (x13056x)) + ((!n_n4361) & (!n_n4370) & (!n_n4275) & (n_n3176) & (!x13056x)) + ((!n_n4361) & (!n_n4370) & (!n_n4275) & (n_n3176) & (x13056x)) + ((!n_n4361) & (!n_n4370) & (n_n4275) & (!n_n3176) & (!x13056x)) + ((!n_n4361) & (!n_n4370) & (n_n4275) & (!n_n3176) & (x13056x)) + ((!n_n4361) & (!n_n4370) & (n_n4275) & (n_n3176) & (!x13056x)) + ((!n_n4361) & (!n_n4370) & (n_n4275) & (n_n3176) & (x13056x)) + ((!n_n4361) & (n_n4370) & (!n_n4275) & (!n_n3176) & (!x13056x)) + ((!n_n4361) & (n_n4370) & (!n_n4275) & (!n_n3176) & (x13056x)) + ((!n_n4361) & (n_n4370) & (!n_n4275) & (n_n3176) & (!x13056x)) + ((!n_n4361) & (n_n4370) & (!n_n4275) & (n_n3176) & (x13056x)) + ((!n_n4361) & (n_n4370) & (n_n4275) & (!n_n3176) & (!x13056x)) + ((!n_n4361) & (n_n4370) & (n_n4275) & (!n_n3176) & (x13056x)) + ((!n_n4361) & (n_n4370) & (n_n4275) & (n_n3176) & (!x13056x)) + ((!n_n4361) & (n_n4370) & (n_n4275) & (n_n3176) & (x13056x)) + ((n_n4361) & (!n_n4370) & (!n_n4275) & (!n_n3176) & (!x13056x)) + ((n_n4361) & (!n_n4370) & (!n_n4275) & (!n_n3176) & (x13056x)) + ((n_n4361) & (!n_n4370) & (!n_n4275) & (n_n3176) & (!x13056x)) + ((n_n4361) & (!n_n4370) & (!n_n4275) & (n_n3176) & (x13056x)) + ((n_n4361) & (!n_n4370) & (n_n4275) & (!n_n3176) & (!x13056x)) + ((n_n4361) & (!n_n4370) & (n_n4275) & (!n_n3176) & (x13056x)) + ((n_n4361) & (!n_n4370) & (n_n4275) & (n_n3176) & (!x13056x)) + ((n_n4361) & (!n_n4370) & (n_n4275) & (n_n3176) & (x13056x)) + ((n_n4361) & (n_n4370) & (!n_n4275) & (!n_n3176) & (!x13056x)) + ((n_n4361) & (n_n4370) & (!n_n4275) & (!n_n3176) & (x13056x)) + ((n_n4361) & (n_n4370) & (!n_n4275) & (n_n3176) & (!x13056x)) + ((n_n4361) & (n_n4370) & (!n_n4275) & (n_n3176) & (x13056x)) + ((n_n4361) & (n_n4370) & (n_n4275) & (!n_n3176) & (!x13056x)) + ((n_n4361) & (n_n4370) & (n_n4275) & (!n_n3176) & (x13056x)) + ((n_n4361) & (n_n4370) & (n_n4275) & (n_n3176) & (!x13056x)) + ((n_n4361) & (n_n4370) & (n_n4275) & (n_n3176) & (x13056x)));
	assign x13064x = (((!n_n4373) & (!n_n4362) & (!n_n4374) & (!n_n4360) & (x27x)) + ((!n_n4373) & (!n_n4362) & (!n_n4374) & (n_n4360) & (!x27x)) + ((!n_n4373) & (!n_n4362) & (!n_n4374) & (n_n4360) & (x27x)) + ((!n_n4373) & (!n_n4362) & (n_n4374) & (!n_n4360) & (!x27x)) + ((!n_n4373) & (!n_n4362) & (n_n4374) & (!n_n4360) & (x27x)) + ((!n_n4373) & (!n_n4362) & (n_n4374) & (n_n4360) & (!x27x)) + ((!n_n4373) & (!n_n4362) & (n_n4374) & (n_n4360) & (x27x)) + ((!n_n4373) & (n_n4362) & (!n_n4374) & (!n_n4360) & (!x27x)) + ((!n_n4373) & (n_n4362) & (!n_n4374) & (!n_n4360) & (x27x)) + ((!n_n4373) & (n_n4362) & (!n_n4374) & (n_n4360) & (!x27x)) + ((!n_n4373) & (n_n4362) & (!n_n4374) & (n_n4360) & (x27x)) + ((!n_n4373) & (n_n4362) & (n_n4374) & (!n_n4360) & (!x27x)) + ((!n_n4373) & (n_n4362) & (n_n4374) & (!n_n4360) & (x27x)) + ((!n_n4373) & (n_n4362) & (n_n4374) & (n_n4360) & (!x27x)) + ((!n_n4373) & (n_n4362) & (n_n4374) & (n_n4360) & (x27x)) + ((n_n4373) & (!n_n4362) & (!n_n4374) & (!n_n4360) & (!x27x)) + ((n_n4373) & (!n_n4362) & (!n_n4374) & (!n_n4360) & (x27x)) + ((n_n4373) & (!n_n4362) & (!n_n4374) & (n_n4360) & (!x27x)) + ((n_n4373) & (!n_n4362) & (!n_n4374) & (n_n4360) & (x27x)) + ((n_n4373) & (!n_n4362) & (n_n4374) & (!n_n4360) & (!x27x)) + ((n_n4373) & (!n_n4362) & (n_n4374) & (!n_n4360) & (x27x)) + ((n_n4373) & (!n_n4362) & (n_n4374) & (n_n4360) & (!x27x)) + ((n_n4373) & (!n_n4362) & (n_n4374) & (n_n4360) & (x27x)) + ((n_n4373) & (n_n4362) & (!n_n4374) & (!n_n4360) & (!x27x)) + ((n_n4373) & (n_n4362) & (!n_n4374) & (!n_n4360) & (x27x)) + ((n_n4373) & (n_n4362) & (!n_n4374) & (n_n4360) & (!x27x)) + ((n_n4373) & (n_n4362) & (!n_n4374) & (n_n4360) & (x27x)) + ((n_n4373) & (n_n4362) & (n_n4374) & (!n_n4360) & (!x27x)) + ((n_n4373) & (n_n4362) & (n_n4374) & (!n_n4360) & (x27x)) + ((n_n4373) & (n_n4362) & (n_n4374) & (n_n4360) & (!x27x)) + ((n_n4373) & (n_n4362) & (n_n4374) & (n_n4360) & (x27x)));
	assign x13074x = (((!n_n4383) & (!n_n4388) & (!n_n4396) & (n_n4395)) + ((!n_n4383) & (!n_n4388) & (n_n4396) & (!n_n4395)) + ((!n_n4383) & (!n_n4388) & (n_n4396) & (n_n4395)) + ((!n_n4383) & (n_n4388) & (!n_n4396) & (!n_n4395)) + ((!n_n4383) & (n_n4388) & (!n_n4396) & (n_n4395)) + ((!n_n4383) & (n_n4388) & (n_n4396) & (!n_n4395)) + ((!n_n4383) & (n_n4388) & (n_n4396) & (n_n4395)) + ((n_n4383) & (!n_n4388) & (!n_n4396) & (!n_n4395)) + ((n_n4383) & (!n_n4388) & (!n_n4396) & (n_n4395)) + ((n_n4383) & (!n_n4388) & (n_n4396) & (!n_n4395)) + ((n_n4383) & (!n_n4388) & (n_n4396) & (n_n4395)) + ((n_n4383) & (n_n4388) & (!n_n4396) & (!n_n4395)) + ((n_n4383) & (n_n4388) & (!n_n4396) & (n_n4395)) + ((n_n4383) & (n_n4388) & (n_n4396) & (!n_n4395)) + ((n_n4383) & (n_n4388) & (n_n4396) & (n_n4395)));
	assign x13075x = (((!n_n4389) & (!n_n4393) & (!n_n4390) & (!n_n4394) & (n_n4386)) + ((!n_n4389) & (!n_n4393) & (!n_n4390) & (n_n4394) & (!n_n4386)) + ((!n_n4389) & (!n_n4393) & (!n_n4390) & (n_n4394) & (n_n4386)) + ((!n_n4389) & (!n_n4393) & (n_n4390) & (!n_n4394) & (!n_n4386)) + ((!n_n4389) & (!n_n4393) & (n_n4390) & (!n_n4394) & (n_n4386)) + ((!n_n4389) & (!n_n4393) & (n_n4390) & (n_n4394) & (!n_n4386)) + ((!n_n4389) & (!n_n4393) & (n_n4390) & (n_n4394) & (n_n4386)) + ((!n_n4389) & (n_n4393) & (!n_n4390) & (!n_n4394) & (!n_n4386)) + ((!n_n4389) & (n_n4393) & (!n_n4390) & (!n_n4394) & (n_n4386)) + ((!n_n4389) & (n_n4393) & (!n_n4390) & (n_n4394) & (!n_n4386)) + ((!n_n4389) & (n_n4393) & (!n_n4390) & (n_n4394) & (n_n4386)) + ((!n_n4389) & (n_n4393) & (n_n4390) & (!n_n4394) & (!n_n4386)) + ((!n_n4389) & (n_n4393) & (n_n4390) & (!n_n4394) & (n_n4386)) + ((!n_n4389) & (n_n4393) & (n_n4390) & (n_n4394) & (!n_n4386)) + ((!n_n4389) & (n_n4393) & (n_n4390) & (n_n4394) & (n_n4386)) + ((n_n4389) & (!n_n4393) & (!n_n4390) & (!n_n4394) & (!n_n4386)) + ((n_n4389) & (!n_n4393) & (!n_n4390) & (!n_n4394) & (n_n4386)) + ((n_n4389) & (!n_n4393) & (!n_n4390) & (n_n4394) & (!n_n4386)) + ((n_n4389) & (!n_n4393) & (!n_n4390) & (n_n4394) & (n_n4386)) + ((n_n4389) & (!n_n4393) & (n_n4390) & (!n_n4394) & (!n_n4386)) + ((n_n4389) & (!n_n4393) & (n_n4390) & (!n_n4394) & (n_n4386)) + ((n_n4389) & (!n_n4393) & (n_n4390) & (n_n4394) & (!n_n4386)) + ((n_n4389) & (!n_n4393) & (n_n4390) & (n_n4394) & (n_n4386)) + ((n_n4389) & (n_n4393) & (!n_n4390) & (!n_n4394) & (!n_n4386)) + ((n_n4389) & (n_n4393) & (!n_n4390) & (!n_n4394) & (n_n4386)) + ((n_n4389) & (n_n4393) & (!n_n4390) & (n_n4394) & (!n_n4386)) + ((n_n4389) & (n_n4393) & (!n_n4390) & (n_n4394) & (n_n4386)) + ((n_n4389) & (n_n4393) & (n_n4390) & (!n_n4394) & (!n_n4386)) + ((n_n4389) & (n_n4393) & (n_n4390) & (!n_n4394) & (n_n4386)) + ((n_n4389) & (n_n4393) & (n_n4390) & (n_n4394) & (!n_n4386)) + ((n_n4389) & (n_n4393) & (n_n4390) & (n_n4394) & (n_n4386)));
	assign x13079x = (((!n_n4401) & (!n_n4400) & (!n_n4407) & (!n_n4405) & (n_n4402)) + ((!n_n4401) & (!n_n4400) & (!n_n4407) & (n_n4405) & (!n_n4402)) + ((!n_n4401) & (!n_n4400) & (!n_n4407) & (n_n4405) & (n_n4402)) + ((!n_n4401) & (!n_n4400) & (n_n4407) & (!n_n4405) & (!n_n4402)) + ((!n_n4401) & (!n_n4400) & (n_n4407) & (!n_n4405) & (n_n4402)) + ((!n_n4401) & (!n_n4400) & (n_n4407) & (n_n4405) & (!n_n4402)) + ((!n_n4401) & (!n_n4400) & (n_n4407) & (n_n4405) & (n_n4402)) + ((!n_n4401) & (n_n4400) & (!n_n4407) & (!n_n4405) & (!n_n4402)) + ((!n_n4401) & (n_n4400) & (!n_n4407) & (!n_n4405) & (n_n4402)) + ((!n_n4401) & (n_n4400) & (!n_n4407) & (n_n4405) & (!n_n4402)) + ((!n_n4401) & (n_n4400) & (!n_n4407) & (n_n4405) & (n_n4402)) + ((!n_n4401) & (n_n4400) & (n_n4407) & (!n_n4405) & (!n_n4402)) + ((!n_n4401) & (n_n4400) & (n_n4407) & (!n_n4405) & (n_n4402)) + ((!n_n4401) & (n_n4400) & (n_n4407) & (n_n4405) & (!n_n4402)) + ((!n_n4401) & (n_n4400) & (n_n4407) & (n_n4405) & (n_n4402)) + ((n_n4401) & (!n_n4400) & (!n_n4407) & (!n_n4405) & (!n_n4402)) + ((n_n4401) & (!n_n4400) & (!n_n4407) & (!n_n4405) & (n_n4402)) + ((n_n4401) & (!n_n4400) & (!n_n4407) & (n_n4405) & (!n_n4402)) + ((n_n4401) & (!n_n4400) & (!n_n4407) & (n_n4405) & (n_n4402)) + ((n_n4401) & (!n_n4400) & (n_n4407) & (!n_n4405) & (!n_n4402)) + ((n_n4401) & (!n_n4400) & (n_n4407) & (!n_n4405) & (n_n4402)) + ((n_n4401) & (!n_n4400) & (n_n4407) & (n_n4405) & (!n_n4402)) + ((n_n4401) & (!n_n4400) & (n_n4407) & (n_n4405) & (n_n4402)) + ((n_n4401) & (n_n4400) & (!n_n4407) & (!n_n4405) & (!n_n4402)) + ((n_n4401) & (n_n4400) & (!n_n4407) & (!n_n4405) & (n_n4402)) + ((n_n4401) & (n_n4400) & (!n_n4407) & (n_n4405) & (!n_n4402)) + ((n_n4401) & (n_n4400) & (!n_n4407) & (n_n4405) & (n_n4402)) + ((n_n4401) & (n_n4400) & (n_n4407) & (!n_n4405) & (!n_n4402)) + ((n_n4401) & (n_n4400) & (n_n4407) & (!n_n4405) & (n_n4402)) + ((n_n4401) & (n_n4400) & (n_n4407) & (n_n4405) & (!n_n4402)) + ((n_n4401) & (n_n4400) & (n_n4407) & (n_n4405) & (n_n4402)));
	assign x13080x = (((!n_n4406) & (!n_n4397) & (!n_n4398) & (!n_n4408) & (x13079x)) + ((!n_n4406) & (!n_n4397) & (!n_n4398) & (n_n4408) & (!x13079x)) + ((!n_n4406) & (!n_n4397) & (!n_n4398) & (n_n4408) & (x13079x)) + ((!n_n4406) & (!n_n4397) & (n_n4398) & (!n_n4408) & (!x13079x)) + ((!n_n4406) & (!n_n4397) & (n_n4398) & (!n_n4408) & (x13079x)) + ((!n_n4406) & (!n_n4397) & (n_n4398) & (n_n4408) & (!x13079x)) + ((!n_n4406) & (!n_n4397) & (n_n4398) & (n_n4408) & (x13079x)) + ((!n_n4406) & (n_n4397) & (!n_n4398) & (!n_n4408) & (!x13079x)) + ((!n_n4406) & (n_n4397) & (!n_n4398) & (!n_n4408) & (x13079x)) + ((!n_n4406) & (n_n4397) & (!n_n4398) & (n_n4408) & (!x13079x)) + ((!n_n4406) & (n_n4397) & (!n_n4398) & (n_n4408) & (x13079x)) + ((!n_n4406) & (n_n4397) & (n_n4398) & (!n_n4408) & (!x13079x)) + ((!n_n4406) & (n_n4397) & (n_n4398) & (!n_n4408) & (x13079x)) + ((!n_n4406) & (n_n4397) & (n_n4398) & (n_n4408) & (!x13079x)) + ((!n_n4406) & (n_n4397) & (n_n4398) & (n_n4408) & (x13079x)) + ((n_n4406) & (!n_n4397) & (!n_n4398) & (!n_n4408) & (!x13079x)) + ((n_n4406) & (!n_n4397) & (!n_n4398) & (!n_n4408) & (x13079x)) + ((n_n4406) & (!n_n4397) & (!n_n4398) & (n_n4408) & (!x13079x)) + ((n_n4406) & (!n_n4397) & (!n_n4398) & (n_n4408) & (x13079x)) + ((n_n4406) & (!n_n4397) & (n_n4398) & (!n_n4408) & (!x13079x)) + ((n_n4406) & (!n_n4397) & (n_n4398) & (!n_n4408) & (x13079x)) + ((n_n4406) & (!n_n4397) & (n_n4398) & (n_n4408) & (!x13079x)) + ((n_n4406) & (!n_n4397) & (n_n4398) & (n_n4408) & (x13079x)) + ((n_n4406) & (n_n4397) & (!n_n4398) & (!n_n4408) & (!x13079x)) + ((n_n4406) & (n_n4397) & (!n_n4398) & (!n_n4408) & (x13079x)) + ((n_n4406) & (n_n4397) & (!n_n4398) & (n_n4408) & (!x13079x)) + ((n_n4406) & (n_n4397) & (!n_n4398) & (n_n4408) & (x13079x)) + ((n_n4406) & (n_n4397) & (n_n4398) & (!n_n4408) & (!x13079x)) + ((n_n4406) & (n_n4397) & (n_n4398) & (!n_n4408) & (x13079x)) + ((n_n4406) & (n_n4397) & (n_n4398) & (n_n4408) & (!x13079x)) + ((n_n4406) & (n_n4397) & (n_n4398) & (n_n4408) & (x13079x)));
	assign x13085x = (((!n_n4339) & (!n_n4344) & (!n_n4343) & (!n_n4342) & (n_n4348)) + ((!n_n4339) & (!n_n4344) & (!n_n4343) & (n_n4342) & (!n_n4348)) + ((!n_n4339) & (!n_n4344) & (!n_n4343) & (n_n4342) & (n_n4348)) + ((!n_n4339) & (!n_n4344) & (n_n4343) & (!n_n4342) & (!n_n4348)) + ((!n_n4339) & (!n_n4344) & (n_n4343) & (!n_n4342) & (n_n4348)) + ((!n_n4339) & (!n_n4344) & (n_n4343) & (n_n4342) & (!n_n4348)) + ((!n_n4339) & (!n_n4344) & (n_n4343) & (n_n4342) & (n_n4348)) + ((!n_n4339) & (n_n4344) & (!n_n4343) & (!n_n4342) & (!n_n4348)) + ((!n_n4339) & (n_n4344) & (!n_n4343) & (!n_n4342) & (n_n4348)) + ((!n_n4339) & (n_n4344) & (!n_n4343) & (n_n4342) & (!n_n4348)) + ((!n_n4339) & (n_n4344) & (!n_n4343) & (n_n4342) & (n_n4348)) + ((!n_n4339) & (n_n4344) & (n_n4343) & (!n_n4342) & (!n_n4348)) + ((!n_n4339) & (n_n4344) & (n_n4343) & (!n_n4342) & (n_n4348)) + ((!n_n4339) & (n_n4344) & (n_n4343) & (n_n4342) & (!n_n4348)) + ((!n_n4339) & (n_n4344) & (n_n4343) & (n_n4342) & (n_n4348)) + ((n_n4339) & (!n_n4344) & (!n_n4343) & (!n_n4342) & (!n_n4348)) + ((n_n4339) & (!n_n4344) & (!n_n4343) & (!n_n4342) & (n_n4348)) + ((n_n4339) & (!n_n4344) & (!n_n4343) & (n_n4342) & (!n_n4348)) + ((n_n4339) & (!n_n4344) & (!n_n4343) & (n_n4342) & (n_n4348)) + ((n_n4339) & (!n_n4344) & (n_n4343) & (!n_n4342) & (!n_n4348)) + ((n_n4339) & (!n_n4344) & (n_n4343) & (!n_n4342) & (n_n4348)) + ((n_n4339) & (!n_n4344) & (n_n4343) & (n_n4342) & (!n_n4348)) + ((n_n4339) & (!n_n4344) & (n_n4343) & (n_n4342) & (n_n4348)) + ((n_n4339) & (n_n4344) & (!n_n4343) & (!n_n4342) & (!n_n4348)) + ((n_n4339) & (n_n4344) & (!n_n4343) & (!n_n4342) & (n_n4348)) + ((n_n4339) & (n_n4344) & (!n_n4343) & (n_n4342) & (!n_n4348)) + ((n_n4339) & (n_n4344) & (!n_n4343) & (n_n4342) & (n_n4348)) + ((n_n4339) & (n_n4344) & (n_n4343) & (!n_n4342) & (!n_n4348)) + ((n_n4339) & (n_n4344) & (n_n4343) & (!n_n4342) & (n_n4348)) + ((n_n4339) & (n_n4344) & (n_n4343) & (n_n4342) & (!n_n4348)) + ((n_n4339) & (n_n4344) & (n_n4343) & (n_n4342) & (n_n4348)));
	assign n_n715 = (((!n_n4598) & (!n_n4593) & (!n_n4594) & (!n_n4600) & (x13102x)) + ((!n_n4598) & (!n_n4593) & (!n_n4594) & (n_n4600) & (!x13102x)) + ((!n_n4598) & (!n_n4593) & (!n_n4594) & (n_n4600) & (x13102x)) + ((!n_n4598) & (!n_n4593) & (n_n4594) & (!n_n4600) & (!x13102x)) + ((!n_n4598) & (!n_n4593) & (n_n4594) & (!n_n4600) & (x13102x)) + ((!n_n4598) & (!n_n4593) & (n_n4594) & (n_n4600) & (!x13102x)) + ((!n_n4598) & (!n_n4593) & (n_n4594) & (n_n4600) & (x13102x)) + ((!n_n4598) & (n_n4593) & (!n_n4594) & (!n_n4600) & (!x13102x)) + ((!n_n4598) & (n_n4593) & (!n_n4594) & (!n_n4600) & (x13102x)) + ((!n_n4598) & (n_n4593) & (!n_n4594) & (n_n4600) & (!x13102x)) + ((!n_n4598) & (n_n4593) & (!n_n4594) & (n_n4600) & (x13102x)) + ((!n_n4598) & (n_n4593) & (n_n4594) & (!n_n4600) & (!x13102x)) + ((!n_n4598) & (n_n4593) & (n_n4594) & (!n_n4600) & (x13102x)) + ((!n_n4598) & (n_n4593) & (n_n4594) & (n_n4600) & (!x13102x)) + ((!n_n4598) & (n_n4593) & (n_n4594) & (n_n4600) & (x13102x)) + ((n_n4598) & (!n_n4593) & (!n_n4594) & (!n_n4600) & (!x13102x)) + ((n_n4598) & (!n_n4593) & (!n_n4594) & (!n_n4600) & (x13102x)) + ((n_n4598) & (!n_n4593) & (!n_n4594) & (n_n4600) & (!x13102x)) + ((n_n4598) & (!n_n4593) & (!n_n4594) & (n_n4600) & (x13102x)) + ((n_n4598) & (!n_n4593) & (n_n4594) & (!n_n4600) & (!x13102x)) + ((n_n4598) & (!n_n4593) & (n_n4594) & (!n_n4600) & (x13102x)) + ((n_n4598) & (!n_n4593) & (n_n4594) & (n_n4600) & (!x13102x)) + ((n_n4598) & (!n_n4593) & (n_n4594) & (n_n4600) & (x13102x)) + ((n_n4598) & (n_n4593) & (!n_n4594) & (!n_n4600) & (!x13102x)) + ((n_n4598) & (n_n4593) & (!n_n4594) & (!n_n4600) & (x13102x)) + ((n_n4598) & (n_n4593) & (!n_n4594) & (n_n4600) & (!x13102x)) + ((n_n4598) & (n_n4593) & (!n_n4594) & (n_n4600) & (x13102x)) + ((n_n4598) & (n_n4593) & (n_n4594) & (!n_n4600) & (!x13102x)) + ((n_n4598) & (n_n4593) & (n_n4594) & (!n_n4600) & (x13102x)) + ((n_n4598) & (n_n4593) & (n_n4594) & (n_n4600) & (!x13102x)) + ((n_n4598) & (n_n4593) & (n_n4594) & (n_n4600) & (x13102x)));
	assign x13108x = (((!n_n4571) & (!n_n4582) & (!n_n4574) & (n_n4580)) + ((!n_n4571) & (!n_n4582) & (n_n4574) & (!n_n4580)) + ((!n_n4571) & (!n_n4582) & (n_n4574) & (n_n4580)) + ((!n_n4571) & (n_n4582) & (!n_n4574) & (!n_n4580)) + ((!n_n4571) & (n_n4582) & (!n_n4574) & (n_n4580)) + ((!n_n4571) & (n_n4582) & (n_n4574) & (!n_n4580)) + ((!n_n4571) & (n_n4582) & (n_n4574) & (n_n4580)) + ((n_n4571) & (!n_n4582) & (!n_n4574) & (!n_n4580)) + ((n_n4571) & (!n_n4582) & (!n_n4574) & (n_n4580)) + ((n_n4571) & (!n_n4582) & (n_n4574) & (!n_n4580)) + ((n_n4571) & (!n_n4582) & (n_n4574) & (n_n4580)) + ((n_n4571) & (n_n4582) & (!n_n4574) & (!n_n4580)) + ((n_n4571) & (n_n4582) & (!n_n4574) & (n_n4580)) + ((n_n4571) & (n_n4582) & (n_n4574) & (!n_n4580)) + ((n_n4571) & (n_n4582) & (n_n4574) & (n_n4580)));
	assign x13109x = (((!n_n4570) & (!n_n881) & (!n_n4569) & (x91x)) + ((!n_n4570) & (!n_n881) & (n_n4569) & (!x91x)) + ((!n_n4570) & (!n_n881) & (n_n4569) & (x91x)) + ((!n_n4570) & (n_n881) & (!n_n4569) & (!x91x)) + ((!n_n4570) & (n_n881) & (!n_n4569) & (x91x)) + ((!n_n4570) & (n_n881) & (n_n4569) & (!x91x)) + ((!n_n4570) & (n_n881) & (n_n4569) & (x91x)) + ((n_n4570) & (!n_n881) & (!n_n4569) & (!x91x)) + ((n_n4570) & (!n_n881) & (!n_n4569) & (x91x)) + ((n_n4570) & (!n_n881) & (n_n4569) & (!x91x)) + ((n_n4570) & (!n_n881) & (n_n4569) & (x91x)) + ((n_n4570) & (n_n881) & (!n_n4569) & (!x91x)) + ((n_n4570) & (n_n881) & (!n_n4569) & (x91x)) + ((n_n4570) & (n_n881) & (n_n4569) & (!x91x)) + ((n_n4570) & (n_n881) & (n_n4569) & (x91x)));
	assign x22133x = (((!n_n4577) & (!n_n4576) & (!x100x) & (!x238x) & (!x222x)));
	assign n_n651 = (((!n_n715) & (!x13108x) & (!x13109x) & (!x22133x)) + ((!n_n715) & (!x13108x) & (x13109x) & (!x22133x)) + ((!n_n715) & (!x13108x) & (x13109x) & (x22133x)) + ((!n_n715) & (x13108x) & (!x13109x) & (!x22133x)) + ((!n_n715) & (x13108x) & (!x13109x) & (x22133x)) + ((!n_n715) & (x13108x) & (x13109x) & (!x22133x)) + ((!n_n715) & (x13108x) & (x13109x) & (x22133x)) + ((n_n715) & (!x13108x) & (!x13109x) & (!x22133x)) + ((n_n715) & (!x13108x) & (!x13109x) & (x22133x)) + ((n_n715) & (!x13108x) & (x13109x) & (!x22133x)) + ((n_n715) & (!x13108x) & (x13109x) & (x22133x)) + ((n_n715) & (x13108x) & (!x13109x) & (!x22133x)) + ((n_n715) & (x13108x) & (!x13109x) & (x22133x)) + ((n_n715) & (x13108x) & (x13109x) & (!x22133x)) + ((n_n715) & (x13108x) & (x13109x) & (x22133x)));
	assign n_n714 = (((!n_n4612) & (!n_n4609) & (!n_n4610) & (!x51x) & (n_n2036)) + ((!n_n4612) & (!n_n4609) & (!n_n4610) & (x51x) & (!n_n2036)) + ((!n_n4612) & (!n_n4609) & (!n_n4610) & (x51x) & (n_n2036)) + ((!n_n4612) & (!n_n4609) & (n_n4610) & (!x51x) & (!n_n2036)) + ((!n_n4612) & (!n_n4609) & (n_n4610) & (!x51x) & (n_n2036)) + ((!n_n4612) & (!n_n4609) & (n_n4610) & (x51x) & (!n_n2036)) + ((!n_n4612) & (!n_n4609) & (n_n4610) & (x51x) & (n_n2036)) + ((!n_n4612) & (n_n4609) & (!n_n4610) & (!x51x) & (!n_n2036)) + ((!n_n4612) & (n_n4609) & (!n_n4610) & (!x51x) & (n_n2036)) + ((!n_n4612) & (n_n4609) & (!n_n4610) & (x51x) & (!n_n2036)) + ((!n_n4612) & (n_n4609) & (!n_n4610) & (x51x) & (n_n2036)) + ((!n_n4612) & (n_n4609) & (n_n4610) & (!x51x) & (!n_n2036)) + ((!n_n4612) & (n_n4609) & (n_n4610) & (!x51x) & (n_n2036)) + ((!n_n4612) & (n_n4609) & (n_n4610) & (x51x) & (!n_n2036)) + ((!n_n4612) & (n_n4609) & (n_n4610) & (x51x) & (n_n2036)) + ((n_n4612) & (!n_n4609) & (!n_n4610) & (!x51x) & (!n_n2036)) + ((n_n4612) & (!n_n4609) & (!n_n4610) & (!x51x) & (n_n2036)) + ((n_n4612) & (!n_n4609) & (!n_n4610) & (x51x) & (!n_n2036)) + ((n_n4612) & (!n_n4609) & (!n_n4610) & (x51x) & (n_n2036)) + ((n_n4612) & (!n_n4609) & (n_n4610) & (!x51x) & (!n_n2036)) + ((n_n4612) & (!n_n4609) & (n_n4610) & (!x51x) & (n_n2036)) + ((n_n4612) & (!n_n4609) & (n_n4610) & (x51x) & (!n_n2036)) + ((n_n4612) & (!n_n4609) & (n_n4610) & (x51x) & (n_n2036)) + ((n_n4612) & (n_n4609) & (!n_n4610) & (!x51x) & (!n_n2036)) + ((n_n4612) & (n_n4609) & (!n_n4610) & (!x51x) & (n_n2036)) + ((n_n4612) & (n_n4609) & (!n_n4610) & (x51x) & (!n_n2036)) + ((n_n4612) & (n_n4609) & (!n_n4610) & (x51x) & (n_n2036)) + ((n_n4612) & (n_n4609) & (n_n4610) & (!x51x) & (!n_n2036)) + ((n_n4612) & (n_n4609) & (n_n4610) & (!x51x) & (n_n2036)) + ((n_n4612) & (n_n4609) & (n_n4610) & (x51x) & (!n_n2036)) + ((n_n4612) & (n_n4609) & (n_n4610) & (x51x) & (n_n2036)));
	assign x13120x = (((!n_n4617) & (!n_n4634) & (!n_n4628) & (n_n4640)) + ((!n_n4617) & (!n_n4634) & (n_n4628) & (!n_n4640)) + ((!n_n4617) & (!n_n4634) & (n_n4628) & (n_n4640)) + ((!n_n4617) & (n_n4634) & (!n_n4628) & (!n_n4640)) + ((!n_n4617) & (n_n4634) & (!n_n4628) & (n_n4640)) + ((!n_n4617) & (n_n4634) & (n_n4628) & (!n_n4640)) + ((!n_n4617) & (n_n4634) & (n_n4628) & (n_n4640)) + ((n_n4617) & (!n_n4634) & (!n_n4628) & (!n_n4640)) + ((n_n4617) & (!n_n4634) & (!n_n4628) & (n_n4640)) + ((n_n4617) & (!n_n4634) & (n_n4628) & (!n_n4640)) + ((n_n4617) & (!n_n4634) & (n_n4628) & (n_n4640)) + ((n_n4617) & (n_n4634) & (!n_n4628) & (!n_n4640)) + ((n_n4617) & (n_n4634) & (!n_n4628) & (n_n4640)) + ((n_n4617) & (n_n4634) & (n_n4628) & (!n_n4640)) + ((n_n4617) & (n_n4634) & (n_n4628) & (n_n4640)));
	assign x13121x = (((!n_n4621) & (!x348x) & (!n_n4632) & (!n_n4622) & (x75x)) + ((!n_n4621) & (!x348x) & (!n_n4632) & (n_n4622) & (!x75x)) + ((!n_n4621) & (!x348x) & (!n_n4632) & (n_n4622) & (x75x)) + ((!n_n4621) & (!x348x) & (n_n4632) & (!n_n4622) & (!x75x)) + ((!n_n4621) & (!x348x) & (n_n4632) & (!n_n4622) & (x75x)) + ((!n_n4621) & (!x348x) & (n_n4632) & (n_n4622) & (!x75x)) + ((!n_n4621) & (!x348x) & (n_n4632) & (n_n4622) & (x75x)) + ((!n_n4621) & (x348x) & (!n_n4632) & (!n_n4622) & (!x75x)) + ((!n_n4621) & (x348x) & (!n_n4632) & (!n_n4622) & (x75x)) + ((!n_n4621) & (x348x) & (!n_n4632) & (n_n4622) & (!x75x)) + ((!n_n4621) & (x348x) & (!n_n4632) & (n_n4622) & (x75x)) + ((!n_n4621) & (x348x) & (n_n4632) & (!n_n4622) & (!x75x)) + ((!n_n4621) & (x348x) & (n_n4632) & (!n_n4622) & (x75x)) + ((!n_n4621) & (x348x) & (n_n4632) & (n_n4622) & (!x75x)) + ((!n_n4621) & (x348x) & (n_n4632) & (n_n4622) & (x75x)) + ((n_n4621) & (!x348x) & (!n_n4632) & (!n_n4622) & (!x75x)) + ((n_n4621) & (!x348x) & (!n_n4632) & (!n_n4622) & (x75x)) + ((n_n4621) & (!x348x) & (!n_n4632) & (n_n4622) & (!x75x)) + ((n_n4621) & (!x348x) & (!n_n4632) & (n_n4622) & (x75x)) + ((n_n4621) & (!x348x) & (n_n4632) & (!n_n4622) & (!x75x)) + ((n_n4621) & (!x348x) & (n_n4632) & (!n_n4622) & (x75x)) + ((n_n4621) & (!x348x) & (n_n4632) & (n_n4622) & (!x75x)) + ((n_n4621) & (!x348x) & (n_n4632) & (n_n4622) & (x75x)) + ((n_n4621) & (x348x) & (!n_n4632) & (!n_n4622) & (!x75x)) + ((n_n4621) & (x348x) & (!n_n4632) & (!n_n4622) & (x75x)) + ((n_n4621) & (x348x) & (!n_n4632) & (n_n4622) & (!x75x)) + ((n_n4621) & (x348x) & (!n_n4632) & (n_n4622) & (x75x)) + ((n_n4621) & (x348x) & (n_n4632) & (!n_n4622) & (!x75x)) + ((n_n4621) & (x348x) & (n_n4632) & (!n_n4622) & (x75x)) + ((n_n4621) & (x348x) & (n_n4632) & (n_n4622) & (!x75x)) + ((n_n4621) & (x348x) & (n_n4632) & (n_n4622) & (x75x)));
	assign x13122x = (((!n_n4629) & (!n_n4630) & (!x271x) & (!x190x) & (x270x)) + ((!n_n4629) & (!n_n4630) & (!x271x) & (x190x) & (!x270x)) + ((!n_n4629) & (!n_n4630) & (!x271x) & (x190x) & (x270x)) + ((!n_n4629) & (!n_n4630) & (x271x) & (!x190x) & (!x270x)) + ((!n_n4629) & (!n_n4630) & (x271x) & (!x190x) & (x270x)) + ((!n_n4629) & (!n_n4630) & (x271x) & (x190x) & (!x270x)) + ((!n_n4629) & (!n_n4630) & (x271x) & (x190x) & (x270x)) + ((!n_n4629) & (n_n4630) & (!x271x) & (!x190x) & (!x270x)) + ((!n_n4629) & (n_n4630) & (!x271x) & (!x190x) & (x270x)) + ((!n_n4629) & (n_n4630) & (!x271x) & (x190x) & (!x270x)) + ((!n_n4629) & (n_n4630) & (!x271x) & (x190x) & (x270x)) + ((!n_n4629) & (n_n4630) & (x271x) & (!x190x) & (!x270x)) + ((!n_n4629) & (n_n4630) & (x271x) & (!x190x) & (x270x)) + ((!n_n4629) & (n_n4630) & (x271x) & (x190x) & (!x270x)) + ((!n_n4629) & (n_n4630) & (x271x) & (x190x) & (x270x)) + ((n_n4629) & (!n_n4630) & (!x271x) & (!x190x) & (!x270x)) + ((n_n4629) & (!n_n4630) & (!x271x) & (!x190x) & (x270x)) + ((n_n4629) & (!n_n4630) & (!x271x) & (x190x) & (!x270x)) + ((n_n4629) & (!n_n4630) & (!x271x) & (x190x) & (x270x)) + ((n_n4629) & (!n_n4630) & (x271x) & (!x190x) & (!x270x)) + ((n_n4629) & (!n_n4630) & (x271x) & (!x190x) & (x270x)) + ((n_n4629) & (!n_n4630) & (x271x) & (x190x) & (!x270x)) + ((n_n4629) & (!n_n4630) & (x271x) & (x190x) & (x270x)) + ((n_n4629) & (n_n4630) & (!x271x) & (!x190x) & (!x270x)) + ((n_n4629) & (n_n4630) & (!x271x) & (!x190x) & (x270x)) + ((n_n4629) & (n_n4630) & (!x271x) & (x190x) & (!x270x)) + ((n_n4629) & (n_n4630) & (!x271x) & (x190x) & (x270x)) + ((n_n4629) & (n_n4630) & (x271x) & (!x190x) & (!x270x)) + ((n_n4629) & (n_n4630) & (x271x) & (!x190x) & (x270x)) + ((n_n4629) & (n_n4630) & (x271x) & (x190x) & (!x270x)) + ((n_n4629) & (n_n4630) & (x271x) & (x190x) & (x270x)));
	assign n_n650 = (((!n_n714) & (!x13120x) & (!x13121x) & (x13122x)) + ((!n_n714) & (!x13120x) & (x13121x) & (!x13122x)) + ((!n_n714) & (!x13120x) & (x13121x) & (x13122x)) + ((!n_n714) & (x13120x) & (!x13121x) & (!x13122x)) + ((!n_n714) & (x13120x) & (!x13121x) & (x13122x)) + ((!n_n714) & (x13120x) & (x13121x) & (!x13122x)) + ((!n_n714) & (x13120x) & (x13121x) & (x13122x)) + ((n_n714) & (!x13120x) & (!x13121x) & (!x13122x)) + ((n_n714) & (!x13120x) & (!x13121x) & (x13122x)) + ((n_n714) & (!x13120x) & (x13121x) & (!x13122x)) + ((n_n714) & (!x13120x) & (x13121x) & (x13122x)) + ((n_n714) & (x13120x) & (!x13121x) & (!x13122x)) + ((n_n714) & (x13120x) & (!x13121x) & (x13122x)) + ((n_n714) & (x13120x) & (x13121x) & (!x13122x)) + ((n_n714) & (x13120x) & (x13121x) & (x13122x)));
	assign x13130x = (((!n_n4561) & (!n_n4532) & (!x178x) & (n_n3875)) + ((!n_n4561) & (!n_n4532) & (x178x) & (!n_n3875)) + ((!n_n4561) & (!n_n4532) & (x178x) & (n_n3875)) + ((!n_n4561) & (n_n4532) & (!x178x) & (!n_n3875)) + ((!n_n4561) & (n_n4532) & (!x178x) & (n_n3875)) + ((!n_n4561) & (n_n4532) & (x178x) & (!n_n3875)) + ((!n_n4561) & (n_n4532) & (x178x) & (n_n3875)) + ((n_n4561) & (!n_n4532) & (!x178x) & (!n_n3875)) + ((n_n4561) & (!n_n4532) & (!x178x) & (n_n3875)) + ((n_n4561) & (!n_n4532) & (x178x) & (!n_n3875)) + ((n_n4561) & (!n_n4532) & (x178x) & (n_n3875)) + ((n_n4561) & (n_n4532) & (!x178x) & (!n_n3875)) + ((n_n4561) & (n_n4532) & (!x178x) & (n_n3875)) + ((n_n4561) & (n_n4532) & (x178x) & (!n_n3875)) + ((n_n4561) & (n_n4532) & (x178x) & (n_n3875)));
	assign x13131x = (((!n_n889) & (!n_n3870) & (!x82x) & (x13126x)) + ((!n_n889) & (!n_n3870) & (x82x) & (!x13126x)) + ((!n_n889) & (!n_n3870) & (x82x) & (x13126x)) + ((!n_n889) & (n_n3870) & (!x82x) & (!x13126x)) + ((!n_n889) & (n_n3870) & (!x82x) & (x13126x)) + ((!n_n889) & (n_n3870) & (x82x) & (!x13126x)) + ((!n_n889) & (n_n3870) & (x82x) & (x13126x)) + ((n_n889) & (!n_n3870) & (!x82x) & (!x13126x)) + ((n_n889) & (!n_n3870) & (!x82x) & (x13126x)) + ((n_n889) & (!n_n3870) & (x82x) & (!x13126x)) + ((n_n889) & (!n_n3870) & (x82x) & (x13126x)) + ((n_n889) & (n_n3870) & (!x82x) & (!x13126x)) + ((n_n889) & (n_n3870) & (!x82x) & (x13126x)) + ((n_n889) & (n_n3870) & (x82x) & (!x13126x)) + ((n_n889) & (n_n3870) & (x82x) & (x13126x)));
	assign x15655x = (((!n_n5281) & (!n_n5272) & (!n_n5279) & (!n_n5283) & (n_n5280)) + ((!n_n5281) & (!n_n5272) & (!n_n5279) & (n_n5283) & (!n_n5280)) + ((!n_n5281) & (!n_n5272) & (!n_n5279) & (n_n5283) & (n_n5280)) + ((!n_n5281) & (!n_n5272) & (n_n5279) & (!n_n5283) & (!n_n5280)) + ((!n_n5281) & (!n_n5272) & (n_n5279) & (!n_n5283) & (n_n5280)) + ((!n_n5281) & (!n_n5272) & (n_n5279) & (n_n5283) & (!n_n5280)) + ((!n_n5281) & (!n_n5272) & (n_n5279) & (n_n5283) & (n_n5280)) + ((!n_n5281) & (n_n5272) & (!n_n5279) & (!n_n5283) & (!n_n5280)) + ((!n_n5281) & (n_n5272) & (!n_n5279) & (!n_n5283) & (n_n5280)) + ((!n_n5281) & (n_n5272) & (!n_n5279) & (n_n5283) & (!n_n5280)) + ((!n_n5281) & (n_n5272) & (!n_n5279) & (n_n5283) & (n_n5280)) + ((!n_n5281) & (n_n5272) & (n_n5279) & (!n_n5283) & (!n_n5280)) + ((!n_n5281) & (n_n5272) & (n_n5279) & (!n_n5283) & (n_n5280)) + ((!n_n5281) & (n_n5272) & (n_n5279) & (n_n5283) & (!n_n5280)) + ((!n_n5281) & (n_n5272) & (n_n5279) & (n_n5283) & (n_n5280)) + ((n_n5281) & (!n_n5272) & (!n_n5279) & (!n_n5283) & (!n_n5280)) + ((n_n5281) & (!n_n5272) & (!n_n5279) & (!n_n5283) & (n_n5280)) + ((n_n5281) & (!n_n5272) & (!n_n5279) & (n_n5283) & (!n_n5280)) + ((n_n5281) & (!n_n5272) & (!n_n5279) & (n_n5283) & (n_n5280)) + ((n_n5281) & (!n_n5272) & (n_n5279) & (!n_n5283) & (!n_n5280)) + ((n_n5281) & (!n_n5272) & (n_n5279) & (!n_n5283) & (n_n5280)) + ((n_n5281) & (!n_n5272) & (n_n5279) & (n_n5283) & (!n_n5280)) + ((n_n5281) & (!n_n5272) & (n_n5279) & (n_n5283) & (n_n5280)) + ((n_n5281) & (n_n5272) & (!n_n5279) & (!n_n5283) & (!n_n5280)) + ((n_n5281) & (n_n5272) & (!n_n5279) & (!n_n5283) & (n_n5280)) + ((n_n5281) & (n_n5272) & (!n_n5279) & (n_n5283) & (!n_n5280)) + ((n_n5281) & (n_n5272) & (!n_n5279) & (n_n5283) & (n_n5280)) + ((n_n5281) & (n_n5272) & (n_n5279) & (!n_n5283) & (!n_n5280)) + ((n_n5281) & (n_n5272) & (n_n5279) & (!n_n5283) & (n_n5280)) + ((n_n5281) & (n_n5272) & (n_n5279) & (n_n5283) & (!n_n5280)) + ((n_n5281) & (n_n5272) & (n_n5279) & (n_n5283) & (n_n5280)));
	assign n_n2939 = (((!x19x) & (!x492x) & (!x572x) & (!x333x) & (x15655x)) + ((!x19x) & (!x492x) & (!x572x) & (x333x) & (!x15655x)) + ((!x19x) & (!x492x) & (!x572x) & (x333x) & (x15655x)) + ((!x19x) & (!x492x) & (x572x) & (!x333x) & (x15655x)) + ((!x19x) & (!x492x) & (x572x) & (x333x) & (!x15655x)) + ((!x19x) & (!x492x) & (x572x) & (x333x) & (x15655x)) + ((!x19x) & (x492x) & (!x572x) & (!x333x) & (x15655x)) + ((!x19x) & (x492x) & (!x572x) & (x333x) & (!x15655x)) + ((!x19x) & (x492x) & (!x572x) & (x333x) & (x15655x)) + ((!x19x) & (x492x) & (x572x) & (!x333x) & (x15655x)) + ((!x19x) & (x492x) & (x572x) & (x333x) & (!x15655x)) + ((!x19x) & (x492x) & (x572x) & (x333x) & (x15655x)) + ((x19x) & (!x492x) & (!x572x) & (!x333x) & (x15655x)) + ((x19x) & (!x492x) & (!x572x) & (x333x) & (!x15655x)) + ((x19x) & (!x492x) & (!x572x) & (x333x) & (x15655x)) + ((x19x) & (!x492x) & (x572x) & (!x333x) & (!x15655x)) + ((x19x) & (!x492x) & (x572x) & (!x333x) & (x15655x)) + ((x19x) & (!x492x) & (x572x) & (x333x) & (!x15655x)) + ((x19x) & (!x492x) & (x572x) & (x333x) & (x15655x)) + ((x19x) & (x492x) & (!x572x) & (!x333x) & (!x15655x)) + ((x19x) & (x492x) & (!x572x) & (!x333x) & (x15655x)) + ((x19x) & (x492x) & (!x572x) & (x333x) & (!x15655x)) + ((x19x) & (x492x) & (!x572x) & (x333x) & (x15655x)) + ((x19x) & (x492x) & (x572x) & (!x333x) & (!x15655x)) + ((x19x) & (x492x) & (x572x) & (!x333x) & (x15655x)) + ((x19x) & (x492x) & (x572x) & (x333x) & (!x15655x)) + ((x19x) & (x492x) & (x572x) & (x333x) & (x15655x)));
	assign x15712x = (((!n_n524) & (!n_n509) & (!x18x) & (!n_n5003) & (x405x)) + ((!n_n524) & (!n_n509) & (!x18x) & (n_n5003) & (!x405x)) + ((!n_n524) & (!n_n509) & (!x18x) & (n_n5003) & (x405x)) + ((!n_n524) & (!n_n509) & (x18x) & (!n_n5003) & (x405x)) + ((!n_n524) & (!n_n509) & (x18x) & (n_n5003) & (!x405x)) + ((!n_n524) & (!n_n509) & (x18x) & (n_n5003) & (x405x)) + ((!n_n524) & (n_n509) & (!x18x) & (!n_n5003) & (x405x)) + ((!n_n524) & (n_n509) & (!x18x) & (n_n5003) & (!x405x)) + ((!n_n524) & (n_n509) & (!x18x) & (n_n5003) & (x405x)) + ((!n_n524) & (n_n509) & (x18x) & (!n_n5003) & (x405x)) + ((!n_n524) & (n_n509) & (x18x) & (n_n5003) & (!x405x)) + ((!n_n524) & (n_n509) & (x18x) & (n_n5003) & (x405x)) + ((n_n524) & (!n_n509) & (!x18x) & (!n_n5003) & (x405x)) + ((n_n524) & (!n_n509) & (!x18x) & (n_n5003) & (!x405x)) + ((n_n524) & (!n_n509) & (!x18x) & (n_n5003) & (x405x)) + ((n_n524) & (!n_n509) & (x18x) & (!n_n5003) & (x405x)) + ((n_n524) & (!n_n509) & (x18x) & (n_n5003) & (!x405x)) + ((n_n524) & (!n_n509) & (x18x) & (n_n5003) & (x405x)) + ((n_n524) & (n_n509) & (!x18x) & (!n_n5003) & (x405x)) + ((n_n524) & (n_n509) & (!x18x) & (n_n5003) & (!x405x)) + ((n_n524) & (n_n509) & (!x18x) & (n_n5003) & (x405x)) + ((n_n524) & (n_n509) & (x18x) & (!n_n5003) & (!x405x)) + ((n_n524) & (n_n509) & (x18x) & (!n_n5003) & (x405x)) + ((n_n524) & (n_n509) & (x18x) & (n_n5003) & (!x405x)) + ((n_n524) & (n_n509) & (x18x) & (n_n5003) & (x405x)));
	assign x15714x = (((!n_n4996) & (!n_n4999) & (!n_n5000) & (!n_n5004) & (x15712x)) + ((!n_n4996) & (!n_n4999) & (!n_n5000) & (n_n5004) & (!x15712x)) + ((!n_n4996) & (!n_n4999) & (!n_n5000) & (n_n5004) & (x15712x)) + ((!n_n4996) & (!n_n4999) & (n_n5000) & (!n_n5004) & (!x15712x)) + ((!n_n4996) & (!n_n4999) & (n_n5000) & (!n_n5004) & (x15712x)) + ((!n_n4996) & (!n_n4999) & (n_n5000) & (n_n5004) & (!x15712x)) + ((!n_n4996) & (!n_n4999) & (n_n5000) & (n_n5004) & (x15712x)) + ((!n_n4996) & (n_n4999) & (!n_n5000) & (!n_n5004) & (!x15712x)) + ((!n_n4996) & (n_n4999) & (!n_n5000) & (!n_n5004) & (x15712x)) + ((!n_n4996) & (n_n4999) & (!n_n5000) & (n_n5004) & (!x15712x)) + ((!n_n4996) & (n_n4999) & (!n_n5000) & (n_n5004) & (x15712x)) + ((!n_n4996) & (n_n4999) & (n_n5000) & (!n_n5004) & (!x15712x)) + ((!n_n4996) & (n_n4999) & (n_n5000) & (!n_n5004) & (x15712x)) + ((!n_n4996) & (n_n4999) & (n_n5000) & (n_n5004) & (!x15712x)) + ((!n_n4996) & (n_n4999) & (n_n5000) & (n_n5004) & (x15712x)) + ((n_n4996) & (!n_n4999) & (!n_n5000) & (!n_n5004) & (!x15712x)) + ((n_n4996) & (!n_n4999) & (!n_n5000) & (!n_n5004) & (x15712x)) + ((n_n4996) & (!n_n4999) & (!n_n5000) & (n_n5004) & (!x15712x)) + ((n_n4996) & (!n_n4999) & (!n_n5000) & (n_n5004) & (x15712x)) + ((n_n4996) & (!n_n4999) & (n_n5000) & (!n_n5004) & (!x15712x)) + ((n_n4996) & (!n_n4999) & (n_n5000) & (!n_n5004) & (x15712x)) + ((n_n4996) & (!n_n4999) & (n_n5000) & (n_n5004) & (!x15712x)) + ((n_n4996) & (!n_n4999) & (n_n5000) & (n_n5004) & (x15712x)) + ((n_n4996) & (n_n4999) & (!n_n5000) & (!n_n5004) & (!x15712x)) + ((n_n4996) & (n_n4999) & (!n_n5000) & (!n_n5004) & (x15712x)) + ((n_n4996) & (n_n4999) & (!n_n5000) & (n_n5004) & (!x15712x)) + ((n_n4996) & (n_n4999) & (!n_n5000) & (n_n5004) & (x15712x)) + ((n_n4996) & (n_n4999) & (n_n5000) & (!n_n5004) & (!x15712x)) + ((n_n4996) & (n_n4999) & (n_n5000) & (!n_n5004) & (x15712x)) + ((n_n4996) & (n_n4999) & (n_n5000) & (n_n5004) & (!x15712x)) + ((n_n4996) & (n_n4999) & (n_n5000) & (n_n5004) & (x15712x)));
	assign x15713x = (((!n_n5006) & (!n_n5007) & (!x247x) & (!x394x) & (x104x)) + ((!n_n5006) & (!n_n5007) & (!x247x) & (x394x) & (!x104x)) + ((!n_n5006) & (!n_n5007) & (!x247x) & (x394x) & (x104x)) + ((!n_n5006) & (!n_n5007) & (x247x) & (!x394x) & (!x104x)) + ((!n_n5006) & (!n_n5007) & (x247x) & (!x394x) & (x104x)) + ((!n_n5006) & (!n_n5007) & (x247x) & (x394x) & (!x104x)) + ((!n_n5006) & (!n_n5007) & (x247x) & (x394x) & (x104x)) + ((!n_n5006) & (n_n5007) & (!x247x) & (!x394x) & (!x104x)) + ((!n_n5006) & (n_n5007) & (!x247x) & (!x394x) & (x104x)) + ((!n_n5006) & (n_n5007) & (!x247x) & (x394x) & (!x104x)) + ((!n_n5006) & (n_n5007) & (!x247x) & (x394x) & (x104x)) + ((!n_n5006) & (n_n5007) & (x247x) & (!x394x) & (!x104x)) + ((!n_n5006) & (n_n5007) & (x247x) & (!x394x) & (x104x)) + ((!n_n5006) & (n_n5007) & (x247x) & (x394x) & (!x104x)) + ((!n_n5006) & (n_n5007) & (x247x) & (x394x) & (x104x)) + ((n_n5006) & (!n_n5007) & (!x247x) & (!x394x) & (!x104x)) + ((n_n5006) & (!n_n5007) & (!x247x) & (!x394x) & (x104x)) + ((n_n5006) & (!n_n5007) & (!x247x) & (x394x) & (!x104x)) + ((n_n5006) & (!n_n5007) & (!x247x) & (x394x) & (x104x)) + ((n_n5006) & (!n_n5007) & (x247x) & (!x394x) & (!x104x)) + ((n_n5006) & (!n_n5007) & (x247x) & (!x394x) & (x104x)) + ((n_n5006) & (!n_n5007) & (x247x) & (x394x) & (!x104x)) + ((n_n5006) & (!n_n5007) & (x247x) & (x394x) & (x104x)) + ((n_n5006) & (n_n5007) & (!x247x) & (!x394x) & (!x104x)) + ((n_n5006) & (n_n5007) & (!x247x) & (!x394x) & (x104x)) + ((n_n5006) & (n_n5007) & (!x247x) & (x394x) & (!x104x)) + ((n_n5006) & (n_n5007) & (!x247x) & (x394x) & (x104x)) + ((n_n5006) & (n_n5007) & (x247x) & (!x394x) & (!x104x)) + ((n_n5006) & (n_n5007) & (x247x) & (!x394x) & (x104x)) + ((n_n5006) & (n_n5007) & (x247x) & (x394x) & (!x104x)) + ((n_n5006) & (n_n5007) & (x247x) & (x394x) & (x104x)));
	assign n_n2917 = (((!x296x) & (!x298x) & (!x15705x) & (!x15714x) & (x15713x)) + ((!x296x) & (!x298x) & (!x15705x) & (x15714x) & (!x15713x)) + ((!x296x) & (!x298x) & (!x15705x) & (x15714x) & (x15713x)) + ((!x296x) & (!x298x) & (x15705x) & (!x15714x) & (!x15713x)) + ((!x296x) & (!x298x) & (x15705x) & (!x15714x) & (x15713x)) + ((!x296x) & (!x298x) & (x15705x) & (x15714x) & (!x15713x)) + ((!x296x) & (!x298x) & (x15705x) & (x15714x) & (x15713x)) + ((!x296x) & (x298x) & (!x15705x) & (!x15714x) & (!x15713x)) + ((!x296x) & (x298x) & (!x15705x) & (!x15714x) & (x15713x)) + ((!x296x) & (x298x) & (!x15705x) & (x15714x) & (!x15713x)) + ((!x296x) & (x298x) & (!x15705x) & (x15714x) & (x15713x)) + ((!x296x) & (x298x) & (x15705x) & (!x15714x) & (!x15713x)) + ((!x296x) & (x298x) & (x15705x) & (!x15714x) & (x15713x)) + ((!x296x) & (x298x) & (x15705x) & (x15714x) & (!x15713x)) + ((!x296x) & (x298x) & (x15705x) & (x15714x) & (x15713x)) + ((x296x) & (!x298x) & (!x15705x) & (!x15714x) & (!x15713x)) + ((x296x) & (!x298x) & (!x15705x) & (!x15714x) & (x15713x)) + ((x296x) & (!x298x) & (!x15705x) & (x15714x) & (!x15713x)) + ((x296x) & (!x298x) & (!x15705x) & (x15714x) & (x15713x)) + ((x296x) & (!x298x) & (x15705x) & (!x15714x) & (!x15713x)) + ((x296x) & (!x298x) & (x15705x) & (!x15714x) & (x15713x)) + ((x296x) & (!x298x) & (x15705x) & (x15714x) & (!x15713x)) + ((x296x) & (!x298x) & (x15705x) & (x15714x) & (x15713x)) + ((x296x) & (x298x) & (!x15705x) & (!x15714x) & (!x15713x)) + ((x296x) & (x298x) & (!x15705x) & (!x15714x) & (x15713x)) + ((x296x) & (x298x) & (!x15705x) & (x15714x) & (!x15713x)) + ((x296x) & (x298x) & (!x15705x) & (x15714x) & (x15713x)) + ((x296x) & (x298x) & (x15705x) & (!x15714x) & (!x15713x)) + ((x296x) & (x298x) & (x15705x) & (!x15714x) & (x15713x)) + ((x296x) & (x298x) & (x15705x) & (x15714x) & (!x15713x)) + ((x296x) & (x298x) & (x15705x) & (x15714x) & (x15713x)));
	assign x15284x = (((!n_n5163) & (!n_n5157) & (!n_n5158) & (!n_n5159) & (n_n5160)) + ((!n_n5163) & (!n_n5157) & (!n_n5158) & (n_n5159) & (!n_n5160)) + ((!n_n5163) & (!n_n5157) & (!n_n5158) & (n_n5159) & (n_n5160)) + ((!n_n5163) & (!n_n5157) & (n_n5158) & (!n_n5159) & (!n_n5160)) + ((!n_n5163) & (!n_n5157) & (n_n5158) & (!n_n5159) & (n_n5160)) + ((!n_n5163) & (!n_n5157) & (n_n5158) & (n_n5159) & (!n_n5160)) + ((!n_n5163) & (!n_n5157) & (n_n5158) & (n_n5159) & (n_n5160)) + ((!n_n5163) & (n_n5157) & (!n_n5158) & (!n_n5159) & (!n_n5160)) + ((!n_n5163) & (n_n5157) & (!n_n5158) & (!n_n5159) & (n_n5160)) + ((!n_n5163) & (n_n5157) & (!n_n5158) & (n_n5159) & (!n_n5160)) + ((!n_n5163) & (n_n5157) & (!n_n5158) & (n_n5159) & (n_n5160)) + ((!n_n5163) & (n_n5157) & (n_n5158) & (!n_n5159) & (!n_n5160)) + ((!n_n5163) & (n_n5157) & (n_n5158) & (!n_n5159) & (n_n5160)) + ((!n_n5163) & (n_n5157) & (n_n5158) & (n_n5159) & (!n_n5160)) + ((!n_n5163) & (n_n5157) & (n_n5158) & (n_n5159) & (n_n5160)) + ((n_n5163) & (!n_n5157) & (!n_n5158) & (!n_n5159) & (!n_n5160)) + ((n_n5163) & (!n_n5157) & (!n_n5158) & (!n_n5159) & (n_n5160)) + ((n_n5163) & (!n_n5157) & (!n_n5158) & (n_n5159) & (!n_n5160)) + ((n_n5163) & (!n_n5157) & (!n_n5158) & (n_n5159) & (n_n5160)) + ((n_n5163) & (!n_n5157) & (n_n5158) & (!n_n5159) & (!n_n5160)) + ((n_n5163) & (!n_n5157) & (n_n5158) & (!n_n5159) & (n_n5160)) + ((n_n5163) & (!n_n5157) & (n_n5158) & (n_n5159) & (!n_n5160)) + ((n_n5163) & (!n_n5157) & (n_n5158) & (n_n5159) & (n_n5160)) + ((n_n5163) & (n_n5157) & (!n_n5158) & (!n_n5159) & (!n_n5160)) + ((n_n5163) & (n_n5157) & (!n_n5158) & (!n_n5159) & (n_n5160)) + ((n_n5163) & (n_n5157) & (!n_n5158) & (n_n5159) & (!n_n5160)) + ((n_n5163) & (n_n5157) & (!n_n5158) & (n_n5159) & (n_n5160)) + ((n_n5163) & (n_n5157) & (n_n5158) & (!n_n5159) & (!n_n5160)) + ((n_n5163) & (n_n5157) & (n_n5158) & (!n_n5159) & (n_n5160)) + ((n_n5163) & (n_n5157) & (n_n5158) & (n_n5159) & (!n_n5160)) + ((n_n5163) & (n_n5157) & (n_n5158) & (n_n5159) & (n_n5160)));
	assign x22158x = (((!n_n4704) & (!n_n4697) & (!n_n4709) & (!n_n4705)));
	assign x11875x = (((!n_n4707) & (!n_n4702) & (!n_n4700) & (!x221x) & (!x22158x)) + ((!n_n4707) & (!n_n4702) & (!n_n4700) & (x221x) & (!x22158x)) + ((!n_n4707) & (!n_n4702) & (!n_n4700) & (x221x) & (x22158x)) + ((!n_n4707) & (!n_n4702) & (n_n4700) & (!x221x) & (!x22158x)) + ((!n_n4707) & (!n_n4702) & (n_n4700) & (!x221x) & (x22158x)) + ((!n_n4707) & (!n_n4702) & (n_n4700) & (x221x) & (!x22158x)) + ((!n_n4707) & (!n_n4702) & (n_n4700) & (x221x) & (x22158x)) + ((!n_n4707) & (n_n4702) & (!n_n4700) & (!x221x) & (!x22158x)) + ((!n_n4707) & (n_n4702) & (!n_n4700) & (!x221x) & (x22158x)) + ((!n_n4707) & (n_n4702) & (!n_n4700) & (x221x) & (!x22158x)) + ((!n_n4707) & (n_n4702) & (!n_n4700) & (x221x) & (x22158x)) + ((!n_n4707) & (n_n4702) & (n_n4700) & (!x221x) & (!x22158x)) + ((!n_n4707) & (n_n4702) & (n_n4700) & (!x221x) & (x22158x)) + ((!n_n4707) & (n_n4702) & (n_n4700) & (x221x) & (!x22158x)) + ((!n_n4707) & (n_n4702) & (n_n4700) & (x221x) & (x22158x)) + ((n_n4707) & (!n_n4702) & (!n_n4700) & (!x221x) & (!x22158x)) + ((n_n4707) & (!n_n4702) & (!n_n4700) & (!x221x) & (x22158x)) + ((n_n4707) & (!n_n4702) & (!n_n4700) & (x221x) & (!x22158x)) + ((n_n4707) & (!n_n4702) & (!n_n4700) & (x221x) & (x22158x)) + ((n_n4707) & (!n_n4702) & (n_n4700) & (!x221x) & (!x22158x)) + ((n_n4707) & (!n_n4702) & (n_n4700) & (!x221x) & (x22158x)) + ((n_n4707) & (!n_n4702) & (n_n4700) & (x221x) & (!x22158x)) + ((n_n4707) & (!n_n4702) & (n_n4700) & (x221x) & (x22158x)) + ((n_n4707) & (n_n4702) & (!n_n4700) & (!x221x) & (!x22158x)) + ((n_n4707) & (n_n4702) & (!n_n4700) & (!x221x) & (x22158x)) + ((n_n4707) & (n_n4702) & (!n_n4700) & (x221x) & (!x22158x)) + ((n_n4707) & (n_n4702) & (!n_n4700) & (x221x) & (x22158x)) + ((n_n4707) & (n_n4702) & (n_n4700) & (!x221x) & (!x22158x)) + ((n_n4707) & (n_n4702) & (n_n4700) & (!x221x) & (x22158x)) + ((n_n4707) & (n_n4702) & (n_n4700) & (x221x) & (!x22158x)) + ((n_n4707) & (n_n4702) & (n_n4700) & (x221x) & (x22158x)));
	assign n_n1032 = (((!n_n1093) & (!x11867x) & (!x11868x) & (x11875x)) + ((!n_n1093) & (!x11867x) & (x11868x) & (!x11875x)) + ((!n_n1093) & (!x11867x) & (x11868x) & (x11875x)) + ((!n_n1093) & (x11867x) & (!x11868x) & (!x11875x)) + ((!n_n1093) & (x11867x) & (!x11868x) & (x11875x)) + ((!n_n1093) & (x11867x) & (x11868x) & (!x11875x)) + ((!n_n1093) & (x11867x) & (x11868x) & (x11875x)) + ((n_n1093) & (!x11867x) & (!x11868x) & (!x11875x)) + ((n_n1093) & (!x11867x) & (!x11868x) & (x11875x)) + ((n_n1093) & (!x11867x) & (x11868x) & (!x11875x)) + ((n_n1093) & (!x11867x) & (x11868x) & (x11875x)) + ((n_n1093) & (x11867x) & (!x11868x) & (!x11875x)) + ((n_n1093) & (x11867x) & (!x11868x) & (x11875x)) + ((n_n1093) & (x11867x) & (x11868x) & (!x11875x)) + ((n_n1093) & (x11867x) & (x11868x) & (x11875x)));
	assign x12791x = (((!n_n4725) & (!n_n4726) & (!n_n4715) & (!n_n4723) & (n_n4721)) + ((!n_n4725) & (!n_n4726) & (!n_n4715) & (n_n4723) & (!n_n4721)) + ((!n_n4725) & (!n_n4726) & (!n_n4715) & (n_n4723) & (n_n4721)) + ((!n_n4725) & (!n_n4726) & (n_n4715) & (!n_n4723) & (!n_n4721)) + ((!n_n4725) & (!n_n4726) & (n_n4715) & (!n_n4723) & (n_n4721)) + ((!n_n4725) & (!n_n4726) & (n_n4715) & (n_n4723) & (!n_n4721)) + ((!n_n4725) & (!n_n4726) & (n_n4715) & (n_n4723) & (n_n4721)) + ((!n_n4725) & (n_n4726) & (!n_n4715) & (!n_n4723) & (!n_n4721)) + ((!n_n4725) & (n_n4726) & (!n_n4715) & (!n_n4723) & (n_n4721)) + ((!n_n4725) & (n_n4726) & (!n_n4715) & (n_n4723) & (!n_n4721)) + ((!n_n4725) & (n_n4726) & (!n_n4715) & (n_n4723) & (n_n4721)) + ((!n_n4725) & (n_n4726) & (n_n4715) & (!n_n4723) & (!n_n4721)) + ((!n_n4725) & (n_n4726) & (n_n4715) & (!n_n4723) & (n_n4721)) + ((!n_n4725) & (n_n4726) & (n_n4715) & (n_n4723) & (!n_n4721)) + ((!n_n4725) & (n_n4726) & (n_n4715) & (n_n4723) & (n_n4721)) + ((n_n4725) & (!n_n4726) & (!n_n4715) & (!n_n4723) & (!n_n4721)) + ((n_n4725) & (!n_n4726) & (!n_n4715) & (!n_n4723) & (n_n4721)) + ((n_n4725) & (!n_n4726) & (!n_n4715) & (n_n4723) & (!n_n4721)) + ((n_n4725) & (!n_n4726) & (!n_n4715) & (n_n4723) & (n_n4721)) + ((n_n4725) & (!n_n4726) & (n_n4715) & (!n_n4723) & (!n_n4721)) + ((n_n4725) & (!n_n4726) & (n_n4715) & (!n_n4723) & (n_n4721)) + ((n_n4725) & (!n_n4726) & (n_n4715) & (n_n4723) & (!n_n4721)) + ((n_n4725) & (!n_n4726) & (n_n4715) & (n_n4723) & (n_n4721)) + ((n_n4725) & (n_n4726) & (!n_n4715) & (!n_n4723) & (!n_n4721)) + ((n_n4725) & (n_n4726) & (!n_n4715) & (!n_n4723) & (n_n4721)) + ((n_n4725) & (n_n4726) & (!n_n4715) & (n_n4723) & (!n_n4721)) + ((n_n4725) & (n_n4726) & (!n_n4715) & (n_n4723) & (n_n4721)) + ((n_n4725) & (n_n4726) & (n_n4715) & (!n_n4723) & (!n_n4721)) + ((n_n4725) & (n_n4726) & (n_n4715) & (!n_n4723) & (n_n4721)) + ((n_n4725) & (n_n4726) & (n_n4715) & (n_n4723) & (!n_n4721)) + ((n_n4725) & (n_n4726) & (n_n4715) & (n_n4723) & (n_n4721)));
	assign x14754x = (((!x11x) & (!n_n535) & (!n_n195) & (!n_n4962) & (n_n4961)) + ((!x11x) & (!n_n535) & (!n_n195) & (n_n4962) & (!n_n4961)) + ((!x11x) & (!n_n535) & (!n_n195) & (n_n4962) & (n_n4961)) + ((!x11x) & (!n_n535) & (n_n195) & (!n_n4962) & (n_n4961)) + ((!x11x) & (!n_n535) & (n_n195) & (n_n4962) & (!n_n4961)) + ((!x11x) & (!n_n535) & (n_n195) & (n_n4962) & (n_n4961)) + ((!x11x) & (n_n535) & (!n_n195) & (!n_n4962) & (n_n4961)) + ((!x11x) & (n_n535) & (!n_n195) & (n_n4962) & (!n_n4961)) + ((!x11x) & (n_n535) & (!n_n195) & (n_n4962) & (n_n4961)) + ((!x11x) & (n_n535) & (n_n195) & (!n_n4962) & (n_n4961)) + ((!x11x) & (n_n535) & (n_n195) & (n_n4962) & (!n_n4961)) + ((!x11x) & (n_n535) & (n_n195) & (n_n4962) & (n_n4961)) + ((x11x) & (!n_n535) & (!n_n195) & (!n_n4962) & (n_n4961)) + ((x11x) & (!n_n535) & (!n_n195) & (n_n4962) & (!n_n4961)) + ((x11x) & (!n_n535) & (!n_n195) & (n_n4962) & (n_n4961)) + ((x11x) & (!n_n535) & (n_n195) & (!n_n4962) & (n_n4961)) + ((x11x) & (!n_n535) & (n_n195) & (n_n4962) & (!n_n4961)) + ((x11x) & (!n_n535) & (n_n195) & (n_n4962) & (n_n4961)) + ((x11x) & (n_n535) & (!n_n195) & (!n_n4962) & (n_n4961)) + ((x11x) & (n_n535) & (!n_n195) & (n_n4962) & (!n_n4961)) + ((x11x) & (n_n535) & (!n_n195) & (n_n4962) & (n_n4961)) + ((x11x) & (n_n535) & (n_n195) & (!n_n4962) & (!n_n4961)) + ((x11x) & (n_n535) & (n_n195) & (!n_n4962) & (n_n4961)) + ((x11x) & (n_n535) & (n_n195) & (n_n4962) & (!n_n4961)) + ((x11x) & (n_n535) & (n_n195) & (n_n4962) & (n_n4961)));
	assign x22109x = (((!n_n4320) & (!n_n4315) & (!n_n4312) & (!n_n4316)));
	assign n_n3740 = (((!n_n4313) & (!n_n4322) & (!n_n4323) & (!x106x) & (!x22109x)) + ((!n_n4313) & (!n_n4322) & (!n_n4323) & (x106x) & (!x22109x)) + ((!n_n4313) & (!n_n4322) & (!n_n4323) & (x106x) & (x22109x)) + ((!n_n4313) & (!n_n4322) & (n_n4323) & (!x106x) & (!x22109x)) + ((!n_n4313) & (!n_n4322) & (n_n4323) & (!x106x) & (x22109x)) + ((!n_n4313) & (!n_n4322) & (n_n4323) & (x106x) & (!x22109x)) + ((!n_n4313) & (!n_n4322) & (n_n4323) & (x106x) & (x22109x)) + ((!n_n4313) & (n_n4322) & (!n_n4323) & (!x106x) & (!x22109x)) + ((!n_n4313) & (n_n4322) & (!n_n4323) & (!x106x) & (x22109x)) + ((!n_n4313) & (n_n4322) & (!n_n4323) & (x106x) & (!x22109x)) + ((!n_n4313) & (n_n4322) & (!n_n4323) & (x106x) & (x22109x)) + ((!n_n4313) & (n_n4322) & (n_n4323) & (!x106x) & (!x22109x)) + ((!n_n4313) & (n_n4322) & (n_n4323) & (!x106x) & (x22109x)) + ((!n_n4313) & (n_n4322) & (n_n4323) & (x106x) & (!x22109x)) + ((!n_n4313) & (n_n4322) & (n_n4323) & (x106x) & (x22109x)) + ((n_n4313) & (!n_n4322) & (!n_n4323) & (!x106x) & (!x22109x)) + ((n_n4313) & (!n_n4322) & (!n_n4323) & (!x106x) & (x22109x)) + ((n_n4313) & (!n_n4322) & (!n_n4323) & (x106x) & (!x22109x)) + ((n_n4313) & (!n_n4322) & (!n_n4323) & (x106x) & (x22109x)) + ((n_n4313) & (!n_n4322) & (n_n4323) & (!x106x) & (!x22109x)) + ((n_n4313) & (!n_n4322) & (n_n4323) & (!x106x) & (x22109x)) + ((n_n4313) & (!n_n4322) & (n_n4323) & (x106x) & (!x22109x)) + ((n_n4313) & (!n_n4322) & (n_n4323) & (x106x) & (x22109x)) + ((n_n4313) & (n_n4322) & (!n_n4323) & (!x106x) & (!x22109x)) + ((n_n4313) & (n_n4322) & (!n_n4323) & (!x106x) & (x22109x)) + ((n_n4313) & (n_n4322) & (!n_n4323) & (x106x) & (!x22109x)) + ((n_n4313) & (n_n4322) & (!n_n4323) & (x106x) & (x22109x)) + ((n_n4313) & (n_n4322) & (n_n4323) & (!x106x) & (!x22109x)) + ((n_n4313) & (n_n4322) & (n_n4323) & (!x106x) & (x22109x)) + ((n_n4313) & (n_n4322) & (n_n4323) & (x106x) & (!x22109x)) + ((n_n4313) & (n_n4322) & (n_n4323) & (x106x) & (x22109x)));
	assign x14486x = (((!n_n4341) & (!n_n4351) & (!n_n4349) & (n_n4334)) + ((!n_n4341) & (!n_n4351) & (n_n4349) & (!n_n4334)) + ((!n_n4341) & (!n_n4351) & (n_n4349) & (n_n4334)) + ((!n_n4341) & (n_n4351) & (!n_n4349) & (!n_n4334)) + ((!n_n4341) & (n_n4351) & (!n_n4349) & (n_n4334)) + ((!n_n4341) & (n_n4351) & (n_n4349) & (!n_n4334)) + ((!n_n4341) & (n_n4351) & (n_n4349) & (n_n4334)) + ((n_n4341) & (!n_n4351) & (!n_n4349) & (!n_n4334)) + ((n_n4341) & (!n_n4351) & (!n_n4349) & (n_n4334)) + ((n_n4341) & (!n_n4351) & (n_n4349) & (!n_n4334)) + ((n_n4341) & (!n_n4351) & (n_n4349) & (n_n4334)) + ((n_n4341) & (n_n4351) & (!n_n4349) & (!n_n4334)) + ((n_n4341) & (n_n4351) & (!n_n4349) & (n_n4334)) + ((n_n4341) & (n_n4351) & (n_n4349) & (!n_n4334)) + ((n_n4341) & (n_n4351) & (n_n4349) & (n_n4334)));
	assign x14488x = (((!n_n4343) & (!x198x) & (!n_n4342) & (x14485x)) + ((!n_n4343) & (!x198x) & (n_n4342) & (!x14485x)) + ((!n_n4343) & (!x198x) & (n_n4342) & (x14485x)) + ((!n_n4343) & (x198x) & (!n_n4342) & (!x14485x)) + ((!n_n4343) & (x198x) & (!n_n4342) & (x14485x)) + ((!n_n4343) & (x198x) & (n_n4342) & (!x14485x)) + ((!n_n4343) & (x198x) & (n_n4342) & (x14485x)) + ((n_n4343) & (!x198x) & (!n_n4342) & (!x14485x)) + ((n_n4343) & (!x198x) & (!n_n4342) & (x14485x)) + ((n_n4343) & (!x198x) & (n_n4342) & (!x14485x)) + ((n_n4343) & (!x198x) & (n_n4342) & (x14485x)) + ((n_n4343) & (x198x) & (!n_n4342) & (!x14485x)) + ((n_n4343) & (x198x) & (!n_n4342) & (x14485x)) + ((n_n4343) & (x198x) & (n_n4342) & (!x14485x)) + ((n_n4343) & (x198x) & (n_n4342) & (x14485x)));
	assign x15657x = (((!x21x) & (!x11x) & (!n_n500) & (!n_n65) & (n_n5266)) + ((!x21x) & (!x11x) & (!n_n500) & (n_n65) & (n_n5266)) + ((!x21x) & (!x11x) & (n_n500) & (!n_n65) & (n_n5266)) + ((!x21x) & (!x11x) & (n_n500) & (n_n65) & (n_n5266)) + ((!x21x) & (x11x) & (!n_n500) & (!n_n65) & (n_n5266)) + ((!x21x) & (x11x) & (!n_n500) & (n_n65) & (n_n5266)) + ((!x21x) & (x11x) & (n_n500) & (!n_n65) & (n_n5266)) + ((!x21x) & (x11x) & (n_n500) & (n_n65) & (!n_n5266)) + ((!x21x) & (x11x) & (n_n500) & (n_n65) & (n_n5266)) + ((x21x) & (!x11x) & (!n_n500) & (!n_n65) & (n_n5266)) + ((x21x) & (!x11x) & (!n_n500) & (n_n65) & (n_n5266)) + ((x21x) & (!x11x) & (n_n500) & (!n_n65) & (n_n5266)) + ((x21x) & (!x11x) & (n_n500) & (n_n65) & (!n_n5266)) + ((x21x) & (!x11x) & (n_n500) & (n_n65) & (n_n5266)) + ((x21x) & (x11x) & (!n_n500) & (!n_n65) & (n_n5266)) + ((x21x) & (x11x) & (!n_n500) & (n_n65) & (n_n5266)) + ((x21x) & (x11x) & (n_n500) & (!n_n65) & (n_n5266)) + ((x21x) & (x11x) & (n_n500) & (n_n65) & (!n_n5266)) + ((x21x) & (x11x) & (n_n500) & (n_n65) & (n_n5266)));
	assign n_n2940 = (((!n_n5268) & (!n_n5271) & (!x205x) & (!x419x) & (x15657x)) + ((!n_n5268) & (!n_n5271) & (!x205x) & (x419x) & (!x15657x)) + ((!n_n5268) & (!n_n5271) & (!x205x) & (x419x) & (x15657x)) + ((!n_n5268) & (!n_n5271) & (x205x) & (!x419x) & (!x15657x)) + ((!n_n5268) & (!n_n5271) & (x205x) & (!x419x) & (x15657x)) + ((!n_n5268) & (!n_n5271) & (x205x) & (x419x) & (!x15657x)) + ((!n_n5268) & (!n_n5271) & (x205x) & (x419x) & (x15657x)) + ((!n_n5268) & (n_n5271) & (!x205x) & (!x419x) & (!x15657x)) + ((!n_n5268) & (n_n5271) & (!x205x) & (!x419x) & (x15657x)) + ((!n_n5268) & (n_n5271) & (!x205x) & (x419x) & (!x15657x)) + ((!n_n5268) & (n_n5271) & (!x205x) & (x419x) & (x15657x)) + ((!n_n5268) & (n_n5271) & (x205x) & (!x419x) & (!x15657x)) + ((!n_n5268) & (n_n5271) & (x205x) & (!x419x) & (x15657x)) + ((!n_n5268) & (n_n5271) & (x205x) & (x419x) & (!x15657x)) + ((!n_n5268) & (n_n5271) & (x205x) & (x419x) & (x15657x)) + ((n_n5268) & (!n_n5271) & (!x205x) & (!x419x) & (!x15657x)) + ((n_n5268) & (!n_n5271) & (!x205x) & (!x419x) & (x15657x)) + ((n_n5268) & (!n_n5271) & (!x205x) & (x419x) & (!x15657x)) + ((n_n5268) & (!n_n5271) & (!x205x) & (x419x) & (x15657x)) + ((n_n5268) & (!n_n5271) & (x205x) & (!x419x) & (!x15657x)) + ((n_n5268) & (!n_n5271) & (x205x) & (!x419x) & (x15657x)) + ((n_n5268) & (!n_n5271) & (x205x) & (x419x) & (!x15657x)) + ((n_n5268) & (!n_n5271) & (x205x) & (x419x) & (x15657x)) + ((n_n5268) & (n_n5271) & (!x205x) & (!x419x) & (!x15657x)) + ((n_n5268) & (n_n5271) & (!x205x) & (!x419x) & (x15657x)) + ((n_n5268) & (n_n5271) & (!x205x) & (x419x) & (!x15657x)) + ((n_n5268) & (n_n5271) & (!x205x) & (x419x) & (x15657x)) + ((n_n5268) & (n_n5271) & (x205x) & (!x419x) & (!x15657x)) + ((n_n5268) & (n_n5271) & (x205x) & (!x419x) & (x15657x)) + ((n_n5268) & (n_n5271) & (x205x) & (x419x) & (!x15657x)) + ((n_n5268) & (n_n5271) & (x205x) & (x419x) & (x15657x)));
	assign x15493x = (((!x15x) & (!n_n390) & (!n_n500) & (!n_n4632) & (n_n1646)) + ((!x15x) & (!n_n390) & (!n_n500) & (n_n4632) & (!n_n1646)) + ((!x15x) & (!n_n390) & (!n_n500) & (n_n4632) & (n_n1646)) + ((!x15x) & (!n_n390) & (n_n500) & (!n_n4632) & (n_n1646)) + ((!x15x) & (!n_n390) & (n_n500) & (n_n4632) & (!n_n1646)) + ((!x15x) & (!n_n390) & (n_n500) & (n_n4632) & (n_n1646)) + ((!x15x) & (n_n390) & (!n_n500) & (!n_n4632) & (n_n1646)) + ((!x15x) & (n_n390) & (!n_n500) & (n_n4632) & (!n_n1646)) + ((!x15x) & (n_n390) & (!n_n500) & (n_n4632) & (n_n1646)) + ((!x15x) & (n_n390) & (n_n500) & (!n_n4632) & (n_n1646)) + ((!x15x) & (n_n390) & (n_n500) & (n_n4632) & (!n_n1646)) + ((!x15x) & (n_n390) & (n_n500) & (n_n4632) & (n_n1646)) + ((x15x) & (!n_n390) & (!n_n500) & (!n_n4632) & (n_n1646)) + ((x15x) & (!n_n390) & (!n_n500) & (n_n4632) & (!n_n1646)) + ((x15x) & (!n_n390) & (!n_n500) & (n_n4632) & (n_n1646)) + ((x15x) & (!n_n390) & (n_n500) & (!n_n4632) & (n_n1646)) + ((x15x) & (!n_n390) & (n_n500) & (n_n4632) & (!n_n1646)) + ((x15x) & (!n_n390) & (n_n500) & (n_n4632) & (n_n1646)) + ((x15x) & (n_n390) & (!n_n500) & (!n_n4632) & (n_n1646)) + ((x15x) & (n_n390) & (!n_n500) & (n_n4632) & (!n_n1646)) + ((x15x) & (n_n390) & (!n_n500) & (n_n4632) & (n_n1646)) + ((x15x) & (n_n390) & (n_n500) & (!n_n4632) & (!n_n1646)) + ((x15x) & (n_n390) & (n_n500) & (!n_n4632) & (n_n1646)) + ((x15x) & (n_n390) & (n_n500) & (n_n4632) & (!n_n1646)) + ((x15x) & (n_n390) & (n_n500) & (n_n4632) & (n_n1646)));
	assign x15719x = (((!n_n4991) & (!n_n4981) & (!n_n4979) & (!n_n4985) & (n_n4978)) + ((!n_n4991) & (!n_n4981) & (!n_n4979) & (n_n4985) & (!n_n4978)) + ((!n_n4991) & (!n_n4981) & (!n_n4979) & (n_n4985) & (n_n4978)) + ((!n_n4991) & (!n_n4981) & (n_n4979) & (!n_n4985) & (!n_n4978)) + ((!n_n4991) & (!n_n4981) & (n_n4979) & (!n_n4985) & (n_n4978)) + ((!n_n4991) & (!n_n4981) & (n_n4979) & (n_n4985) & (!n_n4978)) + ((!n_n4991) & (!n_n4981) & (n_n4979) & (n_n4985) & (n_n4978)) + ((!n_n4991) & (n_n4981) & (!n_n4979) & (!n_n4985) & (!n_n4978)) + ((!n_n4991) & (n_n4981) & (!n_n4979) & (!n_n4985) & (n_n4978)) + ((!n_n4991) & (n_n4981) & (!n_n4979) & (n_n4985) & (!n_n4978)) + ((!n_n4991) & (n_n4981) & (!n_n4979) & (n_n4985) & (n_n4978)) + ((!n_n4991) & (n_n4981) & (n_n4979) & (!n_n4985) & (!n_n4978)) + ((!n_n4991) & (n_n4981) & (n_n4979) & (!n_n4985) & (n_n4978)) + ((!n_n4991) & (n_n4981) & (n_n4979) & (n_n4985) & (!n_n4978)) + ((!n_n4991) & (n_n4981) & (n_n4979) & (n_n4985) & (n_n4978)) + ((n_n4991) & (!n_n4981) & (!n_n4979) & (!n_n4985) & (!n_n4978)) + ((n_n4991) & (!n_n4981) & (!n_n4979) & (!n_n4985) & (n_n4978)) + ((n_n4991) & (!n_n4981) & (!n_n4979) & (n_n4985) & (!n_n4978)) + ((n_n4991) & (!n_n4981) & (!n_n4979) & (n_n4985) & (n_n4978)) + ((n_n4991) & (!n_n4981) & (n_n4979) & (!n_n4985) & (!n_n4978)) + ((n_n4991) & (!n_n4981) & (n_n4979) & (!n_n4985) & (n_n4978)) + ((n_n4991) & (!n_n4981) & (n_n4979) & (n_n4985) & (!n_n4978)) + ((n_n4991) & (!n_n4981) & (n_n4979) & (n_n4985) & (n_n4978)) + ((n_n4991) & (n_n4981) & (!n_n4979) & (!n_n4985) & (!n_n4978)) + ((n_n4991) & (n_n4981) & (!n_n4979) & (!n_n4985) & (n_n4978)) + ((n_n4991) & (n_n4981) & (!n_n4979) & (n_n4985) & (!n_n4978)) + ((n_n4991) & (n_n4981) & (!n_n4979) & (n_n4985) & (n_n4978)) + ((n_n4991) & (n_n4981) & (n_n4979) & (!n_n4985) & (!n_n4978)) + ((n_n4991) & (n_n4981) & (n_n4979) & (!n_n4985) & (n_n4978)) + ((n_n4991) & (n_n4981) & (n_n4979) & (n_n4985) & (!n_n4978)) + ((n_n4991) & (n_n4981) & (n_n4979) & (n_n4985) & (n_n4978)));
	assign n_n2962 = (((!n_n4982) & (!n_n4983) & (!n_n4988) & (!n_n4987) & (x15719x)) + ((!n_n4982) & (!n_n4983) & (!n_n4988) & (n_n4987) & (!x15719x)) + ((!n_n4982) & (!n_n4983) & (!n_n4988) & (n_n4987) & (x15719x)) + ((!n_n4982) & (!n_n4983) & (n_n4988) & (!n_n4987) & (!x15719x)) + ((!n_n4982) & (!n_n4983) & (n_n4988) & (!n_n4987) & (x15719x)) + ((!n_n4982) & (!n_n4983) & (n_n4988) & (n_n4987) & (!x15719x)) + ((!n_n4982) & (!n_n4983) & (n_n4988) & (n_n4987) & (x15719x)) + ((!n_n4982) & (n_n4983) & (!n_n4988) & (!n_n4987) & (!x15719x)) + ((!n_n4982) & (n_n4983) & (!n_n4988) & (!n_n4987) & (x15719x)) + ((!n_n4982) & (n_n4983) & (!n_n4988) & (n_n4987) & (!x15719x)) + ((!n_n4982) & (n_n4983) & (!n_n4988) & (n_n4987) & (x15719x)) + ((!n_n4982) & (n_n4983) & (n_n4988) & (!n_n4987) & (!x15719x)) + ((!n_n4982) & (n_n4983) & (n_n4988) & (!n_n4987) & (x15719x)) + ((!n_n4982) & (n_n4983) & (n_n4988) & (n_n4987) & (!x15719x)) + ((!n_n4982) & (n_n4983) & (n_n4988) & (n_n4987) & (x15719x)) + ((n_n4982) & (!n_n4983) & (!n_n4988) & (!n_n4987) & (!x15719x)) + ((n_n4982) & (!n_n4983) & (!n_n4988) & (!n_n4987) & (x15719x)) + ((n_n4982) & (!n_n4983) & (!n_n4988) & (n_n4987) & (!x15719x)) + ((n_n4982) & (!n_n4983) & (!n_n4988) & (n_n4987) & (x15719x)) + ((n_n4982) & (!n_n4983) & (n_n4988) & (!n_n4987) & (!x15719x)) + ((n_n4982) & (!n_n4983) & (n_n4988) & (!n_n4987) & (x15719x)) + ((n_n4982) & (!n_n4983) & (n_n4988) & (n_n4987) & (!x15719x)) + ((n_n4982) & (!n_n4983) & (n_n4988) & (n_n4987) & (x15719x)) + ((n_n4982) & (n_n4983) & (!n_n4988) & (!n_n4987) & (!x15719x)) + ((n_n4982) & (n_n4983) & (!n_n4988) & (!n_n4987) & (x15719x)) + ((n_n4982) & (n_n4983) & (!n_n4988) & (n_n4987) & (!x15719x)) + ((n_n4982) & (n_n4983) & (!n_n4988) & (n_n4987) & (x15719x)) + ((n_n4982) & (n_n4983) & (n_n4988) & (!n_n4987) & (!x15719x)) + ((n_n4982) & (n_n4983) & (n_n4988) & (!n_n4987) & (x15719x)) + ((n_n4982) & (n_n4983) & (n_n4988) & (n_n4987) & (!x15719x)) + ((n_n4982) & (n_n4983) & (n_n4988) & (n_n4987) & (x15719x)));
	assign x15728x = (((!n_n4953) & (!n_n4956) & (!n_n4965) & (!n_n4955) & (x137x)) + ((!n_n4953) & (!n_n4956) & (!n_n4965) & (n_n4955) & (!x137x)) + ((!n_n4953) & (!n_n4956) & (!n_n4965) & (n_n4955) & (x137x)) + ((!n_n4953) & (!n_n4956) & (n_n4965) & (!n_n4955) & (!x137x)) + ((!n_n4953) & (!n_n4956) & (n_n4965) & (!n_n4955) & (x137x)) + ((!n_n4953) & (!n_n4956) & (n_n4965) & (n_n4955) & (!x137x)) + ((!n_n4953) & (!n_n4956) & (n_n4965) & (n_n4955) & (x137x)) + ((!n_n4953) & (n_n4956) & (!n_n4965) & (!n_n4955) & (!x137x)) + ((!n_n4953) & (n_n4956) & (!n_n4965) & (!n_n4955) & (x137x)) + ((!n_n4953) & (n_n4956) & (!n_n4965) & (n_n4955) & (!x137x)) + ((!n_n4953) & (n_n4956) & (!n_n4965) & (n_n4955) & (x137x)) + ((!n_n4953) & (n_n4956) & (n_n4965) & (!n_n4955) & (!x137x)) + ((!n_n4953) & (n_n4956) & (n_n4965) & (!n_n4955) & (x137x)) + ((!n_n4953) & (n_n4956) & (n_n4965) & (n_n4955) & (!x137x)) + ((!n_n4953) & (n_n4956) & (n_n4965) & (n_n4955) & (x137x)) + ((n_n4953) & (!n_n4956) & (!n_n4965) & (!n_n4955) & (!x137x)) + ((n_n4953) & (!n_n4956) & (!n_n4965) & (!n_n4955) & (x137x)) + ((n_n4953) & (!n_n4956) & (!n_n4965) & (n_n4955) & (!x137x)) + ((n_n4953) & (!n_n4956) & (!n_n4965) & (n_n4955) & (x137x)) + ((n_n4953) & (!n_n4956) & (n_n4965) & (!n_n4955) & (!x137x)) + ((n_n4953) & (!n_n4956) & (n_n4965) & (!n_n4955) & (x137x)) + ((n_n4953) & (!n_n4956) & (n_n4965) & (n_n4955) & (!x137x)) + ((n_n4953) & (!n_n4956) & (n_n4965) & (n_n4955) & (x137x)) + ((n_n4953) & (n_n4956) & (!n_n4965) & (!n_n4955) & (!x137x)) + ((n_n4953) & (n_n4956) & (!n_n4965) & (!n_n4955) & (x137x)) + ((n_n4953) & (n_n4956) & (!n_n4965) & (n_n4955) & (!x137x)) + ((n_n4953) & (n_n4956) & (!n_n4965) & (n_n4955) & (x137x)) + ((n_n4953) & (n_n4956) & (n_n4965) & (!n_n4955) & (!x137x)) + ((n_n4953) & (n_n4956) & (n_n4965) & (!n_n4955) & (x137x)) + ((n_n4953) & (n_n4956) & (n_n4965) & (n_n4955) & (!x137x)) + ((n_n4953) & (n_n4956) & (n_n4965) & (n_n4955) & (x137x)));
	assign x15725x = (((!n_n4958) & (!n_n4947) & (!n_n4966) & (n_n4962)) + ((!n_n4958) & (!n_n4947) & (n_n4966) & (!n_n4962)) + ((!n_n4958) & (!n_n4947) & (n_n4966) & (n_n4962)) + ((!n_n4958) & (n_n4947) & (!n_n4966) & (!n_n4962)) + ((!n_n4958) & (n_n4947) & (!n_n4966) & (n_n4962)) + ((!n_n4958) & (n_n4947) & (n_n4966) & (!n_n4962)) + ((!n_n4958) & (n_n4947) & (n_n4966) & (n_n4962)) + ((n_n4958) & (!n_n4947) & (!n_n4966) & (!n_n4962)) + ((n_n4958) & (!n_n4947) & (!n_n4966) & (n_n4962)) + ((n_n4958) & (!n_n4947) & (n_n4966) & (!n_n4962)) + ((n_n4958) & (!n_n4947) & (n_n4966) & (n_n4962)) + ((n_n4958) & (n_n4947) & (!n_n4966) & (!n_n4962)) + ((n_n4958) & (n_n4947) & (!n_n4966) & (n_n4962)) + ((n_n4958) & (n_n4947) & (n_n4966) & (!n_n4962)) + ((n_n4958) & (n_n4947) & (n_n4966) & (n_n4962)));
	assign n_n2918 = (((!x341x) & (!x317x) & (!n_n2962) & (!x15728x) & (x15725x)) + ((!x341x) & (!x317x) & (!n_n2962) & (x15728x) & (!x15725x)) + ((!x341x) & (!x317x) & (!n_n2962) & (x15728x) & (x15725x)) + ((!x341x) & (!x317x) & (n_n2962) & (!x15728x) & (!x15725x)) + ((!x341x) & (!x317x) & (n_n2962) & (!x15728x) & (x15725x)) + ((!x341x) & (!x317x) & (n_n2962) & (x15728x) & (!x15725x)) + ((!x341x) & (!x317x) & (n_n2962) & (x15728x) & (x15725x)) + ((!x341x) & (x317x) & (!n_n2962) & (!x15728x) & (!x15725x)) + ((!x341x) & (x317x) & (!n_n2962) & (!x15728x) & (x15725x)) + ((!x341x) & (x317x) & (!n_n2962) & (x15728x) & (!x15725x)) + ((!x341x) & (x317x) & (!n_n2962) & (x15728x) & (x15725x)) + ((!x341x) & (x317x) & (n_n2962) & (!x15728x) & (!x15725x)) + ((!x341x) & (x317x) & (n_n2962) & (!x15728x) & (x15725x)) + ((!x341x) & (x317x) & (n_n2962) & (x15728x) & (!x15725x)) + ((!x341x) & (x317x) & (n_n2962) & (x15728x) & (x15725x)) + ((x341x) & (!x317x) & (!n_n2962) & (!x15728x) & (!x15725x)) + ((x341x) & (!x317x) & (!n_n2962) & (!x15728x) & (x15725x)) + ((x341x) & (!x317x) & (!n_n2962) & (x15728x) & (!x15725x)) + ((x341x) & (!x317x) & (!n_n2962) & (x15728x) & (x15725x)) + ((x341x) & (!x317x) & (n_n2962) & (!x15728x) & (!x15725x)) + ((x341x) & (!x317x) & (n_n2962) & (!x15728x) & (x15725x)) + ((x341x) & (!x317x) & (n_n2962) & (x15728x) & (!x15725x)) + ((x341x) & (!x317x) & (n_n2962) & (x15728x) & (x15725x)) + ((x341x) & (x317x) & (!n_n2962) & (!x15728x) & (!x15725x)) + ((x341x) & (x317x) & (!n_n2962) & (!x15728x) & (x15725x)) + ((x341x) & (x317x) & (!n_n2962) & (x15728x) & (!x15725x)) + ((x341x) & (x317x) & (!n_n2962) & (x15728x) & (x15725x)) + ((x341x) & (x317x) & (n_n2962) & (!x15728x) & (!x15725x)) + ((x341x) & (x317x) & (n_n2962) & (!x15728x) & (x15725x)) + ((x341x) & (x317x) & (n_n2962) & (x15728x) & (!x15725x)) + ((x341x) & (x317x) & (n_n2962) & (x15728x) & (x15725x)));
	assign x22204x = (((!n_n5142) & (!n_n5145) & (!n_n5155) & (!n_n5143)));
	assign x13102x = (((!x23x) & (!x583x) & (!x257x) & (!n_n4591) & (n_n4603)) + ((!x23x) & (!x583x) & (!x257x) & (n_n4591) & (!n_n4603)) + ((!x23x) & (!x583x) & (!x257x) & (n_n4591) & (n_n4603)) + ((!x23x) & (!x583x) & (x257x) & (!n_n4591) & (!n_n4603)) + ((!x23x) & (!x583x) & (x257x) & (!n_n4591) & (n_n4603)) + ((!x23x) & (!x583x) & (x257x) & (n_n4591) & (!n_n4603)) + ((!x23x) & (!x583x) & (x257x) & (n_n4591) & (n_n4603)) + ((!x23x) & (x583x) & (!x257x) & (!n_n4591) & (n_n4603)) + ((!x23x) & (x583x) & (!x257x) & (n_n4591) & (!n_n4603)) + ((!x23x) & (x583x) & (!x257x) & (n_n4591) & (n_n4603)) + ((!x23x) & (x583x) & (x257x) & (!n_n4591) & (!n_n4603)) + ((!x23x) & (x583x) & (x257x) & (!n_n4591) & (n_n4603)) + ((!x23x) & (x583x) & (x257x) & (n_n4591) & (!n_n4603)) + ((!x23x) & (x583x) & (x257x) & (n_n4591) & (n_n4603)) + ((x23x) & (!x583x) & (!x257x) & (!n_n4591) & (n_n4603)) + ((x23x) & (!x583x) & (!x257x) & (n_n4591) & (!n_n4603)) + ((x23x) & (!x583x) & (!x257x) & (n_n4591) & (n_n4603)) + ((x23x) & (!x583x) & (x257x) & (!n_n4591) & (!n_n4603)) + ((x23x) & (!x583x) & (x257x) & (!n_n4591) & (n_n4603)) + ((x23x) & (!x583x) & (x257x) & (n_n4591) & (!n_n4603)) + ((x23x) & (!x583x) & (x257x) & (n_n4591) & (n_n4603)) + ((x23x) & (x583x) & (!x257x) & (!n_n4591) & (!n_n4603)) + ((x23x) & (x583x) & (!x257x) & (!n_n4591) & (n_n4603)) + ((x23x) & (x583x) & (!x257x) & (n_n4591) & (!n_n4603)) + ((x23x) & (x583x) & (!x257x) & (n_n4591) & (n_n4603)) + ((x23x) & (x583x) & (x257x) & (!n_n4591) & (!n_n4603)) + ((x23x) & (x583x) & (x257x) & (!n_n4591) & (n_n4603)) + ((x23x) & (x583x) & (x257x) & (n_n4591) & (!n_n4603)) + ((x23x) & (x583x) & (x257x) & (n_n4591) & (n_n4603)));
	assign x14620x = (((!n_n5199) & (!n_n5194) & (!n_n5192) & (x36x)) + ((!n_n5199) & (!n_n5194) & (n_n5192) & (!x36x)) + ((!n_n5199) & (!n_n5194) & (n_n5192) & (x36x)) + ((!n_n5199) & (n_n5194) & (!n_n5192) & (!x36x)) + ((!n_n5199) & (n_n5194) & (!n_n5192) & (x36x)) + ((!n_n5199) & (n_n5194) & (n_n5192) & (!x36x)) + ((!n_n5199) & (n_n5194) & (n_n5192) & (x36x)) + ((n_n5199) & (!n_n5194) & (!n_n5192) & (!x36x)) + ((n_n5199) & (!n_n5194) & (!n_n5192) & (x36x)) + ((n_n5199) & (!n_n5194) & (n_n5192) & (!x36x)) + ((n_n5199) & (!n_n5194) & (n_n5192) & (x36x)) + ((n_n5199) & (n_n5194) & (!n_n5192) & (!x36x)) + ((n_n5199) & (n_n5194) & (!n_n5192) & (x36x)) + ((n_n5199) & (n_n5194) & (n_n5192) & (!x36x)) + ((n_n5199) & (n_n5194) & (n_n5192) & (x36x)));
	assign n_n3670 = (((!n_n5200) & (!n_n5193) & (!x452x) & (x14620x)) + ((!n_n5200) & (!n_n5193) & (x452x) & (!x14620x)) + ((!n_n5200) & (!n_n5193) & (x452x) & (x14620x)) + ((!n_n5200) & (n_n5193) & (!x452x) & (!x14620x)) + ((!n_n5200) & (n_n5193) & (!x452x) & (x14620x)) + ((!n_n5200) & (n_n5193) & (x452x) & (!x14620x)) + ((!n_n5200) & (n_n5193) & (x452x) & (x14620x)) + ((n_n5200) & (!n_n5193) & (!x452x) & (!x14620x)) + ((n_n5200) & (!n_n5193) & (!x452x) & (x14620x)) + ((n_n5200) & (!n_n5193) & (x452x) & (!x14620x)) + ((n_n5200) & (!n_n5193) & (x452x) & (x14620x)) + ((n_n5200) & (n_n5193) & (!x452x) & (!x14620x)) + ((n_n5200) & (n_n5193) & (!x452x) & (x14620x)) + ((n_n5200) & (n_n5193) & (x452x) & (!x14620x)) + ((n_n5200) & (n_n5193) & (x452x) & (x14620x)));
	assign x15531x = (((!i_9_) & (n_n536) & (!n_n532) & (n_n534) & (n_n464)) + ((!i_9_) & (n_n536) & (n_n532) & (!n_n534) & (n_n464)) + ((!i_9_) & (n_n536) & (n_n532) & (n_n534) & (n_n464)) + ((i_9_) & (n_n536) & (n_n532) & (!n_n534) & (n_n464)) + ((i_9_) & (n_n536) & (n_n532) & (n_n534) & (n_n464)));
	assign x22200x = (((!n_n4434) & (!n_n4432) & (!n_n4430) & (!n_n4429)));
	assign x22084x = (((!x19x) & (!n_n5310) & (!x502x) & (!n_n5300) & (!n_n5299)) + ((!x19x) & (!n_n5310) & (x502x) & (!n_n5300) & (!n_n5299)) + ((x19x) & (!n_n5310) & (!x502x) & (!n_n5300) & (!n_n5299)));
	assign n_n2937 = (((!x592x) & (!x23x) & (!n_n5313) & (!n_n3019) & (!x22084x)) + ((!x592x) & (!x23x) & (!n_n5313) & (n_n3019) & (!x22084x)) + ((!x592x) & (!x23x) & (!n_n5313) & (n_n3019) & (x22084x)) + ((!x592x) & (!x23x) & (n_n5313) & (!n_n3019) & (!x22084x)) + ((!x592x) & (!x23x) & (n_n5313) & (!n_n3019) & (x22084x)) + ((!x592x) & (!x23x) & (n_n5313) & (n_n3019) & (!x22084x)) + ((!x592x) & (!x23x) & (n_n5313) & (n_n3019) & (x22084x)) + ((!x592x) & (x23x) & (!n_n5313) & (!n_n3019) & (!x22084x)) + ((!x592x) & (x23x) & (!n_n5313) & (n_n3019) & (!x22084x)) + ((!x592x) & (x23x) & (!n_n5313) & (n_n3019) & (x22084x)) + ((!x592x) & (x23x) & (n_n5313) & (!n_n3019) & (!x22084x)) + ((!x592x) & (x23x) & (n_n5313) & (!n_n3019) & (x22084x)) + ((!x592x) & (x23x) & (n_n5313) & (n_n3019) & (!x22084x)) + ((!x592x) & (x23x) & (n_n5313) & (n_n3019) & (x22084x)) + ((x592x) & (!x23x) & (!n_n5313) & (!n_n3019) & (!x22084x)) + ((x592x) & (!x23x) & (!n_n5313) & (n_n3019) & (!x22084x)) + ((x592x) & (!x23x) & (!n_n5313) & (n_n3019) & (x22084x)) + ((x592x) & (!x23x) & (n_n5313) & (!n_n3019) & (!x22084x)) + ((x592x) & (!x23x) & (n_n5313) & (!n_n3019) & (x22084x)) + ((x592x) & (!x23x) & (n_n5313) & (n_n3019) & (!x22084x)) + ((x592x) & (!x23x) & (n_n5313) & (n_n3019) & (x22084x)) + ((x592x) & (x23x) & (!n_n5313) & (!n_n3019) & (!x22084x)) + ((x592x) & (x23x) & (!n_n5313) & (!n_n3019) & (x22084x)) + ((x592x) & (x23x) & (!n_n5313) & (n_n3019) & (!x22084x)) + ((x592x) & (x23x) & (!n_n5313) & (n_n3019) & (x22084x)) + ((x592x) & (x23x) & (n_n5313) & (!n_n3019) & (!x22084x)) + ((x592x) & (x23x) & (n_n5313) & (!n_n3019) & (x22084x)) + ((x592x) & (x23x) & (n_n5313) & (n_n3019) & (!x22084x)) + ((x592x) & (x23x) & (n_n5313) & (n_n3019) & (x22084x)));
	assign x15433x = (((!i_9_) & (n_n455) & (n_n532) & (!n_n534) & (n_n491)) + ((!i_9_) & (n_n455) & (n_n532) & (n_n534) & (n_n491)) + ((i_9_) & (n_n455) & (!n_n532) & (n_n534) & (n_n491)) + ((i_9_) & (n_n455) & (n_n532) & (n_n534) & (n_n491)));
	assign x15734x = (((!n_n4934) & (!n_n4946) & (!n_n4937) & (!n_n4935) & (n_n4944)) + ((!n_n4934) & (!n_n4946) & (!n_n4937) & (n_n4935) & (!n_n4944)) + ((!n_n4934) & (!n_n4946) & (!n_n4937) & (n_n4935) & (n_n4944)) + ((!n_n4934) & (!n_n4946) & (n_n4937) & (!n_n4935) & (!n_n4944)) + ((!n_n4934) & (!n_n4946) & (n_n4937) & (!n_n4935) & (n_n4944)) + ((!n_n4934) & (!n_n4946) & (n_n4937) & (n_n4935) & (!n_n4944)) + ((!n_n4934) & (!n_n4946) & (n_n4937) & (n_n4935) & (n_n4944)) + ((!n_n4934) & (n_n4946) & (!n_n4937) & (!n_n4935) & (!n_n4944)) + ((!n_n4934) & (n_n4946) & (!n_n4937) & (!n_n4935) & (n_n4944)) + ((!n_n4934) & (n_n4946) & (!n_n4937) & (n_n4935) & (!n_n4944)) + ((!n_n4934) & (n_n4946) & (!n_n4937) & (n_n4935) & (n_n4944)) + ((!n_n4934) & (n_n4946) & (n_n4937) & (!n_n4935) & (!n_n4944)) + ((!n_n4934) & (n_n4946) & (n_n4937) & (!n_n4935) & (n_n4944)) + ((!n_n4934) & (n_n4946) & (n_n4937) & (n_n4935) & (!n_n4944)) + ((!n_n4934) & (n_n4946) & (n_n4937) & (n_n4935) & (n_n4944)) + ((n_n4934) & (!n_n4946) & (!n_n4937) & (!n_n4935) & (!n_n4944)) + ((n_n4934) & (!n_n4946) & (!n_n4937) & (!n_n4935) & (n_n4944)) + ((n_n4934) & (!n_n4946) & (!n_n4937) & (n_n4935) & (!n_n4944)) + ((n_n4934) & (!n_n4946) & (!n_n4937) & (n_n4935) & (n_n4944)) + ((n_n4934) & (!n_n4946) & (n_n4937) & (!n_n4935) & (!n_n4944)) + ((n_n4934) & (!n_n4946) & (n_n4937) & (!n_n4935) & (n_n4944)) + ((n_n4934) & (!n_n4946) & (n_n4937) & (n_n4935) & (!n_n4944)) + ((n_n4934) & (!n_n4946) & (n_n4937) & (n_n4935) & (n_n4944)) + ((n_n4934) & (n_n4946) & (!n_n4937) & (!n_n4935) & (!n_n4944)) + ((n_n4934) & (n_n4946) & (!n_n4937) & (!n_n4935) & (n_n4944)) + ((n_n4934) & (n_n4946) & (!n_n4937) & (n_n4935) & (!n_n4944)) + ((n_n4934) & (n_n4946) & (!n_n4937) & (n_n4935) & (n_n4944)) + ((n_n4934) & (n_n4946) & (n_n4937) & (!n_n4935) & (!n_n4944)) + ((n_n4934) & (n_n4946) & (n_n4937) & (!n_n4935) & (n_n4944)) + ((n_n4934) & (n_n4946) & (n_n4937) & (n_n4935) & (!n_n4944)) + ((n_n4934) & (n_n4946) & (n_n4937) & (n_n4935) & (n_n4944)));
	assign n_n2965 = (((!x15x) & (!x531x) & (!n_n4942) & (!x411x) & (x15734x)) + ((!x15x) & (!x531x) & (!n_n4942) & (x411x) & (!x15734x)) + ((!x15x) & (!x531x) & (!n_n4942) & (x411x) & (x15734x)) + ((!x15x) & (!x531x) & (n_n4942) & (!x411x) & (!x15734x)) + ((!x15x) & (!x531x) & (n_n4942) & (!x411x) & (x15734x)) + ((!x15x) & (!x531x) & (n_n4942) & (x411x) & (!x15734x)) + ((!x15x) & (!x531x) & (n_n4942) & (x411x) & (x15734x)) + ((!x15x) & (x531x) & (!n_n4942) & (!x411x) & (x15734x)) + ((!x15x) & (x531x) & (!n_n4942) & (x411x) & (!x15734x)) + ((!x15x) & (x531x) & (!n_n4942) & (x411x) & (x15734x)) + ((!x15x) & (x531x) & (n_n4942) & (!x411x) & (!x15734x)) + ((!x15x) & (x531x) & (n_n4942) & (!x411x) & (x15734x)) + ((!x15x) & (x531x) & (n_n4942) & (x411x) & (!x15734x)) + ((!x15x) & (x531x) & (n_n4942) & (x411x) & (x15734x)) + ((x15x) & (!x531x) & (!n_n4942) & (!x411x) & (x15734x)) + ((x15x) & (!x531x) & (!n_n4942) & (x411x) & (!x15734x)) + ((x15x) & (!x531x) & (!n_n4942) & (x411x) & (x15734x)) + ((x15x) & (!x531x) & (n_n4942) & (!x411x) & (!x15734x)) + ((x15x) & (!x531x) & (n_n4942) & (!x411x) & (x15734x)) + ((x15x) & (!x531x) & (n_n4942) & (x411x) & (!x15734x)) + ((x15x) & (!x531x) & (n_n4942) & (x411x) & (x15734x)) + ((x15x) & (x531x) & (!n_n4942) & (!x411x) & (!x15734x)) + ((x15x) & (x531x) & (!n_n4942) & (!x411x) & (x15734x)) + ((x15x) & (x531x) & (!n_n4942) & (x411x) & (!x15734x)) + ((x15x) & (x531x) & (!n_n4942) & (x411x) & (x15734x)) + ((x15x) & (x531x) & (n_n4942) & (!x411x) & (!x15734x)) + ((x15x) & (x531x) & (n_n4942) & (!x411x) & (x15734x)) + ((x15x) & (x531x) & (n_n4942) & (x411x) & (!x15734x)) + ((x15x) & (x531x) & (n_n4942) & (x411x) & (x15734x)));
	assign x14561x = (((!n_n5321) & (!n_n5319) & (!n_n5322) & (!n_n5324) & (n_n5328)) + ((!n_n5321) & (!n_n5319) & (!n_n5322) & (n_n5324) & (!n_n5328)) + ((!n_n5321) & (!n_n5319) & (!n_n5322) & (n_n5324) & (n_n5328)) + ((!n_n5321) & (!n_n5319) & (n_n5322) & (!n_n5324) & (!n_n5328)) + ((!n_n5321) & (!n_n5319) & (n_n5322) & (!n_n5324) & (n_n5328)) + ((!n_n5321) & (!n_n5319) & (n_n5322) & (n_n5324) & (!n_n5328)) + ((!n_n5321) & (!n_n5319) & (n_n5322) & (n_n5324) & (n_n5328)) + ((!n_n5321) & (n_n5319) & (!n_n5322) & (!n_n5324) & (!n_n5328)) + ((!n_n5321) & (n_n5319) & (!n_n5322) & (!n_n5324) & (n_n5328)) + ((!n_n5321) & (n_n5319) & (!n_n5322) & (n_n5324) & (!n_n5328)) + ((!n_n5321) & (n_n5319) & (!n_n5322) & (n_n5324) & (n_n5328)) + ((!n_n5321) & (n_n5319) & (n_n5322) & (!n_n5324) & (!n_n5328)) + ((!n_n5321) & (n_n5319) & (n_n5322) & (!n_n5324) & (n_n5328)) + ((!n_n5321) & (n_n5319) & (n_n5322) & (n_n5324) & (!n_n5328)) + ((!n_n5321) & (n_n5319) & (n_n5322) & (n_n5324) & (n_n5328)) + ((n_n5321) & (!n_n5319) & (!n_n5322) & (!n_n5324) & (!n_n5328)) + ((n_n5321) & (!n_n5319) & (!n_n5322) & (!n_n5324) & (n_n5328)) + ((n_n5321) & (!n_n5319) & (!n_n5322) & (n_n5324) & (!n_n5328)) + ((n_n5321) & (!n_n5319) & (!n_n5322) & (n_n5324) & (n_n5328)) + ((n_n5321) & (!n_n5319) & (n_n5322) & (!n_n5324) & (!n_n5328)) + ((n_n5321) & (!n_n5319) & (n_n5322) & (!n_n5324) & (n_n5328)) + ((n_n5321) & (!n_n5319) & (n_n5322) & (n_n5324) & (!n_n5328)) + ((n_n5321) & (!n_n5319) & (n_n5322) & (n_n5324) & (n_n5328)) + ((n_n5321) & (n_n5319) & (!n_n5322) & (!n_n5324) & (!n_n5328)) + ((n_n5321) & (n_n5319) & (!n_n5322) & (!n_n5324) & (n_n5328)) + ((n_n5321) & (n_n5319) & (!n_n5322) & (n_n5324) & (!n_n5328)) + ((n_n5321) & (n_n5319) & (!n_n5322) & (n_n5324) & (n_n5328)) + ((n_n5321) & (n_n5319) & (n_n5322) & (!n_n5324) & (!n_n5328)) + ((n_n5321) & (n_n5319) & (n_n5322) & (!n_n5324) & (n_n5328)) + ((n_n5321) & (n_n5319) & (n_n5322) & (n_n5324) & (!n_n5328)) + ((n_n5321) & (n_n5319) & (n_n5322) & (n_n5324) & (n_n5328)));
	assign x15536x = (((!i_9_) & (!n_n536) & (!n_n524) & (!n_n473) & (x215x)) + ((!i_9_) & (!n_n536) & (!n_n524) & (n_n473) & (x215x)) + ((!i_9_) & (!n_n536) & (n_n524) & (!n_n473) & (x215x)) + ((!i_9_) & (!n_n536) & (n_n524) & (n_n473) & (x215x)) + ((!i_9_) & (n_n536) & (!n_n524) & (!n_n473) & (x215x)) + ((!i_9_) & (n_n536) & (!n_n524) & (n_n473) & (x215x)) + ((!i_9_) & (n_n536) & (n_n524) & (!n_n473) & (x215x)) + ((!i_9_) & (n_n536) & (n_n524) & (n_n473) & (!x215x)) + ((!i_9_) & (n_n536) & (n_n524) & (n_n473) & (x215x)) + ((i_9_) & (!n_n536) & (!n_n524) & (!n_n473) & (x215x)) + ((i_9_) & (!n_n536) & (!n_n524) & (n_n473) & (x215x)) + ((i_9_) & (!n_n536) & (n_n524) & (!n_n473) & (x215x)) + ((i_9_) & (!n_n536) & (n_n524) & (n_n473) & (x215x)) + ((i_9_) & (n_n536) & (!n_n524) & (!n_n473) & (x215x)) + ((i_9_) & (n_n536) & (!n_n524) & (n_n473) & (x215x)) + ((i_9_) & (n_n536) & (n_n524) & (!n_n473) & (x215x)) + ((i_9_) & (n_n536) & (n_n524) & (n_n473) & (!x215x)) + ((i_9_) & (n_n536) & (n_n524) & (n_n473) & (x215x)));
	assign x15668x = (((!x592x) & (!x11x) & (!n_n5289) & (!x208x) & (n_n5285)) + ((!x592x) & (!x11x) & (!n_n5289) & (x208x) & (!n_n5285)) + ((!x592x) & (!x11x) & (!n_n5289) & (x208x) & (n_n5285)) + ((!x592x) & (!x11x) & (n_n5289) & (!x208x) & (!n_n5285)) + ((!x592x) & (!x11x) & (n_n5289) & (!x208x) & (n_n5285)) + ((!x592x) & (!x11x) & (n_n5289) & (x208x) & (!n_n5285)) + ((!x592x) & (!x11x) & (n_n5289) & (x208x) & (n_n5285)) + ((!x592x) & (x11x) & (!n_n5289) & (!x208x) & (n_n5285)) + ((!x592x) & (x11x) & (!n_n5289) & (x208x) & (!n_n5285)) + ((!x592x) & (x11x) & (!n_n5289) & (x208x) & (n_n5285)) + ((!x592x) & (x11x) & (n_n5289) & (!x208x) & (!n_n5285)) + ((!x592x) & (x11x) & (n_n5289) & (!x208x) & (n_n5285)) + ((!x592x) & (x11x) & (n_n5289) & (x208x) & (!n_n5285)) + ((!x592x) & (x11x) & (n_n5289) & (x208x) & (n_n5285)) + ((x592x) & (!x11x) & (!n_n5289) & (!x208x) & (n_n5285)) + ((x592x) & (!x11x) & (!n_n5289) & (x208x) & (!n_n5285)) + ((x592x) & (!x11x) & (!n_n5289) & (x208x) & (n_n5285)) + ((x592x) & (!x11x) & (n_n5289) & (!x208x) & (!n_n5285)) + ((x592x) & (!x11x) & (n_n5289) & (!x208x) & (n_n5285)) + ((x592x) & (!x11x) & (n_n5289) & (x208x) & (!n_n5285)) + ((x592x) & (!x11x) & (n_n5289) & (x208x) & (n_n5285)) + ((x592x) & (x11x) & (!n_n5289) & (!x208x) & (!n_n5285)) + ((x592x) & (x11x) & (!n_n5289) & (!x208x) & (n_n5285)) + ((x592x) & (x11x) & (!n_n5289) & (x208x) & (!n_n5285)) + ((x592x) & (x11x) & (!n_n5289) & (x208x) & (n_n5285)) + ((x592x) & (x11x) & (n_n5289) & (!x208x) & (!n_n5285)) + ((x592x) & (x11x) & (n_n5289) & (!x208x) & (n_n5285)) + ((x592x) & (x11x) & (n_n5289) & (x208x) & (!n_n5285)) + ((x592x) & (x11x) & (n_n5289) & (x208x) & (n_n5285)));
	assign x22080x = (((!n_n4547) & (!n_n4544) & (!n_n4538) & (!n_n4546)));
	assign x15453x = (((!x201x) & (!n_n4549) & (!n_n4545) & (!n_n4550) & (!x22080x)) + ((!x201x) & (!n_n4549) & (!n_n4545) & (n_n4550) & (!x22080x)) + ((!x201x) & (!n_n4549) & (!n_n4545) & (n_n4550) & (x22080x)) + ((!x201x) & (!n_n4549) & (n_n4545) & (!n_n4550) & (!x22080x)) + ((!x201x) & (!n_n4549) & (n_n4545) & (!n_n4550) & (x22080x)) + ((!x201x) & (!n_n4549) & (n_n4545) & (n_n4550) & (!x22080x)) + ((!x201x) & (!n_n4549) & (n_n4545) & (n_n4550) & (x22080x)) + ((!x201x) & (n_n4549) & (!n_n4545) & (!n_n4550) & (!x22080x)) + ((!x201x) & (n_n4549) & (!n_n4545) & (!n_n4550) & (x22080x)) + ((!x201x) & (n_n4549) & (!n_n4545) & (n_n4550) & (!x22080x)) + ((!x201x) & (n_n4549) & (!n_n4545) & (n_n4550) & (x22080x)) + ((!x201x) & (n_n4549) & (n_n4545) & (!n_n4550) & (!x22080x)) + ((!x201x) & (n_n4549) & (n_n4545) & (!n_n4550) & (x22080x)) + ((!x201x) & (n_n4549) & (n_n4545) & (n_n4550) & (!x22080x)) + ((!x201x) & (n_n4549) & (n_n4545) & (n_n4550) & (x22080x)) + ((x201x) & (!n_n4549) & (!n_n4545) & (!n_n4550) & (!x22080x)) + ((x201x) & (!n_n4549) & (!n_n4545) & (!n_n4550) & (x22080x)) + ((x201x) & (!n_n4549) & (!n_n4545) & (n_n4550) & (!x22080x)) + ((x201x) & (!n_n4549) & (!n_n4545) & (n_n4550) & (x22080x)) + ((x201x) & (!n_n4549) & (n_n4545) & (!n_n4550) & (!x22080x)) + ((x201x) & (!n_n4549) & (n_n4545) & (!n_n4550) & (x22080x)) + ((x201x) & (!n_n4549) & (n_n4545) & (n_n4550) & (!x22080x)) + ((x201x) & (!n_n4549) & (n_n4545) & (n_n4550) & (x22080x)) + ((x201x) & (n_n4549) & (!n_n4545) & (!n_n4550) & (!x22080x)) + ((x201x) & (n_n4549) & (!n_n4545) & (!n_n4550) & (x22080x)) + ((x201x) & (n_n4549) & (!n_n4545) & (n_n4550) & (!x22080x)) + ((x201x) & (n_n4549) & (!n_n4545) & (n_n4550) & (x22080x)) + ((x201x) & (n_n4549) & (n_n4545) & (!n_n4550) & (!x22080x)) + ((x201x) & (n_n4549) & (n_n4545) & (!n_n4550) & (x22080x)) + ((x201x) & (n_n4549) & (n_n4545) & (n_n4550) & (!x22080x)) + ((x201x) & (n_n4549) & (n_n4545) & (n_n4550) & (x22080x)));
	assign x15876x = (((!i_5_) & (i_3_) & (!i_4_) & (x15x) & (n_n130)) + ((i_5_) & (!i_3_) & (i_4_) & (x15x) & (n_n130)));
	assign x15879x = (((!n_n5179) & (!n_n5178) & (!n_n5138) & (x15876x)) + ((!n_n5179) & (!n_n5178) & (n_n5138) & (!x15876x)) + ((!n_n5179) & (!n_n5178) & (n_n5138) & (x15876x)) + ((!n_n5179) & (n_n5178) & (!n_n5138) & (!x15876x)) + ((!n_n5179) & (n_n5178) & (!n_n5138) & (x15876x)) + ((!n_n5179) & (n_n5178) & (n_n5138) & (!x15876x)) + ((!n_n5179) & (n_n5178) & (n_n5138) & (x15876x)) + ((n_n5179) & (!n_n5178) & (!n_n5138) & (!x15876x)) + ((n_n5179) & (!n_n5178) & (!n_n5138) & (x15876x)) + ((n_n5179) & (!n_n5178) & (n_n5138) & (!x15876x)) + ((n_n5179) & (!n_n5178) & (n_n5138) & (x15876x)) + ((n_n5179) & (n_n5178) & (!n_n5138) & (!x15876x)) + ((n_n5179) & (n_n5178) & (!n_n5138) & (x15876x)) + ((n_n5179) & (n_n5178) & (n_n5138) & (!x15876x)) + ((n_n5179) & (n_n5178) & (n_n5138) & (x15876x)));
	assign x11682x = (((!n_n4834) & (!n_n4832) & (!n_n4850) & (!n_n4844) & (n_n4833)) + ((!n_n4834) & (!n_n4832) & (!n_n4850) & (n_n4844) & (!n_n4833)) + ((!n_n4834) & (!n_n4832) & (!n_n4850) & (n_n4844) & (n_n4833)) + ((!n_n4834) & (!n_n4832) & (n_n4850) & (!n_n4844) & (!n_n4833)) + ((!n_n4834) & (!n_n4832) & (n_n4850) & (!n_n4844) & (n_n4833)) + ((!n_n4834) & (!n_n4832) & (n_n4850) & (n_n4844) & (!n_n4833)) + ((!n_n4834) & (!n_n4832) & (n_n4850) & (n_n4844) & (n_n4833)) + ((!n_n4834) & (n_n4832) & (!n_n4850) & (!n_n4844) & (!n_n4833)) + ((!n_n4834) & (n_n4832) & (!n_n4850) & (!n_n4844) & (n_n4833)) + ((!n_n4834) & (n_n4832) & (!n_n4850) & (n_n4844) & (!n_n4833)) + ((!n_n4834) & (n_n4832) & (!n_n4850) & (n_n4844) & (n_n4833)) + ((!n_n4834) & (n_n4832) & (n_n4850) & (!n_n4844) & (!n_n4833)) + ((!n_n4834) & (n_n4832) & (n_n4850) & (!n_n4844) & (n_n4833)) + ((!n_n4834) & (n_n4832) & (n_n4850) & (n_n4844) & (!n_n4833)) + ((!n_n4834) & (n_n4832) & (n_n4850) & (n_n4844) & (n_n4833)) + ((n_n4834) & (!n_n4832) & (!n_n4850) & (!n_n4844) & (!n_n4833)) + ((n_n4834) & (!n_n4832) & (!n_n4850) & (!n_n4844) & (n_n4833)) + ((n_n4834) & (!n_n4832) & (!n_n4850) & (n_n4844) & (!n_n4833)) + ((n_n4834) & (!n_n4832) & (!n_n4850) & (n_n4844) & (n_n4833)) + ((n_n4834) & (!n_n4832) & (n_n4850) & (!n_n4844) & (!n_n4833)) + ((n_n4834) & (!n_n4832) & (n_n4850) & (!n_n4844) & (n_n4833)) + ((n_n4834) & (!n_n4832) & (n_n4850) & (n_n4844) & (!n_n4833)) + ((n_n4834) & (!n_n4832) & (n_n4850) & (n_n4844) & (n_n4833)) + ((n_n4834) & (n_n4832) & (!n_n4850) & (!n_n4844) & (!n_n4833)) + ((n_n4834) & (n_n4832) & (!n_n4850) & (!n_n4844) & (n_n4833)) + ((n_n4834) & (n_n4832) & (!n_n4850) & (n_n4844) & (!n_n4833)) + ((n_n4834) & (n_n4832) & (!n_n4850) & (n_n4844) & (n_n4833)) + ((n_n4834) & (n_n4832) & (n_n4850) & (!n_n4844) & (!n_n4833)) + ((n_n4834) & (n_n4832) & (n_n4850) & (!n_n4844) & (n_n4833)) + ((n_n4834) & (n_n4832) & (n_n4850) & (n_n4844) & (!n_n4833)) + ((n_n4834) & (n_n4832) & (n_n4850) & (n_n4844) & (n_n4833)));
	assign x12763x = (((!n_n4784) & (!n_n4788) & (!n_n4780) & (!n_n4783) & (n_n4778)) + ((!n_n4784) & (!n_n4788) & (!n_n4780) & (n_n4783) & (!n_n4778)) + ((!n_n4784) & (!n_n4788) & (!n_n4780) & (n_n4783) & (n_n4778)) + ((!n_n4784) & (!n_n4788) & (n_n4780) & (!n_n4783) & (!n_n4778)) + ((!n_n4784) & (!n_n4788) & (n_n4780) & (!n_n4783) & (n_n4778)) + ((!n_n4784) & (!n_n4788) & (n_n4780) & (n_n4783) & (!n_n4778)) + ((!n_n4784) & (!n_n4788) & (n_n4780) & (n_n4783) & (n_n4778)) + ((!n_n4784) & (n_n4788) & (!n_n4780) & (!n_n4783) & (!n_n4778)) + ((!n_n4784) & (n_n4788) & (!n_n4780) & (!n_n4783) & (n_n4778)) + ((!n_n4784) & (n_n4788) & (!n_n4780) & (n_n4783) & (!n_n4778)) + ((!n_n4784) & (n_n4788) & (!n_n4780) & (n_n4783) & (n_n4778)) + ((!n_n4784) & (n_n4788) & (n_n4780) & (!n_n4783) & (!n_n4778)) + ((!n_n4784) & (n_n4788) & (n_n4780) & (!n_n4783) & (n_n4778)) + ((!n_n4784) & (n_n4788) & (n_n4780) & (n_n4783) & (!n_n4778)) + ((!n_n4784) & (n_n4788) & (n_n4780) & (n_n4783) & (n_n4778)) + ((n_n4784) & (!n_n4788) & (!n_n4780) & (!n_n4783) & (!n_n4778)) + ((n_n4784) & (!n_n4788) & (!n_n4780) & (!n_n4783) & (n_n4778)) + ((n_n4784) & (!n_n4788) & (!n_n4780) & (n_n4783) & (!n_n4778)) + ((n_n4784) & (!n_n4788) & (!n_n4780) & (n_n4783) & (n_n4778)) + ((n_n4784) & (!n_n4788) & (n_n4780) & (!n_n4783) & (!n_n4778)) + ((n_n4784) & (!n_n4788) & (n_n4780) & (!n_n4783) & (n_n4778)) + ((n_n4784) & (!n_n4788) & (n_n4780) & (n_n4783) & (!n_n4778)) + ((n_n4784) & (!n_n4788) & (n_n4780) & (n_n4783) & (n_n4778)) + ((n_n4784) & (n_n4788) & (!n_n4780) & (!n_n4783) & (!n_n4778)) + ((n_n4784) & (n_n4788) & (!n_n4780) & (!n_n4783) & (n_n4778)) + ((n_n4784) & (n_n4788) & (!n_n4780) & (n_n4783) & (!n_n4778)) + ((n_n4784) & (n_n4788) & (!n_n4780) & (n_n4783) & (n_n4778)) + ((n_n4784) & (n_n4788) & (n_n4780) & (!n_n4783) & (!n_n4778)) + ((n_n4784) & (n_n4788) & (n_n4780) & (!n_n4783) & (n_n4778)) + ((n_n4784) & (n_n4788) & (n_n4780) & (n_n4783) & (!n_n4778)) + ((n_n4784) & (n_n4788) & (n_n4780) & (n_n4783) & (n_n4778)));
	assign x14687x = (((!i_9_) & (n_n524) & (!n_n528) & (n_n509) & (n_n260)) + ((!i_9_) & (n_n524) & (n_n528) & (n_n509) & (n_n260)) + ((i_9_) & (!n_n524) & (n_n528) & (n_n509) & (n_n260)) + ((i_9_) & (n_n524) & (n_n528) & (n_n509) & (n_n260)));
	assign x22111x = (((!n_n4843) & (!n_n4845) & (!n_n4848) & (!n_n4842)));
	assign x14548x = (((!i_9_) & (!n_n528) & (!n_n500) & (!n_n65) & (x77x)) + ((!i_9_) & (!n_n528) & (!n_n500) & (n_n65) & (x77x)) + ((!i_9_) & (!n_n528) & (n_n500) & (!n_n65) & (x77x)) + ((!i_9_) & (!n_n528) & (n_n500) & (n_n65) & (x77x)) + ((!i_9_) & (n_n528) & (!n_n500) & (!n_n65) & (x77x)) + ((!i_9_) & (n_n528) & (!n_n500) & (n_n65) & (x77x)) + ((!i_9_) & (n_n528) & (n_n500) & (!n_n65) & (x77x)) + ((!i_9_) & (n_n528) & (n_n500) & (n_n65) & (!x77x)) + ((!i_9_) & (n_n528) & (n_n500) & (n_n65) & (x77x)) + ((i_9_) & (!n_n528) & (!n_n500) & (!n_n65) & (x77x)) + ((i_9_) & (!n_n528) & (!n_n500) & (n_n65) & (x77x)) + ((i_9_) & (!n_n528) & (n_n500) & (!n_n65) & (x77x)) + ((i_9_) & (!n_n528) & (n_n500) & (n_n65) & (x77x)) + ((i_9_) & (n_n528) & (!n_n500) & (!n_n65) & (x77x)) + ((i_9_) & (n_n528) & (!n_n500) & (n_n65) & (x77x)) + ((i_9_) & (n_n528) & (n_n500) & (!n_n65) & (x77x)) + ((i_9_) & (n_n528) & (n_n500) & (n_n65) & (x77x)));
	assign x14506x = (((!i_9_) & (!n_n536) & (!n_n473) & (!n_n532) & (x14504x)) + ((!i_9_) & (!n_n536) & (!n_n473) & (n_n532) & (x14504x)) + ((!i_9_) & (!n_n536) & (n_n473) & (!n_n532) & (x14504x)) + ((!i_9_) & (!n_n536) & (n_n473) & (n_n532) & (x14504x)) + ((!i_9_) & (n_n536) & (!n_n473) & (!n_n532) & (x14504x)) + ((!i_9_) & (n_n536) & (!n_n473) & (n_n532) & (x14504x)) + ((!i_9_) & (n_n536) & (n_n473) & (!n_n532) & (x14504x)) + ((!i_9_) & (n_n536) & (n_n473) & (n_n532) & (!x14504x)) + ((!i_9_) & (n_n536) & (n_n473) & (n_n532) & (x14504x)) + ((i_9_) & (!n_n536) & (!n_n473) & (!n_n532) & (x14504x)) + ((i_9_) & (!n_n536) & (!n_n473) & (n_n532) & (x14504x)) + ((i_9_) & (!n_n536) & (n_n473) & (!n_n532) & (x14504x)) + ((i_9_) & (!n_n536) & (n_n473) & (n_n532) & (x14504x)) + ((i_9_) & (n_n536) & (!n_n473) & (!n_n532) & (x14504x)) + ((i_9_) & (n_n536) & (!n_n473) & (n_n532) & (x14504x)) + ((i_9_) & (n_n536) & (n_n473) & (!n_n532) & (x14504x)) + ((i_9_) & (n_n536) & (n_n473) & (n_n532) & (!x14504x)) + ((i_9_) & (n_n536) & (n_n473) & (n_n532) & (x14504x)));
	assign x15542x = (((!n_n4401) & (!n_n4404) & (!n_n4406) & (!n_n4402) & (n_n4408)) + ((!n_n4401) & (!n_n4404) & (!n_n4406) & (n_n4402) & (!n_n4408)) + ((!n_n4401) & (!n_n4404) & (!n_n4406) & (n_n4402) & (n_n4408)) + ((!n_n4401) & (!n_n4404) & (n_n4406) & (!n_n4402) & (!n_n4408)) + ((!n_n4401) & (!n_n4404) & (n_n4406) & (!n_n4402) & (n_n4408)) + ((!n_n4401) & (!n_n4404) & (n_n4406) & (n_n4402) & (!n_n4408)) + ((!n_n4401) & (!n_n4404) & (n_n4406) & (n_n4402) & (n_n4408)) + ((!n_n4401) & (n_n4404) & (!n_n4406) & (!n_n4402) & (!n_n4408)) + ((!n_n4401) & (n_n4404) & (!n_n4406) & (!n_n4402) & (n_n4408)) + ((!n_n4401) & (n_n4404) & (!n_n4406) & (n_n4402) & (!n_n4408)) + ((!n_n4401) & (n_n4404) & (!n_n4406) & (n_n4402) & (n_n4408)) + ((!n_n4401) & (n_n4404) & (n_n4406) & (!n_n4402) & (!n_n4408)) + ((!n_n4401) & (n_n4404) & (n_n4406) & (!n_n4402) & (n_n4408)) + ((!n_n4401) & (n_n4404) & (n_n4406) & (n_n4402) & (!n_n4408)) + ((!n_n4401) & (n_n4404) & (n_n4406) & (n_n4402) & (n_n4408)) + ((n_n4401) & (!n_n4404) & (!n_n4406) & (!n_n4402) & (!n_n4408)) + ((n_n4401) & (!n_n4404) & (!n_n4406) & (!n_n4402) & (n_n4408)) + ((n_n4401) & (!n_n4404) & (!n_n4406) & (n_n4402) & (!n_n4408)) + ((n_n4401) & (!n_n4404) & (!n_n4406) & (n_n4402) & (n_n4408)) + ((n_n4401) & (!n_n4404) & (n_n4406) & (!n_n4402) & (!n_n4408)) + ((n_n4401) & (!n_n4404) & (n_n4406) & (!n_n4402) & (n_n4408)) + ((n_n4401) & (!n_n4404) & (n_n4406) & (n_n4402) & (!n_n4408)) + ((n_n4401) & (!n_n4404) & (n_n4406) & (n_n4402) & (n_n4408)) + ((n_n4401) & (n_n4404) & (!n_n4406) & (!n_n4402) & (!n_n4408)) + ((n_n4401) & (n_n4404) & (!n_n4406) & (!n_n4402) & (n_n4408)) + ((n_n4401) & (n_n4404) & (!n_n4406) & (n_n4402) & (!n_n4408)) + ((n_n4401) & (n_n4404) & (!n_n4406) & (n_n4402) & (n_n4408)) + ((n_n4401) & (n_n4404) & (n_n4406) & (!n_n4402) & (!n_n4408)) + ((n_n4401) & (n_n4404) & (n_n4406) & (!n_n4402) & (n_n4408)) + ((n_n4401) & (n_n4404) & (n_n4406) & (n_n4402) & (!n_n4408)) + ((n_n4401) & (n_n4404) & (n_n4406) & (n_n4402) & (n_n4408)));
	assign x22223x = (((!n_n4533) & (!n_n4531) & (!n_n4535) & (!n_n4536)));
	assign x22067x = (((!x19x) & (!x572x) & (!n_n5278) & (!n_n5287) & (!n_n5281)) + ((!x19x) & (x572x) & (!n_n5278) & (!n_n5287) & (!n_n5281)) + ((x19x) & (!x572x) & (!n_n5278) & (!n_n5287) & (!n_n5281)));
	assign x16301x = (((!x592x) & (!n_n5296) & (!x21x) & (!x392x) & (n_n5292)) + ((!x592x) & (!n_n5296) & (!x21x) & (x392x) & (!n_n5292)) + ((!x592x) & (!n_n5296) & (!x21x) & (x392x) & (n_n5292)) + ((!x592x) & (!n_n5296) & (x21x) & (!x392x) & (n_n5292)) + ((!x592x) & (!n_n5296) & (x21x) & (x392x) & (!n_n5292)) + ((!x592x) & (!n_n5296) & (x21x) & (x392x) & (n_n5292)) + ((!x592x) & (n_n5296) & (!x21x) & (!x392x) & (!n_n5292)) + ((!x592x) & (n_n5296) & (!x21x) & (!x392x) & (n_n5292)) + ((!x592x) & (n_n5296) & (!x21x) & (x392x) & (!n_n5292)) + ((!x592x) & (n_n5296) & (!x21x) & (x392x) & (n_n5292)) + ((!x592x) & (n_n5296) & (x21x) & (!x392x) & (!n_n5292)) + ((!x592x) & (n_n5296) & (x21x) & (!x392x) & (n_n5292)) + ((!x592x) & (n_n5296) & (x21x) & (x392x) & (!n_n5292)) + ((!x592x) & (n_n5296) & (x21x) & (x392x) & (n_n5292)) + ((x592x) & (!n_n5296) & (!x21x) & (!x392x) & (n_n5292)) + ((x592x) & (!n_n5296) & (!x21x) & (x392x) & (!n_n5292)) + ((x592x) & (!n_n5296) & (!x21x) & (x392x) & (n_n5292)) + ((x592x) & (!n_n5296) & (x21x) & (!x392x) & (!n_n5292)) + ((x592x) & (!n_n5296) & (x21x) & (!x392x) & (n_n5292)) + ((x592x) & (!n_n5296) & (x21x) & (x392x) & (!n_n5292)) + ((x592x) & (!n_n5296) & (x21x) & (x392x) & (n_n5292)) + ((x592x) & (n_n5296) & (!x21x) & (!x392x) & (!n_n5292)) + ((x592x) & (n_n5296) & (!x21x) & (!x392x) & (n_n5292)) + ((x592x) & (n_n5296) & (!x21x) & (x392x) & (!n_n5292)) + ((x592x) & (n_n5296) & (!x21x) & (x392x) & (n_n5292)) + ((x592x) & (n_n5296) & (x21x) & (!x392x) & (!n_n5292)) + ((x592x) & (n_n5296) & (x21x) & (!x392x) & (n_n5292)) + ((x592x) & (n_n5296) & (x21x) & (x392x) & (!n_n5292)) + ((x592x) & (n_n5296) & (x21x) & (x392x) & (n_n5292)));
	assign x16302x = (((!i_9_) & (!n_n532) & (!n_n491) & (!n_n65) & (n_n5271)) + ((!i_9_) & (!n_n532) & (!n_n491) & (n_n65) & (n_n5271)) + ((!i_9_) & (!n_n532) & (n_n491) & (!n_n65) & (n_n5271)) + ((!i_9_) & (!n_n532) & (n_n491) & (n_n65) & (n_n5271)) + ((!i_9_) & (n_n532) & (!n_n491) & (!n_n65) & (n_n5271)) + ((!i_9_) & (n_n532) & (!n_n491) & (n_n65) & (n_n5271)) + ((!i_9_) & (n_n532) & (n_n491) & (!n_n65) & (n_n5271)) + ((!i_9_) & (n_n532) & (n_n491) & (n_n65) & (!n_n5271)) + ((!i_9_) & (n_n532) & (n_n491) & (n_n65) & (n_n5271)) + ((i_9_) & (!n_n532) & (!n_n491) & (!n_n65) & (n_n5271)) + ((i_9_) & (!n_n532) & (!n_n491) & (n_n65) & (n_n5271)) + ((i_9_) & (!n_n532) & (n_n491) & (!n_n65) & (n_n5271)) + ((i_9_) & (!n_n532) & (n_n491) & (n_n65) & (n_n5271)) + ((i_9_) & (n_n532) & (!n_n491) & (!n_n65) & (n_n5271)) + ((i_9_) & (n_n532) & (!n_n491) & (n_n65) & (n_n5271)) + ((i_9_) & (n_n532) & (n_n491) & (!n_n65) & (n_n5271)) + ((i_9_) & (n_n532) & (n_n491) & (n_n65) & (n_n5271)));
	assign x16007x = (((!n_n2059) & (!n_n4465) & (!x11505x) & (!x55x) & (n_n2058)) + ((!n_n2059) & (!n_n4465) & (!x11505x) & (x55x) & (!n_n2058)) + ((!n_n2059) & (!n_n4465) & (!x11505x) & (x55x) & (n_n2058)) + ((!n_n2059) & (!n_n4465) & (x11505x) & (!x55x) & (!n_n2058)) + ((!n_n2059) & (!n_n4465) & (x11505x) & (!x55x) & (n_n2058)) + ((!n_n2059) & (!n_n4465) & (x11505x) & (x55x) & (!n_n2058)) + ((!n_n2059) & (!n_n4465) & (x11505x) & (x55x) & (n_n2058)) + ((!n_n2059) & (n_n4465) & (!x11505x) & (!x55x) & (!n_n2058)) + ((!n_n2059) & (n_n4465) & (!x11505x) & (!x55x) & (n_n2058)) + ((!n_n2059) & (n_n4465) & (!x11505x) & (x55x) & (!n_n2058)) + ((!n_n2059) & (n_n4465) & (!x11505x) & (x55x) & (n_n2058)) + ((!n_n2059) & (n_n4465) & (x11505x) & (!x55x) & (!n_n2058)) + ((!n_n2059) & (n_n4465) & (x11505x) & (!x55x) & (n_n2058)) + ((!n_n2059) & (n_n4465) & (x11505x) & (x55x) & (!n_n2058)) + ((!n_n2059) & (n_n4465) & (x11505x) & (x55x) & (n_n2058)) + ((n_n2059) & (!n_n4465) & (!x11505x) & (!x55x) & (!n_n2058)) + ((n_n2059) & (!n_n4465) & (!x11505x) & (!x55x) & (n_n2058)) + ((n_n2059) & (!n_n4465) & (!x11505x) & (x55x) & (!n_n2058)) + ((n_n2059) & (!n_n4465) & (!x11505x) & (x55x) & (n_n2058)) + ((n_n2059) & (!n_n4465) & (x11505x) & (!x55x) & (!n_n2058)) + ((n_n2059) & (!n_n4465) & (x11505x) & (!x55x) & (n_n2058)) + ((n_n2059) & (!n_n4465) & (x11505x) & (x55x) & (!n_n2058)) + ((n_n2059) & (!n_n4465) & (x11505x) & (x55x) & (n_n2058)) + ((n_n2059) & (n_n4465) & (!x11505x) & (!x55x) & (!n_n2058)) + ((n_n2059) & (n_n4465) & (!x11505x) & (!x55x) & (n_n2058)) + ((n_n2059) & (n_n4465) & (!x11505x) & (x55x) & (!n_n2058)) + ((n_n2059) & (n_n4465) & (!x11505x) & (x55x) & (n_n2058)) + ((n_n2059) & (n_n4465) & (x11505x) & (!x55x) & (!n_n2058)) + ((n_n2059) & (n_n4465) & (x11505x) & (!x55x) & (n_n2058)) + ((n_n2059) & (n_n4465) & (x11505x) & (x55x) & (!n_n2058)) + ((n_n2059) & (n_n4465) & (x11505x) & (x55x) & (n_n2058)));
	assign n_n1889 = (((!n_n4440) & (!n_n4434) & (!n_n4431) & (!n_n4444) & (x16002x)) + ((!n_n4440) & (!n_n4434) & (!n_n4431) & (n_n4444) & (!x16002x)) + ((!n_n4440) & (!n_n4434) & (!n_n4431) & (n_n4444) & (x16002x)) + ((!n_n4440) & (!n_n4434) & (n_n4431) & (!n_n4444) & (!x16002x)) + ((!n_n4440) & (!n_n4434) & (n_n4431) & (!n_n4444) & (x16002x)) + ((!n_n4440) & (!n_n4434) & (n_n4431) & (n_n4444) & (!x16002x)) + ((!n_n4440) & (!n_n4434) & (n_n4431) & (n_n4444) & (x16002x)) + ((!n_n4440) & (n_n4434) & (!n_n4431) & (!n_n4444) & (!x16002x)) + ((!n_n4440) & (n_n4434) & (!n_n4431) & (!n_n4444) & (x16002x)) + ((!n_n4440) & (n_n4434) & (!n_n4431) & (n_n4444) & (!x16002x)) + ((!n_n4440) & (n_n4434) & (!n_n4431) & (n_n4444) & (x16002x)) + ((!n_n4440) & (n_n4434) & (n_n4431) & (!n_n4444) & (!x16002x)) + ((!n_n4440) & (n_n4434) & (n_n4431) & (!n_n4444) & (x16002x)) + ((!n_n4440) & (n_n4434) & (n_n4431) & (n_n4444) & (!x16002x)) + ((!n_n4440) & (n_n4434) & (n_n4431) & (n_n4444) & (x16002x)) + ((n_n4440) & (!n_n4434) & (!n_n4431) & (!n_n4444) & (!x16002x)) + ((n_n4440) & (!n_n4434) & (!n_n4431) & (!n_n4444) & (x16002x)) + ((n_n4440) & (!n_n4434) & (!n_n4431) & (n_n4444) & (!x16002x)) + ((n_n4440) & (!n_n4434) & (!n_n4431) & (n_n4444) & (x16002x)) + ((n_n4440) & (!n_n4434) & (n_n4431) & (!n_n4444) & (!x16002x)) + ((n_n4440) & (!n_n4434) & (n_n4431) & (!n_n4444) & (x16002x)) + ((n_n4440) & (!n_n4434) & (n_n4431) & (n_n4444) & (!x16002x)) + ((n_n4440) & (!n_n4434) & (n_n4431) & (n_n4444) & (x16002x)) + ((n_n4440) & (n_n4434) & (!n_n4431) & (!n_n4444) & (!x16002x)) + ((n_n4440) & (n_n4434) & (!n_n4431) & (!n_n4444) & (x16002x)) + ((n_n4440) & (n_n4434) & (!n_n4431) & (n_n4444) & (!x16002x)) + ((n_n4440) & (n_n4434) & (!n_n4431) & (n_n4444) & (x16002x)) + ((n_n4440) & (n_n4434) & (n_n4431) & (!n_n4444) & (!x16002x)) + ((n_n4440) & (n_n4434) & (n_n4431) & (!n_n4444) & (x16002x)) + ((n_n4440) & (n_n4434) & (n_n4431) & (n_n4444) & (!x16002x)) + ((n_n4440) & (n_n4434) & (n_n4431) & (n_n4444) & (x16002x)));
	assign x16047x = (((!n_n4616) & (!n_n4625) & (!n_n4619) & (!n_n4626) & (n_n4623)) + ((!n_n4616) & (!n_n4625) & (!n_n4619) & (n_n4626) & (!n_n4623)) + ((!n_n4616) & (!n_n4625) & (!n_n4619) & (n_n4626) & (n_n4623)) + ((!n_n4616) & (!n_n4625) & (n_n4619) & (!n_n4626) & (!n_n4623)) + ((!n_n4616) & (!n_n4625) & (n_n4619) & (!n_n4626) & (n_n4623)) + ((!n_n4616) & (!n_n4625) & (n_n4619) & (n_n4626) & (!n_n4623)) + ((!n_n4616) & (!n_n4625) & (n_n4619) & (n_n4626) & (n_n4623)) + ((!n_n4616) & (n_n4625) & (!n_n4619) & (!n_n4626) & (!n_n4623)) + ((!n_n4616) & (n_n4625) & (!n_n4619) & (!n_n4626) & (n_n4623)) + ((!n_n4616) & (n_n4625) & (!n_n4619) & (n_n4626) & (!n_n4623)) + ((!n_n4616) & (n_n4625) & (!n_n4619) & (n_n4626) & (n_n4623)) + ((!n_n4616) & (n_n4625) & (n_n4619) & (!n_n4626) & (!n_n4623)) + ((!n_n4616) & (n_n4625) & (n_n4619) & (!n_n4626) & (n_n4623)) + ((!n_n4616) & (n_n4625) & (n_n4619) & (n_n4626) & (!n_n4623)) + ((!n_n4616) & (n_n4625) & (n_n4619) & (n_n4626) & (n_n4623)) + ((n_n4616) & (!n_n4625) & (!n_n4619) & (!n_n4626) & (!n_n4623)) + ((n_n4616) & (!n_n4625) & (!n_n4619) & (!n_n4626) & (n_n4623)) + ((n_n4616) & (!n_n4625) & (!n_n4619) & (n_n4626) & (!n_n4623)) + ((n_n4616) & (!n_n4625) & (!n_n4619) & (n_n4626) & (n_n4623)) + ((n_n4616) & (!n_n4625) & (n_n4619) & (!n_n4626) & (!n_n4623)) + ((n_n4616) & (!n_n4625) & (n_n4619) & (!n_n4626) & (n_n4623)) + ((n_n4616) & (!n_n4625) & (n_n4619) & (n_n4626) & (!n_n4623)) + ((n_n4616) & (!n_n4625) & (n_n4619) & (n_n4626) & (n_n4623)) + ((n_n4616) & (n_n4625) & (!n_n4619) & (!n_n4626) & (!n_n4623)) + ((n_n4616) & (n_n4625) & (!n_n4619) & (!n_n4626) & (n_n4623)) + ((n_n4616) & (n_n4625) & (!n_n4619) & (n_n4626) & (!n_n4623)) + ((n_n4616) & (n_n4625) & (!n_n4619) & (n_n4626) & (n_n4623)) + ((n_n4616) & (n_n4625) & (n_n4619) & (!n_n4626) & (!n_n4623)) + ((n_n4616) & (n_n4625) & (n_n4619) & (!n_n4626) & (n_n4623)) + ((n_n4616) & (n_n4625) & (n_n4619) & (n_n4626) & (!n_n4623)) + ((n_n4616) & (n_n4625) & (n_n4619) & (n_n4626) & (n_n4623)));
	assign x16064x = (((!x10x) & (!n_n534) & (!n_n491) & (!n_n4635) & (n_n2030)) + ((!x10x) & (!n_n534) & (!n_n491) & (n_n4635) & (!n_n2030)) + ((!x10x) & (!n_n534) & (!n_n491) & (n_n4635) & (n_n2030)) + ((!x10x) & (!n_n534) & (n_n491) & (!n_n4635) & (n_n2030)) + ((!x10x) & (!n_n534) & (n_n491) & (n_n4635) & (!n_n2030)) + ((!x10x) & (!n_n534) & (n_n491) & (n_n4635) & (n_n2030)) + ((!x10x) & (n_n534) & (!n_n491) & (!n_n4635) & (n_n2030)) + ((!x10x) & (n_n534) & (!n_n491) & (n_n4635) & (!n_n2030)) + ((!x10x) & (n_n534) & (!n_n491) & (n_n4635) & (n_n2030)) + ((!x10x) & (n_n534) & (n_n491) & (!n_n4635) & (n_n2030)) + ((!x10x) & (n_n534) & (n_n491) & (n_n4635) & (!n_n2030)) + ((!x10x) & (n_n534) & (n_n491) & (n_n4635) & (n_n2030)) + ((x10x) & (!n_n534) & (!n_n491) & (!n_n4635) & (n_n2030)) + ((x10x) & (!n_n534) & (!n_n491) & (n_n4635) & (!n_n2030)) + ((x10x) & (!n_n534) & (!n_n491) & (n_n4635) & (n_n2030)) + ((x10x) & (!n_n534) & (n_n491) & (!n_n4635) & (n_n2030)) + ((x10x) & (!n_n534) & (n_n491) & (n_n4635) & (!n_n2030)) + ((x10x) & (!n_n534) & (n_n491) & (n_n4635) & (n_n2030)) + ((x10x) & (n_n534) & (!n_n491) & (!n_n4635) & (n_n2030)) + ((x10x) & (n_n534) & (!n_n491) & (n_n4635) & (!n_n2030)) + ((x10x) & (n_n534) & (!n_n491) & (n_n4635) & (n_n2030)) + ((x10x) & (n_n534) & (n_n491) & (!n_n4635) & (!n_n2030)) + ((x10x) & (n_n534) & (n_n491) & (!n_n4635) & (n_n2030)) + ((x10x) & (n_n534) & (n_n491) & (n_n4635) & (!n_n2030)) + ((x10x) & (n_n534) & (n_n491) & (n_n4635) & (n_n2030)));
	assign x16065x = (((!n_n4634) & (!x26x) & (!n_n4633) & (x16064x)) + ((!n_n4634) & (!x26x) & (n_n4633) & (!x16064x)) + ((!n_n4634) & (!x26x) & (n_n4633) & (x16064x)) + ((!n_n4634) & (x26x) & (!n_n4633) & (!x16064x)) + ((!n_n4634) & (x26x) & (!n_n4633) & (x16064x)) + ((!n_n4634) & (x26x) & (n_n4633) & (!x16064x)) + ((!n_n4634) & (x26x) & (n_n4633) & (x16064x)) + ((n_n4634) & (!x26x) & (!n_n4633) & (!x16064x)) + ((n_n4634) & (!x26x) & (!n_n4633) & (x16064x)) + ((n_n4634) & (!x26x) & (n_n4633) & (!x16064x)) + ((n_n4634) & (!x26x) & (n_n4633) & (x16064x)) + ((n_n4634) & (x26x) & (!n_n4633) & (!x16064x)) + ((n_n4634) & (x26x) & (!n_n4633) & (x16064x)) + ((n_n4634) & (x26x) & (n_n4633) & (!x16064x)) + ((n_n4634) & (x26x) & (n_n4633) & (x16064x)));
	assign x16053x = (((!n_n4666) & (!n_n4662) & (!n_n4671) & (n_n4672)) + ((!n_n4666) & (!n_n4662) & (n_n4671) & (!n_n4672)) + ((!n_n4666) & (!n_n4662) & (n_n4671) & (n_n4672)) + ((!n_n4666) & (n_n4662) & (!n_n4671) & (!n_n4672)) + ((!n_n4666) & (n_n4662) & (!n_n4671) & (n_n4672)) + ((!n_n4666) & (n_n4662) & (n_n4671) & (!n_n4672)) + ((!n_n4666) & (n_n4662) & (n_n4671) & (n_n4672)) + ((n_n4666) & (!n_n4662) & (!n_n4671) & (!n_n4672)) + ((n_n4666) & (!n_n4662) & (!n_n4671) & (n_n4672)) + ((n_n4666) & (!n_n4662) & (n_n4671) & (!n_n4672)) + ((n_n4666) & (!n_n4662) & (n_n4671) & (n_n4672)) + ((n_n4666) & (n_n4662) & (!n_n4671) & (!n_n4672)) + ((n_n4666) & (n_n4662) & (!n_n4671) & (n_n4672)) + ((n_n4666) & (n_n4662) & (n_n4671) & (!n_n4672)) + ((n_n4666) & (n_n4662) & (n_n4671) & (n_n4672)));
	assign x16054x = (((!n_n4669) & (!n_n4670) & (!n_n4674) & (!n_n4661) & (n_n4665)) + ((!n_n4669) & (!n_n4670) & (!n_n4674) & (n_n4661) & (!n_n4665)) + ((!n_n4669) & (!n_n4670) & (!n_n4674) & (n_n4661) & (n_n4665)) + ((!n_n4669) & (!n_n4670) & (n_n4674) & (!n_n4661) & (!n_n4665)) + ((!n_n4669) & (!n_n4670) & (n_n4674) & (!n_n4661) & (n_n4665)) + ((!n_n4669) & (!n_n4670) & (n_n4674) & (n_n4661) & (!n_n4665)) + ((!n_n4669) & (!n_n4670) & (n_n4674) & (n_n4661) & (n_n4665)) + ((!n_n4669) & (n_n4670) & (!n_n4674) & (!n_n4661) & (!n_n4665)) + ((!n_n4669) & (n_n4670) & (!n_n4674) & (!n_n4661) & (n_n4665)) + ((!n_n4669) & (n_n4670) & (!n_n4674) & (n_n4661) & (!n_n4665)) + ((!n_n4669) & (n_n4670) & (!n_n4674) & (n_n4661) & (n_n4665)) + ((!n_n4669) & (n_n4670) & (n_n4674) & (!n_n4661) & (!n_n4665)) + ((!n_n4669) & (n_n4670) & (n_n4674) & (!n_n4661) & (n_n4665)) + ((!n_n4669) & (n_n4670) & (n_n4674) & (n_n4661) & (!n_n4665)) + ((!n_n4669) & (n_n4670) & (n_n4674) & (n_n4661) & (n_n4665)) + ((n_n4669) & (!n_n4670) & (!n_n4674) & (!n_n4661) & (!n_n4665)) + ((n_n4669) & (!n_n4670) & (!n_n4674) & (!n_n4661) & (n_n4665)) + ((n_n4669) & (!n_n4670) & (!n_n4674) & (n_n4661) & (!n_n4665)) + ((n_n4669) & (!n_n4670) & (!n_n4674) & (n_n4661) & (n_n4665)) + ((n_n4669) & (!n_n4670) & (n_n4674) & (!n_n4661) & (!n_n4665)) + ((n_n4669) & (!n_n4670) & (n_n4674) & (!n_n4661) & (n_n4665)) + ((n_n4669) & (!n_n4670) & (n_n4674) & (n_n4661) & (!n_n4665)) + ((n_n4669) & (!n_n4670) & (n_n4674) & (n_n4661) & (n_n4665)) + ((n_n4669) & (n_n4670) & (!n_n4674) & (!n_n4661) & (!n_n4665)) + ((n_n4669) & (n_n4670) & (!n_n4674) & (!n_n4661) & (n_n4665)) + ((n_n4669) & (n_n4670) & (!n_n4674) & (n_n4661) & (!n_n4665)) + ((n_n4669) & (n_n4670) & (!n_n4674) & (n_n4661) & (n_n4665)) + ((n_n4669) & (n_n4670) & (n_n4674) & (!n_n4661) & (!n_n4665)) + ((n_n4669) & (n_n4670) & (n_n4674) & (!n_n4661) & (n_n4665)) + ((n_n4669) & (n_n4670) & (n_n4674) & (n_n4661) & (!n_n4665)) + ((n_n4669) & (n_n4670) & (n_n4674) & (n_n4661) & (n_n4665)));
	assign n_n1873 = (((!x309x) & (!n_n4642) & (!n_n4646) & (!n_n4659) & (!x22079x)) + ((!x309x) & (!n_n4642) & (!n_n4646) & (n_n4659) & (!x22079x)) + ((!x309x) & (!n_n4642) & (!n_n4646) & (n_n4659) & (x22079x)) + ((!x309x) & (!n_n4642) & (n_n4646) & (!n_n4659) & (!x22079x)) + ((!x309x) & (!n_n4642) & (n_n4646) & (!n_n4659) & (x22079x)) + ((!x309x) & (!n_n4642) & (n_n4646) & (n_n4659) & (!x22079x)) + ((!x309x) & (!n_n4642) & (n_n4646) & (n_n4659) & (x22079x)) + ((!x309x) & (n_n4642) & (!n_n4646) & (!n_n4659) & (!x22079x)) + ((!x309x) & (n_n4642) & (!n_n4646) & (!n_n4659) & (x22079x)) + ((!x309x) & (n_n4642) & (!n_n4646) & (n_n4659) & (!x22079x)) + ((!x309x) & (n_n4642) & (!n_n4646) & (n_n4659) & (x22079x)) + ((!x309x) & (n_n4642) & (n_n4646) & (!n_n4659) & (!x22079x)) + ((!x309x) & (n_n4642) & (n_n4646) & (!n_n4659) & (x22079x)) + ((!x309x) & (n_n4642) & (n_n4646) & (n_n4659) & (!x22079x)) + ((!x309x) & (n_n4642) & (n_n4646) & (n_n4659) & (x22079x)) + ((x309x) & (!n_n4642) & (!n_n4646) & (!n_n4659) & (!x22079x)) + ((x309x) & (!n_n4642) & (!n_n4646) & (!n_n4659) & (x22079x)) + ((x309x) & (!n_n4642) & (!n_n4646) & (n_n4659) & (!x22079x)) + ((x309x) & (!n_n4642) & (!n_n4646) & (n_n4659) & (x22079x)) + ((x309x) & (!n_n4642) & (n_n4646) & (!n_n4659) & (!x22079x)) + ((x309x) & (!n_n4642) & (n_n4646) & (!n_n4659) & (x22079x)) + ((x309x) & (!n_n4642) & (n_n4646) & (n_n4659) & (!x22079x)) + ((x309x) & (!n_n4642) & (n_n4646) & (n_n4659) & (x22079x)) + ((x309x) & (n_n4642) & (!n_n4646) & (!n_n4659) & (!x22079x)) + ((x309x) & (n_n4642) & (!n_n4646) & (!n_n4659) & (x22079x)) + ((x309x) & (n_n4642) & (!n_n4646) & (n_n4659) & (!x22079x)) + ((x309x) & (n_n4642) & (!n_n4646) & (n_n4659) & (x22079x)) + ((x309x) & (n_n4642) & (n_n4646) & (!n_n4659) & (!x22079x)) + ((x309x) & (n_n4642) & (n_n4646) & (!n_n4659) & (x22079x)) + ((x309x) & (n_n4642) & (n_n4646) & (n_n4659) & (!x22079x)) + ((x309x) & (n_n4642) & (n_n4646) & (n_n4659) & (x22079x)));
	assign x11881x = (((!n_n4652) & (!n_n4656) & (!x140x) & (!n_n4657) & (x431x)) + ((!n_n4652) & (!n_n4656) & (!x140x) & (n_n4657) & (!x431x)) + ((!n_n4652) & (!n_n4656) & (!x140x) & (n_n4657) & (x431x)) + ((!n_n4652) & (!n_n4656) & (x140x) & (!n_n4657) & (!x431x)) + ((!n_n4652) & (!n_n4656) & (x140x) & (!n_n4657) & (x431x)) + ((!n_n4652) & (!n_n4656) & (x140x) & (n_n4657) & (!x431x)) + ((!n_n4652) & (!n_n4656) & (x140x) & (n_n4657) & (x431x)) + ((!n_n4652) & (n_n4656) & (!x140x) & (!n_n4657) & (!x431x)) + ((!n_n4652) & (n_n4656) & (!x140x) & (!n_n4657) & (x431x)) + ((!n_n4652) & (n_n4656) & (!x140x) & (n_n4657) & (!x431x)) + ((!n_n4652) & (n_n4656) & (!x140x) & (n_n4657) & (x431x)) + ((!n_n4652) & (n_n4656) & (x140x) & (!n_n4657) & (!x431x)) + ((!n_n4652) & (n_n4656) & (x140x) & (!n_n4657) & (x431x)) + ((!n_n4652) & (n_n4656) & (x140x) & (n_n4657) & (!x431x)) + ((!n_n4652) & (n_n4656) & (x140x) & (n_n4657) & (x431x)) + ((n_n4652) & (!n_n4656) & (!x140x) & (!n_n4657) & (!x431x)) + ((n_n4652) & (!n_n4656) & (!x140x) & (!n_n4657) & (x431x)) + ((n_n4652) & (!n_n4656) & (!x140x) & (n_n4657) & (!x431x)) + ((n_n4652) & (!n_n4656) & (!x140x) & (n_n4657) & (x431x)) + ((n_n4652) & (!n_n4656) & (x140x) & (!n_n4657) & (!x431x)) + ((n_n4652) & (!n_n4656) & (x140x) & (!n_n4657) & (x431x)) + ((n_n4652) & (!n_n4656) & (x140x) & (n_n4657) & (!x431x)) + ((n_n4652) & (!n_n4656) & (x140x) & (n_n4657) & (x431x)) + ((n_n4652) & (n_n4656) & (!x140x) & (!n_n4657) & (!x431x)) + ((n_n4652) & (n_n4656) & (!x140x) & (!n_n4657) & (x431x)) + ((n_n4652) & (n_n4656) & (!x140x) & (n_n4657) & (!x431x)) + ((n_n4652) & (n_n4656) & (!x140x) & (n_n4657) & (x431x)) + ((n_n4652) & (n_n4656) & (x140x) & (!n_n4657) & (!x431x)) + ((n_n4652) & (n_n4656) & (x140x) & (!n_n4657) & (x431x)) + ((n_n4652) & (n_n4656) & (x140x) & (n_n4657) & (!x431x)) + ((n_n4652) & (n_n4656) & (x140x) & (n_n4657) & (x431x)));
	assign x11882x = (((!n_n4649) & (!n_n4659) & (!x192x) & (n_n1636)) + ((!n_n4649) & (!n_n4659) & (x192x) & (!n_n1636)) + ((!n_n4649) & (!n_n4659) & (x192x) & (n_n1636)) + ((!n_n4649) & (n_n4659) & (!x192x) & (!n_n1636)) + ((!n_n4649) & (n_n4659) & (!x192x) & (n_n1636)) + ((!n_n4649) & (n_n4659) & (x192x) & (!n_n1636)) + ((!n_n4649) & (n_n4659) & (x192x) & (n_n1636)) + ((n_n4649) & (!n_n4659) & (!x192x) & (!n_n1636)) + ((n_n4649) & (!n_n4659) & (!x192x) & (n_n1636)) + ((n_n4649) & (!n_n4659) & (x192x) & (!n_n1636)) + ((n_n4649) & (!n_n4659) & (x192x) & (n_n1636)) + ((n_n4649) & (n_n4659) & (!x192x) & (!n_n1636)) + ((n_n4649) & (n_n4659) & (!x192x) & (n_n1636)) + ((n_n4649) & (n_n4659) & (x192x) & (!n_n1636)) + ((n_n4649) & (n_n4659) & (x192x) & (n_n1636)));
	assign x11884x = (((!x432x) & (!x11859x) & (!x11881x) & (x11882x)) + ((!x432x) & (!x11859x) & (x11881x) & (!x11882x)) + ((!x432x) & (!x11859x) & (x11881x) & (x11882x)) + ((!x432x) & (x11859x) & (!x11881x) & (!x11882x)) + ((!x432x) & (x11859x) & (!x11881x) & (x11882x)) + ((!x432x) & (x11859x) & (x11881x) & (!x11882x)) + ((!x432x) & (x11859x) & (x11881x) & (x11882x)) + ((x432x) & (!x11859x) & (!x11881x) & (!x11882x)) + ((x432x) & (!x11859x) & (!x11881x) & (x11882x)) + ((x432x) & (!x11859x) & (x11881x) & (!x11882x)) + ((x432x) & (!x11859x) & (x11881x) & (x11882x)) + ((x432x) & (x11859x) & (!x11881x) & (!x11882x)) + ((x432x) & (x11859x) & (!x11881x) & (x11882x)) + ((x432x) & (x11859x) & (x11881x) & (!x11882x)) + ((x432x) & (x11859x) & (x11881x) & (x11882x)));
	assign x11850x = (((!n_n4725) & (!n_n4726) & (!x73x) & (!x94x) & (x293x)) + ((!n_n4725) & (!n_n4726) & (!x73x) & (x94x) & (!x293x)) + ((!n_n4725) & (!n_n4726) & (!x73x) & (x94x) & (x293x)) + ((!n_n4725) & (!n_n4726) & (x73x) & (!x94x) & (!x293x)) + ((!n_n4725) & (!n_n4726) & (x73x) & (!x94x) & (x293x)) + ((!n_n4725) & (!n_n4726) & (x73x) & (x94x) & (!x293x)) + ((!n_n4725) & (!n_n4726) & (x73x) & (x94x) & (x293x)) + ((!n_n4725) & (n_n4726) & (!x73x) & (!x94x) & (!x293x)) + ((!n_n4725) & (n_n4726) & (!x73x) & (!x94x) & (x293x)) + ((!n_n4725) & (n_n4726) & (!x73x) & (x94x) & (!x293x)) + ((!n_n4725) & (n_n4726) & (!x73x) & (x94x) & (x293x)) + ((!n_n4725) & (n_n4726) & (x73x) & (!x94x) & (!x293x)) + ((!n_n4725) & (n_n4726) & (x73x) & (!x94x) & (x293x)) + ((!n_n4725) & (n_n4726) & (x73x) & (x94x) & (!x293x)) + ((!n_n4725) & (n_n4726) & (x73x) & (x94x) & (x293x)) + ((n_n4725) & (!n_n4726) & (!x73x) & (!x94x) & (!x293x)) + ((n_n4725) & (!n_n4726) & (!x73x) & (!x94x) & (x293x)) + ((n_n4725) & (!n_n4726) & (!x73x) & (x94x) & (!x293x)) + ((n_n4725) & (!n_n4726) & (!x73x) & (x94x) & (x293x)) + ((n_n4725) & (!n_n4726) & (x73x) & (!x94x) & (!x293x)) + ((n_n4725) & (!n_n4726) & (x73x) & (!x94x) & (x293x)) + ((n_n4725) & (!n_n4726) & (x73x) & (x94x) & (!x293x)) + ((n_n4725) & (!n_n4726) & (x73x) & (x94x) & (x293x)) + ((n_n4725) & (n_n4726) & (!x73x) & (!x94x) & (!x293x)) + ((n_n4725) & (n_n4726) & (!x73x) & (!x94x) & (x293x)) + ((n_n4725) & (n_n4726) & (!x73x) & (x94x) & (!x293x)) + ((n_n4725) & (n_n4726) & (!x73x) & (x94x) & (x293x)) + ((n_n4725) & (n_n4726) & (x73x) & (!x94x) & (!x293x)) + ((n_n4725) & (n_n4726) & (x73x) & (!x94x) & (x293x)) + ((n_n4725) & (n_n4726) & (x73x) & (x94x) & (!x293x)) + ((n_n4725) & (n_n4726) & (x73x) & (x94x) & (x293x)));
	assign x14703x = (((!n_n4806) & (!n_n4810) & (!n_n4805) & (!n_n4813) & (n_n4808)) + ((!n_n4806) & (!n_n4810) & (!n_n4805) & (n_n4813) & (!n_n4808)) + ((!n_n4806) & (!n_n4810) & (!n_n4805) & (n_n4813) & (n_n4808)) + ((!n_n4806) & (!n_n4810) & (n_n4805) & (!n_n4813) & (!n_n4808)) + ((!n_n4806) & (!n_n4810) & (n_n4805) & (!n_n4813) & (n_n4808)) + ((!n_n4806) & (!n_n4810) & (n_n4805) & (n_n4813) & (!n_n4808)) + ((!n_n4806) & (!n_n4810) & (n_n4805) & (n_n4813) & (n_n4808)) + ((!n_n4806) & (n_n4810) & (!n_n4805) & (!n_n4813) & (!n_n4808)) + ((!n_n4806) & (n_n4810) & (!n_n4805) & (!n_n4813) & (n_n4808)) + ((!n_n4806) & (n_n4810) & (!n_n4805) & (n_n4813) & (!n_n4808)) + ((!n_n4806) & (n_n4810) & (!n_n4805) & (n_n4813) & (n_n4808)) + ((!n_n4806) & (n_n4810) & (n_n4805) & (!n_n4813) & (!n_n4808)) + ((!n_n4806) & (n_n4810) & (n_n4805) & (!n_n4813) & (n_n4808)) + ((!n_n4806) & (n_n4810) & (n_n4805) & (n_n4813) & (!n_n4808)) + ((!n_n4806) & (n_n4810) & (n_n4805) & (n_n4813) & (n_n4808)) + ((n_n4806) & (!n_n4810) & (!n_n4805) & (!n_n4813) & (!n_n4808)) + ((n_n4806) & (!n_n4810) & (!n_n4805) & (!n_n4813) & (n_n4808)) + ((n_n4806) & (!n_n4810) & (!n_n4805) & (n_n4813) & (!n_n4808)) + ((n_n4806) & (!n_n4810) & (!n_n4805) & (n_n4813) & (n_n4808)) + ((n_n4806) & (!n_n4810) & (n_n4805) & (!n_n4813) & (!n_n4808)) + ((n_n4806) & (!n_n4810) & (n_n4805) & (!n_n4813) & (n_n4808)) + ((n_n4806) & (!n_n4810) & (n_n4805) & (n_n4813) & (!n_n4808)) + ((n_n4806) & (!n_n4810) & (n_n4805) & (n_n4813) & (n_n4808)) + ((n_n4806) & (n_n4810) & (!n_n4805) & (!n_n4813) & (!n_n4808)) + ((n_n4806) & (n_n4810) & (!n_n4805) & (!n_n4813) & (n_n4808)) + ((n_n4806) & (n_n4810) & (!n_n4805) & (n_n4813) & (!n_n4808)) + ((n_n4806) & (n_n4810) & (!n_n4805) & (n_n4813) & (n_n4808)) + ((n_n4806) & (n_n4810) & (n_n4805) & (!n_n4813) & (!n_n4808)) + ((n_n4806) & (n_n4810) & (n_n4805) & (!n_n4813) & (n_n4808)) + ((n_n4806) & (n_n4810) & (n_n4805) & (n_n4813) & (!n_n4808)) + ((n_n4806) & (n_n4810) & (n_n4805) & (n_n4813) & (n_n4808)));
	assign n_n3701 = (((!n_n4816) & (!n_n4812) & (!n_n4804) & (!n_n4815) & (x14703x)) + ((!n_n4816) & (!n_n4812) & (!n_n4804) & (n_n4815) & (!x14703x)) + ((!n_n4816) & (!n_n4812) & (!n_n4804) & (n_n4815) & (x14703x)) + ((!n_n4816) & (!n_n4812) & (n_n4804) & (!n_n4815) & (!x14703x)) + ((!n_n4816) & (!n_n4812) & (n_n4804) & (!n_n4815) & (x14703x)) + ((!n_n4816) & (!n_n4812) & (n_n4804) & (n_n4815) & (!x14703x)) + ((!n_n4816) & (!n_n4812) & (n_n4804) & (n_n4815) & (x14703x)) + ((!n_n4816) & (n_n4812) & (!n_n4804) & (!n_n4815) & (!x14703x)) + ((!n_n4816) & (n_n4812) & (!n_n4804) & (!n_n4815) & (x14703x)) + ((!n_n4816) & (n_n4812) & (!n_n4804) & (n_n4815) & (!x14703x)) + ((!n_n4816) & (n_n4812) & (!n_n4804) & (n_n4815) & (x14703x)) + ((!n_n4816) & (n_n4812) & (n_n4804) & (!n_n4815) & (!x14703x)) + ((!n_n4816) & (n_n4812) & (n_n4804) & (!n_n4815) & (x14703x)) + ((!n_n4816) & (n_n4812) & (n_n4804) & (n_n4815) & (!x14703x)) + ((!n_n4816) & (n_n4812) & (n_n4804) & (n_n4815) & (x14703x)) + ((n_n4816) & (!n_n4812) & (!n_n4804) & (!n_n4815) & (!x14703x)) + ((n_n4816) & (!n_n4812) & (!n_n4804) & (!n_n4815) & (x14703x)) + ((n_n4816) & (!n_n4812) & (!n_n4804) & (n_n4815) & (!x14703x)) + ((n_n4816) & (!n_n4812) & (!n_n4804) & (n_n4815) & (x14703x)) + ((n_n4816) & (!n_n4812) & (n_n4804) & (!n_n4815) & (!x14703x)) + ((n_n4816) & (!n_n4812) & (n_n4804) & (!n_n4815) & (x14703x)) + ((n_n4816) & (!n_n4812) & (n_n4804) & (n_n4815) & (!x14703x)) + ((n_n4816) & (!n_n4812) & (n_n4804) & (n_n4815) & (x14703x)) + ((n_n4816) & (n_n4812) & (!n_n4804) & (!n_n4815) & (!x14703x)) + ((n_n4816) & (n_n4812) & (!n_n4804) & (!n_n4815) & (x14703x)) + ((n_n4816) & (n_n4812) & (!n_n4804) & (n_n4815) & (!x14703x)) + ((n_n4816) & (n_n4812) & (!n_n4804) & (n_n4815) & (x14703x)) + ((n_n4816) & (n_n4812) & (n_n4804) & (!n_n4815) & (!x14703x)) + ((n_n4816) & (n_n4812) & (n_n4804) & (!n_n4815) & (x14703x)) + ((n_n4816) & (n_n4812) & (n_n4804) & (n_n4815) & (!x14703x)) + ((n_n4816) & (n_n4812) & (n_n4804) & (n_n4815) & (x14703x)));
	assign x14708x = (((!x23x) & (!x530x) & (!n_n4817) & (!n_n4828) & (n_n4820)) + ((!x23x) & (!x530x) & (!n_n4817) & (n_n4828) & (!n_n4820)) + ((!x23x) & (!x530x) & (!n_n4817) & (n_n4828) & (n_n4820)) + ((!x23x) & (!x530x) & (n_n4817) & (!n_n4828) & (!n_n4820)) + ((!x23x) & (!x530x) & (n_n4817) & (!n_n4828) & (n_n4820)) + ((!x23x) & (!x530x) & (n_n4817) & (n_n4828) & (!n_n4820)) + ((!x23x) & (!x530x) & (n_n4817) & (n_n4828) & (n_n4820)) + ((!x23x) & (x530x) & (!n_n4817) & (!n_n4828) & (n_n4820)) + ((!x23x) & (x530x) & (!n_n4817) & (n_n4828) & (!n_n4820)) + ((!x23x) & (x530x) & (!n_n4817) & (n_n4828) & (n_n4820)) + ((!x23x) & (x530x) & (n_n4817) & (!n_n4828) & (!n_n4820)) + ((!x23x) & (x530x) & (n_n4817) & (!n_n4828) & (n_n4820)) + ((!x23x) & (x530x) & (n_n4817) & (n_n4828) & (!n_n4820)) + ((!x23x) & (x530x) & (n_n4817) & (n_n4828) & (n_n4820)) + ((x23x) & (!x530x) & (!n_n4817) & (!n_n4828) & (n_n4820)) + ((x23x) & (!x530x) & (!n_n4817) & (n_n4828) & (!n_n4820)) + ((x23x) & (!x530x) & (!n_n4817) & (n_n4828) & (n_n4820)) + ((x23x) & (!x530x) & (n_n4817) & (!n_n4828) & (!n_n4820)) + ((x23x) & (!x530x) & (n_n4817) & (!n_n4828) & (n_n4820)) + ((x23x) & (!x530x) & (n_n4817) & (n_n4828) & (!n_n4820)) + ((x23x) & (!x530x) & (n_n4817) & (n_n4828) & (n_n4820)) + ((x23x) & (x530x) & (!n_n4817) & (!n_n4828) & (!n_n4820)) + ((x23x) & (x530x) & (!n_n4817) & (!n_n4828) & (n_n4820)) + ((x23x) & (x530x) & (!n_n4817) & (n_n4828) & (!n_n4820)) + ((x23x) & (x530x) & (!n_n4817) & (n_n4828) & (n_n4820)) + ((x23x) & (x530x) & (n_n4817) & (!n_n4828) & (!n_n4820)) + ((x23x) & (x530x) & (n_n4817) & (!n_n4828) & (n_n4820)) + ((x23x) & (x530x) & (n_n4817) & (n_n4828) & (!n_n4820)) + ((x23x) & (x530x) & (n_n4817) & (n_n4828) & (n_n4820)));
	assign x14709x = (((!n_n4826) & (!n_n4821) & (!n_n4822) & (!n_n4818) & (n_n4819)) + ((!n_n4826) & (!n_n4821) & (!n_n4822) & (n_n4818) & (!n_n4819)) + ((!n_n4826) & (!n_n4821) & (!n_n4822) & (n_n4818) & (n_n4819)) + ((!n_n4826) & (!n_n4821) & (n_n4822) & (!n_n4818) & (!n_n4819)) + ((!n_n4826) & (!n_n4821) & (n_n4822) & (!n_n4818) & (n_n4819)) + ((!n_n4826) & (!n_n4821) & (n_n4822) & (n_n4818) & (!n_n4819)) + ((!n_n4826) & (!n_n4821) & (n_n4822) & (n_n4818) & (n_n4819)) + ((!n_n4826) & (n_n4821) & (!n_n4822) & (!n_n4818) & (!n_n4819)) + ((!n_n4826) & (n_n4821) & (!n_n4822) & (!n_n4818) & (n_n4819)) + ((!n_n4826) & (n_n4821) & (!n_n4822) & (n_n4818) & (!n_n4819)) + ((!n_n4826) & (n_n4821) & (!n_n4822) & (n_n4818) & (n_n4819)) + ((!n_n4826) & (n_n4821) & (n_n4822) & (!n_n4818) & (!n_n4819)) + ((!n_n4826) & (n_n4821) & (n_n4822) & (!n_n4818) & (n_n4819)) + ((!n_n4826) & (n_n4821) & (n_n4822) & (n_n4818) & (!n_n4819)) + ((!n_n4826) & (n_n4821) & (n_n4822) & (n_n4818) & (n_n4819)) + ((n_n4826) & (!n_n4821) & (!n_n4822) & (!n_n4818) & (!n_n4819)) + ((n_n4826) & (!n_n4821) & (!n_n4822) & (!n_n4818) & (n_n4819)) + ((n_n4826) & (!n_n4821) & (!n_n4822) & (n_n4818) & (!n_n4819)) + ((n_n4826) & (!n_n4821) & (!n_n4822) & (n_n4818) & (n_n4819)) + ((n_n4826) & (!n_n4821) & (n_n4822) & (!n_n4818) & (!n_n4819)) + ((n_n4826) & (!n_n4821) & (n_n4822) & (!n_n4818) & (n_n4819)) + ((n_n4826) & (!n_n4821) & (n_n4822) & (n_n4818) & (!n_n4819)) + ((n_n4826) & (!n_n4821) & (n_n4822) & (n_n4818) & (n_n4819)) + ((n_n4826) & (n_n4821) & (!n_n4822) & (!n_n4818) & (!n_n4819)) + ((n_n4826) & (n_n4821) & (!n_n4822) & (!n_n4818) & (n_n4819)) + ((n_n4826) & (n_n4821) & (!n_n4822) & (n_n4818) & (!n_n4819)) + ((n_n4826) & (n_n4821) & (!n_n4822) & (n_n4818) & (n_n4819)) + ((n_n4826) & (n_n4821) & (n_n4822) & (!n_n4818) & (!n_n4819)) + ((n_n4826) & (n_n4821) & (n_n4822) & (!n_n4818) & (n_n4819)) + ((n_n4826) & (n_n4821) & (n_n4822) & (n_n4818) & (!n_n4819)) + ((n_n4826) & (n_n4821) & (n_n4822) & (n_n4818) & (n_n4819)));
	assign x22110x = (((!n_n4832) & (!n_n3820) & (!n_n4837) & (!x38x) & (!x303x)));
	assign x14562x = (((!i_9_) & (!n_n524) & (!n_n482) & (!n_n65) & (n_n5302)) + ((!i_9_) & (!n_n524) & (!n_n482) & (n_n65) & (n_n5302)) + ((!i_9_) & (!n_n524) & (n_n482) & (!n_n65) & (n_n5302)) + ((!i_9_) & (!n_n524) & (n_n482) & (n_n65) & (n_n5302)) + ((!i_9_) & (n_n524) & (!n_n482) & (!n_n65) & (n_n5302)) + ((!i_9_) & (n_n524) & (!n_n482) & (n_n65) & (n_n5302)) + ((!i_9_) & (n_n524) & (n_n482) & (!n_n65) & (n_n5302)) + ((!i_9_) & (n_n524) & (n_n482) & (n_n65) & (!n_n5302)) + ((!i_9_) & (n_n524) & (n_n482) & (n_n65) & (n_n5302)) + ((i_9_) & (!n_n524) & (!n_n482) & (!n_n65) & (n_n5302)) + ((i_9_) & (!n_n524) & (!n_n482) & (n_n65) & (n_n5302)) + ((i_9_) & (!n_n524) & (n_n482) & (!n_n65) & (n_n5302)) + ((i_9_) & (!n_n524) & (n_n482) & (n_n65) & (n_n5302)) + ((i_9_) & (n_n524) & (!n_n482) & (!n_n65) & (n_n5302)) + ((i_9_) & (n_n524) & (!n_n482) & (n_n65) & (n_n5302)) + ((i_9_) & (n_n524) & (n_n482) & (!n_n65) & (n_n5302)) + ((i_9_) & (n_n524) & (n_n482) & (n_n65) & (n_n5302)));
	assign x14572x = (((!n_n5240) & (!n_n5238) & (!n_n5244) & (n_n5233)) + ((!n_n5240) & (!n_n5238) & (n_n5244) & (!n_n5233)) + ((!n_n5240) & (!n_n5238) & (n_n5244) & (n_n5233)) + ((!n_n5240) & (n_n5238) & (!n_n5244) & (!n_n5233)) + ((!n_n5240) & (n_n5238) & (!n_n5244) & (n_n5233)) + ((!n_n5240) & (n_n5238) & (n_n5244) & (!n_n5233)) + ((!n_n5240) & (n_n5238) & (n_n5244) & (n_n5233)) + ((n_n5240) & (!n_n5238) & (!n_n5244) & (!n_n5233)) + ((n_n5240) & (!n_n5238) & (!n_n5244) & (n_n5233)) + ((n_n5240) & (!n_n5238) & (n_n5244) & (!n_n5233)) + ((n_n5240) & (!n_n5238) & (n_n5244) & (n_n5233)) + ((n_n5240) & (n_n5238) & (!n_n5244) & (!n_n5233)) + ((n_n5240) & (n_n5238) & (!n_n5244) & (n_n5233)) + ((n_n5240) & (n_n5238) & (n_n5244) & (!n_n5233)) + ((n_n5240) & (n_n5238) & (n_n5244) & (n_n5233)));
	assign x14573x = (((!n_n5241) & (!n_n5242) & (!n_n5229) & (!n_n5235) & (n_n5234)) + ((!n_n5241) & (!n_n5242) & (!n_n5229) & (n_n5235) & (!n_n5234)) + ((!n_n5241) & (!n_n5242) & (!n_n5229) & (n_n5235) & (n_n5234)) + ((!n_n5241) & (!n_n5242) & (n_n5229) & (!n_n5235) & (!n_n5234)) + ((!n_n5241) & (!n_n5242) & (n_n5229) & (!n_n5235) & (n_n5234)) + ((!n_n5241) & (!n_n5242) & (n_n5229) & (n_n5235) & (!n_n5234)) + ((!n_n5241) & (!n_n5242) & (n_n5229) & (n_n5235) & (n_n5234)) + ((!n_n5241) & (n_n5242) & (!n_n5229) & (!n_n5235) & (!n_n5234)) + ((!n_n5241) & (n_n5242) & (!n_n5229) & (!n_n5235) & (n_n5234)) + ((!n_n5241) & (n_n5242) & (!n_n5229) & (n_n5235) & (!n_n5234)) + ((!n_n5241) & (n_n5242) & (!n_n5229) & (n_n5235) & (n_n5234)) + ((!n_n5241) & (n_n5242) & (n_n5229) & (!n_n5235) & (!n_n5234)) + ((!n_n5241) & (n_n5242) & (n_n5229) & (!n_n5235) & (n_n5234)) + ((!n_n5241) & (n_n5242) & (n_n5229) & (n_n5235) & (!n_n5234)) + ((!n_n5241) & (n_n5242) & (n_n5229) & (n_n5235) & (n_n5234)) + ((n_n5241) & (!n_n5242) & (!n_n5229) & (!n_n5235) & (!n_n5234)) + ((n_n5241) & (!n_n5242) & (!n_n5229) & (!n_n5235) & (n_n5234)) + ((n_n5241) & (!n_n5242) & (!n_n5229) & (n_n5235) & (!n_n5234)) + ((n_n5241) & (!n_n5242) & (!n_n5229) & (n_n5235) & (n_n5234)) + ((n_n5241) & (!n_n5242) & (n_n5229) & (!n_n5235) & (!n_n5234)) + ((n_n5241) & (!n_n5242) & (n_n5229) & (!n_n5235) & (n_n5234)) + ((n_n5241) & (!n_n5242) & (n_n5229) & (n_n5235) & (!n_n5234)) + ((n_n5241) & (!n_n5242) & (n_n5229) & (n_n5235) & (n_n5234)) + ((n_n5241) & (n_n5242) & (!n_n5229) & (!n_n5235) & (!n_n5234)) + ((n_n5241) & (n_n5242) & (!n_n5229) & (!n_n5235) & (n_n5234)) + ((n_n5241) & (n_n5242) & (!n_n5229) & (n_n5235) & (!n_n5234)) + ((n_n5241) & (n_n5242) & (!n_n5229) & (n_n5235) & (n_n5234)) + ((n_n5241) & (n_n5242) & (n_n5229) & (!n_n5235) & (!n_n5234)) + ((n_n5241) & (n_n5242) & (n_n5229) & (!n_n5235) & (n_n5234)) + ((n_n5241) & (n_n5242) & (n_n5229) & (n_n5235) & (!n_n5234)) + ((n_n5241) & (n_n5242) & (n_n5229) & (n_n5235) & (n_n5234)));
	assign x14579x = (((!n_n5245) & (!n_n5254) & (!n_n5217) & (n_n5248)) + ((!n_n5245) & (!n_n5254) & (n_n5217) & (!n_n5248)) + ((!n_n5245) & (!n_n5254) & (n_n5217) & (n_n5248)) + ((!n_n5245) & (n_n5254) & (!n_n5217) & (!n_n5248)) + ((!n_n5245) & (n_n5254) & (!n_n5217) & (n_n5248)) + ((!n_n5245) & (n_n5254) & (n_n5217) & (!n_n5248)) + ((!n_n5245) & (n_n5254) & (n_n5217) & (n_n5248)) + ((n_n5245) & (!n_n5254) & (!n_n5217) & (!n_n5248)) + ((n_n5245) & (!n_n5254) & (!n_n5217) & (n_n5248)) + ((n_n5245) & (!n_n5254) & (n_n5217) & (!n_n5248)) + ((n_n5245) & (!n_n5254) & (n_n5217) & (n_n5248)) + ((n_n5245) & (n_n5254) & (!n_n5217) & (!n_n5248)) + ((n_n5245) & (n_n5254) & (!n_n5217) & (n_n5248)) + ((n_n5245) & (n_n5254) & (n_n5217) & (!n_n5248)) + ((n_n5245) & (n_n5254) & (n_n5217) & (n_n5248)));
	assign x14580x = (((!n_n5247) & (!n_n5246) & (!n_n5227) & (n_n761)) + ((!n_n5247) & (!n_n5246) & (n_n5227) & (!n_n761)) + ((!n_n5247) & (!n_n5246) & (n_n5227) & (n_n761)) + ((!n_n5247) & (n_n5246) & (!n_n5227) & (!n_n761)) + ((!n_n5247) & (n_n5246) & (!n_n5227) & (n_n761)) + ((!n_n5247) & (n_n5246) & (n_n5227) & (!n_n761)) + ((!n_n5247) & (n_n5246) & (n_n5227) & (n_n761)) + ((n_n5247) & (!n_n5246) & (!n_n5227) & (!n_n761)) + ((n_n5247) & (!n_n5246) & (!n_n5227) & (n_n761)) + ((n_n5247) & (!n_n5246) & (n_n5227) & (!n_n761)) + ((n_n5247) & (!n_n5246) & (n_n5227) & (n_n761)) + ((n_n5247) & (n_n5246) & (!n_n5227) & (!n_n761)) + ((n_n5247) & (n_n5246) & (!n_n5227) & (n_n761)) + ((n_n5247) & (n_n5246) & (n_n5227) & (!n_n761)) + ((n_n5247) & (n_n5246) & (n_n5227) & (n_n761)));
	assign x14581x = (((!n_n5258) & (!n_n5259) & (!x383x) & (!x183x) & (x434x)) + ((!n_n5258) & (!n_n5259) & (!x383x) & (x183x) & (!x434x)) + ((!n_n5258) & (!n_n5259) & (!x383x) & (x183x) & (x434x)) + ((!n_n5258) & (!n_n5259) & (x383x) & (!x183x) & (!x434x)) + ((!n_n5258) & (!n_n5259) & (x383x) & (!x183x) & (x434x)) + ((!n_n5258) & (!n_n5259) & (x383x) & (x183x) & (!x434x)) + ((!n_n5258) & (!n_n5259) & (x383x) & (x183x) & (x434x)) + ((!n_n5258) & (n_n5259) & (!x383x) & (!x183x) & (!x434x)) + ((!n_n5258) & (n_n5259) & (!x383x) & (!x183x) & (x434x)) + ((!n_n5258) & (n_n5259) & (!x383x) & (x183x) & (!x434x)) + ((!n_n5258) & (n_n5259) & (!x383x) & (x183x) & (x434x)) + ((!n_n5258) & (n_n5259) & (x383x) & (!x183x) & (!x434x)) + ((!n_n5258) & (n_n5259) & (x383x) & (!x183x) & (x434x)) + ((!n_n5258) & (n_n5259) & (x383x) & (x183x) & (!x434x)) + ((!n_n5258) & (n_n5259) & (x383x) & (x183x) & (x434x)) + ((n_n5258) & (!n_n5259) & (!x383x) & (!x183x) & (!x434x)) + ((n_n5258) & (!n_n5259) & (!x383x) & (!x183x) & (x434x)) + ((n_n5258) & (!n_n5259) & (!x383x) & (x183x) & (!x434x)) + ((n_n5258) & (!n_n5259) & (!x383x) & (x183x) & (x434x)) + ((n_n5258) & (!n_n5259) & (x383x) & (!x183x) & (!x434x)) + ((n_n5258) & (!n_n5259) & (x383x) & (!x183x) & (x434x)) + ((n_n5258) & (!n_n5259) & (x383x) & (x183x) & (!x434x)) + ((n_n5258) & (!n_n5259) & (x383x) & (x183x) & (x434x)) + ((n_n5258) & (n_n5259) & (!x383x) & (!x183x) & (!x434x)) + ((n_n5258) & (n_n5259) & (!x383x) & (!x183x) & (x434x)) + ((n_n5258) & (n_n5259) & (!x383x) & (x183x) & (!x434x)) + ((n_n5258) & (n_n5259) & (!x383x) & (x183x) & (x434x)) + ((n_n5258) & (n_n5259) & (x383x) & (!x183x) & (!x434x)) + ((n_n5258) & (n_n5259) & (x383x) & (!x183x) & (x434x)) + ((n_n5258) & (n_n5259) & (x383x) & (x183x) & (!x434x)) + ((n_n5258) & (n_n5259) & (x383x) & (x183x) & (x434x)));
	assign x16267x = (((!n_n5244) & (!n_n5241) & (!n_n5236) & (n_n5237)) + ((!n_n5244) & (!n_n5241) & (n_n5236) & (!n_n5237)) + ((!n_n5244) & (!n_n5241) & (n_n5236) & (n_n5237)) + ((!n_n5244) & (n_n5241) & (!n_n5236) & (!n_n5237)) + ((!n_n5244) & (n_n5241) & (!n_n5236) & (n_n5237)) + ((!n_n5244) & (n_n5241) & (n_n5236) & (!n_n5237)) + ((!n_n5244) & (n_n5241) & (n_n5236) & (n_n5237)) + ((n_n5244) & (!n_n5241) & (!n_n5236) & (!n_n5237)) + ((n_n5244) & (!n_n5241) & (!n_n5236) & (n_n5237)) + ((n_n5244) & (!n_n5241) & (n_n5236) & (!n_n5237)) + ((n_n5244) & (!n_n5241) & (n_n5236) & (n_n5237)) + ((n_n5244) & (n_n5241) & (!n_n5236) & (!n_n5237)) + ((n_n5244) & (n_n5241) & (!n_n5236) & (n_n5237)) + ((n_n5244) & (n_n5241) & (n_n5236) & (!n_n5237)) + ((n_n5244) & (n_n5241) & (n_n5236) & (n_n5237)));
	assign x16268x = (((!n_n5239) & (!n_n5240) & (!n_n5242) & (!n_n5246) & (n_n5234)) + ((!n_n5239) & (!n_n5240) & (!n_n5242) & (n_n5246) & (!n_n5234)) + ((!n_n5239) & (!n_n5240) & (!n_n5242) & (n_n5246) & (n_n5234)) + ((!n_n5239) & (!n_n5240) & (n_n5242) & (!n_n5246) & (!n_n5234)) + ((!n_n5239) & (!n_n5240) & (n_n5242) & (!n_n5246) & (n_n5234)) + ((!n_n5239) & (!n_n5240) & (n_n5242) & (n_n5246) & (!n_n5234)) + ((!n_n5239) & (!n_n5240) & (n_n5242) & (n_n5246) & (n_n5234)) + ((!n_n5239) & (n_n5240) & (!n_n5242) & (!n_n5246) & (!n_n5234)) + ((!n_n5239) & (n_n5240) & (!n_n5242) & (!n_n5246) & (n_n5234)) + ((!n_n5239) & (n_n5240) & (!n_n5242) & (n_n5246) & (!n_n5234)) + ((!n_n5239) & (n_n5240) & (!n_n5242) & (n_n5246) & (n_n5234)) + ((!n_n5239) & (n_n5240) & (n_n5242) & (!n_n5246) & (!n_n5234)) + ((!n_n5239) & (n_n5240) & (n_n5242) & (!n_n5246) & (n_n5234)) + ((!n_n5239) & (n_n5240) & (n_n5242) & (n_n5246) & (!n_n5234)) + ((!n_n5239) & (n_n5240) & (n_n5242) & (n_n5246) & (n_n5234)) + ((n_n5239) & (!n_n5240) & (!n_n5242) & (!n_n5246) & (!n_n5234)) + ((n_n5239) & (!n_n5240) & (!n_n5242) & (!n_n5246) & (n_n5234)) + ((n_n5239) & (!n_n5240) & (!n_n5242) & (n_n5246) & (!n_n5234)) + ((n_n5239) & (!n_n5240) & (!n_n5242) & (n_n5246) & (n_n5234)) + ((n_n5239) & (!n_n5240) & (n_n5242) & (!n_n5246) & (!n_n5234)) + ((n_n5239) & (!n_n5240) & (n_n5242) & (!n_n5246) & (n_n5234)) + ((n_n5239) & (!n_n5240) & (n_n5242) & (n_n5246) & (!n_n5234)) + ((n_n5239) & (!n_n5240) & (n_n5242) & (n_n5246) & (n_n5234)) + ((n_n5239) & (n_n5240) & (!n_n5242) & (!n_n5246) & (!n_n5234)) + ((n_n5239) & (n_n5240) & (!n_n5242) & (!n_n5246) & (n_n5234)) + ((n_n5239) & (n_n5240) & (!n_n5242) & (n_n5246) & (!n_n5234)) + ((n_n5239) & (n_n5240) & (!n_n5242) & (n_n5246) & (n_n5234)) + ((n_n5239) & (n_n5240) & (n_n5242) & (!n_n5246) & (!n_n5234)) + ((n_n5239) & (n_n5240) & (n_n5242) & (!n_n5246) & (n_n5234)) + ((n_n5239) & (n_n5240) & (n_n5242) & (n_n5246) & (!n_n5234)) + ((n_n5239) & (n_n5240) & (n_n5242) & (n_n5246) & (n_n5234)));
	assign x16273x = (((!n_n5226) & (!n_n5225) & (!n_n5224) & (!n_n5227) & (n_n5215)) + ((!n_n5226) & (!n_n5225) & (!n_n5224) & (n_n5227) & (!n_n5215)) + ((!n_n5226) & (!n_n5225) & (!n_n5224) & (n_n5227) & (n_n5215)) + ((!n_n5226) & (!n_n5225) & (n_n5224) & (!n_n5227) & (!n_n5215)) + ((!n_n5226) & (!n_n5225) & (n_n5224) & (!n_n5227) & (n_n5215)) + ((!n_n5226) & (!n_n5225) & (n_n5224) & (n_n5227) & (!n_n5215)) + ((!n_n5226) & (!n_n5225) & (n_n5224) & (n_n5227) & (n_n5215)) + ((!n_n5226) & (n_n5225) & (!n_n5224) & (!n_n5227) & (!n_n5215)) + ((!n_n5226) & (n_n5225) & (!n_n5224) & (!n_n5227) & (n_n5215)) + ((!n_n5226) & (n_n5225) & (!n_n5224) & (n_n5227) & (!n_n5215)) + ((!n_n5226) & (n_n5225) & (!n_n5224) & (n_n5227) & (n_n5215)) + ((!n_n5226) & (n_n5225) & (n_n5224) & (!n_n5227) & (!n_n5215)) + ((!n_n5226) & (n_n5225) & (n_n5224) & (!n_n5227) & (n_n5215)) + ((!n_n5226) & (n_n5225) & (n_n5224) & (n_n5227) & (!n_n5215)) + ((!n_n5226) & (n_n5225) & (n_n5224) & (n_n5227) & (n_n5215)) + ((n_n5226) & (!n_n5225) & (!n_n5224) & (!n_n5227) & (!n_n5215)) + ((n_n5226) & (!n_n5225) & (!n_n5224) & (!n_n5227) & (n_n5215)) + ((n_n5226) & (!n_n5225) & (!n_n5224) & (n_n5227) & (!n_n5215)) + ((n_n5226) & (!n_n5225) & (!n_n5224) & (n_n5227) & (n_n5215)) + ((n_n5226) & (!n_n5225) & (n_n5224) & (!n_n5227) & (!n_n5215)) + ((n_n5226) & (!n_n5225) & (n_n5224) & (!n_n5227) & (n_n5215)) + ((n_n5226) & (!n_n5225) & (n_n5224) & (n_n5227) & (!n_n5215)) + ((n_n5226) & (!n_n5225) & (n_n5224) & (n_n5227) & (n_n5215)) + ((n_n5226) & (n_n5225) & (!n_n5224) & (!n_n5227) & (!n_n5215)) + ((n_n5226) & (n_n5225) & (!n_n5224) & (!n_n5227) & (n_n5215)) + ((n_n5226) & (n_n5225) & (!n_n5224) & (n_n5227) & (!n_n5215)) + ((n_n5226) & (n_n5225) & (!n_n5224) & (n_n5227) & (n_n5215)) + ((n_n5226) & (n_n5225) & (n_n5224) & (!n_n5227) & (!n_n5215)) + ((n_n5226) & (n_n5225) & (n_n5224) & (!n_n5227) & (n_n5215)) + ((n_n5226) & (n_n5225) & (n_n5224) & (n_n5227) & (!n_n5215)) + ((n_n5226) & (n_n5225) & (n_n5224) & (n_n5227) & (n_n5215)));
	assign n_n1829 = (((!n_n5232) & (!n_n5233) & (!n_n5228) & (!n_n5220) & (x16273x)) + ((!n_n5232) & (!n_n5233) & (!n_n5228) & (n_n5220) & (!x16273x)) + ((!n_n5232) & (!n_n5233) & (!n_n5228) & (n_n5220) & (x16273x)) + ((!n_n5232) & (!n_n5233) & (n_n5228) & (!n_n5220) & (!x16273x)) + ((!n_n5232) & (!n_n5233) & (n_n5228) & (!n_n5220) & (x16273x)) + ((!n_n5232) & (!n_n5233) & (n_n5228) & (n_n5220) & (!x16273x)) + ((!n_n5232) & (!n_n5233) & (n_n5228) & (n_n5220) & (x16273x)) + ((!n_n5232) & (n_n5233) & (!n_n5228) & (!n_n5220) & (!x16273x)) + ((!n_n5232) & (n_n5233) & (!n_n5228) & (!n_n5220) & (x16273x)) + ((!n_n5232) & (n_n5233) & (!n_n5228) & (n_n5220) & (!x16273x)) + ((!n_n5232) & (n_n5233) & (!n_n5228) & (n_n5220) & (x16273x)) + ((!n_n5232) & (n_n5233) & (n_n5228) & (!n_n5220) & (!x16273x)) + ((!n_n5232) & (n_n5233) & (n_n5228) & (!n_n5220) & (x16273x)) + ((!n_n5232) & (n_n5233) & (n_n5228) & (n_n5220) & (!x16273x)) + ((!n_n5232) & (n_n5233) & (n_n5228) & (n_n5220) & (x16273x)) + ((n_n5232) & (!n_n5233) & (!n_n5228) & (!n_n5220) & (!x16273x)) + ((n_n5232) & (!n_n5233) & (!n_n5228) & (!n_n5220) & (x16273x)) + ((n_n5232) & (!n_n5233) & (!n_n5228) & (n_n5220) & (!x16273x)) + ((n_n5232) & (!n_n5233) & (!n_n5228) & (n_n5220) & (x16273x)) + ((n_n5232) & (!n_n5233) & (n_n5228) & (!n_n5220) & (!x16273x)) + ((n_n5232) & (!n_n5233) & (n_n5228) & (!n_n5220) & (x16273x)) + ((n_n5232) & (!n_n5233) & (n_n5228) & (n_n5220) & (!x16273x)) + ((n_n5232) & (!n_n5233) & (n_n5228) & (n_n5220) & (x16273x)) + ((n_n5232) & (n_n5233) & (!n_n5228) & (!n_n5220) & (!x16273x)) + ((n_n5232) & (n_n5233) & (!n_n5228) & (!n_n5220) & (x16273x)) + ((n_n5232) & (n_n5233) & (!n_n5228) & (n_n5220) & (!x16273x)) + ((n_n5232) & (n_n5233) & (!n_n5228) & (n_n5220) & (x16273x)) + ((n_n5232) & (n_n5233) & (n_n5228) & (!n_n5220) & (!x16273x)) + ((n_n5232) & (n_n5233) & (n_n5228) & (!n_n5220) & (x16273x)) + ((n_n5232) & (n_n5233) & (n_n5228) & (n_n5220) & (!x16273x)) + ((n_n5232) & (n_n5233) & (n_n5228) & (n_n5220) & (x16273x)));
	assign x16278x = (((!n_n5258) & (!n_n5251) & (!n_n5249) & (n_n5252)) + ((!n_n5258) & (!n_n5251) & (n_n5249) & (!n_n5252)) + ((!n_n5258) & (!n_n5251) & (n_n5249) & (n_n5252)) + ((!n_n5258) & (n_n5251) & (!n_n5249) & (!n_n5252)) + ((!n_n5258) & (n_n5251) & (!n_n5249) & (n_n5252)) + ((!n_n5258) & (n_n5251) & (n_n5249) & (!n_n5252)) + ((!n_n5258) & (n_n5251) & (n_n5249) & (n_n5252)) + ((n_n5258) & (!n_n5251) & (!n_n5249) & (!n_n5252)) + ((n_n5258) & (!n_n5251) & (!n_n5249) & (n_n5252)) + ((n_n5258) & (!n_n5251) & (n_n5249) & (!n_n5252)) + ((n_n5258) & (!n_n5251) & (n_n5249) & (n_n5252)) + ((n_n5258) & (n_n5251) & (!n_n5249) & (!n_n5252)) + ((n_n5258) & (n_n5251) & (!n_n5249) & (n_n5252)) + ((n_n5258) & (n_n5251) & (n_n5249) & (!n_n5252)) + ((n_n5258) & (n_n5251) & (n_n5249) & (n_n5252)));
	assign x16279x = (((!n_n5247) & (!n_n5261) & (!n_n5260) & (!n_n5250) & (n_n5259)) + ((!n_n5247) & (!n_n5261) & (!n_n5260) & (n_n5250) & (!n_n5259)) + ((!n_n5247) & (!n_n5261) & (!n_n5260) & (n_n5250) & (n_n5259)) + ((!n_n5247) & (!n_n5261) & (n_n5260) & (!n_n5250) & (!n_n5259)) + ((!n_n5247) & (!n_n5261) & (n_n5260) & (!n_n5250) & (n_n5259)) + ((!n_n5247) & (!n_n5261) & (n_n5260) & (n_n5250) & (!n_n5259)) + ((!n_n5247) & (!n_n5261) & (n_n5260) & (n_n5250) & (n_n5259)) + ((!n_n5247) & (n_n5261) & (!n_n5260) & (!n_n5250) & (!n_n5259)) + ((!n_n5247) & (n_n5261) & (!n_n5260) & (!n_n5250) & (n_n5259)) + ((!n_n5247) & (n_n5261) & (!n_n5260) & (n_n5250) & (!n_n5259)) + ((!n_n5247) & (n_n5261) & (!n_n5260) & (n_n5250) & (n_n5259)) + ((!n_n5247) & (n_n5261) & (n_n5260) & (!n_n5250) & (!n_n5259)) + ((!n_n5247) & (n_n5261) & (n_n5260) & (!n_n5250) & (n_n5259)) + ((!n_n5247) & (n_n5261) & (n_n5260) & (n_n5250) & (!n_n5259)) + ((!n_n5247) & (n_n5261) & (n_n5260) & (n_n5250) & (n_n5259)) + ((n_n5247) & (!n_n5261) & (!n_n5260) & (!n_n5250) & (!n_n5259)) + ((n_n5247) & (!n_n5261) & (!n_n5260) & (!n_n5250) & (n_n5259)) + ((n_n5247) & (!n_n5261) & (!n_n5260) & (n_n5250) & (!n_n5259)) + ((n_n5247) & (!n_n5261) & (!n_n5260) & (n_n5250) & (n_n5259)) + ((n_n5247) & (!n_n5261) & (n_n5260) & (!n_n5250) & (!n_n5259)) + ((n_n5247) & (!n_n5261) & (n_n5260) & (!n_n5250) & (n_n5259)) + ((n_n5247) & (!n_n5261) & (n_n5260) & (n_n5250) & (!n_n5259)) + ((n_n5247) & (!n_n5261) & (n_n5260) & (n_n5250) & (n_n5259)) + ((n_n5247) & (n_n5261) & (!n_n5260) & (!n_n5250) & (!n_n5259)) + ((n_n5247) & (n_n5261) & (!n_n5260) & (!n_n5250) & (n_n5259)) + ((n_n5247) & (n_n5261) & (!n_n5260) & (n_n5250) & (!n_n5259)) + ((n_n5247) & (n_n5261) & (!n_n5260) & (n_n5250) & (n_n5259)) + ((n_n5247) & (n_n5261) & (n_n5260) & (!n_n5250) & (!n_n5259)) + ((n_n5247) & (n_n5261) & (n_n5260) & (!n_n5250) & (n_n5259)) + ((n_n5247) & (n_n5261) & (n_n5260) & (n_n5250) & (!n_n5259)) + ((n_n5247) & (n_n5261) & (n_n5260) & (n_n5250) & (n_n5259)));
	assign x14494x = (((!i_9_) & (n_n536) & (!n_n524) & (n_n473) & (n_n530)) + ((!i_9_) & (n_n536) & (n_n524) & (n_n473) & (n_n530)) + ((i_9_) & (n_n536) & (!n_n524) & (n_n473) & (n_n530)) + ((i_9_) & (n_n536) & (n_n524) & (n_n473) & (!n_n530)) + ((i_9_) & (n_n536) & (n_n524) & (n_n473) & (n_n530)));
	assign x22108x = (((!n_n4420) & (!n_n4419) & (!n_n4421) & (!n_n4417)));
	assign x14712x = (((!x21x) & (n_n482) & (!n_n473) & (n_n325) & (x23x)) + ((!x21x) & (n_n482) & (n_n473) & (n_n325) & (x23x)) + ((x21x) & (!n_n482) & (n_n473) & (n_n325) & (!x23x)) + ((x21x) & (!n_n482) & (n_n473) & (n_n325) & (x23x)) + ((x21x) & (n_n482) & (!n_n473) & (n_n325) & (x23x)) + ((x21x) & (n_n482) & (n_n473) & (n_n325) & (!x23x)) + ((x21x) & (n_n482) & (n_n473) & (n_n325) & (x23x)));
	assign x14629x = (((!n_n5191) & (!n_n4129) & (!n_n5188) & (!n_n1532) & (n_n3037)) + ((!n_n5191) & (!n_n4129) & (!n_n5188) & (n_n1532) & (!n_n3037)) + ((!n_n5191) & (!n_n4129) & (!n_n5188) & (n_n1532) & (n_n3037)) + ((!n_n5191) & (!n_n4129) & (n_n5188) & (!n_n1532) & (!n_n3037)) + ((!n_n5191) & (!n_n4129) & (n_n5188) & (!n_n1532) & (n_n3037)) + ((!n_n5191) & (!n_n4129) & (n_n5188) & (n_n1532) & (!n_n3037)) + ((!n_n5191) & (!n_n4129) & (n_n5188) & (n_n1532) & (n_n3037)) + ((!n_n5191) & (n_n4129) & (!n_n5188) & (!n_n1532) & (!n_n3037)) + ((!n_n5191) & (n_n4129) & (!n_n5188) & (!n_n1532) & (n_n3037)) + ((!n_n5191) & (n_n4129) & (!n_n5188) & (n_n1532) & (!n_n3037)) + ((!n_n5191) & (n_n4129) & (!n_n5188) & (n_n1532) & (n_n3037)) + ((!n_n5191) & (n_n4129) & (n_n5188) & (!n_n1532) & (!n_n3037)) + ((!n_n5191) & (n_n4129) & (n_n5188) & (!n_n1532) & (n_n3037)) + ((!n_n5191) & (n_n4129) & (n_n5188) & (n_n1532) & (!n_n3037)) + ((!n_n5191) & (n_n4129) & (n_n5188) & (n_n1532) & (n_n3037)) + ((n_n5191) & (!n_n4129) & (!n_n5188) & (!n_n1532) & (!n_n3037)) + ((n_n5191) & (!n_n4129) & (!n_n5188) & (!n_n1532) & (n_n3037)) + ((n_n5191) & (!n_n4129) & (!n_n5188) & (n_n1532) & (!n_n3037)) + ((n_n5191) & (!n_n4129) & (!n_n5188) & (n_n1532) & (n_n3037)) + ((n_n5191) & (!n_n4129) & (n_n5188) & (!n_n1532) & (!n_n3037)) + ((n_n5191) & (!n_n4129) & (n_n5188) & (!n_n1532) & (n_n3037)) + ((n_n5191) & (!n_n4129) & (n_n5188) & (n_n1532) & (!n_n3037)) + ((n_n5191) & (!n_n4129) & (n_n5188) & (n_n1532) & (n_n3037)) + ((n_n5191) & (n_n4129) & (!n_n5188) & (!n_n1532) & (!n_n3037)) + ((n_n5191) & (n_n4129) & (!n_n5188) & (!n_n1532) & (n_n3037)) + ((n_n5191) & (n_n4129) & (!n_n5188) & (n_n1532) & (!n_n3037)) + ((n_n5191) & (n_n4129) & (!n_n5188) & (n_n1532) & (n_n3037)) + ((n_n5191) & (n_n4129) & (n_n5188) & (!n_n1532) & (!n_n3037)) + ((n_n5191) & (n_n4129) & (n_n5188) & (!n_n1532) & (n_n3037)) + ((n_n5191) & (n_n4129) & (n_n5188) & (n_n1532) & (!n_n3037)) + ((n_n5191) & (n_n4129) & (n_n5188) & (n_n1532) & (n_n3037)));
	assign x14625x = (((!n_n5185) & (!n_n5183) & (!n_n5206) & (n_n5204)) + ((!n_n5185) & (!n_n5183) & (n_n5206) & (!n_n5204)) + ((!n_n5185) & (!n_n5183) & (n_n5206) & (n_n5204)) + ((!n_n5185) & (n_n5183) & (!n_n5206) & (!n_n5204)) + ((!n_n5185) & (n_n5183) & (!n_n5206) & (n_n5204)) + ((!n_n5185) & (n_n5183) & (n_n5206) & (!n_n5204)) + ((!n_n5185) & (n_n5183) & (n_n5206) & (n_n5204)) + ((n_n5185) & (!n_n5183) & (!n_n5206) & (!n_n5204)) + ((n_n5185) & (!n_n5183) & (!n_n5206) & (n_n5204)) + ((n_n5185) & (!n_n5183) & (n_n5206) & (!n_n5204)) + ((n_n5185) & (!n_n5183) & (n_n5206) & (n_n5204)) + ((n_n5185) & (n_n5183) & (!n_n5206) & (!n_n5204)) + ((n_n5185) & (n_n5183) & (!n_n5206) & (n_n5204)) + ((n_n5185) & (n_n5183) & (n_n5206) & (!n_n5204)) + ((n_n5185) & (n_n5183) & (n_n5206) & (n_n5204)));
	assign x14670x = (((!i_9_) & (!n_n526) & (n_n534) & (n_n195) & (n_n500)) + ((!i_9_) & (n_n526) & (n_n534) & (n_n195) & (n_n500)) + ((i_9_) & (!n_n526) & (n_n534) & (n_n195) & (n_n500)) + ((i_9_) & (n_n526) & (!n_n534) & (n_n195) & (n_n500)) + ((i_9_) & (n_n526) & (n_n534) & (n_n195) & (n_n500)));
	assign x14748x = (((!n_n4924) & (!n_n4947) & (!n_n4912) & (n_n4918)) + ((!n_n4924) & (!n_n4947) & (n_n4912) & (!n_n4918)) + ((!n_n4924) & (!n_n4947) & (n_n4912) & (n_n4918)) + ((!n_n4924) & (n_n4947) & (!n_n4912) & (!n_n4918)) + ((!n_n4924) & (n_n4947) & (!n_n4912) & (n_n4918)) + ((!n_n4924) & (n_n4947) & (n_n4912) & (!n_n4918)) + ((!n_n4924) & (n_n4947) & (n_n4912) & (n_n4918)) + ((n_n4924) & (!n_n4947) & (!n_n4912) & (!n_n4918)) + ((n_n4924) & (!n_n4947) & (!n_n4912) & (n_n4918)) + ((n_n4924) & (!n_n4947) & (n_n4912) & (!n_n4918)) + ((n_n4924) & (!n_n4947) & (n_n4912) & (n_n4918)) + ((n_n4924) & (n_n4947) & (!n_n4912) & (!n_n4918)) + ((n_n4924) & (n_n4947) & (!n_n4912) & (n_n4918)) + ((n_n4924) & (n_n4947) & (n_n4912) & (!n_n4918)) + ((n_n4924) & (n_n4947) & (n_n4912) & (n_n4918)));
	assign x14749x = (((!n_n4920) & (!n_n4914) & (!n_n4919) & (!n_n4917) & (x42x)) + ((!n_n4920) & (!n_n4914) & (!n_n4919) & (n_n4917) & (!x42x)) + ((!n_n4920) & (!n_n4914) & (!n_n4919) & (n_n4917) & (x42x)) + ((!n_n4920) & (!n_n4914) & (n_n4919) & (!n_n4917) & (!x42x)) + ((!n_n4920) & (!n_n4914) & (n_n4919) & (!n_n4917) & (x42x)) + ((!n_n4920) & (!n_n4914) & (n_n4919) & (n_n4917) & (!x42x)) + ((!n_n4920) & (!n_n4914) & (n_n4919) & (n_n4917) & (x42x)) + ((!n_n4920) & (n_n4914) & (!n_n4919) & (!n_n4917) & (!x42x)) + ((!n_n4920) & (n_n4914) & (!n_n4919) & (!n_n4917) & (x42x)) + ((!n_n4920) & (n_n4914) & (!n_n4919) & (n_n4917) & (!x42x)) + ((!n_n4920) & (n_n4914) & (!n_n4919) & (n_n4917) & (x42x)) + ((!n_n4920) & (n_n4914) & (n_n4919) & (!n_n4917) & (!x42x)) + ((!n_n4920) & (n_n4914) & (n_n4919) & (!n_n4917) & (x42x)) + ((!n_n4920) & (n_n4914) & (n_n4919) & (n_n4917) & (!x42x)) + ((!n_n4920) & (n_n4914) & (n_n4919) & (n_n4917) & (x42x)) + ((n_n4920) & (!n_n4914) & (!n_n4919) & (!n_n4917) & (!x42x)) + ((n_n4920) & (!n_n4914) & (!n_n4919) & (!n_n4917) & (x42x)) + ((n_n4920) & (!n_n4914) & (!n_n4919) & (n_n4917) & (!x42x)) + ((n_n4920) & (!n_n4914) & (!n_n4919) & (n_n4917) & (x42x)) + ((n_n4920) & (!n_n4914) & (n_n4919) & (!n_n4917) & (!x42x)) + ((n_n4920) & (!n_n4914) & (n_n4919) & (!n_n4917) & (x42x)) + ((n_n4920) & (!n_n4914) & (n_n4919) & (n_n4917) & (!x42x)) + ((n_n4920) & (!n_n4914) & (n_n4919) & (n_n4917) & (x42x)) + ((n_n4920) & (n_n4914) & (!n_n4919) & (!n_n4917) & (!x42x)) + ((n_n4920) & (n_n4914) & (!n_n4919) & (!n_n4917) & (x42x)) + ((n_n4920) & (n_n4914) & (!n_n4919) & (n_n4917) & (!x42x)) + ((n_n4920) & (n_n4914) & (!n_n4919) & (n_n4917) & (x42x)) + ((n_n4920) & (n_n4914) & (n_n4919) & (!n_n4917) & (!x42x)) + ((n_n4920) & (n_n4914) & (n_n4919) & (!n_n4917) & (x42x)) + ((n_n4920) & (n_n4914) & (n_n4919) & (n_n4917) & (!x42x)) + ((n_n4920) & (n_n4914) & (n_n4919) & (n_n4917) & (x42x)));
	assign x14764x = (((!n_n4980) & (!n_n4985) & (!n_n4986) & (!n_n4978) & (x229x)) + ((!n_n4980) & (!n_n4985) & (!n_n4986) & (n_n4978) & (!x229x)) + ((!n_n4980) & (!n_n4985) & (!n_n4986) & (n_n4978) & (x229x)) + ((!n_n4980) & (!n_n4985) & (n_n4986) & (!n_n4978) & (!x229x)) + ((!n_n4980) & (!n_n4985) & (n_n4986) & (!n_n4978) & (x229x)) + ((!n_n4980) & (!n_n4985) & (n_n4986) & (n_n4978) & (!x229x)) + ((!n_n4980) & (!n_n4985) & (n_n4986) & (n_n4978) & (x229x)) + ((!n_n4980) & (n_n4985) & (!n_n4986) & (!n_n4978) & (!x229x)) + ((!n_n4980) & (n_n4985) & (!n_n4986) & (!n_n4978) & (x229x)) + ((!n_n4980) & (n_n4985) & (!n_n4986) & (n_n4978) & (!x229x)) + ((!n_n4980) & (n_n4985) & (!n_n4986) & (n_n4978) & (x229x)) + ((!n_n4980) & (n_n4985) & (n_n4986) & (!n_n4978) & (!x229x)) + ((!n_n4980) & (n_n4985) & (n_n4986) & (!n_n4978) & (x229x)) + ((!n_n4980) & (n_n4985) & (n_n4986) & (n_n4978) & (!x229x)) + ((!n_n4980) & (n_n4985) & (n_n4986) & (n_n4978) & (x229x)) + ((n_n4980) & (!n_n4985) & (!n_n4986) & (!n_n4978) & (!x229x)) + ((n_n4980) & (!n_n4985) & (!n_n4986) & (!n_n4978) & (x229x)) + ((n_n4980) & (!n_n4985) & (!n_n4986) & (n_n4978) & (!x229x)) + ((n_n4980) & (!n_n4985) & (!n_n4986) & (n_n4978) & (x229x)) + ((n_n4980) & (!n_n4985) & (n_n4986) & (!n_n4978) & (!x229x)) + ((n_n4980) & (!n_n4985) & (n_n4986) & (!n_n4978) & (x229x)) + ((n_n4980) & (!n_n4985) & (n_n4986) & (n_n4978) & (!x229x)) + ((n_n4980) & (!n_n4985) & (n_n4986) & (n_n4978) & (x229x)) + ((n_n4980) & (n_n4985) & (!n_n4986) & (!n_n4978) & (!x229x)) + ((n_n4980) & (n_n4985) & (!n_n4986) & (!n_n4978) & (x229x)) + ((n_n4980) & (n_n4985) & (!n_n4986) & (n_n4978) & (!x229x)) + ((n_n4980) & (n_n4985) & (!n_n4986) & (n_n4978) & (x229x)) + ((n_n4980) & (n_n4985) & (n_n4986) & (!n_n4978) & (!x229x)) + ((n_n4980) & (n_n4985) & (n_n4986) & (!n_n4978) & (x229x)) + ((n_n4980) & (n_n4985) & (n_n4986) & (n_n4978) & (!x229x)) + ((n_n4980) & (n_n4985) & (n_n4986) & (n_n4978) & (x229x)));
	assign x14763x = (((!n_n4983) & (!n_n4984) & (!n_n4972) & (x14761x)) + ((!n_n4983) & (!n_n4984) & (n_n4972) & (!x14761x)) + ((!n_n4983) & (!n_n4984) & (n_n4972) & (x14761x)) + ((!n_n4983) & (n_n4984) & (!n_n4972) & (!x14761x)) + ((!n_n4983) & (n_n4984) & (!n_n4972) & (x14761x)) + ((!n_n4983) & (n_n4984) & (n_n4972) & (!x14761x)) + ((!n_n4983) & (n_n4984) & (n_n4972) & (x14761x)) + ((n_n4983) & (!n_n4984) & (!n_n4972) & (!x14761x)) + ((n_n4983) & (!n_n4984) & (!n_n4972) & (x14761x)) + ((n_n4983) & (!n_n4984) & (n_n4972) & (!x14761x)) + ((n_n4983) & (!n_n4984) & (n_n4972) & (x14761x)) + ((n_n4983) & (n_n4984) & (!n_n4972) & (!x14761x)) + ((n_n4983) & (n_n4984) & (!n_n4972) & (x14761x)) + ((n_n4983) & (n_n4984) & (n_n4972) & (!x14761x)) + ((n_n4983) & (n_n4984) & (n_n4972) & (x14761x)));
	assign x15740x = (((!n_n4905) & (!n_n4918) & (!x305x) & (!x15735x) & (x15737x)) + ((!n_n4905) & (!n_n4918) & (!x305x) & (x15735x) & (!x15737x)) + ((!n_n4905) & (!n_n4918) & (!x305x) & (x15735x) & (x15737x)) + ((!n_n4905) & (!n_n4918) & (x305x) & (!x15735x) & (!x15737x)) + ((!n_n4905) & (!n_n4918) & (x305x) & (!x15735x) & (x15737x)) + ((!n_n4905) & (!n_n4918) & (x305x) & (x15735x) & (!x15737x)) + ((!n_n4905) & (!n_n4918) & (x305x) & (x15735x) & (x15737x)) + ((!n_n4905) & (n_n4918) & (!x305x) & (!x15735x) & (!x15737x)) + ((!n_n4905) & (n_n4918) & (!x305x) & (!x15735x) & (x15737x)) + ((!n_n4905) & (n_n4918) & (!x305x) & (x15735x) & (!x15737x)) + ((!n_n4905) & (n_n4918) & (!x305x) & (x15735x) & (x15737x)) + ((!n_n4905) & (n_n4918) & (x305x) & (!x15735x) & (!x15737x)) + ((!n_n4905) & (n_n4918) & (x305x) & (!x15735x) & (x15737x)) + ((!n_n4905) & (n_n4918) & (x305x) & (x15735x) & (!x15737x)) + ((!n_n4905) & (n_n4918) & (x305x) & (x15735x) & (x15737x)) + ((n_n4905) & (!n_n4918) & (!x305x) & (!x15735x) & (!x15737x)) + ((n_n4905) & (!n_n4918) & (!x305x) & (!x15735x) & (x15737x)) + ((n_n4905) & (!n_n4918) & (!x305x) & (x15735x) & (!x15737x)) + ((n_n4905) & (!n_n4918) & (!x305x) & (x15735x) & (x15737x)) + ((n_n4905) & (!n_n4918) & (x305x) & (!x15735x) & (!x15737x)) + ((n_n4905) & (!n_n4918) & (x305x) & (!x15735x) & (x15737x)) + ((n_n4905) & (!n_n4918) & (x305x) & (x15735x) & (!x15737x)) + ((n_n4905) & (!n_n4918) & (x305x) & (x15735x) & (x15737x)) + ((n_n4905) & (n_n4918) & (!x305x) & (!x15735x) & (!x15737x)) + ((n_n4905) & (n_n4918) & (!x305x) & (!x15735x) & (x15737x)) + ((n_n4905) & (n_n4918) & (!x305x) & (x15735x) & (!x15737x)) + ((n_n4905) & (n_n4918) & (!x305x) & (x15735x) & (x15737x)) + ((n_n4905) & (n_n4918) & (x305x) & (!x15735x) & (!x15737x)) + ((n_n4905) & (n_n4918) & (x305x) & (!x15735x) & (x15737x)) + ((n_n4905) & (n_n4918) & (x305x) & (x15735x) & (!x15737x)) + ((n_n4905) & (n_n4918) & (x305x) & (x15735x) & (x15737x)));
	assign x15783x = (((!n_n4749) & (!n_n4748) & (!n_n4747) & (!n_n4743) & (n_n4742)) + ((!n_n4749) & (!n_n4748) & (!n_n4747) & (n_n4743) & (!n_n4742)) + ((!n_n4749) & (!n_n4748) & (!n_n4747) & (n_n4743) & (n_n4742)) + ((!n_n4749) & (!n_n4748) & (n_n4747) & (!n_n4743) & (!n_n4742)) + ((!n_n4749) & (!n_n4748) & (n_n4747) & (!n_n4743) & (n_n4742)) + ((!n_n4749) & (!n_n4748) & (n_n4747) & (n_n4743) & (!n_n4742)) + ((!n_n4749) & (!n_n4748) & (n_n4747) & (n_n4743) & (n_n4742)) + ((!n_n4749) & (n_n4748) & (!n_n4747) & (!n_n4743) & (!n_n4742)) + ((!n_n4749) & (n_n4748) & (!n_n4747) & (!n_n4743) & (n_n4742)) + ((!n_n4749) & (n_n4748) & (!n_n4747) & (n_n4743) & (!n_n4742)) + ((!n_n4749) & (n_n4748) & (!n_n4747) & (n_n4743) & (n_n4742)) + ((!n_n4749) & (n_n4748) & (n_n4747) & (!n_n4743) & (!n_n4742)) + ((!n_n4749) & (n_n4748) & (n_n4747) & (!n_n4743) & (n_n4742)) + ((!n_n4749) & (n_n4748) & (n_n4747) & (n_n4743) & (!n_n4742)) + ((!n_n4749) & (n_n4748) & (n_n4747) & (n_n4743) & (n_n4742)) + ((n_n4749) & (!n_n4748) & (!n_n4747) & (!n_n4743) & (!n_n4742)) + ((n_n4749) & (!n_n4748) & (!n_n4747) & (!n_n4743) & (n_n4742)) + ((n_n4749) & (!n_n4748) & (!n_n4747) & (n_n4743) & (!n_n4742)) + ((n_n4749) & (!n_n4748) & (!n_n4747) & (n_n4743) & (n_n4742)) + ((n_n4749) & (!n_n4748) & (n_n4747) & (!n_n4743) & (!n_n4742)) + ((n_n4749) & (!n_n4748) & (n_n4747) & (!n_n4743) & (n_n4742)) + ((n_n4749) & (!n_n4748) & (n_n4747) & (n_n4743) & (!n_n4742)) + ((n_n4749) & (!n_n4748) & (n_n4747) & (n_n4743) & (n_n4742)) + ((n_n4749) & (n_n4748) & (!n_n4747) & (!n_n4743) & (!n_n4742)) + ((n_n4749) & (n_n4748) & (!n_n4747) & (!n_n4743) & (n_n4742)) + ((n_n4749) & (n_n4748) & (!n_n4747) & (n_n4743) & (!n_n4742)) + ((n_n4749) & (n_n4748) & (!n_n4747) & (n_n4743) & (n_n4742)) + ((n_n4749) & (n_n4748) & (n_n4747) & (!n_n4743) & (!n_n4742)) + ((n_n4749) & (n_n4748) & (n_n4747) & (!n_n4743) & (n_n4742)) + ((n_n4749) & (n_n4748) & (n_n4747) & (n_n4743) & (!n_n4742)) + ((n_n4749) & (n_n4748) & (n_n4747) & (n_n4743) & (n_n4742)));
	assign x15786x = (((!n_n2981) & (!x374x) & (!x47x) & (!n_n2982) & (x15783x)) + ((!n_n2981) & (!x374x) & (!x47x) & (n_n2982) & (!x15783x)) + ((!n_n2981) & (!x374x) & (!x47x) & (n_n2982) & (x15783x)) + ((!n_n2981) & (!x374x) & (x47x) & (!n_n2982) & (!x15783x)) + ((!n_n2981) & (!x374x) & (x47x) & (!n_n2982) & (x15783x)) + ((!n_n2981) & (!x374x) & (x47x) & (n_n2982) & (!x15783x)) + ((!n_n2981) & (!x374x) & (x47x) & (n_n2982) & (x15783x)) + ((!n_n2981) & (x374x) & (!x47x) & (!n_n2982) & (!x15783x)) + ((!n_n2981) & (x374x) & (!x47x) & (!n_n2982) & (x15783x)) + ((!n_n2981) & (x374x) & (!x47x) & (n_n2982) & (!x15783x)) + ((!n_n2981) & (x374x) & (!x47x) & (n_n2982) & (x15783x)) + ((!n_n2981) & (x374x) & (x47x) & (!n_n2982) & (!x15783x)) + ((!n_n2981) & (x374x) & (x47x) & (!n_n2982) & (x15783x)) + ((!n_n2981) & (x374x) & (x47x) & (n_n2982) & (!x15783x)) + ((!n_n2981) & (x374x) & (x47x) & (n_n2982) & (x15783x)) + ((n_n2981) & (!x374x) & (!x47x) & (!n_n2982) & (!x15783x)) + ((n_n2981) & (!x374x) & (!x47x) & (!n_n2982) & (x15783x)) + ((n_n2981) & (!x374x) & (!x47x) & (n_n2982) & (!x15783x)) + ((n_n2981) & (!x374x) & (!x47x) & (n_n2982) & (x15783x)) + ((n_n2981) & (!x374x) & (x47x) & (!n_n2982) & (!x15783x)) + ((n_n2981) & (!x374x) & (x47x) & (!n_n2982) & (x15783x)) + ((n_n2981) & (!x374x) & (x47x) & (n_n2982) & (!x15783x)) + ((n_n2981) & (!x374x) & (x47x) & (n_n2982) & (x15783x)) + ((n_n2981) & (x374x) & (!x47x) & (!n_n2982) & (!x15783x)) + ((n_n2981) & (x374x) & (!x47x) & (!n_n2982) & (x15783x)) + ((n_n2981) & (x374x) & (!x47x) & (n_n2982) & (!x15783x)) + ((n_n2981) & (x374x) & (!x47x) & (n_n2982) & (x15783x)) + ((n_n2981) & (x374x) & (x47x) & (!n_n2982) & (!x15783x)) + ((n_n2981) & (x374x) & (x47x) & (!n_n2982) & (x15783x)) + ((n_n2981) & (x374x) & (x47x) & (n_n2982) & (!x15783x)) + ((n_n2981) & (x374x) & (x47x) & (n_n2982) & (x15783x)));
	assign x15798x = (((!n_n4806) & (!n_n4805) & (!n_n4197) & (x390x)) + ((!n_n4806) & (!n_n4805) & (n_n4197) & (!x390x)) + ((!n_n4806) & (!n_n4805) & (n_n4197) & (x390x)) + ((!n_n4806) & (n_n4805) & (!n_n4197) & (!x390x)) + ((!n_n4806) & (n_n4805) & (!n_n4197) & (x390x)) + ((!n_n4806) & (n_n4805) & (n_n4197) & (!x390x)) + ((!n_n4806) & (n_n4805) & (n_n4197) & (x390x)) + ((n_n4806) & (!n_n4805) & (!n_n4197) & (!x390x)) + ((n_n4806) & (!n_n4805) & (!n_n4197) & (x390x)) + ((n_n4806) & (!n_n4805) & (n_n4197) & (!x390x)) + ((n_n4806) & (!n_n4805) & (n_n4197) & (x390x)) + ((n_n4806) & (n_n4805) & (!n_n4197) & (!x390x)) + ((n_n4806) & (n_n4805) & (!n_n4197) & (x390x)) + ((n_n4806) & (n_n4805) & (n_n4197) & (!x390x)) + ((n_n4806) & (n_n4805) & (n_n4197) & (x390x)));
	assign x15797x = (((!n_n4816) & (!n_n4800) & (!x71x) & (!x440x) & (x381x)) + ((!n_n4816) & (!n_n4800) & (!x71x) & (x440x) & (!x381x)) + ((!n_n4816) & (!n_n4800) & (!x71x) & (x440x) & (x381x)) + ((!n_n4816) & (!n_n4800) & (x71x) & (!x440x) & (!x381x)) + ((!n_n4816) & (!n_n4800) & (x71x) & (!x440x) & (x381x)) + ((!n_n4816) & (!n_n4800) & (x71x) & (x440x) & (!x381x)) + ((!n_n4816) & (!n_n4800) & (x71x) & (x440x) & (x381x)) + ((!n_n4816) & (n_n4800) & (!x71x) & (!x440x) & (!x381x)) + ((!n_n4816) & (n_n4800) & (!x71x) & (!x440x) & (x381x)) + ((!n_n4816) & (n_n4800) & (!x71x) & (x440x) & (!x381x)) + ((!n_n4816) & (n_n4800) & (!x71x) & (x440x) & (x381x)) + ((!n_n4816) & (n_n4800) & (x71x) & (!x440x) & (!x381x)) + ((!n_n4816) & (n_n4800) & (x71x) & (!x440x) & (x381x)) + ((!n_n4816) & (n_n4800) & (x71x) & (x440x) & (!x381x)) + ((!n_n4816) & (n_n4800) & (x71x) & (x440x) & (x381x)) + ((n_n4816) & (!n_n4800) & (!x71x) & (!x440x) & (!x381x)) + ((n_n4816) & (!n_n4800) & (!x71x) & (!x440x) & (x381x)) + ((n_n4816) & (!n_n4800) & (!x71x) & (x440x) & (!x381x)) + ((n_n4816) & (!n_n4800) & (!x71x) & (x440x) & (x381x)) + ((n_n4816) & (!n_n4800) & (x71x) & (!x440x) & (!x381x)) + ((n_n4816) & (!n_n4800) & (x71x) & (!x440x) & (x381x)) + ((n_n4816) & (!n_n4800) & (x71x) & (x440x) & (!x381x)) + ((n_n4816) & (!n_n4800) & (x71x) & (x440x) & (x381x)) + ((n_n4816) & (n_n4800) & (!x71x) & (!x440x) & (!x381x)) + ((n_n4816) & (n_n4800) & (!x71x) & (!x440x) & (x381x)) + ((n_n4816) & (n_n4800) & (!x71x) & (x440x) & (!x381x)) + ((n_n4816) & (n_n4800) & (!x71x) & (x440x) & (x381x)) + ((n_n4816) & (n_n4800) & (x71x) & (!x440x) & (!x381x)) + ((n_n4816) & (n_n4800) & (x71x) & (!x440x) & (x381x)) + ((n_n4816) & (n_n4800) & (x71x) & (x440x) & (!x381x)) + ((n_n4816) & (n_n4800) & (x71x) & (x440x) & (x381x)));
	assign x16002x = (((!x20x) & (!x233x) & (!n_n4436) & (n_n4447) & (!x496x)) + ((!x20x) & (!x233x) & (!n_n4436) & (n_n4447) & (x496x)) + ((!x20x) & (!x233x) & (n_n4436) & (!n_n4447) & (!x496x)) + ((!x20x) & (!x233x) & (n_n4436) & (!n_n4447) & (x496x)) + ((!x20x) & (!x233x) & (n_n4436) & (n_n4447) & (!x496x)) + ((!x20x) & (!x233x) & (n_n4436) & (n_n4447) & (x496x)) + ((!x20x) & (x233x) & (!n_n4436) & (!n_n4447) & (!x496x)) + ((!x20x) & (x233x) & (!n_n4436) & (!n_n4447) & (x496x)) + ((!x20x) & (x233x) & (!n_n4436) & (n_n4447) & (!x496x)) + ((!x20x) & (x233x) & (!n_n4436) & (n_n4447) & (x496x)) + ((!x20x) & (x233x) & (n_n4436) & (!n_n4447) & (!x496x)) + ((!x20x) & (x233x) & (n_n4436) & (!n_n4447) & (x496x)) + ((!x20x) & (x233x) & (n_n4436) & (n_n4447) & (!x496x)) + ((!x20x) & (x233x) & (n_n4436) & (n_n4447) & (x496x)) + ((x20x) & (!x233x) & (!n_n4436) & (!n_n4447) & (x496x)) + ((x20x) & (!x233x) & (!n_n4436) & (n_n4447) & (!x496x)) + ((x20x) & (!x233x) & (!n_n4436) & (n_n4447) & (x496x)) + ((x20x) & (!x233x) & (n_n4436) & (!n_n4447) & (!x496x)) + ((x20x) & (!x233x) & (n_n4436) & (!n_n4447) & (x496x)) + ((x20x) & (!x233x) & (n_n4436) & (n_n4447) & (!x496x)) + ((x20x) & (!x233x) & (n_n4436) & (n_n4447) & (x496x)) + ((x20x) & (x233x) & (!n_n4436) & (!n_n4447) & (!x496x)) + ((x20x) & (x233x) & (!n_n4436) & (!n_n4447) & (x496x)) + ((x20x) & (x233x) & (!n_n4436) & (n_n4447) & (!x496x)) + ((x20x) & (x233x) & (!n_n4436) & (n_n4447) & (x496x)) + ((x20x) & (x233x) & (n_n4436) & (!n_n4447) & (!x496x)) + ((x20x) & (x233x) & (n_n4436) & (!n_n4447) & (x496x)) + ((x20x) & (x233x) & (n_n4436) & (n_n4447) & (!x496x)) + ((x20x) & (x233x) & (n_n4436) & (n_n4447) & (x496x)));
	assign x14604x = (((!n_n524) & (!n_n509) & (!x12x) & (!n_n5123) & (n_n5125)) + ((!n_n524) & (!n_n509) & (!x12x) & (n_n5123) & (!n_n5125)) + ((!n_n524) & (!n_n509) & (!x12x) & (n_n5123) & (n_n5125)) + ((!n_n524) & (!n_n509) & (x12x) & (!n_n5123) & (n_n5125)) + ((!n_n524) & (!n_n509) & (x12x) & (n_n5123) & (!n_n5125)) + ((!n_n524) & (!n_n509) & (x12x) & (n_n5123) & (n_n5125)) + ((!n_n524) & (n_n509) & (!x12x) & (!n_n5123) & (n_n5125)) + ((!n_n524) & (n_n509) & (!x12x) & (n_n5123) & (!n_n5125)) + ((!n_n524) & (n_n509) & (!x12x) & (n_n5123) & (n_n5125)) + ((!n_n524) & (n_n509) & (x12x) & (!n_n5123) & (n_n5125)) + ((!n_n524) & (n_n509) & (x12x) & (n_n5123) & (!n_n5125)) + ((!n_n524) & (n_n509) & (x12x) & (n_n5123) & (n_n5125)) + ((n_n524) & (!n_n509) & (!x12x) & (!n_n5123) & (n_n5125)) + ((n_n524) & (!n_n509) & (!x12x) & (n_n5123) & (!n_n5125)) + ((n_n524) & (!n_n509) & (!x12x) & (n_n5123) & (n_n5125)) + ((n_n524) & (!n_n509) & (x12x) & (!n_n5123) & (n_n5125)) + ((n_n524) & (!n_n509) & (x12x) & (n_n5123) & (!n_n5125)) + ((n_n524) & (!n_n509) & (x12x) & (n_n5123) & (n_n5125)) + ((n_n524) & (n_n509) & (!x12x) & (!n_n5123) & (n_n5125)) + ((n_n524) & (n_n509) & (!x12x) & (n_n5123) & (!n_n5125)) + ((n_n524) & (n_n509) & (!x12x) & (n_n5123) & (n_n5125)) + ((n_n524) & (n_n509) & (x12x) & (!n_n5123) & (!n_n5125)) + ((n_n524) & (n_n509) & (x12x) & (!n_n5123) & (n_n5125)) + ((n_n524) & (n_n509) & (x12x) & (n_n5123) & (!n_n5125)) + ((n_n524) & (n_n509) & (x12x) & (n_n5123) & (n_n5125)));
	assign x22105x = (((!n_n5116) & (!n_n5120) & (!n_n5115) & (!n_n5118)));
	assign x22079x = (((!i_7_) & (!i_8_) & (!i_6_) & (!n_n482) & (!x10x)) + ((!i_7_) & (!i_8_) & (!i_6_) & (!n_n482) & (x10x)) + ((!i_7_) & (!i_8_) & (!i_6_) & (n_n482) & (!x10x)) + ((!i_7_) & (!i_8_) & (!i_6_) & (n_n482) & (x10x)) + ((!i_7_) & (!i_8_) & (i_6_) & (!n_n482) & (!x10x)) + ((!i_7_) & (!i_8_) & (i_6_) & (!n_n482) & (x10x)) + ((!i_7_) & (!i_8_) & (i_6_) & (n_n482) & (!x10x)) + ((!i_7_) & (i_8_) & (!i_6_) & (!n_n482) & (!x10x)) + ((!i_7_) & (i_8_) & (!i_6_) & (!n_n482) & (x10x)) + ((!i_7_) & (i_8_) & (!i_6_) & (n_n482) & (!x10x)) + ((!i_7_) & (i_8_) & (i_6_) & (!n_n482) & (!x10x)) + ((!i_7_) & (i_8_) & (i_6_) & (!n_n482) & (x10x)) + ((!i_7_) & (i_8_) & (i_6_) & (n_n482) & (!x10x)) + ((i_7_) & (!i_8_) & (!i_6_) & (!n_n482) & (!x10x)) + ((i_7_) & (!i_8_) & (!i_6_) & (!n_n482) & (x10x)) + ((i_7_) & (!i_8_) & (!i_6_) & (n_n482) & (!x10x)) + ((i_7_) & (!i_8_) & (!i_6_) & (n_n482) & (x10x)) + ((i_7_) & (!i_8_) & (i_6_) & (!n_n482) & (!x10x)) + ((i_7_) & (!i_8_) & (i_6_) & (!n_n482) & (x10x)) + ((i_7_) & (!i_8_) & (i_6_) & (n_n482) & (!x10x)) + ((i_7_) & (i_8_) & (!i_6_) & (!n_n482) & (!x10x)) + ((i_7_) & (i_8_) & (!i_6_) & (!n_n482) & (x10x)) + ((i_7_) & (i_8_) & (!i_6_) & (n_n482) & (!x10x)) + ((i_7_) & (i_8_) & (!i_6_) & (n_n482) & (x10x)) + ((i_7_) & (i_8_) & (i_6_) & (!n_n482) & (!x10x)) + ((i_7_) & (i_8_) & (i_6_) & (!n_n482) & (x10x)) + ((i_7_) & (i_8_) & (i_6_) & (n_n482) & (!x10x)) + ((i_7_) & (i_8_) & (i_6_) & (n_n482) & (x10x)));
	assign x617x = (((i_1_) & (!i_2_) & (i_0_) & (n_n509) & (x20x)));
	assign x11524x = (((n_n536) & (n_n473) & (!x20x) & (x23x)) + ((n_n536) & (n_n473) & (x20x) & (!x23x)) + ((n_n536) & (n_n473) & (x20x) & (x23x)));
	assign x11571x = (((!n_n4578) & (!n_n4582) & (!n_n4569) & (n_n4573)) + ((!n_n4578) & (!n_n4582) & (n_n4569) & (!n_n4573)) + ((!n_n4578) & (!n_n4582) & (n_n4569) & (n_n4573)) + ((!n_n4578) & (n_n4582) & (!n_n4569) & (!n_n4573)) + ((!n_n4578) & (n_n4582) & (!n_n4569) & (n_n4573)) + ((!n_n4578) & (n_n4582) & (n_n4569) & (!n_n4573)) + ((!n_n4578) & (n_n4582) & (n_n4569) & (n_n4573)) + ((n_n4578) & (!n_n4582) & (!n_n4569) & (!n_n4573)) + ((n_n4578) & (!n_n4582) & (!n_n4569) & (n_n4573)) + ((n_n4578) & (!n_n4582) & (n_n4569) & (!n_n4573)) + ((n_n4578) & (!n_n4582) & (n_n4569) & (n_n4573)) + ((n_n4578) & (n_n4582) & (!n_n4569) & (!n_n4573)) + ((n_n4578) & (n_n4582) & (!n_n4569) & (n_n4573)) + ((n_n4578) & (n_n4582) & (n_n4569) & (!n_n4573)) + ((n_n4578) & (n_n4582) & (n_n4569) & (n_n4573)));
	assign x11631x = (((!x198x) & (!n_n4328) & (!n_n4334) & (n_n4322)) + ((!x198x) & (!n_n4328) & (n_n4334) & (!n_n4322)) + ((!x198x) & (!n_n4328) & (n_n4334) & (n_n4322)) + ((!x198x) & (n_n4328) & (!n_n4334) & (!n_n4322)) + ((!x198x) & (n_n4328) & (!n_n4334) & (n_n4322)) + ((!x198x) & (n_n4328) & (n_n4334) & (!n_n4322)) + ((!x198x) & (n_n4328) & (n_n4334) & (n_n4322)) + ((x198x) & (!n_n4328) & (!n_n4334) & (!n_n4322)) + ((x198x) & (!n_n4328) & (!n_n4334) & (n_n4322)) + ((x198x) & (!n_n4328) & (n_n4334) & (!n_n4322)) + ((x198x) & (!n_n4328) & (n_n4334) & (n_n4322)) + ((x198x) & (n_n4328) & (!n_n4334) & (!n_n4322)) + ((x198x) & (n_n4328) & (!n_n4334) & (n_n4322)) + ((x198x) & (n_n4328) & (n_n4334) & (!n_n4322)) + ((x198x) & (n_n4328) & (n_n4334) & (n_n4322)));
	assign x11732x = (((!n_n5302) & (!n_n5289) & (!n_n5335) & (n_n5304)) + ((!n_n5302) & (!n_n5289) & (n_n5335) & (!n_n5304)) + ((!n_n5302) & (!n_n5289) & (n_n5335) & (n_n5304)) + ((!n_n5302) & (n_n5289) & (!n_n5335) & (!n_n5304)) + ((!n_n5302) & (n_n5289) & (!n_n5335) & (n_n5304)) + ((!n_n5302) & (n_n5289) & (n_n5335) & (!n_n5304)) + ((!n_n5302) & (n_n5289) & (n_n5335) & (n_n5304)) + ((n_n5302) & (!n_n5289) & (!n_n5335) & (!n_n5304)) + ((n_n5302) & (!n_n5289) & (!n_n5335) & (n_n5304)) + ((n_n5302) & (!n_n5289) & (n_n5335) & (!n_n5304)) + ((n_n5302) & (!n_n5289) & (n_n5335) & (n_n5304)) + ((n_n5302) & (n_n5289) & (!n_n5335) & (!n_n5304)) + ((n_n5302) & (n_n5289) & (!n_n5335) & (n_n5304)) + ((n_n5302) & (n_n5289) & (n_n5335) & (!n_n5304)) + ((n_n5302) & (n_n5289) & (n_n5335) & (n_n5304)));
	assign x22198x = (((!x19x) & (!x506x) & (!n_n5320) & (!n_n5307) & (!n_n5329)) + ((!x19x) & (x506x) & (!n_n5320) & (!n_n5307) & (!n_n5329)) + ((x19x) & (!x506x) & (!n_n5320) & (!n_n5307) & (!n_n5329)));
	assign x11742x = (((!n_n536) & (!x21x) & (!n_n535) & (!n_n4374) & (n_n1002)) + ((!n_n536) & (!x21x) & (!n_n535) & (n_n4374) & (!n_n1002)) + ((!n_n536) & (!x21x) & (!n_n535) & (n_n4374) & (n_n1002)) + ((!n_n536) & (!x21x) & (n_n535) & (!n_n4374) & (n_n1002)) + ((!n_n536) & (!x21x) & (n_n535) & (n_n4374) & (!n_n1002)) + ((!n_n536) & (!x21x) & (n_n535) & (n_n4374) & (n_n1002)) + ((!n_n536) & (x21x) & (!n_n535) & (!n_n4374) & (n_n1002)) + ((!n_n536) & (x21x) & (!n_n535) & (n_n4374) & (!n_n1002)) + ((!n_n536) & (x21x) & (!n_n535) & (n_n4374) & (n_n1002)) + ((!n_n536) & (x21x) & (n_n535) & (!n_n4374) & (n_n1002)) + ((!n_n536) & (x21x) & (n_n535) & (n_n4374) & (!n_n1002)) + ((!n_n536) & (x21x) & (n_n535) & (n_n4374) & (n_n1002)) + ((n_n536) & (!x21x) & (!n_n535) & (!n_n4374) & (n_n1002)) + ((n_n536) & (!x21x) & (!n_n535) & (n_n4374) & (!n_n1002)) + ((n_n536) & (!x21x) & (!n_n535) & (n_n4374) & (n_n1002)) + ((n_n536) & (!x21x) & (n_n535) & (!n_n4374) & (n_n1002)) + ((n_n536) & (!x21x) & (n_n535) & (n_n4374) & (!n_n1002)) + ((n_n536) & (!x21x) & (n_n535) & (n_n4374) & (n_n1002)) + ((n_n536) & (x21x) & (!n_n535) & (!n_n4374) & (n_n1002)) + ((n_n536) & (x21x) & (!n_n535) & (n_n4374) & (!n_n1002)) + ((n_n536) & (x21x) & (!n_n535) & (n_n4374) & (n_n1002)) + ((n_n536) & (x21x) & (n_n535) & (!n_n4374) & (!n_n1002)) + ((n_n536) & (x21x) & (n_n535) & (!n_n4374) & (n_n1002)) + ((n_n536) & (x21x) & (n_n535) & (n_n4374) & (!n_n1002)) + ((n_n536) & (x21x) & (n_n535) & (n_n4374) & (n_n1002)));
	assign x11743x = (((!n_n4324) & (!n_n4340) & (!n_n4384) & (!n_n4390) & (x11742x)) + ((!n_n4324) & (!n_n4340) & (!n_n4384) & (n_n4390) & (!x11742x)) + ((!n_n4324) & (!n_n4340) & (!n_n4384) & (n_n4390) & (x11742x)) + ((!n_n4324) & (!n_n4340) & (n_n4384) & (!n_n4390) & (!x11742x)) + ((!n_n4324) & (!n_n4340) & (n_n4384) & (!n_n4390) & (x11742x)) + ((!n_n4324) & (!n_n4340) & (n_n4384) & (n_n4390) & (!x11742x)) + ((!n_n4324) & (!n_n4340) & (n_n4384) & (n_n4390) & (x11742x)) + ((!n_n4324) & (n_n4340) & (!n_n4384) & (!n_n4390) & (!x11742x)) + ((!n_n4324) & (n_n4340) & (!n_n4384) & (!n_n4390) & (x11742x)) + ((!n_n4324) & (n_n4340) & (!n_n4384) & (n_n4390) & (!x11742x)) + ((!n_n4324) & (n_n4340) & (!n_n4384) & (n_n4390) & (x11742x)) + ((!n_n4324) & (n_n4340) & (n_n4384) & (!n_n4390) & (!x11742x)) + ((!n_n4324) & (n_n4340) & (n_n4384) & (!n_n4390) & (x11742x)) + ((!n_n4324) & (n_n4340) & (n_n4384) & (n_n4390) & (!x11742x)) + ((!n_n4324) & (n_n4340) & (n_n4384) & (n_n4390) & (x11742x)) + ((n_n4324) & (!n_n4340) & (!n_n4384) & (!n_n4390) & (!x11742x)) + ((n_n4324) & (!n_n4340) & (!n_n4384) & (!n_n4390) & (x11742x)) + ((n_n4324) & (!n_n4340) & (!n_n4384) & (n_n4390) & (!x11742x)) + ((n_n4324) & (!n_n4340) & (!n_n4384) & (n_n4390) & (x11742x)) + ((n_n4324) & (!n_n4340) & (n_n4384) & (!n_n4390) & (!x11742x)) + ((n_n4324) & (!n_n4340) & (n_n4384) & (!n_n4390) & (x11742x)) + ((n_n4324) & (!n_n4340) & (n_n4384) & (n_n4390) & (!x11742x)) + ((n_n4324) & (!n_n4340) & (n_n4384) & (n_n4390) & (x11742x)) + ((n_n4324) & (n_n4340) & (!n_n4384) & (!n_n4390) & (!x11742x)) + ((n_n4324) & (n_n4340) & (!n_n4384) & (!n_n4390) & (x11742x)) + ((n_n4324) & (n_n4340) & (!n_n4384) & (n_n4390) & (!x11742x)) + ((n_n4324) & (n_n4340) & (!n_n4384) & (n_n4390) & (x11742x)) + ((n_n4324) & (n_n4340) & (n_n4384) & (!n_n4390) & (!x11742x)) + ((n_n4324) & (n_n4340) & (n_n4384) & (!n_n4390) & (x11742x)) + ((n_n4324) & (n_n4340) & (n_n4384) & (n_n4390) & (!x11742x)) + ((n_n4324) & (n_n4340) & (n_n4384) & (n_n4390) & (x11742x)));
	assign x11828x = (((!i_7_) & (!i_8_) & (!i_6_) & (x17x) & (n_n491)) + ((!i_7_) & (!i_8_) & (i_6_) & (x17x) & (n_n491)) + ((!i_7_) & (i_8_) & (i_6_) & (x17x) & (n_n491)) + ((i_7_) & (!i_8_) & (!i_6_) & (x17x) & (n_n491)));
	assign x11889x = (((!n_n4782) & (!n_n4779) & (!n_n4786) & (!n_n4780) & (n_n4775)) + ((!n_n4782) & (!n_n4779) & (!n_n4786) & (n_n4780) & (!n_n4775)) + ((!n_n4782) & (!n_n4779) & (!n_n4786) & (n_n4780) & (n_n4775)) + ((!n_n4782) & (!n_n4779) & (n_n4786) & (!n_n4780) & (!n_n4775)) + ((!n_n4782) & (!n_n4779) & (n_n4786) & (!n_n4780) & (n_n4775)) + ((!n_n4782) & (!n_n4779) & (n_n4786) & (n_n4780) & (!n_n4775)) + ((!n_n4782) & (!n_n4779) & (n_n4786) & (n_n4780) & (n_n4775)) + ((!n_n4782) & (n_n4779) & (!n_n4786) & (!n_n4780) & (!n_n4775)) + ((!n_n4782) & (n_n4779) & (!n_n4786) & (!n_n4780) & (n_n4775)) + ((!n_n4782) & (n_n4779) & (!n_n4786) & (n_n4780) & (!n_n4775)) + ((!n_n4782) & (n_n4779) & (!n_n4786) & (n_n4780) & (n_n4775)) + ((!n_n4782) & (n_n4779) & (n_n4786) & (!n_n4780) & (!n_n4775)) + ((!n_n4782) & (n_n4779) & (n_n4786) & (!n_n4780) & (n_n4775)) + ((!n_n4782) & (n_n4779) & (n_n4786) & (n_n4780) & (!n_n4775)) + ((!n_n4782) & (n_n4779) & (n_n4786) & (n_n4780) & (n_n4775)) + ((n_n4782) & (!n_n4779) & (!n_n4786) & (!n_n4780) & (!n_n4775)) + ((n_n4782) & (!n_n4779) & (!n_n4786) & (!n_n4780) & (n_n4775)) + ((n_n4782) & (!n_n4779) & (!n_n4786) & (n_n4780) & (!n_n4775)) + ((n_n4782) & (!n_n4779) & (!n_n4786) & (n_n4780) & (n_n4775)) + ((n_n4782) & (!n_n4779) & (n_n4786) & (!n_n4780) & (!n_n4775)) + ((n_n4782) & (!n_n4779) & (n_n4786) & (!n_n4780) & (n_n4775)) + ((n_n4782) & (!n_n4779) & (n_n4786) & (n_n4780) & (!n_n4775)) + ((n_n4782) & (!n_n4779) & (n_n4786) & (n_n4780) & (n_n4775)) + ((n_n4782) & (n_n4779) & (!n_n4786) & (!n_n4780) & (!n_n4775)) + ((n_n4782) & (n_n4779) & (!n_n4786) & (!n_n4780) & (n_n4775)) + ((n_n4782) & (n_n4779) & (!n_n4786) & (n_n4780) & (!n_n4775)) + ((n_n4782) & (n_n4779) & (!n_n4786) & (n_n4780) & (n_n4775)) + ((n_n4782) & (n_n4779) & (n_n4786) & (!n_n4780) & (!n_n4775)) + ((n_n4782) & (n_n4779) & (n_n4786) & (!n_n4780) & (n_n4775)) + ((n_n4782) & (n_n4779) & (n_n4786) & (n_n4780) & (!n_n4775)) + ((n_n4782) & (n_n4779) & (n_n4786) & (n_n4780) & (n_n4775)));
	assign x11959x = (((!n_n5239) & (!n_n5230) & (!n_n5233) & (!n_n5236) & (n_n5237)) + ((!n_n5239) & (!n_n5230) & (!n_n5233) & (n_n5236) & (!n_n5237)) + ((!n_n5239) & (!n_n5230) & (!n_n5233) & (n_n5236) & (n_n5237)) + ((!n_n5239) & (!n_n5230) & (n_n5233) & (!n_n5236) & (!n_n5237)) + ((!n_n5239) & (!n_n5230) & (n_n5233) & (!n_n5236) & (n_n5237)) + ((!n_n5239) & (!n_n5230) & (n_n5233) & (n_n5236) & (!n_n5237)) + ((!n_n5239) & (!n_n5230) & (n_n5233) & (n_n5236) & (n_n5237)) + ((!n_n5239) & (n_n5230) & (!n_n5233) & (!n_n5236) & (!n_n5237)) + ((!n_n5239) & (n_n5230) & (!n_n5233) & (!n_n5236) & (n_n5237)) + ((!n_n5239) & (n_n5230) & (!n_n5233) & (n_n5236) & (!n_n5237)) + ((!n_n5239) & (n_n5230) & (!n_n5233) & (n_n5236) & (n_n5237)) + ((!n_n5239) & (n_n5230) & (n_n5233) & (!n_n5236) & (!n_n5237)) + ((!n_n5239) & (n_n5230) & (n_n5233) & (!n_n5236) & (n_n5237)) + ((!n_n5239) & (n_n5230) & (n_n5233) & (n_n5236) & (!n_n5237)) + ((!n_n5239) & (n_n5230) & (n_n5233) & (n_n5236) & (n_n5237)) + ((n_n5239) & (!n_n5230) & (!n_n5233) & (!n_n5236) & (!n_n5237)) + ((n_n5239) & (!n_n5230) & (!n_n5233) & (!n_n5236) & (n_n5237)) + ((n_n5239) & (!n_n5230) & (!n_n5233) & (n_n5236) & (!n_n5237)) + ((n_n5239) & (!n_n5230) & (!n_n5233) & (n_n5236) & (n_n5237)) + ((n_n5239) & (!n_n5230) & (n_n5233) & (!n_n5236) & (!n_n5237)) + ((n_n5239) & (!n_n5230) & (n_n5233) & (!n_n5236) & (n_n5237)) + ((n_n5239) & (!n_n5230) & (n_n5233) & (n_n5236) & (!n_n5237)) + ((n_n5239) & (!n_n5230) & (n_n5233) & (n_n5236) & (n_n5237)) + ((n_n5239) & (n_n5230) & (!n_n5233) & (!n_n5236) & (!n_n5237)) + ((n_n5239) & (n_n5230) & (!n_n5233) & (!n_n5236) & (n_n5237)) + ((n_n5239) & (n_n5230) & (!n_n5233) & (n_n5236) & (!n_n5237)) + ((n_n5239) & (n_n5230) & (!n_n5233) & (n_n5236) & (n_n5237)) + ((n_n5239) & (n_n5230) & (n_n5233) & (!n_n5236) & (!n_n5237)) + ((n_n5239) & (n_n5230) & (n_n5233) & (!n_n5236) & (n_n5237)) + ((n_n5239) & (n_n5230) & (n_n5233) & (n_n5236) & (!n_n5237)) + ((n_n5239) & (n_n5230) & (n_n5233) & (n_n5236) & (n_n5237)));
	assign x22192x = (((!n_n5244) & (!n_n5247) & (!n_n5246) & (!n_n5249) & (!n_n1139)));
	assign x12033x = (((!n_n5149) & (!n_n5138) & (!x125x) & (n_n5143)) + ((!n_n5149) & (!n_n5138) & (x125x) & (!n_n5143)) + ((!n_n5149) & (!n_n5138) & (x125x) & (n_n5143)) + ((!n_n5149) & (n_n5138) & (!x125x) & (!n_n5143)) + ((!n_n5149) & (n_n5138) & (!x125x) & (n_n5143)) + ((!n_n5149) & (n_n5138) & (x125x) & (!n_n5143)) + ((!n_n5149) & (n_n5138) & (x125x) & (n_n5143)) + ((n_n5149) & (!n_n5138) & (!x125x) & (!n_n5143)) + ((n_n5149) & (!n_n5138) & (!x125x) & (n_n5143)) + ((n_n5149) & (!n_n5138) & (x125x) & (!n_n5143)) + ((n_n5149) & (!n_n5138) & (x125x) & (n_n5143)) + ((n_n5149) & (n_n5138) & (!x125x) & (!n_n5143)) + ((n_n5149) & (n_n5138) & (!x125x) & (n_n5143)) + ((n_n5149) & (n_n5138) & (x125x) & (!n_n5143)) + ((n_n5149) & (n_n5138) & (x125x) & (n_n5143)));
	assign x12128x = (((!n_n5321) & (!n_n5326) & (!n_n5302) & (!n_n5294) & (n_n5335)) + ((!n_n5321) & (!n_n5326) & (!n_n5302) & (n_n5294) & (!n_n5335)) + ((!n_n5321) & (!n_n5326) & (!n_n5302) & (n_n5294) & (n_n5335)) + ((!n_n5321) & (!n_n5326) & (n_n5302) & (!n_n5294) & (!n_n5335)) + ((!n_n5321) & (!n_n5326) & (n_n5302) & (!n_n5294) & (n_n5335)) + ((!n_n5321) & (!n_n5326) & (n_n5302) & (n_n5294) & (!n_n5335)) + ((!n_n5321) & (!n_n5326) & (n_n5302) & (n_n5294) & (n_n5335)) + ((!n_n5321) & (n_n5326) & (!n_n5302) & (!n_n5294) & (!n_n5335)) + ((!n_n5321) & (n_n5326) & (!n_n5302) & (!n_n5294) & (n_n5335)) + ((!n_n5321) & (n_n5326) & (!n_n5302) & (n_n5294) & (!n_n5335)) + ((!n_n5321) & (n_n5326) & (!n_n5302) & (n_n5294) & (n_n5335)) + ((!n_n5321) & (n_n5326) & (n_n5302) & (!n_n5294) & (!n_n5335)) + ((!n_n5321) & (n_n5326) & (n_n5302) & (!n_n5294) & (n_n5335)) + ((!n_n5321) & (n_n5326) & (n_n5302) & (n_n5294) & (!n_n5335)) + ((!n_n5321) & (n_n5326) & (n_n5302) & (n_n5294) & (n_n5335)) + ((n_n5321) & (!n_n5326) & (!n_n5302) & (!n_n5294) & (!n_n5335)) + ((n_n5321) & (!n_n5326) & (!n_n5302) & (!n_n5294) & (n_n5335)) + ((n_n5321) & (!n_n5326) & (!n_n5302) & (n_n5294) & (!n_n5335)) + ((n_n5321) & (!n_n5326) & (!n_n5302) & (n_n5294) & (n_n5335)) + ((n_n5321) & (!n_n5326) & (n_n5302) & (!n_n5294) & (!n_n5335)) + ((n_n5321) & (!n_n5326) & (n_n5302) & (!n_n5294) & (n_n5335)) + ((n_n5321) & (!n_n5326) & (n_n5302) & (n_n5294) & (!n_n5335)) + ((n_n5321) & (!n_n5326) & (n_n5302) & (n_n5294) & (n_n5335)) + ((n_n5321) & (n_n5326) & (!n_n5302) & (!n_n5294) & (!n_n5335)) + ((n_n5321) & (n_n5326) & (!n_n5302) & (!n_n5294) & (n_n5335)) + ((n_n5321) & (n_n5326) & (!n_n5302) & (n_n5294) & (!n_n5335)) + ((n_n5321) & (n_n5326) & (!n_n5302) & (n_n5294) & (n_n5335)) + ((n_n5321) & (n_n5326) & (n_n5302) & (!n_n5294) & (!n_n5335)) + ((n_n5321) & (n_n5326) & (n_n5302) & (!n_n5294) & (n_n5335)) + ((n_n5321) & (n_n5326) & (n_n5302) & (n_n5294) & (!n_n5335)) + ((n_n5321) & (n_n5326) & (n_n5302) & (n_n5294) & (n_n5335)));
	assign x12146x = (((!n_n4400) & (!n_n4383) & (!n_n4369) & (n_n4372)) + ((!n_n4400) & (!n_n4383) & (n_n4369) & (!n_n4372)) + ((!n_n4400) & (!n_n4383) & (n_n4369) & (n_n4372)) + ((!n_n4400) & (n_n4383) & (!n_n4369) & (!n_n4372)) + ((!n_n4400) & (n_n4383) & (!n_n4369) & (n_n4372)) + ((!n_n4400) & (n_n4383) & (n_n4369) & (!n_n4372)) + ((!n_n4400) & (n_n4383) & (n_n4369) & (n_n4372)) + ((n_n4400) & (!n_n4383) & (!n_n4369) & (!n_n4372)) + ((n_n4400) & (!n_n4383) & (!n_n4369) & (n_n4372)) + ((n_n4400) & (!n_n4383) & (n_n4369) & (!n_n4372)) + ((n_n4400) & (!n_n4383) & (n_n4369) & (n_n4372)) + ((n_n4400) & (n_n4383) & (!n_n4369) & (!n_n4372)) + ((n_n4400) & (n_n4383) & (!n_n4369) & (n_n4372)) + ((n_n4400) & (n_n4383) & (n_n4369) & (!n_n4372)) + ((n_n4400) & (n_n4383) & (n_n4369) & (n_n4372)));
	assign x12147x = (((!n_n4397) & (!n_n4360) & (!x423x) & (n_n4375)) + ((!n_n4397) & (!n_n4360) & (x423x) & (!n_n4375)) + ((!n_n4397) & (!n_n4360) & (x423x) & (n_n4375)) + ((!n_n4397) & (n_n4360) & (!x423x) & (!n_n4375)) + ((!n_n4397) & (n_n4360) & (!x423x) & (n_n4375)) + ((!n_n4397) & (n_n4360) & (x423x) & (!n_n4375)) + ((!n_n4397) & (n_n4360) & (x423x) & (n_n4375)) + ((n_n4397) & (!n_n4360) & (!x423x) & (!n_n4375)) + ((n_n4397) & (!n_n4360) & (!x423x) & (n_n4375)) + ((n_n4397) & (!n_n4360) & (x423x) & (!n_n4375)) + ((n_n4397) & (!n_n4360) & (x423x) & (n_n4375)) + ((n_n4397) & (n_n4360) & (!x423x) & (!n_n4375)) + ((n_n4397) & (n_n4360) & (!x423x) & (n_n4375)) + ((n_n4397) & (n_n4360) & (x423x) & (!n_n4375)) + ((n_n4397) & (n_n4360) & (x423x) & (n_n4375)));
	assign x12196x = (((!n_n4963) & (!n_n4964) & (!n_n4968) & (!n_n4962) & (n_n4973)) + ((!n_n4963) & (!n_n4964) & (!n_n4968) & (n_n4962) & (!n_n4973)) + ((!n_n4963) & (!n_n4964) & (!n_n4968) & (n_n4962) & (n_n4973)) + ((!n_n4963) & (!n_n4964) & (n_n4968) & (!n_n4962) & (!n_n4973)) + ((!n_n4963) & (!n_n4964) & (n_n4968) & (!n_n4962) & (n_n4973)) + ((!n_n4963) & (!n_n4964) & (n_n4968) & (n_n4962) & (!n_n4973)) + ((!n_n4963) & (!n_n4964) & (n_n4968) & (n_n4962) & (n_n4973)) + ((!n_n4963) & (n_n4964) & (!n_n4968) & (!n_n4962) & (!n_n4973)) + ((!n_n4963) & (n_n4964) & (!n_n4968) & (!n_n4962) & (n_n4973)) + ((!n_n4963) & (n_n4964) & (!n_n4968) & (n_n4962) & (!n_n4973)) + ((!n_n4963) & (n_n4964) & (!n_n4968) & (n_n4962) & (n_n4973)) + ((!n_n4963) & (n_n4964) & (n_n4968) & (!n_n4962) & (!n_n4973)) + ((!n_n4963) & (n_n4964) & (n_n4968) & (!n_n4962) & (n_n4973)) + ((!n_n4963) & (n_n4964) & (n_n4968) & (n_n4962) & (!n_n4973)) + ((!n_n4963) & (n_n4964) & (n_n4968) & (n_n4962) & (n_n4973)) + ((n_n4963) & (!n_n4964) & (!n_n4968) & (!n_n4962) & (!n_n4973)) + ((n_n4963) & (!n_n4964) & (!n_n4968) & (!n_n4962) & (n_n4973)) + ((n_n4963) & (!n_n4964) & (!n_n4968) & (n_n4962) & (!n_n4973)) + ((n_n4963) & (!n_n4964) & (!n_n4968) & (n_n4962) & (n_n4973)) + ((n_n4963) & (!n_n4964) & (n_n4968) & (!n_n4962) & (!n_n4973)) + ((n_n4963) & (!n_n4964) & (n_n4968) & (!n_n4962) & (n_n4973)) + ((n_n4963) & (!n_n4964) & (n_n4968) & (n_n4962) & (!n_n4973)) + ((n_n4963) & (!n_n4964) & (n_n4968) & (n_n4962) & (n_n4973)) + ((n_n4963) & (n_n4964) & (!n_n4968) & (!n_n4962) & (!n_n4973)) + ((n_n4963) & (n_n4964) & (!n_n4968) & (!n_n4962) & (n_n4973)) + ((n_n4963) & (n_n4964) & (!n_n4968) & (n_n4962) & (!n_n4973)) + ((n_n4963) & (n_n4964) & (!n_n4968) & (n_n4962) & (n_n4973)) + ((n_n4963) & (n_n4964) & (n_n4968) & (!n_n4962) & (!n_n4973)) + ((n_n4963) & (n_n4964) & (n_n4968) & (!n_n4962) & (n_n4973)) + ((n_n4963) & (n_n4964) & (n_n4968) & (n_n4962) & (!n_n4973)) + ((n_n4963) & (n_n4964) & (n_n4968) & (n_n4962) & (n_n4973)));
	assign x12385x = (((!n_n482) & (!n_n532) & (!x18x) & (!n_n5027) & (x253x)) + ((!n_n482) & (!n_n532) & (!x18x) & (n_n5027) & (!x253x)) + ((!n_n482) & (!n_n532) & (!x18x) & (n_n5027) & (x253x)) + ((!n_n482) & (!n_n532) & (x18x) & (!n_n5027) & (x253x)) + ((!n_n482) & (!n_n532) & (x18x) & (n_n5027) & (!x253x)) + ((!n_n482) & (!n_n532) & (x18x) & (n_n5027) & (x253x)) + ((!n_n482) & (n_n532) & (!x18x) & (!n_n5027) & (x253x)) + ((!n_n482) & (n_n532) & (!x18x) & (n_n5027) & (!x253x)) + ((!n_n482) & (n_n532) & (!x18x) & (n_n5027) & (x253x)) + ((!n_n482) & (n_n532) & (x18x) & (!n_n5027) & (x253x)) + ((!n_n482) & (n_n532) & (x18x) & (n_n5027) & (!x253x)) + ((!n_n482) & (n_n532) & (x18x) & (n_n5027) & (x253x)) + ((n_n482) & (!n_n532) & (!x18x) & (!n_n5027) & (x253x)) + ((n_n482) & (!n_n532) & (!x18x) & (n_n5027) & (!x253x)) + ((n_n482) & (!n_n532) & (!x18x) & (n_n5027) & (x253x)) + ((n_n482) & (!n_n532) & (x18x) & (!n_n5027) & (x253x)) + ((n_n482) & (!n_n532) & (x18x) & (n_n5027) & (!x253x)) + ((n_n482) & (!n_n532) & (x18x) & (n_n5027) & (x253x)) + ((n_n482) & (n_n532) & (!x18x) & (!n_n5027) & (x253x)) + ((n_n482) & (n_n532) & (!x18x) & (n_n5027) & (!x253x)) + ((n_n482) & (n_n532) & (!x18x) & (n_n5027) & (x253x)) + ((n_n482) & (n_n532) & (x18x) & (!n_n5027) & (!x253x)) + ((n_n482) & (n_n532) & (x18x) & (!n_n5027) & (x253x)) + ((n_n482) & (n_n532) & (x18x) & (n_n5027) & (!x253x)) + ((n_n482) & (n_n532) & (x18x) & (n_n5027) & (x253x)));
	assign x12386x = (((!n_n5038) & (!n_n5035) & (!n_n5031) & (!n_n5037) & (n_n5029)) + ((!n_n5038) & (!n_n5035) & (!n_n5031) & (n_n5037) & (!n_n5029)) + ((!n_n5038) & (!n_n5035) & (!n_n5031) & (n_n5037) & (n_n5029)) + ((!n_n5038) & (!n_n5035) & (n_n5031) & (!n_n5037) & (!n_n5029)) + ((!n_n5038) & (!n_n5035) & (n_n5031) & (!n_n5037) & (n_n5029)) + ((!n_n5038) & (!n_n5035) & (n_n5031) & (n_n5037) & (!n_n5029)) + ((!n_n5038) & (!n_n5035) & (n_n5031) & (n_n5037) & (n_n5029)) + ((!n_n5038) & (n_n5035) & (!n_n5031) & (!n_n5037) & (!n_n5029)) + ((!n_n5038) & (n_n5035) & (!n_n5031) & (!n_n5037) & (n_n5029)) + ((!n_n5038) & (n_n5035) & (!n_n5031) & (n_n5037) & (!n_n5029)) + ((!n_n5038) & (n_n5035) & (!n_n5031) & (n_n5037) & (n_n5029)) + ((!n_n5038) & (n_n5035) & (n_n5031) & (!n_n5037) & (!n_n5029)) + ((!n_n5038) & (n_n5035) & (n_n5031) & (!n_n5037) & (n_n5029)) + ((!n_n5038) & (n_n5035) & (n_n5031) & (n_n5037) & (!n_n5029)) + ((!n_n5038) & (n_n5035) & (n_n5031) & (n_n5037) & (n_n5029)) + ((n_n5038) & (!n_n5035) & (!n_n5031) & (!n_n5037) & (!n_n5029)) + ((n_n5038) & (!n_n5035) & (!n_n5031) & (!n_n5037) & (n_n5029)) + ((n_n5038) & (!n_n5035) & (!n_n5031) & (n_n5037) & (!n_n5029)) + ((n_n5038) & (!n_n5035) & (!n_n5031) & (n_n5037) & (n_n5029)) + ((n_n5038) & (!n_n5035) & (n_n5031) & (!n_n5037) & (!n_n5029)) + ((n_n5038) & (!n_n5035) & (n_n5031) & (!n_n5037) & (n_n5029)) + ((n_n5038) & (!n_n5035) & (n_n5031) & (n_n5037) & (!n_n5029)) + ((n_n5038) & (!n_n5035) & (n_n5031) & (n_n5037) & (n_n5029)) + ((n_n5038) & (n_n5035) & (!n_n5031) & (!n_n5037) & (!n_n5029)) + ((n_n5038) & (n_n5035) & (!n_n5031) & (!n_n5037) & (n_n5029)) + ((n_n5038) & (n_n5035) & (!n_n5031) & (n_n5037) & (!n_n5029)) + ((n_n5038) & (n_n5035) & (!n_n5031) & (n_n5037) & (n_n5029)) + ((n_n5038) & (n_n5035) & (n_n5031) & (!n_n5037) & (!n_n5029)) + ((n_n5038) & (n_n5035) & (n_n5031) & (!n_n5037) & (n_n5029)) + ((n_n5038) & (n_n5035) & (n_n5031) & (n_n5037) & (!n_n5029)) + ((n_n5038) & (n_n5035) & (n_n5031) & (n_n5037) & (n_n5029)));
	assign x22170x = (((!n_n518) & (!n_n390) & (!x23x) & (!n_n4601) & (!n_n4600)) + ((!n_n518) & (!n_n390) & (x23x) & (!n_n4601) & (!n_n4600)) + ((!n_n518) & (n_n390) & (!x23x) & (!n_n4601) & (!n_n4600)) + ((!n_n518) & (n_n390) & (x23x) & (!n_n4601) & (!n_n4600)) + ((n_n518) & (!n_n390) & (!x23x) & (!n_n4601) & (!n_n4600)) + ((n_n518) & (!n_n390) & (x23x) & (!n_n4601) & (!n_n4600)) + ((n_n518) & (n_n390) & (!x23x) & (!n_n4601) & (!n_n4600)));
	assign x12669x = (((!n_n491) & (!n_n520) & (!x18x) & (!n_n5027) & (n_n5048)) + ((!n_n491) & (!n_n520) & (!x18x) & (n_n5027) & (!n_n5048)) + ((!n_n491) & (!n_n520) & (!x18x) & (n_n5027) & (n_n5048)) + ((!n_n491) & (!n_n520) & (x18x) & (!n_n5027) & (n_n5048)) + ((!n_n491) & (!n_n520) & (x18x) & (n_n5027) & (!n_n5048)) + ((!n_n491) & (!n_n520) & (x18x) & (n_n5027) & (n_n5048)) + ((!n_n491) & (n_n520) & (!x18x) & (!n_n5027) & (n_n5048)) + ((!n_n491) & (n_n520) & (!x18x) & (n_n5027) & (!n_n5048)) + ((!n_n491) & (n_n520) & (!x18x) & (n_n5027) & (n_n5048)) + ((!n_n491) & (n_n520) & (x18x) & (!n_n5027) & (n_n5048)) + ((!n_n491) & (n_n520) & (x18x) & (n_n5027) & (!n_n5048)) + ((!n_n491) & (n_n520) & (x18x) & (n_n5027) & (n_n5048)) + ((n_n491) & (!n_n520) & (!x18x) & (!n_n5027) & (n_n5048)) + ((n_n491) & (!n_n520) & (!x18x) & (n_n5027) & (!n_n5048)) + ((n_n491) & (!n_n520) & (!x18x) & (n_n5027) & (n_n5048)) + ((n_n491) & (!n_n520) & (x18x) & (!n_n5027) & (n_n5048)) + ((n_n491) & (!n_n520) & (x18x) & (n_n5027) & (!n_n5048)) + ((n_n491) & (!n_n520) & (x18x) & (n_n5027) & (n_n5048)) + ((n_n491) & (n_n520) & (!x18x) & (!n_n5027) & (n_n5048)) + ((n_n491) & (n_n520) & (!x18x) & (n_n5027) & (!n_n5048)) + ((n_n491) & (n_n520) & (!x18x) & (n_n5027) & (n_n5048)) + ((n_n491) & (n_n520) & (x18x) & (!n_n5027) & (!n_n5048)) + ((n_n491) & (n_n520) & (x18x) & (!n_n5027) & (n_n5048)) + ((n_n491) & (n_n520) & (x18x) & (n_n5027) & (!n_n5048)) + ((n_n491) & (n_n520) & (x18x) & (n_n5027) & (n_n5048)));
	assign x12741x = (((!i_7_) & (!i_8_) & (!i_6_) & (x17x) & (n_n535)) + ((!i_7_) & (i_8_) & (!i_6_) & (x17x) & (n_n535)) + ((i_7_) & (!i_8_) & (!i_6_) & (x17x) & (n_n535)));
	assign x12772x = (((!n_n4887) & (!x262x) & (!n_n4880) & (n_n4891)) + ((!n_n4887) & (!x262x) & (n_n4880) & (!n_n4891)) + ((!n_n4887) & (!x262x) & (n_n4880) & (n_n4891)) + ((!n_n4887) & (x262x) & (!n_n4880) & (!n_n4891)) + ((!n_n4887) & (x262x) & (!n_n4880) & (n_n4891)) + ((!n_n4887) & (x262x) & (n_n4880) & (!n_n4891)) + ((!n_n4887) & (x262x) & (n_n4880) & (n_n4891)) + ((n_n4887) & (!x262x) & (!n_n4880) & (!n_n4891)) + ((n_n4887) & (!x262x) & (!n_n4880) & (n_n4891)) + ((n_n4887) & (!x262x) & (n_n4880) & (!n_n4891)) + ((n_n4887) & (!x262x) & (n_n4880) & (n_n4891)) + ((n_n4887) & (x262x) & (!n_n4880) & (!n_n4891)) + ((n_n4887) & (x262x) & (!n_n4880) & (n_n4891)) + ((n_n4887) & (x262x) & (n_n4880) & (!n_n4891)) + ((n_n4887) & (x262x) & (n_n4880) & (n_n4891)));
	assign x22174x = (((!n_n4920) & (!n_n4916) & (!n_n4908) & (!n_n4919)));
	assign x12863x = (((!n_n4912) & (!x351x) & (!n_n4915) & (!n_n4910) & (!x22174x)) + ((!n_n4912) & (!x351x) & (!n_n4915) & (n_n4910) & (!x22174x)) + ((!n_n4912) & (!x351x) & (!n_n4915) & (n_n4910) & (x22174x)) + ((!n_n4912) & (!x351x) & (n_n4915) & (!n_n4910) & (!x22174x)) + ((!n_n4912) & (!x351x) & (n_n4915) & (!n_n4910) & (x22174x)) + ((!n_n4912) & (!x351x) & (n_n4915) & (n_n4910) & (!x22174x)) + ((!n_n4912) & (!x351x) & (n_n4915) & (n_n4910) & (x22174x)) + ((!n_n4912) & (x351x) & (!n_n4915) & (!n_n4910) & (!x22174x)) + ((!n_n4912) & (x351x) & (!n_n4915) & (!n_n4910) & (x22174x)) + ((!n_n4912) & (x351x) & (!n_n4915) & (n_n4910) & (!x22174x)) + ((!n_n4912) & (x351x) & (!n_n4915) & (n_n4910) & (x22174x)) + ((!n_n4912) & (x351x) & (n_n4915) & (!n_n4910) & (!x22174x)) + ((!n_n4912) & (x351x) & (n_n4915) & (!n_n4910) & (x22174x)) + ((!n_n4912) & (x351x) & (n_n4915) & (n_n4910) & (!x22174x)) + ((!n_n4912) & (x351x) & (n_n4915) & (n_n4910) & (x22174x)) + ((n_n4912) & (!x351x) & (!n_n4915) & (!n_n4910) & (!x22174x)) + ((n_n4912) & (!x351x) & (!n_n4915) & (!n_n4910) & (x22174x)) + ((n_n4912) & (!x351x) & (!n_n4915) & (n_n4910) & (!x22174x)) + ((n_n4912) & (!x351x) & (!n_n4915) & (n_n4910) & (x22174x)) + ((n_n4912) & (!x351x) & (n_n4915) & (!n_n4910) & (!x22174x)) + ((n_n4912) & (!x351x) & (n_n4915) & (!n_n4910) & (x22174x)) + ((n_n4912) & (!x351x) & (n_n4915) & (n_n4910) & (!x22174x)) + ((n_n4912) & (!x351x) & (n_n4915) & (n_n4910) & (x22174x)) + ((n_n4912) & (x351x) & (!n_n4915) & (!n_n4910) & (!x22174x)) + ((n_n4912) & (x351x) & (!n_n4915) & (!n_n4910) & (x22174x)) + ((n_n4912) & (x351x) & (!n_n4915) & (n_n4910) & (!x22174x)) + ((n_n4912) & (x351x) & (!n_n4915) & (n_n4910) & (x22174x)) + ((n_n4912) & (x351x) & (n_n4915) & (!n_n4910) & (!x22174x)) + ((n_n4912) & (x351x) & (n_n4915) & (!n_n4910) & (x22174x)) + ((n_n4912) & (x351x) & (n_n4915) & (n_n4910) & (!x22174x)) + ((n_n4912) & (x351x) & (n_n4915) & (n_n4910) & (x22174x)));
	assign x22129x = (((!n_n526) & (!n_n482) & (!n_n195) & (!n_n530)) + ((!n_n526) & (!n_n482) & (!n_n195) & (n_n530)) + ((!n_n526) & (!n_n482) & (n_n195) & (!n_n530)) + ((!n_n526) & (!n_n482) & (n_n195) & (n_n530)) + ((!n_n526) & (n_n482) & (!n_n195) & (!n_n530)) + ((!n_n526) & (n_n482) & (!n_n195) & (n_n530)) + ((!n_n526) & (n_n482) & (n_n195) & (!n_n530)) + ((n_n526) & (!n_n482) & (!n_n195) & (!n_n530)) + ((n_n526) & (!n_n482) & (!n_n195) & (n_n530)) + ((n_n526) & (!n_n482) & (n_n195) & (!n_n530)) + ((n_n526) & (!n_n482) & (n_n195) & (n_n530)) + ((n_n526) & (n_n482) & (!n_n195) & (!n_n530)) + ((n_n526) & (n_n482) & (!n_n195) & (n_n530)));
	assign x12980x = (((!n_n5290) & (!n_n5289) & (!x208x) & (n_n5298)) + ((!n_n5290) & (!n_n5289) & (x208x) & (!n_n5298)) + ((!n_n5290) & (!n_n5289) & (x208x) & (n_n5298)) + ((!n_n5290) & (n_n5289) & (!x208x) & (!n_n5298)) + ((!n_n5290) & (n_n5289) & (!x208x) & (n_n5298)) + ((!n_n5290) & (n_n5289) & (x208x) & (!n_n5298)) + ((!n_n5290) & (n_n5289) & (x208x) & (n_n5298)) + ((n_n5290) & (!n_n5289) & (!x208x) & (!n_n5298)) + ((n_n5290) & (!n_n5289) & (!x208x) & (n_n5298)) + ((n_n5290) & (!n_n5289) & (x208x) & (!n_n5298)) + ((n_n5290) & (!n_n5289) & (x208x) & (n_n5298)) + ((n_n5290) & (n_n5289) & (!x208x) & (!n_n5298)) + ((n_n5290) & (n_n5289) & (!x208x) & (n_n5298)) + ((n_n5290) & (n_n5289) & (x208x) & (!n_n5298)) + ((n_n5290) & (n_n5289) & (x208x) & (n_n5298)));
	assign x12995x = (((!n_n5171) & (!n_n5181) & (!n_n5184) & (n_n5170)) + ((!n_n5171) & (!n_n5181) & (n_n5184) & (!n_n5170)) + ((!n_n5171) & (!n_n5181) & (n_n5184) & (n_n5170)) + ((!n_n5171) & (n_n5181) & (!n_n5184) & (!n_n5170)) + ((!n_n5171) & (n_n5181) & (!n_n5184) & (n_n5170)) + ((!n_n5171) & (n_n5181) & (n_n5184) & (!n_n5170)) + ((!n_n5171) & (n_n5181) & (n_n5184) & (n_n5170)) + ((n_n5171) & (!n_n5181) & (!n_n5184) & (!n_n5170)) + ((n_n5171) & (!n_n5181) & (!n_n5184) & (n_n5170)) + ((n_n5171) & (!n_n5181) & (n_n5184) & (!n_n5170)) + ((n_n5171) & (!n_n5181) & (n_n5184) & (n_n5170)) + ((n_n5171) & (n_n5181) & (!n_n5184) & (!n_n5170)) + ((n_n5171) & (n_n5181) & (!n_n5184) & (n_n5170)) + ((n_n5171) & (n_n5181) & (n_n5184) & (!n_n5170)) + ((n_n5171) & (n_n5181) & (n_n5184) & (n_n5170)));
	assign x12996x = (((!n_n5174) & (!n_n5175) & (!n_n5177) & (!n_n5172) & (n_n5176)) + ((!n_n5174) & (!n_n5175) & (!n_n5177) & (n_n5172) & (!n_n5176)) + ((!n_n5174) & (!n_n5175) & (!n_n5177) & (n_n5172) & (n_n5176)) + ((!n_n5174) & (!n_n5175) & (n_n5177) & (!n_n5172) & (!n_n5176)) + ((!n_n5174) & (!n_n5175) & (n_n5177) & (!n_n5172) & (n_n5176)) + ((!n_n5174) & (!n_n5175) & (n_n5177) & (n_n5172) & (!n_n5176)) + ((!n_n5174) & (!n_n5175) & (n_n5177) & (n_n5172) & (n_n5176)) + ((!n_n5174) & (n_n5175) & (!n_n5177) & (!n_n5172) & (!n_n5176)) + ((!n_n5174) & (n_n5175) & (!n_n5177) & (!n_n5172) & (n_n5176)) + ((!n_n5174) & (n_n5175) & (!n_n5177) & (n_n5172) & (!n_n5176)) + ((!n_n5174) & (n_n5175) & (!n_n5177) & (n_n5172) & (n_n5176)) + ((!n_n5174) & (n_n5175) & (n_n5177) & (!n_n5172) & (!n_n5176)) + ((!n_n5174) & (n_n5175) & (n_n5177) & (!n_n5172) & (n_n5176)) + ((!n_n5174) & (n_n5175) & (n_n5177) & (n_n5172) & (!n_n5176)) + ((!n_n5174) & (n_n5175) & (n_n5177) & (n_n5172) & (n_n5176)) + ((n_n5174) & (!n_n5175) & (!n_n5177) & (!n_n5172) & (!n_n5176)) + ((n_n5174) & (!n_n5175) & (!n_n5177) & (!n_n5172) & (n_n5176)) + ((n_n5174) & (!n_n5175) & (!n_n5177) & (n_n5172) & (!n_n5176)) + ((n_n5174) & (!n_n5175) & (!n_n5177) & (n_n5172) & (n_n5176)) + ((n_n5174) & (!n_n5175) & (n_n5177) & (!n_n5172) & (!n_n5176)) + ((n_n5174) & (!n_n5175) & (n_n5177) & (!n_n5172) & (n_n5176)) + ((n_n5174) & (!n_n5175) & (n_n5177) & (n_n5172) & (!n_n5176)) + ((n_n5174) & (!n_n5175) & (n_n5177) & (n_n5172) & (n_n5176)) + ((n_n5174) & (n_n5175) & (!n_n5177) & (!n_n5172) & (!n_n5176)) + ((n_n5174) & (n_n5175) & (!n_n5177) & (!n_n5172) & (n_n5176)) + ((n_n5174) & (n_n5175) & (!n_n5177) & (n_n5172) & (!n_n5176)) + ((n_n5174) & (n_n5175) & (!n_n5177) & (n_n5172) & (n_n5176)) + ((n_n5174) & (n_n5175) & (n_n5177) & (!n_n5172) & (!n_n5176)) + ((n_n5174) & (n_n5175) & (n_n5177) & (!n_n5172) & (n_n5176)) + ((n_n5174) & (n_n5175) & (n_n5177) & (n_n5172) & (!n_n5176)) + ((n_n5174) & (n_n5175) & (n_n5177) & (n_n5172) & (n_n5176)));
	assign x13126x = (((!i_7_) & (!i_8_) & (i_6_) & (x13x) & (n_n464)) + ((!i_7_) & (i_8_) & (i_6_) & (x13x) & (n_n464)));
	assign x13141x = (((!n_n5305) & (!n_n5293) & (!n_n5296) & (!n_n5284) & (n_n5297)) + ((!n_n5305) & (!n_n5293) & (!n_n5296) & (n_n5284) & (!n_n5297)) + ((!n_n5305) & (!n_n5293) & (!n_n5296) & (n_n5284) & (n_n5297)) + ((!n_n5305) & (!n_n5293) & (n_n5296) & (!n_n5284) & (!n_n5297)) + ((!n_n5305) & (!n_n5293) & (n_n5296) & (!n_n5284) & (n_n5297)) + ((!n_n5305) & (!n_n5293) & (n_n5296) & (n_n5284) & (!n_n5297)) + ((!n_n5305) & (!n_n5293) & (n_n5296) & (n_n5284) & (n_n5297)) + ((!n_n5305) & (n_n5293) & (!n_n5296) & (!n_n5284) & (!n_n5297)) + ((!n_n5305) & (n_n5293) & (!n_n5296) & (!n_n5284) & (n_n5297)) + ((!n_n5305) & (n_n5293) & (!n_n5296) & (n_n5284) & (!n_n5297)) + ((!n_n5305) & (n_n5293) & (!n_n5296) & (n_n5284) & (n_n5297)) + ((!n_n5305) & (n_n5293) & (n_n5296) & (!n_n5284) & (!n_n5297)) + ((!n_n5305) & (n_n5293) & (n_n5296) & (!n_n5284) & (n_n5297)) + ((!n_n5305) & (n_n5293) & (n_n5296) & (n_n5284) & (!n_n5297)) + ((!n_n5305) & (n_n5293) & (n_n5296) & (n_n5284) & (n_n5297)) + ((n_n5305) & (!n_n5293) & (!n_n5296) & (!n_n5284) & (!n_n5297)) + ((n_n5305) & (!n_n5293) & (!n_n5296) & (!n_n5284) & (n_n5297)) + ((n_n5305) & (!n_n5293) & (!n_n5296) & (n_n5284) & (!n_n5297)) + ((n_n5305) & (!n_n5293) & (!n_n5296) & (n_n5284) & (n_n5297)) + ((n_n5305) & (!n_n5293) & (n_n5296) & (!n_n5284) & (!n_n5297)) + ((n_n5305) & (!n_n5293) & (n_n5296) & (!n_n5284) & (n_n5297)) + ((n_n5305) & (!n_n5293) & (n_n5296) & (n_n5284) & (!n_n5297)) + ((n_n5305) & (!n_n5293) & (n_n5296) & (n_n5284) & (n_n5297)) + ((n_n5305) & (n_n5293) & (!n_n5296) & (!n_n5284) & (!n_n5297)) + ((n_n5305) & (n_n5293) & (!n_n5296) & (!n_n5284) & (n_n5297)) + ((n_n5305) & (n_n5293) & (!n_n5296) & (n_n5284) & (!n_n5297)) + ((n_n5305) & (n_n5293) & (!n_n5296) & (n_n5284) & (n_n5297)) + ((n_n5305) & (n_n5293) & (n_n5296) & (!n_n5284) & (!n_n5297)) + ((n_n5305) & (n_n5293) & (n_n5296) & (!n_n5284) & (n_n5297)) + ((n_n5305) & (n_n5293) & (n_n5296) & (n_n5284) & (!n_n5297)) + ((n_n5305) & (n_n5293) & (n_n5296) & (n_n5284) & (n_n5297)));
	assign x13142x = (((!x12700x) & (!x12701x) & (x13141x)) + ((!x12700x) & (x12701x) & (!x13141x)) + ((!x12700x) & (x12701x) & (x13141x)) + ((x12700x) & (!x12701x) & (!x13141x)) + ((x12700x) & (!x12701x) & (x13141x)) + ((x12700x) & (x12701x) & (!x13141x)) + ((x12700x) & (x12701x) & (x13141x)));
	assign x13143x = (((!x12707x) & (!x12708x) & (!x12714x) & (x12715x)) + ((!x12707x) & (!x12708x) & (x12714x) & (!x12715x)) + ((!x12707x) & (!x12708x) & (x12714x) & (x12715x)) + ((!x12707x) & (x12708x) & (!x12714x) & (!x12715x)) + ((!x12707x) & (x12708x) & (!x12714x) & (x12715x)) + ((!x12707x) & (x12708x) & (x12714x) & (!x12715x)) + ((!x12707x) & (x12708x) & (x12714x) & (x12715x)) + ((x12707x) & (!x12708x) & (!x12714x) & (!x12715x)) + ((x12707x) & (!x12708x) & (!x12714x) & (x12715x)) + ((x12707x) & (!x12708x) & (x12714x) & (!x12715x)) + ((x12707x) & (!x12708x) & (x12714x) & (x12715x)) + ((x12707x) & (x12708x) & (!x12714x) & (!x12715x)) + ((x12707x) & (x12708x) & (!x12714x) & (x12715x)) + ((x12707x) & (x12708x) & (x12714x) & (!x12715x)) + ((x12707x) & (x12708x) & (x12714x) & (x12715x)));
	assign x13182x = (((!i_7_) & (!i_8_) & (i_6_) & (n_n482) & (x14x)) + ((i_7_) & (i_8_) & (!i_6_) & (n_n482) & (x14x)));
	assign x13224x = (((!n_n4953) & (!n_n4967) & (!n_n4962) & (n_n4948)) + ((!n_n4953) & (!n_n4967) & (n_n4962) & (!n_n4948)) + ((!n_n4953) & (!n_n4967) & (n_n4962) & (n_n4948)) + ((!n_n4953) & (n_n4967) & (!n_n4962) & (!n_n4948)) + ((!n_n4953) & (n_n4967) & (!n_n4962) & (n_n4948)) + ((!n_n4953) & (n_n4967) & (n_n4962) & (!n_n4948)) + ((!n_n4953) & (n_n4967) & (n_n4962) & (n_n4948)) + ((n_n4953) & (!n_n4967) & (!n_n4962) & (!n_n4948)) + ((n_n4953) & (!n_n4967) & (!n_n4962) & (n_n4948)) + ((n_n4953) & (!n_n4967) & (n_n4962) & (!n_n4948)) + ((n_n4953) & (!n_n4967) & (n_n4962) & (n_n4948)) + ((n_n4953) & (n_n4967) & (!n_n4962) & (!n_n4948)) + ((n_n4953) & (n_n4967) & (!n_n4962) & (n_n4948)) + ((n_n4953) & (n_n4967) & (n_n4962) & (!n_n4948)) + ((n_n4953) & (n_n4967) & (n_n4962) & (n_n4948)));
	assign x22125x = (((!n_n4754) & (!n_n4749) & (!n_n4747) & (!n_n4753)));
	assign x13420x = (((!n_n4988) & (!n_n4989) & (!n_n4980) & (!n_n4985) & (n_n4984)) + ((!n_n4988) & (!n_n4989) & (!n_n4980) & (n_n4985) & (!n_n4984)) + ((!n_n4988) & (!n_n4989) & (!n_n4980) & (n_n4985) & (n_n4984)) + ((!n_n4988) & (!n_n4989) & (n_n4980) & (!n_n4985) & (!n_n4984)) + ((!n_n4988) & (!n_n4989) & (n_n4980) & (!n_n4985) & (n_n4984)) + ((!n_n4988) & (!n_n4989) & (n_n4980) & (n_n4985) & (!n_n4984)) + ((!n_n4988) & (!n_n4989) & (n_n4980) & (n_n4985) & (n_n4984)) + ((!n_n4988) & (n_n4989) & (!n_n4980) & (!n_n4985) & (!n_n4984)) + ((!n_n4988) & (n_n4989) & (!n_n4980) & (!n_n4985) & (n_n4984)) + ((!n_n4988) & (n_n4989) & (!n_n4980) & (n_n4985) & (!n_n4984)) + ((!n_n4988) & (n_n4989) & (!n_n4980) & (n_n4985) & (n_n4984)) + ((!n_n4988) & (n_n4989) & (n_n4980) & (!n_n4985) & (!n_n4984)) + ((!n_n4988) & (n_n4989) & (n_n4980) & (!n_n4985) & (n_n4984)) + ((!n_n4988) & (n_n4989) & (n_n4980) & (n_n4985) & (!n_n4984)) + ((!n_n4988) & (n_n4989) & (n_n4980) & (n_n4985) & (n_n4984)) + ((n_n4988) & (!n_n4989) & (!n_n4980) & (!n_n4985) & (!n_n4984)) + ((n_n4988) & (!n_n4989) & (!n_n4980) & (!n_n4985) & (n_n4984)) + ((n_n4988) & (!n_n4989) & (!n_n4980) & (n_n4985) & (!n_n4984)) + ((n_n4988) & (!n_n4989) & (!n_n4980) & (n_n4985) & (n_n4984)) + ((n_n4988) & (!n_n4989) & (n_n4980) & (!n_n4985) & (!n_n4984)) + ((n_n4988) & (!n_n4989) & (n_n4980) & (!n_n4985) & (n_n4984)) + ((n_n4988) & (!n_n4989) & (n_n4980) & (n_n4985) & (!n_n4984)) + ((n_n4988) & (!n_n4989) & (n_n4980) & (n_n4985) & (n_n4984)) + ((n_n4988) & (n_n4989) & (!n_n4980) & (!n_n4985) & (!n_n4984)) + ((n_n4988) & (n_n4989) & (!n_n4980) & (!n_n4985) & (n_n4984)) + ((n_n4988) & (n_n4989) & (!n_n4980) & (n_n4985) & (!n_n4984)) + ((n_n4988) & (n_n4989) & (!n_n4980) & (n_n4985) & (n_n4984)) + ((n_n4988) & (n_n4989) & (n_n4980) & (!n_n4985) & (!n_n4984)) + ((n_n4988) & (n_n4989) & (n_n4980) & (!n_n4985) & (n_n4984)) + ((n_n4988) & (n_n4989) & (n_n4980) & (n_n4985) & (!n_n4984)) + ((n_n4988) & (n_n4989) & (n_n4980) & (n_n4985) & (n_n4984)));
	assign x13449x = (((!i_9_) & (!n_n528) & (n_n390) & (n_n535) & (n_n530)) + ((!i_9_) & (n_n528) & (n_n390) & (n_n535) & (n_n530)) + ((i_9_) & (!n_n528) & (n_n390) & (n_n535) & (n_n530)) + ((i_9_) & (n_n528) & (n_n390) & (n_n535) & (!n_n530)) + ((i_9_) & (n_n528) & (n_n390) & (n_n535) & (n_n530)));
	assign x13477x = (((!i_9_) & (n_n482) & (n_n455) & (n_n528) & (!n_n520)) + ((!i_9_) & (n_n482) & (n_n455) & (n_n528) & (n_n520)) + ((i_9_) & (n_n482) & (n_n455) & (!n_n528) & (n_n520)) + ((i_9_) & (n_n482) & (n_n455) & (n_n528) & (n_n520)));
	assign x13544x = (((!n_n4360) & (!n_n4370) & (n_n4275)) + ((!n_n4360) & (n_n4370) & (!n_n4275)) + ((!n_n4360) & (n_n4370) & (n_n4275)) + ((n_n4360) & (!n_n4370) & (!n_n4275)) + ((n_n4360) & (!n_n4370) & (n_n4275)) + ((n_n4360) & (n_n4370) & (!n_n4275)) + ((n_n4360) & (n_n4370) & (n_n4275)));
	assign x13551x = (((!n_n4455) & (!n_n3520) & (!n_n4456) & (!n_n4458) & (x55x)) + ((!n_n4455) & (!n_n3520) & (!n_n4456) & (n_n4458) & (!x55x)) + ((!n_n4455) & (!n_n3520) & (!n_n4456) & (n_n4458) & (x55x)) + ((!n_n4455) & (!n_n3520) & (n_n4456) & (!n_n4458) & (!x55x)) + ((!n_n4455) & (!n_n3520) & (n_n4456) & (!n_n4458) & (x55x)) + ((!n_n4455) & (!n_n3520) & (n_n4456) & (n_n4458) & (!x55x)) + ((!n_n4455) & (!n_n3520) & (n_n4456) & (n_n4458) & (x55x)) + ((!n_n4455) & (n_n3520) & (!n_n4456) & (!n_n4458) & (!x55x)) + ((!n_n4455) & (n_n3520) & (!n_n4456) & (!n_n4458) & (x55x)) + ((!n_n4455) & (n_n3520) & (!n_n4456) & (n_n4458) & (!x55x)) + ((!n_n4455) & (n_n3520) & (!n_n4456) & (n_n4458) & (x55x)) + ((!n_n4455) & (n_n3520) & (n_n4456) & (!n_n4458) & (!x55x)) + ((!n_n4455) & (n_n3520) & (n_n4456) & (!n_n4458) & (x55x)) + ((!n_n4455) & (n_n3520) & (n_n4456) & (n_n4458) & (!x55x)) + ((!n_n4455) & (n_n3520) & (n_n4456) & (n_n4458) & (x55x)) + ((n_n4455) & (!n_n3520) & (!n_n4456) & (!n_n4458) & (!x55x)) + ((n_n4455) & (!n_n3520) & (!n_n4456) & (!n_n4458) & (x55x)) + ((n_n4455) & (!n_n3520) & (!n_n4456) & (n_n4458) & (!x55x)) + ((n_n4455) & (!n_n3520) & (!n_n4456) & (n_n4458) & (x55x)) + ((n_n4455) & (!n_n3520) & (n_n4456) & (!n_n4458) & (!x55x)) + ((n_n4455) & (!n_n3520) & (n_n4456) & (!n_n4458) & (x55x)) + ((n_n4455) & (!n_n3520) & (n_n4456) & (n_n4458) & (!x55x)) + ((n_n4455) & (!n_n3520) & (n_n4456) & (n_n4458) & (x55x)) + ((n_n4455) & (n_n3520) & (!n_n4456) & (!n_n4458) & (!x55x)) + ((n_n4455) & (n_n3520) & (!n_n4456) & (!n_n4458) & (x55x)) + ((n_n4455) & (n_n3520) & (!n_n4456) & (n_n4458) & (!x55x)) + ((n_n4455) & (n_n3520) & (!n_n4456) & (n_n4458) & (x55x)) + ((n_n4455) & (n_n3520) & (n_n4456) & (!n_n4458) & (!x55x)) + ((n_n4455) & (n_n3520) & (n_n4456) & (!n_n4458) & (x55x)) + ((n_n4455) & (n_n3520) & (n_n4456) & (n_n4458) & (!x55x)) + ((n_n4455) & (n_n3520) & (n_n4456) & (n_n4458) & (x55x)));
	assign x13615x = (((!x13592x) & (!x13593x) & (!x13599x) & (x13600x)) + ((!x13592x) & (!x13593x) & (x13599x) & (!x13600x)) + ((!x13592x) & (!x13593x) & (x13599x) & (x13600x)) + ((!x13592x) & (x13593x) & (!x13599x) & (!x13600x)) + ((!x13592x) & (x13593x) & (!x13599x) & (x13600x)) + ((!x13592x) & (x13593x) & (x13599x) & (!x13600x)) + ((!x13592x) & (x13593x) & (x13599x) & (x13600x)) + ((x13592x) & (!x13593x) & (!x13599x) & (!x13600x)) + ((x13592x) & (!x13593x) & (!x13599x) & (x13600x)) + ((x13592x) & (!x13593x) & (x13599x) & (!x13600x)) + ((x13592x) & (!x13593x) & (x13599x) & (x13600x)) + ((x13592x) & (x13593x) & (!x13599x) & (!x13600x)) + ((x13592x) & (x13593x) & (!x13599x) & (x13600x)) + ((x13592x) & (x13593x) & (x13599x) & (!x13600x)) + ((x13592x) & (x13593x) & (x13599x) & (x13600x)));
	assign x13681x = (((!x13623x) & (!x13624x) & (!x13672x) & (!x13673x) & (n_n3937)) + ((!x13623x) & (!x13624x) & (!x13672x) & (x13673x) & (!n_n3937)) + ((!x13623x) & (!x13624x) & (!x13672x) & (x13673x) & (n_n3937)) + ((!x13623x) & (!x13624x) & (x13672x) & (!x13673x) & (!n_n3937)) + ((!x13623x) & (!x13624x) & (x13672x) & (!x13673x) & (n_n3937)) + ((!x13623x) & (!x13624x) & (x13672x) & (x13673x) & (!n_n3937)) + ((!x13623x) & (!x13624x) & (x13672x) & (x13673x) & (n_n3937)) + ((!x13623x) & (x13624x) & (!x13672x) & (!x13673x) & (!n_n3937)) + ((!x13623x) & (x13624x) & (!x13672x) & (!x13673x) & (n_n3937)) + ((!x13623x) & (x13624x) & (!x13672x) & (x13673x) & (!n_n3937)) + ((!x13623x) & (x13624x) & (!x13672x) & (x13673x) & (n_n3937)) + ((!x13623x) & (x13624x) & (x13672x) & (!x13673x) & (!n_n3937)) + ((!x13623x) & (x13624x) & (x13672x) & (!x13673x) & (n_n3937)) + ((!x13623x) & (x13624x) & (x13672x) & (x13673x) & (!n_n3937)) + ((!x13623x) & (x13624x) & (x13672x) & (x13673x) & (n_n3937)) + ((x13623x) & (!x13624x) & (!x13672x) & (!x13673x) & (!n_n3937)) + ((x13623x) & (!x13624x) & (!x13672x) & (!x13673x) & (n_n3937)) + ((x13623x) & (!x13624x) & (!x13672x) & (x13673x) & (!n_n3937)) + ((x13623x) & (!x13624x) & (!x13672x) & (x13673x) & (n_n3937)) + ((x13623x) & (!x13624x) & (x13672x) & (!x13673x) & (!n_n3937)) + ((x13623x) & (!x13624x) & (x13672x) & (!x13673x) & (n_n3937)) + ((x13623x) & (!x13624x) & (x13672x) & (x13673x) & (!n_n3937)) + ((x13623x) & (!x13624x) & (x13672x) & (x13673x) & (n_n3937)) + ((x13623x) & (x13624x) & (!x13672x) & (!x13673x) & (!n_n3937)) + ((x13623x) & (x13624x) & (!x13672x) & (!x13673x) & (n_n3937)) + ((x13623x) & (x13624x) & (!x13672x) & (x13673x) & (!n_n3937)) + ((x13623x) & (x13624x) & (!x13672x) & (x13673x) & (n_n3937)) + ((x13623x) & (x13624x) & (x13672x) & (!x13673x) & (!n_n3937)) + ((x13623x) & (x13624x) & (x13672x) & (!x13673x) & (n_n3937)) + ((x13623x) & (x13624x) & (x13672x) & (x13673x) & (!n_n3937)) + ((x13623x) & (x13624x) & (x13672x) & (x13673x) & (n_n3937)));
	assign x13727x = (((!n_n4996) & (!n_n4987) & (!n_n5006) & (!n_n5033) & (n_n5051)) + ((!n_n4996) & (!n_n4987) & (!n_n5006) & (n_n5033) & (!n_n5051)) + ((!n_n4996) & (!n_n4987) & (!n_n5006) & (n_n5033) & (n_n5051)) + ((!n_n4996) & (!n_n4987) & (n_n5006) & (!n_n5033) & (!n_n5051)) + ((!n_n4996) & (!n_n4987) & (n_n5006) & (!n_n5033) & (n_n5051)) + ((!n_n4996) & (!n_n4987) & (n_n5006) & (n_n5033) & (!n_n5051)) + ((!n_n4996) & (!n_n4987) & (n_n5006) & (n_n5033) & (n_n5051)) + ((!n_n4996) & (n_n4987) & (!n_n5006) & (!n_n5033) & (!n_n5051)) + ((!n_n4996) & (n_n4987) & (!n_n5006) & (!n_n5033) & (n_n5051)) + ((!n_n4996) & (n_n4987) & (!n_n5006) & (n_n5033) & (!n_n5051)) + ((!n_n4996) & (n_n4987) & (!n_n5006) & (n_n5033) & (n_n5051)) + ((!n_n4996) & (n_n4987) & (n_n5006) & (!n_n5033) & (!n_n5051)) + ((!n_n4996) & (n_n4987) & (n_n5006) & (!n_n5033) & (n_n5051)) + ((!n_n4996) & (n_n4987) & (n_n5006) & (n_n5033) & (!n_n5051)) + ((!n_n4996) & (n_n4987) & (n_n5006) & (n_n5033) & (n_n5051)) + ((n_n4996) & (!n_n4987) & (!n_n5006) & (!n_n5033) & (!n_n5051)) + ((n_n4996) & (!n_n4987) & (!n_n5006) & (!n_n5033) & (n_n5051)) + ((n_n4996) & (!n_n4987) & (!n_n5006) & (n_n5033) & (!n_n5051)) + ((n_n4996) & (!n_n4987) & (!n_n5006) & (n_n5033) & (n_n5051)) + ((n_n4996) & (!n_n4987) & (n_n5006) & (!n_n5033) & (!n_n5051)) + ((n_n4996) & (!n_n4987) & (n_n5006) & (!n_n5033) & (n_n5051)) + ((n_n4996) & (!n_n4987) & (n_n5006) & (n_n5033) & (!n_n5051)) + ((n_n4996) & (!n_n4987) & (n_n5006) & (n_n5033) & (n_n5051)) + ((n_n4996) & (n_n4987) & (!n_n5006) & (!n_n5033) & (!n_n5051)) + ((n_n4996) & (n_n4987) & (!n_n5006) & (!n_n5033) & (n_n5051)) + ((n_n4996) & (n_n4987) & (!n_n5006) & (n_n5033) & (!n_n5051)) + ((n_n4996) & (n_n4987) & (!n_n5006) & (n_n5033) & (n_n5051)) + ((n_n4996) & (n_n4987) & (n_n5006) & (!n_n5033) & (!n_n5051)) + ((n_n4996) & (n_n4987) & (n_n5006) & (!n_n5033) & (n_n5051)) + ((n_n4996) & (n_n4987) & (n_n5006) & (n_n5033) & (!n_n5051)) + ((n_n4996) & (n_n4987) & (n_n5006) & (n_n5033) & (n_n5051)));
	assign x13728x = (((!n_n4994) & (!n_n5002) & (!n_n5056) & (!n_n5053) & (x13727x)) + ((!n_n4994) & (!n_n5002) & (!n_n5056) & (n_n5053) & (!x13727x)) + ((!n_n4994) & (!n_n5002) & (!n_n5056) & (n_n5053) & (x13727x)) + ((!n_n4994) & (!n_n5002) & (n_n5056) & (!n_n5053) & (!x13727x)) + ((!n_n4994) & (!n_n5002) & (n_n5056) & (!n_n5053) & (x13727x)) + ((!n_n4994) & (!n_n5002) & (n_n5056) & (n_n5053) & (!x13727x)) + ((!n_n4994) & (!n_n5002) & (n_n5056) & (n_n5053) & (x13727x)) + ((!n_n4994) & (n_n5002) & (!n_n5056) & (!n_n5053) & (!x13727x)) + ((!n_n4994) & (n_n5002) & (!n_n5056) & (!n_n5053) & (x13727x)) + ((!n_n4994) & (n_n5002) & (!n_n5056) & (n_n5053) & (!x13727x)) + ((!n_n4994) & (n_n5002) & (!n_n5056) & (n_n5053) & (x13727x)) + ((!n_n4994) & (n_n5002) & (n_n5056) & (!n_n5053) & (!x13727x)) + ((!n_n4994) & (n_n5002) & (n_n5056) & (!n_n5053) & (x13727x)) + ((!n_n4994) & (n_n5002) & (n_n5056) & (n_n5053) & (!x13727x)) + ((!n_n4994) & (n_n5002) & (n_n5056) & (n_n5053) & (x13727x)) + ((n_n4994) & (!n_n5002) & (!n_n5056) & (!n_n5053) & (!x13727x)) + ((n_n4994) & (!n_n5002) & (!n_n5056) & (!n_n5053) & (x13727x)) + ((n_n4994) & (!n_n5002) & (!n_n5056) & (n_n5053) & (!x13727x)) + ((n_n4994) & (!n_n5002) & (!n_n5056) & (n_n5053) & (x13727x)) + ((n_n4994) & (!n_n5002) & (n_n5056) & (!n_n5053) & (!x13727x)) + ((n_n4994) & (!n_n5002) & (n_n5056) & (!n_n5053) & (x13727x)) + ((n_n4994) & (!n_n5002) & (n_n5056) & (n_n5053) & (!x13727x)) + ((n_n4994) & (!n_n5002) & (n_n5056) & (n_n5053) & (x13727x)) + ((n_n4994) & (n_n5002) & (!n_n5056) & (!n_n5053) & (!x13727x)) + ((n_n4994) & (n_n5002) & (!n_n5056) & (!n_n5053) & (x13727x)) + ((n_n4994) & (n_n5002) & (!n_n5056) & (n_n5053) & (!x13727x)) + ((n_n4994) & (n_n5002) & (!n_n5056) & (n_n5053) & (x13727x)) + ((n_n4994) & (n_n5002) & (n_n5056) & (!n_n5053) & (!x13727x)) + ((n_n4994) & (n_n5002) & (n_n5056) & (!n_n5053) & (x13727x)) + ((n_n4994) & (n_n5002) & (n_n5056) & (n_n5053) & (!x13727x)) + ((n_n4994) & (n_n5002) & (n_n5056) & (n_n5053) & (x13727x)));
	assign x13729x = (((!x13696x) & (!x13697x) & (!x13719x) & (x13720x)) + ((!x13696x) & (!x13697x) & (x13719x) & (!x13720x)) + ((!x13696x) & (!x13697x) & (x13719x) & (x13720x)) + ((!x13696x) & (x13697x) & (!x13719x) & (!x13720x)) + ((!x13696x) & (x13697x) & (!x13719x) & (x13720x)) + ((!x13696x) & (x13697x) & (x13719x) & (!x13720x)) + ((!x13696x) & (x13697x) & (x13719x) & (x13720x)) + ((x13696x) & (!x13697x) & (!x13719x) & (!x13720x)) + ((x13696x) & (!x13697x) & (!x13719x) & (x13720x)) + ((x13696x) & (!x13697x) & (x13719x) & (!x13720x)) + ((x13696x) & (!x13697x) & (x13719x) & (x13720x)) + ((x13696x) & (x13697x) & (!x13719x) & (!x13720x)) + ((x13696x) & (x13697x) & (!x13719x) & (x13720x)) + ((x13696x) & (x13697x) & (x13719x) & (!x13720x)) + ((x13696x) & (x13697x) & (x13719x) & (x13720x)));
	assign x13973x = (((!x592x) & (!x24x) & (!x392x) & (!n_n5288) & (n_n5286)) + ((!x592x) & (!x24x) & (!x392x) & (n_n5288) & (!n_n5286)) + ((!x592x) & (!x24x) & (!x392x) & (n_n5288) & (n_n5286)) + ((!x592x) & (!x24x) & (x392x) & (!n_n5288) & (!n_n5286)) + ((!x592x) & (!x24x) & (x392x) & (!n_n5288) & (n_n5286)) + ((!x592x) & (!x24x) & (x392x) & (n_n5288) & (!n_n5286)) + ((!x592x) & (!x24x) & (x392x) & (n_n5288) & (n_n5286)) + ((!x592x) & (x24x) & (!x392x) & (!n_n5288) & (n_n5286)) + ((!x592x) & (x24x) & (!x392x) & (n_n5288) & (!n_n5286)) + ((!x592x) & (x24x) & (!x392x) & (n_n5288) & (n_n5286)) + ((!x592x) & (x24x) & (x392x) & (!n_n5288) & (!n_n5286)) + ((!x592x) & (x24x) & (x392x) & (!n_n5288) & (n_n5286)) + ((!x592x) & (x24x) & (x392x) & (n_n5288) & (!n_n5286)) + ((!x592x) & (x24x) & (x392x) & (n_n5288) & (n_n5286)) + ((x592x) & (!x24x) & (!x392x) & (!n_n5288) & (n_n5286)) + ((x592x) & (!x24x) & (!x392x) & (n_n5288) & (!n_n5286)) + ((x592x) & (!x24x) & (!x392x) & (n_n5288) & (n_n5286)) + ((x592x) & (!x24x) & (x392x) & (!n_n5288) & (!n_n5286)) + ((x592x) & (!x24x) & (x392x) & (!n_n5288) & (n_n5286)) + ((x592x) & (!x24x) & (x392x) & (n_n5288) & (!n_n5286)) + ((x592x) & (!x24x) & (x392x) & (n_n5288) & (n_n5286)) + ((x592x) & (x24x) & (!x392x) & (!n_n5288) & (!n_n5286)) + ((x592x) & (x24x) & (!x392x) & (!n_n5288) & (n_n5286)) + ((x592x) & (x24x) & (!x392x) & (n_n5288) & (!n_n5286)) + ((x592x) & (x24x) & (!x392x) & (n_n5288) & (n_n5286)) + ((x592x) & (x24x) & (x392x) & (!n_n5288) & (!n_n5286)) + ((x592x) & (x24x) & (x392x) & (!n_n5288) & (n_n5286)) + ((x592x) & (x24x) & (x392x) & (n_n5288) & (!n_n5286)) + ((x592x) & (x24x) & (x392x) & (n_n5288) & (n_n5286)));
	assign x14021x = (((!x11x) & (!n_n195) & (!n_n500) & (!n_n3427) & (n_n5008)) + ((!x11x) & (!n_n195) & (!n_n500) & (n_n3427) & (!n_n5008)) + ((!x11x) & (!n_n195) & (!n_n500) & (n_n3427) & (n_n5008)) + ((!x11x) & (!n_n195) & (n_n500) & (!n_n3427) & (n_n5008)) + ((!x11x) & (!n_n195) & (n_n500) & (n_n3427) & (!n_n5008)) + ((!x11x) & (!n_n195) & (n_n500) & (n_n3427) & (n_n5008)) + ((!x11x) & (n_n195) & (!n_n500) & (!n_n3427) & (n_n5008)) + ((!x11x) & (n_n195) & (!n_n500) & (n_n3427) & (!n_n5008)) + ((!x11x) & (n_n195) & (!n_n500) & (n_n3427) & (n_n5008)) + ((!x11x) & (n_n195) & (n_n500) & (!n_n3427) & (n_n5008)) + ((!x11x) & (n_n195) & (n_n500) & (n_n3427) & (!n_n5008)) + ((!x11x) & (n_n195) & (n_n500) & (n_n3427) & (n_n5008)) + ((x11x) & (!n_n195) & (!n_n500) & (!n_n3427) & (n_n5008)) + ((x11x) & (!n_n195) & (!n_n500) & (n_n3427) & (!n_n5008)) + ((x11x) & (!n_n195) & (!n_n500) & (n_n3427) & (n_n5008)) + ((x11x) & (!n_n195) & (n_n500) & (!n_n3427) & (n_n5008)) + ((x11x) & (!n_n195) & (n_n500) & (n_n3427) & (!n_n5008)) + ((x11x) & (!n_n195) & (n_n500) & (n_n3427) & (n_n5008)) + ((x11x) & (n_n195) & (!n_n500) & (!n_n3427) & (n_n5008)) + ((x11x) & (n_n195) & (!n_n500) & (n_n3427) & (!n_n5008)) + ((x11x) & (n_n195) & (!n_n500) & (n_n3427) & (n_n5008)) + ((x11x) & (n_n195) & (n_n500) & (!n_n3427) & (!n_n5008)) + ((x11x) & (n_n195) & (n_n500) & (!n_n3427) & (n_n5008)) + ((x11x) & (n_n195) & (n_n500) & (n_n3427) & (!n_n5008)) + ((x11x) & (n_n195) & (n_n500) & (n_n3427) & (n_n5008)));
	assign x14054x = (((!i_7_) & (i_8_) & (i_6_) & (x12x) & (n_n464)) + ((i_7_) & (!i_8_) & (i_6_) & (x12x) & (n_n464)) + ((i_7_) & (i_8_) & (i_6_) & (x12x) & (n_n464)));
	assign x14059x = (((!n_n524) & (n_n532) & (n_n491) & (x12x) & (!n_n500)) + ((!n_n524) & (n_n532) & (n_n491) & (x12x) & (n_n500)) + ((n_n524) & (!n_n532) & (!n_n491) & (x12x) & (n_n500)) + ((n_n524) & (!n_n532) & (n_n491) & (x12x) & (n_n500)) + ((n_n524) & (n_n532) & (!n_n491) & (x12x) & (n_n500)) + ((n_n524) & (n_n532) & (n_n491) & (x12x) & (!n_n500)) + ((n_n524) & (n_n532) & (n_n491) & (x12x) & (n_n500)));
	assign x14063x = (((!n_n3771) & (!n_n5144) & (!n_n5143) & (!x211x) & (x14059x)) + ((!n_n3771) & (!n_n5144) & (!n_n5143) & (x211x) & (!x14059x)) + ((!n_n3771) & (!n_n5144) & (!n_n5143) & (x211x) & (x14059x)) + ((!n_n3771) & (!n_n5144) & (n_n5143) & (!x211x) & (!x14059x)) + ((!n_n3771) & (!n_n5144) & (n_n5143) & (!x211x) & (x14059x)) + ((!n_n3771) & (!n_n5144) & (n_n5143) & (x211x) & (!x14059x)) + ((!n_n3771) & (!n_n5144) & (n_n5143) & (x211x) & (x14059x)) + ((!n_n3771) & (n_n5144) & (!n_n5143) & (!x211x) & (!x14059x)) + ((!n_n3771) & (n_n5144) & (!n_n5143) & (!x211x) & (x14059x)) + ((!n_n3771) & (n_n5144) & (!n_n5143) & (x211x) & (!x14059x)) + ((!n_n3771) & (n_n5144) & (!n_n5143) & (x211x) & (x14059x)) + ((!n_n3771) & (n_n5144) & (n_n5143) & (!x211x) & (!x14059x)) + ((!n_n3771) & (n_n5144) & (n_n5143) & (!x211x) & (x14059x)) + ((!n_n3771) & (n_n5144) & (n_n5143) & (x211x) & (!x14059x)) + ((!n_n3771) & (n_n5144) & (n_n5143) & (x211x) & (x14059x)) + ((n_n3771) & (!n_n5144) & (!n_n5143) & (!x211x) & (!x14059x)) + ((n_n3771) & (!n_n5144) & (!n_n5143) & (!x211x) & (x14059x)) + ((n_n3771) & (!n_n5144) & (!n_n5143) & (x211x) & (!x14059x)) + ((n_n3771) & (!n_n5144) & (!n_n5143) & (x211x) & (x14059x)) + ((n_n3771) & (!n_n5144) & (n_n5143) & (!x211x) & (!x14059x)) + ((n_n3771) & (!n_n5144) & (n_n5143) & (!x211x) & (x14059x)) + ((n_n3771) & (!n_n5144) & (n_n5143) & (x211x) & (!x14059x)) + ((n_n3771) & (!n_n5144) & (n_n5143) & (x211x) & (x14059x)) + ((n_n3771) & (n_n5144) & (!n_n5143) & (!x211x) & (!x14059x)) + ((n_n3771) & (n_n5144) & (!n_n5143) & (!x211x) & (x14059x)) + ((n_n3771) & (n_n5144) & (!n_n5143) & (x211x) & (!x14059x)) + ((n_n3771) & (n_n5144) & (!n_n5143) & (x211x) & (x14059x)) + ((n_n3771) & (n_n5144) & (n_n5143) & (!x211x) & (!x14059x)) + ((n_n3771) & (n_n5144) & (n_n5143) & (!x211x) & (x14059x)) + ((n_n3771) & (n_n5144) & (n_n5143) & (x211x) & (!x14059x)) + ((n_n3771) & (n_n5144) & (n_n5143) & (x211x) & (x14059x)));
	assign x14143x = (((!n_n4420) & (!n_n4430) & (x84x)) + ((!n_n4420) & (n_n4430) & (!x84x)) + ((!n_n4420) & (n_n4430) & (x84x)) + ((n_n4420) & (!n_n4430) & (!x84x)) + ((n_n4420) & (!n_n4430) & (x84x)) + ((n_n4420) & (n_n4430) & (!x84x)) + ((n_n4420) & (n_n4430) & (x84x)));
	assign x22112x = (((!n_n4338) & (!n_n4337) & (!n_n4345) & (!n_n4341)));
	assign x14218x = (((!x13689x) & (!x13690x) & (!x13735x) & (x13736x)) + ((!x13689x) & (!x13690x) & (x13735x) & (!x13736x)) + ((!x13689x) & (!x13690x) & (x13735x) & (x13736x)) + ((!x13689x) & (x13690x) & (!x13735x) & (!x13736x)) + ((!x13689x) & (x13690x) & (!x13735x) & (x13736x)) + ((!x13689x) & (x13690x) & (x13735x) & (!x13736x)) + ((!x13689x) & (x13690x) & (x13735x) & (x13736x)) + ((x13689x) & (!x13690x) & (!x13735x) & (!x13736x)) + ((x13689x) & (!x13690x) & (!x13735x) & (x13736x)) + ((x13689x) & (!x13690x) & (x13735x) & (!x13736x)) + ((x13689x) & (!x13690x) & (x13735x) & (x13736x)) + ((x13689x) & (x13690x) & (!x13735x) & (!x13736x)) + ((x13689x) & (x13690x) & (!x13735x) & (x13736x)) + ((x13689x) & (x13690x) & (x13735x) & (!x13736x)) + ((x13689x) & (x13690x) & (x13735x) & (x13736x)));
	assign x14273x = (((!n_n5034) & (!n_n4996) & (!n_n5026) & (n_n4988)) + ((!n_n5034) & (!n_n4996) & (n_n5026) & (!n_n4988)) + ((!n_n5034) & (!n_n4996) & (n_n5026) & (n_n4988)) + ((!n_n5034) & (n_n4996) & (!n_n5026) & (!n_n4988)) + ((!n_n5034) & (n_n4996) & (!n_n5026) & (n_n4988)) + ((!n_n5034) & (n_n4996) & (n_n5026) & (!n_n4988)) + ((!n_n5034) & (n_n4996) & (n_n5026) & (n_n4988)) + ((n_n5034) & (!n_n4996) & (!n_n5026) & (!n_n4988)) + ((n_n5034) & (!n_n4996) & (!n_n5026) & (n_n4988)) + ((n_n5034) & (!n_n4996) & (n_n5026) & (!n_n4988)) + ((n_n5034) & (!n_n4996) & (n_n5026) & (n_n4988)) + ((n_n5034) & (n_n4996) & (!n_n5026) & (!n_n4988)) + ((n_n5034) & (n_n4996) & (!n_n5026) & (n_n4988)) + ((n_n5034) & (n_n4996) & (n_n5026) & (!n_n4988)) + ((n_n5034) & (n_n4996) & (n_n5026) & (n_n4988)));
	assign x14338x = (((!x37x) & (!n_n4399) & (!n_n4409) & (n_n4370)) + ((!x37x) & (!n_n4399) & (n_n4409) & (!n_n4370)) + ((!x37x) & (!n_n4399) & (n_n4409) & (n_n4370)) + ((!x37x) & (n_n4399) & (!n_n4409) & (!n_n4370)) + ((!x37x) & (n_n4399) & (!n_n4409) & (n_n4370)) + ((!x37x) & (n_n4399) & (n_n4409) & (!n_n4370)) + ((!x37x) & (n_n4399) & (n_n4409) & (n_n4370)) + ((x37x) & (!n_n4399) & (!n_n4409) & (!n_n4370)) + ((x37x) & (!n_n4399) & (!n_n4409) & (n_n4370)) + ((x37x) & (!n_n4399) & (n_n4409) & (!n_n4370)) + ((x37x) & (!n_n4399) & (n_n4409) & (n_n4370)) + ((x37x) & (n_n4399) & (!n_n4409) & (!n_n4370)) + ((x37x) & (n_n4399) & (!n_n4409) & (n_n4370)) + ((x37x) & (n_n4399) & (n_n4409) & (!n_n4370)) + ((x37x) & (n_n4399) & (n_n4409) & (n_n4370)));
	assign x14339x = (((!n_n4406) & (!n_n4364) & (!n_n4374) & (!n_n4408) & (x14338x)) + ((!n_n4406) & (!n_n4364) & (!n_n4374) & (n_n4408) & (!x14338x)) + ((!n_n4406) & (!n_n4364) & (!n_n4374) & (n_n4408) & (x14338x)) + ((!n_n4406) & (!n_n4364) & (n_n4374) & (!n_n4408) & (!x14338x)) + ((!n_n4406) & (!n_n4364) & (n_n4374) & (!n_n4408) & (x14338x)) + ((!n_n4406) & (!n_n4364) & (n_n4374) & (n_n4408) & (!x14338x)) + ((!n_n4406) & (!n_n4364) & (n_n4374) & (n_n4408) & (x14338x)) + ((!n_n4406) & (n_n4364) & (!n_n4374) & (!n_n4408) & (!x14338x)) + ((!n_n4406) & (n_n4364) & (!n_n4374) & (!n_n4408) & (x14338x)) + ((!n_n4406) & (n_n4364) & (!n_n4374) & (n_n4408) & (!x14338x)) + ((!n_n4406) & (n_n4364) & (!n_n4374) & (n_n4408) & (x14338x)) + ((!n_n4406) & (n_n4364) & (n_n4374) & (!n_n4408) & (!x14338x)) + ((!n_n4406) & (n_n4364) & (n_n4374) & (!n_n4408) & (x14338x)) + ((!n_n4406) & (n_n4364) & (n_n4374) & (n_n4408) & (!x14338x)) + ((!n_n4406) & (n_n4364) & (n_n4374) & (n_n4408) & (x14338x)) + ((n_n4406) & (!n_n4364) & (!n_n4374) & (!n_n4408) & (!x14338x)) + ((n_n4406) & (!n_n4364) & (!n_n4374) & (!n_n4408) & (x14338x)) + ((n_n4406) & (!n_n4364) & (!n_n4374) & (n_n4408) & (!x14338x)) + ((n_n4406) & (!n_n4364) & (!n_n4374) & (n_n4408) & (x14338x)) + ((n_n4406) & (!n_n4364) & (n_n4374) & (!n_n4408) & (!x14338x)) + ((n_n4406) & (!n_n4364) & (n_n4374) & (!n_n4408) & (x14338x)) + ((n_n4406) & (!n_n4364) & (n_n4374) & (n_n4408) & (!x14338x)) + ((n_n4406) & (!n_n4364) & (n_n4374) & (n_n4408) & (x14338x)) + ((n_n4406) & (n_n4364) & (!n_n4374) & (!n_n4408) & (!x14338x)) + ((n_n4406) & (n_n4364) & (!n_n4374) & (!n_n4408) & (x14338x)) + ((n_n4406) & (n_n4364) & (!n_n4374) & (n_n4408) & (!x14338x)) + ((n_n4406) & (n_n4364) & (!n_n4374) & (n_n4408) & (x14338x)) + ((n_n4406) & (n_n4364) & (n_n4374) & (!n_n4408) & (!x14338x)) + ((n_n4406) & (n_n4364) & (n_n4374) & (!n_n4408) & (x14338x)) + ((n_n4406) & (n_n4364) & (n_n4374) & (n_n4408) & (!x14338x)) + ((n_n4406) & (n_n4364) & (n_n4374) & (n_n4408) & (x14338x)));
	assign x14382x = (((!i_9_) & (!n_n524) & (n_n325) & (n_n500) & (n_n530)) + ((!i_9_) & (n_n524) & (n_n325) & (n_n500) & (n_n530)) + ((i_9_) & (n_n524) & (n_n325) & (n_n500) & (!n_n530)) + ((i_9_) & (n_n524) & (n_n325) & (n_n500) & (n_n530)));
	assign x22168x = (((!n_n4607) & (!n_n4612) & (!n_n4606) & (!n_n4611)));
	assign x14485x = (((!i_9_) & (n_n536) & (!n_n532) & (n_n534) & (n_n509)) + ((!i_9_) & (n_n536) & (n_n532) & (!n_n534) & (n_n509)) + ((!i_9_) & (n_n536) & (n_n532) & (n_n534) & (n_n509)) + ((i_9_) & (n_n536) & (!n_n532) & (n_n534) & (n_n509)) + ((i_9_) & (n_n536) & (n_n532) & (!n_n534) & (n_n509)) + ((i_9_) & (n_n536) & (n_n532) & (n_n534) & (n_n509)));
	assign x14504x = (((!i_9_) & (n_n536) & (!n_n524) & (n_n526) & (n_n482)) + ((!i_9_) & (n_n536) & (n_n524) & (!n_n526) & (n_n482)) + ((!i_9_) & (n_n536) & (n_n524) & (n_n526) & (n_n482)) + ((i_9_) & (n_n536) & (n_n524) & (!n_n526) & (n_n482)) + ((i_9_) & (n_n536) & (n_n524) & (n_n526) & (n_n482)));
	assign x14527x = (((!i_7_) & (!i_8_) & (i_6_) & (x13x) & (n_n535)) + ((i_7_) & (!i_8_) & (!i_6_) & (x13x) & (n_n535)) + ((i_7_) & (i_8_) & (i_6_) & (x13x) & (n_n535)));
	assign x14535x = (((!n_n4468) & (!n_n4471) & (!n_n4472) & (!n_n4474) & (n_n4465)) + ((!n_n4468) & (!n_n4471) & (!n_n4472) & (n_n4474) & (!n_n4465)) + ((!n_n4468) & (!n_n4471) & (!n_n4472) & (n_n4474) & (n_n4465)) + ((!n_n4468) & (!n_n4471) & (n_n4472) & (!n_n4474) & (!n_n4465)) + ((!n_n4468) & (!n_n4471) & (n_n4472) & (!n_n4474) & (n_n4465)) + ((!n_n4468) & (!n_n4471) & (n_n4472) & (n_n4474) & (!n_n4465)) + ((!n_n4468) & (!n_n4471) & (n_n4472) & (n_n4474) & (n_n4465)) + ((!n_n4468) & (n_n4471) & (!n_n4472) & (!n_n4474) & (!n_n4465)) + ((!n_n4468) & (n_n4471) & (!n_n4472) & (!n_n4474) & (n_n4465)) + ((!n_n4468) & (n_n4471) & (!n_n4472) & (n_n4474) & (!n_n4465)) + ((!n_n4468) & (n_n4471) & (!n_n4472) & (n_n4474) & (n_n4465)) + ((!n_n4468) & (n_n4471) & (n_n4472) & (!n_n4474) & (!n_n4465)) + ((!n_n4468) & (n_n4471) & (n_n4472) & (!n_n4474) & (n_n4465)) + ((!n_n4468) & (n_n4471) & (n_n4472) & (n_n4474) & (!n_n4465)) + ((!n_n4468) & (n_n4471) & (n_n4472) & (n_n4474) & (n_n4465)) + ((n_n4468) & (!n_n4471) & (!n_n4472) & (!n_n4474) & (!n_n4465)) + ((n_n4468) & (!n_n4471) & (!n_n4472) & (!n_n4474) & (n_n4465)) + ((n_n4468) & (!n_n4471) & (!n_n4472) & (n_n4474) & (!n_n4465)) + ((n_n4468) & (!n_n4471) & (!n_n4472) & (n_n4474) & (n_n4465)) + ((n_n4468) & (!n_n4471) & (n_n4472) & (!n_n4474) & (!n_n4465)) + ((n_n4468) & (!n_n4471) & (n_n4472) & (!n_n4474) & (n_n4465)) + ((n_n4468) & (!n_n4471) & (n_n4472) & (n_n4474) & (!n_n4465)) + ((n_n4468) & (!n_n4471) & (n_n4472) & (n_n4474) & (n_n4465)) + ((n_n4468) & (n_n4471) & (!n_n4472) & (!n_n4474) & (!n_n4465)) + ((n_n4468) & (n_n4471) & (!n_n4472) & (!n_n4474) & (n_n4465)) + ((n_n4468) & (n_n4471) & (!n_n4472) & (n_n4474) & (!n_n4465)) + ((n_n4468) & (n_n4471) & (!n_n4472) & (n_n4474) & (n_n4465)) + ((n_n4468) & (n_n4471) & (n_n4472) & (!n_n4474) & (!n_n4465)) + ((n_n4468) & (n_n4471) & (n_n4472) & (!n_n4474) & (n_n4465)) + ((n_n4468) & (n_n4471) & (n_n4472) & (n_n4474) & (!n_n4465)) + ((n_n4468) & (n_n4471) & (n_n4472) & (n_n4474) & (n_n4465)));
	assign x22107x = (((!x592x) & (!n_n5284) & (!x24x) & (!n_n5281) & (!n_n5288)) + ((!x592x) & (!n_n5284) & (x24x) & (!n_n5281) & (!n_n5288)) + ((x592x) & (!n_n5284) & (!x24x) & (!n_n5281) & (!n_n5288)));
	assign x14635x = (((!n_n5179) & (!n_n5178) & (!n_n5175) & (!n_n5177) & (n_n5170)) + ((!n_n5179) & (!n_n5178) & (!n_n5175) & (n_n5177) & (!n_n5170)) + ((!n_n5179) & (!n_n5178) & (!n_n5175) & (n_n5177) & (n_n5170)) + ((!n_n5179) & (!n_n5178) & (n_n5175) & (!n_n5177) & (!n_n5170)) + ((!n_n5179) & (!n_n5178) & (n_n5175) & (!n_n5177) & (n_n5170)) + ((!n_n5179) & (!n_n5178) & (n_n5175) & (n_n5177) & (!n_n5170)) + ((!n_n5179) & (!n_n5178) & (n_n5175) & (n_n5177) & (n_n5170)) + ((!n_n5179) & (n_n5178) & (!n_n5175) & (!n_n5177) & (!n_n5170)) + ((!n_n5179) & (n_n5178) & (!n_n5175) & (!n_n5177) & (n_n5170)) + ((!n_n5179) & (n_n5178) & (!n_n5175) & (n_n5177) & (!n_n5170)) + ((!n_n5179) & (n_n5178) & (!n_n5175) & (n_n5177) & (n_n5170)) + ((!n_n5179) & (n_n5178) & (n_n5175) & (!n_n5177) & (!n_n5170)) + ((!n_n5179) & (n_n5178) & (n_n5175) & (!n_n5177) & (n_n5170)) + ((!n_n5179) & (n_n5178) & (n_n5175) & (n_n5177) & (!n_n5170)) + ((!n_n5179) & (n_n5178) & (n_n5175) & (n_n5177) & (n_n5170)) + ((n_n5179) & (!n_n5178) & (!n_n5175) & (!n_n5177) & (!n_n5170)) + ((n_n5179) & (!n_n5178) & (!n_n5175) & (!n_n5177) & (n_n5170)) + ((n_n5179) & (!n_n5178) & (!n_n5175) & (n_n5177) & (!n_n5170)) + ((n_n5179) & (!n_n5178) & (!n_n5175) & (n_n5177) & (n_n5170)) + ((n_n5179) & (!n_n5178) & (n_n5175) & (!n_n5177) & (!n_n5170)) + ((n_n5179) & (!n_n5178) & (n_n5175) & (!n_n5177) & (n_n5170)) + ((n_n5179) & (!n_n5178) & (n_n5175) & (n_n5177) & (!n_n5170)) + ((n_n5179) & (!n_n5178) & (n_n5175) & (n_n5177) & (n_n5170)) + ((n_n5179) & (n_n5178) & (!n_n5175) & (!n_n5177) & (!n_n5170)) + ((n_n5179) & (n_n5178) & (!n_n5175) & (!n_n5177) & (n_n5170)) + ((n_n5179) & (n_n5178) & (!n_n5175) & (n_n5177) & (!n_n5170)) + ((n_n5179) & (n_n5178) & (!n_n5175) & (n_n5177) & (n_n5170)) + ((n_n5179) & (n_n5178) & (n_n5175) & (!n_n5177) & (!n_n5170)) + ((n_n5179) & (n_n5178) & (n_n5175) & (!n_n5177) & (n_n5170)) + ((n_n5179) & (n_n5178) & (n_n5175) & (n_n5177) & (!n_n5170)) + ((n_n5179) & (n_n5178) & (n_n5175) & (n_n5177) & (n_n5170)));
	assign x14681x = (((!n_n5021) & (!n_n5010) & (!n_n5012) & (!n_n5011) & (n_n5013)) + ((!n_n5021) & (!n_n5010) & (!n_n5012) & (n_n5011) & (!n_n5013)) + ((!n_n5021) & (!n_n5010) & (!n_n5012) & (n_n5011) & (n_n5013)) + ((!n_n5021) & (!n_n5010) & (n_n5012) & (!n_n5011) & (!n_n5013)) + ((!n_n5021) & (!n_n5010) & (n_n5012) & (!n_n5011) & (n_n5013)) + ((!n_n5021) & (!n_n5010) & (n_n5012) & (n_n5011) & (!n_n5013)) + ((!n_n5021) & (!n_n5010) & (n_n5012) & (n_n5011) & (n_n5013)) + ((!n_n5021) & (n_n5010) & (!n_n5012) & (!n_n5011) & (!n_n5013)) + ((!n_n5021) & (n_n5010) & (!n_n5012) & (!n_n5011) & (n_n5013)) + ((!n_n5021) & (n_n5010) & (!n_n5012) & (n_n5011) & (!n_n5013)) + ((!n_n5021) & (n_n5010) & (!n_n5012) & (n_n5011) & (n_n5013)) + ((!n_n5021) & (n_n5010) & (n_n5012) & (!n_n5011) & (!n_n5013)) + ((!n_n5021) & (n_n5010) & (n_n5012) & (!n_n5011) & (n_n5013)) + ((!n_n5021) & (n_n5010) & (n_n5012) & (n_n5011) & (!n_n5013)) + ((!n_n5021) & (n_n5010) & (n_n5012) & (n_n5011) & (n_n5013)) + ((n_n5021) & (!n_n5010) & (!n_n5012) & (!n_n5011) & (!n_n5013)) + ((n_n5021) & (!n_n5010) & (!n_n5012) & (!n_n5011) & (n_n5013)) + ((n_n5021) & (!n_n5010) & (!n_n5012) & (n_n5011) & (!n_n5013)) + ((n_n5021) & (!n_n5010) & (!n_n5012) & (n_n5011) & (n_n5013)) + ((n_n5021) & (!n_n5010) & (n_n5012) & (!n_n5011) & (!n_n5013)) + ((n_n5021) & (!n_n5010) & (n_n5012) & (!n_n5011) & (n_n5013)) + ((n_n5021) & (!n_n5010) & (n_n5012) & (n_n5011) & (!n_n5013)) + ((n_n5021) & (!n_n5010) & (n_n5012) & (n_n5011) & (n_n5013)) + ((n_n5021) & (n_n5010) & (!n_n5012) & (!n_n5011) & (!n_n5013)) + ((n_n5021) & (n_n5010) & (!n_n5012) & (!n_n5011) & (n_n5013)) + ((n_n5021) & (n_n5010) & (!n_n5012) & (n_n5011) & (!n_n5013)) + ((n_n5021) & (n_n5010) & (!n_n5012) & (n_n5011) & (n_n5013)) + ((n_n5021) & (n_n5010) & (n_n5012) & (!n_n5011) & (!n_n5013)) + ((n_n5021) & (n_n5010) & (n_n5012) & (!n_n5011) & (n_n5013)) + ((n_n5021) & (n_n5010) & (n_n5012) & (n_n5011) & (!n_n5013)) + ((n_n5021) & (n_n5010) & (n_n5012) & (n_n5011) & (n_n5013)));
	assign x14718x = (((!i_9_) & (!n_n526) & (!n_n482) & (!n_n325) & (x313x)) + ((!i_9_) & (!n_n526) & (!n_n482) & (n_n325) & (x313x)) + ((!i_9_) & (!n_n526) & (n_n482) & (!n_n325) & (x313x)) + ((!i_9_) & (!n_n526) & (n_n482) & (n_n325) & (x313x)) + ((!i_9_) & (n_n526) & (!n_n482) & (!n_n325) & (x313x)) + ((!i_9_) & (n_n526) & (!n_n482) & (n_n325) & (x313x)) + ((!i_9_) & (n_n526) & (n_n482) & (!n_n325) & (x313x)) + ((!i_9_) & (n_n526) & (n_n482) & (n_n325) & (!x313x)) + ((!i_9_) & (n_n526) & (n_n482) & (n_n325) & (x313x)) + ((i_9_) & (!n_n526) & (!n_n482) & (!n_n325) & (x313x)) + ((i_9_) & (!n_n526) & (!n_n482) & (n_n325) & (x313x)) + ((i_9_) & (!n_n526) & (n_n482) & (!n_n325) & (x313x)) + ((i_9_) & (!n_n526) & (n_n482) & (n_n325) & (x313x)) + ((i_9_) & (n_n526) & (!n_n482) & (!n_n325) & (x313x)) + ((i_9_) & (n_n526) & (!n_n482) & (n_n325) & (x313x)) + ((i_9_) & (n_n526) & (n_n482) & (!n_n325) & (x313x)) + ((i_9_) & (n_n526) & (n_n482) & (n_n325) & (x313x)));
	assign x14727x = (((!n_n532) & (!n_n509) & (!x17x) & (!n_n4853) & (n_n2727)) + ((!n_n532) & (!n_n509) & (!x17x) & (n_n4853) & (!n_n2727)) + ((!n_n532) & (!n_n509) & (!x17x) & (n_n4853) & (n_n2727)) + ((!n_n532) & (!n_n509) & (x17x) & (!n_n4853) & (n_n2727)) + ((!n_n532) & (!n_n509) & (x17x) & (n_n4853) & (!n_n2727)) + ((!n_n532) & (!n_n509) & (x17x) & (n_n4853) & (n_n2727)) + ((!n_n532) & (n_n509) & (!x17x) & (!n_n4853) & (n_n2727)) + ((!n_n532) & (n_n509) & (!x17x) & (n_n4853) & (!n_n2727)) + ((!n_n532) & (n_n509) & (!x17x) & (n_n4853) & (n_n2727)) + ((!n_n532) & (n_n509) & (x17x) & (!n_n4853) & (n_n2727)) + ((!n_n532) & (n_n509) & (x17x) & (n_n4853) & (!n_n2727)) + ((!n_n532) & (n_n509) & (x17x) & (n_n4853) & (n_n2727)) + ((n_n532) & (!n_n509) & (!x17x) & (!n_n4853) & (n_n2727)) + ((n_n532) & (!n_n509) & (!x17x) & (n_n4853) & (!n_n2727)) + ((n_n532) & (!n_n509) & (!x17x) & (n_n4853) & (n_n2727)) + ((n_n532) & (!n_n509) & (x17x) & (!n_n4853) & (n_n2727)) + ((n_n532) & (!n_n509) & (x17x) & (n_n4853) & (!n_n2727)) + ((n_n532) & (!n_n509) & (x17x) & (n_n4853) & (n_n2727)) + ((n_n532) & (n_n509) & (!x17x) & (!n_n4853) & (n_n2727)) + ((n_n532) & (n_n509) & (!x17x) & (n_n4853) & (!n_n2727)) + ((n_n532) & (n_n509) & (!x17x) & (n_n4853) & (n_n2727)) + ((n_n532) & (n_n509) & (x17x) & (!n_n4853) & (!n_n2727)) + ((n_n532) & (n_n509) & (x17x) & (!n_n4853) & (n_n2727)) + ((n_n532) & (n_n509) & (x17x) & (n_n4853) & (!n_n2727)) + ((n_n532) & (n_n509) & (x17x) & (n_n4853) & (n_n2727)));
	assign x14761x = (((!n_n4976) & (!n_n4977) & (!n_n4981) & (n_n4987)) + ((!n_n4976) & (!n_n4977) & (n_n4981) & (!n_n4987)) + ((!n_n4976) & (!n_n4977) & (n_n4981) & (n_n4987)) + ((!n_n4976) & (n_n4977) & (!n_n4981) & (!n_n4987)) + ((!n_n4976) & (n_n4977) & (!n_n4981) & (n_n4987)) + ((!n_n4976) & (n_n4977) & (n_n4981) & (!n_n4987)) + ((!n_n4976) & (n_n4977) & (n_n4981) & (n_n4987)) + ((n_n4976) & (!n_n4977) & (!n_n4981) & (!n_n4987)) + ((n_n4976) & (!n_n4977) & (!n_n4981) & (n_n4987)) + ((n_n4976) & (!n_n4977) & (n_n4981) & (!n_n4987)) + ((n_n4976) & (!n_n4977) & (n_n4981) & (n_n4987)) + ((n_n4976) & (n_n4977) & (!n_n4981) & (!n_n4987)) + ((n_n4976) & (n_n4977) & (!n_n4981) & (n_n4987)) + ((n_n4976) & (n_n4977) & (n_n4981) & (!n_n4987)) + ((n_n4976) & (n_n4977) & (n_n4981) & (n_n4987)));
	assign x14769x = (((!x17x) & (!n_n522) & (!n_n500) & (!n_n4877) & (n_n3815)) + ((!x17x) & (!n_n522) & (!n_n500) & (n_n4877) & (!n_n3815)) + ((!x17x) & (!n_n522) & (!n_n500) & (n_n4877) & (n_n3815)) + ((!x17x) & (!n_n522) & (n_n500) & (!n_n4877) & (n_n3815)) + ((!x17x) & (!n_n522) & (n_n500) & (n_n4877) & (!n_n3815)) + ((!x17x) & (!n_n522) & (n_n500) & (n_n4877) & (n_n3815)) + ((!x17x) & (n_n522) & (!n_n500) & (!n_n4877) & (n_n3815)) + ((!x17x) & (n_n522) & (!n_n500) & (n_n4877) & (!n_n3815)) + ((!x17x) & (n_n522) & (!n_n500) & (n_n4877) & (n_n3815)) + ((!x17x) & (n_n522) & (n_n500) & (!n_n4877) & (n_n3815)) + ((!x17x) & (n_n522) & (n_n500) & (n_n4877) & (!n_n3815)) + ((!x17x) & (n_n522) & (n_n500) & (n_n4877) & (n_n3815)) + ((x17x) & (!n_n522) & (!n_n500) & (!n_n4877) & (n_n3815)) + ((x17x) & (!n_n522) & (!n_n500) & (n_n4877) & (!n_n3815)) + ((x17x) & (!n_n522) & (!n_n500) & (n_n4877) & (n_n3815)) + ((x17x) & (!n_n522) & (n_n500) & (!n_n4877) & (n_n3815)) + ((x17x) & (!n_n522) & (n_n500) & (n_n4877) & (!n_n3815)) + ((x17x) & (!n_n522) & (n_n500) & (n_n4877) & (n_n3815)) + ((x17x) & (n_n522) & (!n_n500) & (!n_n4877) & (n_n3815)) + ((x17x) & (n_n522) & (!n_n500) & (n_n4877) & (!n_n3815)) + ((x17x) & (n_n522) & (!n_n500) & (n_n4877) & (n_n3815)) + ((x17x) & (n_n522) & (n_n500) & (!n_n4877) & (!n_n3815)) + ((x17x) & (n_n522) & (n_n500) & (!n_n4877) & (n_n3815)) + ((x17x) & (n_n522) & (n_n500) & (n_n4877) & (!n_n3815)) + ((x17x) & (n_n522) & (n_n500) & (n_n4877) & (n_n3815)));
	assign x22190x = (((!n_n5330) & (!n_n5331) & (!n_n3708) & (!n_n3710) & (!x14357x)));
	assign x14846x = (((!x15x) & (!x583x) & (!n_n4557) & (!n_n4533) & (n_n4587)) + ((!x15x) & (!x583x) & (!n_n4557) & (n_n4533) & (!n_n4587)) + ((!x15x) & (!x583x) & (!n_n4557) & (n_n4533) & (n_n4587)) + ((!x15x) & (!x583x) & (n_n4557) & (!n_n4533) & (!n_n4587)) + ((!x15x) & (!x583x) & (n_n4557) & (!n_n4533) & (n_n4587)) + ((!x15x) & (!x583x) & (n_n4557) & (n_n4533) & (!n_n4587)) + ((!x15x) & (!x583x) & (n_n4557) & (n_n4533) & (n_n4587)) + ((!x15x) & (x583x) & (!n_n4557) & (!n_n4533) & (n_n4587)) + ((!x15x) & (x583x) & (!n_n4557) & (n_n4533) & (!n_n4587)) + ((!x15x) & (x583x) & (!n_n4557) & (n_n4533) & (n_n4587)) + ((!x15x) & (x583x) & (n_n4557) & (!n_n4533) & (!n_n4587)) + ((!x15x) & (x583x) & (n_n4557) & (!n_n4533) & (n_n4587)) + ((!x15x) & (x583x) & (n_n4557) & (n_n4533) & (!n_n4587)) + ((!x15x) & (x583x) & (n_n4557) & (n_n4533) & (n_n4587)) + ((x15x) & (!x583x) & (!n_n4557) & (!n_n4533) & (n_n4587)) + ((x15x) & (!x583x) & (!n_n4557) & (n_n4533) & (!n_n4587)) + ((x15x) & (!x583x) & (!n_n4557) & (n_n4533) & (n_n4587)) + ((x15x) & (!x583x) & (n_n4557) & (!n_n4533) & (!n_n4587)) + ((x15x) & (!x583x) & (n_n4557) & (!n_n4533) & (n_n4587)) + ((x15x) & (!x583x) & (n_n4557) & (n_n4533) & (!n_n4587)) + ((x15x) & (!x583x) & (n_n4557) & (n_n4533) & (n_n4587)) + ((x15x) & (x583x) & (!n_n4557) & (!n_n4533) & (!n_n4587)) + ((x15x) & (x583x) & (!n_n4557) & (!n_n4533) & (n_n4587)) + ((x15x) & (x583x) & (!n_n4557) & (n_n4533) & (!n_n4587)) + ((x15x) & (x583x) & (!n_n4557) & (n_n4533) & (n_n4587)) + ((x15x) & (x583x) & (n_n4557) & (!n_n4533) & (!n_n4587)) + ((x15x) & (x583x) & (n_n4557) & (!n_n4533) & (n_n4587)) + ((x15x) & (x583x) & (n_n4557) & (n_n4533) & (!n_n4587)) + ((x15x) & (x583x) & (n_n4557) & (n_n4533) & (n_n4587)));
	assign x14847x = (((!n_n4593) & (!n_n4571) & (!n_n4592) & (!n_n4556) & (n_n4527)) + ((!n_n4593) & (!n_n4571) & (!n_n4592) & (n_n4556) & (!n_n4527)) + ((!n_n4593) & (!n_n4571) & (!n_n4592) & (n_n4556) & (n_n4527)) + ((!n_n4593) & (!n_n4571) & (n_n4592) & (!n_n4556) & (!n_n4527)) + ((!n_n4593) & (!n_n4571) & (n_n4592) & (!n_n4556) & (n_n4527)) + ((!n_n4593) & (!n_n4571) & (n_n4592) & (n_n4556) & (!n_n4527)) + ((!n_n4593) & (!n_n4571) & (n_n4592) & (n_n4556) & (n_n4527)) + ((!n_n4593) & (n_n4571) & (!n_n4592) & (!n_n4556) & (!n_n4527)) + ((!n_n4593) & (n_n4571) & (!n_n4592) & (!n_n4556) & (n_n4527)) + ((!n_n4593) & (n_n4571) & (!n_n4592) & (n_n4556) & (!n_n4527)) + ((!n_n4593) & (n_n4571) & (!n_n4592) & (n_n4556) & (n_n4527)) + ((!n_n4593) & (n_n4571) & (n_n4592) & (!n_n4556) & (!n_n4527)) + ((!n_n4593) & (n_n4571) & (n_n4592) & (!n_n4556) & (n_n4527)) + ((!n_n4593) & (n_n4571) & (n_n4592) & (n_n4556) & (!n_n4527)) + ((!n_n4593) & (n_n4571) & (n_n4592) & (n_n4556) & (n_n4527)) + ((n_n4593) & (!n_n4571) & (!n_n4592) & (!n_n4556) & (!n_n4527)) + ((n_n4593) & (!n_n4571) & (!n_n4592) & (!n_n4556) & (n_n4527)) + ((n_n4593) & (!n_n4571) & (!n_n4592) & (n_n4556) & (!n_n4527)) + ((n_n4593) & (!n_n4571) & (!n_n4592) & (n_n4556) & (n_n4527)) + ((n_n4593) & (!n_n4571) & (n_n4592) & (!n_n4556) & (!n_n4527)) + ((n_n4593) & (!n_n4571) & (n_n4592) & (!n_n4556) & (n_n4527)) + ((n_n4593) & (!n_n4571) & (n_n4592) & (n_n4556) & (!n_n4527)) + ((n_n4593) & (!n_n4571) & (n_n4592) & (n_n4556) & (n_n4527)) + ((n_n4593) & (n_n4571) & (!n_n4592) & (!n_n4556) & (!n_n4527)) + ((n_n4593) & (n_n4571) & (!n_n4592) & (!n_n4556) & (n_n4527)) + ((n_n4593) & (n_n4571) & (!n_n4592) & (n_n4556) & (!n_n4527)) + ((n_n4593) & (n_n4571) & (!n_n4592) & (n_n4556) & (n_n4527)) + ((n_n4593) & (n_n4571) & (n_n4592) & (!n_n4556) & (!n_n4527)) + ((n_n4593) & (n_n4571) & (n_n4592) & (!n_n4556) & (n_n4527)) + ((n_n4593) & (n_n4571) & (n_n4592) & (n_n4556) & (!n_n4527)) + ((n_n4593) & (n_n4571) & (n_n4592) & (n_n4556) & (n_n4527)));
	assign x14887x = (((!n_n4440) & (!n_n4453) & (!n_n4420) & (!n_n4407) & (n_n4444)) + ((!n_n4440) & (!n_n4453) & (!n_n4420) & (n_n4407) & (!n_n4444)) + ((!n_n4440) & (!n_n4453) & (!n_n4420) & (n_n4407) & (n_n4444)) + ((!n_n4440) & (!n_n4453) & (n_n4420) & (!n_n4407) & (!n_n4444)) + ((!n_n4440) & (!n_n4453) & (n_n4420) & (!n_n4407) & (n_n4444)) + ((!n_n4440) & (!n_n4453) & (n_n4420) & (n_n4407) & (!n_n4444)) + ((!n_n4440) & (!n_n4453) & (n_n4420) & (n_n4407) & (n_n4444)) + ((!n_n4440) & (n_n4453) & (!n_n4420) & (!n_n4407) & (!n_n4444)) + ((!n_n4440) & (n_n4453) & (!n_n4420) & (!n_n4407) & (n_n4444)) + ((!n_n4440) & (n_n4453) & (!n_n4420) & (n_n4407) & (!n_n4444)) + ((!n_n4440) & (n_n4453) & (!n_n4420) & (n_n4407) & (n_n4444)) + ((!n_n4440) & (n_n4453) & (n_n4420) & (!n_n4407) & (!n_n4444)) + ((!n_n4440) & (n_n4453) & (n_n4420) & (!n_n4407) & (n_n4444)) + ((!n_n4440) & (n_n4453) & (n_n4420) & (n_n4407) & (!n_n4444)) + ((!n_n4440) & (n_n4453) & (n_n4420) & (n_n4407) & (n_n4444)) + ((n_n4440) & (!n_n4453) & (!n_n4420) & (!n_n4407) & (!n_n4444)) + ((n_n4440) & (!n_n4453) & (!n_n4420) & (!n_n4407) & (n_n4444)) + ((n_n4440) & (!n_n4453) & (!n_n4420) & (n_n4407) & (!n_n4444)) + ((n_n4440) & (!n_n4453) & (!n_n4420) & (n_n4407) & (n_n4444)) + ((n_n4440) & (!n_n4453) & (n_n4420) & (!n_n4407) & (!n_n4444)) + ((n_n4440) & (!n_n4453) & (n_n4420) & (!n_n4407) & (n_n4444)) + ((n_n4440) & (!n_n4453) & (n_n4420) & (n_n4407) & (!n_n4444)) + ((n_n4440) & (!n_n4453) & (n_n4420) & (n_n4407) & (n_n4444)) + ((n_n4440) & (n_n4453) & (!n_n4420) & (!n_n4407) & (!n_n4444)) + ((n_n4440) & (n_n4453) & (!n_n4420) & (!n_n4407) & (n_n4444)) + ((n_n4440) & (n_n4453) & (!n_n4420) & (n_n4407) & (!n_n4444)) + ((n_n4440) & (n_n4453) & (!n_n4420) & (n_n4407) & (n_n4444)) + ((n_n4440) & (n_n4453) & (n_n4420) & (!n_n4407) & (!n_n4444)) + ((n_n4440) & (n_n4453) & (n_n4420) & (!n_n4407) & (n_n4444)) + ((n_n4440) & (n_n4453) & (n_n4420) & (n_n4407) & (!n_n4444)) + ((n_n4440) & (n_n4453) & (n_n4420) & (n_n4407) & (n_n4444)));
	assign x14889x = (((!x14876x) & (!x14877x) & (!x14882x) & (x14883x)) + ((!x14876x) & (!x14877x) & (x14882x) & (!x14883x)) + ((!x14876x) & (!x14877x) & (x14882x) & (x14883x)) + ((!x14876x) & (x14877x) & (!x14882x) & (!x14883x)) + ((!x14876x) & (x14877x) & (!x14882x) & (x14883x)) + ((!x14876x) & (x14877x) & (x14882x) & (!x14883x)) + ((!x14876x) & (x14877x) & (x14882x) & (x14883x)) + ((x14876x) & (!x14877x) & (!x14882x) & (!x14883x)) + ((x14876x) & (!x14877x) & (!x14882x) & (x14883x)) + ((x14876x) & (!x14877x) & (x14882x) & (!x14883x)) + ((x14876x) & (!x14877x) & (x14882x) & (x14883x)) + ((x14876x) & (x14877x) & (!x14882x) & (!x14883x)) + ((x14876x) & (x14877x) & (!x14882x) & (x14883x)) + ((x14876x) & (x14877x) & (x14882x) & (!x14883x)) + ((x14876x) & (x14877x) & (x14882x) & (x14883x)));
	assign x14890x = (((!x323x) & (!n_n4416) & (!n_n4415) & (!x14887x) & (x14889x)) + ((!x323x) & (!n_n4416) & (!n_n4415) & (x14887x) & (!x14889x)) + ((!x323x) & (!n_n4416) & (!n_n4415) & (x14887x) & (x14889x)) + ((!x323x) & (!n_n4416) & (n_n4415) & (!x14887x) & (!x14889x)) + ((!x323x) & (!n_n4416) & (n_n4415) & (!x14887x) & (x14889x)) + ((!x323x) & (!n_n4416) & (n_n4415) & (x14887x) & (!x14889x)) + ((!x323x) & (!n_n4416) & (n_n4415) & (x14887x) & (x14889x)) + ((!x323x) & (n_n4416) & (!n_n4415) & (!x14887x) & (!x14889x)) + ((!x323x) & (n_n4416) & (!n_n4415) & (!x14887x) & (x14889x)) + ((!x323x) & (n_n4416) & (!n_n4415) & (x14887x) & (!x14889x)) + ((!x323x) & (n_n4416) & (!n_n4415) & (x14887x) & (x14889x)) + ((!x323x) & (n_n4416) & (n_n4415) & (!x14887x) & (!x14889x)) + ((!x323x) & (n_n4416) & (n_n4415) & (!x14887x) & (x14889x)) + ((!x323x) & (n_n4416) & (n_n4415) & (x14887x) & (!x14889x)) + ((!x323x) & (n_n4416) & (n_n4415) & (x14887x) & (x14889x)) + ((x323x) & (!n_n4416) & (!n_n4415) & (!x14887x) & (!x14889x)) + ((x323x) & (!n_n4416) & (!n_n4415) & (!x14887x) & (x14889x)) + ((x323x) & (!n_n4416) & (!n_n4415) & (x14887x) & (!x14889x)) + ((x323x) & (!n_n4416) & (!n_n4415) & (x14887x) & (x14889x)) + ((x323x) & (!n_n4416) & (n_n4415) & (!x14887x) & (!x14889x)) + ((x323x) & (!n_n4416) & (n_n4415) & (!x14887x) & (x14889x)) + ((x323x) & (!n_n4416) & (n_n4415) & (x14887x) & (!x14889x)) + ((x323x) & (!n_n4416) & (n_n4415) & (x14887x) & (x14889x)) + ((x323x) & (n_n4416) & (!n_n4415) & (!x14887x) & (!x14889x)) + ((x323x) & (n_n4416) & (!n_n4415) & (!x14887x) & (x14889x)) + ((x323x) & (n_n4416) & (!n_n4415) & (x14887x) & (!x14889x)) + ((x323x) & (n_n4416) & (!n_n4415) & (x14887x) & (x14889x)) + ((x323x) & (n_n4416) & (n_n4415) & (!x14887x) & (!x14889x)) + ((x323x) & (n_n4416) & (n_n4415) & (!x14887x) & (x14889x)) + ((x323x) & (n_n4416) & (n_n4415) & (x14887x) & (!x14889x)) + ((x323x) & (n_n4416) & (n_n4415) & (x14887x) & (x14889x)));
	assign x14891x = (((!x14849x) & (!x14870x) & (!x14871x) & (!x14846x) & (x14847x)) + ((!x14849x) & (!x14870x) & (!x14871x) & (x14846x) & (!x14847x)) + ((!x14849x) & (!x14870x) & (!x14871x) & (x14846x) & (x14847x)) + ((!x14849x) & (!x14870x) & (x14871x) & (!x14846x) & (!x14847x)) + ((!x14849x) & (!x14870x) & (x14871x) & (!x14846x) & (x14847x)) + ((!x14849x) & (!x14870x) & (x14871x) & (x14846x) & (!x14847x)) + ((!x14849x) & (!x14870x) & (x14871x) & (x14846x) & (x14847x)) + ((!x14849x) & (x14870x) & (!x14871x) & (!x14846x) & (!x14847x)) + ((!x14849x) & (x14870x) & (!x14871x) & (!x14846x) & (x14847x)) + ((!x14849x) & (x14870x) & (!x14871x) & (x14846x) & (!x14847x)) + ((!x14849x) & (x14870x) & (!x14871x) & (x14846x) & (x14847x)) + ((!x14849x) & (x14870x) & (x14871x) & (!x14846x) & (!x14847x)) + ((!x14849x) & (x14870x) & (x14871x) & (!x14846x) & (x14847x)) + ((!x14849x) & (x14870x) & (x14871x) & (x14846x) & (!x14847x)) + ((!x14849x) & (x14870x) & (x14871x) & (x14846x) & (x14847x)) + ((x14849x) & (!x14870x) & (!x14871x) & (!x14846x) & (!x14847x)) + ((x14849x) & (!x14870x) & (!x14871x) & (!x14846x) & (x14847x)) + ((x14849x) & (!x14870x) & (!x14871x) & (x14846x) & (!x14847x)) + ((x14849x) & (!x14870x) & (!x14871x) & (x14846x) & (x14847x)) + ((x14849x) & (!x14870x) & (x14871x) & (!x14846x) & (!x14847x)) + ((x14849x) & (!x14870x) & (x14871x) & (!x14846x) & (x14847x)) + ((x14849x) & (!x14870x) & (x14871x) & (x14846x) & (!x14847x)) + ((x14849x) & (!x14870x) & (x14871x) & (x14846x) & (x14847x)) + ((x14849x) & (x14870x) & (!x14871x) & (!x14846x) & (!x14847x)) + ((x14849x) & (x14870x) & (!x14871x) & (!x14846x) & (x14847x)) + ((x14849x) & (x14870x) & (!x14871x) & (x14846x) & (!x14847x)) + ((x14849x) & (x14870x) & (!x14871x) & (x14846x) & (x14847x)) + ((x14849x) & (x14870x) & (x14871x) & (!x14846x) & (!x14847x)) + ((x14849x) & (x14870x) & (x14871x) & (!x14846x) & (x14847x)) + ((x14849x) & (x14870x) & (x14871x) & (x14846x) & (!x14847x)) + ((x14849x) & (x14870x) & (x14871x) & (x14846x) & (x14847x)));
	assign x14932x = (((!n_n524) & (!n_n509) & (!x17x) & (!n_n4863) & (n_n2727)) + ((!n_n524) & (!n_n509) & (!x17x) & (n_n4863) & (!n_n2727)) + ((!n_n524) & (!n_n509) & (!x17x) & (n_n4863) & (n_n2727)) + ((!n_n524) & (!n_n509) & (x17x) & (!n_n4863) & (n_n2727)) + ((!n_n524) & (!n_n509) & (x17x) & (n_n4863) & (!n_n2727)) + ((!n_n524) & (!n_n509) & (x17x) & (n_n4863) & (n_n2727)) + ((!n_n524) & (n_n509) & (!x17x) & (!n_n4863) & (n_n2727)) + ((!n_n524) & (n_n509) & (!x17x) & (n_n4863) & (!n_n2727)) + ((!n_n524) & (n_n509) & (!x17x) & (n_n4863) & (n_n2727)) + ((!n_n524) & (n_n509) & (x17x) & (!n_n4863) & (n_n2727)) + ((!n_n524) & (n_n509) & (x17x) & (n_n4863) & (!n_n2727)) + ((!n_n524) & (n_n509) & (x17x) & (n_n4863) & (n_n2727)) + ((n_n524) & (!n_n509) & (!x17x) & (!n_n4863) & (n_n2727)) + ((n_n524) & (!n_n509) & (!x17x) & (n_n4863) & (!n_n2727)) + ((n_n524) & (!n_n509) & (!x17x) & (n_n4863) & (n_n2727)) + ((n_n524) & (!n_n509) & (x17x) & (!n_n4863) & (n_n2727)) + ((n_n524) & (!n_n509) & (x17x) & (n_n4863) & (!n_n2727)) + ((n_n524) & (!n_n509) & (x17x) & (n_n4863) & (n_n2727)) + ((n_n524) & (n_n509) & (!x17x) & (!n_n4863) & (n_n2727)) + ((n_n524) & (n_n509) & (!x17x) & (n_n4863) & (!n_n2727)) + ((n_n524) & (n_n509) & (!x17x) & (n_n4863) & (n_n2727)) + ((n_n524) & (n_n509) & (x17x) & (!n_n4863) & (!n_n2727)) + ((n_n524) & (n_n509) & (x17x) & (!n_n4863) & (n_n2727)) + ((n_n524) & (n_n509) & (x17x) & (n_n4863) & (!n_n2727)) + ((n_n524) & (n_n509) & (x17x) & (n_n4863) & (n_n2727)));
	assign x15096x = (((!i_9_) & (n_n524) & (n_n482) & (n_n455) & (!n_n528)) + ((!i_9_) & (n_n524) & (n_n482) & (n_n455) & (n_n528)) + ((i_9_) & (!n_n524) & (n_n482) & (n_n455) & (n_n528)) + ((i_9_) & (n_n524) & (n_n482) & (n_n455) & (n_n528)));
	assign x15098x = (((!i_9_) & (n_n482) & (n_n455) & (n_n532) & (!n_n520)) + ((!i_9_) & (n_n482) & (n_n455) & (n_n532) & (n_n520)) + ((i_9_) & (n_n482) & (n_n455) & (!n_n532) & (n_n520)) + ((i_9_) & (n_n482) & (n_n455) & (n_n532) & (!n_n520)) + ((i_9_) & (n_n482) & (n_n455) & (n_n532) & (n_n520)));
	assign x15164x = (((!n_n4340) & (!n_n4353) & (!n_n4354) & (!n_n4350) & (n_n4348)) + ((!n_n4340) & (!n_n4353) & (!n_n4354) & (n_n4350) & (!n_n4348)) + ((!n_n4340) & (!n_n4353) & (!n_n4354) & (n_n4350) & (n_n4348)) + ((!n_n4340) & (!n_n4353) & (n_n4354) & (!n_n4350) & (!n_n4348)) + ((!n_n4340) & (!n_n4353) & (n_n4354) & (!n_n4350) & (n_n4348)) + ((!n_n4340) & (!n_n4353) & (n_n4354) & (n_n4350) & (!n_n4348)) + ((!n_n4340) & (!n_n4353) & (n_n4354) & (n_n4350) & (n_n4348)) + ((!n_n4340) & (n_n4353) & (!n_n4354) & (!n_n4350) & (!n_n4348)) + ((!n_n4340) & (n_n4353) & (!n_n4354) & (!n_n4350) & (n_n4348)) + ((!n_n4340) & (n_n4353) & (!n_n4354) & (n_n4350) & (!n_n4348)) + ((!n_n4340) & (n_n4353) & (!n_n4354) & (n_n4350) & (n_n4348)) + ((!n_n4340) & (n_n4353) & (n_n4354) & (!n_n4350) & (!n_n4348)) + ((!n_n4340) & (n_n4353) & (n_n4354) & (!n_n4350) & (n_n4348)) + ((!n_n4340) & (n_n4353) & (n_n4354) & (n_n4350) & (!n_n4348)) + ((!n_n4340) & (n_n4353) & (n_n4354) & (n_n4350) & (n_n4348)) + ((n_n4340) & (!n_n4353) & (!n_n4354) & (!n_n4350) & (!n_n4348)) + ((n_n4340) & (!n_n4353) & (!n_n4354) & (!n_n4350) & (n_n4348)) + ((n_n4340) & (!n_n4353) & (!n_n4354) & (n_n4350) & (!n_n4348)) + ((n_n4340) & (!n_n4353) & (!n_n4354) & (n_n4350) & (n_n4348)) + ((n_n4340) & (!n_n4353) & (n_n4354) & (!n_n4350) & (!n_n4348)) + ((n_n4340) & (!n_n4353) & (n_n4354) & (!n_n4350) & (n_n4348)) + ((n_n4340) & (!n_n4353) & (n_n4354) & (n_n4350) & (!n_n4348)) + ((n_n4340) & (!n_n4353) & (n_n4354) & (n_n4350) & (n_n4348)) + ((n_n4340) & (n_n4353) & (!n_n4354) & (!n_n4350) & (!n_n4348)) + ((n_n4340) & (n_n4353) & (!n_n4354) & (!n_n4350) & (n_n4348)) + ((n_n4340) & (n_n4353) & (!n_n4354) & (n_n4350) & (!n_n4348)) + ((n_n4340) & (n_n4353) & (!n_n4354) & (n_n4350) & (n_n4348)) + ((n_n4340) & (n_n4353) & (n_n4354) & (!n_n4350) & (!n_n4348)) + ((n_n4340) & (n_n4353) & (n_n4354) & (!n_n4350) & (n_n4348)) + ((n_n4340) & (n_n4353) & (n_n4354) & (n_n4350) & (!n_n4348)) + ((n_n4340) & (n_n4353) & (n_n4354) & (n_n4350) & (n_n4348)));
	assign x15246x = (((!n_n5100) & (!n_n5103) & (!n_n5102) & (n_n5106)) + ((!n_n5100) & (!n_n5103) & (n_n5102) & (!n_n5106)) + ((!n_n5100) & (!n_n5103) & (n_n5102) & (n_n5106)) + ((!n_n5100) & (n_n5103) & (!n_n5102) & (!n_n5106)) + ((!n_n5100) & (n_n5103) & (!n_n5102) & (n_n5106)) + ((!n_n5100) & (n_n5103) & (n_n5102) & (!n_n5106)) + ((!n_n5100) & (n_n5103) & (n_n5102) & (n_n5106)) + ((n_n5100) & (!n_n5103) & (!n_n5102) & (!n_n5106)) + ((n_n5100) & (!n_n5103) & (!n_n5102) & (n_n5106)) + ((n_n5100) & (!n_n5103) & (n_n5102) & (!n_n5106)) + ((n_n5100) & (!n_n5103) & (n_n5102) & (n_n5106)) + ((n_n5100) & (n_n5103) & (!n_n5102) & (!n_n5106)) + ((n_n5100) & (n_n5103) & (!n_n5102) & (n_n5106)) + ((n_n5100) & (n_n5103) & (n_n5102) & (!n_n5106)) + ((n_n5100) & (n_n5103) & (n_n5102) & (n_n5106)));
	assign x22184x = (((!x21x) & (!x11x) & (!n_n130) & (!n_n500) & (!n_n5137)) + ((!x21x) & (!x11x) & (!n_n130) & (n_n500) & (!n_n5137)) + ((!x21x) & (!x11x) & (n_n130) & (!n_n500) & (!n_n5137)) + ((!x21x) & (!x11x) & (n_n130) & (n_n500) & (!n_n5137)) + ((!x21x) & (x11x) & (!n_n130) & (!n_n500) & (!n_n5137)) + ((!x21x) & (x11x) & (!n_n130) & (n_n500) & (!n_n5137)) + ((!x21x) & (x11x) & (n_n130) & (!n_n500) & (!n_n5137)) + ((x21x) & (!x11x) & (!n_n130) & (!n_n500) & (!n_n5137)) + ((x21x) & (!x11x) & (!n_n130) & (n_n500) & (!n_n5137)) + ((x21x) & (!x11x) & (n_n130) & (!n_n500) & (!n_n5137)) + ((x21x) & (x11x) & (!n_n130) & (!n_n500) & (!n_n5137)) + ((x21x) & (x11x) & (!n_n130) & (n_n500) & (!n_n5137)) + ((x21x) & (x11x) & (n_n130) & (!n_n500) & (!n_n5137)));
	assign x15396x = (((!n_n4921) & (!n_n4938) & (!n_n4936) & (n_n4917)) + ((!n_n4921) & (!n_n4938) & (n_n4936) & (!n_n4917)) + ((!n_n4921) & (!n_n4938) & (n_n4936) & (n_n4917)) + ((!n_n4921) & (n_n4938) & (!n_n4936) & (!n_n4917)) + ((!n_n4921) & (n_n4938) & (!n_n4936) & (n_n4917)) + ((!n_n4921) & (n_n4938) & (n_n4936) & (!n_n4917)) + ((!n_n4921) & (n_n4938) & (n_n4936) & (n_n4917)) + ((n_n4921) & (!n_n4938) & (!n_n4936) & (!n_n4917)) + ((n_n4921) & (!n_n4938) & (!n_n4936) & (n_n4917)) + ((n_n4921) & (!n_n4938) & (n_n4936) & (!n_n4917)) + ((n_n4921) & (!n_n4938) & (n_n4936) & (n_n4917)) + ((n_n4921) & (n_n4938) & (!n_n4936) & (!n_n4917)) + ((n_n4921) & (n_n4938) & (!n_n4936) & (n_n4917)) + ((n_n4921) & (n_n4938) & (n_n4936) & (!n_n4917)) + ((n_n4921) & (n_n4938) & (n_n4936) & (n_n4917)));
	assign x22090x = (((!x25x) & (!x523x) & (!n_n4560) & (!n_n4561) & (!n_n4556)) + ((!x25x) & (x523x) & (!n_n4560) & (!n_n4561) & (!n_n4556)) + ((x25x) & (!x523x) & (!n_n4560) & (!n_n4561) & (!n_n4556)));
	assign x15671x = (((!n_n5331) & (!n_n5332) & (!n_n5328) & (!n_n5335) & (n_n5334)) + ((!n_n5331) & (!n_n5332) & (!n_n5328) & (n_n5335) & (!n_n5334)) + ((!n_n5331) & (!n_n5332) & (!n_n5328) & (n_n5335) & (n_n5334)) + ((!n_n5331) & (!n_n5332) & (n_n5328) & (!n_n5335) & (!n_n5334)) + ((!n_n5331) & (!n_n5332) & (n_n5328) & (!n_n5335) & (n_n5334)) + ((!n_n5331) & (!n_n5332) & (n_n5328) & (n_n5335) & (!n_n5334)) + ((!n_n5331) & (!n_n5332) & (n_n5328) & (n_n5335) & (n_n5334)) + ((!n_n5331) & (n_n5332) & (!n_n5328) & (!n_n5335) & (!n_n5334)) + ((!n_n5331) & (n_n5332) & (!n_n5328) & (!n_n5335) & (n_n5334)) + ((!n_n5331) & (n_n5332) & (!n_n5328) & (n_n5335) & (!n_n5334)) + ((!n_n5331) & (n_n5332) & (!n_n5328) & (n_n5335) & (n_n5334)) + ((!n_n5331) & (n_n5332) & (n_n5328) & (!n_n5335) & (!n_n5334)) + ((!n_n5331) & (n_n5332) & (n_n5328) & (!n_n5335) & (n_n5334)) + ((!n_n5331) & (n_n5332) & (n_n5328) & (n_n5335) & (!n_n5334)) + ((!n_n5331) & (n_n5332) & (n_n5328) & (n_n5335) & (n_n5334)) + ((n_n5331) & (!n_n5332) & (!n_n5328) & (!n_n5335) & (!n_n5334)) + ((n_n5331) & (!n_n5332) & (!n_n5328) & (!n_n5335) & (n_n5334)) + ((n_n5331) & (!n_n5332) & (!n_n5328) & (n_n5335) & (!n_n5334)) + ((n_n5331) & (!n_n5332) & (!n_n5328) & (n_n5335) & (n_n5334)) + ((n_n5331) & (!n_n5332) & (n_n5328) & (!n_n5335) & (!n_n5334)) + ((n_n5331) & (!n_n5332) & (n_n5328) & (!n_n5335) & (n_n5334)) + ((n_n5331) & (!n_n5332) & (n_n5328) & (n_n5335) & (!n_n5334)) + ((n_n5331) & (!n_n5332) & (n_n5328) & (n_n5335) & (n_n5334)) + ((n_n5331) & (n_n5332) & (!n_n5328) & (!n_n5335) & (!n_n5334)) + ((n_n5331) & (n_n5332) & (!n_n5328) & (!n_n5335) & (n_n5334)) + ((n_n5331) & (n_n5332) & (!n_n5328) & (n_n5335) & (!n_n5334)) + ((n_n5331) & (n_n5332) & (!n_n5328) & (n_n5335) & (n_n5334)) + ((n_n5331) & (n_n5332) & (n_n5328) & (!n_n5335) & (!n_n5334)) + ((n_n5331) & (n_n5332) & (n_n5328) & (!n_n5335) & (n_n5334)) + ((n_n5331) & (n_n5332) & (n_n5328) & (n_n5335) & (!n_n5334)) + ((n_n5331) & (n_n5332) & (n_n5328) & (n_n5335) & (n_n5334)));
	assign x15735x = (((!i_9_) & (n_n526) & (n_n482) & (n_n260) & (!n_n522)) + ((!i_9_) & (n_n526) & (n_n482) & (n_n260) & (n_n522)) + ((i_9_) & (!n_n526) & (n_n482) & (n_n260) & (n_n522)) + ((i_9_) & (n_n526) & (n_n482) & (n_n260) & (n_n522)));
	assign x15737x = (((!i_7_) & (!i_8_) & (i_6_) & (n_n482) & (x17x)) + ((i_7_) & (!i_8_) & (!i_6_) & (n_n482) & (x17x)) + ((i_7_) & (i_8_) & (!i_6_) & (n_n482) & (x17x)));
	assign x15775x = (((!n_n4712) & (!n_n4685) & (!n_n4695) & (n_n4694)) + ((!n_n4712) & (!n_n4685) & (n_n4695) & (!n_n4694)) + ((!n_n4712) & (!n_n4685) & (n_n4695) & (n_n4694)) + ((!n_n4712) & (n_n4685) & (!n_n4695) & (!n_n4694)) + ((!n_n4712) & (n_n4685) & (!n_n4695) & (n_n4694)) + ((!n_n4712) & (n_n4685) & (n_n4695) & (!n_n4694)) + ((!n_n4712) & (n_n4685) & (n_n4695) & (n_n4694)) + ((n_n4712) & (!n_n4685) & (!n_n4695) & (!n_n4694)) + ((n_n4712) & (!n_n4685) & (!n_n4695) & (n_n4694)) + ((n_n4712) & (!n_n4685) & (n_n4695) & (!n_n4694)) + ((n_n4712) & (!n_n4685) & (n_n4695) & (n_n4694)) + ((n_n4712) & (n_n4685) & (!n_n4695) & (!n_n4694)) + ((n_n4712) & (n_n4685) & (!n_n4695) & (n_n4694)) + ((n_n4712) & (n_n4685) & (n_n4695) & (!n_n4694)) + ((n_n4712) & (n_n4685) & (n_n4695) & (n_n4694)));
	assign x15802x = (((!n_n4882) & (!n_n4878) & (!n_n4875) & (n_n4873)) + ((!n_n4882) & (!n_n4878) & (n_n4875) & (!n_n4873)) + ((!n_n4882) & (!n_n4878) & (n_n4875) & (n_n4873)) + ((!n_n4882) & (n_n4878) & (!n_n4875) & (!n_n4873)) + ((!n_n4882) & (n_n4878) & (!n_n4875) & (n_n4873)) + ((!n_n4882) & (n_n4878) & (n_n4875) & (!n_n4873)) + ((!n_n4882) & (n_n4878) & (n_n4875) & (n_n4873)) + ((n_n4882) & (!n_n4878) & (!n_n4875) & (!n_n4873)) + ((n_n4882) & (!n_n4878) & (!n_n4875) & (n_n4873)) + ((n_n4882) & (!n_n4878) & (n_n4875) & (!n_n4873)) + ((n_n4882) & (!n_n4878) & (n_n4875) & (n_n4873)) + ((n_n4882) & (n_n4878) & (!n_n4875) & (!n_n4873)) + ((n_n4882) & (n_n4878) & (!n_n4875) & (n_n4873)) + ((n_n4882) & (n_n4878) & (n_n4875) & (!n_n4873)) + ((n_n4882) & (n_n4878) & (n_n4875) & (n_n4873)));
	assign x15803x = (((!x17x) & (!n_n522) & (!n_n500) & (!n_n3450) & (n_n4879)) + ((!x17x) & (!n_n522) & (!n_n500) & (n_n3450) & (!n_n4879)) + ((!x17x) & (!n_n522) & (!n_n500) & (n_n3450) & (n_n4879)) + ((!x17x) & (!n_n522) & (n_n500) & (!n_n3450) & (n_n4879)) + ((!x17x) & (!n_n522) & (n_n500) & (n_n3450) & (!n_n4879)) + ((!x17x) & (!n_n522) & (n_n500) & (n_n3450) & (n_n4879)) + ((!x17x) & (n_n522) & (!n_n500) & (!n_n3450) & (n_n4879)) + ((!x17x) & (n_n522) & (!n_n500) & (n_n3450) & (!n_n4879)) + ((!x17x) & (n_n522) & (!n_n500) & (n_n3450) & (n_n4879)) + ((!x17x) & (n_n522) & (n_n500) & (!n_n3450) & (n_n4879)) + ((!x17x) & (n_n522) & (n_n500) & (n_n3450) & (!n_n4879)) + ((!x17x) & (n_n522) & (n_n500) & (n_n3450) & (n_n4879)) + ((x17x) & (!n_n522) & (!n_n500) & (!n_n3450) & (n_n4879)) + ((x17x) & (!n_n522) & (!n_n500) & (n_n3450) & (!n_n4879)) + ((x17x) & (!n_n522) & (!n_n500) & (n_n3450) & (n_n4879)) + ((x17x) & (!n_n522) & (n_n500) & (!n_n3450) & (n_n4879)) + ((x17x) & (!n_n522) & (n_n500) & (n_n3450) & (!n_n4879)) + ((x17x) & (!n_n522) & (n_n500) & (n_n3450) & (n_n4879)) + ((x17x) & (n_n522) & (!n_n500) & (!n_n3450) & (n_n4879)) + ((x17x) & (n_n522) & (!n_n500) & (n_n3450) & (!n_n4879)) + ((x17x) & (n_n522) & (!n_n500) & (n_n3450) & (n_n4879)) + ((x17x) & (n_n522) & (n_n500) & (!n_n3450) & (!n_n4879)) + ((x17x) & (n_n522) & (n_n500) & (!n_n3450) & (n_n4879)) + ((x17x) & (n_n522) & (n_n500) & (n_n3450) & (!n_n4879)) + ((x17x) & (n_n522) & (n_n500) & (n_n3450) & (n_n4879)));
	assign x15811x = (((!x15308x) & (!x15309x) & (!n_n2844) & (n_n2846)) + ((!x15308x) & (!x15309x) & (n_n2844) & (!n_n2846)) + ((!x15308x) & (!x15309x) & (n_n2844) & (n_n2846)) + ((!x15308x) & (x15309x) & (!n_n2844) & (!n_n2846)) + ((!x15308x) & (x15309x) & (!n_n2844) & (n_n2846)) + ((!x15308x) & (x15309x) & (n_n2844) & (!n_n2846)) + ((!x15308x) & (x15309x) & (n_n2844) & (n_n2846)) + ((x15308x) & (!x15309x) & (!n_n2844) & (!n_n2846)) + ((x15308x) & (!x15309x) & (!n_n2844) & (n_n2846)) + ((x15308x) & (!x15309x) & (n_n2844) & (!n_n2846)) + ((x15308x) & (!x15309x) & (n_n2844) & (n_n2846)) + ((x15308x) & (x15309x) & (!n_n2844) & (!n_n2846)) + ((x15308x) & (x15309x) & (!n_n2844) & (n_n2846)) + ((x15308x) & (x15309x) & (n_n2844) & (!n_n2846)) + ((x15308x) & (x15309x) & (n_n2844) & (n_n2846)));
	assign x15898x = (((!x592x) & (!n_n5331) & (!x23x) & (!n_n5325) & (n_n5333)) + ((!x592x) & (!n_n5331) & (!x23x) & (n_n5325) & (!n_n5333)) + ((!x592x) & (!n_n5331) & (!x23x) & (n_n5325) & (n_n5333)) + ((!x592x) & (!n_n5331) & (x23x) & (!n_n5325) & (n_n5333)) + ((!x592x) & (!n_n5331) & (x23x) & (n_n5325) & (!n_n5333)) + ((!x592x) & (!n_n5331) & (x23x) & (n_n5325) & (n_n5333)) + ((!x592x) & (n_n5331) & (!x23x) & (!n_n5325) & (!n_n5333)) + ((!x592x) & (n_n5331) & (!x23x) & (!n_n5325) & (n_n5333)) + ((!x592x) & (n_n5331) & (!x23x) & (n_n5325) & (!n_n5333)) + ((!x592x) & (n_n5331) & (!x23x) & (n_n5325) & (n_n5333)) + ((!x592x) & (n_n5331) & (x23x) & (!n_n5325) & (!n_n5333)) + ((!x592x) & (n_n5331) & (x23x) & (!n_n5325) & (n_n5333)) + ((!x592x) & (n_n5331) & (x23x) & (n_n5325) & (!n_n5333)) + ((!x592x) & (n_n5331) & (x23x) & (n_n5325) & (n_n5333)) + ((x592x) & (!n_n5331) & (!x23x) & (!n_n5325) & (n_n5333)) + ((x592x) & (!n_n5331) & (!x23x) & (n_n5325) & (!n_n5333)) + ((x592x) & (!n_n5331) & (!x23x) & (n_n5325) & (n_n5333)) + ((x592x) & (!n_n5331) & (x23x) & (!n_n5325) & (!n_n5333)) + ((x592x) & (!n_n5331) & (x23x) & (!n_n5325) & (n_n5333)) + ((x592x) & (!n_n5331) & (x23x) & (n_n5325) & (!n_n5333)) + ((x592x) & (!n_n5331) & (x23x) & (n_n5325) & (n_n5333)) + ((x592x) & (n_n5331) & (!x23x) & (!n_n5325) & (!n_n5333)) + ((x592x) & (n_n5331) & (!x23x) & (!n_n5325) & (n_n5333)) + ((x592x) & (n_n5331) & (!x23x) & (n_n5325) & (!n_n5333)) + ((x592x) & (n_n5331) & (!x23x) & (n_n5325) & (n_n5333)) + ((x592x) & (n_n5331) & (x23x) & (!n_n5325) & (!n_n5333)) + ((x592x) & (n_n5331) & (x23x) & (!n_n5325) & (n_n5333)) + ((x592x) & (n_n5331) & (x23x) & (n_n5325) & (!n_n5333)) + ((x592x) & (n_n5331) & (x23x) & (n_n5325) & (n_n5333)));
	assign x15938x = (((!n_n4371) & (!n_n4343) & (!n_n4362) & (!n_n4320) & (n_n4360)) + ((!n_n4371) & (!n_n4343) & (!n_n4362) & (n_n4320) & (!n_n4360)) + ((!n_n4371) & (!n_n4343) & (!n_n4362) & (n_n4320) & (n_n4360)) + ((!n_n4371) & (!n_n4343) & (n_n4362) & (!n_n4320) & (!n_n4360)) + ((!n_n4371) & (!n_n4343) & (n_n4362) & (!n_n4320) & (n_n4360)) + ((!n_n4371) & (!n_n4343) & (n_n4362) & (n_n4320) & (!n_n4360)) + ((!n_n4371) & (!n_n4343) & (n_n4362) & (n_n4320) & (n_n4360)) + ((!n_n4371) & (n_n4343) & (!n_n4362) & (!n_n4320) & (!n_n4360)) + ((!n_n4371) & (n_n4343) & (!n_n4362) & (!n_n4320) & (n_n4360)) + ((!n_n4371) & (n_n4343) & (!n_n4362) & (n_n4320) & (!n_n4360)) + ((!n_n4371) & (n_n4343) & (!n_n4362) & (n_n4320) & (n_n4360)) + ((!n_n4371) & (n_n4343) & (n_n4362) & (!n_n4320) & (!n_n4360)) + ((!n_n4371) & (n_n4343) & (n_n4362) & (!n_n4320) & (n_n4360)) + ((!n_n4371) & (n_n4343) & (n_n4362) & (n_n4320) & (!n_n4360)) + ((!n_n4371) & (n_n4343) & (n_n4362) & (n_n4320) & (n_n4360)) + ((n_n4371) & (!n_n4343) & (!n_n4362) & (!n_n4320) & (!n_n4360)) + ((n_n4371) & (!n_n4343) & (!n_n4362) & (!n_n4320) & (n_n4360)) + ((n_n4371) & (!n_n4343) & (!n_n4362) & (n_n4320) & (!n_n4360)) + ((n_n4371) & (!n_n4343) & (!n_n4362) & (n_n4320) & (n_n4360)) + ((n_n4371) & (!n_n4343) & (n_n4362) & (!n_n4320) & (!n_n4360)) + ((n_n4371) & (!n_n4343) & (n_n4362) & (!n_n4320) & (n_n4360)) + ((n_n4371) & (!n_n4343) & (n_n4362) & (n_n4320) & (!n_n4360)) + ((n_n4371) & (!n_n4343) & (n_n4362) & (n_n4320) & (n_n4360)) + ((n_n4371) & (n_n4343) & (!n_n4362) & (!n_n4320) & (!n_n4360)) + ((n_n4371) & (n_n4343) & (!n_n4362) & (!n_n4320) & (n_n4360)) + ((n_n4371) & (n_n4343) & (!n_n4362) & (n_n4320) & (!n_n4360)) + ((n_n4371) & (n_n4343) & (!n_n4362) & (n_n4320) & (n_n4360)) + ((n_n4371) & (n_n4343) & (n_n4362) & (!n_n4320) & (!n_n4360)) + ((n_n4371) & (n_n4343) & (n_n4362) & (!n_n4320) & (n_n4360)) + ((n_n4371) & (n_n4343) & (n_n4362) & (n_n4320) & (!n_n4360)) + ((n_n4371) & (n_n4343) & (n_n4362) & (n_n4320) & (n_n4360)));
	assign x22069x = (((!n_n5035) & (!n_n5032) & (!n_n5036) & (!n_n5037)));
	assign x16238x = (((!n_n4782) & (!n_n4788) & (!n_n4777) & (!n_n4204) & (n_n3469)) + ((!n_n4782) & (!n_n4788) & (!n_n4777) & (n_n4204) & (!n_n3469)) + ((!n_n4782) & (!n_n4788) & (!n_n4777) & (n_n4204) & (n_n3469)) + ((!n_n4782) & (!n_n4788) & (n_n4777) & (!n_n4204) & (!n_n3469)) + ((!n_n4782) & (!n_n4788) & (n_n4777) & (!n_n4204) & (n_n3469)) + ((!n_n4782) & (!n_n4788) & (n_n4777) & (n_n4204) & (!n_n3469)) + ((!n_n4782) & (!n_n4788) & (n_n4777) & (n_n4204) & (n_n3469)) + ((!n_n4782) & (n_n4788) & (!n_n4777) & (!n_n4204) & (!n_n3469)) + ((!n_n4782) & (n_n4788) & (!n_n4777) & (!n_n4204) & (n_n3469)) + ((!n_n4782) & (n_n4788) & (!n_n4777) & (n_n4204) & (!n_n3469)) + ((!n_n4782) & (n_n4788) & (!n_n4777) & (n_n4204) & (n_n3469)) + ((!n_n4782) & (n_n4788) & (n_n4777) & (!n_n4204) & (!n_n3469)) + ((!n_n4782) & (n_n4788) & (n_n4777) & (!n_n4204) & (n_n3469)) + ((!n_n4782) & (n_n4788) & (n_n4777) & (n_n4204) & (!n_n3469)) + ((!n_n4782) & (n_n4788) & (n_n4777) & (n_n4204) & (n_n3469)) + ((n_n4782) & (!n_n4788) & (!n_n4777) & (!n_n4204) & (!n_n3469)) + ((n_n4782) & (!n_n4788) & (!n_n4777) & (!n_n4204) & (n_n3469)) + ((n_n4782) & (!n_n4788) & (!n_n4777) & (n_n4204) & (!n_n3469)) + ((n_n4782) & (!n_n4788) & (!n_n4777) & (n_n4204) & (n_n3469)) + ((n_n4782) & (!n_n4788) & (n_n4777) & (!n_n4204) & (!n_n3469)) + ((n_n4782) & (!n_n4788) & (n_n4777) & (!n_n4204) & (n_n3469)) + ((n_n4782) & (!n_n4788) & (n_n4777) & (n_n4204) & (!n_n3469)) + ((n_n4782) & (!n_n4788) & (n_n4777) & (n_n4204) & (n_n3469)) + ((n_n4782) & (n_n4788) & (!n_n4777) & (!n_n4204) & (!n_n3469)) + ((n_n4782) & (n_n4788) & (!n_n4777) & (!n_n4204) & (n_n3469)) + ((n_n4782) & (n_n4788) & (!n_n4777) & (n_n4204) & (!n_n3469)) + ((n_n4782) & (n_n4788) & (!n_n4777) & (n_n4204) & (n_n3469)) + ((n_n4782) & (n_n4788) & (n_n4777) & (!n_n4204) & (!n_n3469)) + ((n_n4782) & (n_n4788) & (n_n4777) & (!n_n4204) & (n_n3469)) + ((n_n4782) & (n_n4788) & (n_n4777) & (n_n4204) & (!n_n3469)) + ((n_n4782) & (n_n4788) & (n_n4777) & (n_n4204) & (n_n3469)));
	assign x22077x = (((!n_n5146) & (!n_n5154) & (!n_n5150) & (!n_n5147)));
	assign x22060x = (((!n_n4779) & (!n_n4790) & (!n_n4776) & (!n_n4774)));
	assign x16408x = (((!i_7_) & (i_8_) & (!i_6_) & (n_n482) & (x10x)) + ((i_7_) & (!i_8_) & (!i_6_) & (n_n482) & (x10x)));
	assign x16421x = (((!i_9_) & (!n_n524) & (n_n325) & (n_n522) & (n_n500)) + ((!i_9_) & (n_n524) & (n_n325) & (!n_n522) & (n_n500)) + ((!i_9_) & (n_n524) & (n_n325) & (n_n522) & (n_n500)) + ((i_9_) & (!n_n524) & (n_n325) & (n_n522) & (n_n500)) + ((i_9_) & (n_n524) & (n_n325) & (!n_n522) & (n_n500)) + ((i_9_) & (n_n524) & (n_n325) & (n_n522) & (n_n500)));
	assign x16462x = (((!i_9_) & (!n_n524) & (n_n528) & (n_n535) & (n_n195)) + ((!i_9_) & (n_n524) & (!n_n528) & (n_n535) & (n_n195)) + ((!i_9_) & (n_n524) & (n_n528) & (n_n535) & (n_n195)));
	assign x16466x = (((!n_n4960) & (!n_n4964) & (!n_n3802) & (!x250x) & (x16462x)) + ((!n_n4960) & (!n_n4964) & (!n_n3802) & (x250x) & (!x16462x)) + ((!n_n4960) & (!n_n4964) & (!n_n3802) & (x250x) & (x16462x)) + ((!n_n4960) & (!n_n4964) & (n_n3802) & (!x250x) & (!x16462x)) + ((!n_n4960) & (!n_n4964) & (n_n3802) & (!x250x) & (x16462x)) + ((!n_n4960) & (!n_n4964) & (n_n3802) & (x250x) & (!x16462x)) + ((!n_n4960) & (!n_n4964) & (n_n3802) & (x250x) & (x16462x)) + ((!n_n4960) & (n_n4964) & (!n_n3802) & (!x250x) & (!x16462x)) + ((!n_n4960) & (n_n4964) & (!n_n3802) & (!x250x) & (x16462x)) + ((!n_n4960) & (n_n4964) & (!n_n3802) & (x250x) & (!x16462x)) + ((!n_n4960) & (n_n4964) & (!n_n3802) & (x250x) & (x16462x)) + ((!n_n4960) & (n_n4964) & (n_n3802) & (!x250x) & (!x16462x)) + ((!n_n4960) & (n_n4964) & (n_n3802) & (!x250x) & (x16462x)) + ((!n_n4960) & (n_n4964) & (n_n3802) & (x250x) & (!x16462x)) + ((!n_n4960) & (n_n4964) & (n_n3802) & (x250x) & (x16462x)) + ((n_n4960) & (!n_n4964) & (!n_n3802) & (!x250x) & (!x16462x)) + ((n_n4960) & (!n_n4964) & (!n_n3802) & (!x250x) & (x16462x)) + ((n_n4960) & (!n_n4964) & (!n_n3802) & (x250x) & (!x16462x)) + ((n_n4960) & (!n_n4964) & (!n_n3802) & (x250x) & (x16462x)) + ((n_n4960) & (!n_n4964) & (n_n3802) & (!x250x) & (!x16462x)) + ((n_n4960) & (!n_n4964) & (n_n3802) & (!x250x) & (x16462x)) + ((n_n4960) & (!n_n4964) & (n_n3802) & (x250x) & (!x16462x)) + ((n_n4960) & (!n_n4964) & (n_n3802) & (x250x) & (x16462x)) + ((n_n4960) & (n_n4964) & (!n_n3802) & (!x250x) & (!x16462x)) + ((n_n4960) & (n_n4964) & (!n_n3802) & (!x250x) & (x16462x)) + ((n_n4960) & (n_n4964) & (!n_n3802) & (x250x) & (!x16462x)) + ((n_n4960) & (n_n4964) & (!n_n3802) & (x250x) & (x16462x)) + ((n_n4960) & (n_n4964) & (n_n3802) & (!x250x) & (!x16462x)) + ((n_n4960) & (n_n4964) & (n_n3802) & (!x250x) & (x16462x)) + ((n_n4960) & (n_n4964) & (n_n3802) & (x250x) & (!x16462x)) + ((n_n4960) & (n_n4964) & (n_n3802) & (x250x) & (x16462x)));
	assign x16595x = (((!x13x) & (!n_n522) & (!n_n520) & (!n_n500) & (x387x)) + ((!x13x) & (!n_n522) & (!n_n520) & (n_n500) & (x387x)) + ((!x13x) & (!n_n522) & (n_n520) & (!n_n500) & (x387x)) + ((!x13x) & (!n_n522) & (n_n520) & (n_n500) & (x387x)) + ((!x13x) & (n_n522) & (!n_n520) & (!n_n500) & (x387x)) + ((!x13x) & (n_n522) & (!n_n520) & (n_n500) & (x387x)) + ((!x13x) & (n_n522) & (n_n520) & (!n_n500) & (x387x)) + ((!x13x) & (n_n522) & (n_n520) & (n_n500) & (x387x)) + ((x13x) & (!n_n522) & (!n_n520) & (!n_n500) & (x387x)) + ((x13x) & (!n_n522) & (!n_n520) & (n_n500) & (x387x)) + ((x13x) & (!n_n522) & (n_n520) & (!n_n500) & (x387x)) + ((x13x) & (!n_n522) & (n_n520) & (n_n500) & (!x387x)) + ((x13x) & (!n_n522) & (n_n520) & (n_n500) & (x387x)) + ((x13x) & (n_n522) & (!n_n520) & (!n_n500) & (x387x)) + ((x13x) & (n_n522) & (!n_n520) & (n_n500) & (!x387x)) + ((x13x) & (n_n522) & (!n_n520) & (n_n500) & (x387x)) + ((x13x) & (n_n522) & (n_n520) & (!n_n500) & (x387x)) + ((x13x) & (n_n522) & (n_n520) & (n_n500) & (!x387x)) + ((x13x) & (n_n522) & (n_n520) & (n_n500) & (x387x)));
	assign x16659x = (((!n_n5330) & (!n_n5331) & (!n_n5318) & (!n_n5320) & (n_n2274)) + ((!n_n5330) & (!n_n5331) & (!n_n5318) & (n_n5320) & (!n_n2274)) + ((!n_n5330) & (!n_n5331) & (!n_n5318) & (n_n5320) & (n_n2274)) + ((!n_n5330) & (!n_n5331) & (n_n5318) & (!n_n5320) & (!n_n2274)) + ((!n_n5330) & (!n_n5331) & (n_n5318) & (!n_n5320) & (n_n2274)) + ((!n_n5330) & (!n_n5331) & (n_n5318) & (n_n5320) & (!n_n2274)) + ((!n_n5330) & (!n_n5331) & (n_n5318) & (n_n5320) & (n_n2274)) + ((!n_n5330) & (n_n5331) & (!n_n5318) & (!n_n5320) & (!n_n2274)) + ((!n_n5330) & (n_n5331) & (!n_n5318) & (!n_n5320) & (n_n2274)) + ((!n_n5330) & (n_n5331) & (!n_n5318) & (n_n5320) & (!n_n2274)) + ((!n_n5330) & (n_n5331) & (!n_n5318) & (n_n5320) & (n_n2274)) + ((!n_n5330) & (n_n5331) & (n_n5318) & (!n_n5320) & (!n_n2274)) + ((!n_n5330) & (n_n5331) & (n_n5318) & (!n_n5320) & (n_n2274)) + ((!n_n5330) & (n_n5331) & (n_n5318) & (n_n5320) & (!n_n2274)) + ((!n_n5330) & (n_n5331) & (n_n5318) & (n_n5320) & (n_n2274)) + ((n_n5330) & (!n_n5331) & (!n_n5318) & (!n_n5320) & (!n_n2274)) + ((n_n5330) & (!n_n5331) & (!n_n5318) & (!n_n5320) & (n_n2274)) + ((n_n5330) & (!n_n5331) & (!n_n5318) & (n_n5320) & (!n_n2274)) + ((n_n5330) & (!n_n5331) & (!n_n5318) & (n_n5320) & (n_n2274)) + ((n_n5330) & (!n_n5331) & (n_n5318) & (!n_n5320) & (!n_n2274)) + ((n_n5330) & (!n_n5331) & (n_n5318) & (!n_n5320) & (n_n2274)) + ((n_n5330) & (!n_n5331) & (n_n5318) & (n_n5320) & (!n_n2274)) + ((n_n5330) & (!n_n5331) & (n_n5318) & (n_n5320) & (n_n2274)) + ((n_n5330) & (n_n5331) & (!n_n5318) & (!n_n5320) & (!n_n2274)) + ((n_n5330) & (n_n5331) & (!n_n5318) & (!n_n5320) & (n_n2274)) + ((n_n5330) & (n_n5331) & (!n_n5318) & (n_n5320) & (!n_n2274)) + ((n_n5330) & (n_n5331) & (!n_n5318) & (n_n5320) & (n_n2274)) + ((n_n5330) & (n_n5331) & (n_n5318) & (!n_n5320) & (!n_n2274)) + ((n_n5330) & (n_n5331) & (n_n5318) & (!n_n5320) & (n_n2274)) + ((n_n5330) & (n_n5331) & (n_n5318) & (n_n5320) & (!n_n2274)) + ((n_n5330) & (n_n5331) & (n_n5318) & (n_n5320) & (n_n2274)));
	assign x22058x = (((!n_n5321) & (!n_n5307) & (!n_n5326) & (!n_n5325)));
	assign x16660x = (((!n_n5310) & (!n_n5332) & (!n_n5329) & (!n_n5311) & (!x22058x)) + ((!n_n5310) & (!n_n5332) & (!n_n5329) & (n_n5311) & (!x22058x)) + ((!n_n5310) & (!n_n5332) & (!n_n5329) & (n_n5311) & (x22058x)) + ((!n_n5310) & (!n_n5332) & (n_n5329) & (!n_n5311) & (!x22058x)) + ((!n_n5310) & (!n_n5332) & (n_n5329) & (!n_n5311) & (x22058x)) + ((!n_n5310) & (!n_n5332) & (n_n5329) & (n_n5311) & (!x22058x)) + ((!n_n5310) & (!n_n5332) & (n_n5329) & (n_n5311) & (x22058x)) + ((!n_n5310) & (n_n5332) & (!n_n5329) & (!n_n5311) & (!x22058x)) + ((!n_n5310) & (n_n5332) & (!n_n5329) & (!n_n5311) & (x22058x)) + ((!n_n5310) & (n_n5332) & (!n_n5329) & (n_n5311) & (!x22058x)) + ((!n_n5310) & (n_n5332) & (!n_n5329) & (n_n5311) & (x22058x)) + ((!n_n5310) & (n_n5332) & (n_n5329) & (!n_n5311) & (!x22058x)) + ((!n_n5310) & (n_n5332) & (n_n5329) & (!n_n5311) & (x22058x)) + ((!n_n5310) & (n_n5332) & (n_n5329) & (n_n5311) & (!x22058x)) + ((!n_n5310) & (n_n5332) & (n_n5329) & (n_n5311) & (x22058x)) + ((n_n5310) & (!n_n5332) & (!n_n5329) & (!n_n5311) & (!x22058x)) + ((n_n5310) & (!n_n5332) & (!n_n5329) & (!n_n5311) & (x22058x)) + ((n_n5310) & (!n_n5332) & (!n_n5329) & (n_n5311) & (!x22058x)) + ((n_n5310) & (!n_n5332) & (!n_n5329) & (n_n5311) & (x22058x)) + ((n_n5310) & (!n_n5332) & (n_n5329) & (!n_n5311) & (!x22058x)) + ((n_n5310) & (!n_n5332) & (n_n5329) & (!n_n5311) & (x22058x)) + ((n_n5310) & (!n_n5332) & (n_n5329) & (n_n5311) & (!x22058x)) + ((n_n5310) & (!n_n5332) & (n_n5329) & (n_n5311) & (x22058x)) + ((n_n5310) & (n_n5332) & (!n_n5329) & (!n_n5311) & (!x22058x)) + ((n_n5310) & (n_n5332) & (!n_n5329) & (!n_n5311) & (x22058x)) + ((n_n5310) & (n_n5332) & (!n_n5329) & (n_n5311) & (!x22058x)) + ((n_n5310) & (n_n5332) & (!n_n5329) & (n_n5311) & (x22058x)) + ((n_n5310) & (n_n5332) & (n_n5329) & (!n_n5311) & (!x22058x)) + ((n_n5310) & (n_n5332) & (n_n5329) & (!n_n5311) & (x22058x)) + ((n_n5310) & (n_n5332) & (n_n5329) & (n_n5311) & (!x22058x)) + ((n_n5310) & (n_n5332) & (n_n5329) & (n_n5311) & (x22058x)));
	assign x22059x = (((!n_n5162) & (!n_n5166) & (!n_n5163) & (!n_n5169)));
	assign x16741x = (((!n_n5050) & (!n_n5049) & (!n_n5039) & (!n_n5029) & (x153x)) + ((!n_n5050) & (!n_n5049) & (!n_n5039) & (n_n5029) & (!x153x)) + ((!n_n5050) & (!n_n5049) & (!n_n5039) & (n_n5029) & (x153x)) + ((!n_n5050) & (!n_n5049) & (n_n5039) & (!n_n5029) & (!x153x)) + ((!n_n5050) & (!n_n5049) & (n_n5039) & (!n_n5029) & (x153x)) + ((!n_n5050) & (!n_n5049) & (n_n5039) & (n_n5029) & (!x153x)) + ((!n_n5050) & (!n_n5049) & (n_n5039) & (n_n5029) & (x153x)) + ((!n_n5050) & (n_n5049) & (!n_n5039) & (!n_n5029) & (!x153x)) + ((!n_n5050) & (n_n5049) & (!n_n5039) & (!n_n5029) & (x153x)) + ((!n_n5050) & (n_n5049) & (!n_n5039) & (n_n5029) & (!x153x)) + ((!n_n5050) & (n_n5049) & (!n_n5039) & (n_n5029) & (x153x)) + ((!n_n5050) & (n_n5049) & (n_n5039) & (!n_n5029) & (!x153x)) + ((!n_n5050) & (n_n5049) & (n_n5039) & (!n_n5029) & (x153x)) + ((!n_n5050) & (n_n5049) & (n_n5039) & (n_n5029) & (!x153x)) + ((!n_n5050) & (n_n5049) & (n_n5039) & (n_n5029) & (x153x)) + ((n_n5050) & (!n_n5049) & (!n_n5039) & (!n_n5029) & (!x153x)) + ((n_n5050) & (!n_n5049) & (!n_n5039) & (!n_n5029) & (x153x)) + ((n_n5050) & (!n_n5049) & (!n_n5039) & (n_n5029) & (!x153x)) + ((n_n5050) & (!n_n5049) & (!n_n5039) & (n_n5029) & (x153x)) + ((n_n5050) & (!n_n5049) & (n_n5039) & (!n_n5029) & (!x153x)) + ((n_n5050) & (!n_n5049) & (n_n5039) & (!n_n5029) & (x153x)) + ((n_n5050) & (!n_n5049) & (n_n5039) & (n_n5029) & (!x153x)) + ((n_n5050) & (!n_n5049) & (n_n5039) & (n_n5029) & (x153x)) + ((n_n5050) & (n_n5049) & (!n_n5039) & (!n_n5029) & (!x153x)) + ((n_n5050) & (n_n5049) & (!n_n5039) & (!n_n5029) & (x153x)) + ((n_n5050) & (n_n5049) & (!n_n5039) & (n_n5029) & (!x153x)) + ((n_n5050) & (n_n5049) & (!n_n5039) & (n_n5029) & (x153x)) + ((n_n5050) & (n_n5049) & (n_n5039) & (!n_n5029) & (!x153x)) + ((n_n5050) & (n_n5049) & (n_n5039) & (!n_n5029) & (x153x)) + ((n_n5050) & (n_n5049) & (n_n5039) & (n_n5029) & (!x153x)) + ((n_n5050) & (n_n5049) & (n_n5039) & (n_n5029) & (x153x)));
	assign x16761x = (((!x20x) & (!x23x) & (!n_n464) & (!n_n65) & (n_n5334)) + ((!x20x) & (!x23x) & (!n_n464) & (n_n65) & (n_n5334)) + ((!x20x) & (!x23x) & (n_n464) & (!n_n65) & (n_n5334)) + ((!x20x) & (!x23x) & (n_n464) & (n_n65) & (n_n5334)) + ((!x20x) & (x23x) & (!n_n464) & (!n_n65) & (n_n5334)) + ((!x20x) & (x23x) & (!n_n464) & (n_n65) & (n_n5334)) + ((!x20x) & (x23x) & (n_n464) & (!n_n65) & (n_n5334)) + ((!x20x) & (x23x) & (n_n464) & (n_n65) & (!n_n5334)) + ((!x20x) & (x23x) & (n_n464) & (n_n65) & (n_n5334)) + ((x20x) & (!x23x) & (!n_n464) & (!n_n65) & (n_n5334)) + ((x20x) & (!x23x) & (!n_n464) & (n_n65) & (n_n5334)) + ((x20x) & (!x23x) & (n_n464) & (!n_n65) & (n_n5334)) + ((x20x) & (!x23x) & (n_n464) & (n_n65) & (!n_n5334)) + ((x20x) & (!x23x) & (n_n464) & (n_n65) & (n_n5334)) + ((x20x) & (x23x) & (!n_n464) & (!n_n65) & (n_n5334)) + ((x20x) & (x23x) & (!n_n464) & (n_n65) & (n_n5334)) + ((x20x) & (x23x) & (n_n464) & (!n_n65) & (n_n5334)) + ((x20x) & (x23x) & (n_n464) & (n_n65) & (!n_n5334)) + ((x20x) & (x23x) & (n_n464) & (n_n65) & (n_n5334)));
	assign x16818x = (((!n_n4934) & (!n_n4938) & (!n_n4947) & (n_n4940)) + ((!n_n4934) & (!n_n4938) & (n_n4947) & (!n_n4940)) + ((!n_n4934) & (!n_n4938) & (n_n4947) & (n_n4940)) + ((!n_n4934) & (n_n4938) & (!n_n4947) & (!n_n4940)) + ((!n_n4934) & (n_n4938) & (!n_n4947) & (n_n4940)) + ((!n_n4934) & (n_n4938) & (n_n4947) & (!n_n4940)) + ((!n_n4934) & (n_n4938) & (n_n4947) & (n_n4940)) + ((n_n4934) & (!n_n4938) & (!n_n4947) & (!n_n4940)) + ((n_n4934) & (!n_n4938) & (!n_n4947) & (n_n4940)) + ((n_n4934) & (!n_n4938) & (n_n4947) & (!n_n4940)) + ((n_n4934) & (!n_n4938) & (n_n4947) & (n_n4940)) + ((n_n4934) & (n_n4938) & (!n_n4947) & (!n_n4940)) + ((n_n4934) & (n_n4938) & (!n_n4947) & (n_n4940)) + ((n_n4934) & (n_n4938) & (n_n4947) & (!n_n4940)) + ((n_n4934) & (n_n4938) & (n_n4947) & (n_n4940)));
	assign x16819x = (((!n_n4912) & (!n_n4931) & (!n_n4932) & (!n_n4944) & (n_n4910)) + ((!n_n4912) & (!n_n4931) & (!n_n4932) & (n_n4944) & (!n_n4910)) + ((!n_n4912) & (!n_n4931) & (!n_n4932) & (n_n4944) & (n_n4910)) + ((!n_n4912) & (!n_n4931) & (n_n4932) & (!n_n4944) & (!n_n4910)) + ((!n_n4912) & (!n_n4931) & (n_n4932) & (!n_n4944) & (n_n4910)) + ((!n_n4912) & (!n_n4931) & (n_n4932) & (n_n4944) & (!n_n4910)) + ((!n_n4912) & (!n_n4931) & (n_n4932) & (n_n4944) & (n_n4910)) + ((!n_n4912) & (n_n4931) & (!n_n4932) & (!n_n4944) & (!n_n4910)) + ((!n_n4912) & (n_n4931) & (!n_n4932) & (!n_n4944) & (n_n4910)) + ((!n_n4912) & (n_n4931) & (!n_n4932) & (n_n4944) & (!n_n4910)) + ((!n_n4912) & (n_n4931) & (!n_n4932) & (n_n4944) & (n_n4910)) + ((!n_n4912) & (n_n4931) & (n_n4932) & (!n_n4944) & (!n_n4910)) + ((!n_n4912) & (n_n4931) & (n_n4932) & (!n_n4944) & (n_n4910)) + ((!n_n4912) & (n_n4931) & (n_n4932) & (n_n4944) & (!n_n4910)) + ((!n_n4912) & (n_n4931) & (n_n4932) & (n_n4944) & (n_n4910)) + ((n_n4912) & (!n_n4931) & (!n_n4932) & (!n_n4944) & (!n_n4910)) + ((n_n4912) & (!n_n4931) & (!n_n4932) & (!n_n4944) & (n_n4910)) + ((n_n4912) & (!n_n4931) & (!n_n4932) & (n_n4944) & (!n_n4910)) + ((n_n4912) & (!n_n4931) & (!n_n4932) & (n_n4944) & (n_n4910)) + ((n_n4912) & (!n_n4931) & (n_n4932) & (!n_n4944) & (!n_n4910)) + ((n_n4912) & (!n_n4931) & (n_n4932) & (!n_n4944) & (n_n4910)) + ((n_n4912) & (!n_n4931) & (n_n4932) & (n_n4944) & (!n_n4910)) + ((n_n4912) & (!n_n4931) & (n_n4932) & (n_n4944) & (n_n4910)) + ((n_n4912) & (n_n4931) & (!n_n4932) & (!n_n4944) & (!n_n4910)) + ((n_n4912) & (n_n4931) & (!n_n4932) & (!n_n4944) & (n_n4910)) + ((n_n4912) & (n_n4931) & (!n_n4932) & (n_n4944) & (!n_n4910)) + ((n_n4912) & (n_n4931) & (!n_n4932) & (n_n4944) & (n_n4910)) + ((n_n4912) & (n_n4931) & (n_n4932) & (!n_n4944) & (!n_n4910)) + ((n_n4912) & (n_n4931) & (n_n4932) & (!n_n4944) & (n_n4910)) + ((n_n4912) & (n_n4931) & (n_n4932) & (n_n4944) & (!n_n4910)) + ((n_n4912) & (n_n4931) & (n_n4932) & (n_n4944) & (n_n4910)));
	assign x16821x = (((!x16778x) & (!x16779x) & (n_n2095)) + ((!x16778x) & (x16779x) & (!n_n2095)) + ((!x16778x) & (x16779x) & (n_n2095)) + ((x16778x) & (!x16779x) & (!n_n2095)) + ((x16778x) & (!x16779x) & (n_n2095)) + ((x16778x) & (x16779x) & (!n_n2095)) + ((x16778x) & (x16779x) & (n_n2095)));
	assign x16822x = (((!x16812x) & (!x16813x) & (!x16818x) & (x16819x)) + ((!x16812x) & (!x16813x) & (x16818x) & (!x16819x)) + ((!x16812x) & (!x16813x) & (x16818x) & (x16819x)) + ((!x16812x) & (x16813x) & (!x16818x) & (!x16819x)) + ((!x16812x) & (x16813x) & (!x16818x) & (x16819x)) + ((!x16812x) & (x16813x) & (x16818x) & (!x16819x)) + ((!x16812x) & (x16813x) & (x16818x) & (x16819x)) + ((x16812x) & (!x16813x) & (!x16818x) & (!x16819x)) + ((x16812x) & (!x16813x) & (!x16818x) & (x16819x)) + ((x16812x) & (!x16813x) & (x16818x) & (!x16819x)) + ((x16812x) & (!x16813x) & (x16818x) & (x16819x)) + ((x16812x) & (x16813x) & (!x16818x) & (!x16819x)) + ((x16812x) & (x16813x) & (!x16818x) & (x16819x)) + ((x16812x) & (x16813x) & (x16818x) & (!x16819x)) + ((x16812x) & (x16813x) & (x16818x) & (x16819x)));
	assign x16824x = (((!x16476x) & (!x16477x) & (!x16651x) & (x16652x)) + ((!x16476x) & (!x16477x) & (x16651x) & (!x16652x)) + ((!x16476x) & (!x16477x) & (x16651x) & (x16652x)) + ((!x16476x) & (x16477x) & (!x16651x) & (!x16652x)) + ((!x16476x) & (x16477x) & (!x16651x) & (x16652x)) + ((!x16476x) & (x16477x) & (x16651x) & (!x16652x)) + ((!x16476x) & (x16477x) & (x16651x) & (x16652x)) + ((x16476x) & (!x16477x) & (!x16651x) & (!x16652x)) + ((x16476x) & (!x16477x) & (!x16651x) & (x16652x)) + ((x16476x) & (!x16477x) & (x16651x) & (!x16652x)) + ((x16476x) & (!x16477x) & (x16651x) & (x16652x)) + ((x16476x) & (x16477x) & (!x16651x) & (!x16652x)) + ((x16476x) & (x16477x) & (!x16651x) & (x16652x)) + ((x16476x) & (x16477x) & (x16651x) & (!x16652x)) + ((x16476x) & (x16477x) & (x16651x) & (x16652x)));

endmodule