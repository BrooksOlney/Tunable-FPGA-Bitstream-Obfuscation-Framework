module apex4_qmap_map (sk, i_0_, i_1_, i_2_, i_6_, i_7_, i_8_, i_3_, i_4_, i_5_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_);

	input i_0_;
	input i_1_;
	input i_2_;
	input i_6_;
	input i_7_;
	input i_8_;
	input i_3_;
	input i_4_;
	input i_5_;
	output o_0_;
	output o_1_;
	output o_2_;
	output o_3_;
	output o_4_;
	output o_5_;
	output o_6_;
	output o_7_;
	output o_8_;
	output o_9_;
	output o_10_;
	output o_11_;
	output o_12_;
	output o_13_;
	output o_14_;
	output o_15_;
	output o_16_;
	output o_17_;
	output o_18_;



	wire gnd, g82, g199, g263, g320, g356, g395, g418, g437, g454, g467, g490, g510, g520, g523, g532, g537, g540, g542, g1, g2;
	wire g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23;
	wire g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44;
	wire g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65;
	wire g66, g67, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g79, g80, g81, g83, g84, g85, g86, g87;
	wire g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106, g107, g108;
	wire g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129;
	wire g130, g131, g683, g132, g694, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147, g148;
	wire g149, g150, g151, g152, g670, g153, g154, g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g168;
	wire g169, g170, g171, g172, g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189;
	wire g190, g657, g191, g192, g193, g194, g195, g196, g197, g198, g200, g201, g202, g203, g204, g205, g206, g207, g208, g209, g644;
	wire g210, g211, g212, g213, g214, g215, g216, g217, g218, g219, g220, g221, g222, g223, g224, g225, g226, g227, g228, g229, g230;
	wire g231, g232, g631, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250;
	wire g251, g252, g253, g254, g255, g256, g257, g258, g259, g260, g261, g262, g264, g265, g266, g267, g268, g269, g270, g271, g272;
	wire g273, g274, g275, g276, g277, g278, g279, g280, g281, g282, g283, g284, g285, g286, g287, g288, g289, g290, g291, g292, g293;
	wire g294, g295, g296, g297, g298, g299, g300, g301, g302, g303, g304, g305, g607, g306, g307, g308, g309, g310, g311, g312, g313;
	wire g314, g315, g316, g317, g318, g319, g618, g321, g322, g596, g323, g324, g325, g326, g327, g328, g329, g330, g331, g332, g333;
	wire g334, g335, g336, g337, g338, g339, g340, g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351, g352, g353, g354;
	wire g355, g357, g358, g359, g360, g361, g362, g363, g364, g365, g366, g367, g368, g369, g370, g371, g372, g373, g374, g375, g376;
	wire g377, g378, g379, g380, g381, g382, g383, g384, g385, g386, g387, g388, g389, g390, g391, g392, g583, g393, g394, g396, g397;
	wire g398, g399, g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410, g411, g412, g413, g414, g415, g416, g417, g419;
	wire g420, g421, g422, g572, g423, g424, g425, g426, g427, g428, g429, g430, g431, g432, g433, g434, g435, g436, g438, g439, g440;
	wire g441, g442, g443, g444, g445, g446, g447, g448, g449, g559, g450, g451, g452, g453, g455, g456, g457, g458, g459, g460, g461;
	wire g462, g463, g464, g465, g466, g468, g469, g470, g471, g472, g473, g474, g475, g476, g477, g478, g549, g479, g480, g481, g482;
	wire g483, g484, g485, g486, g487, g488, g489, g491, g492, g493, g494, g495, g496, g497, g498, g499, g500, g501, g502, g503, g504;
	wire g505, g506, g507, g508, g509, g511, g512, g513, g514, g515, g516, g517, g543, g518, g519, g521, g522, g524, g525, g526, g527;
	wire g528, g529, g530, g531, g533, g534, g535, g536, g538, g539, g541, g544, g545, g546, g547, g548, g550, g551, g552, g554, g553;
	wire g555, g556, g557, g558, g560, g561, g562, g565, g563, g564, g568, g569, g566, g567, g570, g571, g573, g574, g575, g578, g576;
	wire g577, g580, g581, g579, g582, g584, g585, g586, g589, g587, g588, g592, g593, g590, g591, g594, g595, g597, g598, g599, g601;
	wire g600, g604, g602, g603, g605, g606, g608, g609, g610, g612, g611, g615, g613, g614, g616, g617, g619, g620, g621, g624, g622;
	wire g623, g627, g628, g625, g626, g629, g630, g632, g633, g634, g637, g635, g636, g640, g641, g638, g639, g642, g643, g645, g646;
	wire g647, g650, g648, g649, g653, g654, g651, g652, g655, g656, g658, g659, g660, g663, g661, g662, g666, g667, g664, g665, g668;
	wire g669, g671, g672, g673, g676, g674, g675, g679, g680, g677, g678, g681, g682, g684, g685, g686, g689, g687, g688, g691, g692;
	wire g690, g693, g695, g696, g697, g699, g698, g702, g700, g701, g703, g704;

	lut_sub lut_4 ({gnd}, o_0_);
	defparam lut_4.LUT_SIZE = 1;
	defparam lut_4.mask = 2'b01;

	lut_sub lut_7 ({g82}, o_1_);
	defparam lut_7.LUT_SIZE = 1;
	defparam lut_7.mask = 2'b10;

	lut_sub lut_11 ({g199}, o_2_);
	defparam lut_11.LUT_SIZE = 1;
	defparam lut_11.mask = 2'b10;

	lut_sub lut_15 ({g263}, o_3_);
	defparam lut_15.LUT_SIZE = 1;
	defparam lut_15.mask = 2'b10;

	lut_sub lut_19 ({g320}, o_4_);
	defparam lut_19.LUT_SIZE = 1;
	defparam lut_19.mask = 2'b10;

	lut_sub lut_23 ({g356}, o_5_);
	defparam lut_23.LUT_SIZE = 1;
	defparam lut_23.mask = 2'b10;

	lut_sub lut_27 ({g395}, o_6_);
	defparam lut_27.LUT_SIZE = 1;
	defparam lut_27.mask = 2'b10;

	lut_sub lut_31 ({g418}, o_7_);
	defparam lut_31.LUT_SIZE = 1;
	defparam lut_31.mask = 2'b10;

	lut_sub lut_35 ({g437}, o_8_);
	defparam lut_35.LUT_SIZE = 1;
	defparam lut_35.mask = 2'b10;

	lut_sub lut_39 ({g454}, o_9_);
	defparam lut_39.LUT_SIZE = 1;
	defparam lut_39.mask = 2'b10;

	lut_sub lut_43 ({g467}, o_10_);
	defparam lut_43.LUT_SIZE = 1;
	defparam lut_43.mask = 2'b10;

	lut_sub lut_47 ({g490}, o_11_);
	defparam lut_47.LUT_SIZE = 1;
	defparam lut_47.mask = 2'b10;

	lut_sub lut_51 ({g510}, o_12_);
	defparam lut_51.LUT_SIZE = 1;
	defparam lut_51.mask = 2'b10;

	lut_sub lut_55 ({g520}, o_13_);
	defparam lut_55.LUT_SIZE = 1;
	defparam lut_55.mask = 2'b10;

	lut_sub lut_59 ({g523}, o_14_);
	defparam lut_59.LUT_SIZE = 1;
	defparam lut_59.mask = 2'b10;

	lut_sub lut_63 ({g532}, o_15_);
	defparam lut_63.LUT_SIZE = 1;
	defparam lut_63.mask = 2'b10;

	lut_sub lut_67 ({g537}, o_16_);
	defparam lut_67.LUT_SIZE = 1;
	defparam lut_67.mask = 2'b10;

	lut_sub lut_71 ({g540}, o_17_);
	defparam lut_71.LUT_SIZE = 1;
	defparam lut_71.mask = 2'b10;

	lut_sub lut_75 ({g542}, o_18_);
	defparam lut_75.LUT_SIZE = 1;
	defparam lut_75.mask = 2'b10;

	lut_sub lut_79 ({i_0_, i_1_, i_2_}, g1);
	defparam lut_79.LUT_SIZE = 3;
	defparam lut_79.mask = 8'hf7;

	lut_sub lut_89 ({i_6_, i_7_, i_8_}, g2);
	defparam lut_89.LUT_SIZE = 3;
	defparam lut_89.mask = 8'h08;

	lut_sub lut_93 ({i_3_, i_4_, i_5_}, g3);
	defparam lut_93.LUT_SIZE = 3;
	defparam lut_93.mask = 8'h20;

	lut_sub lut_99 ({g2, g3}, g4);
	defparam lut_99.LUT_SIZE = 2;
	defparam lut_99.mask = 4'b0001;

	lut_sub lut_103 ({i_3_, i_4_}, g5);
	defparam lut_103.LUT_SIZE = 2;
	defparam lut_103.mask = 4'b0100;

	lut_sub lut_107 ({i_6_, i_7_, i_8_}, g6);
	defparam lut_107.LUT_SIZE = 3;
	defparam lut_107.mask = 8'h04;

	lut_sub lut_113 ({g1, g6}, g7);
	defparam lut_113.LUT_SIZE = 2;
	defparam lut_113.mask = 4'b0100;

	lut_sub lut_117 ({i_6_, i_7_, i_8_}, g8);
	defparam lut_117.LUT_SIZE = 3;
	defparam lut_117.mask = 8'h10;

	lut_sub lut_123 ({g8, g1}, g9);
	defparam lut_123.LUT_SIZE = 2;
	defparam lut_123.mask = 4'b0010;

	lut_sub lut_130 ({i_5_, g5, g7, g9}, g10);
	defparam lut_130.LUT_SIZE = 4;
	defparam lut_130.mask = 16'h0503;

	lut_sub lut_137 ({i_3_, i_4_, i_5_}, g11);
	defparam lut_137.LUT_SIZE = 3;
	defparam lut_137.mask = 8'hbf;

	lut_sub lut_147 ({i_6_, i_7_, i_8_}, g12);
	defparam lut_147.LUT_SIZE = 3;
	defparam lut_147.mask = 8'h20;

	lut_sub lut_151 ({i_0_, i_1_, i_2_}, g13);
	defparam lut_151.LUT_SIZE = 3;
	defparam lut_151.mask = 8'hfd;

	lut_sub lut_161 ({i_7_, i_8_}, g14);
	defparam lut_161.LUT_SIZE = 2;
	defparam lut_161.mask = 4'b0001;

	lut_sub lut_165 ({i_4_, i_5_, i_6_}, g15);
	defparam lut_165.LUT_SIZE = 3;
	defparam lut_165.mask = 8'h02;

	lut_sub lut_171 ({g14, g15}, g16);
	defparam lut_171.LUT_SIZE = 2;
	defparam lut_171.mask = 4'b0001;

	lut_sub lut_175 ({i_3_, i_0_, i_2_}, g17);
	defparam lut_175.LUT_SIZE = 3;
	defparam lut_175.mask = 8'h02;

	lut_sub lut_181 ({g16, g17}, g18);
	defparam lut_181.LUT_SIZE = 2;
	defparam lut_181.mask = 4'b0001;

	lut_sub lut_189 ({g11, g12, g13, g18}, g19);
	defparam lut_189.LUT_SIZE = 4;
	defparam lut_189.mask = 16'ha2aa;

	lut_sub lut_203 ({g1, g4, g10, g19}, g20);
	defparam lut_203.LUT_SIZE = 4;
	defparam lut_203.mask = 16'h4044;

	lut_sub lut_209 ({i_3_, i_4_, i_5_}, g21);
	defparam lut_209.LUT_SIZE = 3;
	defparam lut_209.mask = 8'hfb;

	lut_sub lut_221 ({g21, g2}, g22);
	defparam lut_221.LUT_SIZE = 2;
	defparam lut_221.mask = 4'b0100;

	lut_sub lut_225 ({i_6_, i_7_, i_8_}, g23);
	defparam lut_225.LUT_SIZE = 3;
	defparam lut_225.mask = 8'hfd;

	lut_sub lut_235 ({i_0_, i_1_, i_2_}, g24);
	defparam lut_235.LUT_SIZE = 3;
	defparam lut_235.mask = 8'hef;

	lut_sub lut_245 ({i_0_, i_1_, i_2_}, g25);
	defparam lut_245.LUT_SIZE = 3;
	defparam lut_245.mask = 8'hdf;

	lut_sub lut_257 ({g11, g25}, g26);
	defparam lut_257.LUT_SIZE = 2;
	defparam lut_257.mask = 4'b1000;

	lut_sub lut_261 ({i_0_, i_1_, i_2_}, g27);
	defparam lut_261.LUT_SIZE = 3;
	defparam lut_261.mask = 8'hfe;

	lut_sub lut_271 ({i_6_, i_7_, i_8_}, g28);
	defparam lut_271.LUT_SIZE = 3;
	defparam lut_271.mask = 8'h01;

	lut_sub lut_277 ({g28, g1}, g29);
	defparam lut_277.LUT_SIZE = 2;
	defparam lut_277.mask = 4'b0010;

	lut_sub lut_286 ({g11, g27, g21, g6, g29}, g30);
	defparam lut_286.LUT_SIZE = 5;
	defparam lut_286.mask = 32'h73505050;

	lut_sub lut_305 ({g22, g23, g24, g26, g30}, g31);
	defparam lut_305.LUT_SIZE = 5;
	defparam lut_305.mask = 32'h88aa080a;

	lut_sub lut_317 ({i_3_, i_4_, i_5_}, g32);
	defparam lut_317.LUT_SIZE = 3;
	defparam lut_317.mask = 8'h80;

	lut_sub lut_323 ({g24, g3}, g33);
	defparam lut_323.LUT_SIZE = 2;
	defparam lut_323.mask = 4'b0100;

	lut_sub lut_333 ({g11, g27, g6, g23, g32, g33}, g34);
	defparam lut_333.LUT_SIZE = 6;
	defparam lut_333.mask = 64'hf0f3505050735050;

	lut_sub lut_361 ({i_6_, i_7_, i_8_}, g35);
	defparam lut_361.LUT_SIZE = 3;
	defparam lut_361.mask = 8'h80;

	lut_sub lut_365 ({i_3_, i_4_, i_5_}, g36);
	defparam lut_365.LUT_SIZE = 3;
	defparam lut_365.mask = 8'hf7;

	lut_sub lut_375 ({i_6_, i_7_}, g37);
	defparam lut_375.LUT_SIZE = 2;
	defparam lut_375.mask = 4'b1000;

	lut_sub lut_379 ({i_3_, i_4_, i_5_}, g38);
	defparam lut_379.LUT_SIZE = 3;
	defparam lut_379.mask = 8'hef;

	lut_sub lut_394 ({g11, g27, g2, g37, g38}, g39);
	defparam lut_394.LUT_SIZE = 5;
	defparam lut_394.mask = 32'h2f002200;

	lut_sub lut_408 ({g35, g1, g36, g39}, g40);
	defparam lut_408.LUT_SIZE = 4;
	defparam lut_408.mask = 16'haa2a;

	lut_sub lut_420 ({g27, g35}, g41);
	defparam lut_420.LUT_SIZE = 2;
	defparam lut_420.mask = 4'b0100;

	lut_sub lut_424 ({i_0_, i_1_, i_2_}, g42);
	defparam lut_424.LUT_SIZE = 3;
	defparam lut_424.mask = 8'h04;

	lut_sub lut_431 ({g21, g28, g42}, g43);
	defparam lut_431.LUT_SIZE = 3;
	defparam lut_431.mask = 8'h10;

	lut_sub lut_439 ({g11, g41, g43, g3}, g44);
	defparam lut_439.LUT_SIZE = 4;
	defparam lut_439.mask = 16'hc0c8;

	lut_sub lut_447 ({i_3_, i_4_, i_5_}, g45);
	defparam lut_447.LUT_SIZE = 3;
	defparam lut_447.mask = 8'hfd;

	lut_sub lut_459 ({g25, g45}, g46);
	defparam lut_459.LUT_SIZE = 2;
	defparam lut_459.mask = 4'b1000;

	lut_sub lut_463 ({i_7_, i_8_}, g47);
	defparam lut_463.LUT_SIZE = 2;
	defparam lut_463.mask = 4'b0100;

	lut_sub lut_468 ({i_6_, g47}, g48);
	defparam lut_468.LUT_SIZE = 2;
	defparam lut_468.mask = 4'b0100;

	lut_sub lut_474 ({g32, g13}, g49);
	defparam lut_474.LUT_SIZE = 2;
	defparam lut_474.mask = 4'b0010;

	lut_sub lut_478 ({i_4_, i_5_}, g50);
	defparam lut_478.LUT_SIZE = 2;
	defparam lut_478.mask = 4'b0100;

	lut_sub lut_482 ({i_3_, i_0_, i_2_}, g51);
	defparam lut_482.LUT_SIZE = 3;
	defparam lut_482.mask = 8'h20;

	lut_sub lut_488 ({g50, g51}, g52);
	defparam lut_488.LUT_SIZE = 2;
	defparam lut_488.mask = 4'b0001;

	lut_sub lut_497 ({g8, g46, g48, g49, g52}, g53);
	defparam lut_497.LUT_SIZE = 5;
	defparam lut_497.mask = 32'hf8f8f800;

	lut_sub lut_515 ({i_4_, i_5_, i_6_, i_7_, i_8_}, g54);
	defparam lut_515.LUT_SIZE = 5;
	defparam lut_515.mask = 32'h40422020;

	lut_sub lut_528 ({g50, g42, g1, g12, g22}, g55);
	defparam lut_528.LUT_SIZE = 5;
	defparam lut_528.mask = 32'h00553075;

	lut_sub lut_545 ({i_3_, g1, g54, g55}, g56);
	defparam lut_545.LUT_SIZE = 4;
	defparam lut_545.mask = 16'haa8a;

	lut_sub lut_555 ({i_3_, i_1_, i_2_}, g57);
	defparam lut_555.LUT_SIZE = 3;
	defparam lut_555.mask = 8'h04;

	lut_sub lut_561 ({i_4_, i_5_, g57, g6}, g58);
	defparam lut_561.LUT_SIZE = 4;
	defparam lut_561.mask = 16'h0001;

	lut_sub lut_565 ({i_3_, i_4_, i_5_}, g59);
	defparam lut_565.LUT_SIZE = 3;
	defparam lut_565.mask = 8'hfe;

	lut_sub lut_575 ({i_6_, i_7_}, g60);
	defparam lut_575.LUT_SIZE = 2;
	defparam lut_575.mask = 4'b0001;

	lut_sub lut_584 ({g42, g58, g59, g13, g60}, g61);
	defparam lut_584.LUT_SIZE = 5;
	defparam lut_584.mask = 32'hbf00af00;

	lut_sub lut_605 ({g40, g44, g53, g56, g61}, g62);
	defparam lut_605.LUT_SIZE = 5;
	defparam lut_605.mask = 32'h00000001;

	lut_sub lut_609 ({i_7_, i_8_}, g63);
	defparam lut_609.LUT_SIZE = 2;
	defparam lut_609.mask = 4'b1000;

	lut_sub lut_613 ({i_4_, i_5_, i_6_}, g64);
	defparam lut_613.LUT_SIZE = 3;
	defparam lut_613.mask = 8'h08;

	lut_sub lut_618 ({i_3_, i_0_, i_1_, g64}, g65);
	defparam lut_618.LUT_SIZE = 4;
	defparam lut_618.mask = 16'h0004;

	lut_sub lut_627 ({g42, g45, g23, g36, g29}, g66);
	defparam lut_627.LUT_SIZE = 5;
	defparam lut_627.mask = 32'h4444f444;

	lut_sub lut_643 ({g27, g2}, g67);
	defparam lut_643.LUT_SIZE = 2;
	defparam lut_643.mask = 4'b0100;

	lut_sub lut_652 ({g1, g23, g32, g36, g67}, g68);
	defparam lut_652.LUT_SIZE = 5;
	defparam lut_652.mask = 32'hcd050505;

	lut_sub lut_670 ({g42, g45, g6, g68}, g69);
	defparam lut_670.LUT_SIZE = 4;
	defparam lut_670.mask = 16'haa8a;

	lut_sub lut_682 ({g25, g32}, g70);
	defparam lut_682.LUT_SIZE = 2;
	defparam lut_682.mask = 4'b0100;

	lut_sub lut_688 ({g42, g59}, g71);
	defparam lut_688.LUT_SIZE = 2;
	defparam lut_688.mask = 4'b0010;

	lut_sub lut_697 ({g27, g28, g32, g37, g71}, g72);
	defparam lut_697.LUT_SIZE = 5;
	defparam lut_697.mask = 32'h111f1111;

	lut_sub lut_713 ({g11, g24}, g73);
	defparam lut_713.LUT_SIZE = 2;
	defparam lut_713.mask = 4'b1000;

	lut_sub lut_720 ({g6, g24, g32}, g74);
	defparam lut_720.LUT_SIZE = 3;
	defparam lut_720.mask = 8'h04;

	lut_sub lut_726 ({g24, g59}, g75);
	defparam lut_726.LUT_SIZE = 2;
	defparam lut_726.mask = 4'b1000;

	lut_sub lut_734 ({g23, g73, g74, g75}, g76);
	defparam lut_734.LUT_SIZE = 4;
	defparam lut_734.mask = 16'h80cc;

	lut_sub lut_744 ({g25, g59}, g77);
	defparam lut_744.LUT_SIZE = 2;
	defparam lut_744.mask = 4'b1000;

	lut_sub lut_752 ({g28, g2, g77, g33}, g78);
	defparam lut_752.LUT_SIZE = 4;
	defparam lut_752.mask = 16'h0357;

	lut_sub lut_767 ({g6, g70, g72, g76, g78}, g79);
	defparam lut_767.LUT_SIZE = 5;
	defparam lut_767.mask = 32'h20202000;

	lut_sub lut_778 ({g21, g8, g24, g69, g79}, g80);
	defparam lut_778.LUT_SIZE = 5;
	defparam lut_778.mask = 32'h11011111;

	lut_sub lut_792 ({g63, g65, g66, g80}, g81);
	defparam lut_792.LUT_SIZE = 4;
	defparam lut_792.mask = 16'h4440;

	lut_sub lut_803 ({g20, g31, g34, g62, g81}, g82);
	defparam lut_803.LUT_SIZE = 5;
	defparam lut_803.mask = 32'h00000010;

	lut_sub lut_812 ({g21, g8, g24, g77, g37}, g83);
	defparam lut_812.LUT_SIZE = 5;
	defparam lut_812.mask = 32'h50730033;

	lut_sub lut_828 ({g1, g38}, g84);
	defparam lut_828.LUT_SIZE = 2;
	defparam lut_828.mask = 4'b1000;

	lut_sub lut_832 ({i_4_, i_5_, i_6_}, g85);
	defparam lut_832.LUT_SIZE = 3;
	defparam lut_832.mask = 8'h40;

	lut_sub lut_836 ({i_3_, i_0_, i_2_}, g86);
	defparam lut_836.LUT_SIZE = 3;
	defparam lut_836.mask = 8'h01;

	lut_sub lut_845 ({g63, g8, g84, g85, g86}, g87);
	defparam lut_845.LUT_SIZE = 5;
	defparam lut_845.mask = 32'h000f111f;

	lut_sub lut_861 ({g42, g36}, g88);
	defparam lut_861.LUT_SIZE = 2;
	defparam lut_861.mask = 4'b0010;

	lut_sub lut_869 ({g23, g3, g29, g88}, g89);
	defparam lut_869.LUT_SIZE = 4;
	defparam lut_869.mask = 16'h5703;

	lut_sub lut_883 ({g45, g6, g13, g89}, g90);
	defparam lut_883.LUT_SIZE = 4;
	defparam lut_883.mask = 16'ha2aa;

	lut_sub lut_895 ({g36, g13}, g91);
	defparam lut_895.LUT_SIZE = 2;
	defparam lut_895.mask = 4'b1000;

	lut_sub lut_902 ({g42, g12, g3}, g92);
	defparam lut_902.LUT_SIZE = 3;
	defparam lut_902.mask = 8'h01;

	lut_sub lut_911 ({g41, g45, g48, g91, g92}, g93);
	defparam lut_911.LUT_SIZE = 5;
	defparam lut_911.mask = 32'ha8a800a8;

	lut_sub lut_923 ({i_3_, i_0_, i_1_}, g94);
	defparam lut_923.LUT_SIZE = 3;
	defparam lut_923.mask = 8'h20;

	lut_sub lut_929 ({g47, g94}, g95);
	defparam lut_929.LUT_SIZE = 2;
	defparam lut_929.mask = 4'b0001;

	lut_sub lut_935 ({g85, g95}, g96);
	defparam lut_935.LUT_SIZE = 2;
	defparam lut_935.mask = 4'b0001;

	lut_sub lut_942 ({g27, g23, g32}, g97);
	defparam lut_942.LUT_SIZE = 3;
	defparam lut_942.mask = 8'h40;

	lut_sub lut_948 ({g24, g36}, g98);
	defparam lut_948.LUT_SIZE = 2;
	defparam lut_948.mask = 4'b1000;

	lut_sub lut_954 ({g25, g3}, g99);
	defparam lut_954.LUT_SIZE = 2;
	defparam lut_954.mask = 4'b0100;

	lut_sub lut_960 ({g3, g13}, g100);
	defparam lut_960.LUT_SIZE = 2;
	defparam lut_960.mask = 4'b0010;

	lut_sub lut_967 ({i_6_, i_7_, i_8_, g98, g99, g100}, g101);
	defparam lut_967.LUT_SIZE = 6;
	defparam lut_967.mask = 64'h00330f0f55550000;

	lut_sub lut_994 ({g8, g12, g75, g49}, g102);
	defparam lut_994.LUT_SIZE = 4;
	defparam lut_994.mask = 16'h0537;

	lut_sub lut_1008 ({g28, g42, g45, g24}, g103);
	defparam lut_1008.LUT_SIZE = 4;
	defparam lut_1008.mask = 16'h008c;

	lut_sub lut_1018 ({g21, g25, g12, g103}, g104);
	defparam lut_1018.LUT_SIZE = 4;
	defparam lut_1018.mask = 16'h8aaa;

	lut_sub lut_1030 ({g24, g38}, g105);
	defparam lut_1030.LUT_SIZE = 2;
	defparam lut_1030.mask = 4'b0111;

	lut_sub lut_1040 ({g21, g25, g48, g105}, g106);
	defparam lut_1040.LUT_SIZE = 4;
	defparam lut_1040.mask = 16'h3222;

	lut_sub lut_1053 ({g35, g98, g102, g104, g106}, g107);
	defparam lut_1053.LUT_SIZE = 5;
	defparam lut_1053.mask = 32'h20202000;

	lut_sub lut_1063 ({g96, g97, g101, g107}, g108);
	defparam lut_1063.LUT_SIZE = 4;
	defparam lut_1063.mask = 16'h4000;

	lut_sub lut_1072 ({g83, g87, g90, g93, g108}, g109);
	defparam lut_1072.LUT_SIZE = 5;
	defparam lut_1072.mask = 32'h01000000;

	lut_sub lut_1076 ({i_0_, i_1_, i_2_}, g110);
	defparam lut_1076.LUT_SIZE = 3;
	defparam lut_1076.mask = 8'h40;

	lut_sub lut_1080 ({i_6_, i_7_}, g111);
	defparam lut_1080.LUT_SIZE = 2;
	defparam lut_1080.mask = 4'b0100;

	lut_sub lut_1087 ({g36, g110, g111}, g112);
	defparam lut_1087.LUT_SIZE = 3;
	defparam lut_1087.mask = 8'h10;

	lut_sub lut_1093 ({i_7_, i_8_, g21, g36}, g113);
	defparam lut_1093.LUT_SIZE = 4;
	defparam lut_1093.mask = 16'ha0c0;

	lut_sub lut_1105 ({g5, g36, g110, g111, g113}, g114);
	defparam lut_1105.LUT_SIZE = 5;
	defparam lut_1105.mask = 32'ha8aa8888;

	lut_sub lut_1125 ({g47, g13, g15, g26, g112, g114}, g115);
	defparam lut_1125.LUT_SIZE = 6;
	defparam lut_1125.mask = 64'h5555dddd5000d0c0;

	lut_sub lut_1155 ({i_3_, i_5_}, g116);
	defparam lut_1155.LUT_SIZE = 2;
	defparam lut_1155.mask = 4'b0001;

	lut_sub lut_1161 ({g13, g116}, g117);
	defparam lut_1161.LUT_SIZE = 2;
	defparam lut_1161.mask = 4'b0100;

	lut_sub lut_1170 ({g21, g42, g12, g2, g59}, g118);
	defparam lut_1170.LUT_SIZE = 5;
	defparam lut_1170.mask = 32'h002f0022;

	lut_sub lut_1185 ({g28, g48, g26, g117, g118}, g119);
	defparam lut_1185.LUT_SIZE = 5;
	defparam lut_1185.mask = 32'haa88a080;

	lut_sub lut_1197 ({i_3_, i_4_}, g120);
	defparam lut_1197.LUT_SIZE = 2;
	defparam lut_1197.mask = 4'b0001;

	lut_sub lut_1203 ({g28, g13}, g121);
	defparam lut_1203.LUT_SIZE = 2;
	defparam lut_1203.mask = 4'b0010;

	lut_sub lut_1213 ({g42, g45, g6, g24, g3, g111}, g122);
	defparam lut_1213.LUT_SIZE = 6;
	defparam lut_1213.mask = 64'h5050000050730033;

	lut_sub lut_1233 ({g50, g8}, g123);
	defparam lut_1233.LUT_SIZE = 2;
	defparam lut_1233.mask = 4'b0001;

	lut_sub lut_1240 ({g21, g2, g110}, g124);
	defparam lut_1240.LUT_SIZE = 3;
	defparam lut_1240.mask = 8'h10;

	lut_sub lut_1249 ({g12, g123, g105, g86, g124}, g125);
	defparam lut_1249.LUT_SIZE = 5;
	defparam lut_1249.mask = 32'haa880a08;

	lut_sub lut_1261 ({i_3_, i_4_, i_5_, i_0_, i_1_}, g126);
	defparam lut_1261.LUT_SIZE = 5;
	defparam lut_1261.mask = 32'hddffffbf;

	lut_sub lut_1293 ({i_0_, i_1_}, g127);
	defparam lut_1293.LUT_SIZE = 2;
	defparam lut_1293.mask = 4'b0001;

	lut_sub lut_1298 ({i_3_, i_4_, g127}, g128);
	defparam lut_1298.LUT_SIZE = 3;
	defparam lut_1298.mask = 8'h04;

	lut_sub lut_1304 ({g42, g32}, g129);
	defparam lut_1304.LUT_SIZE = 2;
	defparam lut_1304.mask = 4'b0001;

	lut_sub lut_1313 ({g28, g75, g37, g99, g129}, g130);
	defparam lut_1313.LUT_SIZE = 5;
	defparam lut_1313.mask = 32'hfafa8800;

	lut_sub lut_1335 ({g120, g1, g48, g2, g38}, g131);
	defparam lut_1335.LUT_SIZE = 5;
	defparam lut_1335.mask = 32'h22002f00;

	lut_sub lut_1350 ({g12, g683, g128, g130, g131}, g132);
	defparam lut_1350.LUT_SIZE = 5;
	defparam lut_1350.mask = 32'h00220020;

	lut_sub lut_1360 ({g694, g122, g125, g132}, g133);
	defparam lut_1360.LUT_SIZE = 4;
	defparam lut_1360.mask = 16'h0010;

	lut_sub lut_1364 ({i_4_, i_5_, i_6_}, g134);
	defparam lut_1364.LUT_SIZE = 3;
	defparam lut_1364.mask = 8'h80;

	lut_sub lut_1370 ({i_3_, i_2_, g47, g134}, g135);
	defparam lut_1370.LUT_SIZE = 4;
	defparam lut_1370.mask = 16'h0001;

	lut_sub lut_1377 ({i_3_, i_5_, i_2_, g35, g14, g64}, g136);
	defparam lut_1377.LUT_SIZE = 6;
	defparam lut_1377.mask = 64'h0f00000000110011;

	lut_sub lut_1388 ({i_7_, i_8_}, g137);
	defparam lut_1388.LUT_SIZE = 2;
	defparam lut_1388.mask = 4'b0010;

	lut_sub lut_1394 ({i_3_, i_0_, i_1_, g137, g85}, g138);
	defparam lut_1394.LUT_SIZE = 5;
	defparam lut_1394.mask = 32'h01000000;

	lut_sub lut_1400 ({i_3_, i_5_, g28, g24}, g139);
	defparam lut_1400.LUT_SIZE = 4;
	defparam lut_1400.mask = 16'h0200;

	lut_sub lut_1409 ({g27, g6, g36, g138, g139}, g140);
	defparam lut_1409.LUT_SIZE = 5;
	defparam lut_1409.mask = 32'h88088888;

	lut_sub lut_1421 ({g35, g24}, g141);
	defparam lut_1421.LUT_SIZE = 2;
	defparam lut_1421.mask = 4'b0010;

	lut_sub lut_1429 ({i_3_, g42, g8, g45, g141}, g142);
	defparam lut_1429.LUT_SIZE = 5;
	defparam lut_1429.mask = 32'h444f4444;

	lut_sub lut_1446 ({i_8_, g51, g64, g142}, g143);
	defparam lut_1446.LUT_SIZE = 4;
	defparam lut_1446.mask = 16'ha8aa;

	lut_sub lut_1460 ({i_1_, g135, g136, g140, g143}, g144);
	defparam lut_1460.LUT_SIZE = 5;
	defparam lut_1460.mask = 32'h11111000;

	lut_sub lut_1472 ({i_6_, g137, g51, g33, g85}, g145);
	defparam lut_1472.LUT_SIZE = 5;
	defparam lut_1472.mask = 32'h00370005;

	lut_sub lut_1486 ({g27, i_6_, g47, g24, g3}, g146);
	defparam lut_1486.LUT_SIZE = 5;
	defparam lut_1486.mask = 32'h05050004;

	lut_sub lut_1499 ({g37, g38, g110, g145, g146}, g147);
	defparam lut_1499.LUT_SIZE = 5;
	defparam lut_1499.mask = 32'h88888088;

	lut_sub lut_1514 ({g11, g42, g47, g64, g111}, g148);
	defparam lut_1514.LUT_SIZE = 5;
	defparam lut_1514.mask = 32'h00570003;

	lut_sub lut_1528 ({g21, g23, g7, g100}, g149);
	defparam lut_1528.LUT_SIZE = 4;
	defparam lut_1528.mask = 16'h7350;

	lut_sub lut_1541 ({g12, g59, g13}, g150);
	defparam lut_1541.LUT_SIZE = 3;
	defparam lut_1541.mask = 8'h08;

	lut_sub lut_1549 ({g25, g12, g3, g150}, g151);
	defparam lut_1549.LUT_SIZE = 4;
	defparam lut_1549.mask = 16'ha8aa;

	lut_sub lut_1564 ({g6, g77, g148, g149, g151}, g152);
	defparam lut_1564.LUT_SIZE = 5;
	defparam lut_1564.mask = 32'h40404000;

	lut_sub lut_1573 ({g670, g147, g152}, g153);
	defparam lut_1573.LUT_SIZE = 3;
	defparam lut_1573.mask = 8'h01;

	lut_sub lut_1582 ({g115, g119, g133, g144, g153}, g154);
	defparam lut_1582.LUT_SIZE = 5;
	defparam lut_1582.mask = 32'h00000001;

	lut_sub lut_1589 ({g11, g27, g28}, g155);
	defparam lut_1589.LUT_SIZE = 3;
	defparam lut_1589.mask = 8'h40;

	lut_sub lut_1597 ({g23, g36, g7, g129}, g156);
	defparam lut_1597.LUT_SIZE = 4;
	defparam lut_1597.mask = 16'h7530;

	lut_sub lut_1611 ({g47, g75, g155, g156}, g157);
	defparam lut_1611.LUT_SIZE = 4;
	defparam lut_1611.mask = 16'h8880;

	lut_sub lut_1619 ({g1, g59}, g158);
	defparam lut_1619.LUT_SIZE = 2;
	defparam lut_1619.mask = 4'b1000;

	lut_sub lut_1625 ({g21, g48}, g159);
	defparam lut_1625.LUT_SIZE = 2;
	defparam lut_1625.mask = 4'b0100;

	lut_sub lut_1633 ({g42, g12, g84, g159}, g160);
	defparam lut_1633.LUT_SIZE = 4;
	defparam lut_1633.mask = 16'h0357;

	lut_sub lut_1645 ({g11, g110}, g161);
	defparam lut_1645.LUT_SIZE = 2;
	defparam lut_1645.mask = 4'b0100;

	lut_sub lut_1654 ({g28, g2, g24, g32, g161}, g162);
	defparam lut_1654.LUT_SIZE = 5;
	defparam lut_1654.mask = 32'h00305575;

	lut_sub lut_1671 ({i_7_, i_8_, g45, g13, g88}, g163);
	defparam lut_1671.LUT_SIZE = 5;
	defparam lut_1671.mask = 32'h0000c055;

	lut_sub lut_1685 ({g2, g158, g160, g162, g163}, g164);
	defparam lut_1685.LUT_SIZE = 5;
	defparam lut_1685.mask = 32'h80808000;

	lut_sub lut_1694 ({g27, g59, g60}, g165);
	defparam lut_1694.LUT_SIZE = 3;
	defparam lut_1694.mask = 8'h40;

	lut_sub lut_1701 ({i_5_, g42, g2, g165}, g166);
	defparam lut_1701.LUT_SIZE = 4;
	defparam lut_1701.mask = 16'ha8aa;

	lut_sub lut_1713 ({g14, g134}, g167);
	defparam lut_1713.LUT_SIZE = 2;
	defparam lut_1713.mask = 4'b0001;

	lut_sub lut_1720 ({i_0_, i_2_, g35, g75, g167}, g168);
	defparam lut_1720.LUT_SIZE = 5;
	defparam lut_1720.mask = 32'h03030357;

	lut_sub lut_1737 ({g50, i_6_, g42, g47}, g169);
	defparam lut_1737.LUT_SIZE = 4;
	defparam lut_1737.mask = 16'h0001;

	lut_sub lut_1743 ({i_3_, i_5_, g25, g12}, g170);
	defparam lut_1743.LUT_SIZE = 4;
	defparam lut_1743.mask = 16'h0040;

	lut_sub lut_1749 ({i_3_, i_5_, g2, g13}, g171);
	defparam lut_1749.LUT_SIZE = 4;
	defparam lut_1749.mask = 16'h0200;

	lut_sub lut_1757 ({g32, g121, g170, g171}, g172);
	defparam lut_1757.LUT_SIZE = 4;
	defparam lut_1757.mask = 16'h8880;

	lut_sub lut_1767 ({g127, i_2_, g8, g45, g12}, g173);
	defparam lut_1767.LUT_SIZE = 5;
	defparam lut_1767.mask = 32'h00000c44;

	lut_sub lut_1778 ({g11, g8, g29, g91}, g174);
	defparam lut_1778.LUT_SIZE = 4;
	defparam lut_1778.mask = 16'h3705;

	lut_sub lut_1792 ({g25, g45, g22, g6}, g175);
	defparam lut_1792.LUT_SIZE = 4;
	defparam lut_1792.mask = 16'h7300;

	lut_sub lut_1805 ({g28, g25, g59, g7, g110}, g176);
	defparam lut_1805.LUT_SIZE = 5;
	defparam lut_1805.mask = 32'h3030f070;

	lut_sub lut_1823 ({g173, g174, g175, g176}, g177);
	defparam lut_1823.LUT_SIZE = 4;
	defparam lut_1823.mask = 16'h8000;

	lut_sub lut_1832 ({g11, g9, g169, g172, g177}, g178);
	defparam lut_1832.LUT_SIZE = 5;
	defparam lut_1832.mask = 32'h10001010;

	lut_sub lut_1843 ({g35, g21, g12, g24, g26}, g179);
	defparam lut_1843.LUT_SIZE = 5;
	defparam lut_1843.mask = 32'h0c005d55;

	lut_sub lut_1860 ({i_3_, i_4_, i_5_, g127, g63, g51}, g180);
	defparam lut_1860.LUT_SIZE = 6;
	defparam lut_1860.mask = 64'h0011000000110003;

	lut_sub lut_1871 ({g45, g110}, g181);
	defparam lut_1871.LUT_SIZE = 2;
	defparam lut_1871.mask = 4'b0100;

	lut_sub lut_1878 ({i_6_, i_7_, i_8_, g75, g181, g105}, g182);
	defparam lut_1878.LUT_SIZE = 6;
	defparam lut_1878.mask = 64'h00000f00aa000033;

	lut_sub lut_1896 ({i_3_, i_5_, g127, g28, g123}, g183);
	defparam lut_1896.LUT_SIZE = 5;
	defparam lut_1896.mask = 32'h05050003;

	lut_sub lut_1907 ({g59, g110}, g184);
	defparam lut_1907.LUT_SIZE = 2;
	defparam lut_1907.mask = 4'b0100;

	lut_sub lut_1915 ({g2, g23, g70, g184}, g185);
	defparam lut_1915.LUT_SIZE = 4;
	defparam lut_1915.mask = 16'h5073;

	lut_sub lut_1930 ({g45, g48, g2, g24, g184}, g186);
	defparam lut_1930.LUT_SIZE = 5;
	defparam lut_1930.mask = 32'h05cd0505;

	lut_sub lut_1944 ({i_3_, i_4_, i_5_, i_6_, i_7_, i_8_}, g187);
	defparam lut_1944.LUT_SIZE = 6;
	defparam lut_1944.mask = 64'hff7fff7fbf7faf7f;

	lut_sub lut_2006 ({i_3_, i_5_, g35, g42}, g188);
	defparam lut_2006.LUT_SIZE = 4;
	defparam lut_2006.mask = 16'h0010;

	lut_sub lut_2012 ({g3, g110}, g189);
	defparam lut_2012.LUT_SIZE = 2;
	defparam lut_2012.mask = 4'b0001;

	lut_sub lut_2020 ({i_6_, g63, g188, g181, g189}, g190);
	defparam lut_2020.LUT_SIZE = 5;
	defparam lut_2020.mask = 32'hf0a0f0c0;

	lut_sub lut_2039 ({g185, g186, g657, g190}, g191);
	defparam lut_2039.LUT_SIZE = 4;
	defparam lut_2039.mask = 16'h1000;

	lut_sub lut_2048 ({g179, g180, g182, g183, g191}, g192);
	defparam lut_2048.LUT_SIZE = 5;
	defparam lut_2048.mask = 32'h40000000;

	lut_sub lut_2056 ({g23, g3, g7, g181}, g193);
	defparam lut_2056.LUT_SIZE = 4;
	defparam lut_2056.mask = 16'h5703;

	lut_sub lut_2068 ({g21, g6}, g194);
	defparam lut_2068.LUT_SIZE = 2;
	defparam lut_2068.mask = 4'b0100;

	lut_sub lut_2076 ({g8, g13, g181, g194}, g195);
	defparam lut_2076.LUT_SIZE = 4;
	defparam lut_2076.mask = 16'h5073;

	lut_sub lut_2091 ({g27, g23, g3, g110, g194}, g196);
	defparam lut_2091.LUT_SIZE = 5;
	defparam lut_2091.mask = 32'h1f111111;

	lut_sub lut_2110 ({g47, g73, g193, g195, g196}, g197);
	defparam lut_2110.LUT_SIZE = 5;
	defparam lut_2110.mask = 32'h80808000;

	lut_sub lut_2121 ({g166, g168, g178, g192, g197}, g198);
	defparam lut_2121.LUT_SIZE = 5;
	defparam lut_2121.mask = 32'h00000100;

	lut_sub lut_2130 ({g109, g154, g157, g164, g198}, g199);
	defparam lut_2130.LUT_SIZE = 5;
	defparam lut_2130.mask = 32'h00000001;

	lut_sub lut_2139 ({g27, g45, g23, g36, g121}, g200);
	defparam lut_2139.LUT_SIZE = 5;
	defparam lut_2139.mask = 32'hf4444444;

	lut_sub lut_2157 ({g50, i_6_, g137, g94, g88}, g201);
	defparam lut_2157.LUT_SIZE = 5;
	defparam lut_2157.mask = 32'h05000503;

	lut_sub lut_2170 ({g45, g37, g13, g201}, g202);
	defparam lut_2170.LUT_SIZE = 4;
	defparam lut_2170.mask = 16'ha2aa;

	lut_sub lut_2184 ({i_6_, g63, g21, g13, g84}, g203);
	defparam lut_2184.LUT_SIZE = 5;
	defparam lut_2184.mask = 32'h00c00055;

	lut_sub lut_2196 ({i_6_, i_8_, g32, g105, g141}, g204);
	defparam lut_2196.LUT_SIZE = 5;
	defparam lut_2196.mask = 32'h050505cd;

	lut_sub lut_2213 ({g23, g70, g204}, g205);
	defparam lut_2213.LUT_SIZE = 3;
	defparam lut_2213.mask = 8'h8a;

	lut_sub lut_2224 ({g150, g200, g202, g203, g205}, g206);
	defparam lut_2224.LUT_SIZE = 5;
	defparam lut_2224.mask = 32'h04000000;

	lut_sub lut_2230 ({i_3_, i_5_, g8, g24}, g207);
	defparam lut_2230.LUT_SIZE = 4;
	defparam lut_2230.mask = 16'h2000;

	lut_sub lut_2238 ({i_6_, g42, g46, g47, g38}, g208);
	defparam lut_2238.LUT_SIZE = 5;
	defparam lut_2238.mask = 32'h03030022;

	lut_sub lut_2251 ({g127, i_2_, g8, g22, g59}, g209);
	defparam lut_2251.LUT_SIZE = 5;
	defparam lut_2251.mask = 32'h0000330a;

	lut_sub lut_2265 ({g28, g26, g208, g644, g209}, g210);
	defparam lut_2265.LUT_SIZE = 5;
	defparam lut_2265.mask = 32'h20202000;

	lut_sub lut_2276 ({g1, g47, g64, g207, g210}, g211);
	defparam lut_2276.LUT_SIZE = 5;
	defparam lut_2276.mask = 32'h44404444;

	lut_sub lut_2289 ({g45, g23, g24}, g212);
	defparam lut_2289.LUT_SIZE = 3;
	defparam lut_2289.mask = 8'h80;

	lut_sub lut_2296 ({g50, i_6_, g42, g137}, g213);
	defparam lut_2296.LUT_SIZE = 4;
	defparam lut_2296.mask = 16'h0001;

	lut_sub lut_2305 ({g2, g73, g38, g29, g213}, g214);
	defparam lut_2305.LUT_SIZE = 5;
	defparam lut_2305.mask = 32'h8a8a8a00;

	lut_sub lut_2320 ({i_4_, i_5_, g6, g13, g214}, g215);
	defparam lut_2320.LUT_SIZE = 5;
	defparam lut_2320.mask = 32'h55555551;

	lut_sub lut_2341 ({i_1_, g135, g212, g215}, g216);
	defparam lut_2341.LUT_SIZE = 4;
	defparam lut_2341.mask = 16'h4044;

	lut_sub lut_2347 ({i_3_, i_5_, i_6_}, g217);
	defparam lut_2347.LUT_SIZE = 3;
	defparam lut_2347.mask = 8'h20;

	lut_sub lut_2353 ({g42, g217}, g218);
	defparam lut_2353.LUT_SIZE = 2;
	defparam lut_2353.mask = 4'b0001;

	lut_sub lut_2359 ({g63, g15}, g219);
	defparam lut_2359.LUT_SIZE = 2;
	defparam lut_2359.mask = 4'b0001;

	lut_sub lut_2364 ({i_3_, i_1_, i_2_, g219}, g220);
	defparam lut_2364.LUT_SIZE = 4;
	defparam lut_2364.mask = 16'h0400;

	lut_sub lut_2373 ({g27, g35, g28, g1, g36}, g221);
	defparam lut_2373.LUT_SIZE = 5;
	defparam lut_2373.mask = 32'h0a8a0088;

	lut_sub lut_2388 ({g23, g59, g13, g105, g221}, g222);
	defparam lut_2388.LUT_SIZE = 5;
	defparam lut_2388.mask = 32'h0222aaaa;

	lut_sub lut_2406 ({g27, g43, g23, g3}, g223);
	defparam lut_2406.LUT_SIZE = 4;
	defparam lut_2406.mask = 16'hb0f0;

	lut_sub lut_2420 ({i_7_, g218, g220, g222, g223}, g224);
	defparam lut_2420.LUT_SIZE = 5;
	defparam lut_2420.mask = 32'h10001010;

	lut_sub lut_2426 ({i_3_, i_4_, i_6_}, g225);
	defparam lut_2426.LUT_SIZE = 3;
	defparam lut_2426.mask = 8'h80;

	lut_sub lut_2435 ({g63, g41, g1, g36, g225}, g226);
	defparam lut_2435.LUT_SIZE = 5;
	defparam lut_2435.mask = 32'h00cc50dc;

	lut_sub lut_2451 ({i_6_, i_7_, i_8_, g100, g129}, g227);
	defparam lut_2451.LUT_SIZE = 5;
	defparam lut_2451.mask = 32'h03400000;

	lut_sub lut_2460 ({g186, g226, g227}, g228);
	defparam lut_2460.LUT_SIZE = 3;
	defparam lut_2460.mask = 8'h80;

	lut_sub lut_2467 ({g23, g71, g161}, g229);
	defparam lut_2467.LUT_SIZE = 3;
	defparam lut_2467.mask = 8'h70;

	lut_sub lut_2473 ({i_3_, i_1_, i_2_}, g230);
	defparam lut_2473.LUT_SIZE = 3;
	defparam lut_2473.mask = 8'h10;

	lut_sub lut_2482 ({g50, g8, g12, g57, g230}, g231);
	defparam lut_2482.LUT_SIZE = 5;
	defparam lut_2482.mask = 32'h00000537;

	lut_sub lut_2495 ({i_6_, i_7_, i_8_, g75, g158, g231}, g232);
	defparam lut_2495.LUT_SIZE = 6;
	defparam lut_2495.mask = 64'h88aaa0aaa0aaaaa0;

	lut_sub lut_2527 ({g25, g194, g229, g631, g232}, g233);
	defparam lut_2527.LUT_SIZE = 5;
	defparam lut_2527.mask = 32'h10001010;

	lut_sub lut_2538 ({g30, g216, g224, g228, g233}, g234);
	defparam lut_2538.LUT_SIZE = 5;
	defparam lut_2538.mask = 32'h00010000;

	lut_sub lut_2547 ({g35, g21, g8, g25, g32}, g235);
	defparam lut_2547.LUT_SIZE = 5;
	defparam lut_2547.mask = 32'h0404cc04;

	lut_sub lut_2562 ({g6, g73, g49, g60, g235}, g236);
	defparam lut_2562.LUT_SIZE = 5;
	defparam lut_2562.mask = 32'ha8a8a800;

	lut_sub lut_2578 ({g21, g8, g24, g69}, g237);
	defparam lut_2578.LUT_SIZE = 4;
	defparam lut_2578.mask = 16'h5155;

	lut_sub lut_2593 ({g11, g1, g23, g3, g141}, g238);
	defparam lut_2593.LUT_SIZE = 5;
	defparam lut_2593.mask = 32'h75553000;

	lut_sub lut_2612 ({g11, g45, g2, g23, g13}, g239);
	defparam lut_2612.LUT_SIZE = 5;
	defparam lut_2612.mask = 32'h8a880a00;

	lut_sub lut_2626 ({g25, g120, g12, g181}, g240);
	defparam lut_2626.LUT_SIZE = 4;
	defparam lut_2626.mask = 16'h1311;

	lut_sub lut_2638 ({g59, g29, g239, g240}, g241);
	defparam lut_2638.LUT_SIZE = 4;
	defparam lut_2638.mask = 16'h8088;

	lut_sub lut_2648 ({g6, g88, g238, g241}, g242);
	defparam lut_2648.LUT_SIZE = 4;
	defparam lut_2648.mask = 16'h4440;

	lut_sub lut_2656 ({g25, g36}, g243);
	defparam lut_2656.LUT_SIZE = 2;
	defparam lut_2656.mask = 4'b1000;

	lut_sub lut_2663 ({g63, g51, g134}, g244);
	defparam lut_2663.LUT_SIZE = 3;
	defparam lut_2663.mask = 8'h01;

	lut_sub lut_2671 ({g2, g24, g32, g244}, g245);
	defparam lut_2671.LUT_SIZE = 4;
	defparam lut_2671.mask = 16'haa8a;

	lut_sub lut_2683 ({i_6_, i_8_, g243, g245}, g246);
	defparam lut_2683.LUT_SIZE = 4;
	defparam lut_2683.mask = 16'h5455;

	lut_sub lut_2698 ({g35, g42, g25, g23, g3}, g247);
	defparam lut_2698.LUT_SIZE = 5;
	defparam lut_2698.mask = 32'h40404055;

	lut_sub lut_2712 ({g45, g38, g29, g121}, g248);
	defparam lut_2712.LUT_SIZE = 4;
	defparam lut_2712.mask = 16'h7350;

	lut_sub lut_2727 ({g21, g8, g25, g247, g248}, g249);
	defparam lut_2727.LUT_SIZE = 5;
	defparam lut_2727.mask = 32'h88088888;

	lut_sub lut_2738 ({i_3_, i_4_, g27, i_6_, i_8_}, g250);
	defparam lut_2738.LUT_SIZE = 5;
	defparam lut_2738.mask = 32'h00002000;

	lut_sub lut_2744 ({i_3_, i_0_, i_1_, g219, g250}, g251);
	defparam lut_2744.LUT_SIZE = 5;
	defparam lut_2744.mask = 32'ha8aaaaaa;

	lut_sub lut_2765 ({g27, g28, g45}, g252);
	defparam lut_2765.LUT_SIZE = 3;
	defparam lut_2765.mask = 8'h20;

	lut_sub lut_2774 ({g48, g57, g33, g16, g252}, g253);
	defparam lut_2774.LUT_SIZE = 5;
	defparam lut_2774.mask = 32'haa88a080;

	lut_sub lut_2791 ({g127, g6, g5, g251, g253}, g254);
	defparam lut_2791.LUT_SIZE = 5;
	defparam lut_2791.mask = 32'h11111110;

	lut_sub lut_2806 ({g14, g1, g12, g3, g225}, g255);
	defparam lut_2806.LUT_SIZE = 5;
	defparam lut_2806.mask = 32'h03005700;

	lut_sub lut_2819 ({g25, g120, g23}, g256);
	defparam lut_2819.LUT_SIZE = 3;
	defparam lut_2819.mask = 8'h20;

	lut_sub lut_2828 ({g8, g1, g22, g105, g256}, g257);
	defparam lut_2828.LUT_SIZE = 5;
	defparam lut_2828.mask = 32'ha0aa2022;

	lut_sub lut_2845 ({g28, g70, g189, g167, g230}, g258);
	defparam lut_2845.LUT_SIZE = 5;
	defparam lut_2845.mask = 32'heeeee000;

	lut_sub lut_2867 ({g45, g6, g110, g141}, g259);
	defparam lut_2867.LUT_SIZE = 4;
	defparam lut_2867.mask = 16'h5700;

	lut_sub lut_2880 ({g24, g36, g60, g4, g259}, g260);
	defparam lut_2880.LUT_SIZE = 5;
	defparam lut_2880.mask = 32'h8088aaaa;

	lut_sub lut_2899 ({g83, g255, g257, g258, g260}, g261);
	defparam lut_2899.LUT_SIZE = 5;
	defparam lut_2899.mask = 32'h01000000;

	lut_sub lut_2909 ({g237, g242, g246, g249, g254, g261}, g262);
	defparam lut_2909.LUT_SIZE = 6;
	defparam lut_2909.mask = 64'h0000000000000001;

	lut_sub lut_2919 ({g157, g206, g211, g234, g236, g262}, g263);
	defparam lut_2919.LUT_SIZE = 6;
	defparam lut_2919.mask = 64'h0000000000000001;

	lut_sub lut_2929 ({g11, g42, g23, g13, g60, g38}, g264);
	defparam lut_2929.LUT_SIZE = 6;
	defparam lut_2929.mask = 64'ha000b333a000a000;

	lut_sub lut_2949 ({g27, i_6_, g47}, g265);
	defparam lut_2949.LUT_SIZE = 3;
	defparam lut_2949.mask = 8'h40;

	lut_sub lut_2957 ({g11, g12, g71, g265}, g266);
	defparam lut_2957.LUT_SIZE = 4;
	defparam lut_2957.mask = 16'h5703;

	lut_sub lut_2972 ({g27, g35, g36, g110, g194}, g267);
	defparam lut_2972.LUT_SIZE = 5;
	defparam lut_2972.mask = 32'h55750030;

	lut_sub lut_2988 ({g24, g225}, g268);
	defparam lut_2988.LUT_SIZE = 2;
	defparam lut_2988.mask = 4'b0100;

	lut_sub lut_2995 ({i_7_, g28, g75, g268}, g269);
	defparam lut_2995.LUT_SIZE = 4;
	defparam lut_2995.mask = 16'h0357;

	lut_sub lut_3009 ({g1, g6, g36, g49}, g270);
	defparam lut_3009.LUT_SIZE = 4;
	defparam lut_3009.mask = 16'h0d05;

	lut_sub lut_3023 ({g27, g45, g1, g23, g4, g189}, g271);
	defparam lut_3023.LUT_SIZE = 6;
	defparam lut_3023.mask = 64'hf3737373f0505050;

	lut_sub lut_3061 ({g48, g105, g270, g271}, g272);
	defparam lut_3061.LUT_SIZE = 4;
	defparam lut_3061.mask = 16'h8808;

	lut_sub lut_3072 ({g8, g77, g200, g269, g272}, g273);
	defparam lut_3072.LUT_SIZE = 5;
	defparam lut_3072.mask = 32'h40404000;

	lut_sub lut_3083 ({g264, g266, g267, g215, g273}, g274);
	defparam lut_3083.LUT_SIZE = 5;
	defparam lut_3083.mask = 32'h10000000;

	lut_sub lut_3090 ({g27, i_7_, i_8_, g36, g100}, g275);
	defparam lut_3090.LUT_SIZE = 5;
	defparam lut_3090.mask = 32'h00c50005;

	lut_sub lut_3104 ({g28, g42, g23, g3, g91}, g276);
	defparam lut_3104.LUT_SIZE = 5;
	defparam lut_3104.mask = 32'h50505073;

	lut_sub lut_3123 ({g11, g8, g12, g13, g184}, g277);
	defparam lut_3123.LUT_SIZE = 5;
	defparam lut_3123.mask = 32'h0c5d0055;

	lut_sub lut_3140 ({g35, g46, g158}, g278);
	defparam lut_3140.LUT_SIZE = 3;
	defparam lut_3140.mask = 8'h07;

	lut_sub lut_3150 ({g38, g94, g265, g167}, g279);
	defparam lut_3150.LUT_SIZE = 4;
	defparam lut_3150.mask = 16'h3705;

	lut_sub lut_3165 ({g25, g6, g32, g121, g252}, g280);
	defparam lut_3165.LUT_SIZE = 5;
	defparam lut_3165.mask = 32'ha8a0a8a8;

	lut_sub lut_3183 ({g35, g6, g117, g161}, g281);
	defparam lut_3183.LUT_SIZE = 4;
	defparam lut_3183.mask = 16'h0537;

	lut_sub lut_3198 ({g277, g278, g279, g280, g281}, g282);
	defparam lut_3198.LUT_SIZE = 5;
	defparam lut_3198.mask = 32'h20000000;

	lut_sub lut_3206 ({i_0_, g135, g275, g276, g282}, g283);
	defparam lut_3206.LUT_SIZE = 5;
	defparam lut_3206.mask = 32'h40404000;

	lut_sub lut_3215 ({g27, g137, g15}, g284);
	defparam lut_3215.LUT_SIZE = 3;
	defparam lut_3215.mask = 8'h10;

	lut_sub lut_3221 ({i_6_, i_8_, g1, g32}, g285);
	defparam lut_3221.LUT_SIZE = 4;
	defparam lut_3221.mask = 16'h4000;

	lut_sub lut_3228 ({g2, g26, g155}, g286);
	defparam lut_3228.LUT_SIZE = 3;
	defparam lut_3228.mask = 8'ha8;

	lut_sub lut_3239 ({g25, g194, g212, g285, g286}, g287);
	defparam lut_3239.LUT_SIZE = 5;
	defparam lut_3239.mask = 32'h40004040;

	lut_sub lut_3249 ({g28, g12, g184, g243}, g288);
	defparam lut_3249.LUT_SIZE = 4;
	defparam lut_3249.mask = 16'h0357;

	lut_sub lut_3264 ({g13, g123, g284, g287, g288}, g289);
	defparam lut_3264.LUT_SIZE = 5;
	defparam lut_3264.mask = 32'h20002020;

	lut_sub lut_3273 ({g42, g2, g38}, g290);
	defparam lut_3273.LUT_SIZE = 3;
	defparam lut_3273.mask = 8'h02;

	lut_sub lut_3281 ({g48, g181, g244, g290}, g291);
	defparam lut_3281.LUT_SIZE = 4;
	defparam lut_3281.mask = 16'h8880;

	lut_sub lut_3289 ({g27, i_6_, i_8_, g21}, g292);
	defparam lut_3289.LUT_SIZE = 4;
	defparam lut_3289.mask = 16'h0800;

	lut_sub lut_3298 ({g27, g35, g45, g6, g84}, g293);
	defparam lut_3298.LUT_SIZE = 5;
	defparam lut_3298.mask = 32'h30750055;

	lut_sub lut_3315 ({g28, g45, g24}, g294);
	defparam lut_3315.LUT_SIZE = 3;
	defparam lut_3315.mask = 8'h08;

	lut_sub lut_3324 ({i_5_, g35, g42, g5, g121, g294}, g295);
	defparam lut_3324.LUT_SIZE = 6;
	defparam lut_3324.mask = 64'haaaaaaa0a8a8a8a8;

	lut_sub lut_3355 ({g8, g243}, g296);
	defparam lut_3355.LUT_SIZE = 2;
	defparam lut_3355.mask = 4'b0001;

	lut_sub lut_3362 ({i_3_, i_5_, g35, g14, g85}, g297);
	defparam lut_3362.LUT_SIZE = 5;
	defparam lut_3362.mask = 32'h1f111111;

	lut_sub lut_3381 ({g23, g24, g70, g296, g297}, g298);
	defparam lut_3381.LUT_SIZE = 5;
	defparam lut_3381.mask = 32'h80c088cc;

	lut_sub lut_3397 ({g292, g293, g295, g298}, g299);
	defparam lut_3397.LUT_SIZE = 4;
	defparam lut_3397.mask = 16'h1000;

	lut_sub lut_3406 ({g164, g283, g289, g291, g299}, g300);
	defparam lut_3406.LUT_SIZE = 5;
	defparam lut_3406.mask = 32'h00000001;

	lut_sub lut_3414 ({i_6_, g137, g77, g13, g64}, g301);
	defparam lut_3414.LUT_SIZE = 5;
	defparam lut_3414.mask = 32'h004f0044;

	lut_sub lut_3428 ({i_6_, g21, g1, g137, g59}, g302);
	defparam lut_3428.LUT_SIZE = 5;
	defparam lut_3428.mask = 32'h20203020;

	lut_sub lut_3440 ({g27, g63, g38, g96}, g303);
	defparam lut_3440.LUT_SIZE = 4;
	defparam lut_3440.mask = 16'ha2aa;

	lut_sub lut_3455 ({g35, g45, g13, g4, g243}, g304);
	defparam lut_3455.LUT_SIZE = 5;
	defparam lut_3455.mask = 32'h3030f575;

	lut_sub lut_3477 ({g2, g6, g75, g71}, g305);
	defparam lut_3477.LUT_SIZE = 4;
	defparam lut_3477.mask = 16'h0537;

	lut_sub lut_3492 ({g23, g184, g304, g607, g305}, g306);
	defparam lut_3492.LUT_SIZE = 5;
	defparam lut_3492.mask = 32'h20002020;

	lut_sub lut_3503 ({g11, g67, g302, g303, g306}, g307);
	defparam lut_3503.LUT_SIZE = 5;
	defparam lut_3503.mask = 32'h10001010;

	lut_sub lut_3511 ({i_3_, i_4_, i_0_, i_2_, g12, g219}, g308);
	defparam lut_3511.LUT_SIZE = 6;
	defparam lut_3511.mask = 64'h0505050503000000;

	lut_sub lut_3528 ({g42, g23, g194, g98}, g309);
	defparam lut_3528.LUT_SIZE = 4;
	defparam lut_3528.mask = 16'h5073;

	lut_sub lut_3540 ({i_6_, i_7_, g129, g309}, g310);
	defparam lut_3540.LUT_SIZE = 4;
	defparam lut_3540.mask = 16'haa8a;

	lut_sub lut_3555 ({g2, g23, g59, g13, g84}, g311);
	defparam lut_3555.LUT_SIZE = 5;
	defparam lut_3555.mask = 32'h5500d5c0;

	lut_sub lut_3572 ({i_3_, i_4_, g28, g24, g311}, g312);
	defparam lut_3572.LUT_SIZE = 5;
	defparam lut_3572.mask = 32'haaaaa2aa;

	lut_sub lut_3595 ({g25, g12, g32, g9, g116}, g313);
	defparam lut_3595.LUT_SIZE = 5;
	defparam lut_3595.mask = 32'h111f1111;

	lut_sub lut_3614 ({g11, g48, g24, g32, g9}, g314);
	defparam lut_3614.LUT_SIZE = 5;
	defparam lut_3614.mask = 32'h55750030;

	lut_sub lut_3631 ({g1, g32, g37}, g315);
	defparam lut_3631.LUT_SIZE = 3;
	defparam lut_3631.mask = 8'h10;

	lut_sub lut_3638 ({g6, g105, g315}, g316);
	defparam lut_3638.LUT_SIZE = 3;
	defparam lut_3638.mask = 8'ha2;

	lut_sub lut_3649 ({g48, g313, g314, g52, g316}, g317);
	defparam lut_3649.LUT_SIZE = 5;
	defparam lut_3649.mask = 32'h50004000;

	lut_sub lut_3659 ({g168, g310, g312, g317}, g318);
	defparam lut_3659.LUT_SIZE = 4;
	defparam lut_3659.mask = 16'h0100;

	lut_sub lut_3668 ({g301, g211, g307, g308, g318}, g319);
	defparam lut_3668.LUT_SIZE = 5;
	defparam lut_3668.mask = 32'h00040000;

	lut_sub lut_3678 ({g90, g224, g274, g618, g300, g319}, g320);
	defparam lut_3678.LUT_SIZE = 6;
	defparam lut_3678.mask = 64'h0000000000000001;

	lut_sub lut_3685 ({i_6_, i_7_, i_8_, g26, g243, g268}, g321);
	defparam lut_3685.LUT_SIZE = 6;
	defparam lut_3685.mask = 64'h000033550f003355;

	lut_sub lut_3713 ({g27, g45, g1, g6, g16}, g322);
	defparam lut_3713.LUT_SIZE = 5;
	defparam lut_3713.mask = 32'h73505050;

	lut_sub lut_3732 ({g264, g279, g596, g321, g322}, g323);
	defparam lut_3732.LUT_SIZE = 5;
	defparam lut_3732.mask = 32'h08000000;

	lut_sub lut_3740 ({g28, g48, g189, g184}, g324);
	defparam lut_3740.LUT_SIZE = 4;
	defparam lut_3740.mask = 16'h0537;

	lut_sub lut_3753 ({g137, g134, g230}, g325);
	defparam lut_3753.LUT_SIZE = 3;
	defparam lut_3753.mask = 8'h01;

	lut_sub lut_3762 ({g35, g25, g59, g4, g325}, g326);
	defparam lut_3762.LUT_SIZE = 5;
	defparam lut_3762.mask = 32'h88aa08aa;

	lut_sub lut_3781 ({g35, g181, g276, g324, g326}, g327);
	defparam lut_3781.LUT_SIZE = 5;
	defparam lut_3781.mask = 32'h40404000;

	lut_sub lut_3790 ({i_6_, g14, g26, g99}, g328);
	defparam lut_3790.LUT_SIZE = 4;
	defparam lut_3790.mask = 16'h0305;

	lut_sub lut_3802 ({g45, g6, g24, g67, g91}, g329);
	defparam lut_3802.LUT_SIZE = 5;
	defparam lut_3802.mask = 32'h33f70055;

	lut_sub lut_3825 ({g32, g29, g193, g328, g329}, g330);
	defparam lut_3825.LUT_SIZE = 5;
	defparam lut_3825.mask = 32'h80808000;

	lut_sub lut_3834 ({g14, g64, g230}, g331);
	defparam lut_3834.LUT_SIZE = 3;
	defparam lut_3834.mask = 8'h01;

	lut_sub lut_3843 ({g45, g2, g49, g7, g331}, g332);
	defparam lut_3843.LUT_SIZE = 5;
	defparam lut_3843.mask = 32'h8880aaa0;

	lut_sub lut_3855 ({i_3_, i_4_, i_5_, i_6_, i_7_, i_8_}, g333);
	defparam lut_3855.LUT_SIZE = 6;
	defparam lut_3855.mask = 64'h0000000010000080;

	lut_sub lut_3862 ({i_3_, g27, i_6_, g333}, g334);
	defparam lut_3862.LUT_SIZE = 4;
	defparam lut_3862.mask = 16'h0040;

	lut_sub lut_3872 ({g11, g35, g28, g25, g38, g334}, g335);
	defparam lut_3872.LUT_SIZE = 6;
	defparam lut_3872.mask = 64'haa2a0a0aaa2aaa2a;

	lut_sub lut_3904 ({i_3_, g21, g42, g8, g7}, g336);
	defparam lut_3904.LUT_SIZE = 5;
	defparam lut_3904.mask = 32'h55005703;

	lut_sub lut_3920 ({i_6_, i_7_, i_8_, g70, g184}, g337);
	defparam lut_3920.LUT_SIZE = 5;
	defparam lut_3920.mask = 32'h00503050;

	lut_sub lut_3932 ({g46, g48, g60}, g338);
	defparam lut_3932.LUT_SIZE = 3;
	defparam lut_3932.mask = 8'h07;

	lut_sub lut_3943 ({g2, g98, g252, g337, g338}, g339);
	defparam lut_3943.LUT_SIZE = 5;
	defparam lut_3943.mask = 32'h80808000;

	lut_sub lut_3954 ({g312, g332, g335, g336, g339}, g340);
	defparam lut_3954.LUT_SIZE = 5;
	defparam lut_3954.mask = 32'h00000004;

	lut_sub lut_3963 ({g119, g206, g327, g330, g340}, g341);
	defparam lut_3963.LUT_SIZE = 5;
	defparam lut_3963.mask = 32'h00000001;

	lut_sub lut_3971 ({i_0_, g27, g14, g135, g217}, g342);
	defparam lut_3971.LUT_SIZE = 5;
	defparam lut_3971.mask = 32'h05003733;

	lut_sub lut_3989 ({g27, g23, g36, g285}, g343);
	defparam lut_3989.LUT_SIZE = 4;
	defparam lut_3989.mask = 16'h2aaa;

	lut_sub lut_4004 ({g21, g6, g23, g24, g129}, g344);
	defparam lut_4004.LUT_SIZE = 5;
	defparam lut_4004.mask = 32'hc0d50055;

	lut_sub lut_4019 ({i_5_, i_6_, i_7_, i_8_, g5}, g345);
	defparam lut_4019.LUT_SIZE = 5;
	defparam lut_4019.mask = 32'h00440400;

	lut_sub lut_4031 ({g28, g42, g38, g110, g159, g345}, g346);
	defparam lut_4031.LUT_SIZE = 6;
	defparam lut_4031.mask = 64'h030357570f035f57;

	lut_sub lut_4068 ({i_6_, i_7_, i_8_, g46, g77, g189}, g347);
	defparam lut_4068.LUT_SIZE = 6;
	defparam lut_4068.mask = 64'h0f0000000f770f00;

	lut_sub lut_4089 ({i_3_, i_4_, i_0_, i_1_}, g348);
	defparam lut_4089.LUT_SIZE = 4;
	defparam lut_4089.mask = 16'h0020;

	lut_sub lut_4097 ({g2, g161, g296, g348}, g349);
	defparam lut_4097.LUT_SIZE = 4;
	defparam lut_4097.mask = 16'hcc80;

	lut_sub lut_4110 ({g343, g344, g346, g347, g349}, g350);
	defparam lut_4110.LUT_SIZE = 5;
	defparam lut_4110.mask = 32'h00004000;

	lut_sub lut_4116 ({i_5_, i_2_, g48, g219}, g351);
	defparam lut_4116.LUT_SIZE = 4;
	defparam lut_4116.mask = 16'h8aaa;

	lut_sub lut_4127 ({i_3_, i_0_, i_1_, g351}, g352);
	defparam lut_4127.LUT_SIZE = 4;
	defparam lut_4127.mask = 16'h2000;

	lut_sub lut_4133 ({g50, i_6_, i_7_, g86}, g353);
	defparam lut_4133.LUT_SIZE = 4;
	defparam lut_4133.mask = 16'h0004;

	lut_sub lut_4142 ({g13, g4, g352, g125, g353}, g354);
	defparam lut_4142.LUT_SIZE = 5;
	defparam lut_4142.mask = 32'h20002020;

	lut_sub lut_4153 ({g301, g20, g342, g350, g354}, g355);
	defparam lut_4153.LUT_SIZE = 5;
	defparam lut_4153.mask = 32'h00100000;

	lut_sub lut_4162 ({g178, g234, g323, g341, g355}, g356);
	defparam lut_4162.LUT_SIZE = 5;
	defparam lut_4162.mask = 32'h00000001;

	lut_sub lut_4170 ({g6, g4, g110, g243}, g357);
	defparam lut_4170.LUT_SIZE = 4;
	defparam lut_4170.mask = 16'h0357;

	lut_sub lut_4182 ({i_6_, i_7_, g75, g357}, g358);
	defparam lut_4182.LUT_SIZE = 4;
	defparam lut_4182.mask = 16'haa8a;

	lut_sub lut_4194 ({g21, g110}, g359);
	defparam lut_4194.LUT_SIZE = 2;
	defparam lut_4194.mask = 4'b0100;

	lut_sub lut_4201 ({i_6_, i_7_, i_8_, g73, g184, g359}, g360);
	defparam lut_4201.LUT_SIZE = 6;
	defparam lut_4201.mask = 64'h553f0000000f0000;

	lut_sub lut_4221 ({g127, i_2_, i_6_, g137, g5}, g361);
	defparam lut_4221.LUT_SIZE = 5;
	defparam lut_4221.mask = 32'h00001001;

	lut_sub lut_4231 ({g11, g42, g22, g121, g361}, g362);
	defparam lut_4231.LUT_SIZE = 5;
	defparam lut_4231.mask = 32'h8880aaa0;

	lut_sub lut_4245 ({i_4_, i_5_, g23, g110}, g363);
	defparam lut_4245.LUT_SIZE = 4;
	defparam lut_4245.mask = 16'h0004;

	lut_sub lut_4252 ({g21, g6, g24}, g364);
	defparam lut_4252.LUT_SIZE = 3;
	defparam lut_4252.mask = 8'h20;

	lut_sub lut_4261 ({g21, g38, g7, g265, g364}, g365);
	defparam lut_4261.LUT_SIZE = 5;
	defparam lut_4261.mask = 32'h8088a0aa;

	lut_sub lut_4277 ({g175, g256, g363, g365}, g366);
	defparam lut_4277.LUT_SIZE = 4;
	defparam lut_4277.mask = 16'h4000;

	lut_sub lut_4286 ({g202, g358, g360, g362, g366}, g367);
	defparam lut_4286.LUT_SIZE = 5;
	defparam lut_4286.mask = 32'h00000010;

	lut_sub lut_4294 ({g11, g41, g28, g70}, g368);
	defparam lut_4294.LUT_SIZE = 4;
	defparam lut_4294.mask = 16'h1f11;

	lut_sub lut_4308 ({g50, i_6_, g14, g25, g129}, g369);
	defparam lut_4308.LUT_SIZE = 5;
	defparam lut_4308.mask = 32'h0005000d;

	lut_sub lut_4320 ({i_6_, g45, g1, g47, g110}, g370);
	defparam lut_4320.LUT_SIZE = 5;
	defparam lut_4320.mask = 32'h30001100;

	lut_sub lut_4332 ({g25, g159, g368, g369, g370}, g371);
	defparam lut_4332.LUT_SIZE = 5;
	defparam lut_4332.mask = 32'h80008080;

	lut_sub lut_4340 ({i_6_, i_7_, i_8_, g77, g99}, g372);
	defparam lut_4340.LUT_SIZE = 5;
	defparam lut_4340.mask = 32'h35000300;

	lut_sub lut_4352 ({g67, g116, g290}, g373);
	defparam lut_4352.LUT_SIZE = 3;
	defparam lut_4352.mask = 8'ha8;

	lut_sub lut_4363 ({g173, g294, g145, g140, g373}, g374);
	defparam lut_4363.LUT_SIZE = 5;
	defparam lut_4363.mask = 32'h10000000;

	lut_sub lut_4372 ({g23, g75, g160, g372, g374}, g375);
	defparam lut_4372.LUT_SIZE = 5;
	defparam lut_4372.mask = 32'h40004040;

	lut_sub lut_4383 ({g50, g35, g1, g12, g184}, g376);
	defparam lut_4383.LUT_SIZE = 5;
	defparam lut_4383.mask = 32'h00553075;

	lut_sub lut_4400 ({i_6_, i_7_, i_8_, g24, g64, g26}, g377);
	defparam lut_4400.LUT_SIZE = 6;
	defparam lut_4400.mask = 64'h5500553000000030;

	lut_sub lut_4420 ({g204, g376, g246, g249, g377}, g378);
	defparam lut_4420.LUT_SIZE = 5;
	defparam lut_4420.mask = 32'h02000000;

	lut_sub lut_4426 ({i_0_, i_1_, i_2_, g23, g123}, g379);
	defparam lut_4426.LUT_SIZE = 5;
	defparam lut_4426.mask = 32'h05050c00;

	lut_sub lut_4439 ({i_3_, g195, g379, g90, g618}, g380);
	defparam lut_4439.LUT_SIZE = 5;
	defparam lut_4439.mask = 32'h10001100;

	lut_sub lut_4451 ({g228, g330, g371, g375, g378, g380}, g381);
	defparam lut_4451.LUT_SIZE = 6;
	defparam lut_4451.mask = 64'h0000000000000001;

	lut_sub lut_4460 ({i_6_, g63, g21, g25, g110, g218}, g382);
	defparam lut_4460.LUT_SIZE = 6;
	defparam lut_4460.mask = 64'h0000f55500007755;

	lut_sub lut_4489 ({g27, g45, g6, g251, g287, g382}, g383);
	defparam lut_4489.LUT_SIZE = 6;
	defparam lut_4489.mask = 64'h0200020202020202;

	lut_sub lut_4505 ({g27, g42, g12, g48, g59, g38}, g384);
	defparam lut_4505.LUT_SIZE = 6;
	defparam lut_4505.mask = 64'h00cc0ace00000a0a;

	lut_sub lut_4528 ({g27, g21, g6, g3, g121}, g385);
	defparam lut_4528.LUT_SIZE = 5;
	defparam lut_4528.mask = 32'h57035500;

	lut_sub lut_4548 ({g45, g1, g2, g38, g384, g385}, g386);
	defparam lut_4548.LUT_SIZE = 6;
	defparam lut_4548.mask = 64'h8800888888088888;

	lut_sub lut_4567 ({g63, g42, g134}, g387);
	defparam lut_4567.LUT_SIZE = 3;
	defparam lut_4567.mask = 8'h01;

	lut_sub lut_4575 ({g1, g159, g150, g387}, g388);
	defparam lut_4575.LUT_SIZE = 4;
	defparam lut_4575.mask = 16'h8088;

	lut_sub lut_4585 ({g28, g110, g116, g141}, g389);
	defparam lut_4585.LUT_SIZE = 4;
	defparam lut_4585.mask = 16'h1113;

	lut_sub lut_4596 ({g18, g170, g389}, g390);
	defparam lut_4596.LUT_SIZE = 3;
	defparam lut_4596.mask = 8'h80;

	lut_sub lut_4602 ({g127, i_2_, i_6_, i_7_, i_8_, g3}, g391);
	defparam lut_4602.LUT_SIZE = 6;
	defparam lut_4602.mask = 64'h0000000004540404;

	lut_sub lut_4613 ({i_4_, i_5_, i_0_, i_1_, g8, g117}, g392);
	defparam lut_4613.LUT_SIZE = 6;
	defparam lut_4613.mask = 64'hececeeceeeeeeeee;

	lut_sub lut_4666 ({g344, g388, g390, g391, g583}, g393);
	defparam lut_4666.LUT_SIZE = 5;
	defparam lut_4666.mask = 32'h00040000;

	lut_sub lut_4675 ({g72, g166, g383, g386, g393}, g394);
	defparam lut_4675.LUT_SIZE = 5;
	defparam lut_4675.mask = 32'h00010000;

	lut_sub lut_4684 ({g274, g283, g367, g381, g394}, g395);
	defparam lut_4684.LUT_SIZE = 5;
	defparam lut_4684.mask = 32'h00000001;

	lut_sub lut_4692 ({g8, g32, g99, g265}, g396);
	defparam lut_4692.LUT_SIZE = 4;
	defparam lut_4692.mask = 16'h0537;

	lut_sub lut_4705 ({i_4_, g42, g12, g9}, g397);
	defparam lut_4705.LUT_SIZE = 4;
	defparam lut_4705.mask = 16'h5503;

	lut_sub lut_4716 ({i_3_, i_5_, g396, g397}, g398);
	defparam lut_4716.LUT_SIZE = 4;
	defparam lut_4716.mask = 16'hcc8c;

	lut_sub lut_4731 ({g21, g42, g12, g75, g124}, g399);
	defparam lut_4731.LUT_SIZE = 5;
	defparam lut_4731.mask = 32'ha8a0a8a8;

	lut_sub lut_4750 ({g2, g3, g9, g243, g399}, g400);
	defparam lut_4750.LUT_SIZE = 5;
	defparam lut_4750.mask = 32'h55504440;

	lut_sub lut_4763 ({i_3_, g50, i_0_, i_2_, i_6_}, g401);
	defparam lut_4763.LUT_SIZE = 5;
	defparam lut_4763.mask = 32'h00200000;

	lut_sub lut_4771 ({i_6_, g25, g137, g38, g401}, g402);
	defparam lut_4771.LUT_SIZE = 5;
	defparam lut_4771.mask = 32'h05050d05;

	lut_sub lut_4786 ({i_6_, i_7_, i_8_, g77, g71, g161}, g403);
	defparam lut_4786.LUT_SIZE = 6;
	defparam lut_4786.mask = 64'h003300007700000f;

	lut_sub lut_4807 ({g402, g93, g631, g403}, g404);
	defparam lut_4807.LUT_SIZE = 4;
	defparam lut_4807.mask = 16'h0200;

	lut_sub lut_4816 ({g149, g398, g242, g400, g404}, g405);
	defparam lut_4816.LUT_SIZE = 5;
	defparam lut_4816.mask = 32'h00010000;

	lut_sub lut_4821 ({i_3_, i_0_, i_2_, g85}, g406);
	defparam lut_4821.LUT_SIZE = 4;
	defparam lut_4821.mask = 16'h0010;

	lut_sub lut_4830 ({g50, g48, g88, g111, g230}, g407);
	defparam lut_4830.LUT_SIZE = 5;
	defparam lut_4830.mask = 32'h000f111f;

	lut_sub lut_4849 ({g14, g1, g22, g406, g407}, g408);
	defparam lut_4849.LUT_SIZE = 5;
	defparam lut_4849.mask = 32'ha0aa8088;

	lut_sub lut_4864 ({i_6_, i_7_, i_8_, g33, g184, g401}, g409);
	defparam lut_4864.LUT_SIZE = 6;
	defparam lut_4864.mask = 64'h0055000000550f33;

	lut_sub lut_4887 ({g35, g48, g117, g334}, g410);
	defparam lut_4887.LUT_SIZE = 4;
	defparam lut_4887.mask = 16'ha888;

	lut_sub lut_4896 ({i_4_, i_5_, i_0_, i_1_, g12}, g411);
	defparam lut_4896.LUT_SIZE = 5;
	defparam lut_4896.mask = 32'h10000000;

	lut_sub lut_4905 ({g8, g137, g91, g243, g411}, g412);
	defparam lut_4905.LUT_SIZE = 5;
	defparam lut_4905.mask = 32'haa88a080;

	lut_sub lut_4920 ({g2, g70, g158}, g413);
	defparam lut_4920.LUT_SIZE = 3;
	defparam lut_4920.mask = 8'h07;

	lut_sub lut_4930 ({i_5_, g6, g5, g110, g111}, g414);
	defparam lut_4930.LUT_SIZE = 5;
	defparam lut_4930.mask = 32'h01030003;

	lut_sub lut_4942 ({g23, g359, g413, g414}, g415);
	defparam lut_4942.LUT_SIZE = 4;
	defparam lut_4942.mask = 16'h8088;

	lut_sub lut_4953 ({g87, g346, g410, g412, g415}, g416);
	defparam lut_4953.LUT_SIZE = 5;
	defparam lut_4953.mask = 32'h01000000;

	lut_sub lut_4962 ({g254, g307, g289, g409, g416}, g417);
	defparam lut_4962.LUT_SIZE = 5;
	defparam lut_4962.mask = 32'h00000004;

	lut_sub lut_4970 ({g381, g405, g408, g417}, g418);
	defparam lut_4970.LUT_SIZE = 4;
	defparam lut_4970.mask = 16'h0001;

	lut_sub lut_4976 ({i_6_, i_7_, i_8_, g189, g406}, g419);
	defparam lut_4976.LUT_SIZE = 5;
	defparam lut_4976.mask = 32'h03530050;

	lut_sub lut_4987 ({i_0_, i_1_, i_2_, i_6_, i_7_, i_8_}, g420);
	defparam lut_4987.LUT_SIZE = 6;
	defparam lut_4987.mask = 64'h0010c00000000000;

	lut_sub lut_4995 ({i_0_, i_6_, g38, g420}, g421);
	defparam lut_4995.LUT_SIZE = 4;
	defparam lut_4995.mask = 16'h4000;

	lut_sub lut_5004 ({g28, g42, g45, g1, g32}, g422);
	defparam lut_5004.LUT_SIZE = 5;
	defparam lut_5004.mask = 32'h000044f4;

	lut_sub lut_5019 ({g27, g6, g36, g422, g572}, g423);
	defparam lut_5019.LUT_SIZE = 5;
	defparam lut_5019.mask = 32'h44044444;

	lut_sub lut_5034 ({g2, g38, g110, g421, g423}, g424);
	defparam lut_5034.LUT_SIZE = 5;
	defparam lut_5034.mask = 32'h44444044;

	lut_sub lut_5046 ({i_6_, i_8_, g21, g1}, g425);
	defparam lut_5046.LUT_SIZE = 4;
	defparam lut_5046.mask = 16'h8000;

	lut_sub lut_5053 ({i_6_, g14, g32, g110}, g426);
	defparam lut_5053.LUT_SIZE = 4;
	defparam lut_5053.mask = 16'h0111;

	lut_sub lut_5063 ({g24, g4, g425, g426}, g427);
	defparam lut_5063.LUT_SIZE = 4;
	defparam lut_5063.mask = 16'h8088;

	lut_sub lut_5070 ({i_3_, i_0_, i_2_, g123}, g428);
	defparam lut_5070.LUT_SIZE = 4;
	defparam lut_5070.mask = 16'h0100;

	lut_sub lut_5077 ({g11, g29, g428}, g429);
	defparam lut_5077.LUT_SIZE = 3;
	defparam lut_5077.mask = 8'h8a;

	lut_sub lut_5087 ({g63, g45, g129, g141}, g430);
	defparam lut_5087.LUT_SIZE = 4;
	defparam lut_5087.mask = 16'h5073;

	lut_sub lut_5101 ({g35, g1, g16, g161}, g431);
	defparam lut_5101.LUT_SIZE = 4;
	defparam lut_5101.mask = 16'h3075;

	lut_sub lut_5116 ({i_7_, g8, g25, g32, g97, g217}, g432);
	defparam lut_5116.LUT_SIZE = 6;
	defparam lut_5116.mask = 64'hccccc0cc88cc80cc;

	lut_sub lut_5147 ({i_1_, g6, g33, g38}, g433);
	defparam lut_5147.LUT_SIZE = 4;
	defparam lut_5147.mask = 16'h030b;

	lut_sub lut_5161 ({g35, g189, g229, g431, g432, g433}, g434);
	defparam lut_5161.LUT_SIZE = 6;
	defparam lut_5161.mask = 64'h2000200020000000;

	lut_sub lut_5172 ({g352, g332, g429, g430, g434}, g435);
	defparam lut_5172.LUT_SIZE = 5;
	defparam lut_5172.mask = 32'h00040000;

	lut_sub lut_5181 ({g419, g367, g424, g427, g435}, g436);
	defparam lut_5181.LUT_SIZE = 5;
	defparam lut_5181.mask = 32'h00010000;

	lut_sub lut_5190 ({g31, g300, g371, g405, g436}, g437);
	defparam lut_5190.LUT_SIZE = 5;
	defparam lut_5190.mask = 32'h00000001;

	lut_sub lut_5197 ({g48, g33, g368}, g438);
	defparam lut_5197.LUT_SIZE = 3;
	defparam lut_5197.mask = 8'ha8;

	lut_sub lut_5208 ({g21, g1, g2, g24, g36}, g439);
	defparam lut_5208.LUT_SIZE = 5;
	defparam lut_5208.mask = 32'h0e0c0a00;

	lut_sub lut_5218 ({i_3_, i_1_, i_2_}, g440);
	defparam lut_5218.LUT_SIZE = 3;
	defparam lut_5218.mask = 8'h40;

	lut_sub lut_5225 ({g137, g15, g440}, g441);
	defparam lut_5225.LUT_SIZE = 3;
	defparam lut_5225.mask = 8'h01;

	lut_sub lut_5234 ({g6, g5, g110, g99, g441}, g442);
	defparam lut_5234.LUT_SIZE = 5;
	defparam lut_5234.mask = 32'haaaa8880;

	lut_sub lut_5253 ({g35, g161, g376, g439, g442}, g443);
	defparam lut_5253.LUT_SIZE = 5;
	defparam lut_5253.mask = 32'h40404000;

	lut_sub lut_5262 ({i_8_, g65, g247, g398}, g444);
	defparam lut_5262.LUT_SIZE = 4;
	defparam lut_5262.mask = 16'h4440;

	lut_sub lut_5273 ({g266, g438, g358, g443, g444}, g445);
	defparam lut_5273.LUT_SIZE = 5;
	defparam lut_5273.mask = 32'h00010000;

	lut_sub lut_5278 ({i_3_, i_1_, i_2_, i_7_, g64}, g446);
	defparam lut_5278.LUT_SIZE = 5;
	defparam lut_5278.mask = 32'h00000010;

	lut_sub lut_5287 ({g14, g24, g64, g194, g446}, g447);
	defparam lut_5287.LUT_SIZE = 5;
	defparam lut_5287.mask = 32'h88aa80aa;

	lut_sub lut_5305 ({g25, g2, g38, g110}, g448);
	defparam lut_5305.LUT_SIZE = 4;
	defparam lut_5305.mask = 16'hf3fb;

	lut_sub lut_5325 ({i_5_, g6, g23, g110, g440}, g449);
	defparam lut_5325.LUT_SIZE = 5;
	defparam lut_5325.mask = 32'haf8cffff;

	lut_sub lut_5357 ({g255, g384, g310, g559}, g450);
	defparam lut_5357.LUT_SIZE = 4;
	defparam lut_5357.mask = 16'h1000;

	lut_sub lut_5365 ({g50, i_6_, i_8_, g5, g13, g17}, g451);
	defparam lut_5365.LUT_SIZE = 6;
	defparam lut_5365.mask = 64'h0000000c0055000c;

	lut_sub lut_5381 ({g275, g402, g670, g147, g451}, g452);
	defparam lut_5381.LUT_SIZE = 5;
	defparam lut_5381.mask = 32'h02000000;

	lut_sub lut_5391 ({g80, g291, g383, g427, g450, g452}, g453);
	defparam lut_5391.LUT_SIZE = 6;
	defparam lut_5391.mask = 64'h0000000000000001;

	lut_sub lut_5400 ({g109, g341, g408, g445, g453}, g454);
	defparam lut_5400.LUT_SIZE = 5;
	defparam lut_5400.mask = 32'h00000001;

	lut_sub lut_5408 ({g127, i_2_, g2, g60, g38}, g455);
	defparam lut_5408.LUT_SIZE = 5;
	defparam lut_5408.mask = 32'h00000a22;

	lut_sub lut_5420 ({g23, g66, g189, g455, g315}, g456);
	defparam lut_5420.LUT_SIZE = 5;
	defparam lut_5420.mask = 32'h80008800;

	lut_sub lut_5431 ({g2, g36, g38, g110, g121}, g457);
	defparam lut_5431.LUT_SIZE = 5;
	defparam lut_5431.mask = 32'h50507350;

	lut_sub lut_5448 ({g63, g64, g17}, g458);
	defparam lut_5448.LUT_SIZE = 3;
	defparam lut_5448.mask = 8'h01;

	lut_sub lut_5458 ({g267, g313, g389, g419, g457, g458}, g459);
	defparam lut_5458.LUT_SIZE = 6;
	defparam lut_5458.mask = 64'h8000000000000000;

	lut_sub lut_5463 ({i_4_, i_5_, i_1_, i_2_, i_6_, g14}, g460);
	defparam lut_5463.LUT_SIZE = 6;
	defparam lut_5463.mask = 64'h0000000500000100;

	lut_sub lut_5470 ({i_3_, i_6_, i_8_, g13}, g461);
	defparam lut_5470.LUT_SIZE = 4;
	defparam lut_5470.mask = 16'h8000;

	lut_sub lut_5478 ({g27, g28, g36, g461}, g462);
	defparam lut_5478.LUT_SIZE = 4;
	defparam lut_5478.mask = 16'ha2aa;

	lut_sub lut_5490 ({i_6_, i_7_, i_8_, g71, g26}, g463);
	defparam lut_5490.LUT_SIZE = 5;
	defparam lut_5490.mask = 32'h53500050;

	lut_sub lut_5505 ({g50, g47, g94, g401}, g464);
	defparam lut_5505.LUT_SIZE = 4;
	defparam lut_5505.mask = 16'h0507;

	lut_sub lut_5518 ({g292, g327, g363, g463, g464}, g465);
	defparam lut_5518.LUT_SIZE = 5;
	defparam lut_5518.mask = 32'h00800000;

	lut_sub lut_5527 ({g34, g323, g460, g462, g465}, g466);
	defparam lut_5527.LUT_SIZE = 5;
	defparam lut_5527.mask = 32'h00100000;

	lut_sub lut_5537 ({g154, g216, g445, g456, g459, g466}, g467);
	defparam lut_5537.LUT_SIZE = 6;
	defparam lut_5537.mask = 64'h0000000000000001;

	lut_sub lut_5545 ({g8, g45, g13, g165}, g468);
	defparam lut_5545.LUT_SIZE = 4;
	defparam lut_5545.mask = 16'haa2a;

	lut_sub lut_5560 ({g21, g6, g23, g24, g3}, g469);
	defparam lut_5560.LUT_SIZE = 5;
	defparam lut_5560.mask = 32'hc0c40044;

	lut_sub lut_5575 ({g8, g2, g26, g239, g469}, g470);
	defparam lut_5575.LUT_SIZE = 5;
	defparam lut_5575.mask = 32'h88808080;

	lut_sub lut_5588 ({g102, g208, g278, g40, g470}, g471);
	defparam lut_5588.LUT_SIZE = 5;
	defparam lut_5588.mask = 32'h10000000;

	lut_sub lut_5592 ({i_3_, i_0_, i_1_}, g472);
	defparam lut_5592.LUT_SIZE = 3;
	defparam lut_5592.mask = 8'h80;

	lut_sub lut_5599 ({i_4_, i_6_, g4, g110, g472}, g473);
	defparam lut_5599.LUT_SIZE = 5;
	defparam lut_5599.mask = 32'h57030303;

	lut_sub lut_5617 ({g42, g38, g29, g159}, g474);
	defparam lut_5617.LUT_SIZE = 4;
	defparam lut_5617.mask = 16'h3075;

	lut_sub lut_5632 ({g694, g473, g400, g409, g474}, g475);
	defparam lut_5632.LUT_SIZE = 5;
	defparam lut_5632.mask = 32'h00000800;

	lut_sub lut_5641 ({g36, g121, g468, g471, g475}, g476);
	defparam lut_5641.LUT_SIZE = 5;
	defparam lut_5641.mask = 32'h01000101;

	lut_sub lut_5650 ({g50, i_6_, g63, g440}, g477);
	defparam lut_5650.LUT_SIZE = 4;
	defparam lut_5650.mask = 16'h0001;

	lut_sub lut_5657 ({i_6_, i_7_, i_8_, g181, g105, g359}, g478);
	defparam lut_5657.LUT_SIZE = 6;
	defparam lut_5657.mask = 64'h0000000f0fcc5500;

	lut_sub lut_5681 ({g41, g32, g343, g549, g478}, g479);
	defparam lut_5681.LUT_SIZE = 5;
	defparam lut_5681.mask = 32'h02020200;

	lut_sub lut_5692 ({g43, g92, g257, g477, g479}, g480);
	defparam lut_5692.LUT_SIZE = 5;
	defparam lut_5692.mask = 32'h04000000;

	lut_sub lut_5701 ({g46, g60, g226, g396, g456}, g481);
	defparam lut_5701.LUT_SIZE = 5;
	defparam lut_5701.mask = 32'h40404000;

	lut_sub lut_5712 ({g101, g152, g424, g480, g481}, g482);
	defparam lut_5712.LUT_SIZE = 5;
	defparam lut_5712.mask = 32'h00010000;

	lut_sub lut_5721 ({g21, g12, g6, g13, g110}, g483);
	defparam lut_5721.LUT_SIZE = 5;
	defparam lut_5721.mask = 32'h05cd0000;

	lut_sub lut_5736 ({g28, g25, g12, g32, g36}, g484);
	defparam lut_5736.LUT_SIZE = 5;
	defparam lut_5736.mask = 32'h0300ab00;

	lut_sub lut_5752 ({g11, g27, g45, g48, g2, g24}, g485);
	defparam lut_5752.LUT_SIZE = 6;
	defparam lut_5752.mask = 64'h3b222a223b000a00;

	lut_sub lut_5780 ({g1, g6, g23, g3, g49, g110}, g486);
	defparam lut_5780.LUT_SIZE = 6;
	defparam lut_5780.mask = 64'h0f003f3700003737;

	lut_sub lut_5813 ({g155, g483, g484, g485, g486}, g487);
	defparam lut_5813.LUT_SIZE = 5;
	defparam lut_5813.mask = 32'h80000000;

	lut_sub lut_5819 ({i_6_, i_7_, g188, g129}, g488);
	defparam lut_5819.LUT_SIZE = 4;
	defparam lut_5819.mask = 16'hcc8c;

	lut_sub lut_5833 ({i_6_, g32, g18, g110, g488}, g489);
	defparam lut_5833.LUT_SIZE = 5;
	defparam lut_5833.mask = 32'h50505040;

	lut_sub lut_5847 ({g476, g482, g487, g489}, g490);
	defparam lut_5847.LUT_SIZE = 4;
	defparam lut_5847.mask = 16'h0001;

	lut_sub lut_5853 ({i_5_, g48, g472}, g491);
	defparam lut_5853.LUT_SIZE = 3;
	defparam lut_5853.mask = 8'h10;

	lut_sub lut_5861 ({g1, g12, g3, g290}, g492);
	defparam lut_5861.LUT_SIZE = 4;
	defparam lut_5861.mask = 16'ha8aa;

	lut_sub lut_5876 ({g11, g41, g45, g29, g141}, g493);
	defparam lut_5876.LUT_SIZE = 5;
	defparam lut_5876.mask = 32'h8a0acf0f;

	lut_sub lut_5899 ({g21, g48, g49, g110, g364}, g494);
	defparam lut_5899.LUT_SIZE = 5;
	defparam lut_5899.mask = 32'haa80aaa0;

	lut_sub lut_5918 ({g23, g184, g492, g493, g494}, g495);
	defparam lut_5918.LUT_SIZE = 5;
	defparam lut_5918.mask = 32'h01000101;

	lut_sub lut_5929 ({g23, g91, g296, g491, g495}, g496);
	defparam lut_5929.LUT_SIZE = 5;
	defparam lut_5929.mask = 32'h40004040;

	lut_sub lut_5939 ({g11, i_6_, g2, g32, g110}, g497);
	defparam lut_5939.LUT_SIZE = 5;
	defparam lut_5939.mask = 32'h05150011;

	lut_sub lut_5954 ({g35, g74, g189, g359, g497}, g498);
	defparam lut_5954.LUT_SIZE = 5;
	defparam lut_5954.mask = 32'haa008000;

	lut_sub lut_5963 ({i_0_, i_1_, i_2_, g194}, g499);
	defparam lut_5963.LUT_SIZE = 4;
	defparam lut_5963.mask = 16'hc400;

	lut_sub lut_5974 ({g35, g25, g22, g36, g499}, g500);
	defparam lut_5974.LUT_SIZE = 5;
	defparam lut_5974.mask = 32'ha0aa20aa;

	lut_sub lut_5993 ({g23, g71, g294, g88, g212}, g501);
	defparam lut_5993.LUT_SIZE = 5;
	defparam lut_5993.mask = 32'h8000a0a0;

	lut_sub lut_6006 ({g27, g12, g33, g4, g194}, g502);
	defparam lut_6006.LUT_SIZE = 5;
	defparam lut_6006.mask = 32'h8880fff0;

	lut_sub lut_6029 ({g174, g277, g500, g501, g502}, g503);
	defparam lut_6029.LUT_SIZE = 5;
	defparam lut_6029.mask = 32'h01000000;

	lut_sub lut_6037 ({g6, g59, g88, g265}, g504);
	defparam lut_6037.LUT_SIZE = 4;
	defparam lut_6037.mask = 16'h5073;

	lut_sub lut_6051 ({g37, g129, g386, g504}, g505);
	defparam lut_6051.LUT_SIZE = 4;
	defparam lut_6051.mask = 16'h2220;

	lut_sub lut_6062 ({g179, g438, g498, g503, g505}, g506);
	defparam lut_6062.LUT_SIZE = 5;
	defparam lut_6062.mask = 32'h00010000;

	lut_sub lut_6069 ({g35, g45, g13}, g507);
	defparam lut_6069.LUT_SIZE = 3;
	defparam lut_6069.mask = 8'h08;

	lut_sub lut_6077 ({i_3_, g50, g127, g8, g84}, g508);
	defparam lut_6077.LUT_SIZE = 5;
	defparam lut_6077.mask = 32'h11131111;

	lut_sub lut_6094 ({g63, g6, g129, g507, g508}, g509);
	defparam lut_6094.LUT_SIZE = 5;
	defparam lut_6094.mask = 32'h88808080;

	lut_sub lut_6106 ({g476, g496, g506, g509}, g510);
	defparam lut_6106.LUT_SIZE = 4;
	defparam lut_6106.mask = 16'h0001;

	lut_sub lut_6116 ({g21, g25, g48, g2, g13, g38}, g511);
	defparam lut_6116.LUT_SIZE = 6;
	defparam lut_6116.mask = 64'h0eff0c0c0a0a0000;

	lut_sub lut_6142 ({g42, g12, g59, g7}, g512);
	defparam lut_6142.LUT_SIZE = 4;
	defparam lut_6142.mask = 16'h444c;

	lut_sub lut_6154 ({g27, g45, g23, g512}, g513);
	defparam lut_6154.LUT_SIZE = 4;
	defparam lut_6154.mask = 16'h2aaa;

	lut_sub lut_6169 ({g41, g21, g3, g29, g265}, g514);
	defparam lut_6169.LUT_SIZE = 5;
	defparam lut_6169.mask = 32'ha8f8a0f0;

	lut_sub lut_6191 ({g134, g413, g457, g472, g514}, g515);
	defparam lut_6191.LUT_SIZE = 5;
	defparam lut_6191.mask = 32'h50004000;

	lut_sub lut_6201 ({g28, g32, g67, g181}, g516);
	defparam lut_6201.LUT_SIZE = 4;
	defparam lut_6201.mask = 16'h0357;

	lut_sub lut_6215 ({g314, g293, g236, g516}, g517);
	defparam lut_6215.LUT_SIZE = 4;
	defparam lut_6215.mask = 16'h2000;

	lut_sub lut_6224 ({g122, g511, g513, g543, g517}, g518);
	defparam lut_6224.LUT_SIZE = 5;
	defparam lut_6224.mask = 32'h01000000;

	lut_sub lut_6232 ({g13, g123, g387, g458}, g519);
	defparam lut_6232.LUT_SIZE = 4;
	defparam lut_6232.mask = 16'h8088;

	lut_sub lut_6243 ({g431, g487, g506, g518, g519}, g520);
	defparam lut_6243.LUT_SIZE = 5;
	defparam lut_6243.mask = 32'h00010000;

	lut_sub lut_6250 ({g8, g117, g428}, g521);
	defparam lut_6250.LUT_SIZE = 3;
	defparam lut_6250.mask = 8'ha8;

	lut_sub lut_6260 ({i_4_, i_5_, g63, g65, g472, g521}, g522);
	defparam lut_6260.LUT_SIZE = 6;
	defparam lut_6260.mask = 64'h5540555055505550;

	lut_sub lut_6290 ({g482, g496, g518, g522}, g523);
	defparam lut_6290.LUT_SIZE = 4;
	defparam lut_6290.mask = 16'h0001;

	lut_sub lut_6299 ({g28, g25, g38, g110, g159}, g524);
	defparam lut_6299.LUT_SIZE = 5;
	defparam lut_6299.mask = 32'h1111f111;

	lut_sub lut_6316 ({i_6_, i_7_, i_8_, g45, g3, g110}, g525);
	defparam lut_6316.LUT_SIZE = 6;
	defparam lut_6316.mask = 64'h0000000050505150;

	lut_sub lut_6331 ({i_6_, i_7_, i_8_, g21, g25, g110}, g526);
	defparam lut_6331.LUT_SIZE = 6;
	defparam lut_6331.mask = 64'h0000d0c00000c0c0;

	lut_sub lut_6345 ({i_6_, i_7_, i_8_, g46, g184}, g527);
	defparam lut_6345.LUT_SIZE = 5;
	defparam lut_6345.mask = 32'h75500000;

	lut_sub lut_6359 ({g500, g525, g526, g527}, g528);
	defparam lut_6359.LUT_SIZE = 4;
	defparam lut_6359.mask = 16'h0080;

	lut_sub lut_6365 ({i_6_, i_7_, i_8_, g189, g161}, g529);
	defparam lut_6365.LUT_SIZE = 5;
	defparam lut_6365.mask = 32'h00330755;

	lut_sub lut_6383 ({g25, g23, g38, g491}, g530);
	defparam lut_6383.LUT_SIZE = 4;
	defparam lut_6383.mask = 16'h2aaa;

	lut_sub lut_6397 ({g473, g498, g529, g530}, g531);
	defparam lut_6397.LUT_SIZE = 4;
	defparam lut_6397.mask = 16'h0400;

	lut_sub lut_6404 ({g524, g528, g531}, g532);
	defparam lut_6404.LUT_SIZE = 3;
	defparam lut_6404.mask = 8'h10;

	lut_sub lut_6413 ({g35, g23, g36, g110, g99}, g533);
	defparam lut_6413.LUT_SIZE = 5;
	defparam lut_6413.mask = 32'h55007530;

	lut_sub lut_6429 ({i_0_, i_1_, i_2_, g2, g59}, g534);
	defparam lut_6429.LUT_SIZE = 5;
	defparam lut_6429.mask = 32'hf0200000;

	lut_sub lut_6441 ({g6, g23, g189, g99}, g535);
	defparam lut_6441.LUT_SIZE = 4;
	defparam lut_6441.mask = 16'h3075;

	lut_sub lut_6456 ({g28, g38, g110, g534, g535}, g536);
	defparam lut_6456.LUT_SIZE = 5;
	defparam lut_6456.mask = 32'h88888088;

	lut_sub lut_6469 ({g533, g531, g536}, g537);
	defparam lut_6469.LUT_SIZE = 3;
	defparam lut_6469.mask = 8'h10;

	lut_sub lut_6477 ({g8, g46, g2, g26}, g538);
	defparam lut_6477.LUT_SIZE = 4;
	defparam lut_6477.mask = 16'h111f;

	lut_sub lut_6490 ({i_4_, i_6_, g6, g161, g472}, g539);
	defparam lut_6490.LUT_SIZE = 5;
	defparam lut_6490.mask = 32'h57030303;

	lut_sub lut_6509 ({g497, g524, g538, g536, g539}, g540);
	defparam lut_6509.LUT_SIZE = 5;
	defparam lut_6509.mask = 32'h20000000;

	lut_sub lut_6515 ({i_4_, i_5_, i_6_, g63, g472}, g541);
	defparam lut_6515.LUT_SIZE = 5;
	defparam lut_6515.mask = 32'h51000000;

	lut_sub lut_6525 ({g533, g538, g541, g528}, g542);
	defparam lut_6525.LUT_SIZE = 4;
	defparam lut_6525.mask = 16'h4000;

	lut_sub lut_6531 ({g515, g544}, g543);
	defparam lut_6531.LUT_SIZE = 2;
	defparam lut_6531.mask = 4'b0001;

	lut_sub lut_6537 ({g545, g546}, g544);
	defparam lut_6537.LUT_SIZE = 2;
	defparam lut_6537.mask = 4'b1000;

	lut_sub lut_6542 ({i_6_, g547}, g545);
	defparam lut_6542.LUT_SIZE = 2;
	defparam lut_6542.mask = 4'b0100;

	lut_sub lut_6547 ({i_6_, g548}, g546);
	defparam lut_6547.LUT_SIZE = 2;
	defparam lut_6547.mask = 4'b0001;

	lut_sub lut_6552 ({i_8_, g88, i_7_}, g547);
	defparam lut_6552.LUT_SIZE = 3;
	defparam lut_6552.mask = 8'hed;

	lut_sub lut_6563 ({g98, i_8_, g73, i_7_}, g548);
	defparam lut_6563.LUT_SIZE = 4;
	defparam lut_6563.mask = 16'hefaf;

	lut_sub lut_6581 ({g550, g551}, g549);
	defparam lut_6581.LUT_SIZE = 2;
	defparam lut_6581.mask = 4'b1000;

	lut_sub lut_6586 ({i_0_, g552}, g550);
	defparam lut_6586.LUT_SIZE = 2;
	defparam lut_6586.mask = 4'b0100;

	lut_sub lut_6591 ({i_0_, g554}, g551);
	defparam lut_6591.LUT_SIZE = 2;
	defparam lut_6591.mask = 4'b0001;

	lut_sub lut_6596 ({i_1_, g553}, g552);
	defparam lut_6596.LUT_SIZE = 2;
	defparam lut_6596.mask = 4'b1000;

	lut_sub lut_6600 ({i_1_, i_2_}, g553);
	defparam lut_6600.LUT_SIZE = 2;
	defparam lut_6600.mask = 4'b0100;

	lut_sub lut_6606 ({g555, g556}, g554);
	defparam lut_6606.LUT_SIZE = 2;
	defparam lut_6606.mask = 4'b1000;

	lut_sub lut_6611 ({i_1_, g557}, g555);
	defparam lut_6611.LUT_SIZE = 2;
	defparam lut_6611.mask = 4'b0100;

	lut_sub lut_6616 ({i_1_, g558}, g556);
	defparam lut_6616.LUT_SIZE = 2;
	defparam lut_6616.mask = 4'b0001;

	lut_sub lut_6623 ({g36, g23, g6, i_2_}, g557);
	defparam lut_6623.LUT_SIZE = 4;
	defparam lut_6623.mask = 16'h5dff;

	lut_sub lut_6640 ({g16, i_2_}, g558);
	defparam lut_6640.LUT_SIZE = 2;
	defparam lut_6640.mask = 4'b1101;

	lut_sub lut_6648 ({g560, g561}, g559);
	defparam lut_6648.LUT_SIZE = 2;
	defparam lut_6648.mask = 4'b1000;

	lut_sub lut_6654 ({g243, g562}, g560);
	defparam lut_6654.LUT_SIZE = 2;
	defparam lut_6654.mask = 4'b0100;

	lut_sub lut_6660 ({g243, g565}, g561);
	defparam lut_6660.LUT_SIZE = 2;
	defparam lut_6660.mask = 4'b0001;

	lut_sub lut_6666 ({g563, g564}, g562);
	defparam lut_6666.LUT_SIZE = 2;
	defparam lut_6666.mask = 4'b1000;

	lut_sub lut_6671 ({i_8_, g568}, g563);
	defparam lut_6671.LUT_SIZE = 2;
	defparam lut_6671.mask = 4'b0100;

	lut_sub lut_6676 ({i_8_, g569}, g564);
	defparam lut_6676.LUT_SIZE = 2;
	defparam lut_6676.mask = 4'b0001;

	lut_sub lut_6682 ({g566, g567}, g565);
	defparam lut_6682.LUT_SIZE = 2;
	defparam lut_6682.mask = 4'b1000;

	lut_sub lut_6687 ({i_8_, g570}, g566);
	defparam lut_6687.LUT_SIZE = 2;
	defparam lut_6687.mask = 4'b0100;

	lut_sub lut_6692 ({i_8_, g571}, g567);
	defparam lut_6692.LUT_SIZE = 2;
	defparam lut_6692.mask = 4'b0001;

	lut_sub lut_6699 ({g448, g449, g447}, g568);
	defparam lut_6699.LUT_SIZE = 3;
	defparam lut_6699.mask = 8'h01;

	lut_sub lut_6706 ({g448, g449, g447}, g569);
	defparam lut_6706.LUT_SIZE = 3;
	defparam lut_6706.mask = 8'h01;

	lut_sub lut_6713 ({g448, g449, i_7_, g447}, g570);
	defparam lut_6713.LUT_SIZE = 4;
	defparam lut_6713.mask = 16'h0001;

	lut_sub lut_6720 ({g448, g449, i_6_, g447}, g571);
	defparam lut_6720.LUT_SIZE = 4;
	defparam lut_6720.mask = 16'h0001;

	lut_sub lut_6726 ({g573, g574}, g572);
	defparam lut_6726.LUT_SIZE = 2;
	defparam lut_6726.mask = 4'b1000;

	lut_sub lut_6731 ({i_6_, g575}, g573);
	defparam lut_6731.LUT_SIZE = 2;
	defparam lut_6731.mask = 4'b0100;

	lut_sub lut_6736 ({i_6_, g578}, g574);
	defparam lut_6736.LUT_SIZE = 2;
	defparam lut_6736.mask = 4'b0001;

	lut_sub lut_6742 ({g576, g577}, g575);
	defparam lut_6742.LUT_SIZE = 2;
	defparam lut_6742.mask = 4'b1000;

	lut_sub lut_6747 ({i_8_, g580}, g576);
	defparam lut_6747.LUT_SIZE = 2;
	defparam lut_6747.mask = 4'b0100;

	lut_sub lut_6752 ({i_8_, g581}, g577);
	defparam lut_6752.LUT_SIZE = 2;
	defparam lut_6752.mask = 4'b0001;

	lut_sub lut_6757 ({i_8_, g579}, g578);
	defparam lut_6757.LUT_SIZE = 2;
	defparam lut_6757.mask = 4'b1000;

	lut_sub lut_6762 ({i_8_, g582}, g579);
	defparam lut_6762.LUT_SIZE = 2;
	defparam lut_6762.mask = 4'b0100;

	lut_sub lut_6768 ({g59, g25, i_7_}, g580);
	defparam lut_6768.LUT_SIZE = 3;
	defparam lut_6768.mask = 8'h7f;

	lut_sub lut_6780 ({g59, g13}, g581);
	defparam lut_6780.LUT_SIZE = 2;
	defparam lut_6780.mask = 4'b0111;

	lut_sub lut_6787 ({i_7_, g105}, g582);
	defparam lut_6787.LUT_SIZE = 2;
	defparam lut_6787.mask = 4'b0111;

	lut_sub lut_6795 ({g584, g585}, g583);
	defparam lut_6795.LUT_SIZE = 2;
	defparam lut_6795.mask = 4'b1000;

	lut_sub lut_6801 ({g359, g586}, g584);
	defparam lut_6801.LUT_SIZE = 2;
	defparam lut_6801.mask = 4'b0100;

	lut_sub lut_6807 ({g359, g589}, g585);
	defparam lut_6807.LUT_SIZE = 2;
	defparam lut_6807.mask = 4'b0001;

	lut_sub lut_6813 ({g587, g588}, g586);
	defparam lut_6813.LUT_SIZE = 2;
	defparam lut_6813.mask = 4'b1000;

	lut_sub lut_6818 ({i_6_, g592}, g587);
	defparam lut_6818.LUT_SIZE = 2;
	defparam lut_6818.mask = 4'b0100;

	lut_sub lut_6823 ({i_6_, g593}, g588);
	defparam lut_6823.LUT_SIZE = 2;
	defparam lut_6823.mask = 4'b0001;

	lut_sub lut_6829 ({g590, g591}, g589);
	defparam lut_6829.LUT_SIZE = 2;
	defparam lut_6829.mask = 4'b1000;

	lut_sub lut_6834 ({i_6_, g594}, g590);
	defparam lut_6834.LUT_SIZE = 2;
	defparam lut_6834.mask = 4'b0100;

	lut_sub lut_6839 ({i_6_, g595}, g591);
	defparam lut_6839.LUT_SIZE = 2;
	defparam lut_6839.mask = 4'b0001;

	lut_sub lut_6845 ({i_8_, i_7_, g105, g392}, g592);
	defparam lut_6845.LUT_SIZE = 4;
	defparam lut_6845.mask = 16'h5155;

	lut_sub lut_6857 ({i_8_, i_7_, g98, g392}, g593);
	defparam lut_6857.LUT_SIZE = 4;
	defparam lut_6857.mask = 16'h4454;

	lut_sub lut_6866 ({i_8_, i_7_, g392}, g594);
	defparam lut_6866.LUT_SIZE = 3;
	defparam lut_6866.mask = 8'h45;

	lut_sub lut_6874 ({i_8_, i_7_, g98, g392}, g595);
	defparam lut_6874.LUT_SIZE = 4;
	defparam lut_6874.mask = 16'h4454;

	lut_sub lut_6884 ({g597, g598}, g596);
	defparam lut_6884.LUT_SIZE = 2;
	defparam lut_6884.mask = 4'b1000;

	lut_sub lut_6889 ({i_6_, g599}, g597);
	defparam lut_6889.LUT_SIZE = 2;
	defparam lut_6889.mask = 4'b0100;

	lut_sub lut_6894 ({i_6_, g601}, g598);
	defparam lut_6894.LUT_SIZE = 2;
	defparam lut_6894.mask = 4'b0001;

	lut_sub lut_6899 ({i_7_, g600}, g599);
	defparam lut_6899.LUT_SIZE = 2;
	defparam lut_6899.mask = 4'b1000;

	lut_sub lut_6904 ({i_7_, g604}, g600);
	defparam lut_6904.LUT_SIZE = 2;
	defparam lut_6904.mask = 4'b0100;

	lut_sub lut_6910 ({g602, g603}, g601);
	defparam lut_6910.LUT_SIZE = 2;
	defparam lut_6910.mask = 4'b1000;

	lut_sub lut_6915 ({i_7_, g605}, g602);
	defparam lut_6915.LUT_SIZE = 2;
	defparam lut_6915.mask = 4'b0100;

	lut_sub lut_6920 ({i_7_, g606}, g603);
	defparam lut_6920.LUT_SIZE = 2;
	defparam lut_6920.mask = 4'b0001;

	lut_sub lut_6926 ({g59, g25, i_8_}, g604);
	defparam lut_6926.LUT_SIZE = 3;
	defparam lut_6926.mask = 8'hbf;

	lut_sub lut_6937 ({g98, i_8_}, g605);
	defparam lut_6937.LUT_SIZE = 2;
	defparam lut_6937.mask = 4'b1110;

	lut_sub lut_6945 ({g25, g21}, g606);
	defparam lut_6945.LUT_SIZE = 2;
	defparam lut_6945.mask = 4'b0111;

	lut_sub lut_6953 ({g608, g609}, g607);
	defparam lut_6953.LUT_SIZE = 2;
	defparam lut_6953.mask = 4'b1000;

	lut_sub lut_6959 ({g6, g610}, g608);
	defparam lut_6959.LUT_SIZE = 2;
	defparam lut_6959.mask = 4'b0100;

	lut_sub lut_6965 ({g6, g612}, g609);
	defparam lut_6965.LUT_SIZE = 2;
	defparam lut_6965.mask = 4'b0001;

	lut_sub lut_6971 ({g11, g611}, g610);
	defparam lut_6971.LUT_SIZE = 2;
	defparam lut_6971.mask = 4'b1000;

	lut_sub lut_6977 ({g11, g615}, g611);
	defparam lut_6977.LUT_SIZE = 2;
	defparam lut_6977.mask = 4'b0100;

	lut_sub lut_6983 ({g613, g614}, g612);
	defparam lut_6983.LUT_SIZE = 2;
	defparam lut_6983.mask = 4'b1000;

	lut_sub lut_6989 ({g11, g616}, g613);
	defparam lut_6989.LUT_SIZE = 2;
	defparam lut_6989.mask = 4'b0100;

	lut_sub lut_6995 ({g11, g617}, g614);
	defparam lut_6995.LUT_SIZE = 2;
	defparam lut_6995.mask = 4'b0001;

	lut_sub lut_7001 ({g13, g47}, g615);
	defparam lut_7001.LUT_SIZE = 2;
	defparam lut_7001.mask = 4'b1011;

	lut_sub lut_7011 ({g13, g24, g47, g99}, g616);
	defparam lut_7011.LUT_SIZE = 4;
	defparam lut_7011.mask = 16'h080a;

	lut_sub lut_7020 ({g24, g36, g99}, g617);
	defparam lut_7020.LUT_SIZE = 3;
	defparam lut_7020.mask = 8'h2a;

	lut_sub lut_7028 ({g619, g620}, g618);
	defparam lut_7028.LUT_SIZE = 2;
	defparam lut_7028.mask = 4'b1000;

	lut_sub lut_7034 ({g11, g621}, g619);
	defparam lut_7034.LUT_SIZE = 2;
	defparam lut_7034.mask = 4'b0100;

	lut_sub lut_7040 ({g11, g624}, g620);
	defparam lut_7040.LUT_SIZE = 2;
	defparam lut_7040.mask = 4'b0001;

	lut_sub lut_7046 ({g622, g623}, g621);
	defparam lut_7046.LUT_SIZE = 2;
	defparam lut_7046.mask = 4'b1000;

	lut_sub lut_7051 ({i_8_, g627}, g622);
	defparam lut_7051.LUT_SIZE = 2;
	defparam lut_7051.mask = 4'b0100;

	lut_sub lut_7056 ({i_8_, g628}, g623);
	defparam lut_7056.LUT_SIZE = 2;
	defparam lut_7056.mask = 4'b0001;

	lut_sub lut_7062 ({g625, g626}, g624);
	defparam lut_7062.LUT_SIZE = 2;
	defparam lut_7062.mask = 4'b1000;

	lut_sub lut_7067 ({i_8_, g629}, g625);
	defparam lut_7067.LUT_SIZE = 2;
	defparam lut_7067.mask = 4'b0100;

	lut_sub lut_7072 ({i_8_, g630}, g626);
	defparam lut_7072.LUT_SIZE = 2;
	defparam lut_7072.mask = 4'b0001;

	lut_sub lut_7077 ({i_6_, g46}, g627);
	defparam lut_7077.LUT_SIZE = 2;
	defparam lut_7077.mask = 4'b1110;

	lut_sub lut_7085 ({g77, i_6_, i_7_, g1}, g628);
	defparam lut_7085.LUT_SIZE = 4;
	defparam lut_7085.mask = 16'hf737;

	lut_sub lut_7101 ({i_6_, g46}, g629);
	defparam lut_7101.LUT_SIZE = 2;
	defparam lut_7101.mask = 4'b1110;

	lut_sub lut_7108 ({g77, i_6_, i_7_}, g630);
	defparam lut_7108.LUT_SIZE = 3;
	defparam lut_7108.mask = 8'hf7;

	lut_sub lut_7120 ({g632, g633}, g631);
	defparam lut_7120.LUT_SIZE = 2;
	defparam lut_7120.mask = 4'b1000;

	lut_sub lut_7126 ({g35, g634}, g632);
	defparam lut_7126.LUT_SIZE = 2;
	defparam lut_7126.mask = 4'b0100;

	lut_sub lut_7132 ({g35, g637}, g633);
	defparam lut_7132.LUT_SIZE = 2;
	defparam lut_7132.mask = 4'b0001;

	lut_sub lut_7138 ({g635, g636}, g634);
	defparam lut_7138.LUT_SIZE = 2;
	defparam lut_7138.mask = 4'b1000;

	lut_sub lut_7143 ({i_5_, g640}, g635);
	defparam lut_7143.LUT_SIZE = 2;
	defparam lut_7143.mask = 4'b0100;

	lut_sub lut_7148 ({i_5_, g641}, g636);
	defparam lut_7148.LUT_SIZE = 2;
	defparam lut_7148.mask = 4'b0001;

	lut_sub lut_7154 ({g638, g639}, g637);
	defparam lut_7154.LUT_SIZE = 2;
	defparam lut_7154.mask = 4'b1000;

	lut_sub lut_7159 ({i_5_, g642}, g638);
	defparam lut_7159.LUT_SIZE = 2;
	defparam lut_7159.mask = 4'b0100;

	lut_sub lut_7164 ({i_5_, g643}, g639);
	defparam lut_7164.LUT_SIZE = 2;
	defparam lut_7164.mask = 4'b0001;

	lut_sub lut_7169 ({i_4_, g121}, g640);
	defparam lut_7169.LUT_SIZE = 2;
	defparam lut_7169.mask = 4'b1110;

	lut_sub lut_7176 ({g95, i_4_, i_6_}, g641);
	defparam lut_7176.LUT_SIZE = 3;
	defparam lut_7176.mask = 8'hfd;

	lut_sub lut_7187 ({i_4_, g121}, g642);
	defparam lut_7187.LUT_SIZE = 2;
	defparam lut_7187.mask = 4'b1110;

	lut_sub lut_7195 ({g95, i_4_, i_6_, g42}, g643);
	defparam lut_7195.LUT_SIZE = 4;
	defparam lut_7195.mask = 16'hafa3;

	lut_sub lut_7210 ({g645, g646}, g644);
	defparam lut_7210.LUT_SIZE = 2;
	defparam lut_7210.mask = 4'b1000;

	lut_sub lut_7216 ({g42, g647}, g645);
	defparam lut_7216.LUT_SIZE = 2;
	defparam lut_7216.mask = 4'b0100;

	lut_sub lut_7222 ({g42, g650}, g646);
	defparam lut_7222.LUT_SIZE = 2;
	defparam lut_7222.mask = 4'b0001;

	lut_sub lut_7228 ({g648, g649}, g647);
	defparam lut_7228.LUT_SIZE = 2;
	defparam lut_7228.mask = 4'b1000;

	lut_sub lut_7233 ({i_6_, g653}, g648);
	defparam lut_7233.LUT_SIZE = 2;
	defparam lut_7233.mask = 4'b0100;

	lut_sub lut_7238 ({i_6_, g654}, g649);
	defparam lut_7238.LUT_SIZE = 2;
	defparam lut_7238.mask = 4'b0001;

	lut_sub lut_7244 ({g651, g652}, g650);
	defparam lut_7244.LUT_SIZE = 2;
	defparam lut_7244.mask = 4'b1000;

	lut_sub lut_7249 ({i_6_, g655}, g651);
	defparam lut_7249.LUT_SIZE = 2;
	defparam lut_7249.mask = 4'b0100;

	lut_sub lut_7254 ({i_6_, g656}, g652);
	defparam lut_7254.LUT_SIZE = 2;
	defparam lut_7254.mask = 4'b0001;

	lut_sub lut_7260 ({g24, i_8_, g36, i_7_}, g653);
	defparam lut_7260.LUT_SIZE = 4;
	defparam lut_7260.mask = 16'h7fff;

	lut_sub lut_7280 ({g24, i_8_, g45, i_7_}, g654);
	defparam lut_7280.LUT_SIZE = 4;
	defparam lut_7280.mask = 16'hf7ff;

	lut_sub lut_7300 ({g24, i_8_, g36, i_7_}, g655);
	defparam lut_7300.LUT_SIZE = 4;
	defparam lut_7300.mask = 16'h7fff;

	lut_sub lut_7320 ({g24, i_8_, g45, i_7_}, g656);
	defparam lut_7320.LUT_SIZE = 4;
	defparam lut_7320.mask = 16'h777f;

	lut_sub lut_7338 ({g658, g659}, g657);
	defparam lut_7338.LUT_SIZE = 2;
	defparam lut_7338.mask = 4'b1000;

	lut_sub lut_7344 ({g23, g660}, g658);
	defparam lut_7344.LUT_SIZE = 2;
	defparam lut_7344.mask = 4'b0100;

	lut_sub lut_7350 ({g23, g663}, g659);
	defparam lut_7350.LUT_SIZE = 2;
	defparam lut_7350.mask = 4'b0001;

	lut_sub lut_7356 ({g661, g662}, g660);
	defparam lut_7356.LUT_SIZE = 2;
	defparam lut_7356.mask = 4'b1000;

	lut_sub lut_7361 ({i_2_, g666}, g661);
	defparam lut_7361.LUT_SIZE = 2;
	defparam lut_7361.mask = 4'b0100;

	lut_sub lut_7366 ({i_2_, g667}, g662);
	defparam lut_7366.LUT_SIZE = 2;
	defparam lut_7366.mask = 4'b0001;

	lut_sub lut_7372 ({g664, g665}, g663);
	defparam lut_7372.LUT_SIZE = 2;
	defparam lut_7372.mask = 4'b1000;

	lut_sub lut_7377 ({i_2_, g668}, g664);
	defparam lut_7377.LUT_SIZE = 2;
	defparam lut_7377.mask = 4'b0100;

	lut_sub lut_7382 ({i_2_, g669}, g665);
	defparam lut_7382.LUT_SIZE = 2;
	defparam lut_7382.mask = 4'b0001;

	lut_sub lut_7388 ({i_0_, g187, i_1_, g38}, g666);
	defparam lut_7388.LUT_SIZE = 4;
	defparam lut_7388.mask = 16'hff37;

	lut_sub lut_7405 ({i_0_, i_7_, g38}, g667);
	defparam lut_7405.LUT_SIZE = 3;
	defparam lut_7405.mask = 8'hfd;

	lut_sub lut_7416 ({i_0_, g187, i_1_}, g668);
	defparam lut_7416.LUT_SIZE = 3;
	defparam lut_7416.mask = 8'hf7;

	lut_sub lut_7427 ({i_0_, i_7_, g38}, g669);
	defparam lut_7427.LUT_SIZE = 3;
	defparam lut_7427.mask = 8'hfd;

	lut_sub lut_7439 ({g671, g672}, g670);
	defparam lut_7439.LUT_SIZE = 2;
	defparam lut_7439.mask = 4'b1000;

	lut_sub lut_7445 ({g41, g673}, g671);
	defparam lut_7445.LUT_SIZE = 2;
	defparam lut_7445.mask = 4'b0100;

	lut_sub lut_7451 ({g41, g676}, g672);
	defparam lut_7451.LUT_SIZE = 2;
	defparam lut_7451.mask = 4'b0001;

	lut_sub lut_7457 ({g674, g675}, g673);
	defparam lut_7457.LUT_SIZE = 2;
	defparam lut_7457.mask = 4'b1000;

	lut_sub lut_7462 ({i_4_, g679}, g674);
	defparam lut_7462.LUT_SIZE = 2;
	defparam lut_7462.mask = 4'b0100;

	lut_sub lut_7467 ({i_4_, g680}, g675);
	defparam lut_7467.LUT_SIZE = 2;
	defparam lut_7467.mask = 4'b0001;

	lut_sub lut_7473 ({g677, g678}, g676);
	defparam lut_7473.LUT_SIZE = 2;
	defparam lut_7473.mask = 4'b1000;

	lut_sub lut_7478 ({i_4_, g681}, g677);
	defparam lut_7478.LUT_SIZE = 2;
	defparam lut_7478.mask = 4'b0100;

	lut_sub lut_7483 ({i_4_, g682}, g678);
	defparam lut_7483.LUT_SIZE = 2;
	defparam lut_7483.mask = 4'b0001;

	lut_sub lut_7489 ({g1, i_5_, g12, i_3_}, g679);
	defparam lut_7489.LUT_SIZE = 4;
	defparam lut_7489.mask = 16'hefff;

	lut_sub lut_7509 ({g1, i_5_, g28, i_3_}, g680);
	defparam lut_7509.LUT_SIZE = 4;
	defparam lut_7509.mask = 16'hefff;

	lut_sub lut_7529 ({g1, i_5_, g12, i_3_}, g681);
	defparam lut_7529.LUT_SIZE = 4;
	defparam lut_7529.mask = 16'h4f5f;

	lut_sub lut_7545 ({g1, i_5_, g28, i_3_}, g682);
	defparam lut_7545.LUT_SIZE = 4;
	defparam lut_7545.mask = 16'hefff;

	lut_sub lut_7565 ({g684, g685}, g683);
	defparam lut_7565.LUT_SIZE = 2;
	defparam lut_7565.mask = 4'b1000;

	lut_sub lut_7571 ({g27, g686}, g684);
	defparam lut_7571.LUT_SIZE = 2;
	defparam lut_7571.mask = 4'b0100;

	lut_sub lut_7577 ({g27, g689}, g685);
	defparam lut_7577.LUT_SIZE = 2;
	defparam lut_7577.mask = 4'b0001;

	lut_sub lut_7583 ({g687, g688}, g686);
	defparam lut_7583.LUT_SIZE = 2;
	defparam lut_7583.mask = 4'b1000;

	lut_sub lut_7588 ({i_8_, g691}, g687);
	defparam lut_7588.LUT_SIZE = 2;
	defparam lut_7588.mask = 4'b0100;

	lut_sub lut_7593 ({i_8_, g692}, g688);
	defparam lut_7593.LUT_SIZE = 2;
	defparam lut_7593.mask = 4'b0001;

	lut_sub lut_7598 ({i_8_, g690}, g689);
	defparam lut_7598.LUT_SIZE = 2;
	defparam lut_7598.mask = 4'b1000;

	lut_sub lut_7603 ({i_8_, g693}, g690);
	defparam lut_7603.LUT_SIZE = 2;
	defparam lut_7603.mask = 4'b0100;

	lut_sub lut_7609 ({g116, i_7_, g126, i_6_}, g691);
	defparam lut_7609.LUT_SIZE = 4;
	defparam lut_7609.mask = 16'hbf1f;

	lut_sub lut_7626 ({g116, i_7_, g5, i_6_}, g692);
	defparam lut_7626.LUT_SIZE = 4;
	defparam lut_7626.mask = 16'hfe5e;

	lut_sub lut_7642 ({i_7_, g126, i_6_}, g693);
	defparam lut_7642.LUT_SIZE = 3;
	defparam lut_7642.mask = 8'hbf;

	lut_sub lut_7654 ({g695, g696}, g694);
	defparam lut_7654.LUT_SIZE = 2;
	defparam lut_7654.mask = 4'b1000;

	lut_sub lut_7660 ({g47, g697}, g695);
	defparam lut_7660.LUT_SIZE = 2;
	defparam lut_7660.mask = 4'b0100;

	lut_sub lut_7666 ({g47, g699}, g696);
	defparam lut_7666.LUT_SIZE = 2;
	defparam lut_7666.mask = 4'b0001;

	lut_sub lut_7671 ({i_4_, g698}, g697);
	defparam lut_7671.LUT_SIZE = 2;
	defparam lut_7671.mask = 4'b1000;

	lut_sub lut_7676 ({i_4_, g702}, g698);
	defparam lut_7676.LUT_SIZE = 2;
	defparam lut_7676.mask = 4'b0100;

	lut_sub lut_7682 ({g700, g701}, g699);
	defparam lut_7682.LUT_SIZE = 2;
	defparam lut_7682.mask = 4'b1000;

	lut_sub lut_7687 ({i_4_, g703}, g700);
	defparam lut_7687.LUT_SIZE = 2;
	defparam lut_7687.mask = 4'b0100;

	lut_sub lut_7692 ({i_4_, g704}, g701);
	defparam lut_7692.LUT_SIZE = 2;
	defparam lut_7692.mask = 4'b0001;

	lut_sub lut_7697 ({i_5_, g121, i_3_}, g702);
	defparam lut_7697.LUT_SIZE = 3;
	defparam lut_7697.mask = 8'hfd;

	lut_sub lut_7708 ({i_5_, g121, i_3_}, g703);
	defparam lut_7708.LUT_SIZE = 3;
	defparam lut_7708.mask = 8'hfd;

	lut_sub lut_7719 ({i_6_, i_5_, g27, i_3_}, g704);
	defparam lut_7719.LUT_SIZE = 4;
	defparam lut_7719.mask = 16'hbffb;

	lut_sub lut_7734 ({}, gnd);
	defparam lut_7734.LUT_SIZE = 0;
	defparam lut_7734.mask = 1'b0;


endmodule