module apex4x5_map (i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_, o_1_, o_2_, o_12_, o_11_, o_14_, o_13_, o_16_, o_15_, o_18_, o_17_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

	input i_7_;
	input i_8_;
	input i_5_;
	input i_6_;
	input i_3_;
	input i_4_;
	input i_1_;
	input i_2_;
	input i_0_;
	output o_1_;
	output o_2_;
	output o_12_;
	output o_11_;
	output o_14_;
	output o_13_;
	output o_16_;
	output o_15_;
	output o_18_;
	output o_17_;
	output o_10_;
	output o_9_;
	output o_7_;
	output o_8_;
	output o_5_;
	output o_6_;
	output o_3_;
	output o_4_;



	wire x4869x, x4838x, x4839x, x4865x, x4991x, x4992x, x5048x, x5010x, x5011x, x5029x, x5030x, n_n722, n_n724, x5108x, x6347x, x5168x, x5139x, x5140x, x5164x, x5165x, x5221x;
	wire x5218x, x5219x, x5232x, x178x, x258x, x310x, x5230x, x5250x, x188x, x114x, x5246x, x5265x, x5260x, x5261x, x5270x, x187x, x259x, x294x, x261x, x5373x, x5315x;
	wire x5316x, x5369x, x5370x, x5490x, x5485x, x5486x, x5488x, n_n444, n_n450, x5586x, x5587x, x5588x, x5685x, n_n517, x5654x, x5655x, x5656x, x5781x, x5732x, n_n305, x5731x;
	wire x5877x, n_n377, x5818x, x5819x, x5820x, x5942x, x5937x, x5938x, x6028x, x6029x, x4855x, x4856x, x4861x, x4862x, x4864x, n_n78, x42x, n_n1120, x355x, n_n1156, n_n86;
	wire n_n1021, x4837x, n_n80, x337x, x1589x, x4848x, x4860x, x4928x, x4929x, x232x, x4984x, x4987x, n_n131, x4919x, x4920x, x4985x, x4986x, x5038x, x5039x, x5040x, x5041x;
	wire x5046x, n_n73, x21x, x256x, x299x, x5006x, x190x, x265x, x5003x, x5004x, x5005x, x135x, n_n949, x97x, x204x, x5025x, x195x, x151x, x5021x, x5023x, x5024x;
	wire x5060x, x5061x, x5062x, x5063x, x5064x, x5076x, x5077x, x5078x, x5079x, n_n1324, n_n1092, x5087x, x5099x, x5104x, x257x, x5093x, x5100x, x5101x, x5103x, n_n846, x5154x;
	wire x5155x, x5156x, x5157x, n_n38, x52x, x306x, x1480x, x5135x, x141x, x279x, x5131x, x5133x, x5134x, x64x, n_n82, x342x, x5148x, x5159x, x123x, x183x, x5150x;
	wire x5151x, x5152x, x5185x, x5186x, x5202x, x5203x, x1413x, x1414x, x5208x, x5214x, x1285x, x186x, x5217x, x6355x, n_n1369, n_n1176, x76x, x43x, n_n91, n_n92, n_n74;
	wire n_n90, n_n1297, n_n1283, n_n1312, x326x, n_n93, n_n1074, n_n1294, x136x, x230x, x5242x, x5248x, n_n101, x325x, n_n1047, n_n94, n_n1042, n_n1281, n_n1279, x5259x, x5262x;
	wire n_n1169, n_n942, n_n1057, n_n1125, n_n1128, n_n1286, n_n63, x49x, x248x, x341x, n_n95, x36x, x31x, x54x, n_n1132, x131x, x5012x, x39x, n_n941, x5331x, x5332x;
	wire x5333x, x5334x, x5371x, x5273x, x5274x, x5306x, x5307x, x5298x, x5309x, x5310x, x6345x, n_n1082, x1487x, x90x, x298x, x5364x, n_n958, x5358x, x5359x, x6344x, x6351x;
	wire x5388x, x5389x, x5403x, x5404x, x5484x, x5450x, x335x, x1440x, x5446x, x5482x, x5454x, x263x, x91x, x5478x, x5479x, x5421x, x5422x, x5440x, x5441x, x5539x, x5513x;
	wire x5508x, x5509x, x5538x, x5550x, x5551x, x5552x, x5553x, x5554x, x5571x, x5580x, x5573x, x5574x, x5575x, x5576x, x168x, x5568x, x5579x, x6358x, n_n514, x5676x, x5677x;
	wire x5680x, x5682x, x5616x, x5617x, x5618x, x5619x, x5620x, x94x, x223x, x101x, x5648x, x5641x, x5642x, x5643x, x5644x, x125x, x5645x, x5646x, x6340x, n_n308, x5773x;
	wire x5774x, x5776x, x5778x, n_n1160, x617x, x5717x, x5726x, x5729x, x5699x, x5700x, x5703x, x5704x, x5706x, x160x, x166x, x281x, x121x, x5727x, n_n376, x5869x, x5870x;
	wire x5872x, x5874x, x5791x, x5792x, x5793x, x6333x, x215x, x153x, x103x, n_n959, x5814x, n_n944, n_n939, x5399x, x5808x, x6357x, x303x, n_n652, x5809x, x5810x, x5812x;
	wire x5896x, x5897x, x5934x, x5935x, x5936x, x5901x, n_n984, x5899x, x5933x, x5904x, x5907x, x5908x, n_n952, x5953x, x5954x, x5955x, x5956x, x6026x, x5987x, x5985x, x5986x;
	wire x6024x, x6025x, x57x, x113x, x132x, x27x, x208x, x34x, n_n83, n_n102, x4852x, n_n58, x26x, x87x, x104x, n_n1185, x227x, x4858x, x111x, x41x, x4927x;
	wire n_n67, x1479x, x4971x, x4972x, x4973x, x4974x, x4943x, x4950x, x4951x, n_n1215, x4899x, x4891x, x4892x, x4898x, x292x, n_n882, x4910x, x4913x, x4914x, x4917x, x4975x;
	wire x4976x, x4982x, n_n137, x4936x, x231x, x4935x, x32x, n_n77, x346x, x343x, x255x, x48x, n_n1204, x25x, x53x, x5035x, x61x, x301x, x5037x, x296x, x5121x;
	wire x5123x, x5124x, x206x, x72x, n_n1193, n_n1330, n_n1267, x5176x, x5181x, x254x, x88x, x5178x, x5179x, x5180x, x5193x, x5198x, x5196x, x5197x, x5200x, x351x, x37x;
	wire x333x, x278x, n_n1259, n_n1032, x5244x, x189x, n_n1046, x75x, n_n1028, n_n1018, n_n1040, n_n1011, x59x, x1085x, x201x, x164x, x288x, x203x, n_n999, n_n1009, x156x;
	wire x5321x, x5322x, x5360x, x5362x, n_n980, n_n983, n_n986, x5384x, n_n1001, n_n1004, x5383x, x5386x, n_n953, x5393x, x5400x, x282x, x285x, x5472x, x5474x, x5475x, x119x;
	wire x5524x, x5532x, x5536x, x102x, x5504x, x5505x, x5507x, x5493x, n_n1130, n_n1164, x246x, x1082x, x262x, n_n1163, x220x, x5526x, x5528x, x5529x, x5599x, x5600x, x5601x;
	wire x5602x, x5603x, x66x, n_n71, x5668x, x224x, x1384x, x670x, x67x, x5664x, x6342x, n_n211, x120x, x139x, x5672x, x5673x, x5743x, x5744x, x5746x, x6339x, n_n1091;
	wire n_n982, x268x, x5751x, x5753x, n_n84, x6338x, x6350x, x162x, x266x, x5763x, x6337x, x5769x, x5770x, x5841x, x5842x, x5844x, x6334x, x158x, x159x, x5848x, x340x;
	wire x5850x, x5852x, x5853x, x5858x, x5859x, x5860x, x5826x, x5827x, x5854x, x5855x, x5866x, x138x, x5886x, x5892x, n_n1014, x152x, x5889x, x5895x, x5927x, x92x, x155x;
	wire x307x, x5919x, x226x, x267x, x5921x, x5922x, x5924x, n_n1079, x753x, x5609x, x287x, n_n1030, x98x, x154x, n_n1087, x280x, x5944x, x5946x, x5990x, x5991x, x6018x;
	wire x350x, x5964x, x5975x, x5984x, x23x, x5910x, x5514x, x6360x, x225x, x5971x, x5972x, x5974x, x6009x, x6010x, x6011x, x6012x, x6013x, x6014x, x6015x, x6016x, n_n75;
	wire n_n81, n_n64, n_n52, x175x, n_n100, x108x, x128x, n_n85, n_n70, n_n54, n_n1134, n_n103, n_n97, x45x, x55x, x58x, n_n1217, x112x, x56x, x318x, x63x;
	wire x172x, x235x, x252x, x311x, x329x, n_n1036, x107x, x110x, x4887x, x249x, x4888x, x22x, x324x, x327x, x4889x, n_n1052, x70x, x237x, n_n1013, x4885x, x6348x;
	wire n_n76, x146x, n_n973, n_n975, x29x, x1557x, n_n943, n_n976, n_n1006, n_n978, n_n967, x202x, n_n1172, n_n1078, x245x, x38x, x239x, x30x, x339x, x118x, x6352x;
	wire x354x, x62x, x4934x, n_n1153, x44x, n_n87, x4938x, x304x, n_n1103, x319x, x4944x, n_n1105, n_n1108, n_n1100, x19x, x105x, x109x, x127x, x207x, x1483x, x1484x;
	wire x35x, x251x, x321x, x328x, n_n1085, n_n1095, x20x, n_n1088, n_n1181, n_n1146, n_n1022, x322x, n_n1060, x28x, n_n951, x79x, n_n969, n_n1188, x1518x, x1519x, x46x;
	wire x5031x, n_n1039, x78x, n_n1216, n_n1170, x5056x, x5059x, n_n954, x147x, n_n1010, n_n981, x272x, n_n1093, n_n1331, n_n40, x1359x, n_n66, x353x, x117x, n_n1058, x133x;
	wire x148x, x173x, x177x, x323x, x1352x, x233x, x5083x, x1348x, x5085x, x271x, n_n966, x145x, x270x, x5114x, x83x, n_n1177, n_n1158, x65x, x1291x, x1292x, x348x;
	wire x194x, n_n1184, x274x, x185x, x352x, n_n1109, n_n937, x217x, x290x, x6349x, x1143x, x5283x, x6346x, x332x, x5288x, x5289x, x5290x, x71x, x5291x, x5292x, x5305x;
	wire x234x, x320x, n_n989, n_n1121, n_n53, x1588x, x330x, n_n962, x5338x, x236x, n_n1118, x275x, x238x, x313x, n_n987, n_n994, x163x, x200x, x1017x, x5392x, n_n1045;
	wire n_n1043, x1153x, x5407x, x309x, x289x, x5417x, x5413x, x210x, x5414x, x5415x, x5411x, x5416x, x33x, x5429x, x5436x, x5432x, x122x, x5433x, x5434x, x5435x, x5442x;
	wire n_n1101, x6359x, n_n1059, x334x, x142x, x944x, x150x, x85x, x331x, x5068x, n_n971, n_n1037, x903x, x5492x, x242x, x877x, x835x, x5519x, x5531x, n_n947, x829x;
	wire x212x, n_n1026, x68x, x805x, x1008x, x5595x, x869x, x6353x, x5715x, x6336x, n_n1002, n_n296, x129x, x161x, x218x, x526x, x5835x, x6335x, x247x, x316x, x344x;
	wire x827x, x5880x, x5881x, x5882x, x615x, x6361x, x157x, x174x, x662x, x663x, x336x, x130x, x5686x, x5687x, x5965x, x5966x, x5967x, x5968x, x312x, x345x, x1583x;
	wire x4876x, x1581x, x900x, x5499x, x876x, x5697x, x5693x, x5694x, x5695x, x1508x, x5828x, x1108x, x1442x, x1446x, x4849x, x4961x, x4967x, x4968x, x4969x, x4970x, x5205x;
	wire x5206x, x6356x, x5293x, x5342x, x5351x, x5460x, x5467x, x5468x, x6343x, x5518x, x5522x, x6341x, x5758x, x5798x, x5856x, x5914x, x5915x, x5918x, x5926x, x5969x, x5996x;
	wire x6006x;

	assign o_1_ = (((x4869x) & (!x4838x) & (!x4839x) & (!x4865x)) + ((!x4869x) & (x4838x) & (!x4839x) & (!x4865x)) + ((!x4869x) & (!x4838x) & (x4839x) & (!x4865x)) + ((!x4869x) & (!x4838x) & (!x4839x) & (x4865x)));
	assign o_2_ = (((x4991x) & (!x4992x)) + ((!x4991x) & (x4992x)));
	assign o_12_ = (((x5048x) & (!x5010x) & (!x5011x) & (!x5029x) & (!x5030x)) + ((!x5048x) & (x5010x) & (!x5011x) & (!x5029x) & (!x5030x)) + ((!x5048x) & (!x5010x) & (x5011x) & (!x5029x) & (!x5030x)) + ((!x5048x) & (!x5010x) & (!x5011x) & (x5029x) & (!x5030x)) + ((!x5048x) & (!x5010x) & (!x5011x) & (!x5029x) & (x5030x)));
	assign o_11_ = (((n_n722) & (!n_n724) & (!x5108x) & (!x6347x)) + ((!n_n722) & (n_n724) & (!x5108x) & (!x6347x)) + ((!n_n722) & (!n_n724) & (x5108x) & (!x6347x)) + ((!n_n722) & (!n_n724) & (!x5108x) & (!x6347x)));
	assign o_14_ = (((x5168x) & (!x5139x) & (!x5140x) & (!x5164x) & (!x5165x)) + ((!x5168x) & (x5139x) & (!x5140x) & (!x5164x) & (!x5165x)) + ((!x5168x) & (!x5139x) & (x5140x) & (!x5164x) & (!x5165x)) + ((!x5168x) & (!x5139x) & (!x5140x) & (x5164x) & (!x5165x)) + ((!x5168x) & (!x5139x) & (!x5140x) & (!x5164x) & (x5165x)));
	assign o_13_ = (((x5221x) & (!x5218x) & (!x5219x)) + ((!x5221x) & (x5218x) & (!x5219x)) + ((!x5221x) & (!x5218x) & (x5219x)));
	assign o_16_ = (((x5232x) & (!x178x) & (!x258x) & (!x310x) & (!x5230x)) + ((!x5232x) & (x178x) & (!x258x) & (!x310x) & (!x5230x)) + ((!x5232x) & (!x178x) & (x258x) & (!x310x) & (!x5230x)) + ((!x5232x) & (!x178x) & (!x258x) & (x310x) & (!x5230x)) + ((!x5232x) & (!x178x) & (!x258x) & (!x310x) & (x5230x)));
	assign o_15_ = (((x5250x) & (!x310x) & (!x188x) & (!x114x) & (!x5246x)) + ((!x5250x) & (x310x) & (!x188x) & (!x114x) & (!x5246x)) + ((!x5250x) & (!x310x) & (x188x) & (!x114x) & (!x5246x)) + ((!x5250x) & (!x310x) & (!x188x) & (x114x) & (!x5246x)) + ((!x5250x) & (!x310x) & (!x188x) & (!x114x) & (x5246x)));
	assign o_18_ = (((x5265x) & (!x5260x) & (!x5261x)) + ((!x5265x) & (x5260x) & (!x5261x)) + ((!x5265x) & (!x5260x) & (x5261x)));
	assign o_17_ = (((x5270x) & (!x187x) & (!x259x) & (!x294x) & (!x261x)) + ((!x5270x) & (x187x) & (!x259x) & (!x294x) & (!x261x)) + ((!x5270x) & (!x187x) & (x259x) & (!x294x) & (!x261x)) + ((!x5270x) & (!x187x) & (!x259x) & (x294x) & (!x261x)) + ((!x5270x) & (!x187x) & (!x259x) & (!x294x) & (x261x)));
	assign o_10_ = (((x5373x) & (!x5315x) & (!x5316x) & (!x5369x) & (!x5370x)) + ((!x5373x) & (x5315x) & (!x5316x) & (!x5369x) & (!x5370x)) + ((!x5373x) & (!x5315x) & (x5316x) & (!x5369x) & (!x5370x)) + ((!x5373x) & (!x5315x) & (!x5316x) & (x5369x) & (!x5370x)) + ((!x5373x) & (!x5315x) & (!x5316x) & (!x5369x) & (x5370x)));
	assign o_9_ = (((x5490x) & (!x5485x) & (!x5486x) & (!x5488x)) + ((!x5490x) & (x5485x) & (!x5486x) & (!x5488x)) + ((!x5490x) & (!x5485x) & (x5486x) & (!x5488x)) + ((!x5490x) & (!x5485x) & (!x5486x) & (x5488x)));
	assign o_7_ = (((n_n444) & (!n_n450) & (!x5586x) & (!x5587x) & (!x5588x)) + ((!n_n444) & (n_n450) & (!x5586x) & (!x5587x) & (!x5588x)) + ((!n_n444) & (!n_n450) & (x5586x) & (!x5587x) & (!x5588x)) + ((!n_n444) & (!n_n450) & (!x5586x) & (x5587x) & (!x5588x)) + ((!n_n444) & (!n_n450) & (!x5586x) & (!x5587x) & (x5588x)));
	assign o_8_ = (((x5685x) & (!n_n517) & (!x5654x) & (!x5655x) & (!x5656x)) + ((!x5685x) & (n_n517) & (!x5654x) & (!x5655x) & (!x5656x)) + ((!x5685x) & (!n_n517) & (x5654x) & (!x5655x) & (!x5656x)) + ((!x5685x) & (!n_n517) & (!x5654x) & (x5655x) & (!x5656x)) + ((!x5685x) & (!n_n517) & (!x5654x) & (!x5655x) & (x5656x)));
	assign o_5_ = (((x5781x) & (!x5732x) & (!n_n305) & (!x5731x)) + ((!x5781x) & (x5732x) & (!n_n305) & (!x5731x)) + ((!x5781x) & (!x5732x) & (n_n305) & (!x5731x)) + ((!x5781x) & (!x5732x) & (!n_n305) & (x5731x)));
	assign o_6_ = (((x5877x) & (!n_n377) & (!x5818x) & (!x5819x) & (!x5820x)) + ((!x5877x) & (n_n377) & (!x5818x) & (!x5819x) & (!x5820x)) + ((!x5877x) & (!n_n377) & (x5818x) & (!x5819x) & (!x5820x)) + ((!x5877x) & (!n_n377) & (!x5818x) & (x5819x) & (!x5820x)) + ((!x5877x) & (!n_n377) & (!x5818x) & (!x5819x) & (x5820x)));
	assign o_3_ = (((x5942x) & (!x5937x) & (!x5938x)) + ((!x5942x) & (x5937x) & (!x5938x)) + ((!x5942x) & (!x5937x) & (x5938x)));
	assign o_4_ = (((x6028x) & (!x6029x)) + ((!x6028x) & (x6029x)));
	assign x4869x = (((x4855x) & (!x4856x) & (!x4861x) & (!x4862x) & (!x4864x)) + ((!x4855x) & (x4856x) & (!x4861x) & (!x4862x) & (!x4864x)) + ((!x4855x) & (!x4856x) & (x4861x) & (!x4862x) & (!x4864x)) + ((!x4855x) & (!x4856x) & (!x4861x) & (x4862x) & (!x4864x)) + ((!x4855x) & (!x4856x) & (!x4861x) & (!x4862x) & (x4864x)));
	assign x4838x = (((!n_n78) & (!x42x) & (n_n1120) & (!x355x) & (!n_n1156)) + ((!n_n78) & (!x42x) & (!n_n1120) & (x355x) & (!n_n1156)) + ((!n_n78) & (!x42x) & (!n_n1120) & (!x355x) & (n_n1156)) + ((n_n78) & (x42x) & (!n_n1120) & (!x355x) & (!n_n1156)));
	assign x4839x = (((!i_6_) & (!n_n86) & (!x42x) & (n_n1021) & (!x4837x)) + ((!i_6_) & (!n_n86) & (!x42x) & (!n_n1021) & (x4837x)) + ((i_6_) & (n_n86) & (x42x) & (!n_n1021) & (!x4837x)));
	assign x4865x = (((!n_n80) & (!x337x) & (x1589x) & (!x4848x) & (!x4860x)) + ((!n_n80) & (!x337x) & (!x1589x) & (x4848x) & (!x4860x)) + ((!n_n80) & (!x337x) & (!x1589x) & (!x4848x) & (x4860x)) + ((n_n80) & (x337x) & (!x1589x) & (!x4848x) & (!x4860x)));
	assign x4991x = (((x4928x) & (!x4929x) & (!x232x) & (!x4984x) & (!x4987x)) + ((!x4928x) & (x4929x) & (!x232x) & (!x4984x) & (!x4987x)) + ((!x4928x) & (!x4929x) & (x232x) & (!x4984x) & (!x4987x)) + ((!x4928x) & (!x4929x) & (!x232x) & (x4984x) & (!x4987x)) + ((!x4928x) & (!x4929x) & (!x232x) & (!x4984x) & (x4987x)));
	assign x4992x = (((n_n131) & (!x4919x) & (!x4920x) & (!x4985x) & (!x4986x)) + ((!n_n131) & (x4919x) & (!x4920x) & (!x4985x) & (!x4986x)) + ((!n_n131) & (!x4919x) & (x4920x) & (!x4985x) & (!x4986x)) + ((!n_n131) & (!x4919x) & (!x4920x) & (x4985x) & (!x4986x)) + ((!n_n131) & (!x4919x) & (!x4920x) & (!x4985x) & (x4986x)));
	assign x5048x = (((x5038x) & (!x5039x) & (!x5040x) & (!x5041x) & (!x5046x)) + ((!x5038x) & (x5039x) & (!x5040x) & (!x5041x) & (!x5046x)) + ((!x5038x) & (!x5039x) & (x5040x) & (!x5041x) & (!x5046x)) + ((!x5038x) & (!x5039x) & (!x5040x) & (x5041x) & (!x5046x)) + ((!x5038x) & (!x5039x) & (!x5040x) & (!x5041x) & (x5046x)));
	assign x5010x = (((!n_n73) & (!x21x) & (x256x) & (!x299x) & (!x5006x)) + ((!n_n73) & (!x21x) & (!x256x) & (x299x) & (!x5006x)) + ((!n_n73) & (!x21x) & (!x256x) & (!x299x) & (x5006x)) + ((n_n73) & (x21x) & (!x256x) & (!x299x) & (!x5006x)));
	assign x5011x = (((x190x) & (!x265x) & (!x5003x) & (!x5004x) & (!x5005x)) + ((!x190x) & (x265x) & (!x5003x) & (!x5004x) & (!x5005x)) + ((!x190x) & (!x265x) & (x5003x) & (!x5004x) & (!x5005x)) + ((!x190x) & (!x265x) & (!x5003x) & (x5004x) & (!x5005x)) + ((!x190x) & (!x265x) & (!x5003x) & (!x5004x) & (x5005x)));
	assign x5029x = (((x135x) & (!n_n949) & (!x97x) & (!x204x) & (!x5025x)) + ((!x135x) & (n_n949) & (!x97x) & (!x204x) & (!x5025x)) + ((!x135x) & (!n_n949) & (x97x) & (!x204x) & (!x5025x)) + ((!x135x) & (!n_n949) & (!x97x) & (x204x) & (!x5025x)) + ((!x135x) & (!n_n949) & (!x97x) & (!x204x) & (x5025x)));
	assign x5030x = (((x195x) & (!x151x) & (!x5021x) & (!x5023x) & (!x5024x)) + ((!x195x) & (x151x) & (!x5021x) & (!x5023x) & (!x5024x)) + ((!x195x) & (!x151x) & (x5021x) & (!x5023x) & (!x5024x)) + ((!x195x) & (!x151x) & (!x5021x) & (x5023x) & (!x5024x)) + ((!x195x) & (!x151x) & (!x5021x) & (!x5023x) & (x5024x)));
	assign n_n722 = (((x5060x) & (!x5061x) & (!x5062x) & (!x5063x) & (!x5064x)) + ((!x5060x) & (x5061x) & (!x5062x) & (!x5063x) & (!x5064x)) + ((!x5060x) & (!x5061x) & (x5062x) & (!x5063x) & (!x5064x)) + ((!x5060x) & (!x5061x) & (!x5062x) & (x5063x) & (!x5064x)) + ((!x5060x) & (!x5061x) & (!x5062x) & (!x5063x) & (x5064x)));
	assign n_n724 = (((x5076x) & (!x5077x) & (!x5078x) & (!x5079x)) + ((!x5076x) & (x5077x) & (!x5078x) & (!x5079x)) + ((!x5076x) & (!x5077x) & (x5078x) & (!x5079x)) + ((!x5076x) & (!x5077x) & (!x5078x) & (x5079x)));
	assign x5108x = (((n_n1324) & (!n_n1092) & (!x5087x) & (!x5099x) & (!x5104x)) + ((!n_n1324) & (n_n1092) & (!x5087x) & (!x5099x) & (!x5104x)) + ((!n_n1324) & (!n_n1092) & (x5087x) & (!x5099x) & (!x5104x)) + ((!n_n1324) & (!n_n1092) & (!x5087x) & (x5099x) & (!x5104x)) + ((!n_n1324) & (!n_n1092) & (!x5087x) & (!x5099x) & (x5104x)));
	assign x6347x = (((!x257x) & (!x5093x) & (!x5100x) & (!x5101x) & (!x5103x)));
	assign x5168x = (((n_n846) & (!x5154x) & (!x5155x) & (!x5156x) & (!x5157x)) + ((!n_n846) & (x5154x) & (!x5155x) & (!x5156x) & (!x5157x)) + ((!n_n846) & (!x5154x) & (x5155x) & (!x5156x) & (!x5157x)) + ((!n_n846) & (!x5154x) & (!x5155x) & (x5156x) & (!x5157x)) + ((!n_n846) & (!x5154x) & (!x5155x) & (!x5156x) & (x5157x)));
	assign x5139x = (((!n_n38) & (!x52x) & (x306x) & (!x1480x) & (!x5135x)) + ((!n_n38) & (!x52x) & (!x306x) & (x1480x) & (!x5135x)) + ((!n_n38) & (!x52x) & (!x306x) & (!x1480x) & (x5135x)) + ((n_n38) & (x52x) & (!x306x) & (!x1480x) & (!x5135x)));
	assign x5140x = (((x141x) & (!x279x) & (!x5131x) & (!x5133x) & (!x5134x)) + ((!x141x) & (x279x) & (!x5131x) & (!x5133x) & (!x5134x)) + ((!x141x) & (!x279x) & (x5131x) & (!x5133x) & (!x5134x)) + ((!x141x) & (!x279x) & (!x5131x) & (x5133x) & (!x5134x)) + ((!x141x) & (!x279x) & (!x5131x) & (!x5133x) & (x5134x)));
	assign x5164x = (((!x64x) & (!n_n82) & (x342x) & (!x5148x) & (!x5159x)) + ((!x64x) & (!n_n82) & (!x342x) & (x5148x) & (!x5159x)) + ((!x64x) & (!n_n82) & (!x342x) & (!x5148x) & (x5159x)) + ((x64x) & (n_n82) & (!x342x) & (!x5148x) & (!x5159x)));
	assign x5165x = (((x123x) & (!x183x) & (!x5150x) & (!x5151x) & (!x5152x)) + ((!x123x) & (x183x) & (!x5150x) & (!x5151x) & (!x5152x)) + ((!x123x) & (!x183x) & (x5150x) & (!x5151x) & (!x5152x)) + ((!x123x) & (!x183x) & (!x5150x) & (x5151x) & (!x5152x)) + ((!x123x) & (!x183x) & (!x5150x) & (!x5151x) & (x5152x)));
	assign x5221x = (((x5185x) & (!x5186x) & (!x5202x) & (!x5203x)) + ((!x5185x) & (x5186x) & (!x5202x) & (!x5203x)) + ((!x5185x) & (!x5186x) & (x5202x) & (!x5203x)) + ((!x5185x) & (!x5186x) & (!x5202x) & (x5203x)));
	assign x5218x = (((x178x) & (!x1413x) & (!x1414x) & (!x5208x) & (!x5214x)) + ((!x178x) & (x1413x) & (!x1414x) & (!x5208x) & (!x5214x)) + ((!x178x) & (!x1413x) & (x1414x) & (!x5208x) & (!x5214x)) + ((!x178x) & (!x1413x) & (!x1414x) & (x5208x) & (!x5214x)) + ((!x178x) & (!x1413x) & (!x1414x) & (!x5208x) & (x5214x)));
	assign x5219x = (((x1285x) & (!x186x) & (!x5217x) & (!x6355x)) + ((!x1285x) & (x186x) & (!x5217x) & (!x6355x)) + ((!x1285x) & (!x186x) & (x5217x) & (!x6355x)) + ((!x1285x) & (!x186x) & (!x5217x) & (!x6355x)));
	assign x5232x = (((n_n1369) & (!n_n1176) & (!x187x) & (!x259x) & (!x294x)) + ((!n_n1369) & (n_n1176) & (!x187x) & (!x259x) & (!x294x)) + ((!n_n1369) & (!n_n1176) & (x187x) & (!x259x) & (!x294x)) + ((!n_n1369) & (!n_n1176) & (!x187x) & (x259x) & (!x294x)) + ((!n_n1369) & (!n_n1176) & (!x187x) & (!x259x) & (x294x)));
	assign x178x = (((!i_7_) & (i_8_) & (i_6_) & (x76x) & (!x43x)) + ((!i_7_) & (!i_8_) & (!i_6_) & (!x76x) & (x43x)));
	assign x258x = (((n_n78) & (!n_n91) & (n_n92) & (!n_n74) & (n_n90)) + ((!n_n78) & (n_n91) & (!n_n92) & (n_n74) & (n_n90)));
	assign x310x = (((n_n1297) & (!n_n1283) & (!n_n1312) & (!x326x)) + ((!n_n1297) & (n_n1283) & (!n_n1312) & (!x326x)) + ((!n_n1297) & (!n_n1283) & (n_n1312) & (!x326x)) + ((!n_n1297) & (!n_n1283) & (!n_n1312) & (x326x)));
	assign x5230x = (((!n_n38) & (!n_n93) & (!x43x) & (n_n1074) & (!n_n1294)) + ((!n_n38) & (!n_n93) & (!x43x) & (!n_n1074) & (n_n1294)) + ((n_n38) & (!n_n93) & (x43x) & (!n_n1074) & (!n_n1294)) + ((!n_n38) & (n_n93) & (x43x) & (!n_n1074) & (!n_n1294)));
	assign x5250x = (((x136x) & (!x230x) & (!x5242x) & (!x5248x)) + ((!x136x) & (x230x) & (!x5242x) & (!x5248x)) + ((!x136x) & (!x230x) & (x5242x) & (!x5248x)) + ((!x136x) & (!x230x) & (!x5242x) & (x5248x)));
	assign x188x = (((!i_3_) & (!n_n101) & (!x325x) & (!n_n90) & (n_n1047)) + ((i_3_) & (n_n101) & (x325x) & (n_n90) & (!n_n1047)));
	assign x114x = (((!i_3_) & (!n_n78) & (!n_n94) & (!x325x) & (n_n1042)) + ((i_3_) & (n_n78) & (n_n94) & (x325x) & (!n_n1042)));
	assign x5246x = (((n_n1281) & (!n_n1279) & (!x258x) & (!x259x) & (!x294x)) + ((!n_n1281) & (n_n1279) & (!x258x) & (!x259x) & (!x294x)) + ((!n_n1281) & (!n_n1279) & (x258x) & (!x259x) & (!x294x)) + ((!n_n1281) & (!n_n1279) & (!x258x) & (x259x) & (!x294x)) + ((!n_n1281) & (!n_n1279) & (!x258x) & (!x259x) & (x294x)));
	assign x5265x = (((x230x) & (!x261x) & (!x5259x) & (!x5262x)) + ((!x230x) & (x261x) & (!x5259x) & (!x5262x)) + ((!x230x) & (!x261x) & (x5259x) & (!x5262x)) + ((!x230x) & (!x261x) & (!x5259x) & (x5262x)));
	assign x5260x = (((n_n1294) & (!n_n1169) & (!n_n942) & (!n_n1057)) + ((!n_n1294) & (n_n1169) & (!n_n942) & (!n_n1057)) + ((!n_n1294) & (!n_n1169) & (n_n942) & (!n_n1057)) + ((!n_n1294) & (!n_n1169) & (!n_n942) & (n_n1057)));
	assign x5261x = (((!n_n101) & (!x43x) & (n_n1125) & (!n_n1128) & (!n_n1286)) + ((!n_n101) & (!x43x) & (!n_n1125) & (n_n1128) & (!n_n1286)) + ((!n_n101) & (!x43x) & (!n_n1125) & (!n_n1128) & (n_n1286)) + ((n_n101) & (x43x) & (!n_n1125) & (!n_n1128) & (!n_n1286)));
	assign x5270x = (((!n_n63) & (!x49x) & (n_n1176) & (!x248x) & (!n_n1283)) + ((!n_n63) & (!x49x) & (!n_n1176) & (x248x) & (!n_n1283)) + ((!n_n63) & (!x49x) & (!n_n1176) & (!x248x) & (n_n1283)) + ((n_n63) & (x49x) & (!n_n1176) & (!x248x) & (!n_n1283)));
	assign x187x = (((!i_3_) & (!x341x) & (n_n95) & (x36x) & (!x31x)) + ((i_3_) & (x341x) & (!n_n95) & (!x36x) & (x31x)));
	assign x259x = (((!i_5_) & (!n_n101) & (!x54x) & (!n_n90) & (n_n1132)) + ((!i_5_) & (n_n101) & (x54x) & (n_n90) & (!n_n1132)));
	assign x294x = (((!i_1_) & (!i_2_) & (!i_0_) & (!x131x) & (!x5012x)) + ((!i_1_) & (!i_2_) & (!i_0_) & (x131x) & (!x5012x)) + ((!i_1_) & (!i_2_) & (!i_0_) & (!x131x) & (x5012x)));
	assign x261x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x39x) & (n_n941)) + ((i_7_) & (i_8_) & (!i_6_) & (x39x) & (!n_n941)));
	assign x5373x = (((x5331x) & (!x5332x) & (!x5333x) & (!x5334x) & (!x5371x)) + ((!x5331x) & (x5332x) & (!x5333x) & (!x5334x) & (!x5371x)) + ((!x5331x) & (!x5332x) & (x5333x) & (!x5334x) & (!x5371x)) + ((!x5331x) & (!x5332x) & (!x5333x) & (x5334x) & (!x5371x)) + ((!x5331x) & (!x5332x) & (!x5333x) & (!x5334x) & (x5371x)));
	assign x5315x = (((x5273x) & (!x5274x) & (!x5306x) & (!x5307x)) + ((!x5273x) & (x5274x) & (!x5306x) & (!x5307x)) + ((!x5273x) & (!x5274x) & (x5306x) & (!x5307x)) + ((!x5273x) & (!x5274x) & (!x5306x) & (x5307x)));
	assign x5316x = (((x5298x) & (!x5309x) & (!x5310x) & (!x6345x)) + ((!x5298x) & (x5309x) & (!x5310x) & (!x6345x)) + ((!x5298x) & (!x5309x) & (x5310x) & (!x6345x)) + ((!x5298x) & (!x5309x) & (!x5310x) & (!x6345x)));
	assign x5369x = (((n_n1082) & (!x1487x) & (!x90x) & (!x298x) & (!x5364x)) + ((!n_n1082) & (x1487x) & (!x90x) & (!x298x) & (!x5364x)) + ((!n_n1082) & (!x1487x) & (x90x) & (!x298x) & (!x5364x)) + ((!n_n1082) & (!x1487x) & (!x90x) & (x298x) & (!x5364x)) + ((!n_n1082) & (!x1487x) & (!x90x) & (!x298x) & (x5364x)));
	assign x5370x = (((n_n958) & (!x5358x) & (!x5359x) & (!x6344x) & (!x6351x)) + ((!n_n958) & (x5358x) & (!x5359x) & (!x6344x) & (!x6351x)) + ((!n_n958) & (!x5358x) & (x5359x) & (!x6344x) & (!x6351x)) + ((!n_n958) & (!x5358x) & (!x5359x) & (!x6344x) & (!x6351x)) + ((!n_n958) & (!x5358x) & (!x5359x) & (!x6344x) & (!x6351x)));
	assign x5490x = (((x5388x) & (!x5389x) & (!x5403x) & (!x5404x) & (!x5484x)) + ((!x5388x) & (x5389x) & (!x5403x) & (!x5404x) & (!x5484x)) + ((!x5388x) & (!x5389x) & (x5403x) & (!x5404x) & (!x5484x)) + ((!x5388x) & (!x5389x) & (!x5403x) & (x5404x) & (!x5484x)) + ((!x5388x) & (!x5389x) & (!x5403x) & (!x5404x) & (x5484x)));
	assign x5485x = (((x5450x) & (!x335x) & (!x1440x) & (!x5446x) & (!x5482x)) + ((!x5450x) & (x335x) & (!x1440x) & (!x5446x) & (!x5482x)) + ((!x5450x) & (!x335x) & (x1440x) & (!x5446x) & (!x5482x)) + ((!x5450x) & (!x335x) & (!x1440x) & (x5446x) & (!x5482x)) + ((!x5450x) & (!x335x) & (!x1440x) & (!x5446x) & (x5482x)));
	assign x5486x = (((x5454x) & (!x263x) & (!x91x) & (!x5478x) & (!x5479x)) + ((!x5454x) & (x263x) & (!x91x) & (!x5478x) & (!x5479x)) + ((!x5454x) & (!x263x) & (x91x) & (!x5478x) & (!x5479x)) + ((!x5454x) & (!x263x) & (!x91x) & (x5478x) & (!x5479x)) + ((!x5454x) & (!x263x) & (!x91x) & (!x5478x) & (x5479x)));
	assign x5488x = (((x5421x) & (!x5422x) & (!x5440x) & (!x5441x)) + ((!x5421x) & (x5422x) & (!x5440x) & (!x5441x)) + ((!x5421x) & (!x5422x) & (x5440x) & (!x5441x)) + ((!x5421x) & (!x5422x) & (!x5440x) & (x5441x)));
	assign n_n444 = (((x5539x) & (!x5513x) & (!x5508x) & (!x5509x) & (!x5538x)) + ((!x5539x) & (x5513x) & (!x5508x) & (!x5509x) & (!x5538x)) + ((!x5539x) & (!x5513x) & (x5508x) & (!x5509x) & (!x5538x)) + ((!x5539x) & (!x5513x) & (!x5508x) & (x5509x) & (!x5538x)) + ((!x5539x) & (!x5513x) & (!x5508x) & (!x5509x) & (x5538x)));
	assign n_n450 = (((x5550x) & (!x5551x) & (!x5552x) & (!x5553x) & (!x5554x)) + ((!x5550x) & (x5551x) & (!x5552x) & (!x5553x) & (!x5554x)) + ((!x5550x) & (!x5551x) & (x5552x) & (!x5553x) & (!x5554x)) + ((!x5550x) & (!x5551x) & (!x5552x) & (x5553x) & (!x5554x)) + ((!x5550x) & (!x5551x) & (!x5552x) & (!x5553x) & (x5554x)));
	assign x5586x = (((x204x) & (!x263x) & (!x5571x) & (!x5580x)) + ((!x204x) & (x263x) & (!x5571x) & (!x5580x)) + ((!x204x) & (!x263x) & (x5571x) & (!x5580x)) + ((!x204x) & (!x263x) & (!x5571x) & (x5580x)));
	assign x5587x = (((x5573x) & (!x5574x) & (!x5575x) & (!x5576x)) + ((!x5573x) & (x5574x) & (!x5575x) & (!x5576x)) + ((!x5573x) & (!x5574x) & (x5575x) & (!x5576x)) + ((!x5573x) & (!x5574x) & (!x5575x) & (x5576x)));
	assign x5588x = (((x168x) & (!x5568x) & (!x5579x) & (!x6358x)) + ((!x168x) & (x5568x) & (!x5579x) & (!x6358x)) + ((!x168x) & (!x5568x) & (x5579x) & (!x6358x)) + ((!x168x) & (!x5568x) & (!x5579x) & (!x6358x)));
	assign x5685x = (((n_n514) & (!x5676x) & (!x5677x) & (!x5680x) & (!x5682x)) + ((!n_n514) & (x5676x) & (!x5677x) & (!x5680x) & (!x5682x)) + ((!n_n514) & (!x5676x) & (x5677x) & (!x5680x) & (!x5682x)) + ((!n_n514) & (!x5676x) & (!x5677x) & (x5680x) & (!x5682x)) + ((!n_n514) & (!x5676x) & (!x5677x) & (!x5680x) & (x5682x)));
	assign n_n517 = (((x5616x) & (!x5617x) & (!x5618x) & (!x5619x) & (!x5620x)) + ((!x5616x) & (x5617x) & (!x5618x) & (!x5619x) & (!x5620x)) + ((!x5616x) & (!x5617x) & (x5618x) & (!x5619x) & (!x5620x)) + ((!x5616x) & (!x5617x) & (!x5618x) & (x5619x) & (!x5620x)) + ((!x5616x) & (!x5617x) & (!x5618x) & (!x5619x) & (x5620x)));
	assign x5654x = (((x94x) & (!x195x) & (!x223x) & (!x101x) & (!x5648x)) + ((!x94x) & (x195x) & (!x223x) & (!x101x) & (!x5648x)) + ((!x94x) & (!x195x) & (x223x) & (!x101x) & (!x5648x)) + ((!x94x) & (!x195x) & (!x223x) & (x101x) & (!x5648x)) + ((!x94x) & (!x195x) & (!x223x) & (!x101x) & (x5648x)));
	assign x5655x = (((x5641x) & (!x5642x) & (!x5643x) & (!x5644x)) + ((!x5641x) & (x5642x) & (!x5643x) & (!x5644x)) + ((!x5641x) & (!x5642x) & (x5643x) & (!x5644x)) + ((!x5641x) & (!x5642x) & (!x5643x) & (x5644x)));
	assign x5656x = (((x97x) & (!x125x) & (!x5645x) & (!x5646x) & (!x6340x)) + ((!x97x) & (x125x) & (!x5645x) & (!x5646x) & (!x6340x)) + ((!x97x) & (!x125x) & (x5645x) & (!x5646x) & (!x6340x)) + ((!x97x) & (!x125x) & (!x5645x) & (x5646x) & (!x6340x)) + ((!x97x) & (!x125x) & (!x5645x) & (!x5646x) & (!x6340x)));
	assign x5781x = (((n_n308) & (!x5773x) & (!x5774x) & (!x5776x) & (!x5778x)) + ((!n_n308) & (x5773x) & (!x5774x) & (!x5776x) & (!x5778x)) + ((!n_n308) & (!x5773x) & (x5774x) & (!x5776x) & (!x5778x)) + ((!n_n308) & (!x5773x) & (!x5774x) & (x5776x) & (!x5778x)) + ((!n_n308) & (!x5773x) & (!x5774x) & (!x5776x) & (x5778x)));
	assign x5732x = (((n_n1160) & (!x617x) & (!x5717x) & (!x5726x) & (!x5729x)) + ((!n_n1160) & (x617x) & (!x5717x) & (!x5726x) & (!x5729x)) + ((!n_n1160) & (!x617x) & (x5717x) & (!x5726x) & (!x5729x)) + ((!n_n1160) & (!x617x) & (!x5717x) & (x5726x) & (!x5729x)) + ((!n_n1160) & (!x617x) & (!x5717x) & (!x5726x) & (x5729x)));
	assign n_n305 = (((x5699x) & (!x5700x) & (!x5703x) & (!x5704x) & (!x5706x)) + ((!x5699x) & (x5700x) & (!x5703x) & (!x5704x) & (!x5706x)) + ((!x5699x) & (!x5700x) & (x5703x) & (!x5704x) & (!x5706x)) + ((!x5699x) & (!x5700x) & (!x5703x) & (x5704x) & (!x5706x)) + ((!x5699x) & (!x5700x) & (!x5703x) & (!x5704x) & (x5706x)));
	assign x5731x = (((x160x) & (!x166x) & (!x281x) & (!x121x) & (!x5727x)) + ((!x160x) & (x166x) & (!x281x) & (!x121x) & (!x5727x)) + ((!x160x) & (!x166x) & (x281x) & (!x121x) & (!x5727x)) + ((!x160x) & (!x166x) & (!x281x) & (x121x) & (!x5727x)) + ((!x160x) & (!x166x) & (!x281x) & (!x121x) & (x5727x)));
	assign x5877x = (((n_n376) & (!x5869x) & (!x5870x) & (!x5872x) & (!x5874x)) + ((!n_n376) & (x5869x) & (!x5870x) & (!x5872x) & (!x5874x)) + ((!n_n376) & (!x5869x) & (x5870x) & (!x5872x) & (!x5874x)) + ((!n_n376) & (!x5869x) & (!x5870x) & (x5872x) & (!x5874x)) + ((!n_n376) & (!x5869x) & (!x5870x) & (!x5872x) & (x5874x)));
	assign n_n377 = (((x5791x) & (!x5792x) & (!x5793x) & (!x6333x)) + ((!x5791x) & (x5792x) & (!x5793x) & (!x6333x)) + ((!x5791x) & (!x5792x) & (x5793x) & (!x6333x)) + ((!x5791x) & (!x5792x) & (!x5793x) & (!x6333x)));
	assign x5818x = (((x215x) & (!x153x) & (!x103x) & (!n_n959) & (!x5814x)) + ((!x215x) & (x153x) & (!x103x) & (!n_n959) & (!x5814x)) + ((!x215x) & (!x153x) & (x103x) & (!n_n959) & (!x5814x)) + ((!x215x) & (!x153x) & (!x103x) & (n_n959) & (!x5814x)) + ((!x215x) & (!x153x) & (!x103x) & (!n_n959) & (x5814x)));
	assign x5819x = (((n_n944) & (!n_n939) & (!x5399x) & (!x5808x) & (!x6357x)) + ((!n_n944) & (n_n939) & (!x5399x) & (!x5808x) & (!x6357x)) + ((!n_n944) & (!n_n939) & (x5399x) & (!x5808x) & (!x6357x)) + ((!n_n944) & (!n_n939) & (!x5399x) & (x5808x) & (!x6357x)) + ((!n_n944) & (!n_n939) & (!x5399x) & (!x5808x) & (!x6357x)));
	assign x5820x = (((x303x) & (!n_n652) & (!x5809x) & (!x5810x) & (!x5812x)) + ((!x303x) & (n_n652) & (!x5809x) & (!x5810x) & (!x5812x)) + ((!x303x) & (!n_n652) & (x5809x) & (!x5810x) & (!x5812x)) + ((!x303x) & (!n_n652) & (!x5809x) & (x5810x) & (!x5812x)) + ((!x303x) & (!n_n652) & (!x5809x) & (!x5810x) & (x5812x)));
	assign x5942x = (((x5896x) & (!x5897x) & (!x5934x) & (!x5935x) & (!x5936x)) + ((!x5896x) & (x5897x) & (!x5934x) & (!x5935x) & (!x5936x)) + ((!x5896x) & (!x5897x) & (x5934x) & (!x5935x) & (!x5936x)) + ((!x5896x) & (!x5897x) & (!x5934x) & (x5935x) & (!x5936x)) + ((!x5896x) & (!x5897x) & (!x5934x) & (!x5935x) & (x5936x)));
	assign x5937x = (((x103x) & (!x5901x) & (!n_n984) & (!x5899x) & (!x5933x)) + ((!x103x) & (x5901x) & (!n_n984) & (!x5899x) & (!x5933x)) + ((!x103x) & (!x5901x) & (n_n984) & (!x5899x) & (!x5933x)) + ((!x103x) & (!x5901x) & (!n_n984) & (x5899x) & (!x5933x)) + ((!x103x) & (!x5901x) & (!n_n984) & (!x5899x) & (x5933x)));
	assign x5938x = (((x153x) & (!x5904x) & (!x5907x) & (!x5908x) & (!n_n952)) + ((!x153x) & (x5904x) & (!x5907x) & (!x5908x) & (!n_n952)) + ((!x153x) & (!x5904x) & (x5907x) & (!x5908x) & (!n_n952)) + ((!x153x) & (!x5904x) & (!x5907x) & (x5908x) & (!n_n952)) + ((!x153x) & (!x5904x) & (!x5907x) & (!x5908x) & (n_n952)));
	assign x6028x = (((x5953x) & (!x5954x) & (!x5955x) & (!x5956x) & (!x6026x)) + ((!x5953x) & (x5954x) & (!x5955x) & (!x5956x) & (!x6026x)) + ((!x5953x) & (!x5954x) & (x5955x) & (!x5956x) & (!x6026x)) + ((!x5953x) & (!x5954x) & (!x5955x) & (x5956x) & (!x6026x)) + ((!x5953x) & (!x5954x) & (!x5955x) & (!x5956x) & (x6026x)));
	assign x6029x = (((x5987x) & (!x5985x) & (!x5986x) & (!x6024x) & (!x6025x)) + ((!x5987x) & (x5985x) & (!x5986x) & (!x6024x) & (!x6025x)) + ((!x5987x) & (!x5985x) & (x5986x) & (!x6024x) & (!x6025x)) + ((!x5987x) & (!x5985x) & (!x5986x) & (x6024x) & (!x6025x)) + ((!x5987x) & (!x5985x) & (!x5986x) & (!x6024x) & (x6025x)));
	assign x4855x = (((!x57x) & (!n_n92) & (x113x) & (!n_n95) & (!x132x)) + ((x57x) & (!n_n92) & (!x113x) & (n_n95) & (!x132x)) + ((!x57x) & (n_n92) & (!x113x) & (!n_n95) & (x132x)));
	assign x4856x = (((!x27x) & (!n_n63) & (x208x) & (!n_n95) & (!x34x)) + ((x27x) & (!n_n63) & (!x208x) & (n_n95) & (!x34x)) + ((!x27x) & (n_n63) & (!x208x) & (!n_n95) & (x34x)));
	assign x4861x = (((!n_n101) & (!n_n91) & (!n_n83) & (!n_n102) & (x4852x)) + ((n_n101) & (!n_n91) & (n_n83) & (n_n102) & (!x4852x)) + ((!n_n101) & (n_n91) & (n_n83) & (n_n102) & (!x4852x)));
	assign x4862x = (((!n_n58) & (!x26x) & (!x39x) & (x87x) & (!x104x)) + ((!n_n58) & (!x26x) & (!x39x) & (!x87x) & (x104x)) + ((n_n58) & (x26x) & (!x39x) & (!x87x) & (!x104x)) + ((n_n58) & (!x26x) & (x39x) & (!x87x) & (!x104x)));
	assign x4864x = (((!n_n91) & (!x76x) & (n_n1185) & (!x227x) & (!x4858x)) + ((!n_n91) & (!x76x) & (!n_n1185) & (x227x) & (!x4858x)) + ((!n_n91) & (!x76x) & (!n_n1185) & (!x227x) & (x4858x)) + ((n_n91) & (x76x) & (!n_n1185) & (!x227x) & (!x4858x)));
	assign x4928x = (((!n_n91) & (!x49x) & (!x111x) & (!x41x) & (x136x)) + ((n_n91) & (x49x) & (!x111x) & (!x41x) & (!x136x)) + ((!n_n91) & (!x49x) & (x111x) & (x41x) & (!x136x)));
	assign x4929x = (((!x27x) & (!x26x) & (!n_n63) & (!n_n82) & (x4927x)) + ((x27x) & (!x26x) & (n_n63) & (!n_n82) & (!x4927x)) + ((!x27x) & (x26x) & (!n_n63) & (n_n82) & (!x4927x)));
	assign x232x = (((!i_4_) & (!n_n93) & (!n_n67) & (x1479x) & (!x1480x)) + ((!i_4_) & (!n_n93) & (!n_n67) & (!x1479x) & (x1480x)) + ((!i_4_) & (n_n93) & (n_n67) & (!x1479x) & (!x1480x)));
	assign x4984x = (((x4971x) & (!x4972x) & (!x4973x) & (!x4974x)) + ((!x4971x) & (x4972x) & (!x4973x) & (!x4974x)) + ((!x4971x) & (!x4972x) & (x4973x) & (!x4974x)) + ((!x4971x) & (!x4972x) & (!x4973x) & (x4974x)));
	assign x4987x = (((x4943x) & (!x4950x) & (!x4951x) & (!n_n1215) & (!x121x)) + ((!x4943x) & (x4950x) & (!x4951x) & (!n_n1215) & (!x121x)) + ((!x4943x) & (!x4950x) & (x4951x) & (!n_n1215) & (!x121x)) + ((!x4943x) & (!x4950x) & (!x4951x) & (n_n1215) & (!x121x)) + ((!x4943x) & (!x4950x) & (!x4951x) & (!n_n1215) & (x121x)));
	assign n_n131 = (((x4899x) & (!x4891x) & (!x4892x) & (!x4898x)) + ((!x4899x) & (x4891x) & (!x4892x) & (!x4898x)) + ((!x4899x) & (!x4891x) & (x4892x) & (!x4898x)) + ((!x4899x) & (!x4891x) & (!x4892x) & (x4898x)));
	assign x4919x = (((x298x) & (!x292x) & (!n_n882) & (!x4910x)) + ((!x298x) & (x292x) & (!n_n882) & (!x4910x)) + ((!x298x) & (!x292x) & (n_n882) & (!x4910x)) + ((!x298x) & (!x292x) & (!n_n882) & (x4910x)));
	assign x4920x = (((x4913x) & (!x4914x) & (!x4917x)) + ((!x4913x) & (x4914x) & (!x4917x)) + ((!x4913x) & (!x4914x) & (x4917x)));
	assign x4985x = (((x4975x) & (!x4976x) & (!x4982x)) + ((!x4975x) & (x4976x) & (!x4982x)) + ((!x4975x) & (!x4976x) & (x4982x)));
	assign x4986x = (((n_n137) & (!x4936x) & (!x231x) & (!x4935x)) + ((!n_n137) & (x4936x) & (!x231x) & (!x4935x)) + ((!n_n137) & (!x4936x) & (x231x) & (!x4935x)) + ((!n_n137) & (!x4936x) & (!x231x) & (x4935x)));
	assign x5038x = (((!x32x) & (!n_n77) & (x346x) & (!x1413x) & (!x1414x)) + ((!x32x) & (!n_n77) & (!x346x) & (x1413x) & (!x1414x)) + ((!x32x) & (!n_n77) & (!x346x) & (!x1413x) & (x1414x)) + ((x32x) & (n_n77) & (!x346x) & (!x1413x) & (!x1414x)));
	assign x5039x = (((!i_5_) & (!x54x) & (x343x) & (!x255x) & (!x48x)) + ((!i_5_) & (!x54x) & (!x343x) & (x255x) & (!x48x)) + ((i_5_) & (x54x) & (!x343x) & (!x255x) & (x48x)));
	assign x5040x = (((!n_n78) & (!n_n63) & (!x49x) & (n_n1204) & (!n_n1369)) + ((!n_n78) & (!n_n63) & (!x49x) & (!n_n1204) & (n_n1369)) + ((n_n78) & (!n_n63) & (x49x) & (!n_n1204) & (!n_n1369)) + ((!n_n78) & (n_n63) & (x49x) & (!n_n1204) & (!n_n1369)));
	assign x5041x = (((!n_n58) & (!n_n78) & (!x25x) & (!x53x) & (x5035x)) + ((n_n58) & (!n_n78) & (x25x) & (!x53x) & (!x5035x)) + ((!n_n58) & (n_n78) & (!x25x) & (x53x) & (!x5035x)));
	assign x5046x = (((x87x) & (!x61x) & (!x231x) & (!x301x) & (!x5037x)) + ((!x87x) & (x61x) & (!x231x) & (!x301x) & (!x5037x)) + ((!x87x) & (!x61x) & (x231x) & (!x301x) & (!x5037x)) + ((!x87x) & (!x61x) & (!x231x) & (x301x) & (!x5037x)) + ((!x87x) & (!x61x) & (!x231x) & (!x301x) & (x5037x)));
	assign n_n846 = (((n_n882) & (!x296x) & (!x5121x) & (!x5123x) & (!x5124x)) + ((!n_n882) & (x296x) & (!x5121x) & (!x5123x) & (!x5124x)) + ((!n_n882) & (!x296x) & (x5121x) & (!x5123x) & (!x5124x)) + ((!n_n882) & (!x296x) & (!x5121x) & (x5123x) & (!x5124x)) + ((!n_n882) & (!x296x) & (!x5121x) & (!x5123x) & (x5124x)));
	assign x5154x = (((!i_5_) & (!x54x) & (x1285x) & (!x186x) & (!x31x)) + ((!i_5_) & (!x54x) & (!x1285x) & (x186x) & (!x31x)) + ((i_5_) & (x54x) & (!x1285x) & (!x186x) & (x31x)));
	assign x5155x = (((!i_7_) & (!i_6_) & (!x34x) & (x206x) & (!n_n1215)) + ((!i_7_) & (!i_6_) & (!x34x) & (!x206x) & (n_n1215)) + ((i_7_) & (i_6_) & (x34x) & (!x206x) & (!n_n1215)));
	assign x5156x = (((!i_1_) & (!n_n86) & (n_n1324) & (!n_n1369) & (!x72x)) + ((!i_1_) & (!n_n86) & (!n_n1324) & (n_n1369) & (!x72x)) + ((!i_1_) & (n_n86) & (!n_n1324) & (!n_n1369) & (x72x)));
	assign x5157x = (((!n_n63) & (!x49x) & (n_n1193) & (!n_n1330) & (!n_n1267)) + ((!n_n63) & (!x49x) & (!n_n1193) & (n_n1330) & (!n_n1267)) + ((!n_n63) & (!x49x) & (!n_n1193) & (!n_n1330) & (n_n1267)) + ((n_n63) & (x49x) & (!n_n1193) & (!n_n1330) & (!n_n1267)));
	assign x5185x = (((x306x) & (!x5176x) & (!x5181x)) + ((!x306x) & (x5176x) & (!x5181x)) + ((!x306x) & (!x5176x) & (x5181x)));
	assign x5186x = (((x254x) & (!x88x) & (!x5178x) & (!x5179x) & (!x5180x)) + ((!x254x) & (x88x) & (!x5178x) & (!x5179x) & (!x5180x)) + ((!x254x) & (!x88x) & (x5178x) & (!x5179x) & (!x5180x)) + ((!x254x) & (!x88x) & (!x5178x) & (x5179x) & (!x5180x)) + ((!x254x) & (!x88x) & (!x5178x) & (!x5179x) & (x5180x)));
	assign x5202x = (((x125x) & (!x5193x) & (!x5198x)) + ((!x125x) & (x5193x) & (!x5198x)) + ((!x125x) & (!x5193x) & (x5198x)));
	assign x5203x = (((x5196x) & (!x5197x) & (!x5200x)) + ((!x5196x) & (x5197x) & (!x5200x)) + ((!x5196x) & (!x5197x) & (x5200x)));
	assign n_n1369 = (((!i_7_) & (i_8_) & (!i_5_) & (!i_6_) & (x351x)));
	assign n_n1176 = (((i_1_) & (!i_2_) & (!i_0_) & (n_n91) & (n_n74)));
	assign x136x = (((!i_5_) & (!i_3_) & (!i_4_) & (!x37x) & (n_n1330)) + ((i_5_) & (i_3_) & (!i_4_) & (x37x) & (!n_n1330)));
	assign x230x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x49x) & (x333x)) + ((i_7_) & (!i_8_) & (!i_6_) & (x49x) & (!x333x)));
	assign x5242x = (((!n_n93) & (!n_n102) & (n_n1369) & (!n_n90) & (!x278x)) + ((!n_n93) & (!n_n102) & (!n_n1369) & (!n_n90) & (x278x)) + ((n_n93) & (n_n102) & (!n_n1369) & (n_n90) & (!x278x)));
	assign x5248x = (((n_n1259) & (!n_n1032) & (!n_n1169) & (!n_n942) & (!x5244x)) + ((!n_n1259) & (n_n1032) & (!n_n1169) & (!n_n942) & (!x5244x)) + ((!n_n1259) & (!n_n1032) & (n_n1169) & (!n_n942) & (!x5244x)) + ((!n_n1259) & (!n_n1032) & (!n_n1169) & (n_n942) & (!x5244x)) + ((!n_n1259) & (!n_n1032) & (!n_n1169) & (!n_n942) & (x5244x)));
	assign x5259x = (((!i_1_) & (!n_n86) & (n_n1324) & (!x72x) & (!n_n1074)) + ((!i_1_) & (!n_n86) & (!n_n1324) & (!x72x) & (n_n1074)) + ((!i_1_) & (n_n86) & (!n_n1324) & (x72x) & (!n_n1074)));
	assign x5262x = (((x136x) & (!x114x) & (!x189x) & (!n_n1046) & (!n_n1047)) + ((!x136x) & (x114x) & (!x189x) & (!n_n1046) & (!n_n1047)) + ((!x136x) & (!x114x) & (x189x) & (!n_n1046) & (!n_n1047)) + ((!x136x) & (!x114x) & (!x189x) & (n_n1046) & (!n_n1047)) + ((!x136x) & (!x114x) & (!x189x) & (!n_n1046) & (n_n1047)));
	assign n_n63 = (((!i_7_) & (i_8_) & (!i_6_)));
	assign x49x = (((i_5_) & (i_3_) & (!i_4_) & (!i_0_) & (x75x)));
	assign x248x = (((i_1_) & (!i_2_) & (!i_0_) & (n_n95) & (n_n77)));
	assign n_n1283 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n91) & (n_n90)));
	assign x5331x = (((!x57x) & (!n_n63) & (n_n1047) & (!n_n1028) & (!n_n1018)) + ((!x57x) & (!n_n63) & (!n_n1047) & (n_n1028) & (!n_n1018)) + ((!x57x) & (!n_n63) & (!n_n1047) & (!n_n1028) & (n_n1018)) + ((x57x) & (n_n63) & (!n_n1047) & (!n_n1028) & (!n_n1018)));
	assign x5332x = (((n_n1032) & (!n_n1040) & (!n_n1011) & (!x59x) & (!x1085x)) + ((!n_n1032) & (n_n1040) & (!n_n1011) & (!x59x) & (!x1085x)) + ((!n_n1032) & (!n_n1040) & (n_n1011) & (!x59x) & (!x1085x)) + ((!n_n1032) & (!n_n1040) & (!n_n1011) & (x59x) & (!x1085x)) + ((!n_n1032) & (!n_n1040) & (!n_n1011) & (!x59x) & (x1085x)));
	assign x5333x = (((x201x) & (!x164x) & (!x288x) & (!x203x)) + ((!x201x) & (x164x) & (!x288x) & (!x203x)) + ((!x201x) & (!x164x) & (x288x) & (!x203x)) + ((!x201x) & (!x164x) & (!x288x) & (x203x)));
	assign x5334x = (((n_n999) & (!n_n1009) & (!x156x) & (!x5321x) & (!x5322x)) + ((!n_n999) & (n_n1009) & (!x156x) & (!x5321x) & (!x5322x)) + ((!n_n999) & (!n_n1009) & (x156x) & (!x5321x) & (!x5322x)) + ((!n_n999) & (!n_n1009) & (!x156x) & (x5321x) & (!x5322x)) + ((!n_n999) & (!n_n1009) & (!x156x) & (!x5321x) & (x5322x)));
	assign x5371x = (((x232x) & (!x257x) & (!x168x) & (!x5360x) & (!x5362x)) + ((!x232x) & (x257x) & (!x168x) & (!x5360x) & (!x5362x)) + ((!x232x) & (!x257x) & (x168x) & (!x5360x) & (!x5362x)) + ((!x232x) & (!x257x) & (!x168x) & (x5360x) & (!x5362x)) + ((!x232x) & (!x257x) & (!x168x) & (!x5360x) & (x5362x)));
	assign x5388x = (((n_n980) & (!n_n983) & (!n_n882) & (!n_n986) & (!x5384x)) + ((!n_n980) & (n_n983) & (!n_n882) & (!n_n986) & (!x5384x)) + ((!n_n980) & (!n_n983) & (n_n882) & (!n_n986) & (!x5384x)) + ((!n_n980) & (!n_n983) & (!n_n882) & (n_n986) & (!x5384x)) + ((!n_n980) & (!n_n983) & (!n_n882) & (!n_n986) & (x5384x)));
	assign x5389x = (((n_n1001) & (!n_n1004) & (!x223x) & (!x5383x) & (!x5386x)) + ((!n_n1001) & (n_n1004) & (!x223x) & (!x5383x) & (!x5386x)) + ((!n_n1001) & (!n_n1004) & (x223x) & (!x5383x) & (!x5386x)) + ((!n_n1001) & (!n_n1004) & (!x223x) & (x5383x) & (!x5386x)) + ((!n_n1001) & (!n_n1004) & (!x223x) & (!x5383x) & (x5386x)));
	assign x5403x = (((x168x) & (!n_n953) & (!n_n652) & (!x195x)) + ((!x168x) & (n_n953) & (!n_n652) & (!x195x)) + ((!x168x) & (!n_n953) & (n_n652) & (!x195x)) + ((!x168x) & (!n_n953) & (!n_n652) & (x195x)));
	assign x5404x = (((x97x) & (!x125x) & (!x303x) & (!x5393x) & (!x5400x)) + ((!x97x) & (x125x) & (!x303x) & (!x5393x) & (!x5400x)) + ((!x97x) & (!x125x) & (x303x) & (!x5393x) & (!x5400x)) + ((!x97x) & (!x125x) & (!x303x) & (x5393x) & (!x5400x)) + ((!x97x) & (!x125x) & (!x303x) & (!x5393x) & (x5400x)));
	assign x5484x = (((x282x) & (!x285x) & (!x5472x) & (!x5474x) & (!x5475x)) + ((!x282x) & (x285x) & (!x5472x) & (!x5474x) & (!x5475x)) + ((!x282x) & (!x285x) & (x5472x) & (!x5474x) & (!x5475x)) + ((!x282x) & (!x285x) & (!x5472x) & (x5474x) & (!x5475x)) + ((!x282x) & (!x285x) & (!x5472x) & (!x5474x) & (x5475x)));
	assign x5539x = (((x119x) & (!x160x) & (!x5524x) & (!x5532x) & (!x5536x)) + ((!x119x) & (x160x) & (!x5524x) & (!x5532x) & (!x5536x)) + ((!x119x) & (!x160x) & (x5524x) & (!x5532x) & (!x5536x)) + ((!x119x) & (!x160x) & (!x5524x) & (x5532x) & (!x5536x)) + ((!x119x) & (!x160x) & (!x5524x) & (!x5532x) & (x5536x)));
	assign x5513x = (((x101x) & (!x102x) & (!x5504x) & (!x5505x) & (!x5507x)) + ((!x101x) & (x102x) & (!x5504x) & (!x5505x) & (!x5507x)) + ((!x101x) & (!x102x) & (x5504x) & (!x5505x) & (!x5507x)) + ((!x101x) & (!x102x) & (!x5504x) & (x5505x) & (!x5507x)) + ((!x101x) & (!x102x) & (!x5504x) & (!x5505x) & (x5507x)));
	assign x5508x = (((!n_n94) & (!x5493x) & (n_n1130) & (!n_n1164) & (!x246x)) + ((!n_n94) & (!x5493x) & (!n_n1130) & (n_n1164) & (!x246x)) + ((!n_n94) & (!x5493x) & (!n_n1130) & (!n_n1164) & (x246x)) + ((n_n94) & (x5493x) & (!n_n1130) & (!n_n1164) & (!x246x)));
	assign x5509x = (((n_n1125) & (!x1082x) & (!x262x) & (!n_n1163) & (!x265x)) + ((!n_n1125) & (x1082x) & (!x262x) & (!n_n1163) & (!x265x)) + ((!n_n1125) & (!x1082x) & (x262x) & (!n_n1163) & (!x265x)) + ((!n_n1125) & (!x1082x) & (!x262x) & (n_n1163) & (!x265x)) + ((!n_n1125) & (!x1082x) & (!x262x) & (!n_n1163) & (x265x)));
	assign x5538x = (((x220x) & (!x281x) & (!x5526x) & (!x5528x) & (!x5529x)) + ((!x220x) & (x281x) & (!x5526x) & (!x5528x) & (!x5529x)) + ((!x220x) & (!x281x) & (x5526x) & (!x5528x) & (!x5529x)) + ((!x220x) & (!x281x) & (!x5526x) & (x5528x) & (!x5529x)) + ((!x220x) & (!x281x) & (!x5526x) & (!x5528x) & (x5529x)));
	assign n_n514 = (((x5599x) & (!x5600x) & (!x5601x) & (!x5602x) & (!x5603x)) + ((!x5599x) & (x5600x) & (!x5601x) & (!x5602x) & (!x5603x)) + ((!x5599x) & (!x5600x) & (x5601x) & (!x5602x) & (!x5603x)) + ((!x5599x) & (!x5600x) & (!x5601x) & (x5602x) & (!x5603x)) + ((!x5599x) & (!x5600x) & (!x5601x) & (!x5602x) & (x5603x)));
	assign x5676x = (((!n_n92) & (!x66x) & (!x132x) & (!n_n71) & (x5668x)) + ((n_n92) & (!x66x) & (x132x) & (!n_n71) & (!x5668x)) + ((!n_n92) & (x66x) & (!x132x) & (n_n71) & (!x5668x)));
	assign x5677x = (((!n_n58) & (!x36x) & (x224x) & (!x1384x) & (!x670x)) + ((!n_n58) & (!x36x) & (!x224x) & (x1384x) & (!x670x)) + ((!n_n58) & (!x36x) & (!x224x) & (!x1384x) & (x670x)) + ((n_n58) & (x36x) & (!x224x) & (!x1384x) & (!x670x)));
	assign x5680x = (((!n_n95) & (!x67x) & (n_n1169) & (!x5664x) & (!x6342x)) + ((!n_n95) & (!x67x) & (!n_n1169) & (x5664x) & (!x6342x)) + ((!n_n95) & (!x67x) & (!n_n1169) & (!x5664x) & (!x6342x)) + ((n_n95) & (x67x) & (!n_n1169) & (!x5664x) & (!x6342x)));
	assign x5682x = (((n_n211) & (!x120x) & (!x139x) & (!x5672x) & (!x5673x)) + ((!n_n211) & (x120x) & (!x139x) & (!x5672x) & (!x5673x)) + ((!n_n211) & (!x120x) & (x139x) & (!x5672x) & (!x5673x)) + ((!n_n211) & (!x120x) & (!x139x) & (x5672x) & (!x5673x)) + ((!n_n211) & (!x120x) & (!x139x) & (!x5672x) & (x5673x)));
	assign n_n308 = (((x5743x) & (!x5744x) & (!x5746x) & (!x6339x)) + ((!x5743x) & (x5744x) & (!x5746x) & (!x6339x)) + ((!x5743x) & (!x5744x) & (x5746x) & (!x6339x)) + ((!x5743x) & (!x5744x) & (!x5746x) & (!x6339x)));
	assign x5773x = (((n_n1091) & (!n_n982) & (!x268x) & (!x5751x) & (!x5753x)) + ((!n_n1091) & (n_n982) & (!x268x) & (!x5751x) & (!x5753x)) + ((!n_n1091) & (!n_n982) & (x268x) & (!x5751x) & (!x5753x)) + ((!n_n1091) & (!n_n982) & (!x268x) & (x5751x) & (!x5753x)) + ((!n_n1091) & (!n_n982) & (!x268x) & (!x5751x) & (x5753x)));
	assign x5774x = (((!n_n84) & (!n_n83) & (!n_n82) & (!x6338x) & (!x6350x)) + ((!n_n84) & (!n_n83) & (!n_n82) & (!x6338x) & (!x6350x)) + ((n_n84) & (n_n83) & (n_n82) & (!x6338x) & (!x6350x)));
	assign x5776x = (((x162x) & (!x266x) & (!x5763x) & (!x6337x)) + ((!x162x) & (x266x) & (!x5763x) & (!x6337x)) + ((!x162x) & (!x266x) & (x5763x) & (!x6337x)) + ((!x162x) & (!x266x) & (!x5763x) & (!x6337x)));
	assign x5778x = (((x303x) & (!x5393x) & (!x5769x) & (!x5770x)) + ((!x303x) & (x5393x) & (!x5769x) & (!x5770x)) + ((!x303x) & (!x5393x) & (x5769x) & (!x5770x)) + ((!x303x) & (!x5393x) & (!x5769x) & (x5770x)));
	assign n_n376 = (((x5841x) & (!x5842x) & (!x5844x) & (!x6334x)) + ((!x5841x) & (x5842x) & (!x5844x) & (!x6334x)) + ((!x5841x) & (!x5842x) & (x5844x) & (!x6334x)) + ((!x5841x) & (!x5842x) & (!x5844x) & (!x6334x)));
	assign x5869x = (((n_n1286) & (!n_n1283) & (!x158x) & (!x159x) & (!x5848x)) + ((!n_n1286) & (n_n1283) & (!x158x) & (!x159x) & (!x5848x)) + ((!n_n1286) & (!n_n1283) & (x158x) & (!x159x) & (!x5848x)) + ((!n_n1286) & (!n_n1283) & (!x158x) & (x159x) & (!x5848x)) + ((!n_n1286) & (!n_n1283) & (!x158x) & (!x159x) & (x5848x)));
	assign x5870x = (((x335x) & (!x340x) & (!x5850x) & (!x5852x) & (!x5853x)) + ((!x335x) & (x340x) & (!x5850x) & (!x5852x) & (!x5853x)) + ((!x335x) & (!x340x) & (x5850x) & (!x5852x) & (!x5853x)) + ((!x335x) & (!x340x) & (!x5850x) & (x5852x) & (!x5853x)) + ((!x335x) & (!x340x) & (!x5850x) & (!x5852x) & (x5853x)));
	assign x5872x = (((x301x) & (!x5858x) & (!x5859x) & (!x5860x)) + ((!x301x) & (x5858x) & (!x5859x) & (!x5860x)) + ((!x301x) & (!x5858x) & (x5859x) & (!x5860x)) + ((!x301x) & (!x5858x) & (!x5859x) & (x5860x)));
	assign x5874x = (((x5826x) & (!x5827x) & (!x5854x) & (!x5855x) & (!x5866x)) + ((!x5826x) & (x5827x) & (!x5854x) & (!x5855x) & (!x5866x)) + ((!x5826x) & (!x5827x) & (x5854x) & (!x5855x) & (!x5866x)) + ((!x5826x) & (!x5827x) & (!x5854x) & (x5855x) & (!x5866x)) + ((!x5826x) & (!x5827x) & (!x5854x) & (!x5855x) & (x5866x)));
	assign x5896x = (((x138x) & (!x268x) & (!x5886x) & (!x5892x)) + ((!x138x) & (x268x) & (!x5886x) & (!x5892x)) + ((!x138x) & (!x268x) & (x5886x) & (!x5892x)) + ((!x138x) & (!x268x) & (!x5886x) & (x5892x)));
	assign x5897x = (((n_n1014) & (!x152x) & (!n_n1018) & (!x5889x) & (!x5895x)) + ((!n_n1014) & (x152x) & (!n_n1018) & (!x5889x) & (!x5895x)) + ((!n_n1014) & (!x152x) & (n_n1018) & (!x5889x) & (!x5895x)) + ((!n_n1014) & (!x152x) & (!n_n1018) & (x5889x) & (!x5895x)) + ((!n_n1014) & (!x152x) & (!n_n1018) & (!x5889x) & (x5895x)));
	assign x5934x = (((x168x) & (!n_n211) & (!x5927x)) + ((!x168x) & (n_n211) & (!x5927x)) + ((!x168x) & (!n_n211) & (x5927x)));
	assign x5935x = (((x303x) & (!x92x) & (!x155x) & (!x307x) & (!x5919x)) + ((!x303x) & (x92x) & (!x155x) & (!x307x) & (!x5919x)) + ((!x303x) & (!x92x) & (x155x) & (!x307x) & (!x5919x)) + ((!x303x) & (!x92x) & (!x155x) & (x307x) & (!x5919x)) + ((!x303x) & (!x92x) & (!x155x) & (!x307x) & (x5919x)));
	assign x5936x = (((x226x) & (!x267x) & (!x5921x) & (!x5922x) & (!x5924x)) + ((!x226x) & (x267x) & (!x5921x) & (!x5922x) & (!x5924x)) + ((!x226x) & (!x267x) & (x5921x) & (!x5922x) & (!x5924x)) + ((!x226x) & (!x267x) & (!x5921x) & (x5922x) & (!x5924x)) + ((!x226x) & (!x267x) & (!x5921x) & (!x5922x) & (x5924x)));
	assign x5953x = (((!n_n95) & (n_n1079) & (!x34x) & (!x753x) & (!x5609x)) + ((!n_n95) & (!n_n1079) & (!x34x) & (x753x) & (!x5609x)) + ((!n_n95) & (!n_n1079) & (!x34x) & (!x753x) & (x5609x)) + ((n_n95) & (!n_n1079) & (x34x) & (!x753x) & (!x5609x)));
	assign x5954x = (((!n_n102) & (!n_n94) & (!n_n63) & (x282x) & (!x287x)) + ((!n_n102) & (!n_n94) & (!n_n63) & (!x282x) & (x287x)) + ((n_n102) & (n_n94) & (n_n63) & (!x282x) & (!x287x)));
	assign x5955x = (((n_n1030) & (!n_n1021) & (!x151x) & (!x98x) & (!x154x)) + ((!n_n1030) & (n_n1021) & (!x151x) & (!x98x) & (!x154x)) + ((!n_n1030) & (!n_n1021) & (x151x) & (!x98x) & (!x154x)) + ((!n_n1030) & (!n_n1021) & (!x151x) & (x98x) & (!x154x)) + ((!n_n1030) & (!n_n1021) & (!x151x) & (!x98x) & (x154x)));
	assign x5956x = (((n_n1057) & (!n_n1087) & (!x280x) & (!x5944x) & (!x5946x)) + ((!n_n1057) & (n_n1087) & (!x280x) & (!x5944x) & (!x5946x)) + ((!n_n1057) & (!n_n1087) & (x280x) & (!x5944x) & (!x5946x)) + ((!n_n1057) & (!n_n1087) & (!x280x) & (x5944x) & (!x5946x)) + ((!n_n1057) & (!n_n1087) & (!x280x) & (!x5944x) & (x5946x)));
	assign x6026x = (((x125x) & (!n_n652) & (!x5990x) & (!x5991x) & (!x6018x)) + ((!x125x) & (n_n652) & (!x5990x) & (!x5991x) & (!x6018x)) + ((!x125x) & (!n_n652) & (x5990x) & (!x5991x) & (!x6018x)) + ((!x125x) & (!n_n652) & (!x5990x) & (x5991x) & (!x6018x)) + ((!x125x) & (!n_n652) & (!x5990x) & (!x5991x) & (x6018x)));
	assign x5987x = (((n_n1215) & (!x350x) & (!x5964x) & (!x5975x) & (!x5984x)) + ((!n_n1215) & (x350x) & (!x5964x) & (!x5975x) & (!x5984x)) + ((!n_n1215) & (!x350x) & (x5964x) & (!x5975x) & (!x5984x)) + ((!n_n1215) & (!x350x) & (!x5964x) & (x5975x) & (!x5984x)) + ((!n_n1215) & (!x350x) & (!x5964x) & (!x5975x) & (x5984x)));
	assign x5985x = (((!n_n58) & (!x23x) & (x5910x) & (!x5514x) & (!x6360x)) + ((!n_n58) & (!x23x) & (!x5910x) & (x5514x) & (!x6360x)) + ((!n_n58) & (!x23x) & (!x5910x) & (!x5514x) & (!x6360x)) + ((n_n58) & (x23x) & (!x5910x) & (!x5514x) & (!x6360x)));
	assign x5986x = (((x155x) & (!x225x) & (!x5971x) & (!x5972x) & (!x5974x)) + ((!x155x) & (x225x) & (!x5971x) & (!x5972x) & (!x5974x)) + ((!x155x) & (!x225x) & (x5971x) & (!x5972x) & (!x5974x)) + ((!x155x) & (!x225x) & (!x5971x) & (x5972x) & (!x5974x)) + ((!x155x) & (!x225x) & (!x5971x) & (!x5972x) & (x5974x)));
	assign x6024x = (((x6009x) & (!x6010x) & (!x6011x) & (!x6012x)) + ((!x6009x) & (x6010x) & (!x6011x) & (!x6012x)) + ((!x6009x) & (!x6010x) & (x6011x) & (!x6012x)) + ((!x6009x) & (!x6010x) & (!x6011x) & (x6012x)));
	assign x6025x = (((x6013x) & (!x6014x) & (!x6015x) & (!x6016x)) + ((!x6013x) & (x6014x) & (!x6015x) & (!x6016x)) + ((!x6013x) & (!x6014x) & (x6015x) & (!x6016x)) + ((!x6013x) & (!x6014x) & (!x6015x) & (x6016x)));
	assign n_n80 = (((!i_3_) & (!i_2_) & (i_0_)));
	assign n_n75 = (((!i_7_) & (i_8_)));
	assign x341x = (((i_5_) & (i_4_)));
	assign n_n81 = (((i_5_) & (i_3_) & (i_4_)));
	assign n_n38 = (((i_7_) & (!i_6_)));
	assign n_n64 = (((i_7_) & (i_8_)));
	assign n_n58 = (((i_7_) & (i_8_) & (!i_6_)));
	assign n_n52 = (((i_7_) & (i_6_)));
	assign n_n101 = (((i_7_) & (!i_8_) & (i_6_)));
	assign n_n86 = (((!i_7_) & (!i_8_)));
	assign n_n93 = (((!i_7_) & (!i_8_) & (i_6_)));
	assign n_n73 = (((!i_7_) & (!i_6_)));
	assign n_n78 = (((!i_7_) & (!i_8_) & (!i_6_)));
	assign n_n91 = (((!i_7_) & (i_8_) & (i_6_)));
	assign x175x = (((i_1_) & (!i_0_)));
	assign x76x = (((!i_5_) & (!i_3_) & (!i_4_) & (i_2_) & (x175x)));
	assign n_n1281 = (((!i_7_) & (i_8_) & (i_6_) & (x76x)));
	assign n_n100 = (((!i_1_) & (!i_2_) & (i_0_)));
	assign x27x = (((!i_5_) & (i_3_) & (!i_4_) & (n_n100)));
	assign n_n1185 = (((!i_5_) & (i_3_) & (!i_4_) & (n_n78) & (n_n100)));
	assign x42x = (((i_5_) & (!i_3_) & (!i_4_) & (i_2_) & (x108x)));
	assign n_n1120 = (((i_5_) & (i_3_) & (!i_4_) & (n_n83) & (n_n95)));
	assign x355x = (((!i_7_) & (!i_6_) & (i_3_) & (x341x) & (n_n83)));
	assign n_n1156 = (((!i_7_) & (i_8_) & (i_6_) & (x128x)));
	assign n_n1021 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n85) & (n_n82)));
	assign x4837x = (((!n_n100) & (!n_n70) & (!n_n54) & (n_n1134) & (!n_n1091)) + ((!n_n100) & (!n_n70) & (!n_n54) & (!n_n1134) & (n_n1091)) + ((n_n100) & (n_n70) & (n_n54) & (!n_n1134) & (!n_n1091)));
	assign x108x = (((i_1_) & (i_0_)));
	assign x57x = (((!i_5_) & (!i_3_) & (!i_4_) & (i_2_) & (x108x)));
	assign n_n92 = (((i_5_) & (i_3_) & (!i_4_)));
	assign n_n103 = (((i_1_) & (i_2_) & (!i_0_)));
	assign x26x = (((i_5_) & (i_3_) & (!i_4_) & (i_2_) & (x175x)));
	assign n_n84 = (((!i_5_) & (i_3_) & (!i_4_)));
	assign n_n83 = (((!i_1_) & (i_2_) & (i_0_)));
	assign x32x = (((!i_1_) & (i_2_) & (i_0_) & (n_n91)));
	assign n_n102 = (((!i_5_) & (i_3_) & (i_4_)));
	assign n_n94 = (((i_1_) & (!i_2_) & (!i_0_)));
	assign x39x = (((!i_5_) & (i_3_) & (i_4_) & (!i_2_) & (x175x)));
	assign n_n74 = (((!i_5_) & (!i_3_) & (i_4_)));
	assign n_n97 = (((i_1_) & (i_2_) & (i_0_)));
	assign x45x = (((i_5_) & (i_3_) & (!i_4_) & (n_n100)));
	assign x55x = (((i_5_) & (!i_3_) & (!i_4_) & (!i_2_) & (x175x)));
	assign x325x = (((!i_5_) & (i_4_)));
	assign x58x = (((i_3_) & (!i_1_) & (i_2_) & (i_0_) & (x325x)));
	assign x64x = (((!i_5_) & (!i_3_) & (i_4_) & (n_n100)));
	assign x75x = (((!i_1_) & (i_2_)));
	assign n_n1217 = (((i_1_) & (i_2_) & (!i_0_) & (n_n101) & (n_n74)));
	assign n_n77 = (((i_5_) & (!i_3_) & (i_4_)));
	assign x87x = (((!i_7_) & (!i_6_) & (!n_n97) & (n_n1217) & (!n_n77)) + ((!i_7_) & (!i_6_) & (n_n97) & (!n_n1217) & (n_n77)));
	assign n_n95 = (((i_7_) & (i_8_) & (i_6_)));
	assign x104x = (((!n_n91) & (n_n92) & (n_n100) & (n_n95) & (!n_n77)) + ((n_n91) & (!n_n92) & (n_n100) & (!n_n95) & (n_n77)));
	assign x112x = (((i_5_) & (i_3_) & (i_4_) & (i_0_) & (x75x)));
	assign x56x = (((i_3_) & (i_0_)));
	assign x318x = (((!i_7_) & (!i_8_) & (!i_5_) & (!i_6_) & (i_4_)));
	assign x63x = (((i_5_) & (!i_3_) & (!i_4_) & (i_2_) & (x175x)));
	assign x113x = (((!i_1_) & (n_n101) & (!x56x) & (!x318x) & (x63x)) + ((!i_1_) & (!n_n101) & (x56x) & (x318x) & (!x63x)));
	assign n_n70 = (((i_7_) & (!i_8_)));
	assign x172x = (((i_7_) & (!i_8_) & (i_4_)));
	assign x31x = (((!i_7_) & (!i_8_) & (i_6_) & (!i_2_) & (x175x)));
	assign x208x = (((n_n81) & (!n_n103) & (!n_n74) & (!n_n95) & (x31x)) + ((!n_n81) & (n_n103) & (n_n74) & (n_n95) & (!x31x)));
	assign x227x = (((!i_7_) & (i_8_) & (i_6_) & (x57x) & (!x42x)) + ((i_7_) & (!i_8_) & (i_6_) & (!x57x) & (x42x)));
	assign x235x = (((!i_7_) & (i_8_) & (i_6_) & (x42x)));
	assign x252x = (((!i_7_) & (!i_8_) & (i_6_) & (n_n92) & (n_n103)));
	assign n_n85 = (((i_1_) & (!i_2_) & (i_0_)));
	assign x311x = (((!i_6_) & (i_3_) & (!i_1_) & (!i_2_) & (i_0_)));
	assign x25x = (((i_5_) & (i_3_) & (i_4_) & (i_2_) & (x175x)));
	assign x329x = (((i_5_) & (i_3_) & (i_4_) & (n_n101) & (n_n103)));
	assign n_n54 = (((i_5_) & (!i_6_) & (!i_4_)));
	assign x337x = (((!i_7_) & (i_8_) & (i_5_) & (!i_6_) & (!i_4_)));
	assign x201x = (((!i_5_) & (!i_3_) & (!i_4_) & (n_n1036) & (!x107x)) + ((!i_5_) & (!i_3_) & (i_4_) & (!n_n1036) & (x107x)));
	assign x164x = (((!i_3_) & (n_n58) & (n_n83) & (!n_n95) & (!x110x)) + ((!i_3_) & (!n_n58) & (n_n83) & (n_n95) & (x110x)));
	assign x4887x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x34x) & (n_n1040)) + ((i_7_) & (i_8_) & (i_6_) & (x34x) & (!n_n1040)));
	assign x4888x = (((!i_6_) & (!n_n91) & (!x110x) & (!n_n67) & (x249x)) + ((i_6_) & (n_n91) & (x110x) & (n_n67) & (!x249x)));
	assign x4889x = (((!i_7_) & (!i_6_) & (!x22x) & (x324x) & (x327x)) + ((i_7_) & (!i_6_) & (x22x) & (!x324x) & (!x327x)));
	assign x4899x = (((x201x) & (!x164x) & (!x4887x) & (!x4888x) & (!x4889x)) + ((!x201x) & (x164x) & (!x4887x) & (!x4888x) & (!x4889x)) + ((!x201x) & (!x164x) & (x4887x) & (!x4888x) & (!x4889x)) + ((!x201x) & (!x164x) & (!x4887x) & (x4888x) & (!x4889x)) + ((!x201x) & (!x164x) & (!x4887x) & (!x4888x) & (x4889x)));
	assign x4891x = (((!i_5_) & (!n_n93) & (!n_n83) & (n_n1046) & (!x288x)) + ((!i_5_) & (!n_n93) & (!n_n83) & (!n_n1046) & (x288x)) + ((!i_5_) & (n_n93) & (n_n83) & (!n_n1046) & (!x288x)));
	assign x4892x = (((!i_8_) & (!n_n58) & (!x53x) & (n_n1052) & (!x70x)) + ((!i_8_) & (n_n58) & (x53x) & (!n_n1052) & (!x70x)) + ((!i_8_) & (!n_n58) & (!x53x) & (!n_n1052) & (x70x)));
	assign x4898x = (((!n_n82) & (!x237x) & (n_n1013) & (!x4885x) & (!x6348x)) + ((!n_n82) & (!x237x) & (!n_n1013) & (x4885x) & (!x6348x)) + ((!n_n82) & (!x237x) & (!n_n1013) & (!x4885x) & (!x6348x)) + ((n_n82) & (x237x) & (!n_n1013) & (!x4885x) & (!x6348x)));
	assign x298x = (((!i_2_) & (!n_n75) & (!x108x) & (!n_n76) & (x146x)) + ((!i_2_) & (n_n75) & (x108x) & (n_n76) & (!x146x)));
	assign x292x = (((!n_n80) & (!n_n70) & (n_n973) & (!n_n71) & (!n_n975)) + ((!n_n80) & (!n_n70) & (!n_n973) & (!n_n71) & (n_n975)) + ((n_n80) & (n_n70) & (!n_n973) & (n_n71) & (!n_n975)));
	assign n_n882 = (((!n_n78) & (!x64x) & (!n_n95) & (!x29x) & (x1557x)) + ((!n_n78) & (x64x) & (n_n95) & (!x29x) & (!x1557x)) + ((n_n78) & (!x64x) & (!n_n95) & (x29x) & (!x1557x)));
	assign x4910x = (((!i_7_) & (!i_0_) & (!n_n80) & (!n_n77) & (n_n943)) + ((i_7_) & (i_0_) & (!n_n80) & (n_n77) & (!n_n943)));
	assign x4913x = (((!n_n95) & (!x41x) & (n_n952) & (!n_n976) & (!n_n986)) + ((!n_n95) & (!x41x) & (!n_n952) & (n_n976) & (!n_n986)) + ((!n_n95) & (!x41x) & (!n_n952) & (!n_n976) & (n_n986)) + ((n_n95) & (x41x) & (!n_n952) & (!n_n976) & (!n_n986)));
	assign x4914x = (((!x42x) & (!n_n95) & (n_n984) & (!n_n1006) & (!n_n978)) + ((!x42x) & (!n_n95) & (!n_n984) & (n_n1006) & (!n_n978)) + ((!x42x) & (!n_n95) & (!n_n984) & (!n_n1006) & (n_n978)) + ((x42x) & (n_n95) & (!n_n984) & (!n_n1006) & (!n_n978)));
	assign x4917x = (((n_n982) & (!n_n967) & (!x204x) & (!x202x) & (!x203x)) + ((!n_n982) & (n_n967) & (!x204x) & (!x202x) & (!x203x)) + ((!n_n982) & (!n_n967) & (x204x) & (!x202x) & (!x203x)) + ((!n_n982) & (!n_n967) & (!x204x) & (x202x) & (!x203x)) + ((!n_n982) & (!n_n967) & (!x204x) & (!x202x) & (x203x)));
	assign x54x = (((!i_3_) & (i_4_)));
	assign n_n82 = (((i_7_) & (!i_8_) & (!i_6_)));
	assign n_n90 = (((!i_1_) & (i_2_) & (!i_0_)));
	assign n_n1172 = (((i_5_) & (i_3_) & (i_4_) & (n_n95) & (n_n90)));
	assign n_n1078 = (((!i_5_) & (!i_3_) & (!i_4_) & (n_n78) & (n_n97)));
	assign x245x = (((i_3_) & (i_2_) & (i_0_)));
	assign x38x = (((i_7_) & (i_8_) & (i_5_) & (!i_6_) & (!i_4_)));
	assign x43x = (((!i_5_) & (!i_3_) & (i_4_) & (!i_0_) & (x75x)));
	assign n_n1279 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n78) & (n_n90)));
	assign x61x = (((!i_7_) & (i_8_) & (!i_6_) & (x29x) & (!x23x)) + ((!i_7_) & (i_8_) & (i_6_) & (!x29x) & (x23x)));
	assign x139x = (((!i_3_) & (!x341x) & (!n_n94) & (n_n95) & (x239x)) + ((i_3_) & (x341x) & (n_n94) & (n_n95) & (!x239x)));
	assign x118x = (((!i_1_) & (n_n78) & (x52x) & (!x30x) & (!x339x)) + ((i_1_) & (!n_n78) & (!x52x) & (x30x) & (x339x)));
	assign x6352x = (((!n_n78) & (!n_n91) & (!x39x) & (!x55x) & (!x22x)) + ((!n_n78) & (!n_n91) & (!x39x) & (!x55x) & (!x22x)) + ((!n_n78) & (!n_n91) & (!x39x) & (!x55x) & (!x22x)) + ((!n_n78) & (!n_n91) & (!x39x) & (!x55x) & (!x22x)));
	assign n_n137 = (((x61x) & (!x139x) & (!x118x) & (!x6352x)) + ((!x61x) & (x139x) & (!x118x) & (!x6352x)) + ((!x61x) & (!x139x) & (x118x) & (!x6352x)) + ((!x61x) & (!x139x) & (!x118x) & (!x6352x)));
	assign x111x = (((i_8_) & (!i_6_)));
	assign x41x = (((!i_5_) & (i_3_) & (i_4_) & (n_n100)));
	assign x4927x = (((!i_7_) & (!i_8_) & (!i_6_) & (x25x) & (!x21x)) + ((i_7_) & (!i_8_) & (i_6_) & (!x25x) & (x21x)));
	assign x340x = (((i_5_) & (i_3_) & (!i_4_) & (n_n91) & (n_n85)));
	assign x4934x = (((!n_n93) & (!n_n102) & (!x175x) & (x354x) & (x62x)) + ((n_n93) & (n_n102) & (x175x) & (!x354x) & (!x62x)));
	assign x4936x = (((!i_4_) & (!n_n75) & (!x311x) & (x340x) & (!x4934x)) + ((!i_4_) & (!n_n75) & (!x311x) & (!x340x) & (x4934x)) + ((i_4_) & (n_n75) & (x311x) & (!x340x) & (!x4934x)));
	assign n_n1153 = (((!i_5_) & (i_3_) & (i_4_) & (n_n58) & (n_n90)));
	assign x44x = (((!i_5_) & (i_3_) & (!i_4_) & (!i_2_) & (x108x)));
	assign x4938x = (((i_7_) & (!i_8_) & (n_n92) & (n_n85) & (!n_n87)) + ((!i_7_) & (i_8_) & (!n_n92) & (n_n85) & (n_n87)));
	assign x304x = (((!n_n58) & (!n_n101) & (!x57x) & (!x25x) & (x350x)) + ((!n_n58) & (n_n101) & (x57x) & (!x25x) & (!x350x)) + ((n_n58) & (!n_n101) & (!x57x) & (x25x) & (!x350x)));
	assign x4943x = (((!i_7_) & (!i_8_) & (!x44x) & (x4938x) & (!x304x)) + ((!i_7_) & (!i_8_) & (!x44x) & (!x4938x) & (x304x)) + ((!i_7_) & (!i_8_) & (x44x) & (!x4938x) & (!x304x)));
	assign n_n1297 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n95) & (n_n90)));
	assign n_n1324 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n102) & (n_n90)));
	assign n_n1092 = (((!i_5_) & (i_3_) & (!i_4_) & (n_n91) & (n_n100)));
	assign n_n1103 = (((!i_1_) & (i_2_) & (i_0_) & (n_n102) & (n_n95)));
	assign x319x = (((!i_7_) & (i_5_) & (!i_6_) & (x54x) & (n_n90)));
	assign n_n1130 = (((i_7_) & (i_8_) & (!i_6_) & (n_n84) & (n_n85)));
	assign x354x = (((!i_5_) & (!i_6_) & (i_3_)));
	assign x4944x = (((i_7_) & (!i_8_) & (i_1_) & (!i_2_) & (!i_0_)));
	assign x4950x = (((n_n1103) & (!x319x) & (!n_n1130) & (!x354x) & (!x4944x)) + ((!n_n1103) & (x319x) & (!n_n1130) & (!x354x) & (!x4944x)) + ((!n_n1103) & (!x319x) & (n_n1130) & (!x354x) & (!x4944x)) + ((!n_n1103) & (!x319x) & (!n_n1130) & (x354x) & (x4944x)));
	assign n_n1105 = (((i_5_) & (i_3_) & (i_4_) & (n_n58) & (n_n94)));
	assign n_n1108 = (((i_5_) & (i_3_) & (i_4_) & (n_n93) & (n_n90)));
	assign x94x = (((!i_7_) & (!i_8_) & (!n_n84) & (!n_n83) & (n_n1100)) + ((i_7_) & (i_8_) & (n_n84) & (n_n83) & (!n_n1100)));
	assign x4951x = (((!n_n63) & (!x44x) & (n_n1105) & (!n_n1108) & (!x94x)) + ((!n_n63) & (!x44x) & (!n_n1105) & (n_n1108) & (!x94x)) + ((!n_n63) & (!x44x) & (!n_n1105) & (!n_n1108) & (x94x)) + ((n_n63) & (x44x) & (!n_n1105) & (!n_n1108) & (!x94x)));
	assign x19x = (((i_5_) & (i_1_) & (i_2_) & (!i_0_) & (x54x)));
	assign x29x = (((!i_5_) & (i_3_) & (i_4_) & (i_2_) & (x108x)));
	assign x37x = (((i_1_) & (!i_2_) & (!i_0_) & (n_n38) & (n_n70)));
	assign x105x = (((n_n81) & (n_n91) & (n_n100) & (!n_n83) & (!n_n74)) + ((!n_n81) & (n_n91) & (!n_n100) & (n_n83) & (n_n74)));
	assign x109x = (((i_5_) & (!i_4_)));
	assign x127x = (((i_6_) & (!i_3_) & (i_4_)));
	assign n_n1082 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n97) & (n_n63)));
	assign x110x = (((!i_5_) & (!i_4_)));
	assign x1487x = (((!i_7_) & (!i_6_) & (!i_3_) & (n_n83) & (x110x)));
	assign x207x = (((n_n75) & (!n_n38) & (!n_n84) & (x55x) & (!n_n90)) + ((!n_n75) & (n_n38) & (n_n84) & (!x55x) & (n_n90)));
	assign x1483x = (((!i_7_) & (i_8_) & (!i_3_) & (n_n103) & (x109x)));
	assign x1484x = (((i_7_) & (!i_8_) & (i_3_) & (n_n85) & (x325x)));
	assign n_n67 = (((!i_3_) & (!i_1_) & (i_0_)));
	assign x1479x = (((i_7_) & (!i_6_) & (i_2_) & (n_n102) & (x175x)));
	assign x1480x = (((!i_1_) & (i_2_) & (i_0_) & (x35x)));
	assign x251x = (((!i_7_) & (i_8_) & (!i_6_) & (n_n103) & (n_n77)));
	assign n_n1079 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n81) & (n_n100)));
	assign x254x = (((!i_5_) & (!i_3_) & (!i_4_) & (n_n1079) & (!x31x)) + ((!i_5_) & (!i_3_) & (!i_4_) & (!n_n1079) & (x31x)));
	assign x321x = (((!i_5_) & (!i_3_) & (i_4_) & (n_n101) & (n_n97)));
	assign x328x = (((i_7_) & (i_8_) & (i_1_) & (i_2_) & (i_0_)));
	assign n_n1259 = (((!i_7_) & (i_8_) & (!i_6_) & (n_n92) & (n_n90)));
	assign x239x = (((i_5_) & (!i_3_) & (!i_4_) & (n_n100)));
	assign n_n1204 = (((i_7_) & (i_8_) & (i_6_) & (x239x)));
	assign x351x = (((!i_3_) & (!i_1_) & (!i_0_)));
	assign x21x = (((!i_5_) & (!i_3_) & (!i_4_) & (i_0_) & (x75x)));
	assign x256x = (((!i_3_) & (!n_n58) & (!n_n94) & (!x109x) & (n_n1085)) + ((!i_3_) & (n_n58) & (n_n94) & (x109x) & (!n_n1085)));
	assign x299x = (((!i_6_) & (!n_n86) & (!x43x) & (n_n1040) & (!x114x)) + ((!i_6_) & (!n_n86) & (!x43x) & (!n_n1040) & (x114x)) + ((i_6_) & (n_n86) & (x43x) & (!n_n1040) & (!x114x)));
	assign x5006x = (((!n_n102) & (n_n1095) & (!x20x) & (!n_n1088) & (!n_n1181)) + ((!n_n102) & (!n_n1095) & (!x20x) & (n_n1088) & (!n_n1181)) + ((!n_n102) & (!n_n1095) & (!x20x) & (!n_n1088) & (n_n1181)) + ((n_n102) & (!n_n1095) & (x20x) & (!n_n1088) & (!n_n1181)));
	assign x190x = (((!i_5_) & (!i_3_) & (!i_4_) & (!x32x) & (n_n1160)) + ((!i_5_) & (i_3_) & (!i_4_) & (x32x) & (!n_n1160)));
	assign x265x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x63x) & (n_n1146)) + ((!i_7_) & (!i_8_) & (!i_6_) & (x63x) & (!n_n1146)));
	assign x5003x = (((!n_n58) & (!x64x) & (n_n1132) & (!x335x) & (!x1440x)) + ((!n_n58) & (!x64x) & (!n_n1132) & (x335x) & (!x1440x)) + ((!n_n58) & (!x64x) & (!n_n1132) & (!x335x) & (x1440x)) + ((n_n58) & (x64x) & (!n_n1132) & (!x335x) & (!x1440x)));
	assign x5004x = (((!x337x) & (n_n1172) & (!n_n1022) & (!x322x) & (!n_n1128)) + ((!x337x) & (!n_n1172) & (n_n1022) & (!x322x) & (!n_n1128)) + ((!x337x) & (!n_n1172) & (!n_n1022) & (!x322x) & (n_n1128)) + ((x337x) & (!n_n1172) & (!n_n1022) & (x322x) & (!n_n1128)));
	assign x5005x = (((!n_n58) & (n_n1036) & (!x44x) & (!n_n1060) & (!n_n1164)) + ((!n_n58) & (!n_n1036) & (!x44x) & (n_n1060) & (!n_n1164)) + ((!n_n58) & (!n_n1036) & (!x44x) & (!n_n1060) & (n_n1164)) + ((n_n58) & (!n_n1036) & (x44x) & (!n_n1060) & (!n_n1164)));
	assign x135x = (((!i_4_) & (!i_1_) & (!i_2_) & (!i_0_) & (!x28x)) + ((!i_4_) & (!i_1_) & (!i_2_) & (!i_0_) & (x28x)));
	assign n_n949 = (((!i_5_) & (i_3_) & (!i_4_) & (n_n101) & (n_n85)));
	assign x97x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x49x) & (n_n941)) + ((!i_7_) & (!i_8_) & (i_6_) & (x49x) & (!n_n941)));
	assign x204x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x52x) & (n_n951)) + ((i_7_) & (i_8_) & (i_6_) & (x52x) & (!n_n951)));
	assign x5025x = (((!x25x) & (!n_n82) & (n_n1021) & (!x249x) & (!n_n978)) + ((!x25x) & (!n_n82) & (!n_n1021) & (x249x) & (!n_n978)) + ((!x25x) & (!n_n82) & (!n_n1021) & (!x249x) & (n_n978)) + ((x25x) & (n_n82) & (!n_n1021) & (!x249x) & (!n_n978)));
	assign x195x = (((!i_0_) & (n_n78) & (!x75x) & (x42x) & (!x5012x)) + ((!i_0_) & (!n_n78) & (x75x) & (!x42x) & (x5012x)));
	assign x151x = (((!i_3_) & (!x341x) & (!n_n78) & (!n_n100) & (n_n1018)) + ((i_3_) & (x341x) & (n_n78) & (n_n100) & (!n_n1018)));
	assign x5021x = (((!n_n103) & (!n_n74) & (!n_n82) & (x79x) & (!n_n975)) + ((!n_n103) & (!n_n74) & (!n_n82) & (!x79x) & (n_n975)) + ((n_n103) & (n_n74) & (n_n82) & (!x79x) & (!n_n975)));
	assign x5023x = (((!n_n78) & (!x29x) & (n_n967) & (!n_n969) & (!x1557x)) + ((!n_n78) & (!x29x) & (!n_n967) & (n_n969) & (!x1557x)) + ((!n_n78) & (!x29x) & (!n_n967) & (!n_n969) & (x1557x)) + ((n_n78) & (x29x) & (!n_n967) & (!n_n969) & (!x1557x)));
	assign x5024x = (((!n_n95) & (!x41x) & (!x128x) & (!x44x) & (n_n1004)) + ((n_n95) & (x41x) & (!x128x) & (!x44x) & (!n_n1004)) + ((n_n95) & (!x41x) & (x128x) & (!x44x) & (!n_n1004)) + ((n_n95) & (!x41x) & (!x128x) & (x44x) & (!n_n1004)));
	assign x34x = (((!i_5_) & (!i_3_) & (!i_4_) & (!i_2_) & (x108x)));
	assign x23x = (((i_5_) & (i_3_) & (i_4_) & (i_2_) & (x108x)));
	assign n_n1188 = (((i_5_) & (i_3_) & (i_4_) & (n_n58) & (n_n90)));
	assign x88x = (((!i_6_) & (!n_n86) & (!n_n74) & (!n_n97) & (n_n1188)) + ((i_6_) & (n_n86) & (n_n74) & (n_n97) & (!n_n1188)));
	assign x346x = (((!i_5_) & (!i_3_) & (i_4_) & (n_n100) & (n_n82)));
	assign x1413x = (((i_5_) & (i_3_) & (!i_4_) & (n_n103) & (n_n82)));
	assign x1414x = (((!i_7_) & (i_8_) & (!i_6_) & (n_n81) & (n_n97)));
	assign x343x = (((i_5_) & (i_3_) & (!i_4_) & (n_n101) & (n_n103)));
	assign x1518x = (((i_7_) & (!i_8_) & (!i_6_) & (x34x)));
	assign x1519x = (((i_5_) & (!i_3_) & (i_4_) & (n_n58) & (n_n100)));
	assign x231x = (((!i_3_) & (!x38x) & (!x108x) & (x1518x) & (!x1519x)) + ((!i_3_) & (!x38x) & (!x108x) & (!x1518x) & (x1519x)) + ((!i_3_) & (x38x) & (x108x) & (!x1518x) & (!x1519x)));
	assign n_n1193 = (((i_7_) & (i_8_) & (!i_6_) & (n_n84) & (n_n94)));
	assign x255x = (((!n_n58) & (n_n78) & (n_n100) & (n_n84) & (!n_n94)) + ((n_n58) & (!n_n78) & (!n_n100) & (n_n84) & (n_n94)));
	assign x46x = (((i_5_) & (i_3_) & (!i_4_) & (!i_2_) & (x108x)));
	assign x5031x = (((i_7_) & (i_8_) & (i_6_) & (x46x) & (!x41x)) + ((!i_7_) & (!i_8_) & (i_6_) & (!x46x) & (x41x)));
	assign x301x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x21x) & (x5031x)) + ((!i_7_) & (i_8_) & (i_6_) & (x21x) & (!x5031x)));
	assign x53x = (((!i_5_) & (i_3_) & (i_4_) & (!i_2_) & (x108x)));
	assign n_n1022 = (((i_7_) & (i_8_) & (!i_6_) & (n_n102) & (n_n85)));
	assign n_n1134 = (((i_7_) & (i_8_) & (!i_6_) & (n_n100) & (n_n74)));
	assign n_n1039 = (((!i_5_) & (i_3_) & (i_4_) & (n_n78) & (n_n94)));
	assign x78x = (((i_7_) & (i_8_) & (i_5_) & (!i_6_) & (i_4_)));
	assign n_n87 = (((i_5_) & (!i_6_) & (i_4_)));
	assign n_n1091 = (((i_3_) & (!i_2_) & (i_0_) & (n_n64) & (n_n87)));
	assign x5060x = (((!n_n58) & (!x25x) & (n_n1153) & (!n_n1267) & (!x342x)) + ((!n_n58) & (!x25x) & (!n_n1153) & (n_n1267) & (!x342x)) + ((!n_n58) & (!x25x) & (!n_n1153) & (!n_n1267) & (x342x)) + ((n_n58) & (x25x) & (!n_n1153) & (!n_n1267) & (!x342x)));
	assign x5061x = (((!n_n95) & (!x67x) & (n_n1216) & (!n_n1146) & (!n_n1164)) + ((!n_n95) & (!x67x) & (!n_n1216) & (n_n1146) & (!n_n1164)) + ((!n_n95) & (!x67x) & (!n_n1216) & (!n_n1146) & (n_n1164)) + ((n_n95) & (x67x) & (!n_n1216) & (!n_n1146) & (!n_n1164)));
	assign x5062x = (((!n_n101) & (!n_n92) & (!n_n103) & (n_n1170) & (!x5056x)) + ((!n_n101) & (!n_n92) & (!n_n103) & (!n_n1170) & (x5056x)) + ((n_n101) & (n_n92) & (n_n103) & (!n_n1170) & (!x5056x)));
	assign x5063x = (((x87x) & (!x61x) & (!x224x) & (!x1384x)) + ((!x87x) & (x61x) & (!x224x) & (!x1384x)) + ((!x87x) & (!x61x) & (x224x) & (!x1384x)) + ((!x87x) & (!x61x) & (!x224x) & (x1384x)));
	assign x5064x = (((x206x) & (!x225x) & (!x5059x)) + ((!x206x) & (x225x) & (!x5059x)) + ((!x206x) & (!x225x) & (x5059x)));
	assign x5076x = (((!x42x) & (!n_n95) & (n_n983) & (!n_n999) & (!x249x)) + ((!x42x) & (!n_n95) & (!n_n983) & (n_n999) & (!x249x)) + ((!x42x) & (!n_n95) & (!n_n983) & (!n_n999) & (x249x)) + ((x42x) & (n_n95) & (!n_n983) & (!n_n999) & (!x249x)));
	assign x5077x = (((n_n951) & (!n_n954) & (!n_n952) & (!x147x) & (!x202x)) + ((!n_n951) & (n_n954) & (!n_n952) & (!x147x) & (!x202x)) + ((!n_n951) & (!n_n954) & (n_n952) & (!x147x) & (!x202x)) + ((!n_n951) & (!n_n954) & (!n_n952) & (x147x) & (!x202x)) + ((!n_n951) & (!n_n954) & (!n_n952) & (!x147x) & (x202x)));
	assign x5078x = (((x294x) & (!x146x) & (!n_n1001) & (!n_n1010) & (!n_n978)) + ((!x294x) & (x146x) & (!n_n1001) & (!n_n1010) & (!n_n978)) + ((!x294x) & (!x146x) & (n_n1001) & (!n_n1010) & (!n_n978)) + ((!x294x) & (!x146x) & (!n_n1001) & (n_n1010) & (!n_n978)) + ((!x294x) & (!x146x) & (!n_n1001) & (!n_n1010) & (n_n978)));
	assign x5079x = (((x97x) & (!n_n939) & (!n_n981) & (!x272x) & (!x151x)) + ((!x97x) & (n_n939) & (!n_n981) & (!x272x) & (!x151x)) + ((!x97x) & (!n_n939) & (n_n981) & (!x272x) & (!x151x)) + ((!x97x) & (!n_n939) & (!n_n981) & (x272x) & (!x151x)) + ((!x97x) & (!n_n939) & (!n_n981) & (!x272x) & (x151x)));
	assign x322x = (((!i_3_) & (i_2_) & (!i_0_)));
	assign n_n1093 = (((!i_7_) & (i_8_) & (!i_6_) & (x109x) & (x322x)));
	assign n_n1052 = (((i_1_) & (!i_2_) & (!i_0_) & (n_n74) & (n_n63)));
	assign n_n1331 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n91) & (n_n90)));
	assign n_n40 = (((!i_5_) & (!i_6_) & (i_4_)));
	assign x35x = (((!i_3_) & (n_n75) & (!n_n38) & (!x109x) & (n_n40)) + ((!i_3_) & (!n_n75) & (n_n38) & (x109x) & (!n_n40)));
	assign x1359x = (((!i_5_) & (!i_3_) & (i_4_) & (n_n94) & (n_n82)));
	assign n_n66 = (((i_5_) & (i_6_) & (!i_4_)));
	assign x20x = (((!i_7_) & (!i_8_) & (i_6_) & (!i_2_) & (x108x)));
	assign x353x = (((!i_3_) & (!i_1_) & (i_2_)));
	assign x117x = (((!n_n86) & (n_n77) & (!n_n66) & (x20x) & (!x353x)) + ((n_n86) & (!n_n77) & (n_n66) & (!x20x) & (x353x)));
	assign n_n1058 = (((i_1_) & (!i_2_) & (!i_0_) & (n_n58) & (n_n74)));
	assign x133x = (((!i_7_) & (!i_6_) & (!n_n103) & (!n_n84) & (n_n1058)) + ((i_7_) & (!i_6_) & (n_n103) & (n_n84) & (!n_n1058)));
	assign n_n1032 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n74) & (n_n90)));
	assign n_n1040 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n85) & (n_n95)));
	assign x148x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x43x) & (n_n1040)) + ((!i_7_) & (!i_8_) & (i_6_) & (x43x) & (!n_n1040)));
	assign x173x = (((!i_7_) & (i_6_)));
	assign x177x = (((!i_7_) & (i_8_) & (i_6_)) + ((i_7_) & (!i_8_) & (i_6_)));
	assign x323x = (((!i_5_) & (!i_3_) & (!i_4_) & (n_n94) & (n_n82)));
	assign x1352x = (((!i_5_) & (i_3_) & (!i_4_) & (n_n100) & (n_n95)));
	assign n_n1036 = (((i_1_) & (i_2_) & (!i_0_) & (n_n91) & (n_n74)));
	assign x107x = (((i_1_) & (!i_2_) & (i_0_) & (n_n101)));
	assign x233x = (((n_n58) & (!n_n91) & (n_n103) & (n_n77) & (!n_n90)) + ((!n_n58) & (n_n91) & (n_n103) & (n_n77) & (!n_n90)) + ((n_n58) & (!n_n91) & (!n_n103) & (n_n77) & (n_n90)));
	assign n_n1085 = (((!i_5_) & (i_3_) & (i_4_) & (n_n94) & (n_n63)));
	assign x5083x = (((!i_7_) & (!i_6_) & (!n_n97) & (n_n1078) & (!n_n77)) + ((i_7_) & (i_6_) & (n_n97) & (!n_n1078) & (n_n77)));
	assign x1348x = (((!i_7_) & (!i_6_) & (!i_3_) & (n_n100) & (x110x)));
	assign x257x = (((!n_n101) & (!n_n74) & (!n_n90) & (x5083x) & (!x1348x)) + ((!n_n101) & (!n_n74) & (!n_n90) & (!x5083x) & (x1348x)) + ((n_n101) & (n_n74) & (n_n90) & (!x5083x) & (!x1348x)));
	assign x237x = (((!i_5_) & (!i_1_) & (i_2_) & (i_0_) & (x54x)));
	assign x5085x = (((i_7_) & (!i_8_) & (i_6_) & (i_3_) & (i_4_)));
	assign x271x = (((!i_2_) & (n_n82) & (!x175x) & (x237x) & (!x5085x)) + ((!i_2_) & (!n_n82) & (x175x) & (!x237x) & (x5085x)));
	assign x296x = (((!n_n84) & (!n_n83) & (!n_n82) & (n_n983) & (!n_n986)) + ((!n_n84) & (!n_n83) & (!n_n82) & (!n_n983) & (n_n986)) + ((n_n84) & (n_n83) & (n_n82) & (!n_n983) & (!n_n986)));
	assign x5121x = (((!n_n95) & (!x41x) & (n_n949) & (!n_n969) & (!n_n966)) + ((!n_n95) & (!x41x) & (!n_n949) & (n_n969) & (!n_n966)) + ((!n_n95) & (!x41x) & (!n_n949) & (!n_n969) & (n_n966)) + ((n_n95) & (x41x) & (!n_n949) & (!n_n969) & (!n_n966)));
	assign x5123x = (((x271x) & (!n_n944) & (!x145x) & (!x146x) & (!n_n939)) + ((!x271x) & (n_n944) & (!x145x) & (!x146x) & (!n_n939)) + ((!x271x) & (!n_n944) & (x145x) & (!x146x) & (!n_n939)) + ((!x271x) & (!n_n944) & (!x145x) & (x146x) & (!n_n939)) + ((!x271x) & (!n_n944) & (!x145x) & (!x146x) & (n_n939)));
	assign x5124x = (((x189x) & (!n_n958) & (!x270x) & (!x272x) & (!x5114x)) + ((!x189x) & (n_n958) & (!x270x) & (!x272x) & (!x5114x)) + ((!x189x) & (!n_n958) & (x270x) & (!x272x) & (!x5114x)) + ((!x189x) & (!n_n958) & (!x270x) & (x272x) & (!x5114x)) + ((!x189x) & (!n_n958) & (!x270x) & (!x272x) & (x5114x)));
	assign x52x = (((i_3_) & (i_1_) & (i_2_) & (!i_0_) & (x325x)));
	assign x306x = (((!n_n93) & (!x57x) & (!n_n63) & (!x83x) & (n_n1177)) + ((n_n93) & (x57x) & (!n_n63) & (!x83x) & (!n_n1177)) + ((!n_n93) & (!x57x) & (n_n63) & (x83x) & (!n_n1177)));
	assign x5135x = (((!i_6_) & (!n_n86) & (x257x) & (!n_n1158) & (!x65x)) + ((!i_6_) & (!n_n86) & (!x257x) & (n_n1158) & (!x65x)) + ((i_6_) & (n_n86) & (!x257x) & (!n_n1158) & (x65x)));
	assign x141x = (((!i_3_) & (n_n52) & (x39x) & (!x110x) & (!x31x)) + ((!i_3_) & (!n_n52) & (!x39x) & (x110x) & (x31x)));
	assign x279x = (((!i_0_) & (!n_n102) & (!x75x) & (!n_n95) & (n_n1095)) + ((i_0_) & (n_n102) & (x75x) & (n_n95) & (!n_n1095)));
	assign x5131x = (((!i_8_) & (!i_6_) & (!n_n81) & (!n_n85) & (x133x)) + ((i_8_) & (!i_6_) & (n_n81) & (n_n85) & (!x133x)));
	assign x5133x = (((!n_n91) & (!n_n100) & (!n_n84) & (n_n1153) & (!x267x)) + ((!n_n91) & (!n_n100) & (!n_n84) & (!n_n1153) & (x267x)) + ((n_n91) & (n_n100) & (n_n84) & (!n_n1153) & (!x267x)));
	assign x5134x = (((!n_n74) & (n_n1082) & (!n_n1120) & (!n_n1052) & (!x107x)) + ((!n_n74) & (!n_n1082) & (n_n1120) & (!n_n1052) & (!x107x)) + ((!n_n74) & (!n_n1082) & (!n_n1120) & (n_n1052) & (!x107x)) + ((n_n74) & (!n_n1082) & (!n_n1120) & (!n_n1052) & (x107x)));
	assign x67x = (((!i_5_) & (i_3_) & (!i_4_) & (!i_2_) & (x175x)));
	assign n_n1330 = (((!i_5_) & (i_3_) & (i_4_) & (n_n95) & (n_n90)));
	assign n_n1267 = (((!i_5_) & (i_3_) & (!i_4_) & (n_n101) & (n_n100)));
	assign x36x = (((i_5_) & (!i_3_) & (i_4_) & (!i_0_) & (x75x)));
	assign x48x = (((!i_1_) & (i_2_) & (i_0_) & (n_n73) & (x111x)));
	assign x72x = (((i_7_) & (!i_5_) & (!i_3_) & (!i_4_) & (!i_0_)) + ((!i_7_) & (!i_5_) & (!i_3_) & (!i_4_) & (!i_0_)));
	assign x1291x = (((i_1_) & (i_2_) & (!i_0_) & (n_n101) & (n_n84)));
	assign x1292x = (((i_5_) & (i_3_) & (!i_4_) & (n_n93) & (n_n85)));
	assign x327x = (((i_2_) & (i_0_)));
	assign x123x = (((!i_3_) & (n_n93) & (!x38x) & (x19x) & (!x327x)) + ((!i_3_) & (!n_n93) & (x38x) & (!x19x) & (x327x)));
	assign x183x = (((!n_n93) & (x76x) & (!n_n84) & (n_n63) & (!n_n90)) + ((n_n93) & (!x76x) & (n_n84) & (!n_n63) & (n_n90)));
	assign x1285x = (((!i_5_) & (!i_3_) & (i_4_) & (n_n78) & (n_n97)));
	assign x348x = (((i_5_) & (!i_3_) & (i_4_) & (n_n78) & (n_n100)));
	assign x128x = (((!i_5_) & (!i_3_) & (!i_4_) & (!i_2_) & (x175x)));
	assign x186x = (((!i_7_) & (!i_8_) & (!i_6_) & (x348x) & (!x128x)) + ((i_7_) & (i_8_) & (!i_6_) & (!x348x) & (x128x)));
	assign x206x = (((!i_2_) & (!n_n101) & (!n_n84) & (x108x) & (x78x)) + ((i_2_) & (n_n101) & (n_n84) & (x108x) & (!x78x)));
	assign n_n76 = (((i_5_) & (!i_6_) & (i_3_)));
	assign n_n1215 = (((i_7_) & (i_8_) & (!i_6_) & (x239x)));
	assign x342x = (((!i_7_) & (!i_6_) & (!i_2_) & (n_n77) & (x175x)));
	assign x5176x = (((!i_7_) & (!i_6_) & (n_n1082) & (!x21x) & (!x52x)) + ((!i_7_) & (!i_6_) & (!n_n1082) & (x21x) & (!x52x)) + ((i_7_) & (!i_6_) & (!n_n1082) & (!x21x) & (x52x)));
	assign x5181x = (((!x48x) & (n_n1216) & (!n_n1088) & (!n_n1181) & (!x194x)) + ((!x48x) & (!n_n1216) & (n_n1088) & (!n_n1181) & (!x194x)) + ((!x48x) & (!n_n1216) & (!n_n1088) & (n_n1181) & (!x194x)) + ((x48x) & (!n_n1216) & (!n_n1088) & (!n_n1181) & (x194x)));
	assign x5178x = (((!i_7_) & (!i_6_) & (!x34x) & (n_n1215) & (!x190x)) + ((!i_7_) & (!i_6_) & (!x34x) & (!n_n1215) & (x190x)) + ((i_7_) & (i_6_) & (x34x) & (!n_n1215) & (!x190x)));
	assign x5179x = (((!n_n100) & (n_n1204) & (!x78x) & (!n_n1128) & (!n_n1184)) + ((!n_n100) & (!n_n1204) & (!x78x) & (n_n1128) & (!n_n1184)) + ((!n_n100) & (!n_n1204) & (!x78x) & (!n_n1128) & (n_n1184)) + ((n_n100) & (!n_n1204) & (x78x) & (!n_n1128) & (!n_n1184)));
	assign x5180x = (((!n_n91) & (!x63x) & (n_n1132) & (!n_n1130) & (!x335x)) + ((!n_n91) & (!x63x) & (!n_n1132) & (n_n1130) & (!x335x)) + ((!n_n91) & (!x63x) & (!n_n1132) & (!n_n1130) & (x335x)) + ((n_n91) & (x63x) & (!n_n1132) & (!n_n1130) & (!x335x)));
	assign x125x = (((!n_n101) & (!x42x) & (!n_n95) & (n_n942) & (!x52x)) + ((!n_n101) & (x42x) & (n_n95) & (!n_n942) & (!x52x)) + ((n_n101) & (!x42x) & (!n_n95) & (!n_n942) & (x52x)));
	assign x5193x = (((!i_2_) & (!x38x) & (!x108x) & (n_n973) & (!n_n975)) + ((!i_2_) & (!x38x) & (!x108x) & (!n_n973) & (n_n975)) + ((!i_2_) & (x38x) & (x108x) & (!n_n973) & (!n_n975)));
	assign x5198x = (((!n_n95) & (!x52x) & (!x128x) & (n_n986) & (!n_n1042)) + ((!n_n95) & (!x52x) & (!x128x) & (!n_n986) & (n_n1042)) + ((n_n95) & (x52x) & (!x128x) & (!n_n986) & (!n_n1042)) + ((n_n95) & (!x52x) & (x128x) & (!n_n986) & (!n_n1042)));
	assign x5196x = (((!n_n91) & (!x29x) & (x189x) & (!n_n958) & (!n_n1060)) + ((!n_n91) & (!x29x) & (!x189x) & (n_n958) & (!n_n1060)) + ((!n_n91) & (!x29x) & (!x189x) & (!n_n958) & (n_n1060)) + ((n_n91) & (x29x) & (!x189x) & (!n_n958) & (!n_n1060)));
	assign x5197x = (((!x64x) & (!n_n95) & (n_n980) & (!n_n999) & (!n_n1004)) + ((!x64x) & (!n_n95) & (!n_n980) & (n_n999) & (!n_n1004)) + ((!x64x) & (!n_n95) & (!n_n980) & (!n_n999) & (n_n1004)) + ((x64x) & (n_n95) & (!n_n980) & (!n_n999) & (!n_n1004)));
	assign x5200x = (((n_n967) & (!n_n966) & (!x147x) & (!x195x) & (!x274x)) + ((!n_n967) & (n_n966) & (!x147x) & (!x195x) & (!x274x)) + ((!n_n967) & (!n_n966) & (x147x) & (!x195x) & (!x274x)) + ((!n_n967) & (!n_n966) & (!x147x) & (x195x) & (!x274x)) + ((!n_n967) & (!n_n966) & (!x147x) & (!x195x) & (x274x)));
	assign x62x = (((!i_7_) & (!i_8_) & (!i_1_) & (i_2_) & (i_0_)));
	assign x185x = (((!i_6_) & (n_n91) & (x34x) & (!x110x) & (!x62x)) + ((!i_6_) & (!n_n91) & (!x34x) & (x110x) & (x62x)));
	assign x352x = (((i_5_) & (!i_3_) & (!i_4_) & (n_n78) & (n_n90)));
	assign n_n1074 = (((i_1_) & (!i_2_) & (!i_0_) & (n_n101) & (n_n74)));
	assign n_n1294 = (((!i_5_) & (i_3_) & (!i_4_) & (n_n78) & (n_n90)));
	assign n_n1109 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n101) & (n_n90)));
	assign n_n1132 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n93) & (n_n90)));
	assign x28x = (((!i_6_) & (!i_3_)));
	assign x131x = (((!i_6_) & (!i_3_) & (!i_4_)));
	assign x5012x = (((!i_5_) & (i_6_) & (!i_3_) & (!i_4_)));
	assign n_n1312 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n101) & (n_n90)));
	assign x326x = (((i_1_) & (!i_2_) & (!i_0_) & (n_n101) & (n_n77)));
	assign n_n1169 = (((!i_5_) & (i_3_) & (i_4_) & (n_n91) & (n_n90)));
	assign n_n942 = (((i_5_) & (i_3_) & (!i_4_) & (n_n91) & (n_n94)));
	assign n_n1057 = (((i_5_) & (i_3_) & (i_4_) & (n_n82) & (n_n90)));
	assign n_n1125 = (((i_5_) & (i_3_) & (i_4_) & (n_n78) & (n_n90)));
	assign n_n1128 = (((!i_5_) & (i_3_) & (!i_4_) & (n_n78) & (n_n94)));
	assign x333x = (((i_7_) & (i_6_) & (i_3_) & (n_n94) & (x109x)));
	assign n_n1286 = (((i_5_) & (i_3_) & (!i_4_) & (n_n58) & (n_n94)));
	assign x278x = (((!i_7_) & (!i_6_) & (!n_n74) & (!n_n90) & (n_n1286)) + ((i_7_) & (!i_6_) & (n_n74) & (n_n90) & (!n_n1286)));
	assign n_n1047 = (((i_5_) & (i_3_) & (i_4_) & (n_n63) & (n_n90)));
	assign n_n1042 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n92) & (n_n94)));
	assign n_n937 = (((!i_1_) & (!i_2_) & (!i_0_)));
	assign x189x = (((!i_5_) & (!i_6_) & (!i_4_) & (!x351x) & (n_n937)) + ((!i_5_) & (!i_6_) & (!i_4_) & (x351x) & (!n_n937)));
	assign n_n941 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n93) & (n_n94)));
	assign n_n1087 = (((i_5_) & (i_3_) & (i_4_) & (n_n94) & (n_n63)));
	assign x5273x = (((!n_n101) & (!n_n83) & (!n_n102) & (x1359x) & (!x217x)) + ((!n_n101) & (!n_n83) & (!n_n102) & (!x1359x) & (x217x)) + ((n_n101) & (n_n83) & (n_n102) & (!x1359x) & (!x217x)));
	assign x5274x = (((!i_2_) & (!x56x) & (!x318x) & (n_n1294) & (!x290x)) + ((!i_2_) & (!x56x) & (!x318x) & (!n_n1294) & (x290x)) + ((!i_2_) & (x56x) & (x318x) & (!n_n1294) & (!x290x)));
	assign x5306x = (((!i_6_) & (!n_n86) & (!x27x) & (x4938x) & (!x6349x)) + ((!i_6_) & (!n_n86) & (!x27x) & (!x4938x) & (!x6349x)) + ((i_6_) & (n_n86) & (x27x) & (!x4938x) & (!x6349x)));
	assign x5307x = (((x227x) & (!n_n77) & (!x207x) & (!x61x) & (!x20x)) + ((!x227x) & (!n_n77) & (x207x) & (!x61x) & (!x20x)) + ((!x227x) & (!n_n77) & (!x207x) & (x61x) & (!x20x)) + ((!x227x) & (n_n77) & (!x207x) & (!x61x) & (x20x)));
	assign x5298x = (((!n_n101) & (!x55x) & (x323x) & (!x1352x) & (!x1143x)) + ((!n_n101) & (!x55x) & (!x323x) & (x1352x) & (!x1143x)) + ((!n_n101) & (!x55x) & (!x323x) & (!x1352x) & (x1143x)) + ((n_n101) & (x55x) & (!x323x) & (!x1352x) & (!x1143x)));
	assign x5309x = (((x352x) & (!n_n1176) & (!x5283x) & (!x6346x)) + ((!x352x) & (n_n1176) & (!x5283x) & (!x6346x)) + ((!x352x) & (!n_n1176) & (x5283x) & (!x6346x)) + ((!x352x) & (!n_n1176) & (!x5283x) & (!x6346x)));
	assign x5310x = (((x333x) & (!x332x) & (!x5288x) & (!x5289x) & (!x5290x)) + ((!x333x) & (x332x) & (!x5288x) & (!x5289x) & (!x5290x)) + ((!x333x) & (!x332x) & (x5288x) & (!x5289x) & (!x5290x)) + ((!x333x) & (!x332x) & (!x5288x) & (x5289x) & (!x5290x)) + ((!x333x) & (!x332x) & (!x5288x) & (!x5289x) & (x5290x)));
	assign x6345x = (((!x71x) & (!x118x) & (!x5291x) & (!x5292x) & (!x5305x)));
	assign x234x = (((i_7_) & (!i_8_) & (!i_5_) & (i_6_) & (!i_4_)));
	assign n_n958 = (((i_1_) & (!i_2_) & (i_0_) & (n_n95) & (n_n77)));
	assign x320x = (((i_7_) & (!i_8_) & (i_5_) & (i_6_) & (!i_4_)));
	assign n_n973 = (((i_1_) & (i_2_) & (!i_0_) & (n_n74) & (n_n82)));
	assign n_n989 = (((i_5_) & (i_3_) & (i_4_) & (n_n91) & (n_n94)));
	assign n_n944 = (((!i_5_) & (i_3_) & (i_4_) & (n_n91) & (n_n97)));
	assign n_n982 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n81) & (n_n83)));
	assign n_n967 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n100) & (n_n77)));
	assign n_n1121 = (((i_5_) & (i_6_) & (i_4_) & (n_n70) & (n_n90)));
	assign n_n53 = (((!i_3_) & (i_1_) & (i_2_)));
	assign x1588x = (((!i_5_) & (!i_6_) & (i_4_) & (n_n80)));
	assign x330x = (((i_1_) & (!i_2_)));
	assign x70x = (((!i_5_) & (!i_3_) & (!n_n73) & (x1588x) & (!x330x)) + ((!i_5_) & (!i_3_) & (n_n73) & (!x1588x) & (x330x)));
	assign x83x = (((i_5_) & (i_3_) & (!i_4_) & (i_2_) & (x108x)));
	assign x1082x = (((!i_8_) & (!i_6_) & (!i_3_) & (n_n94) & (x109x)));
	assign x90x = (((!i_8_) & (!i_6_) & (!x55x) & (n_n1125)) + ((!i_8_) & (!i_6_) & (x55x) & (!n_n1125)));
	assign n_n962 = (((!i_1_) & (i_2_) & (i_0_) & (n_n78) & (n_n74)));
	assign x168x = (((!n_n64) & (!n_n52) & (!x41x) & (!x128x) & (n_n962)) + ((n_n64) & (n_n52) & (x41x) & (!x128x) & (!n_n962)) + ((n_n64) & (n_n52) & (!x41x) & (x128x) & (!n_n962)));
	assign x5338x = (((i_5_) & (i_6_) & (i_4_)));
	assign x324x = (((i_7_) & (i_8_) & (!i_5_) & (!i_6_) & (!i_4_)));
	assign x215x = (((!n_n75) & (!n_n85) & (!x5338x) & (x324x) & (n_n67)) + ((n_n75) & (n_n85) & (x5338x) & (!x324x) & (!n_n67)));
	assign x236x = (((i_7_) & (i_8_) & (!i_6_) & (x341x) & (n_n100)));
	assign n_n1118 = (((!i_7_) & (i_8_) & (i_6_) & (x54x) & (n_n90)));
	assign x262x = (((!i_7_) & (!i_8_) & (!n_n84) & (!n_n94) & (n_n1118)) + ((i_7_) & (!i_8_) & (n_n84) & (n_n94) & (!n_n1118)));
	assign x275x = (((!i_7_) & (!i_8_) & (i_6_) & (x25x) & (!x237x)) + ((i_7_) & (i_8_) & (i_6_) & (!x25x) & (x237x)));
	assign n_n952 = (((i_5_) & (i_3_) & (i_4_) & (n_n85) & (n_n82)));
	assign x145x = (((!i_3_) & (!x341x) & (!n_n78) & (!n_n94) & (n_n952)) + ((i_3_) & (x341x) & (n_n78) & (n_n94) & (!n_n952)));
	assign n_n951 = (((i_5_) & (i_3_) & (!i_4_) & (n_n83) & (n_n82)));
	assign n_n959 = (((!i_5_) & (i_3_) & (!i_4_) & (n_n91) & (n_n97)));
	assign x146x = (((!i_3_) & (!n_n91) & (!n_n100) & (!x109x) & (n_n959)) + ((i_3_) & (n_n91) & (n_n100) & (x109x) & (!n_n959)));
	assign n_n980 = (((!i_5_) & (i_3_) & (!i_4_) & (n_n83) & (n_n82)));
	assign n_n983 = (((!i_5_) & (!i_3_) & (!i_4_) & (n_n100) & (n_n95)));
	assign n_n986 = (((i_5_) & (i_3_) & (!i_4_) & (n_n94) & (n_n63)));
	assign x5384x = (((!i_3_) & (!n_n64) & (x292x) & (!x238x) & (!x313x)) + ((!i_3_) & (n_n64) & (!x292x) & (x238x) & (!x313x)) + ((i_3_) & (!n_n64) & (!x292x) & (!x238x) & (x313x)));
	assign n_n1001 = (((!i_7_) & (i_8_) & (!i_6_) & (x57x)));
	assign n_n1004 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n91) & (n_n97)));
	assign x223x = (((!i_7_) & (!i_8_) & (n_n969) & (!n_n66) & (!n_n67)) + ((i_7_) & (!i_8_) & (!n_n969) & (n_n66) & (n_n67)));
	assign x5383x = (((!n_n82) & (!x237x) & (n_n976) & (!n_n987) & (!n_n994)) + ((!n_n82) & (!x237x) & (!n_n976) & (n_n987) & (!n_n994)) + ((!n_n82) & (!x237x) & (!n_n976) & (!n_n987) & (n_n994)) + ((n_n82) & (x237x) & (!n_n976) & (!n_n987) & (!n_n994)));
	assign x5386x = (((x275x) & (!x59x) & (!x163x) & (!x200x)) + ((!x275x) & (x59x) & (!x163x) & (!x200x)) + ((!x275x) & (!x59x) & (x163x) & (!x200x)) + ((!x275x) & (!x59x) & (!x163x) & (x200x)));
	assign n_n953 = (((!i_7_) & (!i_8_) & (!i_6_) & (n_n80) & (x110x)));
	assign n_n652 = (((!n_n103) & (!n_n102) & (!n_n97) & (!n_n95) & (n_n949)) + ((n_n103) & (n_n102) & (!n_n97) & (n_n95) & (!n_n949)) + ((!n_n103) & (n_n102) & (n_n97) & (n_n95) & (!n_n949)));
	assign x303x = (((!n_n73) & (!x53x) & (n_n967) & (!n_n966) & (!x1017x)) + ((!n_n73) & (!x53x) & (!n_n967) & (n_n966) & (!x1017x)) + ((!n_n73) & (!x53x) & (!n_n967) & (!n_n966) & (x1017x)) + ((n_n73) & (x53x) & (!n_n967) & (!n_n966) & (!x1017x)));
	assign x5393x = (((n_n951) & (!n_n954) & (!n_n952) & (!x5392x)) + ((!n_n951) & (n_n954) & (!n_n952) & (!x5392x)) + ((!n_n951) & (!n_n954) & (n_n952) & (!x5392x)) + ((!n_n951) & (!n_n954) & (!n_n952) & (x5392x)));
	assign x5400x = (((!n_n91) & (!n_n102) & (!n_n97) & (n_n939) & (!x5399x)) + ((!n_n91) & (!n_n102) & (!n_n97) & (!n_n939) & (x5399x)) + ((n_n91) & (n_n102) & (n_n97) & (!n_n939) & (!x5399x)));
	assign n_n1045 = (((i_8_) & (!i_6_) & (i_3_) & (n_n94) & (x110x)));
	assign n_n1043 = (((!i_5_) & (i_3_) & (i_4_) & (n_n91) & (n_n85)));
	assign x290x = (((!x27x) & (!n_n74) & (!n_n82) & (!x31x) & (x1153x)) + ((x27x) & (!n_n74) & (n_n82) & (!x31x) & (!x1153x)) + ((!x27x) & (n_n74) & (!n_n82) & (x31x) & (!x1153x)));
	assign x309x = (((!n_n93) & (!n_n103) & (!n_n74) & (x352x) & (!x5407x)) + ((!n_n93) & (!n_n103) & (!n_n74) & (!x352x) & (x5407x)) + ((n_n93) & (n_n103) & (n_n74) & (!x352x) & (!x5407x)));
	assign x5417x = (((!n_n92) & (!x32x) & (!n_n77) & (!x31x) & (x289x)) + ((n_n92) & (x32x) & (!n_n77) & (!x31x) & (!x289x)) + ((!n_n92) & (!x32x) & (n_n77) & (x31x) & (!x289x)));
	assign x5421x = (((x290x) & (!x309x) & (!x5417x)) + ((!x290x) & (x309x) & (!x5417x)) + ((!x290x) & (!x309x) & (x5417x)));
	assign x5413x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x27x) & (x208x)) + ((!i_7_) & (!i_8_) & (i_6_) & (x27x) & (!x208x)));
	assign x5414x = (((!n_n58) & (!x26x) & (!x32x) & (!n_n102) & (x210x)) + ((n_n58) & (x26x) & (!x32x) & (!n_n102) & (!x210x)) + ((!n_n58) & (!x26x) & (x32x) & (n_n102) & (!x210x)));
	assign x5415x = (((!n_n101) & (n_n1281) & (!x346x) & (!x63x) & (!x248x)) + ((!n_n101) & (!n_n1281) & (x346x) & (!x63x) & (!x248x)) + ((!n_n101) & (!n_n1281) & (!x346x) & (!x63x) & (x248x)) + ((n_n101) & (!n_n1281) & (!x346x) & (x63x) & (!x248x)));
	assign x5416x = (((!n_n64) & (!n_n52) & (!x57x) & (x326x) & (!x5411x)) + ((!n_n64) & (!n_n52) & (!x57x) & (!x326x) & (x5411x)) + ((n_n64) & (n_n52) & (x57x) & (!x326x) & (!x5411x)));
	assign x5422x = (((x5413x) & (!x5414x) & (!x5415x) & (!x5416x)) + ((!x5413x) & (x5414x) & (!x5415x) & (!x5416x)) + ((!x5413x) & (!x5414x) & (x5415x) & (!x5416x)) + ((!x5413x) & (!x5414x) & (!x5415x) & (x5416x)));
	assign x22x = (((i_3_) & (i_1_) & (i_2_) & (!i_0_) & (x110x)));
	assign x158x = (((!i_5_) & (n_n91) & (x67x) & (!x28x) & (!x62x)) + ((i_5_) & (!n_n91) & (!x67x) & (x28x) & (x62x)));
	assign x5436x = (((!n_n58) & (!n_n78) & (!x23x) & (!x33x) & (x5429x)) + ((!n_n58) & (n_n78) & (x23x) & (!x33x) & (!x5429x)) + ((n_n58) & (!n_n78) & (!x23x) & (x33x) & (!x5429x)));
	assign x5440x = (((!n_n101) & (!x22x) & (x158x) & (!x304x) & (!x5436x)) + ((!n_n101) & (!x22x) & (!x158x) & (x304x) & (!x5436x)) + ((!n_n101) & (!x22x) & (!x158x) & (!x304x) & (x5436x)) + ((n_n101) & (x22x) & (!x158x) & (!x304x) & (!x5436x)));
	assign x5432x = (((!n_n38) & (!n_n70) & (!x34x) & (x119x) & (!x1519x)) + ((!n_n38) & (!n_n70) & (!x34x) & (!x119x) & (x1519x)) + ((n_n38) & (n_n70) & (x34x) & (!x119x) & (!x1519x)));
	assign x5433x = (((!i_6_) & (!n_n86) & (!x57x) & (n_n1177) & (!x122x)) + ((!i_6_) & (!n_n86) & (!x57x) & (!n_n1177) & (x122x)) + ((i_6_) & (n_n86) & (x57x) & (!n_n1177) & (!x122x)));
	assign x5434x = (((!n_n93) & (!x26x) & (x329x) & (!n_n1176) & (!x22x)) + ((!n_n93) & (!x26x) & (!x329x) & (n_n1176) & (!x22x)) + ((n_n93) & (x26x) & (!x329x) & (!n_n1176) & (!x22x)) + ((n_n93) & (!x26x) & (!x329x) & (!n_n1176) & (x22x)));
	assign x5435x = (((!n_n78) & (!x55x) & (!x22x) & (x332x) & (!n_n1170)) + ((!n_n78) & (!x55x) & (!x22x) & (!x332x) & (n_n1170)) + ((n_n78) & (x55x) & (!x22x) & (!x332x) & (!n_n1170)) + ((n_n78) & (!x55x) & (x22x) & (!x332x) & (!n_n1170)));
	assign x5441x = (((x5432x) & (!x5433x) & (!x5434x) & (!x5435x)) + ((!x5432x) & (x5433x) & (!x5434x) & (!x5435x)) + ((!x5432x) & (!x5433x) & (x5434x) & (!x5435x)) + ((!x5432x) & (!x5433x) & (!x5434x) & (x5435x)));
	assign n_n1030 = (((i_5_) & (i_3_) & (i_4_) & (n_n83) & (n_n82)));
	assign x66x = (((i_7_) & (i_8_) & (i_1_) & (i_2_) & (!i_0_)));
	assign x5442x = (((i_6_) & (i_3_) & (!i_4_)));
	assign n_n1101 = (((i_7_) & (!i_8_) & (!i_6_) & (x109x) & (x322x)));
	assign x6359x = (((i_5_) & (!n_n101) & (!x58x) & (!n_n82) & (!x353x)) + ((!i_5_) & (!n_n101) & (!x58x) & (!n_n82) & (!x353x)) + ((i_5_) & (!n_n101) & (!x58x) & (!n_n82) & (!x353x)) + ((!i_5_) & (!n_n101) & (!x58x) & (!n_n82) & (!x353x)) + ((!i_5_) & (!n_n101) & (!x58x) & (!n_n82) & (!x353x)) + ((!i_5_) & (!n_n101) & (!x58x) & (!n_n82) & (!x353x)));
	assign x5450x = (((!n_n63) & (n_n1128) & (!x44x) & (!n_n1156) & (!x6359x)) + ((!n_n63) & (!n_n1128) & (!x44x) & (n_n1156) & (!x6359x)) + ((!n_n63) & (!n_n1128) & (!x44x) & (!n_n1156) & (!x6359x)) + ((n_n63) & (!n_n1128) & (x44x) & (!n_n1156) & (!x6359x)));
	assign n_n1059 = (((!i_7_) & (!i_8_) & (i_0_) & (n_n71) & (x30x)));
	assign x156x = (((!i_8_) & (!i_1_) & (!x56x) & (!n_n40) & (n_n1060)) + ((i_8_) & (!i_1_) & (x56x) & (n_n40) & (!n_n1060)));
	assign x5454x = (((!n_n38) & (n_n1058) & (!n_n1059) & (!x22x) & (!x156x)) + ((!n_n38) & (!n_n1058) & (n_n1059) & (!x22x) & (!x156x)) + ((!n_n38) & (!n_n1058) & (!n_n1059) & (!x22x) & (x156x)) + ((n_n38) & (!n_n1058) & (!n_n1059) & (x22x) & (!x156x)));
	assign x334x = (((!i_7_) & (!i_8_) & (!i_6_) & (x76x)));
	assign x142x = (((!i_6_) & (!n_n70) & (!x110x) & (!n_n53) & (x334x)) + ((!i_6_) & (n_n70) & (x110x) & (n_n53) & (!x334x)));
	assign x944x = (((!i_7_) & (i_8_) & (!i_6_) & (x42x)));
	assign x150x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x42x) & (n_n1105)) + ((!i_7_) & (i_8_) & (!i_6_) & (x42x) & (!n_n1105)));
	assign n_n1046 = (((!i_5_) & (i_3_) & (i_4_) & (n_n101) & (n_n90)));
	assign n_n1095 = (((i_5_) & (i_3_) & (!i_4_) & (n_n91) & (n_n103)));
	assign x85x = (((!i_7_) & (i_8_) & (!i_3_) & (!i_1_) & (i_0_)));
	assign x282x = (((!i_6_) & (x55x) & (n_n95) & (!x110x) & (!x85x)) + ((i_6_) & (!x55x) & (!n_n95) & (x110x) & (x85x)));
	assign x285x = (((!i_5_) & (!n_n91) & (!n_n100) & (!x54x) & (n_n1074)) + ((!i_5_) & (n_n91) & (n_n100) & (x54x) & (!n_n1074)));
	assign n_n1060 = (((i_1_) & (i_2_) & (!i_0_) & (n_n74) & (n_n63)));
	assign n_n1100 = (((i_5_) & (!i_3_) & (i_4_) & (n_n100) & (n_n82)));
	assign x132x = (((!i_7_) & (!i_8_) & (i_6_) & (i_0_) & (x75x)));
	assign n_n969 = (((i_5_) & (!i_3_) & (i_4_) & (n_n93) & (n_n83)));
	assign n_n954 = (((i_5_) & (i_3_) & (i_4_) & (n_n78) & (n_n94)));
	assign x331x = (((!i_8_) & (!i_6_)));
	assign n_n939 = (((!i_5_) & (!i_3_) & (!i_4_) & (n_n100) & (x331x)));
	assign x5068x = (((!i_7_) & (!i_8_) & (!i_1_) & (!i_2_) & (i_0_)));
	assign n_n971 = (((!i_6_) & (!i_3_) & (!i_4_) & (n_n86) & (n_n100)));
	assign n_n1037 = (((!i_8_) & (i_6_) & (i_3_) & (n_n94) & (x325x)));
	assign x903x = (((!i_5_) & (!i_6_) & (i_4_) & (n_n64) & (n_n103)));
	assign x5492x = (((!i_7_) & (!i_8_) & (!i_6_) & (x76x) & (!x21x)) + ((i_7_) & (i_8_) & (i_6_) & (!x76x) & (x21x)));
	assign x119x = (((n_n38) & (n_n64) & (x27x) & (!n_n71) & (!x242x)) + ((!n_n38) & (n_n64) & (!x27x) & (n_n71) & (x242x)));
	assign x160x = (((!i_7_) & (!i_8_) & (i_6_) & (x237x) & (!x33x)) + ((i_7_) & (i_8_) & (!i_6_) & (!x237x) & (x33x)));
	assign x5524x = (((!i_6_) & (!n_n86) & (!x25x) & (x267x) & (!x877x)) + ((!i_6_) & (!n_n86) & (!x25x) & (!x267x) & (x877x)) + ((i_6_) & (n_n86) & (x25x) & (!x267x) & (!x877x)));
	assign x5532x = (((!n_n81) & (!x32x) & (x278x) & (!x159x) & (!x5514x)) + ((!n_n81) & (!x32x) & (!x278x) & (x159x) & (!x5514x)) + ((!n_n81) & (!x32x) & (!x278x) & (!x159x) & (x5514x)) + ((n_n81) & (x32x) & (!x278x) & (!x159x) & (!x5514x)));
	assign x5536x = (((!n_n101) & (!x49x) & (x835x) & (!x5519x) & (!x5531x)) + ((!n_n101) & (!x49x) & (!x835x) & (x5519x) & (!x5531x)) + ((!n_n101) & (!x49x) & (!x835x) & (!x5519x) & (x5531x)) + ((n_n101) & (x49x) & (!x835x) & (!x5519x) & (!x5531x)));
	assign n_n947 = (((!i_3_) & (i_1_) & (!i_0_) & (n_n86) & (n_n87)));
	assign x162x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x29x) & (n_n947)) + ((i_7_) & (i_8_) & (i_6_) & (x29x) & (!n_n947)));
	assign x829x = (((!i_8_) & (i_6_) & (i_3_) & (!i_4_) & (n_n97)));
	assign x5550x = (((!n_n92) & (!n_n94) & (!n_n63) & (n_n983) & (!x212x)) + ((!n_n92) & (!n_n94) & (!n_n63) & (!n_n983) & (x212x)) + ((n_n92) & (n_n94) & (n_n63) & (!n_n983) & (!x212x)));
	assign x5551x = (((!n_n82) & (!x237x) & (n_n994) & (!n_n1013) & (!n_n978)) + ((!n_n82) & (!x237x) & (!n_n994) & (n_n1013) & (!n_n978)) + ((!n_n82) & (!x237x) & (!n_n994) & (!n_n1013) & (n_n978)) + ((n_n82) & (x237x) & (!n_n994) & (!n_n1013) & (!n_n978)));
	assign x5552x = (((!n_n86) & (!n_n85) & (!n_n76) & (n_n882) & (!n_n1026)) + ((!n_n86) & (!n_n85) & (!n_n76) & (!n_n882) & (n_n1026)) + ((n_n86) & (n_n85) & (n_n76) & (!n_n882) & (!n_n1026)));
	assign x5553x = (((n_n987) & (!n_n984) & (!n_n1011) & (!x59x) & (!x202x)) + ((!n_n987) & (n_n984) & (!n_n1011) & (!x59x) & (!x202x)) + ((!n_n987) & (!n_n984) & (n_n1011) & (!x59x) & (!x202x)) + ((!n_n987) & (!n_n984) & (!n_n1011) & (x59x) & (!x202x)) + ((!n_n987) & (!n_n984) & (!n_n1011) & (!x59x) & (x202x)));
	assign x5554x = (((!n_n71) & (x270x) & (!x85x) & (!x200x) & (!x152x)) + ((!n_n71) & (!x270x) & (!x85x) & (x200x) & (!x152x)) + ((!n_n71) & (!x270x) & (!x85x) & (!x200x) & (x152x)) + ((n_n71) & (!x270x) & (x85x) & (!x200x) & (!x152x)));
	assign n_n71 = (((!i_5_) & (i_6_) & (!i_4_)));
	assign x30x = (((i_3_) & (i_2_)));
	assign x68x = (((!i_2_) & (!n_n70) & (x38x) & (x108x) & (!n_n87)) + ((i_2_) & (n_n70) & (!x38x) & (x108x) & (n_n87)));
	assign x138x = (((!n_n91) & (!x54x) & (!x108x) & (n_n87) & (x85x)) + ((n_n91) & (x54x) & (x108x) & (!n_n87) & (!x85x)));
	assign x805x = (((i_7_) & (!i_8_) & (!i_6_) & (n_n102) & (n_n97)));
	assign x153x = (((!i_2_) & (!n_n95) & (!n_n77) & (!x108x) & (n_n953)) + ((!i_2_) & (n_n95) & (n_n77) & (x108x) & (!n_n953)));
	assign x263x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x55x) & (n_n1052)) + ((i_7_) & (i_8_) & (!i_6_) & (x55x) & (!n_n1052)));
	assign n_n975 = (((!i_5_) & (i_3_) & (!i_4_) & (n_n101) & (n_n83)));
	assign n_n1184 = (((i_7_) & (i_8_) & (i_6_) & (n_n84) & (n_n94)));
	assign x5493x = (((i_7_) & (!i_8_) & (!i_6_) & (i_3_) & (i_4_)));
	assign x224x = (((n_n93) & (n_n84) & (!n_n102) & (n_n94) & (!n_n85)) + ((n_n93) & (!n_n84) & (n_n102) & (!n_n94) & (n_n85)));
	assign x1384x = (((i_8_) & (!i_6_) & (i_3_) & (x341x) & (n_n85)));
	assign x5599x = (((!n_n91) & (!n_n100) & (!n_n102) & (x122x) & (!x1008x)) + ((!n_n91) & (!n_n100) & (!n_n102) & (!x122x) & (x1008x)) + ((n_n91) & (n_n100) & (n_n102) & (!x122x) & (!x1008x)));
	assign x5600x = (((!n_n78) & (x252x) & (!x43x) & (!x49x) & (!x348x)) + ((!n_n78) & (!x252x) & (!x43x) & (!x49x) & (x348x)) + ((n_n78) & (!x252x) & (x43x) & (!x49x) & (!x348x)) + ((n_n78) & (!x252x) & (!x43x) & (x49x) & (!x348x)));
	assign x5601x = (((!n_n63) & (!x41x) & (!x234x) & (!x242x) & (x5595x)) + ((n_n63) & (x41x) & (!x234x) & (!x242x) & (!x5595x)) + ((!n_n63) & (!x41x) & (x234x) & (x242x) & (!x5595x)));
	assign x5602x = (((n_n1297) & (!n_n1283) & (!n_n1312) & (!x309x) & (!x326x)) + ((!n_n1297) & (n_n1283) & (!n_n1312) & (!x309x) & (!x326x)) + ((!n_n1297) & (!n_n1283) & (n_n1312) & (!x309x) & (!x326x)) + ((!n_n1297) & (!n_n1283) & (!n_n1312) & (x309x) & (!x326x)) + ((!n_n1297) & (!n_n1283) & (!n_n1312) & (!x309x) & (x326x)));
	assign x5603x = (((!n_n86) & (x104x) & (!x21x) & (!x123x) & (!x217x)) + ((!n_n86) & (!x104x) & (!x21x) & (x123x) & (!x217x)) + ((!n_n86) & (!x104x) & (!x21x) & (!x123x) & (x217x)) + ((n_n86) & (!x104x) & (x21x) & (!x123x) & (!x217x)));
	assign x65x = (((i_5_) & (i_3_) & (i_4_) & (n_n100)));
	assign x869x = (((!i_5_) & (i_3_) & (i_4_) & (n_n82) & (n_n90)));
	assign n_n211 = (((!n_n58) & (!n_n95) & (!x128x) & (!x65x) & (x869x)) + ((n_n58) & (!n_n95) & (x128x) & (!x65x) & (!x869x)) + ((!n_n58) & (n_n95) & (!x128x) & (x65x) & (!x869x)));
	assign x120x = (((!x172x) & (n_n63) & (!n_n85) & (x83x) & (!x28x)) + ((x172x) & (!n_n63) & (n_n85) & (!x83x) & (x28x)));
	assign n_n1163 = (((!i_5_) & (i_3_) & (!i_4_) & (n_n91) & (n_n83)));
	assign n_n1160 = (((i_5_) & (i_3_) & (i_4_) & (n_n101) & (n_n83)));
	assign x1143x = (((i_7_) & (i_8_) & (!i_6_) & (n_n100) & (n_n84)));
	assign n_n1216 = (((!i_5_) & (!i_3_) & (i_4_) & (n_n101) & (n_n100)));
	assign n_n1158 = (((!i_7_) & (!i_8_) & (!i_6_) & (x63x)));
	assign n_n1146 = (((i_5_) & (!i_3_) & (!i_4_) & (n_n101) & (n_n85)));
	assign n_n981 = (((i_7_) & (i_8_) & (i_6_) & (n_n84) & (n_n85)));
	assign x617x = (((i_3_) & (!i_4_) & (!i_1_) & (i_0_) & (n_n93)));
	assign x5717x = (((n_n74) & (!n_n70) & (n_n63) & (n_n85) & (!n_n40)) + ((!n_n74) & (n_n70) & (!n_n63) & (n_n85) & (n_n40)));
	assign x5726x = (((!i_3_) & (!x341x) & (!x37x) & (x139x) & (!x6353x)) + ((!i_3_) & (!x341x) & (!x37x) & (!x139x) & (!x6353x)) + ((i_3_) & (x341x) & (x37x) & (!x139x) & (!x6353x)));
	assign x5729x = (((!n_n91) & (!x22x) & (n_n1181) & (!x5715x) & (!x6336x)) + ((!n_n91) & (!x22x) & (!n_n1181) & (x5715x) & (!x6336x)) + ((!n_n91) & (!x22x) & (!n_n1181) & (!x5715x) & (!x6336x)) + ((n_n91) & (x22x) & (!n_n1181) & (!x5715x) & (!x6336x)));
	assign x5743x = (((!n_n95) & (n_n1022) & (!x237x) & (!n_n1021) & (!n_n994)) + ((!n_n95) & (!n_n1022) & (!x237x) & (n_n1021) & (!n_n994)) + ((!n_n95) & (!n_n1022) & (!x237x) & (!n_n1021) & (n_n994)) + ((n_n95) & (!n_n1022) & (x237x) & (!n_n1021) & (!n_n994)));
	assign x5744x = (((!i_3_) & (n_n1010) & (!n_n1006) & (!x313x) & (!n_n1002)) + ((!i_3_) & (!n_n1010) & (n_n1006) & (!x313x) & (!n_n1002)) + ((!i_3_) & (!n_n1010) & (!n_n1006) & (!x313x) & (n_n1002)) + ((i_3_) & (!n_n1010) & (!n_n1006) & (x313x) & (!n_n1002)));
	assign x5746x = (((n_n987) & (!n_n984) & (!x152x) & (!x151x) & (!x202x)) + ((!n_n987) & (n_n984) & (!x152x) & (!x151x) & (!x202x)) + ((!n_n987) & (!n_n984) & (x152x) & (!x151x) & (!x202x)) + ((!n_n987) & (!n_n984) & (!x152x) & (x151x) & (!x202x)) + ((!n_n987) & (!n_n984) & (!x152x) & (!x151x) & (x202x)));
	assign x6339x = (((!x188x) & (!x114x) & (!n_n296) & (!x98x) & (!x280x)));
	assign n_n966 = (((!i_5_) & (i_3_) & (i_4_) & (n_n101) & (n_n97)));
	assign x1017x = (((i_8_) & (i_6_) & (i_2_) & (n_n77) & (x175x)));
	assign x5392x = (((!n_n91) & (!n_n92) & (!n_n100) & (n_n76) & (x129x)) + ((n_n91) & (n_n92) & (n_n100) & (!n_n76) & (!x129x)));
	assign x79x = (((!i_2_) & (!n_n101) & (!n_n102) & (n_n942) & (!x175x)) + ((i_2_) & (n_n101) & (n_n102) & (!n_n942) & (x175x)));
	assign x91x = (((!i_7_) & (!i_8_) & (!n_n40) & (n_n1057) & (!n_n53)) + ((i_7_) & (i_8_) & (n_n40) & (!n_n1057) & (n_n53)));
	assign x103x = (((!i_3_) & (!i_1_) & (!i_2_) & (i_0_) & (x320x)) + ((!i_3_) & (!i_1_) & (i_2_) & (i_0_) & (x320x)));
	assign x161x = (((!i_3_) & (!n_n91) & (!n_n85) & (!x110x) & (n_n1108)) + ((i_3_) & (n_n91) & (n_n85) & (x110x) & (!n_n1108)));
	assign x266x = (((!i_6_) & (!x341x) & (n_n95) & (x34x) & (!x85x)) + ((!i_6_) & (x341x) & (!n_n95) & (!x34x) & (x85x)));
	assign x268x = (((!i_7_) & (!i_8_) & (!i_6_) & (n_n1120) & (!x128x)) + ((i_7_) & (!i_8_) & (i_6_) & (!n_n1120) & (x128x)));
	assign n_n1177 = (((i_5_) & (i_3_) & (!i_4_) & (n_n78) & (n_n94)));
	assign x218x = (((!i_7_) & (!i_8_) & (!n_n97) & (!x127x) & (n_n1121)) + ((i_7_) & (!i_8_) & (n_n97) & (x127x) & (!n_n1121)));
	assign x5826x = (((!n_n103) & (!n_n82) & (!n_n77) & (!x107x) & (x218x)) + ((!n_n103) & (!n_n82) & (n_n77) & (x107x) & (!x218x)) + ((n_n103) & (n_n82) & (n_n77) & (!x107x) & (!x218x)));
	assign x526x = (((!i_6_) & (!i_1_) & (i_0_) & (n_n58) & (x109x)));
	assign x5827x = (((!n_n63) & (n_n1153) & (!x19x) & (!x90x) & (!x526x)) + ((!n_n63) & (!n_n1153) & (!x19x) & (x90x) & (!x526x)) + ((!n_n63) & (!n_n1153) & (!x19x) & (!x90x) & (x526x)) + ((n_n63) & (!n_n1153) & (x19x) & (!x90x) & (!x526x)));
	assign x5841x = (((!n_n64) & (!n_n52) & (!x34x) & (n_n1047) & (!x5835x)) + ((!n_n64) & (!n_n52) & (!x34x) & (!n_n1047) & (x5835x)) + ((n_n64) & (n_n52) & (x34x) & (!n_n1047) & (!x5835x)));
	assign x5842x = (((n_n1105) & (!x944x) & (!x285x) & (!x903x) & (!x5492x)) + ((!n_n1105) & (x944x) & (!x285x) & (!x903x) & (!x5492x)) + ((!n_n1105) & (!x944x) & (x285x) & (!x903x) & (!x5492x)) + ((!n_n1105) & (!x944x) & (!x285x) & (x903x) & (!x5492x)) + ((!n_n1105) & (!x944x) & (!x285x) & (!x903x) & (x5492x)));
	assign x5844x = (((n_n1109) & (!n_n1095) & (!x355x) & (!n_n1088) & (!x6335x)) + ((!n_n1109) & (n_n1095) & (!x355x) & (!n_n1088) & (!x6335x)) + ((!n_n1109) & (!n_n1095) & (x355x) & (!n_n1088) & (!x6335x)) + ((!n_n1109) & (!n_n1095) & (!x355x) & (n_n1088) & (!x6335x)) + ((!n_n1109) & (!n_n1095) & (!x355x) & (!n_n1088) & (!x6335x)));
	assign x6334x = (((!n_n1087) & (!x805x) & (!x263x) & (!x161x) & (!x102x)));
	assign x238x = (((!i_5_) & (!i_3_) & (i_4_) & (!i_2_) & (x108x)));
	assign x92x = (((!i_7_) & (!i_8_) & (!i_6_) & (n_n1169) & (!x238x)) + ((!i_7_) & (i_8_) & (!i_6_) & (!n_n1169) & (x238x)));
	assign x159x = (((!n_n81) & (!n_n101) & (!n_n103) & (x38x) & (x322x)) + ((n_n81) & (n_n101) & (n_n103) & (!x38x) & (!x322x)));
	assign x247x = (((!i_7_) & (!i_8_) & (i_1_) & (i_2_) & (!i_0_)));
	assign x316x = (((i_7_) & (i_8_) & (!i_1_) & (i_2_) & (!i_0_)));
	assign x335x = (((i_7_) & (!i_8_) & (!i_6_) & (n_n81) & (n_n97)));
	assign x344x = (((!i_7_) & (!i_8_) & (i_6_) & (n_n103) & (n_n84)));
	assign x5886x = (((!n_n73) & (!x26x) & (!n_n102) & (n_n1085) & (!x20x)) + ((n_n73) & (x26x) & (!n_n102) & (!n_n1085) & (!x20x)) + ((!n_n73) & (!x26x) & (n_n102) & (!n_n1085) & (x20x)));
	assign x5892x = (((!n_n94) & (x334x) & (!n_n1105) & (!n_n1108) & (!x5085x)) + ((!n_n94) & (!x334x) & (n_n1105) & (!n_n1108) & (!x5085x)) + ((!n_n94) & (!x334x) & (!n_n1105) & (n_n1108) & (!x5085x)) + ((n_n94) & (!x334x) & (!n_n1105) & (!n_n1108) & (x5085x)));
	assign n_n1014 = (((i_5_) & (i_3_) & (i_4_) & (n_n78) & (n_n100)));
	assign x152x = (((!i_6_) & (!n_n64) & (!n_n85) & (!x325x) & (x827x)) + ((i_6_) & (n_n64) & (n_n85) & (x325x) & (!x827x)));
	assign n_n1018 = (((i_5_) & (!i_3_) & (i_4_) & (n_n100) & (n_n95)));
	assign x5889x = (((!n_n91) & (!x27x) & (n_n1074) & (!n_n1045) & (!n_n1060)) + ((!n_n91) & (!x27x) & (!n_n1074) & (n_n1045) & (!n_n1060)) + ((!n_n91) & (!x27x) & (!n_n1074) & (!n_n1045) & (n_n1060)) + ((n_n91) & (x27x) & (!n_n1074) & (!n_n1045) & (!n_n1060)));
	assign x5895x = (((n_n1146) & (!n_n1010) & (!x5880x) & (!x5881x) & (!x5882x)) + ((!n_n1146) & (n_n1010) & (!x5880x) & (!x5881x) & (!x5882x)) + ((!n_n1146) & (!n_n1010) & (x5880x) & (!x5881x) & (!x5882x)) + ((!n_n1146) & (!n_n1010) & (!x5880x) & (x5881x) & (!x5882x)) + ((!n_n1146) & (!n_n1010) & (!x5880x) & (!x5881x) & (x5882x)));
	assign n_n999 = (((!i_7_) & (!i_8_) & (i_6_) & (x63x)));
	assign x615x = (((!i_7_) & (i_5_) & (!i_6_) & (!i_3_) & (n_n83)));
	assign x5901x = (((!n_n95) & (!x44x) & (n_n980) & (!n_n999) & (!x615x)) + ((!n_n95) & (!x44x) & (!n_n980) & (n_n999) & (!x615x)) + ((!n_n95) & (!x44x) & (!n_n980) & (!n_n999) & (x615x)) + ((n_n95) & (x44x) & (!n_n980) & (!n_n999) & (!x615x)));
	assign x5904x = (((!n_n95) & (!x29x) & (x829x) & (!x125x) & (!n_n947)) + ((!n_n95) & (!x29x) & (!x829x) & (x125x) & (!n_n947)) + ((!n_n95) & (!x29x) & (!x829x) & (!x125x) & (n_n947)) + ((n_n95) & (x29x) & (!x829x) & (!x125x) & (!n_n947)));
	assign x129x = (((!i_7_) & (i_8_) & (i_1_) & (!i_2_) & (i_0_)));
	assign x877x = (((i_7_) & (!i_8_) & (!i_6_) & (x21x)));
	assign x5907x = (((!n_n93) & (!x57x) & (!x25x) & (n_n1177) & (!x877x)) + ((!n_n93) & (!x57x) & (!x25x) & (!n_n1177) & (x877x)) + ((n_n93) & (x57x) & (!x25x) & (!n_n1177) & (!x877x)) + ((n_n93) & (!x57x) & (x25x) & (!n_n1177) & (!x877x)));
	assign x6361x = (((n_n52) & (!n_n78) & (x34x) & (!x52x) & (!x22x)) + ((!n_n52) & (n_n78) & (!x34x) & (x52x) & (!x22x)) + ((!n_n52) & (n_n78) & (!x34x) & (!x52x) & (x22x)));
	assign x5908x = (((!n_n78) & (!n_n100) & (!n_n84) & (n_n1216) & (!x6361x)) + ((!n_n78) & (!n_n100) & (!n_n84) & (!n_n1216) & (x6361x)) + ((n_n78) & (n_n100) & (n_n84) & (!n_n1216) & (!x6361x)));
	assign x155x = (((!n_n75) & (n_n81) & (!n_n100) & (!n_n40) & (x107x)) + ((n_n75) & (!n_n81) & (n_n100) & (n_n40) & (!x107x)));
	assign x332x = (((i_7_) & (i_8_) & (i_6_) & (n_n74) & (n_n90)));
	assign x157x = (((!i_7_) & (!i_8_) & (!n_n54) & (!n_n53) & (x332x)) + ((i_7_) & (!i_8_) & (n_n54) & (n_n53) & (!x332x)));
	assign x174x = (((i_3_) & (!i_1_) & (i_2_)));
	assign x210x = (((!i_7_) & (!i_8_) & (!n_n100) & (n_n1267) & (!x131x)) + ((i_7_) & (i_8_) & (n_n100) & (!n_n1267) & (x131x)));
	assign x662x = (((i_5_) & (i_3_) & (!i_4_) & (n_n78) & (n_n85)));
	assign x663x = (((i_1_) & (i_2_) & (!i_0_) & (n_n101) & (n_n77)));
	assign x336x = (((i_7_) & (i_8_) & (i_6_) & (n_n84) & (n_n97)));
	assign x33x = (((!i_5_) & (i_3_) & (!i_4_) & (i_2_) & (x108x)));
	assign x226x = (((!i_7_) & (!i_8_) & (!i_6_) & (x321x) & (!x33x)) + ((i_7_) & (i_8_) & (i_6_) & (!x321x) & (x33x)));
	assign n_n1170 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n92) & (n_n100)));
	assign x267x = (((!i_7_) & (!i_8_) & (i_6_) & (x45x) & (!x63x)) + ((!i_7_) & (i_8_) & (i_6_) & (!x45x) & (x63x)));
	assign x130x = (((!i_5_) & (!i_6_) & (!i_3_)));
	assign x5910x = (((!n_n93) & (!n_n83) & (!n_n102) & (x66x) & (x130x)) + ((n_n93) & (n_n83) & (n_n102) & (!x66x) & (!x130x)));
	assign x307x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x23x) & (x5910x)) + ((i_7_) & (i_8_) & (!i_6_) & (x23x) & (!x5910x)));
	assign x5686x = (((!i_7_) & (!i_8_) & (!i_3_)));
	assign x5687x = (((i_5_) & (!i_6_) & (i_4_) & (i_1_) & (!i_2_)));
	assign n_n1164 = (((!i_7_) & (!i_8_) & (i_6_) & (x42x)));
	assign n_n1088 = (((i_5_) & (i_3_) & (!i_4_) & (n_n91) & (n_n97)));
	assign x350x = (((i_5_) & (!i_3_) & (i_4_) & (n_n101) & (n_n100)));
	assign x5964x = (((!i_7_) & (!i_8_) & (!n_n85) & (x348x) & (!n_n40)) + ((i_7_) & (!i_8_) & (n_n85) & (!x348x) & (n_n40)));
	assign x5975x = (((!n_n78) & (x323x) & (!n_n1294) & (!n_n1283) & (!x22x)) + ((!n_n78) & (!x323x) & (n_n1294) & (!n_n1283) & (!x22x)) + ((!n_n78) & (!x323x) & (!n_n1294) & (n_n1283) & (!x22x)) + ((n_n78) & (!x323x) & (!n_n1294) & (!n_n1283) & (x22x)));
	assign x5984x = (((x5965x) & (!x5966x) & (!x5967x) & (!x5968x)) + ((!x5965x) & (x5966x) & (!x5967x) & (!x5968x)) + ((!x5965x) & (!x5966x) & (x5967x) & (!x5968x)) + ((!x5965x) & (!x5966x) & (!x5967x) & (x5968x)));
	assign x163x = (((i_2_) & (n_n84) & (n_n70) & (!n_n95) & (x108x)) + ((!i_2_) & (n_n84) & (!n_n70) & (n_n95) & (x108x)));
	assign n_n978 = (((i_5_) & (i_3_) & (!i_4_) & (n_n83) & (n_n63)));
	assign x5990x = (((!n_n91) & (!n_n103) & (!n_n102) & (x163x) & (!n_n978)) + ((!n_n91) & (!n_n103) & (!n_n102) & (!x163x) & (n_n978)) + ((n_n91) & (n_n103) & (n_n102) & (!x163x) & (!n_n978)));
	assign n_n296 = (((!n_n81) & (!n_n101) & (!n_n90) & (n_n999) & (!x615x)) + ((!n_n81) & (!n_n101) & (!n_n90) & (!n_n999) & (x615x)) + ((n_n81) & (n_n101) & (n_n90) & (!n_n999) & (!x615x)));
	assign x5991x = (((!n_n100) & (!n_n83) & (!n_n74) & (!n_n95) & (n_n296)) + ((n_n100) & (!n_n83) & (n_n74) & (n_n95) & (!n_n296)) + ((!n_n100) & (n_n83) & (n_n74) & (n_n95) & (!n_n296)));
	assign x242x = (((i_3_) & (i_2_) & (!i_0_)));
	assign x246x = (((i_1_) & (i_2_) & (!i_0_) & (n_n91) & (n_n84)));
	assign x1557x = (((i_5_) & (i_3_) & (i_4_) & (n_n101) & (n_n90)));
	assign n_n1010 = (((!i_5_) & (i_3_) & (!i_4_) & (n_n78) & (n_n97)));
	assign x270x = (((!i_7_) & (i_8_) & (!i_6_) & (x57x) & (!x33x)) + ((!i_7_) & (!i_8_) & (!i_6_) & (!x57x) & (x33x)));
	assign n_n976 = (((!i_7_) & (!i_5_) & (i_6_) & (n_n85) & (x54x)));
	assign x272x = (((!i_6_) & (!i_3_) & (!i_4_) & (!x5068x) & (n_n976)) + ((!i_6_) & (!i_3_) & (!i_4_) & (x5068x) & (!n_n976)));
	assign n_n1181 = (((!i_7_) & (!i_8_) & (!i_6_) & (x55x)));
	assign x194x = (((i_5_) & (!i_3_) & (i_4_)) + ((!i_5_) & (i_3_) & (!i_4_)));
	assign n_n987 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n102) & (n_n97)));
	assign n_n984 = (((!i_7_) & (i_8_) & (!i_6_) & (n_n103) & (n_n102)));
	assign x147x = (((!i_7_) & (!i_8_) & (i_6_) & (x29x) & (!x52x)) + ((!i_7_) & (i_8_) & (!i_6_) & (!x29x) & (x52x)));
	assign x274x = (((!i_3_) & (!x341x) & (!n_n83) & (!n_n82) & (n_n1021)) + ((i_3_) & (x341x) & (n_n83) & (n_n82) & (!n_n1021)));
	assign n_n1009 = (((i_5_) & (i_3_) & (i_4_) & (n_n103) & (n_n95)));
	assign n_n1011 = (((i_5_) & (i_6_) & (!i_3_) & (n_n64) & (n_n103)));
	assign x339x = (((!i_7_) & (i_8_) & (!i_5_) & (!i_6_) & (!i_4_)));
	assign x217x = (((!i_8_) & (!i_6_) & (n_n81) & (!x43x) & (x48x)) + ((i_8_) & (!i_6_) & (!n_n81) & (x43x) & (!x48x)));
	assign x71x = (((i_5_) & (!n_n103) & (x54x) & (!n_n82) & (x107x)) + ((i_5_) & (n_n103) & (x54x) & (n_n82) & (!x107x)));
	assign n_n994 = (((i_1_) & (i_2_) & (!i_0_) & (n_n91) & (n_n102)));
	assign n_n1006 = (((i_1_) & (!i_2_) & (!i_0_) & (n_n74) & (n_n95)));
	assign x59x = (((!i_7_) & (!i_8_) & (!n_n100) & (!n_n54) & (n_n1006)) + ((i_7_) & (!i_8_) & (n_n100) & (n_n54) & (!n_n1006)));
	assign x200x = (((!i_7_) & (!i_6_) & (!x109x) & (n_n982) & (!n_n53)) + ((i_7_) & (!i_6_) & (x109x) & (!n_n982) & (n_n53)));
	assign x313x = (((!i_1_) & (i_2_) & (i_0_) & (n_n38) & (n_n64)));
	assign x5399x = (((!i_8_) & (!i_6_) & (!n_n97) & (n_n947) & (!x312x)) + ((!i_8_) & (i_6_) & (n_n97) & (!n_n947) & (x312x)));
	assign n_n1013 = (((!i_7_) & (!i_8_) & (i_6_) & (x76x)));
	assign n_n1028 = (((i_1_) & (i_2_) & (i_0_) & (n_n63) & (n_n77)));
	assign x827x = (((i_5_) & (!i_6_) & (!i_4_) & (n_n86) & (n_n83)));
	assign x753x = (((!i_7_) & (!i_8_) & (!i_2_) & (x108x) & (n_n76)));
	assign n_n1002 = (((i_3_) & (i_2_) & (i_0_) & (x339x)));
	assign x5609x = (((!i_7_) & (!i_8_) & (!n_n74) & (!n_n85) & (n_n1002)) + ((i_7_) & (i_8_) & (n_n74) & (n_n85) & (!n_n1002)));
	assign x5616x = (((!i_6_) & (!n_n86) & (!x112x) & (n_n1001) & (!x152x)) + ((!i_6_) & (!n_n86) & (!x112x) & (!n_n1001) & (x152x)) + ((i_6_) & (n_n86) & (x112x) & (!n_n1001) & (!x152x)));
	assign x5617x = (((!x25x) & (!n_n82) & (n_n1047) & (!n_n1013) & (!n_n1014)) + ((!x25x) & (!n_n82) & (!n_n1047) & (n_n1013) & (!n_n1014)) + ((!x25x) & (!n_n82) & (!n_n1047) & (!n_n1013) & (n_n1014)) + ((x25x) & (n_n82) & (!n_n1047) & (!n_n1013) & (!n_n1014)));
	assign x5618x = (((n_n980) & (!n_n983) & (!n_n986) & (!n_n1021) & (!n_n1028)) + ((!n_n980) & (n_n983) & (!n_n986) & (!n_n1021) & (!n_n1028)) + ((!n_n980) & (!n_n983) & (n_n986) & (!n_n1021) & (!n_n1028)) + ((!n_n980) & (!n_n983) & (!n_n986) & (n_n1021) & (!n_n1028)) + ((!n_n980) & (!n_n983) & (!n_n986) & (!n_n1021) & (n_n1028)));
	assign x5619x = (((!n_n86) & (!n_n85) & (!n_n76) & (x5609x) & (!x299x)) + ((!n_n86) & (!n_n85) & (!n_n76) & (!x5609x) & (x299x)) + ((n_n86) & (n_n85) & (n_n76) & (!x5609x) & (!x299x)));
	assign x5620x = (((!n_n78) & (!x29x) & (x201x) & (!x271x) & (!x275x)) + ((!n_n78) & (!x29x) & (!x201x) & (x271x) & (!x275x)) + ((!n_n78) & (!x29x) & (!x201x) & (!x271x) & (x275x)) + ((n_n78) & (x29x) & (!x201x) & (!x271x) & (!x275x)));
	assign x345x = (((i_7_) & (i_8_) & (i_6_) & (x21x)));
	assign x249x = (((i_7_) & (i_6_) & (i_3_) & (x341x) & (n_n97)));
	assign x1583x = (((!i_7_) & (!i_8_) & (!i_5_) & (i_6_) & (n_n83)));
	assign n_n1026 = (((!i_3_) & (i_1_) & (!i_0_) & (n_n70) & (n_n71)));
	assign x4876x = (((i_7_) & (!i_8_) & (!i_6_) & (!i_4_)));
	assign x1581x = (((i_7_) & (!i_6_) & (!i_3_) & (i_4_) & (n_n85)));
	assign x288x = (((!i_1_) & (!x56x) & (n_n1026) & (!x4876x) & (!x1581x)) + ((!i_1_) & (!x56x) & (!n_n1026) & (!x4876x) & (x1581x)) + ((i_1_) & (x56x) & (!n_n1026) & (x4876x) & (!x1581x)));
	assign n_n943 = (((!i_7_) & (!i_8_) & (i_6_) & (n_n92) & (n_n90)));
	assign x202x = (((!i_2_) & (n_n81) & (n_n91) & (!n_n82) & (x175x)) + ((i_2_) & (n_n81) & (!n_n91) & (n_n82) & (x175x)));
	assign x203x = (((!i_7_) & (!i_2_) & (!x108x) & (!n_n76) & (n_n1004)) + ((!i_7_) & (i_2_) & (x108x) & (n_n76) & (!n_n1004)));
	assign x225x = (((!i_0_) & (n_n91) & (!x75x) & (!n_n77) & (x34x)) + ((i_0_) & (n_n91) & (x75x) & (n_n77) & (!x34x)));
	assign x1008x = (((!i_5_) & (!i_3_) & (!i_4_) & (n_n93) & (n_n85)));
	assign x289x = (((!n_n81) & (!n_n91) & (!x41x) & (!x20x) & (x1008x)) + ((!n_n81) & (n_n91) & (x41x) & (!x20x) & (!x1008x)) + ((n_n81) & (!n_n91) & (!x41x) & (x20x) & (!x1008x)));
	assign x1153x = (((!i_5_) & (i_3_) & (i_4_) & (n_n78) & (n_n90)));
	assign x5407x = (((!n_n93) & (n_n102) & (n_n63) & (!n_n77) & (n_n90)) + ((n_n93) & (!n_n102) & (!n_n63) & (n_n77) & (n_n90)));
	assign x98x = (((!i_3_) & (!n_n52) & (!n_n83) & (!x109x) & (n_n1009)) + ((!i_3_) & (n_n52) & (n_n83) & (x109x) & (!n_n1009)));
	assign x154x = (((!i_3_) & (!i_4_) & (!n_n38) & (!n_n103) & (n_n1043)) + ((!i_3_) & (!i_4_) & (n_n38) & (n_n103) & (!n_n1043)));
	assign x212x = (((!i_3_) & (!i_0_) & (!n_n101) & (!x75x) & (n_n1022)) + ((!i_3_) & (i_0_) & (n_n101) & (x75x) & (!n_n1022)));
	assign x280x = (((!i_8_) & (!i_6_) & (!n_n102) & (!n_n94) & (n_n1028)) + ((!i_8_) & (i_6_) & (n_n102) & (n_n94) & (!n_n1028)));
	assign x5791x = (((!n_n94) & (n_n1010) & (!x5085x) & (!x249x) & (!n_n1026)) + ((!n_n94) & (!n_n1010) & (!x5085x) & (x249x) & (!n_n1026)) + ((!n_n94) & (!n_n1010) & (!x5085x) & (!x249x) & (n_n1026)) + ((n_n94) & (!n_n1010) & (x5085x) & (!x249x) & (!n_n1026)));
	assign x5792x = (((n_n1032) & (!n_n1040) & (!x114x) & (!n_n1011) & (!x59x)) + ((!n_n1032) & (n_n1040) & (!x114x) & (!n_n1011) & (!x59x)) + ((!n_n1032) & (!n_n1040) & (x114x) & (!n_n1011) & (!x59x)) + ((!n_n1032) & (!n_n1040) & (!x114x) & (n_n1011) & (!x59x)) + ((!n_n1032) & (!n_n1040) & (!x114x) & (!n_n1011) & (x59x)));
	assign x5793x = (((n_n1046) & (!x274x) & (!x151x) & (!x1583x) & (!x98x)) + ((!n_n1046) & (x274x) & (!x151x) & (!x1583x) & (!x98x)) + ((!n_n1046) & (!x274x) & (x151x) & (!x1583x) & (!x98x)) + ((!n_n1046) & (!x274x) & (!x151x) & (x1583x) & (!x98x)) + ((!n_n1046) & (!x274x) & (!x151x) & (!x1583x) & (x98x)));
	assign x6333x = (((!n_n1045) & (!n_n1013) & (!x154x) & (!x212x) & (!x280x)));
	assign x101x = (((i_7_) & (!i_8_) & (!i_6_) & (x58x) & (!x44x)) + ((!i_7_) & (i_8_) & (!i_6_) & (!x58x) & (x44x)));
	assign x102x = (((!i_5_) & (!i_3_) & (!n_n93) & (!n_n97) & (x900x)) + ((i_5_) & (i_3_) & (n_n93) & (n_n97) & (!x900x)));
	assign x5504x = (((!n_n91) & (!n_n84) & (!n_n85) & (n_n1108) & (!x92x)) + ((!n_n91) & (!n_n84) & (!n_n85) & (!n_n1108) & (x92x)) + ((n_n91) & (n_n84) & (n_n85) & (!n_n1108) & (!x92x)));
	assign x5505x = (((!n_n86) & (!n_n97) & (!n_n77) & (n_n1128) & (!x224x)) + ((!n_n86) & (!n_n97) & (!n_n77) & (!n_n1128) & (x224x)) + ((n_n86) & (n_n97) & (n_n77) & (!n_n1128) & (!x224x)));
	assign x5507x = (((!n_n38) & (!n_n64) & (!x64x) & (n_n1132) & (!x5499x)) + ((!n_n38) & (!n_n64) & (!x64x) & (!n_n1132) & (x5499x)) + ((n_n38) & (n_n64) & (x64x) & (!n_n1132) & (!x5499x)));
	assign x876x = (((!i_7_) & (!i_8_) & (i_6_) & (n_n81) & (n_n103)));
	assign x166x = (((i_0_) & (x75x) & (n_n82) & (!n_n95) & (n_n77)) + ((!i_0_) & (x75x) & (!n_n82) & (n_n95) & (n_n77)));
	assign x220x = (((!i_7_) & (!i_8_) & (n_n74) & (x20x) & (!x65x)) + ((i_7_) & (!i_8_) & (!n_n74) & (!x20x) & (x65x)));
	assign x281x = (((!i_3_) & (!x341x) & (!n_n78) & (!n_n97) & (n_n1172)) + ((i_3_) & (x341x) & (n_n78) & (n_n97) & (!n_n1172)));
	assign x5514x = (((i_7_) & (!i_8_) & (i_6_) & (x45x) & (!x239x)) + ((!i_7_) & (i_8_) & (i_6_) & (!x45x) & (x239x)));
	assign x5699x = (((!n_n74) & (x662x) & (!x663x) & (!x31x) & (!x1153x)) + ((!n_n74) & (!x662x) & (x663x) & (!x31x) & (!x1153x)) + ((!n_n74) & (!x662x) & (!x663x) & (!x31x) & (x1153x)) + ((n_n74) & (!x662x) & (!x663x) & (x31x) & (!x1153x)));
	assign x5700x = (((!n_n91) & (!x42x) & (n_n1259) & (!x344x) & (!n_n1312)) + ((!n_n91) & (!x42x) & (!n_n1259) & (x344x) & (!n_n1312)) + ((!n_n91) & (!x42x) & (!n_n1259) & (!x344x) & (n_n1312)) + ((n_n91) & (x42x) & (!n_n1259) & (!x344x) & (!n_n1312)));
	assign x5703x = (((!n_n101) & (!n_n91) & (!x33x) & (!x65x) & (x5697x)) + ((n_n101) & (!n_n91) & (x33x) & (!x65x) & (!x5697x)) + ((!n_n101) & (n_n91) & (!x33x) & (x65x) & (!x5697x)));
	assign x5704x = (((x104x) & (!x157x) & (!x289x)) + ((!x104x) & (x157x) & (!x289x)) + ((!x104x) & (!x157x) & (x289x)));
	assign x5706x = (((x343x) & (!n_n1215) & (!x5693x) & (!x5694x) & (!x5695x)) + ((!x343x) & (n_n1215) & (!x5693x) & (!x5694x) & (!x5695x)) + ((!x343x) & (!n_n1215) & (x5693x) & (!x5694x) & (!x5695x)) + ((!x343x) & (!n_n1215) & (!x5693x) & (x5694x) & (!x5695x)) + ((!x343x) & (!n_n1215) & (!x5693x) & (!x5694x) & (x5695x)));
	assign x1508x = (((!i_7_) & (i_8_) & (i_0_) & (x75x) & (n_n66)));
	assign x121x = (((!i_5_) & (!i_3_) & (!n_n93) & (!n_n85) & (x1508x)) + ((i_5_) & (!i_3_) & (n_n93) & (n_n85) & (!x1508x)));
	assign x287x = (((!i_8_) & (!i_6_) & (!n_n92) & (!n_n97) & (x68x)) + ((!i_8_) & (i_6_) & (n_n92) & (n_n97) & (!x68x)));
	assign x122x = (((!i_3_) & (x45x) & (!x110x) & (x331x) & (!x316x)) + ((!i_3_) & (!x45x) & (x110x) & (!x331x) & (x316x)));
	assign x900x = (((i_7_) & (i_8_) & (!i_2_) & (x175x) & (n_n66)));
	assign x1440x = (((!i_5_) & (i_3_) & (!i_4_) & (n_n93) & (n_n94)));
	assign x312x = (((i_3_) & (!i_4_)));
	assign x5828x = (((i_7_) & (!i_8_) & (i_0_)));
	assign x670x = (((i_7_) & (!i_8_) & (i_6_) & (x57x)));
	assign x835x = (((i_5_) & (i_3_) & (i_4_) & (n_n94) & (n_n95)));
	assign x1085x = (((i_7_) & (i_6_) & (!i_3_) & (n_n83) & (x109x)));
	assign x1108x = (((i_5_) & (i_6_) & (i_3_) & (n_n64) & (n_n90)));
	assign x1442x = (((i_8_) & (i_5_) & (i_1_) & (n_n52) & (x56x)));
	assign x1446x = (((!i_7_) & (!i_8_) & (i_5_) & (!i_6_) & (n_n100)));
	assign x1589x = (((!i_7_) & (i_8_) & (i_6_) & (n_n81) & (x75x)));
	assign x4848x = (((!n_n81) & (!n_n52) & (x172x) & (!n_n85) & (x311x)) + ((n_n81) & (n_n52) & (!x172x) & (n_n85) & (!x311x)));
	assign x4849x = (((i_7_) & (!i_8_) & (i_6_) & (x27x) & (!x45x)) + ((!i_7_) & (i_8_) & (!i_6_) & (x27x) & (!x45x)) + ((i_7_) & (!i_8_) & (i_6_) & (!x27x) & (x45x)) + ((!i_7_) & (i_8_) & (!i_6_) & (!x27x) & (x45x)));
	assign x4852x = (((n_n101) & (!n_n78) & (!n_n74) & (!n_n97) & (x55x)) + ((!n_n101) & (n_n78) & (n_n74) & (n_n97) & (!x55x)));
	assign x4858x = (((!n_n93) & (!x57x) & (!x26x) & (x235x) & (!x329x)) + ((!n_n93) & (!x57x) & (!x26x) & (!x235x) & (x329x)) + ((n_n93) & (x57x) & (!x26x) & (!x235x) & (!x329x)) + ((n_n93) & (!x57x) & (x26x) & (!x235x) & (!x329x)));
	assign x4860x = (((!n_n52) & (!n_n93) & (!x64x) & (!x112x) & (x4849x)) + ((!n_n52) & (n_n93) & (x64x) & (!x112x) & (!x4849x)) + ((n_n52) & (!n_n93) & (!x64x) & (x112x) & (!x4849x)));
	assign x4885x = (((!n_n81) & (!n_n64) & (!n_n52) & (!n_n103) & (n_n1011)) + ((n_n81) & (n_n64) & (n_n52) & (n_n103) & (!n_n1011)));
	assign x6348x = (((!x55x) & (!n_n95) & (!n_n1043) & (!n_n1059) & (!n_n1042)) + ((!x55x) & (!n_n95) & (!n_n1043) & (!n_n1059) & (!n_n1042)));
	assign x4935x = (((n_n75) & (n_n81) & (!n_n93) & (n_n103) & (!n_n77)) + ((!n_n75) & (!n_n81) & (n_n93) & (n_n103) & (n_n77)));
	assign x4961x = (((!n_n81) & (!n_n86) & (n_n91) & (x64x) & (!x108x)) + ((n_n81) & (n_n86) & (!n_n91) & (!x64x) & (x108x)));
	assign x4967x = (((!i_1_) & (!i_2_) & (!n_n58) & (!n_n102) & (x1446x)) + ((i_1_) & (i_2_) & (n_n58) & (n_n102) & (!x1446x)));
	assign x4968x = (((!i_5_) & (!i_6_) & (x54x) & (x37x) & (!x328x)) + ((!i_5_) & (i_6_) & (x54x) & (!x37x) & (x328x)));
	assign x4969x = (((!i_3_) & (x27x) & (!n_n97) & (n_n82) & (!x325x)) + ((i_3_) & (!x27x) & (n_n97) & (n_n82) & (x325x)));
	assign x4970x = (((n_n73) & (n_n92) & (n_n103) & (!n_n82) & (!n_n77)) + ((!n_n73) & (!n_n92) & (n_n103) & (n_n82) & (n_n77)));
	assign x4971x = (((!n_n80) & (!n_n86) & (x105x) & (!x109x) & (!x1442x)) + ((!n_n80) & (!n_n86) & (!x105x) & (!x109x) & (x1442x)) + ((n_n80) & (n_n86) & (!x105x) & (x109x) & (!x1442x)));
	assign x4972x = (((!i_7_) & (!i_6_) & (n_n1082) & (!x207x) & (!x21x)) + ((!i_7_) & (!i_6_) & (!n_n1082) & (x207x) & (!x21x)) + ((!i_7_) & (!i_6_) & (!n_n1082) & (!x207x) & (x21x)));
	assign x4973x = (((!i_7_) & (!i_8_) & (x254x) & (!x53x) & (!x63x)) + ((i_7_) & (!i_8_) & (!x254x) & (x53x) & (!x63x)) + ((!i_7_) & (i_8_) & (!x254x) & (!x53x) & (x63x)));
	assign x4974x = (((!n_n81) & (!n_n95) & (n_n1078) & (!n_n90) & (!x4961x)) + ((!n_n81) & (!n_n95) & (!n_n1078) & (!n_n90) & (x4961x)) + ((n_n81) & (n_n95) & (!n_n1078) & (n_n90) & (!x4961x)));
	assign x4975x = (((!x245x) & (!x38x) & (n_n1279) & (!n_n1153) & (!n_n1297)) + ((!x245x) & (!x38x) & (!n_n1279) & (n_n1153) & (!n_n1297)) + ((!x245x) & (!x38x) & (!n_n1279) & (!n_n1153) & (n_n1297)) + ((x245x) & (x38x) & (!n_n1279) & (!n_n1153) & (!n_n1297)));
	assign x4976x = (((!n_n91) & (!x27x) & (n_n1324) & (!x251x) & (!x321x)) + ((!n_n91) & (!x27x) & (!n_n1324) & (x251x) & (!x321x)) + ((!n_n91) & (!x27x) & (!n_n1324) & (!x251x) & (x321x)) + ((n_n91) & (x27x) & (!n_n1324) & (!x251x) & (!x321x)));
	assign x4982x = (((x4967x) & (!x4968x) & (!x4969x) & (!x4970x)) + ((!x4967x) & (x4968x) & (!x4969x) & (!x4970x)) + ((!x4967x) & (!x4968x) & (x4969x) & (!x4970x)) + ((!x4967x) & (!x4968x) & (!x4969x) & (x4970x)));
	assign x5035x = (((!i_7_) & (!i_8_) & (!i_6_) & (x21x) & (!x34x)) + ((!i_7_) & (i_8_) & (!i_6_) & (!x21x) & (x34x)));
	assign x5037x = (((!n_n93) & (!n_n74) & (!n_n97) & (n_n1188) & (!x178x)) + ((!n_n93) & (!n_n74) & (!n_n97) & (!n_n1188) & (x178x)) + ((n_n93) & (n_n74) & (n_n97) & (!n_n1188) & (!x178x)));
	assign x5056x = (((!n_n38) & (!n_n70) & (!x34x) & (x354x) & (x62x)) + ((n_n38) & (n_n70) & (x34x) & (!x354x) & (!x62x)));
	assign x5059x = (((!n_n93) & (n_n1185) & (!n_n1172) & (!x19x) & (!x36x)) + ((!n_n93) & (!n_n1185) & (n_n1172) & (!x19x) & (!x36x)) + ((n_n93) & (!n_n1185) & (!n_n1172) & (x19x) & (!x36x)) + ((n_n93) & (!n_n1185) & (!n_n1172) & (!x19x) & (x36x)));
	assign x5087x = (((i_7_) & (i_8_) & (!i_6_) & (x64x) & (!x53x)) + ((i_7_) & (i_8_) & (!i_6_) & (!x64x) & (x53x)));
	assign x5093x = (((!n_n52) & (!n_n101) & (!x39x) & (!x58x) & (x1359x)) + ((n_n52) & (!n_n101) & (x39x) & (!x58x) & (!x1359x)) + ((!n_n52) & (n_n101) & (!x39x) & (x58x) & (!x1359x)));
	assign x5099x = (((!x337x) & (n_n1039) & (!n_n1091) & (!x322x) & (!n_n1103)) + ((!x337x) & (!n_n1039) & (n_n1091) & (!x322x) & (!n_n1103)) + ((!x337x) & (!n_n1039) & (!n_n1091) & (!x322x) & (n_n1103)) + ((x337x) & (!n_n1039) & (!n_n1091) & (x322x) & (!n_n1103)));
	assign x5100x = (((!x49x) & (n_n1120) & (!n_n1052) & (!n_n1331) & (!x177x)) + ((!x49x) & (!n_n1120) & (n_n1052) & (!n_n1331) & (!x177x)) + ((!x49x) & (!n_n1120) & (!n_n1052) & (n_n1331) & (!x177x)) + ((x49x) & (!n_n1120) & (!n_n1052) & (!n_n1331) & (x177x)));
	assign x5101x = (((!n_n82) & (!x21x) & (!x46x) & (!x173x) & (x233x)) + ((n_n82) & (!x21x) & (x46x) & (!x173x) & (!x233x)) + ((!n_n82) & (x21x) & (!x46x) & (x173x) & (!x233x)));
	assign x5103x = (((x117x) & (!x133x) & (!x148x) & (!x323x) & (!x1352x)) + ((!x117x) & (x133x) & (!x148x) & (!x323x) & (!x1352x)) + ((!x117x) & (!x133x) & (x148x) & (!x323x) & (!x1352x)) + ((!x117x) & (!x133x) & (!x148x) & (x323x) & (!x1352x)) + ((!x117x) & (!x133x) & (!x148x) & (!x323x) & (x1352x)));
	assign x5104x = (((!n_n83) & (!x35x) & (x201x) & (!x256x) & (!x271x)) + ((!n_n83) & (!x35x) & (!x201x) & (x256x) & (!x271x)) + ((!n_n83) & (!x35x) & (!x201x) & (!x256x) & (x271x)) + ((n_n83) & (x35x) & (!x201x) & (!x256x) & (!x271x)));
	assign x5114x = (((!i_3_) & (!x341x) & (!n_n83) & (!n_n82) & (n_n989)) + ((i_3_) & (x341x) & (n_n83) & (n_n82) & (!n_n989)));
	assign x5148x = (((!n_n64) & (n_n101) & (!n_n85) & (x49x) & (!n_n76)) + ((n_n64) & (!n_n101) & (n_n85) & (!x49x) & (n_n76)));
	assign x5150x = (((!x27x) & (x113x) & (!n_n63) & (!n_n95) & (!x34x)) + ((x27x) & (!x113x) & (!n_n63) & (n_n95) & (!x34x)) + ((!x27x) & (!x113x) & (n_n63) & (!n_n95) & (x34x)));
	assign x5151x = (((!n_n101) & (!n_n83) & (!n_n102) & (x105x) & (!x1359x)) + ((!n_n101) & (!n_n83) & (!n_n102) & (!x105x) & (x1359x)) + ((n_n101) & (n_n83) & (n_n102) & (!x105x) & (!x1359x)));
	assign x5152x = (((!n_n101) & (!n_n103) & (!n_n84) & (x117x) & (!x1292x)) + ((!n_n101) & (!n_n103) & (!n_n84) & (!x117x) & (x1292x)) + ((n_n101) & (n_n103) & (n_n84) & (!x117x) & (!x1292x)));
	assign x5159x = (((!n_n93) & (!n_n84) & (x233x) & (!x36x) & (!x48x)) + ((n_n93) & (!n_n84) & (!x233x) & (x36x) & (!x48x)) + ((!n_n93) & (n_n84) & (!x233x) & (!x36x) & (x48x)));
	assign x5205x = (((!i_7_) & (!i_8_) & (!i_6_) & (x352x) & (!x63x)) + ((i_7_) & (!i_8_) & (i_6_) & (!x352x) & (x63x)));
	assign x5206x = (((!i_2_) & (n_n91) & (!x56x) & (x49x) & (!x318x)) + ((!i_2_) & (!n_n91) & (x56x) & (!x49x) & (x318x)));
	assign x5208x = (((!i_7_) & (!i_8_) & (!i_6_) & (x105x) & (!x41x)) + ((!i_7_) & (!i_8_) & (i_6_) & (!x105x) & (x41x)));
	assign x5214x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x46x) & (x5206x)) + ((i_7_) & (i_8_) & (i_6_) & (x46x) & (!x5206x)) + ((i_7_) & (!i_8_) & (!i_6_) & (x46x) & (!x5206x)));
	assign x5217x = (((x323x) & (!n_n1330) & (!x185x) & (!x258x) & (!x5205x)) + ((!x323x) & (n_n1330) & (!x185x) & (!x258x) & (!x5205x)) + ((!x323x) & (!n_n1330) & (x185x) & (!x258x) & (!x5205x)) + ((!x323x) & (!n_n1330) & (!x185x) & (x258x) & (!x5205x)) + ((!x323x) & (!n_n1330) & (!x185x) & (!x258x) & (x5205x)));
	assign x6355x = (((!n_n77) & (!x1291x) & (!x1292x) & (!x183x) & (!x31x)) + ((!n_n77) & (!x1291x) & (!x1292x) & (!x183x) & (!x31x)));
	assign x5244x = (((!n_n78) & (!x67x) & (n_n1057) & (!n_n1125) & (!x248x)) + ((!n_n78) & (!x67x) & (!n_n1057) & (n_n1125) & (!x248x)) + ((!n_n78) & (!x67x) & (!n_n1057) & (!n_n1125) & (x248x)) + ((n_n78) & (x67x) & (!n_n1057) & (!n_n1125) & (!x248x)));
	assign x5283x = (((!i_8_) & (!x341x) & (!n_n52) & (!x75x) & (x252x)) + ((i_8_) & (x341x) & (n_n52) & (x75x) & (!x252x)));
	assign x5288x = (((!i_1_) & (!n_n64) & (!n_n40) & (!x30x) & (x1108x)) + ((i_1_) & (n_n64) & (n_n40) & (x30x) & (!x1108x)));
	assign x6356x = (((i_1_) & (!i_2_) & (!n_n70) & (!n_n77) & (!n_n87)) + ((!i_1_) & (!i_2_) & (!n_n70) & (!n_n77) & (!n_n87)) + ((!i_1_) & (!i_2_) & (!n_n70) & (!n_n77) & (!n_n87)) + ((!i_1_) & (!i_2_) & (!n_n70) & (!n_n77) & (!n_n87)) + ((!i_1_) & (!i_2_) & (!n_n70) & (!n_n77) & (!n_n87)));
	assign x5289x = (((!i_7_) & (!i_8_) & (!i_4_) & (!x311x) & (!x6356x)) + ((!i_7_) & (i_8_) & (i_4_) & (x311x) & (!x6356x)));
	assign x5290x = (((!n_n93) & (!n_n102) & (x127x) & (x328x) & (!x175x)) + ((n_n93) & (n_n102) & (!x127x) & (!x328x) & (x175x)));
	assign x5291x = (((!i_7_) & (!i_8_) & (n_n103) & (!n_n100) & (n_n76)) + ((i_7_) & (i_8_) & (!n_n103) & (n_n100) & (n_n76)));
	assign x5292x = (((!i_4_) & (x234x) & (!x66x) & (x242x) & (!x28x)) + ((!i_4_) & (!x234x) & (x66x) & (!x242x) & (x28x)));
	assign x5293x = (((!n_n93) & (!n_n84) & (x109x) & (!n_n90) & (x85x)) + ((n_n93) & (n_n84) & (!x109x) & (n_n90) & (!x85x)));
	assign x5305x = (((!n_n91) & (!x58x) & (!n_n82) & (!x67x) & (x5293x)) + ((!n_n91) & (x58x) & (n_n82) & (!x67x) & (!x5293x)) + ((n_n91) & (!x58x) & (!n_n82) & (x67x) & (!x5293x)));
	assign x6349x = (((i_7_) & (!i_8_) & (!x32x) & (!n_n74) & (!x44x)) + ((!i_7_) & (i_8_) & (!x32x) & (!n_n74) & (!x44x)) + ((i_7_) & (!i_8_) & (!x32x) & (!n_n74) & (!x44x)) + ((!i_7_) & (i_8_) & (!x32x) & (!n_n74) & (!x44x)) + ((!i_7_) & (!i_8_) & (!x32x) & (!n_n74) & (!x44x)) + ((!i_7_) & (!i_8_) & (!x32x) & (!n_n74) & (!x44x)));
	assign x6346x = (((!n_n1217) & (!x174x) & (!x336x) & (!x246x) & (!x339x)) + ((!n_n1217) & (!x174x) & (!x336x) & (!x246x) & (!x339x)));
	assign x5321x = (((!i_8_) & (!i_6_) & (!i_3_) & (!n_n85) & (n_n1030)) + ((!i_8_) & (!i_6_) & (!i_3_) & (n_n85) & (!n_n1030)));
	assign x5322x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x55x) & (n_n1058)) + ((i_7_) & (i_8_) & (i_6_) & (x55x) & (!n_n1058)));
	assign x5342x = (((!i_1_) & (!i_2_) & (!n_n64) & (!x109x) & (x83x)) + ((i_1_) & (i_2_) & (n_n64) & (x109x) & (!x83x)));
	assign x5351x = (((!i_6_) & (!n_n70) & (!x110x) & (!n_n53) & (x319x)) + ((!i_6_) & (n_n70) & (x110x) & (n_n53) & (!x319x)));
	assign x5358x = (((!n_n101) & (n_n989) & (!x52x) & (!n_n944) & (!n_n982)) + ((!n_n101) & (!n_n989) & (!x52x) & (n_n944) & (!n_n982)) + ((!n_n101) & (!n_n989) & (!x52x) & (!n_n944) & (n_n982)) + ((n_n101) & (!n_n989) & (x52x) & (!n_n944) & (!n_n982)));
	assign x5359x = (((!n_n78) & (!x42x) & (n_n967) & (!n_n1121) & (!x236x)) + ((!n_n78) & (!x42x) & (!n_n967) & (n_n1121) & (!x236x)) + ((!n_n78) & (!x42x) & (!n_n967) & (!n_n1121) & (x236x)) + ((n_n78) & (x42x) & (!n_n967) & (!n_n1121) & (!x236x)));
	assign x5360x = (((!n_n73) & (!x42x) & (!x111x) & (x5342x) & (!x5351x)) + ((!n_n73) & (!x42x) & (!x111x) & (!x5342x) & (x5351x)) + ((n_n73) & (x42x) & (x111x) & (!x5342x) & (!x5351x)));
	assign x5362x = (((!n_n101) & (x97x) & (!x145x) & (!n_n951) & (!x44x)) + ((!n_n101) & (!x97x) & (x145x) & (!n_n951) & (!x44x)) + ((!n_n101) & (!x97x) & (!x145x) & (n_n951) & (!x44x)) + ((n_n101) & (!x97x) & (!x145x) & (!n_n951) & (x44x)));
	assign x5364x = (((!i_8_) & (!x70x) & (x215x) & (!x262x) & (!x275x)) + ((!i_8_) & (!x70x) & (!x215x) & (x262x) & (!x275x)) + ((!i_8_) & (!x70x) & (!x215x) & (!x262x) & (x275x)) + ((!i_8_) & (x70x) & (!x215x) & (!x262x) & (!x275x)));
	assign x6344x = (((!x245x) & (!x38x) & (!n_n1093) & (!n_n1074) & (!n_n1087)) + ((!x245x) & (!x38x) & (!n_n1093) & (!n_n1074) & (!n_n1087)));
	assign x6351x = (((!n_n80) & (!n_n83) & (!x234x) & (!x320x) & (!n_n973)) + ((!n_n80) & (!n_n83) & (!x234x) & (!x320x) & (!n_n973)) + ((!n_n80) & (!n_n83) & (!x234x) & (!x320x) & (!n_n973)) + ((!n_n80) & (!n_n83) & (!x234x) & (!x320x) & (!n_n973)));
	assign x5411x = (((i_3_) & (!n_n78) & (!n_n85) & (x37x) & (x109x)) + ((i_3_) & (n_n78) & (n_n85) & (!x37x) & (x109x)));
	assign x5429x = (((!n_n70) & (x48x) & (!n_n87) & (x194x) & (!x353x)) + ((n_n70) & (!x48x) & (n_n87) & (!x194x) & (x353x)));
	assign x5446x = (((!i_5_) & (!i_6_) & (!n_n75) & (x251x) & (!n_n90)) + ((!i_5_) & (i_6_) & (n_n75) & (!x251x) & (n_n90)));
	assign x5460x = (((!i_7_) & (!i_3_) & (n_n1078) & (!n_n40) & (!x330x)) + ((i_7_) & (i_3_) & (!n_n1078) & (n_n40) & (x330x)));
	assign x5467x = (((!i_8_) & (!i_2_) & (!n_n54) & (!x56x) & (x355x)) + ((i_8_) & (!i_2_) & (n_n54) & (x56x) & (!x355x)));
	assign x5468x = (((!i_8_) & (!n_n85) & (!x127x) & (x21x) & (x173x)) + ((i_8_) & (n_n85) & (x127x) & (!x21x) & (!x173x)));
	assign x5472x = (((!i_7_) & (!i_6_) & (!x26x) & (n_n1085) & (!x279x)) + ((!i_7_) & (!i_6_) & (!x26x) & (!n_n1085) & (x279x)) + ((!i_7_) & (!i_6_) & (x26x) & (!n_n1085) & (!x279x)));
	assign x5474x = (((!i_6_) & (!n_n86) & (!x43x) & (n_n1125) & (!x5460x)) + ((!i_6_) & (!n_n86) & (!x43x) & (!n_n1125) & (x5460x)) + ((i_6_) & (n_n86) & (x43x) & (!n_n1125) & (!x5460x)));
	assign x5475x = (((!n_n73) & (n_n1082) & (!x36x) & (!n_n1045) & (!n_n1043)) + ((!n_n73) & (!n_n1082) & (!x36x) & (n_n1045) & (!n_n1043)) + ((!n_n73) & (!n_n1082) & (!x36x) & (!n_n1045) & (n_n1043)) + ((n_n73) & (!n_n1082) & (x36x) & (!n_n1045) & (!n_n1043)));
	assign x5478x = (((!n_n91) & (!n_n40) & (!x66x) & (!x44x) & (x5468x)) + ((!n_n91) & (n_n40) & (x66x) & (!x44x) & (!x5468x)) + ((n_n91) & (!n_n40) & (!x66x) & (x44x) & (!x5468x)));
	assign x5479x = (((x141x) & (!x142x) & (!x150x) & (!n_n1046) & (!n_n1047)) + ((!x141x) & (x142x) & (!x150x) & (!n_n1046) & (!n_n1047)) + ((!x141x) & (!x142x) & (x150x) & (!n_n1046) & (!n_n1047)) + ((!x141x) & (!x142x) & (!x150x) & (n_n1046) & (!n_n1047)) + ((!x141x) & (!x142x) & (!x150x) & (!n_n1046) & (n_n1047)));
	assign x6343x = (((!n_n1118) & (!n_n1030) & (!x66x) & (!x5442x) & (!n_n1101)) + ((!n_n1118) & (!n_n1030) & (!x66x) & (!x5442x) & (!n_n1101)));
	assign x5482x = (((!n_n101) & (n_n1036) & (!x128x) & (!x5467x) & (!x6343x)) + ((!n_n101) & (!n_n1036) & (!x128x) & (x5467x) & (!x6343x)) + ((!n_n101) & (!n_n1036) & (!x128x) & (!x5467x) & (!x6343x)) + ((n_n101) & (!n_n1036) & (x128x) & (!x5467x) & (!x6343x)));
	assign x5499x = (((!i_8_) & (!n_n38) & (n_n1153) & (!x110x) & (!x175x)) + ((!i_8_) & (n_n38) & (!n_n1153) & (x110x) & (x175x)));
	assign x5518x = (((!i_5_) & (i_2_) & (n_n101) & (x54x) & (x175x)) + ((i_5_) & (!i_2_) & (n_n101) & (x54x) & (x175x)));
	assign x5519x = (((!i_3_) & (!x109x) & (x78x) & (!x129x) & (x174x)) + ((!i_3_) & (x109x) & (!x78x) & (x129x) & (!x174x)));
	assign x5522x = (((!n_n58) & (n_n100) & (n_n102) & (n_n63) & (!n_n77)) + ((n_n58) & (n_n100) & (!n_n102) & (!n_n63) & (n_n77)));
	assign x5526x = (((!n_n64) & (!n_n52) & (!x65x) & (x166x) & (!x869x)) + ((!n_n64) & (!n_n52) & (!x65x) & (!x166x) & (x869x)) + ((n_n64) & (n_n52) & (x65x) & (!x166x) & (!x869x)));
	assign x5528x = (((!n_n78) & (n_n1259) & (!x53x) & (!n_n1176) & (!n_n1184)) + ((!n_n78) & (!n_n1259) & (!x53x) & (n_n1176) & (!n_n1184)) + ((!n_n78) & (!n_n1259) & (!x53x) & (!n_n1176) & (n_n1184)) + ((n_n78) & (!n_n1259) & (x53x) & (!n_n1176) & (!n_n1184)));
	assign x5529x = (((!n_n101) & (!n_n100) & (!n_n74) & (x340x) & (!x5518x)) + ((!n_n101) & (!n_n100) & (!n_n74) & (!x340x) & (x5518x)) + ((n_n101) & (n_n100) & (n_n74) & (!x340x) & (!x5518x)));
	assign x5531x = (((!i_5_) & (!i_3_) & (!i_4_) & (!x48x) & (x5522x)) + ((i_5_) & (i_3_) & (i_4_) & (x48x) & (!x5522x)) + ((!i_5_) & (i_3_) & (!i_4_) & (x48x) & (!x5522x)));
	assign x5568x = (((!i_8_) & (!i_6_) & (!n_n103) & (!n_n77) & (n_n1059)) + ((i_8_) & (i_6_) & (n_n103) & (n_n77) & (!n_n1059)));
	assign x5571x = (((!n_n38) & (!n_n70) & (!x29x) & (n_n1087) & (!x153x)) + ((!n_n38) & (!n_n70) & (!x29x) & (!n_n1087) & (x153x)) + ((n_n38) & (n_n70) & (x29x) & (!n_n1087) & (!x153x)));
	assign x5573x = (((!n_n78) & (!x42x) & (n_n1093) & (!n_n1057) & (!n_n1045)) + ((!n_n78) & (!x42x) & (!n_n1093) & (n_n1057) & (!n_n1045)) + ((!n_n78) & (!x42x) & (!n_n1093) & (!n_n1057) & (n_n1045)) + ((n_n78) & (x42x) & (!n_n1093) & (!n_n1057) & (!n_n1045)));
	assign x5574x = (((!n_n91) & (!x53x) & (n_n1101) & (!n_n1060) & (!n_n1100)) + ((!n_n91) & (!x53x) & (!n_n1101) & (n_n1060) & (!n_n1100)) + ((!n_n91) & (!x53x) & (!n_n1101) & (!n_n1060) & (n_n1100)) + ((n_n91) & (x53x) & (!n_n1101) & (!n_n1060) & (!n_n1100)));
	assign x5575x = (((!n_n77) & (n_n1046) & (!x132x) & (!n_n954) & (!n_n939)) + ((!n_n77) & (!n_n1046) & (!x132x) & (n_n954) & (!n_n939)) + ((!n_n77) & (!n_n1046) & (!x132x) & (!n_n954) & (n_n939)) + ((n_n77) & (!n_n1046) & (x132x) & (!n_n954) & (!n_n939)));
	assign x5576x = (((!n_n74) & (n_n1058) & (!n_n971) & (!x107x) & (!n_n1037)) + ((!n_n74) & (!n_n1058) & (n_n971) & (!x107x) & (!n_n1037)) + ((!n_n74) & (!n_n1058) & (!n_n971) & (!x107x) & (n_n1037)) + ((n_n74) & (!n_n1058) & (!n_n971) & (x107x) & (!n_n1037)));
	assign x5579x = (((!n_n95) & (!x29x) & (x829x) & (!x292x) & (!n_n947)) + ((!n_n95) & (!x29x) & (!x829x) & (x292x) & (!n_n947)) + ((!n_n95) & (!x29x) & (!x829x) & (!x292x) & (n_n947)) + ((n_n95) & (x29x) & (!x829x) & (!x292x) & (!n_n947)));
	assign x5580x = (((x254x) & (!x285x) & (!x68x) & (!x138x)) + ((!x254x) & (x285x) & (!x68x) & (!x138x)) + ((!x254x) & (!x285x) & (x68x) & (!x138x)) + ((!x254x) & (!x285x) & (!x68x) & (x138x)));
	assign x6358x = (((!x97x) & (!x298x) & (!x903x) & (!x5492x) & (!x125x)));
	assign x5595x = (((!i_7_) & (!i_8_) & (i_2_) & (x175x) & (x130x)) + ((!i_7_) & (i_8_) & (!i_2_) & (x175x) & (x130x)));
	assign x5641x = (((!n_n95) & (n_n1134) & (!n_n1132) & (!x128x) & (!n_n962)) + ((!n_n95) & (!n_n1134) & (n_n1132) & (!x128x) & (!n_n962)) + ((!n_n95) & (!n_n1134) & (!n_n1132) & (!x128x) & (n_n962)) + ((n_n95) & (!n_n1134) & (!n_n1132) & (x128x) & (!n_n962)));
	assign x5642x = (((!n_n101) & (!n_n100) & (!x78x) & (!x128x) & (x218x)) + ((!n_n101) & (n_n100) & (x78x) & (!x128x) & (!x218x)) + ((n_n101) & (!n_n100) & (!x78x) & (x128x) & (!x218x)));
	assign x5643x = (((!n_n101) & (n_n1058) & (!n_n1101) & (!x44x) & (!n_n954)) + ((!n_n101) & (!n_n1058) & (n_n1101) & (!x44x) & (!n_n954)) + ((!n_n101) & (!n_n1058) & (!n_n1101) & (!x44x) & (n_n954)) + ((n_n101) & (!n_n1058) & (!n_n1101) & (x44x) & (!n_n954)));
	assign x5644x = (((n_n1079) & (!x324x) & (!n_n67) & (!x345x) & (!n_n978)) + ((!n_n1079) & (!x324x) & (!n_n67) & (x345x) & (!n_n978)) + ((!n_n1079) & (!x324x) & (!n_n67) & (!x345x) & (n_n978)) + ((!n_n1079) & (x324x) & (n_n67) & (!x345x) & (!n_n978)));
	assign x6341x = (((!i_1_) & (!n_n91) & (!x45x) & (!n_n77) & (!n_n959)) + ((!i_1_) & (!n_n91) & (!x45x) & (!n_n77) & (!n_n959)) + ((!i_1_) & (!n_n91) & (!x45x) & (!n_n77) & (!n_n959)));
	assign x5645x = (((!i_7_) & (!i_8_) & (!n_n94) & (!n_n66) & (!x6341x)) + ((i_7_) & (i_8_) & (n_n94) & (n_n66) & (!x6341x)));
	assign x5646x = (((!n_n73) & (!n_n70) & (!x53x) & (!x33x) & (x287x)) + ((n_n73) & (!n_n70) & (x53x) & (!x33x) & (!x287x)) + ((!n_n73) & (n_n70) & (!x53x) & (x33x) & (!x287x)));
	assign x5648x = (((n_n944) & (!n_n939) & (!x162x) & (!x91x) & (!x266x)) + ((!n_n944) & (n_n939) & (!x162x) & (!x91x) & (!x266x)) + ((!n_n944) & (!n_n939) & (x162x) & (!x91x) & (!x266x)) + ((!n_n944) & (!n_n939) & (!x162x) & (x91x) & (!x266x)) + ((!n_n944) & (!n_n939) & (!x162x) & (!x91x) & (x266x)));
	assign x6340x = (((!x1483x) & (!x1484x) & (!x279x) & (!x153x) & (!x204x)));
	assign x5664x = (((!i_5_) & (!i_3_) & (!n_n38) & (!n_n94) & (x235x)) + ((i_5_) & (!i_3_) & (n_n38) & (n_n94) & (!x235x)));
	assign x5668x = (((!i_5_) & (i_3_) & (!i_4_) & (n_n91) & (n_n94)) + ((!i_5_) & (!i_3_) & (!i_4_) & (n_n91) & (n_n94)));
	assign x5672x = (((!n_n101) & (!x55x) & (!x112x) & (n_n1163) & (!x1143x)) + ((!n_n101) & (!x55x) & (!x112x) & (!n_n1163) & (x1143x)) + ((n_n101) & (x55x) & (!x112x) & (!n_n1163) & (!x1143x)) + ((n_n101) & (!x55x) & (x112x) & (!n_n1163) & (!x1143x)));
	assign x5673x = (((!n_n78) & (!x63x) & (!x52x) & (n_n1216) & (!n_n1146)) + ((!n_n78) & (!x63x) & (!x52x) & (!n_n1216) & (n_n1146)) + ((n_n78) & (x63x) & (!x52x) & (!n_n1216) & (!n_n1146)) + ((n_n78) & (!x63x) & (x52x) & (!n_n1216) & (!n_n1146)));
	assign x6342x = (((!n_n94) & (!n_n1188) & (!n_n1193) & (!x342x) & (!x5493x)) + ((!n_n94) & (!n_n1188) & (!n_n1193) & (!x342x) & (!x5493x)));
	assign x5693x = (((!i_5_) & (!i_6_) & (!i_3_) & (!x328x) & (x350x)) + ((i_5_) & (!i_6_) & (!i_3_) & (x328x) & (!x350x)));
	assign x5694x = (((!n_n75) & (!n_n94) & (x38x) & (x174x) & (!x130x)) + ((n_n75) & (n_n94) & (!x38x) & (!x174x) & (x130x)));
	assign x5695x = (((!i_3_) & (!x341x) & (x66x) & (x131x) & (!x107x)) + ((i_3_) & (x341x) & (!x66x) & (!x131x) & (x107x)));
	assign x5697x = (((!i_5_) & (n_n91) & (!x54x) & (x21x) & (!x20x)) + ((!i_5_) & (!n_n91) & (x54x) & (!x21x) & (x20x)));
	assign x5715x = (((!i_3_) & (!i_1_) & (!i_2_) & (x333x) & (!x339x)) + ((i_3_) & (!i_1_) & (i_2_) & (!x333x) & (x339x)));
	assign x6353x = (((i_7_) & (!i_8_) & (!i_6_) & (!x39x) & (!x64x)) + ((!i_7_) & (!i_8_) & (!i_6_) & (!x39x) & (!x64x)) + ((!i_7_) & (i_8_) & (!i_6_) & (!x39x) & (!x64x)) + ((!i_7_) & (!i_8_) & (!i_6_) & (!x39x) & (!x64x)));
	assign x5727x = (((x255x) & (!x226x) & (!x71x) & (!x876x) & (!x877x)) + ((!x255x) & (x226x) & (!x71x) & (!x876x) & (!x877x)) + ((!x255x) & (!x226x) & (x71x) & (!x876x) & (!x877x)) + ((!x255x) & (!x226x) & (!x71x) & (x876x) & (!x877x)) + ((!x255x) & (!x226x) & (!x71x) & (!x876x) & (x877x)));
	assign x6336x = (((!n_n1134) & (!n_n1331) & (!x248x) & (!x5686x) & (!x5687x)) + ((!n_n1134) & (!n_n1331) & (!x248x) & (!x5686x) & (!x5687x)));
	assign x5751x = (((!i_0_) & (n_n91) & (x64x) & (!x38x) & (!x30x)) + ((i_0_) & (!n_n91) & (!x64x) & (x38x) & (x30x)));
	assign x5753x = (((!i_6_) & (!i_3_) & (!i_4_) & (x236x) & (!x66x)) + ((i_6_) & (i_3_) & (!i_4_) & (!x236x) & (x66x)));
	assign x5758x = (((i_7_) & (!i_8_) & (!x245x) & (x67x) & (!n_n66)) + ((!i_7_) & (!i_8_) & (x245x) & (!x67x) & (n_n66)));
	assign x5763x = (((!n_n91) & (!n_n102) & (!n_n97) & (n_n939) & (!x161x)) + ((!n_n91) & (!n_n102) & (!n_n97) & (!n_n939) & (x161x)) + ((n_n91) & (n_n102) & (n_n97) & (!n_n939) & (!x161x)));
	assign x5769x = (((!n_n101) & (!n_n84) & (!n_n85) & (x97x) & (!x5758x)) + ((!n_n101) & (!n_n84) & (!n_n85) & (!x97x) & (x5758x)) + ((n_n101) & (n_n84) & (n_n85) & (!x97x) & (!x5758x)));
	assign x5770x = (((x256x) & (!x215x) & (!x141x) & (!x142x)) + ((!x256x) & (x215x) & (!x141x) & (!x142x)) + ((!x256x) & (!x215x) & (x141x) & (!x142x)) + ((!x256x) & (!x215x) & (!x141x) & (x142x)));
	assign x6338x = (((!n_n58) & (!n_n95) & (!n_n1132) & (!x44x) & (!n_n971)) + ((!n_n58) & (!n_n95) & (!n_n1132) & (!x44x) & (!n_n971)));
	assign x6350x = (((!x55x) & (!n_n95) & (!n_n983) & (!x354x) & (!x4944x)) + ((!x55x) & (!n_n95) & (!n_n983) & (!x354x) & (!x4944x)) + ((!x55x) & (!n_n95) & (!n_n983) & (!x354x) & (!x4944x)) + ((!x55x) & (!n_n95) & (!n_n983) & (!x354x) & (!x4944x)));
	assign x6337x = (((!n_n1087) & (!x805x) & (!x79x) & (!x91x) & (!x103x)));
	assign x5798x = (((!i_1_) & (n_n80) & (!n_n58) & (!x110x) & (x234x)) + ((i_1_) & (!n_n80) & (n_n58) & (x110x) & (!x234x)));
	assign x5808x = (((!n_n78) & (!x42x) & (n_n989) & (!x5798x)) + ((!n_n78) & (!x42x) & (!n_n989) & (x5798x)) + ((n_n78) & (x42x) & (!n_n989) & (!x5798x)));
	assign x5809x = (((!x64x) & (!n_n95) & (n_n969) & (!n_n999) & (!n_n1004)) + ((!x64x) & (!n_n95) & (!n_n969) & (n_n999) & (!n_n1004)) + ((!x64x) & (!n_n95) & (!n_n969) & (!n_n999) & (n_n1004)) + ((x64x) & (n_n95) & (!n_n969) & (!n_n999) & (!n_n1004)));
	assign x5810x = (((!x25x) & (!n_n95) & (!x173x) & (x168x) & (!x237x)) + ((x25x) & (!n_n95) & (x173x) & (!x168x) & (!x237x)) + ((!x25x) & (n_n95) & (!x173x) & (!x168x) & (x237x)));
	assign x5812x = (((n_n980) & (!n_n983) & (!n_n986) & (!x753x) & (!x5609x)) + ((!n_n980) & (n_n983) & (!n_n986) & (!x753x) & (!x5609x)) + ((!n_n980) & (!n_n983) & (n_n986) & (!x753x) & (!x5609x)) + ((!n_n980) & (!n_n983) & (!n_n986) & (x753x) & (!x5609x)) + ((!n_n980) & (!n_n983) & (!n_n986) & (!x753x) & (x5609x)));
	assign x5814x = (((n_n973) & (!x145x) & (!n_n975) & (!x272x) & (!x147x)) + ((!n_n973) & (x145x) & (!n_n975) & (!x272x) & (!x147x)) + ((!n_n973) & (!x145x) & (n_n975) & (!x272x) & (!x147x)) + ((!n_n973) & (!x145x) & (!n_n975) & (x272x) & (!x147x)) + ((!n_n973) & (!x145x) & (!n_n975) & (!x272x) & (x147x)));
	assign x6357x = (((!x97x) & (!x125x) & (!n_n994) & (!x163x) & (!n_n978)));
	assign x5835x = (((n_n75) & (!n_n74) & (x63x) & (!n_n67) & (!x5828x)) + ((!n_n75) & (n_n74) & (!x63x) & (!n_n67) & (x5828x)));
	assign x6335x = (((!n_n1092) & (!n_n1091) & (!n_n1100) & (!x354x) & (!x4944x)) + ((!n_n1092) & (!n_n1091) & (!n_n1100) & (!x354x) & (!x4944x)));
	assign x5848x = (((!i_5_) & (i_3_) & (!i_4_) & (n_n78) & (n_n90)));
	assign x5850x = (((!i_7_) & (!i_8_) & (!i_6_) & (!x128x) & (n_n1177)) + ((!i_7_) & (i_8_) & (i_6_) & (x128x) & (!n_n1177)));
	assign x5852x = (((!i_5_) & (!i_6_) & (!i_3_) & (!x316x) & (x344x)) + ((i_5_) & (i_6_) & (i_3_) & (x316x) & (!x344x)));
	assign x5853x = (((!i_7_) & (!i_8_) & (n_n103) & (!n_n85) & (n_n76)) + ((i_7_) & (i_8_) & (!n_n103) & (n_n85) & (n_n76)));
	assign x5854x = (((!i_7_) & (i_8_) & (i_6_) & (x239x) & (!x41x)) + ((i_7_) & (!i_8_) & (i_6_) & (!x239x) & (x41x)) + ((!i_7_) & (i_8_) & (!i_6_) & (!x239x) & (x41x)));
	assign x5855x = (((!i_7_) & (i_8_) & (!i_6_) & (x45x) & (!x49x)) + ((i_7_) & (!i_8_) & (!i_6_) & (!x45x) & (x49x)));
	assign x5856x = (((!i_5_) & (n_n91) & (!n_n100) & (x39x) & (!x54x)) + ((i_5_) & (n_n91) & (n_n100) & (!x39x) & (x54x)));
	assign x5858x = (((!x57x) & (!n_n92) & (!n_n95) & (x88x) & (!x132x)) + ((x57x) & (!n_n92) & (n_n95) & (!x88x) & (!x132x)) + ((!x57x) & (n_n92) & (!n_n95) & (!x88x) & (x132x)));
	assign x5859x = (((!i_5_) & (!x54x) & (x343x) & (!x48x) & (!x185x)) + ((!i_5_) & (!x54x) & (!x343x) & (!x48x) & (x185x)) + ((i_5_) & (x54x) & (!x343x) & (x48x) & (!x185x)));
	assign x5860x = (((!n_n73) & (!x111x) & (n_n1169) & (!x120x) & (!x238x)) + ((!n_n73) & (!x111x) & (!n_n1169) & (x120x) & (!x238x)) + ((n_n73) & (x111x) & (!n_n1169) & (!x120x) & (x238x)));
	assign x5866x = (((!n_n52) & (!n_n82) & (!x21x) & (!x22x) & (x5856x)) + ((!n_n52) & (n_n82) & (x21x) & (!x22x) & (!x5856x)) + ((n_n52) & (!n_n82) & (!x21x) & (x22x) & (!x5856x)));
	assign x5880x = (((!i_2_) & (x55x) & (n_n95) & (!x5493x) & (!x175x)) + ((!i_2_) & (!x55x) & (!n_n95) & (x5493x) & (x175x)));
	assign x5881x = (((!i_7_) & (!i_8_) & (!i_3_) & (!x5687x) & (n_n1009)) + ((!i_7_) & (!i_8_) & (!i_3_) & (x5687x) & (!n_n1009)));
	assign x5882x = (((!i_3_) & (!i_1_) & (!i_2_) & (!x339x) & (n_n1013)) + ((i_3_) & (!i_1_) & (i_2_) & (x339x) & (!n_n1013)));
	assign x5899x = (((!n_n81) & (n_n91) & (n_n103) & (n_n102) & (!n_n82)) + ((n_n81) & (!n_n91) & (n_n103) & (!n_n102) & (n_n82)));
	assign x5914x = (((i_3_) & (!i_1_) & (i_2_) & (x78x) & (!x324x)) + ((!i_3_) & (i_1_) & (i_2_) & (!x78x) & (x324x)));
	assign x5915x = (((!n_n93) & (!n_n103) & (!n_n74) & (x38x) & (x174x)) + ((n_n93) & (n_n103) & (n_n74) & (!x38x) & (!x174x)));
	assign x5918x = (((!i_3_) & (n_n58) & (x19x) & (!x109x) & (!x20x)) + ((i_3_) & (!n_n58) & (!x19x) & (x109x) & (x20x)));
	assign x5919x = (((!i_5_) & (!x32x) & (!x54x) & (x346x) & (!x190x)) + ((!i_5_) & (!x32x) & (!x54x) & (!x346x) & (x190x)) + ((i_5_) & (x32x) & (x54x) & (!x346x) & (!x190x)));
	assign x5921x = (((!n_n58) & (!x26x) & (!x32x) & (!n_n102) & (x157x)) + ((n_n58) & (x26x) & (!x32x) & (!n_n102) & (!x157x)) + ((!n_n58) & (!x26x) & (x32x) & (n_n102) & (!x157x)));
	assign x5922x = (((!n_n78) & (!n_n92) & (!n_n85) & (x210x) & (!x663x)) + ((!n_n78) & (!n_n92) & (!n_n85) & (!x210x) & (x663x)) + ((n_n78) & (n_n92) & (n_n85) & (!x210x) & (!x663x)));
	assign x5924x = (((x235x) & (!n_n1286) & (!x131x) & (!x5068x) & (!n_n1158)) + ((!x235x) & (n_n1286) & (!x131x) & (!x5068x) & (!n_n1158)) + ((!x235x) & (!n_n1286) & (!x131x) & (!x5068x) & (n_n1158)) + ((!x235x) & (!n_n1286) & (x131x) & (x5068x) & (!n_n1158)));
	assign x5926x = (((!n_n75) & (!x45x) & (!x25x) & (!n_n95) & (x5915x)) + ((n_n75) & (!x45x) & (x25x) & (!n_n95) & (!x5915x)) + ((!n_n75) & (x45x) & (!x25x) & (n_n95) & (!x5915x)));
	assign x5927x = (((!n_n52) & (!n_n101) & (!x21x) & (!x22x) & (x5918x)) + ((!n_n52) & (n_n101) & (x21x) & (!x22x) & (!x5918x)) + ((n_n52) & (!n_n101) & (!x21x) & (x22x) & (!x5918x)));
	assign x5933x = (((n_n1312) & (!x129x) & (!x5338x) & (!x5914x) & (!x5926x)) + ((!n_n1312) & (!x129x) & (!x5338x) & (x5914x) & (!x5926x)) + ((!n_n1312) & (!x129x) & (!x5338x) & (!x5914x) & (x5926x)) + ((!n_n1312) & (x129x) & (x5338x) & (!x5914x) & (!x5926x)));
	assign x5944x = (((!i_5_) & (!i_4_) & (!n_n58) & (n_n1039) & (!x327x)) + ((!i_5_) & (!i_4_) & (n_n58) & (!n_n1039) & (x327x)));
	assign x5946x = (((!i_6_) & (!i_3_) & (!i_4_) & (!x66x) & (n_n1013)) + ((i_6_) & (i_3_) & (!i_4_) & (x66x) & (!n_n1013)));
	assign x5965x = (((!i_5_) & (n_n80) & (x337x) & (!x247x) & (!x28x)) + ((!i_5_) & (!n_n80) & (!x337x) & (x247x) & (x28x)));
	assign x5966x = (((!n_n64) & (!n_n100) & (x25x) & (!n_n76) & (x247x)) + ((n_n64) & (n_n100) & (!x25x) & (n_n76) & (!x247x)));
	assign x5967x = (((!i_3_) & (x19x) & (!x109x) & (x177x) & (!x129x)) + ((!i_3_) & (!x19x) & (x109x) & (!x177x) & (x129x)));
	assign x5968x = (((!i_6_) & (x76x) & (n_n63) & (!x110x) & (!x66x)) + ((i_6_) & (!x76x) & (!n_n63) & (x110x) & (x66x)));
	assign x5969x = (((n_n101) & (n_n100) & (n_n102) & (!n_n63) & (!n_n90)) + ((!n_n101) & (!n_n100) & (n_n102) & (n_n63) & (n_n90)));
	assign x5971x = (((!i_5_) & (!i_3_) & (!i_4_) & (x88x) & (!x20x)) + ((i_5_) & (i_3_) & (i_4_) & (!x88x) & (x20x)));
	assign x5972x = (((!n_n78) & (!x27x) & (n_n1193) & (!x1291x) & (!x1292x)) + ((!n_n78) & (!x27x) & (!n_n1193) & (x1291x) & (!x1292x)) + ((!n_n78) & (!x27x) & (!n_n1193) & (!x1291x) & (x1292x)) + ((n_n78) & (x27x) & (!n_n1193) & (!x1291x) & (!x1292x)));
	assign x5974x = (((!n_n78) & (!n_n102) & (!n_n85) & (n_n1297) & (!x220x)) + ((!n_n78) & (!n_n102) & (!n_n85) & (!n_n1297) & (x220x)) + ((n_n78) & (n_n102) & (n_n85) & (!n_n1297) & (!x220x)));
	assign x6360x = (((!n_n81) & (!n_n92) & (!x32x) & (!x37x) & (!x5969x)) + ((!n_n81) & (!n_n92) & (!x32x) & (!x37x) & (!x5969x)) + ((!n_n81) & (!n_n92) & (!x32x) & (!x37x) & (!x5969x)));
	assign x5996x = (((!i_8_) & (!i_4_) & (!n_n38) & (n_n1092) & (!x242x)) + ((!i_8_) & (!i_4_) & (n_n38) & (!n_n1092) & (x242x)));
	assign x6006x = (((i_2_) & (!n_n101) & (n_n78) & (n_n77) & (!x108x)) + ((!i_2_) & (n_n101) & (!n_n78) & (n_n77) & (x108x)));
	assign x6009x = (((!n_n91) & (!n_n102) & (!n_n97) & (n_n939) & (!x268x)) + ((!n_n91) & (!n_n102) & (!n_n97) & (!n_n939) & (x268x)) + ((n_n91) & (n_n102) & (n_n97) & (!n_n939) & (!x268x)));
	assign x6010x = (((!n_n101) & (!n_n74) & (!n_n90) & (x94x) & (!x1348x)) + ((!n_n101) & (!n_n74) & (!n_n90) & (!x94x) & (x1348x)) + ((n_n101) & (n_n74) & (n_n90) & (!x94x) & (!x1348x)));
	assign x6011x = (((!n_n86) & (!n_n97) & (!n_n77) & (n_n1128) & (!x5996x)) + ((!n_n86) & (!n_n97) & (!n_n77) & (!n_n1128) & (x5996x)) + ((n_n86) & (n_n97) & (n_n77) & (!n_n1128) & (!x5996x)));
	assign x6012x = (((!n_n83) & (x251x) & (!x321x) & (!n_n1176) & (!x320x)) + ((!n_n83) & (!x251x) & (x321x) & (!n_n1176) & (!x320x)) + ((!n_n83) & (!x251x) & (!x321x) & (n_n1176) & (!x320x)) + ((n_n83) & (!x251x) & (!x321x) & (!n_n1176) & (x320x)));
	assign x6013x = (((n_n969) & (!n_n1184) & (!n_n1156) & (!x5686x) & (!x5687x)) + ((!n_n969) & (n_n1184) & (!n_n1156) & (!x5686x) & (!x5687x)) + ((!n_n969) & (!n_n1184) & (n_n1156) & (!x5686x) & (!x5687x)) + ((!n_n969) & (!n_n1184) & (!n_n1156) & (x5686x) & (x5687x)));
	assign x6014x = (((!n_n78) & (n_n941) & (!x237x) & (!n_n1164) & (!n_n975)) + ((!n_n78) & (!n_n941) & (!x237x) & (n_n1164) & (!n_n975)) + ((!n_n78) & (!n_n941) & (!x237x) & (!n_n1164) & (n_n975)) + ((n_n78) & (!n_n941) & (x237x) & (!n_n1164) & (!n_n975)));
	assign x6015x = (((!n_n91) & (!x63x) & (!x83x) & (!x22x) & (n_n966)) + ((n_n91) & (x63x) & (!x83x) & (!x22x) & (!n_n966)) + ((n_n91) & (!x63x) & (x83x) & (!x22x) & (!n_n966)) + ((n_n91) & (!x63x) & (!x83x) & (x22x) & (!n_n966)));
	assign x6016x = (((!i_7_) & (!i_6_) & (!x21x) & (x336x) & (!x6006x)) + ((!i_7_) & (!i_6_) & (!x21x) & (!x336x) & (x6006x)) + ((!i_7_) & (i_6_) & (x21x) & (!x336x) & (!x6006x)));
	assign x6018x = (((!n_n70) & (!x53x) & (x215x) & (!x150x) & (!x153x)) + ((!n_n70) & (!x53x) & (!x215x) & (x150x) & (!x153x)) + ((!n_n70) & (!x53x) & (!x215x) & (!x150x) & (x153x)) + ((n_n70) & (x53x) & (!x215x) & (!x150x) & (!x153x)));

endmodule