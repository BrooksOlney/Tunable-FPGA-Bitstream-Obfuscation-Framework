module dsip (
	key<254>, key<253>, key<252>, key<251>, key<250>, key<249>, key<248>, key<246>, 
	key<245>, key<244>, key<243>, key<242>, key<241>, key<240>, key<238>, key<237>, key<235>, key<234>, 
	key<233>, key<232>, key<230>, key<229>, key<228>, key<227>, key<226>, key<225>, key<224>, key<222>, 
	key<221>, key<220>, key<219>, key<218>, key<217>, key<216>, key<214>, key<213>, key<212>, key<211>, 
	key<210>, key<209>, key<208>, key<206>, key<205>, key<204>, key<203>, key<202>, key<201>, key<200>, 
	key<198>, key<197>, key<196>, key<195>, key<194>, key<193>, key<192>, key<190>, key<189>, key<188>, 
	key<187>, key<186>, key<185>, key<184>, key<182>, key<181>, key<180>, key<179>, key<178>, key<177>, 
	key<176>, key<174>, key<173>, key<172>, key<171>, key<170>, key<169>, key<168>, key<166>, key<165>, 
	key<164>, key<163>, key<162>, key<161>, key<160>, key<158>, key<157>, key<156>, key<155>, key<154>, 
	key<153>, key<152>, key<150>, key<149>, key<148>, key<147>, key<146>, key<145>, key<144>, key<142>, 
	key<141>, key<140>, key<139>, key<138>, key<137>, key<136>, key<134>, key<133>, key<132>, key<131>, 
	key<130>, key<129>, key<128>, key<126>, key<125>, key<124>, key<123>, key<122>, key<121>, key<120>, 
	key<118>, key<117>, key<116>, key<115>, key<114>, key<113>, key<112>, key<110>, key<109>, key<107>, 
	key<106>, key<105>, key<104>, key<102>, key<101>, key<100>, key<99>, key<98>, key<97>, key<96>, 
	key<94>, key<93>, key<92>, key<91>, key<90>, key<89>, key<88>, key<86>, key<85>, key<84>, 
	key<83>, key<82>, key<81>, key<80>, key<78>, key<77>, key<76>, key<75>, key<74>, key<73>, 
	key<72>, key<70>, key<69>, key<68>, key<67>, key<66>, key<65>, key<64>, key<62>, key<61>, 
	key<60>, key<59>, key<58>, key<57>, key<56>, key<54>, key<53>, key<52>, key<51>, key<50>, 
	key<49>, key<48>, key<46>, key<45>, key<44>, key<43>, key<42>, key<41>, key<40>, key<38>, 
	key<37>, key<36>, key<35>, key<34>, key<33>, key<32>, key<30>, key<29>, key<28>, key<27>, 
	key<26>, key<25>, key<24>, key<22>, key<21>, key<20>, key<19>, key<18>, key<17>, key<16>, 
	key<14>, key<13>, key<12>, key<11>, key<10>, key<9>, key<8>, key<6>, key<5>, key<4>, 
	key<3>, key<2>, key<1>, key<0>, count<3>, count<2>, count<1>, count<0>, encrypt<0>, start<0>, 
	KSi<191>, KSi<190>, KSi<189>, KSi<188>, KSi<187>, KSi<186>, KSi<185>, KSi<184>, KSi<183>, KSi<182>, 
	KSi<181>, KSi<180>, KSi<179>, KSi<178>, KSi<177>, KSi<176>, KSi<175>, KSi<174>, KSi<173>, KSi<172>, 
	KSi<171>, KSi<170>, KSi<169>, KSi<168>, KSi<167>, KSi<166>, KSi<165>, KSi<164>, KSi<163>, KSi<162>, 
	KSi<161>, KSi<160>, KSi<159>, KSi<158>, KSi<157>, KSi<156>, KSi<155>, KSi<154>, KSi<153>, KSi<152>, 
	KSi<151>, KSi<150>, KSi<149>, KSi<148>, KSi<147>, KSi<146>, KSi<145>, KSi<144>, KSi<143>, KSi<142>, 
	KSi<141>, KSi<140>, KSi<139>, KSi<138>, KSi<137>, KSi<136>, KSi<135>, KSi<134>, KSi<133>, KSi<132>, 
	KSi<131>, KSi<130>, KSi<129>, KSi<128>, KSi<127>, KSi<126>, KSi<125>, KSi<124>, KSi<123>, KSi<122>, 
	KSi<121>, KSi<120>, KSi<119>, KSi<118>, KSi<117>, KSi<116>, KSi<115>, KSi<114>, KSi<113>, KSi<112>, 
	KSi<111>, KSi<110>, KSi<109>, KSi<108>, KSi<107>, KSi<106>, KSi<105>, KSi<104>, KSi<103>, KSi<102>, 
	KSi<101>, KSi<100>, KSi<99>, KSi<98>, KSi<97>, KSi<96>, KSi<95>, KSi<94>, KSi<93>, KSi<92>, 
	KSi<91>, KSi<90>, KSi<89>, KSi<88>, KSi<87>, KSi<86>, KSi<85>, KSi<84>, KSi<83>, KSi<82>, 
	KSi<81>, KSi<80>, KSi<79>, KSi<78>, KSi<77>, KSi<76>, KSi<75>, KSi<74>, KSi<73>, KSi<72>, 
	KSi<71>, KSi<70>, KSi<69>, KSi<68>, KSi<67>, KSi<66>, KSi<65>, KSi<64>, KSi<63>, KSi<62>, 
	KSi<61>, KSi<60>, KSi<59>, KSi<58>, KSi<57>, KSi<56>, KSi<55>, KSi<54>, KSi<53>, KSi<52>, 
	KSi<51>, KSi<50>, KSi<49>, KSi<48>, KSi<47>, KSi<46>, KSi<45>, KSi<44>, KSi<43>, KSi<42>, 
	KSi<41>, KSi<40>, KSi<39>, KSi<38>, KSi<37>, KSi<36>, KSi<35>, KSi<34>, KSi<33>, KSi<32>, 
	KSi<31>, KSi<30>, KSi<29>, KSi<28>, KSi<27>, KSi<26>, KSi<25>, KSi<24>, KSi<23>, KSi<22>, 
	KSi<21>, KSi<20>, KSi<19>, KSi<18>, KSi<17>, KSi<16>, KSi<15>, KSi<14>, KSi<13>, KSi<12>, 
	KSi<11>, KSi<10>, KSi<9>, KSi<8>, KSi<7>, KSi<6>, KSi<5>, KSi<4>, KSi<3>, KSi<2>, 
	KSi<1>, KSi<0>, new_count<3>, new_count<2>, new_count<1>, new_count<0>, data_ready<0>);

input key<254>, key<253>, key<252>, key<251>, key<250>, key<249>, key<248>, key<246>, key<245>, key<244>, key<243>, key<242>, key<241>, key<240>, key<238>, key<237>, key<235>, key<234>, key<233>, key<232>, key<230>, key<229>, key<228>, key<227>, key<226>, key<225>, key<224>, key<222>, key<221>, key<220>, key<219>, key<218>, key<217>, key<216>, key<214>, key<213>, key<212>, key<211>, key<210>, key<209>, key<208>, key<206>, key<205>, key<204>, key<203>, key<202>, key<201>, key<200>, key<198>, key<197>, key<196>, key<195>, key<194>, key<193>, key<192>, key<190>, key<189>, key<188>, key<187>, key<186>, key<185>, key<184>, key<182>, key<181>, key<180>, key<179>, key<178>, key<177>, key<176>, key<174>, key<173>, key<172>, key<171>, key<170>, key<169>, key<168>, key<166>, key<165>, key<164>, key<163>, key<162>, key<161>, key<160>, key<158>, key<157>, key<156>, key<155>, key<154>, key<153>, key<152>, key<150>, key<149>, key<148>, key<147>, key<146>, key<145>, key<144>, key<142>, key<141>, key<140>, key<139>, key<138>, key<137>, key<136>, key<134>, key<133>, key<132>, key<131>, key<130>, key<129>, key<128>, key<126>, key<125>, key<124>, key<123>, key<122>, key<121>, key<120>, key<118>, key<117>, key<116>, key<115>, key<114>, key<113>, key<112>, key<110>, key<109>, key<107>, key<106>, key<105>, key<104>, key<102>, key<101>, key<100>, key<99>, key<98>, key<97>, key<96>, key<94>, key<93>, key<92>, key<91>, key<90>, key<89>, key<88>, key<86>, key<85>, key<84>, key<83>, key<82>, key<81>, key<80>, key<78>, key<77>, key<76>, key<75>, key<74>, key<73>, key<72>, key<70>, key<69>, key<68>, key<67>, key<66>, key<65>, key<64>, key<62>, key<61>, key<60>, key<59>, key<58>, key<57>, key<56>, key<54>, key<53>, key<52>, key<51>, key<50>, key<49>, key<48>, key<46>, key<45>, key<44>, key<43>, key<42>, key<41>, key<40>, key<38>, key<37>, key<36>, key<35>, key<34>, key<33>, key<32>, key<30>, key<29>, key<28>, key<27>, key<26>, key<25>, key<24>, key<22>, key<21>, key<20>, key<19>, key<18>, key<17>, key<16>, key<14>, key<13>, key<12>, key<11>, key<10>, key<9>, key<8>, key<6>, key<5>, key<4>, key<3>, key<2>, key<1>, key<0>, count<3>, count<2>, count<1>, count<0>, encrypt<0>, start<0>;

output KSi<191>, KSi<190>, KSi<189>, KSi<188>, KSi<187>, KSi<186>, KSi<185>, KSi<184>, KSi<183>, KSi<182>, KSi<181>, KSi<180>, KSi<179>, KSi<178>, KSi<177>, KSi<176>, KSi<175>, KSi<174>, KSi<173>, KSi<172>, KSi<171>, KSi<170>, KSi<169>, KSi<168>, KSi<167>, KSi<166>, KSi<165>, KSi<164>, KSi<163>, KSi<162>, KSi<161>, KSi<160>, KSi<159>, KSi<158>, KSi<157>, KSi<156>, KSi<155>, KSi<154>, KSi<153>, KSi<152>, KSi<151>, KSi<150>, KSi<149>, KSi<148>, KSi<147>, KSi<146>, KSi<145>, KSi<144>, KSi<143>, KSi<142>, KSi<141>, KSi<140>, KSi<139>, KSi<138>, KSi<137>, KSi<136>, KSi<135>, KSi<134>, KSi<133>, KSi<132>, KSi<131>, KSi<130>, KSi<129>, KSi<128>, KSi<127>, KSi<126>, KSi<125>, KSi<124>, KSi<123>, KSi<122>, KSi<121>, KSi<120>, KSi<119>, KSi<118>, KSi<117>, KSi<116>, KSi<115>, KSi<114>, KSi<113>, KSi<112>, KSi<111>, KSi<110>, KSi<109>, KSi<108>, KSi<107>, KSi<106>, KSi<105>, KSi<104>, KSi<103>, KSi<102>, KSi<101>, KSi<100>, KSi<99>, KSi<98>, KSi<97>, KSi<96>, KSi<95>, KSi<94>, KSi<93>, KSi<92>, KSi<91>, KSi<90>, KSi<89>, KSi<88>, KSi<87>, KSi<86>, KSi<85>, KSi<84>, KSi<83>, KSi<82>, KSi<81>, KSi<80>, KSi<79>, KSi<78>, KSi<77>, KSi<76>, KSi<75>, KSi<74>, KSi<73>, KSi<72>, KSi<71>, KSi<70>, KSi<69>, KSi<68>, KSi<67>, KSi<66>, KSi<65>, KSi<64>, KSi<63>, KSi<62>, KSi<61>, KSi<60>, KSi<59>, KSi<58>, KSi<57>, KSi<56>, KSi<55>, KSi<54>, KSi<53>, KSi<52>, KSi<51>, KSi<50>, KSi<49>, KSi<48>, KSi<47>, KSi<46>, KSi<45>, KSi<44>, KSi<43>, KSi<42>, KSi<41>, KSi<40>, KSi<39>, KSi<38>, KSi<37>, KSi<36>, KSi<35>, KSi<34>, KSi<33>, KSi<32>, KSi<31>, KSi<30>, KSi<29>, KSi<28>, KSi<27>, KSi<26>, KSi<25>, KSi<24>, KSi<23>, KSi<22>, KSi<21>, KSi<20>, KSi<19>, KSi<18>, KSi<17>, KSi<16>, KSi<15>, KSi<14>, KSi<13>, KSi<12>, KSi<11>, KSi<10>, KSi<9>, KSi<8>, KSi<7>, KSi<6>, KSi<5>, KSi<4>, KSi<3>, KSi<2>, KSi<1>, KSi<0>, new_count<3>, new_count<2>, new_count<1>, new_count<0>, data_ready<0>;

wire wire7572, wire17163, wire7573, wire7574, wire7568, wire7575, I199, I200, wire7576, wire11699, main/$MINUS_4_1/c<0>8, wire7577, I205, main/$MINUS_4_1/c<0>8, wire17165, I208, wire7565, wire7580, wire17167, wire7566, wire7581, wire17157, wire17159, wire17161, wire7571, wire7586, wire14444, wire7587, I223, I224, I226, wire194, I228, I229, wire7541, wire7569, wire17145, wire17147, wire7591, wire7600, wire2074, wire7475, wire2079, wire7292, wire7284, I242, I243, wire7595, wire7597, wire7473, wire7598, wire7599, I249, I250, wire7606, wire2077, wire7560, wire7602, wire7603, wire7604, wire7605, I258, I259, new_C<111>, wire2068, wire7608, wire7609, I264, I265, wire7612, wire2071, wire7485, wire7611, I270, I271, new_C<110>, wire2062, wire7489, wire7614, I276, I277, wire7617, wire2065, wire7616, I281, I282, new_C<109>, wire2056, wire7480, wire7619, I287, I288, wire7622, wire2059, wire7621, I292, I293, new_C<108>, wire2050, wire7624, wire7625, I298, I299, wire7628, wire2053, wire7627, I303, I304, new_C<107>, wire2044, wire7482, wire7630, I309, I310, wire7633, wire2047, wire7632, I314, I315, new_C<106>, wire2038, wire7472, wire7635, I320, I321, wire7638, wire2041, wire7637, I325, I326, new_C<105>, wire2032, wire7479, wire7640, I331, I332, wire7643, wire2035, wire7642, I336, I337, new_C<104>, wire2026, wire7645, wire7646, I342, I343, wire7649, wire2029, wire7648, I347, I348, new_C<103>, wire2020, wire7491, wire7651, I353, I354, wire7654, wire2023, wire7653, I358, I359, new_C<102>, wire2014, wire7656, wire7657, I364, I365, wire7660, wire2017, wire7659, I369, I370, new_C<101>, wire2008, wire7484, wire7662, I375, I376, wire7665, wire2011, wire7664, I380, I381, new_C<100>, wire2002, wire7492, wire7667, I386, I387, wire7670, wire2005, wire7669, I391, I392, new_C<99>, wire1996, wire7471, wire7672, I397, I398, wire7675, wire1999, wire7674, I402, I403, new_C<98>, wire1990, wire7478, wire7677, I408, I409, wire7680, wire1993, wire7679, I413, I414, new_C<97>, wire1984, wire7490, wire7682, I419, I420, wire7685, wire1987, wire7684, I424, I425, new_C<96>, wire1978, wire7481, wire7687, I430, I431, wire7690, wire1981, wire7689, I435, I436, new_C<95>, wire1972, wire7692, wire7693, I441, I442, wire7696, wire1975, wire7695, I446, I447, new_C<94>, wire1966, wire7476, wire7698, I452, I453, wire7701, wire1969, wire7700, I457, I458, new_C<93>, wire1960, wire7474, wire7703, I463, I464, wire7706, wire1963, wire7705, I468, I469, new_C<92>, wire1954, wire7483, wire7708, I474, I475, wire7711, wire1957, wire7710, I479, I480, new_C<91>, wire1948, wire7487, wire7713, I485, I486, wire7716, wire1951, wire7715, I490, I491, new_C<90>, wire1942, wire7477, wire7718, I496, I497, wire7721, wire1945, wire7720, I501, I502, new_C<89>, wire1936, wire7486, wire7723, I507, I508, wire7726, wire1939, wire7725, I512, I513, new_C<88>, wire1930, wire7470, wire7728, I518, I519, wire7731, wire1933, wire7730, I523, I524, new_C<87>, wire1924, wire7488, wire7733, I529, I530, wire7736, wire1927, wire7735, I534, I535, new_C<86>, wire1918, wire7509, wire7738, I540, I541, wire7741, wire1921, wire7740, I545, I546, new_C<85>, wire1912, wire7496, wire7743, I551, I552, wire7746, wire1915, wire7745, I556, I557, new_C<84>, wire1906, wire7500, wire7748, I562, I563, wire7751, wire1909, wire7750, I567, I568, new_C<83>, wire1900, wire7753, wire7754, I573, I574, wire7757, wire1903, wire7756, I578, I579, new_C<82>, wire1894, wire7513, wire7759, I584, I585, wire7762, wire1897, wire7761, I589, I590, new_C<81>, wire1888, wire7504, wire7764, I595, I596, wire7767, wire1891, wire7766, I600, I601, new_C<80>, wire1882, wire7769, wire7770, I606, I607, wire7773, wire1885, wire7772, I611, I612, new_C<79>, wire1876, wire7506, wire7775, I617, I618, wire7778, wire1879, wire7777, I622, I623, new_C<78>, wire1870, wire7495, wire7780, I628, I629, wire7783, wire1873, wire7782, I633, I634, new_C<77>, wire1864, wire7503, wire7785, I639, I640, wire7788, wire1867, wire7787, I644, I645, new_C<76>, wire1858, wire7790, wire7791, I650, I651, wire7794, wire1861, wire7793, I655, I656, new_C<75>, wire1852, wire7515, wire7796, I661, I662, wire7799, wire1855, wire7798, I666, I667, new_C<74>, wire1846, wire7498, wire7801, I672, I673, wire7804, wire1849, wire7803, I677, I678, new_C<73>, wire1840, wire7508, wire7806, I683, I684, wire7809, wire1843, wire7808, I688, I689, new_C<72>, wire1834, wire7516, wire7811, I694, I695, wire7814, wire1837, wire7813, I699, I700, new_C<71>, wire1828, wire7494, wire7816, I705, I706, wire7819, wire1831, wire7818, I710, I711, new_C<70>, wire1822, wire7502, wire7821, I716, I717, wire7824, wire1825, wire7823, I721, I722, new_C<69>, wire1816, wire7514, wire7826, I727, I728, wire7829, wire1819, wire7828, I732, I733, new_C<68>, wire1810, wire7505, wire7831, I738, I739, wire7834, wire1813, wire7833, I743, I744, new_C<67>, wire1804, wire7836, wire7837, I749, I750, wire7840, wire1807, wire7839, I754, I755, new_C<66>, wire1798, wire7499, wire7842, I760, I761, wire7845, wire1801, wire7844, I765, I766, new_C<65>, wire1792, wire7497, wire7847, I771, I772, wire7850, wire1795, wire7849, I776, I777, new_C<64>, wire1786, wire7507, wire7852, I782, I783, wire7855, wire1789, wire7854, I787, I788, new_C<63>, wire1780, wire7511, wire7857, I793, I794, wire7860, wire1783, wire7859, I798, I799, new_C<62>, wire1774, wire7501, wire7862, I804, I805, wire7865, wire1777, wire7864, I809, I810, new_C<61>, wire1768, wire7510, wire7867, I815, I816, wire7870, wire1771, wire7869, I820, I821, new_C<60>, wire1762, wire7493, wire7872, I826, I827, wire7875, wire1765, wire7874, I831, I832, new_C<59>, wire1756, wire7512, wire7877, I837, I838, wire7880, wire1759, wire7879, I842, I843, new_C<58>, wire1750, wire7533, wire7882, I848, I849, wire7885, wire1753, wire7884, I853, I854, new_C<57>, wire1744, wire7520, wire7887, I859, I860, wire7890, wire1747, wire7889, I864, I865, new_C<56>, wire1738, wire7524, wire7892, I870, I871, wire7895, wire1741, wire7894, I875, I876, new_C<55>, wire1732, wire7897, wire7898, I881, I882, wire7901, wire1735, wire7900, I886, I887, new_C<54>, wire1726, wire7537, wire7903, I892, I893, wire7906, wire1729, wire7905, I897, I898, new_C<53>, wire1720, wire7528, wire7908, I903, I904, wire7911, wire1723, wire7910, I908, I909, new_C<52>, wire1714, wire7913, wire7914, I914, I915, wire7917, wire1717, wire7916, I919, I920, new_C<51>, wire1708, wire7530, wire7919, I925, I926, wire7922, wire1711, wire7921, I930, I931, new_C<50>, wire1702, wire7519, wire7924, I936, I937, wire7927, wire1705, wire7926, I941, I942, new_C<49>, wire1696, wire7527, wire7929, I947, I948, wire7932, wire1699, wire7931, I952, I953, new_C<48>, wire1690, wire7934, wire7935, I958, I959, wire7938, wire1693, wire7937, I963, I964, new_C<47>, wire1684, wire7539, wire7940, I969, I970, wire7943, wire1687, wire7942, I974, I975, new_C<46>, wire1678, wire7522, wire7945, I980, I981, wire7948, wire1681, wire7947, I985, I986, new_C<45>, wire1672, wire7532, wire7950, I991, I992, wire7953, wire1675, wire7952, I996, I997, new_C<44>, wire1666, wire7540, wire7955, I1002, I1003, wire7958, wire1669, wire7957, I1007, I1008, new_C<43>, wire1660, wire7518, wire7960, I1013, I1014, wire7963, wire1663, wire7962, I1018, I1019, new_C<42>, wire1654, wire7526, wire7965, I1024, I1025, wire7968, wire1657, wire7967, I1029, I1030, new_C<41>, wire1648, wire7538, wire7970, I1035, I1036, wire7973, wire1651, wire7972, I1040, I1041, new_C<40>, wire1642, wire7529, wire7975, I1046, I1047, wire7978, wire1645, wire7977, I1051, I1052, new_C<39>, wire1636, wire7980, wire7981, I1057, I1058, wire7984, wire1639, wire7983, I1062, I1063, new_C<38>, wire1630, wire7523, wire7986, I1068, I1069, wire7989, wire1633, wire7988, I1073, I1074, new_C<37>, wire1624, wire7521, wire7991, I1079, I1080, wire7994, wire1627, wire7993, I1084, I1085, new_C<36>, wire1618, wire7531, wire7996, I1090, I1091, wire7999, wire1621, wire7998, I1095, I1096, new_C<35>, wire1612, wire7535, wire8001, I1101, I1102, wire8004, wire1615, wire8003, I1106, I1107, new_C<34>, wire1606, wire7525, wire8006, I1112, I1113, wire8009, wire1609, wire8008, I1117, I1118, new_C<33>, wire1600, wire7534, wire8011, I1123, I1124, wire8014, wire1603, wire8013, I1128, I1129, new_C<32>, wire1594, wire7517, wire8016, I1134, I1135, wire8019, wire1597, wire8018, I1139, I1140, new_C<31>, wire1588, wire7536, wire8021, I1145, I1146, wire8024, wire1591, wire8023, I1150, I1151, new_C<30>, wire1582, wire7557, wire8026, I1156, I1157, wire8029, wire1585, wire8028, I1161, I1162, new_C<29>, wire1576, wire7544, wire8031, I1167, I1168, wire8034, wire1579, wire8033, I1172, I1173, new_C<28>, wire1570, wire7548, wire8036, I1178, I1179, wire8039, wire1573, wire8038, I1183, I1184, new_C<27>, wire1564, wire8041, wire8042, I1189, I1190, wire8045, wire1567, wire8044, I1194, I1195, new_C<26>, wire1558, wire7561, wire8047, I1200, I1201, wire8050, wire1561, wire8049, I1205, I1206, new_C<25>, wire1552, wire7552, wire8052, I1211, I1212, wire8055, wire1555, wire8054, I1216, I1217, new_C<24>, wire1546, wire8057, wire8058, I1222, I1223, wire8061, wire1549, wire8060, I1227, I1228, new_C<23>, wire1540, wire7554, wire8063, I1233, I1234, wire8066, wire1543, wire8065, I1238, I1239, new_C<22>, wire1534, wire7543, wire8068, I1244, I1245, wire8071, wire1537, wire8070, I1249, I1250, new_C<21>, wire1528, wire7551, wire8073, I1255, I1256, wire8076, wire1531, wire8075, I1260, I1261, new_C<20>, wire1522, wire8078, wire8079, I1266, I1267, wire8082, wire1525, wire8081, I1271, I1272, new_C<19>, wire1516, wire7563, wire8084, I1277, I1278, wire8087, wire1519, wire8086, I1282, I1283, new_C<18>, wire1510, wire7546, wire8089, I1288, I1289, wire8092, wire1513, wire8091, I1293, I1294, new_C<17>, wire1504, wire7556, wire8094, I1299, I1300, wire8097, wire1507, wire8096, I1304, I1305, new_C<16>, wire1498, wire7564, wire8099, I1310, I1311, wire8102, wire1501, wire8101, I1315, I1316, new_C<15>, wire1492, wire7542, wire8104, I1321, I1322, wire8107, wire1495, wire8106, I1326, I1327, new_C<14>, wire1486, wire7550, wire8109, I1332, I1333, wire8112, wire1489, wire8111, I1337, I1338, new_C<13>, wire1480, wire7562, wire8114, I1343, I1344, wire8117, wire1483, wire8116, I1348, I1349, new_C<12>, wire1474, wire7553, wire8119, I1354, I1355, wire8122, wire1477, wire8121, I1359, I1360, new_C<11>, wire1468, wire8124, wire8125, I1365, I1366, wire8128, wire1471, wire8127, I1370, I1371, new_C<10>, wire1462, wire7547, wire8130, I1376, I1377, wire8133, wire1465, wire8132, I1381, I1382, new_C<9>, wire1456, wire7545, wire8135, I1387, I1388, wire8138, wire1459, wire8137, I1392, I1393, new_C<8>, wire1450, wire7555, wire8140, I1398, I1399, wire8143, wire1453, wire8142, I1403, I1404, new_C<7>, wire1444, wire7559, wire8145, I1409, I1410, wire8148, wire1447, wire8147, I1414, I1415, new_C<6>, wire1438, wire7549, wire8150, I1420, I1421, wire8153, wire1441, wire8152, I1425, I1426, new_C<5>, wire1432, wire7558, wire8155, I1431, I1432, wire8158, wire1435, wire8157, I1436, I1437, new_C<4>, wire1426, wire8160, I1441, I1442, wire8163, wire1429, wire8162, I1446, I1447, new_C<3>, wire1420, wire8165, I1451, I1452, wire8168, wire1423, wire8167, I1456, I1457, new_C<2>, wire1414, wire8170, I1461, I1462, wire8173, wire1417, wire8172, I1466, I1467, new_C<1>, wire1408, wire8175, I1471, I1472, wire1411, wire8177, I1475, I1476, new_C<0>, wire7463, wire1402, wire8179, wire7394, wire8180, I1483, I1484, wire8184, wire1405, wire7447, wire8182, wire8183, I1490, I1491, new_D<111>, wire1396, wire7382, wire8186, I1496, I1497, wire8189, wire1399, wire7384, wire8188, I1502, I1503, new_D<110>, wire1390, wire7398, wire8191, I1508, I1509, wire8194, wire1393, wire8193, I1513, I1514, new_D<109>, wire1384, wire7391, wire8196, I1519, I1520, wire8199, wire1387, wire8198, I1524, I1525, new_D<108>, wire1378, wire7380, wire8201, I1530, I1531, wire8204, wire1381, wire8203, I1535, I1536, new_D<107>, wire1372, wire7386, wire8206, I1541, I1542, wire8209, wire1375, wire8208, I1546, I1547, new_D<106>, wire1366, wire7388, wire8211, I1552, I1553, wire8214, wire1369, wire8213, I1557, I1558, new_D<105>, wire1360, wire7395, wire8216, I1563, I1564, wire8219, wire1363, wire8218, I1568, I1569, new_D<104>, wire1354, wire7381, wire8221, I1574, I1575, wire8224, wire1357, wire8223, I1579, I1580, new_D<103>, wire1348, wire7390, wire8226, I1585, I1586, wire8229, wire1351, wire8228, I1590, I1591, new_D<102>, wire1342, wire7387, wire8231, I1596, I1597, wire8234, wire1345, wire8233, I1601, I1602, new_D<101>, wire1336, wire8236, wire8237, I1607, I1608, wire8240, wire1339, wire8239, I1612, I1613, new_D<100>, wire1330, wire8242, wire8243, I1618, I1619, wire8246, wire1333, wire8245, I1623, I1624, new_D<99>, wire1324, wire8248, wire8249, I1629, I1630, wire8252, wire1327, wire8251, I1634, I1635, new_D<98>, wire1318, wire7392, wire8254, I1640, I1641, wire8257, wire1321, wire8256, I1645, I1646, new_D<97>, wire1312, wire7385, wire8259, I1651, I1652, wire8262, wire1315, wire8261, I1656, I1657, new_D<96>, wire1306, wire8264, wire8265, I1662, I1663, wire8268, wire1309, wire8267, I1667, I1668, new_D<95>, wire1300, wire7396, wire8270, I1673, I1674, wire8273, wire1303, wire8272, I1678, I1679, new_D<94>, wire1294, wire7379, wire8275, I1684, I1685, wire8278, wire1297, wire8277, I1689, I1690, new_D<93>, wire1288, wire8280, wire8281, I1695, I1696, wire8284, wire1291, wire8283, I1700, I1701, new_D<92>, wire1282, wire7383, wire8286, I1706, I1707, wire8289, wire1285, wire8288, I1711, I1712, new_D<91>, wire1276, wire7389, wire8291, I1717, I1718, wire8294, wire1279, wire8293, I1722, I1723, new_D<90>, wire1270, wire7377, wire8296, I1728, I1729, wire8299, wire1273, wire8298, I1733, I1734, new_D<89>, wire1264, wire7397, wire8301, I1739, I1740, wire8304, wire1267, wire8303, I1744, I1745, new_D<88>, wire1258, wire7393, wire8306, I1750, I1751, wire8309, wire1261, wire8308, I1755, I1756, new_D<87>, wire1252, wire7378, wire8311, I1761, I1762, wire8314, wire1255, wire8313, I1766, I1767, new_D<86>, wire1246, wire7407, wire8316, I1772, I1773, wire8319, wire1249, wire8318, I1777, I1778, new_D<85>, wire1240, wire7417, wire8321, I1783, I1784, wire8324, wire1243, wire8323, I1788, I1789, new_D<84>, wire1234, wire8326, wire8327, I1794, I1795, wire8330, wire1237, wire8329, I1799, I1800, new_D<83>, wire1228, wire7405, wire8332, I1805, I1806, wire8335, wire1231, wire8334, I1810, I1811, new_D<82>, wire1222, wire7421, wire8337, I1816, I1817, wire8340, wire1225, wire8339, I1821, I1822, new_D<81>, wire1216, wire7414, wire8342, I1827, I1828, wire8345, wire1219, wire8344, I1832, I1833, new_D<80>, wire1210, wire7402, wire8347, I1838, I1839, wire8350, wire1213, wire8349, I1843, I1844, new_D<79>, wire1204, wire7409, wire8352, I1849, I1850, wire8355, wire1207, wire8354, I1854, I1855, new_D<78>, wire1198, wire7411, wire8357, I1860, I1861, wire8360, wire1201, wire8359, I1865, I1866, new_D<77>, wire1192, wire7418, wire8362, I1871, I1872, wire8365, wire1195, wire8364, I1876, I1877, new_D<76>, wire1186, wire7404, wire8367, I1882, I1883, wire8370, wire1189, wire8369, I1887, I1888, new_D<75>, wire1180, wire8372, wire8373, I1893, I1894, wire1183, wire8375, I1897, I1898, new_D<74>, wire1174, wire7410, wire8377, I1903, I1904, wire8380, wire1177, wire8379, I1908, I1909, new_D<73>, wire1168, wire7413, wire8382, I1914, I1915, wire8385, wire1171, wire8384, I1919, I1920, new_D<72>, wire1162, wire7403, wire8387, I1925, I1926, wire8390, wire1165, wire8389, I1930, I1931, new_D<71>, wire1156, wire7422, wire8392, I1936, I1937, wire8395, wire1159, wire8394, I1941, I1942, new_D<70>, wire1150, wire7415, wire8397, I1947, I1948, wire8400, wire1153, wire8399, I1952, I1953, new_D<69>, wire1144, wire7408, wire8402, I1958, I1959, wire8405, wire1147, wire8404, I1963, I1964, new_D<68>, wire1138, wire8407, wire8408, I1969, I1970, wire8411, wire1141, wire8410, I1974, I1975, new_D<67>, wire1132, wire7419, wire8413, I1980, I1981, wire8416, wire1135, wire8415, I1985, I1986, new_D<66>, wire1126, wire7401, wire8418, I1991, I1992, wire8421, wire1129, wire8420, I1996, I1997, new_D<65>, wire1120, wire8423, wire8424, I2002, I2003, wire8427, wire1123, wire8426, I2007, I2008, new_D<64>, wire1114, wire7406, wire8429, I2013, I2014, wire8432, wire1117, wire8431, I2018, I2019, new_D<63>, wire1108, wire7412, wire8434, I2024, I2025, wire8437, wire1111, wire8436, I2029, I2030, new_D<62>, wire1102, wire7399, wire8439, I2035, I2036, wire8442, wire1105, wire8441, I2040, I2041, new_D<61>, wire1096, wire7420, wire8444, I2046, I2047, wire8447, wire1099, wire8446, I2051, I2052, new_D<60>, wire1090, wire7416, wire8449, I2057, I2058, wire8452, wire1093, wire8451, I2062, I2063, new_D<59>, wire1084, wire7400, wire8454, I2068, I2069, wire8457, wire1087, wire8456, I2073, I2074, new_D<58>, wire1078, wire7430, wire8459, I2079, I2080, wire8462, wire1081, wire8461, I2084, I2085, new_D<57>, wire1072, wire7440, wire8464, I2090, I2091, wire8467, wire1075, wire8466, I2095, I2096, new_D<56>, wire1066, wire8469, wire8470, I2101, I2102, wire8473, wire1069, wire8472, I2106, I2107, new_D<55>, wire1060, wire7428, wire8475, I2112, I2113, wire8478, wire1063, wire8477, I2117, I2118, new_D<54>, wire1054, wire7444, wire8480, I2123, I2124, wire8483, wire1057, wire8482, I2128, I2129, new_D<53>, wire1048, wire7437, wire8485, I2134, I2135, wire8488, wire1051, wire8487, I2139, I2140, new_D<52>, wire1042, wire7426, wire8490, I2145, I2146, wire8493, wire1045, wire8492, I2150, I2151, new_D<51>, wire1036, wire7432, wire8495, I2156, I2157, wire8498, wire1039, wire8497, I2161, I2162, new_D<50>, wire1030, wire7434, wire8500, I2167, I2168, wire8503, wire1033, wire8502, I2172, I2173, new_D<49>, wire1024, wire7441, wire8505, I2178, I2179, wire8508, wire1027, wire8507, I2183, I2184, new_D<48>, wire1018, wire7427, wire8510, I2189, I2190, wire8513, wire1021, wire8512, I2194, I2195, new_D<47>, wire1012, wire7436, wire8515, I2200, I2201, wire8518, wire1015, wire8517, I2205, I2206, new_D<46>, wire1006, wire7433, wire8520, I2211, I2212, wire8523, wire1009, wire8522, I2216, I2217, new_D<45>, wire1000, wire8525, wire8526, I2222, I2223, wire8529, wire1003, wire8528, I2227, I2228, new_D<44>, wire994, wire8531, wire8532, I2233, I2234, wire8535, wire997, wire8534, I2238, I2239, new_D<43>, wire988, wire7445, wire8537, I2244, I2245, wire8540, wire991, wire8539, I2249, I2250, new_D<42>, wire982, wire7438, wire8542, I2255, I2256, wire8545, wire985, wire8544, I2260, I2261, new_D<41>, wire976, wire7431, wire8547, I2266, I2267, wire8550, wire979, wire8549, I2271, I2272, new_D<40>, wire970, wire8552, wire8553, I2277, I2278, wire8556, wire973, wire8555, I2282, I2283, new_D<39>, wire964, wire7442, wire8558, I2288, I2289, wire8561, wire967, wire8560, I2293, I2294, new_D<38>, wire958, wire7425, wire8563, I2299, I2300, wire8566, wire961, wire8565, I2304, I2305, new_D<37>, wire952, wire8568, wire8569, I2310, I2311, wire8572, wire955, wire8571, I2315, I2316, new_D<36>, wire946, wire7429, wire8574, I2321, I2322, wire8577, wire949, wire8576, I2326, I2327, new_D<35>, wire940, wire7435, wire8579, I2332, I2333, wire8582, wire943, wire8581, I2337, I2338, new_D<34>, wire934, wire7423, wire8584, I2343, I2344, wire8587, wire937, wire8586, I2348, I2349, new_D<33>, wire928, wire7443, wire8589, I2354, I2355, wire8592, wire931, wire8591, I2359, I2360, new_D<32>, wire922, wire7439, wire8594, I2365, I2366, wire8597, wire925, wire8596, I2370, I2371, new_D<31>, wire916, wire7424, wire8599, I2376, I2377, wire8602, wire919, wire8601, I2381, I2382, new_D<30>, wire910, wire7454, wire8604, I2387, I2388, wire8607, wire913, wire8606, I2392, I2393, new_D<29>, wire904, wire7464, wire8609, I2398, I2399, wire8612, wire907, wire8611, I2403, I2404, new_D<28>, wire898, wire8614, wire8615, I2409, I2410, wire8618, wire901, wire8617, I2414, I2415, new_D<27>, wire892, wire7452, wire8620, I2420, I2421, wire8623, wire895, wire8622, I2425, I2426, new_D<26>, wire886, wire7468, wire8625, I2431, I2432, wire8628, wire889, wire8627, I2436, I2437, new_D<25>, wire880, wire7461, wire8630, I2442, I2443, wire8633, wire883, wire8632, I2447, I2448, new_D<24>, wire874, wire7449, wire8635, I2453, I2454, wire8638, wire877, wire8637, I2458, I2459, new_D<23>, wire868, wire7456, wire8640, I2464, I2465, wire8643, wire871, wire8642, I2469, I2470, new_D<22>, wire862, wire7458, wire8645, I2475, I2476, wire8648, wire865, wire8647, I2480, I2481, new_D<21>, wire856, wire7465, wire8650, I2486, I2487, wire8653, wire859, wire8652, I2491, I2492, new_D<20>, wire850, wire7451, wire8655, I2497, I2498, wire8658, wire853, wire8657, I2502, I2503, new_D<19>, wire844, wire7460, wire8660, I2508, I2509, wire847, wire8662, I2512, I2513, new_D<18>, wire838, wire7457, wire8664, I2518, I2519, wire8667, wire841, wire8666, I2523, I2524, new_D<17>, wire832, wire8669, wire8670, I2529, I2530, wire8673, wire835, wire8672, I2534, I2535, new_D<16>, wire826, wire7450, wire8675, I2540, I2541, wire8678, wire829, wire8677, I2545, I2546, new_D<15>, wire820, wire7469, wire8680, I2551, I2552, wire8683, wire823, wire8682, I2556, I2557, new_D<14>, wire814, wire7462, wire8685, I2562, I2563, wire8688, wire817, wire8687, I2567, I2568, new_D<13>, wire808, wire7455, wire8690, I2573, I2574, wire8693, wire811, wire8692, I2578, I2579, new_D<12>, wire802, wire8695, wire8696, I2584, I2585, wire8699, wire805, wire8698, I2589, I2590, new_D<11>, wire796, wire7466, wire8701, I2595, I2596, wire8704, wire799, wire8703, I2600, I2601, new_D<10>, wire790, wire7448, wire8706, I2606, I2607, wire8709, wire793, wire8708, I2611, I2612, new_D<9>, wire784, wire8711, wire8712, I2617, I2618, wire8715, wire787, wire8714, I2622, I2623, new_D<8>, wire778, wire7453, wire8717, I2628, I2629, wire8720, wire781, wire8719, I2633, I2634, new_D<7>, wire772, wire7459, wire8722, I2639, I2640, wire8725, wire775, wire8724, I2644, I2645, new_D<6>, wire766, wire7446, wire8727, I2650, I2651, wire8730, wire769, wire8729, I2655, I2656, new_D<5>, wire760, wire7467, wire8732, I2661, I2662, wire8735, wire763, wire8734, I2666, I2667, new_D<4>, wire754, wire8737, I2671, I2672, wire8740, wire757, wire8739, I2676, I2677, new_D<3>, wire748, wire8742, I2681, I2682, wire8745, wire751, wire8744, I2686, I2687, new_D<2>, wire742, wire8747, I2691, I2692, wire8750, wire745, wire8749, I2696, I2697, new_D<1>, wire736, wire8752, I2701, I2702, wire739, wire8754, I2705, I2706, new_D<0>, wire7596, wire7570, wire8756, wire8757, I2713, I2714, start<0>*, wire7573*, encrypt<0>*, count<2>*, wire7574*, wire7568*, count<0>*, count<1>*, wire7576*, wire11699*, main/$MINUS_4_1/c<0>8, count<3>*, wire7575*, wire7577*, wire7565*, wire7566*, wire17163*, wire17165*, wire17167*, wire7581*, wire17157*, wire17159*, wire17161*, wire7571*, wire7586*, wire14444*, wire7587*, new_count<0>*, wire194*, C<1>*, wire7569*, wire7580*, wire17145*, wire17147*, wire7541*, wire7600*, C<109>*, wire7591*, wire2079*, wire7292*, wire7572*, wire7284*, C<110>*, wire7595*, wire7475*, wire7597*, wire7473*, wire7598*, key<227>*, wire7606*, C<0>*, key<56>*, wire7560*, wire7602*, wire7603*, wire7604*, C<108>*, wire7608*, key<235>*, wire7612*, C<111>*, wire7485*, C<107>*, wire7489*, key<243>*, wire7617*, C<106>*, wire7480*, key<251>*, wire7622*, C<105>*, wire7624*, key<194>*, wire7628*, C<104>*, wire7482*, key<202>*, wire7633*, C<103>*, wire7472*, key<210>*, wire7638*, C<102>*, wire7479*, key<218>*, wire7643*, C<101>*, wire7645*, key<226>*, wire7649*, C<100>*, wire7491*, key<234>*, wire7654*, C<99>*, wire7656*, key<242>*, wire7660*, C<98>*, wire7484*, key<250>*, wire7665*, C<97>*, wire7492*, key<193>*, wire7670*, C<96>*, wire7471*, key<201>*, wire7675*, C<95>*, wire7478*, key<209>*, wire7680*, C<94>*, wire7490*, key<217>*, wire7685*, C<93>*, wire7481*, key<225>*, wire7690*, C<92>*, wire7692*, key<233>*, wire7696*, C<91>*, wire7476*, key<241>*, wire7701*, C<90>*, wire7474*, key<249>*, wire7706*, C<89>*, wire7483*, key<192>*, wire7711*, C<88>*, wire7487*, key<200>*, wire7716*, C<87>*, wire7477*, key<208>*, wire7721*, C<86>*, wire7486*, key<216>*, wire7726*, C<85>*, wire7470*, key<224>*, wire7731*, C<84>*, wire7488*, key<232>*, wire7736*, C<83>*, wire7509*, key<240>*, wire7741*, C<82>*, wire7496*, key<248>*, wire7746*, C<81>*, wire7500*, key<163>*, wire7751*, C<80>*, wire7753*, key<171>*, wire7757*, C<79>*, wire7513*, key<179>*, wire7762*, C<78>*, wire7504*, key<187>*, wire7767*, C<77>*, wire7769*, key<130>*, wire7773*, C<76>*, wire7506*, key<138>*, wire7778*, C<75>*, wire7495*, key<146>*, wire7783*, C<74>*, wire7503*, key<154>*, wire7788*, C<73>*, wire7790*, key<162>*, wire7794*, C<72>*, wire7515*, key<170>*, wire7799*, C<71>*, wire7498*, key<178>*, wire7804*, C<70>*, wire7508*, key<186>*, wire7809*, C<69>*, wire7516*, key<129>*, wire7814*, C<68>*, wire7494*, key<137>*, wire7819*, C<67>*, wire7502*, key<145>*, wire7824*, C<66>*, wire7514*, key<153>*, wire7829*, C<65>*, wire7505*, key<161>*, wire7834*, C<64>*, wire7836*, key<169>*, wire7840*, C<63>*, wire7499*, key<177>*, wire7845*, C<62>*, wire7497*, key<185>*, wire7850*, C<61>*, wire7507*, key<128>*, wire7855*, C<60>*, wire7511*, key<136>*, wire7860*, C<59>*, wire7501*, key<144>*, wire7865*, C<58>*, wire7510*, key<152>*, wire7870*, C<57>*, wire7493*, key<160>*, wire7875*, C<56>*, wire7512*, key<168>*, wire7880*, C<55>*, wire7533*, key<176>*, wire7885*, C<54>*, wire7520*, key<184>*, wire7890*, C<53>*, wire7524*, key<99>*, wire7895*, C<52>*, wire7897*, key<107>*, wire7901*, C<51>*, wire7537*, key<115>*, wire7906*, C<50>*, wire7528*, key<123>*, wire7911*, C<49>*, wire7913*, key<66>*, wire7917*, C<48>*, wire7530*, key<74>*, wire7922*, C<47>*, wire7519*, key<82>*, wire7927*, C<46>*, wire7527*, key<90>*, wire7932*, C<45>*, wire7934*, key<98>*, wire7938*, C<44>*, wire7539*, key<106>*, wire7943*, C<43>*, wire7522*, key<114>*, wire7948*, C<42>*, wire7532*, key<122>*, wire7953*, C<41>*, wire7540*, key<65>*, wire7958*, C<40>*, wire7518*, key<73>*, wire7963*, C<39>*, wire7526*, key<81>*, wire7968*, C<38>*, wire7538*, key<89>*, wire7973*, C<37>*, wire7529*, key<97>*, wire7978*, C<36>*, wire7980*, key<105>*, wire7984*, C<35>*, wire7523*, key<113>*, wire7989*, C<34>*, wire7521*, key<121>*, wire7994*, C<33>*, wire7531*, key<64>*, wire7999*, C<32>*, wire7535*, key<72>*, wire8004*, C<31>*, wire7525*, key<80>*, wire8009*, C<30>*, wire7534*, key<88>*, wire8014*, C<29>*, wire7517*, key<96>*, wire8019*, C<28>*, wire7536*, key<104>*, wire8024*, C<27>*, wire7557*, key<112>*, wire8029*, C<26>*, wire7544*, key<120>*, wire8034*, C<25>*, wire7548*, key<35>*, wire8039*, C<24>*, wire8041*, key<43>*, wire8045*, C<23>*, wire7561*, key<51>*, wire8050*, C<22>*, wire7552*, key<59>*, wire8055*, C<21>*, wire8057*, key<2>*, wire8061*, C<20>*, wire7554*, key<10>*, wire8066*, C<19>*, wire7543*, key<18>*, wire8071*, C<18>*, wire7551*, key<26>*, wire8076*, C<17>*, wire8078*, key<34>*, wire8082*, C<16>*, wire7563*, key<42>*, wire8087*, C<15>*, wire7546*, key<50>*, wire8092*, C<14>*, wire7556*, key<58>*, wire8097*, C<13>*, wire7564*, key<1>*, wire8102*, C<12>*, wire7542*, key<9>*, wire8107*, C<11>*, wire7550*, key<17>*, wire8112*, C<10>*, wire7562*, key<25>*, wire8117*, C<9>*, wire7553*, key<33>*, wire8122*, C<8>*, wire8124*, key<41>*, wire8128*, C<7>*, wire7547*, key<49>*, wire8133*, C<6>*, wire7545*, key<57>*, wire8138*, C<5>*, wire7555*, key<0>*, wire8143*, C<4>*, wire7559*, key<8>*, wire8148*, C<3>*, wire7549*, key<16>*, wire8153*, C<2>*, wire7558*, key<24>*, wire8158*, key<32>*, wire8163*, key<40>*, wire8168*, key<48>*, wire8173*, D<1>*, wire7463*, D<109>*, D<110>*, wire8179*, wire7394*, key<195>*, wire8184*, D<0>*, key<62>*, wire7447*, wire8182*, D<108>*, wire7382*, key<203>*, wire8189*, D<111>*, wire7384*, D<107>*, wire7398*, key<211>*, wire8194*, D<106>*, wire7391*, key<219>*, wire8199*, D<105>*, wire7380*, key<196>*, wire8204*, D<104>*, wire7386*, key<204>*, wire8209*, D<103>*, wire7388*, key<212>*, wire8214*, D<102>*, wire7395*, key<220>*, wire8219*, D<101>*, wire7381*, key<228>*, wire8224*, D<100>*, wire7390*, key<172>*, wire8229*, D<99>*, wire7387*, key<244>*, wire8234*, D<98>*, wire8236*, key<252>*, wire8240*, D<97>*, wire8242*, key<197>*, wire8246*, D<96>*, wire8248*, key<205>*, wire8252*, D<95>*, wire7392*, key<213>*, wire8257*, D<94>*, wire7385*, key<221>*, wire8262*, D<93>*, wire8264*, key<229>*, wire8268*, D<92>*, wire7396*, key<237>*, wire8273*, D<91>*, wire7379*, key<245>*, wire8278*, D<90>*, wire8280*, key<253>*, wire8284*, D<89>*, wire7383*, key<198>*, wire8289*, D<88>*, wire7389*, key<206>*, wire8294*, D<87>*, wire7377*, key<214>*, wire8299*, D<86>*, wire7397*, key<222>*, wire8304*, D<85>*, wire7393*, key<230>*, wire8309*, D<84>*, wire7378*, key<238>*, wire8314*, D<83>*, wire7407*, key<246>*, wire8319*, D<82>*, wire7417*, key<254>*, wire8324*, D<81>*, wire8326*, key<131>*, wire8330*, D<80>*, wire7405*, key<139>*, wire8335*, D<79>*, wire7421*, key<147>*, wire8340*, D<78>*, wire7414*, key<155>*, wire8345*, D<77>*, wire7402*, key<132>*, wire8350*, D<76>*, wire7409*, key<140>*, wire8355*, D<75>*, wire7411*, key<148>*, wire8360*, D<74>*, wire7418*, key<156>*, wire8365*, D<73>*, wire7404*, key<164>*, wire8370*, D<72>*, wire8372*, D<71>*, wire7410*, key<180>*, wire8380*, D<70>*, wire7413*, key<188>*, wire8385*, D<69>*, wire7403*, key<133>*, wire8390*, D<68>*, wire7422*, key<141>*, wire8395*, D<67>*, wire7415*, key<149>*, wire8400*, D<66>*, wire7408*, key<157>*, wire8405*, D<65>*, wire8407*, key<165>*, wire8411*, D<64>*, wire7419*, key<173>*, wire8416*, D<63>*, wire7401*, key<181>*, wire8421*, D<62>*, wire8423*, key<189>*, wire8427*, D<61>*, wire7406*, key<134>*, wire8432*, D<60>*, wire7412*, key<142>*, wire8437*, D<59>*, wire7399*, key<150>*, wire8442*, D<58>*, wire7420*, key<158>*, wire8447*, D<57>*, wire7416*, key<166>*, wire8452*, D<56>*, wire7400*, key<174>*, wire8457*, D<55>*, wire7430*, key<182>*, wire8462*, D<54>*, wire7440*, key<190>*, wire8467*, D<53>*, wire8469*, key<67>*, wire8473*, D<52>*, wire7428*, key<75>*, wire8478*, D<51>*, wire7444*, key<83>*, wire8483*, D<50>*, wire7437*, key<91>*, wire8488*, D<49>*, wire7426*, key<68>*, wire8493*, D<48>*, wire7432*, key<76>*, wire8498*, D<47>*, wire7434*, key<84>*, wire8503*, D<46>*, wire7441*, key<92>*, wire8508*, D<45>*, wire7427*, key<100>*, wire8513*, D<44>*, wire7436*, key<44>*, wire8518*, D<43>*, wire7433*, key<116>*, wire8523*, D<42>*, wire8525*, key<124>*, wire8529*, D<41>*, wire8531*, key<69>*, wire8535*, D<40>*, wire7445*, key<77>*, wire8540*, D<39>*, wire7438*, key<85>*, wire8545*, D<38>*, wire7431*, key<93>*, wire8550*, D<37>*, wire8552*, key<101>*, wire8556*, D<36>*, wire7442*, key<109>*, wire8561*, D<35>*, wire7425*, key<117>*, wire8566*, D<34>*, wire8568*, key<125>*, wire8572*, D<33>*, wire7429*, key<70>*, wire8577*, D<32>*, wire7435*, key<78>*, wire8582*, D<31>*, wire7423*, key<86>*, wire8587*, D<30>*, wire7443*, key<94>*, wire8592*, D<29>*, wire7439*, key<102>*, wire8597*, D<28>*, wire7424*, key<110>*, wire8602*, D<27>*, wire7454*, key<118>*, wire8607*, D<26>*, wire7464*, key<126>*, wire8612*, D<25>*, wire8614*, key<3>*, wire8618*, D<24>*, wire7452*, key<11>*, wire8623*, D<23>*, wire7468*, key<19>*, wire8628*, D<22>*, wire7461*, key<27>*, wire8633*, D<21>*, wire7449*, key<4>*, wire8638*, D<20>*, wire7456*, key<12>*, wire8643*, D<19>*, wire7458*, key<20>*, wire8648*, D<18>*, wire7465*, key<28>*, wire8653*, D<17>*, wire7451*, key<36>*, wire8658*, D<16>*, wire7460*, D<15>*, wire7457*, key<52>*, wire8667*, D<14>*, wire8669*, key<60>*, wire8673*, D<13>*, wire7450*, key<5>*, wire8678*, D<12>*, wire7469*, key<13>*, wire8683*, D<11>*, wire7462*, key<21>*, wire8688*, D<10>*, wire7455*, key<29>*, wire8693*, D<9>*, wire8695*, key<37>*, wire8699*, D<8>*, wire7466*, key<45>*, wire8704*, D<7>*, wire7448*, key<53>*, wire8709*, D<6>*, wire8711*, key<61>*, wire8715*, D<5>*, wire7453*, key<6>*, wire8720*, D<4>*, wire7459*, key<14>*, wire8725*, D<3>*, wire7446*, key<22>*, wire8730*, D<2>*, wire7467*, key<30>*, wire8735*, key<38>*, wire8740*, key<46>*, wire8745*, key<54>*, wire8750*, wire7570*, wire7596*, wire8756*, wire8757*;

reg C<111>, C<110>, C<109>, C<108>, C<107>, C<106>, C<105>, C<104>, C<103>, C<102>, C<101>, C<100>, C<99>, C<98>, C<97>, C<96>, C<95>, C<94>, C<93>, C<92>, C<91>, C<90>, C<89>, C<88>, C<87>, C<86>, C<85>, C<84>, C<83>, C<82>, C<81>, C<80>, C<79>, C<78>, C<77>, C<76>, C<75>, C<74>, C<73>, C<72>, C<71>, C<70>, C<69>, C<68>, C<67>, C<66>, C<65>, C<64>, C<63>, C<62>, C<61>, C<60>, C<59>, C<58>, C<57>, C<56>, C<55>, C<54>, C<53>, C<52>, C<51>, C<50>, C<49>, C<48>, C<47>, C<46>, C<45>, C<44>, C<43>, C<42>, C<41>, C<40>, C<39>, C<38>, C<37>, C<36>, C<35>, C<34>, C<33>, C<32>, C<31>, C<30>, C<29>, C<28>, C<27>, C<26>, C<25>, C<24>, C<23>, C<22>, C<21>, C<20>, C<19>, C<18>, C<17>, C<16>, C<15>, C<14>, C<13>, C<12>, C<11>, C<10>, C<9>, C<8>, C<7>, C<6>, C<5>, C<4>, C<3>, C<2>, C<1>, C<0>, D<111>, D<110>, D<109>, D<108>, D<107>, D<106>, D<105>, D<104>, D<103>, D<102>, D<101>, D<100>, D<99>, D<98>, D<97>, D<96>, D<95>, D<94>, D<93>, D<92>, D<91>, D<90>, D<89>, D<88>, D<87>, D<86>, D<85>, D<84>, D<83>, D<82>, D<81>, D<80>, D<79>, D<78>, D<77>, D<76>, D<75>, D<74>, D<73>, D<72>, D<71>, D<70>, D<69>, D<68>, D<67>, D<66>, D<65>, D<64>, D<63>, D<62>, D<61>, D<60>, D<59>, D<58>, D<57>, D<56>, D<55>, D<54>, D<53>, D<52>, D<51>, D<50>, D<49>, D<48>, D<47>, D<46>, D<45>, D<44>, D<43>, D<42>, D<41>, D<40>, D<39>, D<38>, D<37>, D<36>, D<35>, D<34>, D<33>, D<32>, D<31>, D<30>, D<29>, D<28>, D<27>, D<26>, D<25>, D<24>, D<23>, D<22>, D<21>, D<20>, D<19>, D<18>, D<17>, D<16>, D<15>, D<14>, D<13>, D<12>, D<11>, D<10>, D<9>, D<8>, D<7>, D<6>, D<5>, D<4>, D<3>, D<2>, D<1>, D<0>;

initial
begin
	C<111> = 0;
	C<110> = 0;
	C<109> = 0;
	C<108> = 0;
	C<107> = 0;
	C<106> = 0;
	C<105> = 0;
	C<104> = 0;
	C<103> = 0;
	C<102> = 0;
	C<101> = 0;
	C<100> = 0;
	C<99> = 0;
	C<98> = 0;
	C<97> = 0;
	C<96> = 0;
	C<95> = 0;
	C<94> = 0;
	C<93> = 0;
	C<92> = 0;
	C<91> = 0;
	C<90> = 0;
	C<89> = 0;
	C<88> = 0;
	C<87> = 0;
	C<86> = 0;
	C<85> = 0;
	C<84> = 0;
	C<83> = 0;
	C<82> = 0;
	C<81> = 0;
	C<80> = 0;
	C<79> = 0;
	C<78> = 0;
	C<77> = 0;
	C<76> = 0;
	C<75> = 0;
	C<74> = 0;
	C<73> = 0;
	C<72> = 0;
	C<71> = 0;
	C<70> = 0;
	C<69> = 0;
	C<68> = 0;
	C<67> = 0;
	C<66> = 0;
	C<65> = 0;
	C<64> = 0;
	C<63> = 0;
	C<62> = 0;
	C<61> = 0;
	C<60> = 0;
	C<59> = 0;
	C<58> = 0;
	C<57> = 0;
	C<56> = 0;
	C<55> = 0;
	C<54> = 0;
	C<53> = 0;
	C<52> = 0;
	C<51> = 0;
	C<50> = 0;
	C<49> = 0;
	C<48> = 0;
	C<47> = 0;
	C<46> = 0;
	C<45> = 0;
	C<44> = 0;
	C<43> = 0;
	C<42> = 0;
	C<41> = 0;
	C<40> = 0;
	C<39> = 0;
	C<38> = 0;
	C<37> = 0;
	C<36> = 0;
	C<35> = 0;
	C<34> = 0;
	C<33> = 0;
	C<32> = 0;
	C<31> = 0;
	C<30> = 0;
	C<29> = 0;
	C<28> = 0;
	C<27> = 0;
	C<26> = 0;
	C<25> = 0;
	C<24> = 0;
	C<23> = 0;
	C<22> = 0;
	C<21> = 0;
	C<20> = 0;
	C<19> = 0;
	C<18> = 0;
	C<17> = 0;
	C<16> = 0;
	C<15> = 0;
	C<14> = 0;
	C<13> = 0;
	C<12> = 0;
	C<11> = 0;
	C<10> = 0;
	C<9> = 0;
	C<8> = 0;
	C<7> = 0;
	C<6> = 0;
	C<5> = 0;
	C<4> = 0;
	C<3> = 0;
	C<2> = 0;
	C<1> = 0;
	C<0> = 0;
	D<111> = 0;
	D<110> = 0;
	D<109> = 0;
	D<108> = 0;
	D<107> = 0;
	D<106> = 0;
	D<105> = 0;
	D<104> = 0;
	D<103> = 0;
	D<102> = 0;
	D<101> = 0;
	D<100> = 0;
	D<99> = 0;
	D<98> = 0;
	D<97> = 0;
	D<96> = 0;
	D<95> = 0;
	D<94> = 0;
	D<93> = 0;
	D<92> = 0;
	D<91> = 0;
	D<90> = 0;
	D<89> = 0;
	D<88> = 0;
	D<87> = 0;
	D<86> = 0;
	D<85> = 0;
	D<84> = 0;
	D<83> = 0;
	D<82> = 0;
	D<81> = 0;
	D<80> = 0;
	D<79> = 0;
	D<78> = 0;
	D<77> = 0;
	D<76> = 0;
	D<75> = 0;
	D<74> = 0;
	D<73> = 0;
	D<72> = 0;
	D<71> = 0;
	D<70> = 0;
	D<69> = 0;
	D<68> = 0;
	D<67> = 0;
	D<66> = 0;
	D<65> = 0;
	D<64> = 0;
	D<63> = 0;
	D<62> = 0;
	D<61> = 0;
	D<60> = 0;
	D<59> = 0;
	D<58> = 0;
	D<57> = 0;
	D<56> = 0;
	D<55> = 0;
	D<54> = 0;
	D<53> = 0;
	D<52> = 0;
	D<51> = 0;
	D<50> = 0;
	D<49> = 0;
	D<48> = 0;
	D<47> = 0;
	D<46> = 0;
	D<45> = 0;
	D<44> = 0;
	D<43> = 0;
	D<42> = 0;
	D<41> = 0;
	D<40> = 0;
	D<39> = 0;
	D<38> = 0;
	D<37> = 0;
	D<36> = 0;
	D<35> = 0;
	D<34> = 0;
	D<33> = 0;
	D<32> = 0;
	D<31> = 0;
	D<30> = 0;
	D<29> = 0;
	D<28> = 0;
	D<27> = 0;
	D<26> = 0;
	D<25> = 0;
	D<24> = 0;
	D<23> = 0;
	D<22> = 0;
	D<21> = 0;
	D<20> = 0;
	D<19> = 0;
	D<18> = 0;
	D<17> = 0;
	D<16> = 0;
	D<15> = 0;
	D<14> = 0;
	D<13> = 0;
	D<12> = 0;
	D<11> = 0;
	D<10> = 0;
	D<9> = 0;
	D<8> = 0;
	D<7> = 0;
	D<6> = 0;
	D<5> = 0;
	D<4> = 0;
	D<3> = 0;
	D<2> = 0;
	D<1> = 0;
	D<0> = 0;
end

always @(new_C<111>)
	C<111><=new_C<111>;

 always @(new_C<110>)
	C<110><=new_C<110>;

 always @(new_C<109>)
	C<109><=new_C<109>;

 always @(new_C<108>)
	C<108><=new_C<108>;

 always @(new_C<107>)
	C<107><=new_C<107>;

 always @(new_C<106>)
	C<106><=new_C<106>;

 always @(new_C<105>)
	C<105><=new_C<105>;

 always @(new_C<104>)
	C<104><=new_C<104>;

 always @(new_C<103>)
	C<103><=new_C<103>;

 always @(new_C<102>)
	C<102><=new_C<102>;

 always @(new_C<101>)
	C<101><=new_C<101>;

 always @(new_C<100>)
	C<100><=new_C<100>;

 always @(new_C<99>)
	C<99><=new_C<99>;

 always @(new_C<98>)
	C<98><=new_C<98>;

 always @(new_C<97>)
	C<97><=new_C<97>;

 always @(new_C<96>)
	C<96><=new_C<96>;

 always @(new_C<95>)
	C<95><=new_C<95>;

 always @(new_C<94>)
	C<94><=new_C<94>;

 always @(new_C<93>)
	C<93><=new_C<93>;

 always @(new_C<92>)
	C<92><=new_C<92>;

 always @(new_C<91>)
	C<91><=new_C<91>;

 always @(new_C<90>)
	C<90><=new_C<90>;

 always @(new_C<89>)
	C<89><=new_C<89>;

 always @(new_C<88>)
	C<88><=new_C<88>;

 always @(new_C<87>)
	C<87><=new_C<87>;

 always @(new_C<86>)
	C<86><=new_C<86>;

 always @(new_C<85>)
	C<85><=new_C<85>;

 always @(new_C<84>)
	C<84><=new_C<84>;

 always @(new_C<83>)
	C<83><=new_C<83>;

 always @(new_C<82>)
	C<82><=new_C<82>;

 always @(new_C<81>)
	C<81><=new_C<81>;

 always @(new_C<80>)
	C<80><=new_C<80>;

 always @(new_C<79>)
	C<79><=new_C<79>;

 always @(new_C<78>)
	C<78><=new_C<78>;

 always @(new_C<77>)
	C<77><=new_C<77>;

 always @(new_C<76>)
	C<76><=new_C<76>;

 always @(new_C<75>)
	C<75><=new_C<75>;

 always @(new_C<74>)
	C<74><=new_C<74>;

 always @(new_C<73>)
	C<73><=new_C<73>;

 always @(new_C<72>)
	C<72><=new_C<72>;

 always @(new_C<71>)
	C<71><=new_C<71>;

 always @(new_C<70>)
	C<70><=new_C<70>;

 always @(new_C<69>)
	C<69><=new_C<69>;

 always @(new_C<68>)
	C<68><=new_C<68>;

 always @(new_C<67>)
	C<67><=new_C<67>;

 always @(new_C<66>)
	C<66><=new_C<66>;

 always @(new_C<65>)
	C<65><=new_C<65>;

 always @(new_C<64>)
	C<64><=new_C<64>;

 always @(new_C<63>)
	C<63><=new_C<63>;

 always @(new_C<62>)
	C<62><=new_C<62>;

 always @(new_C<61>)
	C<61><=new_C<61>;

 always @(new_C<60>)
	C<60><=new_C<60>;

 always @(new_C<59>)
	C<59><=new_C<59>;

 always @(new_C<58>)
	C<58><=new_C<58>;

 always @(new_C<57>)
	C<57><=new_C<57>;

 always @(new_C<56>)
	C<56><=new_C<56>;

 always @(new_C<55>)
	C<55><=new_C<55>;

 always @(new_C<54>)
	C<54><=new_C<54>;

 always @(new_C<53>)
	C<53><=new_C<53>;

 always @(new_C<52>)
	C<52><=new_C<52>;

 always @(new_C<51>)
	C<51><=new_C<51>;

 always @(new_C<50>)
	C<50><=new_C<50>;

 always @(new_C<49>)
	C<49><=new_C<49>;

 always @(new_C<48>)
	C<48><=new_C<48>;

 always @(new_C<47>)
	C<47><=new_C<47>;

 always @(new_C<46>)
	C<46><=new_C<46>;

 always @(new_C<45>)
	C<45><=new_C<45>;

 always @(new_C<44>)
	C<44><=new_C<44>;

 always @(new_C<43>)
	C<43><=new_C<43>;

 always @(new_C<42>)
	C<42><=new_C<42>;

 always @(new_C<41>)
	C<41><=new_C<41>;

 always @(new_C<40>)
	C<40><=new_C<40>;

 always @(new_C<39>)
	C<39><=new_C<39>;

 always @(new_C<38>)
	C<38><=new_C<38>;

 always @(new_C<37>)
	C<37><=new_C<37>;

 always @(new_C<36>)
	C<36><=new_C<36>;

 always @(new_C<35>)
	C<35><=new_C<35>;

 always @(new_C<34>)
	C<34><=new_C<34>;

 always @(new_C<33>)
	C<33><=new_C<33>;

 always @(new_C<32>)
	C<32><=new_C<32>;

 always @(new_C<31>)
	C<31><=new_C<31>;

 always @(new_C<30>)
	C<30><=new_C<30>;

 always @(new_C<29>)
	C<29><=new_C<29>;

 always @(new_C<28>)
	C<28><=new_C<28>;

 always @(new_C<27>)
	C<27><=new_C<27>;

 always @(new_C<26>)
	C<26><=new_C<26>;

 always @(new_C<25>)
	C<25><=new_C<25>;

 always @(new_C<24>)
	C<24><=new_C<24>;

 always @(new_C<23>)
	C<23><=new_C<23>;

 always @(new_C<22>)
	C<22><=new_C<22>;

 always @(new_C<21>)
	C<21><=new_C<21>;

 always @(new_C<20>)
	C<20><=new_C<20>;

 always @(new_C<19>)
	C<19><=new_C<19>;

 always @(new_C<18>)
	C<18><=new_C<18>;

 always @(new_C<17>)
	C<17><=new_C<17>;

 always @(new_C<16>)
	C<16><=new_C<16>;

 always @(new_C<15>)
	C<15><=new_C<15>;

 always @(new_C<14>)
	C<14><=new_C<14>;

 always @(new_C<13>)
	C<13><=new_C<13>;

 always @(new_C<12>)
	C<12><=new_C<12>;

 always @(new_C<11>)
	C<11><=new_C<11>;

 always @(new_C<10>)
	C<10><=new_C<10>;

 always @(new_C<9>)
	C<9><=new_C<9>;

 always @(new_C<8>)
	C<8><=new_C<8>;

 always @(new_C<7>)
	C<7><=new_C<7>;

 always @(new_C<6>)
	C<6><=new_C<6>;

 always @(new_C<5>)
	C<5><=new_C<5>;

 always @(new_C<4>)
	C<4><=new_C<4>;

 always @(new_C<3>)
	C<3><=new_C<3>;

 always @(new_C<2>)
	C<2><=new_C<2>;

 always @(new_C<1>)
	C<1><=new_C<1>;

 always @(new_C<0>)
	C<0><=new_C<0>;

 always @(new_D<111>)
	D<111><=new_D<111>;

 always @(new_D<110>)
	D<110><=new_D<110>;

 always @(new_D<109>)
	D<109><=new_D<109>;

 always @(new_D<108>)
	D<108><=new_D<108>;

 always @(new_D<107>)
	D<107><=new_D<107>;

 always @(new_D<106>)
	D<106><=new_D<106>;

 always @(new_D<105>)
	D<105><=new_D<105>;

 always @(new_D<104>)
	D<104><=new_D<104>;

 always @(new_D<103>)
	D<103><=new_D<103>;

 always @(new_D<102>)
	D<102><=new_D<102>;

 always @(new_D<101>)
	D<101><=new_D<101>;

 always @(new_D<100>)
	D<100><=new_D<100>;

 always @(new_D<99>)
	D<99><=new_D<99>;

 always @(new_D<98>)
	D<98><=new_D<98>;

 always @(new_D<97>)
	D<97><=new_D<97>;

 always @(new_D<96>)
	D<96><=new_D<96>;

 always @(new_D<95>)
	D<95><=new_D<95>;

 always @(new_D<94>)
	D<94><=new_D<94>;

 always @(new_D<93>)
	D<93><=new_D<93>;

 always @(new_D<92>)
	D<92><=new_D<92>;

 always @(new_D<91>)
	D<91><=new_D<91>;

 always @(new_D<90>)
	D<90><=new_D<90>;

 always @(new_D<89>)
	D<89><=new_D<89>;

 always @(new_D<88>)
	D<88><=new_D<88>;

 always @(new_D<87>)
	D<87><=new_D<87>;

 always @(new_D<86>)
	D<86><=new_D<86>;

 always @(new_D<85>)
	D<85><=new_D<85>;

 always @(new_D<84>)
	D<84><=new_D<84>;

 always @(new_D<83>)
	D<83><=new_D<83>;

 always @(new_D<82>)
	D<82><=new_D<82>;

 always @(new_D<81>)
	D<81><=new_D<81>;

 always @(new_D<80>)
	D<80><=new_D<80>;

 always @(new_D<79>)
	D<79><=new_D<79>;

 always @(new_D<78>)
	D<78><=new_D<78>;

 always @(new_D<77>)
	D<77><=new_D<77>;

 always @(new_D<76>)
	D<76><=new_D<76>;

 always @(new_D<75>)
	D<75><=new_D<75>;

 always @(new_D<74>)
	D<74><=new_D<74>;

 always @(new_D<73>)
	D<73><=new_D<73>;

 always @(new_D<72>)
	D<72><=new_D<72>;

 always @(new_D<71>)
	D<71><=new_D<71>;

 always @(new_D<70>)
	D<70><=new_D<70>;

 always @(new_D<69>)
	D<69><=new_D<69>;

 always @(new_D<68>)
	D<68><=new_D<68>;

 always @(new_D<67>)
	D<67><=new_D<67>;

 always @(new_D<66>)
	D<66><=new_D<66>;

 always @(new_D<65>)
	D<65><=new_D<65>;

 always @(new_D<64>)
	D<64><=new_D<64>;

 always @(new_D<63>)
	D<63><=new_D<63>;

 always @(new_D<62>)
	D<62><=new_D<62>;

 always @(new_D<61>)
	D<61><=new_D<61>;

 always @(new_D<60>)
	D<60><=new_D<60>;

 always @(new_D<59>)
	D<59><=new_D<59>;

 always @(new_D<58>)
	D<58><=new_D<58>;

 always @(new_D<57>)
	D<57><=new_D<57>;

 always @(new_D<56>)
	D<56><=new_D<56>;

 always @(new_D<55>)
	D<55><=new_D<55>;

 always @(new_D<54>)
	D<54><=new_D<54>;

 always @(new_D<53>)
	D<53><=new_D<53>;

 always @(new_D<52>)
	D<52><=new_D<52>;

 always @(new_D<51>)
	D<51><=new_D<51>;

 always @(new_D<50>)
	D<50><=new_D<50>;

 always @(new_D<49>)
	D<49><=new_D<49>;

 always @(new_D<48>)
	D<48><=new_D<48>;

 always @(new_D<47>)
	D<47><=new_D<47>;

 always @(new_D<46>)
	D<46><=new_D<46>;

 always @(new_D<45>)
	D<45><=new_D<45>;

 always @(new_D<44>)
	D<44><=new_D<44>;

 always @(new_D<43>)
	D<43><=new_D<43>;

 always @(new_D<42>)
	D<42><=new_D<42>;

 always @(new_D<41>)
	D<41><=new_D<41>;

 always @(new_D<40>)
	D<40><=new_D<40>;

 always @(new_D<39>)
	D<39><=new_D<39>;

 always @(new_D<38>)
	D<38><=new_D<38>;

 always @(new_D<37>)
	D<37><=new_D<37>;

 always @(new_D<36>)
	D<36><=new_D<36>;

 always @(new_D<35>)
	D<35><=new_D<35>;

 always @(new_D<34>)
	D<34><=new_D<34>;

 always @(new_D<33>)
	D<33><=new_D<33>;

 always @(new_D<32>)
	D<32><=new_D<32>;

 always @(new_D<31>)
	D<31><=new_D<31>;

 always @(new_D<30>)
	D<30><=new_D<30>;

 always @(new_D<29>)
	D<29><=new_D<29>;

 always @(new_D<28>)
	D<28><=new_D<28>;

 always @(new_D<27>)
	D<27><=new_D<27>;

 always @(new_D<26>)
	D<26><=new_D<26>;

 always @(new_D<25>)
	D<25><=new_D<25>;

 always @(new_D<24>)
	D<24><=new_D<24>;

 always @(new_D<23>)
	D<23><=new_D<23>;

 always @(new_D<22>)
	D<22><=new_D<22>;

 always @(new_D<21>)
	D<21><=new_D<21>;

 always @(new_D<20>)
	D<20><=new_D<20>;

 always @(new_D<19>)
	D<19><=new_D<19>;

 always @(new_D<18>)
	D<18><=new_D<18>;

 always @(new_D<17>)
	D<17><=new_D<17>;

 always @(new_D<16>)
	D<16><=new_D<16>;

 always @(new_D<15>)
	D<15><=new_D<15>;

 always @(new_D<14>)
	D<14><=new_D<14>;

 always @(new_D<13>)
	D<13><=new_D<13>;

 always @(new_D<12>)
	D<12><=new_D<12>;

 always @(new_D<11>)
	D<11><=new_D<11>;

 always @(new_D<10>)
	D<10><=new_D<10>;

 always @(new_D<9>)
	D<9><=new_D<9>;

 always @(new_D<8>)
	D<8><=new_D<8>;

 always @(new_D<7>)
	D<7><=new_D<7>;

 always @(new_D<6>)
	D<6><=new_D<6>;

 always @(new_D<5>)
	D<5><=new_D<5>;

 always @(new_D<4>)
	D<4><=new_D<4>;

 always @(new_D<3>)
	D<3><=new_D<3>;

 always @(new_D<2>)
	D<2><=new_D<2>;

 always @(new_D<1>)
	D<1><=new_D<1>;

 always @(new_D<0>)
	D<0><=new_D<0>;

 assign KSi<191> = ( D<87> ) ;
 assign KSi<190> = ( D<84> ) ;
 assign KSi<189> = ( D<91> ) ;
 assign KSi<188> = ( D<105> ) ;
 assign KSi<187> = ( D<87> ) ;
 assign KSi<186> = ( D<101> ) ;
 assign KSi<185> = ( D<108> ) ;
 assign KSi<184> = ( D<89> ) ;
 assign KSi<183> = ( D<111> ) ;
 assign KSi<182> = ( D<94> ) ;
 assign KSi<181> = ( D<104> ) ;
 assign KSi<180> = ( D<99> ) ;
 assign KSi<179> = ( D<103> ) ;
 assign KSi<178> = ( D<88> ) ;
 assign KSi<177> = ( D<100> ) ;
 assign KSi<176> = ( D<106> ) ;
 assign KSi<175> = ( D<95> ) ;
 assign KSi<174> = ( D<85> ) ;
 assign KSi<173> = ( D<110> ) ;
 assign KSi<172> = ( D<102> ) ;
 assign KSi<171> = ( D<92> ) ;
 assign KSi<170> = ( D<86> ) ;
 assign KSi<169> = ( D<107> ) ;
 assign KSi<168> = ( D<104> ) ;
 assign KSi<167> = ( D<59> ) ;
 assign KSi<166> = ( D<56> ) ;
 assign KSi<165> = ( D<63> ) ;
 assign KSi<164> = ( D<77> ) ;
 assign KSi<163> = ( D<69> ) ;
 assign KSi<162> = ( D<73> ) ;
 assign KSi<161> = ( D<80> ) ;
 assign KSi<160> = ( D<61> ) ;
 assign KSi<159> = ( D<83> ) ;
 assign KSi<158> = ( D<66> ) ;
 assign KSi<157> = ( D<76> ) ;
 assign KSi<156> = ( D<71> ) ;
 assign KSi<155> = ( D<75> ) ;
 assign KSi<154> = ( D<60> ) ;
 assign KSi<153> = ( D<70> ) ;
 assign KSi<152> = ( D<78> ) ;
 assign KSi<151> = ( D<67> ) ;
 assign KSi<150> = ( D<57> ) ;
 assign KSi<149> = ( D<82> ) ;
 assign KSi<148> = ( D<74> ) ;
 assign KSi<147> = ( D<64> ) ;
 assign KSi<146> = ( D<58> ) ;
 assign KSi<145> = ( D<79> ) ;
 assign KSi<144> = ( D<68> ) ;
 assign KSi<143> = ( D<31> ) ;
 assign KSi<142> = ( D<28> ) ;
 assign KSi<141> = ( D<35> ) ;
 assign KSi<140> = ( D<49> ) ;
 assign KSi<139> = ( D<31> ) ;
 assign KSi<138> = ( D<45> ) ;
 assign KSi<137> = ( D<52> ) ;
 assign KSi<136> = ( D<33> ) ;
 assign KSi<135> = ( D<55> ) ;
 assign KSi<134> = ( D<38> ) ;
 assign KSi<133> = ( D<48> ) ;
 assign KSi<132> = ( D<43> ) ;
 assign KSi<131> = ( D<47> ) ;
 assign KSi<130> = ( D<32> ) ;
 assign KSi<129> = ( D<44> ) ;
 assign KSi<128> = ( D<50> ) ;
 assign KSi<127> = ( D<39> ) ;
 assign KSi<126> = ( D<29> ) ;
 assign KSi<125> = ( D<54> ) ;
 assign KSi<124> = ( D<46> ) ;
 assign KSi<123> = ( D<36> ) ;
 assign KSi<122> = ( D<30> ) ;
 assign KSi<121> = ( D<51> ) ;
 assign KSi<120> = ( D<40> ) ;
 assign KSi<119> = ( D<3> ) ;
 assign KSi<118> = ( D<0> ) ;
 assign KSi<117> = ( D<7> ) ;
 assign KSi<116> = ( D<21> ) ;
 assign KSi<115> = ( D<13> ) ;
 assign KSi<114> = ( D<17> ) ;
 assign KSi<113> = ( D<24> ) ;
 assign KSi<112> = ( D<5> ) ;
 assign KSi<111> = ( D<27> ) ;
 assign KSi<110> = ( D<10> ) ;
 assign KSi<109> = ( D<20> ) ;
 assign KSi<108> = ( D<15> ) ;
 assign KSi<107> = ( D<19> ) ;
 assign KSi<106> = ( D<4> ) ;
 assign KSi<105> = ( D<16> ) ;
 assign KSi<104> = ( D<22> ) ;
 assign KSi<103> = ( D<11> ) ;
 assign KSi<102> = ( D<1> ) ;
 assign KSi<101> = ( D<26> ) ;
 assign KSi<100> = ( D<18> ) ;
 assign KSi<99> = ( D<8> ) ;
 assign KSi<98> = ( D<2> ) ;
 assign KSi<97> = ( D<23> ) ;
 assign KSi<96> = ( D<12> ) ;
 assign KSi<95> = ( C<85> ) ;
 assign KSi<94> = ( C<96> ) ;
 assign KSi<93> = ( C<103> ) ;
 assign KSi<92> = ( C<110> ) ;
 assign KSi<91> = ( C<90> ) ;
 assign KSi<90> = ( C<109> ) ;
 assign KSi<89> = ( C<91> ) ;
 assign KSi<88> = ( C<109> ) ;
 assign KSi<87> = ( C<87> ) ;
 assign KSi<86> = ( C<95> ) ;
 assign KSi<85> = ( C<102> ) ;
 assign KSi<84> = ( C<106> ) ;
 assign KSi<83> = ( C<93> ) ;
 assign KSi<82> = ( C<104> ) ;
 assign KSi<81> = ( C<89> ) ;
 assign KSi<80> = ( C<98> ) ;
 assign KSi<79> = ( C<111> ) ;
 assign KSi<78> = ( C<86> ) ;
 assign KSi<77> = ( C<88> ) ;
 assign KSi<76> = ( C<84> ) ;
 assign KSi<75> = ( C<107> ) ;
 assign KSi<74> = ( C<94> ) ;
 assign KSi<73> = ( C<100> ) ;
 assign KSi<72> = ( C<97> ) ;
 assign KSi<71> = ( C<57> ) ;
 assign KSi<70> = ( C<68> ) ;
 assign KSi<69> = ( C<75> ) ;
 assign KSi<68> = ( C<82> ) ;
 assign KSi<67> = ( C<62> ) ;
 assign KSi<66> = ( C<71> ) ;
 assign KSi<65> = ( C<63> ) ;
 assign KSi<64> = ( C<81> ) ;
 assign KSi<63> = ( C<59> ) ;
 assign KSi<62> = ( C<67> ) ;
 assign KSi<61> = ( C<74> ) ;
 assign KSi<60> = ( C<78> ) ;
 assign KSi<59> = ( C<65> ) ;
 assign KSi<58> = ( C<76> ) ;
 assign KSi<57> = ( C<61> ) ;
 assign KSi<56> = ( C<70> ) ;
 assign KSi<55> = ( C<83> ) ;
 assign KSi<54> = ( C<58> ) ;
 assign KSi<53> = ( C<60> ) ;
 assign KSi<52> = ( C<56> ) ;
 assign KSi<51> = ( C<79> ) ;
 assign KSi<50> = ( C<66> ) ;
 assign KSi<49> = ( C<72> ) ;
 assign KSi<48> = ( C<69> ) ;
 assign KSi<47> = ( C<29> ) ;
 assign KSi<46> = ( C<40> ) ;
 assign KSi<45> = ( C<47> ) ;
 assign KSi<44> = ( C<54> ) ;
 assign KSi<43> = ( C<34> ) ;
 assign KSi<42> = ( C<43> ) ;
 assign KSi<41> = ( C<35> ) ;
 assign KSi<40> = ( C<53> ) ;
 assign KSi<39> = ( C<31> ) ;
 assign KSi<38> = ( C<39> ) ;
 assign KSi<37> = ( C<46> ) ;
 assign KSi<36> = ( C<50> ) ;
 assign KSi<35> = ( C<37> ) ;
 assign KSi<34> = ( C<48> ) ;
 assign KSi<33> = ( C<33> ) ;
 assign KSi<32> = ( C<42> ) ;
 assign KSi<31> = ( C<55> ) ;
 assign KSi<30> = ( C<30> ) ;
 assign KSi<29> = ( C<32> ) ;
 assign KSi<28> = ( C<28> ) ;
 assign KSi<27> = ( C<51> ) ;
 assign KSi<26> = ( C<38> ) ;
 assign KSi<25> = ( C<44> ) ;
 assign KSi<24> = ( C<41> ) ;
 assign KSi<23> = ( C<1> ) ;
 assign KSi<22> = ( C<12> ) ;
 assign KSi<21> = ( C<19> ) ;
 assign KSi<20> = ( C<26> ) ;
 assign KSi<19> = ( C<6> ) ;
 assign KSi<18> = ( C<15> ) ;
 assign KSi<17> = ( C<7> ) ;
 assign KSi<16> = ( C<25> ) ;
 assign KSi<15> = ( C<3> ) ;
 assign KSi<14> = ( C<11> ) ;
 assign KSi<13> = ( C<18> ) ;
 assign KSi<12> = ( C<22> ) ;
 assign KSi<11> = ( C<9> ) ;
 assign KSi<10> = ( C<20> ) ;
 assign KSi<9> = ( C<5> ) ;
 assign KSi<8> = ( C<14> ) ;
 assign KSi<7> = ( C<27> ) ;
 assign KSi<6> = ( C<2> ) ;
 assign KSi<5> = ( C<4> ) ;
 assign KSi<4> = ( C<0> ) ;
 assign KSi<3> = ( C<23> ) ;
 assign KSi<2> = ( C<10> ) ;
 assign KSi<1> = ( C<16> ) ;
 assign KSi<0> = ( C<13> ) ;
 assign wire7572 = ( count<1> ) | ( count<0> ) | ( count<2> ) ;
 assign wire17163 = ( encrypt<0> ) | ( count<3> ) | ( wire7572 ) ;
 assign wire7573 = ( start<0>* ) ;
 assign wire7574 = ( encrypt<0>* ) | ( wire7573* ) ;
 assign wire7568 = ( count<2>* ) ;
 assign wire7575 = ( I200 ) | ( I199 ) ;
 assign I199 = ( wire7574*  &  count<2>* ) ;
 assign I200 = ( wire7568*  &  encrypt<0>* ) ;
 assign wire7576 = ( count<1>* ) | ( count<0>* ) ;
 assign wire11699 = ( wire7576* ) ;
 assign main/$MINUS_4_1/c<0>8 =((~ key<254>) & key<254>);
 assign wire7577 = ( I206 ) | ( I205 ) ;
 assign I205 = ( wire7574*  &  wire11699* ) ;
 assign main/$MINUS_4_1/c<0>8 =((~ key<254>) & key<254>);
 assign wire17165 = ( I208 ) | ( count<3>* ) ;
 assign I208 = ( wire7577*  &  wire7575* ) ;
 assign wire7565 = ( count<3>* ) ;
 assign wire7580 = ( count<2>* ) | ( wire7565* ) | ( wire11699* ) ;
 assign wire17167 = ( wire7580 ) | ( wire7574 ) ;
 assign wire7566 = ( encrypt<0>* ) ;
 assign wire7581 = ( start<0>* ) | ( wire7566* ) ;
 assign new_count<3> = ( wire7581* ) | ( wire17167* ) | ( wire17165* ) | ( wire17163* ) ;
 assign wire17157 = ( wire11699* ) | ( wire7568* ) | ( encrypt<0>* ) | ( wire7573* ) ;
 assign wire17159 = ( wire7572 ) | ( encrypt<0> ) ;
 assign wire17161 = ( count<2>* ) | ( wire7577* ) ;
 assign new_count<2> = ( wire7581* ) | ( wire17161* ) | ( wire17159* ) | ( wire17157* ) ;
 assign wire7571 = ( count<1> ) | ( count<0> ) ;
 assign wire7586 = ( wire7571* ) | ( wire7576* ) ;
 assign wire14444 = ( wire7586* ) ;
 assign wire7587 = ( I224 ) | ( I223 ) ;
 assign I223 = ( wire7586*  &  wire7574* ) ;
 assign I224 = ( wire14444*  &  encrypt<0>* ) ;
 assign new_count<0> = ( I226 ) | ( wire7581* ) ;
 assign I226 = ( start<0>*  &  count<0>* ) ;
 assign wire194 = ( I229 ) | ( I228 ) ;
 assign I228 = ( new_count<0>*  &  wire7587* ) ;
 assign I229 = ( start<0>*  &  wire7587* ) ;
 assign new_count<1> = ( wire194* ) ;
 assign wire7541 = ( C<1>* ) ;
 assign wire7569 = ( count<0>* ) ;
 assign wire17145 = ( count<1>* ) | ( wire7569* ) | ( count<2>* ) | ( count<3>* ) ;
 assign wire17147 = ( wire7572 ) | ( count<3> ) ;
 assign wire7591 = ( wire17147* ) | ( wire17145* ) | ( wire7580* ) ;
 assign wire7600 = ( wire7591 ) | ( wire7574 ) ;
 assign wire2074 = ( wire7600*  &  wire7541* ) ;
 assign wire7475 = ( C<109>* ) ;
 assign wire2079 = ( count<2>*  &  count<3>*  &  count<1>* ) ;
 assign wire7292 = ( wire7591*  &  wire7568* ) ;
 assign wire7284 = ( I243 ) | ( I242 ) ;
 assign I242 = ( wire11699*  &  wire2079* ) ;
 assign I243 = ( wire7292*  &  wire2079* ) ;
 assign wire7595 = ( wire7284* ) | ( wire7572* ) ;
 assign wire7597 = ( start<0> ) | ( encrypt<0> ) | ( wire7595 ) ;
 assign wire7473 = ( C<110>* ) ;
 assign wire7598 = ( wire7573* ) | ( wire7566* ) | ( wire7595* ) ;
 assign wire7599 = ( I250 ) | ( I249 ) ;
 assign I249 = ( wire7597*  &  wire7475* ) ;
 assign I250 = ( wire7598*  &  wire7473* ) ;
 assign wire7606 = ( key<227>* ) ;
 assign wire2077 = ( wire7606*  &  wire7581* ) ;
 assign wire7560 = ( C<0>* ) ;
 assign wire7602 = ( encrypt<0>* ) | ( wire7573* ) | ( wire7591* ) ;
 assign wire7603 = ( key<56>* ) ;
 assign wire7604 = ( start<0>* ) | ( encrypt<0>* ) ;
 assign wire7605 = ( I259 ) | ( I258 ) ;
 assign I258 = ( wire7602*  &  wire7560* ) ;
 assign I259 = ( wire7604*  &  wire7603* ) ;
 assign new_C<111> = ( wire7605 ) | ( wire2077 ) | ( wire7599 ) | ( wire2074 ) ;
 assign wire2068 = ( wire7600*  &  wire7560* ) ;
 assign wire7608 = ( C<108>* ) ;
 assign wire7609 = ( I265 ) | ( I264 ) ;
 assign I264 = ( wire7608*  &  wire7597* ) ;
 assign I265 = ( wire7598*  &  wire7475* ) ;
 assign wire7612 = ( key<235>* ) ;
 assign wire2071 = ( wire7612*  &  wire7581* ) ;
 assign wire7485 = ( C<111>* ) ;
 assign wire7611 = ( I271 ) | ( I270 ) ;
 assign I270 = ( wire7602*  &  wire7485* ) ;
 assign I271 = ( wire7606*  &  wire7604* ) ;
 assign new_C<110> = ( wire7611 ) | ( wire2071 ) | ( wire7609 ) | ( wire2068 ) ;
 assign wire2062 = ( wire7600*  &  wire7485* ) ;
 assign wire7489 = ( C<107>* ) ;
 assign wire7614 = ( I277 ) | ( I276 ) ;
 assign I276 = ( wire7597*  &  wire7489* ) ;
 assign I277 = ( wire7608*  &  wire7598* ) ;
 assign wire7617 = ( key<243>* ) ;
 assign wire2065 = ( wire7617*  &  wire7581* ) ;
 assign wire7616 = ( I282 ) | ( I281 ) ;
 assign I281 = ( wire7602*  &  wire7473* ) ;
 assign I282 = ( wire7612*  &  wire7604* ) ;
 assign new_C<109> = ( wire7616 ) | ( wire2065 ) | ( wire7614 ) | ( wire2062 ) ;
 assign wire2056 = ( wire7600*  &  wire7473* ) ;
 assign wire7480 = ( C<106>* ) ;
 assign wire7619 = ( I288 ) | ( I287 ) ;
 assign I287 = ( wire7597*  &  wire7480* ) ;
 assign I288 = ( wire7598*  &  wire7489* ) ;
 assign wire7622 = ( key<251>* ) ;
 assign wire2059 = ( wire7622*  &  wire7581* ) ;
 assign wire7621 = ( I293 ) | ( I292 ) ;
 assign I292 = ( wire7602*  &  wire7475* ) ;
 assign I293 = ( wire7617*  &  wire7604* ) ;
 assign new_C<108> = ( wire7621 ) | ( wire2059 ) | ( wire7619 ) | ( wire2056 ) ;
 assign wire2050 = ( wire7600*  &  wire7475* ) ;
 assign wire7624 = ( C<105>* ) ;
 assign wire7625 = ( I299 ) | ( I298 ) ;
 assign I298 = ( wire7624*  &  wire7597* ) ;
 assign I299 = ( wire7598*  &  wire7480* ) ;
 assign wire7628 = ( key<194>* ) ;
 assign wire2053 = ( wire7628*  &  wire7581* ) ;
 assign wire7627 = ( I304 ) | ( I303 ) ;
 assign I303 = ( wire7608*  &  wire7602* ) ;
 assign I304 = ( wire7622*  &  wire7604* ) ;
 assign new_C<107> = ( wire7627 ) | ( wire2053 ) | ( wire7625 ) | ( wire2050 ) ;
 assign wire2044 = ( wire7608*  &  wire7600* ) ;
 assign wire7482 = ( C<104>* ) ;
 assign wire7630 = ( I310 ) | ( I309 ) ;
 assign I309 = ( wire7597*  &  wire7482* ) ;
 assign I310 = ( wire7624*  &  wire7598* ) ;
 assign wire7633 = ( key<202>* ) ;
 assign wire2047 = ( wire7633*  &  wire7581* ) ;
 assign wire7632 = ( I315 ) | ( I314 ) ;
 assign I314 = ( wire7602*  &  wire7489* ) ;
 assign I315 = ( wire7628*  &  wire7604* ) ;
 assign new_C<106> = ( wire7632 ) | ( wire2047 ) | ( wire7630 ) | ( wire2044 ) ;
 assign wire2038 = ( wire7600*  &  wire7489* ) ;
 assign wire7472 = ( C<103>* ) ;
 assign wire7635 = ( I321 ) | ( I320 ) ;
 assign I320 = ( wire7597*  &  wire7472* ) ;
 assign I321 = ( wire7598*  &  wire7482* ) ;
 assign wire7638 = ( key<210>* ) ;
 assign wire2041 = ( wire7638*  &  wire7581* ) ;
 assign wire7637 = ( I326 ) | ( I325 ) ;
 assign I325 = ( wire7602*  &  wire7480* ) ;
 assign I326 = ( wire7633*  &  wire7604* ) ;
 assign new_C<105> = ( wire7637 ) | ( wire2041 ) | ( wire7635 ) | ( wire2038 ) ;
 assign wire2032 = ( wire7600*  &  wire7480* ) ;
 assign wire7479 = ( C<102>* ) ;
 assign wire7640 = ( I332 ) | ( I331 ) ;
 assign I331 = ( wire7597*  &  wire7479* ) ;
 assign I332 = ( wire7598*  &  wire7472* ) ;
 assign wire7643 = ( key<218>* ) ;
 assign wire2035 = ( wire7643*  &  wire7581* ) ;
 assign wire7642 = ( I337 ) | ( I336 ) ;
 assign I336 = ( wire7624*  &  wire7602* ) ;
 assign I337 = ( wire7638*  &  wire7604* ) ;
 assign new_C<104> = ( wire7642 ) | ( wire2035 ) | ( wire7640 ) | ( wire2032 ) ;
 assign wire2026 = ( wire7624*  &  wire7600* ) ;
 assign wire7645 = ( C<101>* ) ;
 assign wire7646 = ( I343 ) | ( I342 ) ;
 assign I342 = ( wire7645*  &  wire7597* ) ;
 assign I343 = ( wire7598*  &  wire7479* ) ;
 assign wire7649 = ( key<226>* ) ;
 assign wire2029 = ( wire7649*  &  wire7581* ) ;
 assign wire7648 = ( I348 ) | ( I347 ) ;
 assign I347 = ( wire7602*  &  wire7482* ) ;
 assign I348 = ( wire7643*  &  wire7604* ) ;
 assign new_C<103> = ( wire7648 ) | ( wire2029 ) | ( wire7646 ) | ( wire2026 ) ;
 assign wire2020 = ( wire7600*  &  wire7482* ) ;
 assign wire7491 = ( C<100>* ) ;
 assign wire7651 = ( I354 ) | ( I353 ) ;
 assign I353 = ( wire7597*  &  wire7491* ) ;
 assign I354 = ( wire7645*  &  wire7598* ) ;
 assign wire7654 = ( key<234>* ) ;
 assign wire2023 = ( wire7654*  &  wire7581* ) ;
 assign wire7653 = ( I359 ) | ( I358 ) ;
 assign I358 = ( wire7602*  &  wire7472* ) ;
 assign I359 = ( wire7649*  &  wire7604* ) ;
 assign new_C<102> = ( wire7653 ) | ( wire2023 ) | ( wire7651 ) | ( wire2020 ) ;
 assign wire2014 = ( wire7600*  &  wire7472* ) ;
 assign wire7656 = ( C<99>* ) ;
 assign wire7657 = ( I365 ) | ( I364 ) ;
 assign I364 = ( wire7656*  &  wire7597* ) ;
 assign I365 = ( wire7598*  &  wire7491* ) ;
 assign wire7660 = ( key<242>* ) ;
 assign wire2017 = ( wire7660*  &  wire7581* ) ;
 assign wire7659 = ( I370 ) | ( I369 ) ;
 assign I369 = ( wire7602*  &  wire7479* ) ;
 assign I370 = ( wire7654*  &  wire7604* ) ;
 assign new_C<101> = ( wire7659 ) | ( wire2017 ) | ( wire7657 ) | ( wire2014 ) ;
 assign wire2008 = ( wire7600*  &  wire7479* ) ;
 assign wire7484 = ( C<98>* ) ;
 assign wire7662 = ( I376 ) | ( I375 ) ;
 assign I375 = ( wire7597*  &  wire7484* ) ;
 assign I376 = ( wire7656*  &  wire7598* ) ;
 assign wire7665 = ( key<250>* ) ;
 assign wire2011 = ( wire7665*  &  wire7581* ) ;
 assign wire7664 = ( I381 ) | ( I380 ) ;
 assign I380 = ( wire7645*  &  wire7602* ) ;
 assign I381 = ( wire7660*  &  wire7604* ) ;
 assign new_C<100> = ( wire7664 ) | ( wire2011 ) | ( wire7662 ) | ( wire2008 ) ;
 assign wire2002 = ( wire7645*  &  wire7600* ) ;
 assign wire7492 = ( C<97>* ) ;
 assign wire7667 = ( I387 ) | ( I386 ) ;
 assign I386 = ( wire7597*  &  wire7492* ) ;
 assign I387 = ( wire7598*  &  wire7484* ) ;
 assign wire7670 = ( key<193>* ) ;
 assign wire2005 = ( wire7670*  &  wire7581* ) ;
 assign wire7669 = ( I392 ) | ( I391 ) ;
 assign I391 = ( wire7602*  &  wire7491* ) ;
 assign I392 = ( wire7665*  &  wire7604* ) ;
 assign new_C<99> = ( wire7669 ) | ( wire2005 ) | ( wire7667 ) | ( wire2002 ) ;
 assign wire1996 = ( wire7600*  &  wire7491* ) ;
 assign wire7471 = ( C<96>* ) ;
 assign wire7672 = ( I398 ) | ( I397 ) ;
 assign I397 = ( wire7597*  &  wire7471* ) ;
 assign I398 = ( wire7598*  &  wire7492* ) ;
 assign wire7675 = ( key<201>* ) ;
 assign wire1999 = ( wire7675*  &  wire7581* ) ;
 assign wire7674 = ( I403 ) | ( I402 ) ;
 assign I402 = ( wire7656*  &  wire7602* ) ;
 assign I403 = ( wire7670*  &  wire7604* ) ;
 assign new_C<98> = ( wire7674 ) | ( wire1999 ) | ( wire7672 ) | ( wire1996 ) ;
 assign wire1990 = ( wire7656*  &  wire7600* ) ;
 assign wire7478 = ( C<95>* ) ;
 assign wire7677 = ( I409 ) | ( I408 ) ;
 assign I408 = ( wire7597*  &  wire7478* ) ;
 assign I409 = ( wire7598*  &  wire7471* ) ;
 assign wire7680 = ( key<209>* ) ;
 assign wire1993 = ( wire7680*  &  wire7581* ) ;
 assign wire7679 = ( I414 ) | ( I413 ) ;
 assign I413 = ( wire7602*  &  wire7484* ) ;
 assign I414 = ( wire7675*  &  wire7604* ) ;
 assign new_C<97> = ( wire7679 ) | ( wire1993 ) | ( wire7677 ) | ( wire1990 ) ;
 assign wire1984 = ( wire7600*  &  wire7484* ) ;
 assign wire7490 = ( C<94>* ) ;
 assign wire7682 = ( I420 ) | ( I419 ) ;
 assign I419 = ( wire7597*  &  wire7490* ) ;
 assign I420 = ( wire7598*  &  wire7478* ) ;
 assign wire7685 = ( key<217>* ) ;
 assign wire1987 = ( wire7685*  &  wire7581* ) ;
 assign wire7684 = ( I425 ) | ( I424 ) ;
 assign I424 = ( wire7602*  &  wire7492* ) ;
 assign I425 = ( wire7680*  &  wire7604* ) ;
 assign new_C<96> = ( wire7684 ) | ( wire1987 ) | ( wire7682 ) | ( wire1984 ) ;
 assign wire1978 = ( wire7600*  &  wire7492* ) ;
 assign wire7481 = ( C<93>* ) ;
 assign wire7687 = ( I431 ) | ( I430 ) ;
 assign I430 = ( wire7597*  &  wire7481* ) ;
 assign I431 = ( wire7598*  &  wire7490* ) ;
 assign wire7690 = ( key<225>* ) ;
 assign wire1981 = ( wire7690*  &  wire7581* ) ;
 assign wire7689 = ( I436 ) | ( I435 ) ;
 assign I435 = ( wire7602*  &  wire7471* ) ;
 assign I436 = ( wire7685*  &  wire7604* ) ;
 assign new_C<95> = ( wire7689 ) | ( wire1981 ) | ( wire7687 ) | ( wire1978 ) ;
 assign wire1972 = ( wire7600*  &  wire7471* ) ;
 assign wire7692 = ( C<92>* ) ;
 assign wire7693 = ( I442 ) | ( I441 ) ;
 assign I441 = ( wire7692*  &  wire7597* ) ;
 assign I442 = ( wire7598*  &  wire7481* ) ;
 assign wire7696 = ( key<233>* ) ;
 assign wire1975 = ( wire7696*  &  wire7581* ) ;
 assign wire7695 = ( I447 ) | ( I446 ) ;
 assign I446 = ( wire7602*  &  wire7478* ) ;
 assign I447 = ( wire7690*  &  wire7604* ) ;
 assign new_C<94> = ( wire7695 ) | ( wire1975 ) | ( wire7693 ) | ( wire1972 ) ;
 assign wire1966 = ( wire7600*  &  wire7478* ) ;
 assign wire7476 = ( C<91>* ) ;
 assign wire7698 = ( I453 ) | ( I452 ) ;
 assign I452 = ( wire7597*  &  wire7476* ) ;
 assign I453 = ( wire7692*  &  wire7598* ) ;
 assign wire7701 = ( key<241>* ) ;
 assign wire1969 = ( wire7701*  &  wire7581* ) ;
 assign wire7700 = ( I458 ) | ( I457 ) ;
 assign I457 = ( wire7602*  &  wire7490* ) ;
 assign I458 = ( wire7696*  &  wire7604* ) ;
 assign new_C<93> = ( wire7700 ) | ( wire1969 ) | ( wire7698 ) | ( wire1966 ) ;
 assign wire1960 = ( wire7600*  &  wire7490* ) ;
 assign wire7474 = ( C<90>* ) ;
 assign wire7703 = ( I464 ) | ( I463 ) ;
 assign I463 = ( wire7597*  &  wire7474* ) ;
 assign I464 = ( wire7598*  &  wire7476* ) ;
 assign wire7706 = ( key<249>* ) ;
 assign wire1963 = ( wire7706*  &  wire7581* ) ;
 assign wire7705 = ( I469 ) | ( I468 ) ;
 assign I468 = ( wire7602*  &  wire7481* ) ;
 assign I469 = ( wire7701*  &  wire7604* ) ;
 assign new_C<92> = ( wire7705 ) | ( wire1963 ) | ( wire7703 ) | ( wire1960 ) ;
 assign wire1954 = ( wire7600*  &  wire7481* ) ;
 assign wire7483 = ( C<89>* ) ;
 assign wire7708 = ( I475 ) | ( I474 ) ;
 assign I474 = ( wire7597*  &  wire7483* ) ;
 assign I475 = ( wire7598*  &  wire7474* ) ;
 assign wire7711 = ( key<192>* ) ;
 assign wire1957 = ( wire7711*  &  wire7581* ) ;
 assign wire7710 = ( I480 ) | ( I479 ) ;
 assign I479 = ( wire7692*  &  wire7602* ) ;
 assign I480 = ( wire7706*  &  wire7604* ) ;
 assign new_C<91> = ( wire7710 ) | ( wire1957 ) | ( wire7708 ) | ( wire1954 ) ;
 assign wire1948 = ( wire7692*  &  wire7600* ) ;
 assign wire7487 = ( C<88>* ) ;
 assign wire7713 = ( I486 ) | ( I485 ) ;
 assign I485 = ( wire7597*  &  wire7487* ) ;
 assign I486 = ( wire7598*  &  wire7483* ) ;
 assign wire7716 = ( key<200>* ) ;
 assign wire1951 = ( wire7716*  &  wire7581* ) ;
 assign wire7715 = ( I491 ) | ( I490 ) ;
 assign I490 = ( wire7602*  &  wire7476* ) ;
 assign I491 = ( wire7711*  &  wire7604* ) ;
 assign new_C<90> = ( wire7715 ) | ( wire1951 ) | ( wire7713 ) | ( wire1948 ) ;
 assign wire1942 = ( wire7600*  &  wire7476* ) ;
 assign wire7477 = ( C<87>* ) ;
 assign wire7718 = ( I497 ) | ( I496 ) ;
 assign I496 = ( wire7597*  &  wire7477* ) ;
 assign I497 = ( wire7598*  &  wire7487* ) ;
 assign wire7721 = ( key<208>* ) ;
 assign wire1945 = ( wire7721*  &  wire7581* ) ;
 assign wire7720 = ( I502 ) | ( I501 ) ;
 assign I501 = ( wire7602*  &  wire7474* ) ;
 assign I502 = ( wire7716*  &  wire7604* ) ;
 assign new_C<89> = ( wire7720 ) | ( wire1945 ) | ( wire7718 ) | ( wire1942 ) ;
 assign wire1936 = ( wire7600*  &  wire7474* ) ;
 assign wire7486 = ( C<86>* ) ;
 assign wire7723 = ( I508 ) | ( I507 ) ;
 assign I507 = ( wire7597*  &  wire7486* ) ;
 assign I508 = ( wire7598*  &  wire7477* ) ;
 assign wire7726 = ( key<216>* ) ;
 assign wire1939 = ( wire7726*  &  wire7581* ) ;
 assign wire7725 = ( I513 ) | ( I512 ) ;
 assign I512 = ( wire7602*  &  wire7483* ) ;
 assign I513 = ( wire7721*  &  wire7604* ) ;
 assign new_C<88> = ( wire7725 ) | ( wire1939 ) | ( wire7723 ) | ( wire1936 ) ;
 assign wire1930 = ( wire7600*  &  wire7483* ) ;
 assign wire7470 = ( C<85>* ) ;
 assign wire7728 = ( I519 ) | ( I518 ) ;
 assign I518 = ( wire7597*  &  wire7470* ) ;
 assign I519 = ( wire7598*  &  wire7486* ) ;
 assign wire7731 = ( key<224>* ) ;
 assign wire1933 = ( wire7731*  &  wire7581* ) ;
 assign wire7730 = ( I524 ) | ( I523 ) ;
 assign I523 = ( wire7602*  &  wire7487* ) ;
 assign I524 = ( wire7726*  &  wire7604* ) ;
 assign new_C<87> = ( wire7730 ) | ( wire1933 ) | ( wire7728 ) | ( wire1930 ) ;
 assign wire1924 = ( wire7600*  &  wire7487* ) ;
 assign wire7488 = ( C<84>* ) ;
 assign wire7733 = ( I530 ) | ( I529 ) ;
 assign I529 = ( wire7597*  &  wire7488* ) ;
 assign I530 = ( wire7598*  &  wire7470* ) ;
 assign wire7736 = ( key<232>* ) ;
 assign wire1927 = ( wire7736*  &  wire7581* ) ;
 assign wire7735 = ( I535 ) | ( I534 ) ;
 assign I534 = ( wire7602*  &  wire7477* ) ;
 assign I535 = ( wire7731*  &  wire7604* ) ;
 assign new_C<86> = ( wire7735 ) | ( wire1927 ) | ( wire7733 ) | ( wire1924 ) ;
 assign wire1918 = ( wire7600*  &  wire7477* ) ;
 assign wire7509 = ( C<83>* ) ;
 assign wire7738 = ( I541 ) | ( I540 ) ;
 assign I540 = ( wire7597*  &  wire7509* ) ;
 assign I541 = ( wire7598*  &  wire7488* ) ;
 assign wire7741 = ( key<240>* ) ;
 assign wire1921 = ( wire7741*  &  wire7581* ) ;
 assign wire7740 = ( I546 ) | ( I545 ) ;
 assign I545 = ( wire7602*  &  wire7486* ) ;
 assign I546 = ( wire7736*  &  wire7604* ) ;
 assign new_C<85> = ( wire7740 ) | ( wire1921 ) | ( wire7738 ) | ( wire1918 ) ;
 assign wire1912 = ( wire7600*  &  wire7486* ) ;
 assign wire7496 = ( C<82>* ) ;
 assign wire7743 = ( I552 ) | ( I551 ) ;
 assign I551 = ( wire7597*  &  wire7496* ) ;
 assign I552 = ( wire7598*  &  wire7509* ) ;
 assign wire7746 = ( key<248>* ) ;
 assign wire1915 = ( wire7746*  &  wire7581* ) ;
 assign wire7745 = ( I557 ) | ( I556 ) ;
 assign I556 = ( wire7602*  &  wire7470* ) ;
 assign I557 = ( wire7741*  &  wire7604* ) ;
 assign new_C<84> = ( wire7745 ) | ( wire1915 ) | ( wire7743 ) | ( wire1912 ) ;
 assign wire1906 = ( wire7600*  &  wire7470* ) ;
 assign wire7500 = ( C<81>* ) ;
 assign wire7748 = ( I563 ) | ( I562 ) ;
 assign I562 = ( wire7597*  &  wire7500* ) ;
 assign I563 = ( wire7598*  &  wire7496* ) ;
 assign wire7751 = ( key<163>* ) ;
 assign wire1909 = ( wire7751*  &  wire7581* ) ;
 assign wire7750 = ( I568 ) | ( I567 ) ;
 assign I567 = ( wire7602*  &  wire7488* ) ;
 assign I568 = ( wire7746*  &  wire7604* ) ;
 assign new_C<83> = ( wire7750 ) | ( wire1909 ) | ( wire7748 ) | ( wire1906 ) ;
 assign wire1900 = ( wire7600*  &  wire7488* ) ;
 assign wire7753 = ( C<80>* ) ;
 assign wire7754 = ( I574 ) | ( I573 ) ;
 assign I573 = ( wire7753*  &  wire7597* ) ;
 assign I574 = ( wire7598*  &  wire7500* ) ;
 assign wire7757 = ( key<171>* ) ;
 assign wire1903 = ( wire7757*  &  wire7581* ) ;
 assign wire7756 = ( I579 ) | ( I578 ) ;
 assign I578 = ( wire7602*  &  wire7509* ) ;
 assign I579 = ( wire7751*  &  wire7604* ) ;
 assign new_C<82> = ( wire7756 ) | ( wire1903 ) | ( wire7754 ) | ( wire1900 ) ;
 assign wire1894 = ( wire7600*  &  wire7509* ) ;
 assign wire7513 = ( C<79>* ) ;
 assign wire7759 = ( I585 ) | ( I584 ) ;
 assign I584 = ( wire7597*  &  wire7513* ) ;
 assign I585 = ( wire7753*  &  wire7598* ) ;
 assign wire7762 = ( key<179>* ) ;
 assign wire1897 = ( wire7762*  &  wire7581* ) ;
 assign wire7761 = ( I590 ) | ( I589 ) ;
 assign I589 = ( wire7602*  &  wire7496* ) ;
 assign I590 = ( wire7757*  &  wire7604* ) ;
 assign new_C<81> = ( wire7761 ) | ( wire1897 ) | ( wire7759 ) | ( wire1894 ) ;
 assign wire1888 = ( wire7600*  &  wire7496* ) ;
 assign wire7504 = ( C<78>* ) ;
 assign wire7764 = ( I596 ) | ( I595 ) ;
 assign I595 = ( wire7597*  &  wire7504* ) ;
 assign I596 = ( wire7598*  &  wire7513* ) ;
 assign wire7767 = ( key<187>* ) ;
 assign wire1891 = ( wire7767*  &  wire7581* ) ;
 assign wire7766 = ( I601 ) | ( I600 ) ;
 assign I600 = ( wire7602*  &  wire7500* ) ;
 assign I601 = ( wire7762*  &  wire7604* ) ;
 assign new_C<80> = ( wire7766 ) | ( wire1891 ) | ( wire7764 ) | ( wire1888 ) ;
 assign wire1882 = ( wire7600*  &  wire7500* ) ;
 assign wire7769 = ( C<77>* ) ;
 assign wire7770 = ( I607 ) | ( I606 ) ;
 assign I606 = ( wire7769*  &  wire7597* ) ;
 assign I607 = ( wire7598*  &  wire7504* ) ;
 assign wire7773 = ( key<130>* ) ;
 assign wire1885 = ( wire7773*  &  wire7581* ) ;
 assign wire7772 = ( I612 ) | ( I611 ) ;
 assign I611 = ( wire7753*  &  wire7602* ) ;
 assign I612 = ( wire7767*  &  wire7604* ) ;
 assign new_C<79> = ( wire7772 ) | ( wire1885 ) | ( wire7770 ) | ( wire1882 ) ;
 assign wire1876 = ( wire7753*  &  wire7600* ) ;
 assign wire7506 = ( C<76>* ) ;
 assign wire7775 = ( I618 ) | ( I617 ) ;
 assign I617 = ( wire7597*  &  wire7506* ) ;
 assign I618 = ( wire7769*  &  wire7598* ) ;
 assign wire7778 = ( key<138>* ) ;
 assign wire1879 = ( wire7778*  &  wire7581* ) ;
 assign wire7777 = ( I623 ) | ( I622 ) ;
 assign I622 = ( wire7602*  &  wire7513* ) ;
 assign I623 = ( wire7773*  &  wire7604* ) ;
 assign new_C<78> = ( wire7777 ) | ( wire1879 ) | ( wire7775 ) | ( wire1876 ) ;
 assign wire1870 = ( wire7600*  &  wire7513* ) ;
 assign wire7495 = ( C<75>* ) ;
 assign wire7780 = ( I629 ) | ( I628 ) ;
 assign I628 = ( wire7597*  &  wire7495* ) ;
 assign I629 = ( wire7598*  &  wire7506* ) ;
 assign wire7783 = ( key<146>* ) ;
 assign wire1873 = ( wire7783*  &  wire7581* ) ;
 assign wire7782 = ( I634 ) | ( I633 ) ;
 assign I633 = ( wire7602*  &  wire7504* ) ;
 assign I634 = ( wire7778*  &  wire7604* ) ;
 assign new_C<77> = ( wire7782 ) | ( wire1873 ) | ( wire7780 ) | ( wire1870 ) ;
 assign wire1864 = ( wire7600*  &  wire7504* ) ;
 assign wire7503 = ( C<74>* ) ;
 assign wire7785 = ( I640 ) | ( I639 ) ;
 assign I639 = ( wire7597*  &  wire7503* ) ;
 assign I640 = ( wire7598*  &  wire7495* ) ;
 assign wire7788 = ( key<154>* ) ;
 assign wire1867 = ( wire7788*  &  wire7581* ) ;
 assign wire7787 = ( I645 ) | ( I644 ) ;
 assign I644 = ( wire7769*  &  wire7602* ) ;
 assign I645 = ( wire7783*  &  wire7604* ) ;
 assign new_C<76> = ( wire7787 ) | ( wire1867 ) | ( wire7785 ) | ( wire1864 ) ;
 assign wire1858 = ( wire7769*  &  wire7600* ) ;
 assign wire7790 = ( C<73>* ) ;
 assign wire7791 = ( I651 ) | ( I650 ) ;
 assign I650 = ( wire7790*  &  wire7597* ) ;
 assign I651 = ( wire7598*  &  wire7503* ) ;
 assign wire7794 = ( key<162>* ) ;
 assign wire1861 = ( wire7794*  &  wire7581* ) ;
 assign wire7793 = ( I656 ) | ( I655 ) ;
 assign I655 = ( wire7602*  &  wire7506* ) ;
 assign I656 = ( wire7788*  &  wire7604* ) ;
 assign new_C<75> = ( wire7793 ) | ( wire1861 ) | ( wire7791 ) | ( wire1858 ) ;
 assign wire1852 = ( wire7600*  &  wire7506* ) ;
 assign wire7515 = ( C<72>* ) ;
 assign wire7796 = ( I662 ) | ( I661 ) ;
 assign I661 = ( wire7597*  &  wire7515* ) ;
 assign I662 = ( wire7790*  &  wire7598* ) ;
 assign wire7799 = ( key<170>* ) ;
 assign wire1855 = ( wire7799*  &  wire7581* ) ;
 assign wire7798 = ( I667 ) | ( I666 ) ;
 assign I666 = ( wire7602*  &  wire7495* ) ;
 assign I667 = ( wire7794*  &  wire7604* ) ;
 assign new_C<74> = ( wire7798 ) | ( wire1855 ) | ( wire7796 ) | ( wire1852 ) ;
 assign wire1846 = ( wire7600*  &  wire7495* ) ;
 assign wire7498 = ( C<71>* ) ;
 assign wire7801 = ( I673 ) | ( I672 ) ;
 assign I672 = ( wire7597*  &  wire7498* ) ;
 assign I673 = ( wire7598*  &  wire7515* ) ;
 assign wire7804 = ( key<178>* ) ;
 assign wire1849 = ( wire7804*  &  wire7581* ) ;
 assign wire7803 = ( I678 ) | ( I677 ) ;
 assign I677 = ( wire7602*  &  wire7503* ) ;
 assign I678 = ( wire7799*  &  wire7604* ) ;
 assign new_C<73> = ( wire7803 ) | ( wire1849 ) | ( wire7801 ) | ( wire1846 ) ;
 assign wire1840 = ( wire7600*  &  wire7503* ) ;
 assign wire7508 = ( C<70>* ) ;
 assign wire7806 = ( I684 ) | ( I683 ) ;
 assign I683 = ( wire7597*  &  wire7508* ) ;
 assign I684 = ( wire7598*  &  wire7498* ) ;
 assign wire7809 = ( key<186>* ) ;
 assign wire1843 = ( wire7809*  &  wire7581* ) ;
 assign wire7808 = ( I689 ) | ( I688 ) ;
 assign I688 = ( wire7790*  &  wire7602* ) ;
 assign I689 = ( wire7804*  &  wire7604* ) ;
 assign new_C<72> = ( wire7808 ) | ( wire1843 ) | ( wire7806 ) | ( wire1840 ) ;
 assign wire1834 = ( wire7790*  &  wire7600* ) ;
 assign wire7516 = ( C<69>* ) ;
 assign wire7811 = ( I695 ) | ( I694 ) ;
 assign I694 = ( wire7597*  &  wire7516* ) ;
 assign I695 = ( wire7598*  &  wire7508* ) ;
 assign wire7814 = ( key<129>* ) ;
 assign wire1837 = ( wire7814*  &  wire7581* ) ;
 assign wire7813 = ( I700 ) | ( I699 ) ;
 assign I699 = ( wire7602*  &  wire7515* ) ;
 assign I700 = ( wire7809*  &  wire7604* ) ;
 assign new_C<71> = ( wire7813 ) | ( wire1837 ) | ( wire7811 ) | ( wire1834 ) ;
 assign wire1828 = ( wire7600*  &  wire7515* ) ;
 assign wire7494 = ( C<68>* ) ;
 assign wire7816 = ( I706 ) | ( I705 ) ;
 assign I705 = ( wire7597*  &  wire7494* ) ;
 assign I706 = ( wire7598*  &  wire7516* ) ;
 assign wire7819 = ( key<137>* ) ;
 assign wire1831 = ( wire7819*  &  wire7581* ) ;
 assign wire7818 = ( I711 ) | ( I710 ) ;
 assign I710 = ( wire7602*  &  wire7498* ) ;
 assign I711 = ( wire7814*  &  wire7604* ) ;
 assign new_C<70> = ( wire7818 ) | ( wire1831 ) | ( wire7816 ) | ( wire1828 ) ;
 assign wire1822 = ( wire7600*  &  wire7498* ) ;
 assign wire7502 = ( C<67>* ) ;
 assign wire7821 = ( I717 ) | ( I716 ) ;
 assign I716 = ( wire7597*  &  wire7502* ) ;
 assign I717 = ( wire7598*  &  wire7494* ) ;
 assign wire7824 = ( key<145>* ) ;
 assign wire1825 = ( wire7824*  &  wire7581* ) ;
 assign wire7823 = ( I722 ) | ( I721 ) ;
 assign I721 = ( wire7602*  &  wire7508* ) ;
 assign I722 = ( wire7819*  &  wire7604* ) ;
 assign new_C<69> = ( wire7823 ) | ( wire1825 ) | ( wire7821 ) | ( wire1822 ) ;
 assign wire1816 = ( wire7600*  &  wire7508* ) ;
 assign wire7514 = ( C<66>* ) ;
 assign wire7826 = ( I728 ) | ( I727 ) ;
 assign I727 = ( wire7597*  &  wire7514* ) ;
 assign I728 = ( wire7598*  &  wire7502* ) ;
 assign wire7829 = ( key<153>* ) ;
 assign wire1819 = ( wire7829*  &  wire7581* ) ;
 assign wire7828 = ( I733 ) | ( I732 ) ;
 assign I732 = ( wire7602*  &  wire7516* ) ;
 assign I733 = ( wire7824*  &  wire7604* ) ;
 assign new_C<68> = ( wire7828 ) | ( wire1819 ) | ( wire7826 ) | ( wire1816 ) ;
 assign wire1810 = ( wire7600*  &  wire7516* ) ;
 assign wire7505 = ( C<65>* ) ;
 assign wire7831 = ( I739 ) | ( I738 ) ;
 assign I738 = ( wire7597*  &  wire7505* ) ;
 assign I739 = ( wire7598*  &  wire7514* ) ;
 assign wire7834 = ( key<161>* ) ;
 assign wire1813 = ( wire7834*  &  wire7581* ) ;
 assign wire7833 = ( I744 ) | ( I743 ) ;
 assign I743 = ( wire7602*  &  wire7494* ) ;
 assign I744 = ( wire7829*  &  wire7604* ) ;
 assign new_C<67> = ( wire7833 ) | ( wire1813 ) | ( wire7831 ) | ( wire1810 ) ;
 assign wire1804 = ( wire7600*  &  wire7494* ) ;
 assign wire7836 = ( C<64>* ) ;
 assign wire7837 = ( I750 ) | ( I749 ) ;
 assign I749 = ( wire7836*  &  wire7597* ) ;
 assign I750 = ( wire7598*  &  wire7505* ) ;
 assign wire7840 = ( key<169>* ) ;
 assign wire1807 = ( wire7840*  &  wire7581* ) ;
 assign wire7839 = ( I755 ) | ( I754 ) ;
 assign I754 = ( wire7602*  &  wire7502* ) ;
 assign I755 = ( wire7834*  &  wire7604* ) ;
 assign new_C<66> = ( wire7839 ) | ( wire1807 ) | ( wire7837 ) | ( wire1804 ) ;
 assign wire1798 = ( wire7600*  &  wire7502* ) ;
 assign wire7499 = ( C<63>* ) ;
 assign wire7842 = ( I761 ) | ( I760 ) ;
 assign I760 = ( wire7597*  &  wire7499* ) ;
 assign I761 = ( wire7836*  &  wire7598* ) ;
 assign wire7845 = ( key<177>* ) ;
 assign wire1801 = ( wire7845*  &  wire7581* ) ;
 assign wire7844 = ( I766 ) | ( I765 ) ;
 assign I765 = ( wire7602*  &  wire7514* ) ;
 assign I766 = ( wire7840*  &  wire7604* ) ;
 assign new_C<65> = ( wire7844 ) | ( wire1801 ) | ( wire7842 ) | ( wire1798 ) ;
 assign wire1792 = ( wire7600*  &  wire7514* ) ;
 assign wire7497 = ( C<62>* ) ;
 assign wire7847 = ( I772 ) | ( I771 ) ;
 assign I771 = ( wire7597*  &  wire7497* ) ;
 assign I772 = ( wire7598*  &  wire7499* ) ;
 assign wire7850 = ( key<185>* ) ;
 assign wire1795 = ( wire7850*  &  wire7581* ) ;
 assign wire7849 = ( I777 ) | ( I776 ) ;
 assign I776 = ( wire7602*  &  wire7505* ) ;
 assign I777 = ( wire7845*  &  wire7604* ) ;
 assign new_C<64> = ( wire7849 ) | ( wire1795 ) | ( wire7847 ) | ( wire1792 ) ;
 assign wire1786 = ( wire7600*  &  wire7505* ) ;
 assign wire7507 = ( C<61>* ) ;
 assign wire7852 = ( I783 ) | ( I782 ) ;
 assign I782 = ( wire7597*  &  wire7507* ) ;
 assign I783 = ( wire7598*  &  wire7497* ) ;
 assign wire7855 = ( key<128>* ) ;
 assign wire1789 = ( wire7855*  &  wire7581* ) ;
 assign wire7854 = ( I788 ) | ( I787 ) ;
 assign I787 = ( wire7836*  &  wire7602* ) ;
 assign I788 = ( wire7850*  &  wire7604* ) ;
 assign new_C<63> = ( wire7854 ) | ( wire1789 ) | ( wire7852 ) | ( wire1786 ) ;
 assign wire1780 = ( wire7836*  &  wire7600* ) ;
 assign wire7511 = ( C<60>* ) ;
 assign wire7857 = ( I794 ) | ( I793 ) ;
 assign I793 = ( wire7597*  &  wire7511* ) ;
 assign I794 = ( wire7598*  &  wire7507* ) ;
 assign wire7860 = ( key<136>* ) ;
 assign wire1783 = ( wire7860*  &  wire7581* ) ;
 assign wire7859 = ( I799 ) | ( I798 ) ;
 assign I798 = ( wire7602*  &  wire7499* ) ;
 assign I799 = ( wire7855*  &  wire7604* ) ;
 assign new_C<62> = ( wire7859 ) | ( wire1783 ) | ( wire7857 ) | ( wire1780 ) ;
 assign wire1774 = ( wire7600*  &  wire7499* ) ;
 assign wire7501 = ( C<59>* ) ;
 assign wire7862 = ( I805 ) | ( I804 ) ;
 assign I804 = ( wire7597*  &  wire7501* ) ;
 assign I805 = ( wire7598*  &  wire7511* ) ;
 assign wire7865 = ( key<144>* ) ;
 assign wire1777 = ( wire7865*  &  wire7581* ) ;
 assign wire7864 = ( I810 ) | ( I809 ) ;
 assign I809 = ( wire7602*  &  wire7497* ) ;
 assign I810 = ( wire7860*  &  wire7604* ) ;
 assign new_C<61> = ( wire7864 ) | ( wire1777 ) | ( wire7862 ) | ( wire1774 ) ;
 assign wire1768 = ( wire7600*  &  wire7497* ) ;
 assign wire7510 = ( C<58>* ) ;
 assign wire7867 = ( I816 ) | ( I815 ) ;
 assign I815 = ( wire7597*  &  wire7510* ) ;
 assign I816 = ( wire7598*  &  wire7501* ) ;
 assign wire7870 = ( key<152>* ) ;
 assign wire1771 = ( wire7870*  &  wire7581* ) ;
 assign wire7869 = ( I821 ) | ( I820 ) ;
 assign I820 = ( wire7602*  &  wire7507* ) ;
 assign I821 = ( wire7865*  &  wire7604* ) ;
 assign new_C<60> = ( wire7869 ) | ( wire1771 ) | ( wire7867 ) | ( wire1768 ) ;
 assign wire1762 = ( wire7600*  &  wire7507* ) ;
 assign wire7493 = ( C<57>* ) ;
 assign wire7872 = ( I827 ) | ( I826 ) ;
 assign I826 = ( wire7597*  &  wire7493* ) ;
 assign I827 = ( wire7598*  &  wire7510* ) ;
 assign wire7875 = ( key<160>* ) ;
 assign wire1765 = ( wire7875*  &  wire7581* ) ;
 assign wire7874 = ( I832 ) | ( I831 ) ;
 assign I831 = ( wire7602*  &  wire7511* ) ;
 assign I832 = ( wire7870*  &  wire7604* ) ;
 assign new_C<59> = ( wire7874 ) | ( wire1765 ) | ( wire7872 ) | ( wire1762 ) ;
 assign wire1756 = ( wire7600*  &  wire7511* ) ;
 assign wire7512 = ( C<56>* ) ;
 assign wire7877 = ( I838 ) | ( I837 ) ;
 assign I837 = ( wire7597*  &  wire7512* ) ;
 assign I838 = ( wire7598*  &  wire7493* ) ;
 assign wire7880 = ( key<168>* ) ;
 assign wire1759 = ( wire7880*  &  wire7581* ) ;
 assign wire7879 = ( I843 ) | ( I842 ) ;
 assign I842 = ( wire7602*  &  wire7501* ) ;
 assign I843 = ( wire7875*  &  wire7604* ) ;
 assign new_C<58> = ( wire7879 ) | ( wire1759 ) | ( wire7877 ) | ( wire1756 ) ;
 assign wire1750 = ( wire7600*  &  wire7501* ) ;
 assign wire7533 = ( C<55>* ) ;
 assign wire7882 = ( I849 ) | ( I848 ) ;
 assign I848 = ( wire7597*  &  wire7533* ) ;
 assign I849 = ( wire7598*  &  wire7512* ) ;
 assign wire7885 = ( key<176>* ) ;
 assign wire1753 = ( wire7885*  &  wire7581* ) ;
 assign wire7884 = ( I854 ) | ( I853 ) ;
 assign I853 = ( wire7602*  &  wire7510* ) ;
 assign I854 = ( wire7880*  &  wire7604* ) ;
 assign new_C<57> = ( wire7884 ) | ( wire1753 ) | ( wire7882 ) | ( wire1750 ) ;
 assign wire1744 = ( wire7600*  &  wire7510* ) ;
 assign wire7520 = ( C<54>* ) ;
 assign wire7887 = ( I860 ) | ( I859 ) ;
 assign I859 = ( wire7597*  &  wire7520* ) ;
 assign I860 = ( wire7598*  &  wire7533* ) ;
 assign wire7890 = ( key<184>* ) ;
 assign wire1747 = ( wire7890*  &  wire7581* ) ;
 assign wire7889 = ( I865 ) | ( I864 ) ;
 assign I864 = ( wire7602*  &  wire7493* ) ;
 assign I865 = ( wire7885*  &  wire7604* ) ;
 assign new_C<56> = ( wire7889 ) | ( wire1747 ) | ( wire7887 ) | ( wire1744 ) ;
 assign wire1738 = ( wire7600*  &  wire7493* ) ;
 assign wire7524 = ( C<53>* ) ;
 assign wire7892 = ( I871 ) | ( I870 ) ;
 assign I870 = ( wire7597*  &  wire7524* ) ;
 assign I871 = ( wire7598*  &  wire7520* ) ;
 assign wire7895 = ( key<99>* ) ;
 assign wire1741 = ( wire7895*  &  wire7581* ) ;
 assign wire7894 = ( I876 ) | ( I875 ) ;
 assign I875 = ( wire7602*  &  wire7512* ) ;
 assign I876 = ( wire7890*  &  wire7604* ) ;
 assign new_C<55> = ( wire7894 ) | ( wire1741 ) | ( wire7892 ) | ( wire1738 ) ;
 assign wire1732 = ( wire7600*  &  wire7512* ) ;
 assign wire7897 = ( C<52>* ) ;
 assign wire7898 = ( I882 ) | ( I881 ) ;
 assign I881 = ( wire7897*  &  wire7597* ) ;
 assign I882 = ( wire7598*  &  wire7524* ) ;
 assign wire7901 = ( key<107>* ) ;
 assign wire1735 = ( wire7901*  &  wire7581* ) ;
 assign wire7900 = ( I887 ) | ( I886 ) ;
 assign I886 = ( wire7602*  &  wire7533* ) ;
 assign I887 = ( wire7895*  &  wire7604* ) ;
 assign new_C<54> = ( wire7900 ) | ( wire1735 ) | ( wire7898 ) | ( wire1732 ) ;
 assign wire1726 = ( wire7600*  &  wire7533* ) ;
 assign wire7537 = ( C<51>* ) ;
 assign wire7903 = ( I893 ) | ( I892 ) ;
 assign I892 = ( wire7597*  &  wire7537* ) ;
 assign I893 = ( wire7897*  &  wire7598* ) ;
 assign wire7906 = ( key<115>* ) ;
 assign wire1729 = ( wire7906*  &  wire7581* ) ;
 assign wire7905 = ( I898 ) | ( I897 ) ;
 assign I897 = ( wire7602*  &  wire7520* ) ;
 assign I898 = ( wire7901*  &  wire7604* ) ;
 assign new_C<53> = ( wire7905 ) | ( wire1729 ) | ( wire7903 ) | ( wire1726 ) ;
 assign wire1720 = ( wire7600*  &  wire7520* ) ;
 assign wire7528 = ( C<50>* ) ;
 assign wire7908 = ( I904 ) | ( I903 ) ;
 assign I903 = ( wire7597*  &  wire7528* ) ;
 assign I904 = ( wire7598*  &  wire7537* ) ;
 assign wire7911 = ( key<123>* ) ;
 assign wire1723 = ( wire7911*  &  wire7581* ) ;
 assign wire7910 = ( I909 ) | ( I908 ) ;
 assign I908 = ( wire7602*  &  wire7524* ) ;
 assign I909 = ( wire7906*  &  wire7604* ) ;
 assign new_C<52> = ( wire7910 ) | ( wire1723 ) | ( wire7908 ) | ( wire1720 ) ;
 assign wire1714 = ( wire7600*  &  wire7524* ) ;
 assign wire7913 = ( C<49>* ) ;
 assign wire7914 = ( I915 ) | ( I914 ) ;
 assign I914 = ( wire7913*  &  wire7597* ) ;
 assign I915 = ( wire7598*  &  wire7528* ) ;
 assign wire7917 = ( key<66>* ) ;
 assign wire1717 = ( wire7917*  &  wire7581* ) ;
 assign wire7916 = ( I920 ) | ( I919 ) ;
 assign I919 = ( wire7897*  &  wire7602* ) ;
 assign I920 = ( wire7911*  &  wire7604* ) ;
 assign new_C<51> = ( wire7916 ) | ( wire1717 ) | ( wire7914 ) | ( wire1714 ) ;
 assign wire1708 = ( wire7897*  &  wire7600* ) ;
 assign wire7530 = ( C<48>* ) ;
 assign wire7919 = ( I926 ) | ( I925 ) ;
 assign I925 = ( wire7597*  &  wire7530* ) ;
 assign I926 = ( wire7913*  &  wire7598* ) ;
 assign wire7922 = ( key<74>* ) ;
 assign wire1711 = ( wire7922*  &  wire7581* ) ;
 assign wire7921 = ( I931 ) | ( I930 ) ;
 assign I930 = ( wire7602*  &  wire7537* ) ;
 assign I931 = ( wire7917*  &  wire7604* ) ;
 assign new_C<50> = ( wire7921 ) | ( wire1711 ) | ( wire7919 ) | ( wire1708 ) ;
 assign wire1702 = ( wire7600*  &  wire7537* ) ;
 assign wire7519 = ( C<47>* ) ;
 assign wire7924 = ( I937 ) | ( I936 ) ;
 assign I936 = ( wire7597*  &  wire7519* ) ;
 assign I937 = ( wire7598*  &  wire7530* ) ;
 assign wire7927 = ( key<82>* ) ;
 assign wire1705 = ( wire7927*  &  wire7581* ) ;
 assign wire7926 = ( I942 ) | ( I941 ) ;
 assign I941 = ( wire7602*  &  wire7528* ) ;
 assign I942 = ( wire7922*  &  wire7604* ) ;
 assign new_C<49> = ( wire7926 ) | ( wire1705 ) | ( wire7924 ) | ( wire1702 ) ;
 assign wire1696 = ( wire7600*  &  wire7528* ) ;
 assign wire7527 = ( C<46>* ) ;
 assign wire7929 = ( I948 ) | ( I947 ) ;
 assign I947 = ( wire7597*  &  wire7527* ) ;
 assign I948 = ( wire7598*  &  wire7519* ) ;
 assign wire7932 = ( key<90>* ) ;
 assign wire1699 = ( wire7932*  &  wire7581* ) ;
 assign wire7931 = ( I953 ) | ( I952 ) ;
 assign I952 = ( wire7913*  &  wire7602* ) ;
 assign I953 = ( wire7927*  &  wire7604* ) ;
 assign new_C<48> = ( wire7931 ) | ( wire1699 ) | ( wire7929 ) | ( wire1696 ) ;
 assign wire1690 = ( wire7913*  &  wire7600* ) ;
 assign wire7934 = ( C<45>* ) ;
 assign wire7935 = ( I959 ) | ( I958 ) ;
 assign I958 = ( wire7934*  &  wire7597* ) ;
 assign I959 = ( wire7598*  &  wire7527* ) ;
 assign wire7938 = ( key<98>* ) ;
 assign wire1693 = ( wire7938*  &  wire7581* ) ;
 assign wire7937 = ( I964 ) | ( I963 ) ;
 assign I963 = ( wire7602*  &  wire7530* ) ;
 assign I964 = ( wire7932*  &  wire7604* ) ;
 assign new_C<47> = ( wire7937 ) | ( wire1693 ) | ( wire7935 ) | ( wire1690 ) ;
 assign wire1684 = ( wire7600*  &  wire7530* ) ;
 assign wire7539 = ( C<44>* ) ;
 assign wire7940 = ( I970 ) | ( I969 ) ;
 assign I969 = ( wire7597*  &  wire7539* ) ;
 assign I970 = ( wire7934*  &  wire7598* ) ;
 assign wire7943 = ( key<106>* ) ;
 assign wire1687 = ( wire7943*  &  wire7581* ) ;
 assign wire7942 = ( I975 ) | ( I974 ) ;
 assign I974 = ( wire7602*  &  wire7519* ) ;
 assign I975 = ( wire7938*  &  wire7604* ) ;
 assign new_C<46> = ( wire7942 ) | ( wire1687 ) | ( wire7940 ) | ( wire1684 ) ;
 assign wire1678 = ( wire7600*  &  wire7519* ) ;
 assign wire7522 = ( C<43>* ) ;
 assign wire7945 = ( I981 ) | ( I980 ) ;
 assign I980 = ( wire7597*  &  wire7522* ) ;
 assign I981 = ( wire7598*  &  wire7539* ) ;
 assign wire7948 = ( key<114>* ) ;
 assign wire1681 = ( wire7948*  &  wire7581* ) ;
 assign wire7947 = ( I986 ) | ( I985 ) ;
 assign I985 = ( wire7602*  &  wire7527* ) ;
 assign I986 = ( wire7943*  &  wire7604* ) ;
 assign new_C<45> = ( wire7947 ) | ( wire1681 ) | ( wire7945 ) | ( wire1678 ) ;
 assign wire1672 = ( wire7600*  &  wire7527* ) ;
 assign wire7532 = ( C<42>* ) ;
 assign wire7950 = ( I992 ) | ( I991 ) ;
 assign I991 = ( wire7597*  &  wire7532* ) ;
 assign I992 = ( wire7598*  &  wire7522* ) ;
 assign wire7953 = ( key<122>* ) ;
 assign wire1675 = ( wire7953*  &  wire7581* ) ;
 assign wire7952 = ( I997 ) | ( I996 ) ;
 assign I996 = ( wire7934*  &  wire7602* ) ;
 assign I997 = ( wire7948*  &  wire7604* ) ;
 assign new_C<44> = ( wire7952 ) | ( wire1675 ) | ( wire7950 ) | ( wire1672 ) ;
 assign wire1666 = ( wire7934*  &  wire7600* ) ;
 assign wire7540 = ( C<41>* ) ;
 assign wire7955 = ( I1003 ) | ( I1002 ) ;
 assign I1002 = ( wire7597*  &  wire7540* ) ;
 assign I1003 = ( wire7598*  &  wire7532* ) ;
 assign wire7958 = ( key<65>* ) ;
 assign wire1669 = ( wire7958*  &  wire7581* ) ;
 assign wire7957 = ( I1008 ) | ( I1007 ) ;
 assign I1007 = ( wire7602*  &  wire7539* ) ;
 assign I1008 = ( wire7953*  &  wire7604* ) ;
 assign new_C<43> = ( wire7957 ) | ( wire1669 ) | ( wire7955 ) | ( wire1666 ) ;
 assign wire1660 = ( wire7600*  &  wire7539* ) ;
 assign wire7518 = ( C<40>* ) ;
 assign wire7960 = ( I1014 ) | ( I1013 ) ;
 assign I1013 = ( wire7597*  &  wire7518* ) ;
 assign I1014 = ( wire7598*  &  wire7540* ) ;
 assign wire7963 = ( key<73>* ) ;
 assign wire1663 = ( wire7963*  &  wire7581* ) ;
 assign wire7962 = ( I1019 ) | ( I1018 ) ;
 assign I1018 = ( wire7602*  &  wire7522* ) ;
 assign I1019 = ( wire7958*  &  wire7604* ) ;
 assign new_C<42> = ( wire7962 ) | ( wire1663 ) | ( wire7960 ) | ( wire1660 ) ;
 assign wire1654 = ( wire7600*  &  wire7522* ) ;
 assign wire7526 = ( C<39>* ) ;
 assign wire7965 = ( I1025 ) | ( I1024 ) ;
 assign I1024 = ( wire7597*  &  wire7526* ) ;
 assign I1025 = ( wire7598*  &  wire7518* ) ;
 assign wire7968 = ( key<81>* ) ;
 assign wire1657 = ( wire7968*  &  wire7581* ) ;
 assign wire7967 = ( I1030 ) | ( I1029 ) ;
 assign I1029 = ( wire7602*  &  wire7532* ) ;
 assign I1030 = ( wire7963*  &  wire7604* ) ;
 assign new_C<41> = ( wire7967 ) | ( wire1657 ) | ( wire7965 ) | ( wire1654 ) ;
 assign wire1648 = ( wire7600*  &  wire7532* ) ;
 assign wire7538 = ( C<38>* ) ;
 assign wire7970 = ( I1036 ) | ( I1035 ) ;
 assign I1035 = ( wire7597*  &  wire7538* ) ;
 assign I1036 = ( wire7598*  &  wire7526* ) ;
 assign wire7973 = ( key<89>* ) ;
 assign wire1651 = ( wire7973*  &  wire7581* ) ;
 assign wire7972 = ( I1041 ) | ( I1040 ) ;
 assign I1040 = ( wire7602*  &  wire7540* ) ;
 assign I1041 = ( wire7968*  &  wire7604* ) ;
 assign new_C<40> = ( wire7972 ) | ( wire1651 ) | ( wire7970 ) | ( wire1648 ) ;
 assign wire1642 = ( wire7600*  &  wire7540* ) ;
 assign wire7529 = ( C<37>* ) ;
 assign wire7975 = ( I1047 ) | ( I1046 ) ;
 assign I1046 = ( wire7597*  &  wire7529* ) ;
 assign I1047 = ( wire7598*  &  wire7538* ) ;
 assign wire7978 = ( key<97>* ) ;
 assign wire1645 = ( wire7978*  &  wire7581* ) ;
 assign wire7977 = ( I1052 ) | ( I1051 ) ;
 assign I1051 = ( wire7602*  &  wire7518* ) ;
 assign I1052 = ( wire7973*  &  wire7604* ) ;
 assign new_C<39> = ( wire7977 ) | ( wire1645 ) | ( wire7975 ) | ( wire1642 ) ;
 assign wire1636 = ( wire7600*  &  wire7518* ) ;
 assign wire7980 = ( C<36>* ) ;
 assign wire7981 = ( I1058 ) | ( I1057 ) ;
 assign I1057 = ( wire7980*  &  wire7597* ) ;
 assign I1058 = ( wire7598*  &  wire7529* ) ;
 assign wire7984 = ( key<105>* ) ;
 assign wire1639 = ( wire7984*  &  wire7581* ) ;
 assign wire7983 = ( I1063 ) | ( I1062 ) ;
 assign I1062 = ( wire7602*  &  wire7526* ) ;
 assign I1063 = ( wire7978*  &  wire7604* ) ;
 assign new_C<38> = ( wire7983 ) | ( wire1639 ) | ( wire7981 ) | ( wire1636 ) ;
 assign wire1630 = ( wire7600*  &  wire7526* ) ;
 assign wire7523 = ( C<35>* ) ;
 assign wire7986 = ( I1069 ) | ( I1068 ) ;
 assign I1068 = ( wire7597*  &  wire7523* ) ;
 assign I1069 = ( wire7980*  &  wire7598* ) ;
 assign wire7989 = ( key<113>* ) ;
 assign wire1633 = ( wire7989*  &  wire7581* ) ;
 assign wire7988 = ( I1074 ) | ( I1073 ) ;
 assign I1073 = ( wire7602*  &  wire7538* ) ;
 assign I1074 = ( wire7984*  &  wire7604* ) ;
 assign new_C<37> = ( wire7988 ) | ( wire1633 ) | ( wire7986 ) | ( wire1630 ) ;
 assign wire1624 = ( wire7600*  &  wire7538* ) ;
 assign wire7521 = ( C<34>* ) ;
 assign wire7991 = ( I1080 ) | ( I1079 ) ;
 assign I1079 = ( wire7597*  &  wire7521* ) ;
 assign I1080 = ( wire7598*  &  wire7523* ) ;
 assign wire7994 = ( key<121>* ) ;
 assign wire1627 = ( wire7994*  &  wire7581* ) ;
 assign wire7993 = ( I1085 ) | ( I1084 ) ;
 assign I1084 = ( wire7602*  &  wire7529* ) ;
 assign I1085 = ( wire7989*  &  wire7604* ) ;
 assign new_C<36> = ( wire7993 ) | ( wire1627 ) | ( wire7991 ) | ( wire1624 ) ;
 assign wire1618 = ( wire7600*  &  wire7529* ) ;
 assign wire7531 = ( C<33>* ) ;
 assign wire7996 = ( I1091 ) | ( I1090 ) ;
 assign I1090 = ( wire7597*  &  wire7531* ) ;
 assign I1091 = ( wire7598*  &  wire7521* ) ;
 assign wire7999 = ( key<64>* ) ;
 assign wire1621 = ( wire7999*  &  wire7581* ) ;
 assign wire7998 = ( I1096 ) | ( I1095 ) ;
 assign I1095 = ( wire7980*  &  wire7602* ) ;
 assign I1096 = ( wire7994*  &  wire7604* ) ;
 assign new_C<35> = ( wire7998 ) | ( wire1621 ) | ( wire7996 ) | ( wire1618 ) ;
 assign wire1612 = ( wire7980*  &  wire7600* ) ;
 assign wire7535 = ( C<32>* ) ;
 assign wire8001 = ( I1102 ) | ( I1101 ) ;
 assign I1101 = ( wire7597*  &  wire7535* ) ;
 assign I1102 = ( wire7598*  &  wire7531* ) ;
 assign wire8004 = ( key<72>* ) ;
 assign wire1615 = ( wire8004*  &  wire7581* ) ;
 assign wire8003 = ( I1107 ) | ( I1106 ) ;
 assign I1106 = ( wire7602*  &  wire7523* ) ;
 assign I1107 = ( wire7999*  &  wire7604* ) ;
 assign new_C<34> = ( wire8003 ) | ( wire1615 ) | ( wire8001 ) | ( wire1612 ) ;
 assign wire1606 = ( wire7600*  &  wire7523* ) ;
 assign wire7525 = ( C<31>* ) ;
 assign wire8006 = ( I1113 ) | ( I1112 ) ;
 assign I1112 = ( wire7597*  &  wire7525* ) ;
 assign I1113 = ( wire7598*  &  wire7535* ) ;
 assign wire8009 = ( key<80>* ) ;
 assign wire1609 = ( wire8009*  &  wire7581* ) ;
 assign wire8008 = ( I1118 ) | ( I1117 ) ;
 assign I1117 = ( wire7602*  &  wire7521* ) ;
 assign I1118 = ( wire8004*  &  wire7604* ) ;
 assign new_C<33> = ( wire8008 ) | ( wire1609 ) | ( wire8006 ) | ( wire1606 ) ;
 assign wire1600 = ( wire7600*  &  wire7521* ) ;
 assign wire7534 = ( C<30>* ) ;
 assign wire8011 = ( I1124 ) | ( I1123 ) ;
 assign I1123 = ( wire7597*  &  wire7534* ) ;
 assign I1124 = ( wire7598*  &  wire7525* ) ;
 assign wire8014 = ( key<88>* ) ;
 assign wire1603 = ( wire8014*  &  wire7581* ) ;
 assign wire8013 = ( I1129 ) | ( I1128 ) ;
 assign I1128 = ( wire7602*  &  wire7531* ) ;
 assign I1129 = ( wire8009*  &  wire7604* ) ;
 assign new_C<32> = ( wire8013 ) | ( wire1603 ) | ( wire8011 ) | ( wire1600 ) ;
 assign wire1594 = ( wire7600*  &  wire7531* ) ;
 assign wire7517 = ( C<29>* ) ;
 assign wire8016 = ( I1135 ) | ( I1134 ) ;
 assign I1134 = ( wire7597*  &  wire7517* ) ;
 assign I1135 = ( wire7598*  &  wire7534* ) ;
 assign wire8019 = ( key<96>* ) ;
 assign wire1597 = ( wire8019*  &  wire7581* ) ;
 assign wire8018 = ( I1140 ) | ( I1139 ) ;
 assign I1139 = ( wire7602*  &  wire7535* ) ;
 assign I1140 = ( wire8014*  &  wire7604* ) ;
 assign new_C<31> = ( wire8018 ) | ( wire1597 ) | ( wire8016 ) | ( wire1594 ) ;
 assign wire1588 = ( wire7600*  &  wire7535* ) ;
 assign wire7536 = ( C<28>* ) ;
 assign wire8021 = ( I1146 ) | ( I1145 ) ;
 assign I1145 = ( wire7597*  &  wire7536* ) ;
 assign I1146 = ( wire7598*  &  wire7517* ) ;
 assign wire8024 = ( key<104>* ) ;
 assign wire1591 = ( wire8024*  &  wire7581* ) ;
 assign wire8023 = ( I1151 ) | ( I1150 ) ;
 assign I1150 = ( wire7602*  &  wire7525* ) ;
 assign I1151 = ( wire8019*  &  wire7604* ) ;
 assign new_C<30> = ( wire8023 ) | ( wire1591 ) | ( wire8021 ) | ( wire1588 ) ;
 assign wire1582 = ( wire7600*  &  wire7525* ) ;
 assign wire7557 = ( C<27>* ) ;
 assign wire8026 = ( I1157 ) | ( I1156 ) ;
 assign I1156 = ( wire7597*  &  wire7557* ) ;
 assign I1157 = ( wire7598*  &  wire7536* ) ;
 assign wire8029 = ( key<112>* ) ;
 assign wire1585 = ( wire8029*  &  wire7581* ) ;
 assign wire8028 = ( I1162 ) | ( I1161 ) ;
 assign I1161 = ( wire7602*  &  wire7534* ) ;
 assign I1162 = ( wire8024*  &  wire7604* ) ;
 assign new_C<29> = ( wire8028 ) | ( wire1585 ) | ( wire8026 ) | ( wire1582 ) ;
 assign wire1576 = ( wire7600*  &  wire7534* ) ;
 assign wire7544 = ( C<26>* ) ;
 assign wire8031 = ( I1168 ) | ( I1167 ) ;
 assign I1167 = ( wire7597*  &  wire7544* ) ;
 assign I1168 = ( wire7598*  &  wire7557* ) ;
 assign wire8034 = ( key<120>* ) ;
 assign wire1579 = ( wire8034*  &  wire7581* ) ;
 assign wire8033 = ( I1173 ) | ( I1172 ) ;
 assign I1172 = ( wire7602*  &  wire7517* ) ;
 assign I1173 = ( wire8029*  &  wire7604* ) ;
 assign new_C<28> = ( wire8033 ) | ( wire1579 ) | ( wire8031 ) | ( wire1576 ) ;
 assign wire1570 = ( wire7600*  &  wire7517* ) ;
 assign wire7548 = ( C<25>* ) ;
 assign wire8036 = ( I1179 ) | ( I1178 ) ;
 assign I1178 = ( wire7597*  &  wire7548* ) ;
 assign I1179 = ( wire7598*  &  wire7544* ) ;
 assign wire8039 = ( key<35>* ) ;
 assign wire1573 = ( wire8039*  &  wire7581* ) ;
 assign wire8038 = ( I1184 ) | ( I1183 ) ;
 assign I1183 = ( wire7602*  &  wire7536* ) ;
 assign I1184 = ( wire8034*  &  wire7604* ) ;
 assign new_C<27> = ( wire8038 ) | ( wire1573 ) | ( wire8036 ) | ( wire1570 ) ;
 assign wire1564 = ( wire7600*  &  wire7536* ) ;
 assign wire8041 = ( C<24>* ) ;
 assign wire8042 = ( I1190 ) | ( I1189 ) ;
 assign I1189 = ( wire8041*  &  wire7597* ) ;
 assign I1190 = ( wire7598*  &  wire7548* ) ;
 assign wire8045 = ( key<43>* ) ;
 assign wire1567 = ( wire8045*  &  wire7581* ) ;
 assign wire8044 = ( I1195 ) | ( I1194 ) ;
 assign I1194 = ( wire7602*  &  wire7557* ) ;
 assign I1195 = ( wire8039*  &  wire7604* ) ;
 assign new_C<26> = ( wire8044 ) | ( wire1567 ) | ( wire8042 ) | ( wire1564 ) ;
 assign wire1558 = ( wire7600*  &  wire7557* ) ;
 assign wire7561 = ( C<23>* ) ;
 assign wire8047 = ( I1201 ) | ( I1200 ) ;
 assign I1200 = ( wire7597*  &  wire7561* ) ;
 assign I1201 = ( wire8041*  &  wire7598* ) ;
 assign wire8050 = ( key<51>* ) ;
 assign wire1561 = ( wire8050*  &  wire7581* ) ;
 assign wire8049 = ( I1206 ) | ( I1205 ) ;
 assign I1205 = ( wire7602*  &  wire7544* ) ;
 assign I1206 = ( wire8045*  &  wire7604* ) ;
 assign new_C<25> = ( wire8049 ) | ( wire1561 ) | ( wire8047 ) | ( wire1558 ) ;
 assign wire1552 = ( wire7600*  &  wire7544* ) ;
 assign wire7552 = ( C<22>* ) ;
 assign wire8052 = ( I1212 ) | ( I1211 ) ;
 assign I1211 = ( wire7597*  &  wire7552* ) ;
 assign I1212 = ( wire7598*  &  wire7561* ) ;
 assign wire8055 = ( key<59>* ) ;
 assign wire1555 = ( wire8055*  &  wire7581* ) ;
 assign wire8054 = ( I1217 ) | ( I1216 ) ;
 assign I1216 = ( wire7602*  &  wire7548* ) ;
 assign I1217 = ( wire8050*  &  wire7604* ) ;
 assign new_C<24> = ( wire8054 ) | ( wire1555 ) | ( wire8052 ) | ( wire1552 ) ;
 assign wire1546 = ( wire7600*  &  wire7548* ) ;
 assign wire8057 = ( C<21>* ) ;
 assign wire8058 = ( I1223 ) | ( I1222 ) ;
 assign I1222 = ( wire8057*  &  wire7597* ) ;
 assign I1223 = ( wire7598*  &  wire7552* ) ;
 assign wire8061 = ( key<2>* ) ;
 assign wire1549 = ( wire8061*  &  wire7581* ) ;
 assign wire8060 = ( I1228 ) | ( I1227 ) ;
 assign I1227 = ( wire8041*  &  wire7602* ) ;
 assign I1228 = ( wire8055*  &  wire7604* ) ;
 assign new_C<23> = ( wire8060 ) | ( wire1549 ) | ( wire8058 ) | ( wire1546 ) ;
 assign wire1540 = ( wire8041*  &  wire7600* ) ;
 assign wire7554 = ( C<20>* ) ;
 assign wire8063 = ( I1234 ) | ( I1233 ) ;
 assign I1233 = ( wire7597*  &  wire7554* ) ;
 assign I1234 = ( wire8057*  &  wire7598* ) ;
 assign wire8066 = ( key<10>* ) ;
 assign wire1543 = ( wire8066*  &  wire7581* ) ;
 assign wire8065 = ( I1239 ) | ( I1238 ) ;
 assign I1238 = ( wire7602*  &  wire7561* ) ;
 assign I1239 = ( wire8061*  &  wire7604* ) ;
 assign new_C<22> = ( wire8065 ) | ( wire1543 ) | ( wire8063 ) | ( wire1540 ) ;
 assign wire1534 = ( wire7600*  &  wire7561* ) ;
 assign wire7543 = ( C<19>* ) ;
 assign wire8068 = ( I1245 ) | ( I1244 ) ;
 assign I1244 = ( wire7597*  &  wire7543* ) ;
 assign I1245 = ( wire7598*  &  wire7554* ) ;
 assign wire8071 = ( key<18>* ) ;
 assign wire1537 = ( wire8071*  &  wire7581* ) ;
 assign wire8070 = ( I1250 ) | ( I1249 ) ;
 assign I1249 = ( wire7602*  &  wire7552* ) ;
 assign I1250 = ( wire8066*  &  wire7604* ) ;
 assign new_C<21> = ( wire8070 ) | ( wire1537 ) | ( wire8068 ) | ( wire1534 ) ;
 assign wire1528 = ( wire7600*  &  wire7552* ) ;
 assign wire7551 = ( C<18>* ) ;
 assign wire8073 = ( I1256 ) | ( I1255 ) ;
 assign I1255 = ( wire7597*  &  wire7551* ) ;
 assign I1256 = ( wire7598*  &  wire7543* ) ;
 assign wire8076 = ( key<26>* ) ;
 assign wire1531 = ( wire8076*  &  wire7581* ) ;
 assign wire8075 = ( I1261 ) | ( I1260 ) ;
 assign I1260 = ( wire8057*  &  wire7602* ) ;
 assign I1261 = ( wire8071*  &  wire7604* ) ;
 assign new_C<20> = ( wire8075 ) | ( wire1531 ) | ( wire8073 ) | ( wire1528 ) ;
 assign wire1522 = ( wire8057*  &  wire7600* ) ;
 assign wire8078 = ( C<17>* ) ;
 assign wire8079 = ( I1267 ) | ( I1266 ) ;
 assign I1266 = ( wire8078*  &  wire7597* ) ;
 assign I1267 = ( wire7598*  &  wire7551* ) ;
 assign wire8082 = ( key<34>* ) ;
 assign wire1525 = ( wire8082*  &  wire7581* ) ;
 assign wire8081 = ( I1272 ) | ( I1271 ) ;
 assign I1271 = ( wire7602*  &  wire7554* ) ;
 assign I1272 = ( wire8076*  &  wire7604* ) ;
 assign new_C<19> = ( wire8081 ) | ( wire1525 ) | ( wire8079 ) | ( wire1522 ) ;
 assign wire1516 = ( wire7600*  &  wire7554* ) ;
 assign wire7563 = ( C<16>* ) ;
 assign wire8084 = ( I1278 ) | ( I1277 ) ;
 assign I1277 = ( wire7597*  &  wire7563* ) ;
 assign I1278 = ( wire8078*  &  wire7598* ) ;
 assign wire8087 = ( key<42>* ) ;
 assign wire1519 = ( wire8087*  &  wire7581* ) ;
 assign wire8086 = ( I1283 ) | ( I1282 ) ;
 assign I1282 = ( wire7602*  &  wire7543* ) ;
 assign I1283 = ( wire8082*  &  wire7604* ) ;
 assign new_C<18> = ( wire8086 ) | ( wire1519 ) | ( wire8084 ) | ( wire1516 ) ;
 assign wire1510 = ( wire7600*  &  wire7543* ) ;
 assign wire7546 = ( C<15>* ) ;
 assign wire8089 = ( I1289 ) | ( I1288 ) ;
 assign I1288 = ( wire7597*  &  wire7546* ) ;
 assign I1289 = ( wire7598*  &  wire7563* ) ;
 assign wire8092 = ( key<50>* ) ;
 assign wire1513 = ( wire8092*  &  wire7581* ) ;
 assign wire8091 = ( I1294 ) | ( I1293 ) ;
 assign I1293 = ( wire7602*  &  wire7551* ) ;
 assign I1294 = ( wire8087*  &  wire7604* ) ;
 assign new_C<17> = ( wire8091 ) | ( wire1513 ) | ( wire8089 ) | ( wire1510 ) ;
 assign wire1504 = ( wire7600*  &  wire7551* ) ;
 assign wire7556 = ( C<14>* ) ;
 assign wire8094 = ( I1300 ) | ( I1299 ) ;
 assign I1299 = ( wire7597*  &  wire7556* ) ;
 assign I1300 = ( wire7598*  &  wire7546* ) ;
 assign wire8097 = ( key<58>* ) ;
 assign wire1507 = ( wire8097*  &  wire7581* ) ;
 assign wire8096 = ( I1305 ) | ( I1304 ) ;
 assign I1304 = ( wire8078*  &  wire7602* ) ;
 assign I1305 = ( wire8092*  &  wire7604* ) ;
 assign new_C<16> = ( wire8096 ) | ( wire1507 ) | ( wire8094 ) | ( wire1504 ) ;
 assign wire1498 = ( wire8078*  &  wire7600* ) ;
 assign wire7564 = ( C<13>* ) ;
 assign wire8099 = ( I1311 ) | ( I1310 ) ;
 assign I1310 = ( wire7597*  &  wire7564* ) ;
 assign I1311 = ( wire7598*  &  wire7556* ) ;
 assign wire8102 = ( key<1>* ) ;
 assign wire1501 = ( wire8102*  &  wire7581* ) ;
 assign wire8101 = ( I1316 ) | ( I1315 ) ;
 assign I1315 = ( wire7602*  &  wire7563* ) ;
 assign I1316 = ( wire8097*  &  wire7604* ) ;
 assign new_C<15> = ( wire8101 ) | ( wire1501 ) | ( wire8099 ) | ( wire1498 ) ;
 assign wire1492 = ( wire7600*  &  wire7563* ) ;
 assign wire7542 = ( C<12>* ) ;
 assign wire8104 = ( I1322 ) | ( I1321 ) ;
 assign I1321 = ( wire7597*  &  wire7542* ) ;
 assign I1322 = ( wire7598*  &  wire7564* ) ;
 assign wire8107 = ( key<9>* ) ;
 assign wire1495 = ( wire8107*  &  wire7581* ) ;
 assign wire8106 = ( I1327 ) | ( I1326 ) ;
 assign I1326 = ( wire7602*  &  wire7546* ) ;
 assign I1327 = ( wire8102*  &  wire7604* ) ;
 assign new_C<14> = ( wire8106 ) | ( wire1495 ) | ( wire8104 ) | ( wire1492 ) ;
 assign wire1486 = ( wire7600*  &  wire7546* ) ;
 assign wire7550 = ( C<11>* ) ;
 assign wire8109 = ( I1333 ) | ( I1332 ) ;
 assign I1332 = ( wire7597*  &  wire7550* ) ;
 assign I1333 = ( wire7598*  &  wire7542* ) ;
 assign wire8112 = ( key<17>* ) ;
 assign wire1489 = ( wire8112*  &  wire7581* ) ;
 assign wire8111 = ( I1338 ) | ( I1337 ) ;
 assign I1337 = ( wire7602*  &  wire7556* ) ;
 assign I1338 = ( wire8107*  &  wire7604* ) ;
 assign new_C<13> = ( wire8111 ) | ( wire1489 ) | ( wire8109 ) | ( wire1486 ) ;
 assign wire1480 = ( wire7600*  &  wire7556* ) ;
 assign wire7562 = ( C<10>* ) ;
 assign wire8114 = ( I1344 ) | ( I1343 ) ;
 assign I1343 = ( wire7597*  &  wire7562* ) ;
 assign I1344 = ( wire7598*  &  wire7550* ) ;
 assign wire8117 = ( key<25>* ) ;
 assign wire1483 = ( wire8117*  &  wire7581* ) ;
 assign wire8116 = ( I1349 ) | ( I1348 ) ;
 assign I1348 = ( wire7602*  &  wire7564* ) ;
 assign I1349 = ( wire8112*  &  wire7604* ) ;
 assign new_C<12> = ( wire8116 ) | ( wire1483 ) | ( wire8114 ) | ( wire1480 ) ;
 assign wire1474 = ( wire7600*  &  wire7564* ) ;
 assign wire7553 = ( C<9>* ) ;
 assign wire8119 = ( I1355 ) | ( I1354 ) ;
 assign I1354 = ( wire7597*  &  wire7553* ) ;
 assign I1355 = ( wire7598*  &  wire7562* ) ;
 assign wire8122 = ( key<33>* ) ;
 assign wire1477 = ( wire8122*  &  wire7581* ) ;
 assign wire8121 = ( I1360 ) | ( I1359 ) ;
 assign I1359 = ( wire7602*  &  wire7542* ) ;
 assign I1360 = ( wire8117*  &  wire7604* ) ;
 assign new_C<11> = ( wire8121 ) | ( wire1477 ) | ( wire8119 ) | ( wire1474 ) ;
 assign wire1468 = ( wire7600*  &  wire7542* ) ;
 assign wire8124 = ( C<8>* ) ;
 assign wire8125 = ( I1366 ) | ( I1365 ) ;
 assign I1365 = ( wire8124*  &  wire7597* ) ;
 assign I1366 = ( wire7598*  &  wire7553* ) ;
 assign wire8128 = ( key<41>* ) ;
 assign wire1471 = ( wire8128*  &  wire7581* ) ;
 assign wire8127 = ( I1371 ) | ( I1370 ) ;
 assign I1370 = ( wire7602*  &  wire7550* ) ;
 assign I1371 = ( wire8122*  &  wire7604* ) ;
 assign new_C<10> = ( wire8127 ) | ( wire1471 ) | ( wire8125 ) | ( wire1468 ) ;
 assign wire1462 = ( wire7600*  &  wire7550* ) ;
 assign wire7547 = ( C<7>* ) ;
 assign wire8130 = ( I1377 ) | ( I1376 ) ;
 assign I1376 = ( wire7597*  &  wire7547* ) ;
 assign I1377 = ( wire8124*  &  wire7598* ) ;
 assign wire8133 = ( key<49>* ) ;
 assign wire1465 = ( wire8133*  &  wire7581* ) ;
 assign wire8132 = ( I1382 ) | ( I1381 ) ;
 assign I1381 = ( wire7602*  &  wire7562* ) ;
 assign I1382 = ( wire8128*  &  wire7604* ) ;
 assign new_C<9> = ( wire8132 ) | ( wire1465 ) | ( wire8130 ) | ( wire1462 ) ;
 assign wire1456 = ( wire7600*  &  wire7562* ) ;
 assign wire7545 = ( C<6>* ) ;
 assign wire8135 = ( I1388 ) | ( I1387 ) ;
 assign I1387 = ( wire7597*  &  wire7545* ) ;
 assign I1388 = ( wire7598*  &  wire7547* ) ;
 assign wire8138 = ( key<57>* ) ;
 assign wire1459 = ( wire8138*  &  wire7581* ) ;
 assign wire8137 = ( I1393 ) | ( I1392 ) ;
 assign I1392 = ( wire7602*  &  wire7553* ) ;
 assign I1393 = ( wire8133*  &  wire7604* ) ;
 assign new_C<8> = ( wire8137 ) | ( wire1459 ) | ( wire8135 ) | ( wire1456 ) ;
 assign wire1450 = ( wire7600*  &  wire7553* ) ;
 assign wire7555 = ( C<5>* ) ;
 assign wire8140 = ( I1399 ) | ( I1398 ) ;
 assign I1398 = ( wire7597*  &  wire7555* ) ;
 assign I1399 = ( wire7598*  &  wire7545* ) ;
 assign wire8143 = ( key<0>* ) ;
 assign wire1453 = ( wire8143*  &  wire7581* ) ;
 assign wire8142 = ( I1404 ) | ( I1403 ) ;
 assign I1403 = ( wire8124*  &  wire7602* ) ;
 assign I1404 = ( wire8138*  &  wire7604* ) ;
 assign new_C<7> = ( wire8142 ) | ( wire1453 ) | ( wire8140 ) | ( wire1450 ) ;
 assign wire1444 = ( wire8124*  &  wire7600* ) ;
 assign wire7559 = ( C<4>* ) ;
 assign wire8145 = ( I1410 ) | ( I1409 ) ;
 assign I1409 = ( wire7597*  &  wire7559* ) ;
 assign I1410 = ( wire7598*  &  wire7555* ) ;
 assign wire8148 = ( key<8>* ) ;
 assign wire1447 = ( wire8148*  &  wire7581* ) ;
 assign wire8147 = ( I1415 ) | ( I1414 ) ;
 assign I1414 = ( wire7602*  &  wire7547* ) ;
 assign I1415 = ( wire8143*  &  wire7604* ) ;
 assign new_C<6> = ( wire8147 ) | ( wire1447 ) | ( wire8145 ) | ( wire1444 ) ;
 assign wire1438 = ( wire7600*  &  wire7547* ) ;
 assign wire7549 = ( C<3>* ) ;
 assign wire8150 = ( I1421 ) | ( I1420 ) ;
 assign I1420 = ( wire7597*  &  wire7549* ) ;
 assign I1421 = ( wire7598*  &  wire7559* ) ;
 assign wire8153 = ( key<16>* ) ;
 assign wire1441 = ( wire8153*  &  wire7581* ) ;
 assign wire8152 = ( I1426 ) | ( I1425 ) ;
 assign I1425 = ( wire7602*  &  wire7545* ) ;
 assign I1426 = ( wire8148*  &  wire7604* ) ;
 assign new_C<5> = ( wire8152 ) | ( wire1441 ) | ( wire8150 ) | ( wire1438 ) ;
 assign wire1432 = ( wire7600*  &  wire7545* ) ;
 assign wire7558 = ( C<2>* ) ;
 assign wire8155 = ( I1432 ) | ( I1431 ) ;
 assign I1431 = ( wire7597*  &  wire7558* ) ;
 assign I1432 = ( wire7598*  &  wire7549* ) ;
 assign wire8158 = ( key<24>* ) ;
 assign wire1435 = ( wire8158*  &  wire7581* ) ;
 assign wire8157 = ( I1437 ) | ( I1436 ) ;
 assign I1436 = ( wire7602*  &  wire7555* ) ;
 assign I1437 = ( wire8153*  &  wire7604* ) ;
 assign new_C<4> = ( wire8157 ) | ( wire1435 ) | ( wire8155 ) | ( wire1432 ) ;
 assign wire1426 = ( wire7600*  &  wire7555* ) ;
 assign wire8160 = ( I1442 ) | ( I1441 ) ;
 assign I1441 = ( wire7597*  &  wire7541* ) ;
 assign I1442 = ( wire7598*  &  wire7558* ) ;
 assign wire8163 = ( key<32>* ) ;
 assign wire1429 = ( wire8163*  &  wire7581* ) ;
 assign wire8162 = ( I1447 ) | ( I1446 ) ;
 assign I1446 = ( wire7602*  &  wire7559* ) ;
 assign I1447 = ( wire8158*  &  wire7604* ) ;
 assign new_C<3> = ( wire8162 ) | ( wire1429 ) | ( wire8160 ) | ( wire1426 ) ;
 assign wire1420 = ( wire7600*  &  wire7559* ) ;
 assign wire8165 = ( I1452 ) | ( I1451 ) ;
 assign I1451 = ( wire7597*  &  wire7560* ) ;
 assign I1452 = ( wire7598*  &  wire7541* ) ;
 assign wire8168 = ( key<40>* ) ;
 assign wire1423 = ( wire8168*  &  wire7581* ) ;
 assign wire8167 = ( I1457 ) | ( I1456 ) ;
 assign I1456 = ( wire7602*  &  wire7549* ) ;
 assign I1457 = ( wire8163*  &  wire7604* ) ;
 assign new_C<2> = ( wire8167 ) | ( wire1423 ) | ( wire8165 ) | ( wire1420 ) ;
 assign wire1414 = ( wire7600*  &  wire7549* ) ;
 assign wire8170 = ( I1462 ) | ( I1461 ) ;
 assign I1461 = ( wire7597*  &  wire7485* ) ;
 assign I1462 = ( wire7598*  &  wire7560* ) ;
 assign wire8173 = ( key<48>* ) ;
 assign wire1417 = ( wire8173*  &  wire7581* ) ;
 assign wire8172 = ( I1467 ) | ( I1466 ) ;
 assign I1466 = ( wire7602*  &  wire7558* ) ;
 assign I1467 = ( wire8168*  &  wire7604* ) ;
 assign new_C<1> = ( wire8172 ) | ( wire1417 ) | ( wire8170 ) | ( wire1414 ) ;
 assign wire1408 = ( wire7600*  &  wire7558* ) ;
 assign wire8175 = ( I1472 ) | ( I1471 ) ;
 assign I1471 = ( wire7597*  &  wire7473* ) ;
 assign I1472 = ( wire7598*  &  wire7485* ) ;
 assign wire1411 = ( wire7603*  &  wire7581* ) ;
 assign wire8177 = ( I1476 ) | ( I1475 ) ;
 assign I1475 = ( wire7602*  &  wire7541* ) ;
 assign I1476 = ( wire8173*  &  wire7604* ) ;
 assign new_C<0> = ( wire8177 ) | ( wire1411 ) | ( wire8175 ) | ( wire1408 ) ;
 assign wire7463 = ( D<1>* ) ;
 assign wire1402 = ( wire7600*  &  wire7463* ) ;
 assign wire8179 = ( D<109>* ) ;
 assign wire7394 = ( D<110>* ) ;
 assign wire8180 = ( I1484 ) | ( I1483 ) ;
 assign I1483 = ( wire8179*  &  wire7597* ) ;
 assign I1484 = ( wire7598*  &  wire7394* ) ;
 assign wire8184 = ( key<195>* ) ;
 assign wire1405 = ( wire8184*  &  wire7581* ) ;
 assign wire7447 = ( D<0>* ) ;
 assign wire8182 = ( key<62>* ) ;
 assign wire8183 = ( I1491 ) | ( I1490 ) ;
 assign I1490 = ( wire7602*  &  wire7447* ) ;
 assign I1491 = ( wire8182*  &  wire7604* ) ;
 assign new_D<111> = ( wire8183 ) | ( wire1405 ) | ( wire8180 ) | ( wire1402 ) ;
 assign wire1396 = ( wire7600*  &  wire7447* ) ;
 assign wire7382 = ( D<108>* ) ;
 assign wire8186 = ( I1497 ) | ( I1496 ) ;
 assign I1496 = ( wire7597*  &  wire7382* ) ;
 assign I1497 = ( wire8179*  &  wire7598* ) ;
 assign wire8189 = ( key<203>* ) ;
 assign wire1399 = ( wire8189*  &  wire7581* ) ;
 assign wire7384 = ( D<111>* ) ;
 assign wire8188 = ( I1503 ) | ( I1502 ) ;
 assign I1502 = ( wire7602*  &  wire7384* ) ;
 assign I1503 = ( wire8184*  &  wire7604* ) ;
 assign new_D<110> = ( wire8188 ) | ( wire1399 ) | ( wire8186 ) | ( wire1396 ) ;
 assign wire1390 = ( wire7600*  &  wire7384* ) ;
 assign wire7398 = ( D<107>* ) ;
 assign wire8191 = ( I1509 ) | ( I1508 ) ;
 assign I1508 = ( wire7597*  &  wire7398* ) ;
 assign I1509 = ( wire7598*  &  wire7382* ) ;
 assign wire8194 = ( key<211>* ) ;
 assign wire1393 = ( wire8194*  &  wire7581* ) ;
 assign wire8193 = ( I1514 ) | ( I1513 ) ;
 assign I1513 = ( wire7602*  &  wire7394* ) ;
 assign I1514 = ( wire8189*  &  wire7604* ) ;
 assign new_D<109> = ( wire8193 ) | ( wire1393 ) | ( wire8191 ) | ( wire1390 ) ;
 assign wire1384 = ( wire7600*  &  wire7394* ) ;
 assign wire7391 = ( D<106>* ) ;
 assign wire8196 = ( I1520 ) | ( I1519 ) ;
 assign I1519 = ( wire7597*  &  wire7391* ) ;
 assign I1520 = ( wire7598*  &  wire7398* ) ;
 assign wire8199 = ( key<219>* ) ;
 assign wire1387 = ( wire8199*  &  wire7581* ) ;
 assign wire8198 = ( I1525 ) | ( I1524 ) ;
 assign I1524 = ( wire8179*  &  wire7602* ) ;
 assign I1525 = ( wire8194*  &  wire7604* ) ;
 assign new_D<108> = ( wire8198 ) | ( wire1387 ) | ( wire8196 ) | ( wire1384 ) ;
 assign wire1378 = ( wire8179*  &  wire7600* ) ;
 assign wire7380 = ( D<105>* ) ;
 assign wire8201 = ( I1531 ) | ( I1530 ) ;
 assign I1530 = ( wire7597*  &  wire7380* ) ;
 assign I1531 = ( wire7598*  &  wire7391* ) ;
 assign wire8204 = ( key<196>* ) ;
 assign wire1381 = ( wire8204*  &  wire7581* ) ;
 assign wire8203 = ( I1536 ) | ( I1535 ) ;
 assign I1535 = ( wire7602*  &  wire7382* ) ;
 assign I1536 = ( wire8199*  &  wire7604* ) ;
 assign new_D<107> = ( wire8203 ) | ( wire1381 ) | ( wire8201 ) | ( wire1378 ) ;
 assign wire1372 = ( wire7600*  &  wire7382* ) ;
 assign wire7386 = ( D<104>* ) ;
 assign wire8206 = ( I1542 ) | ( I1541 ) ;
 assign I1541 = ( wire7597*  &  wire7386* ) ;
 assign I1542 = ( wire7598*  &  wire7380* ) ;
 assign wire8209 = ( key<204>* ) ;
 assign wire1375 = ( wire8209*  &  wire7581* ) ;
 assign wire8208 = ( I1547 ) | ( I1546 ) ;
 assign I1546 = ( wire7602*  &  wire7398* ) ;
 assign I1547 = ( wire8204*  &  wire7604* ) ;
 assign new_D<106> = ( wire8208 ) | ( wire1375 ) | ( wire8206 ) | ( wire1372 ) ;
 assign wire1366 = ( wire7600*  &  wire7398* ) ;
 assign wire7388 = ( D<103>* ) ;
 assign wire8211 = ( I1553 ) | ( I1552 ) ;
 assign I1552 = ( wire7597*  &  wire7388* ) ;
 assign I1553 = ( wire7598*  &  wire7386* ) ;
 assign wire8214 = ( key<212>* ) ;
 assign wire1369 = ( wire8214*  &  wire7581* ) ;
 assign wire8213 = ( I1558 ) | ( I1557 ) ;
 assign I1557 = ( wire7602*  &  wire7391* ) ;
 assign I1558 = ( wire8209*  &  wire7604* ) ;
 assign new_D<105> = ( wire8213 ) | ( wire1369 ) | ( wire8211 ) | ( wire1366 ) ;
 assign wire1360 = ( wire7600*  &  wire7391* ) ;
 assign wire7395 = ( D<102>* ) ;
 assign wire8216 = ( I1564 ) | ( I1563 ) ;
 assign I1563 = ( wire7597*  &  wire7395* ) ;
 assign I1564 = ( wire7598*  &  wire7388* ) ;
 assign wire8219 = ( key<220>* ) ;
 assign wire1363 = ( wire8219*  &  wire7581* ) ;
 assign wire8218 = ( I1569 ) | ( I1568 ) ;
 assign I1568 = ( wire7602*  &  wire7380* ) ;
 assign I1569 = ( wire8214*  &  wire7604* ) ;
 assign new_D<104> = ( wire8218 ) | ( wire1363 ) | ( wire8216 ) | ( wire1360 ) ;
 assign wire1354 = ( wire7600*  &  wire7380* ) ;
 assign wire7381 = ( D<101>* ) ;
 assign wire8221 = ( I1575 ) | ( I1574 ) ;
 assign I1574 = ( wire7597*  &  wire7381* ) ;
 assign I1575 = ( wire7598*  &  wire7395* ) ;
 assign wire8224 = ( key<228>* ) ;
 assign wire1357 = ( wire8224*  &  wire7581* ) ;
 assign wire8223 = ( I1580 ) | ( I1579 ) ;
 assign I1579 = ( wire7602*  &  wire7386* ) ;
 assign I1580 = ( wire8219*  &  wire7604* ) ;
 assign new_D<103> = ( wire8223 ) | ( wire1357 ) | ( wire8221 ) | ( wire1354 ) ;
 assign wire1348 = ( wire7600*  &  wire7386* ) ;
 assign wire7390 = ( D<100>* ) ;
 assign wire8226 = ( I1586 ) | ( I1585 ) ;
 assign I1585 = ( wire7597*  &  wire7390* ) ;
 assign I1586 = ( wire7598*  &  wire7381* ) ;
 assign wire8229 = ( key<172>* ) ;
 assign wire1351 = ( wire8229*  &  wire7581* ) ;
 assign wire8228 = ( I1591 ) | ( I1590 ) ;
 assign I1590 = ( wire7602*  &  wire7388* ) ;
 assign I1591 = ( wire8224*  &  wire7604* ) ;
 assign new_D<102> = ( wire8228 ) | ( wire1351 ) | ( wire8226 ) | ( wire1348 ) ;
 assign wire1342 = ( wire7600*  &  wire7388* ) ;
 assign wire7387 = ( D<99>* ) ;
 assign wire8231 = ( I1597 ) | ( I1596 ) ;
 assign I1596 = ( wire7597*  &  wire7387* ) ;
 assign I1597 = ( wire7598*  &  wire7390* ) ;
 assign wire8234 = ( key<244>* ) ;
 assign wire1345 = ( wire8234*  &  wire7581* ) ;
 assign wire8233 = ( I1602 ) | ( I1601 ) ;
 assign I1601 = ( wire7602*  &  wire7395* ) ;
 assign I1602 = ( wire8229*  &  wire7604* ) ;
 assign new_D<101> = ( wire8233 ) | ( wire1345 ) | ( wire8231 ) | ( wire1342 ) ;
 assign wire1336 = ( wire7600*  &  wire7395* ) ;
 assign wire8236 = ( D<98>* ) ;
 assign wire8237 = ( I1608 ) | ( I1607 ) ;
 assign I1607 = ( wire8236*  &  wire7597* ) ;
 assign I1608 = ( wire7598*  &  wire7387* ) ;
 assign wire8240 = ( key<252>* ) ;
 assign wire1339 = ( wire8240*  &  wire7581* ) ;
 assign wire8239 = ( I1613 ) | ( I1612 ) ;
 assign I1612 = ( wire7602*  &  wire7381* ) ;
 assign I1613 = ( wire8234*  &  wire7604* ) ;
 assign new_D<100> = ( wire8239 ) | ( wire1339 ) | ( wire8237 ) | ( wire1336 ) ;
 assign wire1330 = ( wire7600*  &  wire7381* ) ;
 assign wire8242 = ( D<97>* ) ;
 assign wire8243 = ( I1619 ) | ( I1618 ) ;
 assign I1618 = ( wire8242*  &  wire7597* ) ;
 assign I1619 = ( wire8236*  &  wire7598* ) ;
 assign wire8246 = ( key<197>* ) ;
 assign wire1333 = ( wire8246*  &  wire7581* ) ;
 assign wire8245 = ( I1624 ) | ( I1623 ) ;
 assign I1623 = ( wire7602*  &  wire7390* ) ;
 assign I1624 = ( wire8240*  &  wire7604* ) ;
 assign new_D<99> = ( wire8245 ) | ( wire1333 ) | ( wire8243 ) | ( wire1330 ) ;
 assign wire1324 = ( wire7600*  &  wire7390* ) ;
 assign wire8248 = ( D<96>* ) ;
 assign wire8249 = ( I1630 ) | ( I1629 ) ;
 assign I1629 = ( wire8248*  &  wire7597* ) ;
 assign I1630 = ( wire8242*  &  wire7598* ) ;
 assign wire8252 = ( key<205>* ) ;
 assign wire1327 = ( wire8252*  &  wire7581* ) ;
 assign wire8251 = ( I1635 ) | ( I1634 ) ;
 assign I1634 = ( wire7602*  &  wire7387* ) ;
 assign I1635 = ( wire8246*  &  wire7604* ) ;
 assign new_D<98> = ( wire8251 ) | ( wire1327 ) | ( wire8249 ) | ( wire1324 ) ;
 assign wire1318 = ( wire7600*  &  wire7387* ) ;
 assign wire7392 = ( D<95>* ) ;
 assign wire8254 = ( I1641 ) | ( I1640 ) ;
 assign I1640 = ( wire7597*  &  wire7392* ) ;
 assign I1641 = ( wire8248*  &  wire7598* ) ;
 assign wire8257 = ( key<213>* ) ;
 assign wire1321 = ( wire8257*  &  wire7581* ) ;
 assign wire8256 = ( I1646 ) | ( I1645 ) ;
 assign I1645 = ( wire8236*  &  wire7602* ) ;
 assign I1646 = ( wire8252*  &  wire7604* ) ;
 assign new_D<97> = ( wire8256 ) | ( wire1321 ) | ( wire8254 ) | ( wire1318 ) ;
 assign wire1312 = ( wire8236*  &  wire7600* ) ;
 assign wire7385 = ( D<94>* ) ;
 assign wire8259 = ( I1652 ) | ( I1651 ) ;
 assign I1651 = ( wire7597*  &  wire7385* ) ;
 assign I1652 = ( wire7598*  &  wire7392* ) ;
 assign wire8262 = ( key<221>* ) ;
 assign wire1315 = ( wire8262*  &  wire7581* ) ;
 assign wire8261 = ( I1657 ) | ( I1656 ) ;
 assign I1656 = ( wire8242*  &  wire7602* ) ;
 assign I1657 = ( wire8257*  &  wire7604* ) ;
 assign new_D<96> = ( wire8261 ) | ( wire1315 ) | ( wire8259 ) | ( wire1312 ) ;
 assign wire1306 = ( wire8242*  &  wire7600* ) ;
 assign wire8264 = ( D<93>* ) ;
 assign wire8265 = ( I1663 ) | ( I1662 ) ;
 assign I1662 = ( wire8264*  &  wire7597* ) ;
 assign I1663 = ( wire7598*  &  wire7385* ) ;
 assign wire8268 = ( key<229>* ) ;
 assign wire1309 = ( wire8268*  &  wire7581* ) ;
 assign wire8267 = ( I1668 ) | ( I1667 ) ;
 assign I1667 = ( wire8248*  &  wire7602* ) ;
 assign I1668 = ( wire8262*  &  wire7604* ) ;
 assign new_D<95> = ( wire8267 ) | ( wire1309 ) | ( wire8265 ) | ( wire1306 ) ;
 assign wire1300 = ( wire8248*  &  wire7600* ) ;
 assign wire7396 = ( D<92>* ) ;
 assign wire8270 = ( I1674 ) | ( I1673 ) ;
 assign I1673 = ( wire7597*  &  wire7396* ) ;
 assign I1674 = ( wire8264*  &  wire7598* ) ;
 assign wire8273 = ( key<237>* ) ;
 assign wire1303 = ( wire8273*  &  wire7581* ) ;
 assign wire8272 = ( I1679 ) | ( I1678 ) ;
 assign I1678 = ( wire7602*  &  wire7392* ) ;
 assign I1679 = ( wire8268*  &  wire7604* ) ;
 assign new_D<94> = ( wire8272 ) | ( wire1303 ) | ( wire8270 ) | ( wire1300 ) ;
 assign wire1294 = ( wire7600*  &  wire7392* ) ;
 assign wire7379 = ( D<91>* ) ;
 assign wire8275 = ( I1685 ) | ( I1684 ) ;
 assign I1684 = ( wire7597*  &  wire7379* ) ;
 assign I1685 = ( wire7598*  &  wire7396* ) ;
 assign wire8278 = ( key<245>* ) ;
 assign wire1297 = ( wire8278*  &  wire7581* ) ;
 assign wire8277 = ( I1690 ) | ( I1689 ) ;
 assign I1689 = ( wire7602*  &  wire7385* ) ;
 assign I1690 = ( wire8273*  &  wire7604* ) ;
 assign new_D<93> = ( wire8277 ) | ( wire1297 ) | ( wire8275 ) | ( wire1294 ) ;
 assign wire1288 = ( wire7600*  &  wire7385* ) ;
 assign wire8280 = ( D<90>* ) ;
 assign wire8281 = ( I1696 ) | ( I1695 ) ;
 assign I1695 = ( wire8280*  &  wire7597* ) ;
 assign I1696 = ( wire7598*  &  wire7379* ) ;
 assign wire8284 = ( key<253>* ) ;
 assign wire1291 = ( wire8284*  &  wire7581* ) ;
 assign wire8283 = ( I1701 ) | ( I1700 ) ;
 assign I1700 = ( wire8264*  &  wire7602* ) ;
 assign I1701 = ( wire8278*  &  wire7604* ) ;
 assign new_D<92> = ( wire8283 ) | ( wire1291 ) | ( wire8281 ) | ( wire1288 ) ;
 assign wire1282 = ( wire8264*  &  wire7600* ) ;
 assign wire7383 = ( D<89>* ) ;
 assign wire8286 = ( I1707 ) | ( I1706 ) ;
 assign I1706 = ( wire7597*  &  wire7383* ) ;
 assign I1707 = ( wire8280*  &  wire7598* ) ;
 assign wire8289 = ( key<198>* ) ;
 assign wire1285 = ( wire8289*  &  wire7581* ) ;
 assign wire8288 = ( I1712 ) | ( I1711 ) ;
 assign I1711 = ( wire7602*  &  wire7396* ) ;
 assign I1712 = ( wire8284*  &  wire7604* ) ;
 assign new_D<91> = ( wire8288 ) | ( wire1285 ) | ( wire8286 ) | ( wire1282 ) ;
 assign wire1276 = ( wire7600*  &  wire7396* ) ;
 assign wire7389 = ( D<88>* ) ;
 assign wire8291 = ( I1718 ) | ( I1717 ) ;
 assign I1717 = ( wire7597*  &  wire7389* ) ;
 assign I1718 = ( wire7598*  &  wire7383* ) ;
 assign wire8294 = ( key<206>* ) ;
 assign wire1279 = ( wire8294*  &  wire7581* ) ;
 assign wire8293 = ( I1723 ) | ( I1722 ) ;
 assign I1722 = ( wire7602*  &  wire7379* ) ;
 assign I1723 = ( wire8289*  &  wire7604* ) ;
 assign new_D<90> = ( wire8293 ) | ( wire1279 ) | ( wire8291 ) | ( wire1276 ) ;
 assign wire1270 = ( wire7600*  &  wire7379* ) ;
 assign wire7377 = ( D<87>* ) ;
 assign wire8296 = ( I1729 ) | ( I1728 ) ;
 assign I1728 = ( wire7597*  &  wire7377* ) ;
 assign I1729 = ( wire7598*  &  wire7389* ) ;
 assign wire8299 = ( key<214>* ) ;
 assign wire1273 = ( wire8299*  &  wire7581* ) ;
 assign wire8298 = ( I1734 ) | ( I1733 ) ;
 assign I1733 = ( wire8280*  &  wire7602* ) ;
 assign I1734 = ( wire8294*  &  wire7604* ) ;
 assign new_D<89> = ( wire8298 ) | ( wire1273 ) | ( wire8296 ) | ( wire1270 ) ;
 assign wire1264 = ( wire8280*  &  wire7600* ) ;
 assign wire7397 = ( D<86>* ) ;
 assign wire8301 = ( I1740 ) | ( I1739 ) ;
 assign I1739 = ( wire7597*  &  wire7397* ) ;
 assign I1740 = ( wire7598*  &  wire7377* ) ;
 assign wire8304 = ( key<222>* ) ;
 assign wire1267 = ( wire8304*  &  wire7581* ) ;
 assign wire8303 = ( I1745 ) | ( I1744 ) ;
 assign I1744 = ( wire7602*  &  wire7383* ) ;
 assign I1745 = ( wire8299*  &  wire7604* ) ;
 assign new_D<88> = ( wire8303 ) | ( wire1267 ) | ( wire8301 ) | ( wire1264 ) ;
 assign wire1258 = ( wire7600*  &  wire7383* ) ;
 assign wire7393 = ( D<85>* ) ;
 assign wire8306 = ( I1751 ) | ( I1750 ) ;
 assign I1750 = ( wire7597*  &  wire7393* ) ;
 assign I1751 = ( wire7598*  &  wire7397* ) ;
 assign wire8309 = ( key<230>* ) ;
 assign wire1261 = ( wire8309*  &  wire7581* ) ;
 assign wire8308 = ( I1756 ) | ( I1755 ) ;
 assign I1755 = ( wire7602*  &  wire7389* ) ;
 assign I1756 = ( wire8304*  &  wire7604* ) ;
 assign new_D<87> = ( wire8308 ) | ( wire1261 ) | ( wire8306 ) | ( wire1258 ) ;
 assign wire1252 = ( wire7600*  &  wire7389* ) ;
 assign wire7378 = ( D<84>* ) ;
 assign wire8311 = ( I1762 ) | ( I1761 ) ;
 assign I1761 = ( wire7597*  &  wire7378* ) ;
 assign I1762 = ( wire7598*  &  wire7393* ) ;
 assign wire8314 = ( key<238>* ) ;
 assign wire1255 = ( wire8314*  &  wire7581* ) ;
 assign wire8313 = ( I1767 ) | ( I1766 ) ;
 assign I1766 = ( wire7602*  &  wire7377* ) ;
 assign I1767 = ( wire8309*  &  wire7604* ) ;
 assign new_D<86> = ( wire8313 ) | ( wire1255 ) | ( wire8311 ) | ( wire1252 ) ;
 assign wire1246 = ( wire7600*  &  wire7377* ) ;
 assign wire7407 = ( D<83>* ) ;
 assign wire8316 = ( I1773 ) | ( I1772 ) ;
 assign I1772 = ( wire7597*  &  wire7407* ) ;
 assign I1773 = ( wire7598*  &  wire7378* ) ;
 assign wire8319 = ( key<246>* ) ;
 assign wire1249 = ( wire8319*  &  wire7581* ) ;
 assign wire8318 = ( I1778 ) | ( I1777 ) ;
 assign I1777 = ( wire7602*  &  wire7397* ) ;
 assign I1778 = ( wire8314*  &  wire7604* ) ;
 assign new_D<85> = ( wire8318 ) | ( wire1249 ) | ( wire8316 ) | ( wire1246 ) ;
 assign wire1240 = ( wire7600*  &  wire7397* ) ;
 assign wire7417 = ( D<82>* ) ;
 assign wire8321 = ( I1784 ) | ( I1783 ) ;
 assign I1783 = ( wire7597*  &  wire7417* ) ;
 assign I1784 = ( wire7598*  &  wire7407* ) ;
 assign wire8324 = ( key<254>* ) ;
 assign wire1243 = ( wire8324*  &  wire7581* ) ;
 assign wire8323 = ( I1789 ) | ( I1788 ) ;
 assign I1788 = ( wire7602*  &  wire7393* ) ;
 assign I1789 = ( wire8319*  &  wire7604* ) ;
 assign new_D<84> = ( wire8323 ) | ( wire1243 ) | ( wire8321 ) | ( wire1240 ) ;
 assign wire1234 = ( wire7600*  &  wire7393* ) ;
 assign wire8326 = ( D<81>* ) ;
 assign wire8327 = ( I1795 ) | ( I1794 ) ;
 assign I1794 = ( wire8326*  &  wire7597* ) ;
 assign I1795 = ( wire7598*  &  wire7417* ) ;
 assign wire8330 = ( key<131>* ) ;
 assign wire1237 = ( wire8330*  &  wire7581* ) ;
 assign wire8329 = ( I1800 ) | ( I1799 ) ;
 assign I1799 = ( wire7602*  &  wire7378* ) ;
 assign I1800 = ( wire8324*  &  wire7604* ) ;
 assign new_D<83> = ( wire8329 ) | ( wire1237 ) | ( wire8327 ) | ( wire1234 ) ;
 assign wire1228 = ( wire7600*  &  wire7378* ) ;
 assign wire7405 = ( D<80>* ) ;
 assign wire8332 = ( I1806 ) | ( I1805 ) ;
 assign I1805 = ( wire7597*  &  wire7405* ) ;
 assign I1806 = ( wire8326*  &  wire7598* ) ;
 assign wire8335 = ( key<139>* ) ;
 assign wire1231 = ( wire8335*  &  wire7581* ) ;
 assign wire8334 = ( I1811 ) | ( I1810 ) ;
 assign I1810 = ( wire7602*  &  wire7407* ) ;
 assign I1811 = ( wire8330*  &  wire7604* ) ;
 assign new_D<82> = ( wire8334 ) | ( wire1231 ) | ( wire8332 ) | ( wire1228 ) ;
 assign wire1222 = ( wire7600*  &  wire7407* ) ;
 assign wire7421 = ( D<79>* ) ;
 assign wire8337 = ( I1817 ) | ( I1816 ) ;
 assign I1816 = ( wire7597*  &  wire7421* ) ;
 assign I1817 = ( wire7598*  &  wire7405* ) ;
 assign wire8340 = ( key<147>* ) ;
 assign wire1225 = ( wire8340*  &  wire7581* ) ;
 assign wire8339 = ( I1822 ) | ( I1821 ) ;
 assign I1821 = ( wire7602*  &  wire7417* ) ;
 assign I1822 = ( wire8335*  &  wire7604* ) ;
 assign new_D<81> = ( wire8339 ) | ( wire1225 ) | ( wire8337 ) | ( wire1222 ) ;
 assign wire1216 = ( wire7600*  &  wire7417* ) ;
 assign wire7414 = ( D<78>* ) ;
 assign wire8342 = ( I1828 ) | ( I1827 ) ;
 assign I1827 = ( wire7597*  &  wire7414* ) ;
 assign I1828 = ( wire7598*  &  wire7421* ) ;
 assign wire8345 = ( key<155>* ) ;
 assign wire1219 = ( wire8345*  &  wire7581* ) ;
 assign wire8344 = ( I1833 ) | ( I1832 ) ;
 assign I1832 = ( wire8326*  &  wire7602* ) ;
 assign I1833 = ( wire8340*  &  wire7604* ) ;
 assign new_D<80> = ( wire8344 ) | ( wire1219 ) | ( wire8342 ) | ( wire1216 ) ;
 assign wire1210 = ( wire8326*  &  wire7600* ) ;
 assign wire7402 = ( D<77>* ) ;
 assign wire8347 = ( I1839 ) | ( I1838 ) ;
 assign I1838 = ( wire7597*  &  wire7402* ) ;
 assign I1839 = ( wire7598*  &  wire7414* ) ;
 assign wire8350 = ( key<132>* ) ;
 assign wire1213 = ( wire8350*  &  wire7581* ) ;
 assign wire8349 = ( I1844 ) | ( I1843 ) ;
 assign I1843 = ( wire7602*  &  wire7405* ) ;
 assign I1844 = ( wire8345*  &  wire7604* ) ;
 assign new_D<79> = ( wire8349 ) | ( wire1213 ) | ( wire8347 ) | ( wire1210 ) ;
 assign wire1204 = ( wire7600*  &  wire7405* ) ;
 assign wire7409 = ( D<76>* ) ;
 assign wire8352 = ( I1850 ) | ( I1849 ) ;
 assign I1849 = ( wire7597*  &  wire7409* ) ;
 assign I1850 = ( wire7598*  &  wire7402* ) ;
 assign wire8355 = ( key<140>* ) ;
 assign wire1207 = ( wire8355*  &  wire7581* ) ;
 assign wire8354 = ( I1855 ) | ( I1854 ) ;
 assign I1854 = ( wire7602*  &  wire7421* ) ;
 assign I1855 = ( wire8350*  &  wire7604* ) ;
 assign new_D<78> = ( wire8354 ) | ( wire1207 ) | ( wire8352 ) | ( wire1204 ) ;
 assign wire1198 = ( wire7600*  &  wire7421* ) ;
 assign wire7411 = ( D<75>* ) ;
 assign wire8357 = ( I1861 ) | ( I1860 ) ;
 assign I1860 = ( wire7597*  &  wire7411* ) ;
 assign I1861 = ( wire7598*  &  wire7409* ) ;
 assign wire8360 = ( key<148>* ) ;
 assign wire1201 = ( wire8360*  &  wire7581* ) ;
 assign wire8359 = ( I1866 ) | ( I1865 ) ;
 assign I1865 = ( wire7602*  &  wire7414* ) ;
 assign I1866 = ( wire8355*  &  wire7604* ) ;
 assign new_D<77> = ( wire8359 ) | ( wire1201 ) | ( wire8357 ) | ( wire1198 ) ;
 assign wire1192 = ( wire7600*  &  wire7414* ) ;
 assign wire7418 = ( D<74>* ) ;
 assign wire8362 = ( I1872 ) | ( I1871 ) ;
 assign I1871 = ( wire7597*  &  wire7418* ) ;
 assign I1872 = ( wire7598*  &  wire7411* ) ;
 assign wire8365 = ( key<156>* ) ;
 assign wire1195 = ( wire8365*  &  wire7581* ) ;
 assign wire8364 = ( I1877 ) | ( I1876 ) ;
 assign I1876 = ( wire7602*  &  wire7402* ) ;
 assign I1877 = ( wire8360*  &  wire7604* ) ;
 assign new_D<76> = ( wire8364 ) | ( wire1195 ) | ( wire8362 ) | ( wire1192 ) ;
 assign wire1186 = ( wire7600*  &  wire7402* ) ;
 assign wire7404 = ( D<73>* ) ;
 assign wire8367 = ( I1883 ) | ( I1882 ) ;
 assign I1882 = ( wire7597*  &  wire7404* ) ;
 assign I1883 = ( wire7598*  &  wire7418* ) ;
 assign wire8370 = ( key<164>* ) ;
 assign wire1189 = ( wire8370*  &  wire7581* ) ;
 assign wire8369 = ( I1888 ) | ( I1887 ) ;
 assign I1887 = ( wire7602*  &  wire7409* ) ;
 assign I1888 = ( wire8365*  &  wire7604* ) ;
 assign new_D<75> = ( wire8369 ) | ( wire1189 ) | ( wire8367 ) | ( wire1186 ) ;
 assign wire1180 = ( wire7600*  &  wire7409* ) ;
 assign wire8372 = ( D<72>* ) ;
 assign wire8373 = ( I1894 ) | ( I1893 ) ;
 assign I1893 = ( wire8372*  &  wire7597* ) ;
 assign I1894 = ( wire7598*  &  wire7404* ) ;
 assign wire1183 = ( wire8229*  &  wire7581* ) ;
 assign wire8375 = ( I1898 ) | ( I1897 ) ;
 assign I1897 = ( wire7602*  &  wire7411* ) ;
 assign I1898 = ( wire8370*  &  wire7604* ) ;
 assign new_D<74> = ( wire8375 ) | ( wire1183 ) | ( wire8373 ) | ( wire1180 ) ;
 assign wire1174 = ( wire7600*  &  wire7411* ) ;
 assign wire7410 = ( D<71>* ) ;
 assign wire8377 = ( I1904 ) | ( I1903 ) ;
 assign I1903 = ( wire7597*  &  wire7410* ) ;
 assign I1904 = ( wire8372*  &  wire7598* ) ;
 assign wire8380 = ( key<180>* ) ;
 assign wire1177 = ( wire8380*  &  wire7581* ) ;
 assign wire8379 = ( I1909 ) | ( I1908 ) ;
 assign I1908 = ( wire7602*  &  wire7418* ) ;
 assign I1909 = ( wire8229*  &  wire7604* ) ;
 assign new_D<73> = ( wire8379 ) | ( wire1177 ) | ( wire8377 ) | ( wire1174 ) ;
 assign wire1168 = ( wire7600*  &  wire7418* ) ;
 assign wire7413 = ( D<70>* ) ;
 assign wire8382 = ( I1915 ) | ( I1914 ) ;
 assign I1914 = ( wire7597*  &  wire7413* ) ;
 assign I1915 = ( wire7598*  &  wire7410* ) ;
 assign wire8385 = ( key<188>* ) ;
 assign wire1171 = ( wire8385*  &  wire7581* ) ;
 assign wire8384 = ( I1920 ) | ( I1919 ) ;
 assign I1919 = ( wire7602*  &  wire7404* ) ;
 assign I1920 = ( wire8380*  &  wire7604* ) ;
 assign new_D<72> = ( wire8384 ) | ( wire1171 ) | ( wire8382 ) | ( wire1168 ) ;
 assign wire1162 = ( wire7600*  &  wire7404* ) ;
 assign wire7403 = ( D<69>* ) ;
 assign wire8387 = ( I1926 ) | ( I1925 ) ;
 assign I1925 = ( wire7597*  &  wire7403* ) ;
 assign I1926 = ( wire7598*  &  wire7413* ) ;
 assign wire8390 = ( key<133>* ) ;
 assign wire1165 = ( wire8390*  &  wire7581* ) ;
 assign wire8389 = ( I1931 ) | ( I1930 ) ;
 assign I1930 = ( wire8372*  &  wire7602* ) ;
 assign I1931 = ( wire8385*  &  wire7604* ) ;
 assign new_D<71> = ( wire8389 ) | ( wire1165 ) | ( wire8387 ) | ( wire1162 ) ;
 assign wire1156 = ( wire8372*  &  wire7600* ) ;
 assign wire7422 = ( D<68>* ) ;
 assign wire8392 = ( I1937 ) | ( I1936 ) ;
 assign I1936 = ( wire7597*  &  wire7422* ) ;
 assign I1937 = ( wire7598*  &  wire7403* ) ;
 assign wire8395 = ( key<141>* ) ;
 assign wire1159 = ( wire8395*  &  wire7581* ) ;
 assign wire8394 = ( I1942 ) | ( I1941 ) ;
 assign I1941 = ( wire7602*  &  wire7410* ) ;
 assign I1942 = ( wire8390*  &  wire7604* ) ;
 assign new_D<70> = ( wire8394 ) | ( wire1159 ) | ( wire8392 ) | ( wire1156 ) ;
 assign wire1150 = ( wire7600*  &  wire7410* ) ;
 assign wire7415 = ( D<67>* ) ;
 assign wire8397 = ( I1948 ) | ( I1947 ) ;
 assign I1947 = ( wire7597*  &  wire7415* ) ;
 assign I1948 = ( wire7598*  &  wire7422* ) ;
 assign wire8400 = ( key<149>* ) ;
 assign wire1153 = ( wire8400*  &  wire7581* ) ;
 assign wire8399 = ( I1953 ) | ( I1952 ) ;
 assign I1952 = ( wire7602*  &  wire7413* ) ;
 assign I1953 = ( wire8395*  &  wire7604* ) ;
 assign new_D<69> = ( wire8399 ) | ( wire1153 ) | ( wire8397 ) | ( wire1150 ) ;
 assign wire1144 = ( wire7600*  &  wire7413* ) ;
 assign wire7408 = ( D<66>* ) ;
 assign wire8402 = ( I1959 ) | ( I1958 ) ;
 assign I1958 = ( wire7597*  &  wire7408* ) ;
 assign I1959 = ( wire7598*  &  wire7415* ) ;
 assign wire8405 = ( key<157>* ) ;
 assign wire1147 = ( wire8405*  &  wire7581* ) ;
 assign wire8404 = ( I1964 ) | ( I1963 ) ;
 assign I1963 = ( wire7602*  &  wire7403* ) ;
 assign I1964 = ( wire8400*  &  wire7604* ) ;
 assign new_D<68> = ( wire8404 ) | ( wire1147 ) | ( wire8402 ) | ( wire1144 ) ;
 assign wire1138 = ( wire7600*  &  wire7403* ) ;
 assign wire8407 = ( D<65>* ) ;
 assign wire8408 = ( I1970 ) | ( I1969 ) ;
 assign I1969 = ( wire8407*  &  wire7597* ) ;
 assign I1970 = ( wire7598*  &  wire7408* ) ;
 assign wire8411 = ( key<165>* ) ;
 assign wire1141 = ( wire8411*  &  wire7581* ) ;
 assign wire8410 = ( I1975 ) | ( I1974 ) ;
 assign I1974 = ( wire7602*  &  wire7422* ) ;
 assign I1975 = ( wire8405*  &  wire7604* ) ;
 assign new_D<67> = ( wire8410 ) | ( wire1141 ) | ( wire8408 ) | ( wire1138 ) ;
 assign wire1132 = ( wire7600*  &  wire7422* ) ;
 assign wire7419 = ( D<64>* ) ;
 assign wire8413 = ( I1981 ) | ( I1980 ) ;
 assign I1980 = ( wire7597*  &  wire7419* ) ;
 assign I1981 = ( wire8407*  &  wire7598* ) ;
 assign wire8416 = ( key<173>* ) ;
 assign wire1135 = ( wire8416*  &  wire7581* ) ;
 assign wire8415 = ( I1986 ) | ( I1985 ) ;
 assign I1985 = ( wire7602*  &  wire7415* ) ;
 assign I1986 = ( wire8411*  &  wire7604* ) ;
 assign new_D<66> = ( wire8415 ) | ( wire1135 ) | ( wire8413 ) | ( wire1132 ) ;
 assign wire1126 = ( wire7600*  &  wire7415* ) ;
 assign wire7401 = ( D<63>* ) ;
 assign wire8418 = ( I1992 ) | ( I1991 ) ;
 assign I1991 = ( wire7597*  &  wire7401* ) ;
 assign I1992 = ( wire7598*  &  wire7419* ) ;
 assign wire8421 = ( key<181>* ) ;
 assign wire1129 = ( wire8421*  &  wire7581* ) ;
 assign wire8420 = ( I1997 ) | ( I1996 ) ;
 assign I1996 = ( wire7602*  &  wire7408* ) ;
 assign I1997 = ( wire8416*  &  wire7604* ) ;
 assign new_D<65> = ( wire8420 ) | ( wire1129 ) | ( wire8418 ) | ( wire1126 ) ;
 assign wire1120 = ( wire7600*  &  wire7408* ) ;
 assign wire8423 = ( D<62>* ) ;
 assign wire8424 = ( I2003 ) | ( I2002 ) ;
 assign I2002 = ( wire8423*  &  wire7597* ) ;
 assign I2003 = ( wire7598*  &  wire7401* ) ;
 assign wire8427 = ( key<189>* ) ;
 assign wire1123 = ( wire8427*  &  wire7581* ) ;
 assign wire8426 = ( I2008 ) | ( I2007 ) ;
 assign I2007 = ( wire8407*  &  wire7602* ) ;
 assign I2008 = ( wire8421*  &  wire7604* ) ;
 assign new_D<64> = ( wire8426 ) | ( wire1123 ) | ( wire8424 ) | ( wire1120 ) ;
 assign wire1114 = ( wire8407*  &  wire7600* ) ;
 assign wire7406 = ( D<61>* ) ;
 assign wire8429 = ( I2014 ) | ( I2013 ) ;
 assign I2013 = ( wire7597*  &  wire7406* ) ;
 assign I2014 = ( wire8423*  &  wire7598* ) ;
 assign wire8432 = ( key<134>* ) ;
 assign wire1117 = ( wire8432*  &  wire7581* ) ;
 assign wire8431 = ( I2019 ) | ( I2018 ) ;
 assign I2018 = ( wire7602*  &  wire7419* ) ;
 assign I2019 = ( wire8427*  &  wire7604* ) ;
 assign new_D<63> = ( wire8431 ) | ( wire1117 ) | ( wire8429 ) | ( wire1114 ) ;
 assign wire1108 = ( wire7600*  &  wire7419* ) ;
 assign wire7412 = ( D<60>* ) ;
 assign wire8434 = ( I2025 ) | ( I2024 ) ;
 assign I2024 = ( wire7597*  &  wire7412* ) ;
 assign I2025 = ( wire7598*  &  wire7406* ) ;
 assign wire8437 = ( key<142>* ) ;
 assign wire1111 = ( wire8437*  &  wire7581* ) ;
 assign wire8436 = ( I2030 ) | ( I2029 ) ;
 assign I2029 = ( wire7602*  &  wire7401* ) ;
 assign I2030 = ( wire8432*  &  wire7604* ) ;
 assign new_D<62> = ( wire8436 ) | ( wire1111 ) | ( wire8434 ) | ( wire1108 ) ;
 assign wire1102 = ( wire7600*  &  wire7401* ) ;
 assign wire7399 = ( D<59>* ) ;
 assign wire8439 = ( I2036 ) | ( I2035 ) ;
 assign I2035 = ( wire7597*  &  wire7399* ) ;
 assign I2036 = ( wire7598*  &  wire7412* ) ;
 assign wire8442 = ( key<150>* ) ;
 assign wire1105 = ( wire8442*  &  wire7581* ) ;
 assign wire8441 = ( I2041 ) | ( I2040 ) ;
 assign I2040 = ( wire8423*  &  wire7602* ) ;
 assign I2041 = ( wire8437*  &  wire7604* ) ;
 assign new_D<61> = ( wire8441 ) | ( wire1105 ) | ( wire8439 ) | ( wire1102 ) ;
 assign wire1096 = ( wire8423*  &  wire7600* ) ;
 assign wire7420 = ( D<58>* ) ;
 assign wire8444 = ( I2047 ) | ( I2046 ) ;
 assign I2046 = ( wire7597*  &  wire7420* ) ;
 assign I2047 = ( wire7598*  &  wire7399* ) ;
 assign wire8447 = ( key<158>* ) ;
 assign wire1099 = ( wire8447*  &  wire7581* ) ;
 assign wire8446 = ( I2052 ) | ( I2051 ) ;
 assign I2051 = ( wire7602*  &  wire7406* ) ;
 assign I2052 = ( wire8442*  &  wire7604* ) ;
 assign new_D<60> = ( wire8446 ) | ( wire1099 ) | ( wire8444 ) | ( wire1096 ) ;
 assign wire1090 = ( wire7600*  &  wire7406* ) ;
 assign wire7416 = ( D<57>* ) ;
 assign wire8449 = ( I2058 ) | ( I2057 ) ;
 assign I2057 = ( wire7597*  &  wire7416* ) ;
 assign I2058 = ( wire7598*  &  wire7420* ) ;
 assign wire8452 = ( key<166>* ) ;
 assign wire1093 = ( wire8452*  &  wire7581* ) ;
 assign wire8451 = ( I2063 ) | ( I2062 ) ;
 assign I2062 = ( wire7602*  &  wire7412* ) ;
 assign I2063 = ( wire8447*  &  wire7604* ) ;
 assign new_D<59> = ( wire8451 ) | ( wire1093 ) | ( wire8449 ) | ( wire1090 ) ;
 assign wire1084 = ( wire7600*  &  wire7412* ) ;
 assign wire7400 = ( D<56>* ) ;
 assign wire8454 = ( I2069 ) | ( I2068 ) ;
 assign I2068 = ( wire7597*  &  wire7400* ) ;
 assign I2069 = ( wire7598*  &  wire7416* ) ;
 assign wire8457 = ( key<174>* ) ;
 assign wire1087 = ( wire8457*  &  wire7581* ) ;
 assign wire8456 = ( I2074 ) | ( I2073 ) ;
 assign I2073 = ( wire7602*  &  wire7399* ) ;
 assign I2074 = ( wire8452*  &  wire7604* ) ;
 assign new_D<58> = ( wire8456 ) | ( wire1087 ) | ( wire8454 ) | ( wire1084 ) ;
 assign wire1078 = ( wire7600*  &  wire7399* ) ;
 assign wire7430 = ( D<55>* ) ;
 assign wire8459 = ( I2080 ) | ( I2079 ) ;
 assign I2079 = ( wire7597*  &  wire7430* ) ;
 assign I2080 = ( wire7598*  &  wire7400* ) ;
 assign wire8462 = ( key<182>* ) ;
 assign wire1081 = ( wire8462*  &  wire7581* ) ;
 assign wire8461 = ( I2085 ) | ( I2084 ) ;
 assign I2084 = ( wire7602*  &  wire7420* ) ;
 assign I2085 = ( wire8457*  &  wire7604* ) ;
 assign new_D<57> = ( wire8461 ) | ( wire1081 ) | ( wire8459 ) | ( wire1078 ) ;
 assign wire1072 = ( wire7600*  &  wire7420* ) ;
 assign wire7440 = ( D<54>* ) ;
 assign wire8464 = ( I2091 ) | ( I2090 ) ;
 assign I2090 = ( wire7597*  &  wire7440* ) ;
 assign I2091 = ( wire7598*  &  wire7430* ) ;
 assign wire8467 = ( key<190>* ) ;
 assign wire1075 = ( wire8467*  &  wire7581* ) ;
 assign wire8466 = ( I2096 ) | ( I2095 ) ;
 assign I2095 = ( wire7602*  &  wire7416* ) ;
 assign I2096 = ( wire8462*  &  wire7604* ) ;
 assign new_D<56> = ( wire8466 ) | ( wire1075 ) | ( wire8464 ) | ( wire1072 ) ;
 assign wire1066 = ( wire7600*  &  wire7416* ) ;
 assign wire8469 = ( D<53>* ) ;
 assign wire8470 = ( I2102 ) | ( I2101 ) ;
 assign I2101 = ( wire8469*  &  wire7597* ) ;
 assign I2102 = ( wire7598*  &  wire7440* ) ;
 assign wire8473 = ( key<67>* ) ;
 assign wire1069 = ( wire8473*  &  wire7581* ) ;
 assign wire8472 = ( I2107 ) | ( I2106 ) ;
 assign I2106 = ( wire7602*  &  wire7400* ) ;
 assign I2107 = ( wire8467*  &  wire7604* ) ;
 assign new_D<55> = ( wire8472 ) | ( wire1069 ) | ( wire8470 ) | ( wire1066 ) ;
 assign wire1060 = ( wire7600*  &  wire7400* ) ;
 assign wire7428 = ( D<52>* ) ;
 assign wire8475 = ( I2113 ) | ( I2112 ) ;
 assign I2112 = ( wire7597*  &  wire7428* ) ;
 assign I2113 = ( wire8469*  &  wire7598* ) ;
 assign wire8478 = ( key<75>* ) ;
 assign wire1063 = ( wire8478*  &  wire7581* ) ;
 assign wire8477 = ( I2118 ) | ( I2117 ) ;
 assign I2117 = ( wire7602*  &  wire7430* ) ;
 assign I2118 = ( wire8473*  &  wire7604* ) ;
 assign new_D<54> = ( wire8477 ) | ( wire1063 ) | ( wire8475 ) | ( wire1060 ) ;
 assign wire1054 = ( wire7600*  &  wire7430* ) ;
 assign wire7444 = ( D<51>* ) ;
 assign wire8480 = ( I2124 ) | ( I2123 ) ;
 assign I2123 = ( wire7597*  &  wire7444* ) ;
 assign I2124 = ( wire7598*  &  wire7428* ) ;
 assign wire8483 = ( key<83>* ) ;
 assign wire1057 = ( wire8483*  &  wire7581* ) ;
 assign wire8482 = ( I2129 ) | ( I2128 ) ;
 assign I2128 = ( wire7602*  &  wire7440* ) ;
 assign I2129 = ( wire8478*  &  wire7604* ) ;
 assign new_D<53> = ( wire8482 ) | ( wire1057 ) | ( wire8480 ) | ( wire1054 ) ;
 assign wire1048 = ( wire7600*  &  wire7440* ) ;
 assign wire7437 = ( D<50>* ) ;
 assign wire8485 = ( I2135 ) | ( I2134 ) ;
 assign I2134 = ( wire7597*  &  wire7437* ) ;
 assign I2135 = ( wire7598*  &  wire7444* ) ;
 assign wire8488 = ( key<91>* ) ;
 assign wire1051 = ( wire8488*  &  wire7581* ) ;
 assign wire8487 = ( I2140 ) | ( I2139 ) ;
 assign I2139 = ( wire8469*  &  wire7602* ) ;
 assign I2140 = ( wire8483*  &  wire7604* ) ;
 assign new_D<52> = ( wire8487 ) | ( wire1051 ) | ( wire8485 ) | ( wire1048 ) ;
 assign wire1042 = ( wire8469*  &  wire7600* ) ;
 assign wire7426 = ( D<49>* ) ;
 assign wire8490 = ( I2146 ) | ( I2145 ) ;
 assign I2145 = ( wire7597*  &  wire7426* ) ;
 assign I2146 = ( wire7598*  &  wire7437* ) ;
 assign wire8493 = ( key<68>* ) ;
 assign wire1045 = ( wire8493*  &  wire7581* ) ;
 assign wire8492 = ( I2151 ) | ( I2150 ) ;
 assign I2150 = ( wire7602*  &  wire7428* ) ;
 assign I2151 = ( wire8488*  &  wire7604* ) ;
 assign new_D<51> = ( wire8492 ) | ( wire1045 ) | ( wire8490 ) | ( wire1042 ) ;
 assign wire1036 = ( wire7600*  &  wire7428* ) ;
 assign wire7432 = ( D<48>* ) ;
 assign wire8495 = ( I2157 ) | ( I2156 ) ;
 assign I2156 = ( wire7597*  &  wire7432* ) ;
 assign I2157 = ( wire7598*  &  wire7426* ) ;
 assign wire8498 = ( key<76>* ) ;
 assign wire1039 = ( wire8498*  &  wire7581* ) ;
 assign wire8497 = ( I2162 ) | ( I2161 ) ;
 assign I2161 = ( wire7602*  &  wire7444* ) ;
 assign I2162 = ( wire8493*  &  wire7604* ) ;
 assign new_D<50> = ( wire8497 ) | ( wire1039 ) | ( wire8495 ) | ( wire1036 ) ;
 assign wire1030 = ( wire7600*  &  wire7444* ) ;
 assign wire7434 = ( D<47>* ) ;
 assign wire8500 = ( I2168 ) | ( I2167 ) ;
 assign I2167 = ( wire7597*  &  wire7434* ) ;
 assign I2168 = ( wire7598*  &  wire7432* ) ;
 assign wire8503 = ( key<84>* ) ;
 assign wire1033 = ( wire8503*  &  wire7581* ) ;
 assign wire8502 = ( I2173 ) | ( I2172 ) ;
 assign I2172 = ( wire7602*  &  wire7437* ) ;
 assign I2173 = ( wire8498*  &  wire7604* ) ;
 assign new_D<49> = ( wire8502 ) | ( wire1033 ) | ( wire8500 ) | ( wire1030 ) ;
 assign wire1024 = ( wire7600*  &  wire7437* ) ;
 assign wire7441 = ( D<46>* ) ;
 assign wire8505 = ( I2179 ) | ( I2178 ) ;
 assign I2178 = ( wire7597*  &  wire7441* ) ;
 assign I2179 = ( wire7598*  &  wire7434* ) ;
 assign wire8508 = ( key<92>* ) ;
 assign wire1027 = ( wire8508*  &  wire7581* ) ;
 assign wire8507 = ( I2184 ) | ( I2183 ) ;
 assign I2183 = ( wire7602*  &  wire7426* ) ;
 assign I2184 = ( wire8503*  &  wire7604* ) ;
 assign new_D<48> = ( wire8507 ) | ( wire1027 ) | ( wire8505 ) | ( wire1024 ) ;
 assign wire1018 = ( wire7600*  &  wire7426* ) ;
 assign wire7427 = ( D<45>* ) ;
 assign wire8510 = ( I2190 ) | ( I2189 ) ;
 assign I2189 = ( wire7597*  &  wire7427* ) ;
 assign I2190 = ( wire7598*  &  wire7441* ) ;
 assign wire8513 = ( key<100>* ) ;
 assign wire1021 = ( wire8513*  &  wire7581* ) ;
 assign wire8512 = ( I2195 ) | ( I2194 ) ;
 assign I2194 = ( wire7602*  &  wire7432* ) ;
 assign I2195 = ( wire8508*  &  wire7604* ) ;
 assign new_D<47> = ( wire8512 ) | ( wire1021 ) | ( wire8510 ) | ( wire1018 ) ;
 assign wire1012 = ( wire7600*  &  wire7432* ) ;
 assign wire7436 = ( D<44>* ) ;
 assign wire8515 = ( I2201 ) | ( I2200 ) ;
 assign I2200 = ( wire7597*  &  wire7436* ) ;
 assign I2201 = ( wire7598*  &  wire7427* ) ;
 assign wire8518 = ( key<44>* ) ;
 assign wire1015 = ( wire8518*  &  wire7581* ) ;
 assign wire8517 = ( I2206 ) | ( I2205 ) ;
 assign I2205 = ( wire7602*  &  wire7434* ) ;
 assign I2206 = ( wire8513*  &  wire7604* ) ;
 assign new_D<46> = ( wire8517 ) | ( wire1015 ) | ( wire8515 ) | ( wire1012 ) ;
 assign wire1006 = ( wire7600*  &  wire7434* ) ;
 assign wire7433 = ( D<43>* ) ;
 assign wire8520 = ( I2212 ) | ( I2211 ) ;
 assign I2211 = ( wire7597*  &  wire7433* ) ;
 assign I2212 = ( wire7598*  &  wire7436* ) ;
 assign wire8523 = ( key<116>* ) ;
 assign wire1009 = ( wire8523*  &  wire7581* ) ;
 assign wire8522 = ( I2217 ) | ( I2216 ) ;
 assign I2216 = ( wire7602*  &  wire7441* ) ;
 assign I2217 = ( wire8518*  &  wire7604* ) ;
 assign new_D<45> = ( wire8522 ) | ( wire1009 ) | ( wire8520 ) | ( wire1006 ) ;
 assign wire1000 = ( wire7600*  &  wire7441* ) ;
 assign wire8525 = ( D<42>* ) ;
 assign wire8526 = ( I2223 ) | ( I2222 ) ;
 assign I2222 = ( wire8525*  &  wire7597* ) ;
 assign I2223 = ( wire7598*  &  wire7433* ) ;
 assign wire8529 = ( key<124>* ) ;
 assign wire1003 = ( wire8529*  &  wire7581* ) ;
 assign wire8528 = ( I2228 ) | ( I2227 ) ;
 assign I2227 = ( wire7602*  &  wire7427* ) ;
 assign I2228 = ( wire8523*  &  wire7604* ) ;
 assign new_D<44> = ( wire8528 ) | ( wire1003 ) | ( wire8526 ) | ( wire1000 ) ;
 assign wire994 = ( wire7600*  &  wire7427* ) ;
 assign wire8531 = ( D<41>* ) ;
 assign wire8532 = ( I2234 ) | ( I2233 ) ;
 assign I2233 = ( wire8531*  &  wire7597* ) ;
 assign I2234 = ( wire8525*  &  wire7598* ) ;
 assign wire8535 = ( key<69>* ) ;
 assign wire997 = ( wire8535*  &  wire7581* ) ;
 assign wire8534 = ( I2239 ) | ( I2238 ) ;
 assign I2238 = ( wire7602*  &  wire7436* ) ;
 assign I2239 = ( wire8529*  &  wire7604* ) ;
 assign new_D<43> = ( wire8534 ) | ( wire997 ) | ( wire8532 ) | ( wire994 ) ;
 assign wire988 = ( wire7600*  &  wire7436* ) ;
 assign wire7445 = ( D<40>* ) ;
 assign wire8537 = ( I2245 ) | ( I2244 ) ;
 assign I2244 = ( wire7597*  &  wire7445* ) ;
 assign I2245 = ( wire8531*  &  wire7598* ) ;
 assign wire8540 = ( key<77>* ) ;
 assign wire991 = ( wire8540*  &  wire7581* ) ;
 assign wire8539 = ( I2250 ) | ( I2249 ) ;
 assign I2249 = ( wire7602*  &  wire7433* ) ;
 assign I2250 = ( wire8535*  &  wire7604* ) ;
 assign new_D<42> = ( wire8539 ) | ( wire991 ) | ( wire8537 ) | ( wire988 ) ;
 assign wire982 = ( wire7600*  &  wire7433* ) ;
 assign wire7438 = ( D<39>* ) ;
 assign wire8542 = ( I2256 ) | ( I2255 ) ;
 assign I2255 = ( wire7597*  &  wire7438* ) ;
 assign I2256 = ( wire7598*  &  wire7445* ) ;
 assign wire8545 = ( key<85>* ) ;
 assign wire985 = ( wire8545*  &  wire7581* ) ;
 assign wire8544 = ( I2261 ) | ( I2260 ) ;
 assign I2260 = ( wire8525*  &  wire7602* ) ;
 assign I2261 = ( wire8540*  &  wire7604* ) ;
 assign new_D<41> = ( wire8544 ) | ( wire985 ) | ( wire8542 ) | ( wire982 ) ;
 assign wire976 = ( wire8525*  &  wire7600* ) ;
 assign wire7431 = ( D<38>* ) ;
 assign wire8547 = ( I2267 ) | ( I2266 ) ;
 assign I2266 = ( wire7597*  &  wire7431* ) ;
 assign I2267 = ( wire7598*  &  wire7438* ) ;
 assign wire8550 = ( key<93>* ) ;
 assign wire979 = ( wire8550*  &  wire7581* ) ;
 assign wire8549 = ( I2272 ) | ( I2271 ) ;
 assign I2271 = ( wire8531*  &  wire7602* ) ;
 assign I2272 = ( wire8545*  &  wire7604* ) ;
 assign new_D<40> = ( wire8549 ) | ( wire979 ) | ( wire8547 ) | ( wire976 ) ;
 assign wire970 = ( wire8531*  &  wire7600* ) ;
 assign wire8552 = ( D<37>* ) ;
 assign wire8553 = ( I2278 ) | ( I2277 ) ;
 assign I2277 = ( wire8552*  &  wire7597* ) ;
 assign I2278 = ( wire7598*  &  wire7431* ) ;
 assign wire8556 = ( key<101>* ) ;
 assign wire973 = ( wire8556*  &  wire7581* ) ;
 assign wire8555 = ( I2283 ) | ( I2282 ) ;
 assign I2282 = ( wire7602*  &  wire7445* ) ;
 assign I2283 = ( wire8550*  &  wire7604* ) ;
 assign new_D<39> = ( wire8555 ) | ( wire973 ) | ( wire8553 ) | ( wire970 ) ;
 assign wire964 = ( wire7600*  &  wire7445* ) ;
 assign wire7442 = ( D<36>* ) ;
 assign wire8558 = ( I2289 ) | ( I2288 ) ;
 assign I2288 = ( wire7597*  &  wire7442* ) ;
 assign I2289 = ( wire8552*  &  wire7598* ) ;
 assign wire8561 = ( key<109>* ) ;
 assign wire967 = ( wire8561*  &  wire7581* ) ;
 assign wire8560 = ( I2294 ) | ( I2293 ) ;
 assign I2293 = ( wire7602*  &  wire7438* ) ;
 assign I2294 = ( wire8556*  &  wire7604* ) ;
 assign new_D<38> = ( wire8560 ) | ( wire967 ) | ( wire8558 ) | ( wire964 ) ;
 assign wire958 = ( wire7600*  &  wire7438* ) ;
 assign wire7425 = ( D<35>* ) ;
 assign wire8563 = ( I2300 ) | ( I2299 ) ;
 assign I2299 = ( wire7597*  &  wire7425* ) ;
 assign I2300 = ( wire7598*  &  wire7442* ) ;
 assign wire8566 = ( key<117>* ) ;
 assign wire961 = ( wire8566*  &  wire7581* ) ;
 assign wire8565 = ( I2305 ) | ( I2304 ) ;
 assign I2304 = ( wire7602*  &  wire7431* ) ;
 assign I2305 = ( wire8561*  &  wire7604* ) ;
 assign new_D<37> = ( wire8565 ) | ( wire961 ) | ( wire8563 ) | ( wire958 ) ;
 assign wire952 = ( wire7600*  &  wire7431* ) ;
 assign wire8568 = ( D<34>* ) ;
 assign wire8569 = ( I2311 ) | ( I2310 ) ;
 assign I2310 = ( wire8568*  &  wire7597* ) ;
 assign I2311 = ( wire7598*  &  wire7425* ) ;
 assign wire8572 = ( key<125>* ) ;
 assign wire955 = ( wire8572*  &  wire7581* ) ;
 assign wire8571 = ( I2316 ) | ( I2315 ) ;
 assign I2315 = ( wire8552*  &  wire7602* ) ;
 assign I2316 = ( wire8566*  &  wire7604* ) ;
 assign new_D<36> = ( wire8571 ) | ( wire955 ) | ( wire8569 ) | ( wire952 ) ;
 assign wire946 = ( wire8552*  &  wire7600* ) ;
 assign wire7429 = ( D<33>* ) ;
 assign wire8574 = ( I2322 ) | ( I2321 ) ;
 assign I2321 = ( wire7597*  &  wire7429* ) ;
 assign I2322 = ( wire8568*  &  wire7598* ) ;
 assign wire8577 = ( key<70>* ) ;
 assign wire949 = ( wire8577*  &  wire7581* ) ;
 assign wire8576 = ( I2327 ) | ( I2326 ) ;
 assign I2326 = ( wire7602*  &  wire7442* ) ;
 assign I2327 = ( wire8572*  &  wire7604* ) ;
 assign new_D<35> = ( wire8576 ) | ( wire949 ) | ( wire8574 ) | ( wire946 ) ;
 assign wire940 = ( wire7600*  &  wire7442* ) ;
 assign wire7435 = ( D<32>* ) ;
 assign wire8579 = ( I2333 ) | ( I2332 ) ;
 assign I2332 = ( wire7597*  &  wire7435* ) ;
 assign I2333 = ( wire7598*  &  wire7429* ) ;
 assign wire8582 = ( key<78>* ) ;
 assign wire943 = ( wire8582*  &  wire7581* ) ;
 assign wire8581 = ( I2338 ) | ( I2337 ) ;
 assign I2337 = ( wire7602*  &  wire7425* ) ;
 assign I2338 = ( wire8577*  &  wire7604* ) ;
 assign new_D<34> = ( wire8581 ) | ( wire943 ) | ( wire8579 ) | ( wire940 ) ;
 assign wire934 = ( wire7600*  &  wire7425* ) ;
 assign wire7423 = ( D<31>* ) ;
 assign wire8584 = ( I2344 ) | ( I2343 ) ;
 assign I2343 = ( wire7597*  &  wire7423* ) ;
 assign I2344 = ( wire7598*  &  wire7435* ) ;
 assign wire8587 = ( key<86>* ) ;
 assign wire937 = ( wire8587*  &  wire7581* ) ;
 assign wire8586 = ( I2349 ) | ( I2348 ) ;
 assign I2348 = ( wire8568*  &  wire7602* ) ;
 assign I2349 = ( wire8582*  &  wire7604* ) ;
 assign new_D<33> = ( wire8586 ) | ( wire937 ) | ( wire8584 ) | ( wire934 ) ;
 assign wire928 = ( wire8568*  &  wire7600* ) ;
 assign wire7443 = ( D<30>* ) ;
 assign wire8589 = ( I2355 ) | ( I2354 ) ;
 assign I2354 = ( wire7597*  &  wire7443* ) ;
 assign I2355 = ( wire7598*  &  wire7423* ) ;
 assign wire8592 = ( key<94>* ) ;
 assign wire931 = ( wire8592*  &  wire7581* ) ;
 assign wire8591 = ( I2360 ) | ( I2359 ) ;
 assign I2359 = ( wire7602*  &  wire7429* ) ;
 assign I2360 = ( wire8587*  &  wire7604* ) ;
 assign new_D<32> = ( wire8591 ) | ( wire931 ) | ( wire8589 ) | ( wire928 ) ;
 assign wire922 = ( wire7600*  &  wire7429* ) ;
 assign wire7439 = ( D<29>* ) ;
 assign wire8594 = ( I2366 ) | ( I2365 ) ;
 assign I2365 = ( wire7597*  &  wire7439* ) ;
 assign I2366 = ( wire7598*  &  wire7443* ) ;
 assign wire8597 = ( key<102>* ) ;
 assign wire925 = ( wire8597*  &  wire7581* ) ;
 assign wire8596 = ( I2371 ) | ( I2370 ) ;
 assign I2370 = ( wire7602*  &  wire7435* ) ;
 assign I2371 = ( wire8592*  &  wire7604* ) ;
 assign new_D<31> = ( wire8596 ) | ( wire925 ) | ( wire8594 ) | ( wire922 ) ;
 assign wire916 = ( wire7600*  &  wire7435* ) ;
 assign wire7424 = ( D<28>* ) ;
 assign wire8599 = ( I2377 ) | ( I2376 ) ;
 assign I2376 = ( wire7597*  &  wire7424* ) ;
 assign I2377 = ( wire7598*  &  wire7439* ) ;
 assign wire8602 = ( key<110>* ) ;
 assign wire919 = ( wire8602*  &  wire7581* ) ;
 assign wire8601 = ( I2382 ) | ( I2381 ) ;
 assign I2381 = ( wire7602*  &  wire7423* ) ;
 assign I2382 = ( wire8597*  &  wire7604* ) ;
 assign new_D<30> = ( wire8601 ) | ( wire919 ) | ( wire8599 ) | ( wire916 ) ;
 assign wire910 = ( wire7600*  &  wire7423* ) ;
 assign wire7454 = ( D<27>* ) ;
 assign wire8604 = ( I2388 ) | ( I2387 ) ;
 assign I2387 = ( wire7597*  &  wire7454* ) ;
 assign I2388 = ( wire7598*  &  wire7424* ) ;
 assign wire8607 = ( key<118>* ) ;
 assign wire913 = ( wire8607*  &  wire7581* ) ;
 assign wire8606 = ( I2393 ) | ( I2392 ) ;
 assign I2392 = ( wire7602*  &  wire7443* ) ;
 assign I2393 = ( wire8602*  &  wire7604* ) ;
 assign new_D<29> = ( wire8606 ) | ( wire913 ) | ( wire8604 ) | ( wire910 ) ;
 assign wire904 = ( wire7600*  &  wire7443* ) ;
 assign wire7464 = ( D<26>* ) ;
 assign wire8609 = ( I2399 ) | ( I2398 ) ;
 assign I2398 = ( wire7597*  &  wire7464* ) ;
 assign I2399 = ( wire7598*  &  wire7454* ) ;
 assign wire8612 = ( key<126>* ) ;
 assign wire907 = ( wire8612*  &  wire7581* ) ;
 assign wire8611 = ( I2404 ) | ( I2403 ) ;
 assign I2403 = ( wire7602*  &  wire7439* ) ;
 assign I2404 = ( wire8607*  &  wire7604* ) ;
 assign new_D<28> = ( wire8611 ) | ( wire907 ) | ( wire8609 ) | ( wire904 ) ;
 assign wire898 = ( wire7600*  &  wire7439* ) ;
 assign wire8614 = ( D<25>* ) ;
 assign wire8615 = ( I2410 ) | ( I2409 ) ;
 assign I2409 = ( wire8614*  &  wire7597* ) ;
 assign I2410 = ( wire7598*  &  wire7464* ) ;
 assign wire8618 = ( key<3>* ) ;
 assign wire901 = ( wire8618*  &  wire7581* ) ;
 assign wire8617 = ( I2415 ) | ( I2414 ) ;
 assign I2414 = ( wire7602*  &  wire7424* ) ;
 assign I2415 = ( wire8612*  &  wire7604* ) ;
 assign new_D<27> = ( wire8617 ) | ( wire901 ) | ( wire8615 ) | ( wire898 ) ;
 assign wire892 = ( wire7600*  &  wire7424* ) ;
 assign wire7452 = ( D<24>* ) ;
 assign wire8620 = ( I2421 ) | ( I2420 ) ;
 assign I2420 = ( wire7597*  &  wire7452* ) ;
 assign I2421 = ( wire8614*  &  wire7598* ) ;
 assign wire8623 = ( key<11>* ) ;
 assign wire895 = ( wire8623*  &  wire7581* ) ;
 assign wire8622 = ( I2426 ) | ( I2425 ) ;
 assign I2425 = ( wire7602*  &  wire7454* ) ;
 assign I2426 = ( wire8618*  &  wire7604* ) ;
 assign new_D<26> = ( wire8622 ) | ( wire895 ) | ( wire8620 ) | ( wire892 ) ;
 assign wire886 = ( wire7600*  &  wire7454* ) ;
 assign wire7468 = ( D<23>* ) ;
 assign wire8625 = ( I2432 ) | ( I2431 ) ;
 assign I2431 = ( wire7597*  &  wire7468* ) ;
 assign I2432 = ( wire7598*  &  wire7452* ) ;
 assign wire8628 = ( key<19>* ) ;
 assign wire889 = ( wire8628*  &  wire7581* ) ;
 assign wire8627 = ( I2437 ) | ( I2436 ) ;
 assign I2436 = ( wire7602*  &  wire7464* ) ;
 assign I2437 = ( wire8623*  &  wire7604* ) ;
 assign new_D<25> = ( wire8627 ) | ( wire889 ) | ( wire8625 ) | ( wire886 ) ;
 assign wire880 = ( wire7600*  &  wire7464* ) ;
 assign wire7461 = ( D<22>* ) ;
 assign wire8630 = ( I2443 ) | ( I2442 ) ;
 assign I2442 = ( wire7597*  &  wire7461* ) ;
 assign I2443 = ( wire7598*  &  wire7468* ) ;
 assign wire8633 = ( key<27>* ) ;
 assign wire883 = ( wire8633*  &  wire7581* ) ;
 assign wire8632 = ( I2448 ) | ( I2447 ) ;
 assign I2447 = ( wire8614*  &  wire7602* ) ;
 assign I2448 = ( wire8628*  &  wire7604* ) ;
 assign new_D<24> = ( wire8632 ) | ( wire883 ) | ( wire8630 ) | ( wire880 ) ;
 assign wire874 = ( wire8614*  &  wire7600* ) ;
 assign wire7449 = ( D<21>* ) ;
 assign wire8635 = ( I2454 ) | ( I2453 ) ;
 assign I2453 = ( wire7597*  &  wire7449* ) ;
 assign I2454 = ( wire7598*  &  wire7461* ) ;
 assign wire8638 = ( key<4>* ) ;
 assign wire877 = ( wire8638*  &  wire7581* ) ;
 assign wire8637 = ( I2459 ) | ( I2458 ) ;
 assign I2458 = ( wire7602*  &  wire7452* ) ;
 assign I2459 = ( wire8633*  &  wire7604* ) ;
 assign new_D<23> = ( wire8637 ) | ( wire877 ) | ( wire8635 ) | ( wire874 ) ;
 assign wire868 = ( wire7600*  &  wire7452* ) ;
 assign wire7456 = ( D<20>* ) ;
 assign wire8640 = ( I2465 ) | ( I2464 ) ;
 assign I2464 = ( wire7597*  &  wire7456* ) ;
 assign I2465 = ( wire7598*  &  wire7449* ) ;
 assign wire8643 = ( key<12>* ) ;
 assign wire871 = ( wire8643*  &  wire7581* ) ;
 assign wire8642 = ( I2470 ) | ( I2469 ) ;
 assign I2469 = ( wire7602*  &  wire7468* ) ;
 assign I2470 = ( wire8638*  &  wire7604* ) ;
 assign new_D<22> = ( wire8642 ) | ( wire871 ) | ( wire8640 ) | ( wire868 ) ;
 assign wire862 = ( wire7600*  &  wire7468* ) ;
 assign wire7458 = ( D<19>* ) ;
 assign wire8645 = ( I2476 ) | ( I2475 ) ;
 assign I2475 = ( wire7597*  &  wire7458* ) ;
 assign I2476 = ( wire7598*  &  wire7456* ) ;
 assign wire8648 = ( key<20>* ) ;
 assign wire865 = ( wire8648*  &  wire7581* ) ;
 assign wire8647 = ( I2481 ) | ( I2480 ) ;
 assign I2480 = ( wire7602*  &  wire7461* ) ;
 assign I2481 = ( wire8643*  &  wire7604* ) ;
 assign new_D<21> = ( wire8647 ) | ( wire865 ) | ( wire8645 ) | ( wire862 ) ;
 assign wire856 = ( wire7600*  &  wire7461* ) ;
 assign wire7465 = ( D<18>* ) ;
 assign wire8650 = ( I2487 ) | ( I2486 ) ;
 assign I2486 = ( wire7597*  &  wire7465* ) ;
 assign I2487 = ( wire7598*  &  wire7458* ) ;
 assign wire8653 = ( key<28>* ) ;
 assign wire859 = ( wire8653*  &  wire7581* ) ;
 assign wire8652 = ( I2492 ) | ( I2491 ) ;
 assign I2491 = ( wire7602*  &  wire7449* ) ;
 assign I2492 = ( wire8648*  &  wire7604* ) ;
 assign new_D<20> = ( wire8652 ) | ( wire859 ) | ( wire8650 ) | ( wire856 ) ;
 assign wire850 = ( wire7600*  &  wire7449* ) ;
 assign wire7451 = ( D<17>* ) ;
 assign wire8655 = ( I2498 ) | ( I2497 ) ;
 assign I2497 = ( wire7597*  &  wire7451* ) ;
 assign I2498 = ( wire7598*  &  wire7465* ) ;
 assign wire8658 = ( key<36>* ) ;
 assign wire853 = ( wire8658*  &  wire7581* ) ;
 assign wire8657 = ( I2503 ) | ( I2502 ) ;
 assign I2502 = ( wire7602*  &  wire7456* ) ;
 assign I2503 = ( wire8653*  &  wire7604* ) ;
 assign new_D<19> = ( wire8657 ) | ( wire853 ) | ( wire8655 ) | ( wire850 ) ;
 assign wire844 = ( wire7600*  &  wire7456* ) ;
 assign wire7460 = ( D<16>* ) ;
 assign wire8660 = ( I2509 ) | ( I2508 ) ;
 assign I2508 = ( wire7597*  &  wire7460* ) ;
 assign I2509 = ( wire7598*  &  wire7451* ) ;
 assign wire847 = ( wire8518*  &  wire7581* ) ;
 assign wire8662 = ( I2513 ) | ( I2512 ) ;
 assign I2512 = ( wire7602*  &  wire7458* ) ;
 assign I2513 = ( wire8658*  &  wire7604* ) ;
 assign new_D<18> = ( wire8662 ) | ( wire847 ) | ( wire8660 ) | ( wire844 ) ;
 assign wire838 = ( wire7600*  &  wire7458* ) ;
 assign wire7457 = ( D<15>* ) ;
 assign wire8664 = ( I2519 ) | ( I2518 ) ;
 assign I2518 = ( wire7597*  &  wire7457* ) ;
 assign I2519 = ( wire7598*  &  wire7460* ) ;
 assign wire8667 = ( key<52>* ) ;
 assign wire841 = ( wire8667*  &  wire7581* ) ;
 assign wire8666 = ( I2524 ) | ( I2523 ) ;
 assign I2523 = ( wire7602*  &  wire7465* ) ;
 assign I2524 = ( wire8518*  &  wire7604* ) ;
 assign new_D<17> = ( wire8666 ) | ( wire841 ) | ( wire8664 ) | ( wire838 ) ;
 assign wire832 = ( wire7600*  &  wire7465* ) ;
 assign wire8669 = ( D<14>* ) ;
 assign wire8670 = ( I2530 ) | ( I2529 ) ;
 assign I2529 = ( wire8669*  &  wire7597* ) ;
 assign I2530 = ( wire7598*  &  wire7457* ) ;
 assign wire8673 = ( key<60>* ) ;
 assign wire835 = ( wire8673*  &  wire7581* ) ;
 assign wire8672 = ( I2535 ) | ( I2534 ) ;
 assign I2534 = ( wire7602*  &  wire7451* ) ;
 assign I2535 = ( wire8667*  &  wire7604* ) ;
 assign new_D<16> = ( wire8672 ) | ( wire835 ) | ( wire8670 ) | ( wire832 ) ;
 assign wire826 = ( wire7600*  &  wire7451* ) ;
 assign wire7450 = ( D<13>* ) ;
 assign wire8675 = ( I2541 ) | ( I2540 ) ;
 assign I2540 = ( wire7597*  &  wire7450* ) ;
 assign I2541 = ( wire8669*  &  wire7598* ) ;
 assign wire8678 = ( key<5>* ) ;
 assign wire829 = ( wire8678*  &  wire7581* ) ;
 assign wire8677 = ( I2546 ) | ( I2545 ) ;
 assign I2545 = ( wire7602*  &  wire7460* ) ;
 assign I2546 = ( wire8673*  &  wire7604* ) ;
 assign new_D<15> = ( wire8677 ) | ( wire829 ) | ( wire8675 ) | ( wire826 ) ;
 assign wire820 = ( wire7600*  &  wire7460* ) ;
 assign wire7469 = ( D<12>* ) ;
 assign wire8680 = ( I2552 ) | ( I2551 ) ;
 assign I2551 = ( wire7597*  &  wire7469* ) ;
 assign I2552 = ( wire7598*  &  wire7450* ) ;
 assign wire8683 = ( key<13>* ) ;
 assign wire823 = ( wire8683*  &  wire7581* ) ;
 assign wire8682 = ( I2557 ) | ( I2556 ) ;
 assign I2556 = ( wire7602*  &  wire7457* ) ;
 assign I2557 = ( wire8678*  &  wire7604* ) ;
 assign new_D<14> = ( wire8682 ) | ( wire823 ) | ( wire8680 ) | ( wire820 ) ;
 assign wire814 = ( wire7600*  &  wire7457* ) ;
 assign wire7462 = ( D<11>* ) ;
 assign wire8685 = ( I2563 ) | ( I2562 ) ;
 assign I2562 = ( wire7597*  &  wire7462* ) ;
 assign I2563 = ( wire7598*  &  wire7469* ) ;
 assign wire8688 = ( key<21>* ) ;
 assign wire817 = ( wire8688*  &  wire7581* ) ;
 assign wire8687 = ( I2568 ) | ( I2567 ) ;
 assign I2567 = ( wire8669*  &  wire7602* ) ;
 assign I2568 = ( wire8683*  &  wire7604* ) ;
 assign new_D<13> = ( wire8687 ) | ( wire817 ) | ( wire8685 ) | ( wire814 ) ;
 assign wire808 = ( wire8669*  &  wire7600* ) ;
 assign wire7455 = ( D<10>* ) ;
 assign wire8690 = ( I2574 ) | ( I2573 ) ;
 assign I2573 = ( wire7597*  &  wire7455* ) ;
 assign I2574 = ( wire7598*  &  wire7462* ) ;
 assign wire8693 = ( key<29>* ) ;
 assign wire811 = ( wire8693*  &  wire7581* ) ;
 assign wire8692 = ( I2579 ) | ( I2578 ) ;
 assign I2578 = ( wire7602*  &  wire7450* ) ;
 assign I2579 = ( wire8688*  &  wire7604* ) ;
 assign new_D<12> = ( wire8692 ) | ( wire811 ) | ( wire8690 ) | ( wire808 ) ;
 assign wire802 = ( wire7600*  &  wire7450* ) ;
 assign wire8695 = ( D<9>* ) ;
 assign wire8696 = ( I2585 ) | ( I2584 ) ;
 assign I2584 = ( wire8695*  &  wire7597* ) ;
 assign I2585 = ( wire7598*  &  wire7455* ) ;
 assign wire8699 = ( key<37>* ) ;
 assign wire805 = ( wire8699*  &  wire7581* ) ;
 assign wire8698 = ( I2590 ) | ( I2589 ) ;
 assign I2589 = ( wire7602*  &  wire7469* ) ;
 assign I2590 = ( wire8693*  &  wire7604* ) ;
 assign new_D<11> = ( wire8698 ) | ( wire805 ) | ( wire8696 ) | ( wire802 ) ;
 assign wire796 = ( wire7600*  &  wire7469* ) ;
 assign wire7466 = ( D<8>* ) ;
 assign wire8701 = ( I2596 ) | ( I2595 ) ;
 assign I2595 = ( wire7597*  &  wire7466* ) ;
 assign I2596 = ( wire8695*  &  wire7598* ) ;
 assign wire8704 = ( key<45>* ) ;
 assign wire799 = ( wire8704*  &  wire7581* ) ;
 assign wire8703 = ( I2601 ) | ( I2600 ) ;
 assign I2600 = ( wire7602*  &  wire7462* ) ;
 assign I2601 = ( wire8699*  &  wire7604* ) ;
 assign new_D<10> = ( wire8703 ) | ( wire799 ) | ( wire8701 ) | ( wire796 ) ;
 assign wire790 = ( wire7600*  &  wire7462* ) ;
 assign wire7448 = ( D<7>* ) ;
 assign wire8706 = ( I2607 ) | ( I2606 ) ;
 assign I2606 = ( wire7597*  &  wire7448* ) ;
 assign I2607 = ( wire7598*  &  wire7466* ) ;
 assign wire8709 = ( key<53>* ) ;
 assign wire793 = ( wire8709*  &  wire7581* ) ;
 assign wire8708 = ( I2612 ) | ( I2611 ) ;
 assign I2611 = ( wire7602*  &  wire7455* ) ;
 assign I2612 = ( wire8704*  &  wire7604* ) ;
 assign new_D<9> = ( wire8708 ) | ( wire793 ) | ( wire8706 ) | ( wire790 ) ;
 assign wire784 = ( wire7600*  &  wire7455* ) ;
 assign wire8711 = ( D<6>* ) ;
 assign wire8712 = ( I2618 ) | ( I2617 ) ;
 assign I2617 = ( wire8711*  &  wire7597* ) ;
 assign I2618 = ( wire7598*  &  wire7448* ) ;
 assign wire8715 = ( key<61>* ) ;
 assign wire787 = ( wire8715*  &  wire7581* ) ;
 assign wire8714 = ( I2623 ) | ( I2622 ) ;
 assign I2622 = ( wire8695*  &  wire7602* ) ;
 assign I2623 = ( wire8709*  &  wire7604* ) ;
 assign new_D<8> = ( wire8714 ) | ( wire787 ) | ( wire8712 ) | ( wire784 ) ;
 assign wire778 = ( wire8695*  &  wire7600* ) ;
 assign wire7453 = ( D<5>* ) ;
 assign wire8717 = ( I2629 ) | ( I2628 ) ;
 assign I2628 = ( wire7597*  &  wire7453* ) ;
 assign I2629 = ( wire8711*  &  wire7598* ) ;
 assign wire8720 = ( key<6>* ) ;
 assign wire781 = ( wire8720*  &  wire7581* ) ;
 assign wire8719 = ( I2634 ) | ( I2633 ) ;
 assign I2633 = ( wire7602*  &  wire7466* ) ;
 assign I2634 = ( wire8715*  &  wire7604* ) ;
 assign new_D<7> = ( wire8719 ) | ( wire781 ) | ( wire8717 ) | ( wire778 ) ;
 assign wire772 = ( wire7600*  &  wire7466* ) ;
 assign wire7459 = ( D<4>* ) ;
 assign wire8722 = ( I2640 ) | ( I2639 ) ;
 assign I2639 = ( wire7597*  &  wire7459* ) ;
 assign I2640 = ( wire7598*  &  wire7453* ) ;
 assign wire8725 = ( key<14>* ) ;
 assign wire775 = ( wire8725*  &  wire7581* ) ;
 assign wire8724 = ( I2645 ) | ( I2644 ) ;
 assign I2644 = ( wire7602*  &  wire7448* ) ;
 assign I2645 = ( wire8720*  &  wire7604* ) ;
 assign new_D<6> = ( wire8724 ) | ( wire775 ) | ( wire8722 ) | ( wire772 ) ;
 assign wire766 = ( wire7600*  &  wire7448* ) ;
 assign wire7446 = ( D<3>* ) ;
 assign wire8727 = ( I2651 ) | ( I2650 ) ;
 assign I2650 = ( wire7597*  &  wire7446* ) ;
 assign I2651 = ( wire7598*  &  wire7459* ) ;
 assign wire8730 = ( key<22>* ) ;
 assign wire769 = ( wire8730*  &  wire7581* ) ;
 assign wire8729 = ( I2656 ) | ( I2655 ) ;
 assign I2655 = ( wire8711*  &  wire7602* ) ;
 assign I2656 = ( wire8725*  &  wire7604* ) ;
 assign new_D<5> = ( wire8729 ) | ( wire769 ) | ( wire8727 ) | ( wire766 ) ;
 assign wire760 = ( wire8711*  &  wire7600* ) ;
 assign wire7467 = ( D<2>* ) ;
 assign wire8732 = ( I2662 ) | ( I2661 ) ;
 assign I2661 = ( wire7597*  &  wire7467* ) ;
 assign I2662 = ( wire7598*  &  wire7446* ) ;
 assign wire8735 = ( key<30>* ) ;
 assign wire763 = ( wire8735*  &  wire7581* ) ;
 assign wire8734 = ( I2667 ) | ( I2666 ) ;
 assign I2666 = ( wire7602*  &  wire7453* ) ;
 assign I2667 = ( wire8730*  &  wire7604* ) ;
 assign new_D<4> = ( wire8734 ) | ( wire763 ) | ( wire8732 ) | ( wire760 ) ;
 assign wire754 = ( wire7600*  &  wire7453* ) ;
 assign wire8737 = ( I2672 ) | ( I2671 ) ;
 assign I2671 = ( wire7597*  &  wire7463* ) ;
 assign I2672 = ( wire7598*  &  wire7467* ) ;
 assign wire8740 = ( key<38>* ) ;
 assign wire757 = ( wire8740*  &  wire7581* ) ;
 assign wire8739 = ( I2677 ) | ( I2676 ) ;
 assign I2676 = ( wire7602*  &  wire7459* ) ;
 assign I2677 = ( wire8735*  &  wire7604* ) ;
 assign new_D<3> = ( wire8739 ) | ( wire757 ) | ( wire8737 ) | ( wire754 ) ;
 assign wire748 = ( wire7600*  &  wire7459* ) ;
 assign wire8742 = ( I2682 ) | ( I2681 ) ;
 assign I2681 = ( wire7597*  &  wire7447* ) ;
 assign I2682 = ( wire7598*  &  wire7463* ) ;
 assign wire8745 = ( key<46>* ) ;
 assign wire751 = ( wire8745*  &  wire7581* ) ;
 assign wire8744 = ( I2687 ) | ( I2686 ) ;
 assign I2686 = ( wire7602*  &  wire7446* ) ;
 assign I2687 = ( wire8740*  &  wire7604* ) ;
 assign new_D<2> = ( wire8744 ) | ( wire751 ) | ( wire8742 ) | ( wire748 ) ;
 assign wire742 = ( wire7600*  &  wire7446* ) ;
 assign wire8747 = ( I2692 ) | ( I2691 ) ;
 assign I2691 = ( wire7597*  &  wire7384* ) ;
 assign I2692 = ( wire7598*  &  wire7447* ) ;
 assign wire8750 = ( key<54>* ) ;
 assign wire745 = ( wire8750*  &  wire7581* ) ;
 assign wire8749 = ( I2697 ) | ( I2696 ) ;
 assign I2696 = ( wire7602*  &  wire7467* ) ;
 assign I2697 = ( wire8745*  &  wire7604* ) ;
 assign new_D<1> = ( wire8749 ) | ( wire745 ) | ( wire8747 ) | ( wire742 ) ;
 assign wire736 = ( wire7600*  &  wire7467* ) ;
 assign wire8752 = ( I2702 ) | ( I2701 ) ;
 assign I2701 = ( wire7597*  &  wire7394* ) ;
 assign I2702 = ( wire7598*  &  wire7384* ) ;
 assign wire739 = ( wire8182*  &  wire7581* ) ;
 assign wire8754 = ( I2706 ) | ( I2705 ) ;
 assign I2705 = ( wire7602*  &  wire7463* ) ;
 assign I2706 = ( wire8750*  &  wire7604* ) ;
 assign new_D<0> = ( wire8754 ) | ( wire739 ) | ( wire8752 ) | ( wire736 ) ;
 assign wire7596 = ( wire7573* ) | ( wire7566* ) ;
 assign wire7570 = ( count<1>* ) ;
 assign wire8756 = ( wire7570* ) | ( wire7569* ) | ( wire7591* ) ;
 assign wire8757 = ( wire11699* ) | ( wire7595* ) ;
 assign data_ready<0> = ( I2714 ) | ( I2713 ) ;
 assign I2713 = ( wire8756*  &  wire7596* ) ;
 assign I2714 = ( wire8757*  &  wire7574* ) ;
 assign start<0>* = ( (~ start<0>) ) ;
 assign wire7573* = ( (~ wire7573) ) ;
 assign encrypt<0>* = ( (~ encrypt<0>) ) ;
 assign count<2>* = ( (~ count<2>) ) ;
 assign wire7574* = ( (~ wire7574) ) ;
 assign wire7568* = ( (~ wire7568) ) ;
 assign count<0>* = ( (~ count<0>) ) ;
 assign count<1>* = ( (~ count<1>) ) ;
 assign wire7576* = ( (~ wire7576) ) ;
 assign wire11699* = ( (~ wire11699) ) ;
 assign main/$MINUS_4_1/c<0>8 =((~ key<254>) & key<254>);
 assign count<3>* = ( (~ count<3>) ) ;
 assign wire7575* = ( (~ wire7575) ) ;
 assign wire7577* = ( (~ wire7577) ) ;
 assign wire7565* = ( (~ wire7565) ) ;
 assign wire7566* = ( (~ wire7566) ) ;
 assign wire17163* = ( (~ wire17163) ) ;
 assign wire17165* = ( (~ wire17165) ) ;
 assign wire17167* = ( (~ wire17167) ) ;
 assign wire7581* = ( (~ wire7581) ) ;
 assign wire17157* = ( (~ wire17157) ) ;
 assign wire17159* = ( (~ wire17159) ) ;
 assign wire17161* = ( (~ wire17161) ) ;
 assign wire7571* = ( (~ wire7571) ) ;
 assign wire7586* = ( (~ wire7586) ) ;
 assign wire14444* = ( (~ wire14444) ) ;
 assign wire7587* = ( (~ wire7587) ) ;
 assign new_count<0>* = ( (~ new_count<0>) ) ;
 assign wire194* = ( (~ wire194) ) ;
 assign C<1>* = ( (~ C<1>) ) ;
 assign wire7569* = ( (~ wire7569) ) ;
 assign wire7580* = ( (~ wire7580) ) ;
 assign wire17145* = ( (~ wire17145) ) ;
 assign wire17147* = ( (~ wire17147) ) ;
 assign wire7541* = ( (~ wire7541) ) ;
 assign wire7600* = ( (~ wire7600) ) ;
 assign C<109>* = ( (~ C<109>) ) ;
 assign wire7591* = ( (~ wire7591) ) ;
 assign wire2079* = ( (~ wire2079) ) ;
 assign wire7292* = ( (~ wire7292) ) ;
 assign wire7572* = ( (~ wire7572) ) ;
 assign wire7284* = ( (~ wire7284) ) ;
 assign C<110>* = ( (~ C<110>) ) ;
 assign wire7595* = ( (~ wire7595) ) ;
 assign wire7475* = ( (~ wire7475) ) ;
 assign wire7597* = ( (~ wire7597) ) ;
 assign wire7473* = ( (~ wire7473) ) ;
 assign wire7598* = ( (~ wire7598) ) ;
 assign key<227>* = ( (~ key<227>) ) ;
 assign wire7606* = ( (~ wire7606) ) ;
 assign C<0>* = ( (~ C<0>) ) ;
 assign key<56>* = ( (~ key<56>) ) ;
 assign wire7560* = ( (~ wire7560) ) ;
 assign wire7602* = ( (~ wire7602) ) ;
 assign wire7603* = ( (~ wire7603) ) ;
 assign wire7604* = ( (~ wire7604) ) ;
 assign C<108>* = ( (~ C<108>) ) ;
 assign wire7608* = ( (~ wire7608) ) ;
 assign key<235>* = ( (~ key<235>) ) ;
 assign wire7612* = ( (~ wire7612) ) ;
 assign C<111>* = ( (~ C<111>) ) ;
 assign wire7485* = ( (~ wire7485) ) ;
 assign C<107>* = ( (~ C<107>) ) ;
 assign wire7489* = ( (~ wire7489) ) ;
 assign key<243>* = ( (~ key<243>) ) ;
 assign wire7617* = ( (~ wire7617) ) ;
 assign C<106>* = ( (~ C<106>) ) ;
 assign wire7480* = ( (~ wire7480) ) ;
 assign key<251>* = ( (~ key<251>) ) ;
 assign wire7622* = ( (~ wire7622) ) ;
 assign C<105>* = ( (~ C<105>) ) ;
 assign wire7624* = ( (~ wire7624) ) ;
 assign key<194>* = ( (~ key<194>) ) ;
 assign wire7628* = ( (~ wire7628) ) ;
 assign C<104>* = ( (~ C<104>) ) ;
 assign wire7482* = ( (~ wire7482) ) ;
 assign key<202>* = ( (~ key<202>) ) ;
 assign wire7633* = ( (~ wire7633) ) ;
 assign C<103>* = ( (~ C<103>) ) ;
 assign wire7472* = ( (~ wire7472) ) ;
 assign key<210>* = ( (~ key<210>) ) ;
 assign wire7638* = ( (~ wire7638) ) ;
 assign C<102>* = ( (~ C<102>) ) ;
 assign wire7479* = ( (~ wire7479) ) ;
 assign key<218>* = ( (~ key<218>) ) ;
 assign wire7643* = ( (~ wire7643) ) ;
 assign C<101>* = ( (~ C<101>) ) ;
 assign wire7645* = ( (~ wire7645) ) ;
 assign key<226>* = ( (~ key<226>) ) ;
 assign wire7649* = ( (~ wire7649) ) ;
 assign C<100>* = ( (~ C<100>) ) ;
 assign wire7491* = ( (~ wire7491) ) ;
 assign key<234>* = ( (~ key<234>) ) ;
 assign wire7654* = ( (~ wire7654) ) ;
 assign C<99>* = ( (~ C<99>) ) ;
 assign wire7656* = ( (~ wire7656) ) ;
 assign key<242>* = ( (~ key<242>) ) ;
 assign wire7660* = ( (~ wire7660) ) ;
 assign C<98>* = ( (~ C<98>) ) ;
 assign wire7484* = ( (~ wire7484) ) ;
 assign key<250>* = ( (~ key<250>) ) ;
 assign wire7665* = ( (~ wire7665) ) ;
 assign C<97>* = ( (~ C<97>) ) ;
 assign wire7492* = ( (~ wire7492) ) ;
 assign key<193>* = ( (~ key<193>) ) ;
 assign wire7670* = ( (~ wire7670) ) ;
 assign C<96>* = ( (~ C<96>) ) ;
 assign wire7471* = ( (~ wire7471) ) ;
 assign key<201>* = ( (~ key<201>) ) ;
 assign wire7675* = ( (~ wire7675) ) ;
 assign C<95>* = ( (~ C<95>) ) ;
 assign wire7478* = ( (~ wire7478) ) ;
 assign key<209>* = ( (~ key<209>) ) ;
 assign wire7680* = ( (~ wire7680) ) ;
 assign C<94>* = ( (~ C<94>) ) ;
 assign wire7490* = ( (~ wire7490) ) ;
 assign key<217>* = ( (~ key<217>) ) ;
 assign wire7685* = ( (~ wire7685) ) ;
 assign C<93>* = ( (~ C<93>) ) ;
 assign wire7481* = ( (~ wire7481) ) ;
 assign key<225>* = ( (~ key<225>) ) ;
 assign wire7690* = ( (~ wire7690) ) ;
 assign C<92>* = ( (~ C<92>) ) ;
 assign wire7692* = ( (~ wire7692) ) ;
 assign key<233>* = ( (~ key<233>) ) ;
 assign wire7696* = ( (~ wire7696) ) ;
 assign C<91>* = ( (~ C<91>) ) ;
 assign wire7476* = ( (~ wire7476) ) ;
 assign key<241>* = ( (~ key<241>) ) ;
 assign wire7701* = ( (~ wire7701) ) ;
 assign C<90>* = ( (~ C<90>) ) ;
 assign wire7474* = ( (~ wire7474) ) ;
 assign key<249>* = ( (~ key<249>) ) ;
 assign wire7706* = ( (~ wire7706) ) ;
 assign C<89>* = ( (~ C<89>) ) ;
 assign wire7483* = ( (~ wire7483) ) ;
 assign key<192>* = ( (~ key<192>) ) ;
 assign wire7711* = ( (~ wire7711) ) ;
 assign C<88>* = ( (~ C<88>) ) ;
 assign wire7487* = ( (~ wire7487) ) ;
 assign key<200>* = ( (~ key<200>) ) ;
 assign wire7716* = ( (~ wire7716) ) ;
 assign C<87>* = ( (~ C<87>) ) ;
 assign wire7477* = ( (~ wire7477) ) ;
 assign key<208>* = ( (~ key<208>) ) ;
 assign wire7721* = ( (~ wire7721) ) ;
 assign C<86>* = ( (~ C<86>) ) ;
 assign wire7486* = ( (~ wire7486) ) ;
 assign key<216>* = ( (~ key<216>) ) ;
 assign wire7726* = ( (~ wire7726) ) ;
 assign C<85>* = ( (~ C<85>) ) ;
 assign wire7470* = ( (~ wire7470) ) ;
 assign key<224>* = ( (~ key<224>) ) ;
 assign wire7731* = ( (~ wire7731) ) ;
 assign C<84>* = ( (~ C<84>) ) ;
 assign wire7488* = ( (~ wire7488) ) ;
 assign key<232>* = ( (~ key<232>) ) ;
 assign wire7736* = ( (~ wire7736) ) ;
 assign C<83>* = ( (~ C<83>) ) ;
 assign wire7509* = ( (~ wire7509) ) ;
 assign key<240>* = ( (~ key<240>) ) ;
 assign wire7741* = ( (~ wire7741) ) ;
 assign C<82>* = ( (~ C<82>) ) ;
 assign wire7496* = ( (~ wire7496) ) ;
 assign key<248>* = ( (~ key<248>) ) ;
 assign wire7746* = ( (~ wire7746) ) ;
 assign C<81>* = ( (~ C<81>) ) ;
 assign wire7500* = ( (~ wire7500) ) ;
 assign key<163>* = ( (~ key<163>) ) ;
 assign wire7751* = ( (~ wire7751) ) ;
 assign C<80>* = ( (~ C<80>) ) ;
 assign wire7753* = ( (~ wire7753) ) ;
 assign key<171>* = ( (~ key<171>) ) ;
 assign wire7757* = ( (~ wire7757) ) ;
 assign C<79>* = ( (~ C<79>) ) ;
 assign wire7513* = ( (~ wire7513) ) ;
 assign key<179>* = ( (~ key<179>) ) ;
 assign wire7762* = ( (~ wire7762) ) ;
 assign C<78>* = ( (~ C<78>) ) ;
 assign wire7504* = ( (~ wire7504) ) ;
 assign key<187>* = ( (~ key<187>) ) ;
 assign wire7767* = ( (~ wire7767) ) ;
 assign C<77>* = ( (~ C<77>) ) ;
 assign wire7769* = ( (~ wire7769) ) ;
 assign key<130>* = ( (~ key<130>) ) ;
 assign wire7773* = ( (~ wire7773) ) ;
 assign C<76>* = ( (~ C<76>) ) ;
 assign wire7506* = ( (~ wire7506) ) ;
 assign key<138>* = ( (~ key<138>) ) ;
 assign wire7778* = ( (~ wire7778) ) ;
 assign C<75>* = ( (~ C<75>) ) ;
 assign wire7495* = ( (~ wire7495) ) ;
 assign key<146>* = ( (~ key<146>) ) ;
 assign wire7783* = ( (~ wire7783) ) ;
 assign C<74>* = ( (~ C<74>) ) ;
 assign wire7503* = ( (~ wire7503) ) ;
 assign key<154>* = ( (~ key<154>) ) ;
 assign wire7788* = ( (~ wire7788) ) ;
 assign C<73>* = ( (~ C<73>) ) ;
 assign wire7790* = ( (~ wire7790) ) ;
 assign key<162>* = ( (~ key<162>) ) ;
 assign wire7794* = ( (~ wire7794) ) ;
 assign C<72>* = ( (~ C<72>) ) ;
 assign wire7515* = ( (~ wire7515) ) ;
 assign key<170>* = ( (~ key<170>) ) ;
 assign wire7799* = ( (~ wire7799) ) ;
 assign C<71>* = ( (~ C<71>) ) ;
 assign wire7498* = ( (~ wire7498) ) ;
 assign key<178>* = ( (~ key<178>) ) ;
 assign wire7804* = ( (~ wire7804) ) ;
 assign C<70>* = ( (~ C<70>) ) ;
 assign wire7508* = ( (~ wire7508) ) ;
 assign key<186>* = ( (~ key<186>) ) ;
 assign wire7809* = ( (~ wire7809) ) ;
 assign C<69>* = ( (~ C<69>) ) ;
 assign wire7516* = ( (~ wire7516) ) ;
 assign key<129>* = ( (~ key<129>) ) ;
 assign wire7814* = ( (~ wire7814) ) ;
 assign C<68>* = ( (~ C<68>) ) ;
 assign wire7494* = ( (~ wire7494) ) ;
 assign key<137>* = ( (~ key<137>) ) ;
 assign wire7819* = ( (~ wire7819) ) ;
 assign C<67>* = ( (~ C<67>) ) ;
 assign wire7502* = ( (~ wire7502) ) ;
 assign key<145>* = ( (~ key<145>) ) ;
 assign wire7824* = ( (~ wire7824) ) ;
 assign C<66>* = ( (~ C<66>) ) ;
 assign wire7514* = ( (~ wire7514) ) ;
 assign key<153>* = ( (~ key<153>) ) ;
 assign wire7829* = ( (~ wire7829) ) ;
 assign C<65>* = ( (~ C<65>) ) ;
 assign wire7505* = ( (~ wire7505) ) ;
 assign key<161>* = ( (~ key<161>) ) ;
 assign wire7834* = ( (~ wire7834) ) ;
 assign C<64>* = ( (~ C<64>) ) ;
 assign wire7836* = ( (~ wire7836) ) ;
 assign key<169>* = ( (~ key<169>) ) ;
 assign wire7840* = ( (~ wire7840) ) ;
 assign C<63>* = ( (~ C<63>) ) ;
 assign wire7499* = ( (~ wire7499) ) ;
 assign key<177>* = ( (~ key<177>) ) ;
 assign wire7845* = ( (~ wire7845) ) ;
 assign C<62>* = ( (~ C<62>) ) ;
 assign wire7497* = ( (~ wire7497) ) ;
 assign key<185>* = ( (~ key<185>) ) ;
 assign wire7850* = ( (~ wire7850) ) ;
 assign C<61>* = ( (~ C<61>) ) ;
 assign wire7507* = ( (~ wire7507) ) ;
 assign key<128>* = ( (~ key<128>) ) ;
 assign wire7855* = ( (~ wire7855) ) ;
 assign C<60>* = ( (~ C<60>) ) ;
 assign wire7511* = ( (~ wire7511) ) ;
 assign key<136>* = ( (~ key<136>) ) ;
 assign wire7860* = ( (~ wire7860) ) ;
 assign C<59>* = ( (~ C<59>) ) ;
 assign wire7501* = ( (~ wire7501) ) ;
 assign key<144>* = ( (~ key<144>) ) ;
 assign wire7865* = ( (~ wire7865) ) ;
 assign C<58>* = ( (~ C<58>) ) ;
 assign wire7510* = ( (~ wire7510) ) ;
 assign key<152>* = ( (~ key<152>) ) ;
 assign wire7870* = ( (~ wire7870) ) ;
 assign C<57>* = ( (~ C<57>) ) ;
 assign wire7493* = ( (~ wire7493) ) ;
 assign key<160>* = ( (~ key<160>) ) ;
 assign wire7875* = ( (~ wire7875) ) ;
 assign C<56>* = ( (~ C<56>) ) ;
 assign wire7512* = ( (~ wire7512) ) ;
 assign key<168>* = ( (~ key<168>) ) ;
 assign wire7880* = ( (~ wire7880) ) ;
 assign C<55>* = ( (~ C<55>) ) ;
 assign wire7533* = ( (~ wire7533) ) ;
 assign key<176>* = ( (~ key<176>) ) ;
 assign wire7885* = ( (~ wire7885) ) ;
 assign C<54>* = ( (~ C<54>) ) ;
 assign wire7520* = ( (~ wire7520) ) ;
 assign key<184>* = ( (~ key<184>) ) ;
 assign wire7890* = ( (~ wire7890) ) ;
 assign C<53>* = ( (~ C<53>) ) ;
 assign wire7524* = ( (~ wire7524) ) ;
 assign key<99>* = ( (~ key<99>) ) ;
 assign wire7895* = ( (~ wire7895) ) ;
 assign C<52>* = ( (~ C<52>) ) ;
 assign wire7897* = ( (~ wire7897) ) ;
 assign key<107>* = ( (~ key<107>) ) ;
 assign wire7901* = ( (~ wire7901) ) ;
 assign C<51>* = ( (~ C<51>) ) ;
 assign wire7537* = ( (~ wire7537) ) ;
 assign key<115>* = ( (~ key<115>) ) ;
 assign wire7906* = ( (~ wire7906) ) ;
 assign C<50>* = ( (~ C<50>) ) ;
 assign wire7528* = ( (~ wire7528) ) ;
 assign key<123>* = ( (~ key<123>) ) ;
 assign wire7911* = ( (~ wire7911) ) ;
 assign C<49>* = ( (~ C<49>) ) ;
 assign wire7913* = ( (~ wire7913) ) ;
 assign key<66>* = ( (~ key<66>) ) ;
 assign wire7917* = ( (~ wire7917) ) ;
 assign C<48>* = ( (~ C<48>) ) ;
 assign wire7530* = ( (~ wire7530) ) ;
 assign key<74>* = ( (~ key<74>) ) ;
 assign wire7922* = ( (~ wire7922) ) ;
 assign C<47>* = ( (~ C<47>) ) ;
 assign wire7519* = ( (~ wire7519) ) ;
 assign key<82>* = ( (~ key<82>) ) ;
 assign wire7927* = ( (~ wire7927) ) ;
 assign C<46>* = ( (~ C<46>) ) ;
 assign wire7527* = ( (~ wire7527) ) ;
 assign key<90>* = ( (~ key<90>) ) ;
 assign wire7932* = ( (~ wire7932) ) ;
 assign C<45>* = ( (~ C<45>) ) ;
 assign wire7934* = ( (~ wire7934) ) ;
 assign key<98>* = ( (~ key<98>) ) ;
 assign wire7938* = ( (~ wire7938) ) ;
 assign C<44>* = ( (~ C<44>) ) ;
 assign wire7539* = ( (~ wire7539) ) ;
 assign key<106>* = ( (~ key<106>) ) ;
 assign wire7943* = ( (~ wire7943) ) ;
 assign C<43>* = ( (~ C<43>) ) ;
 assign wire7522* = ( (~ wire7522) ) ;
 assign key<114>* = ( (~ key<114>) ) ;
 assign wire7948* = ( (~ wire7948) ) ;
 assign C<42>* = ( (~ C<42>) ) ;
 assign wire7532* = ( (~ wire7532) ) ;
 assign key<122>* = ( (~ key<122>) ) ;
 assign wire7953* = ( (~ wire7953) ) ;
 assign C<41>* = ( (~ C<41>) ) ;
 assign wire7540* = ( (~ wire7540) ) ;
 assign key<65>* = ( (~ key<65>) ) ;
 assign wire7958* = ( (~ wire7958) ) ;
 assign C<40>* = ( (~ C<40>) ) ;
 assign wire7518* = ( (~ wire7518) ) ;
 assign key<73>* = ( (~ key<73>) ) ;
 assign wire7963* = ( (~ wire7963) ) ;
 assign C<39>* = ( (~ C<39>) ) ;
 assign wire7526* = ( (~ wire7526) ) ;
 assign key<81>* = ( (~ key<81>) ) ;
 assign wire7968* = ( (~ wire7968) ) ;
 assign C<38>* = ( (~ C<38>) ) ;
 assign wire7538* = ( (~ wire7538) ) ;
 assign key<89>* = ( (~ key<89>) ) ;
 assign wire7973* = ( (~ wire7973) ) ;
 assign C<37>* = ( (~ C<37>) ) ;
 assign wire7529* = ( (~ wire7529) ) ;
 assign key<97>* = ( (~ key<97>) ) ;
 assign wire7978* = ( (~ wire7978) ) ;
 assign C<36>* = ( (~ C<36>) ) ;
 assign wire7980* = ( (~ wire7980) ) ;
 assign key<105>* = ( (~ key<105>) ) ;
 assign wire7984* = ( (~ wire7984) ) ;
 assign C<35>* = ( (~ C<35>) ) ;
 assign wire7523* = ( (~ wire7523) ) ;
 assign key<113>* = ( (~ key<113>) ) ;
 assign wire7989* = ( (~ wire7989) ) ;
 assign C<34>* = ( (~ C<34>) ) ;
 assign wire7521* = ( (~ wire7521) ) ;
 assign key<121>* = ( (~ key<121>) ) ;
 assign wire7994* = ( (~ wire7994) ) ;
 assign C<33>* = ( (~ C<33>) ) ;
 assign wire7531* = ( (~ wire7531) ) ;
 assign key<64>* = ( (~ key<64>) ) ;
 assign wire7999* = ( (~ wire7999) ) ;
 assign C<32>* = ( (~ C<32>) ) ;
 assign wire7535* = ( (~ wire7535) ) ;
 assign key<72>* = ( (~ key<72>) ) ;
 assign wire8004* = ( (~ wire8004) ) ;
 assign C<31>* = ( (~ C<31>) ) ;
 assign wire7525* = ( (~ wire7525) ) ;
 assign key<80>* = ( (~ key<80>) ) ;
 assign wire8009* = ( (~ wire8009) ) ;
 assign C<30>* = ( (~ C<30>) ) ;
 assign wire7534* = ( (~ wire7534) ) ;
 assign key<88>* = ( (~ key<88>) ) ;
 assign wire8014* = ( (~ wire8014) ) ;
 assign C<29>* = ( (~ C<29>) ) ;
 assign wire7517* = ( (~ wire7517) ) ;
 assign key<96>* = ( (~ key<96>) ) ;
 assign wire8019* = ( (~ wire8019) ) ;
 assign C<28>* = ( (~ C<28>) ) ;
 assign wire7536* = ( (~ wire7536) ) ;
 assign key<104>* = ( (~ key<104>) ) ;
 assign wire8024* = ( (~ wire8024) ) ;
 assign C<27>* = ( (~ C<27>) ) ;
 assign wire7557* = ( (~ wire7557) ) ;
 assign key<112>* = ( (~ key<112>) ) ;
 assign wire8029* = ( (~ wire8029) ) ;
 assign C<26>* = ( (~ C<26>) ) ;
 assign wire7544* = ( (~ wire7544) ) ;
 assign key<120>* = ( (~ key<120>) ) ;
 assign wire8034* = ( (~ wire8034) ) ;
 assign C<25>* = ( (~ C<25>) ) ;
 assign wire7548* = ( (~ wire7548) ) ;
 assign key<35>* = ( (~ key<35>) ) ;
 assign wire8039* = ( (~ wire8039) ) ;
 assign C<24>* = ( (~ C<24>) ) ;
 assign wire8041* = ( (~ wire8041) ) ;
 assign key<43>* = ( (~ key<43>) ) ;
 assign wire8045* = ( (~ wire8045) ) ;
 assign C<23>* = ( (~ C<23>) ) ;
 assign wire7561* = ( (~ wire7561) ) ;
 assign key<51>* = ( (~ key<51>) ) ;
 assign wire8050* = ( (~ wire8050) ) ;
 assign C<22>* = ( (~ C<22>) ) ;
 assign wire7552* = ( (~ wire7552) ) ;
 assign key<59>* = ( (~ key<59>) ) ;
 assign wire8055* = ( (~ wire8055) ) ;
 assign C<21>* = ( (~ C<21>) ) ;
 assign wire8057* = ( (~ wire8057) ) ;
 assign key<2>* = ( (~ key<2>) ) ;
 assign wire8061* = ( (~ wire8061) ) ;
 assign C<20>* = ( (~ C<20>) ) ;
 assign wire7554* = ( (~ wire7554) ) ;
 assign key<10>* = ( (~ key<10>) ) ;
 assign wire8066* = ( (~ wire8066) ) ;
 assign C<19>* = ( (~ C<19>) ) ;
 assign wire7543* = ( (~ wire7543) ) ;
 assign key<18>* = ( (~ key<18>) ) ;
 assign wire8071* = ( (~ wire8071) ) ;
 assign C<18>* = ( (~ C<18>) ) ;
 assign wire7551* = ( (~ wire7551) ) ;
 assign key<26>* = ( (~ key<26>) ) ;
 assign wire8076* = ( (~ wire8076) ) ;
 assign C<17>* = ( (~ C<17>) ) ;
 assign wire8078* = ( (~ wire8078) ) ;
 assign key<34>* = ( (~ key<34>) ) ;
 assign wire8082* = ( (~ wire8082) ) ;
 assign C<16>* = ( (~ C<16>) ) ;
 assign wire7563* = ( (~ wire7563) ) ;
 assign key<42>* = ( (~ key<42>) ) ;
 assign wire8087* = ( (~ wire8087) ) ;
 assign C<15>* = ( (~ C<15>) ) ;
 assign wire7546* = ( (~ wire7546) ) ;
 assign key<50>* = ( (~ key<50>) ) ;
 assign wire8092* = ( (~ wire8092) ) ;
 assign C<14>* = ( (~ C<14>) ) ;
 assign wire7556* = ( (~ wire7556) ) ;
 assign key<58>* = ( (~ key<58>) ) ;
 assign wire8097* = ( (~ wire8097) ) ;
 assign C<13>* = ( (~ C<13>) ) ;
 assign wire7564* = ( (~ wire7564) ) ;
 assign key<1>* = ( (~ key<1>) ) ;
 assign wire8102* = ( (~ wire8102) ) ;
 assign C<12>* = ( (~ C<12>) ) ;
 assign wire7542* = ( (~ wire7542) ) ;
 assign key<9>* = ( (~ key<9>) ) ;
 assign wire8107* = ( (~ wire8107) ) ;
 assign C<11>* = ( (~ C<11>) ) ;
 assign wire7550* = ( (~ wire7550) ) ;
 assign key<17>* = ( (~ key<17>) ) ;
 assign wire8112* = ( (~ wire8112) ) ;
 assign C<10>* = ( (~ C<10>) ) ;
 assign wire7562* = ( (~ wire7562) ) ;
 assign key<25>* = ( (~ key<25>) ) ;
 assign wire8117* = ( (~ wire8117) ) ;
 assign C<9>* = ( (~ C<9>) ) ;
 assign wire7553* = ( (~ wire7553) ) ;
 assign key<33>* = ( (~ key<33>) ) ;
 assign wire8122* = ( (~ wire8122) ) ;
 assign C<8>* = ( (~ C<8>) ) ;
 assign wire8124* = ( (~ wire8124) ) ;
 assign key<41>* = ( (~ key<41>) ) ;
 assign wire8128* = ( (~ wire8128) ) ;
 assign C<7>* = ( (~ C<7>) ) ;
 assign wire7547* = ( (~ wire7547) ) ;
 assign key<49>* = ( (~ key<49>) ) ;
 assign wire8133* = ( (~ wire8133) ) ;
 assign C<6>* = ( (~ C<6>) ) ;
 assign wire7545* = ( (~ wire7545) ) ;
 assign key<57>* = ( (~ key<57>) ) ;
 assign wire8138* = ( (~ wire8138) ) ;
 assign C<5>* = ( (~ C<5>) ) ;
 assign wire7555* = ( (~ wire7555) ) ;
 assign key<0>* = ( (~ key<0>) ) ;
 assign wire8143* = ( (~ wire8143) ) ;
 assign C<4>* = ( (~ C<4>) ) ;
 assign wire7559* = ( (~ wire7559) ) ;
 assign key<8>* = ( (~ key<8>) ) ;
 assign wire8148* = ( (~ wire8148) ) ;
 assign C<3>* = ( (~ C<3>) ) ;
 assign wire7549* = ( (~ wire7549) ) ;
 assign key<16>* = ( (~ key<16>) ) ;
 assign wire8153* = ( (~ wire8153) ) ;
 assign C<2>* = ( (~ C<2>) ) ;
 assign wire7558* = ( (~ wire7558) ) ;
 assign key<24>* = ( (~ key<24>) ) ;
 assign wire8158* = ( (~ wire8158) ) ;
 assign key<32>* = ( (~ key<32>) ) ;
 assign wire8163* = ( (~ wire8163) ) ;
 assign key<40>* = ( (~ key<40>) ) ;
 assign wire8168* = ( (~ wire8168) ) ;
 assign key<48>* = ( (~ key<48>) ) ;
 assign wire8173* = ( (~ wire8173) ) ;
 assign D<1>* = ( (~ D<1>) ) ;
 assign wire7463* = ( (~ wire7463) ) ;
 assign D<109>* = ( (~ D<109>) ) ;
 assign D<110>* = ( (~ D<110>) ) ;
 assign wire8179* = ( (~ wire8179) ) ;
 assign wire7394* = ( (~ wire7394) ) ;
 assign key<195>* = ( (~ key<195>) ) ;
 assign wire8184* = ( (~ wire8184) ) ;
 assign D<0>* = ( (~ D<0>) ) ;
 assign key<62>* = ( (~ key<62>) ) ;
 assign wire7447* = ( (~ wire7447) ) ;
 assign wire8182* = ( (~ wire8182) ) ;
 assign D<108>* = ( (~ D<108>) ) ;
 assign wire7382* = ( (~ wire7382) ) ;
 assign key<203>* = ( (~ key<203>) ) ;
 assign wire8189* = ( (~ wire8189) ) ;
 assign D<111>* = ( (~ D<111>) ) ;
 assign wire7384* = ( (~ wire7384) ) ;
 assign D<107>* = ( (~ D<107>) ) ;
 assign wire7398* = ( (~ wire7398) ) ;
 assign key<211>* = ( (~ key<211>) ) ;
 assign wire8194* = ( (~ wire8194) ) ;
 assign D<106>* = ( (~ D<106>) ) ;
 assign wire7391* = ( (~ wire7391) ) ;
 assign key<219>* = ( (~ key<219>) ) ;
 assign wire8199* = ( (~ wire8199) ) ;
 assign D<105>* = ( (~ D<105>) ) ;
 assign wire7380* = ( (~ wire7380) ) ;
 assign key<196>* = ( (~ key<196>) ) ;
 assign wire8204* = ( (~ wire8204) ) ;
 assign D<104>* = ( (~ D<104>) ) ;
 assign wire7386* = ( (~ wire7386) ) ;
 assign key<204>* = ( (~ key<204>) ) ;
 assign wire8209* = ( (~ wire8209) ) ;
 assign D<103>* = ( (~ D<103>) ) ;
 assign wire7388* = ( (~ wire7388) ) ;
 assign key<212>* = ( (~ key<212>) ) ;
 assign wire8214* = ( (~ wire8214) ) ;
 assign D<102>* = ( (~ D<102>) ) ;
 assign wire7395* = ( (~ wire7395) ) ;
 assign key<220>* = ( (~ key<220>) ) ;
 assign wire8219* = ( (~ wire8219) ) ;
 assign D<101>* = ( (~ D<101>) ) ;
 assign wire7381* = ( (~ wire7381) ) ;
 assign key<228>* = ( (~ key<228>) ) ;
 assign wire8224* = ( (~ wire8224) ) ;
 assign D<100>* = ( (~ D<100>) ) ;
 assign wire7390* = ( (~ wire7390) ) ;
 assign key<172>* = ( (~ key<172>) ) ;
 assign wire8229* = ( (~ wire8229) ) ;
 assign D<99>* = ( (~ D<99>) ) ;
 assign wire7387* = ( (~ wire7387) ) ;
 assign key<244>* = ( (~ key<244>) ) ;
 assign wire8234* = ( (~ wire8234) ) ;
 assign D<98>* = ( (~ D<98>) ) ;
 assign wire8236* = ( (~ wire8236) ) ;
 assign key<252>* = ( (~ key<252>) ) ;
 assign wire8240* = ( (~ wire8240) ) ;
 assign D<97>* = ( (~ D<97>) ) ;
 assign wire8242* = ( (~ wire8242) ) ;
 assign key<197>* = ( (~ key<197>) ) ;
 assign wire8246* = ( (~ wire8246) ) ;
 assign D<96>* = ( (~ D<96>) ) ;
 assign wire8248* = ( (~ wire8248) ) ;
 assign key<205>* = ( (~ key<205>) ) ;
 assign wire8252* = ( (~ wire8252) ) ;
 assign D<95>* = ( (~ D<95>) ) ;
 assign wire7392* = ( (~ wire7392) ) ;
 assign key<213>* = ( (~ key<213>) ) ;
 assign wire8257* = ( (~ wire8257) ) ;
 assign D<94>* = ( (~ D<94>) ) ;
 assign wire7385* = ( (~ wire7385) ) ;
 assign key<221>* = ( (~ key<221>) ) ;
 assign wire8262* = ( (~ wire8262) ) ;
 assign D<93>* = ( (~ D<93>) ) ;
 assign wire8264* = ( (~ wire8264) ) ;
 assign key<229>* = ( (~ key<229>) ) ;
 assign wire8268* = ( (~ wire8268) ) ;
 assign D<92>* = ( (~ D<92>) ) ;
 assign wire7396* = ( (~ wire7396) ) ;
 assign key<237>* = ( (~ key<237>) ) ;
 assign wire8273* = ( (~ wire8273) ) ;
 assign D<91>* = ( (~ D<91>) ) ;
 assign wire7379* = ( (~ wire7379) ) ;
 assign key<245>* = ( (~ key<245>) ) ;
 assign wire8278* = ( (~ wire8278) ) ;
 assign D<90>* = ( (~ D<90>) ) ;
 assign wire8280* = ( (~ wire8280) ) ;
 assign key<253>* = ( (~ key<253>) ) ;
 assign wire8284* = ( (~ wire8284) ) ;
 assign D<89>* = ( (~ D<89>) ) ;
 assign wire7383* = ( (~ wire7383) ) ;
 assign key<198>* = ( (~ key<198>) ) ;
 assign wire8289* = ( (~ wire8289) ) ;
 assign D<88>* = ( (~ D<88>) ) ;
 assign wire7389* = ( (~ wire7389) ) ;
 assign key<206>* = ( (~ key<206>) ) ;
 assign wire8294* = ( (~ wire8294) ) ;
 assign D<87>* = ( (~ D<87>) ) ;
 assign wire7377* = ( (~ wire7377) ) ;
 assign key<214>* = ( (~ key<214>) ) ;
 assign wire8299* = ( (~ wire8299) ) ;
 assign D<86>* = ( (~ D<86>) ) ;
 assign wire7397* = ( (~ wire7397) ) ;
 assign key<222>* = ( (~ key<222>) ) ;
 assign wire8304* = ( (~ wire8304) ) ;
 assign D<85>* = ( (~ D<85>) ) ;
 assign wire7393* = ( (~ wire7393) ) ;
 assign key<230>* = ( (~ key<230>) ) ;
 assign wire8309* = ( (~ wire8309) ) ;
 assign D<84>* = ( (~ D<84>) ) ;
 assign wire7378* = ( (~ wire7378) ) ;
 assign key<238>* = ( (~ key<238>) ) ;
 assign wire8314* = ( (~ wire8314) ) ;
 assign D<83>* = ( (~ D<83>) ) ;
 assign wire7407* = ( (~ wire7407) ) ;
 assign key<246>* = ( (~ key<246>) ) ;
 assign wire8319* = ( (~ wire8319) ) ;
 assign D<82>* = ( (~ D<82>) ) ;
 assign wire7417* = ( (~ wire7417) ) ;
 assign key<254>* = ( (~ key<254>) ) ;
 assign wire8324* = ( (~ wire8324) ) ;
 assign D<81>* = ( (~ D<81>) ) ;
 assign wire8326* = ( (~ wire8326) ) ;
 assign key<131>* = ( (~ key<131>) ) ;
 assign wire8330* = ( (~ wire8330) ) ;
 assign D<80>* = ( (~ D<80>) ) ;
 assign wire7405* = ( (~ wire7405) ) ;
 assign key<139>* = ( (~ key<139>) ) ;
 assign wire8335* = ( (~ wire8335) ) ;
 assign D<79>* = ( (~ D<79>) ) ;
 assign wire7421* = ( (~ wire7421) ) ;
 assign key<147>* = ( (~ key<147>) ) ;
 assign wire8340* = ( (~ wire8340) ) ;
 assign D<78>* = ( (~ D<78>) ) ;
 assign wire7414* = ( (~ wire7414) ) ;
 assign key<155>* = ( (~ key<155>) ) ;
 assign wire8345* = ( (~ wire8345) ) ;
 assign D<77>* = ( (~ D<77>) ) ;
 assign wire7402* = ( (~ wire7402) ) ;
 assign key<132>* = ( (~ key<132>) ) ;
 assign wire8350* = ( (~ wire8350) ) ;
 assign D<76>* = ( (~ D<76>) ) ;
 assign wire7409* = ( (~ wire7409) ) ;
 assign key<140>* = ( (~ key<140>) ) ;
 assign wire8355* = ( (~ wire8355) ) ;
 assign D<75>* = ( (~ D<75>) ) ;
 assign wire7411* = ( (~ wire7411) ) ;
 assign key<148>* = ( (~ key<148>) ) ;
 assign wire8360* = ( (~ wire8360) ) ;
 assign D<74>* = ( (~ D<74>) ) ;
 assign wire7418* = ( (~ wire7418) ) ;
 assign key<156>* = ( (~ key<156>) ) ;
 assign wire8365* = ( (~ wire8365) ) ;
 assign D<73>* = ( (~ D<73>) ) ;
 assign wire7404* = ( (~ wire7404) ) ;
 assign key<164>* = ( (~ key<164>) ) ;
 assign wire8370* = ( (~ wire8370) ) ;
 assign D<72>* = ( (~ D<72>) ) ;
 assign wire8372* = ( (~ wire8372) ) ;
 assign D<71>* = ( (~ D<71>) ) ;
 assign wire7410* = ( (~ wire7410) ) ;
 assign key<180>* = ( (~ key<180>) ) ;
 assign wire8380* = ( (~ wire8380) ) ;
 assign D<70>* = ( (~ D<70>) ) ;
 assign wire7413* = ( (~ wire7413) ) ;
 assign key<188>* = ( (~ key<188>) ) ;
 assign wire8385* = ( (~ wire8385) ) ;
 assign D<69>* = ( (~ D<69>) ) ;
 assign wire7403* = ( (~ wire7403) ) ;
 assign key<133>* = ( (~ key<133>) ) ;
 assign wire8390* = ( (~ wire8390) ) ;
 assign D<68>* = ( (~ D<68>) ) ;
 assign wire7422* = ( (~ wire7422) ) ;
 assign key<141>* = ( (~ key<141>) ) ;
 assign wire8395* = ( (~ wire8395) ) ;
 assign D<67>* = ( (~ D<67>) ) ;
 assign wire7415* = ( (~ wire7415) ) ;
 assign key<149>* = ( (~ key<149>) ) ;
 assign wire8400* = ( (~ wire8400) ) ;
 assign D<66>* = ( (~ D<66>) ) ;
 assign wire7408* = ( (~ wire7408) ) ;
 assign key<157>* = ( (~ key<157>) ) ;
 assign wire8405* = ( (~ wire8405) ) ;
 assign D<65>* = ( (~ D<65>) ) ;
 assign wire8407* = ( (~ wire8407) ) ;
 assign key<165>* = ( (~ key<165>) ) ;
 assign wire8411* = ( (~ wire8411) ) ;
 assign D<64>* = ( (~ D<64>) ) ;
 assign wire7419* = ( (~ wire7419) ) ;
 assign key<173>* = ( (~ key<173>) ) ;
 assign wire8416* = ( (~ wire8416) ) ;
 assign D<63>* = ( (~ D<63>) ) ;
 assign wire7401* = ( (~ wire7401) ) ;
 assign key<181>* = ( (~ key<181>) ) ;
 assign wire8421* = ( (~ wire8421) ) ;
 assign D<62>* = ( (~ D<62>) ) ;
 assign wire8423* = ( (~ wire8423) ) ;
 assign key<189>* = ( (~ key<189>) ) ;
 assign wire8427* = ( (~ wire8427) ) ;
 assign D<61>* = ( (~ D<61>) ) ;
 assign wire7406* = ( (~ wire7406) ) ;
 assign key<134>* = ( (~ key<134>) ) ;
 assign wire8432* = ( (~ wire8432) ) ;
 assign D<60>* = ( (~ D<60>) ) ;
 assign wire7412* = ( (~ wire7412) ) ;
 assign key<142>* = ( (~ key<142>) ) ;
 assign wire8437* = ( (~ wire8437) ) ;
 assign D<59>* = ( (~ D<59>) ) ;
 assign wire7399* = ( (~ wire7399) ) ;
 assign key<150>* = ( (~ key<150>) ) ;
 assign wire8442* = ( (~ wire8442) ) ;
 assign D<58>* = ( (~ D<58>) ) ;
 assign wire7420* = ( (~ wire7420) ) ;
 assign key<158>* = ( (~ key<158>) ) ;
 assign wire8447* = ( (~ wire8447) ) ;
 assign D<57>* = ( (~ D<57>) ) ;
 assign wire7416* = ( (~ wire7416) ) ;
 assign key<166>* = ( (~ key<166>) ) ;
 assign wire8452* = ( (~ wire8452) ) ;
 assign D<56>* = ( (~ D<56>) ) ;
 assign wire7400* = ( (~ wire7400) ) ;
 assign key<174>* = ( (~ key<174>) ) ;
 assign wire8457* = ( (~ wire8457) ) ;
 assign D<55>* = ( (~ D<55>) ) ;
 assign wire7430* = ( (~ wire7430) ) ;
 assign key<182>* = ( (~ key<182>) ) ;
 assign wire8462* = ( (~ wire8462) ) ;
 assign D<54>* = ( (~ D<54>) ) ;
 assign wire7440* = ( (~ wire7440) ) ;
 assign key<190>* = ( (~ key<190>) ) ;
 assign wire8467* = ( (~ wire8467) ) ;
 assign D<53>* = ( (~ D<53>) ) ;
 assign wire8469* = ( (~ wire8469) ) ;
 assign key<67>* = ( (~ key<67>) ) ;
 assign wire8473* = ( (~ wire8473) ) ;
 assign D<52>* = ( (~ D<52>) ) ;
 assign wire7428* = ( (~ wire7428) ) ;
 assign key<75>* = ( (~ key<75>) ) ;
 assign wire8478* = ( (~ wire8478) ) ;
 assign D<51>* = ( (~ D<51>) ) ;
 assign wire7444* = ( (~ wire7444) ) ;
 assign key<83>* = ( (~ key<83>) ) ;
 assign wire8483* = ( (~ wire8483) ) ;
 assign D<50>* = ( (~ D<50>) ) ;
 assign wire7437* = ( (~ wire7437) ) ;
 assign key<91>* = ( (~ key<91>) ) ;
 assign wire8488* = ( (~ wire8488) ) ;
 assign D<49>* = ( (~ D<49>) ) ;
 assign wire7426* = ( (~ wire7426) ) ;
 assign key<68>* = ( (~ key<68>) ) ;
 assign wire8493* = ( (~ wire8493) ) ;
 assign D<48>* = ( (~ D<48>) ) ;
 assign wire7432* = ( (~ wire7432) ) ;
 assign key<76>* = ( (~ key<76>) ) ;
 assign wire8498* = ( (~ wire8498) ) ;
 assign D<47>* = ( (~ D<47>) ) ;
 assign wire7434* = ( (~ wire7434) ) ;
 assign key<84>* = ( (~ key<84>) ) ;
 assign wire8503* = ( (~ wire8503) ) ;
 assign D<46>* = ( (~ D<46>) ) ;
 assign wire7441* = ( (~ wire7441) ) ;
 assign key<92>* = ( (~ key<92>) ) ;
 assign wire8508* = ( (~ wire8508) ) ;
 assign D<45>* = ( (~ D<45>) ) ;
 assign wire7427* = ( (~ wire7427) ) ;
 assign key<100>* = ( (~ key<100>) ) ;
 assign wire8513* = ( (~ wire8513) ) ;
 assign D<44>* = ( (~ D<44>) ) ;
 assign wire7436* = ( (~ wire7436) ) ;
 assign key<44>* = ( (~ key<44>) ) ;
 assign wire8518* = ( (~ wire8518) ) ;
 assign D<43>* = ( (~ D<43>) ) ;
 assign wire7433* = ( (~ wire7433) ) ;
 assign key<116>* = ( (~ key<116>) ) ;
 assign wire8523* = ( (~ wire8523) ) ;
 assign D<42>* = ( (~ D<42>) ) ;
 assign wire8525* = ( (~ wire8525) ) ;
 assign key<124>* = ( (~ key<124>) ) ;
 assign wire8529* = ( (~ wire8529) ) ;
 assign D<41>* = ( (~ D<41>) ) ;
 assign wire8531* = ( (~ wire8531) ) ;
 assign key<69>* = ( (~ key<69>) ) ;
 assign wire8535* = ( (~ wire8535) ) ;
 assign D<40>* = ( (~ D<40>) ) ;
 assign wire7445* = ( (~ wire7445) ) ;
 assign key<77>* = ( (~ key<77>) ) ;
 assign wire8540* = ( (~ wire8540) ) ;
 assign D<39>* = ( (~ D<39>) ) ;
 assign wire7438* = ( (~ wire7438) ) ;
 assign key<85>* = ( (~ key<85>) ) ;
 assign wire8545* = ( (~ wire8545) ) ;
 assign D<38>* = ( (~ D<38>) ) ;
 assign wire7431* = ( (~ wire7431) ) ;
 assign key<93>* = ( (~ key<93>) ) ;
 assign wire8550* = ( (~ wire8550) ) ;
 assign D<37>* = ( (~ D<37>) ) ;
 assign wire8552* = ( (~ wire8552) ) ;
 assign key<101>* = ( (~ key<101>) ) ;
 assign wire8556* = ( (~ wire8556) ) ;
 assign D<36>* = ( (~ D<36>) ) ;
 assign wire7442* = ( (~ wire7442) ) ;
 assign key<109>* = ( (~ key<109>) ) ;
 assign wire8561* = ( (~ wire8561) ) ;
 assign D<35>* = ( (~ D<35>) ) ;
 assign wire7425* = ( (~ wire7425) ) ;
 assign key<117>* = ( (~ key<117>) ) ;
 assign wire8566* = ( (~ wire8566) ) ;
 assign D<34>* = ( (~ D<34>) ) ;
 assign wire8568* = ( (~ wire8568) ) ;
 assign key<125>* = ( (~ key<125>) ) ;
 assign wire8572* = ( (~ wire8572) ) ;
 assign D<33>* = ( (~ D<33>) ) ;
 assign wire7429* = ( (~ wire7429) ) ;
 assign key<70>* = ( (~ key<70>) ) ;
 assign wire8577* = ( (~ wire8577) ) ;
 assign D<32>* = ( (~ D<32>) ) ;
 assign wire7435* = ( (~ wire7435) ) ;
 assign key<78>* = ( (~ key<78>) ) ;
 assign wire8582* = ( (~ wire8582) ) ;
 assign D<31>* = ( (~ D<31>) ) ;
 assign wire7423* = ( (~ wire7423) ) ;
 assign key<86>* = ( (~ key<86>) ) ;
 assign wire8587* = ( (~ wire8587) ) ;
 assign D<30>* = ( (~ D<30>) ) ;
 assign wire7443* = ( (~ wire7443) ) ;
 assign key<94>* = ( (~ key<94>) ) ;
 assign wire8592* = ( (~ wire8592) ) ;
 assign D<29>* = ( (~ D<29>) ) ;
 assign wire7439* = ( (~ wire7439) ) ;
 assign key<102>* = ( (~ key<102>) ) ;
 assign wire8597* = ( (~ wire8597) ) ;
 assign D<28>* = ( (~ D<28>) ) ;
 assign wire7424* = ( (~ wire7424) ) ;
 assign key<110>* = ( (~ key<110>) ) ;
 assign wire8602* = ( (~ wire8602) ) ;
 assign D<27>* = ( (~ D<27>) ) ;
 assign wire7454* = ( (~ wire7454) ) ;
 assign key<118>* = ( (~ key<118>) ) ;
 assign wire8607* = ( (~ wire8607) ) ;
 assign D<26>* = ( (~ D<26>) ) ;
 assign wire7464* = ( (~ wire7464) ) ;
 assign key<126>* = ( (~ key<126>) ) ;
 assign wire8612* = ( (~ wire8612) ) ;
 assign D<25>* = ( (~ D<25>) ) ;
 assign wire8614* = ( (~ wire8614) ) ;
 assign key<3>* = ( (~ key<3>) ) ;
 assign wire8618* = ( (~ wire8618) ) ;
 assign D<24>* = ( (~ D<24>) ) ;
 assign wire7452* = ( (~ wire7452) ) ;
 assign key<11>* = ( (~ key<11>) ) ;
 assign wire8623* = ( (~ wire8623) ) ;
 assign D<23>* = ( (~ D<23>) ) ;
 assign wire7468* = ( (~ wire7468) ) ;
 assign key<19>* = ( (~ key<19>) ) ;
 assign wire8628* = ( (~ wire8628) ) ;
 assign D<22>* = ( (~ D<22>) ) ;
 assign wire7461* = ( (~ wire7461) ) ;
 assign key<27>* = ( (~ key<27>) ) ;
 assign wire8633* = ( (~ wire8633) ) ;
 assign D<21>* = ( (~ D<21>) ) ;
 assign wire7449* = ( (~ wire7449) ) ;
 assign key<4>* = ( (~ key<4>) ) ;
 assign wire8638* = ( (~ wire8638) ) ;
 assign D<20>* = ( (~ D<20>) ) ;
 assign wire7456* = ( (~ wire7456) ) ;
 assign key<12>* = ( (~ key<12>) ) ;
 assign wire8643* = ( (~ wire8643) ) ;
 assign D<19>* = ( (~ D<19>) ) ;
 assign wire7458* = ( (~ wire7458) ) ;
 assign key<20>* = ( (~ key<20>) ) ;
 assign wire8648* = ( (~ wire8648) ) ;
 assign D<18>* = ( (~ D<18>) ) ;
 assign wire7465* = ( (~ wire7465) ) ;
 assign key<28>* = ( (~ key<28>) ) ;
 assign wire8653* = ( (~ wire8653) ) ;
 assign D<17>* = ( (~ D<17>) ) ;
 assign wire7451* = ( (~ wire7451) ) ;
 assign key<36>* = ( (~ key<36>) ) ;
 assign wire8658* = ( (~ wire8658) ) ;
 assign D<16>* = ( (~ D<16>) ) ;
 assign wire7460* = ( (~ wire7460) ) ;
 assign D<15>* = ( (~ D<15>) ) ;
 assign wire7457* = ( (~ wire7457) ) ;
 assign key<52>* = ( (~ key<52>) ) ;
 assign wire8667* = ( (~ wire8667) ) ;
 assign D<14>* = ( (~ D<14>) ) ;
 assign wire8669* = ( (~ wire8669) ) ;
 assign key<60>* = ( (~ key<60>) ) ;
 assign wire8673* = ( (~ wire8673) ) ;
 assign D<13>* = ( (~ D<13>) ) ;
 assign wire7450* = ( (~ wire7450) ) ;
 assign key<5>* = ( (~ key<5>) ) ;
 assign wire8678* = ( (~ wire8678) ) ;
 assign D<12>* = ( (~ D<12>) ) ;
 assign wire7469* = ( (~ wire7469) ) ;
 assign key<13>* = ( (~ key<13>) ) ;
 assign wire8683* = ( (~ wire8683) ) ;
 assign D<11>* = ( (~ D<11>) ) ;
 assign wire7462* = ( (~ wire7462) ) ;
 assign key<21>* = ( (~ key<21>) ) ;
 assign wire8688* = ( (~ wire8688) ) ;
 assign D<10>* = ( (~ D<10>) ) ;
 assign wire7455* = ( (~ wire7455) ) ;
 assign key<29>* = ( (~ key<29>) ) ;
 assign wire8693* = ( (~ wire8693) ) ;
 assign D<9>* = ( (~ D<9>) ) ;
 assign wire8695* = ( (~ wire8695) ) ;
 assign key<37>* = ( (~ key<37>) ) ;
 assign wire8699* = ( (~ wire8699) ) ;
 assign D<8>* = ( (~ D<8>) ) ;
 assign wire7466* = ( (~ wire7466) ) ;
 assign key<45>* = ( (~ key<45>) ) ;
 assign wire8704* = ( (~ wire8704) ) ;
 assign D<7>* = ( (~ D<7>) ) ;
 assign wire7448* = ( (~ wire7448) ) ;
 assign key<53>* = ( (~ key<53>) ) ;
 assign wire8709* = ( (~ wire8709) ) ;
 assign D<6>* = ( (~ D<6>) ) ;
 assign wire8711* = ( (~ wire8711) ) ;
 assign key<61>* = ( (~ key<61>) ) ;
 assign wire8715* = ( (~ wire8715) ) ;
 assign D<5>* = ( (~ D<5>) ) ;
 assign wire7453* = ( (~ wire7453) ) ;
 assign key<6>* = ( (~ key<6>) ) ;
 assign wire8720* = ( (~ wire8720) ) ;
 assign D<4>* = ( (~ D<4>) ) ;
 assign wire7459* = ( (~ wire7459) ) ;
 assign key<14>* = ( (~ key<14>) ) ;
 assign wire8725* = ( (~ wire8725) ) ;
 assign D<3>* = ( (~ D<3>) ) ;
 assign wire7446* = ( (~ wire7446) ) ;
 assign key<22>* = ( (~ key<22>) ) ;
 assign wire8730* = ( (~ wire8730) ) ;
 assign D<2>* = ( (~ D<2>) ) ;
 assign wire7467* = ( (~ wire7467) ) ;
 assign key<30>* = ( (~ key<30>) ) ;
 assign wire8735* = ( (~ wire8735) ) ;
 assign key<38>* = ( (~ key<38>) ) ;
 assign wire8740* = ( (~ wire8740) ) ;
 assign key<46>* = ( (~ key<46>) ) ;
 assign wire8745* = ( (~ wire8745) ) ;
 assign key<54>* = ( (~ key<54>) ) ;
 assign wire8750* = ( (~ wire8750) ) ;
 assign wire7570* = ( (~ wire7570) ) ;
 assign wire7596* = ( (~ wire7596) ) ;
 assign wire8756* = ( (~ wire8756) ) ;
 assign wire8757* = ( (~ wire8757) ) ;


endmodule

