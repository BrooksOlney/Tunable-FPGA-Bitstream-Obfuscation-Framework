module ks_pdc_qmap_map (sk, i_5_, i_3_, i_4_, i_1_, i_0_, i_2_, i_8_, i_7_, i_6_, i_9_, i_10_, i_11_, i_15_, i_14_, i_12_, i_13_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_);

	input i_5_;
	input i_3_;
	input i_4_;
	input i_1_;
	input i_0_;
	input i_2_;
	input i_8_;
	input i_7_;
	input i_6_;
	input i_9_;
	input i_10_;
	input i_11_;
	input i_15_;
	input i_14_;
	input i_12_;
	input i_13_;
	output o_0_;
	output o_1_;
	output o_2_;
	output o_3_;
	output o_4_;
	output o_5_;
	output o_6_;
	output o_7_;
	output o_8_;
	output o_9_;
	output o_10_;
	output o_11_;
	output o_12_;
	output o_13_;
	output o_14_;
	output o_15_;
	output o_16_;
	output o_17_;
	output o_18_;
	output o_19_;
	output o_20_;
	output o_21_;
	output o_22_;
	output o_23_;
	output o_24_;
	output o_25_;
	output o_26_;
	output o_27_;
	output o_28_;
	output o_29_;
	output o_30_;
	output o_31_;
	output o_32_;
	output o_33_;
	output o_34_;
	output o_35_;
	output o_36_;
	output o_37_;
	output o_38_;
	output o_39_;

	input [127 : 0] sk /* synthesis noprune */;


	wire g854, g68, g874, g1029, g1640, g1094, g1137, g29, g1138, g1437, g1467, g1469, g1476, g1477, g1491, g1503, g1506, g1509, g1530, g1, g2;
	wire g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23;
	wire g24, g25, g26, g27, g28, g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44, g45;
	wire g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66;
	wire g67, g69, g70, g71, g72, g73, g75, g76, g77, g78, g79, g80, g81, g82, g1544, g83, g85, g87, g88, g89, g90;
	wire g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111;
	wire g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g132;
	wire g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153;
	wire g154, g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g1775, g168, g1782, g169, g170, g171, g172;
	wire g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193;
	wire g194, g195, g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207, g208, g209, g210, g211, g212, g213, g214;
	wire g215, g216, g217, g218, g219, g220, g221, g222, g223, g224, g225, g226, g227, g228, g229, g230, g231, g232, g233, g234, g1543;
	wire g235, g236, g237, g238, g239, g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250, g251, g252, g253, g254, g255;
	wire g256, g257, g258, g259, g260, g261, g262, g263, g264, g265, g266, g267, g268, g269, g270, g271, g272, g273, g274, g275, g276;
	wire g277, g278, g279, g280, g281, g282, g283, g284, g285, g286, g287, g288, g289, g290, g291, g292, g293, g294, g295, g296, g297;
	wire g298, g299, g300, g301, g302, g303, g304, g305, g306, g307, g308, g309, g310, g311, g312, g313, g314, g315, g316, g317, g318;
	wire g319, g320, g321, g1768, g322, g323, g324, g325, g326, g327, g328, g329, g330, g331, g332, g333, g334, g1761, g335, g336, g337;
	wire g338, g339, g340, g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351, g352, g353, g354, g355, g356, g357, g358;
	wire g359, g360, g361, g362, g363, g364, g365, g366, g367, g368, g369, g370, g371, g372, g373, g1754, g374, g375, g376, g377, g378;
	wire g379, g380, g381, g382, g383, g384, g385, g386, g387, g388, g389, g390, g391, g392, g393, g394, g395, g396, g397, g398, g399;
	wire g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410, g1747, g411, g412, g413, g414, g415, g416, g417, g418, g419;
	wire g420, g421, g422, g423, g424, g425, g426, g427, g428, g429, g430, g431, g432, g433, g434, g435, g436, g437, g438, g439, g440;
	wire g441, g442, g443, g444, g445, g446, g447, g448, g449, g450, g451, g452, g453, g454, g455, g456, g457, g458, g460, g461, g462;
	wire g463, g464, g465, g466, g467, g468, g469, g470, g471, g472, g473, g474, g475, g476, g477, g478, g479, g480, g481, g482, g483;
	wire g484, g485, g486, g487, g488, g489, g490, g491, g492, g493, g494, g495, g496, g497, g498, g499, g500, g501, g502, g503, g504;
	wire g505, g506, g507, g508, g509, g510, g511, g512, g513, g514, g515, g516, g517, g518, g519, g520, g1737, g1728, g521, g522, g523;
	wire g524, g525, g526, g527, g528, g529, g530, g531, g532, g533, g534, g535, g536, g537, g538, g539, g540, g541, g542, g1721, g543;
	wire g544, g545, g546, g547, g548, g549, g550, g551, g552, g553, g554, g555, g556, g557, g558, g559, g560, g561, g562, g563, g564;
	wire g565, g566, g567, g1708, g568, g569, g570, g571, g572, g573, g574, g575, g576, g577, g578, g579, g580, g581, g582, g583, g584;
	wire g585, g586, g587, g588, g589, g590, g591, g592, g593, g594, g595, g596, g597, g598, g599, g600, g601, g602, g603, g604, g605;
	wire g606, g1695, g607, g608, g609, g610, g611, g612, g613, g614, g615, g616, g617, g618, g619, g620, g621, g622, g623, g624, g625;
	wire g626, g627, g628, g629, g630, g631, g632, g1686, g633, g634, g635, g636, g637, g638, g639, g640, g641, g642, g643, g644, g645;
	wire g646, g647, g648, g649, g650, g651, g652, g653, g654, g655, g656, g657, g658, g659, g660, g661, g662, g663, g664, g666, g667;
	wire g668, g669, g670, g671, g672, g673, g674, g675, g676, g677, g678, g679, g680, g681, g682, g683, g684, g685, g686, g687, g688;
	wire g689, g690, g691, g692, g693, g694, g695, g696, g697, g698, g699, g700, g701, g702, g703, g704, g705, g706, g707, g708, g709;
	wire g710, g711, g712, g713, g714, g715, g716, g717, g718, g719, g720, g721, g722, g723, g724, g725, g726, g727, g728, g729, g730;
	wire g731, g732, g733, g734, g735, g736, g737, g738, g739, g740, g741, g742, g743, g744, g745, g746, g747, g748, g749, g750, g751;
	wire g752, g753, g754, g755, g756, g757, g758, g759, g760, g761, g762, g763, g764, g765, g766, g767, g768, g769, g770, g771, g772;
	wire g773, g774, g775, g776, g777, g778, g779, g780, g781, g782, g783, g784, g785, g786, g787, g788, g789, g790, g791, g792, g793;
	wire g794, g795, g796, g797, g798, g799, g800, g801, g802, g803, g804, g805, g806, g807, g808, g809, g810, g811, g812, g813, g814;
	wire g815, g1673, g1666, g816, g817, g818, g819, g820, g821, g822, g823, g824, g825, g826, g827, g828, g829, g830, g831, g832, g833;
	wire g834, g835, g836, g837, g838, g839, g840, g1653, g841, g842, g843, g844, g845, g846, g847, g848, g849, g850, g851, g852, g853;
	wire g855, g857, g858, g859, g860, g861, g862, g863, g864, g865, g866, g867, g868, g869, g870, g871, g872, g873, g875, g876, g877;
	wire g878, g879, g880, g881, g882, g883, g884, g885, g886, g887, g888, g889, g890, g891, g892, g893, g894, g895, g896, g897, g898;
	wire g899, g900, g901, g902, g903, g904, g905, g906, g907, g908, g909, g910, g911, g912, g913, g914, g915, g916, g917, g918, g919;
	wire g920, g921, g922, g923, g924, g925, g926, g927, g928, g929, g930, g931, g932, g933, g934, g935, g936, g937, g938, g939, g940;
	wire g941, g942, g943, g944, g945, g946, g947, g948, g949, g950, g951, g952, g953, g954, g955, g956, g957, g958, g959, g960, g961;
	wire g962, g963, g964, g965, g966, g967, g968, g970, g971, g972, g973, g974, g975, g976, g977, g978, g979, g980, g981, g982, g983;
	wire g984, g985, g986, g987, g988, g989, g990, g991, g992, g993, g994, g995, g996, g997, g998, g999, g1000, g1001, g1002, g1003, g1004;
	wire g1005, g1006, g1007, g1008, g1009, g1010, g1011, g1012, g1013, g1014, g1015, g1016, g1017, g1018, g1019, g1020, g1021, g1022, g1023, g1024, g1025;
	wire g1026, g1027, g1542, g1028, g1030, g1031, g1032, g1033, g1034, g1035, g1036, g1037, g1038, g1039, g1040, g1041, g1042, g1043, g1044, g1045, g1046;
	wire g1047, g1048, g1049, g1050, g1051, g1052, g1053, g1054, g1055, g1056, g1057, g1058, g1059, g1060, g1061, g1062, g1063, g1064, g1065, g1066, g1067;
	wire g1068, g1069, g1070, g1071, g1072, g1073, g1074, g1075, g1076, g1077, g1078, g1079, g1080, g1081, g1082, g1083, g1084, g1085, g1086, g1087, g1088;
	wire g1089, g1090, g1091, g1092, g1093, g1095, g1096, g1097, g1098, g1099, g1100, g1541, g1101, g1102, g1103, g1104, g1628, g1622, g1105, g1106, g1107;
	wire g1108, g1109, g1110, g1111, g1112, g1113, g1114, g1115, g1116, g1117, g1118, g1616, g1119, g1120, g1121, g1122, g1123, g1124, g1125, g1126, g1127;
	wire g1128, g1129, g1130, g1131, g1132, g1133, g1134, g1135, g1136, g1139, g1140, g1141, g1142, g1143, g1144, g1145, g1146, g1147, g1148, g1149, g1150;
	wire g1151, g1152, g1153, g1154, g1155, g1156, g1157, g1158, g1159, g1160, g1161, g1162, g1163, g1164, g1165, g1166, g1167, g1168, g1169, g1170, g1171;
	wire g1172, g1173, g1174, g1175, g1176, g1177, g1178, g1179, g1180, g1181, g1182, g1183, g1184, g1185, g1186, g1187, g1188, g1189, g1191, g1192, g1193;
	wire g1194, g1195, g1196, g1197, g1198, g1199, g1200, g1201, g1202, g1203, g1204, g1205, g1206, g1207, g1208, g1209, g1210, g1211, g1212, g1213, g1214;
	wire g1215, g1216, g1607, g1217, g1218, g1219, g1220, g1221, g1222, g1223, g1224, g1225, g1226, g1227, g1228, g1229, g1230, g1231, g1232, g1233, g1234;
	wire g1235, g1236, g1237, g1238, g1239, g1240, g1241, g1242, g1243, g1244, g1245, g1246, g1247, g1248, g1249, g1250, g1251, g1252, g1253, g1254, g1255;
	wire g1256, g1257, g1258, g1259, g1260, g1261, g1262, g1263, g1264, g1265, g1266, g1267, g1268, g1269, g1270, g1271, g1272, g1273, g1274, g1275, g1276;
	wire g1277, g1278, g1279, g1280, g1281, g1282, g1283, g1284, g1285, g1286, g1287, g1288, g1289, g1290, g1291, g1292, g1293, g1294, g1295, g1296, g1297;
	wire g1298, g1299, g1596, g1300, g1301, g1303, g1304, g1305, g1306, g1307, g1308, g1309, g1310, g1311, g1312, g1313, g1314, g1315, g1316, g1317, g1318;
	wire g1319, g1320, g1321, g1322, g1323, g1324, g1325, g1326, g1327, g1328, g1329, g1589, g1330, g1331, g1332, g1333, g1334, g1335, g1336, g1337, g1338;
	wire g1339, g1340, g1341, g1342, g1343, g1344, g1345, g1346, g1347, g1348, g1349, g1350, g1351, g1352, g1353, g1354, g1355, g1356, g1357, g1358, g1359;
	wire g1360, g1361, g1362, g1363, g1364, g1365, g1366, g1367, g1368, g1369, g1370, g1371, g1372, g1580, g1373, g1374, g1375, g1376, g1377, g1378, g1379;
	wire g1380, g1381, g1382, g1384, g1385, g1386, g1387, g1388, g1389, g1390, g1391, g1538, g1392, g1393, g1394, g1395, g1396, g1397, g1398, g1399, g1400;
	wire g1401, g1402, g1403, g1404, g1405, g1406, g1407, g1408, g1409, g1410, g1411, g1558, g1412, g1413, g1568, g1415, g1416, g1417, g1418, g1419, g1420;
	wire g1421, g1422, g1423, g1424, g1425, g1426, g1427, g1428, g1429, g1430, g1431, g1432, g1433, g1434, g1435, g1438, g1439, g1441, g1442, g1443, g1444;
	wire g1445, g1446, g1447, g1448, g1449, g1450, g1451, g1545, g1452, g1453, g1454, g1455, g1456, g1457, g1458, g1459, g1460, g1461, g1462, g1463, g1464;
	wire g1465, g1466, g1468, g1470, g1471, g1472, g1473, g1474, g1475, g1479, g1480, g1481, g1482, g1483, g1484, g1485, g1486, g1487, g1488, g1489, g1490;
	wire g1492, g1493, g1494, g1495, g1496, g1497, g1498, g1499, g1501, g1502, g1504, g1507, g1508, g1510, g1511, g1512, g1513, g1514, g1515, g1516, g1517;
	wire g1518, g1519, g1520, g1521, g1522, g1524, g1526, g1527, g1528, g1529, g1531, g1532, g1536, g1537, g1539, g1540, g1546, g1547, g1548, g1551, g1549;
	wire g1550, g1554, g1555, g1552, g1553, g1556, g1557, g1559, g1560, g1561, g1564, g1562, g1563, g1566, g1565, g1567, g1569, g1570, g1571, g1574, g1572;
	wire g1573, g1577, g1578, g1575, g1576, g1579, g1581, g1582, g1583, g1585, g1584, g1587, g1586, g1588, g1590, g1591, g1592, g1593, g1594, g1595, g1597;
	wire g1598, g1599, g1601, g1600, g1604, g1602, g1603, g1605, g1606, g1608, g1609, g1610, g1613, g1611, g1612, g1614, g1615, g1617, g1618, g1619, g1620;
	wire g1621, g1623, g1624, g1625, g1626, g1627, g1629, g1630, g1631, g1634, g1632, g1633, g1637, g1635, g1636, g1638, g1639, g1641, g1642, g1643, g1646;
	wire g1644, g1645, g1649, g1650, g1647, g1648, g1651, g1652, g1654, g1655, g1656, g1659, g1657, g1658, g1662, g1663, g1660, g1661, g1664, g1665, g1667;
	wire g1668, g1669, g1670, g1671, g1672, g1674, g1675, g1676, g1679, g1677, g1678, g1682, g1683, g1680, g1681, g1684, g1685, g1687, g1688, g1689, g1691;
	wire g1690, g1693, g1692, g1694, g1696, g1697, g1698, g1701, g1699, g1700, g1704, g1705, g1702, g1703, g1706, g1707, g1709, g1710, g1711, g1714, g1712;
	wire g1713, g1717, g1718, g1715, g1716, g1719, g1720, g1722, g1723, g1724, g1725, g1726, g1727, g1729, g1730, g1731, g1732, g1733, g1734, g1735, g1736;
	wire g1738, g1739, g1740, g1741, g1744, g1742, g1743, g1745, g1746, g1748, g1749, g1750, g1751, g1752, g1753, g1755, g1756, g1757, g1758, g1759, g1760;
	wire g1762, g1763, g1764, g1765, g1766, g1767, g1769, g1770, g1771, g1772, g1773, g1774, g1776, g1777, g1778, g1779, g1780, g1781, g1783, g1784, g1785;
	wire g1786, g1789, g1787, g1788, g1790, g1791;

	assign o_5_ = (((sk[0]) & (!g854)));
	assign o_6_ = (((sk[1]) & (!g68)));
	assign o_8_ = (((sk[2]) & (!g874)));
	assign o_10_ = (((sk[3]) & (!g1029)));
	assign o_11_ = (((sk[4]) & (!g1640)));
	assign o_12_ = (((sk[5]) & (!g1094)));
	assign o_13_ = (((sk[6]) & (!g1137)));
	assign o_14_ = (((sk[7]) & (g29)));
	assign o_15_ = (((sk[8]) & (!g1138)));
	assign o_21_ = (((sk[9]) & (!g1437)));
	assign o_23_ = (((sk[10]) & (!g1467)));
	assign o_24_ = (((sk[11]) & (!g1469)));
	assign o_25_ = (((sk[12]) & (!g1476)));
	assign o_26_ = (((sk[13]) & (!g1477)));
	assign o_28_ = (((sk[14]) & (!g1491)));
	assign o_30_ = (((sk[15]) & (!g1503)));
	assign o_32_ = (((sk[16]) & (!g1506)));
	assign o_33_ = (((sk[17]) & (!g1509)));
	assign o_36_ = (((sk[18]) & (!g1530)));
	assign g1 = (((!sk[19]) & (!i_1_) & (!i_0_) & (i_2_)) + ((!sk[19]) & (!i_1_) & (i_0_) & (i_2_)) + ((!sk[19]) & (i_1_) & (!i_0_) & (!i_2_)) + ((!sk[19]) & (i_1_) & (!i_0_) & (i_2_)) + ((!sk[19]) & (i_1_) & (i_0_) & (!i_2_)) + ((!sk[19]) & (i_1_) & (i_0_) & (i_2_)) + ((sk[19]) & (i_1_) & (!i_0_) & (!i_2_)));
	assign g2 = (((!i_5_) & (!sk[20]) & (!i_3_) & (!i_4_) & (g1)) + ((!i_5_) & (!sk[20]) & (!i_3_) & (i_4_) & (!g1)) + ((!i_5_) & (!sk[20]) & (!i_3_) & (i_4_) & (g1)) + ((!i_5_) & (!sk[20]) & (i_3_) & (!i_4_) & (g1)) + ((!i_5_) & (!sk[20]) & (i_3_) & (i_4_) & (!g1)) + ((!i_5_) & (!sk[20]) & (i_3_) & (i_4_) & (g1)) + ((!i_5_) & (sk[20]) & (!i_3_) & (!i_4_) & (g1)) + ((i_5_) & (!sk[20]) & (!i_3_) & (!i_4_) & (g1)) + ((i_5_) & (!sk[20]) & (!i_3_) & (i_4_) & (!g1)) + ((i_5_) & (!sk[20]) & (!i_3_) & (i_4_) & (g1)) + ((i_5_) & (!sk[20]) & (i_3_) & (!i_4_) & (g1)) + ((i_5_) & (!sk[20]) & (i_3_) & (i_4_) & (!g1)) + ((i_5_) & (!sk[20]) & (i_3_) & (i_4_) & (g1)));
	assign g3 = (((!sk[21]) & (!g2) & (!i_8_) & (i_7_)) + ((!sk[21]) & (!g2) & (i_8_) & (i_7_)) + ((!sk[21]) & (g2) & (!i_8_) & (!i_7_)) + ((!sk[21]) & (g2) & (!i_8_) & (i_7_)) + ((!sk[21]) & (g2) & (i_8_) & (!i_7_)) + ((!sk[21]) & (g2) & (i_8_) & (i_7_)) + ((sk[21]) & (g2) & (i_8_) & (!i_7_)));
	assign g4 = (((!sk[22]) & (!i_6_) & (i_7_)) + ((!sk[22]) & (i_6_) & (i_7_)) + ((sk[22]) & (i_6_) & (i_7_)));
	assign g5 = (((!i_9_) & (!sk[23]) & (i_10_)) + ((!i_9_) & (sk[23]) & (!i_10_)) + ((i_9_) & (!sk[23]) & (i_10_)));
	assign g6 = (((!i_11_) & (!i_9_) & (!sk[24]) & (i_10_)) + ((!i_11_) & (i_9_) & (!sk[24]) & (i_10_)) + ((!i_11_) & (i_9_) & (sk[24]) & (!i_10_)) + ((i_11_) & (!i_9_) & (!sk[24]) & (!i_10_)) + ((i_11_) & (!i_9_) & (!sk[24]) & (i_10_)) + ((i_11_) & (i_9_) & (!sk[24]) & (!i_10_)) + ((i_11_) & (i_9_) & (!sk[24]) & (i_10_)));
	assign g7 = (((!i_14_) & (!i_12_) & (!sk[25]) & (i_13_)) + ((!i_14_) & (!i_12_) & (sk[25]) & (!i_13_)) + ((!i_14_) & (i_12_) & (!sk[25]) & (i_13_)) + ((i_14_) & (!i_12_) & (!sk[25]) & (!i_13_)) + ((i_14_) & (!i_12_) & (!sk[25]) & (i_13_)) + ((i_14_) & (i_12_) & (!sk[25]) & (!i_13_)) + ((i_14_) & (i_12_) & (!sk[25]) & (i_13_)));
	assign g8 = (((!g6) & (!sk[26]) & (!i_15_) & (g7)) + ((!g6) & (!sk[26]) & (i_15_) & (g7)) + ((!g6) & (sk[26]) & (!i_15_) & (!g7)) + ((!g6) & (sk[26]) & (!i_15_) & (g7)) + ((!g6) & (sk[26]) & (i_15_) & (!g7)) + ((!g6) & (sk[26]) & (i_15_) & (g7)) + ((g6) & (!sk[26]) & (!i_15_) & (!g7)) + ((g6) & (!sk[26]) & (!i_15_) & (g7)) + ((g6) & (!sk[26]) & (i_15_) & (!g7)) + ((g6) & (!sk[26]) & (i_15_) & (g7)) + ((g6) & (sk[26]) & (!i_15_) & (!g7)) + ((g6) & (sk[26]) & (!i_15_) & (g7)) + ((g6) & (sk[26]) & (i_15_) & (!g7)));
	assign g9 = (((!i_14_) & (!i_12_) & (!sk[27]) & (i_13_)) + ((!i_14_) & (!i_12_) & (sk[27]) & (i_13_)) + ((!i_14_) & (i_12_) & (!sk[27]) & (i_13_)) + ((i_14_) & (!i_12_) & (!sk[27]) & (!i_13_)) + ((i_14_) & (!i_12_) & (!sk[27]) & (i_13_)) + ((i_14_) & (i_12_) & (!sk[27]) & (!i_13_)) + ((i_14_) & (i_12_) & (!sk[27]) & (i_13_)));
	assign g10 = (((!g6) & (!sk[28]) & (!i_15_) & (g9)) + ((!g6) & (!sk[28]) & (i_15_) & (g9)) + ((g6) & (!sk[28]) & (!i_15_) & (!g9)) + ((g6) & (!sk[28]) & (!i_15_) & (g9)) + ((g6) & (!sk[28]) & (i_15_) & (!g9)) + ((g6) & (!sk[28]) & (i_15_) & (g9)) + ((g6) & (sk[28]) & (!i_15_) & (g9)));
	assign g11 = (((!i_11_) & (!i_9_) & (!i_10_) & (!sk[29]) & (i_15_)) + ((!i_11_) & (!i_9_) & (i_10_) & (!sk[29]) & (!i_15_)) + ((!i_11_) & (!i_9_) & (i_10_) & (!sk[29]) & (i_15_)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[29]) & (i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[29]) & (!i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[29]) & (i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (sk[29]) & (!i_15_)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[29]) & (i_15_)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[29]) & (!i_15_)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[29]) & (i_15_)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[29]) & (i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[29]) & (!i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[29]) & (i_15_)));
	assign g12 = (((!sk[30]) & (!g11) & (g9)) + ((!sk[30]) & (g11) & (g9)) + ((sk[30]) & (g11) & (g9)));
	assign g13 = (((!sk[31]) & (!i_14_) & (!i_12_) & (i_13_)) + ((!sk[31]) & (!i_14_) & (i_12_) & (i_13_)) + ((!sk[31]) & (i_14_) & (!i_12_) & (!i_13_)) + ((!sk[31]) & (i_14_) & (!i_12_) & (i_13_)) + ((!sk[31]) & (i_14_) & (i_12_) & (!i_13_)) + ((!sk[31]) & (i_14_) & (i_12_) & (i_13_)) + ((sk[31]) & (i_14_) & (!i_12_) & (!i_13_)));
	assign g14 = (((!g6) & (!i_15_) & (!sk[32]) & (g13)) + ((!g6) & (i_15_) & (!sk[32]) & (g13)) + ((g6) & (!i_15_) & (!sk[32]) & (!g13)) + ((g6) & (!i_15_) & (!sk[32]) & (g13)) + ((g6) & (!i_15_) & (sk[32]) & (g13)) + ((g6) & (i_15_) & (!sk[32]) & (!g13)) + ((g6) & (i_15_) & (!sk[32]) & (g13)));
	assign g15 = (((!i_11_) & (!i_9_) & (!sk[33]) & (!i_10_) & (i_15_)) + ((!i_11_) & (!i_9_) & (!sk[33]) & (i_10_) & (!i_15_)) + ((!i_11_) & (!i_9_) & (!sk[33]) & (i_10_) & (i_15_)) + ((!i_11_) & (!i_9_) & (sk[33]) & (!i_10_) & (!i_15_)) + ((!i_11_) & (!i_9_) & (sk[33]) & (!i_10_) & (i_15_)) + ((!i_11_) & (!i_9_) & (sk[33]) & (i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (!sk[33]) & (!i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (!sk[33]) & (i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (!sk[33]) & (i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (sk[33]) & (!i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (sk[33]) & (!i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (sk[33]) & (i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (sk[33]) & (i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (!sk[33]) & (!i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (!sk[33]) & (i_10_) & (!i_15_)) + ((i_11_) & (!i_9_) & (!sk[33]) & (i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (sk[33]) & (!i_10_) & (!i_15_)) + ((i_11_) & (!i_9_) & (sk[33]) & (!i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (sk[33]) & (i_10_) & (!i_15_)) + ((i_11_) & (!i_9_) & (sk[33]) & (i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (!sk[33]) & (!i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (!sk[33]) & (i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (!sk[33]) & (i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (sk[33]) & (!i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (sk[33]) & (!i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (sk[33]) & (i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (sk[33]) & (i_10_) & (i_15_)));
	assign g16 = (((!sk[34]) & (!g15) & (g9)) + ((!sk[34]) & (g15) & (g9)) + ((sk[34]) & (!g15) & (!g9)) + ((sk[34]) & (g15) & (!g9)) + ((sk[34]) & (g15) & (g9)));
	assign g17 = (((!g12) & (!g14) & (!sk[35]) & (g16)) + ((!g12) & (!g14) & (sk[35]) & (g16)) + ((!g12) & (g14) & (!sk[35]) & (g16)) + ((g12) & (!g14) & (!sk[35]) & (!g16)) + ((g12) & (!g14) & (!sk[35]) & (g16)) + ((g12) & (g14) & (!sk[35]) & (!g16)) + ((g12) & (g14) & (!sk[35]) & (g16)));
	assign g18 = (((!i_11_) & (!sk[36]) & (!i_9_) & (!i_10_) & (i_15_)) + ((!i_11_) & (!sk[36]) & (!i_9_) & (i_10_) & (!i_15_)) + ((!i_11_) & (!sk[36]) & (!i_9_) & (i_10_) & (i_15_)) + ((!i_11_) & (!sk[36]) & (i_9_) & (!i_10_) & (i_15_)) + ((!i_11_) & (!sk[36]) & (i_9_) & (i_10_) & (!i_15_)) + ((!i_11_) & (!sk[36]) & (i_9_) & (i_10_) & (i_15_)) + ((!i_11_) & (sk[36]) & (!i_9_) & (!i_10_) & (!i_15_)) + ((!i_11_) & (sk[36]) & (!i_9_) & (!i_10_) & (i_15_)) + ((!i_11_) & (sk[36]) & (!i_9_) & (i_10_) & (!i_15_)) + ((!i_11_) & (sk[36]) & (i_9_) & (!i_10_) & (!i_15_)) + ((!i_11_) & (sk[36]) & (i_9_) & (!i_10_) & (i_15_)) + ((!i_11_) & (sk[36]) & (i_9_) & (i_10_) & (!i_15_)) + ((!i_11_) & (sk[36]) & (i_9_) & (i_10_) & (i_15_)) + ((i_11_) & (!sk[36]) & (!i_9_) & (!i_10_) & (i_15_)) + ((i_11_) & (!sk[36]) & (!i_9_) & (i_10_) & (!i_15_)) + ((i_11_) & (!sk[36]) & (!i_9_) & (i_10_) & (i_15_)) + ((i_11_) & (!sk[36]) & (i_9_) & (!i_10_) & (i_15_)) + ((i_11_) & (!sk[36]) & (i_9_) & (i_10_) & (!i_15_)) + ((i_11_) & (!sk[36]) & (i_9_) & (i_10_) & (i_15_)) + ((i_11_) & (sk[36]) & (!i_9_) & (!i_10_) & (!i_15_)) + ((i_11_) & (sk[36]) & (!i_9_) & (!i_10_) & (i_15_)) + ((i_11_) & (sk[36]) & (!i_9_) & (i_10_) & (!i_15_)) + ((i_11_) & (sk[36]) & (!i_9_) & (i_10_) & (i_15_)) + ((i_11_) & (sk[36]) & (i_9_) & (!i_10_) & (!i_15_)) + ((i_11_) & (sk[36]) & (i_9_) & (!i_10_) & (i_15_)) + ((i_11_) & (sk[36]) & (i_9_) & (i_10_) & (!i_15_)) + ((i_11_) & (sk[36]) & (i_9_) & (i_10_) & (i_15_)));
	assign g19 = (((!g7) & (!sk[37]) & (g18)) + ((g7) & (!sk[37]) & (g18)) + ((g7) & (sk[37]) & (!g18)));
	assign g20 = (((!g15) & (!sk[38]) & (g13)) + ((!g15) & (sk[38]) & (!g13)) + ((g15) & (!sk[38]) & (g13)) + ((g15) & (sk[38]) & (!g13)) + ((g15) & (sk[38]) & (g13)));
	assign g21 = (((!sk[39]) & (!g13) & (g11)) + ((!sk[39]) & (g13) & (g11)) + ((sk[39]) & (g13) & (g11)));
	assign g22 = (((!sk[40]) & (!i_11_) & (!i_9_) & (!i_10_) & (i_15_)) + ((!sk[40]) & (!i_11_) & (!i_9_) & (i_10_) & (!i_15_)) + ((!sk[40]) & (!i_11_) & (!i_9_) & (i_10_) & (i_15_)) + ((!sk[40]) & (!i_11_) & (i_9_) & (!i_10_) & (i_15_)) + ((!sk[40]) & (!i_11_) & (i_9_) & (i_10_) & (!i_15_)) + ((!sk[40]) & (!i_11_) & (i_9_) & (i_10_) & (i_15_)) + ((!sk[40]) & (i_11_) & (!i_9_) & (!i_10_) & (i_15_)) + ((!sk[40]) & (i_11_) & (!i_9_) & (i_10_) & (!i_15_)) + ((!sk[40]) & (i_11_) & (!i_9_) & (i_10_) & (i_15_)) + ((!sk[40]) & (i_11_) & (i_9_) & (!i_10_) & (i_15_)) + ((!sk[40]) & (i_11_) & (i_9_) & (i_10_) & (!i_15_)) + ((!sk[40]) & (i_11_) & (i_9_) & (i_10_) & (i_15_)) + ((sk[40]) & (!i_11_) & (i_9_) & (i_10_) & (i_15_)));
	assign g23 = (((g7) & (!sk[41]) & (!g22)) + ((g7) & (!sk[41]) & (g22)) + ((g7) & (sk[41]) & (g22)));
	assign g24 = (((!sk[42]) & (!g19) & (g20) & (g21) & (!g23)) + ((!sk[42]) & (!g19) & (g20) & (g21) & (g23)) + ((!sk[42]) & (g19) & (!g20) & (!g21) & (!g23)) + ((!sk[42]) & (g19) & (!g20) & (!g21) & (g23)) + ((!sk[42]) & (g19) & (!g20) & (g21) & (!g23)) + ((!sk[42]) & (g19) & (!g20) & (g21) & (g23)) + ((!sk[42]) & (g19) & (g20) & (!g21) & (!g23)) + ((!sk[42]) & (g19) & (g20) & (!g21) & (g23)) + ((!sk[42]) & (g19) & (g20) & (g21) & (!g23)) + ((!sk[42]) & (g19) & (g20) & (g21) & (g23)) + ((sk[42]) & (!g19) & (g20) & (!g21) & (!g23)));
	assign g25 = (((!g8) & (g10) & (!sk[43]) & (g17) & (!g24)) + ((!g8) & (g10) & (!sk[43]) & (g17) & (g24)) + ((g8) & (!g10) & (!sk[43]) & (!g17) & (!g24)) + ((g8) & (!g10) & (!sk[43]) & (!g17) & (g24)) + ((g8) & (!g10) & (!sk[43]) & (g17) & (!g24)) + ((g8) & (!g10) & (!sk[43]) & (g17) & (g24)) + ((g8) & (!g10) & (sk[43]) & (g17) & (g24)) + ((g8) & (g10) & (!sk[43]) & (!g17) & (!g24)) + ((g8) & (g10) & (!sk[43]) & (!g17) & (g24)) + ((g8) & (g10) & (!sk[43]) & (g17) & (!g24)) + ((g8) & (g10) & (!sk[43]) & (g17) & (g24)));
	assign g26 = (((!g5) & (sk[44]) & (g25)) + ((g5) & (!sk[44]) & (!g25)) + ((g5) & (!sk[44]) & (g25)));
	assign g27 = (((!i_8_) & (sk[45]) & (i_6_) & (!i_7_)) + ((i_8_) & (!sk[45]) & (!i_6_) & (!i_7_)) + ((i_8_) & (!sk[45]) & (!i_6_) & (i_7_)) + ((i_8_) & (!sk[45]) & (i_6_) & (!i_7_)) + ((i_8_) & (!sk[45]) & (i_6_) & (i_7_)));
	assign g28 = (((!g2) & (g4) & (!sk[46]) & (g26) & (!g27)) + ((!g2) & (g4) & (!sk[46]) & (g26) & (g27)) + ((g2) & (!g4) & (!sk[46]) & (!g26) & (!g27)) + ((g2) & (!g4) & (!sk[46]) & (!g26) & (g27)) + ((g2) & (!g4) & (!sk[46]) & (g26) & (!g27)) + ((g2) & (!g4) & (!sk[46]) & (g26) & (g27)) + ((g2) & (!g4) & (sk[46]) & (!g26) & (g27)) + ((g2) & (g4) & (!sk[46]) & (!g26) & (!g27)) + ((g2) & (g4) & (!sk[46]) & (!g26) & (g27)) + ((g2) & (g4) & (!sk[46]) & (g26) & (!g27)) + ((g2) & (g4) & (!sk[46]) & (g26) & (g27)) + ((g2) & (g4) & (sk[46]) & (!g26) & (!g27)) + ((g2) & (g4) & (sk[46]) & (!g26) & (g27)) + ((g2) & (g4) & (sk[46]) & (g26) & (!g27)) + ((g2) & (g4) & (sk[46]) & (g26) & (g27)));
	assign g29 = (((!i_1_) & (sk[47]) & (i_0_)) + ((i_1_) & (!sk[47]) & (!i_0_)) + ((i_1_) & (!sk[47]) & (i_0_)));
	assign g30 = (((!sk[48]) & (i_6_) & (!i_7_)) + ((!sk[48]) & (i_6_) & (i_7_)) + ((sk[48]) & (!i_6_) & (!i_7_)));
	assign g31 = (((!sk[49]) & (i_8_) & (!g30)) + ((!sk[49]) & (i_8_) & (g30)) + ((sk[49]) & (!i_8_) & (g30)));
	assign g32 = (((g2) & (!sk[50]) & (!g31)) + ((g2) & (!sk[50]) & (g31)) + ((g2) & (sk[50]) & (g31)));
	assign g33 = (((!g10) & (!g23) & (sk[51]) & (g17) & (!g5)) + ((!g10) & (g23) & (!sk[51]) & (g17) & (!g5)) + ((!g10) & (g23) & (!sk[51]) & (g17) & (g5)) + ((g10) & (!g23) & (!sk[51]) & (!g17) & (!g5)) + ((g10) & (!g23) & (!sk[51]) & (!g17) & (g5)) + ((g10) & (!g23) & (!sk[51]) & (g17) & (!g5)) + ((g10) & (!g23) & (!sk[51]) & (g17) & (g5)) + ((g10) & (g23) & (!sk[51]) & (!g17) & (!g5)) + ((g10) & (g23) & (!sk[51]) & (!g17) & (g5)) + ((g10) & (g23) & (!sk[51]) & (g17) & (!g5)) + ((g10) & (g23) & (!sk[51]) & (g17) & (g5)));
	assign g34 = (((!sk[52]) & (i_6_) & (!i_7_)) + ((!sk[52]) & (i_6_) & (i_7_)) + ((sk[52]) & (!i_6_) & (i_7_)));
	assign g35 = (((!sk[53]) & (!g8) & (!g2) & (!g31) & (!g19) & (g34)) + ((!sk[53]) & (!g8) & (!g2) & (!g31) & (g19) & (g34)) + ((!sk[53]) & (!g8) & (!g2) & (g31) & (!g19) & (g34)) + ((!sk[53]) & (!g8) & (!g2) & (g31) & (g19) & (g34)) + ((!sk[53]) & (!g8) & (g2) & (!g31) & (!g19) & (g34)) + ((!sk[53]) & (!g8) & (g2) & (!g31) & (g19) & (g34)) + ((!sk[53]) & (!g8) & (g2) & (g31) & (!g19) & (g34)) + ((!sk[53]) & (!g8) & (g2) & (g31) & (g19) & (g34)) + ((!sk[53]) & (g8) & (!g2) & (!g31) & (!g19) & (!g34)) + ((!sk[53]) & (g8) & (!g2) & (!g31) & (!g19) & (g34)) + ((!sk[53]) & (g8) & (!g2) & (!g31) & (g19) & (!g34)) + ((!sk[53]) & (g8) & (!g2) & (!g31) & (g19) & (g34)) + ((!sk[53]) & (g8) & (!g2) & (g31) & (!g19) & (!g34)) + ((!sk[53]) & (g8) & (!g2) & (g31) & (!g19) & (g34)) + ((!sk[53]) & (g8) & (!g2) & (g31) & (g19) & (!g34)) + ((!sk[53]) & (g8) & (!g2) & (g31) & (g19) & (g34)) + ((!sk[53]) & (g8) & (g2) & (!g31) & (!g19) & (!g34)) + ((!sk[53]) & (g8) & (g2) & (!g31) & (!g19) & (g34)) + ((!sk[53]) & (g8) & (g2) & (!g31) & (g19) & (!g34)) + ((!sk[53]) & (g8) & (g2) & (!g31) & (g19) & (g34)) + ((!sk[53]) & (g8) & (g2) & (g31) & (!g19) & (!g34)) + ((!sk[53]) & (g8) & (g2) & (g31) & (!g19) & (g34)) + ((!sk[53]) & (g8) & (g2) & (g31) & (g19) & (!g34)) + ((!sk[53]) & (g8) & (g2) & (g31) & (g19) & (g34)) + ((sk[53]) & (!g8) & (g2) & (!g31) & (!g19) & (g34)) + ((sk[53]) & (!g8) & (g2) & (!g31) & (g19) & (g34)) + ((sk[53]) & (!g8) & (g2) & (g31) & (!g19) & (!g34)) + ((sk[53]) & (!g8) & (g2) & (g31) & (!g19) & (g34)) + ((sk[53]) & (!g8) & (g2) & (g31) & (g19) & (!g34)) + ((sk[53]) & (!g8) & (g2) & (g31) & (g19) & (g34)) + ((sk[53]) & (g8) & (g2) & (!g31) & (!g19) & (g34)) + ((sk[53]) & (g8) & (g2) & (!g31) & (g19) & (g34)) + ((sk[53]) & (g8) & (g2) & (g31) & (!g19) & (g34)) + ((sk[53]) & (g8) & (g2) & (g31) & (g19) & (!g34)) + ((sk[53]) & (g8) & (g2) & (g31) & (g19) & (g34)));
	assign g36 = (((!g32) & (!g20) & (!g21) & (!g33) & (!sk[54]) & (g35)) + ((!g32) & (!g20) & (!g21) & (!g33) & (sk[54]) & (!g35)) + ((!g32) & (!g20) & (!g21) & (g33) & (!sk[54]) & (g35)) + ((!g32) & (!g20) & (!g21) & (g33) & (sk[54]) & (!g35)) + ((!g32) & (!g20) & (g21) & (!g33) & (!sk[54]) & (g35)) + ((!g32) & (!g20) & (g21) & (!g33) & (sk[54]) & (!g35)) + ((!g32) & (!g20) & (g21) & (g33) & (!sk[54]) & (g35)) + ((!g32) & (!g20) & (g21) & (g33) & (sk[54]) & (!g35)) + ((!g32) & (g20) & (!g21) & (!g33) & (!sk[54]) & (g35)) + ((!g32) & (g20) & (!g21) & (!g33) & (sk[54]) & (!g35)) + ((!g32) & (g20) & (!g21) & (g33) & (!sk[54]) & (g35)) + ((!g32) & (g20) & (!g21) & (g33) & (sk[54]) & (!g35)) + ((!g32) & (g20) & (g21) & (!g33) & (!sk[54]) & (g35)) + ((!g32) & (g20) & (g21) & (!g33) & (sk[54]) & (!g35)) + ((!g32) & (g20) & (g21) & (g33) & (!sk[54]) & (g35)) + ((!g32) & (g20) & (g21) & (g33) & (sk[54]) & (!g35)) + ((g32) & (!g20) & (!g21) & (!g33) & (!sk[54]) & (!g35)) + ((g32) & (!g20) & (!g21) & (!g33) & (!sk[54]) & (g35)) + ((g32) & (!g20) & (!g21) & (g33) & (!sk[54]) & (!g35)) + ((g32) & (!g20) & (!g21) & (g33) & (!sk[54]) & (g35)) + ((g32) & (!g20) & (g21) & (!g33) & (!sk[54]) & (!g35)) + ((g32) & (!g20) & (g21) & (!g33) & (!sk[54]) & (g35)) + ((g32) & (!g20) & (g21) & (g33) & (!sk[54]) & (!g35)) + ((g32) & (!g20) & (g21) & (g33) & (!sk[54]) & (g35)) + ((g32) & (g20) & (!g21) & (!g33) & (!sk[54]) & (!g35)) + ((g32) & (g20) & (!g21) & (!g33) & (!sk[54]) & (g35)) + ((g32) & (g20) & (!g21) & (g33) & (!sk[54]) & (!g35)) + ((g32) & (g20) & (!g21) & (g33) & (!sk[54]) & (g35)) + ((g32) & (g20) & (!g21) & (g33) & (sk[54]) & (!g35)) + ((g32) & (g20) & (g21) & (!g33) & (!sk[54]) & (!g35)) + ((g32) & (g20) & (g21) & (!g33) & (!sk[54]) & (g35)) + ((g32) & (g20) & (g21) & (g33) & (!sk[54]) & (!g35)) + ((g32) & (g20) & (g21) & (g33) & (!sk[54]) & (g35)));
	assign g37 = (((!i_3_) & (!i_4_) & (!sk[55]) & (!g28) & (!g29) & (g36)) + ((!i_3_) & (!i_4_) & (!sk[55]) & (!g28) & (g29) & (g36)) + ((!i_3_) & (!i_4_) & (!sk[55]) & (g28) & (!g29) & (g36)) + ((!i_3_) & (!i_4_) & (!sk[55]) & (g28) & (g29) & (g36)) + ((!i_3_) & (!i_4_) & (sk[55]) & (!g28) & (!g29) & (g36)) + ((!i_3_) & (i_4_) & (!sk[55]) & (!g28) & (!g29) & (g36)) + ((!i_3_) & (i_4_) & (!sk[55]) & (!g28) & (g29) & (g36)) + ((!i_3_) & (i_4_) & (!sk[55]) & (g28) & (!g29) & (g36)) + ((!i_3_) & (i_4_) & (!sk[55]) & (g28) & (g29) & (g36)) + ((!i_3_) & (i_4_) & (sk[55]) & (!g28) & (!g29) & (g36)) + ((!i_3_) & (i_4_) & (sk[55]) & (!g28) & (g29) & (g36)) + ((i_3_) & (!i_4_) & (!sk[55]) & (!g28) & (!g29) & (!g36)) + ((i_3_) & (!i_4_) & (!sk[55]) & (!g28) & (!g29) & (g36)) + ((i_3_) & (!i_4_) & (!sk[55]) & (!g28) & (g29) & (!g36)) + ((i_3_) & (!i_4_) & (!sk[55]) & (!g28) & (g29) & (g36)) + ((i_3_) & (!i_4_) & (!sk[55]) & (g28) & (!g29) & (!g36)) + ((i_3_) & (!i_4_) & (!sk[55]) & (g28) & (!g29) & (g36)) + ((i_3_) & (!i_4_) & (!sk[55]) & (g28) & (g29) & (!g36)) + ((i_3_) & (!i_4_) & (!sk[55]) & (g28) & (g29) & (g36)) + ((i_3_) & (!i_4_) & (sk[55]) & (!g28) & (!g29) & (g36)) + ((i_3_) & (!i_4_) & (sk[55]) & (!g28) & (g29) & (g36)) + ((i_3_) & (i_4_) & (!sk[55]) & (!g28) & (!g29) & (!g36)) + ((i_3_) & (i_4_) & (!sk[55]) & (!g28) & (!g29) & (g36)) + ((i_3_) & (i_4_) & (!sk[55]) & (!g28) & (g29) & (!g36)) + ((i_3_) & (i_4_) & (!sk[55]) & (!g28) & (g29) & (g36)) + ((i_3_) & (i_4_) & (!sk[55]) & (g28) & (!g29) & (!g36)) + ((i_3_) & (i_4_) & (!sk[55]) & (g28) & (!g29) & (g36)) + ((i_3_) & (i_4_) & (!sk[55]) & (g28) & (g29) & (!g36)) + ((i_3_) & (i_4_) & (!sk[55]) & (g28) & (g29) & (g36)) + ((i_3_) & (i_4_) & (sk[55]) & (!g28) & (!g29) & (g36)) + ((i_3_) & (i_4_) & (sk[55]) & (!g28) & (g29) & (g36)));
	assign g38 = (((!sk[56]) & (i_8_) & (!g4)) + ((!sk[56]) & (i_8_) & (g4)) + ((sk[56]) & (!i_8_) & (g4)));
	assign g39 = (((!i_5_) & (sk[57]) & (!i_3_) & (i_4_)) + ((i_5_) & (!sk[57]) & (!i_3_) & (!i_4_)) + ((i_5_) & (!sk[57]) & (!i_3_) & (i_4_)) + ((i_5_) & (!sk[57]) & (i_3_) & (!i_4_)) + ((i_5_) & (!sk[57]) & (i_3_) & (i_4_)));
	assign g40 = (((!sk[58]) & (g1) & (!g39)) + ((!sk[58]) & (g1) & (g39)) + ((sk[58]) & (g1) & (g39)));
	assign g41 = (((!sk[59]) & (i_8_) & (!i_7_) & (!g40)) + ((!sk[59]) & (i_8_) & (!i_7_) & (g40)) + ((!sk[59]) & (i_8_) & (i_7_) & (!g40)) + ((!sk[59]) & (i_8_) & (i_7_) & (g40)) + ((sk[59]) & (!i_8_) & (!i_7_) & (g40)));
	assign g42 = (((!sk[60]) & (i_5_) & (!i_3_) & (!g1)) + ((!sk[60]) & (i_5_) & (!i_3_) & (g1)) + ((!sk[60]) & (i_5_) & (i_3_) & (!g1)) + ((!sk[60]) & (i_5_) & (i_3_) & (g1)) + ((sk[60]) & (i_5_) & (!i_3_) & (g1)));
	assign g43 = (((!sk[61]) & (g7) & (!g15)) + ((!sk[61]) & (g7) & (g15)) + ((sk[61]) & (g7) & (!g15)));
	assign g44 = (((!sk[62]) & (g18) & (!g9)) + ((!sk[62]) & (g18) & (g9)) + ((sk[62]) & (!g18) & (g9)));
	assign g45 = (((g6) & (!i_15_) & (!sk[63]) & (!g13)) + ((g6) & (!i_15_) & (!sk[63]) & (g13)) + ((g6) & (i_15_) & (!sk[63]) & (!g13)) + ((g6) & (i_15_) & (!sk[63]) & (g13)) + ((g6) & (i_15_) & (sk[63]) & (g13)));
	assign g46 = (((g6) & (!sk[64]) & (!i_15_) & (!g9)) + ((g6) & (!sk[64]) & (!i_15_) & (g9)) + ((g6) & (!sk[64]) & (i_15_) & (!g9)) + ((g6) & (!sk[64]) & (i_15_) & (g9)) + ((g6) & (sk[64]) & (i_15_) & (g9)));
	assign g47 = (((!g18) & (sk[65]) & (g13)) + ((g18) & (!sk[65]) & (!g13)) + ((g18) & (!sk[65]) & (g13)));
	assign g48 = (((!sk[66]) & (i_14_) & (!i_12_) & (!i_13_)) + ((!sk[66]) & (i_14_) & (!i_12_) & (i_13_)) + ((!sk[66]) & (i_14_) & (i_12_) & (!i_13_)) + ((!sk[66]) & (i_14_) & (i_12_) & (i_13_)) + ((sk[66]) & (!i_14_) & (!i_12_) & (!i_13_)) + ((sk[66]) & (!i_14_) & (!i_12_) & (i_13_)) + ((sk[66]) & (!i_14_) & (i_12_) & (!i_13_)) + ((sk[66]) & (!i_14_) & (i_12_) & (i_13_)) + ((sk[66]) & (i_14_) & (!i_12_) & (!i_13_)) + ((sk[66]) & (i_14_) & (i_12_) & (!i_13_)) + ((sk[66]) & (i_14_) & (i_12_) & (i_13_)));
	assign g49 = (((!i_11_) & (!i_9_) & (!i_10_) & (!i_12_) & (!sk[67]) & (g48)) + ((!i_11_) & (!i_9_) & (!i_10_) & (i_12_) & (!sk[67]) & (g48)) + ((!i_11_) & (!i_9_) & (i_10_) & (!i_12_) & (!sk[67]) & (g48)) + ((!i_11_) & (!i_9_) & (i_10_) & (!i_12_) & (sk[67]) & (!g48)) + ((!i_11_) & (!i_9_) & (i_10_) & (i_12_) & (!sk[67]) & (g48)) + ((!i_11_) & (!i_9_) & (i_10_) & (i_12_) & (sk[67]) & (!g48)) + ((!i_11_) & (!i_9_) & (i_10_) & (i_12_) & (sk[67]) & (g48)) + ((!i_11_) & (i_9_) & (!i_10_) & (!i_12_) & (!sk[67]) & (g48)) + ((!i_11_) & (i_9_) & (!i_10_) & (!i_12_) & (sk[67]) & (!g48)) + ((!i_11_) & (i_9_) & (!i_10_) & (i_12_) & (!sk[67]) & (g48)) + ((!i_11_) & (i_9_) & (!i_10_) & (i_12_) & (sk[67]) & (!g48)) + ((!i_11_) & (i_9_) & (!i_10_) & (i_12_) & (sk[67]) & (g48)) + ((!i_11_) & (i_9_) & (i_10_) & (!i_12_) & (!sk[67]) & (g48)) + ((!i_11_) & (i_9_) & (i_10_) & (i_12_) & (!sk[67]) & (g48)) + ((i_11_) & (!i_9_) & (!i_10_) & (!i_12_) & (!sk[67]) & (!g48)) + ((i_11_) & (!i_9_) & (!i_10_) & (!i_12_) & (!sk[67]) & (g48)) + ((i_11_) & (!i_9_) & (!i_10_) & (i_12_) & (!sk[67]) & (!g48)) + ((i_11_) & (!i_9_) & (!i_10_) & (i_12_) & (!sk[67]) & (g48)) + ((i_11_) & (!i_9_) & (i_10_) & (!i_12_) & (!sk[67]) & (!g48)) + ((i_11_) & (!i_9_) & (i_10_) & (!i_12_) & (!sk[67]) & (g48)) + ((i_11_) & (!i_9_) & (i_10_) & (!i_12_) & (sk[67]) & (!g48)) + ((i_11_) & (!i_9_) & (i_10_) & (!i_12_) & (sk[67]) & (g48)) + ((i_11_) & (!i_9_) & (i_10_) & (i_12_) & (!sk[67]) & (!g48)) + ((i_11_) & (!i_9_) & (i_10_) & (i_12_) & (!sk[67]) & (g48)) + ((i_11_) & (!i_9_) & (i_10_) & (i_12_) & (sk[67]) & (!g48)) + ((i_11_) & (!i_9_) & (i_10_) & (i_12_) & (sk[67]) & (g48)) + ((i_11_) & (i_9_) & (!i_10_) & (!i_12_) & (!sk[67]) & (!g48)) + ((i_11_) & (i_9_) & (!i_10_) & (!i_12_) & (!sk[67]) & (g48)) + ((i_11_) & (i_9_) & (!i_10_) & (!i_12_) & (sk[67]) & (!g48)) + ((i_11_) & (i_9_) & (!i_10_) & (!i_12_) & (sk[67]) & (g48)) + ((i_11_) & (i_9_) & (!i_10_) & (i_12_) & (!sk[67]) & (!g48)) + ((i_11_) & (i_9_) & (!i_10_) & (i_12_) & (!sk[67]) & (g48)) + ((i_11_) & (i_9_) & (!i_10_) & (i_12_) & (sk[67]) & (!g48)) + ((i_11_) & (i_9_) & (!i_10_) & (i_12_) & (sk[67]) & (g48)) + ((i_11_) & (i_9_) & (i_10_) & (!i_12_) & (!sk[67]) & (!g48)) + ((i_11_) & (i_9_) & (i_10_) & (!i_12_) & (!sk[67]) & (g48)) + ((i_11_) & (i_9_) & (i_10_) & (i_12_) & (!sk[67]) & (!g48)) + ((i_11_) & (i_9_) & (i_10_) & (i_12_) & (!sk[67]) & (g48)));
	assign g50 = (((!sk[68]) & (!g44) & (!g45) & (!g46) & (!g47) & (g49)) + ((!sk[68]) & (!g44) & (!g45) & (!g46) & (g47) & (g49)) + ((!sk[68]) & (!g44) & (!g45) & (g46) & (!g47) & (g49)) + ((!sk[68]) & (!g44) & (!g45) & (g46) & (g47) & (g49)) + ((!sk[68]) & (!g44) & (g45) & (!g46) & (!g47) & (g49)) + ((!sk[68]) & (!g44) & (g45) & (!g46) & (g47) & (g49)) + ((!sk[68]) & (!g44) & (g45) & (g46) & (!g47) & (g49)) + ((!sk[68]) & (!g44) & (g45) & (g46) & (g47) & (g49)) + ((!sk[68]) & (g44) & (!g45) & (!g46) & (!g47) & (!g49)) + ((!sk[68]) & (g44) & (!g45) & (!g46) & (!g47) & (g49)) + ((!sk[68]) & (g44) & (!g45) & (!g46) & (g47) & (!g49)) + ((!sk[68]) & (g44) & (!g45) & (!g46) & (g47) & (g49)) + ((!sk[68]) & (g44) & (!g45) & (g46) & (!g47) & (!g49)) + ((!sk[68]) & (g44) & (!g45) & (g46) & (!g47) & (g49)) + ((!sk[68]) & (g44) & (!g45) & (g46) & (g47) & (!g49)) + ((!sk[68]) & (g44) & (!g45) & (g46) & (g47) & (g49)) + ((!sk[68]) & (g44) & (g45) & (!g46) & (!g47) & (!g49)) + ((!sk[68]) & (g44) & (g45) & (!g46) & (!g47) & (g49)) + ((!sk[68]) & (g44) & (g45) & (!g46) & (g47) & (!g49)) + ((!sk[68]) & (g44) & (g45) & (!g46) & (g47) & (g49)) + ((!sk[68]) & (g44) & (g45) & (g46) & (!g47) & (!g49)) + ((!sk[68]) & (g44) & (g45) & (g46) & (!g47) & (g49)) + ((!sk[68]) & (g44) & (g45) & (g46) & (g47) & (!g49)) + ((!sk[68]) & (g44) & (g45) & (g46) & (g47) & (g49)) + ((sk[68]) & (!g44) & (!g45) & (!g46) & (!g47) & (!g49)));
	assign g51 = (((!g38) & (!g41) & (!sk[69]) & (!g42) & (!g43) & (g50)) + ((!g38) & (!g41) & (!sk[69]) & (!g42) & (g43) & (g50)) + ((!g38) & (!g41) & (!sk[69]) & (g42) & (!g43) & (g50)) + ((!g38) & (!g41) & (!sk[69]) & (g42) & (g43) & (g50)) + ((!g38) & (g41) & (!sk[69]) & (!g42) & (!g43) & (g50)) + ((!g38) & (g41) & (!sk[69]) & (!g42) & (g43) & (g50)) + ((!g38) & (g41) & (!sk[69]) & (g42) & (!g43) & (g50)) + ((!g38) & (g41) & (!sk[69]) & (g42) & (g43) & (g50)) + ((!g38) & (g41) & (sk[69]) & (!g42) & (!g43) & (!g50)) + ((!g38) & (g41) & (sk[69]) & (!g42) & (g43) & (!g50)) + ((!g38) & (g41) & (sk[69]) & (!g42) & (g43) & (g50)) + ((!g38) & (g41) & (sk[69]) & (g42) & (!g43) & (!g50)) + ((!g38) & (g41) & (sk[69]) & (g42) & (g43) & (!g50)) + ((!g38) & (g41) & (sk[69]) & (g42) & (g43) & (g50)) + ((g38) & (!g41) & (!sk[69]) & (!g42) & (!g43) & (!g50)) + ((g38) & (!g41) & (!sk[69]) & (!g42) & (!g43) & (g50)) + ((g38) & (!g41) & (!sk[69]) & (!g42) & (g43) & (!g50)) + ((g38) & (!g41) & (!sk[69]) & (!g42) & (g43) & (g50)) + ((g38) & (!g41) & (!sk[69]) & (g42) & (!g43) & (!g50)) + ((g38) & (!g41) & (!sk[69]) & (g42) & (!g43) & (g50)) + ((g38) & (!g41) & (!sk[69]) & (g42) & (g43) & (!g50)) + ((g38) & (!g41) & (!sk[69]) & (g42) & (g43) & (g50)) + ((g38) & (!g41) & (sk[69]) & (g42) & (!g43) & (!g50)) + ((g38) & (!g41) & (sk[69]) & (g42) & (g43) & (!g50)) + ((g38) & (!g41) & (sk[69]) & (g42) & (g43) & (g50)) + ((g38) & (g41) & (!sk[69]) & (!g42) & (!g43) & (!g50)) + ((g38) & (g41) & (!sk[69]) & (!g42) & (!g43) & (g50)) + ((g38) & (g41) & (!sk[69]) & (!g42) & (g43) & (!g50)) + ((g38) & (g41) & (!sk[69]) & (!g42) & (g43) & (g50)) + ((g38) & (g41) & (!sk[69]) & (g42) & (!g43) & (!g50)) + ((g38) & (g41) & (!sk[69]) & (g42) & (!g43) & (g50)) + ((g38) & (g41) & (!sk[69]) & (g42) & (g43) & (!g50)) + ((g38) & (g41) & (!sk[69]) & (g42) & (g43) & (g50)) + ((g38) & (g41) & (sk[69]) & (!g42) & (!g43) & (!g50)) + ((g38) & (g41) & (sk[69]) & (!g42) & (g43) & (!g50)) + ((g38) & (g41) & (sk[69]) & (!g42) & (g43) & (g50)) + ((g38) & (g41) & (sk[69]) & (g42) & (!g43) & (!g50)) + ((g38) & (g41) & (sk[69]) & (g42) & (g43) & (!g50)) + ((g38) & (g41) & (sk[69]) & (g42) & (g43) & (g50)));
	assign g52 = (((i_5_) & (!i_3_) & (!sk[70]) & (!i_4_)) + ((i_5_) & (!i_3_) & (!sk[70]) & (i_4_)) + ((i_5_) & (!i_3_) & (sk[70]) & (!i_4_)) + ((i_5_) & (i_3_) & (!sk[70]) & (!i_4_)) + ((i_5_) & (i_3_) & (!sk[70]) & (i_4_)));
	assign g53 = (((!sk[71]) & (i_11_) & (!i_15_)) + ((!sk[71]) & (i_11_) & (i_15_)) + ((sk[71]) & (!i_11_) & (!i_15_)));
	assign g54 = (((!i_9_) & (!i_10_) & (!g7) & (!i_4_) & (!sk[72]) & (g53)) + ((!i_9_) & (!i_10_) & (!g7) & (i_4_) & (!sk[72]) & (g53)) + ((!i_9_) & (!i_10_) & (g7) & (!i_4_) & (!sk[72]) & (g53)) + ((!i_9_) & (!i_10_) & (g7) & (!i_4_) & (sk[72]) & (g53)) + ((!i_9_) & (!i_10_) & (g7) & (i_4_) & (!sk[72]) & (g53)) + ((!i_9_) & (i_10_) & (!g7) & (!i_4_) & (!sk[72]) & (g53)) + ((!i_9_) & (i_10_) & (!g7) & (i_4_) & (!sk[72]) & (g53)) + ((!i_9_) & (i_10_) & (g7) & (!i_4_) & (!sk[72]) & (g53)) + ((!i_9_) & (i_10_) & (g7) & (!i_4_) & (sk[72]) & (g53)) + ((!i_9_) & (i_10_) & (g7) & (i_4_) & (!sk[72]) & (g53)) + ((!i_9_) & (i_10_) & (g7) & (i_4_) & (sk[72]) & (g53)) + ((i_9_) & (!i_10_) & (!g7) & (!i_4_) & (!sk[72]) & (!g53)) + ((i_9_) & (!i_10_) & (!g7) & (!i_4_) & (!sk[72]) & (g53)) + ((i_9_) & (!i_10_) & (!g7) & (i_4_) & (!sk[72]) & (!g53)) + ((i_9_) & (!i_10_) & (!g7) & (i_4_) & (!sk[72]) & (g53)) + ((i_9_) & (!i_10_) & (g7) & (!i_4_) & (!sk[72]) & (!g53)) + ((i_9_) & (!i_10_) & (g7) & (!i_4_) & (!sk[72]) & (g53)) + ((i_9_) & (!i_10_) & (g7) & (!i_4_) & (sk[72]) & (g53)) + ((i_9_) & (!i_10_) & (g7) & (i_4_) & (!sk[72]) & (!g53)) + ((i_9_) & (!i_10_) & (g7) & (i_4_) & (!sk[72]) & (g53)) + ((i_9_) & (!i_10_) & (g7) & (i_4_) & (sk[72]) & (g53)) + ((i_9_) & (i_10_) & (!g7) & (!i_4_) & (!sk[72]) & (!g53)) + ((i_9_) & (i_10_) & (!g7) & (!i_4_) & (!sk[72]) & (g53)) + ((i_9_) & (i_10_) & (!g7) & (i_4_) & (!sk[72]) & (!g53)) + ((i_9_) & (i_10_) & (!g7) & (i_4_) & (!sk[72]) & (g53)) + ((i_9_) & (i_10_) & (g7) & (!i_4_) & (!sk[72]) & (!g53)) + ((i_9_) & (i_10_) & (g7) & (!i_4_) & (!sk[72]) & (g53)) + ((i_9_) & (i_10_) & (g7) & (i_4_) & (!sk[72]) & (!g53)) + ((i_9_) & (i_10_) & (g7) & (i_4_) & (!sk[72]) & (g53)));
	assign g55 = (((!i_5_) & (!sk[73]) & (i_3_) & (i_8_) & (!i_7_)) + ((!i_5_) & (!sk[73]) & (i_3_) & (i_8_) & (i_7_)) + ((!i_5_) & (sk[73]) & (!i_3_) & (i_8_) & (!i_7_)) + ((i_5_) & (!sk[73]) & (!i_3_) & (!i_8_) & (!i_7_)) + ((i_5_) & (!sk[73]) & (!i_3_) & (!i_8_) & (i_7_)) + ((i_5_) & (!sk[73]) & (!i_3_) & (i_8_) & (!i_7_)) + ((i_5_) & (!sk[73]) & (!i_3_) & (i_8_) & (i_7_)) + ((i_5_) & (!sk[73]) & (i_3_) & (!i_8_) & (!i_7_)) + ((i_5_) & (!sk[73]) & (i_3_) & (!i_8_) & (i_7_)) + ((i_5_) & (!sk[73]) & (i_3_) & (i_8_) & (!i_7_)) + ((i_5_) & (!sk[73]) & (i_3_) & (i_8_) & (i_7_)));
	assign g56 = (((!sk[74]) & (!i_0_) & (g52) & (g54) & (!g55)) + ((!sk[74]) & (!i_0_) & (g52) & (g54) & (g55)) + ((!sk[74]) & (i_0_) & (!g52) & (!g54) & (!g55)) + ((!sk[74]) & (i_0_) & (!g52) & (!g54) & (g55)) + ((!sk[74]) & (i_0_) & (!g52) & (g54) & (!g55)) + ((!sk[74]) & (i_0_) & (!g52) & (g54) & (g55)) + ((!sk[74]) & (i_0_) & (g52) & (!g54) & (!g55)) + ((!sk[74]) & (i_0_) & (g52) & (!g54) & (g55)) + ((!sk[74]) & (i_0_) & (g52) & (g54) & (!g55)) + ((!sk[74]) & (i_0_) & (g52) & (g54) & (g55)) + ((sk[74]) & (!i_0_) & (!g52) & (!g54) & (g55)) + ((sk[74]) & (!i_0_) & (g52) & (!g54) & (g55)) + ((sk[74]) & (i_0_) & (!g52) & (!g54) & (!g55)) + ((sk[74]) & (i_0_) & (!g52) & (!g54) & (g55)) + ((sk[74]) & (i_0_) & (!g52) & (g54) & (!g55)) + ((sk[74]) & (i_0_) & (!g52) & (g54) & (g55)) + ((sk[74]) & (i_0_) & (g52) & (!g54) & (g55)));
	assign g57 = (((!i_1_) & (sk[75]) & (!i_0_) & (!i_2_)) + ((i_1_) & (!sk[75]) & (!i_0_) & (!i_2_)) + ((i_1_) & (!sk[75]) & (!i_0_) & (i_2_)) + ((i_1_) & (!sk[75]) & (i_0_) & (!i_2_)) + ((i_1_) & (!sk[75]) & (i_0_) & (i_2_)));
	assign g58 = (((!i_5_) & (!i_3_) & (!i_4_) & (sk[76]) & (g57)) + ((!i_5_) & (i_3_) & (i_4_) & (!sk[76]) & (!g57)) + ((!i_5_) & (i_3_) & (i_4_) & (!sk[76]) & (g57)) + ((i_5_) & (!i_3_) & (!i_4_) & (!sk[76]) & (!g57)) + ((i_5_) & (!i_3_) & (!i_4_) & (!sk[76]) & (g57)) + ((i_5_) & (!i_3_) & (i_4_) & (!sk[76]) & (!g57)) + ((i_5_) & (!i_3_) & (i_4_) & (!sk[76]) & (g57)) + ((i_5_) & (i_3_) & (!i_4_) & (!sk[76]) & (!g57)) + ((i_5_) & (i_3_) & (!i_4_) & (!sk[76]) & (g57)) + ((i_5_) & (i_3_) & (i_4_) & (!sk[76]) & (!g57)) + ((i_5_) & (i_3_) & (i_4_) & (!sk[76]) & (g57)));
	assign g59 = (((g58) & (!sk[77]) & (!g38)) + ((g58) & (!sk[77]) & (g38)) + ((g58) & (sk[77]) & (g38)));
	assign g60 = (((!sk[78]) & (!i_11_) & (i_12_) & (g59) & (!g41)) + ((!sk[78]) & (!i_11_) & (i_12_) & (g59) & (g41)) + ((!sk[78]) & (i_11_) & (!i_12_) & (!g59) & (!g41)) + ((!sk[78]) & (i_11_) & (!i_12_) & (!g59) & (g41)) + ((!sk[78]) & (i_11_) & (!i_12_) & (g59) & (!g41)) + ((!sk[78]) & (i_11_) & (!i_12_) & (g59) & (g41)) + ((!sk[78]) & (i_11_) & (i_12_) & (!g59) & (!g41)) + ((!sk[78]) & (i_11_) & (i_12_) & (!g59) & (g41)) + ((!sk[78]) & (i_11_) & (i_12_) & (g59) & (!g41)) + ((!sk[78]) & (i_11_) & (i_12_) & (g59) & (g41)) + ((sk[78]) & (!i_11_) & (!i_12_) & (!g59) & (!g41)) + ((sk[78]) & (!i_11_) & (!i_12_) & (!g59) & (g41)) + ((sk[78]) & (!i_11_) & (i_12_) & (!g59) & (!g41)) + ((sk[78]) & (i_11_) & (!i_12_) & (!g59) & (!g41)) + ((sk[78]) & (i_11_) & (!i_12_) & (!g59) & (g41)) + ((sk[78]) & (i_11_) & (i_12_) & (!g59) & (!g41)) + ((sk[78]) & (i_11_) & (i_12_) & (!g59) & (g41)));
	assign g61 = (((!i_5_) & (!sk[79]) & (i_3_) & (i_4_) & (!g1)) + ((!i_5_) & (!sk[79]) & (i_3_) & (i_4_) & (g1)) + ((!i_5_) & (sk[79]) & (i_3_) & (i_4_) & (g1)) + ((i_5_) & (!sk[79]) & (!i_3_) & (!i_4_) & (!g1)) + ((i_5_) & (!sk[79]) & (!i_3_) & (!i_4_) & (g1)) + ((i_5_) & (!sk[79]) & (!i_3_) & (i_4_) & (!g1)) + ((i_5_) & (!sk[79]) & (!i_3_) & (i_4_) & (g1)) + ((i_5_) & (!sk[79]) & (i_3_) & (!i_4_) & (!g1)) + ((i_5_) & (!sk[79]) & (i_3_) & (!i_4_) & (g1)) + ((i_5_) & (!sk[79]) & (i_3_) & (i_4_) & (!g1)) + ((i_5_) & (!sk[79]) & (i_3_) & (i_4_) & (g1)));
	assign g62 = (((!i_5_) & (!sk[80]) & (i_3_) & (i_4_) & (!g1)) + ((!i_5_) & (!sk[80]) & (i_3_) & (i_4_) & (g1)) + ((!i_5_) & (sk[80]) & (i_3_) & (!i_4_) & (g1)) + ((i_5_) & (!sk[80]) & (!i_3_) & (!i_4_) & (!g1)) + ((i_5_) & (!sk[80]) & (!i_3_) & (!i_4_) & (g1)) + ((i_5_) & (!sk[80]) & (!i_3_) & (i_4_) & (!g1)) + ((i_5_) & (!sk[80]) & (!i_3_) & (i_4_) & (g1)) + ((i_5_) & (!sk[80]) & (i_3_) & (!i_4_) & (!g1)) + ((i_5_) & (!sk[80]) & (i_3_) & (!i_4_) & (g1)) + ((i_5_) & (!sk[80]) & (i_3_) & (i_4_) & (!g1)) + ((i_5_) & (!sk[80]) & (i_3_) & (i_4_) & (g1)));
	assign g63 = (((g31) & (!sk[81]) & (!g61) & (!g62)) + ((g31) & (!sk[81]) & (!g61) & (g62)) + ((g31) & (!sk[81]) & (g61) & (!g62)) + ((g31) & (!sk[81]) & (g61) & (g62)) + ((g31) & (sk[81]) & (!g61) & (g62)) + ((g31) & (sk[81]) & (g61) & (!g62)) + ((g31) & (sk[81]) & (g61) & (g62)));
	assign g64 = (((!i_5_) & (i_3_) & (!sk[82]) & (i_4_) & (!g1)) + ((!i_5_) & (i_3_) & (!sk[82]) & (i_4_) & (g1)) + ((i_5_) & (!i_3_) & (!sk[82]) & (!i_4_) & (!g1)) + ((i_5_) & (!i_3_) & (!sk[82]) & (!i_4_) & (g1)) + ((i_5_) & (!i_3_) & (!sk[82]) & (i_4_) & (!g1)) + ((i_5_) & (!i_3_) & (!sk[82]) & (i_4_) & (g1)) + ((i_5_) & (!i_3_) & (sk[82]) & (i_4_) & (g1)) + ((i_5_) & (i_3_) & (!sk[82]) & (!i_4_) & (!g1)) + ((i_5_) & (i_3_) & (!sk[82]) & (!i_4_) & (g1)) + ((i_5_) & (i_3_) & (!sk[82]) & (i_4_) & (!g1)) + ((i_5_) & (i_3_) & (!sk[82]) & (i_4_) & (g1)));
	assign g65 = (((!sk[83]) & (g1) & (!g52)) + ((!sk[83]) & (g1) & (g52)) + ((sk[83]) & (g1) & (g52)));
	assign g66 = (((!sk[84]) & (g6) & (!i_15_) & (!g7)) + ((!sk[84]) & (g6) & (!i_15_) & (g7)) + ((!sk[84]) & (g6) & (i_15_) & (!g7)) + ((!sk[84]) & (g6) & (i_15_) & (g7)) + ((sk[84]) & (g6) & (!i_15_) & (g7)));
	assign g67 = (((!i_9_) & (i_10_) & (sk[85]) & (!g66)) + ((i_9_) & (!i_10_) & (!sk[85]) & (!g66)) + ((i_9_) & (!i_10_) & (!sk[85]) & (g66)) + ((i_9_) & (!i_10_) & (sk[85]) & (!g66)) + ((i_9_) & (i_10_) & (!sk[85]) & (!g66)) + ((i_9_) & (i_10_) & (!sk[85]) & (g66)));
	assign g68 = (((!sk[86]) & (i_3_) & (!i_1_) & (!i_0_)) + ((!sk[86]) & (i_3_) & (!i_1_) & (i_0_)) + ((!sk[86]) & (i_3_) & (i_1_) & (!i_0_)) + ((!sk[86]) & (i_3_) & (i_1_) & (i_0_)) + ((sk[86]) & (!i_3_) & (!i_1_) & (!i_0_)) + ((sk[86]) & (!i_3_) & (!i_1_) & (i_0_)) + ((sk[86]) & (!i_3_) & (i_1_) & (!i_0_)) + ((sk[86]) & (!i_3_) & (i_1_) & (i_0_)) + ((sk[86]) & (i_3_) & (!i_1_) & (i_0_)) + ((sk[86]) & (i_3_) & (i_1_) & (!i_0_)) + ((sk[86]) & (i_3_) & (i_1_) & (i_0_)));
	assign g69 = (((!i_8_) & (!i_6_) & (!g64) & (!g65) & (!sk[87]) & (g68)) + ((!i_8_) & (!i_6_) & (!g64) & (!g65) & (sk[87]) & (g68)) + ((!i_8_) & (!i_6_) & (!g64) & (g65) & (!sk[87]) & (g68)) + ((!i_8_) & (!i_6_) & (!g64) & (g65) & (sk[87]) & (g68)) + ((!i_8_) & (!i_6_) & (g64) & (!g65) & (!sk[87]) & (g68)) + ((!i_8_) & (!i_6_) & (g64) & (!g65) & (sk[87]) & (g68)) + ((!i_8_) & (!i_6_) & (g64) & (g65) & (!sk[87]) & (g68)) + ((!i_8_) & (!i_6_) & (g64) & (g65) & (sk[87]) & (g68)) + ((!i_8_) & (i_6_) & (!g64) & (!g65) & (!sk[87]) & (g68)) + ((!i_8_) & (i_6_) & (!g64) & (!g65) & (sk[87]) & (g68)) + ((!i_8_) & (i_6_) & (!g64) & (g65) & (!sk[87]) & (g68)) + ((!i_8_) & (i_6_) & (!g64) & (g65) & (sk[87]) & (g68)) + ((!i_8_) & (i_6_) & (g64) & (!g65) & (!sk[87]) & (g68)) + ((!i_8_) & (i_6_) & (g64) & (!g65) & (sk[87]) & (g68)) + ((!i_8_) & (i_6_) & (g64) & (g65) & (!sk[87]) & (g68)) + ((!i_8_) & (i_6_) & (g64) & (g65) & (sk[87]) & (g68)) + ((i_8_) & (!i_6_) & (!g64) & (!g65) & (!sk[87]) & (!g68)) + ((i_8_) & (!i_6_) & (!g64) & (!g65) & (!sk[87]) & (g68)) + ((i_8_) & (!i_6_) & (!g64) & (!g65) & (sk[87]) & (g68)) + ((i_8_) & (!i_6_) & (!g64) & (g65) & (!sk[87]) & (!g68)) + ((i_8_) & (!i_6_) & (!g64) & (g65) & (!sk[87]) & (g68)) + ((i_8_) & (!i_6_) & (!g64) & (g65) & (sk[87]) & (g68)) + ((i_8_) & (!i_6_) & (g64) & (!g65) & (!sk[87]) & (!g68)) + ((i_8_) & (!i_6_) & (g64) & (!g65) & (!sk[87]) & (g68)) + ((i_8_) & (!i_6_) & (g64) & (!g65) & (sk[87]) & (g68)) + ((i_8_) & (!i_6_) & (g64) & (g65) & (!sk[87]) & (!g68)) + ((i_8_) & (!i_6_) & (g64) & (g65) & (!sk[87]) & (g68)) + ((i_8_) & (!i_6_) & (g64) & (g65) & (sk[87]) & (g68)) + ((i_8_) & (i_6_) & (!g64) & (!g65) & (!sk[87]) & (!g68)) + ((i_8_) & (i_6_) & (!g64) & (!g65) & (!sk[87]) & (g68)) + ((i_8_) & (i_6_) & (!g64) & (!g65) & (sk[87]) & (g68)) + ((i_8_) & (i_6_) & (!g64) & (g65) & (!sk[87]) & (!g68)) + ((i_8_) & (i_6_) & (!g64) & (g65) & (!sk[87]) & (g68)) + ((i_8_) & (i_6_) & (g64) & (!g65) & (!sk[87]) & (!g68)) + ((i_8_) & (i_6_) & (g64) & (!g65) & (!sk[87]) & (g68)) + ((i_8_) & (i_6_) & (g64) & (g65) & (!sk[87]) & (!g68)) + ((i_8_) & (i_6_) & (g64) & (g65) & (!sk[87]) & (g68)));
	assign g70 = (((!i_11_) & (!i_9_) & (!i_10_) & (sk[88]) & (!g59) & (g69)) + ((!i_11_) & (!i_9_) & (!i_10_) & (sk[88]) & (g59) & (g69)) + ((!i_11_) & (!i_9_) & (i_10_) & (sk[88]) & (!g59) & (g69)) + ((!i_11_) & (!i_9_) & (i_10_) & (sk[88]) & (g59) & (g69)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[88]) & (!g59) & (g69)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[88]) & (g59) & (g69)) + ((!i_11_) & (i_9_) & (!i_10_) & (sk[88]) & (!g59) & (g69)) + ((!i_11_) & (i_9_) & (!i_10_) & (sk[88]) & (g59) & (g69)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[88]) & (!g59) & (!g69)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[88]) & (!g59) & (g69)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[88]) & (g59) & (!g69)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[88]) & (g59) & (g69)) + ((!i_11_) & (i_9_) & (i_10_) & (sk[88]) & (!g59) & (g69)) + ((!i_11_) & (i_9_) & (i_10_) & (sk[88]) & (g59) & (g69)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[88]) & (g59) & (!g69)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[88]) & (g59) & (g69)) + ((i_11_) & (!i_9_) & (!i_10_) & (sk[88]) & (!g59) & (g69)) + ((i_11_) & (!i_9_) & (!i_10_) & (sk[88]) & (g59) & (g69)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[88]) & (g59) & (!g69)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[88]) & (g59) & (g69)) + ((i_11_) & (!i_9_) & (i_10_) & (sk[88]) & (!g59) & (g69)) + ((i_11_) & (!i_9_) & (i_10_) & (sk[88]) & (g59) & (g69)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[88]) & (!g59) & (g69)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[88]) & (g59) & (!g69)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[88]) & (g59) & (g69)) + ((i_11_) & (i_9_) & (!i_10_) & (sk[88]) & (!g59) & (g69)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[88]) & (!g59) & (!g69)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[88]) & (!g59) & (g69)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[88]) & (g59) & (!g69)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[88]) & (g59) & (g69)) + ((i_11_) & (i_9_) & (i_10_) & (sk[88]) & (!g59) & (g69)) + ((i_11_) & (i_9_) & (i_10_) & (sk[88]) & (g59) & (g69)));
	assign g71 = (((!g38) & (!g64) & (!g65) & (sk[89]) & (!g67) & (g70)) + ((!g38) & (!g64) & (!g65) & (sk[89]) & (g67) & (g70)) + ((!g38) & (!g64) & (g65) & (sk[89]) & (!g67) & (g70)) + ((!g38) & (!g64) & (g65) & (sk[89]) & (g67) & (g70)) + ((!g38) & (g64) & (!g65) & (!sk[89]) & (!g67) & (g70)) + ((!g38) & (g64) & (!g65) & (!sk[89]) & (g67) & (g70)) + ((!g38) & (g64) & (!g65) & (sk[89]) & (!g67) & (g70)) + ((!g38) & (g64) & (!g65) & (sk[89]) & (g67) & (g70)) + ((!g38) & (g64) & (g65) & (!sk[89]) & (!g67) & (!g70)) + ((!g38) & (g64) & (g65) & (!sk[89]) & (!g67) & (g70)) + ((!g38) & (g64) & (g65) & (!sk[89]) & (g67) & (!g70)) + ((!g38) & (g64) & (g65) & (!sk[89]) & (g67) & (g70)) + ((!g38) & (g64) & (g65) & (sk[89]) & (!g67) & (g70)) + ((!g38) & (g64) & (g65) & (sk[89]) & (g67) & (g70)) + ((g38) & (!g64) & (!g65) & (!sk[89]) & (g67) & (!g70)) + ((g38) & (!g64) & (!g65) & (!sk[89]) & (g67) & (g70)) + ((g38) & (!g64) & (!g65) & (sk[89]) & (!g67) & (g70)) + ((g38) & (!g64) & (!g65) & (sk[89]) & (g67) & (g70)) + ((g38) & (!g64) & (g65) & (!sk[89]) & (g67) & (!g70)) + ((g38) & (!g64) & (g65) & (!sk[89]) & (g67) & (g70)) + ((g38) & (!g64) & (g65) & (sk[89]) & (g67) & (g70)) + ((g38) & (g64) & (!g65) & (!sk[89]) & (!g67) & (g70)) + ((g38) & (g64) & (!g65) & (!sk[89]) & (g67) & (!g70)) + ((g38) & (g64) & (!g65) & (!sk[89]) & (g67) & (g70)) + ((g38) & (g64) & (!g65) & (sk[89]) & (g67) & (g70)) + ((g38) & (g64) & (g65) & (!sk[89]) & (!g67) & (!g70)) + ((g38) & (g64) & (g65) & (!sk[89]) & (!g67) & (g70)) + ((g38) & (g64) & (g65) & (!sk[89]) & (g67) & (!g70)) + ((g38) & (g64) & (g65) & (!sk[89]) & (g67) & (g70)) + ((g38) & (g64) & (g65) & (sk[89]) & (g67) & (g70)));
	assign g72 = (((!i_9_) & (!i_10_) & (!sk[90]) & (!g60) & (g63) & (!g71)) + ((!i_9_) & (!i_10_) & (!sk[90]) & (!g60) & (g63) & (g71)) + ((!i_9_) & (!i_10_) & (!sk[90]) & (g60) & (!g63) & (!g71)) + ((!i_9_) & (!i_10_) & (!sk[90]) & (g60) & (!g63) & (g71)) + ((!i_9_) & (!i_10_) & (!sk[90]) & (g60) & (g63) & (!g71)) + ((!i_9_) & (!i_10_) & (!sk[90]) & (g60) & (g63) & (g71)) + ((!i_9_) & (!i_10_) & (sk[90]) & (!g60) & (!g63) & (g71)) + ((!i_9_) & (!i_10_) & (sk[90]) & (g60) & (!g63) & (g71)) + ((!i_9_) & (i_10_) & (!sk[90]) & (!g60) & (!g63) & (!g71)) + ((!i_9_) & (i_10_) & (!sk[90]) & (!g60) & (!g63) & (g71)) + ((!i_9_) & (i_10_) & (!sk[90]) & (!g60) & (g63) & (!g71)) + ((!i_9_) & (i_10_) & (!sk[90]) & (!g60) & (g63) & (g71)) + ((!i_9_) & (i_10_) & (!sk[90]) & (g60) & (!g63) & (!g71)) + ((!i_9_) & (i_10_) & (!sk[90]) & (g60) & (!g63) & (g71)) + ((!i_9_) & (i_10_) & (!sk[90]) & (g60) & (g63) & (!g71)) + ((!i_9_) & (i_10_) & (!sk[90]) & (g60) & (g63) & (g71)) + ((!i_9_) & (i_10_) & (sk[90]) & (!g60) & (!g63) & (g71)) + ((!i_9_) & (i_10_) & (sk[90]) & (!g60) & (g63) & (g71)) + ((!i_9_) & (i_10_) & (sk[90]) & (g60) & (!g63) & (g71)) + ((!i_9_) & (i_10_) & (sk[90]) & (g60) & (g63) & (g71)) + ((i_9_) & (!i_10_) & (!sk[90]) & (!g60) & (!g63) & (!g71)) + ((i_9_) & (!i_10_) & (!sk[90]) & (!g60) & (!g63) & (g71)) + ((i_9_) & (!i_10_) & (!sk[90]) & (!g60) & (g63) & (!g71)) + ((i_9_) & (!i_10_) & (!sk[90]) & (!g60) & (g63) & (g71)) + ((i_9_) & (!i_10_) & (!sk[90]) & (g60) & (!g63) & (!g71)) + ((i_9_) & (!i_10_) & (!sk[90]) & (g60) & (!g63) & (g71)) + ((i_9_) & (!i_10_) & (!sk[90]) & (g60) & (g63) & (!g71)) + ((i_9_) & (!i_10_) & (!sk[90]) & (g60) & (g63) & (g71)) + ((i_9_) & (!i_10_) & (sk[90]) & (!g60) & (!g63) & (g71)) + ((i_9_) & (!i_10_) & (sk[90]) & (!g60) & (g63) & (g71)) + ((i_9_) & (!i_10_) & (sk[90]) & (g60) & (!g63) & (g71)) + ((i_9_) & (!i_10_) & (sk[90]) & (g60) & (g63) & (g71)) + ((i_9_) & (i_10_) & (!sk[90]) & (!g60) & (!g63) & (!g71)) + ((i_9_) & (i_10_) & (!sk[90]) & (!g60) & (!g63) & (g71)) + ((i_9_) & (i_10_) & (!sk[90]) & (!g60) & (g63) & (!g71)) + ((i_9_) & (i_10_) & (!sk[90]) & (!g60) & (g63) & (g71)) + ((i_9_) & (i_10_) & (!sk[90]) & (g60) & (!g63) & (!g71)) + ((i_9_) & (i_10_) & (!sk[90]) & (g60) & (!g63) & (g71)) + ((i_9_) & (i_10_) & (!sk[90]) & (g60) & (g63) & (!g71)) + ((i_9_) & (i_10_) & (!sk[90]) & (g60) & (g63) & (g71)) + ((i_9_) & (i_10_) & (sk[90]) & (g60) & (!g63) & (g71)));
	assign g73 = (((!i_1_) & (!i_2_) & (!g51) & (!sk[91]) & (g56) & (!g72)) + ((!i_1_) & (!i_2_) & (!g51) & (!sk[91]) & (g56) & (g72)) + ((!i_1_) & (!i_2_) & (!g51) & (sk[91]) & (!g56) & (g72)) + ((!i_1_) & (!i_2_) & (!g51) & (sk[91]) & (g56) & (g72)) + ((!i_1_) & (!i_2_) & (g51) & (!sk[91]) & (!g56) & (!g72)) + ((!i_1_) & (!i_2_) & (g51) & (!sk[91]) & (!g56) & (g72)) + ((!i_1_) & (!i_2_) & (g51) & (!sk[91]) & (g56) & (!g72)) + ((!i_1_) & (!i_2_) & (g51) & (!sk[91]) & (g56) & (g72)) + ((!i_1_) & (i_2_) & (!g51) & (!sk[91]) & (!g56) & (!g72)) + ((!i_1_) & (i_2_) & (!g51) & (!sk[91]) & (!g56) & (g72)) + ((!i_1_) & (i_2_) & (!g51) & (!sk[91]) & (g56) & (!g72)) + ((!i_1_) & (i_2_) & (!g51) & (!sk[91]) & (g56) & (g72)) + ((!i_1_) & (i_2_) & (!g51) & (sk[91]) & (!g56) & (g72)) + ((!i_1_) & (i_2_) & (!g51) & (sk[91]) & (g56) & (g72)) + ((!i_1_) & (i_2_) & (g51) & (!sk[91]) & (!g56) & (!g72)) + ((!i_1_) & (i_2_) & (g51) & (!sk[91]) & (!g56) & (g72)) + ((!i_1_) & (i_2_) & (g51) & (!sk[91]) & (g56) & (!g72)) + ((!i_1_) & (i_2_) & (g51) & (!sk[91]) & (g56) & (g72)) + ((i_1_) & (!i_2_) & (!g51) & (!sk[91]) & (!g56) & (!g72)) + ((i_1_) & (!i_2_) & (!g51) & (!sk[91]) & (!g56) & (g72)) + ((i_1_) & (!i_2_) & (!g51) & (!sk[91]) & (g56) & (!g72)) + ((i_1_) & (!i_2_) & (!g51) & (!sk[91]) & (g56) & (g72)) + ((i_1_) & (!i_2_) & (!g51) & (sk[91]) & (!g56) & (g72)) + ((i_1_) & (!i_2_) & (g51) & (!sk[91]) & (!g56) & (!g72)) + ((i_1_) & (!i_2_) & (g51) & (!sk[91]) & (!g56) & (g72)) + ((i_1_) & (!i_2_) & (g51) & (!sk[91]) & (g56) & (!g72)) + ((i_1_) & (!i_2_) & (g51) & (!sk[91]) & (g56) & (g72)) + ((i_1_) & (i_2_) & (!g51) & (!sk[91]) & (!g56) & (!g72)) + ((i_1_) & (i_2_) & (!g51) & (!sk[91]) & (!g56) & (g72)) + ((i_1_) & (i_2_) & (!g51) & (!sk[91]) & (g56) & (!g72)) + ((i_1_) & (i_2_) & (!g51) & (!sk[91]) & (g56) & (g72)) + ((i_1_) & (i_2_) & (!g51) & (sk[91]) & (!g56) & (g72)) + ((i_1_) & (i_2_) & (!g51) & (sk[91]) & (g56) & (g72)) + ((i_1_) & (i_2_) & (g51) & (!sk[91]) & (!g56) & (!g72)) + ((i_1_) & (i_2_) & (g51) & (!sk[91]) & (!g56) & (g72)) + ((i_1_) & (i_2_) & (g51) & (!sk[91]) & (g56) & (!g72)) + ((i_1_) & (i_2_) & (g51) & (!sk[91]) & (g56) & (g72)));
	assign o_0_ = (((!g3) & (!sk[92]) & (g37) & (!g73)) + ((!g3) & (!sk[92]) & (g37) & (g73)) + ((!g3) & (sk[92]) & (!g37) & (g73)) + ((g3) & (!sk[92]) & (!g37) & (!g73)) + ((g3) & (!sk[92]) & (!g37) & (g73)) + ((g3) & (!sk[92]) & (g37) & (!g73)) + ((g3) & (!sk[92]) & (g37) & (g73)) + ((g3) & (sk[92]) & (!g37) & (g73)) + ((g3) & (sk[92]) & (g37) & (g73)));
	assign g75 = (((!g27) & (!sk[93]) & (g40)) + ((g27) & (!sk[93]) & (g40)) + ((g27) & (sk[93]) & (g40)));
	assign g76 = (((!g21) & (!sk[94]) & (!g23) & (!g4) & (g27) & (!g40)) + ((!g21) & (!sk[94]) & (!g23) & (!g4) & (g27) & (g40)) + ((!g21) & (!sk[94]) & (!g23) & (g4) & (!g27) & (!g40)) + ((!g21) & (!sk[94]) & (!g23) & (g4) & (!g27) & (g40)) + ((!g21) & (!sk[94]) & (!g23) & (g4) & (g27) & (!g40)) + ((!g21) & (!sk[94]) & (!g23) & (g4) & (g27) & (g40)) + ((!g21) & (!sk[94]) & (g23) & (!g4) & (!g27) & (!g40)) + ((!g21) & (!sk[94]) & (g23) & (!g4) & (!g27) & (g40)) + ((!g21) & (!sk[94]) & (g23) & (!g4) & (g27) & (!g40)) + ((!g21) & (!sk[94]) & (g23) & (!g4) & (g27) & (g40)) + ((!g21) & (!sk[94]) & (g23) & (g4) & (!g27) & (!g40)) + ((!g21) & (!sk[94]) & (g23) & (g4) & (!g27) & (g40)) + ((!g21) & (!sk[94]) & (g23) & (g4) & (g27) & (!g40)) + ((!g21) & (!sk[94]) & (g23) & (g4) & (g27) & (g40)) + ((!g21) & (sk[94]) & (!g23) & (g4) & (!g27) & (g40)) + ((!g21) & (sk[94]) & (!g23) & (g4) & (g27) & (g40)) + ((!g21) & (sk[94]) & (g23) & (!g4) & (g27) & (g40)) + ((!g21) & (sk[94]) & (g23) & (g4) & (!g27) & (g40)) + ((!g21) & (sk[94]) & (g23) & (g4) & (g27) & (g40)) + ((g21) & (!sk[94]) & (!g23) & (!g4) & (!g27) & (!g40)) + ((g21) & (!sk[94]) & (!g23) & (!g4) & (!g27) & (g40)) + ((g21) & (!sk[94]) & (!g23) & (!g4) & (g27) & (!g40)) + ((g21) & (!sk[94]) & (!g23) & (!g4) & (g27) & (g40)) + ((g21) & (!sk[94]) & (!g23) & (g4) & (!g27) & (!g40)) + ((g21) & (!sk[94]) & (!g23) & (g4) & (!g27) & (g40)) + ((g21) & (!sk[94]) & (!g23) & (g4) & (g27) & (!g40)) + ((g21) & (!sk[94]) & (!g23) & (g4) & (g27) & (g40)) + ((g21) & (!sk[94]) & (g23) & (!g4) & (!g27) & (!g40)) + ((g21) & (!sk[94]) & (g23) & (!g4) & (!g27) & (g40)) + ((g21) & (!sk[94]) & (g23) & (!g4) & (g27) & (!g40)) + ((g21) & (!sk[94]) & (g23) & (!g4) & (g27) & (g40)) + ((g21) & (!sk[94]) & (g23) & (g4) & (!g27) & (!g40)) + ((g21) & (!sk[94]) & (g23) & (g4) & (!g27) & (g40)) + ((g21) & (!sk[94]) & (g23) & (g4) & (g27) & (!g40)) + ((g21) & (!sk[94]) & (g23) & (g4) & (g27) & (g40)) + ((g21) & (sk[94]) & (!g23) & (!g4) & (g27) & (g40)) + ((g21) & (sk[94]) & (!g23) & (g4) & (!g27) & (g40)) + ((g21) & (sk[94]) & (!g23) & (g4) & (g27) & (g40)) + ((g21) & (sk[94]) & (g23) & (!g4) & (g27) & (g40)) + ((g21) & (sk[94]) & (g23) & (g4) & (!g27) & (g40)) + ((g21) & (sk[94]) & (g23) & (g4) & (g27) & (g40)));
	assign g77 = (((!i_5_) & (!i_3_) & (!i_4_) & (!sk[95]) & (g29)) + ((!i_5_) & (!i_3_) & (i_4_) & (!sk[95]) & (g29)) + ((!i_5_) & (i_3_) & (!i_4_) & (!sk[95]) & (g29)) + ((!i_5_) & (i_3_) & (i_4_) & (!sk[95]) & (g29)) + ((i_5_) & (!i_3_) & (!i_4_) & (!sk[95]) & (!g29)) + ((i_5_) & (!i_3_) & (!i_4_) & (!sk[95]) & (g29)) + ((i_5_) & (!i_3_) & (i_4_) & (!sk[95]) & (!g29)) + ((i_5_) & (!i_3_) & (i_4_) & (!sk[95]) & (g29)) + ((i_5_) & (!i_3_) & (i_4_) & (sk[95]) & (g29)) + ((i_5_) & (i_3_) & (!i_4_) & (!sk[95]) & (!g29)) + ((i_5_) & (i_3_) & (!i_4_) & (!sk[95]) & (g29)) + ((i_5_) & (i_3_) & (i_4_) & (!sk[95]) & (!g29)) + ((i_5_) & (i_3_) & (i_4_) & (!sk[95]) & (g29)));
	assign g78 = (((!sk[96]) & (!g31) & (g40)) + ((!sk[96]) & (g31) & (g40)) + ((sk[96]) & (g31) & (g40)));
	assign g79 = (((!g21) & (!sk[97]) & (!g10) & (!g23) & (g12)) + ((!g21) & (!sk[97]) & (!g10) & (g23) & (g12)) + ((!g21) & (!sk[97]) & (g10) & (!g23) & (g12)) + ((!g21) & (!sk[97]) & (g10) & (g23) & (g12)) + ((!g21) & (sk[97]) & (!g10) & (!g23) & (!g12)) + ((g21) & (!sk[97]) & (!g10) & (!g23) & (!g12)) + ((g21) & (!sk[97]) & (!g10) & (!g23) & (g12)) + ((g21) & (!sk[97]) & (!g10) & (g23) & (!g12)) + ((g21) & (!sk[97]) & (!g10) & (g23) & (g12)) + ((g21) & (!sk[97]) & (g10) & (!g23) & (!g12)) + ((g21) & (!sk[97]) & (g10) & (!g23) & (g12)) + ((g21) & (!sk[97]) & (g10) & (g23) & (!g12)) + ((g21) & (!sk[97]) & (g10) & (g23) & (g12)));
	assign g80 = (((!i_8_) & (!i_6_) & (!i_7_) & (!g19) & (!g20) & (g40)) + ((!i_8_) & (!i_6_) & (!i_7_) & (g19) & (!g20) & (g40)) + ((!i_8_) & (!i_6_) & (!i_7_) & (g19) & (g20) & (g40)) + ((!i_8_) & (!i_6_) & (i_7_) & (!g19) & (!g20) & (g40)) + ((!i_8_) & (!i_6_) & (i_7_) & (!g19) & (g20) & (g40)) + ((!i_8_) & (!i_6_) & (i_7_) & (g19) & (!g20) & (g40)) + ((!i_8_) & (!i_6_) & (i_7_) & (g19) & (g20) & (g40)) + ((i_8_) & (!i_6_) & (i_7_) & (!g19) & (!g20) & (g40)) + ((i_8_) & (!i_6_) & (i_7_) & (!g19) & (g20) & (g40)) + ((i_8_) & (!i_6_) & (i_7_) & (g19) & (!g20) & (g40)) + ((i_8_) & (!i_6_) & (i_7_) & (g19) & (g20) & (g40)));
	assign g81 = (((!sk[99]) & (!g8) & (!g14) & (!g16) & (g78) & (!g80)) + ((!sk[99]) & (!g8) & (!g14) & (!g16) & (g78) & (g80)) + ((!sk[99]) & (!g8) & (!g14) & (g16) & (!g78) & (!g80)) + ((!sk[99]) & (!g8) & (!g14) & (g16) & (!g78) & (g80)) + ((!sk[99]) & (!g8) & (!g14) & (g16) & (g78) & (!g80)) + ((!sk[99]) & (!g8) & (!g14) & (g16) & (g78) & (g80)) + ((!sk[99]) & (!g8) & (g14) & (!g16) & (!g78) & (!g80)) + ((!sk[99]) & (!g8) & (g14) & (!g16) & (!g78) & (g80)) + ((!sk[99]) & (!g8) & (g14) & (!g16) & (g78) & (!g80)) + ((!sk[99]) & (!g8) & (g14) & (!g16) & (g78) & (g80)) + ((!sk[99]) & (!g8) & (g14) & (g16) & (!g78) & (!g80)) + ((!sk[99]) & (!g8) & (g14) & (g16) & (!g78) & (g80)) + ((!sk[99]) & (!g8) & (g14) & (g16) & (g78) & (!g80)) + ((!sk[99]) & (!g8) & (g14) & (g16) & (g78) & (g80)) + ((!sk[99]) & (g8) & (!g14) & (!g16) & (!g78) & (!g80)) + ((!sk[99]) & (g8) & (!g14) & (!g16) & (!g78) & (g80)) + ((!sk[99]) & (g8) & (!g14) & (!g16) & (g78) & (!g80)) + ((!sk[99]) & (g8) & (!g14) & (!g16) & (g78) & (g80)) + ((!sk[99]) & (g8) & (!g14) & (g16) & (!g78) & (!g80)) + ((!sk[99]) & (g8) & (!g14) & (g16) & (!g78) & (g80)) + ((!sk[99]) & (g8) & (!g14) & (g16) & (g78) & (!g80)) + ((!sk[99]) & (g8) & (!g14) & (g16) & (g78) & (g80)) + ((!sk[99]) & (g8) & (g14) & (!g16) & (!g78) & (!g80)) + ((!sk[99]) & (g8) & (g14) & (!g16) & (!g78) & (g80)) + ((!sk[99]) & (g8) & (g14) & (!g16) & (g78) & (!g80)) + ((!sk[99]) & (g8) & (g14) & (!g16) & (g78) & (g80)) + ((!sk[99]) & (g8) & (g14) & (g16) & (!g78) & (!g80)) + ((!sk[99]) & (g8) & (g14) & (g16) & (!g78) & (g80)) + ((!sk[99]) & (g8) & (g14) & (g16) & (g78) & (!g80)) + ((!sk[99]) & (g8) & (g14) & (g16) & (g78) & (g80)) + ((sk[99]) & (!g8) & (!g14) & (!g16) & (!g78) & (!g80)) + ((sk[99]) & (!g8) & (!g14) & (g16) & (!g78) & (!g80)) + ((sk[99]) & (!g8) & (g14) & (!g16) & (!g78) & (!g80)) + ((sk[99]) & (!g8) & (g14) & (g16) & (!g78) & (!g80)) + ((sk[99]) & (g8) & (!g14) & (!g16) & (!g78) & (!g80)) + ((sk[99]) & (g8) & (!g14) & (g16) & (!g78) & (!g80)) + ((sk[99]) & (g8) & (!g14) & (g16) & (g78) & (!g80)) + ((sk[99]) & (g8) & (g14) & (!g16) & (!g78) & (!g80)) + ((sk[99]) & (g8) & (g14) & (g16) & (!g78) & (!g80)));
	assign g82 = (((!g29) & (!g39) & (!g78) & (!g79) & (sk[100]) & (g81)) + ((!g29) & (!g39) & (!g78) & (g79) & (!sk[100]) & (!g81)) + ((!g29) & (!g39) & (!g78) & (g79) & (!sk[100]) & (g81)) + ((!g29) & (!g39) & (!g78) & (g79) & (sk[100]) & (g81)) + ((!g29) & (!g39) & (g78) & (!g79) & (!sk[100]) & (!g81)) + ((!g29) & (!g39) & (g78) & (!g79) & (!sk[100]) & (g81)) + ((!g29) & (!g39) & (g78) & (g79) & (!sk[100]) & (!g81)) + ((!g29) & (!g39) & (g78) & (g79) & (!sk[100]) & (g81)) + ((!g29) & (!g39) & (g78) & (g79) & (sk[100]) & (g81)) + ((!g29) & (g39) & (!g78) & (!g79) & (!sk[100]) & (!g81)) + ((!g29) & (g39) & (!g78) & (!g79) & (!sk[100]) & (g81)) + ((!g29) & (g39) & (!g78) & (!g79) & (sk[100]) & (g81)) + ((!g29) & (g39) & (!g78) & (g79) & (!sk[100]) & (!g81)) + ((!g29) & (g39) & (!g78) & (g79) & (!sk[100]) & (g81)) + ((!g29) & (g39) & (!g78) & (g79) & (sk[100]) & (g81)) + ((!g29) & (g39) & (g78) & (!g79) & (!sk[100]) & (!g81)) + ((!g29) & (g39) & (g78) & (!g79) & (!sk[100]) & (g81)) + ((!g29) & (g39) & (g78) & (g79) & (!sk[100]) & (!g81)) + ((!g29) & (g39) & (g78) & (g79) & (!sk[100]) & (g81)) + ((!g29) & (g39) & (g78) & (g79) & (sk[100]) & (g81)) + ((g29) & (!g39) & (!g78) & (!g79) & (!sk[100]) & (!g81)) + ((g29) & (!g39) & (!g78) & (!g79) & (!sk[100]) & (g81)) + ((g29) & (!g39) & (!g78) & (!g79) & (sk[100]) & (g81)) + ((g29) & (!g39) & (!g78) & (g79) & (!sk[100]) & (!g81)) + ((g29) & (!g39) & (!g78) & (g79) & (!sk[100]) & (g81)) + ((g29) & (!g39) & (!g78) & (g79) & (sk[100]) & (g81)) + ((g29) & (!g39) & (g78) & (!g79) & (!sk[100]) & (!g81)) + ((g29) & (!g39) & (g78) & (!g79) & (!sk[100]) & (g81)) + ((g29) & (!g39) & (g78) & (g79) & (!sk[100]) & (!g81)) + ((g29) & (!g39) & (g78) & (g79) & (!sk[100]) & (g81)) + ((g29) & (!g39) & (g78) & (g79) & (sk[100]) & (g81)) + ((g29) & (g39) & (!g78) & (!g79) & (!sk[100]) & (!g81)) + ((g29) & (g39) & (!g78) & (!g79) & (!sk[100]) & (g81)) + ((g29) & (g39) & (!g78) & (g79) & (!sk[100]) & (!g81)) + ((g29) & (g39) & (!g78) & (g79) & (!sk[100]) & (g81)) + ((g29) & (g39) & (g78) & (!g79) & (!sk[100]) & (!g81)) + ((g29) & (g39) & (g78) & (!g79) & (!sk[100]) & (g81)) + ((g29) & (g39) & (g78) & (g79) & (!sk[100]) & (!g81)) + ((g29) & (g39) & (g78) & (g79) & (!sk[100]) & (g81)));
	assign g83 = (((!g17) & (!g75) & (!sk[101]) & (!g76) & (g1544) & (!g82)) + ((!g17) & (!g75) & (!sk[101]) & (!g76) & (g1544) & (g82)) + ((!g17) & (!g75) & (!sk[101]) & (g76) & (!g1544) & (!g82)) + ((!g17) & (!g75) & (!sk[101]) & (g76) & (!g1544) & (g82)) + ((!g17) & (!g75) & (!sk[101]) & (g76) & (g1544) & (!g82)) + ((!g17) & (!g75) & (!sk[101]) & (g76) & (g1544) & (g82)) + ((!g17) & (!g75) & (sk[101]) & (!g76) & (g1544) & (g82)) + ((!g17) & (g75) & (!sk[101]) & (!g76) & (!g1544) & (!g82)) + ((!g17) & (g75) & (!sk[101]) & (!g76) & (!g1544) & (g82)) + ((!g17) & (g75) & (!sk[101]) & (!g76) & (g1544) & (!g82)) + ((!g17) & (g75) & (!sk[101]) & (!g76) & (g1544) & (g82)) + ((!g17) & (g75) & (!sk[101]) & (g76) & (!g1544) & (!g82)) + ((!g17) & (g75) & (!sk[101]) & (g76) & (!g1544) & (g82)) + ((!g17) & (g75) & (!sk[101]) & (g76) & (g1544) & (!g82)) + ((!g17) & (g75) & (!sk[101]) & (g76) & (g1544) & (g82)) + ((g17) & (!g75) & (!sk[101]) & (!g76) & (!g1544) & (!g82)) + ((g17) & (!g75) & (!sk[101]) & (!g76) & (!g1544) & (g82)) + ((g17) & (!g75) & (!sk[101]) & (!g76) & (g1544) & (!g82)) + ((g17) & (!g75) & (!sk[101]) & (!g76) & (g1544) & (g82)) + ((g17) & (!g75) & (!sk[101]) & (g76) & (!g1544) & (!g82)) + ((g17) & (!g75) & (!sk[101]) & (g76) & (!g1544) & (g82)) + ((g17) & (!g75) & (!sk[101]) & (g76) & (g1544) & (!g82)) + ((g17) & (!g75) & (!sk[101]) & (g76) & (g1544) & (g82)) + ((g17) & (!g75) & (sk[101]) & (!g76) & (g1544) & (g82)) + ((g17) & (g75) & (!sk[101]) & (!g76) & (!g1544) & (!g82)) + ((g17) & (g75) & (!sk[101]) & (!g76) & (!g1544) & (g82)) + ((g17) & (g75) & (!sk[101]) & (!g76) & (g1544) & (!g82)) + ((g17) & (g75) & (!sk[101]) & (!g76) & (g1544) & (g82)) + ((g17) & (g75) & (!sk[101]) & (g76) & (!g1544) & (!g82)) + ((g17) & (g75) & (!sk[101]) & (g76) & (!g1544) & (g82)) + ((g17) & (g75) & (!sk[101]) & (g76) & (g1544) & (!g82)) + ((g17) & (g75) & (!sk[101]) & (g76) & (g1544) & (g82)) + ((g17) & (g75) & (sk[101]) & (!g76) & (g1544) & (g82)));
	assign o_1_ = (((!i_8_) & (!i_7_) & (!g5) & (!g40) & (g73) & (!g83)) + ((!i_8_) & (!i_7_) & (!g5) & (g40) & (g73) & (!g83)) + ((!i_8_) & (!i_7_) & (g5) & (!g40) & (g73) & (!g83)) + ((!i_8_) & (!i_7_) & (g5) & (g40) & (g73) & (!g83)) + ((!i_8_) & (!i_7_) & (g5) & (g40) & (g73) & (g83)) + ((!i_8_) & (i_7_) & (!g5) & (!g40) & (g73) & (!g83)) + ((!i_8_) & (i_7_) & (!g5) & (g40) & (g73) & (!g83)) + ((!i_8_) & (i_7_) & (g5) & (!g40) & (g73) & (!g83)) + ((!i_8_) & (i_7_) & (g5) & (g40) & (g73) & (!g83)) + ((i_8_) & (!i_7_) & (!g5) & (!g40) & (g73) & (!g83)) + ((i_8_) & (!i_7_) & (!g5) & (g40) & (g73) & (!g83)) + ((i_8_) & (!i_7_) & (!g5) & (g40) & (g73) & (g83)) + ((i_8_) & (!i_7_) & (g5) & (!g40) & (g73) & (!g83)) + ((i_8_) & (!i_7_) & (g5) & (g40) & (g73) & (!g83)) + ((i_8_) & (!i_7_) & (g5) & (g40) & (g73) & (g83)) + ((i_8_) & (i_7_) & (!g5) & (!g40) & (g73) & (!g83)) + ((i_8_) & (i_7_) & (!g5) & (g40) & (g73) & (!g83)) + ((i_8_) & (i_7_) & (g5) & (!g40) & (g73) & (!g83)) + ((i_8_) & (i_7_) & (g5) & (g40) & (g73) & (!g83)));
	assign g85 = (((!g2) & (!i_8_) & (!sk[103]) & (!i_6_) & (i_7_)) + ((!g2) & (!i_8_) & (!sk[103]) & (i_6_) & (i_7_)) + ((!g2) & (i_8_) & (!sk[103]) & (!i_6_) & (i_7_)) + ((!g2) & (i_8_) & (!sk[103]) & (i_6_) & (i_7_)) + ((g2) & (!i_8_) & (!sk[103]) & (!i_6_) & (!i_7_)) + ((g2) & (!i_8_) & (!sk[103]) & (!i_6_) & (i_7_)) + ((g2) & (!i_8_) & (!sk[103]) & (i_6_) & (!i_7_)) + ((g2) & (!i_8_) & (!sk[103]) & (i_6_) & (i_7_)) + ((g2) & (i_8_) & (!sk[103]) & (!i_6_) & (!i_7_)) + ((g2) & (i_8_) & (!sk[103]) & (!i_6_) & (i_7_)) + ((g2) & (i_8_) & (!sk[103]) & (i_6_) & (!i_7_)) + ((g2) & (i_8_) & (!sk[103]) & (i_6_) & (i_7_)) + ((g2) & (i_8_) & (sk[103]) & (i_6_) & (!i_7_)));
	assign o_2_ = (((!g28) & (!g52) & (!g29) & (!sk[104]) & (g73) & (!g85)) + ((!g28) & (!g52) & (!g29) & (!sk[104]) & (g73) & (g85)) + ((!g28) & (!g52) & (!g29) & (sk[104]) & (g73) & (g85)) + ((!g28) & (!g52) & (g29) & (!sk[104]) & (!g73) & (!g85)) + ((!g28) & (!g52) & (g29) & (!sk[104]) & (!g73) & (g85)) + ((!g28) & (!g52) & (g29) & (!sk[104]) & (g73) & (!g85)) + ((!g28) & (!g52) & (g29) & (!sk[104]) & (g73) & (g85)) + ((!g28) & (!g52) & (g29) & (sk[104]) & (g73) & (g85)) + ((!g28) & (g52) & (!g29) & (!sk[104]) & (!g73) & (!g85)) + ((!g28) & (g52) & (!g29) & (!sk[104]) & (!g73) & (g85)) + ((!g28) & (g52) & (!g29) & (!sk[104]) & (g73) & (!g85)) + ((!g28) & (g52) & (!g29) & (!sk[104]) & (g73) & (g85)) + ((!g28) & (g52) & (!g29) & (sk[104]) & (g73) & (g85)) + ((!g28) & (g52) & (g29) & (!sk[104]) & (!g73) & (!g85)) + ((!g28) & (g52) & (g29) & (!sk[104]) & (!g73) & (g85)) + ((!g28) & (g52) & (g29) & (!sk[104]) & (g73) & (!g85)) + ((!g28) & (g52) & (g29) & (!sk[104]) & (g73) & (g85)) + ((!g28) & (g52) & (g29) & (sk[104]) & (g73) & (!g85)) + ((!g28) & (g52) & (g29) & (sk[104]) & (g73) & (g85)) + ((g28) & (!g52) & (!g29) & (!sk[104]) & (!g73) & (!g85)) + ((g28) & (!g52) & (!g29) & (!sk[104]) & (!g73) & (g85)) + ((g28) & (!g52) & (!g29) & (!sk[104]) & (g73) & (!g85)) + ((g28) & (!g52) & (!g29) & (!sk[104]) & (g73) & (g85)) + ((g28) & (!g52) & (!g29) & (sk[104]) & (g73) & (!g85)) + ((g28) & (!g52) & (!g29) & (sk[104]) & (g73) & (g85)) + ((g28) & (!g52) & (g29) & (!sk[104]) & (!g73) & (!g85)) + ((g28) & (!g52) & (g29) & (!sk[104]) & (!g73) & (g85)) + ((g28) & (!g52) & (g29) & (!sk[104]) & (g73) & (!g85)) + ((g28) & (!g52) & (g29) & (!sk[104]) & (g73) & (g85)) + ((g28) & (!g52) & (g29) & (sk[104]) & (g73) & (!g85)) + ((g28) & (!g52) & (g29) & (sk[104]) & (g73) & (g85)) + ((g28) & (g52) & (!g29) & (!sk[104]) & (!g73) & (!g85)) + ((g28) & (g52) & (!g29) & (!sk[104]) & (!g73) & (g85)) + ((g28) & (g52) & (!g29) & (!sk[104]) & (g73) & (!g85)) + ((g28) & (g52) & (!g29) & (!sk[104]) & (g73) & (g85)) + ((g28) & (g52) & (!g29) & (sk[104]) & (g73) & (!g85)) + ((g28) & (g52) & (!g29) & (sk[104]) & (g73) & (g85)) + ((g28) & (g52) & (g29) & (!sk[104]) & (!g73) & (!g85)) + ((g28) & (g52) & (g29) & (!sk[104]) & (!g73) & (g85)) + ((g28) & (g52) & (g29) & (!sk[104]) & (g73) & (!g85)) + ((g28) & (g52) & (g29) & (!sk[104]) & (g73) & (g85)) + ((g28) & (g52) & (g29) & (sk[104]) & (g73) & (!g85)) + ((g28) & (g52) & (g29) & (sk[104]) & (g73) & (g85)));
	assign g87 = (((!g57) & (!sk[105]) & (g39)) + ((g57) & (!sk[105]) & (g39)) + ((g57) & (sk[105]) & (g39)));
	assign g88 = (((!sk[106]) & (!g34) & (g87)) + ((!sk[106]) & (g34) & (g87)) + ((sk[106]) & (g34) & (g87)));
	assign g89 = (((!sk[107]) & (!i_8_) & (g88)) + ((!sk[107]) & (i_8_) & (g88)) + ((sk[107]) & (!i_8_) & (!g88)) + ((sk[107]) & (i_8_) & (!g88)) + ((sk[107]) & (i_8_) & (g88)));
	assign g90 = (((!g6) & (!sk[108]) & (i_15_) & (!g48)) + ((!g6) & (!sk[108]) & (i_15_) & (g48)) + ((!g6) & (sk[108]) & (!i_15_) & (!g48)) + ((!g6) & (sk[108]) & (!i_15_) & (g48)) + ((!g6) & (sk[108]) & (i_15_) & (!g48)) + ((!g6) & (sk[108]) & (i_15_) & (g48)) + ((g6) & (!sk[108]) & (!i_15_) & (!g48)) + ((g6) & (!sk[108]) & (!i_15_) & (g48)) + ((g6) & (!sk[108]) & (i_15_) & (!g48)) + ((g6) & (!sk[108]) & (i_15_) & (g48)) + ((g6) & (sk[108]) & (!i_15_) & (g48)) + ((g6) & (sk[108]) & (i_15_) & (!g48)) + ((g6) & (sk[108]) & (i_15_) & (g48)));
	assign g91 = (((!i_14_) & (!i_12_) & (sk[109]) & (!i_13_)) + ((!i_14_) & (!i_12_) & (sk[109]) & (i_13_)) + ((!i_14_) & (i_12_) & (!sk[109]) & (!i_13_)) + ((!i_14_) & (i_12_) & (!sk[109]) & (i_13_)) + ((!i_14_) & (i_12_) & (sk[109]) & (i_13_)) + ((i_14_) & (!i_12_) & (!sk[109]) & (!i_13_)) + ((i_14_) & (!i_12_) & (!sk[109]) & (i_13_)) + ((i_14_) & (!i_12_) & (sk[109]) & (!i_13_)) + ((i_14_) & (!i_12_) & (sk[109]) & (i_13_)) + ((i_14_) & (i_12_) & (!sk[109]) & (!i_13_)) + ((i_14_) & (i_12_) & (!sk[109]) & (i_13_)) + ((i_14_) & (i_12_) & (sk[109]) & (!i_13_)) + ((i_14_) & (i_12_) & (sk[109]) & (i_13_)));
	assign g92 = (((!g6) & (!i_15_) & (sk[110]) & (!g91)) + ((!g6) & (!i_15_) & (sk[110]) & (g91)) + ((!g6) & (i_15_) & (!sk[110]) & (!g91)) + ((!g6) & (i_15_) & (!sk[110]) & (g91)) + ((!g6) & (i_15_) & (sk[110]) & (!g91)) + ((!g6) & (i_15_) & (sk[110]) & (g91)) + ((g6) & (!i_15_) & (!sk[110]) & (!g91)) + ((g6) & (!i_15_) & (!sk[110]) & (g91)) + ((g6) & (!i_15_) & (sk[110]) & (!g91)) + ((g6) & (!i_15_) & (sk[110]) & (g91)) + ((g6) & (i_15_) & (!sk[110]) & (!g91)) + ((g6) & (i_15_) & (!sk[110]) & (g91)) + ((g6) & (i_15_) & (sk[110]) & (g91)));
	assign g93 = (((!i_11_) & (!sk[111]) & (!i_9_) & (!i_10_) & (i_15_)) + ((!i_11_) & (!sk[111]) & (!i_9_) & (i_10_) & (i_15_)) + ((!i_11_) & (!sk[111]) & (i_9_) & (!i_10_) & (i_15_)) + ((!i_11_) & (!sk[111]) & (i_9_) & (i_10_) & (i_15_)) + ((!i_11_) & (sk[111]) & (!i_9_) & (!i_10_) & (!i_15_)) + ((!i_11_) & (sk[111]) & (!i_9_) & (!i_10_) & (i_15_)) + ((!i_11_) & (sk[111]) & (!i_9_) & (i_10_) & (!i_15_)) + ((!i_11_) & (sk[111]) & (!i_9_) & (i_10_) & (i_15_)) + ((!i_11_) & (sk[111]) & (i_9_) & (!i_10_) & (!i_15_)) + ((!i_11_) & (sk[111]) & (i_9_) & (!i_10_) & (i_15_)) + ((!i_11_) & (sk[111]) & (i_9_) & (i_10_) & (!i_15_)) + ((!i_11_) & (sk[111]) & (i_9_) & (i_10_) & (i_15_)) + ((i_11_) & (!sk[111]) & (!i_9_) & (!i_10_) & (!i_15_)) + ((i_11_) & (!sk[111]) & (!i_9_) & (!i_10_) & (i_15_)) + ((i_11_) & (!sk[111]) & (!i_9_) & (i_10_) & (!i_15_)) + ((i_11_) & (!sk[111]) & (!i_9_) & (i_10_) & (i_15_)) + ((i_11_) & (!sk[111]) & (i_9_) & (!i_10_) & (!i_15_)) + ((i_11_) & (!sk[111]) & (i_9_) & (!i_10_) & (i_15_)) + ((i_11_) & (!sk[111]) & (i_9_) & (i_10_) & (!i_15_)) + ((i_11_) & (!sk[111]) & (i_9_) & (i_10_) & (i_15_)) + ((i_11_) & (sk[111]) & (!i_9_) & (!i_10_) & (!i_15_)) + ((i_11_) & (sk[111]) & (!i_9_) & (i_10_) & (!i_15_)) + ((i_11_) & (sk[111]) & (!i_9_) & (i_10_) & (i_15_)) + ((i_11_) & (sk[111]) & (i_9_) & (!i_10_) & (!i_15_)) + ((i_11_) & (sk[111]) & (i_9_) & (!i_10_) & (i_15_)) + ((i_11_) & (sk[111]) & (i_9_) & (i_10_) & (!i_15_)) + ((i_11_) & (sk[111]) & (i_9_) & (i_10_) & (i_15_)));
	assign g94 = (((!g91) & (!sk[112]) & (g93)) + ((!g91) & (sk[112]) & (!g93)) + ((g91) & (!sk[112]) & (g93)));
	assign g95 = (((!i_11_) & (!sk[113]) & (!i_9_) & (!i_10_) & (i_15_)) + ((!i_11_) & (!sk[113]) & (!i_9_) & (i_10_) & (i_15_)) + ((!i_11_) & (!sk[113]) & (i_9_) & (!i_10_) & (i_15_)) + ((!i_11_) & (!sk[113]) & (i_9_) & (i_10_) & (i_15_)) + ((i_11_) & (!sk[113]) & (!i_9_) & (!i_10_) & (!i_15_)) + ((i_11_) & (!sk[113]) & (!i_9_) & (!i_10_) & (i_15_)) + ((i_11_) & (!sk[113]) & (!i_9_) & (i_10_) & (!i_15_)) + ((i_11_) & (!sk[113]) & (!i_9_) & (i_10_) & (i_15_)) + ((i_11_) & (!sk[113]) & (i_9_) & (!i_10_) & (!i_15_)) + ((i_11_) & (!sk[113]) & (i_9_) & (!i_10_) & (i_15_)) + ((i_11_) & (!sk[113]) & (i_9_) & (i_10_) & (!i_15_)) + ((i_11_) & (!sk[113]) & (i_9_) & (i_10_) & (i_15_)) + ((i_11_) & (sk[113]) & (!i_9_) & (!i_10_) & (!i_15_)));
	assign g96 = (((!sk[114]) & (!g48) & (g95)) + ((!sk[114]) & (g48) & (g95)) + ((sk[114]) & (!g48) & (!g95)) + ((sk[114]) & (g48) & (!g95)) + ((sk[114]) & (g48) & (g95)));
	assign g97 = (((!g89) & (!g94) & (sk[115]) & (!g96)) + ((!g89) & (g94) & (!sk[115]) & (!g96)) + ((!g89) & (g94) & (!sk[115]) & (g96)) + ((!g89) & (g94) & (sk[115]) & (!g96)) + ((!g89) & (g94) & (sk[115]) & (g96)) + ((g89) & (!g94) & (!sk[115]) & (!g96)) + ((g89) & (!g94) & (!sk[115]) & (g96)) + ((g89) & (g94) & (!sk[115]) & (!g96)) + ((g89) & (g94) & (!sk[115]) & (g96)));
	assign g98 = (((!i_5_) & (!i_3_) & (!i_4_) & (!sk[116]) & (g57)) + ((!i_5_) & (!i_3_) & (i_4_) & (!sk[116]) & (g57)) + ((!i_5_) & (i_3_) & (!i_4_) & (!sk[116]) & (g57)) + ((!i_5_) & (i_3_) & (i_4_) & (!sk[116]) & (g57)) + ((i_5_) & (!i_3_) & (!i_4_) & (!sk[116]) & (!g57)) + ((i_5_) & (!i_3_) & (!i_4_) & (!sk[116]) & (g57)) + ((i_5_) & (!i_3_) & (i_4_) & (!sk[116]) & (!g57)) + ((i_5_) & (!i_3_) & (i_4_) & (!sk[116]) & (g57)) + ((i_5_) & (!i_3_) & (i_4_) & (sk[116]) & (g57)) + ((i_5_) & (i_3_) & (!i_4_) & (!sk[116]) & (!g57)) + ((i_5_) & (i_3_) & (!i_4_) & (!sk[116]) & (g57)) + ((i_5_) & (i_3_) & (i_4_) & (!sk[116]) & (!g57)) + ((i_5_) & (i_3_) & (i_4_) & (!sk[116]) & (g57)));
	assign g99 = (((!g38) & (!sk[117]) & (g98)) + ((g38) & (!sk[117]) & (g98)) + ((g38) & (sk[117]) & (g98)));
	assign g100 = (((!g4) & (!sk[118]) & (g98)) + ((g4) & (!sk[118]) & (g98)) + ((g4) & (sk[118]) & (g98)));
	assign g101 = (((!sk[119]) & (!i_8_) & (g100)) + ((!sk[119]) & (i_8_) & (g100)) + ((sk[119]) & (i_8_) & (g100)));
	assign g102 = (((!i_11_) & (!i_9_) & (!i_10_) & (!sk[120]) & (i_15_)) + ((!i_11_) & (!i_9_) & (!i_10_) & (sk[120]) & (!i_15_)) + ((!i_11_) & (!i_9_) & (!i_10_) & (sk[120]) & (i_15_)) + ((!i_11_) & (!i_9_) & (i_10_) & (!sk[120]) & (i_15_)) + ((!i_11_) & (!i_9_) & (i_10_) & (sk[120]) & (!i_15_)) + ((!i_11_) & (!i_9_) & (i_10_) & (sk[120]) & (i_15_)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[120]) & (i_15_)) + ((!i_11_) & (i_9_) & (!i_10_) & (sk[120]) & (!i_15_)) + ((!i_11_) & (i_9_) & (!i_10_) & (sk[120]) & (i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[120]) & (i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (sk[120]) & (!i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (sk[120]) & (i_15_)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[120]) & (!i_15_)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[120]) & (i_15_)) + ((i_11_) & (!i_9_) & (!i_10_) & (sk[120]) & (!i_15_)) + ((i_11_) & (!i_9_) & (!i_10_) & (sk[120]) & (i_15_)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[120]) & (!i_15_)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[120]) & (i_15_)) + ((i_11_) & (!i_9_) & (i_10_) & (sk[120]) & (i_15_)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[120]) & (!i_15_)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[120]) & (i_15_)) + ((i_11_) & (i_9_) & (!i_10_) & (sk[120]) & (!i_15_)) + ((i_11_) & (i_9_) & (!i_10_) & (sk[120]) & (i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[120]) & (!i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[120]) & (i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (sk[120]) & (!i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (sk[120]) & (i_15_)));
	assign g103 = (((!g48) & (sk[121]) & (g102)) + ((g48) & (!sk[121]) & (!g102)) + ((g48) & (!sk[121]) & (g102)) + ((g48) & (sk[121]) & (!g102)) + ((g48) & (sk[121]) & (g102)));
	assign g104 = (((!i_11_) & (!i_9_) & (i_10_) & (!sk[122]) & (i_15_)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[122]) & (!i_15_)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[122]) & (i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[122]) & (!i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[122]) & (i_15_)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[122]) & (!i_15_)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[122]) & (i_15_)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[122]) & (!i_15_)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[122]) & (i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[122]) & (!i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[122]) & (i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (sk[122]) & (!i_15_)));
	assign g105 = (((!sk[123]) & (g48) & (!g104)) + ((!sk[123]) & (g48) & (g104)) + ((sk[123]) & (!g48) & (g104)));
	assign g106 = (((!sk[124]) & (!g99) & (!g101) & (!g103) & (!g90) & (g105)) + ((!sk[124]) & (!g99) & (!g101) & (!g103) & (g90) & (g105)) + ((!sk[124]) & (!g99) & (!g101) & (g103) & (!g90) & (g105)) + ((!sk[124]) & (!g99) & (!g101) & (g103) & (g90) & (g105)) + ((!sk[124]) & (!g99) & (g101) & (!g103) & (!g90) & (g105)) + ((!sk[124]) & (!g99) & (g101) & (!g103) & (g90) & (g105)) + ((!sk[124]) & (!g99) & (g101) & (g103) & (!g90) & (g105)) + ((!sk[124]) & (!g99) & (g101) & (g103) & (g90) & (g105)) + ((!sk[124]) & (g99) & (!g101) & (!g103) & (!g90) & (!g105)) + ((!sk[124]) & (g99) & (!g101) & (!g103) & (!g90) & (g105)) + ((!sk[124]) & (g99) & (!g101) & (!g103) & (g90) & (!g105)) + ((!sk[124]) & (g99) & (!g101) & (!g103) & (g90) & (g105)) + ((!sk[124]) & (g99) & (!g101) & (g103) & (!g90) & (!g105)) + ((!sk[124]) & (g99) & (!g101) & (g103) & (!g90) & (g105)) + ((!sk[124]) & (g99) & (!g101) & (g103) & (g90) & (!g105)) + ((!sk[124]) & (g99) & (!g101) & (g103) & (g90) & (g105)) + ((!sk[124]) & (g99) & (g101) & (!g103) & (!g90) & (!g105)) + ((!sk[124]) & (g99) & (g101) & (!g103) & (!g90) & (g105)) + ((!sk[124]) & (g99) & (g101) & (!g103) & (g90) & (!g105)) + ((!sk[124]) & (g99) & (g101) & (!g103) & (g90) & (g105)) + ((!sk[124]) & (g99) & (g101) & (g103) & (!g90) & (!g105)) + ((!sk[124]) & (g99) & (g101) & (g103) & (!g90) & (g105)) + ((!sk[124]) & (g99) & (g101) & (g103) & (g90) & (!g105)) + ((!sk[124]) & (g99) & (g101) & (g103) & (g90) & (g105)) + ((sk[124]) & (!g99) & (!g101) & (!g103) & (!g90) & (!g105)) + ((sk[124]) & (!g99) & (!g101) & (!g103) & (!g90) & (g105)) + ((sk[124]) & (!g99) & (!g101) & (!g103) & (g90) & (!g105)) + ((sk[124]) & (!g99) & (!g101) & (!g103) & (g90) & (g105)) + ((sk[124]) & (!g99) & (!g101) & (g103) & (!g90) & (!g105)) + ((sk[124]) & (!g99) & (!g101) & (g103) & (!g90) & (g105)) + ((sk[124]) & (!g99) & (!g101) & (g103) & (g90) & (!g105)) + ((sk[124]) & (!g99) & (!g101) & (g103) & (g90) & (g105)) + ((sk[124]) & (!g99) & (g101) & (!g103) & (g90) & (!g105)) + ((sk[124]) & (!g99) & (g101) & (g103) & (g90) & (!g105)) + ((sk[124]) & (g99) & (!g101) & (g103) & (!g90) & (!g105)) + ((sk[124]) & (g99) & (!g101) & (g103) & (g90) & (!g105)) + ((sk[124]) & (g99) & (g101) & (g103) & (g90) & (!g105)));
	assign g107 = (((!g89) & (!sk[125]) & (!g90) & (!g92) & (!g97) & (g106)) + ((!g89) & (!sk[125]) & (!g90) & (!g92) & (g97) & (g106)) + ((!g89) & (!sk[125]) & (!g90) & (g92) & (!g97) & (g106)) + ((!g89) & (!sk[125]) & (!g90) & (g92) & (g97) & (g106)) + ((!g89) & (!sk[125]) & (g90) & (!g92) & (!g97) & (g106)) + ((!g89) & (!sk[125]) & (g90) & (!g92) & (g97) & (g106)) + ((!g89) & (!sk[125]) & (g90) & (g92) & (!g97) & (g106)) + ((!g89) & (!sk[125]) & (g90) & (g92) & (g97) & (g106)) + ((!g89) & (sk[125]) & (g90) & (g92) & (!g97) & (g106)) + ((g89) & (!sk[125]) & (!g90) & (!g92) & (!g97) & (!g106)) + ((g89) & (!sk[125]) & (!g90) & (!g92) & (!g97) & (g106)) + ((g89) & (!sk[125]) & (!g90) & (!g92) & (g97) & (!g106)) + ((g89) & (!sk[125]) & (!g90) & (!g92) & (g97) & (g106)) + ((g89) & (!sk[125]) & (!g90) & (g92) & (!g97) & (!g106)) + ((g89) & (!sk[125]) & (!g90) & (g92) & (!g97) & (g106)) + ((g89) & (!sk[125]) & (!g90) & (g92) & (g97) & (!g106)) + ((g89) & (!sk[125]) & (!g90) & (g92) & (g97) & (g106)) + ((g89) & (!sk[125]) & (g90) & (!g92) & (!g97) & (!g106)) + ((g89) & (!sk[125]) & (g90) & (!g92) & (!g97) & (g106)) + ((g89) & (!sk[125]) & (g90) & (!g92) & (g97) & (!g106)) + ((g89) & (!sk[125]) & (g90) & (!g92) & (g97) & (g106)) + ((g89) & (!sk[125]) & (g90) & (g92) & (!g97) & (!g106)) + ((g89) & (!sk[125]) & (g90) & (g92) & (!g97) & (g106)) + ((g89) & (!sk[125]) & (g90) & (g92) & (g97) & (!g106)) + ((g89) & (!sk[125]) & (g90) & (g92) & (g97) & (g106)) + ((g89) & (sk[125]) & (!g90) & (!g92) & (!g97) & (g106)) + ((g89) & (sk[125]) & (!g90) & (g92) & (!g97) & (g106)) + ((g89) & (sk[125]) & (g90) & (!g92) & (!g97) & (g106)) + ((g89) & (sk[125]) & (g90) & (g92) & (!g97) & (g106)));
	assign g108 = (((g34) & (!sk[126]) & (!g98)) + ((g34) & (!sk[126]) & (g98)) + ((g34) & (sk[126]) & (g98)));
	assign g109 = (((!sk[127]) & (i_8_) & (!g108)) + ((!sk[127]) & (i_8_) & (g108)) + ((sk[127]) & (!i_8_) & (g108)));
	assign g110 = (((!sk[0]) & (g52) & (!g57)) + ((!sk[0]) & (g52) & (g57)) + ((sk[0]) & (g52) & (g57)));
	assign g111 = (((!sk[1]) & (i_8_) & (!g30)) + ((!sk[1]) & (i_8_) & (g30)) + ((sk[1]) & (i_8_) & (g30)));
	assign g112 = (((!sk[2]) & (g110) & (!g111)) + ((!sk[2]) & (g110) & (g111)) + ((sk[2]) & (g110) & (g111)));
	assign g113 = (((!sk[3]) & (i_9_) & (!i_10_)) + ((!sk[3]) & (i_9_) & (i_10_)) + ((sk[3]) & (i_9_) & (i_10_)));
	assign g114 = (((!sk[4]) & (g53) & (!g113) & (!g48)) + ((!sk[4]) & (g53) & (!g113) & (g48)) + ((!sk[4]) & (g53) & (g113) & (!g48)) + ((!sk[4]) & (g53) & (g113) & (g48)) + ((sk[4]) & (g53) & (g113) & (!g48)));
	assign g115 = (((!i_11_) & (!i_9_) & (!sk[5]) & (i_10_) & (i_15_)) + ((!i_11_) & (!i_9_) & (sk[5]) & (!i_10_) & (!i_15_)) + ((!i_11_) & (!i_9_) & (sk[5]) & (!i_10_) & (i_15_)) + ((!i_11_) & (!i_9_) & (sk[5]) & (i_10_) & (!i_15_)) + ((!i_11_) & (!i_9_) & (sk[5]) & (i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (!sk[5]) & (!i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (!sk[5]) & (!i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (!sk[5]) & (i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (!sk[5]) & (i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (sk[5]) & (!i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (sk[5]) & (!i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (sk[5]) & (i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (sk[5]) & (i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (!sk[5]) & (i_10_) & (!i_15_)) + ((i_11_) & (!i_9_) & (!sk[5]) & (i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (sk[5]) & (!i_10_) & (!i_15_)) + ((i_11_) & (!i_9_) & (sk[5]) & (!i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (sk[5]) & (i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (!sk[5]) & (!i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (!sk[5]) & (!i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (!sk[5]) & (i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (!sk[5]) & (i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (sk[5]) & (!i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (sk[5]) & (!i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (sk[5]) & (i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (sk[5]) & (i_10_) & (i_15_)));
	assign g116 = (((!g91) & (sk[6]) & (!g115)) + ((g91) & (!sk[6]) & (!g115)) + ((g91) & (!sk[6]) & (g115)));
	assign g117 = (((!sk[7]) & (g18) & (!g91)) + ((!sk[7]) & (g18) & (g91)) + ((sk[7]) & (!g18) & (!g91)));
	assign g118 = (((g31) & (!sk[8]) & (!g110)) + ((g31) & (!sk[8]) & (g110)) + ((g31) & (sk[8]) & (g110)));
	assign g119 = (((!i_11_) & (!i_9_) & (!sk[9]) & (i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (!sk[9]) & (!i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (!sk[9]) & (!i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (!sk[9]) & (i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (!sk[9]) & (i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (!sk[9]) & (i_10_) & (!i_15_)) + ((i_11_) & (!i_9_) & (!sk[9]) & (i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (!sk[9]) & (!i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (!sk[9]) & (!i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (!sk[9]) & (i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (!sk[9]) & (i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (sk[9]) & (!i_10_) & (!i_15_)));
	assign g120 = (((!g48) & (sk[10]) & (!g119)) + ((g48) & (!sk[10]) & (!g119)) + ((g48) & (!sk[10]) & (g119)) + ((g48) & (sk[10]) & (!g119)) + ((g48) & (sk[10]) & (g119)));
	assign g121 = (((g118) & (!g120) & (!sk[11]) & (!g90)) + ((g118) & (!g120) & (!sk[11]) & (g90)) + ((g118) & (!g120) & (sk[11]) & (!g90)) + ((g118) & (!g120) & (sk[11]) & (g90)) + ((g118) & (g120) & (!sk[11]) & (!g90)) + ((g118) & (g120) & (!sk[11]) & (g90)) + ((g118) & (g120) & (sk[11]) & (!g90)));
	assign g122 = (((!i_11_) & (!i_9_) & (!sk[12]) & (i_10_) & (i_15_)) + ((!i_11_) & (!i_9_) & (sk[12]) & (!i_10_) & (!i_15_)) + ((!i_11_) & (!i_9_) & (sk[12]) & (!i_10_) & (i_15_)) + ((!i_11_) & (!i_9_) & (sk[12]) & (i_10_) & (!i_15_)) + ((!i_11_) & (!i_9_) & (sk[12]) & (i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (!sk[12]) & (!i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (!sk[12]) & (!i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (!sk[12]) & (i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (!sk[12]) & (i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (sk[12]) & (!i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (sk[12]) & (!i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (sk[12]) & (i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (sk[12]) & (i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (!sk[12]) & (i_10_) & (!i_15_)) + ((i_11_) & (!i_9_) & (!sk[12]) & (i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (sk[12]) & (!i_10_) & (!i_15_)) + ((i_11_) & (!i_9_) & (sk[12]) & (!i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (sk[12]) & (i_10_) & (!i_15_)) + ((i_11_) & (!i_9_) & (sk[12]) & (i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (!sk[12]) & (!i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (!sk[12]) & (!i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (!sk[12]) & (i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (!sk[12]) & (i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (sk[12]) & (!i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (sk[12]) & (i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (sk[12]) & (i_10_) & (i_15_)));
	assign g123 = (((!g91) & (sk[13]) & (!g122)) + ((g91) & (!sk[13]) & (!g122)) + ((g91) & (!sk[13]) & (g122)));
	assign g124 = (((!sk[14]) & (!i_11_) & (!i_9_) & (i_10_) & (i_15_)) + ((!sk[14]) & (!i_11_) & (i_9_) & (!i_10_) & (!i_15_)) + ((!sk[14]) & (!i_11_) & (i_9_) & (!i_10_) & (i_15_)) + ((!sk[14]) & (!i_11_) & (i_9_) & (i_10_) & (!i_15_)) + ((!sk[14]) & (!i_11_) & (i_9_) & (i_10_) & (i_15_)) + ((!sk[14]) & (i_11_) & (!i_9_) & (i_10_) & (!i_15_)) + ((!sk[14]) & (i_11_) & (!i_9_) & (i_10_) & (i_15_)) + ((!sk[14]) & (i_11_) & (i_9_) & (!i_10_) & (!i_15_)) + ((!sk[14]) & (i_11_) & (i_9_) & (!i_10_) & (i_15_)) + ((!sk[14]) & (i_11_) & (i_9_) & (i_10_) & (!i_15_)) + ((!sk[14]) & (i_11_) & (i_9_) & (i_10_) & (i_15_)) + ((sk[14]) & (i_11_) & (i_9_) & (i_10_) & (i_15_)));
	assign g125 = (((!sk[15]) & (g91) & (!g124)) + ((!sk[15]) & (g91) & (g124)) + ((sk[15]) & (!g91) & (g124)));
	assign g126 = (((!g118) & (!g112) & (!g123) & (sk[16]) & (!g125)) + ((!g118) & (!g112) & (!g123) & (sk[16]) & (g125)) + ((!g118) & (!g112) & (g123) & (!sk[16]) & (g125)) + ((!g118) & (!g112) & (g123) & (sk[16]) & (!g125)) + ((!g118) & (!g112) & (g123) & (sk[16]) & (g125)) + ((!g118) & (g112) & (!g123) & (!sk[16]) & (!g125)) + ((!g118) & (g112) & (!g123) & (!sk[16]) & (g125)) + ((!g118) & (g112) & (!g123) & (sk[16]) & (!g125)) + ((!g118) & (g112) & (g123) & (!sk[16]) & (!g125)) + ((!g118) & (g112) & (g123) & (!sk[16]) & (g125)) + ((g118) & (!g112) & (!g123) & (sk[16]) & (!g125)) + ((g118) & (!g112) & (g123) & (!sk[16]) & (!g125)) + ((g118) & (!g112) & (g123) & (!sk[16]) & (g125)) + ((g118) & (!g112) & (g123) & (sk[16]) & (!g125)) + ((g118) & (g112) & (!g123) & (!sk[16]) & (!g125)) + ((g118) & (g112) & (!g123) & (!sk[16]) & (g125)) + ((g118) & (g112) & (!g123) & (sk[16]) & (!g125)) + ((g118) & (g112) & (g123) & (!sk[16]) & (!g125)) + ((g118) & (g112) & (g123) & (!sk[16]) & (g125)));
	assign g127 = (((!sk[17]) & (g22) & (!g91)) + ((!sk[17]) & (g22) & (g91)) + ((sk[17]) & (!g22) & (!g91)) + ((sk[17]) & (!g22) & (g91)) + ((sk[17]) & (g22) & (g91)));
	assign g128 = (((!sk[18]) & (g88) & (!g127) & (!g125)) + ((!sk[18]) & (g88) & (!g127) & (g125)) + ((!sk[18]) & (g88) & (g127) & (!g125)) + ((!sk[18]) & (g88) & (g127) & (g125)) + ((sk[18]) & (g88) & (!g127) & (!g125)) + ((sk[18]) & (g88) & (!g127) & (g125)) + ((sk[18]) & (g88) & (g127) & (g125)));
	assign g129 = (((!g89) & (!g116) & (!g117) & (!g121) & (g126) & (!g128)) + ((g89) & (!g116) & (!g117) & (!g121) & (g126) & (!g128)) + ((g89) & (!g116) & (g117) & (!g121) & (g126) & (!g128)) + ((g89) & (g116) & (!g117) & (!g121) & (g126) & (!g128)) + ((g89) & (g116) & (g117) & (!g121) & (g126) & (!g128)));
	assign g130 = (((!g99) & (!g101) & (!g109) & (!g112) & (!g114) & (g129)) + ((!g99) & (!g101) & (!g109) & (!g112) & (g114) & (g129)) + ((!g99) & (!g101) & (!g109) & (g112) & (!g114) & (g129)) + ((!g99) & (!g101) & (g109) & (!g112) & (!g114) & (g129)) + ((!g99) & (!g101) & (g109) & (g112) & (!g114) & (g129)) + ((!g99) & (g101) & (!g109) & (!g112) & (!g114) & (g129)) + ((!g99) & (g101) & (!g109) & (g112) & (!g114) & (g129)) + ((!g99) & (g101) & (g109) & (!g112) & (!g114) & (g129)) + ((!g99) & (g101) & (g109) & (g112) & (!g114) & (g129)) + ((g99) & (!g101) & (!g109) & (!g112) & (!g114) & (g129)) + ((g99) & (!g101) & (!g109) & (g112) & (!g114) & (g129)) + ((g99) & (!g101) & (g109) & (!g112) & (!g114) & (g129)) + ((g99) & (!g101) & (g109) & (g112) & (!g114) & (g129)) + ((g99) & (g101) & (!g109) & (!g112) & (!g114) & (g129)) + ((g99) & (g101) & (!g109) & (g112) & (!g114) & (g129)) + ((g99) & (g101) & (g109) & (!g112) & (!g114) & (g129)) + ((g99) & (g101) & (g109) & (g112) & (!g114) & (g129)));
	assign g131 = (((!sk[21]) & (g53) & (!g5)) + ((!sk[21]) & (g53) & (g5)) + ((sk[21]) & (g53) & (g5)));
	assign g132 = (((!sk[22]) & (g48) & (!g131)) + ((!sk[22]) & (g48) & (g131)) + ((sk[22]) & (!g48) & (!g131)) + ((sk[22]) & (g48) & (!g131)) + ((sk[22]) & (g48) & (g131)));
	assign g133 = (((!i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (!g91) & (!g109)) + ((!i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (!g91) & (g109)) + ((!i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (g91) & (!g109)) + ((!i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (g91) & (g109)) + ((!i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (!g91) & (!g109)) + ((!i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (g91) & (!g109)) + ((!i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (g91) & (g109)) + ((!i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (!g91) & (!g109)) + ((!i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (!g91) & (g109)) + ((!i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (g91) & (!g109)) + ((!i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (g91) & (g109)) + ((!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!g91) & (!g109)) + ((!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!g91) & (g109)) + ((!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g91) & (!g109)) + ((!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g91) & (g109)) + ((!i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (!g91) & (!g109)) + ((!i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (!g91) & (g109)) + ((!i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (g91) & (!g109)) + ((!i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (g91) & (g109)) + ((!i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!g91) & (!g109)) + ((!i_11_) & (i_9_) & (!i_10_) & (i_15_) & (g91) & (!g109)) + ((!i_11_) & (i_9_) & (!i_10_) & (i_15_) & (g91) & (g109)) + ((!i_11_) & (i_9_) & (i_10_) & (!i_15_) & (!g91) & (!g109)) + ((!i_11_) & (i_9_) & (i_10_) & (!i_15_) & (!g91) & (g109)) + ((!i_11_) & (i_9_) & (i_10_) & (!i_15_) & (g91) & (!g109)) + ((!i_11_) & (i_9_) & (i_10_) & (!i_15_) & (g91) & (g109)) + ((!i_11_) & (i_9_) & (i_10_) & (i_15_) & (!g91) & (!g109)) + ((!i_11_) & (i_9_) & (i_10_) & (i_15_) & (g91) & (!g109)) + ((!i_11_) & (i_9_) & (i_10_) & (i_15_) & (g91) & (g109)) + ((i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (!g91) & (!g109)) + ((i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (!g91) & (g109)) + ((i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (g91) & (!g109)) + ((i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (g91) & (g109)) + ((i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (!g91) & (!g109)) + ((i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (g91) & (!g109)) + ((i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (g91) & (g109)) + ((i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (!g91) & (!g109)) + ((i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (!g91) & (g109)) + ((i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (g91) & (!g109)) + ((i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (g91) & (g109)) + ((i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!g91) & (!g109)) + ((i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g91) & (!g109)) + ((i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g91) & (g109)) + ((i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (!g91) & (!g109)) + ((i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (!g91) & (g109)) + ((i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (g91) & (!g109)) + ((i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (g91) & (g109)) + ((i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!g91) & (!g109)) + ((i_11_) & (i_9_) & (!i_10_) & (i_15_) & (g91) & (!g109)) + ((i_11_) & (i_9_) & (!i_10_) & (i_15_) & (g91) & (g109)) + ((i_11_) & (i_9_) & (i_10_) & (!i_15_) & (!g91) & (!g109)) + ((i_11_) & (i_9_) & (i_10_) & (!i_15_) & (!g91) & (g109)) + ((i_11_) & (i_9_) & (i_10_) & (!i_15_) & (g91) & (!g109)) + ((i_11_) & (i_9_) & (i_10_) & (!i_15_) & (g91) & (g109)) + ((i_11_) & (i_9_) & (i_10_) & (i_15_) & (!g91) & (!g109)) + ((i_11_) & (i_9_) & (i_10_) & (i_15_) & (!g91) & (g109)) + ((i_11_) & (i_9_) & (i_10_) & (i_15_) & (g91) & (!g109)) + ((i_11_) & (i_9_) & (i_10_) & (i_15_) & (g91) & (g109)));
	assign g134 = (((g27) & (!sk[24]) & (!g58)) + ((g27) & (!sk[24]) & (g58)) + ((g27) & (sk[24]) & (g58)));
	assign g135 = (((i_6_) & (!i_7_) & (!sk[25]) & (!g58)) + ((i_6_) & (!i_7_) & (!sk[25]) & (g58)) + ((i_6_) & (!i_7_) & (sk[25]) & (g58)) + ((i_6_) & (i_7_) & (!sk[25]) & (!g58)) + ((i_6_) & (i_7_) & (!sk[25]) & (g58)));
	assign g136 = (((i_8_) & (!sk[26]) & (!g135)) + ((i_8_) & (!sk[26]) & (g135)) + ((i_8_) & (sk[26]) & (g135)));
	assign g137 = (((!g134) & (!g136) & (!g120) & (!g103) & (!g116) & (!g123)) + ((!g134) & (!g136) & (!g120) & (!g103) & (!g116) & (g123)) + ((!g134) & (!g136) & (!g120) & (!g103) & (g116) & (!g123)) + ((!g134) & (!g136) & (!g120) & (!g103) & (g116) & (g123)) + ((!g134) & (!g136) & (!g120) & (g103) & (!g116) & (!g123)) + ((!g134) & (!g136) & (!g120) & (g103) & (!g116) & (g123)) + ((!g134) & (!g136) & (!g120) & (g103) & (g116) & (!g123)) + ((!g134) & (!g136) & (!g120) & (g103) & (g116) & (g123)) + ((!g134) & (!g136) & (g120) & (!g103) & (!g116) & (!g123)) + ((!g134) & (!g136) & (g120) & (!g103) & (!g116) & (g123)) + ((!g134) & (!g136) & (g120) & (!g103) & (g116) & (!g123)) + ((!g134) & (!g136) & (g120) & (!g103) & (g116) & (g123)) + ((!g134) & (!g136) & (g120) & (g103) & (!g116) & (!g123)) + ((!g134) & (!g136) & (g120) & (g103) & (!g116) & (g123)) + ((!g134) & (!g136) & (g120) & (g103) & (g116) & (!g123)) + ((!g134) & (!g136) & (g120) & (g103) & (g116) & (g123)) + ((!g134) & (g136) & (g120) & (g103) & (!g116) & (!g123)) + ((!g134) & (g136) & (g120) & (g103) & (!g116) & (g123)) + ((g134) & (!g136) & (!g120) & (!g103) & (!g116) & (!g123)) + ((g134) & (!g136) & (!g120) & (!g103) & (g116) & (!g123)) + ((g134) & (!g136) & (!g120) & (g103) & (!g116) & (!g123)) + ((g134) & (!g136) & (!g120) & (g103) & (g116) & (!g123)) + ((g134) & (!g136) & (g120) & (!g103) & (!g116) & (!g123)) + ((g134) & (!g136) & (g120) & (!g103) & (g116) & (!g123)) + ((g134) & (!g136) & (g120) & (g103) & (!g116) & (!g123)) + ((g134) & (!g136) & (g120) & (g103) & (g116) & (!g123)) + ((g134) & (g136) & (g120) & (g103) & (!g116) & (!g123)));
	assign g138 = (((!g118) & (!sk[28]) & (!g94) & (g92) & (g116)) + ((!g118) & (!sk[28]) & (g94) & (!g92) & (!g116)) + ((!g118) & (!sk[28]) & (g94) & (!g92) & (g116)) + ((!g118) & (!sk[28]) & (g94) & (g92) & (!g116)) + ((!g118) & (!sk[28]) & (g94) & (g92) & (g116)) + ((g118) & (!sk[28]) & (!g94) & (g92) & (!g116)) + ((g118) & (!sk[28]) & (!g94) & (g92) & (g116)) + ((g118) & (!sk[28]) & (g94) & (!g92) & (!g116)) + ((g118) & (!sk[28]) & (g94) & (!g92) & (g116)) + ((g118) & (!sk[28]) & (g94) & (g92) & (!g116)) + ((g118) & (!sk[28]) & (g94) & (g92) & (g116)) + ((g118) & (sk[28]) & (!g94) & (!g92) & (!g116)) + ((g118) & (sk[28]) & (!g94) & (!g92) & (g116)) + ((g118) & (sk[28]) & (!g94) & (g92) & (g116)) + ((g118) & (sk[28]) & (g94) & (!g92) & (!g116)) + ((g118) & (sk[28]) & (g94) & (!g92) & (g116)) + ((g118) & (sk[28]) & (g94) & (g92) & (!g116)) + ((g118) & (sk[28]) & (g94) & (g92) & (g116)));
	assign g139 = (((!sk[29]) & (!g134) & (!g103) & (g96) & (g105)) + ((!sk[29]) & (!g134) & (g103) & (!g96) & (!g105)) + ((!sk[29]) & (!g134) & (g103) & (!g96) & (g105)) + ((!sk[29]) & (!g134) & (g103) & (g96) & (!g105)) + ((!sk[29]) & (!g134) & (g103) & (g96) & (g105)) + ((!sk[29]) & (g134) & (!g103) & (g96) & (!g105)) + ((!sk[29]) & (g134) & (!g103) & (g96) & (g105)) + ((!sk[29]) & (g134) & (g103) & (!g96) & (!g105)) + ((!sk[29]) & (g134) & (g103) & (!g96) & (g105)) + ((!sk[29]) & (g134) & (g103) & (g96) & (!g105)) + ((!sk[29]) & (g134) & (g103) & (g96) & (g105)) + ((sk[29]) & (g134) & (!g103) & (!g96) & (!g105)) + ((sk[29]) & (g134) & (!g103) & (!g96) & (g105)) + ((sk[29]) & (g134) & (!g103) & (g96) & (!g105)) + ((sk[29]) & (g134) & (!g103) & (g96) & (g105)) + ((sk[29]) & (g134) & (g103) & (!g96) & (!g105)) + ((sk[29]) & (g134) & (g103) & (!g96) & (g105)) + ((sk[29]) & (g134) & (g103) & (g96) & (g105)));
	assign g140 = (((!g134) & (!sk[30]) & (!g94) & (g116) & (g125)) + ((!g134) & (!sk[30]) & (g94) & (!g116) & (!g125)) + ((!g134) & (!sk[30]) & (g94) & (!g116) & (g125)) + ((!g134) & (!sk[30]) & (g94) & (g116) & (!g125)) + ((!g134) & (!sk[30]) & (g94) & (g116) & (g125)) + ((g134) & (!sk[30]) & (!g94) & (g116) & (!g125)) + ((g134) & (!sk[30]) & (!g94) & (g116) & (g125)) + ((g134) & (!sk[30]) & (g94) & (!g116) & (!g125)) + ((g134) & (!sk[30]) & (g94) & (!g116) & (g125)) + ((g134) & (!sk[30]) & (g94) & (g116) & (!g125)) + ((g134) & (!sk[30]) & (g94) & (g116) & (g125)) + ((g134) & (sk[30]) & (!g94) & (!g116) & (g125)) + ((g134) & (sk[30]) & (!g94) & (g116) & (!g125)) + ((g134) & (sk[30]) & (!g94) & (g116) & (g125)) + ((g134) & (sk[30]) & (g94) & (!g116) & (!g125)) + ((g134) & (sk[30]) & (g94) & (!g116) & (g125)) + ((g134) & (sk[30]) & (g94) & (g116) & (!g125)) + ((g134) & (sk[30]) & (g94) & (g116) & (g125)));
	assign g141 = (((!sk[31]) & (i_9_) & (!i_10_)) + ((!sk[31]) & (i_9_) & (i_10_)) + ((sk[31]) & (!i_9_) & (i_10_)));
	assign g142 = (((!sk[32]) & (!i_11_) & (!i_15_) & (g141) & (g48)) + ((!sk[32]) & (!i_11_) & (i_15_) & (!g141) & (!g48)) + ((!sk[32]) & (!i_11_) & (i_15_) & (!g141) & (g48)) + ((!sk[32]) & (!i_11_) & (i_15_) & (g141) & (!g48)) + ((!sk[32]) & (!i_11_) & (i_15_) & (g141) & (g48)) + ((!sk[32]) & (i_11_) & (!i_15_) & (g141) & (!g48)) + ((!sk[32]) & (i_11_) & (!i_15_) & (g141) & (g48)) + ((!sk[32]) & (i_11_) & (i_15_) & (!g141) & (!g48)) + ((!sk[32]) & (i_11_) & (i_15_) & (!g141) & (g48)) + ((!sk[32]) & (i_11_) & (i_15_) & (g141) & (!g48)) + ((!sk[32]) & (i_11_) & (i_15_) & (g141) & (g48)) + ((sk[32]) & (!i_11_) & (!i_15_) & (g141) & (!g48)));
	assign g143 = (((!sk[33]) & (!g59) & (!g134) & (!g99) & (!g142) & (g90)) + ((!sk[33]) & (!g59) & (!g134) & (!g99) & (g142) & (g90)) + ((!sk[33]) & (!g59) & (!g134) & (g99) & (!g142) & (g90)) + ((!sk[33]) & (!g59) & (!g134) & (g99) & (g142) & (g90)) + ((!sk[33]) & (!g59) & (g134) & (!g99) & (!g142) & (g90)) + ((!sk[33]) & (!g59) & (g134) & (!g99) & (g142) & (g90)) + ((!sk[33]) & (!g59) & (g134) & (g99) & (!g142) & (g90)) + ((!sk[33]) & (!g59) & (g134) & (g99) & (g142) & (g90)) + ((!sk[33]) & (g59) & (!g134) & (!g99) & (!g142) & (!g90)) + ((!sk[33]) & (g59) & (!g134) & (!g99) & (!g142) & (g90)) + ((!sk[33]) & (g59) & (!g134) & (!g99) & (g142) & (!g90)) + ((!sk[33]) & (g59) & (!g134) & (!g99) & (g142) & (g90)) + ((!sk[33]) & (g59) & (!g134) & (g99) & (!g142) & (!g90)) + ((!sk[33]) & (g59) & (!g134) & (g99) & (!g142) & (g90)) + ((!sk[33]) & (g59) & (!g134) & (g99) & (g142) & (!g90)) + ((!sk[33]) & (g59) & (!g134) & (g99) & (g142) & (g90)) + ((!sk[33]) & (g59) & (g134) & (!g99) & (!g142) & (!g90)) + ((!sk[33]) & (g59) & (g134) & (!g99) & (!g142) & (g90)) + ((!sk[33]) & (g59) & (g134) & (!g99) & (g142) & (!g90)) + ((!sk[33]) & (g59) & (g134) & (!g99) & (g142) & (g90)) + ((!sk[33]) & (g59) & (g134) & (g99) & (!g142) & (!g90)) + ((!sk[33]) & (g59) & (g134) & (g99) & (!g142) & (g90)) + ((!sk[33]) & (g59) & (g134) & (g99) & (g142) & (!g90)) + ((!sk[33]) & (g59) & (g134) & (g99) & (g142) & (g90)) + ((sk[33]) & (!g59) & (!g134) & (!g99) & (!g142) & (!g90)) + ((sk[33]) & (!g59) & (!g134) & (!g99) & (!g142) & (g90)) + ((sk[33]) & (!g59) & (!g134) & (!g99) & (g142) & (!g90)) + ((sk[33]) & (!g59) & (!g134) & (!g99) & (g142) & (g90)) + ((sk[33]) & (!g59) & (!g134) & (g99) & (!g142) & (g90)) + ((sk[33]) & (!g59) & (!g134) & (g99) & (g142) & (g90)) + ((sk[33]) & (!g59) & (g134) & (!g99) & (!g142) & (g90)) + ((sk[33]) & (!g59) & (g134) & (g99) & (!g142) & (g90)) + ((sk[33]) & (g59) & (!g134) & (!g99) & (!g142) & (g90)) + ((sk[33]) & (g59) & (!g134) & (g99) & (!g142) & (g90)) + ((sk[33]) & (g59) & (g134) & (!g99) & (!g142) & (g90)) + ((sk[33]) & (g59) & (g134) & (g99) & (!g142) & (g90)));
	assign g144 = (((!g138) & (!g139) & (!sk[34]) & (g140) & (g143)) + ((!g138) & (!g139) & (sk[34]) & (!g140) & (g143)) + ((!g138) & (g139) & (!sk[34]) & (!g140) & (!g143)) + ((!g138) & (g139) & (!sk[34]) & (!g140) & (g143)) + ((!g138) & (g139) & (!sk[34]) & (g140) & (!g143)) + ((!g138) & (g139) & (!sk[34]) & (g140) & (g143)) + ((g138) & (!g139) & (!sk[34]) & (g140) & (!g143)) + ((g138) & (!g139) & (!sk[34]) & (g140) & (g143)) + ((g138) & (g139) & (!sk[34]) & (!g140) & (!g143)) + ((g138) & (g139) & (!sk[34]) & (!g140) & (g143)) + ((g138) & (g139) & (!sk[34]) & (g140) & (!g143)) + ((g138) & (g139) & (!sk[34]) & (g140) & (g143)));
	assign g145 = (((!sk[35]) & (i_8_) & (!g108)) + ((!sk[35]) & (i_8_) & (g108)) + ((sk[35]) & (i_8_) & (g108)));
	assign g146 = (((!i_8_) & (!g88) & (sk[36]) & (!g112)) + ((!i_8_) & (g88) & (sk[36]) & (!g112)) + ((i_8_) & (!g88) & (!sk[36]) & (!g112)) + ((i_8_) & (!g88) & (!sk[36]) & (g112)) + ((i_8_) & (!g88) & (sk[36]) & (!g112)) + ((i_8_) & (g88) & (!sk[36]) & (!g112)) + ((i_8_) & (g88) & (!sk[36]) & (g112)));
	assign g147 = (((!g145) & (!g146) & (!g127) & (!g125) & (!g114) & (!g105)) + ((!g145) & (!g146) & (!g127) & (!g125) & (g114) & (!g105)) + ((!g145) & (!g146) & (!g127) & (g125) & (!g114) & (!g105)) + ((!g145) & (!g146) & (!g127) & (g125) & (g114) & (!g105)) + ((!g145) & (!g146) & (g127) & (!g125) & (!g114) & (!g105)) + ((!g145) & (!g146) & (g127) & (!g125) & (g114) & (!g105)) + ((!g145) & (!g146) & (g127) & (g125) & (!g114) & (!g105)) + ((!g145) & (!g146) & (g127) & (g125) & (g114) & (!g105)) + ((!g145) & (g146) & (!g127) & (!g125) & (!g114) & (!g105)) + ((!g145) & (g146) & (!g127) & (!g125) & (!g114) & (g105)) + ((!g145) & (g146) & (!g127) & (!g125) & (g114) & (!g105)) + ((!g145) & (g146) & (!g127) & (!g125) & (g114) & (g105)) + ((!g145) & (g146) & (!g127) & (g125) & (!g114) & (!g105)) + ((!g145) & (g146) & (!g127) & (g125) & (!g114) & (g105)) + ((!g145) & (g146) & (!g127) & (g125) & (g114) & (!g105)) + ((!g145) & (g146) & (!g127) & (g125) & (g114) & (g105)) + ((!g145) & (g146) & (g127) & (!g125) & (!g114) & (!g105)) + ((!g145) & (g146) & (g127) & (!g125) & (!g114) & (g105)) + ((!g145) & (g146) & (g127) & (!g125) & (g114) & (!g105)) + ((!g145) & (g146) & (g127) & (!g125) & (g114) & (g105)) + ((!g145) & (g146) & (g127) & (g125) & (!g114) & (!g105)) + ((!g145) & (g146) & (g127) & (g125) & (!g114) & (g105)) + ((!g145) & (g146) & (g127) & (g125) & (g114) & (!g105)) + ((!g145) & (g146) & (g127) & (g125) & (g114) & (g105)) + ((g145) & (!g146) & (g127) & (!g125) & (!g114) & (!g105)) + ((g145) & (g146) & (g127) & (!g125) & (!g114) & (!g105)));
	assign g148 = (((!g118) & (!g127) & (!g117) & (g137) & (g144) & (g147)) + ((!g118) & (!g127) & (g117) & (g137) & (g144) & (g147)) + ((!g118) & (g127) & (!g117) & (g137) & (g144) & (g147)) + ((!g118) & (g127) & (g117) & (g137) & (g144) & (g147)) + ((g118) & (g127) & (!g117) & (g137) & (g144) & (g147)));
	assign g149 = (((!sk[39]) & (g27) & (!g98)) + ((!sk[39]) & (g27) & (g98)) + ((sk[39]) & (g27) & (g98)));
	assign g150 = (((!sk[40]) & (g149) & (!g127) & (!g114)) + ((!sk[40]) & (g149) & (!g127) & (g114)) + ((!sk[40]) & (g149) & (g127) & (!g114)) + ((!sk[40]) & (g149) & (g127) & (g114)) + ((sk[40]) & (g149) & (!g127) & (!g114)) + ((sk[40]) & (g149) & (!g127) & (g114)) + ((sk[40]) & (g149) & (g127) & (g114)));
	assign g151 = (((!sk[41]) & (i_8_) & (!g88)) + ((!sk[41]) & (i_8_) & (g88)) + ((sk[41]) & (i_8_) & (g88)));
	assign g152 = (((g99) & (!g142) & (!sk[42]) & (!g117)) + ((g99) & (!g142) & (!sk[42]) & (g117)) + ((g99) & (!g142) & (sk[42]) & (g117)) + ((g99) & (g142) & (!sk[42]) & (!g117)) + ((g99) & (g142) & (!sk[42]) & (g117)) + ((g99) & (g142) & (sk[42]) & (!g117)) + ((g99) & (g142) & (sk[42]) & (g117)));
	assign g153 = (((g134) & (!g127) & (!sk[43]) & (!g114)) + ((g134) & (!g127) & (!sk[43]) & (g114)) + ((g134) & (!g127) & (sk[43]) & (!g114)) + ((g134) & (!g127) & (sk[43]) & (g114)) + ((g134) & (g127) & (!sk[43]) & (!g114)) + ((g134) & (g127) & (!sk[43]) & (g114)) + ((g134) & (g127) & (sk[43]) & (g114)));
	assign g154 = (((!g136) & (!sk[44]) & (!g151) & (!g114) & (!g152) & (g153)) + ((!g136) & (!sk[44]) & (!g151) & (!g114) & (g152) & (g153)) + ((!g136) & (!sk[44]) & (!g151) & (g114) & (!g152) & (g153)) + ((!g136) & (!sk[44]) & (!g151) & (g114) & (g152) & (g153)) + ((!g136) & (!sk[44]) & (g151) & (!g114) & (!g152) & (g153)) + ((!g136) & (!sk[44]) & (g151) & (!g114) & (g152) & (g153)) + ((!g136) & (!sk[44]) & (g151) & (g114) & (!g152) & (g153)) + ((!g136) & (!sk[44]) & (g151) & (g114) & (g152) & (g153)) + ((!g136) & (sk[44]) & (!g151) & (!g114) & (!g152) & (!g153)) + ((!g136) & (sk[44]) & (!g151) & (g114) & (!g152) & (!g153)) + ((!g136) & (sk[44]) & (g151) & (!g114) & (!g152) & (!g153)) + ((g136) & (!sk[44]) & (!g151) & (!g114) & (!g152) & (!g153)) + ((g136) & (!sk[44]) & (!g151) & (!g114) & (!g152) & (g153)) + ((g136) & (!sk[44]) & (!g151) & (!g114) & (g152) & (!g153)) + ((g136) & (!sk[44]) & (!g151) & (!g114) & (g152) & (g153)) + ((g136) & (!sk[44]) & (!g151) & (g114) & (!g152) & (!g153)) + ((g136) & (!sk[44]) & (!g151) & (g114) & (!g152) & (g153)) + ((g136) & (!sk[44]) & (!g151) & (g114) & (g152) & (!g153)) + ((g136) & (!sk[44]) & (!g151) & (g114) & (g152) & (g153)) + ((g136) & (!sk[44]) & (g151) & (!g114) & (!g152) & (!g153)) + ((g136) & (!sk[44]) & (g151) & (!g114) & (!g152) & (g153)) + ((g136) & (!sk[44]) & (g151) & (!g114) & (g152) & (!g153)) + ((g136) & (!sk[44]) & (g151) & (!g114) & (g152) & (g153)) + ((g136) & (!sk[44]) & (g151) & (g114) & (!g152) & (!g153)) + ((g136) & (!sk[44]) & (g151) & (g114) & (!g152) & (g153)) + ((g136) & (!sk[44]) & (g151) & (g114) & (g152) & (!g153)) + ((g136) & (!sk[44]) & (g151) & (g114) & (g152) & (g153)) + ((g136) & (sk[44]) & (!g151) & (!g114) & (!g152) & (!g153)) + ((g136) & (sk[44]) & (g151) & (!g114) & (!g152) & (!g153)));
	assign g155 = (((!i_8_) & (!g100) & (!g108) & (!g142) & (!sk[45]) & (g117)) + ((!i_8_) & (!g100) & (!g108) & (g142) & (!sk[45]) & (g117)) + ((!i_8_) & (!g100) & (g108) & (!g142) & (!sk[45]) & (g117)) + ((!i_8_) & (!g100) & (g108) & (!g142) & (sk[45]) & (g117)) + ((!i_8_) & (!g100) & (g108) & (g142) & (!sk[45]) & (g117)) + ((!i_8_) & (!g100) & (g108) & (g142) & (sk[45]) & (!g117)) + ((!i_8_) & (!g100) & (g108) & (g142) & (sk[45]) & (g117)) + ((!i_8_) & (g100) & (!g108) & (!g142) & (!sk[45]) & (g117)) + ((!i_8_) & (g100) & (!g108) & (g142) & (!sk[45]) & (g117)) + ((!i_8_) & (g100) & (g108) & (!g142) & (!sk[45]) & (g117)) + ((!i_8_) & (g100) & (g108) & (!g142) & (sk[45]) & (g117)) + ((!i_8_) & (g100) & (g108) & (g142) & (!sk[45]) & (g117)) + ((!i_8_) & (g100) & (g108) & (g142) & (sk[45]) & (!g117)) + ((!i_8_) & (g100) & (g108) & (g142) & (sk[45]) & (g117)) + ((i_8_) & (!g100) & (!g108) & (!g142) & (!sk[45]) & (!g117)) + ((i_8_) & (!g100) & (!g108) & (!g142) & (!sk[45]) & (g117)) + ((i_8_) & (!g100) & (!g108) & (g142) & (!sk[45]) & (!g117)) + ((i_8_) & (!g100) & (!g108) & (g142) & (!sk[45]) & (g117)) + ((i_8_) & (!g100) & (g108) & (!g142) & (!sk[45]) & (!g117)) + ((i_8_) & (!g100) & (g108) & (!g142) & (!sk[45]) & (g117)) + ((i_8_) & (!g100) & (g108) & (g142) & (!sk[45]) & (!g117)) + ((i_8_) & (!g100) & (g108) & (g142) & (!sk[45]) & (g117)) + ((i_8_) & (g100) & (!g108) & (!g142) & (!sk[45]) & (!g117)) + ((i_8_) & (g100) & (!g108) & (!g142) & (!sk[45]) & (g117)) + ((i_8_) & (g100) & (!g108) & (g142) & (!sk[45]) & (!g117)) + ((i_8_) & (g100) & (!g108) & (g142) & (!sk[45]) & (g117)) + ((i_8_) & (g100) & (!g108) & (g142) & (sk[45]) & (!g117)) + ((i_8_) & (g100) & (!g108) & (g142) & (sk[45]) & (g117)) + ((i_8_) & (g100) & (g108) & (!g142) & (!sk[45]) & (!g117)) + ((i_8_) & (g100) & (g108) & (!g142) & (!sk[45]) & (g117)) + ((i_8_) & (g100) & (g108) & (g142) & (!sk[45]) & (!g117)) + ((i_8_) & (g100) & (g108) & (g142) & (!sk[45]) & (g117)) + ((i_8_) & (g100) & (g108) & (g142) & (sk[45]) & (!g117)) + ((i_8_) & (g100) & (g108) & (g142) & (sk[45]) & (g117)));
	assign g156 = (((!g109) & (!g136) & (!g125) & (!sk[46]) & (!g105) & (g155)) + ((!g109) & (!g136) & (!g125) & (!sk[46]) & (g105) & (g155)) + ((!g109) & (!g136) & (!g125) & (sk[46]) & (!g105) & (!g155)) + ((!g109) & (!g136) & (!g125) & (sk[46]) & (g105) & (!g155)) + ((!g109) & (!g136) & (g125) & (!sk[46]) & (!g105) & (g155)) + ((!g109) & (!g136) & (g125) & (!sk[46]) & (g105) & (g155)) + ((!g109) & (!g136) & (g125) & (sk[46]) & (!g105) & (!g155)) + ((!g109) & (!g136) & (g125) & (sk[46]) & (g105) & (!g155)) + ((!g109) & (g136) & (!g125) & (!sk[46]) & (!g105) & (g155)) + ((!g109) & (g136) & (!g125) & (!sk[46]) & (g105) & (g155)) + ((!g109) & (g136) & (!g125) & (sk[46]) & (!g105) & (!g155)) + ((!g109) & (g136) & (g125) & (!sk[46]) & (!g105) & (g155)) + ((!g109) & (g136) & (g125) & (!sk[46]) & (g105) & (g155)) + ((!g109) & (g136) & (g125) & (sk[46]) & (!g105) & (!g155)) + ((g109) & (!g136) & (!g125) & (!sk[46]) & (!g105) & (!g155)) + ((g109) & (!g136) & (!g125) & (!sk[46]) & (!g105) & (g155)) + ((g109) & (!g136) & (!g125) & (!sk[46]) & (g105) & (!g155)) + ((g109) & (!g136) & (!g125) & (!sk[46]) & (g105) & (g155)) + ((g109) & (!g136) & (!g125) & (sk[46]) & (!g105) & (!g155)) + ((g109) & (!g136) & (g125) & (!sk[46]) & (!g105) & (!g155)) + ((g109) & (!g136) & (g125) & (!sk[46]) & (!g105) & (g155)) + ((g109) & (!g136) & (g125) & (!sk[46]) & (g105) & (!g155)) + ((g109) & (!g136) & (g125) & (!sk[46]) & (g105) & (g155)) + ((g109) & (g136) & (!g125) & (!sk[46]) & (!g105) & (!g155)) + ((g109) & (g136) & (!g125) & (!sk[46]) & (!g105) & (g155)) + ((g109) & (g136) & (!g125) & (!sk[46]) & (g105) & (!g155)) + ((g109) & (g136) & (!g125) & (!sk[46]) & (g105) & (g155)) + ((g109) & (g136) & (!g125) & (sk[46]) & (!g105) & (!g155)) + ((g109) & (g136) & (g125) & (!sk[46]) & (!g105) & (!g155)) + ((g109) & (g136) & (g125) & (!sk[46]) & (!g105) & (g155)) + ((g109) & (g136) & (g125) & (!sk[46]) & (g105) & (!g155)) + ((g109) & (g136) & (g125) & (!sk[46]) & (g105) & (g155)));
	assign g157 = (((!g136) & (!g125) & (!g150) & (!g154) & (!sk[47]) & (g156)) + ((!g136) & (!g125) & (!g150) & (g154) & (!sk[47]) & (g156)) + ((!g136) & (!g125) & (!g150) & (g154) & (sk[47]) & (g156)) + ((!g136) & (!g125) & (g150) & (!g154) & (!sk[47]) & (g156)) + ((!g136) & (!g125) & (g150) & (g154) & (!sk[47]) & (g156)) + ((!g136) & (g125) & (!g150) & (!g154) & (!sk[47]) & (g156)) + ((!g136) & (g125) & (!g150) & (g154) & (!sk[47]) & (g156)) + ((!g136) & (g125) & (!g150) & (g154) & (sk[47]) & (g156)) + ((!g136) & (g125) & (g150) & (!g154) & (!sk[47]) & (g156)) + ((!g136) & (g125) & (g150) & (g154) & (!sk[47]) & (g156)) + ((g136) & (!g125) & (!g150) & (!g154) & (!sk[47]) & (!g156)) + ((g136) & (!g125) & (!g150) & (!g154) & (!sk[47]) & (g156)) + ((g136) & (!g125) & (!g150) & (g154) & (!sk[47]) & (!g156)) + ((g136) & (!g125) & (!g150) & (g154) & (!sk[47]) & (g156)) + ((g136) & (!g125) & (!g150) & (g154) & (sk[47]) & (g156)) + ((g136) & (!g125) & (g150) & (!g154) & (!sk[47]) & (!g156)) + ((g136) & (!g125) & (g150) & (!g154) & (!sk[47]) & (g156)) + ((g136) & (!g125) & (g150) & (g154) & (!sk[47]) & (!g156)) + ((g136) & (!g125) & (g150) & (g154) & (!sk[47]) & (g156)) + ((g136) & (g125) & (!g150) & (!g154) & (!sk[47]) & (!g156)) + ((g136) & (g125) & (!g150) & (!g154) & (!sk[47]) & (g156)) + ((g136) & (g125) & (!g150) & (g154) & (!sk[47]) & (!g156)) + ((g136) & (g125) & (!g150) & (g154) & (!sk[47]) & (g156)) + ((g136) & (g125) & (g150) & (!g154) & (!sk[47]) & (!g156)) + ((g136) & (g125) & (g150) & (!g154) & (!sk[47]) & (g156)) + ((g136) & (g125) & (g150) & (g154) & (!sk[47]) & (!g156)) + ((g136) & (g125) & (g150) & (g154) & (!sk[47]) & (g156)));
	assign g158 = (((!i_11_) & (!i_9_) & (!i_10_) & (sk[48]) & (i_15_)) + ((!i_11_) & (!i_9_) & (i_10_) & (!sk[48]) & (i_15_)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[48]) & (!i_15_)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[48]) & (i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[48]) & (!i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[48]) & (i_15_)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[48]) & (!i_15_)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[48]) & (i_15_)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[48]) & (!i_15_)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[48]) & (i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[48]) & (!i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[48]) & (i_15_)));
	assign g159 = (((!sk[49]) & (g91) & (!g158)) + ((!sk[49]) & (g91) & (g158)) + ((sk[49]) & (!g91) & (g158)));
	assign g160 = (((!g134) & (!g118) & (!g145) & (!g151) & (!g159) & (!g96)) + ((!g134) & (!g118) & (!g145) & (!g151) & (!g159) & (g96)) + ((!g134) & (!g118) & (!g145) & (!g151) & (g159) & (!g96)) + ((!g134) & (!g118) & (!g145) & (!g151) & (g159) & (g96)) + ((!g134) & (!g118) & (!g145) & (g151) & (!g159) & (g96)) + ((!g134) & (!g118) & (!g145) & (g151) & (g159) & (g96)) + ((!g134) & (!g118) & (g145) & (!g151) & (!g159) & (!g96)) + ((!g134) & (!g118) & (g145) & (!g151) & (!g159) & (g96)) + ((!g134) & (!g118) & (g145) & (g151) & (!g159) & (g96)) + ((!g134) & (g118) & (!g145) & (!g151) & (!g159) & (g96)) + ((!g134) & (g118) & (!g145) & (!g151) & (g159) & (g96)) + ((!g134) & (g118) & (!g145) & (g151) & (!g159) & (g96)) + ((!g134) & (g118) & (!g145) & (g151) & (g159) & (g96)) + ((!g134) & (g118) & (g145) & (!g151) & (!g159) & (g96)) + ((!g134) & (g118) & (g145) & (g151) & (!g159) & (g96)) + ((g134) & (!g118) & (!g145) & (!g151) & (!g159) & (!g96)) + ((g134) & (!g118) & (!g145) & (!g151) & (!g159) & (g96)) + ((g134) & (!g118) & (!g145) & (g151) & (!g159) & (g96)) + ((g134) & (!g118) & (g145) & (!g151) & (!g159) & (!g96)) + ((g134) & (!g118) & (g145) & (!g151) & (!g159) & (g96)) + ((g134) & (!g118) & (g145) & (g151) & (!g159) & (g96)) + ((g134) & (g118) & (!g145) & (!g151) & (!g159) & (g96)) + ((g134) & (g118) & (!g145) & (g151) & (!g159) & (g96)) + ((g134) & (g118) & (g145) & (!g151) & (!g159) & (g96)) + ((g134) & (g118) & (g145) & (g151) & (!g159) & (g96)));
	assign g161 = (((!i_8_) & (!g135) & (!sk[51]) & (g92) & (g123)) + ((!i_8_) & (g135) & (!sk[51]) & (!g92) & (!g123)) + ((!i_8_) & (g135) & (!sk[51]) & (!g92) & (g123)) + ((!i_8_) & (g135) & (!sk[51]) & (g92) & (!g123)) + ((!i_8_) & (g135) & (!sk[51]) & (g92) & (g123)) + ((!i_8_) & (g135) & (sk[51]) & (!g92) & (!g123)) + ((!i_8_) & (g135) & (sk[51]) & (!g92) & (g123)) + ((i_8_) & (!g135) & (!sk[51]) & (g92) & (!g123)) + ((i_8_) & (!g135) & (!sk[51]) & (g92) & (g123)) + ((i_8_) & (g135) & (!sk[51]) & (!g92) & (!g123)) + ((i_8_) & (g135) & (!sk[51]) & (!g92) & (g123)) + ((i_8_) & (g135) & (!sk[51]) & (g92) & (!g123)) + ((i_8_) & (g135) & (!sk[51]) & (g92) & (g123)) + ((i_8_) & (g135) & (sk[51]) & (!g92) & (!g123)) + ((i_8_) & (g135) & (sk[51]) & (!g92) & (g123)) + ((i_8_) & (g135) & (sk[51]) & (g92) & (g123)));
	assign g162 = (((!i_11_) & (!i_9_) & (!i_10_) & (!sk[52]) & (!i_15_) & (g48)) + ((!i_11_) & (!i_9_) & (!i_10_) & (!sk[52]) & (i_15_) & (g48)) + ((!i_11_) & (!i_9_) & (!i_10_) & (sk[52]) & (!i_15_) & (!g48)) + ((!i_11_) & (!i_9_) & (i_10_) & (!sk[52]) & (!i_15_) & (g48)) + ((!i_11_) & (!i_9_) & (i_10_) & (!sk[52]) & (i_15_) & (g48)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[52]) & (!i_15_) & (g48)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[52]) & (i_15_) & (g48)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[52]) & (!i_15_) & (g48)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[52]) & (i_15_) & (g48)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[52]) & (!i_15_) & (!g48)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[52]) & (!i_15_) & (g48)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[52]) & (i_15_) & (!g48)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[52]) & (i_15_) & (g48)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[52]) & (!i_15_) & (!g48)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[52]) & (!i_15_) & (g48)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[52]) & (i_15_) & (!g48)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[52]) & (i_15_) & (g48)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[52]) & (!i_15_) & (!g48)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[52]) & (!i_15_) & (g48)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[52]) & (i_15_) & (!g48)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[52]) & (i_15_) & (g48)) + ((i_11_) & (i_9_) & (!i_10_) & (sk[52]) & (!i_15_) & (!g48)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[52]) & (!i_15_) & (!g48)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[52]) & (!i_15_) & (g48)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[52]) & (i_15_) & (!g48)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[52]) & (i_15_) & (g48)));
	assign g163 = (((!i_8_) & (!g88) & (!sk[53]) & (g108) & (g90)) + ((!i_8_) & (!g88) & (sk[53]) & (g108) & (!g90)) + ((!i_8_) & (g88) & (!sk[53]) & (!g108) & (!g90)) + ((!i_8_) & (g88) & (!sk[53]) & (!g108) & (g90)) + ((!i_8_) & (g88) & (!sk[53]) & (g108) & (!g90)) + ((!i_8_) & (g88) & (!sk[53]) & (g108) & (g90)) + ((!i_8_) & (g88) & (sk[53]) & (g108) & (!g90)) + ((i_8_) & (!g88) & (!sk[53]) & (g108) & (!g90)) + ((i_8_) & (!g88) & (!sk[53]) & (g108) & (g90)) + ((i_8_) & (!g88) & (sk[53]) & (g108) & (!g90)) + ((i_8_) & (g88) & (!sk[53]) & (!g108) & (!g90)) + ((i_8_) & (g88) & (!sk[53]) & (!g108) & (g90)) + ((i_8_) & (g88) & (!sk[53]) & (g108) & (!g90)) + ((i_8_) & (g88) & (!sk[53]) & (g108) & (g90)) + ((i_8_) & (g88) & (sk[53]) & (!g108) & (!g90)) + ((i_8_) & (g88) & (sk[53]) & (g108) & (!g90)));
	assign g164 = (((!sk[54]) & (i_15_) & (!g141)) + ((!sk[54]) & (i_15_) & (g141)) + ((sk[54]) & (i_15_) & (g141)));
	assign g165 = (((!g91) & (sk[55]) & (g164)) + ((g91) & (!sk[55]) & (!g164)) + ((g91) & (!sk[55]) & (g164)));
	assign g166 = (((!g100) & (!g112) & (!sk[56]) & (g127) & (g165)) + ((!g100) & (!g112) & (sk[56]) & (!g127) & (!g165)) + ((!g100) & (!g112) & (sk[56]) & (!g127) & (g165)) + ((!g100) & (!g112) & (sk[56]) & (g127) & (!g165)) + ((!g100) & (!g112) & (sk[56]) & (g127) & (g165)) + ((!g100) & (g112) & (!sk[56]) & (!g127) & (!g165)) + ((!g100) & (g112) & (!sk[56]) & (!g127) & (g165)) + ((!g100) & (g112) & (!sk[56]) & (g127) & (!g165)) + ((!g100) & (g112) & (!sk[56]) & (g127) & (g165)) + ((!g100) & (g112) & (sk[56]) & (g127) & (!g165)) + ((g100) & (!g112) & (!sk[56]) & (g127) & (!g165)) + ((g100) & (!g112) & (!sk[56]) & (g127) & (g165)) + ((g100) & (!g112) & (sk[56]) & (g127) & (!g165)) + ((g100) & (!g112) & (sk[56]) & (g127) & (g165)) + ((g100) & (g112) & (!sk[56]) & (!g127) & (!g165)) + ((g100) & (g112) & (!sk[56]) & (!g127) & (g165)) + ((g100) & (g112) & (!sk[56]) & (g127) & (!g165)) + ((g100) & (g112) & (!sk[56]) & (g127) & (g165)) + ((g100) & (g112) & (sk[56]) & (g127) & (!g165)));
	assign g167 = (((!g134) & (!g117) & (!sk[57]) & (!g162) & (!g163) & (g166)) + ((!g134) & (!g117) & (!sk[57]) & (!g162) & (g163) & (g166)) + ((!g134) & (!g117) & (!sk[57]) & (g162) & (!g163) & (g166)) + ((!g134) & (!g117) & (!sk[57]) & (g162) & (g163) & (g166)) + ((!g134) & (!g117) & (sk[57]) & (!g162) & (!g163) & (g166)) + ((!g134) & (!g117) & (sk[57]) & (g162) & (!g163) & (g166)) + ((!g134) & (g117) & (!sk[57]) & (!g162) & (!g163) & (g166)) + ((!g134) & (g117) & (!sk[57]) & (!g162) & (g163) & (g166)) + ((!g134) & (g117) & (!sk[57]) & (g162) & (!g163) & (g166)) + ((!g134) & (g117) & (!sk[57]) & (g162) & (g163) & (g166)) + ((!g134) & (g117) & (sk[57]) & (!g162) & (!g163) & (g166)) + ((!g134) & (g117) & (sk[57]) & (g162) & (!g163) & (g166)) + ((g134) & (!g117) & (!sk[57]) & (!g162) & (!g163) & (!g166)) + ((g134) & (!g117) & (!sk[57]) & (!g162) & (!g163) & (g166)) + ((g134) & (!g117) & (!sk[57]) & (!g162) & (g163) & (!g166)) + ((g134) & (!g117) & (!sk[57]) & (!g162) & (g163) & (g166)) + ((g134) & (!g117) & (!sk[57]) & (g162) & (!g163) & (!g166)) + ((g134) & (!g117) & (!sk[57]) & (g162) & (!g163) & (g166)) + ((g134) & (!g117) & (!sk[57]) & (g162) & (g163) & (!g166)) + ((g134) & (!g117) & (!sk[57]) & (g162) & (g163) & (g166)) + ((g134) & (!g117) & (sk[57]) & (!g162) & (!g163) & (g166)) + ((g134) & (g117) & (!sk[57]) & (!g162) & (!g163) & (!g166)) + ((g134) & (g117) & (!sk[57]) & (!g162) & (!g163) & (g166)) + ((g134) & (g117) & (!sk[57]) & (!g162) & (g163) & (!g166)) + ((g134) & (g117) & (!sk[57]) & (!g162) & (g163) & (g166)) + ((g134) & (g117) & (!sk[57]) & (g162) & (!g163) & (!g166)) + ((g134) & (g117) & (!sk[57]) & (g162) & (!g163) & (g166)) + ((g134) & (g117) & (!sk[57]) & (g162) & (g163) & (!g166)) + ((g134) & (g117) & (!sk[57]) & (g162) & (g163) & (g166)));
	assign g168 = (((!g160) & (!g1775) & (g161) & (!sk[58]) & (g167)) + ((!g160) & (g1775) & (!g161) & (!sk[58]) & (!g167)) + ((!g160) & (g1775) & (!g161) & (!sk[58]) & (g167)) + ((!g160) & (g1775) & (g161) & (!sk[58]) & (!g167)) + ((!g160) & (g1775) & (g161) & (!sk[58]) & (g167)) + ((g160) & (!g1775) & (g161) & (!sk[58]) & (!g167)) + ((g160) & (!g1775) & (g161) & (!sk[58]) & (g167)) + ((g160) & (g1775) & (!g161) & (!sk[58]) & (!g167)) + ((g160) & (g1775) & (!g161) & (!sk[58]) & (g167)) + ((g160) & (g1775) & (!g161) & (sk[58]) & (g167)) + ((g160) & (g1775) & (g161) & (!sk[58]) & (!g167)) + ((g160) & (g1775) & (g161) & (!sk[58]) & (g167)));
	assign g169 = (((g107) & (g130) & (g1782) & (g148) & (g157) & (g168)));
	assign g170 = (((!i_14_) & (!sk[60]) & (!i_12_) & (!i_13_) & (!g102) & (g119)) + ((!i_14_) & (!sk[60]) & (!i_12_) & (!i_13_) & (g102) & (g119)) + ((!i_14_) & (!sk[60]) & (!i_12_) & (i_13_) & (!g102) & (g119)) + ((!i_14_) & (!sk[60]) & (!i_12_) & (i_13_) & (g102) & (g119)) + ((!i_14_) & (!sk[60]) & (i_12_) & (!i_13_) & (!g102) & (g119)) + ((!i_14_) & (!sk[60]) & (i_12_) & (!i_13_) & (g102) & (g119)) + ((!i_14_) & (!sk[60]) & (i_12_) & (i_13_) & (!g102) & (g119)) + ((!i_14_) & (!sk[60]) & (i_12_) & (i_13_) & (g102) & (g119)) + ((i_14_) & (!sk[60]) & (!i_12_) & (!i_13_) & (!g102) & (!g119)) + ((i_14_) & (!sk[60]) & (!i_12_) & (!i_13_) & (!g102) & (g119)) + ((i_14_) & (!sk[60]) & (!i_12_) & (!i_13_) & (g102) & (!g119)) + ((i_14_) & (!sk[60]) & (!i_12_) & (!i_13_) & (g102) & (g119)) + ((i_14_) & (!sk[60]) & (!i_12_) & (i_13_) & (!g102) & (!g119)) + ((i_14_) & (!sk[60]) & (!i_12_) & (i_13_) & (!g102) & (g119)) + ((i_14_) & (!sk[60]) & (!i_12_) & (i_13_) & (g102) & (!g119)) + ((i_14_) & (!sk[60]) & (!i_12_) & (i_13_) & (g102) & (g119)) + ((i_14_) & (!sk[60]) & (i_12_) & (!i_13_) & (!g102) & (!g119)) + ((i_14_) & (!sk[60]) & (i_12_) & (!i_13_) & (!g102) & (g119)) + ((i_14_) & (!sk[60]) & (i_12_) & (!i_13_) & (g102) & (!g119)) + ((i_14_) & (!sk[60]) & (i_12_) & (!i_13_) & (g102) & (g119)) + ((i_14_) & (!sk[60]) & (i_12_) & (i_13_) & (!g102) & (!g119)) + ((i_14_) & (!sk[60]) & (i_12_) & (i_13_) & (!g102) & (g119)) + ((i_14_) & (!sk[60]) & (i_12_) & (i_13_) & (g102) & (!g119)) + ((i_14_) & (!sk[60]) & (i_12_) & (i_13_) & (g102) & (g119)) + ((i_14_) & (sk[60]) & (!i_12_) & (!i_13_) & (!g102) & (!g119)) + ((i_14_) & (sk[60]) & (!i_12_) & (!i_13_) & (!g102) & (g119)) + ((i_14_) & (sk[60]) & (!i_12_) & (!i_13_) & (g102) & (g119)) + ((i_14_) & (sk[60]) & (!i_12_) & (i_13_) & (!g102) & (!g119)) + ((i_14_) & (sk[60]) & (!i_12_) & (i_13_) & (!g102) & (g119)) + ((i_14_) & (sk[60]) & (!i_12_) & (i_13_) & (g102) & (g119)) + ((i_14_) & (sk[60]) & (i_12_) & (i_13_) & (!g102) & (g119)) + ((i_14_) & (sk[60]) & (i_12_) & (i_13_) & (g102) & (g119)));
	assign g171 = (((!i_14_) & (sk[61]) & (!i_12_) & (!i_13_)) + ((!i_14_) & (sk[61]) & (!i_12_) & (i_13_)) + ((!i_14_) & (sk[61]) & (i_12_) & (!i_13_)) + ((!i_14_) & (sk[61]) & (i_12_) & (i_13_)) + ((i_14_) & (!sk[61]) & (!i_12_) & (!i_13_)) + ((i_14_) & (!sk[61]) & (!i_12_) & (i_13_)) + ((i_14_) & (!sk[61]) & (i_12_) & (!i_13_)) + ((i_14_) & (!sk[61]) & (i_12_) & (i_13_)) + ((i_14_) & (sk[61]) & (!i_12_) & (!i_13_)) + ((i_14_) & (sk[61]) & (!i_12_) & (i_13_)) + ((i_14_) & (sk[61]) & (i_12_) & (!i_13_)));
	assign g172 = (((!g15) & (sk[62]) & (!g171)) + ((g15) & (!sk[62]) & (!g171)) + ((g15) & (!sk[62]) & (g171)));
	assign g173 = (((!sk[63]) & (g102) & (!g171)) + ((!sk[63]) & (g102) & (g171)) + ((sk[63]) & (!g102) & (!g171)));
	assign g174 = (((!g20) & (!g172) & (!sk[64]) & (g142) & (g173)) + ((!g20) & (g172) & (!sk[64]) & (!g142) & (!g173)) + ((!g20) & (g172) & (!sk[64]) & (!g142) & (g173)) + ((!g20) & (g172) & (!sk[64]) & (g142) & (!g173)) + ((!g20) & (g172) & (!sk[64]) & (g142) & (g173)) + ((g20) & (!g172) & (!sk[64]) & (g142) & (!g173)) + ((g20) & (!g172) & (!sk[64]) & (g142) & (g173)) + ((g20) & (!g172) & (sk[64]) & (!g142) & (!g173)) + ((g20) & (g172) & (!sk[64]) & (!g142) & (!g173)) + ((g20) & (g172) & (!sk[64]) & (!g142) & (g173)) + ((g20) & (g172) & (!sk[64]) & (g142) & (!g173)) + ((g20) & (g172) & (!sk[64]) & (g142) & (g173)));
	assign g175 = (((!i_14_) & (!sk[65]) & (!i_12_) & (!i_13_) & (!g119) & (g131)) + ((!i_14_) & (!sk[65]) & (!i_12_) & (!i_13_) & (g119) & (g131)) + ((!i_14_) & (!sk[65]) & (!i_12_) & (i_13_) & (!g119) & (g131)) + ((!i_14_) & (!sk[65]) & (!i_12_) & (i_13_) & (g119) & (g131)) + ((!i_14_) & (!sk[65]) & (i_12_) & (!i_13_) & (!g119) & (g131)) + ((!i_14_) & (!sk[65]) & (i_12_) & (!i_13_) & (g119) & (g131)) + ((!i_14_) & (!sk[65]) & (i_12_) & (i_13_) & (!g119) & (g131)) + ((!i_14_) & (!sk[65]) & (i_12_) & (i_13_) & (g119) & (g131)) + ((i_14_) & (!sk[65]) & (!i_12_) & (!i_13_) & (!g119) & (!g131)) + ((i_14_) & (!sk[65]) & (!i_12_) & (!i_13_) & (!g119) & (g131)) + ((i_14_) & (!sk[65]) & (!i_12_) & (!i_13_) & (g119) & (!g131)) + ((i_14_) & (!sk[65]) & (!i_12_) & (!i_13_) & (g119) & (g131)) + ((i_14_) & (!sk[65]) & (!i_12_) & (i_13_) & (!g119) & (!g131)) + ((i_14_) & (!sk[65]) & (!i_12_) & (i_13_) & (!g119) & (g131)) + ((i_14_) & (!sk[65]) & (!i_12_) & (i_13_) & (g119) & (!g131)) + ((i_14_) & (!sk[65]) & (!i_12_) & (i_13_) & (g119) & (g131)) + ((i_14_) & (!sk[65]) & (i_12_) & (!i_13_) & (!g119) & (!g131)) + ((i_14_) & (!sk[65]) & (i_12_) & (!i_13_) & (!g119) & (g131)) + ((i_14_) & (!sk[65]) & (i_12_) & (!i_13_) & (g119) & (!g131)) + ((i_14_) & (!sk[65]) & (i_12_) & (!i_13_) & (g119) & (g131)) + ((i_14_) & (!sk[65]) & (i_12_) & (i_13_) & (!g119) & (!g131)) + ((i_14_) & (!sk[65]) & (i_12_) & (i_13_) & (!g119) & (g131)) + ((i_14_) & (!sk[65]) & (i_12_) & (i_13_) & (g119) & (!g131)) + ((i_14_) & (!sk[65]) & (i_12_) & (i_13_) & (g119) & (g131)) + ((i_14_) & (sk[65]) & (!i_12_) & (!i_13_) & (!g119) & (g131)) + ((i_14_) & (sk[65]) & (!i_12_) & (!i_13_) & (g119) & (!g131)) + ((i_14_) & (sk[65]) & (!i_12_) & (!i_13_) & (g119) & (g131)) + ((i_14_) & (sk[65]) & (!i_12_) & (i_13_) & (!g119) & (g131)) + ((i_14_) & (sk[65]) & (!i_12_) & (i_13_) & (g119) & (!g131)) + ((i_14_) & (sk[65]) & (!i_12_) & (i_13_) & (g119) & (g131)) + ((i_14_) & (sk[65]) & (i_12_) & (i_13_) & (!g119) & (g131)) + ((i_14_) & (sk[65]) & (i_12_) & (i_13_) & (g119) & (!g131)) + ((i_14_) & (sk[65]) & (i_12_) & (i_13_) & (g119) & (g131)));
	assign g176 = (((!i_8_) & (!g88) & (!g170) & (!g174) & (!sk[66]) & (g175)) + ((!i_8_) & (!g88) & (!g170) & (g174) & (!sk[66]) & (g175)) + ((!i_8_) & (!g88) & (g170) & (!g174) & (!sk[66]) & (g175)) + ((!i_8_) & (!g88) & (g170) & (g174) & (!sk[66]) & (g175)) + ((!i_8_) & (g88) & (!g170) & (!g174) & (!sk[66]) & (g175)) + ((!i_8_) & (g88) & (!g170) & (!g174) & (sk[66]) & (g175)) + ((!i_8_) & (g88) & (!g170) & (g174) & (!sk[66]) & (g175)) + ((!i_8_) & (g88) & (!g170) & (g174) & (sk[66]) & (g175)) + ((!i_8_) & (g88) & (g170) & (!g174) & (!sk[66]) & (g175)) + ((!i_8_) & (g88) & (g170) & (!g174) & (sk[66]) & (g175)) + ((!i_8_) & (g88) & (g170) & (g174) & (!sk[66]) & (g175)) + ((!i_8_) & (g88) & (g170) & (g174) & (sk[66]) & (g175)) + ((i_8_) & (!g88) & (!g170) & (!g174) & (!sk[66]) & (!g175)) + ((i_8_) & (!g88) & (!g170) & (!g174) & (!sk[66]) & (g175)) + ((i_8_) & (!g88) & (!g170) & (g174) & (!sk[66]) & (!g175)) + ((i_8_) & (!g88) & (!g170) & (g174) & (!sk[66]) & (g175)) + ((i_8_) & (!g88) & (g170) & (!g174) & (!sk[66]) & (!g175)) + ((i_8_) & (!g88) & (g170) & (!g174) & (!sk[66]) & (g175)) + ((i_8_) & (!g88) & (g170) & (g174) & (!sk[66]) & (!g175)) + ((i_8_) & (!g88) & (g170) & (g174) & (!sk[66]) & (g175)) + ((i_8_) & (g88) & (!g170) & (!g174) & (!sk[66]) & (!g175)) + ((i_8_) & (g88) & (!g170) & (!g174) & (!sk[66]) & (g175)) + ((i_8_) & (g88) & (!g170) & (!g174) & (sk[66]) & (!g175)) + ((i_8_) & (g88) & (!g170) & (!g174) & (sk[66]) & (g175)) + ((i_8_) & (g88) & (!g170) & (g174) & (!sk[66]) & (!g175)) + ((i_8_) & (g88) & (!g170) & (g174) & (!sk[66]) & (g175)) + ((i_8_) & (g88) & (g170) & (!g174) & (!sk[66]) & (!g175)) + ((i_8_) & (g88) & (g170) & (!g174) & (!sk[66]) & (g175)) + ((i_8_) & (g88) & (g170) & (!g174) & (sk[66]) & (!g175)) + ((i_8_) & (g88) & (g170) & (!g174) & (sk[66]) & (g175)) + ((i_8_) & (g88) & (g170) & (g174) & (!sk[66]) & (!g175)) + ((i_8_) & (g88) & (g170) & (g174) & (!sk[66]) & (g175)) + ((i_8_) & (g88) & (g170) & (g174) & (sk[66]) & (!g175)) + ((i_8_) & (g88) & (g170) & (g174) & (sk[66]) & (g175)));
	assign g177 = (((g11) & (!sk[67]) & (!g171)) + ((g11) & (!sk[67]) & (g171)) + ((g11) & (sk[67]) & (!g171)));
	assign g178 = (((!sk[68]) & (i_11_) & (!i_9_) & (!i_10_)) + ((!sk[68]) & (i_11_) & (!i_9_) & (i_10_)) + ((!sk[68]) & (i_11_) & (i_9_) & (!i_10_)) + ((!sk[68]) & (i_11_) & (i_9_) & (i_10_)) + ((sk[68]) & (!i_11_) & (i_9_) & (!i_10_)) + ((sk[68]) & (i_11_) & (!i_9_) & (!i_10_)));
	assign g179 = (((!sk[69]) & (i_15_) & (!g171) & (!g178)) + ((!sk[69]) & (i_15_) & (!g171) & (g178)) + ((!sk[69]) & (i_15_) & (g171) & (!g178)) + ((!sk[69]) & (i_15_) & (g171) & (g178)) + ((sk[69]) & (!i_15_) & (!g171) & (g178)));
	assign g180 = (((!i_14_) & (!sk[70]) & (!i_12_) & (!i_13_) & (!g59) & (g95)) + ((!i_14_) & (!sk[70]) & (!i_12_) & (!i_13_) & (g59) & (g95)) + ((!i_14_) & (!sk[70]) & (!i_12_) & (i_13_) & (!g59) & (g95)) + ((!i_14_) & (!sk[70]) & (!i_12_) & (i_13_) & (g59) & (g95)) + ((!i_14_) & (!sk[70]) & (i_12_) & (!i_13_) & (!g59) & (g95)) + ((!i_14_) & (!sk[70]) & (i_12_) & (!i_13_) & (g59) & (g95)) + ((!i_14_) & (!sk[70]) & (i_12_) & (i_13_) & (!g59) & (g95)) + ((!i_14_) & (!sk[70]) & (i_12_) & (i_13_) & (g59) & (g95)) + ((i_14_) & (!sk[70]) & (!i_12_) & (!i_13_) & (!g59) & (!g95)) + ((i_14_) & (!sk[70]) & (!i_12_) & (!i_13_) & (!g59) & (g95)) + ((i_14_) & (!sk[70]) & (!i_12_) & (!i_13_) & (g59) & (!g95)) + ((i_14_) & (!sk[70]) & (!i_12_) & (!i_13_) & (g59) & (g95)) + ((i_14_) & (!sk[70]) & (!i_12_) & (i_13_) & (!g59) & (!g95)) + ((i_14_) & (!sk[70]) & (!i_12_) & (i_13_) & (!g59) & (g95)) + ((i_14_) & (!sk[70]) & (!i_12_) & (i_13_) & (g59) & (!g95)) + ((i_14_) & (!sk[70]) & (!i_12_) & (i_13_) & (g59) & (g95)) + ((i_14_) & (!sk[70]) & (i_12_) & (!i_13_) & (!g59) & (!g95)) + ((i_14_) & (!sk[70]) & (i_12_) & (!i_13_) & (!g59) & (g95)) + ((i_14_) & (!sk[70]) & (i_12_) & (!i_13_) & (g59) & (!g95)) + ((i_14_) & (!sk[70]) & (i_12_) & (!i_13_) & (g59) & (g95)) + ((i_14_) & (!sk[70]) & (i_12_) & (i_13_) & (!g59) & (!g95)) + ((i_14_) & (!sk[70]) & (i_12_) & (i_13_) & (!g59) & (g95)) + ((i_14_) & (!sk[70]) & (i_12_) & (i_13_) & (g59) & (!g95)) + ((i_14_) & (!sk[70]) & (i_12_) & (i_13_) & (g59) & (g95)) + ((i_14_) & (sk[70]) & (!i_12_) & (!i_13_) & (g59) & (g95)) + ((i_14_) & (sk[70]) & (!i_12_) & (i_13_) & (g59) & (g95)) + ((i_14_) & (sk[70]) & (i_12_) & (i_13_) & (g59) & (g95)));
	assign g181 = (((!g91) & (sk[71]) & (g119)) + ((g91) & (!sk[71]) & (!g119)) + ((g91) & (!sk[71]) & (g119)));
	assign g182 = (((!sk[72]) & (i_14_) & (!i_12_) & (!i_13_)) + ((!sk[72]) & (i_14_) & (!i_12_) & (i_13_)) + ((!sk[72]) & (i_14_) & (i_12_) & (!i_13_)) + ((!sk[72]) & (i_14_) & (i_12_) & (i_13_)) + ((sk[72]) & (i_14_) & (i_12_) & (!i_13_)));
	assign g183 = (((g119) & (!sk[73]) & (!g182)) + ((g119) & (!sk[73]) & (g182)) + ((g119) & (sk[73]) & (g182)));
	assign g184 = (((!g181) & (!g118) & (g112) & (!sk[74]) & (g183)) + ((!g181) & (g118) & (!g112) & (!sk[74]) & (!g183)) + ((!g181) & (g118) & (!g112) & (!sk[74]) & (g183)) + ((!g181) & (g118) & (!g112) & (sk[74]) & (g183)) + ((!g181) & (g118) & (g112) & (!sk[74]) & (!g183)) + ((!g181) & (g118) & (g112) & (!sk[74]) & (g183)) + ((!g181) & (g118) & (g112) & (sk[74]) & (g183)) + ((g181) & (!g118) & (g112) & (!sk[74]) & (!g183)) + ((g181) & (!g118) & (g112) & (!sk[74]) & (g183)) + ((g181) & (!g118) & (g112) & (sk[74]) & (!g183)) + ((g181) & (!g118) & (g112) & (sk[74]) & (g183)) + ((g181) & (g118) & (!g112) & (!sk[74]) & (!g183)) + ((g181) & (g118) & (!g112) & (!sk[74]) & (g183)) + ((g181) & (g118) & (!g112) & (sk[74]) & (g183)) + ((g181) & (g118) & (g112) & (!sk[74]) & (!g183)) + ((g181) & (g118) & (g112) & (!sk[74]) & (g183)) + ((g181) & (g118) & (g112) & (sk[74]) & (!g183)) + ((g181) & (g118) & (g112) & (sk[74]) & (g183)));
	assign g185 = (((!sk[75]) & (g104) & (!g91)) + ((!sk[75]) & (g104) & (g91)) + ((sk[75]) & (!g104) & (!g91)) + ((sk[75]) & (!g104) & (g91)) + ((sk[75]) & (g104) & (g91)));
	assign g186 = (((!g31) & (sk[76]) & (g34) & (g87)) + ((g31) & (!sk[76]) & (!g34) & (!g87)) + ((g31) & (!sk[76]) & (!g34) & (g87)) + ((g31) & (!sk[76]) & (g34) & (!g87)) + ((g31) & (!sk[76]) & (g34) & (g87)) + ((g31) & (sk[76]) & (!g34) & (g87)) + ((g31) & (sk[76]) & (g34) & (g87)));
	assign g187 = (((g104) & (!sk[77]) & (!g182)) + ((g104) & (!sk[77]) & (g182)) + ((g104) & (sk[77]) & (g182)));
	assign g188 = (((!g134) & (!g118) & (!g185) & (!sk[78]) & (!g186) & (g187)) + ((!g134) & (!g118) & (!g185) & (!sk[78]) & (g186) & (g187)) + ((!g134) & (!g118) & (!g185) & (sk[78]) & (!g186) & (!g187)) + ((!g134) & (!g118) & (!g185) & (sk[78]) & (!g186) & (g187)) + ((!g134) & (!g118) & (!g185) & (sk[78]) & (g186) & (!g187)) + ((!g134) & (!g118) & (g185) & (!sk[78]) & (!g186) & (g187)) + ((!g134) & (!g118) & (g185) & (!sk[78]) & (g186) & (g187)) + ((!g134) & (!g118) & (g185) & (sk[78]) & (!g186) & (!g187)) + ((!g134) & (!g118) & (g185) & (sk[78]) & (!g186) & (g187)) + ((!g134) & (!g118) & (g185) & (sk[78]) & (g186) & (!g187)) + ((!g134) & (g118) & (!g185) & (!sk[78]) & (!g186) & (g187)) + ((!g134) & (g118) & (!g185) & (!sk[78]) & (g186) & (g187)) + ((!g134) & (g118) & (!g185) & (sk[78]) & (!g186) & (!g187)) + ((!g134) & (g118) & (!g185) & (sk[78]) & (g186) & (!g187)) + ((!g134) & (g118) & (g185) & (!sk[78]) & (!g186) & (g187)) + ((!g134) & (g118) & (g185) & (!sk[78]) & (g186) & (g187)) + ((!g134) & (g118) & (g185) & (sk[78]) & (!g186) & (!g187)) + ((!g134) & (g118) & (g185) & (sk[78]) & (g186) & (!g187)) + ((g134) & (!g118) & (!g185) & (!sk[78]) & (!g186) & (!g187)) + ((g134) & (!g118) & (!g185) & (!sk[78]) & (!g186) & (g187)) + ((g134) & (!g118) & (!g185) & (!sk[78]) & (g186) & (!g187)) + ((g134) & (!g118) & (!g185) & (!sk[78]) & (g186) & (g187)) + ((g134) & (!g118) & (g185) & (!sk[78]) & (!g186) & (!g187)) + ((g134) & (!g118) & (g185) & (!sk[78]) & (!g186) & (g187)) + ((g134) & (!g118) & (g185) & (!sk[78]) & (g186) & (!g187)) + ((g134) & (!g118) & (g185) & (!sk[78]) & (g186) & (g187)) + ((g134) & (!g118) & (g185) & (sk[78]) & (!g186) & (!g187)) + ((g134) & (!g118) & (g185) & (sk[78]) & (!g186) & (g187)) + ((g134) & (!g118) & (g185) & (sk[78]) & (g186) & (!g187)) + ((g134) & (g118) & (!g185) & (!sk[78]) & (!g186) & (!g187)) + ((g134) & (g118) & (!g185) & (!sk[78]) & (!g186) & (g187)) + ((g134) & (g118) & (!g185) & (!sk[78]) & (g186) & (!g187)) + ((g134) & (g118) & (!g185) & (!sk[78]) & (g186) & (g187)) + ((g134) & (g118) & (g185) & (!sk[78]) & (!g186) & (!g187)) + ((g134) & (g118) & (g185) & (!sk[78]) & (!g186) & (g187)) + ((g134) & (g118) & (g185) & (!sk[78]) & (g186) & (!g187)) + ((g134) & (g118) & (g185) & (!sk[78]) & (g186) & (g187)) + ((g134) & (g118) & (g185) & (sk[78]) & (!g186) & (!g187)) + ((g134) & (g118) & (g185) & (sk[78]) & (g186) & (!g187)));
	assign g189 = (((!g151) & (!g177) & (!g179) & (!g180) & (!g184) & (g188)) + ((!g151) & (!g177) & (g179) & (!g180) & (!g184) & (g188)) + ((!g151) & (g177) & (!g179) & (!g180) & (!g184) & (g188)) + ((!g151) & (g177) & (g179) & (!g180) & (!g184) & (g188)) + ((g151) & (!g177) & (!g179) & (!g180) & (!g184) & (g188)));
	assign g190 = (((!sk[80]) & (i_14_) & (!g99) & (!g131)) + ((!sk[80]) & (i_14_) & (!g99) & (g131)) + ((!sk[80]) & (i_14_) & (g99) & (!g131)) + ((!sk[80]) & (i_14_) & (g99) & (g131)) + ((sk[80]) & (i_14_) & (g99) & (g131)));
	assign g191 = (((!sk[81]) & (g15) & (!g182)) + ((!sk[81]) & (g15) & (g182)) + ((sk[81]) & (!g15) & (g182)));
	assign g192 = (((!i_8_) & (!i_6_) & (i_7_) & (!g58) & (g98) & (g191)) + ((!i_8_) & (!i_6_) & (i_7_) & (g58) & (g98) & (g191)) + ((!i_8_) & (i_6_) & (!i_7_) & (!g58) & (g98) & (g191)) + ((!i_8_) & (i_6_) & (!i_7_) & (g58) & (g98) & (g191)) + ((!i_8_) & (i_6_) & (i_7_) & (!g58) & (g98) & (g191)) + ((!i_8_) & (i_6_) & (i_7_) & (g58) & (!g98) & (g191)) + ((!i_8_) & (i_6_) & (i_7_) & (g58) & (g98) & (g191)) + ((i_8_) & (!i_6_) & (i_7_) & (!g58) & (g98) & (g191)) + ((i_8_) & (!i_6_) & (i_7_) & (g58) & (g98) & (g191)));
	assign g193 = (((!sk[83]) & (g102) & (!g182)) + ((!sk[83]) & (g102) & (g182)) + ((sk[83]) & (!g102) & (g182)));
	assign g194 = (((!i_8_) & (!g108) & (!sk[84]) & (g183) & (g193)) + ((!i_8_) & (g108) & (!sk[84]) & (!g183) & (!g193)) + ((!i_8_) & (g108) & (!sk[84]) & (!g183) & (g193)) + ((!i_8_) & (g108) & (!sk[84]) & (g183) & (!g193)) + ((!i_8_) & (g108) & (!sk[84]) & (g183) & (g193)) + ((!i_8_) & (g108) & (sk[84]) & (!g183) & (g193)) + ((!i_8_) & (g108) & (sk[84]) & (g183) & (g193)) + ((i_8_) & (!g108) & (!sk[84]) & (g183) & (!g193)) + ((i_8_) & (!g108) & (!sk[84]) & (g183) & (g193)) + ((i_8_) & (g108) & (!sk[84]) & (!g183) & (!g193)) + ((i_8_) & (g108) & (!sk[84]) & (!g183) & (g193)) + ((i_8_) & (g108) & (!sk[84]) & (g183) & (!g193)) + ((i_8_) & (g108) & (!sk[84]) & (g183) & (g193)) + ((i_8_) & (g108) & (sk[84]) & (!g183) & (g193)) + ((i_8_) & (g108) & (sk[84]) & (g183) & (!g193)) + ((i_8_) & (g108) & (sk[84]) & (g183) & (g193)));
	assign g195 = (((!sk[85]) & (g104) & (!g171)) + ((!sk[85]) & (g104) & (g171)) + ((sk[85]) & (g104) & (!g171)));
	assign g196 = (((!i_8_) & (!g108) & (!sk[86]) & (!g185) & (!g195) & (g187)) + ((!i_8_) & (!g108) & (!sk[86]) & (!g185) & (g195) & (g187)) + ((!i_8_) & (!g108) & (!sk[86]) & (g185) & (!g195) & (g187)) + ((!i_8_) & (!g108) & (!sk[86]) & (g185) & (g195) & (g187)) + ((!i_8_) & (g108) & (!sk[86]) & (!g185) & (!g195) & (g187)) + ((!i_8_) & (g108) & (!sk[86]) & (!g185) & (g195) & (g187)) + ((!i_8_) & (g108) & (!sk[86]) & (g185) & (!g195) & (g187)) + ((!i_8_) & (g108) & (!sk[86]) & (g185) & (g195) & (g187)) + ((!i_8_) & (g108) & (sk[86]) & (!g185) & (!g195) & (!g187)) + ((!i_8_) & (g108) & (sk[86]) & (!g185) & (!g195) & (g187)) + ((!i_8_) & (g108) & (sk[86]) & (!g185) & (g195) & (!g187)) + ((!i_8_) & (g108) & (sk[86]) & (!g185) & (g195) & (g187)) + ((!i_8_) & (g108) & (sk[86]) & (g185) & (!g195) & (g187)) + ((!i_8_) & (g108) & (sk[86]) & (g185) & (g195) & (!g187)) + ((!i_8_) & (g108) & (sk[86]) & (g185) & (g195) & (g187)) + ((i_8_) & (!g108) & (!sk[86]) & (!g185) & (!g195) & (!g187)) + ((i_8_) & (!g108) & (!sk[86]) & (!g185) & (!g195) & (g187)) + ((i_8_) & (!g108) & (!sk[86]) & (!g185) & (g195) & (!g187)) + ((i_8_) & (!g108) & (!sk[86]) & (!g185) & (g195) & (g187)) + ((i_8_) & (!g108) & (!sk[86]) & (g185) & (!g195) & (!g187)) + ((i_8_) & (!g108) & (!sk[86]) & (g185) & (!g195) & (g187)) + ((i_8_) & (!g108) & (!sk[86]) & (g185) & (g195) & (!g187)) + ((i_8_) & (!g108) & (!sk[86]) & (g185) & (g195) & (g187)) + ((i_8_) & (g108) & (!sk[86]) & (!g185) & (!g195) & (!g187)) + ((i_8_) & (g108) & (!sk[86]) & (!g185) & (!g195) & (g187)) + ((i_8_) & (g108) & (!sk[86]) & (!g185) & (g195) & (!g187)) + ((i_8_) & (g108) & (!sk[86]) & (!g185) & (g195) & (g187)) + ((i_8_) & (g108) & (!sk[86]) & (g185) & (!g195) & (!g187)) + ((i_8_) & (g108) & (!sk[86]) & (g185) & (!g195) & (g187)) + ((i_8_) & (g108) & (!sk[86]) & (g185) & (g195) & (!g187)) + ((i_8_) & (g108) & (!sk[86]) & (g185) & (g195) & (g187)) + ((i_8_) & (g108) & (sk[86]) & (!g185) & (g195) & (!g187)) + ((i_8_) & (g108) & (sk[86]) & (!g185) & (g195) & (g187)) + ((i_8_) & (g108) & (sk[86]) & (g185) & (g195) & (!g187)) + ((i_8_) & (g108) & (sk[86]) & (g185) & (g195) & (g187)));
	assign g197 = (((g6) & (!sk[87]) & (!i_15_) & (!g171)) + ((g6) & (!sk[87]) & (!i_15_) & (g171)) + ((g6) & (!sk[87]) & (i_15_) & (!g171)) + ((g6) & (!sk[87]) & (i_15_) & (g171)) + ((g6) & (sk[87]) & (!i_15_) & (!g171)));
	assign g198 = (((!sk[88]) & (!i_8_) & (!g108) & (g197) & (g177)) + ((!sk[88]) & (!i_8_) & (g108) & (!g197) & (!g177)) + ((!sk[88]) & (!i_8_) & (g108) & (!g197) & (g177)) + ((!sk[88]) & (!i_8_) & (g108) & (g197) & (!g177)) + ((!sk[88]) & (!i_8_) & (g108) & (g197) & (g177)) + ((!sk[88]) & (i_8_) & (!g108) & (g197) & (!g177)) + ((!sk[88]) & (i_8_) & (!g108) & (g197) & (g177)) + ((!sk[88]) & (i_8_) & (g108) & (!g197) & (!g177)) + ((!sk[88]) & (i_8_) & (g108) & (!g197) & (g177)) + ((!sk[88]) & (i_8_) & (g108) & (g197) & (!g177)) + ((!sk[88]) & (i_8_) & (g108) & (g197) & (g177)) + ((sk[88]) & (!i_8_) & (g108) & (!g197) & (g177)) + ((sk[88]) & (!i_8_) & (g108) & (g197) & (g177)) + ((sk[88]) & (i_8_) & (g108) & (!g197) & (g177)) + ((sk[88]) & (i_8_) & (g108) & (g197) & (!g177)) + ((sk[88]) & (i_8_) & (g108) & (g197) & (g177)));
	assign g199 = (((g119) & (!sk[89]) & (!g171)) + ((g119) & (!sk[89]) & (g171)) + ((g119) & (sk[89]) & (!g171)));
	assign g200 = (((!i_8_) & (!sk[90]) & (!g181) & (g135) & (g199)) + ((!i_8_) & (!sk[90]) & (g181) & (!g135) & (!g199)) + ((!i_8_) & (!sk[90]) & (g181) & (!g135) & (g199)) + ((!i_8_) & (!sk[90]) & (g181) & (g135) & (!g199)) + ((!i_8_) & (!sk[90]) & (g181) & (g135) & (g199)) + ((i_8_) & (!sk[90]) & (!g181) & (g135) & (!g199)) + ((i_8_) & (!sk[90]) & (!g181) & (g135) & (g199)) + ((i_8_) & (!sk[90]) & (g181) & (!g135) & (!g199)) + ((i_8_) & (!sk[90]) & (g181) & (!g135) & (g199)) + ((i_8_) & (!sk[90]) & (g181) & (g135) & (!g199)) + ((i_8_) & (!sk[90]) & (g181) & (g135) & (g199)) + ((i_8_) & (sk[90]) & (!g181) & (g135) & (g199)) + ((i_8_) & (sk[90]) & (g181) & (g135) & (!g199)) + ((i_8_) & (sk[90]) & (g181) & (g135) & (g199)));
	assign g201 = (((!sk[91]) & (g11) & (!g182)) + ((!sk[91]) & (g11) & (g182)) + ((sk[91]) & (!g11) & (!g182)) + ((sk[91]) & (!g11) & (g182)) + ((sk[91]) & (g11) & (!g182)));
	assign g202 = (((!i_8_) & (!i_6_) & (!i_7_) & (!g98) & (!sk[92]) & (g201)) + ((!i_8_) & (!i_6_) & (!i_7_) & (g98) & (!sk[92]) & (g201)) + ((!i_8_) & (!i_6_) & (i_7_) & (!g98) & (!sk[92]) & (g201)) + ((!i_8_) & (!i_6_) & (i_7_) & (g98) & (!sk[92]) & (g201)) + ((!i_8_) & (i_6_) & (!i_7_) & (!g98) & (!sk[92]) & (g201)) + ((!i_8_) & (i_6_) & (!i_7_) & (g98) & (!sk[92]) & (g201)) + ((!i_8_) & (i_6_) & (!i_7_) & (g98) & (sk[92]) & (!g201)) + ((!i_8_) & (i_6_) & (i_7_) & (!g98) & (!sk[92]) & (g201)) + ((!i_8_) & (i_6_) & (i_7_) & (g98) & (!sk[92]) & (g201)) + ((!i_8_) & (i_6_) & (i_7_) & (g98) & (sk[92]) & (!g201)) + ((i_8_) & (!i_6_) & (!i_7_) & (!g98) & (!sk[92]) & (!g201)) + ((i_8_) & (!i_6_) & (!i_7_) & (!g98) & (!sk[92]) & (g201)) + ((i_8_) & (!i_6_) & (!i_7_) & (g98) & (!sk[92]) & (!g201)) + ((i_8_) & (!i_6_) & (!i_7_) & (g98) & (!sk[92]) & (g201)) + ((i_8_) & (!i_6_) & (i_7_) & (!g98) & (!sk[92]) & (!g201)) + ((i_8_) & (!i_6_) & (i_7_) & (!g98) & (!sk[92]) & (g201)) + ((i_8_) & (!i_6_) & (i_7_) & (g98) & (!sk[92]) & (!g201)) + ((i_8_) & (!i_6_) & (i_7_) & (g98) & (!sk[92]) & (g201)) + ((i_8_) & (!i_6_) & (i_7_) & (g98) & (sk[92]) & (!g201)) + ((i_8_) & (i_6_) & (!i_7_) & (!g98) & (!sk[92]) & (!g201)) + ((i_8_) & (i_6_) & (!i_7_) & (!g98) & (!sk[92]) & (g201)) + ((i_8_) & (i_6_) & (!i_7_) & (g98) & (!sk[92]) & (!g201)) + ((i_8_) & (i_6_) & (!i_7_) & (g98) & (!sk[92]) & (g201)) + ((i_8_) & (i_6_) & (i_7_) & (!g98) & (!sk[92]) & (!g201)) + ((i_8_) & (i_6_) & (i_7_) & (!g98) & (!sk[92]) & (g201)) + ((i_8_) & (i_6_) & (i_7_) & (g98) & (!sk[92]) & (!g201)) + ((i_8_) & (i_6_) & (i_7_) & (g98) & (!sk[92]) & (g201)));
	assign g203 = (((g182) & (!sk[93]) & (!g93)) + ((g182) & (!sk[93]) & (g93)) + ((g182) & (sk[93]) & (!g93)));
	assign g204 = (((!g182) & (sk[94]) & (!g158)) + ((!g182) & (sk[94]) & (g158)) + ((g182) & (!sk[94]) & (!g158)) + ((g182) & (!sk[94]) & (g158)) + ((g182) & (sk[94]) & (!g158)));
	assign g205 = (((!i_8_) & (!g100) & (!sk[95]) & (g203) & (g204)) + ((!i_8_) & (g100) & (!sk[95]) & (!g203) & (!g204)) + ((!i_8_) & (g100) & (!sk[95]) & (!g203) & (g204)) + ((!i_8_) & (g100) & (!sk[95]) & (g203) & (!g204)) + ((!i_8_) & (g100) & (!sk[95]) & (g203) & (g204)) + ((i_8_) & (!g100) & (!sk[95]) & (g203) & (!g204)) + ((i_8_) & (!g100) & (!sk[95]) & (g203) & (g204)) + ((i_8_) & (g100) & (!sk[95]) & (!g203) & (!g204)) + ((i_8_) & (g100) & (!sk[95]) & (!g203) & (g204)) + ((i_8_) & (g100) & (!sk[95]) & (g203) & (!g204)) + ((i_8_) & (g100) & (!sk[95]) & (g203) & (g204)) + ((i_8_) & (g100) & (sk[95]) & (!g203) & (!g204)) + ((i_8_) & (g100) & (sk[95]) & (g203) & (!g204)) + ((i_8_) & (g100) & (sk[95]) & (g203) & (g204)));
	assign g206 = (((!sk[96]) & (g11) & (!g91)) + ((!sk[96]) & (g11) & (g91)) + ((sk[96]) & (!g11) & (!g91)) + ((sk[96]) & (!g11) & (g91)) + ((sk[96]) & (g11) & (g91)));
	assign g207 = (((!sk[97]) & (g91) & (!g131)) + ((!sk[97]) & (g91) & (g131)) + ((sk[97]) & (!g91) & (g131)));
	assign g208 = (((!i_8_) & (!g4) & (!sk[98]) & (!g206) & (!g98) & (g207)) + ((!i_8_) & (!g4) & (!sk[98]) & (!g206) & (g98) & (g207)) + ((!i_8_) & (!g4) & (!sk[98]) & (g206) & (!g98) & (g207)) + ((!i_8_) & (!g4) & (!sk[98]) & (g206) & (g98) & (g207)) + ((!i_8_) & (g4) & (!sk[98]) & (!g206) & (!g98) & (g207)) + ((!i_8_) & (g4) & (!sk[98]) & (!g206) & (g98) & (g207)) + ((!i_8_) & (g4) & (!sk[98]) & (g206) & (!g98) & (g207)) + ((!i_8_) & (g4) & (!sk[98]) & (g206) & (g98) & (g207)) + ((!i_8_) & (g4) & (sk[98]) & (!g206) & (g98) & (!g207)) + ((!i_8_) & (g4) & (sk[98]) & (!g206) & (g98) & (g207)) + ((i_8_) & (!g4) & (!sk[98]) & (!g206) & (!g98) & (!g207)) + ((i_8_) & (!g4) & (!sk[98]) & (!g206) & (!g98) & (g207)) + ((i_8_) & (!g4) & (!sk[98]) & (!g206) & (g98) & (!g207)) + ((i_8_) & (!g4) & (!sk[98]) & (!g206) & (g98) & (g207)) + ((i_8_) & (!g4) & (!sk[98]) & (g206) & (!g98) & (!g207)) + ((i_8_) & (!g4) & (!sk[98]) & (g206) & (!g98) & (g207)) + ((i_8_) & (!g4) & (!sk[98]) & (g206) & (g98) & (!g207)) + ((i_8_) & (!g4) & (!sk[98]) & (g206) & (g98) & (g207)) + ((i_8_) & (g4) & (!sk[98]) & (!g206) & (!g98) & (!g207)) + ((i_8_) & (g4) & (!sk[98]) & (!g206) & (!g98) & (g207)) + ((i_8_) & (g4) & (!sk[98]) & (!g206) & (g98) & (!g207)) + ((i_8_) & (g4) & (!sk[98]) & (!g206) & (g98) & (g207)) + ((i_8_) & (g4) & (!sk[98]) & (g206) & (!g98) & (!g207)) + ((i_8_) & (g4) & (!sk[98]) & (g206) & (!g98) & (g207)) + ((i_8_) & (g4) & (!sk[98]) & (g206) & (g98) & (!g207)) + ((i_8_) & (g4) & (!sk[98]) & (g206) & (g98) & (g207)) + ((i_8_) & (g4) & (sk[98]) & (!g206) & (g98) & (!g207)) + ((i_8_) & (g4) & (sk[98]) & (!g206) & (g98) & (g207)) + ((i_8_) & (g4) & (sk[98]) & (g206) & (g98) & (g207)));
	assign g209 = (((g6) & (!i_15_) & (!sk[99]) & (!g182)) + ((g6) & (!i_15_) & (!sk[99]) & (g182)) + ((g6) & (!i_15_) & (sk[99]) & (g182)) + ((g6) & (i_15_) & (!sk[99]) & (!g182)) + ((g6) & (i_15_) & (!sk[99]) & (g182)));
	assign g210 = (((!i_8_) & (!g100) & (!sk[100]) & (g183) & (g209)) + ((!i_8_) & (g100) & (!sk[100]) & (!g183) & (!g209)) + ((!i_8_) & (g100) & (!sk[100]) & (!g183) & (g209)) + ((!i_8_) & (g100) & (!sk[100]) & (g183) & (!g209)) + ((!i_8_) & (g100) & (!sk[100]) & (g183) & (g209)) + ((i_8_) & (!g100) & (!sk[100]) & (g183) & (!g209)) + ((i_8_) & (!g100) & (!sk[100]) & (g183) & (g209)) + ((i_8_) & (g100) & (!sk[100]) & (!g183) & (!g209)) + ((i_8_) & (g100) & (!sk[100]) & (!g183) & (g209)) + ((i_8_) & (g100) & (!sk[100]) & (g183) & (!g209)) + ((i_8_) & (g100) & (!sk[100]) & (g183) & (g209)) + ((i_8_) & (g100) & (sk[100]) & (!g183) & (g209)) + ((i_8_) & (g100) & (sk[100]) & (g183) & (!g209)) + ((i_8_) & (g100) & (sk[100]) & (g183) & (g209)));
	assign g211 = (((!g198) & (!g200) & (!g202) & (!g205) & (!g208) & (!g210)));
	assign g212 = (((!i_8_) & (!sk[102]) & (!g59) & (!g108) & (!g112) & (g135)) + ((!i_8_) & (!sk[102]) & (!g59) & (!g108) & (g112) & (g135)) + ((!i_8_) & (!sk[102]) & (!g59) & (g108) & (!g112) & (g135)) + ((!i_8_) & (!sk[102]) & (!g59) & (g108) & (g112) & (g135)) + ((!i_8_) & (!sk[102]) & (g59) & (!g108) & (!g112) & (g135)) + ((!i_8_) & (!sk[102]) & (g59) & (!g108) & (g112) & (g135)) + ((!i_8_) & (!sk[102]) & (g59) & (g108) & (!g112) & (g135)) + ((!i_8_) & (!sk[102]) & (g59) & (g108) & (g112) & (g135)) + ((!i_8_) & (sk[102]) & (!g59) & (!g108) & (!g112) & (!g135)) + ((i_8_) & (!sk[102]) & (!g59) & (!g108) & (!g112) & (!g135)) + ((i_8_) & (!sk[102]) & (!g59) & (!g108) & (!g112) & (g135)) + ((i_8_) & (!sk[102]) & (!g59) & (!g108) & (g112) & (!g135)) + ((i_8_) & (!sk[102]) & (!g59) & (!g108) & (g112) & (g135)) + ((i_8_) & (!sk[102]) & (!g59) & (g108) & (!g112) & (!g135)) + ((i_8_) & (!sk[102]) & (!g59) & (g108) & (!g112) & (g135)) + ((i_8_) & (!sk[102]) & (!g59) & (g108) & (g112) & (!g135)) + ((i_8_) & (!sk[102]) & (!g59) & (g108) & (g112) & (g135)) + ((i_8_) & (!sk[102]) & (g59) & (!g108) & (!g112) & (!g135)) + ((i_8_) & (!sk[102]) & (g59) & (!g108) & (!g112) & (g135)) + ((i_8_) & (!sk[102]) & (g59) & (!g108) & (g112) & (!g135)) + ((i_8_) & (!sk[102]) & (g59) & (!g108) & (g112) & (g135)) + ((i_8_) & (!sk[102]) & (g59) & (g108) & (!g112) & (!g135)) + ((i_8_) & (!sk[102]) & (g59) & (g108) & (!g112) & (g135)) + ((i_8_) & (!sk[102]) & (g59) & (g108) & (g112) & (!g135)) + ((i_8_) & (!sk[102]) & (g59) & (g108) & (g112) & (g135)) + ((i_8_) & (sk[102]) & (!g59) & (!g108) & (!g112) & (!g135)) + ((i_8_) & (sk[102]) & (!g59) & (g108) & (!g112) & (!g135)));
	assign g213 = (((g95) & (!sk[103]) & (!g182)) + ((g95) & (!sk[103]) & (g182)) + ((g95) & (sk[103]) & (g182)));
	assign g214 = (((!sk[104]) & (i_8_) & (!i_6_) & (!g87)) + ((!sk[104]) & (i_8_) & (!i_6_) & (g87)) + ((!sk[104]) & (i_8_) & (i_6_) & (!g87)) + ((!sk[104]) & (i_8_) & (i_6_) & (g87)) + ((sk[104]) & (!i_8_) & (!i_6_) & (g87)));
	assign g215 = (((!g118) & (sk[105]) & (!g214)) + ((g118) & (!sk[105]) & (!g214)) + ((g118) & (!sk[105]) & (g214)));
	assign g216 = (((g13) & (!sk[106]) & (!g119)) + ((g13) & (!sk[106]) & (g119)) + ((g13) & (sk[106]) & (g119)));
	assign g217 = (((!g112) & (!g216) & (!sk[107]) & (g199) & (g120)) + ((!g112) & (g216) & (!sk[107]) & (!g199) & (!g120)) + ((!g112) & (g216) & (!sk[107]) & (!g199) & (g120)) + ((!g112) & (g216) & (!sk[107]) & (g199) & (!g120)) + ((!g112) & (g216) & (!sk[107]) & (g199) & (g120)) + ((g112) & (!g216) & (!sk[107]) & (g199) & (!g120)) + ((g112) & (!g216) & (!sk[107]) & (g199) & (g120)) + ((g112) & (!g216) & (sk[107]) & (!g199) & (!g120)) + ((g112) & (!g216) & (sk[107]) & (g199) & (!g120)) + ((g112) & (!g216) & (sk[107]) & (g199) & (g120)) + ((g112) & (g216) & (!sk[107]) & (!g199) & (!g120)) + ((g112) & (g216) & (!sk[107]) & (!g199) & (g120)) + ((g112) & (g216) & (!sk[107]) & (g199) & (!g120)) + ((g112) & (g216) & (!sk[107]) & (g199) & (g120)) + ((g112) & (g216) & (sk[107]) & (!g199) & (!g120)) + ((g112) & (g216) & (sk[107]) & (!g199) & (g120)) + ((g112) & (g216) & (sk[107]) & (g199) & (!g120)) + ((g112) & (g216) & (sk[107]) & (g199) & (g120)));
	assign g218 = (((!sk[108]) & (!g212) & (!g213) & (g215) & (g217)) + ((!sk[108]) & (!g212) & (g213) & (!g215) & (!g217)) + ((!sk[108]) & (!g212) & (g213) & (!g215) & (g217)) + ((!sk[108]) & (!g212) & (g213) & (g215) & (!g217)) + ((!sk[108]) & (!g212) & (g213) & (g215) & (g217)) + ((!sk[108]) & (g212) & (!g213) & (g215) & (!g217)) + ((!sk[108]) & (g212) & (!g213) & (g215) & (g217)) + ((!sk[108]) & (g212) & (g213) & (!g215) & (!g217)) + ((!sk[108]) & (g212) & (g213) & (!g215) & (g217)) + ((!sk[108]) & (g212) & (g213) & (g215) & (!g217)) + ((!sk[108]) & (g212) & (g213) & (g215) & (g217)) + ((sk[108]) & (!g212) & (!g213) & (!g215) & (!g217)) + ((sk[108]) & (!g212) & (!g213) & (g215) & (!g217)) + ((sk[108]) & (g212) & (!g213) & (!g215) & (!g217)) + ((sk[108]) & (g212) & (!g213) & (g215) & (!g217)) + ((sk[108]) & (g212) & (g213) & (g215) & (!g217)));
	assign g219 = (((!sk[109]) & (!g134) & (!g183) & (g187) & (g193)) + ((!sk[109]) & (!g134) & (g183) & (!g187) & (!g193)) + ((!sk[109]) & (!g134) & (g183) & (!g187) & (g193)) + ((!sk[109]) & (!g134) & (g183) & (g187) & (!g193)) + ((!sk[109]) & (!g134) & (g183) & (g187) & (g193)) + ((!sk[109]) & (g134) & (!g183) & (g187) & (!g193)) + ((!sk[109]) & (g134) & (!g183) & (g187) & (g193)) + ((!sk[109]) & (g134) & (g183) & (!g187) & (!g193)) + ((!sk[109]) & (g134) & (g183) & (!g187) & (g193)) + ((!sk[109]) & (g134) & (g183) & (g187) & (!g193)) + ((!sk[109]) & (g134) & (g183) & (g187) & (g193)) + ((sk[109]) & (g134) & (!g183) & (!g187) & (g193)) + ((sk[109]) & (g134) & (!g183) & (g187) & (!g193)) + ((sk[109]) & (g134) & (!g183) & (g187) & (g193)) + ((sk[109]) & (g134) & (g183) & (!g187) & (!g193)) + ((sk[109]) & (g134) & (g183) & (!g187) & (g193)) + ((sk[109]) & (g134) & (g183) & (g187) & (!g193)) + ((sk[109]) & (g134) & (g183) & (g187) & (g193)));
	assign g220 = (((!g91) & (sk[110]) & (!g102)) + ((g91) & (!sk[110]) & (!g102)) + ((g91) & (!sk[110]) & (g102)));
	assign g221 = (((!g6) & (!i_15_) & (sk[111]) & (!g91)) + ((!g6) & (!i_15_) & (sk[111]) & (g91)) + ((!g6) & (i_15_) & (sk[111]) & (!g91)) + ((!g6) & (i_15_) & (sk[111]) & (g91)) + ((g6) & (!i_15_) & (!sk[111]) & (!g91)) + ((g6) & (!i_15_) & (!sk[111]) & (g91)) + ((g6) & (!i_15_) & (sk[111]) & (g91)) + ((g6) & (i_15_) & (!sk[111]) & (!g91)) + ((g6) & (i_15_) & (!sk[111]) & (g91)) + ((g6) & (i_15_) & (sk[111]) & (!g91)) + ((g6) & (i_15_) & (sk[111]) & (g91)));
	assign g222 = (((!sk[112]) & (g15) & (!g91)) + ((!sk[112]) & (g15) & (g91)) + ((sk[112]) & (!g15) & (!g91)));
	assign g223 = (((!g99) & (!g220) & (!sk[113]) & (g221) & (g222)) + ((!g99) & (g220) & (!sk[113]) & (!g221) & (!g222)) + ((!g99) & (g220) & (!sk[113]) & (!g221) & (g222)) + ((!g99) & (g220) & (!sk[113]) & (g221) & (!g222)) + ((!g99) & (g220) & (!sk[113]) & (g221) & (g222)) + ((g99) & (!g220) & (!sk[113]) & (g221) & (!g222)) + ((g99) & (!g220) & (!sk[113]) & (g221) & (g222)) + ((g99) & (!g220) & (sk[113]) & (!g221) & (!g222)) + ((g99) & (!g220) & (sk[113]) & (!g221) & (g222)) + ((g99) & (!g220) & (sk[113]) & (g221) & (g222)) + ((g99) & (g220) & (!sk[113]) & (!g221) & (!g222)) + ((g99) & (g220) & (!sk[113]) & (!g221) & (g222)) + ((g99) & (g220) & (!sk[113]) & (g221) & (!g222)) + ((g99) & (g220) & (!sk[113]) & (g221) & (g222)) + ((g99) & (g220) & (sk[113]) & (!g221) & (!g222)) + ((g99) & (g220) & (sk[113]) & (!g221) & (g222)) + ((g99) & (g220) & (sk[113]) & (g221) & (!g222)) + ((g99) & (g220) & (sk[113]) & (g221) & (g222)));
	assign g224 = (((g6) & (!sk[114]) & (!i_15_) & (!g182)) + ((g6) & (!sk[114]) & (!i_15_) & (g182)) + ((g6) & (!sk[114]) & (i_15_) & (!g182)) + ((g6) & (!sk[114]) & (i_15_) & (g182)) + ((g6) & (sk[114]) & (i_15_) & (g182)));
	assign g225 = (((!g99) & (!g183) & (g224) & (!sk[115]) & (g213)) + ((!g99) & (g183) & (!g224) & (!sk[115]) & (!g213)) + ((!g99) & (g183) & (!g224) & (!sk[115]) & (g213)) + ((!g99) & (g183) & (g224) & (!sk[115]) & (!g213)) + ((!g99) & (g183) & (g224) & (!sk[115]) & (g213)) + ((g99) & (!g183) & (!g224) & (sk[115]) & (g213)) + ((g99) & (!g183) & (g224) & (!sk[115]) & (!g213)) + ((g99) & (!g183) & (g224) & (!sk[115]) & (g213)) + ((g99) & (!g183) & (g224) & (sk[115]) & (!g213)) + ((g99) & (!g183) & (g224) & (sk[115]) & (g213)) + ((g99) & (g183) & (!g224) & (!sk[115]) & (!g213)) + ((g99) & (g183) & (!g224) & (!sk[115]) & (g213)) + ((g99) & (g183) & (!g224) & (sk[115]) & (!g213)) + ((g99) & (g183) & (!g224) & (sk[115]) & (g213)) + ((g99) & (g183) & (g224) & (!sk[115]) & (!g213)) + ((g99) & (g183) & (g224) & (!sk[115]) & (g213)) + ((g99) & (g183) & (g224) & (sk[115]) & (!g213)) + ((g99) & (g183) & (g224) & (sk[115]) & (g213)));
	assign g226 = (((!sk[116]) & (g22) & (!g182)) + ((!sk[116]) & (g22) & (g182)) + ((sk[116]) & (!g22) & (!g182)) + ((sk[116]) & (!g22) & (g182)) + ((sk[116]) & (g22) & (!g182)));
	assign g227 = (((g38) & (!sk[117]) & (!g87)) + ((g38) & (!sk[117]) & (g87)) + ((g38) & (sk[117]) & (g87)));
	assign g228 = (((!i_11_) & (!i_9_) & (i_10_) & (!sk[118]) & (i_15_)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[118]) & (!i_15_)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[118]) & (i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[118]) & (!i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[118]) & (i_15_)) + ((!i_11_) & (i_9_) & (i_10_) & (sk[118]) & (i_15_)) + ((i_11_) & (!i_9_) & (!i_10_) & (sk[118]) & (i_15_)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[118]) & (!i_15_)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[118]) & (i_15_)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[118]) & (!i_15_)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[118]) & (i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[118]) & (!i_15_)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[118]) & (i_15_)));
	assign g229 = (((!i_3_) & (i_4_) & (g57) & (g38) & (g182) & (g228)));
	assign g230 = (((!sk[120]) & (!g99) & (!g226) & (!g203) & (!g227) & (g229)) + ((!sk[120]) & (!g99) & (!g226) & (!g203) & (g227) & (g229)) + ((!sk[120]) & (!g99) & (!g226) & (g203) & (!g227) & (g229)) + ((!sk[120]) & (!g99) & (!g226) & (g203) & (g227) & (g229)) + ((!sk[120]) & (!g99) & (g226) & (!g203) & (!g227) & (g229)) + ((!sk[120]) & (!g99) & (g226) & (!g203) & (g227) & (g229)) + ((!sk[120]) & (!g99) & (g226) & (g203) & (!g227) & (g229)) + ((!sk[120]) & (!g99) & (g226) & (g203) & (g227) & (g229)) + ((!sk[120]) & (g99) & (!g226) & (!g203) & (!g227) & (!g229)) + ((!sk[120]) & (g99) & (!g226) & (!g203) & (!g227) & (g229)) + ((!sk[120]) & (g99) & (!g226) & (!g203) & (g227) & (!g229)) + ((!sk[120]) & (g99) & (!g226) & (!g203) & (g227) & (g229)) + ((!sk[120]) & (g99) & (!g226) & (g203) & (!g227) & (!g229)) + ((!sk[120]) & (g99) & (!g226) & (g203) & (!g227) & (g229)) + ((!sk[120]) & (g99) & (!g226) & (g203) & (g227) & (!g229)) + ((!sk[120]) & (g99) & (!g226) & (g203) & (g227) & (g229)) + ((!sk[120]) & (g99) & (g226) & (!g203) & (!g227) & (!g229)) + ((!sk[120]) & (g99) & (g226) & (!g203) & (!g227) & (g229)) + ((!sk[120]) & (g99) & (g226) & (!g203) & (g227) & (!g229)) + ((!sk[120]) & (g99) & (g226) & (!g203) & (g227) & (g229)) + ((!sk[120]) & (g99) & (g226) & (g203) & (!g227) & (!g229)) + ((!sk[120]) & (g99) & (g226) & (g203) & (!g227) & (g229)) + ((!sk[120]) & (g99) & (g226) & (g203) & (g227) & (!g229)) + ((!sk[120]) & (g99) & (g226) & (g203) & (g227) & (g229)) + ((sk[120]) & (!g99) & (!g226) & (!g203) & (g227) & (g229)) + ((sk[120]) & (!g99) & (!g226) & (g203) & (!g227) & (g229)) + ((sk[120]) & (!g99) & (!g226) & (g203) & (g227) & (g229)) + ((sk[120]) & (g99) & (!g226) & (!g203) & (g227) & (g229)) + ((sk[120]) & (g99) & (!g226) & (g203) & (!g227) & (g229)) + ((sk[120]) & (g99) & (!g226) & (g203) & (g227) & (g229)) + ((sk[120]) & (g99) & (g226) & (!g203) & (g227) & (g229)) + ((sk[120]) & (g99) & (g226) & (g203) & (!g227) & (g229)) + ((sk[120]) & (g99) & (g226) & (g203) & (g227) & (g229)));
	assign g231 = (((!sk[121]) & (g182) & (!g124)) + ((!sk[121]) & (g182) & (g124)) + ((sk[121]) & (!g182) & (!g124)) + ((sk[121]) & (!g182) & (g124)) + ((sk[121]) & (g182) & (!g124)));
	assign g232 = (((g182) & (!sk[122]) & (!g115)) + ((g182) & (!sk[122]) & (g115)) + ((g182) & (sk[122]) & (!g115)));
	assign g233 = (((!g99) & (!g193) & (g231) & (!sk[123]) & (g232)) + ((!g99) & (g193) & (!g231) & (!sk[123]) & (!g232)) + ((!g99) & (g193) & (!g231) & (!sk[123]) & (g232)) + ((!g99) & (g193) & (g231) & (!sk[123]) & (!g232)) + ((!g99) & (g193) & (g231) & (!sk[123]) & (g232)) + ((g99) & (!g193) & (!g231) & (sk[123]) & (!g232)) + ((g99) & (!g193) & (!g231) & (sk[123]) & (g232)) + ((g99) & (!g193) & (g231) & (!sk[123]) & (!g232)) + ((g99) & (!g193) & (g231) & (!sk[123]) & (g232)) + ((g99) & (!g193) & (g231) & (sk[123]) & (g232)) + ((g99) & (g193) & (!g231) & (!sk[123]) & (!g232)) + ((g99) & (g193) & (!g231) & (!sk[123]) & (g232)) + ((g99) & (g193) & (!g231) & (sk[123]) & (!g232)) + ((g99) & (g193) & (!g231) & (sk[123]) & (g232)) + ((g99) & (g193) & (g231) & (!sk[123]) & (!g232)) + ((g99) & (g193) & (g231) & (!sk[123]) & (g232)) + ((g99) & (g193) & (g231) & (sk[123]) & (!g232)) + ((g99) & (g193) & (g231) & (sk[123]) & (g232)));
	assign g234 = (((!sk[124]) & (!g219) & (!g223) & (!g225) & (!g230) & (g233)) + ((!sk[124]) & (!g219) & (!g223) & (!g225) & (g230) & (g233)) + ((!sk[124]) & (!g219) & (!g223) & (g225) & (!g230) & (g233)) + ((!sk[124]) & (!g219) & (!g223) & (g225) & (g230) & (g233)) + ((!sk[124]) & (!g219) & (g223) & (!g225) & (!g230) & (g233)) + ((!sk[124]) & (!g219) & (g223) & (!g225) & (g230) & (g233)) + ((!sk[124]) & (!g219) & (g223) & (g225) & (!g230) & (g233)) + ((!sk[124]) & (!g219) & (g223) & (g225) & (g230) & (g233)) + ((!sk[124]) & (g219) & (!g223) & (!g225) & (!g230) & (!g233)) + ((!sk[124]) & (g219) & (!g223) & (!g225) & (!g230) & (g233)) + ((!sk[124]) & (g219) & (!g223) & (!g225) & (g230) & (!g233)) + ((!sk[124]) & (g219) & (!g223) & (!g225) & (g230) & (g233)) + ((!sk[124]) & (g219) & (!g223) & (g225) & (!g230) & (!g233)) + ((!sk[124]) & (g219) & (!g223) & (g225) & (!g230) & (g233)) + ((!sk[124]) & (g219) & (!g223) & (g225) & (g230) & (!g233)) + ((!sk[124]) & (g219) & (!g223) & (g225) & (g230) & (g233)) + ((!sk[124]) & (g219) & (g223) & (!g225) & (!g230) & (!g233)) + ((!sk[124]) & (g219) & (g223) & (!g225) & (!g230) & (g233)) + ((!sk[124]) & (g219) & (g223) & (!g225) & (g230) & (!g233)) + ((!sk[124]) & (g219) & (g223) & (!g225) & (g230) & (g233)) + ((!sk[124]) & (g219) & (g223) & (g225) & (!g230) & (!g233)) + ((!sk[124]) & (g219) & (g223) & (g225) & (!g230) & (g233)) + ((!sk[124]) & (g219) & (g223) & (g225) & (g230) & (!g233)) + ((!sk[124]) & (g219) & (g223) & (g225) & (g230) & (g233)) + ((sk[124]) & (!g219) & (!g223) & (!g225) & (!g230) & (!g233)));
	assign g235 = (((!g176) & (g189) & (g1543) & (g211) & (g218) & (g234)));
	assign g236 = (((!sk[126]) & (i_8_) & (!g34) & (!g110)) + ((!sk[126]) & (i_8_) & (!g34) & (g110)) + ((!sk[126]) & (i_8_) & (g34) & (!g110)) + ((!sk[126]) & (i_8_) & (g34) & (g110)) + ((sk[126]) & (!i_8_) & (g34) & (g110)));
	assign g237 = (((g6) & (!sk[127]) & (!g236)) + ((g6) & (!sk[127]) & (g236)) + ((g6) & (sk[127]) & (g236)));
	assign g238 = (((g31) & (!sk[0]) & (!g98)) + ((g31) & (!sk[0]) & (g98)) + ((g31) & (sk[0]) & (g98)));
	assign g239 = (((!sk[1]) & (g227) & (!g224)) + ((!sk[1]) & (g227) & (g224)) + ((sk[1]) & (g227) & (g224)));
	assign g240 = (((g99) & (!g187) & (!sk[2]) & (!g209)) + ((g99) & (!g187) & (!sk[2]) & (g209)) + ((g99) & (!g187) & (sk[2]) & (g209)) + ((g99) & (g187) & (!sk[2]) & (!g209)) + ((g99) & (g187) & (!sk[2]) & (g209)) + ((g99) & (g187) & (sk[2]) & (!g209)) + ((g99) & (g187) & (sk[2]) & (g209)));
	assign g241 = (((!sk[3]) & (!i_8_) & (!g108) & (g183) & (g201)) + ((!sk[3]) & (!i_8_) & (g108) & (!g183) & (!g201)) + ((!sk[3]) & (!i_8_) & (g108) & (!g183) & (g201)) + ((!sk[3]) & (!i_8_) & (g108) & (g183) & (!g201)) + ((!sk[3]) & (!i_8_) & (g108) & (g183) & (g201)) + ((!sk[3]) & (i_8_) & (!g108) & (g183) & (!g201)) + ((!sk[3]) & (i_8_) & (!g108) & (g183) & (g201)) + ((!sk[3]) & (i_8_) & (g108) & (!g183) & (!g201)) + ((!sk[3]) & (i_8_) & (g108) & (!g183) & (g201)) + ((!sk[3]) & (i_8_) & (g108) & (g183) & (!g201)) + ((!sk[3]) & (i_8_) & (g108) & (g183) & (g201)) + ((sk[3]) & (!i_8_) & (g108) & (!g183) & (!g201)) + ((sk[3]) & (!i_8_) & (g108) & (g183) & (!g201)) + ((sk[3]) & (!i_8_) & (g108) & (g183) & (g201)));
	assign g242 = (((!g14) & (!g237) & (!g238) & (!g239) & (!g240) & (!g241)) + ((!g14) & (!g237) & (g238) & (!g239) & (!g240) & (!g241)) + ((g14) & (!g237) & (!g238) & (!g239) & (!g240) & (!g241)));
	assign g243 = (((!sk[5]) & (g30) & (!g87)) + ((!sk[5]) & (g30) & (g87)) + ((sk[5]) & (g30) & (g87)));
	assign g244 = (((!i_15_) & (sk[6]) & (!g91)) + ((i_15_) & (!sk[6]) & (!g91)) + ((i_15_) & (!sk[6]) & (g91)));
	assign g245 = (((!i_11_) & (!i_9_) & (!sk[7]) & (i_10_) & (g244)) + ((!i_11_) & (i_9_) & (!sk[7]) & (!i_10_) & (!g244)) + ((!i_11_) & (i_9_) & (!sk[7]) & (!i_10_) & (g244)) + ((!i_11_) & (i_9_) & (!sk[7]) & (i_10_) & (!g244)) + ((!i_11_) & (i_9_) & (!sk[7]) & (i_10_) & (g244)) + ((!i_11_) & (i_9_) & (sk[7]) & (i_10_) & (g244)) + ((i_11_) & (!i_9_) & (!sk[7]) & (i_10_) & (!g244)) + ((i_11_) & (!i_9_) & (!sk[7]) & (i_10_) & (g244)) + ((i_11_) & (i_9_) & (!sk[7]) & (!i_10_) & (!g244)) + ((i_11_) & (i_9_) & (!sk[7]) & (!i_10_) & (g244)) + ((i_11_) & (i_9_) & (!sk[7]) & (i_10_) & (!g244)) + ((i_11_) & (i_9_) & (!sk[7]) & (i_10_) & (g244)) + ((i_11_) & (i_9_) & (sk[7]) & (!i_10_) & (g244)));
	assign g246 = (((!i_14_) & (!i_12_) & (i_13_) & (!sk[8]) & (g131)) + ((!i_14_) & (i_12_) & (!i_13_) & (!sk[8]) & (!g131)) + ((!i_14_) & (i_12_) & (!i_13_) & (!sk[8]) & (g131)) + ((!i_14_) & (i_12_) & (i_13_) & (!sk[8]) & (!g131)) + ((!i_14_) & (i_12_) & (i_13_) & (!sk[8]) & (g131)) + ((i_14_) & (!i_12_) & (!i_13_) & (sk[8]) & (g131)) + ((i_14_) & (!i_12_) & (i_13_) & (!sk[8]) & (!g131)) + ((i_14_) & (!i_12_) & (i_13_) & (!sk[8]) & (g131)) + ((i_14_) & (!i_12_) & (i_13_) & (sk[8]) & (g131)) + ((i_14_) & (i_12_) & (!i_13_) & (!sk[8]) & (!g131)) + ((i_14_) & (i_12_) & (!i_13_) & (!sk[8]) & (g131)) + ((i_14_) & (i_12_) & (i_13_) & (!sk[8]) & (!g131)) + ((i_14_) & (i_12_) & (i_13_) & (!sk[8]) & (g131)) + ((i_14_) & (i_12_) & (i_13_) & (sk[8]) & (g131)));
	assign g247 = (((!g221) & (!g183) & (!sk[9]) & (g199) & (g197)) + ((!g221) & (g183) & (!sk[9]) & (!g199) & (!g197)) + ((!g221) & (g183) & (!sk[9]) & (!g199) & (g197)) + ((!g221) & (g183) & (!sk[9]) & (g199) & (!g197)) + ((!g221) & (g183) & (!sk[9]) & (g199) & (g197)) + ((g221) & (!g183) & (!sk[9]) & (g199) & (!g197)) + ((g221) & (!g183) & (!sk[9]) & (g199) & (g197)) + ((g221) & (!g183) & (sk[9]) & (!g199) & (!g197)) + ((g221) & (g183) & (!sk[9]) & (!g199) & (!g197)) + ((g221) & (g183) & (!sk[9]) & (!g199) & (g197)) + ((g221) & (g183) & (!sk[9]) & (g199) & (!g197)) + ((g221) & (g183) & (!sk[9]) & (g199) & (g197)));
	assign g248 = (((!g245) & (!sk[10]) & (!g185) & (!g246) & (!g120) & (g247)) + ((!g245) & (!sk[10]) & (!g185) & (!g246) & (g120) & (g247)) + ((!g245) & (!sk[10]) & (!g185) & (g246) & (!g120) & (g247)) + ((!g245) & (!sk[10]) & (!g185) & (g246) & (g120) & (g247)) + ((!g245) & (!sk[10]) & (g185) & (!g246) & (!g120) & (g247)) + ((!g245) & (!sk[10]) & (g185) & (!g246) & (g120) & (g247)) + ((!g245) & (!sk[10]) & (g185) & (g246) & (!g120) & (g247)) + ((!g245) & (!sk[10]) & (g185) & (g246) & (g120) & (g247)) + ((!g245) & (sk[10]) & (g185) & (!g246) & (g120) & (g247)) + ((g245) & (!sk[10]) & (!g185) & (!g246) & (!g120) & (!g247)) + ((g245) & (!sk[10]) & (!g185) & (!g246) & (!g120) & (g247)) + ((g245) & (!sk[10]) & (!g185) & (!g246) & (g120) & (!g247)) + ((g245) & (!sk[10]) & (!g185) & (!g246) & (g120) & (g247)) + ((g245) & (!sk[10]) & (!g185) & (g246) & (!g120) & (!g247)) + ((g245) & (!sk[10]) & (!g185) & (g246) & (!g120) & (g247)) + ((g245) & (!sk[10]) & (!g185) & (g246) & (g120) & (!g247)) + ((g245) & (!sk[10]) & (!g185) & (g246) & (g120) & (g247)) + ((g245) & (!sk[10]) & (g185) & (!g246) & (!g120) & (!g247)) + ((g245) & (!sk[10]) & (g185) & (!g246) & (!g120) & (g247)) + ((g245) & (!sk[10]) & (g185) & (!g246) & (g120) & (!g247)) + ((g245) & (!sk[10]) & (g185) & (!g246) & (g120) & (g247)) + ((g245) & (!sk[10]) & (g185) & (g246) & (!g120) & (!g247)) + ((g245) & (!sk[10]) & (g185) & (g246) & (!g120) & (g247)) + ((g245) & (!sk[10]) & (g185) & (g246) & (g120) & (!g247)) + ((g245) & (!sk[10]) & (g185) & (g246) & (g120) & (g247)));
	assign g249 = (((!i_14_) & (!sk[11]) & (!i_12_) & (!i_13_) & (!g100) & (g108)) + ((!i_14_) & (!sk[11]) & (!i_12_) & (!i_13_) & (g100) & (g108)) + ((!i_14_) & (!sk[11]) & (!i_12_) & (i_13_) & (!g100) & (g108)) + ((!i_14_) & (!sk[11]) & (!i_12_) & (i_13_) & (g100) & (g108)) + ((!i_14_) & (!sk[11]) & (i_12_) & (!i_13_) & (!g100) & (g108)) + ((!i_14_) & (!sk[11]) & (i_12_) & (!i_13_) & (g100) & (g108)) + ((!i_14_) & (!sk[11]) & (i_12_) & (i_13_) & (!g100) & (g108)) + ((!i_14_) & (!sk[11]) & (i_12_) & (i_13_) & (g100) & (g108)) + ((!i_14_) & (sk[11]) & (i_12_) & (!i_13_) & (g100) & (!g108)) + ((!i_14_) & (sk[11]) & (i_12_) & (!i_13_) & (g100) & (g108)) + ((i_14_) & (!sk[11]) & (!i_12_) & (!i_13_) & (!g100) & (!g108)) + ((i_14_) & (!sk[11]) & (!i_12_) & (!i_13_) & (!g100) & (g108)) + ((i_14_) & (!sk[11]) & (!i_12_) & (!i_13_) & (g100) & (!g108)) + ((i_14_) & (!sk[11]) & (!i_12_) & (!i_13_) & (g100) & (g108)) + ((i_14_) & (!sk[11]) & (!i_12_) & (i_13_) & (!g100) & (!g108)) + ((i_14_) & (!sk[11]) & (!i_12_) & (i_13_) & (!g100) & (g108)) + ((i_14_) & (!sk[11]) & (!i_12_) & (i_13_) & (g100) & (!g108)) + ((i_14_) & (!sk[11]) & (!i_12_) & (i_13_) & (g100) & (g108)) + ((i_14_) & (!sk[11]) & (i_12_) & (!i_13_) & (!g100) & (!g108)) + ((i_14_) & (!sk[11]) & (i_12_) & (!i_13_) & (!g100) & (g108)) + ((i_14_) & (!sk[11]) & (i_12_) & (!i_13_) & (g100) & (!g108)) + ((i_14_) & (!sk[11]) & (i_12_) & (!i_13_) & (g100) & (g108)) + ((i_14_) & (!sk[11]) & (i_12_) & (i_13_) & (!g100) & (!g108)) + ((i_14_) & (!sk[11]) & (i_12_) & (i_13_) & (!g100) & (g108)) + ((i_14_) & (!sk[11]) & (i_12_) & (i_13_) & (g100) & (!g108)) + ((i_14_) & (!sk[11]) & (i_12_) & (i_13_) & (g100) & (g108)) + ((i_14_) & (sk[11]) & (i_12_) & (i_13_) & (!g100) & (g108)) + ((i_14_) & (sk[11]) & (i_12_) & (i_13_) & (g100) & (g108)));
	assign g250 = (((!sk[12]) & (!g119) & (!g243) & (g248) & (g249)) + ((!sk[12]) & (!g119) & (g243) & (!g248) & (!g249)) + ((!sk[12]) & (!g119) & (g243) & (!g248) & (g249)) + ((!sk[12]) & (!g119) & (g243) & (g248) & (!g249)) + ((!sk[12]) & (!g119) & (g243) & (g248) & (g249)) + ((!sk[12]) & (g119) & (!g243) & (g248) & (!g249)) + ((!sk[12]) & (g119) & (!g243) & (g248) & (g249)) + ((!sk[12]) & (g119) & (g243) & (!g248) & (!g249)) + ((!sk[12]) & (g119) & (g243) & (!g248) & (g249)) + ((!sk[12]) & (g119) & (g243) & (g248) & (!g249)) + ((!sk[12]) & (g119) & (g243) & (g248) & (g249)) + ((sk[12]) & (!g119) & (g243) & (!g248) & (!g249)) + ((sk[12]) & (!g119) & (g243) & (!g248) & (g249)) + ((sk[12]) & (g119) & (!g243) & (!g248) & (g249)) + ((sk[12]) & (g119) & (!g243) & (g248) & (g249)) + ((sk[12]) & (g119) & (g243) & (!g248) & (!g249)) + ((sk[12]) & (g119) & (g243) & (!g248) & (g249)) + ((sk[12]) & (g119) & (g243) & (g248) & (g249)));
	assign g251 = (((!i_8_) & (!g88) & (!g118) & (sk[13]) & (g243)) + ((!i_8_) & (!g88) & (g118) & (!sk[13]) & (g243)) + ((!i_8_) & (!g88) & (g118) & (sk[13]) & (!g243)) + ((!i_8_) & (!g88) & (g118) & (sk[13]) & (g243)) + ((!i_8_) & (g88) & (!g118) & (!sk[13]) & (!g243)) + ((!i_8_) & (g88) & (!g118) & (!sk[13]) & (g243)) + ((!i_8_) & (g88) & (!g118) & (sk[13]) & (!g243)) + ((!i_8_) & (g88) & (!g118) & (sk[13]) & (g243)) + ((!i_8_) & (g88) & (g118) & (!sk[13]) & (!g243)) + ((!i_8_) & (g88) & (g118) & (!sk[13]) & (g243)) + ((!i_8_) & (g88) & (g118) & (sk[13]) & (!g243)) + ((!i_8_) & (g88) & (g118) & (sk[13]) & (g243)) + ((i_8_) & (!g88) & (!g118) & (sk[13]) & (g243)) + ((i_8_) & (!g88) & (g118) & (!sk[13]) & (!g243)) + ((i_8_) & (!g88) & (g118) & (!sk[13]) & (g243)) + ((i_8_) & (!g88) & (g118) & (sk[13]) & (!g243)) + ((i_8_) & (!g88) & (g118) & (sk[13]) & (g243)) + ((i_8_) & (g88) & (!g118) & (!sk[13]) & (!g243)) + ((i_8_) & (g88) & (!g118) & (!sk[13]) & (g243)) + ((i_8_) & (g88) & (!g118) & (sk[13]) & (g243)) + ((i_8_) & (g88) & (g118) & (!sk[13]) & (!g243)) + ((i_8_) & (g88) & (g118) & (!sk[13]) & (g243)) + ((i_8_) & (g88) & (g118) & (sk[13]) & (!g243)) + ((i_8_) & (g88) & (g118) & (sk[13]) & (g243)));
	assign g252 = (((!i_11_) & (!i_9_) & (!sk[14]) & (!i_10_) & (!i_15_) & (g171)) + ((!i_11_) & (!i_9_) & (!sk[14]) & (!i_10_) & (i_15_) & (g171)) + ((!i_11_) & (!i_9_) & (!sk[14]) & (i_10_) & (!i_15_) & (g171)) + ((!i_11_) & (!i_9_) & (!sk[14]) & (i_10_) & (i_15_) & (g171)) + ((!i_11_) & (i_9_) & (!sk[14]) & (!i_10_) & (!i_15_) & (g171)) + ((!i_11_) & (i_9_) & (!sk[14]) & (!i_10_) & (i_15_) & (g171)) + ((!i_11_) & (i_9_) & (!sk[14]) & (i_10_) & (!i_15_) & (g171)) + ((!i_11_) & (i_9_) & (!sk[14]) & (i_10_) & (i_15_) & (g171)) + ((i_11_) & (!i_9_) & (!sk[14]) & (!i_10_) & (!i_15_) & (!g171)) + ((i_11_) & (!i_9_) & (!sk[14]) & (!i_10_) & (!i_15_) & (g171)) + ((i_11_) & (!i_9_) & (!sk[14]) & (!i_10_) & (i_15_) & (!g171)) + ((i_11_) & (!i_9_) & (!sk[14]) & (!i_10_) & (i_15_) & (g171)) + ((i_11_) & (!i_9_) & (!sk[14]) & (i_10_) & (!i_15_) & (!g171)) + ((i_11_) & (!i_9_) & (!sk[14]) & (i_10_) & (!i_15_) & (g171)) + ((i_11_) & (!i_9_) & (!sk[14]) & (i_10_) & (i_15_) & (!g171)) + ((i_11_) & (!i_9_) & (!sk[14]) & (i_10_) & (i_15_) & (g171)) + ((i_11_) & (!i_9_) & (sk[14]) & (!i_10_) & (!i_15_) & (!g171)) + ((i_11_) & (i_9_) & (!sk[14]) & (!i_10_) & (!i_15_) & (!g171)) + ((i_11_) & (i_9_) & (!sk[14]) & (!i_10_) & (!i_15_) & (g171)) + ((i_11_) & (i_9_) & (!sk[14]) & (!i_10_) & (i_15_) & (!g171)) + ((i_11_) & (i_9_) & (!sk[14]) & (!i_10_) & (i_15_) & (g171)) + ((i_11_) & (i_9_) & (!sk[14]) & (i_10_) & (!i_15_) & (!g171)) + ((i_11_) & (i_9_) & (!sk[14]) & (i_10_) & (!i_15_) & (g171)) + ((i_11_) & (i_9_) & (!sk[14]) & (i_10_) & (i_15_) & (!g171)) + ((i_11_) & (i_9_) & (!sk[14]) & (i_10_) & (i_15_) & (g171)) + ((i_11_) & (i_9_) & (sk[14]) & (i_10_) & (!i_15_) & (!g171)));
	assign g253 = (((g131) & (!sk[15]) & (!g182)) + ((g131) & (!sk[15]) & (g182)) + ((g131) & (sk[15]) & (g182)));
	assign g254 = (((!i_15_) & (g141) & (sk[16]) & (!g171)) + ((i_15_) & (!g141) & (!sk[16]) & (!g171)) + ((i_15_) & (!g141) & (!sk[16]) & (g171)) + ((i_15_) & (g141) & (!sk[16]) & (!g171)) + ((i_15_) & (g141) & (!sk[16]) & (g171)));
	assign g255 = (((!sk[17]) & (g141) & (!g244)) + ((!sk[17]) & (g141) & (g244)) + ((sk[17]) & (g141) & (g244)));
	assign g256 = (((!g193) & (!sk[18]) & (!g177) & (!g253) & (!g254) & (g255)) + ((!g193) & (!sk[18]) & (!g177) & (!g253) & (g254) & (g255)) + ((!g193) & (!sk[18]) & (!g177) & (g253) & (!g254) & (g255)) + ((!g193) & (!sk[18]) & (!g177) & (g253) & (g254) & (g255)) + ((!g193) & (!sk[18]) & (g177) & (!g253) & (!g254) & (g255)) + ((!g193) & (!sk[18]) & (g177) & (!g253) & (g254) & (g255)) + ((!g193) & (!sk[18]) & (g177) & (g253) & (!g254) & (g255)) + ((!g193) & (!sk[18]) & (g177) & (g253) & (g254) & (g255)) + ((!g193) & (sk[18]) & (!g177) & (!g253) & (!g254) & (!g255)) + ((g193) & (!sk[18]) & (!g177) & (!g253) & (!g254) & (!g255)) + ((g193) & (!sk[18]) & (!g177) & (!g253) & (!g254) & (g255)) + ((g193) & (!sk[18]) & (!g177) & (!g253) & (g254) & (!g255)) + ((g193) & (!sk[18]) & (!g177) & (!g253) & (g254) & (g255)) + ((g193) & (!sk[18]) & (!g177) & (g253) & (!g254) & (!g255)) + ((g193) & (!sk[18]) & (!g177) & (g253) & (!g254) & (g255)) + ((g193) & (!sk[18]) & (!g177) & (g253) & (g254) & (!g255)) + ((g193) & (!sk[18]) & (!g177) & (g253) & (g254) & (g255)) + ((g193) & (!sk[18]) & (g177) & (!g253) & (!g254) & (!g255)) + ((g193) & (!sk[18]) & (g177) & (!g253) & (!g254) & (g255)) + ((g193) & (!sk[18]) & (g177) & (!g253) & (g254) & (!g255)) + ((g193) & (!sk[18]) & (g177) & (!g253) & (g254) & (g255)) + ((g193) & (!sk[18]) & (g177) & (g253) & (!g254) & (!g255)) + ((g193) & (!sk[18]) & (g177) & (g253) & (!g254) & (g255)) + ((g193) & (!sk[18]) & (g177) & (g253) & (g254) & (!g255)) + ((g193) & (!sk[18]) & (g177) & (g253) & (g254) & (g255)));
	assign g257 = (((!g6) & (!sk[19]) & (!i_15_) & (i_14_) & (i_12_)) + ((!g6) & (!sk[19]) & (i_15_) & (!i_14_) & (!i_12_)) + ((!g6) & (!sk[19]) & (i_15_) & (!i_14_) & (i_12_)) + ((!g6) & (!sk[19]) & (i_15_) & (i_14_) & (!i_12_)) + ((!g6) & (!sk[19]) & (i_15_) & (i_14_) & (i_12_)) + ((g6) & (!sk[19]) & (!i_15_) & (i_14_) & (!i_12_)) + ((g6) & (!sk[19]) & (!i_15_) & (i_14_) & (i_12_)) + ((g6) & (!sk[19]) & (i_15_) & (!i_14_) & (!i_12_)) + ((g6) & (!sk[19]) & (i_15_) & (!i_14_) & (i_12_)) + ((g6) & (!sk[19]) & (i_15_) & (i_14_) & (!i_12_)) + ((g6) & (!sk[19]) & (i_15_) & (i_14_) & (i_12_)) + ((g6) & (sk[19]) & (!i_15_) & (i_14_) & (i_12_)));
	assign g258 = (((!g212) & (!g251) & (!g252) & (!g256) & (!sk[20]) & (g257)) + ((!g212) & (!g251) & (!g252) & (!g256) & (sk[20]) & (!g257)) + ((!g212) & (!g251) & (!g252) & (g256) & (!sk[20]) & (g257)) + ((!g212) & (!g251) & (!g252) & (g256) & (sk[20]) & (!g257)) + ((!g212) & (!g251) & (g252) & (!g256) & (!sk[20]) & (g257)) + ((!g212) & (!g251) & (g252) & (!g256) & (sk[20]) & (!g257)) + ((!g212) & (!g251) & (g252) & (g256) & (!sk[20]) & (g257)) + ((!g212) & (!g251) & (g252) & (g256) & (sk[20]) & (!g257)) + ((!g212) & (g251) & (!g252) & (!g256) & (!sk[20]) & (g257)) + ((!g212) & (g251) & (!g252) & (g256) & (!sk[20]) & (g257)) + ((!g212) & (g251) & (!g252) & (g256) & (sk[20]) & (!g257)) + ((!g212) & (g251) & (g252) & (!g256) & (!sk[20]) & (g257)) + ((!g212) & (g251) & (g252) & (g256) & (!sk[20]) & (g257)) + ((g212) & (!g251) & (!g252) & (!g256) & (!sk[20]) & (!g257)) + ((g212) & (!g251) & (!g252) & (!g256) & (!sk[20]) & (g257)) + ((g212) & (!g251) & (!g252) & (!g256) & (sk[20]) & (!g257)) + ((g212) & (!g251) & (!g252) & (!g256) & (sk[20]) & (g257)) + ((g212) & (!g251) & (!g252) & (g256) & (!sk[20]) & (!g257)) + ((g212) & (!g251) & (!g252) & (g256) & (!sk[20]) & (g257)) + ((g212) & (!g251) & (!g252) & (g256) & (sk[20]) & (!g257)) + ((g212) & (!g251) & (!g252) & (g256) & (sk[20]) & (g257)) + ((g212) & (!g251) & (g252) & (!g256) & (!sk[20]) & (!g257)) + ((g212) & (!g251) & (g252) & (!g256) & (!sk[20]) & (g257)) + ((g212) & (!g251) & (g252) & (!g256) & (sk[20]) & (!g257)) + ((g212) & (!g251) & (g252) & (!g256) & (sk[20]) & (g257)) + ((g212) & (!g251) & (g252) & (g256) & (!sk[20]) & (!g257)) + ((g212) & (!g251) & (g252) & (g256) & (!sk[20]) & (g257)) + ((g212) & (!g251) & (g252) & (g256) & (sk[20]) & (!g257)) + ((g212) & (!g251) & (g252) & (g256) & (sk[20]) & (g257)) + ((g212) & (g251) & (!g252) & (!g256) & (!sk[20]) & (!g257)) + ((g212) & (g251) & (!g252) & (!g256) & (!sk[20]) & (g257)) + ((g212) & (g251) & (!g252) & (g256) & (!sk[20]) & (!g257)) + ((g212) & (g251) & (!g252) & (g256) & (!sk[20]) & (g257)) + ((g212) & (g251) & (!g252) & (g256) & (sk[20]) & (!g257)) + ((g212) & (g251) & (!g252) & (g256) & (sk[20]) & (g257)) + ((g212) & (g251) & (g252) & (!g256) & (!sk[20]) & (!g257)) + ((g212) & (g251) & (g252) & (!g256) & (!sk[20]) & (g257)) + ((g212) & (g251) & (g252) & (g256) & (!sk[20]) & (!g257)) + ((g212) & (g251) & (g252) & (g256) & (!sk[20]) & (g257)));
	assign g259 = (((!g207) & (sk[21]) & (g204)) + ((g207) & (!sk[21]) & (!g204)) + ((g207) & (!sk[21]) & (g204)));
	assign g260 = (((!i_11_) & (g113) & (sk[22]) & (g236)) + ((i_11_) & (!g113) & (!sk[22]) & (!g236)) + ((i_11_) & (!g113) & (!sk[22]) & (g236)) + ((i_11_) & (g113) & (!sk[22]) & (!g236)) + ((i_11_) & (g113) & (!sk[22]) & (g236)));
	assign g261 = (((!sk[23]) & (i_8_) & (!g88) & (!g231)) + ((!sk[23]) & (i_8_) & (!g88) & (g231)) + ((!sk[23]) & (i_8_) & (g88) & (!g231)) + ((!sk[23]) & (i_8_) & (g88) & (g231)) + ((sk[23]) & (i_8_) & (g88) & (!g231)));
	assign g262 = (((!i_8_) & (!g30) & (!g20) & (!sk[24]) & (!g21) & (g98)) + ((!i_8_) & (!g30) & (!g20) & (!sk[24]) & (g21) & (g98)) + ((!i_8_) & (!g30) & (g20) & (!sk[24]) & (!g21) & (g98)) + ((!i_8_) & (!g30) & (g20) & (!sk[24]) & (g21) & (g98)) + ((!i_8_) & (g30) & (!g20) & (!sk[24]) & (!g21) & (g98)) + ((!i_8_) & (g30) & (!g20) & (!sk[24]) & (g21) & (g98)) + ((!i_8_) & (g30) & (!g20) & (sk[24]) & (g21) & (g98)) + ((!i_8_) & (g30) & (g20) & (!sk[24]) & (!g21) & (g98)) + ((!i_8_) & (g30) & (g20) & (!sk[24]) & (g21) & (g98)) + ((!i_8_) & (g30) & (g20) & (sk[24]) & (g21) & (g98)) + ((i_8_) & (!g30) & (!g20) & (!sk[24]) & (!g21) & (!g98)) + ((i_8_) & (!g30) & (!g20) & (!sk[24]) & (!g21) & (g98)) + ((i_8_) & (!g30) & (!g20) & (!sk[24]) & (g21) & (!g98)) + ((i_8_) & (!g30) & (!g20) & (!sk[24]) & (g21) & (g98)) + ((i_8_) & (!g30) & (g20) & (!sk[24]) & (!g21) & (!g98)) + ((i_8_) & (!g30) & (g20) & (!sk[24]) & (!g21) & (g98)) + ((i_8_) & (!g30) & (g20) & (!sk[24]) & (g21) & (!g98)) + ((i_8_) & (!g30) & (g20) & (!sk[24]) & (g21) & (g98)) + ((i_8_) & (g30) & (!g20) & (!sk[24]) & (!g21) & (!g98)) + ((i_8_) & (g30) & (!g20) & (!sk[24]) & (!g21) & (g98)) + ((i_8_) & (g30) & (!g20) & (!sk[24]) & (g21) & (!g98)) + ((i_8_) & (g30) & (!g20) & (!sk[24]) & (g21) & (g98)) + ((i_8_) & (g30) & (!g20) & (sk[24]) & (!g21) & (g98)) + ((i_8_) & (g30) & (!g20) & (sk[24]) & (g21) & (g98)) + ((i_8_) & (g30) & (g20) & (!sk[24]) & (!g21) & (!g98)) + ((i_8_) & (g30) & (g20) & (!sk[24]) & (!g21) & (g98)) + ((i_8_) & (g30) & (g20) & (!sk[24]) & (g21) & (!g98)) + ((i_8_) & (g30) & (g20) & (!sk[24]) & (g21) & (g98)));
	assign g263 = (((!g99) & (!g251) & (!g259) & (!g260) & (!g261) & (!g262)) + ((!g99) & (!g251) & (g259) & (!g260) & (!g261) & (!g262)) + ((!g99) & (g251) & (g259) & (!g260) & (!g261) & (!g262)) + ((g99) & (!g251) & (g259) & (!g260) & (!g261) & (!g262)) + ((g99) & (g251) & (g259) & (!g260) & (!g261) & (!g262)));
	assign g264 = (((!sk[26]) & (g13) & (!g102)) + ((!sk[26]) & (g13) & (g102)) + ((sk[26]) & (g13) & (!g102)));
	assign g265 = (((!g185) & (!g216) & (g120) & (!sk[27]) & (g173)) + ((!g185) & (g216) & (!g120) & (!sk[27]) & (!g173)) + ((!g185) & (g216) & (!g120) & (!sk[27]) & (g173)) + ((!g185) & (g216) & (g120) & (!sk[27]) & (!g173)) + ((!g185) & (g216) & (g120) & (!sk[27]) & (g173)) + ((g185) & (!g216) & (g120) & (!sk[27]) & (!g173)) + ((g185) & (!g216) & (g120) & (!sk[27]) & (g173)) + ((g185) & (!g216) & (g120) & (sk[27]) & (!g173)) + ((g185) & (g216) & (!g120) & (!sk[27]) & (!g173)) + ((g185) & (g216) & (!g120) & (!sk[27]) & (g173)) + ((g185) & (g216) & (g120) & (!sk[27]) & (!g173)) + ((g185) & (g216) & (g120) & (!sk[27]) & (g173)));
	assign g266 = (((!sk[28]) & (!i_8_) & (!g4) & (!g98) & (!g221) & (g185)) + ((!sk[28]) & (!i_8_) & (!g4) & (!g98) & (g221) & (g185)) + ((!sk[28]) & (!i_8_) & (!g4) & (g98) & (!g221) & (g185)) + ((!sk[28]) & (!i_8_) & (!g4) & (g98) & (g221) & (g185)) + ((!sk[28]) & (!i_8_) & (g4) & (!g98) & (!g221) & (g185)) + ((!sk[28]) & (!i_8_) & (g4) & (!g98) & (g221) & (g185)) + ((!sk[28]) & (!i_8_) & (g4) & (g98) & (!g221) & (g185)) + ((!sk[28]) & (!i_8_) & (g4) & (g98) & (g221) & (g185)) + ((!sk[28]) & (i_8_) & (!g4) & (!g98) & (!g221) & (!g185)) + ((!sk[28]) & (i_8_) & (!g4) & (!g98) & (!g221) & (g185)) + ((!sk[28]) & (i_8_) & (!g4) & (!g98) & (g221) & (!g185)) + ((!sk[28]) & (i_8_) & (!g4) & (!g98) & (g221) & (g185)) + ((!sk[28]) & (i_8_) & (!g4) & (g98) & (!g221) & (!g185)) + ((!sk[28]) & (i_8_) & (!g4) & (g98) & (!g221) & (g185)) + ((!sk[28]) & (i_8_) & (!g4) & (g98) & (g221) & (!g185)) + ((!sk[28]) & (i_8_) & (!g4) & (g98) & (g221) & (g185)) + ((!sk[28]) & (i_8_) & (g4) & (!g98) & (!g221) & (!g185)) + ((!sk[28]) & (i_8_) & (g4) & (!g98) & (!g221) & (g185)) + ((!sk[28]) & (i_8_) & (g4) & (!g98) & (g221) & (!g185)) + ((!sk[28]) & (i_8_) & (g4) & (!g98) & (g221) & (g185)) + ((!sk[28]) & (i_8_) & (g4) & (g98) & (!g221) & (!g185)) + ((!sk[28]) & (i_8_) & (g4) & (g98) & (!g221) & (g185)) + ((!sk[28]) & (i_8_) & (g4) & (g98) & (g221) & (!g185)) + ((!sk[28]) & (i_8_) & (g4) & (g98) & (g221) & (g185)) + ((sk[28]) & (!i_8_) & (g4) & (g98) & (!g221) & (!g185)) + ((sk[28]) & (!i_8_) & (g4) & (g98) & (g221) & (!g185)) + ((sk[28]) & (i_8_) & (g4) & (g98) & (!g221) & (!g185)) + ((sk[28]) & (i_8_) & (g4) & (g98) & (!g221) & (g185)));
	assign g267 = (((!g264) & (!g101) & (!g199) & (!g265) & (!g103) & (!g266)) + ((!g264) & (!g101) & (!g199) & (!g265) & (g103) & (!g266)) + ((!g264) & (!g101) & (!g199) & (g265) & (!g103) & (!g266)) + ((!g264) & (!g101) & (!g199) & (g265) & (g103) & (!g266)) + ((!g264) & (!g101) & (g199) & (!g265) & (!g103) & (!g266)) + ((!g264) & (!g101) & (g199) & (!g265) & (g103) & (!g266)) + ((!g264) & (!g101) & (g199) & (g265) & (!g103) & (!g266)) + ((!g264) & (!g101) & (g199) & (g265) & (g103) & (!g266)) + ((!g264) & (g101) & (!g199) & (g265) & (g103) & (!g266)) + ((g264) & (!g101) & (!g199) & (!g265) & (!g103) & (!g266)) + ((g264) & (!g101) & (!g199) & (!g265) & (g103) & (!g266)) + ((g264) & (!g101) & (!g199) & (g265) & (!g103) & (!g266)) + ((g264) & (!g101) & (!g199) & (g265) & (g103) & (!g266)) + ((g264) & (!g101) & (g199) & (!g265) & (!g103) & (!g266)) + ((g264) & (!g101) & (g199) & (!g265) & (g103) & (!g266)) + ((g264) & (!g101) & (g199) & (g265) & (!g103) & (!g266)) + ((g264) & (!g101) & (g199) & (g265) & (g103) & (!g266)));
	assign g268 = (((!sk[30]) & (g95) & (!g171)) + ((!sk[30]) & (g95) & (g171)) + ((sk[30]) & (g95) & (!g171)));
	assign g269 = (((!sk[31]) & (!i_14_) & (!i_12_) & (i_13_) & (g102)) + ((!sk[31]) & (!i_14_) & (i_12_) & (!i_13_) & (!g102)) + ((!sk[31]) & (!i_14_) & (i_12_) & (!i_13_) & (g102)) + ((!sk[31]) & (!i_14_) & (i_12_) & (i_13_) & (!g102)) + ((!sk[31]) & (!i_14_) & (i_12_) & (i_13_) & (g102)) + ((!sk[31]) & (i_14_) & (!i_12_) & (i_13_) & (!g102)) + ((!sk[31]) & (i_14_) & (!i_12_) & (i_13_) & (g102)) + ((!sk[31]) & (i_14_) & (i_12_) & (!i_13_) & (!g102)) + ((!sk[31]) & (i_14_) & (i_12_) & (!i_13_) & (g102)) + ((!sk[31]) & (i_14_) & (i_12_) & (i_13_) & (!g102)) + ((!sk[31]) & (i_14_) & (i_12_) & (i_13_) & (g102)) + ((sk[31]) & (i_14_) & (!i_12_) & (!i_13_) & (!g102)) + ((sk[31]) & (i_14_) & (!i_12_) & (i_13_) & (!g102)) + ((sk[31]) & (i_14_) & (i_12_) & (i_13_) & (!g102)));
	assign g270 = (((!g91) & (sk[32]) & (!g95)) + ((g91) & (!sk[32]) & (!g95)) + ((g91) & (!sk[32]) & (g95)) + ((g91) & (sk[32]) & (!g95)) + ((g91) & (sk[32]) & (g95)));
	assign g271 = (((!i_8_) & (!g4) & (!g98) & (!sk[33]) & (!g270) & (g255)) + ((!i_8_) & (!g4) & (!g98) & (!sk[33]) & (g270) & (g255)) + ((!i_8_) & (!g4) & (g98) & (!sk[33]) & (!g270) & (g255)) + ((!i_8_) & (!g4) & (g98) & (!sk[33]) & (g270) & (g255)) + ((!i_8_) & (g4) & (!g98) & (!sk[33]) & (!g270) & (g255)) + ((!i_8_) & (g4) & (!g98) & (!sk[33]) & (g270) & (g255)) + ((!i_8_) & (g4) & (g98) & (!sk[33]) & (!g270) & (g255)) + ((!i_8_) & (g4) & (g98) & (!sk[33]) & (g270) & (g255)) + ((!i_8_) & (g4) & (g98) & (sk[33]) & (!g270) & (!g255)) + ((!i_8_) & (g4) & (g98) & (sk[33]) & (!g270) & (g255)) + ((i_8_) & (!g4) & (!g98) & (!sk[33]) & (!g270) & (!g255)) + ((i_8_) & (!g4) & (!g98) & (!sk[33]) & (!g270) & (g255)) + ((i_8_) & (!g4) & (!g98) & (!sk[33]) & (g270) & (!g255)) + ((i_8_) & (!g4) & (!g98) & (!sk[33]) & (g270) & (g255)) + ((i_8_) & (!g4) & (g98) & (!sk[33]) & (!g270) & (!g255)) + ((i_8_) & (!g4) & (g98) & (!sk[33]) & (!g270) & (g255)) + ((i_8_) & (!g4) & (g98) & (!sk[33]) & (g270) & (!g255)) + ((i_8_) & (!g4) & (g98) & (!sk[33]) & (g270) & (g255)) + ((i_8_) & (g4) & (!g98) & (!sk[33]) & (!g270) & (!g255)) + ((i_8_) & (g4) & (!g98) & (!sk[33]) & (!g270) & (g255)) + ((i_8_) & (g4) & (!g98) & (!sk[33]) & (g270) & (!g255)) + ((i_8_) & (g4) & (!g98) & (!sk[33]) & (g270) & (g255)) + ((i_8_) & (g4) & (g98) & (!sk[33]) & (!g270) & (!g255)) + ((i_8_) & (g4) & (g98) & (!sk[33]) & (!g270) & (g255)) + ((i_8_) & (g4) & (g98) & (!sk[33]) & (g270) & (!g255)) + ((i_8_) & (g4) & (g98) & (!sk[33]) & (g270) & (g255)) + ((i_8_) & (g4) & (g98) & (sk[33]) & (!g270) & (!g255)) + ((i_8_) & (g4) & (g98) & (sk[33]) & (!g270) & (g255)) + ((i_8_) & (g4) & (g98) & (sk[33]) & (g270) & (g255)));
	assign g272 = (((!g134) & (!sk[34]) & (!g118) & (!g201) & (!g209) & (g246)) + ((!g134) & (!sk[34]) & (!g118) & (!g201) & (g209) & (g246)) + ((!g134) & (!sk[34]) & (!g118) & (g201) & (!g209) & (g246)) + ((!g134) & (!sk[34]) & (!g118) & (g201) & (g209) & (g246)) + ((!g134) & (!sk[34]) & (g118) & (!g201) & (!g209) & (g246)) + ((!g134) & (!sk[34]) & (g118) & (!g201) & (g209) & (g246)) + ((!g134) & (!sk[34]) & (g118) & (g201) & (!g209) & (g246)) + ((!g134) & (!sk[34]) & (g118) & (g201) & (g209) & (g246)) + ((!g134) & (sk[34]) & (!g118) & (!g201) & (!g209) & (!g246)) + ((!g134) & (sk[34]) & (!g118) & (!g201) & (!g209) & (g246)) + ((!g134) & (sk[34]) & (!g118) & (!g201) & (g209) & (!g246)) + ((!g134) & (sk[34]) & (!g118) & (!g201) & (g209) & (g246)) + ((!g134) & (sk[34]) & (!g118) & (g201) & (!g209) & (!g246)) + ((!g134) & (sk[34]) & (!g118) & (g201) & (!g209) & (g246)) + ((!g134) & (sk[34]) & (!g118) & (g201) & (g209) & (!g246)) + ((!g134) & (sk[34]) & (!g118) & (g201) & (g209) & (g246)) + ((!g134) & (sk[34]) & (g118) & (g201) & (!g209) & (!g246)) + ((g134) & (!sk[34]) & (!g118) & (!g201) & (!g209) & (!g246)) + ((g134) & (!sk[34]) & (!g118) & (!g201) & (!g209) & (g246)) + ((g134) & (!sk[34]) & (!g118) & (!g201) & (g209) & (!g246)) + ((g134) & (!sk[34]) & (!g118) & (!g201) & (g209) & (g246)) + ((g134) & (!sk[34]) & (!g118) & (g201) & (!g209) & (!g246)) + ((g134) & (!sk[34]) & (!g118) & (g201) & (!g209) & (g246)) + ((g134) & (!sk[34]) & (!g118) & (g201) & (g209) & (!g246)) + ((g134) & (!sk[34]) & (!g118) & (g201) & (g209) & (g246)) + ((g134) & (!sk[34]) & (g118) & (!g201) & (!g209) & (!g246)) + ((g134) & (!sk[34]) & (g118) & (!g201) & (!g209) & (g246)) + ((g134) & (!sk[34]) & (g118) & (!g201) & (g209) & (!g246)) + ((g134) & (!sk[34]) & (g118) & (!g201) & (g209) & (g246)) + ((g134) & (!sk[34]) & (g118) & (g201) & (!g209) & (!g246)) + ((g134) & (!sk[34]) & (g118) & (g201) & (!g209) & (g246)) + ((g134) & (!sk[34]) & (g118) & (g201) & (g209) & (!g246)) + ((g134) & (!sk[34]) & (g118) & (g201) & (g209) & (g246)) + ((g134) & (sk[34]) & (!g118) & (g201) & (!g209) & (!g246)) + ((g134) & (sk[34]) & (!g118) & (g201) & (!g209) & (g246)) + ((g134) & (sk[34]) & (!g118) & (g201) & (g209) & (!g246)) + ((g134) & (sk[34]) & (!g118) & (g201) & (g209) & (g246)) + ((g134) & (sk[34]) & (g118) & (g201) & (!g209) & (!g246)));
	assign g273 = (((!g145) & (!g268) & (!g172) & (!g269) & (!g271) & (g272)) + ((!g145) & (!g268) & (!g172) & (g269) & (!g271) & (g272)) + ((!g145) & (!g268) & (g172) & (!g269) & (!g271) & (g272)) + ((!g145) & (!g268) & (g172) & (g269) & (!g271) & (g272)) + ((!g145) & (g268) & (!g172) & (!g269) & (!g271) & (g272)) + ((!g145) & (g268) & (!g172) & (g269) & (!g271) & (g272)) + ((!g145) & (g268) & (g172) & (!g269) & (!g271) & (g272)) + ((!g145) & (g268) & (g172) & (g269) & (!g271) & (g272)) + ((g145) & (!g268) & (!g172) & (!g269) & (!g271) & (g272)));
	assign g274 = (((g242) & (!g250) & (g258) & (g263) & (g267) & (g273)));
	assign g275 = (((g235) & (!sk[37]) & (!g274)) + ((g235) & (!sk[37]) & (g274)) + ((g235) & (sk[37]) & (g274)));
	assign g276 = (((!g17) & (!g75) & (!sk[38]) & (g76) & (g1544)) + ((!g17) & (!g75) & (sk[38]) & (!g76) & (g1544)) + ((!g17) & (g75) & (!sk[38]) & (!g76) & (!g1544)) + ((!g17) & (g75) & (!sk[38]) & (!g76) & (g1544)) + ((!g17) & (g75) & (!sk[38]) & (g76) & (!g1544)) + ((!g17) & (g75) & (!sk[38]) & (g76) & (g1544)) + ((g17) & (!g75) & (!sk[38]) & (g76) & (!g1544)) + ((g17) & (!g75) & (!sk[38]) & (g76) & (g1544)) + ((g17) & (!g75) & (sk[38]) & (!g76) & (g1544)) + ((g17) & (g75) & (!sk[38]) & (!g76) & (!g1544)) + ((g17) & (g75) & (!sk[38]) & (!g76) & (g1544)) + ((g17) & (g75) & (!sk[38]) & (g76) & (!g1544)) + ((g17) & (g75) & (!sk[38]) & (g76) & (g1544)) + ((g17) & (g75) & (sk[38]) & (!g76) & (g1544)));
	assign g277 = (((!g134) & (sk[39]) & (!g118)) + ((g134) & (!sk[39]) & (!g118)) + ((g134) & (!sk[39]) & (g118)));
	assign g278 = (((!sk[40]) & (g191) & (!g277) & (!g214)) + ((!sk[40]) & (g191) & (!g277) & (g214)) + ((!sk[40]) & (g191) & (g277) & (!g214)) + ((!sk[40]) & (g191) & (g277) & (g214)) + ((sk[40]) & (g191) & (!g277) & (!g214)) + ((sk[40]) & (g191) & (!g277) & (g214)) + ((sk[40]) & (g191) & (g277) & (g214)));
	assign g279 = (((g131) & (!sk[41]) & (!g171)) + ((g131) & (!sk[41]) & (g171)) + ((g131) & (sk[41]) & (!g171)));
	assign g280 = (((i_9_) & (!g53) & (!sk[42]) & (!g182)) + ((i_9_) & (!g53) & (!sk[42]) & (g182)) + ((i_9_) & (g53) & (!sk[42]) & (!g182)) + ((i_9_) & (g53) & (!sk[42]) & (g182)) + ((i_9_) & (g53) & (sk[42]) & (g182)));
	assign g281 = (((!g142) & (!g103) & (g114) & (!sk[43]) & (g105)) + ((!g142) & (g103) & (!g114) & (!sk[43]) & (!g105)) + ((!g142) & (g103) & (!g114) & (!sk[43]) & (g105)) + ((!g142) & (g103) & (!g114) & (sk[43]) & (!g105)) + ((!g142) & (g103) & (g114) & (!sk[43]) & (!g105)) + ((!g142) & (g103) & (g114) & (!sk[43]) & (g105)) + ((g142) & (!g103) & (g114) & (!sk[43]) & (!g105)) + ((g142) & (!g103) & (g114) & (!sk[43]) & (g105)) + ((g142) & (g103) & (!g114) & (!sk[43]) & (!g105)) + ((g142) & (g103) & (!g114) & (!sk[43]) & (g105)) + ((g142) & (g103) & (g114) & (!sk[43]) & (!g105)) + ((g142) & (g103) & (g114) & (!sk[43]) & (g105)));
	assign g282 = (((!i_8_) & (!g88) & (!g118) & (!g216) & (!g243) & (!g281)) + ((!i_8_) & (!g88) & (!g118) & (!g216) & (!g243) & (g281)) + ((!i_8_) & (!g88) & (!g118) & (!g216) & (g243) & (g281)) + ((!i_8_) & (!g88) & (!g118) & (g216) & (!g243) & (!g281)) + ((!i_8_) & (!g88) & (!g118) & (g216) & (!g243) & (g281)) + ((!i_8_) & (!g88) & (!g118) & (g216) & (g243) & (g281)) + ((!i_8_) & (!g88) & (g118) & (!g216) & (!g243) & (g281)) + ((!i_8_) & (!g88) & (g118) & (!g216) & (g243) & (g281)) + ((!i_8_) & (g88) & (!g118) & (!g216) & (!g243) & (g281)) + ((!i_8_) & (g88) & (!g118) & (!g216) & (g243) & (g281)) + ((!i_8_) & (g88) & (!g118) & (g216) & (!g243) & (g281)) + ((!i_8_) & (g88) & (!g118) & (g216) & (g243) & (g281)) + ((!i_8_) & (g88) & (g118) & (!g216) & (!g243) & (g281)) + ((!i_8_) & (g88) & (g118) & (!g216) & (g243) & (g281)) + ((i_8_) & (!g88) & (!g118) & (!g216) & (!g243) & (!g281)) + ((i_8_) & (!g88) & (!g118) & (!g216) & (!g243) & (g281)) + ((i_8_) & (!g88) & (!g118) & (!g216) & (g243) & (g281)) + ((i_8_) & (!g88) & (!g118) & (g216) & (!g243) & (!g281)) + ((i_8_) & (!g88) & (!g118) & (g216) & (!g243) & (g281)) + ((i_8_) & (!g88) & (!g118) & (g216) & (g243) & (g281)) + ((i_8_) & (!g88) & (g118) & (!g216) & (!g243) & (g281)) + ((i_8_) & (!g88) & (g118) & (!g216) & (g243) & (g281)) + ((i_8_) & (g88) & (!g118) & (!g216) & (!g243) & (!g281)) + ((i_8_) & (g88) & (!g118) & (!g216) & (!g243) & (g281)) + ((i_8_) & (g88) & (!g118) & (!g216) & (g243) & (g281)) + ((i_8_) & (g88) & (!g118) & (g216) & (!g243) & (!g281)) + ((i_8_) & (g88) & (!g118) & (g216) & (!g243) & (g281)) + ((i_8_) & (g88) & (!g118) & (g216) & (g243) & (g281)) + ((i_8_) & (g88) & (g118) & (!g216) & (!g243) & (g281)) + ((i_8_) & (g88) & (g118) & (!g216) & (g243) & (g281)));
	assign g283 = (((!g145) & (!sk[45]) & (!g279) & (!g214) & (!g280) & (g282)) + ((!g145) & (!sk[45]) & (!g279) & (!g214) & (g280) & (g282)) + ((!g145) & (!sk[45]) & (!g279) & (g214) & (!g280) & (g282)) + ((!g145) & (!sk[45]) & (!g279) & (g214) & (g280) & (g282)) + ((!g145) & (!sk[45]) & (g279) & (!g214) & (!g280) & (g282)) + ((!g145) & (!sk[45]) & (g279) & (!g214) & (g280) & (g282)) + ((!g145) & (!sk[45]) & (g279) & (g214) & (!g280) & (g282)) + ((!g145) & (!sk[45]) & (g279) & (g214) & (g280) & (g282)) + ((!g145) & (sk[45]) & (!g279) & (!g214) & (!g280) & (g282)) + ((!g145) & (sk[45]) & (!g279) & (!g214) & (g280) & (g282)) + ((!g145) & (sk[45]) & (!g279) & (g214) & (!g280) & (g282)) + ((!g145) & (sk[45]) & (g279) & (!g214) & (!g280) & (g282)) + ((!g145) & (sk[45]) & (g279) & (!g214) & (g280) & (g282)) + ((!g145) & (sk[45]) & (g279) & (g214) & (!g280) & (g282)) + ((g145) & (!sk[45]) & (!g279) & (!g214) & (!g280) & (!g282)) + ((g145) & (!sk[45]) & (!g279) & (!g214) & (!g280) & (g282)) + ((g145) & (!sk[45]) & (!g279) & (!g214) & (g280) & (!g282)) + ((g145) & (!sk[45]) & (!g279) & (!g214) & (g280) & (g282)) + ((g145) & (!sk[45]) & (!g279) & (g214) & (!g280) & (!g282)) + ((g145) & (!sk[45]) & (!g279) & (g214) & (!g280) & (g282)) + ((g145) & (!sk[45]) & (!g279) & (g214) & (g280) & (!g282)) + ((g145) & (!sk[45]) & (!g279) & (g214) & (g280) & (g282)) + ((g145) & (!sk[45]) & (g279) & (!g214) & (!g280) & (!g282)) + ((g145) & (!sk[45]) & (g279) & (!g214) & (!g280) & (g282)) + ((g145) & (!sk[45]) & (g279) & (!g214) & (g280) & (!g282)) + ((g145) & (!sk[45]) & (g279) & (!g214) & (g280) & (g282)) + ((g145) & (!sk[45]) & (g279) & (g214) & (!g280) & (!g282)) + ((g145) & (!sk[45]) & (g279) & (g214) & (!g280) & (g282)) + ((g145) & (!sk[45]) & (g279) & (g214) & (g280) & (!g282)) + ((g145) & (!sk[45]) & (g279) & (g214) & (g280) & (g282)) + ((g145) & (sk[45]) & (!g279) & (!g214) & (!g280) & (g282)) + ((g145) & (sk[45]) & (!g279) & (!g214) & (g280) & (g282)) + ((g145) & (sk[45]) & (!g279) & (g214) & (!g280) & (g282)));
	assign g284 = (((!sk[46]) & (i_8_) & (!g4) & (!g58)) + ((!sk[46]) & (i_8_) & (!g4) & (g58)) + ((!sk[46]) & (i_8_) & (g4) & (!g58)) + ((!sk[46]) & (i_8_) & (g4) & (g58)) + ((sk[46]) & (i_8_) & (g4) & (g58)));
	assign g285 = (((!i_8_) & (!g134) & (sk[47]) & (!g108)) + ((i_8_) & (!g134) & (!sk[47]) & (!g108)) + ((i_8_) & (!g134) & (!sk[47]) & (g108)) + ((i_8_) & (!g134) & (sk[47]) & (!g108)) + ((i_8_) & (!g134) & (sk[47]) & (g108)) + ((i_8_) & (g134) & (!sk[47]) & (!g108)) + ((i_8_) & (g134) & (!sk[47]) & (g108)));
	assign g286 = (((!g100) & (!g251) & (!g253) & (!g284) & (!g159) & (!g285)) + ((!g100) & (!g251) & (!g253) & (!g284) & (!g159) & (g285)) + ((!g100) & (!g251) & (!g253) & (!g284) & (g159) & (!g285)) + ((!g100) & (!g251) & (!g253) & (!g284) & (g159) & (g285)) + ((!g100) & (!g251) & (!g253) & (g284) & (!g159) & (!g285)) + ((!g100) & (!g251) & (!g253) & (g284) & (!g159) & (g285)) + ((!g100) & (!g251) & (g253) & (!g284) & (!g159) & (g285)) + ((!g100) & (!g251) & (g253) & (!g284) & (g159) & (g285)) + ((!g100) & (!g251) & (g253) & (g284) & (!g159) & (g285)) + ((!g100) & (g251) & (!g253) & (!g284) & (!g159) & (!g285)) + ((!g100) & (g251) & (!g253) & (!g284) & (!g159) & (g285)) + ((!g100) & (g251) & (!g253) & (g284) & (!g159) & (!g285)) + ((!g100) & (g251) & (!g253) & (g284) & (!g159) & (g285)) + ((!g100) & (g251) & (g253) & (!g284) & (!g159) & (g285)) + ((!g100) & (g251) & (g253) & (g284) & (!g159) & (g285)) + ((g100) & (!g251) & (!g253) & (!g284) & (!g159) & (!g285)) + ((g100) & (!g251) & (!g253) & (!g284) & (!g159) & (g285)) + ((g100) & (!g251) & (!g253) & (g284) & (!g159) & (!g285)) + ((g100) & (!g251) & (!g253) & (g284) & (!g159) & (g285)) + ((g100) & (!g251) & (g253) & (!g284) & (!g159) & (g285)) + ((g100) & (!g251) & (g253) & (g284) & (!g159) & (g285)) + ((g100) & (g251) & (!g253) & (!g284) & (!g159) & (!g285)) + ((g100) & (g251) & (!g253) & (!g284) & (!g159) & (g285)) + ((g100) & (g251) & (!g253) & (g284) & (!g159) & (!g285)) + ((g100) & (g251) & (!g253) & (g284) & (!g159) & (g285)) + ((g100) & (g251) & (g253) & (!g284) & (!g159) & (g285)) + ((g100) & (g251) & (g253) & (g284) & (!g159) & (g285)));
	assign g287 = (((!sk[49]) & (g99) & (!g94) & (!g116)) + ((!sk[49]) & (g99) & (!g94) & (g116)) + ((!sk[49]) & (g99) & (g94) & (!g116)) + ((!sk[49]) & (g99) & (g94) & (g116)) + ((sk[49]) & (g99) & (!g94) & (g116)) + ((sk[49]) & (g99) & (g94) & (!g116)) + ((sk[49]) & (g99) & (g94) & (g116)));
	assign g288 = (((!i_8_) & (!sk[50]) & (!i_6_) & (!i_7_) & (!g5) & (g40)) + ((!i_8_) & (!sk[50]) & (!i_6_) & (!i_7_) & (g5) & (g40)) + ((!i_8_) & (!sk[50]) & (!i_6_) & (i_7_) & (!g5) & (g40)) + ((!i_8_) & (!sk[50]) & (!i_6_) & (i_7_) & (g5) & (g40)) + ((!i_8_) & (!sk[50]) & (i_6_) & (!i_7_) & (!g5) & (g40)) + ((!i_8_) & (!sk[50]) & (i_6_) & (!i_7_) & (g5) & (g40)) + ((!i_8_) & (!sk[50]) & (i_6_) & (i_7_) & (!g5) & (g40)) + ((!i_8_) & (!sk[50]) & (i_6_) & (i_7_) & (g5) & (g40)) + ((!i_8_) & (sk[50]) & (i_6_) & (!i_7_) & (g5) & (g40)) + ((i_8_) & (!sk[50]) & (!i_6_) & (!i_7_) & (!g5) & (!g40)) + ((i_8_) & (!sk[50]) & (!i_6_) & (!i_7_) & (!g5) & (g40)) + ((i_8_) & (!sk[50]) & (!i_6_) & (!i_7_) & (g5) & (!g40)) + ((i_8_) & (!sk[50]) & (!i_6_) & (!i_7_) & (g5) & (g40)) + ((i_8_) & (!sk[50]) & (!i_6_) & (i_7_) & (!g5) & (!g40)) + ((i_8_) & (!sk[50]) & (!i_6_) & (i_7_) & (!g5) & (g40)) + ((i_8_) & (!sk[50]) & (!i_6_) & (i_7_) & (g5) & (!g40)) + ((i_8_) & (!sk[50]) & (!i_6_) & (i_7_) & (g5) & (g40)) + ((i_8_) & (!sk[50]) & (i_6_) & (!i_7_) & (!g5) & (!g40)) + ((i_8_) & (!sk[50]) & (i_6_) & (!i_7_) & (!g5) & (g40)) + ((i_8_) & (!sk[50]) & (i_6_) & (!i_7_) & (g5) & (!g40)) + ((i_8_) & (!sk[50]) & (i_6_) & (!i_7_) & (g5) & (g40)) + ((i_8_) & (!sk[50]) & (i_6_) & (i_7_) & (!g5) & (!g40)) + ((i_8_) & (!sk[50]) & (i_6_) & (i_7_) & (!g5) & (g40)) + ((i_8_) & (!sk[50]) & (i_6_) & (i_7_) & (g5) & (!g40)) + ((i_8_) & (!sk[50]) & (i_6_) & (i_7_) & (g5) & (g40)) + ((i_8_) & (sk[50]) & (i_6_) & (!i_7_) & (!g5) & (g40)) + ((i_8_) & (sk[50]) & (i_6_) & (!i_7_) & (g5) & (g40)));
	assign g289 = (((i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!g91) & (!g100)) + ((i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!g91) & (g100)) + ((i_11_) & (i_9_) & (i_10_) & (i_15_) & (!g91) & (g100)));
	assign g290 = (((!i_8_) & (!g4) & (!g98) & (!sk[52]) & (!g92) & (g165)) + ((!i_8_) & (!g4) & (!g98) & (!sk[52]) & (g92) & (g165)) + ((!i_8_) & (!g4) & (g98) & (!sk[52]) & (!g92) & (g165)) + ((!i_8_) & (!g4) & (g98) & (!sk[52]) & (g92) & (g165)) + ((!i_8_) & (g4) & (!g98) & (!sk[52]) & (!g92) & (g165)) + ((!i_8_) & (g4) & (!g98) & (!sk[52]) & (g92) & (g165)) + ((!i_8_) & (g4) & (g98) & (!sk[52]) & (!g92) & (g165)) + ((!i_8_) & (g4) & (g98) & (!sk[52]) & (g92) & (g165)) + ((!i_8_) & (g4) & (g98) & (sk[52]) & (!g92) & (!g165)) + ((!i_8_) & (g4) & (g98) & (sk[52]) & (!g92) & (g165)) + ((i_8_) & (!g4) & (!g98) & (!sk[52]) & (!g92) & (!g165)) + ((i_8_) & (!g4) & (!g98) & (!sk[52]) & (!g92) & (g165)) + ((i_8_) & (!g4) & (!g98) & (!sk[52]) & (g92) & (!g165)) + ((i_8_) & (!g4) & (!g98) & (!sk[52]) & (g92) & (g165)) + ((i_8_) & (!g4) & (g98) & (!sk[52]) & (!g92) & (!g165)) + ((i_8_) & (!g4) & (g98) & (!sk[52]) & (!g92) & (g165)) + ((i_8_) & (!g4) & (g98) & (!sk[52]) & (g92) & (!g165)) + ((i_8_) & (!g4) & (g98) & (!sk[52]) & (g92) & (g165)) + ((i_8_) & (g4) & (!g98) & (!sk[52]) & (!g92) & (!g165)) + ((i_8_) & (g4) & (!g98) & (!sk[52]) & (!g92) & (g165)) + ((i_8_) & (g4) & (!g98) & (!sk[52]) & (g92) & (!g165)) + ((i_8_) & (g4) & (!g98) & (!sk[52]) & (g92) & (g165)) + ((i_8_) & (g4) & (g98) & (!sk[52]) & (!g92) & (!g165)) + ((i_8_) & (g4) & (g98) & (!sk[52]) & (!g92) & (g165)) + ((i_8_) & (g4) & (g98) & (!sk[52]) & (g92) & (!g165)) + ((i_8_) & (g4) & (g98) & (!sk[52]) & (g92) & (g165)) + ((i_8_) & (g4) & (g98) & (sk[52]) & (!g92) & (!g165)) + ((i_8_) & (g4) & (g98) & (sk[52]) & (!g92) & (g165)) + ((i_8_) & (g4) & (g98) & (sk[52]) & (g92) & (g165)));
	assign g291 = (((!g100) & (!g251) & (!g287) & (!g288) & (!g289) & (!g290)) + ((!g100) & (!g251) & (!g287) & (!g288) & (g289) & (!g290)) + ((!g100) & (g251) & (!g287) & (!g288) & (!g289) & (!g290)) + ((g100) & (!g251) & (!g287) & (!g288) & (!g289) & (!g290)) + ((g100) & (g251) & (!g287) & (!g288) & (!g289) & (!g290)));
	assign g292 = (((!sk[54]) & (!g127) & (!g90) & (g116) & (g125)) + ((!sk[54]) & (!g127) & (g90) & (!g116) & (!g125)) + ((!sk[54]) & (!g127) & (g90) & (!g116) & (g125)) + ((!sk[54]) & (!g127) & (g90) & (g116) & (!g125)) + ((!sk[54]) & (!g127) & (g90) & (g116) & (g125)) + ((!sk[54]) & (g127) & (!g90) & (g116) & (!g125)) + ((!sk[54]) & (g127) & (!g90) & (g116) & (g125)) + ((!sk[54]) & (g127) & (g90) & (!g116) & (!g125)) + ((!sk[54]) & (g127) & (g90) & (!g116) & (g125)) + ((!sk[54]) & (g127) & (g90) & (g116) & (!g125)) + ((!sk[54]) & (g127) & (g90) & (g116) & (g125)) + ((sk[54]) & (g127) & (g90) & (!g116) & (!g125)));
	assign g293 = (((!i_8_) & (!g48) & (!g91) & (!g95) & (!sk[55]) & (g216)) + ((!i_8_) & (!g48) & (!g91) & (!g95) & (sk[55]) & (!g216)) + ((!i_8_) & (!g48) & (!g91) & (g95) & (!sk[55]) & (g216)) + ((!i_8_) & (!g48) & (g91) & (!g95) & (!sk[55]) & (g216)) + ((!i_8_) & (!g48) & (g91) & (!g95) & (sk[55]) & (!g216)) + ((!i_8_) & (!g48) & (g91) & (g95) & (!sk[55]) & (g216)) + ((!i_8_) & (g48) & (!g91) & (!g95) & (!sk[55]) & (g216)) + ((!i_8_) & (g48) & (!g91) & (!g95) & (sk[55]) & (!g216)) + ((!i_8_) & (g48) & (!g91) & (g95) & (!sk[55]) & (g216)) + ((!i_8_) & (g48) & (g91) & (!g95) & (!sk[55]) & (g216)) + ((!i_8_) & (g48) & (g91) & (!g95) & (sk[55]) & (!g216)) + ((!i_8_) & (g48) & (g91) & (g95) & (!sk[55]) & (g216)) + ((!i_8_) & (g48) & (g91) & (g95) & (sk[55]) & (!g216)) + ((i_8_) & (!g48) & (!g91) & (!g95) & (!sk[55]) & (!g216)) + ((i_8_) & (!g48) & (!g91) & (!g95) & (!sk[55]) & (g216)) + ((i_8_) & (!g48) & (!g91) & (!g95) & (sk[55]) & (!g216)) + ((i_8_) & (!g48) & (!g91) & (g95) & (!sk[55]) & (!g216)) + ((i_8_) & (!g48) & (!g91) & (g95) & (!sk[55]) & (g216)) + ((i_8_) & (!g48) & (!g91) & (g95) & (sk[55]) & (!g216)) + ((i_8_) & (!g48) & (g91) & (!g95) & (!sk[55]) & (!g216)) + ((i_8_) & (!g48) & (g91) & (!g95) & (!sk[55]) & (g216)) + ((i_8_) & (!g48) & (g91) & (!g95) & (sk[55]) & (!g216)) + ((i_8_) & (!g48) & (g91) & (g95) & (!sk[55]) & (!g216)) + ((i_8_) & (!g48) & (g91) & (g95) & (!sk[55]) & (g216)) + ((i_8_) & (!g48) & (g91) & (g95) & (sk[55]) & (!g216)) + ((i_8_) & (g48) & (!g91) & (!g95) & (!sk[55]) & (!g216)) + ((i_8_) & (g48) & (!g91) & (!g95) & (!sk[55]) & (g216)) + ((i_8_) & (g48) & (!g91) & (!g95) & (sk[55]) & (!g216)) + ((i_8_) & (g48) & (!g91) & (g95) & (!sk[55]) & (!g216)) + ((i_8_) & (g48) & (!g91) & (g95) & (!sk[55]) & (g216)) + ((i_8_) & (g48) & (!g91) & (g95) & (sk[55]) & (!g216)) + ((i_8_) & (g48) & (g91) & (!g95) & (!sk[55]) & (!g216)) + ((i_8_) & (g48) & (g91) & (!g95) & (!sk[55]) & (g216)) + ((i_8_) & (g48) & (g91) & (!g95) & (sk[55]) & (!g216)) + ((i_8_) & (g48) & (g91) & (g95) & (!sk[55]) & (!g216)) + ((i_8_) & (g48) & (g91) & (g95) & (!sk[55]) & (g216)) + ((i_8_) & (g48) & (g91) & (g95) & (sk[55]) & (!g216)));
	assign g294 = (((!i_11_) & (!i_9_) & (!sk[56]) & (!i_10_) & (!i_15_) & (g91)) + ((!i_11_) & (!i_9_) & (!sk[56]) & (!i_10_) & (i_15_) & (g91)) + ((!i_11_) & (!i_9_) & (!sk[56]) & (i_10_) & (!i_15_) & (g91)) + ((!i_11_) & (!i_9_) & (!sk[56]) & (i_10_) & (i_15_) & (g91)) + ((!i_11_) & (!i_9_) & (sk[56]) & (i_10_) & (i_15_) & (!g91)) + ((!i_11_) & (i_9_) & (!sk[56]) & (!i_10_) & (!i_15_) & (g91)) + ((!i_11_) & (i_9_) & (!sk[56]) & (!i_10_) & (i_15_) & (g91)) + ((!i_11_) & (i_9_) & (!sk[56]) & (i_10_) & (!i_15_) & (g91)) + ((!i_11_) & (i_9_) & (!sk[56]) & (i_10_) & (i_15_) & (g91)) + ((!i_11_) & (i_9_) & (sk[56]) & (!i_10_) & (i_15_) & (!g91)) + ((i_11_) & (!i_9_) & (!sk[56]) & (!i_10_) & (!i_15_) & (!g91)) + ((i_11_) & (!i_9_) & (!sk[56]) & (!i_10_) & (!i_15_) & (g91)) + ((i_11_) & (!i_9_) & (!sk[56]) & (!i_10_) & (i_15_) & (!g91)) + ((i_11_) & (!i_9_) & (!sk[56]) & (!i_10_) & (i_15_) & (g91)) + ((i_11_) & (!i_9_) & (!sk[56]) & (i_10_) & (!i_15_) & (!g91)) + ((i_11_) & (!i_9_) & (!sk[56]) & (i_10_) & (!i_15_) & (g91)) + ((i_11_) & (!i_9_) & (!sk[56]) & (i_10_) & (i_15_) & (!g91)) + ((i_11_) & (!i_9_) & (!sk[56]) & (i_10_) & (i_15_) & (g91)) + ((i_11_) & (!i_9_) & (sk[56]) & (!i_10_) & (i_15_) & (!g91)) + ((i_11_) & (i_9_) & (!sk[56]) & (!i_10_) & (!i_15_) & (!g91)) + ((i_11_) & (i_9_) & (!sk[56]) & (!i_10_) & (!i_15_) & (g91)) + ((i_11_) & (i_9_) & (!sk[56]) & (!i_10_) & (i_15_) & (!g91)) + ((i_11_) & (i_9_) & (!sk[56]) & (!i_10_) & (i_15_) & (g91)) + ((i_11_) & (i_9_) & (!sk[56]) & (i_10_) & (!i_15_) & (!g91)) + ((i_11_) & (i_9_) & (!sk[56]) & (i_10_) & (!i_15_) & (g91)) + ((i_11_) & (i_9_) & (!sk[56]) & (i_10_) & (i_15_) & (!g91)) + ((i_11_) & (i_9_) & (!sk[56]) & (i_10_) & (i_15_) & (g91)));
	assign g295 = (((!sk[57]) & (!g59) & (!g243) & (!g292) & (!g293) & (g294)) + ((!sk[57]) & (!g59) & (!g243) & (!g292) & (g293) & (g294)) + ((!sk[57]) & (!g59) & (!g243) & (g292) & (!g293) & (g294)) + ((!sk[57]) & (!g59) & (!g243) & (g292) & (g293) & (g294)) + ((!sk[57]) & (!g59) & (g243) & (!g292) & (!g293) & (g294)) + ((!sk[57]) & (!g59) & (g243) & (!g292) & (g293) & (g294)) + ((!sk[57]) & (!g59) & (g243) & (g292) & (!g293) & (g294)) + ((!sk[57]) & (!g59) & (g243) & (g292) & (g293) & (g294)) + ((!sk[57]) & (g59) & (!g243) & (!g292) & (!g293) & (!g294)) + ((!sk[57]) & (g59) & (!g243) & (!g292) & (!g293) & (g294)) + ((!sk[57]) & (g59) & (!g243) & (!g292) & (g293) & (!g294)) + ((!sk[57]) & (g59) & (!g243) & (!g292) & (g293) & (g294)) + ((!sk[57]) & (g59) & (!g243) & (g292) & (!g293) & (!g294)) + ((!sk[57]) & (g59) & (!g243) & (g292) & (!g293) & (g294)) + ((!sk[57]) & (g59) & (!g243) & (g292) & (g293) & (!g294)) + ((!sk[57]) & (g59) & (!g243) & (g292) & (g293) & (g294)) + ((!sk[57]) & (g59) & (g243) & (!g292) & (!g293) & (!g294)) + ((!sk[57]) & (g59) & (g243) & (!g292) & (!g293) & (g294)) + ((!sk[57]) & (g59) & (g243) & (!g292) & (g293) & (!g294)) + ((!sk[57]) & (g59) & (g243) & (!g292) & (g293) & (g294)) + ((!sk[57]) & (g59) & (g243) & (g292) & (!g293) & (!g294)) + ((!sk[57]) & (g59) & (g243) & (g292) & (!g293) & (g294)) + ((!sk[57]) & (g59) & (g243) & (g292) & (g293) & (!g294)) + ((!sk[57]) & (g59) & (g243) & (g292) & (g293) & (g294)) + ((sk[57]) & (!g59) & (!g243) & (!g292) & (!g293) & (!g294)) + ((sk[57]) & (!g59) & (!g243) & (!g292) & (!g293) & (g294)) + ((sk[57]) & (!g59) & (!g243) & (!g292) & (g293) & (!g294)) + ((sk[57]) & (!g59) & (!g243) & (!g292) & (g293) & (g294)) + ((sk[57]) & (!g59) & (!g243) & (g292) & (!g293) & (!g294)) + ((sk[57]) & (!g59) & (!g243) & (g292) & (!g293) & (g294)) + ((sk[57]) & (!g59) & (!g243) & (g292) & (g293) & (!g294)) + ((sk[57]) & (!g59) & (!g243) & (g292) & (g293) & (g294)) + ((sk[57]) & (!g59) & (g243) & (g292) & (g293) & (!g294)) + ((sk[57]) & (g59) & (!g243) & (!g292) & (!g293) & (!g294)) + ((sk[57]) & (g59) & (!g243) & (!g292) & (g293) & (!g294)) + ((sk[57]) & (g59) & (!g243) & (g292) & (!g293) & (!g294)) + ((sk[57]) & (g59) & (!g243) & (g292) & (g293) & (!g294)) + ((sk[57]) & (g59) & (g243) & (g292) & (g293) & (!g294)));
	assign g296 = (((!g134) & (!g252) & (g283) & (g286) & (g291) & (g295)) + ((!g134) & (g252) & (g283) & (g286) & (g291) & (g295)) + ((g134) & (!g252) & (g283) & (g286) & (g291) & (g295)));
	assign g297 = (((!sk[59]) & (g13) & (!g104)) + ((!sk[59]) & (g13) & (g104)) + ((sk[59]) & (g13) & (g104)));
	assign g298 = (((!i_11_) & (!i_9_) & (!sk[60]) & (!i_10_) & (!g59) & (g244)) + ((!i_11_) & (!i_9_) & (!sk[60]) & (!i_10_) & (g59) & (g244)) + ((!i_11_) & (!i_9_) & (!sk[60]) & (i_10_) & (!g59) & (g244)) + ((!i_11_) & (!i_9_) & (!sk[60]) & (i_10_) & (g59) & (g244)) + ((!i_11_) & (!i_9_) & (sk[60]) & (i_10_) & (g59) & (g244)) + ((!i_11_) & (i_9_) & (!sk[60]) & (!i_10_) & (!g59) & (g244)) + ((!i_11_) & (i_9_) & (!sk[60]) & (!i_10_) & (g59) & (g244)) + ((!i_11_) & (i_9_) & (!sk[60]) & (i_10_) & (!g59) & (g244)) + ((!i_11_) & (i_9_) & (!sk[60]) & (i_10_) & (g59) & (g244)) + ((i_11_) & (!i_9_) & (!sk[60]) & (!i_10_) & (!g59) & (!g244)) + ((i_11_) & (!i_9_) & (!sk[60]) & (!i_10_) & (!g59) & (g244)) + ((i_11_) & (!i_9_) & (!sk[60]) & (!i_10_) & (g59) & (!g244)) + ((i_11_) & (!i_9_) & (!sk[60]) & (!i_10_) & (g59) & (g244)) + ((i_11_) & (!i_9_) & (!sk[60]) & (i_10_) & (!g59) & (!g244)) + ((i_11_) & (!i_9_) & (!sk[60]) & (i_10_) & (!g59) & (g244)) + ((i_11_) & (!i_9_) & (!sk[60]) & (i_10_) & (g59) & (!g244)) + ((i_11_) & (!i_9_) & (!sk[60]) & (i_10_) & (g59) & (g244)) + ((i_11_) & (!i_9_) & (sk[60]) & (!i_10_) & (g59) & (g244)) + ((i_11_) & (i_9_) & (!sk[60]) & (!i_10_) & (!g59) & (!g244)) + ((i_11_) & (i_9_) & (!sk[60]) & (!i_10_) & (!g59) & (g244)) + ((i_11_) & (i_9_) & (!sk[60]) & (!i_10_) & (g59) & (!g244)) + ((i_11_) & (i_9_) & (!sk[60]) & (!i_10_) & (g59) & (g244)) + ((i_11_) & (i_9_) & (!sk[60]) & (i_10_) & (!g59) & (!g244)) + ((i_11_) & (i_9_) & (!sk[60]) & (i_10_) & (!g59) & (g244)) + ((i_11_) & (i_9_) & (!sk[60]) & (i_10_) & (g59) & (!g244)) + ((i_11_) & (i_9_) & (!sk[60]) & (i_10_) & (g59) & (g244)));
	assign g299 = (((!i_8_) & (!g20) & (!g4) & (!sk[61]) & (!g98) & (g216)) + ((!i_8_) & (!g20) & (!g4) & (!sk[61]) & (g98) & (g216)) + ((!i_8_) & (!g20) & (g4) & (!sk[61]) & (!g98) & (g216)) + ((!i_8_) & (!g20) & (g4) & (!sk[61]) & (g98) & (g216)) + ((!i_8_) & (!g20) & (g4) & (sk[61]) & (g98) & (g216)) + ((!i_8_) & (g20) & (!g4) & (!sk[61]) & (!g98) & (g216)) + ((!i_8_) & (g20) & (!g4) & (!sk[61]) & (g98) & (g216)) + ((!i_8_) & (g20) & (g4) & (!sk[61]) & (!g98) & (g216)) + ((!i_8_) & (g20) & (g4) & (!sk[61]) & (g98) & (g216)) + ((!i_8_) & (g20) & (g4) & (sk[61]) & (g98) & (g216)) + ((i_8_) & (!g20) & (!g4) & (!sk[61]) & (!g98) & (!g216)) + ((i_8_) & (!g20) & (!g4) & (!sk[61]) & (!g98) & (g216)) + ((i_8_) & (!g20) & (!g4) & (!sk[61]) & (g98) & (!g216)) + ((i_8_) & (!g20) & (!g4) & (!sk[61]) & (g98) & (g216)) + ((i_8_) & (!g20) & (g4) & (!sk[61]) & (!g98) & (!g216)) + ((i_8_) & (!g20) & (g4) & (!sk[61]) & (!g98) & (g216)) + ((i_8_) & (!g20) & (g4) & (!sk[61]) & (g98) & (!g216)) + ((i_8_) & (!g20) & (g4) & (!sk[61]) & (g98) & (g216)) + ((i_8_) & (!g20) & (g4) & (sk[61]) & (g98) & (!g216)) + ((i_8_) & (!g20) & (g4) & (sk[61]) & (g98) & (g216)) + ((i_8_) & (g20) & (!g4) & (!sk[61]) & (!g98) & (!g216)) + ((i_8_) & (g20) & (!g4) & (!sk[61]) & (!g98) & (g216)) + ((i_8_) & (g20) & (!g4) & (!sk[61]) & (g98) & (!g216)) + ((i_8_) & (g20) & (!g4) & (!sk[61]) & (g98) & (g216)) + ((i_8_) & (g20) & (g4) & (!sk[61]) & (!g98) & (!g216)) + ((i_8_) & (g20) & (g4) & (!sk[61]) & (!g98) & (g216)) + ((i_8_) & (g20) & (g4) & (!sk[61]) & (g98) & (!g216)) + ((i_8_) & (g20) & (g4) & (!sk[61]) & (g98) & (g216)));
	assign g300 = (((!g14) & (!g4) & (!g98) & (!g118) & (!sk[62]) & (g299)) + ((!g14) & (!g4) & (!g98) & (!g118) & (sk[62]) & (!g299)) + ((!g14) & (!g4) & (!g98) & (g118) & (!sk[62]) & (g299)) + ((!g14) & (!g4) & (!g98) & (g118) & (sk[62]) & (!g299)) + ((!g14) & (!g4) & (g98) & (!g118) & (!sk[62]) & (g299)) + ((!g14) & (!g4) & (g98) & (!g118) & (sk[62]) & (!g299)) + ((!g14) & (!g4) & (g98) & (g118) & (!sk[62]) & (g299)) + ((!g14) & (!g4) & (g98) & (g118) & (sk[62]) & (!g299)) + ((!g14) & (g4) & (!g98) & (!g118) & (!sk[62]) & (g299)) + ((!g14) & (g4) & (!g98) & (!g118) & (sk[62]) & (!g299)) + ((!g14) & (g4) & (!g98) & (g118) & (!sk[62]) & (g299)) + ((!g14) & (g4) & (!g98) & (g118) & (sk[62]) & (!g299)) + ((!g14) & (g4) & (g98) & (!g118) & (!sk[62]) & (g299)) + ((!g14) & (g4) & (g98) & (!g118) & (sk[62]) & (!g299)) + ((!g14) & (g4) & (g98) & (g118) & (!sk[62]) & (g299)) + ((!g14) & (g4) & (g98) & (g118) & (sk[62]) & (!g299)) + ((g14) & (!g4) & (!g98) & (!g118) & (!sk[62]) & (!g299)) + ((g14) & (!g4) & (!g98) & (!g118) & (!sk[62]) & (g299)) + ((g14) & (!g4) & (!g98) & (!g118) & (sk[62]) & (!g299)) + ((g14) & (!g4) & (!g98) & (g118) & (!sk[62]) & (!g299)) + ((g14) & (!g4) & (!g98) & (g118) & (!sk[62]) & (g299)) + ((g14) & (!g4) & (g98) & (!g118) & (!sk[62]) & (!g299)) + ((g14) & (!g4) & (g98) & (!g118) & (!sk[62]) & (g299)) + ((g14) & (!g4) & (g98) & (!g118) & (sk[62]) & (!g299)) + ((g14) & (!g4) & (g98) & (g118) & (!sk[62]) & (!g299)) + ((g14) & (!g4) & (g98) & (g118) & (!sk[62]) & (g299)) + ((g14) & (g4) & (!g98) & (!g118) & (!sk[62]) & (!g299)) + ((g14) & (g4) & (!g98) & (!g118) & (!sk[62]) & (g299)) + ((g14) & (g4) & (!g98) & (!g118) & (sk[62]) & (!g299)) + ((g14) & (g4) & (!g98) & (g118) & (!sk[62]) & (!g299)) + ((g14) & (g4) & (!g98) & (g118) & (!sk[62]) & (g299)) + ((g14) & (g4) & (g98) & (!g118) & (!sk[62]) & (!g299)) + ((g14) & (g4) & (g98) & (!g118) & (!sk[62]) & (g299)) + ((g14) & (g4) & (g98) & (g118) & (!sk[62]) & (!g299)) + ((g14) & (g4) & (g98) & (g118) & (!sk[62]) & (g299)));
	assign g301 = (((!g297) & (!g89) & (!g245) & (!g136) & (!g298) & (g300)) + ((!g297) & (!g89) & (!g245) & (g136) & (!g298) & (g300)) + ((!g297) & (g89) & (!g245) & (!g136) & (!g298) & (g300)) + ((!g297) & (g89) & (!g245) & (g136) & (!g298) & (g300)) + ((!g297) & (g89) & (g245) & (!g136) & (!g298) & (g300)) + ((!g297) & (g89) & (g245) & (g136) & (!g298) & (g300)) + ((g297) & (!g89) & (!g245) & (!g136) & (!g298) & (g300)) + ((g297) & (g89) & (!g245) & (!g136) & (!g298) & (g300)) + ((g297) & (g89) & (g245) & (!g136) & (!g298) & (g300)));
	assign g302 = (((!sk[64]) & (!i_8_) & (!g220) & (g264) & (g135)) + ((!sk[64]) & (!i_8_) & (g220) & (!g264) & (!g135)) + ((!sk[64]) & (!i_8_) & (g220) & (!g264) & (g135)) + ((!sk[64]) & (!i_8_) & (g220) & (g264) & (!g135)) + ((!sk[64]) & (!i_8_) & (g220) & (g264) & (g135)) + ((!sk[64]) & (i_8_) & (!g220) & (g264) & (!g135)) + ((!sk[64]) & (i_8_) & (!g220) & (g264) & (g135)) + ((!sk[64]) & (i_8_) & (g220) & (!g264) & (!g135)) + ((!sk[64]) & (i_8_) & (g220) & (!g264) & (g135)) + ((!sk[64]) & (i_8_) & (g220) & (g264) & (!g135)) + ((!sk[64]) & (i_8_) & (g220) & (g264) & (g135)) + ((sk[64]) & (i_8_) & (!g220) & (g264) & (g135)) + ((sk[64]) & (i_8_) & (g220) & (!g264) & (g135)) + ((sk[64]) & (i_8_) & (g220) & (g264) & (g135)));
	assign g303 = (((!i_8_) & (!g297) & (!sk[65]) & (g264) & (g108)) + ((!i_8_) & (!g297) & (sk[65]) & (g264) & (g108)) + ((!i_8_) & (g297) & (!sk[65]) & (!g264) & (!g108)) + ((!i_8_) & (g297) & (!sk[65]) & (!g264) & (g108)) + ((!i_8_) & (g297) & (!sk[65]) & (g264) & (!g108)) + ((!i_8_) & (g297) & (!sk[65]) & (g264) & (g108)) + ((!i_8_) & (g297) & (sk[65]) & (!g264) & (g108)) + ((!i_8_) & (g297) & (sk[65]) & (g264) & (g108)) + ((i_8_) & (!g297) & (!sk[65]) & (g264) & (!g108)) + ((i_8_) & (!g297) & (!sk[65]) & (g264) & (g108)) + ((i_8_) & (g297) & (!sk[65]) & (!g264) & (!g108)) + ((i_8_) & (g297) & (!sk[65]) & (!g264) & (g108)) + ((i_8_) & (g297) & (!sk[65]) & (g264) & (!g108)) + ((i_8_) & (g297) & (!sk[65]) & (g264) & (g108)) + ((i_8_) & (g297) & (sk[65]) & (!g264) & (g108)) + ((i_8_) & (g297) & (sk[65]) & (g264) & (g108)));
	assign g304 = (((!sk[66]) & (g13) & (!g95)) + ((!sk[66]) & (g13) & (g95)) + ((sk[66]) & (g13) & (g95)));
	assign g305 = (((!i_8_) & (!g59) & (!g221) & (g88) & (!g304) & (!g270)) + ((!i_8_) & (!g59) & (!g221) & (g88) & (!g304) & (g270)) + ((!i_8_) & (!g59) & (!g221) & (g88) & (g304) & (!g270)) + ((!i_8_) & (!g59) & (!g221) & (g88) & (g304) & (g270)) + ((!i_8_) & (!g59) & (g221) & (g88) & (!g304) & (!g270)) + ((!i_8_) & (!g59) & (g221) & (g88) & (g304) & (!g270)) + ((!i_8_) & (!g59) & (g221) & (g88) & (g304) & (g270)) + ((!i_8_) & (g59) & (!g221) & (!g88) & (!g304) & (!g270)) + ((!i_8_) & (g59) & (!g221) & (!g88) & (!g304) & (g270)) + ((!i_8_) & (g59) & (!g221) & (!g88) & (g304) & (!g270)) + ((!i_8_) & (g59) & (!g221) & (!g88) & (g304) & (g270)) + ((!i_8_) & (g59) & (!g221) & (g88) & (!g304) & (!g270)) + ((!i_8_) & (g59) & (!g221) & (g88) & (!g304) & (g270)) + ((!i_8_) & (g59) & (!g221) & (g88) & (g304) & (!g270)) + ((!i_8_) & (g59) & (!g221) & (g88) & (g304) & (g270)) + ((!i_8_) & (g59) & (g221) & (g88) & (!g304) & (!g270)) + ((!i_8_) & (g59) & (g221) & (g88) & (g304) & (!g270)) + ((!i_8_) & (g59) & (g221) & (g88) & (g304) & (g270)) + ((i_8_) & (g59) & (!g221) & (!g88) & (!g304) & (!g270)) + ((i_8_) & (g59) & (!g221) & (!g88) & (!g304) & (g270)) + ((i_8_) & (g59) & (!g221) & (!g88) & (g304) & (!g270)) + ((i_8_) & (g59) & (!g221) & (!g88) & (g304) & (g270)) + ((i_8_) & (g59) & (!g221) & (g88) & (!g304) & (!g270)) + ((i_8_) & (g59) & (!g221) & (g88) & (!g304) & (g270)) + ((i_8_) & (g59) & (!g221) & (g88) & (g304) & (!g270)) + ((i_8_) & (g59) & (!g221) & (g88) & (g304) & (g270)));
	assign g306 = (((!sk[68]) & (!g89) & (!g185) & (!g302) & (!g303) & (g305)) + ((!sk[68]) & (!g89) & (!g185) & (!g302) & (g303) & (g305)) + ((!sk[68]) & (!g89) & (!g185) & (g302) & (!g303) & (g305)) + ((!sk[68]) & (!g89) & (!g185) & (g302) & (g303) & (g305)) + ((!sk[68]) & (!g89) & (g185) & (!g302) & (!g303) & (g305)) + ((!sk[68]) & (!g89) & (g185) & (!g302) & (g303) & (g305)) + ((!sk[68]) & (!g89) & (g185) & (g302) & (!g303) & (g305)) + ((!sk[68]) & (!g89) & (g185) & (g302) & (g303) & (g305)) + ((!sk[68]) & (g89) & (!g185) & (!g302) & (!g303) & (!g305)) + ((!sk[68]) & (g89) & (!g185) & (!g302) & (!g303) & (g305)) + ((!sk[68]) & (g89) & (!g185) & (!g302) & (g303) & (!g305)) + ((!sk[68]) & (g89) & (!g185) & (!g302) & (g303) & (g305)) + ((!sk[68]) & (g89) & (!g185) & (g302) & (!g303) & (!g305)) + ((!sk[68]) & (g89) & (!g185) & (g302) & (!g303) & (g305)) + ((!sk[68]) & (g89) & (!g185) & (g302) & (g303) & (!g305)) + ((!sk[68]) & (g89) & (!g185) & (g302) & (g303) & (g305)) + ((!sk[68]) & (g89) & (g185) & (!g302) & (!g303) & (!g305)) + ((!sk[68]) & (g89) & (g185) & (!g302) & (!g303) & (g305)) + ((!sk[68]) & (g89) & (g185) & (!g302) & (g303) & (!g305)) + ((!sk[68]) & (g89) & (g185) & (!g302) & (g303) & (g305)) + ((!sk[68]) & (g89) & (g185) & (g302) & (!g303) & (!g305)) + ((!sk[68]) & (g89) & (g185) & (g302) & (!g303) & (g305)) + ((!sk[68]) & (g89) & (g185) & (g302) & (g303) & (!g305)) + ((!sk[68]) & (g89) & (g185) & (g302) & (g303) & (g305)) + ((sk[68]) & (!g89) & (g185) & (!g302) & (!g303) & (!g305)) + ((sk[68]) & (g89) & (!g185) & (!g302) & (!g303) & (!g305)) + ((sk[68]) & (g89) & (g185) & (!g302) & (!g303) & (!g305)));
	assign g307 = (((!sk[69]) & (!g206) & (!g118) & (g112) & (g185)) + ((!sk[69]) & (!g206) & (g118) & (!g112) & (!g185)) + ((!sk[69]) & (!g206) & (g118) & (!g112) & (g185)) + ((!sk[69]) & (!g206) & (g118) & (g112) & (!g185)) + ((!sk[69]) & (!g206) & (g118) & (g112) & (g185)) + ((!sk[69]) & (g206) & (!g118) & (g112) & (!g185)) + ((!sk[69]) & (g206) & (!g118) & (g112) & (g185)) + ((!sk[69]) & (g206) & (g118) & (!g112) & (!g185)) + ((!sk[69]) & (g206) & (g118) & (!g112) & (g185)) + ((!sk[69]) & (g206) & (g118) & (g112) & (!g185)) + ((!sk[69]) & (g206) & (g118) & (g112) & (g185)) + ((sk[69]) & (!g206) & (!g118) & (!g112) & (!g185)) + ((sk[69]) & (!g206) & (!g118) & (!g112) & (g185)) + ((sk[69]) & (g206) & (!g118) & (!g112) & (!g185)) + ((sk[69]) & (g206) & (!g118) & (!g112) & (g185)) + ((sk[69]) & (g206) & (!g118) & (g112) & (g185)) + ((sk[69]) & (g206) & (g118) & (!g112) & (g185)) + ((sk[69]) & (g206) & (g118) & (g112) & (g185)));
	assign g308 = (((g21) & (!g149) & (!sk[70]) & (!g108)) + ((g21) & (!g149) & (!sk[70]) & (g108)) + ((g21) & (!g149) & (sk[70]) & (g108)) + ((g21) & (g149) & (!sk[70]) & (!g108)) + ((g21) & (g149) & (!sk[70]) & (g108)) + ((g21) & (g149) & (sk[70]) & (!g108)) + ((g21) & (g149) & (sk[70]) & (g108)));
	assign g309 = (((!g221) & (!sk[71]) & (!g181) & (g118) & (g270)) + ((!g221) & (!sk[71]) & (g181) & (!g118) & (!g270)) + ((!g221) & (!sk[71]) & (g181) & (!g118) & (g270)) + ((!g221) & (!sk[71]) & (g181) & (g118) & (!g270)) + ((!g221) & (!sk[71]) & (g181) & (g118) & (g270)) + ((!g221) & (sk[71]) & (!g181) & (g118) & (!g270)) + ((!g221) & (sk[71]) & (!g181) & (g118) & (g270)) + ((!g221) & (sk[71]) & (g181) & (g118) & (!g270)) + ((!g221) & (sk[71]) & (g181) & (g118) & (g270)) + ((g221) & (!sk[71]) & (!g181) & (g118) & (!g270)) + ((g221) & (!sk[71]) & (!g181) & (g118) & (g270)) + ((g221) & (!sk[71]) & (g181) & (!g118) & (!g270)) + ((g221) & (!sk[71]) & (g181) & (!g118) & (g270)) + ((g221) & (!sk[71]) & (g181) & (g118) & (!g270)) + ((g221) & (!sk[71]) & (g181) & (g118) & (g270)) + ((g221) & (sk[71]) & (!g181) & (g118) & (!g270)) + ((g221) & (sk[71]) & (g181) & (g118) & (!g270)) + ((g221) & (sk[71]) & (g181) & (g118) & (g270)));
	assign g310 = (((!g20) & (!sk[72]) & (!g99) & (g304) & (g264)) + ((!g20) & (!sk[72]) & (g99) & (!g304) & (!g264)) + ((!g20) & (!sk[72]) & (g99) & (!g304) & (g264)) + ((!g20) & (!sk[72]) & (g99) & (g304) & (!g264)) + ((!g20) & (!sk[72]) & (g99) & (g304) & (g264)) + ((!g20) & (sk[72]) & (g99) & (!g304) & (!g264)) + ((!g20) & (sk[72]) & (g99) & (!g304) & (g264)) + ((!g20) & (sk[72]) & (g99) & (g304) & (!g264)) + ((!g20) & (sk[72]) & (g99) & (g304) & (g264)) + ((g20) & (!sk[72]) & (!g99) & (g304) & (!g264)) + ((g20) & (!sk[72]) & (!g99) & (g304) & (g264)) + ((g20) & (!sk[72]) & (g99) & (!g304) & (!g264)) + ((g20) & (!sk[72]) & (g99) & (!g304) & (g264)) + ((g20) & (!sk[72]) & (g99) & (g304) & (!g264)) + ((g20) & (!sk[72]) & (g99) & (g304) & (g264)) + ((g20) & (sk[72]) & (g99) & (!g304) & (g264)) + ((g20) & (sk[72]) & (g99) & (g304) & (!g264)) + ((g20) & (sk[72]) & (g99) & (g304) & (g264)));
	assign g311 = (((!g21) & (!sk[73]) & (!g297) & (g134) & (g304)) + ((!g21) & (!sk[73]) & (g297) & (!g134) & (!g304)) + ((!g21) & (!sk[73]) & (g297) & (!g134) & (g304)) + ((!g21) & (!sk[73]) & (g297) & (g134) & (!g304)) + ((!g21) & (!sk[73]) & (g297) & (g134) & (g304)) + ((!g21) & (sk[73]) & (!g297) & (g134) & (g304)) + ((!g21) & (sk[73]) & (g297) & (g134) & (!g304)) + ((!g21) & (sk[73]) & (g297) & (g134) & (g304)) + ((g21) & (!sk[73]) & (!g297) & (g134) & (!g304)) + ((g21) & (!sk[73]) & (!g297) & (g134) & (g304)) + ((g21) & (!sk[73]) & (g297) & (!g134) & (!g304)) + ((g21) & (!sk[73]) & (g297) & (!g134) & (g304)) + ((g21) & (!sk[73]) & (g297) & (g134) & (!g304)) + ((g21) & (!sk[73]) & (g297) & (g134) & (g304)) + ((g21) & (sk[73]) & (!g297) & (g134) & (!g304)) + ((g21) & (sk[73]) & (!g297) & (g134) & (g304)) + ((g21) & (sk[73]) & (g297) & (g134) & (!g304)) + ((g21) & (sk[73]) & (g297) & (g134) & (g304)));
	assign g312 = (((!g134) & (!g220) & (!sk[74]) & (g221) & (g181)) + ((!g134) & (g220) & (!sk[74]) & (!g221) & (!g181)) + ((!g134) & (g220) & (!sk[74]) & (!g221) & (g181)) + ((!g134) & (g220) & (!sk[74]) & (g221) & (!g181)) + ((!g134) & (g220) & (!sk[74]) & (g221) & (g181)) + ((g134) & (!g220) & (!sk[74]) & (g221) & (!g181)) + ((g134) & (!g220) & (!sk[74]) & (g221) & (g181)) + ((g134) & (!g220) & (sk[74]) & (!g221) & (!g181)) + ((g134) & (!g220) & (sk[74]) & (!g221) & (g181)) + ((g134) & (!g220) & (sk[74]) & (g221) & (g181)) + ((g134) & (g220) & (!sk[74]) & (!g221) & (!g181)) + ((g134) & (g220) & (!sk[74]) & (!g221) & (g181)) + ((g134) & (g220) & (!sk[74]) & (g221) & (!g181)) + ((g134) & (g220) & (!sk[74]) & (g221) & (g181)) + ((g134) & (g220) & (sk[74]) & (!g221) & (!g181)) + ((g134) & (g220) & (sk[74]) & (!g221) & (g181)) + ((g134) & (g220) & (sk[74]) & (g221) & (!g181)) + ((g134) & (g220) & (sk[74]) & (g221) & (g181)));
	assign g313 = (((g307) & (!g308) & (!g309) & (!g310) & (!g311) & (!g312)));
	assign g314 = (((!i_8_) & (!g20) & (g108) & (!sk[76]) & (g222)) + ((!i_8_) & (!g20) & (g108) & (sk[76]) & (!g222)) + ((!i_8_) & (!g20) & (g108) & (sk[76]) & (g222)) + ((!i_8_) & (g20) & (!g108) & (!sk[76]) & (!g222)) + ((!i_8_) & (g20) & (!g108) & (!sk[76]) & (g222)) + ((!i_8_) & (g20) & (g108) & (!sk[76]) & (!g222)) + ((!i_8_) & (g20) & (g108) & (!sk[76]) & (g222)) + ((!i_8_) & (g20) & (g108) & (sk[76]) & (g222)) + ((i_8_) & (!g20) & (g108) & (!sk[76]) & (!g222)) + ((i_8_) & (!g20) & (g108) & (!sk[76]) & (g222)) + ((i_8_) & (g20) & (!g108) & (!sk[76]) & (!g222)) + ((i_8_) & (g20) & (!g108) & (!sk[76]) & (g222)) + ((i_8_) & (g20) & (g108) & (!sk[76]) & (!g222)) + ((i_8_) & (g20) & (g108) & (!sk[76]) & (g222)));
	assign g315 = (((!i_8_) & (!sk[77]) & (!g304) & (g108) & (g270)) + ((!i_8_) & (!sk[77]) & (g304) & (!g108) & (!g270)) + ((!i_8_) & (!sk[77]) & (g304) & (!g108) & (g270)) + ((!i_8_) & (!sk[77]) & (g304) & (g108) & (!g270)) + ((!i_8_) & (!sk[77]) & (g304) & (g108) & (g270)) + ((!i_8_) & (sk[77]) & (!g304) & (g108) & (!g270)) + ((!i_8_) & (sk[77]) & (g304) & (g108) & (!g270)) + ((!i_8_) & (sk[77]) & (g304) & (g108) & (g270)) + ((i_8_) & (!sk[77]) & (!g304) & (g108) & (!g270)) + ((i_8_) & (!sk[77]) & (!g304) & (g108) & (g270)) + ((i_8_) & (!sk[77]) & (g304) & (!g108) & (!g270)) + ((i_8_) & (!sk[77]) & (g304) & (!g108) & (g270)) + ((i_8_) & (!sk[77]) & (g304) & (g108) & (!g270)) + ((i_8_) & (!sk[77]) & (g304) & (g108) & (g270)));
	assign g316 = (((!sk[78]) & (g13) & (!g131)) + ((!sk[78]) & (g13) & (g131)) + ((sk[78]) & (g13) & (g131)));
	assign g317 = (((!i_8_) & (!sk[79]) & (!g108) & (g316) & (g216)) + ((!i_8_) & (!sk[79]) & (g108) & (!g316) & (!g216)) + ((!i_8_) & (!sk[79]) & (g108) & (!g316) & (g216)) + ((!i_8_) & (!sk[79]) & (g108) & (g316) & (!g216)) + ((!i_8_) & (!sk[79]) & (g108) & (g316) & (g216)) + ((!i_8_) & (sk[79]) & (g108) & (!g316) & (g216)) + ((!i_8_) & (sk[79]) & (g108) & (g316) & (!g216)) + ((!i_8_) & (sk[79]) & (g108) & (g316) & (g216)) + ((i_8_) & (!sk[79]) & (!g108) & (g316) & (!g216)) + ((i_8_) & (!sk[79]) & (!g108) & (g316) & (g216)) + ((i_8_) & (!sk[79]) & (g108) & (!g316) & (!g216)) + ((i_8_) & (!sk[79]) & (g108) & (!g316) & (g216)) + ((i_8_) & (!sk[79]) & (g108) & (g316) & (!g216)) + ((i_8_) & (!sk[79]) & (g108) & (g316) & (g216)));
	assign g318 = (((!sk[80]) & (!i_8_) & (!g206) & (g181) & (g108)) + ((!sk[80]) & (!i_8_) & (g206) & (!g181) & (!g108)) + ((!sk[80]) & (!i_8_) & (g206) & (!g181) & (g108)) + ((!sk[80]) & (!i_8_) & (g206) & (g181) & (!g108)) + ((!sk[80]) & (!i_8_) & (g206) & (g181) & (g108)) + ((!sk[80]) & (i_8_) & (!g206) & (g181) & (!g108)) + ((!sk[80]) & (i_8_) & (!g206) & (g181) & (g108)) + ((!sk[80]) & (i_8_) & (g206) & (!g181) & (!g108)) + ((!sk[80]) & (i_8_) & (g206) & (!g181) & (g108)) + ((!sk[80]) & (i_8_) & (g206) & (g181) & (!g108)) + ((!sk[80]) & (i_8_) & (g206) & (g181) & (g108)) + ((sk[80]) & (!i_8_) & (!g206) & (!g181) & (g108)) + ((sk[80]) & (!i_8_) & (!g206) & (g181) & (g108)) + ((sk[80]) & (!i_8_) & (g206) & (g181) & (g108)));
	assign g319 = (((!i_8_) & (!g220) & (!sk[81]) & (g221) & (g108)) + ((!i_8_) & (!g220) & (sk[81]) & (!g221) & (g108)) + ((!i_8_) & (g220) & (!sk[81]) & (!g221) & (!g108)) + ((!i_8_) & (g220) & (!sk[81]) & (!g221) & (g108)) + ((!i_8_) & (g220) & (!sk[81]) & (g221) & (!g108)) + ((!i_8_) & (g220) & (!sk[81]) & (g221) & (g108)) + ((!i_8_) & (g220) & (sk[81]) & (!g221) & (g108)) + ((!i_8_) & (g220) & (sk[81]) & (g221) & (g108)) + ((i_8_) & (!g220) & (!sk[81]) & (g221) & (!g108)) + ((i_8_) & (!g220) & (!sk[81]) & (g221) & (g108)) + ((i_8_) & (g220) & (!sk[81]) & (!g221) & (!g108)) + ((i_8_) & (g220) & (!sk[81]) & (!g221) & (g108)) + ((i_8_) & (g220) & (!sk[81]) & (g221) & (!g108)) + ((i_8_) & (g220) & (!sk[81]) & (g221) & (g108)));
	assign g320 = (((!g134) & (!g206) & (!g149) & (sk[82]) & (!g222)) + ((!g134) & (!g206) & (!g149) & (sk[82]) & (g222)) + ((!g134) & (!g206) & (g149) & (!sk[82]) & (g222)) + ((!g134) & (g206) & (!g149) & (!sk[82]) & (!g222)) + ((!g134) & (g206) & (!g149) & (!sk[82]) & (g222)) + ((!g134) & (g206) & (!g149) & (sk[82]) & (!g222)) + ((!g134) & (g206) & (!g149) & (sk[82]) & (g222)) + ((!g134) & (g206) & (g149) & (!sk[82]) & (!g222)) + ((!g134) & (g206) & (g149) & (!sk[82]) & (g222)) + ((!g134) & (g206) & (g149) & (sk[82]) & (!g222)) + ((!g134) & (g206) & (g149) & (sk[82]) & (g222)) + ((g134) & (!g206) & (g149) & (!sk[82]) & (!g222)) + ((g134) & (!g206) & (g149) & (!sk[82]) & (g222)) + ((g134) & (g206) & (!g149) & (!sk[82]) & (!g222)) + ((g134) & (g206) & (!g149) & (!sk[82]) & (g222)) + ((g134) & (g206) & (!g149) & (sk[82]) & (!g222)) + ((g134) & (g206) & (g149) & (!sk[82]) & (!g222)) + ((g134) & (g206) & (g149) & (!sk[82]) & (g222)) + ((g134) & (g206) & (g149) & (sk[82]) & (!g222)));
	assign g321 = (((!g314) & (!g315) & (!g317) & (!g318) & (!g319) & (g320)));
	assign g322 = (((!g301) & (!g1768) & (!g306) & (!g313) & (!sk[84]) & (g321)) + ((!g301) & (!g1768) & (!g306) & (g313) & (!sk[84]) & (g321)) + ((!g301) & (!g1768) & (g306) & (!g313) & (!sk[84]) & (g321)) + ((!g301) & (!g1768) & (g306) & (g313) & (!sk[84]) & (g321)) + ((!g301) & (g1768) & (!g306) & (!g313) & (!sk[84]) & (g321)) + ((!g301) & (g1768) & (!g306) & (g313) & (!sk[84]) & (g321)) + ((!g301) & (g1768) & (g306) & (!g313) & (!sk[84]) & (g321)) + ((!g301) & (g1768) & (g306) & (g313) & (!sk[84]) & (g321)) + ((g301) & (!g1768) & (!g306) & (!g313) & (!sk[84]) & (!g321)) + ((g301) & (!g1768) & (!g306) & (!g313) & (!sk[84]) & (g321)) + ((g301) & (!g1768) & (!g306) & (g313) & (!sk[84]) & (!g321)) + ((g301) & (!g1768) & (!g306) & (g313) & (!sk[84]) & (g321)) + ((g301) & (!g1768) & (g306) & (!g313) & (!sk[84]) & (!g321)) + ((g301) & (!g1768) & (g306) & (!g313) & (!sk[84]) & (g321)) + ((g301) & (!g1768) & (g306) & (g313) & (!sk[84]) & (!g321)) + ((g301) & (!g1768) & (g306) & (g313) & (!sk[84]) & (g321)) + ((g301) & (g1768) & (!g306) & (!g313) & (!sk[84]) & (!g321)) + ((g301) & (g1768) & (!g306) & (!g313) & (!sk[84]) & (g321)) + ((g301) & (g1768) & (!g306) & (g313) & (!sk[84]) & (!g321)) + ((g301) & (g1768) & (!g306) & (g313) & (!sk[84]) & (g321)) + ((g301) & (g1768) & (g306) & (!g313) & (!sk[84]) & (!g321)) + ((g301) & (g1768) & (g306) & (!g313) & (!sk[84]) & (g321)) + ((g301) & (g1768) & (g306) & (g313) & (!sk[84]) & (!g321)) + ((g301) & (g1768) & (g306) & (g313) & (!sk[84]) & (g321)) + ((g301) & (g1768) & (g306) & (g313) & (sk[84]) & (g321)));
	assign g323 = (((!sk[85]) & (g87) & (!g111)) + ((!sk[85]) & (g87) & (g111)) + ((sk[85]) & (g87) & (g111)));
	assign g324 = (((!i_8_) & (!sk[86]) & (!g297) & (g100) & (g316)) + ((!i_8_) & (!sk[86]) & (g297) & (!g100) & (!g316)) + ((!i_8_) & (!sk[86]) & (g297) & (!g100) & (g316)) + ((!i_8_) & (!sk[86]) & (g297) & (g100) & (!g316)) + ((!i_8_) & (!sk[86]) & (g297) & (g100) & (g316)) + ((!i_8_) & (sk[86]) & (g297) & (g100) & (!g316)) + ((!i_8_) & (sk[86]) & (g297) & (g100) & (g316)) + ((i_8_) & (!sk[86]) & (!g297) & (g100) & (!g316)) + ((i_8_) & (!sk[86]) & (!g297) & (g100) & (g316)) + ((i_8_) & (!sk[86]) & (g297) & (!g100) & (!g316)) + ((i_8_) & (!sk[86]) & (g297) & (!g100) & (g316)) + ((i_8_) & (!sk[86]) & (g297) & (g100) & (!g316)) + ((i_8_) & (!sk[86]) & (g297) & (g100) & (g316)) + ((i_8_) & (sk[86]) & (!g297) & (g100) & (g316)) + ((i_8_) & (sk[86]) & (g297) & (g100) & (!g316)) + ((i_8_) & (sk[86]) & (g297) & (g100) & (g316)));
	assign g325 = (((!g14) & (!g145) & (!g323) & (!g186) & (!g212) & (!g324)) + ((!g14) & (!g145) & (!g323) & (!g186) & (g212) & (!g324)) + ((!g14) & (!g145) & (!g323) & (g186) & (!g212) & (!g324)) + ((!g14) & (!g145) & (!g323) & (g186) & (g212) & (!g324)) + ((!g14) & (!g145) & (g323) & (!g186) & (!g212) & (!g324)) + ((!g14) & (!g145) & (g323) & (!g186) & (g212) & (!g324)) + ((!g14) & (!g145) & (g323) & (g186) & (!g212) & (!g324)) + ((!g14) & (!g145) & (g323) & (g186) & (g212) & (!g324)) + ((!g14) & (g145) & (!g323) & (!g186) & (!g212) & (!g324)) + ((!g14) & (g145) & (!g323) & (!g186) & (g212) & (!g324)) + ((!g14) & (g145) & (!g323) & (g186) & (!g212) & (!g324)) + ((!g14) & (g145) & (!g323) & (g186) & (g212) & (!g324)) + ((!g14) & (g145) & (g323) & (!g186) & (!g212) & (!g324)) + ((!g14) & (g145) & (g323) & (!g186) & (g212) & (!g324)) + ((!g14) & (g145) & (g323) & (g186) & (!g212) & (!g324)) + ((!g14) & (g145) & (g323) & (g186) & (g212) & (!g324)) + ((g14) & (!g145) & (!g323) & (!g186) & (g212) & (!g324)));
	assign g326 = (((!i_15_) & (sk[88]) & (g13)) + ((i_15_) & (!sk[88]) & (!g13)) + ((i_15_) & (!sk[88]) & (g13)));
	assign g327 = (((i_10_) & (!g326) & (!sk[89]) & (!g251)) + ((i_10_) & (!g326) & (!sk[89]) & (g251)) + ((i_10_) & (g326) & (!sk[89]) & (!g251)) + ((i_10_) & (g326) & (!sk[89]) & (g251)) + ((i_10_) & (g326) & (sk[89]) & (g251)));
	assign g328 = (((!g270) & (!sk[90]) & (!g316) & (g216) & (g207)) + ((!g270) & (!sk[90]) & (g316) & (!g216) & (!g207)) + ((!g270) & (!sk[90]) & (g316) & (!g216) & (g207)) + ((!g270) & (!sk[90]) & (g316) & (g216) & (!g207)) + ((!g270) & (!sk[90]) & (g316) & (g216) & (g207)) + ((g270) & (!sk[90]) & (!g316) & (g216) & (!g207)) + ((g270) & (!sk[90]) & (!g316) & (g216) & (g207)) + ((g270) & (!sk[90]) & (g316) & (!g216) & (!g207)) + ((g270) & (!sk[90]) & (g316) & (!g216) & (g207)) + ((g270) & (!sk[90]) & (g316) & (g216) & (!g207)) + ((g270) & (!sk[90]) & (g316) & (g216) & (g207)) + ((g270) & (sk[90]) & (!g316) & (!g216) & (!g207)));
	assign g329 = (((!g297) & (!g134) & (!sk[91]) & (!g264) & (!g328) & (g146)) + ((!g297) & (!g134) & (!sk[91]) & (!g264) & (g328) & (g146)) + ((!g297) & (!g134) & (!sk[91]) & (g264) & (!g328) & (g146)) + ((!g297) & (!g134) & (!sk[91]) & (g264) & (g328) & (g146)) + ((!g297) & (!g134) & (sk[91]) & (!g264) & (!g328) & (!g146)) + ((!g297) & (!g134) & (sk[91]) & (!g264) & (!g328) & (g146)) + ((!g297) & (!g134) & (sk[91]) & (!g264) & (g328) & (!g146)) + ((!g297) & (!g134) & (sk[91]) & (!g264) & (g328) & (g146)) + ((!g297) & (!g134) & (sk[91]) & (g264) & (!g328) & (!g146)) + ((!g297) & (!g134) & (sk[91]) & (g264) & (!g328) & (g146)) + ((!g297) & (!g134) & (sk[91]) & (g264) & (g328) & (!g146)) + ((!g297) & (!g134) & (sk[91]) & (g264) & (g328) & (g146)) + ((!g297) & (g134) & (!sk[91]) & (!g264) & (!g328) & (g146)) + ((!g297) & (g134) & (!sk[91]) & (!g264) & (g328) & (g146)) + ((!g297) & (g134) & (!sk[91]) & (g264) & (!g328) & (g146)) + ((!g297) & (g134) & (!sk[91]) & (g264) & (g328) & (g146)) + ((!g297) & (g134) & (sk[91]) & (!g264) & (g328) & (!g146)) + ((!g297) & (g134) & (sk[91]) & (!g264) & (g328) & (g146)) + ((g297) & (!g134) & (!sk[91]) & (!g264) & (!g328) & (!g146)) + ((g297) & (!g134) & (!sk[91]) & (!g264) & (!g328) & (g146)) + ((g297) & (!g134) & (!sk[91]) & (!g264) & (g328) & (!g146)) + ((g297) & (!g134) & (!sk[91]) & (!g264) & (g328) & (g146)) + ((g297) & (!g134) & (!sk[91]) & (g264) & (!g328) & (!g146)) + ((g297) & (!g134) & (!sk[91]) & (g264) & (!g328) & (g146)) + ((g297) & (!g134) & (!sk[91]) & (g264) & (g328) & (!g146)) + ((g297) & (!g134) & (!sk[91]) & (g264) & (g328) & (g146)) + ((g297) & (!g134) & (sk[91]) & (!g264) & (!g328) & (g146)) + ((g297) & (!g134) & (sk[91]) & (!g264) & (g328) & (g146)) + ((g297) & (!g134) & (sk[91]) & (g264) & (!g328) & (g146)) + ((g297) & (!g134) & (sk[91]) & (g264) & (g328) & (g146)) + ((g297) & (g134) & (!sk[91]) & (!g264) & (!g328) & (!g146)) + ((g297) & (g134) & (!sk[91]) & (!g264) & (!g328) & (g146)) + ((g297) & (g134) & (!sk[91]) & (!g264) & (g328) & (!g146)) + ((g297) & (g134) & (!sk[91]) & (!g264) & (g328) & (g146)) + ((g297) & (g134) & (!sk[91]) & (g264) & (!g328) & (!g146)) + ((g297) & (g134) & (!sk[91]) & (g264) & (!g328) & (g146)) + ((g297) & (g134) & (!sk[91]) & (g264) & (g328) & (!g146)) + ((g297) & (g134) & (!sk[91]) & (g264) & (g328) & (g146)) + ((g297) & (g134) & (sk[91]) & (!g264) & (g328) & (g146)));
	assign g330 = (((!g59) & (!g112) & (sk[92]) & (!g135)) + ((g59) & (!g112) & (!sk[92]) & (!g135)) + ((g59) & (!g112) & (!sk[92]) & (g135)) + ((g59) & (g112) & (!sk[92]) & (!g135)) + ((g59) & (g112) & (!sk[92]) & (g135)));
	assign g331 = (((!i_9_) & (!i_10_) & (g53) & (g13) & (g145) & (!g330)) + ((!i_9_) & (!i_10_) & (g53) & (g13) & (g145) & (g330)) + ((!i_9_) & (i_10_) & (g53) & (g13) & (!g145) & (!g330)) + ((!i_9_) & (i_10_) & (g53) & (g13) & (g145) & (!g330)));
	assign g332 = (((!sk[94]) & (!g21) & (!g304) & (g118) & (g112)) + ((!sk[94]) & (!g21) & (g304) & (!g118) & (!g112)) + ((!sk[94]) & (!g21) & (g304) & (!g118) & (g112)) + ((!sk[94]) & (!g21) & (g304) & (g118) & (!g112)) + ((!sk[94]) & (!g21) & (g304) & (g118) & (g112)) + ((!sk[94]) & (g21) & (!g304) & (g118) & (!g112)) + ((!sk[94]) & (g21) & (!g304) & (g118) & (g112)) + ((!sk[94]) & (g21) & (g304) & (!g118) & (!g112)) + ((!sk[94]) & (g21) & (g304) & (!g118) & (g112)) + ((!sk[94]) & (g21) & (g304) & (g118) & (!g112)) + ((!sk[94]) & (g21) & (g304) & (g118) & (g112)) + ((sk[94]) & (!g21) & (g304) & (g118) & (!g112)) + ((sk[94]) & (!g21) & (g304) & (g118) & (g112)) + ((sk[94]) & (g21) & (!g304) & (!g118) & (g112)) + ((sk[94]) & (g21) & (!g304) & (g118) & (g112)) + ((sk[94]) & (g21) & (g304) & (!g118) & (g112)) + ((sk[94]) & (g21) & (g304) & (g118) & (!g112)) + ((sk[94]) & (g21) & (g304) & (g118) & (g112)));
	assign g333 = (((!i_8_) & (g21) & (g4) & (g98) & (!g135) & (!g216)) + ((!i_8_) & (g21) & (g4) & (g98) & (!g135) & (g216)) + ((!i_8_) & (g21) & (g4) & (g98) & (g135) & (!g216)) + ((!i_8_) & (g21) & (g4) & (g98) & (g135) & (g216)) + ((i_8_) & (!g21) & (!g4) & (!g98) & (g135) & (g216)) + ((i_8_) & (!g21) & (!g4) & (g98) & (g135) & (g216)) + ((i_8_) & (!g21) & (g4) & (!g98) & (g135) & (g216)) + ((i_8_) & (!g21) & (g4) & (g98) & (g135) & (g216)) + ((i_8_) & (g21) & (!g4) & (!g98) & (g135) & (!g216)) + ((i_8_) & (g21) & (!g4) & (!g98) & (g135) & (g216)) + ((i_8_) & (g21) & (!g4) & (g98) & (g135) & (!g216)) + ((i_8_) & (g21) & (!g4) & (g98) & (g135) & (g216)) + ((i_8_) & (g21) & (g4) & (!g98) & (g135) & (!g216)) + ((i_8_) & (g21) & (g4) & (!g98) & (g135) & (g216)) + ((i_8_) & (g21) & (g4) & (g98) & (!g135) & (!g216)) + ((i_8_) & (g21) & (g4) & (g98) & (!g135) & (g216)) + ((i_8_) & (g21) & (g4) & (g98) & (g135) & (!g216)) + ((i_8_) & (g21) & (g4) & (g98) & (g135) & (g216)));
	assign g334 = (((!g304) & (!sk[96]) & (!g136) & (!g151) & (!g243) & (g333)) + ((!g304) & (!sk[96]) & (!g136) & (!g151) & (g243) & (g333)) + ((!g304) & (!sk[96]) & (!g136) & (g151) & (!g243) & (g333)) + ((!g304) & (!sk[96]) & (!g136) & (g151) & (g243) & (g333)) + ((!g304) & (!sk[96]) & (g136) & (!g151) & (!g243) & (g333)) + ((!g304) & (!sk[96]) & (g136) & (!g151) & (g243) & (g333)) + ((!g304) & (!sk[96]) & (g136) & (g151) & (!g243) & (g333)) + ((!g304) & (!sk[96]) & (g136) & (g151) & (g243) & (g333)) + ((!g304) & (sk[96]) & (!g136) & (!g151) & (!g243) & (!g333)) + ((!g304) & (sk[96]) & (!g136) & (!g151) & (g243) & (!g333)) + ((!g304) & (sk[96]) & (!g136) & (g151) & (!g243) & (!g333)) + ((!g304) & (sk[96]) & (!g136) & (g151) & (g243) & (!g333)) + ((!g304) & (sk[96]) & (g136) & (!g151) & (!g243) & (!g333)) + ((!g304) & (sk[96]) & (g136) & (!g151) & (g243) & (!g333)) + ((!g304) & (sk[96]) & (g136) & (g151) & (!g243) & (!g333)) + ((!g304) & (sk[96]) & (g136) & (g151) & (g243) & (!g333)) + ((g304) & (!sk[96]) & (!g136) & (!g151) & (!g243) & (!g333)) + ((g304) & (!sk[96]) & (!g136) & (!g151) & (!g243) & (g333)) + ((g304) & (!sk[96]) & (!g136) & (!g151) & (g243) & (!g333)) + ((g304) & (!sk[96]) & (!g136) & (!g151) & (g243) & (g333)) + ((g304) & (!sk[96]) & (!g136) & (g151) & (!g243) & (!g333)) + ((g304) & (!sk[96]) & (!g136) & (g151) & (!g243) & (g333)) + ((g304) & (!sk[96]) & (!g136) & (g151) & (g243) & (!g333)) + ((g304) & (!sk[96]) & (!g136) & (g151) & (g243) & (g333)) + ((g304) & (!sk[96]) & (g136) & (!g151) & (!g243) & (!g333)) + ((g304) & (!sk[96]) & (g136) & (!g151) & (!g243) & (g333)) + ((g304) & (!sk[96]) & (g136) & (!g151) & (g243) & (!g333)) + ((g304) & (!sk[96]) & (g136) & (!g151) & (g243) & (g333)) + ((g304) & (!sk[96]) & (g136) & (g151) & (!g243) & (!g333)) + ((g304) & (!sk[96]) & (g136) & (g151) & (!g243) & (g333)) + ((g304) & (!sk[96]) & (g136) & (g151) & (g243) & (!g333)) + ((g304) & (!sk[96]) & (g136) & (g151) & (g243) & (g333)) + ((g304) & (sk[96]) & (!g136) & (!g151) & (!g243) & (!g333)));
	assign g335 = (((!g327) & (g329) & (!g331) & (g1761) & (!g332) & (g334)));
	assign g336 = (((g276) & (!g278) & (g296) & (g322) & (g325) & (g335)));
	assign g337 = (((g136) & (!g204) & (!sk[99]) & (!g279)) + ((g136) & (!g204) & (!sk[99]) & (g279)) + ((g136) & (!g204) & (sk[99]) & (!g279)) + ((g136) & (!g204) & (sk[99]) & (g279)) + ((g136) & (g204) & (!sk[99]) & (!g279)) + ((g136) & (g204) & (!sk[99]) & (g279)) + ((g136) & (g204) & (sk[99]) & (g279)));
	assign g338 = (((!i_8_) & (!i_6_) & (!sk[100]) & (i_7_) & (g98)) + ((!i_8_) & (!i_6_) & (sk[100]) & (!i_7_) & (!g98)) + ((!i_8_) & (!i_6_) & (sk[100]) & (!i_7_) & (g98)) + ((!i_8_) & (!i_6_) & (sk[100]) & (i_7_) & (!g98)) + ((!i_8_) & (!i_6_) & (sk[100]) & (i_7_) & (g98)) + ((!i_8_) & (i_6_) & (!sk[100]) & (!i_7_) & (!g98)) + ((!i_8_) & (i_6_) & (!sk[100]) & (!i_7_) & (g98)) + ((!i_8_) & (i_6_) & (!sk[100]) & (i_7_) & (!g98)) + ((!i_8_) & (i_6_) & (!sk[100]) & (i_7_) & (g98)) + ((!i_8_) & (i_6_) & (sk[100]) & (!i_7_) & (!g98)) + ((!i_8_) & (i_6_) & (sk[100]) & (!i_7_) & (g98)) + ((!i_8_) & (i_6_) & (sk[100]) & (i_7_) & (!g98)) + ((!i_8_) & (i_6_) & (sk[100]) & (i_7_) & (g98)) + ((i_8_) & (!i_6_) & (!sk[100]) & (i_7_) & (!g98)) + ((i_8_) & (!i_6_) & (!sk[100]) & (i_7_) & (g98)) + ((i_8_) & (!i_6_) & (sk[100]) & (!i_7_) & (!g98)) + ((i_8_) & (!i_6_) & (sk[100]) & (!i_7_) & (g98)) + ((i_8_) & (!i_6_) & (sk[100]) & (i_7_) & (!g98)) + ((i_8_) & (!i_6_) & (sk[100]) & (i_7_) & (g98)) + ((i_8_) & (i_6_) & (!sk[100]) & (!i_7_) & (!g98)) + ((i_8_) & (i_6_) & (!sk[100]) & (!i_7_) & (g98)) + ((i_8_) & (i_6_) & (!sk[100]) & (i_7_) & (!g98)) + ((i_8_) & (i_6_) & (!sk[100]) & (i_7_) & (g98)) + ((i_8_) & (i_6_) & (sk[100]) & (!i_7_) & (!g98)) + ((i_8_) & (i_6_) & (sk[100]) & (i_7_) & (!g98)) + ((i_8_) & (i_6_) & (sk[100]) & (i_7_) & (g98)));
	assign g339 = (((!sk[101]) & (g18) & (!g182)) + ((!sk[101]) & (g18) & (g182)) + ((sk[101]) & (!g18) & (g182)));
	assign g340 = (((!g172) & (!g338) & (sk[102]) & (g339)) + ((g172) & (!g338) & (!sk[102]) & (!g339)) + ((g172) & (!g338) & (!sk[102]) & (g339)) + ((g172) & (!g338) & (sk[102]) & (!g339)) + ((g172) & (!g338) & (sk[102]) & (g339)) + ((g172) & (g338) & (!sk[102]) & (!g339)) + ((g172) & (g338) & (!sk[102]) & (g339)));
	assign g341 = (((!sk[103]) & (g203) & (!g268) & (!g338)) + ((!sk[103]) & (g203) & (!g268) & (g338)) + ((!sk[103]) & (g203) & (g268) & (!g338)) + ((!sk[103]) & (g203) & (g268) & (g338)) + ((sk[103]) & (!g203) & (g268) & (!g338)) + ((sk[103]) & (g203) & (!g268) & (!g338)) + ((sk[103]) & (g203) & (g268) & (!g338)));
	assign g342 = (((!sk[104]) & (!g112) & (!g203) & (g224) & (g254)) + ((!sk[104]) & (!g112) & (g203) & (!g224) & (!g254)) + ((!sk[104]) & (!g112) & (g203) & (!g224) & (g254)) + ((!sk[104]) & (!g112) & (g203) & (g224) & (!g254)) + ((!sk[104]) & (!g112) & (g203) & (g224) & (g254)) + ((!sk[104]) & (g112) & (!g203) & (g224) & (!g254)) + ((!sk[104]) & (g112) & (!g203) & (g224) & (g254)) + ((!sk[104]) & (g112) & (g203) & (!g224) & (!g254)) + ((!sk[104]) & (g112) & (g203) & (!g224) & (g254)) + ((!sk[104]) & (g112) & (g203) & (g224) & (!g254)) + ((!sk[104]) & (g112) & (g203) & (g224) & (g254)) + ((sk[104]) & (g112) & (!g203) & (!g224) & (g254)) + ((sk[104]) & (g112) & (!g203) & (g224) & (!g254)) + ((sk[104]) & (g112) & (!g203) & (g224) & (g254)) + ((sk[104]) & (g112) & (g203) & (!g224) & (!g254)) + ((sk[104]) & (g112) & (g203) & (!g224) & (g254)) + ((sk[104]) & (g112) & (g203) & (g224) & (!g254)) + ((sk[104]) & (g112) & (g203) & (g224) & (g254)));
	assign g343 = (((!g112) & (!sk[105]) & (!g323) & (g226) & (g231)) + ((!g112) & (!sk[105]) & (g323) & (!g226) & (!g231)) + ((!g112) & (!sk[105]) & (g323) & (!g226) & (g231)) + ((!g112) & (!sk[105]) & (g323) & (g226) & (!g231)) + ((!g112) & (!sk[105]) & (g323) & (g226) & (g231)) + ((!g112) & (sk[105]) & (!g323) & (!g226) & (!g231)) + ((!g112) & (sk[105]) & (!g323) & (!g226) & (g231)) + ((!g112) & (sk[105]) & (!g323) & (g226) & (!g231)) + ((!g112) & (sk[105]) & (!g323) & (g226) & (g231)) + ((!g112) & (sk[105]) & (g323) & (g226) & (!g231)) + ((!g112) & (sk[105]) & (g323) & (g226) & (g231)) + ((g112) & (!sk[105]) & (!g323) & (g226) & (!g231)) + ((g112) & (!sk[105]) & (!g323) & (g226) & (g231)) + ((g112) & (!sk[105]) & (g323) & (!g226) & (!g231)) + ((g112) & (!sk[105]) & (g323) & (!g226) & (g231)) + ((g112) & (!sk[105]) & (g323) & (g226) & (!g231)) + ((g112) & (!sk[105]) & (g323) & (g226) & (g231)) + ((g112) & (sk[105]) & (!g323) & (g226) & (g231)) + ((g112) & (sk[105]) & (g323) & (g226) & (g231)));
	assign g344 = (((i_8_) & (g100) & (!g226) & (!g268) & (!g279) & (!g339)) + ((i_8_) & (g100) & (!g226) & (!g268) & (!g279) & (g339)) + ((i_8_) & (g100) & (!g226) & (!g268) & (g279) & (!g339)) + ((i_8_) & (g100) & (!g226) & (!g268) & (g279) & (g339)) + ((i_8_) & (g100) & (!g226) & (g268) & (!g279) & (!g339)) + ((i_8_) & (g100) & (!g226) & (g268) & (!g279) & (g339)) + ((i_8_) & (g100) & (!g226) & (g268) & (g279) & (!g339)) + ((i_8_) & (g100) & (!g226) & (g268) & (g279) & (g339)) + ((i_8_) & (g100) & (g226) & (!g268) & (!g279) & (g339)) + ((i_8_) & (g100) & (g226) & (!g268) & (g279) & (!g339)) + ((i_8_) & (g100) & (g226) & (!g268) & (g279) & (g339)) + ((i_8_) & (g100) & (g226) & (g268) & (!g279) & (!g339)) + ((i_8_) & (g100) & (g226) & (g268) & (!g279) & (g339)) + ((i_8_) & (g100) & (g226) & (g268) & (g279) & (!g339)) + ((i_8_) & (g100) & (g226) & (g268) & (g279) & (g339)));
	assign g345 = (((!g340) & (!g341) & (!g342) & (!sk[107]) & (!g343) & (g344)) + ((!g340) & (!g341) & (!g342) & (!sk[107]) & (g343) & (g344)) + ((!g340) & (!g341) & (!g342) & (sk[107]) & (g343) & (!g344)) + ((!g340) & (!g341) & (g342) & (!sk[107]) & (!g343) & (g344)) + ((!g340) & (!g341) & (g342) & (!sk[107]) & (g343) & (g344)) + ((!g340) & (g341) & (!g342) & (!sk[107]) & (!g343) & (g344)) + ((!g340) & (g341) & (!g342) & (!sk[107]) & (g343) & (g344)) + ((!g340) & (g341) & (g342) & (!sk[107]) & (!g343) & (g344)) + ((!g340) & (g341) & (g342) & (!sk[107]) & (g343) & (g344)) + ((g340) & (!g341) & (!g342) & (!sk[107]) & (!g343) & (!g344)) + ((g340) & (!g341) & (!g342) & (!sk[107]) & (!g343) & (g344)) + ((g340) & (!g341) & (!g342) & (!sk[107]) & (g343) & (!g344)) + ((g340) & (!g341) & (!g342) & (!sk[107]) & (g343) & (g344)) + ((g340) & (!g341) & (g342) & (!sk[107]) & (!g343) & (!g344)) + ((g340) & (!g341) & (g342) & (!sk[107]) & (!g343) & (g344)) + ((g340) & (!g341) & (g342) & (!sk[107]) & (g343) & (!g344)) + ((g340) & (!g341) & (g342) & (!sk[107]) & (g343) & (g344)) + ((g340) & (g341) & (!g342) & (!sk[107]) & (!g343) & (!g344)) + ((g340) & (g341) & (!g342) & (!sk[107]) & (!g343) & (g344)) + ((g340) & (g341) & (!g342) & (!sk[107]) & (g343) & (!g344)) + ((g340) & (g341) & (!g342) & (!sk[107]) & (g343) & (g344)) + ((g340) & (g341) & (g342) & (!sk[107]) & (!g343) & (!g344)) + ((g340) & (g341) & (g342) & (!sk[107]) & (!g343) & (g344)) + ((g340) & (g341) & (g342) & (!sk[107]) & (g343) & (!g344)) + ((g340) & (g341) & (g342) & (!sk[107]) & (g343) & (g344)));
	assign g346 = (((!sk[108]) & (!i_8_) & (!g88) & (g224) & (g232)) + ((!sk[108]) & (!i_8_) & (g88) & (!g224) & (!g232)) + ((!sk[108]) & (!i_8_) & (g88) & (!g224) & (g232)) + ((!sk[108]) & (!i_8_) & (g88) & (g224) & (!g232)) + ((!sk[108]) & (!i_8_) & (g88) & (g224) & (g232)) + ((!sk[108]) & (i_8_) & (!g88) & (g224) & (!g232)) + ((!sk[108]) & (i_8_) & (!g88) & (g224) & (g232)) + ((!sk[108]) & (i_8_) & (g88) & (!g224) & (!g232)) + ((!sk[108]) & (i_8_) & (g88) & (!g224) & (g232)) + ((!sk[108]) & (i_8_) & (g88) & (g224) & (!g232)) + ((!sk[108]) & (i_8_) & (g88) & (g224) & (g232)) + ((sk[108]) & (i_8_) & (g88) & (!g224) & (g232)) + ((sk[108]) & (i_8_) & (g88) & (g224) & (!g232)) + ((sk[108]) & (i_8_) & (g88) & (g224) & (g232)));
	assign g347 = (((!g112) & (!g151) & (!g204) & (!g279) & (!g284) & (!g346)) + ((!g112) & (!g151) & (!g204) & (g279) & (!g284) & (!g346)) + ((!g112) & (!g151) & (g204) & (!g279) & (!g284) & (!g346)) + ((!g112) & (!g151) & (g204) & (!g279) & (g284) & (!g346)) + ((!g112) & (!g151) & (g204) & (g279) & (!g284) & (!g346)) + ((!g112) & (g151) & (g204) & (!g279) & (!g284) & (!g346)) + ((!g112) & (g151) & (g204) & (!g279) & (g284) & (!g346)) + ((g112) & (!g151) & (g204) & (!g279) & (!g284) & (!g346)) + ((g112) & (!g151) & (g204) & (!g279) & (g284) & (!g346)) + ((g112) & (g151) & (g204) & (!g279) & (!g284) & (!g346)) + ((g112) & (g151) & (g204) & (!g279) & (g284) & (!g346)));
	assign g348 = (((!g323) & (!g224) & (g232) & (!sk[110]) & (g339)) + ((!g323) & (g224) & (!g232) & (!sk[110]) & (!g339)) + ((!g323) & (g224) & (!g232) & (!sk[110]) & (g339)) + ((!g323) & (g224) & (g232) & (!sk[110]) & (!g339)) + ((!g323) & (g224) & (g232) & (!sk[110]) & (g339)) + ((g323) & (!g224) & (!g232) & (sk[110]) & (g339)) + ((g323) & (!g224) & (g232) & (!sk[110]) & (!g339)) + ((g323) & (!g224) & (g232) & (!sk[110]) & (g339)) + ((g323) & (!g224) & (g232) & (sk[110]) & (!g339)) + ((g323) & (!g224) & (g232) & (sk[110]) & (g339)) + ((g323) & (g224) & (!g232) & (!sk[110]) & (!g339)) + ((g323) & (g224) & (!g232) & (!sk[110]) & (g339)) + ((g323) & (g224) & (!g232) & (sk[110]) & (!g339)) + ((g323) & (g224) & (!g232) & (sk[110]) & (g339)) + ((g323) & (g224) & (g232) & (!sk[110]) & (!g339)) + ((g323) & (g224) & (g232) & (!sk[110]) & (g339)) + ((g323) & (g224) & (g232) & (sk[110]) & (!g339)) + ((g323) & (g224) & (g232) & (sk[110]) & (g339)));
	assign g349 = (((!sk[111]) & (g182) & (!g122)) + ((!sk[111]) & (g182) & (g122)) + ((sk[111]) & (g182) & (!g122)));
	assign g350 = (((!g112) & (!g232) & (g349) & (!sk[112]) & (g339)) + ((!g112) & (g232) & (!g349) & (!sk[112]) & (!g339)) + ((!g112) & (g232) & (!g349) & (!sk[112]) & (g339)) + ((!g112) & (g232) & (g349) & (!sk[112]) & (!g339)) + ((!g112) & (g232) & (g349) & (!sk[112]) & (g339)) + ((g112) & (!g232) & (!g349) & (sk[112]) & (g339)) + ((g112) & (!g232) & (g349) & (!sk[112]) & (!g339)) + ((g112) & (!g232) & (g349) & (!sk[112]) & (g339)) + ((g112) & (!g232) & (g349) & (sk[112]) & (!g339)) + ((g112) & (!g232) & (g349) & (sk[112]) & (g339)) + ((g112) & (g232) & (!g349) & (!sk[112]) & (!g339)) + ((g112) & (g232) & (!g349) & (!sk[112]) & (g339)) + ((g112) & (g232) & (!g349) & (sk[112]) & (!g339)) + ((g112) & (g232) & (!g349) & (sk[112]) & (g339)) + ((g112) & (g232) & (g349) & (!sk[112]) & (!g339)) + ((g112) & (g232) & (g349) & (!sk[112]) & (g339)) + ((g112) & (g232) & (g349) & (sk[112]) & (!g339)) + ((g112) & (g232) & (g349) & (sk[112]) & (g339)));
	assign g351 = (((!sk[113]) & (!i_8_) & (!g135) & (g231) & (g349)) + ((!sk[113]) & (!i_8_) & (g135) & (!g231) & (!g349)) + ((!sk[113]) & (!i_8_) & (g135) & (!g231) & (g349)) + ((!sk[113]) & (!i_8_) & (g135) & (g231) & (!g349)) + ((!sk[113]) & (!i_8_) & (g135) & (g231) & (g349)) + ((!sk[113]) & (i_8_) & (!g135) & (g231) & (!g349)) + ((!sk[113]) & (i_8_) & (!g135) & (g231) & (g349)) + ((!sk[113]) & (i_8_) & (g135) & (!g231) & (!g349)) + ((!sk[113]) & (i_8_) & (g135) & (!g231) & (g349)) + ((!sk[113]) & (i_8_) & (g135) & (g231) & (!g349)) + ((!sk[113]) & (i_8_) & (g135) & (g231) & (g349)) + ((sk[113]) & (i_8_) & (g135) & (!g231) & (!g349)) + ((sk[113]) & (i_8_) & (g135) & (!g231) & (g349)) + ((sk[113]) & (i_8_) & (g135) & (g231) & (g349)));
	assign g352 = (((i_8_) & (g135) & (!g226) & (!g224) & (!g232) & (!g339)) + ((i_8_) & (g135) & (!g226) & (!g224) & (!g232) & (g339)) + ((i_8_) & (g135) & (!g226) & (!g224) & (g232) & (!g339)) + ((i_8_) & (g135) & (!g226) & (!g224) & (g232) & (g339)) + ((i_8_) & (g135) & (!g226) & (g224) & (!g232) & (!g339)) + ((i_8_) & (g135) & (!g226) & (g224) & (!g232) & (g339)) + ((i_8_) & (g135) & (!g226) & (g224) & (g232) & (!g339)) + ((i_8_) & (g135) & (!g226) & (g224) & (g232) & (g339)) + ((i_8_) & (g135) & (g226) & (!g224) & (!g232) & (g339)) + ((i_8_) & (g135) & (g226) & (!g224) & (g232) & (!g339)) + ((i_8_) & (g135) & (g226) & (!g224) & (g232) & (g339)) + ((i_8_) & (g135) & (g226) & (g224) & (!g232) & (!g339)) + ((i_8_) & (g135) & (g226) & (g224) & (!g232) & (g339)) + ((i_8_) & (g135) & (g226) & (g224) & (g232) & (!g339)) + ((i_8_) & (g135) & (g226) & (g224) & (g232) & (g339)));
	assign g353 = (((!g136) & (!g203) & (!g348) & (!g350) & (!g351) & (!g352)) + ((!g136) & (g203) & (!g348) & (!g350) & (!g351) & (!g352)) + ((g136) & (!g203) & (!g348) & (!g350) & (!g351) & (!g352)));
	assign g354 = (((g151) & (!sk[116]) & (!g226) & (!g339)) + ((g151) & (!sk[116]) & (!g226) & (g339)) + ((g151) & (!sk[116]) & (g226) & (!g339)) + ((g151) & (!sk[116]) & (g226) & (g339)) + ((g151) & (sk[116]) & (!g226) & (!g339)) + ((g151) & (sk[116]) & (!g226) & (g339)) + ((g151) & (sk[116]) & (g226) & (g339)));
	assign g355 = (((!i_8_) & (!g108) & (g203) & (!sk[117]) & (g204)) + ((!i_8_) & (g108) & (!g203) & (!sk[117]) & (!g204)) + ((!i_8_) & (g108) & (!g203) & (!sk[117]) & (g204)) + ((!i_8_) & (g108) & (g203) & (!sk[117]) & (!g204)) + ((!i_8_) & (g108) & (g203) & (!sk[117]) & (g204)) + ((i_8_) & (!g108) & (g203) & (!sk[117]) & (!g204)) + ((i_8_) & (!g108) & (g203) & (!sk[117]) & (g204)) + ((i_8_) & (g108) & (!g203) & (!sk[117]) & (!g204)) + ((i_8_) & (g108) & (!g203) & (!sk[117]) & (g204)) + ((i_8_) & (g108) & (!g203) & (sk[117]) & (!g204)) + ((i_8_) & (g108) & (g203) & (!sk[117]) & (!g204)) + ((i_8_) & (g108) & (g203) & (!sk[117]) & (g204)) + ((i_8_) & (g108) & (g203) & (sk[117]) & (!g204)) + ((i_8_) & (g108) & (g203) & (sk[117]) & (g204)));
	assign g356 = (((i_8_) & (g108) & (!g226) & (!g224) & (!g231) & (!g232)) + ((i_8_) & (g108) & (!g226) & (!g224) & (!g231) & (g232)) + ((i_8_) & (g108) & (!g226) & (!g224) & (g231) & (!g232)) + ((i_8_) & (g108) & (!g226) & (!g224) & (g231) & (g232)) + ((i_8_) & (g108) & (!g226) & (g224) & (!g231) & (!g232)) + ((i_8_) & (g108) & (!g226) & (g224) & (!g231) & (g232)) + ((i_8_) & (g108) & (!g226) & (g224) & (g231) & (!g232)) + ((i_8_) & (g108) & (!g226) & (g224) & (g231) & (g232)) + ((i_8_) & (g108) & (g226) & (!g224) & (!g231) & (!g232)) + ((i_8_) & (g108) & (g226) & (!g224) & (!g231) & (g232)) + ((i_8_) & (g108) & (g226) & (!g224) & (g231) & (g232)) + ((i_8_) & (g108) & (g226) & (g224) & (!g231) & (!g232)) + ((i_8_) & (g108) & (g226) & (g224) & (!g231) & (g232)) + ((i_8_) & (g108) & (g226) & (g224) & (g231) & (!g232)) + ((i_8_) & (g108) & (g226) & (g224) & (g231) & (g232)));
	assign g357 = (((!g323) & (!g151) & (!g203) & (!g349) & (!g355) & (!g356)) + ((!g323) & (!g151) & (!g203) & (g349) & (!g355) & (!g356)) + ((!g323) & (!g151) & (g203) & (!g349) & (!g355) & (!g356)) + ((!g323) & (!g151) & (g203) & (g349) & (!g355) & (!g356)) + ((!g323) & (g151) & (!g203) & (!g349) & (!g355) & (!g356)) + ((g323) & (!g151) & (!g203) & (!g349) & (!g355) & (!g356)) + ((g323) & (g151) & (!g203) & (!g349) & (!g355) & (!g356)));
	assign g358 = (((!g337) & (g345) & (g347) & (g353) & (!g354) & (g357)));
	assign g359 = (((!g244) & (!g112) & (!g136) & (!g222) & (!sk[121]) & (g178)) + ((!g244) & (!g112) & (!g136) & (g222) & (!sk[121]) & (g178)) + ((!g244) & (!g112) & (g136) & (!g222) & (!sk[121]) & (g178)) + ((!g244) & (!g112) & (g136) & (g222) & (!sk[121]) & (g178)) + ((!g244) & (!g112) & (g136) & (g222) & (sk[121]) & (!g178)) + ((!g244) & (!g112) & (g136) & (g222) & (sk[121]) & (g178)) + ((!g244) & (g112) & (!g136) & (!g222) & (!sk[121]) & (g178)) + ((!g244) & (g112) & (!g136) & (g222) & (!sk[121]) & (g178)) + ((!g244) & (g112) & (!g136) & (g222) & (sk[121]) & (!g178)) + ((!g244) & (g112) & (!g136) & (g222) & (sk[121]) & (g178)) + ((!g244) & (g112) & (g136) & (!g222) & (!sk[121]) & (g178)) + ((!g244) & (g112) & (g136) & (g222) & (!sk[121]) & (g178)) + ((!g244) & (g112) & (g136) & (g222) & (sk[121]) & (!g178)) + ((!g244) & (g112) & (g136) & (g222) & (sk[121]) & (g178)) + ((g244) & (!g112) & (!g136) & (!g222) & (!sk[121]) & (!g178)) + ((g244) & (!g112) & (!g136) & (!g222) & (!sk[121]) & (g178)) + ((g244) & (!g112) & (!g136) & (g222) & (!sk[121]) & (!g178)) + ((g244) & (!g112) & (!g136) & (g222) & (!sk[121]) & (g178)) + ((g244) & (!g112) & (g136) & (!g222) & (!sk[121]) & (!g178)) + ((g244) & (!g112) & (g136) & (!g222) & (!sk[121]) & (g178)) + ((g244) & (!g112) & (g136) & (g222) & (!sk[121]) & (!g178)) + ((g244) & (!g112) & (g136) & (g222) & (!sk[121]) & (g178)) + ((g244) & (!g112) & (g136) & (g222) & (sk[121]) & (!g178)) + ((g244) & (!g112) & (g136) & (g222) & (sk[121]) & (g178)) + ((g244) & (g112) & (!g136) & (!g222) & (!sk[121]) & (!g178)) + ((g244) & (g112) & (!g136) & (!g222) & (!sk[121]) & (g178)) + ((g244) & (g112) & (!g136) & (!g222) & (sk[121]) & (g178)) + ((g244) & (g112) & (!g136) & (g222) & (!sk[121]) & (!g178)) + ((g244) & (g112) & (!g136) & (g222) & (!sk[121]) & (g178)) + ((g244) & (g112) & (!g136) & (g222) & (sk[121]) & (!g178)) + ((g244) & (g112) & (!g136) & (g222) & (sk[121]) & (g178)) + ((g244) & (g112) & (g136) & (!g222) & (!sk[121]) & (!g178)) + ((g244) & (g112) & (g136) & (!g222) & (!sk[121]) & (g178)) + ((g244) & (g112) & (g136) & (!g222) & (sk[121]) & (g178)) + ((g244) & (g112) & (g136) & (g222) & (!sk[121]) & (!g178)) + ((g244) & (g112) & (g136) & (g222) & (!sk[121]) & (g178)) + ((g244) & (g112) & (g136) & (g222) & (sk[121]) & (!g178)) + ((g244) & (g112) & (g136) & (g222) & (sk[121]) & (g178)));
	assign g360 = (((!g145) & (!g112) & (!g136) & (!g222) & (!g151) & (!g284)) + ((!g145) & (!g112) & (!g136) & (g222) & (!g151) & (!g284)) + ((!g145) & (!g112) & (g136) & (!g222) & (!g151) & (!g284)));
	assign g361 = (((!sk[123]) & (!i_14_) & (!i_12_) & (!i_13_) & (!g15) & (g338)) + ((!sk[123]) & (!i_14_) & (!i_12_) & (!i_13_) & (g15) & (g338)) + ((!sk[123]) & (!i_14_) & (!i_12_) & (i_13_) & (!g15) & (g338)) + ((!sk[123]) & (!i_14_) & (!i_12_) & (i_13_) & (g15) & (g338)) + ((!sk[123]) & (!i_14_) & (i_12_) & (!i_13_) & (!g15) & (g338)) + ((!sk[123]) & (!i_14_) & (i_12_) & (!i_13_) & (g15) & (g338)) + ((!sk[123]) & (!i_14_) & (i_12_) & (i_13_) & (!g15) & (g338)) + ((!sk[123]) & (!i_14_) & (i_12_) & (i_13_) & (g15) & (g338)) + ((!sk[123]) & (i_14_) & (!i_12_) & (!i_13_) & (!g15) & (!g338)) + ((!sk[123]) & (i_14_) & (!i_12_) & (!i_13_) & (!g15) & (g338)) + ((!sk[123]) & (i_14_) & (!i_12_) & (!i_13_) & (g15) & (!g338)) + ((!sk[123]) & (i_14_) & (!i_12_) & (!i_13_) & (g15) & (g338)) + ((!sk[123]) & (i_14_) & (!i_12_) & (i_13_) & (!g15) & (!g338)) + ((!sk[123]) & (i_14_) & (!i_12_) & (i_13_) & (!g15) & (g338)) + ((!sk[123]) & (i_14_) & (!i_12_) & (i_13_) & (g15) & (!g338)) + ((!sk[123]) & (i_14_) & (!i_12_) & (i_13_) & (g15) & (g338)) + ((!sk[123]) & (i_14_) & (i_12_) & (!i_13_) & (!g15) & (!g338)) + ((!sk[123]) & (i_14_) & (i_12_) & (!i_13_) & (!g15) & (g338)) + ((!sk[123]) & (i_14_) & (i_12_) & (!i_13_) & (g15) & (!g338)) + ((!sk[123]) & (i_14_) & (i_12_) & (!i_13_) & (g15) & (g338)) + ((!sk[123]) & (i_14_) & (i_12_) & (i_13_) & (!g15) & (!g338)) + ((!sk[123]) & (i_14_) & (i_12_) & (i_13_) & (!g15) & (g338)) + ((!sk[123]) & (i_14_) & (i_12_) & (i_13_) & (g15) & (!g338)) + ((!sk[123]) & (i_14_) & (i_12_) & (i_13_) & (g15) & (g338)) + ((sk[123]) & (!i_14_) & (i_12_) & (!i_13_) & (!g15) & (!g338)) + ((sk[123]) & (i_14_) & (!i_12_) & (!i_13_) & (!g15) & (!g338)));
	assign g362 = (((!sk[124]) & (g220) & (!g145) & (!g361)) + ((!sk[124]) & (g220) & (!g145) & (g361)) + ((!sk[124]) & (g220) & (g145) & (!g361)) + ((!sk[124]) & (g220) & (g145) & (g361)) + ((sk[124]) & (!g220) & (!g145) & (!g361)) + ((sk[124]) & (!g220) & (g145) & (!g361)) + ((sk[124]) & (g220) & (!g145) & (!g361)));
	assign g363 = (((!i_8_) & (!g20) & (g108) & (!sk[125]) & (g222)) + ((!i_8_) & (g20) & (!g108) & (!sk[125]) & (!g222)) + ((!i_8_) & (g20) & (!g108) & (!sk[125]) & (g222)) + ((!i_8_) & (g20) & (g108) & (!sk[125]) & (!g222)) + ((!i_8_) & (g20) & (g108) & (!sk[125]) & (g222)) + ((i_8_) & (!g20) & (g108) & (!sk[125]) & (!g222)) + ((i_8_) & (!g20) & (g108) & (!sk[125]) & (g222)) + ((i_8_) & (!g20) & (g108) & (sk[125]) & (!g222)) + ((i_8_) & (!g20) & (g108) & (sk[125]) & (g222)) + ((i_8_) & (g20) & (!g108) & (!sk[125]) & (!g222)) + ((i_8_) & (g20) & (!g108) & (!sk[125]) & (g222)) + ((i_8_) & (g20) & (g108) & (!sk[125]) & (!g222)) + ((i_8_) & (g20) & (g108) & (!sk[125]) & (g222)) + ((i_8_) & (g20) & (g108) & (sk[125]) & (g222)));
	assign g364 = (((!i_8_) & (!g221) & (!sk[126]) & (g88) & (g270)) + ((!i_8_) & (g221) & (!sk[126]) & (!g88) & (!g270)) + ((!i_8_) & (g221) & (!sk[126]) & (!g88) & (g270)) + ((!i_8_) & (g221) & (!sk[126]) & (g88) & (!g270)) + ((!i_8_) & (g221) & (!sk[126]) & (g88) & (g270)) + ((i_8_) & (!g221) & (!sk[126]) & (g88) & (!g270)) + ((i_8_) & (!g221) & (!sk[126]) & (g88) & (g270)) + ((i_8_) & (!g221) & (sk[126]) & (g88) & (!g270)) + ((i_8_) & (!g221) & (sk[126]) & (g88) & (g270)) + ((i_8_) & (g221) & (!sk[126]) & (!g88) & (!g270)) + ((i_8_) & (g221) & (!sk[126]) & (!g88) & (g270)) + ((i_8_) & (g221) & (!sk[126]) & (g88) & (!g270)) + ((i_8_) & (g221) & (!sk[126]) & (g88) & (g270)) + ((i_8_) & (g221) & (sk[126]) & (g88) & (!g270)));
	assign g365 = (((!i_8_) & (!g206) & (g88) & (!sk[127]) & (g181)) + ((!i_8_) & (g206) & (!g88) & (!sk[127]) & (!g181)) + ((!i_8_) & (g206) & (!g88) & (!sk[127]) & (g181)) + ((!i_8_) & (g206) & (g88) & (!sk[127]) & (!g181)) + ((!i_8_) & (g206) & (g88) & (!sk[127]) & (g181)) + ((i_8_) & (!g206) & (g88) & (!sk[127]) & (!g181)) + ((i_8_) & (!g206) & (g88) & (!sk[127]) & (g181)) + ((i_8_) & (!g206) & (g88) & (sk[127]) & (!g181)) + ((i_8_) & (!g206) & (g88) & (sk[127]) & (g181)) + ((i_8_) & (g206) & (!g88) & (!sk[127]) & (!g181)) + ((i_8_) & (g206) & (!g88) & (!sk[127]) & (g181)) + ((i_8_) & (g206) & (g88) & (!sk[127]) & (!g181)) + ((i_8_) & (g206) & (g88) & (!sk[127]) & (g181)) + ((i_8_) & (g206) & (g88) & (sk[127]) & (g181)));
	assign g366 = (((!i_8_) & (!g206) & (g108) & (!sk[0]) & (g185)) + ((!i_8_) & (g206) & (!g108) & (!sk[0]) & (!g185)) + ((!i_8_) & (g206) & (!g108) & (!sk[0]) & (g185)) + ((!i_8_) & (g206) & (g108) & (!sk[0]) & (!g185)) + ((!i_8_) & (g206) & (g108) & (!sk[0]) & (g185)) + ((i_8_) & (!g206) & (g108) & (!sk[0]) & (!g185)) + ((i_8_) & (!g206) & (g108) & (!sk[0]) & (g185)) + ((i_8_) & (!g206) & (g108) & (sk[0]) & (!g185)) + ((i_8_) & (!g206) & (g108) & (sk[0]) & (g185)) + ((i_8_) & (g206) & (!g108) & (!sk[0]) & (!g185)) + ((i_8_) & (g206) & (!g108) & (!sk[0]) & (g185)) + ((i_8_) & (g206) & (g108) & (!sk[0]) & (!g185)) + ((i_8_) & (g206) & (g108) & (!sk[0]) & (g185)) + ((i_8_) & (g206) & (g108) & (sk[0]) & (!g185)));
	assign g367 = (((!i_8_) & (!g304) & (!g108) & (!g270) & (!sk[1]) & (g216)) + ((!i_8_) & (!g304) & (!g108) & (g270) & (!sk[1]) & (g216)) + ((!i_8_) & (!g304) & (g108) & (!g270) & (!sk[1]) & (g216)) + ((!i_8_) & (!g304) & (g108) & (g270) & (!sk[1]) & (g216)) + ((!i_8_) & (g304) & (!g108) & (!g270) & (!sk[1]) & (g216)) + ((!i_8_) & (g304) & (!g108) & (g270) & (!sk[1]) & (g216)) + ((!i_8_) & (g304) & (g108) & (!g270) & (!sk[1]) & (g216)) + ((!i_8_) & (g304) & (g108) & (g270) & (!sk[1]) & (g216)) + ((i_8_) & (!g304) & (!g108) & (!g270) & (!sk[1]) & (!g216)) + ((i_8_) & (!g304) & (!g108) & (!g270) & (!sk[1]) & (g216)) + ((i_8_) & (!g304) & (!g108) & (g270) & (!sk[1]) & (!g216)) + ((i_8_) & (!g304) & (!g108) & (g270) & (!sk[1]) & (g216)) + ((i_8_) & (!g304) & (g108) & (!g270) & (!sk[1]) & (!g216)) + ((i_8_) & (!g304) & (g108) & (!g270) & (!sk[1]) & (g216)) + ((i_8_) & (!g304) & (g108) & (!g270) & (sk[1]) & (!g216)) + ((i_8_) & (!g304) & (g108) & (!g270) & (sk[1]) & (g216)) + ((i_8_) & (!g304) & (g108) & (g270) & (!sk[1]) & (!g216)) + ((i_8_) & (!g304) & (g108) & (g270) & (!sk[1]) & (g216)) + ((i_8_) & (!g304) & (g108) & (g270) & (sk[1]) & (g216)) + ((i_8_) & (g304) & (!g108) & (!g270) & (!sk[1]) & (!g216)) + ((i_8_) & (g304) & (!g108) & (!g270) & (!sk[1]) & (g216)) + ((i_8_) & (g304) & (!g108) & (g270) & (!sk[1]) & (!g216)) + ((i_8_) & (g304) & (!g108) & (g270) & (!sk[1]) & (g216)) + ((i_8_) & (g304) & (g108) & (!g270) & (!sk[1]) & (!g216)) + ((i_8_) & (g304) & (g108) & (!g270) & (!sk[1]) & (g216)) + ((i_8_) & (g304) & (g108) & (!g270) & (sk[1]) & (!g216)) + ((i_8_) & (g304) & (g108) & (!g270) & (sk[1]) & (g216)) + ((i_8_) & (g304) & (g108) & (g270) & (!sk[1]) & (!g216)) + ((i_8_) & (g304) & (g108) & (g270) & (!sk[1]) & (g216)) + ((i_8_) & (g304) & (g108) & (g270) & (sk[1]) & (!g216)) + ((i_8_) & (g304) & (g108) & (g270) & (sk[1]) & (g216)));
	assign g368 = (((!g363) & (!sk[2]) & (!g364) & (!g365) & (!g366) & (g367)) + ((!g363) & (!sk[2]) & (!g364) & (!g365) & (g366) & (g367)) + ((!g363) & (!sk[2]) & (!g364) & (g365) & (!g366) & (g367)) + ((!g363) & (!sk[2]) & (!g364) & (g365) & (g366) & (g367)) + ((!g363) & (!sk[2]) & (g364) & (!g365) & (!g366) & (g367)) + ((!g363) & (!sk[2]) & (g364) & (!g365) & (g366) & (g367)) + ((!g363) & (!sk[2]) & (g364) & (g365) & (!g366) & (g367)) + ((!g363) & (!sk[2]) & (g364) & (g365) & (g366) & (g367)) + ((!g363) & (sk[2]) & (!g364) & (!g365) & (!g366) & (!g367)) + ((g363) & (!sk[2]) & (!g364) & (!g365) & (!g366) & (!g367)) + ((g363) & (!sk[2]) & (!g364) & (!g365) & (!g366) & (g367)) + ((g363) & (!sk[2]) & (!g364) & (!g365) & (g366) & (!g367)) + ((g363) & (!sk[2]) & (!g364) & (!g365) & (g366) & (g367)) + ((g363) & (!sk[2]) & (!g364) & (g365) & (!g366) & (!g367)) + ((g363) & (!sk[2]) & (!g364) & (g365) & (!g366) & (g367)) + ((g363) & (!sk[2]) & (!g364) & (g365) & (g366) & (!g367)) + ((g363) & (!sk[2]) & (!g364) & (g365) & (g366) & (g367)) + ((g363) & (!sk[2]) & (g364) & (!g365) & (!g366) & (!g367)) + ((g363) & (!sk[2]) & (g364) & (!g365) & (!g366) & (g367)) + ((g363) & (!sk[2]) & (g364) & (!g365) & (g366) & (!g367)) + ((g363) & (!sk[2]) & (g364) & (!g365) & (g366) & (g367)) + ((g363) & (!sk[2]) & (g364) & (g365) & (!g366) & (!g367)) + ((g363) & (!sk[2]) & (g364) & (g365) & (!g366) & (g367)) + ((g363) & (!sk[2]) & (g364) & (g365) & (g366) & (!g367)) + ((g363) & (!sk[2]) & (g364) & (g365) & (g366) & (g367)));
	assign g369 = (((i_8_) & (!sk[3]) & (!g304) & (!g100)) + ((i_8_) & (!sk[3]) & (!g304) & (g100)) + ((i_8_) & (!sk[3]) & (g304) & (!g100)) + ((i_8_) & (!sk[3]) & (g304) & (g100)) + ((i_8_) & (sk[3]) & (g304) & (g100)));
	assign g370 = (((!sk[4]) & (!i_8_) & (!g206) & (g221) & (g135)) + ((!sk[4]) & (!i_8_) & (g206) & (!g221) & (!g135)) + ((!sk[4]) & (!i_8_) & (g206) & (!g221) & (g135)) + ((!sk[4]) & (!i_8_) & (g206) & (g221) & (!g135)) + ((!sk[4]) & (!i_8_) & (g206) & (g221) & (g135)) + ((!sk[4]) & (i_8_) & (!g206) & (g221) & (!g135)) + ((!sk[4]) & (i_8_) & (!g206) & (g221) & (g135)) + ((!sk[4]) & (i_8_) & (g206) & (!g221) & (!g135)) + ((!sk[4]) & (i_8_) & (g206) & (!g221) & (g135)) + ((!sk[4]) & (i_8_) & (g206) & (g221) & (!g135)) + ((!sk[4]) & (i_8_) & (g206) & (g221) & (g135)) + ((sk[4]) & (i_8_) & (!g206) & (!g221) & (g135)) + ((sk[4]) & (i_8_) & (!g206) & (g221) & (g135)) + ((sk[4]) & (i_8_) & (g206) & (!g221) & (g135)));
	assign g371 = (((!sk[5]) & (g220) & (!g112) & (!g316)) + ((!sk[5]) & (g220) & (!g112) & (g316)) + ((!sk[5]) & (g220) & (g112) & (!g316)) + ((!sk[5]) & (g220) & (g112) & (g316)) + ((sk[5]) & (!g220) & (g112) & (g316)) + ((sk[5]) & (g220) & (g112) & (!g316)) + ((sk[5]) & (g220) & (g112) & (g316)));
	assign g372 = (((!i_8_) & (!g88) & (!g135) & (!g316) & (!sk[6]) & (g284)) + ((!i_8_) & (!g88) & (!g135) & (g316) & (!sk[6]) & (g284)) + ((!i_8_) & (!g88) & (!g135) & (g316) & (sk[6]) & (g284)) + ((!i_8_) & (!g88) & (g135) & (!g316) & (!sk[6]) & (g284)) + ((!i_8_) & (!g88) & (g135) & (g316) & (!sk[6]) & (g284)) + ((!i_8_) & (!g88) & (g135) & (g316) & (sk[6]) & (g284)) + ((!i_8_) & (g88) & (!g135) & (!g316) & (!sk[6]) & (g284)) + ((!i_8_) & (g88) & (!g135) & (g316) & (!sk[6]) & (g284)) + ((!i_8_) & (g88) & (!g135) & (g316) & (sk[6]) & (g284)) + ((!i_8_) & (g88) & (g135) & (!g316) & (!sk[6]) & (g284)) + ((!i_8_) & (g88) & (g135) & (g316) & (!sk[6]) & (g284)) + ((!i_8_) & (g88) & (g135) & (g316) & (sk[6]) & (g284)) + ((i_8_) & (!g88) & (!g135) & (!g316) & (!sk[6]) & (!g284)) + ((i_8_) & (!g88) & (!g135) & (!g316) & (!sk[6]) & (g284)) + ((i_8_) & (!g88) & (!g135) & (g316) & (!sk[6]) & (!g284)) + ((i_8_) & (!g88) & (!g135) & (g316) & (!sk[6]) & (g284)) + ((i_8_) & (!g88) & (!g135) & (g316) & (sk[6]) & (g284)) + ((i_8_) & (!g88) & (g135) & (!g316) & (!sk[6]) & (!g284)) + ((i_8_) & (!g88) & (g135) & (!g316) & (!sk[6]) & (g284)) + ((i_8_) & (!g88) & (g135) & (g316) & (!sk[6]) & (!g284)) + ((i_8_) & (!g88) & (g135) & (g316) & (!sk[6]) & (g284)) + ((i_8_) & (!g88) & (g135) & (g316) & (sk[6]) & (!g284)) + ((i_8_) & (!g88) & (g135) & (g316) & (sk[6]) & (g284)) + ((i_8_) & (g88) & (!g135) & (!g316) & (!sk[6]) & (!g284)) + ((i_8_) & (g88) & (!g135) & (!g316) & (!sk[6]) & (g284)) + ((i_8_) & (g88) & (!g135) & (g316) & (!sk[6]) & (!g284)) + ((i_8_) & (g88) & (!g135) & (g316) & (!sk[6]) & (g284)) + ((i_8_) & (g88) & (!g135) & (g316) & (sk[6]) & (!g284)) + ((i_8_) & (g88) & (!g135) & (g316) & (sk[6]) & (g284)) + ((i_8_) & (g88) & (g135) & (!g316) & (!sk[6]) & (!g284)) + ((i_8_) & (g88) & (g135) & (!g316) & (!sk[6]) & (g284)) + ((i_8_) & (g88) & (g135) & (g316) & (!sk[6]) & (!g284)) + ((i_8_) & (g88) & (g135) & (g316) & (!sk[6]) & (g284)) + ((i_8_) & (g88) & (g135) & (g316) & (sk[6]) & (!g284)) + ((i_8_) & (g88) & (g135) & (g316) & (sk[6]) & (g284)));
	assign g373 = (((!g270) & (!g136) & (!g369) & (!g370) & (!g371) & (!g372)) + ((g270) & (!g136) & (!g369) & (!g370) & (!g371) & (!g372)) + ((g270) & (g136) & (!g369) & (!g370) & (!g371) & (!g372)));
	assign g374 = (((!g359) & (!g1754) & (g360) & (g362) & (g368) & (g373)) + ((!g359) & (g1754) & (!g360) & (g362) & (g368) & (g373)) + ((!g359) & (g1754) & (g360) & (g362) & (g368) & (g373)) + ((g359) & (!g1754) & (g360) & (g362) & (g368) & (g373)) + ((g359) & (g1754) & (g360) & (g362) & (g368) & (g373)));
	assign g375 = (((!i_8_) & (!sk[9]) & (!g4) & (g87) & (g182)) + ((!i_8_) & (!sk[9]) & (g4) & (!g87) & (!g182)) + ((!i_8_) & (!sk[9]) & (g4) & (!g87) & (g182)) + ((!i_8_) & (!sk[9]) & (g4) & (g87) & (!g182)) + ((!i_8_) & (!sk[9]) & (g4) & (g87) & (g182)) + ((i_8_) & (!sk[9]) & (!g4) & (g87) & (!g182)) + ((i_8_) & (!sk[9]) & (!g4) & (g87) & (g182)) + ((i_8_) & (!sk[9]) & (g4) & (!g87) & (!g182)) + ((i_8_) & (!sk[9]) & (g4) & (!g87) & (g182)) + ((i_8_) & (!sk[9]) & (g4) & (g87) & (!g182)) + ((i_8_) & (!sk[9]) & (g4) & (g87) & (g182)) + ((i_8_) & (sk[9]) & (g4) & (g87) & (g182)));
	assign g376 = (((!i_11_) & (!sk[10]) & (!i_9_) & (i_15_) & (g375)) + ((!i_11_) & (!sk[10]) & (i_9_) & (!i_15_) & (!g375)) + ((!i_11_) & (!sk[10]) & (i_9_) & (!i_15_) & (g375)) + ((!i_11_) & (!sk[10]) & (i_9_) & (i_15_) & (!g375)) + ((!i_11_) & (!sk[10]) & (i_9_) & (i_15_) & (g375)) + ((!i_11_) & (sk[10]) & (!i_9_) & (i_15_) & (g375)) + ((i_11_) & (!sk[10]) & (!i_9_) & (i_15_) & (!g375)) + ((i_11_) & (!sk[10]) & (!i_9_) & (i_15_) & (g375)) + ((i_11_) & (!sk[10]) & (i_9_) & (!i_15_) & (!g375)) + ((i_11_) & (!sk[10]) & (i_9_) & (!i_15_) & (g375)) + ((i_11_) & (!sk[10]) & (i_9_) & (i_15_) & (!g375)) + ((i_11_) & (!sk[10]) & (i_9_) & (i_15_) & (g375)));
	assign g377 = (((i_8_) & (!sk[11]) & (!g34) & (!g110)) + ((i_8_) & (!sk[11]) & (!g34) & (g110)) + ((i_8_) & (!sk[11]) & (g34) & (!g110)) + ((i_8_) & (!sk[11]) & (g34) & (g110)) + ((i_8_) & (sk[11]) & (g34) & (g110)));
	assign g378 = (((!sk[12]) & (i_11_) & (!g141) & (!g377)) + ((!sk[12]) & (i_11_) & (!g141) & (g377)) + ((!sk[12]) & (i_11_) & (g141) & (!g377)) + ((!sk[12]) & (i_11_) & (g141) & (g377)) + ((sk[12]) & (!i_11_) & (g141) & (g377)));
	assign g379 = (((!sk[13]) & (!g112) & (!g323) & (g191) & (g201)) + ((!sk[13]) & (!g112) & (g323) & (!g191) & (!g201)) + ((!sk[13]) & (!g112) & (g323) & (!g191) & (g201)) + ((!sk[13]) & (!g112) & (g323) & (g191) & (!g201)) + ((!sk[13]) & (!g112) & (g323) & (g191) & (g201)) + ((!sk[13]) & (g112) & (!g323) & (g191) & (!g201)) + ((!sk[13]) & (g112) & (!g323) & (g191) & (g201)) + ((!sk[13]) & (g112) & (g323) & (!g191) & (!g201)) + ((!sk[13]) & (g112) & (g323) & (!g191) & (g201)) + ((!sk[13]) & (g112) & (g323) & (g191) & (!g201)) + ((!sk[13]) & (g112) & (g323) & (g191) & (g201)) + ((sk[13]) & (!g112) & (g323) & (g191) & (!g201)) + ((sk[13]) & (!g112) & (g323) & (g191) & (g201)) + ((sk[13]) & (g112) & (!g323) & (!g191) & (!g201)) + ((sk[13]) & (g112) & (!g323) & (g191) & (!g201)) + ((sk[13]) & (g112) & (g323) & (!g191) & (!g201)) + ((sk[13]) & (g112) & (g323) & (g191) & (!g201)) + ((sk[13]) & (g112) & (g323) & (g191) & (g201)));
	assign g380 = (((!g145) & (!g151) & (!g213) & (!g209) & (!g378) & (!g379)) + ((!g145) & (!g151) & (!g213) & (g209) & (!g378) & (!g379)) + ((!g145) & (!g151) & (g213) & (!g209) & (!g378) & (!g379)) + ((!g145) & (!g151) & (g213) & (g209) & (!g378) & (!g379)) + ((!g145) & (g151) & (!g213) & (!g209) & (!g378) & (!g379)) + ((!g145) & (g151) & (!g213) & (g209) & (!g378) & (!g379)) + ((g145) & (!g151) & (!g213) & (!g209) & (!g378) & (!g379)) + ((g145) & (!g151) & (g213) & (!g209) & (!g378) & (!g379)) + ((g145) & (g151) & (!g213) & (!g209) & (!g378) & (!g379)));
	assign g381 = (((!i_11_) & (!g5) & (!sk[15]) & (!g112) & (!g253) & (g377)) + ((!i_11_) & (!g5) & (!sk[15]) & (!g112) & (g253) & (g377)) + ((!i_11_) & (!g5) & (!sk[15]) & (g112) & (!g253) & (g377)) + ((!i_11_) & (!g5) & (!sk[15]) & (g112) & (g253) & (g377)) + ((!i_11_) & (!g5) & (sk[15]) & (g112) & (g253) & (!g377)) + ((!i_11_) & (!g5) & (sk[15]) & (g112) & (g253) & (g377)) + ((!i_11_) & (g5) & (!sk[15]) & (!g112) & (!g253) & (g377)) + ((!i_11_) & (g5) & (!sk[15]) & (!g112) & (g253) & (g377)) + ((!i_11_) & (g5) & (!sk[15]) & (g112) & (!g253) & (g377)) + ((!i_11_) & (g5) & (!sk[15]) & (g112) & (g253) & (g377)) + ((!i_11_) & (g5) & (sk[15]) & (!g112) & (!g253) & (g377)) + ((!i_11_) & (g5) & (sk[15]) & (!g112) & (g253) & (g377)) + ((!i_11_) & (g5) & (sk[15]) & (g112) & (!g253) & (g377)) + ((!i_11_) & (g5) & (sk[15]) & (g112) & (g253) & (!g377)) + ((!i_11_) & (g5) & (sk[15]) & (g112) & (g253) & (g377)) + ((i_11_) & (!g5) & (!sk[15]) & (!g112) & (!g253) & (!g377)) + ((i_11_) & (!g5) & (!sk[15]) & (!g112) & (!g253) & (g377)) + ((i_11_) & (!g5) & (!sk[15]) & (!g112) & (g253) & (!g377)) + ((i_11_) & (!g5) & (!sk[15]) & (!g112) & (g253) & (g377)) + ((i_11_) & (!g5) & (!sk[15]) & (g112) & (!g253) & (!g377)) + ((i_11_) & (!g5) & (!sk[15]) & (g112) & (!g253) & (g377)) + ((i_11_) & (!g5) & (!sk[15]) & (g112) & (g253) & (!g377)) + ((i_11_) & (!g5) & (!sk[15]) & (g112) & (g253) & (g377)) + ((i_11_) & (!g5) & (sk[15]) & (g112) & (g253) & (!g377)) + ((i_11_) & (!g5) & (sk[15]) & (g112) & (g253) & (g377)) + ((i_11_) & (g5) & (!sk[15]) & (!g112) & (!g253) & (!g377)) + ((i_11_) & (g5) & (!sk[15]) & (!g112) & (!g253) & (g377)) + ((i_11_) & (g5) & (!sk[15]) & (!g112) & (g253) & (!g377)) + ((i_11_) & (g5) & (!sk[15]) & (!g112) & (g253) & (g377)) + ((i_11_) & (g5) & (!sk[15]) & (g112) & (!g253) & (!g377)) + ((i_11_) & (g5) & (!sk[15]) & (g112) & (!g253) & (g377)) + ((i_11_) & (g5) & (!sk[15]) & (g112) & (g253) & (!g377)) + ((i_11_) & (g5) & (!sk[15]) & (g112) & (g253) & (g377)) + ((i_11_) & (g5) & (sk[15]) & (g112) & (g253) & (!g377)) + ((i_11_) & (g5) & (sk[15]) & (g112) & (g253) & (g377)));
	assign g382 = (((!i_5_) & (!i_3_) & (!sk[16]) & (g57) & (g111)) + ((!i_5_) & (i_3_) & (!sk[16]) & (!g57) & (!g111)) + ((!i_5_) & (i_3_) & (!sk[16]) & (!g57) & (g111)) + ((!i_5_) & (i_3_) & (!sk[16]) & (g57) & (!g111)) + ((!i_5_) & (i_3_) & (!sk[16]) & (g57) & (g111)) + ((i_5_) & (!i_3_) & (!sk[16]) & (g57) & (!g111)) + ((i_5_) & (!i_3_) & (!sk[16]) & (g57) & (g111)) + ((i_5_) & (!i_3_) & (sk[16]) & (g57) & (g111)) + ((i_5_) & (i_3_) & (!sk[16]) & (!g57) & (!g111)) + ((i_5_) & (i_3_) & (!sk[16]) & (!g57) & (g111)) + ((i_5_) & (i_3_) & (!sk[16]) & (g57) & (!g111)) + ((i_5_) & (i_3_) & (!sk[16]) & (g57) & (g111)));
	assign g383 = (((!g98) & (!g112) & (!g316) & (!g268) & (!g381) & (!g382)) + ((!g98) & (!g112) & (!g316) & (!g268) & (!g381) & (g382)) + ((!g98) & (!g112) & (!g316) & (g268) & (!g381) & (!g382)) + ((!g98) & (!g112) & (!g316) & (g268) & (!g381) & (g382)) + ((!g98) & (!g112) & (g316) & (!g268) & (!g381) & (!g382)) + ((!g98) & (!g112) & (g316) & (!g268) & (!g381) & (g382)) + ((!g98) & (!g112) & (g316) & (g268) & (!g381) & (!g382)) + ((!g98) & (g112) & (!g316) & (!g268) & (!g381) & (!g382)) + ((!g98) & (g112) & (!g316) & (!g268) & (!g381) & (g382)) + ((!g98) & (g112) & (!g316) & (g268) & (!g381) & (!g382)) + ((!g98) & (g112) & (g316) & (!g268) & (!g381) & (!g382)) + ((!g98) & (g112) & (g316) & (!g268) & (!g381) & (g382)) + ((!g98) & (g112) & (g316) & (g268) & (!g381) & (!g382)) + ((g98) & (!g112) & (!g316) & (!g268) & (!g381) & (!g382)) + ((g98) & (!g112) & (!g316) & (!g268) & (!g381) & (g382)) + ((g98) & (!g112) & (!g316) & (g268) & (!g381) & (!g382)) + ((g98) & (!g112) & (!g316) & (g268) & (!g381) & (g382)) + ((g98) & (!g112) & (g316) & (!g268) & (!g381) & (!g382)) + ((g98) & (!g112) & (g316) & (g268) & (!g381) & (!g382)) + ((g98) & (g112) & (!g316) & (!g268) & (!g381) & (!g382)) + ((g98) & (g112) & (!g316) & (!g268) & (!g381) & (g382)) + ((g98) & (g112) & (!g316) & (g268) & (!g381) & (!g382)) + ((g98) & (g112) & (g316) & (!g268) & (!g381) & (!g382)) + ((g98) & (g112) & (g316) & (g268) & (!g381) & (!g382)));
	assign g384 = (((!i_9_) & (!i_10_) & (!g53) & (!sk[18]) & (!g323) & (g182)) + ((!i_9_) & (!i_10_) & (!g53) & (!sk[18]) & (g323) & (g182)) + ((!i_9_) & (!i_10_) & (g53) & (!sk[18]) & (!g323) & (g182)) + ((!i_9_) & (!i_10_) & (g53) & (!sk[18]) & (g323) & (g182)) + ((!i_9_) & (!i_10_) & (g53) & (sk[18]) & (!g323) & (g182)) + ((!i_9_) & (!i_10_) & (g53) & (sk[18]) & (g323) & (g182)) + ((!i_9_) & (i_10_) & (!g53) & (!sk[18]) & (!g323) & (g182)) + ((!i_9_) & (i_10_) & (!g53) & (!sk[18]) & (g323) & (g182)) + ((!i_9_) & (i_10_) & (g53) & (!sk[18]) & (!g323) & (g182)) + ((!i_9_) & (i_10_) & (g53) & (!sk[18]) & (g323) & (g182)) + ((i_9_) & (!i_10_) & (!g53) & (!sk[18]) & (!g323) & (!g182)) + ((i_9_) & (!i_10_) & (!g53) & (!sk[18]) & (!g323) & (g182)) + ((i_9_) & (!i_10_) & (!g53) & (!sk[18]) & (g323) & (!g182)) + ((i_9_) & (!i_10_) & (!g53) & (!sk[18]) & (g323) & (g182)) + ((i_9_) & (!i_10_) & (g53) & (!sk[18]) & (!g323) & (!g182)) + ((i_9_) & (!i_10_) & (g53) & (!sk[18]) & (!g323) & (g182)) + ((i_9_) & (!i_10_) & (g53) & (!sk[18]) & (g323) & (!g182)) + ((i_9_) & (!i_10_) & (g53) & (!sk[18]) & (g323) & (g182)) + ((i_9_) & (!i_10_) & (g53) & (sk[18]) & (g323) & (g182)) + ((i_9_) & (i_10_) & (!g53) & (!sk[18]) & (!g323) & (!g182)) + ((i_9_) & (i_10_) & (!g53) & (!sk[18]) & (!g323) & (g182)) + ((i_9_) & (i_10_) & (!g53) & (!sk[18]) & (g323) & (!g182)) + ((i_9_) & (i_10_) & (!g53) & (!sk[18]) & (g323) & (g182)) + ((i_9_) & (i_10_) & (g53) & (!sk[18]) & (!g323) & (!g182)) + ((i_9_) & (i_10_) & (g53) & (!sk[18]) & (!g323) & (g182)) + ((i_9_) & (i_10_) & (g53) & (!sk[18]) & (g323) & (!g182)) + ((i_9_) & (i_10_) & (g53) & (!sk[18]) & (g323) & (g182)));
	assign g385 = (((!sk[19]) & (!g323) & (!g151) & (!g209) & (!g284) & (g384)) + ((!sk[19]) & (!g323) & (!g151) & (!g209) & (g284) & (g384)) + ((!sk[19]) & (!g323) & (!g151) & (g209) & (!g284) & (g384)) + ((!sk[19]) & (!g323) & (!g151) & (g209) & (g284) & (g384)) + ((!sk[19]) & (!g323) & (g151) & (!g209) & (!g284) & (g384)) + ((!sk[19]) & (!g323) & (g151) & (!g209) & (g284) & (g384)) + ((!sk[19]) & (!g323) & (g151) & (g209) & (!g284) & (g384)) + ((!sk[19]) & (!g323) & (g151) & (g209) & (g284) & (g384)) + ((!sk[19]) & (g323) & (!g151) & (!g209) & (!g284) & (!g384)) + ((!sk[19]) & (g323) & (!g151) & (!g209) & (!g284) & (g384)) + ((!sk[19]) & (g323) & (!g151) & (!g209) & (g284) & (!g384)) + ((!sk[19]) & (g323) & (!g151) & (!g209) & (g284) & (g384)) + ((!sk[19]) & (g323) & (!g151) & (g209) & (!g284) & (!g384)) + ((!sk[19]) & (g323) & (!g151) & (g209) & (!g284) & (g384)) + ((!sk[19]) & (g323) & (!g151) & (g209) & (g284) & (!g384)) + ((!sk[19]) & (g323) & (!g151) & (g209) & (g284) & (g384)) + ((!sk[19]) & (g323) & (g151) & (!g209) & (!g284) & (!g384)) + ((!sk[19]) & (g323) & (g151) & (!g209) & (!g284) & (g384)) + ((!sk[19]) & (g323) & (g151) & (!g209) & (g284) & (!g384)) + ((!sk[19]) & (g323) & (g151) & (!g209) & (g284) & (g384)) + ((!sk[19]) & (g323) & (g151) & (g209) & (!g284) & (!g384)) + ((!sk[19]) & (g323) & (g151) & (g209) & (!g284) & (g384)) + ((!sk[19]) & (g323) & (g151) & (g209) & (g284) & (!g384)) + ((!sk[19]) & (g323) & (g151) & (g209) & (g284) & (g384)) + ((sk[19]) & (!g323) & (!g151) & (!g209) & (g284) & (g384)) + ((sk[19]) & (!g323) & (!g151) & (g209) & (g284) & (g384)) + ((sk[19]) & (!g323) & (g151) & (!g209) & (!g284) & (g384)) + ((sk[19]) & (!g323) & (g151) & (!g209) & (g284) & (g384)) + ((sk[19]) & (!g323) & (g151) & (g209) & (!g284) & (g384)) + ((sk[19]) & (!g323) & (g151) & (g209) & (g284) & (g384)) + ((sk[19]) & (g323) & (!g151) & (!g209) & (g284) & (g384)) + ((sk[19]) & (g323) & (!g151) & (g209) & (!g284) & (g384)) + ((sk[19]) & (g323) & (!g151) & (g209) & (g284) & (g384)) + ((sk[19]) & (g323) & (g151) & (!g209) & (!g284) & (g384)) + ((sk[19]) & (g323) & (g151) & (!g209) & (g284) & (g384)) + ((sk[19]) & (g323) & (g151) & (g209) & (!g284) & (g384)) + ((sk[19]) & (g323) & (g151) & (g209) & (g284) & (g384)));
	assign g386 = (((!i_8_) & (!g100) & (g191) & (!sk[20]) & (g201)) + ((!i_8_) & (g100) & (!g191) & (!sk[20]) & (!g201)) + ((!i_8_) & (g100) & (!g191) & (!sk[20]) & (g201)) + ((!i_8_) & (g100) & (g191) & (!sk[20]) & (!g201)) + ((!i_8_) & (g100) & (g191) & (!sk[20]) & (g201)) + ((i_8_) & (!g100) & (g191) & (!sk[20]) & (!g201)) + ((i_8_) & (!g100) & (g191) & (!sk[20]) & (g201)) + ((i_8_) & (g100) & (!g191) & (!sk[20]) & (!g201)) + ((i_8_) & (g100) & (!g191) & (!sk[20]) & (g201)) + ((i_8_) & (g100) & (!g191) & (sk[20]) & (!g201)) + ((i_8_) & (g100) & (g191) & (!sk[20]) & (!g201)) + ((i_8_) & (g100) & (g191) & (!sk[20]) & (g201)) + ((i_8_) & (g100) & (g191) & (sk[20]) & (!g201)) + ((i_8_) & (g100) & (g191) & (sk[20]) & (g201)));
	assign g387 = (((!i_8_) & (!g100) & (!sk[21]) & (g193) & (g232)) + ((!i_8_) & (g100) & (!sk[21]) & (!g193) & (!g232)) + ((!i_8_) & (g100) & (!sk[21]) & (!g193) & (g232)) + ((!i_8_) & (g100) & (!sk[21]) & (g193) & (!g232)) + ((!i_8_) & (g100) & (!sk[21]) & (g193) & (g232)) + ((i_8_) & (!g100) & (!sk[21]) & (g193) & (!g232)) + ((i_8_) & (!g100) & (!sk[21]) & (g193) & (g232)) + ((i_8_) & (g100) & (!sk[21]) & (!g193) & (!g232)) + ((i_8_) & (g100) & (!sk[21]) & (!g193) & (g232)) + ((i_8_) & (g100) & (!sk[21]) & (g193) & (!g232)) + ((i_8_) & (g100) & (!sk[21]) & (g193) & (g232)) + ((i_8_) & (g100) & (sk[21]) & (!g193) & (g232)) + ((i_8_) & (g100) & (sk[21]) & (g193) & (!g232)) + ((i_8_) & (g100) & (sk[21]) & (g193) & (g232)));
	assign g388 = (((!i_8_) & (!sk[22]) & (!g135) & (g187) & (g193)) + ((!i_8_) & (!sk[22]) & (g135) & (!g187) & (!g193)) + ((!i_8_) & (!sk[22]) & (g135) & (!g187) & (g193)) + ((!i_8_) & (!sk[22]) & (g135) & (g187) & (!g193)) + ((!i_8_) & (!sk[22]) & (g135) & (g187) & (g193)) + ((i_8_) & (!sk[22]) & (!g135) & (g187) & (!g193)) + ((i_8_) & (!sk[22]) & (!g135) & (g187) & (g193)) + ((i_8_) & (!sk[22]) & (g135) & (!g187) & (!g193)) + ((i_8_) & (!sk[22]) & (g135) & (!g187) & (g193)) + ((i_8_) & (!sk[22]) & (g135) & (g187) & (!g193)) + ((i_8_) & (!sk[22]) & (g135) & (g187) & (g193)) + ((i_8_) & (sk[22]) & (g135) & (!g187) & (g193)) + ((i_8_) & (sk[22]) & (g135) & (g187) & (!g193)) + ((i_8_) & (sk[22]) & (g135) & (g187) & (g193)));
	assign g389 = (((!g112) & (!g183) & (!sk[23]) & (g187) & (g193)) + ((!g112) & (g183) & (!sk[23]) & (!g187) & (!g193)) + ((!g112) & (g183) & (!sk[23]) & (!g187) & (g193)) + ((!g112) & (g183) & (!sk[23]) & (g187) & (!g193)) + ((!g112) & (g183) & (!sk[23]) & (g187) & (g193)) + ((g112) & (!g183) & (!sk[23]) & (g187) & (!g193)) + ((g112) & (!g183) & (!sk[23]) & (g187) & (g193)) + ((g112) & (!g183) & (sk[23]) & (!g187) & (g193)) + ((g112) & (!g183) & (sk[23]) & (g187) & (!g193)) + ((g112) & (!g183) & (sk[23]) & (g187) & (g193)) + ((g112) & (g183) & (!sk[23]) & (!g187) & (!g193)) + ((g112) & (g183) & (!sk[23]) & (!g187) & (g193)) + ((g112) & (g183) & (!sk[23]) & (g187) & (!g193)) + ((g112) & (g183) & (!sk[23]) & (g187) & (g193)) + ((g112) & (g183) & (sk[23]) & (!g187) & (!g193)) + ((g112) & (g183) & (sk[23]) & (!g187) & (g193)) + ((g112) & (g183) & (sk[23]) & (g187) & (!g193)) + ((g112) & (g183) & (sk[23]) & (g187) & (g193)));
	assign g390 = (((!i_8_) & (!g108) & (!g323) & (!g187) & (!g201) & (!g213)) + ((!i_8_) & (!g108) & (!g323) & (!g187) & (!g201) & (g213)) + ((!i_8_) & (!g108) & (!g323) & (!g187) & (g201) & (!g213)) + ((!i_8_) & (!g108) & (!g323) & (!g187) & (g201) & (g213)) + ((!i_8_) & (!g108) & (!g323) & (g187) & (!g201) & (!g213)) + ((!i_8_) & (!g108) & (!g323) & (g187) & (!g201) & (g213)) + ((!i_8_) & (!g108) & (!g323) & (g187) & (g201) & (!g213)) + ((!i_8_) & (!g108) & (!g323) & (g187) & (g201) & (g213)) + ((!i_8_) & (!g108) & (g323) & (!g187) & (g201) & (!g213)) + ((!i_8_) & (g108) & (!g323) & (!g187) & (!g201) & (!g213)) + ((!i_8_) & (g108) & (!g323) & (!g187) & (!g201) & (g213)) + ((!i_8_) & (g108) & (!g323) & (!g187) & (g201) & (!g213)) + ((!i_8_) & (g108) & (!g323) & (!g187) & (g201) & (g213)) + ((!i_8_) & (g108) & (!g323) & (g187) & (!g201) & (!g213)) + ((!i_8_) & (g108) & (!g323) & (g187) & (!g201) & (g213)) + ((!i_8_) & (g108) & (!g323) & (g187) & (g201) & (!g213)) + ((!i_8_) & (g108) & (!g323) & (g187) & (g201) & (g213)) + ((!i_8_) & (g108) & (g323) & (!g187) & (g201) & (!g213)) + ((i_8_) & (!g108) & (!g323) & (!g187) & (!g201) & (!g213)) + ((i_8_) & (!g108) & (!g323) & (!g187) & (!g201) & (g213)) + ((i_8_) & (!g108) & (!g323) & (!g187) & (g201) & (!g213)) + ((i_8_) & (!g108) & (!g323) & (!g187) & (g201) & (g213)) + ((i_8_) & (!g108) & (!g323) & (g187) & (!g201) & (!g213)) + ((i_8_) & (!g108) & (!g323) & (g187) & (!g201) & (g213)) + ((i_8_) & (!g108) & (!g323) & (g187) & (g201) & (!g213)) + ((i_8_) & (!g108) & (!g323) & (g187) & (g201) & (g213)) + ((i_8_) & (!g108) & (g323) & (!g187) & (g201) & (!g213)) + ((i_8_) & (g108) & (!g323) & (!g187) & (!g201) & (!g213)) + ((i_8_) & (g108) & (!g323) & (!g187) & (g201) & (!g213)) + ((i_8_) & (g108) & (g323) & (!g187) & (g201) & (!g213)));
	assign g391 = (((!g386) & (!g387) & (!g388) & (!sk[25]) & (!g389) & (g390)) + ((!g386) & (!g387) & (!g388) & (!sk[25]) & (g389) & (g390)) + ((!g386) & (!g387) & (!g388) & (sk[25]) & (!g389) & (g390)) + ((!g386) & (!g387) & (g388) & (!sk[25]) & (!g389) & (g390)) + ((!g386) & (!g387) & (g388) & (!sk[25]) & (g389) & (g390)) + ((!g386) & (g387) & (!g388) & (!sk[25]) & (!g389) & (g390)) + ((!g386) & (g387) & (!g388) & (!sk[25]) & (g389) & (g390)) + ((!g386) & (g387) & (g388) & (!sk[25]) & (!g389) & (g390)) + ((!g386) & (g387) & (g388) & (!sk[25]) & (g389) & (g390)) + ((g386) & (!g387) & (!g388) & (!sk[25]) & (!g389) & (!g390)) + ((g386) & (!g387) & (!g388) & (!sk[25]) & (!g389) & (g390)) + ((g386) & (!g387) & (!g388) & (!sk[25]) & (g389) & (!g390)) + ((g386) & (!g387) & (!g388) & (!sk[25]) & (g389) & (g390)) + ((g386) & (!g387) & (g388) & (!sk[25]) & (!g389) & (!g390)) + ((g386) & (!g387) & (g388) & (!sk[25]) & (!g389) & (g390)) + ((g386) & (!g387) & (g388) & (!sk[25]) & (g389) & (!g390)) + ((g386) & (!g387) & (g388) & (!sk[25]) & (g389) & (g390)) + ((g386) & (g387) & (!g388) & (!sk[25]) & (!g389) & (!g390)) + ((g386) & (g387) & (!g388) & (!sk[25]) & (!g389) & (g390)) + ((g386) & (g387) & (!g388) & (!sk[25]) & (g389) & (!g390)) + ((g386) & (g387) & (!g388) & (!sk[25]) & (g389) & (g390)) + ((g386) & (g387) & (g388) & (!sk[25]) & (!g389) & (!g390)) + ((g386) & (g387) & (g388) & (!sk[25]) & (!g389) & (g390)) + ((g386) & (g387) & (g388) & (!sk[25]) & (g389) & (!g390)) + ((g386) & (g387) & (g388) & (!sk[25]) & (g389) & (g390)));
	assign g392 = (((!i_8_) & (!g88) & (g193) & (!sk[26]) & (g255)) + ((!i_8_) & (g88) & (!g193) & (!sk[26]) & (!g255)) + ((!i_8_) & (g88) & (!g193) & (!sk[26]) & (g255)) + ((!i_8_) & (g88) & (g193) & (!sk[26]) & (!g255)) + ((!i_8_) & (g88) & (g193) & (!sk[26]) & (g255)) + ((i_8_) & (!g88) & (g193) & (!sk[26]) & (!g255)) + ((i_8_) & (!g88) & (g193) & (!sk[26]) & (g255)) + ((i_8_) & (g88) & (!g193) & (!sk[26]) & (!g255)) + ((i_8_) & (g88) & (!g193) & (!sk[26]) & (g255)) + ((i_8_) & (g88) & (!g193) & (sk[26]) & (g255)) + ((i_8_) & (g88) & (g193) & (!sk[26]) & (!g255)) + ((i_8_) & (g88) & (g193) & (!sk[26]) & (g255)) + ((i_8_) & (g88) & (g193) & (sk[26]) & (!g255)) + ((i_8_) & (g88) & (g193) & (sk[26]) & (g255)));
	assign g393 = (((!i_8_) & (!g100) & (!sk[27]) & (g213) & (g253)) + ((!i_8_) & (g100) & (!sk[27]) & (!g213) & (!g253)) + ((!i_8_) & (g100) & (!sk[27]) & (!g213) & (g253)) + ((!i_8_) & (g100) & (!sk[27]) & (g213) & (!g253)) + ((!i_8_) & (g100) & (!sk[27]) & (g213) & (g253)) + ((i_8_) & (!g100) & (!sk[27]) & (g213) & (!g253)) + ((i_8_) & (!g100) & (!sk[27]) & (g213) & (g253)) + ((i_8_) & (g100) & (!sk[27]) & (!g213) & (!g253)) + ((i_8_) & (g100) & (!sk[27]) & (!g213) & (g253)) + ((i_8_) & (g100) & (!sk[27]) & (g213) & (!g253)) + ((i_8_) & (g100) & (!sk[27]) & (g213) & (g253)) + ((i_8_) & (g100) & (sk[27]) & (!g213) & (g253)) + ((i_8_) & (g100) & (sk[27]) & (g213) & (!g253)) + ((i_8_) & (g100) & (sk[27]) & (g213) & (g253)));
	assign g394 = (((!i_8_) & (!g100) & (!sk[28]) & (g187) & (g231)) + ((!i_8_) & (g100) & (!sk[28]) & (!g187) & (!g231)) + ((!i_8_) & (g100) & (!sk[28]) & (!g187) & (g231)) + ((!i_8_) & (g100) & (!sk[28]) & (g187) & (!g231)) + ((!i_8_) & (g100) & (!sk[28]) & (g187) & (g231)) + ((i_8_) & (!g100) & (!sk[28]) & (g187) & (!g231)) + ((i_8_) & (!g100) & (!sk[28]) & (g187) & (g231)) + ((i_8_) & (g100) & (!sk[28]) & (!g187) & (!g231)) + ((i_8_) & (g100) & (!sk[28]) & (!g187) & (g231)) + ((i_8_) & (g100) & (!sk[28]) & (g187) & (!g231)) + ((i_8_) & (g100) & (!sk[28]) & (g187) & (g231)) + ((i_8_) & (g100) & (sk[28]) & (!g187) & (!g231)) + ((i_8_) & (g100) & (sk[28]) & (g187) & (!g231)) + ((i_8_) & (g100) & (sk[28]) & (g187) & (g231)));
	assign g395 = (((!sk[29]) & (!i_8_) & (!g100) & (g224) & (g349)) + ((!sk[29]) & (!i_8_) & (g100) & (!g224) & (!g349)) + ((!sk[29]) & (!i_8_) & (g100) & (!g224) & (g349)) + ((!sk[29]) & (!i_8_) & (g100) & (g224) & (!g349)) + ((!sk[29]) & (!i_8_) & (g100) & (g224) & (g349)) + ((!sk[29]) & (i_8_) & (!g100) & (g224) & (!g349)) + ((!sk[29]) & (i_8_) & (!g100) & (g224) & (g349)) + ((!sk[29]) & (i_8_) & (g100) & (!g224) & (!g349)) + ((!sk[29]) & (i_8_) & (g100) & (!g224) & (g349)) + ((!sk[29]) & (i_8_) & (g100) & (g224) & (!g349)) + ((!sk[29]) & (i_8_) & (g100) & (g224) & (g349)) + ((sk[29]) & (i_8_) & (g100) & (!g224) & (g349)) + ((sk[29]) & (i_8_) & (g100) & (g224) & (!g349)) + ((sk[29]) & (i_8_) & (g100) & (g224) & (g349)));
	assign g396 = (((!i_8_) & (!g135) & (!g183) & (!g191) & (!g201) & (!g338)) + ((!i_8_) & (!g135) & (!g183) & (g191) & (!g201) & (!g338)) + ((!i_8_) & (!g135) & (!g183) & (g191) & (g201) & (!g338)) + ((!i_8_) & (!g135) & (g183) & (!g191) & (!g201) & (!g338)) + ((!i_8_) & (!g135) & (g183) & (g191) & (!g201) & (!g338)) + ((!i_8_) & (!g135) & (g183) & (g191) & (g201) & (!g338)) + ((!i_8_) & (g135) & (!g183) & (!g191) & (!g201) & (!g338)) + ((!i_8_) & (g135) & (!g183) & (g191) & (!g201) & (!g338)) + ((!i_8_) & (g135) & (!g183) & (g191) & (g201) & (!g338)) + ((!i_8_) & (g135) & (g183) & (!g191) & (!g201) & (!g338)) + ((!i_8_) & (g135) & (g183) & (g191) & (!g201) & (!g338)) + ((!i_8_) & (g135) & (g183) & (g191) & (g201) & (!g338)) + ((i_8_) & (!g135) & (!g183) & (!g191) & (!g201) & (!g338)) + ((i_8_) & (!g135) & (!g183) & (g191) & (!g201) & (!g338)) + ((i_8_) & (!g135) & (!g183) & (g191) & (g201) & (!g338)) + ((i_8_) & (!g135) & (g183) & (!g191) & (!g201) & (!g338)) + ((i_8_) & (!g135) & (g183) & (g191) & (!g201) & (!g338)) + ((i_8_) & (!g135) & (g183) & (g191) & (g201) & (!g338)) + ((i_8_) & (g135) & (!g183) & (!g191) & (!g201) & (!g338)) + ((i_8_) & (g135) & (!g183) & (!g191) & (!g201) & (g338)) + ((i_8_) & (g135) & (!g183) & (g191) & (!g201) & (!g338)) + ((i_8_) & (g135) & (!g183) & (g191) & (!g201) & (g338)) + ((i_8_) & (g135) & (!g183) & (g191) & (g201) & (!g338)) + ((i_8_) & (g135) & (g183) & (!g191) & (!g201) & (!g338)) + ((i_8_) & (g135) & (g183) & (!g191) & (!g201) & (g338)) + ((i_8_) & (g135) & (g183) & (!g191) & (g201) & (!g338)) + ((i_8_) & (g135) & (g183) & (!g191) & (g201) & (g338)) + ((i_8_) & (g135) & (g183) & (g191) & (!g201) & (!g338)) + ((i_8_) & (g135) & (g183) & (g191) & (!g201) & (g338)) + ((i_8_) & (g135) & (g183) & (g191) & (g201) & (!g338)) + ((i_8_) & (g135) & (g183) & (g191) & (g201) & (g338)));
	assign g397 = (((!g392) & (!sk[31]) & (!g393) & (!g394) & (!g395) & (g396)) + ((!g392) & (!sk[31]) & (!g393) & (!g394) & (g395) & (g396)) + ((!g392) & (!sk[31]) & (!g393) & (g394) & (!g395) & (g396)) + ((!g392) & (!sk[31]) & (!g393) & (g394) & (g395) & (g396)) + ((!g392) & (!sk[31]) & (g393) & (!g394) & (!g395) & (g396)) + ((!g392) & (!sk[31]) & (g393) & (!g394) & (g395) & (g396)) + ((!g392) & (!sk[31]) & (g393) & (g394) & (!g395) & (g396)) + ((!g392) & (!sk[31]) & (g393) & (g394) & (g395) & (g396)) + ((!g392) & (sk[31]) & (!g393) & (!g394) & (!g395) & (!g396)) + ((g392) & (!sk[31]) & (!g393) & (!g394) & (!g395) & (!g396)) + ((g392) & (!sk[31]) & (!g393) & (!g394) & (!g395) & (g396)) + ((g392) & (!sk[31]) & (!g393) & (!g394) & (g395) & (!g396)) + ((g392) & (!sk[31]) & (!g393) & (!g394) & (g395) & (g396)) + ((g392) & (!sk[31]) & (!g393) & (g394) & (!g395) & (!g396)) + ((g392) & (!sk[31]) & (!g393) & (g394) & (!g395) & (g396)) + ((g392) & (!sk[31]) & (!g393) & (g394) & (g395) & (!g396)) + ((g392) & (!sk[31]) & (!g393) & (g394) & (g395) & (g396)) + ((g392) & (!sk[31]) & (g393) & (!g394) & (!g395) & (!g396)) + ((g392) & (!sk[31]) & (g393) & (!g394) & (!g395) & (g396)) + ((g392) & (!sk[31]) & (g393) & (!g394) & (g395) & (!g396)) + ((g392) & (!sk[31]) & (g393) & (!g394) & (g395) & (g396)) + ((g392) & (!sk[31]) & (g393) & (g394) & (!g395) & (!g396)) + ((g392) & (!sk[31]) & (g393) & (g394) & (!g395) & (g396)) + ((g392) & (!sk[31]) & (g393) & (g394) & (g395) & (!g396)) + ((g392) & (!sk[31]) & (g393) & (g394) & (g395) & (g396)));
	assign g398 = (((!g376) & (g380) & (g383) & (!g385) & (g391) & (g397)));
	assign g399 = (((!g142) & (sk[33]) & (!g117)) + ((g142) & (!sk[33]) & (!g117)) + ((g142) & (!sk[33]) & (g117)));
	assign g400 = (((i_6_) & (!sk[34]) & (!g58)) + ((i_6_) & (!sk[34]) & (g58)) + ((i_6_) & (sk[34]) & (g58)));
	assign g401 = (((i_8_) & (!g88) & (!g132) & (!g94) & (!g165) & (g400)) + ((i_8_) & (!g88) & (!g132) & (!g94) & (g165) & (g400)) + ((i_8_) & (!g88) & (!g132) & (g94) & (!g165) & (g400)) + ((i_8_) & (!g88) & (!g132) & (g94) & (g165) & (g400)) + ((i_8_) & (g88) & (!g132) & (!g94) & (!g165) & (!g400)) + ((i_8_) & (g88) & (!g132) & (!g94) & (!g165) & (g400)) + ((i_8_) & (g88) & (!g132) & (!g94) & (g165) & (!g400)) + ((i_8_) & (g88) & (!g132) & (!g94) & (g165) & (g400)) + ((i_8_) & (g88) & (!g132) & (g94) & (!g165) & (!g400)) + ((i_8_) & (g88) & (!g132) & (g94) & (!g165) & (g400)) + ((i_8_) & (g88) & (!g132) & (g94) & (g165) & (!g400)) + ((i_8_) & (g88) & (!g132) & (g94) & (g165) & (g400)) + ((i_8_) & (g88) & (g132) & (!g94) & (g165) & (!g400)) + ((i_8_) & (g88) & (g132) & (!g94) & (g165) & (g400)) + ((i_8_) & (g88) & (g132) & (g94) & (!g165) & (!g400)) + ((i_8_) & (g88) & (g132) & (g94) & (!g165) & (g400)) + ((i_8_) & (g88) & (g132) & (g94) & (g165) & (!g400)) + ((i_8_) & (g88) & (g132) & (g94) & (g165) & (g400)));
	assign g402 = (((!g136) & (!g399) & (sk[36]) & (!g401)) + ((!g136) & (g399) & (sk[36]) & (!g401)) + ((g136) & (!g399) & (!sk[36]) & (!g401)) + ((g136) & (!g399) & (!sk[36]) & (g401)) + ((g136) & (g399) & (!sk[36]) & (!g401)) + ((g136) & (g399) & (!sk[36]) & (g401)) + ((g136) & (g399) & (sk[36]) & (!g401)));
	assign g403 = (((i_8_) & (!g88) & (g135) & (!g159) & (!g92) & (!g96)) + ((i_8_) & (!g88) & (g135) & (!g159) & (g92) & (!g96)) + ((i_8_) & (!g88) & (g135) & (g159) & (!g92) & (!g96)) + ((i_8_) & (!g88) & (g135) & (g159) & (!g92) & (g96)) + ((i_8_) & (!g88) & (g135) & (g159) & (g92) & (!g96)) + ((i_8_) & (!g88) & (g135) & (g159) & (g92) & (g96)) + ((i_8_) & (g88) & (!g135) & (!g159) & (!g92) & (!g96)) + ((i_8_) & (g88) & (!g135) & (!g159) & (!g92) & (g96)) + ((i_8_) & (g88) & (!g135) & (g159) & (!g92) & (!g96)) + ((i_8_) & (g88) & (!g135) & (g159) & (!g92) & (g96)) + ((i_8_) & (g88) & (!g135) & (g159) & (g92) & (!g96)) + ((i_8_) & (g88) & (!g135) & (g159) & (g92) & (g96)) + ((i_8_) & (g88) & (g135) & (!g159) & (!g92) & (!g96)) + ((i_8_) & (g88) & (g135) & (!g159) & (!g92) & (g96)) + ((i_8_) & (g88) & (g135) & (!g159) & (g92) & (!g96)) + ((i_8_) & (g88) & (g135) & (g159) & (!g92) & (!g96)) + ((i_8_) & (g88) & (g135) & (g159) & (!g92) & (g96)) + ((i_8_) & (g88) & (g135) & (g159) & (g92) & (!g96)) + ((i_8_) & (g88) & (g135) & (g159) & (g92) & (g96)));
	assign g404 = (((!sk[38]) & (!g101) & (!g112) & (!g103) & (!g96) & (g403)) + ((!sk[38]) & (!g101) & (!g112) & (!g103) & (g96) & (g403)) + ((!sk[38]) & (!g101) & (!g112) & (g103) & (!g96) & (g403)) + ((!sk[38]) & (!g101) & (!g112) & (g103) & (g96) & (g403)) + ((!sk[38]) & (!g101) & (g112) & (!g103) & (!g96) & (g403)) + ((!sk[38]) & (!g101) & (g112) & (!g103) & (g96) & (g403)) + ((!sk[38]) & (!g101) & (g112) & (g103) & (!g96) & (g403)) + ((!sk[38]) & (!g101) & (g112) & (g103) & (g96) & (g403)) + ((!sk[38]) & (g101) & (!g112) & (!g103) & (!g96) & (!g403)) + ((!sk[38]) & (g101) & (!g112) & (!g103) & (!g96) & (g403)) + ((!sk[38]) & (g101) & (!g112) & (!g103) & (g96) & (!g403)) + ((!sk[38]) & (g101) & (!g112) & (!g103) & (g96) & (g403)) + ((!sk[38]) & (g101) & (!g112) & (g103) & (!g96) & (!g403)) + ((!sk[38]) & (g101) & (!g112) & (g103) & (!g96) & (g403)) + ((!sk[38]) & (g101) & (!g112) & (g103) & (g96) & (!g403)) + ((!sk[38]) & (g101) & (!g112) & (g103) & (g96) & (g403)) + ((!sk[38]) & (g101) & (g112) & (!g103) & (!g96) & (!g403)) + ((!sk[38]) & (g101) & (g112) & (!g103) & (!g96) & (g403)) + ((!sk[38]) & (g101) & (g112) & (!g103) & (g96) & (!g403)) + ((!sk[38]) & (g101) & (g112) & (!g103) & (g96) & (g403)) + ((!sk[38]) & (g101) & (g112) & (g103) & (!g96) & (!g403)) + ((!sk[38]) & (g101) & (g112) & (g103) & (!g96) & (g403)) + ((!sk[38]) & (g101) & (g112) & (g103) & (g96) & (!g403)) + ((!sk[38]) & (g101) & (g112) & (g103) & (g96) & (g403)) + ((sk[38]) & (!g101) & (!g112) & (!g103) & (!g96) & (!g403)) + ((sk[38]) & (!g101) & (!g112) & (!g103) & (g96) & (!g403)) + ((sk[38]) & (!g101) & (!g112) & (g103) & (!g96) & (!g403)) + ((sk[38]) & (!g101) & (!g112) & (g103) & (g96) & (!g403)) + ((sk[38]) & (!g101) & (g112) & (g103) & (!g96) & (!g403)) + ((sk[38]) & (!g101) & (g112) & (g103) & (g96) & (!g403)) + ((sk[38]) & (g101) & (!g112) & (!g103) & (g96) & (!g403)) + ((sk[38]) & (g101) & (!g112) & (g103) & (g96) & (!g403)) + ((sk[38]) & (g101) & (g112) & (g103) & (g96) & (!g403)));
	assign g405 = (((!sk[39]) & (g112) & (!g132) & (!g159)) + ((!sk[39]) & (g112) & (!g132) & (g159)) + ((!sk[39]) & (g112) & (g132) & (!g159)) + ((!sk[39]) & (g112) & (g132) & (g159)) + ((sk[39]) & (g112) & (!g132) & (!g159)) + ((sk[39]) & (g112) & (!g132) & (g159)) + ((sk[39]) & (g112) & (g132) & (g159)));
	assign g406 = (((!sk[40]) & (!i_8_) & (!g108) & (g94) & (g116)) + ((!sk[40]) & (!i_8_) & (g108) & (!g94) & (!g116)) + ((!sk[40]) & (!i_8_) & (g108) & (!g94) & (g116)) + ((!sk[40]) & (!i_8_) & (g108) & (g94) & (!g116)) + ((!sk[40]) & (!i_8_) & (g108) & (g94) & (g116)) + ((!sk[40]) & (i_8_) & (!g108) & (g94) & (!g116)) + ((!sk[40]) & (i_8_) & (!g108) & (g94) & (g116)) + ((!sk[40]) & (i_8_) & (g108) & (!g94) & (!g116)) + ((!sk[40]) & (i_8_) & (g108) & (!g94) & (g116)) + ((!sk[40]) & (i_8_) & (g108) & (g94) & (!g116)) + ((!sk[40]) & (i_8_) & (g108) & (g94) & (g116)) + ((sk[40]) & (i_8_) & (g108) & (!g94) & (g116)) + ((sk[40]) & (i_8_) & (g108) & (g94) & (!g116)) + ((sk[40]) & (i_8_) & (g108) & (g94) & (g116)));
	assign g407 = (((!i_8_) & (!sk[41]) & (!g100) & (g108) & (g132)) + ((!i_8_) & (!sk[41]) & (g100) & (!g108) & (!g132)) + ((!i_8_) & (!sk[41]) & (g100) & (!g108) & (g132)) + ((!i_8_) & (!sk[41]) & (g100) & (g108) & (!g132)) + ((!i_8_) & (!sk[41]) & (g100) & (g108) & (g132)) + ((i_8_) & (!sk[41]) & (!g100) & (g108) & (!g132)) + ((i_8_) & (!sk[41]) & (!g100) & (g108) & (g132)) + ((i_8_) & (!sk[41]) & (g100) & (!g108) & (!g132)) + ((i_8_) & (!sk[41]) & (g100) & (!g108) & (g132)) + ((i_8_) & (!sk[41]) & (g100) & (g108) & (!g132)) + ((i_8_) & (!sk[41]) & (g100) & (g108) & (g132)) + ((i_8_) & (sk[41]) & (!g100) & (g108) & (!g132)) + ((i_8_) & (sk[41]) & (g100) & (!g108) & (!g132)) + ((i_8_) & (sk[41]) & (g100) & (g108) & (!g132)));
	assign g408 = (((g112) & (!sk[42]) & (!g94) & (!g92)) + ((g112) & (!sk[42]) & (!g94) & (g92)) + ((g112) & (!sk[42]) & (g94) & (!g92)) + ((g112) & (!sk[42]) & (g94) & (g92)) + ((g112) & (sk[42]) & (!g94) & (!g92)) + ((g112) & (sk[42]) & (g94) & (!g92)) + ((g112) & (sk[42]) & (g94) & (g92)));
	assign g409 = (((!sk[43]) & (!i_8_) & (!g112) & (!g135) & (!g142) & (g90)) + ((!sk[43]) & (!i_8_) & (!g112) & (!g135) & (g142) & (g90)) + ((!sk[43]) & (!i_8_) & (!g112) & (g135) & (!g142) & (g90)) + ((!sk[43]) & (!i_8_) & (!g112) & (g135) & (g142) & (g90)) + ((!sk[43]) & (!i_8_) & (g112) & (!g135) & (!g142) & (g90)) + ((!sk[43]) & (!i_8_) & (g112) & (!g135) & (g142) & (g90)) + ((!sk[43]) & (!i_8_) & (g112) & (g135) & (!g142) & (g90)) + ((!sk[43]) & (!i_8_) & (g112) & (g135) & (g142) & (g90)) + ((!sk[43]) & (i_8_) & (!g112) & (!g135) & (!g142) & (!g90)) + ((!sk[43]) & (i_8_) & (!g112) & (!g135) & (!g142) & (g90)) + ((!sk[43]) & (i_8_) & (!g112) & (!g135) & (g142) & (!g90)) + ((!sk[43]) & (i_8_) & (!g112) & (!g135) & (g142) & (g90)) + ((!sk[43]) & (i_8_) & (!g112) & (g135) & (!g142) & (!g90)) + ((!sk[43]) & (i_8_) & (!g112) & (g135) & (!g142) & (g90)) + ((!sk[43]) & (i_8_) & (!g112) & (g135) & (g142) & (!g90)) + ((!sk[43]) & (i_8_) & (!g112) & (g135) & (g142) & (g90)) + ((!sk[43]) & (i_8_) & (g112) & (!g135) & (!g142) & (!g90)) + ((!sk[43]) & (i_8_) & (g112) & (!g135) & (!g142) & (g90)) + ((!sk[43]) & (i_8_) & (g112) & (!g135) & (g142) & (!g90)) + ((!sk[43]) & (i_8_) & (g112) & (!g135) & (g142) & (g90)) + ((!sk[43]) & (i_8_) & (g112) & (g135) & (!g142) & (!g90)) + ((!sk[43]) & (i_8_) & (g112) & (g135) & (!g142) & (g90)) + ((!sk[43]) & (i_8_) & (g112) & (g135) & (g142) & (!g90)) + ((!sk[43]) & (i_8_) & (g112) & (g135) & (g142) & (g90)) + ((sk[43]) & (!i_8_) & (g112) & (!g135) & (!g142) & (!g90)) + ((sk[43]) & (!i_8_) & (g112) & (!g135) & (g142) & (!g90)) + ((sk[43]) & (!i_8_) & (g112) & (!g135) & (g142) & (g90)) + ((sk[43]) & (!i_8_) & (g112) & (g135) & (!g142) & (!g90)) + ((sk[43]) & (!i_8_) & (g112) & (g135) & (g142) & (!g90)) + ((sk[43]) & (!i_8_) & (g112) & (g135) & (g142) & (g90)) + ((sk[43]) & (i_8_) & (!g112) & (g135) & (!g142) & (!g90)) + ((sk[43]) & (i_8_) & (!g112) & (g135) & (g142) & (!g90)) + ((sk[43]) & (i_8_) & (g112) & (!g135) & (!g142) & (!g90)) + ((sk[43]) & (i_8_) & (g112) & (!g135) & (g142) & (!g90)) + ((sk[43]) & (i_8_) & (g112) & (!g135) & (g142) & (g90)) + ((sk[43]) & (i_8_) & (g112) & (g135) & (!g142) & (!g90)) + ((sk[43]) & (i_8_) & (g112) & (g135) & (g142) & (!g90)) + ((sk[43]) & (i_8_) & (g112) & (g135) & (g142) & (g90)));
	assign g410 = (((!g405) & (!g406) & (!g407) & (!g408) & (!sk[44]) & (g409)) + ((!g405) & (!g406) & (!g407) & (!g408) & (sk[44]) & (!g409)) + ((!g405) & (!g406) & (!g407) & (g408) & (!sk[44]) & (g409)) + ((!g405) & (!g406) & (g407) & (!g408) & (!sk[44]) & (g409)) + ((!g405) & (!g406) & (g407) & (g408) & (!sk[44]) & (g409)) + ((!g405) & (g406) & (!g407) & (!g408) & (!sk[44]) & (g409)) + ((!g405) & (g406) & (!g407) & (g408) & (!sk[44]) & (g409)) + ((!g405) & (g406) & (g407) & (!g408) & (!sk[44]) & (g409)) + ((!g405) & (g406) & (g407) & (g408) & (!sk[44]) & (g409)) + ((g405) & (!g406) & (!g407) & (!g408) & (!sk[44]) & (!g409)) + ((g405) & (!g406) & (!g407) & (!g408) & (!sk[44]) & (g409)) + ((g405) & (!g406) & (!g407) & (g408) & (!sk[44]) & (!g409)) + ((g405) & (!g406) & (!g407) & (g408) & (!sk[44]) & (g409)) + ((g405) & (!g406) & (g407) & (!g408) & (!sk[44]) & (!g409)) + ((g405) & (!g406) & (g407) & (!g408) & (!sk[44]) & (g409)) + ((g405) & (!g406) & (g407) & (g408) & (!sk[44]) & (!g409)) + ((g405) & (!g406) & (g407) & (g408) & (!sk[44]) & (g409)) + ((g405) & (g406) & (!g407) & (!g408) & (!sk[44]) & (!g409)) + ((g405) & (g406) & (!g407) & (!g408) & (!sk[44]) & (g409)) + ((g405) & (g406) & (!g407) & (g408) & (!sk[44]) & (!g409)) + ((g405) & (g406) & (!g407) & (g408) & (!sk[44]) & (g409)) + ((g405) & (g406) & (g407) & (!g408) & (!sk[44]) & (!g409)) + ((g405) & (g406) & (g407) & (!g408) & (!sk[44]) & (g409)) + ((g405) & (g406) & (g407) & (g408) & (!sk[44]) & (!g409)) + ((g405) & (g406) & (g407) & (g408) & (!sk[44]) & (g409)));
	assign g411 = (((!g338) & (g399) & (g402) & (g404) & (g410) & (g1747)) + ((g338) & (!g399) & (g402) & (g404) & (g410) & (g1747)) + ((g338) & (g399) & (g402) & (g404) & (g410) & (g1747)));
	assign g412 = (((!g15) & (!g91) & (!g131) & (!g182) & (!sk[46]) & (g268)) + ((!g15) & (!g91) & (!g131) & (!g182) & (sk[46]) & (!g268)) + ((!g15) & (!g91) & (!g131) & (g182) & (!sk[46]) & (g268)) + ((!g15) & (!g91) & (g131) & (!g182) & (!sk[46]) & (g268)) + ((!g15) & (!g91) & (g131) & (g182) & (!sk[46]) & (g268)) + ((!g15) & (g91) & (!g131) & (!g182) & (!sk[46]) & (g268)) + ((!g15) & (g91) & (!g131) & (!g182) & (sk[46]) & (!g268)) + ((!g15) & (g91) & (!g131) & (g182) & (!sk[46]) & (g268)) + ((!g15) & (g91) & (g131) & (!g182) & (!sk[46]) & (g268)) + ((!g15) & (g91) & (g131) & (!g182) & (sk[46]) & (!g268)) + ((!g15) & (g91) & (g131) & (g182) & (!sk[46]) & (g268)) + ((g15) & (!g91) & (!g131) & (!g182) & (!sk[46]) & (!g268)) + ((g15) & (!g91) & (!g131) & (!g182) & (!sk[46]) & (g268)) + ((g15) & (!g91) & (!g131) & (!g182) & (sk[46]) & (!g268)) + ((g15) & (!g91) & (!g131) & (g182) & (!sk[46]) & (!g268)) + ((g15) & (!g91) & (!g131) & (g182) & (!sk[46]) & (g268)) + ((g15) & (!g91) & (!g131) & (g182) & (sk[46]) & (!g268)) + ((g15) & (!g91) & (g131) & (!g182) & (!sk[46]) & (!g268)) + ((g15) & (!g91) & (g131) & (!g182) & (!sk[46]) & (g268)) + ((g15) & (!g91) & (g131) & (g182) & (!sk[46]) & (!g268)) + ((g15) & (!g91) & (g131) & (g182) & (!sk[46]) & (g268)) + ((g15) & (g91) & (!g131) & (!g182) & (!sk[46]) & (!g268)) + ((g15) & (g91) & (!g131) & (!g182) & (!sk[46]) & (g268)) + ((g15) & (g91) & (!g131) & (!g182) & (sk[46]) & (!g268)) + ((g15) & (g91) & (!g131) & (g182) & (!sk[46]) & (!g268)) + ((g15) & (g91) & (!g131) & (g182) & (!sk[46]) & (g268)) + ((g15) & (g91) & (!g131) & (g182) & (sk[46]) & (!g268)) + ((g15) & (g91) & (g131) & (!g182) & (!sk[46]) & (!g268)) + ((g15) & (g91) & (g131) & (!g182) & (!sk[46]) & (g268)) + ((g15) & (g91) & (g131) & (!g182) & (sk[46]) & (!g268)) + ((g15) & (g91) & (g131) & (g182) & (!sk[46]) & (!g268)) + ((g15) & (g91) & (g131) & (g182) & (!sk[46]) & (g268)));
	assign g413 = (((!sk[47]) & (i_8_) & (!g135) & (!g172)) + ((!sk[47]) & (i_8_) & (!g135) & (g172)) + ((!sk[47]) & (i_8_) & (g135) & (!g172)) + ((!sk[47]) & (i_8_) & (g135) & (g172)) + ((sk[47]) & (i_8_) & (g135) & (g172)));
	assign g414 = (((!sk[48]) & (!i_8_) & (!g108) & (g349) & (g339)) + ((!sk[48]) & (!i_8_) & (g108) & (!g349) & (!g339)) + ((!sk[48]) & (!i_8_) & (g108) & (!g349) & (g339)) + ((!sk[48]) & (!i_8_) & (g108) & (g349) & (!g339)) + ((!sk[48]) & (!i_8_) & (g108) & (g349) & (g339)) + ((!sk[48]) & (i_8_) & (!g108) & (g349) & (!g339)) + ((!sk[48]) & (i_8_) & (!g108) & (g349) & (g339)) + ((!sk[48]) & (i_8_) & (g108) & (!g349) & (!g339)) + ((!sk[48]) & (i_8_) & (g108) & (!g349) & (g339)) + ((!sk[48]) & (i_8_) & (g108) & (g349) & (!g339)) + ((!sk[48]) & (i_8_) & (g108) & (g349) & (g339)) + ((sk[48]) & (i_8_) & (g108) & (!g349) & (g339)) + ((sk[48]) & (i_8_) & (g108) & (g349) & (!g339)) + ((sk[48]) & (i_8_) & (g108) & (g349) & (g339)));
	assign g415 = (((!i_14_) & (i_12_) & (!i_13_) & (g95) & (!g112) & (g323)) + ((!i_14_) & (i_12_) & (!i_13_) & (g95) & (g112) & (g323)) + ((i_14_) & (!i_12_) & (!i_13_) & (g95) & (g112) & (!g323)) + ((i_14_) & (!i_12_) & (!i_13_) & (g95) & (g112) & (g323)) + ((i_14_) & (!i_12_) & (i_13_) & (g95) & (!g112) & (g323)) + ((i_14_) & (!i_12_) & (i_13_) & (g95) & (g112) & (!g323)) + ((i_14_) & (!i_12_) & (i_13_) & (g95) & (g112) & (g323)));
	assign g416 = (((!i_8_) & (!g100) & (!g135) & (!g94) & (!sk[50]) & (g127)) + ((!i_8_) & (!g100) & (!g135) & (g94) & (!sk[50]) & (g127)) + ((!i_8_) & (!g100) & (g135) & (!g94) & (!sk[50]) & (g127)) + ((!i_8_) & (!g100) & (g135) & (g94) & (!sk[50]) & (g127)) + ((!i_8_) & (g100) & (!g135) & (!g94) & (!sk[50]) & (g127)) + ((!i_8_) & (g100) & (!g135) & (g94) & (!sk[50]) & (g127)) + ((!i_8_) & (g100) & (g135) & (!g94) & (!sk[50]) & (g127)) + ((!i_8_) & (g100) & (g135) & (g94) & (!sk[50]) & (g127)) + ((i_8_) & (!g100) & (!g135) & (!g94) & (!sk[50]) & (!g127)) + ((i_8_) & (!g100) & (!g135) & (!g94) & (!sk[50]) & (g127)) + ((i_8_) & (!g100) & (!g135) & (g94) & (!sk[50]) & (!g127)) + ((i_8_) & (!g100) & (!g135) & (g94) & (!sk[50]) & (g127)) + ((i_8_) & (!g100) & (g135) & (!g94) & (!sk[50]) & (!g127)) + ((i_8_) & (!g100) & (g135) & (!g94) & (!sk[50]) & (g127)) + ((i_8_) & (!g100) & (g135) & (!g94) & (sk[50]) & (!g127)) + ((i_8_) & (!g100) & (g135) & (g94) & (!sk[50]) & (!g127)) + ((i_8_) & (!g100) & (g135) & (g94) & (!sk[50]) & (g127)) + ((i_8_) & (!g100) & (g135) & (g94) & (sk[50]) & (!g127)) + ((i_8_) & (g100) & (!g135) & (!g94) & (!sk[50]) & (!g127)) + ((i_8_) & (g100) & (!g135) & (!g94) & (!sk[50]) & (g127)) + ((i_8_) & (g100) & (!g135) & (g94) & (!sk[50]) & (!g127)) + ((i_8_) & (g100) & (!g135) & (g94) & (!sk[50]) & (g127)) + ((i_8_) & (g100) & (!g135) & (g94) & (sk[50]) & (!g127)) + ((i_8_) & (g100) & (!g135) & (g94) & (sk[50]) & (g127)) + ((i_8_) & (g100) & (g135) & (!g94) & (!sk[50]) & (!g127)) + ((i_8_) & (g100) & (g135) & (!g94) & (!sk[50]) & (g127)) + ((i_8_) & (g100) & (g135) & (!g94) & (sk[50]) & (!g127)) + ((i_8_) & (g100) & (g135) & (g94) & (!sk[50]) & (!g127)) + ((i_8_) & (g100) & (g135) & (g94) & (!sk[50]) & (g127)) + ((i_8_) & (g100) & (g135) & (g94) & (sk[50]) & (!g127)) + ((i_8_) & (g100) & (g135) & (g94) & (sk[50]) & (g127)));
	assign g417 = (((!g151) & (!g280) & (!g413) & (!g414) & (!g415) & (!g416)) + ((!g151) & (g280) & (!g413) & (!g414) & (!g415) & (!g416)) + ((g151) & (!g280) & (!g413) & (!g414) & (!g415) & (!g416)));
	assign g418 = (((!i_9_) & (!i_10_) & (g53) & (g145) & (!g146) & (g182)) + ((!i_9_) & (!i_10_) & (g53) & (g145) & (g146) & (g182)) + ((!i_9_) & (i_10_) & (g53) & (!g145) & (!g146) & (g182)) + ((!i_9_) & (i_10_) & (g53) & (g145) & (!g146) & (g182)));
	assign g419 = (((!g136) & (!g412) & (!sk[53]) & (g417) & (g418)) + ((!g136) & (!g412) & (sk[53]) & (g417) & (!g418)) + ((!g136) & (g412) & (!sk[53]) & (!g417) & (!g418)) + ((!g136) & (g412) & (!sk[53]) & (!g417) & (g418)) + ((!g136) & (g412) & (!sk[53]) & (g417) & (!g418)) + ((!g136) & (g412) & (!sk[53]) & (g417) & (g418)) + ((!g136) & (g412) & (sk[53]) & (g417) & (!g418)) + ((g136) & (!g412) & (!sk[53]) & (g417) & (!g418)) + ((g136) & (!g412) & (!sk[53]) & (g417) & (g418)) + ((g136) & (g412) & (!sk[53]) & (!g417) & (!g418)) + ((g136) & (g412) & (!sk[53]) & (!g417) & (g418)) + ((g136) & (g412) & (!sk[53]) & (g417) & (!g418)) + ((g136) & (g412) & (!sk[53]) & (g417) & (g418)) + ((g136) & (g412) & (sk[53]) & (g417) & (!g418)));
	assign g420 = (((!sk[54]) & (!g358) & (!g374) & (!g398) & (!g411) & (g419)) + ((!sk[54]) & (!g358) & (!g374) & (!g398) & (g411) & (g419)) + ((!sk[54]) & (!g358) & (!g374) & (g398) & (!g411) & (g419)) + ((!sk[54]) & (!g358) & (!g374) & (g398) & (g411) & (g419)) + ((!sk[54]) & (!g358) & (g374) & (!g398) & (!g411) & (g419)) + ((!sk[54]) & (!g358) & (g374) & (!g398) & (g411) & (g419)) + ((!sk[54]) & (!g358) & (g374) & (g398) & (!g411) & (g419)) + ((!sk[54]) & (!g358) & (g374) & (g398) & (g411) & (g419)) + ((!sk[54]) & (g358) & (!g374) & (!g398) & (!g411) & (!g419)) + ((!sk[54]) & (g358) & (!g374) & (!g398) & (!g411) & (g419)) + ((!sk[54]) & (g358) & (!g374) & (!g398) & (g411) & (!g419)) + ((!sk[54]) & (g358) & (!g374) & (!g398) & (g411) & (g419)) + ((!sk[54]) & (g358) & (!g374) & (g398) & (!g411) & (!g419)) + ((!sk[54]) & (g358) & (!g374) & (g398) & (!g411) & (g419)) + ((!sk[54]) & (g358) & (!g374) & (g398) & (g411) & (!g419)) + ((!sk[54]) & (g358) & (!g374) & (g398) & (g411) & (g419)) + ((!sk[54]) & (g358) & (g374) & (!g398) & (!g411) & (!g419)) + ((!sk[54]) & (g358) & (g374) & (!g398) & (!g411) & (g419)) + ((!sk[54]) & (g358) & (g374) & (!g398) & (g411) & (!g419)) + ((!sk[54]) & (g358) & (g374) & (!g398) & (g411) & (g419)) + ((!sk[54]) & (g358) & (g374) & (g398) & (!g411) & (!g419)) + ((!sk[54]) & (g358) & (g374) & (g398) & (!g411) & (g419)) + ((!sk[54]) & (g358) & (g374) & (g398) & (g411) & (!g419)) + ((!sk[54]) & (g358) & (g374) & (g398) & (g411) & (g419)) + ((sk[54]) & (g358) & (g374) & (g398) & (g411) & (g419)));
	assign g421 = (((!g203) & (!g199) & (!g224) & (!g177) & (!sk[55]) & (g339)) + ((!g203) & (!g199) & (!g224) & (!g177) & (sk[55]) & (!g339)) + ((!g203) & (!g199) & (!g224) & (g177) & (!sk[55]) & (g339)) + ((!g203) & (!g199) & (g224) & (!g177) & (!sk[55]) & (g339)) + ((!g203) & (!g199) & (g224) & (g177) & (!sk[55]) & (g339)) + ((!g203) & (g199) & (!g224) & (!g177) & (!sk[55]) & (g339)) + ((!g203) & (g199) & (!g224) & (g177) & (!sk[55]) & (g339)) + ((!g203) & (g199) & (g224) & (!g177) & (!sk[55]) & (g339)) + ((!g203) & (g199) & (g224) & (g177) & (!sk[55]) & (g339)) + ((g203) & (!g199) & (!g224) & (!g177) & (!sk[55]) & (!g339)) + ((g203) & (!g199) & (!g224) & (!g177) & (!sk[55]) & (g339)) + ((g203) & (!g199) & (!g224) & (g177) & (!sk[55]) & (!g339)) + ((g203) & (!g199) & (!g224) & (g177) & (!sk[55]) & (g339)) + ((g203) & (!g199) & (g224) & (!g177) & (!sk[55]) & (!g339)) + ((g203) & (!g199) & (g224) & (!g177) & (!sk[55]) & (g339)) + ((g203) & (!g199) & (g224) & (g177) & (!sk[55]) & (!g339)) + ((g203) & (!g199) & (g224) & (g177) & (!sk[55]) & (g339)) + ((g203) & (g199) & (!g224) & (!g177) & (!sk[55]) & (!g339)) + ((g203) & (g199) & (!g224) & (!g177) & (!sk[55]) & (g339)) + ((g203) & (g199) & (!g224) & (g177) & (!sk[55]) & (!g339)) + ((g203) & (g199) & (!g224) & (g177) & (!sk[55]) & (g339)) + ((g203) & (g199) & (g224) & (!g177) & (!sk[55]) & (!g339)) + ((g203) & (g199) & (g224) & (!g177) & (!sk[55]) & (g339)) + ((g203) & (g199) & (g224) & (g177) & (!sk[55]) & (!g339)) + ((g203) & (g199) & (g224) & (g177) & (!sk[55]) & (g339)));
	assign g422 = (((!g134) & (!sk[56]) & (!g109) & (!g172) & (!g349) & (g421)) + ((!g134) & (!sk[56]) & (!g109) & (!g172) & (g349) & (g421)) + ((!g134) & (!sk[56]) & (!g109) & (g172) & (!g349) & (g421)) + ((!g134) & (!sk[56]) & (!g109) & (g172) & (g349) & (g421)) + ((!g134) & (!sk[56]) & (g109) & (!g172) & (!g349) & (g421)) + ((!g134) & (!sk[56]) & (g109) & (!g172) & (g349) & (g421)) + ((!g134) & (!sk[56]) & (g109) & (g172) & (!g349) & (g421)) + ((!g134) & (!sk[56]) & (g109) & (g172) & (g349) & (g421)) + ((!g134) & (sk[56]) & (!g109) & (!g172) & (!g349) & (!g421)) + ((!g134) & (sk[56]) & (!g109) & (!g172) & (!g349) & (g421)) + ((!g134) & (sk[56]) & (!g109) & (!g172) & (g349) & (!g421)) + ((!g134) & (sk[56]) & (!g109) & (!g172) & (g349) & (g421)) + ((!g134) & (sk[56]) & (!g109) & (g172) & (!g349) & (!g421)) + ((!g134) & (sk[56]) & (!g109) & (g172) & (!g349) & (g421)) + ((!g134) & (sk[56]) & (!g109) & (g172) & (g349) & (!g421)) + ((!g134) & (sk[56]) & (!g109) & (g172) & (g349) & (g421)) + ((!g134) & (sk[56]) & (g109) & (!g172) & (!g349) & (!g421)) + ((!g134) & (sk[56]) & (g109) & (!g172) & (!g349) & (g421)) + ((!g134) & (sk[56]) & (g109) & (g172) & (!g349) & (!g421)) + ((!g134) & (sk[56]) & (g109) & (g172) & (!g349) & (g421)) + ((g134) & (!sk[56]) & (!g109) & (!g172) & (!g349) & (!g421)) + ((g134) & (!sk[56]) & (!g109) & (!g172) & (!g349) & (g421)) + ((g134) & (!sk[56]) & (!g109) & (!g172) & (g349) & (!g421)) + ((g134) & (!sk[56]) & (!g109) & (!g172) & (g349) & (g421)) + ((g134) & (!sk[56]) & (!g109) & (g172) & (!g349) & (!g421)) + ((g134) & (!sk[56]) & (!g109) & (g172) & (!g349) & (g421)) + ((g134) & (!sk[56]) & (!g109) & (g172) & (g349) & (!g421)) + ((g134) & (!sk[56]) & (!g109) & (g172) & (g349) & (g421)) + ((g134) & (!sk[56]) & (g109) & (!g172) & (!g349) & (!g421)) + ((g134) & (!sk[56]) & (g109) & (!g172) & (!g349) & (g421)) + ((g134) & (!sk[56]) & (g109) & (!g172) & (g349) & (!g421)) + ((g134) & (!sk[56]) & (g109) & (!g172) & (g349) & (g421)) + ((g134) & (!sk[56]) & (g109) & (g172) & (!g349) & (!g421)) + ((g134) & (!sk[56]) & (g109) & (g172) & (!g349) & (g421)) + ((g134) & (!sk[56]) & (g109) & (g172) & (g349) & (!g421)) + ((g134) & (!sk[56]) & (g109) & (g172) & (g349) & (g421)) + ((g134) & (sk[56]) & (!g109) & (!g172) & (!g349) & (g421)) + ((g134) & (sk[56]) & (!g109) & (!g172) & (g349) & (g421)) + ((g134) & (sk[56]) & (g109) & (!g172) & (!g349) & (g421)));
	assign g423 = (((!sk[57]) & (g31) & (!g87)) + ((!sk[57]) & (g31) & (g87)) + ((sk[57]) & (g31) & (g87)));
	assign g424 = (((i_15_) & (!g113) & (!sk[58]) & (!g182)) + ((i_15_) & (!g113) & (!sk[58]) & (g182)) + ((i_15_) & (g113) & (!sk[58]) & (!g182)) + ((i_15_) & (g113) & (!sk[58]) & (g182)) + ((i_15_) & (g113) & (sk[58]) & (g182)));
	assign g425 = (((g423) & (!sk[59]) & (!g424)) + ((g423) & (!sk[59]) & (g424)) + ((g423) & (sk[59]) & (g424)));
	assign g426 = (((!g204) & (!g279) & (sk[60]) & (!g285)) + ((!g204) & (g279) & (sk[60]) & (!g285)) + ((g204) & (!g279) & (!sk[60]) & (!g285)) + ((g204) & (!g279) & (!sk[60]) & (g285)) + ((g204) & (g279) & (!sk[60]) & (!g285)) + ((g204) & (g279) & (!sk[60]) & (g285)) + ((g204) & (g279) & (sk[60]) & (!g285)));
	assign g427 = (((!sk[61]) & (g203) & (!g214)) + ((!sk[61]) & (g203) & (g214)) + ((sk[61]) & (g203) & (g214)));
	assign g428 = (((!i_5_) & (!i_3_) & (i_4_) & (!sk[62]) & (g57)) + ((!i_5_) & (!i_3_) & (i_4_) & (sk[62]) & (g57)) + ((!i_5_) & (i_3_) & (!i_4_) & (!sk[62]) & (!g57)) + ((!i_5_) & (i_3_) & (!i_4_) & (!sk[62]) & (g57)) + ((!i_5_) & (i_3_) & (i_4_) & (!sk[62]) & (!g57)) + ((!i_5_) & (i_3_) & (i_4_) & (!sk[62]) & (g57)) + ((i_5_) & (!i_3_) & (!i_4_) & (sk[62]) & (g57)) + ((i_5_) & (!i_3_) & (i_4_) & (!sk[62]) & (!g57)) + ((i_5_) & (!i_3_) & (i_4_) & (!sk[62]) & (g57)) + ((i_5_) & (i_3_) & (!i_4_) & (!sk[62]) & (!g57)) + ((i_5_) & (i_3_) & (!i_4_) & (!sk[62]) & (g57)) + ((i_5_) & (i_3_) & (i_4_) & (!sk[62]) & (!g57)) + ((i_5_) & (i_3_) & (i_4_) & (!sk[62]) & (g57)));
	assign g429 = (((!sk[63]) & (g31) & (!g428)) + ((!sk[63]) & (g31) & (g428)) + ((sk[63]) & (g31) & (g428)));
	assign g430 = (((g110) & (!g111) & (!sk[64]) & (!g177)) + ((g110) & (!g111) & (!sk[64]) & (g177)) + ((g110) & (g111) & (!sk[64]) & (!g177)) + ((g110) & (g111) & (!sk[64]) & (g177)) + ((g110) & (g111) & (sk[64]) & (g177)));
	assign g431 = (((g31) & (!sk[65]) & (!g110) & (!g199)) + ((g31) & (!sk[65]) & (!g110) & (g199)) + ((g31) & (!sk[65]) & (g110) & (!g199)) + ((g31) & (!sk[65]) & (g110) & (g199)) + ((g31) & (sk[65]) & (g110) & (g199)));
	assign g432 = (((!g59) & (!g99) & (!g172) & (!g339) & (!g430) & (!g431)) + ((!g59) & (!g99) & (!g172) & (g339) & (!g430) & (!g431)) + ((!g59) & (!g99) & (g172) & (!g339) & (!g430) & (!g431)) + ((!g59) & (!g99) & (g172) & (g339) & (!g430) & (!g431)) + ((!g59) & (g99) & (!g172) & (!g339) & (!g430) & (!g431)) + ((g59) & (!g99) & (!g172) & (!g339) & (!g430) & (!g431)) + ((g59) & (g99) & (!g172) & (!g339) & (!g430) & (!g431)));
	assign g433 = (((!g277) & (!g232) & (!g339) & (!g427) & (!g429) & (g432)) + ((!g277) & (!g232) & (!g339) & (!g427) & (g429) & (g432)) + ((!g277) & (!g232) & (g339) & (!g427) & (!g429) & (g432)) + ((g277) & (!g232) & (!g339) & (!g427) & (!g429) & (g432)) + ((g277) & (!g232) & (!g339) & (!g427) & (g429) & (g432)) + ((g277) & (!g232) & (g339) & (!g427) & (!g429) & (g432)) + ((g277) & (g232) & (!g339) & (!g427) & (!g429) & (g432)) + ((g277) & (g232) & (!g339) & (!g427) & (g429) & (g432)) + ((g277) & (g232) & (g339) & (!g427) & (!g429) & (g432)));
	assign g434 = (((!sk[68]) & (g134) & (!g118) & (!g231)) + ((!sk[68]) & (g134) & (!g118) & (g231)) + ((!sk[68]) & (g134) & (g118) & (!g231)) + ((!sk[68]) & (g134) & (g118) & (g231)) + ((sk[68]) & (!g134) & (g118) & (!g231)) + ((sk[68]) & (g134) & (!g118) & (!g231)) + ((sk[68]) & (g134) & (g118) & (!g231)));
	assign g435 = (((!sk[69]) & (g118) & (!g224) & (!g197)) + ((!sk[69]) & (g118) & (!g224) & (g197)) + ((!sk[69]) & (g118) & (g224) & (!g197)) + ((!sk[69]) & (g118) & (g224) & (g197)) + ((sk[69]) & (g118) & (!g224) & (g197)) + ((sk[69]) & (g118) & (g224) & (!g197)) + ((sk[69]) & (g118) & (g224) & (g197)));
	assign g436 = (((!i_8_) & (!g134) & (!g135) & (!g177) & (!sk[70]) & (g173)) + ((!i_8_) & (!g134) & (!g135) & (g177) & (!sk[70]) & (g173)) + ((!i_8_) & (!g134) & (g135) & (!g177) & (!sk[70]) & (g173)) + ((!i_8_) & (!g134) & (g135) & (g177) & (!sk[70]) & (g173)) + ((!i_8_) & (g134) & (!g135) & (!g177) & (!sk[70]) & (g173)) + ((!i_8_) & (g134) & (!g135) & (!g177) & (sk[70]) & (g173)) + ((!i_8_) & (g134) & (!g135) & (g177) & (!sk[70]) & (g173)) + ((!i_8_) & (g134) & (!g135) & (g177) & (sk[70]) & (g173)) + ((!i_8_) & (g134) & (g135) & (!g177) & (!sk[70]) & (g173)) + ((!i_8_) & (g134) & (g135) & (!g177) & (sk[70]) & (g173)) + ((!i_8_) & (g134) & (g135) & (g177) & (!sk[70]) & (g173)) + ((!i_8_) & (g134) & (g135) & (g177) & (sk[70]) & (g173)) + ((i_8_) & (!g134) & (!g135) & (!g177) & (!sk[70]) & (!g173)) + ((i_8_) & (!g134) & (!g135) & (!g177) & (!sk[70]) & (g173)) + ((i_8_) & (!g134) & (!g135) & (g177) & (!sk[70]) & (!g173)) + ((i_8_) & (!g134) & (!g135) & (g177) & (!sk[70]) & (g173)) + ((i_8_) & (!g134) & (g135) & (!g177) & (!sk[70]) & (!g173)) + ((i_8_) & (!g134) & (g135) & (!g177) & (!sk[70]) & (g173)) + ((i_8_) & (!g134) & (g135) & (!g177) & (sk[70]) & (g173)) + ((i_8_) & (!g134) & (g135) & (g177) & (!sk[70]) & (!g173)) + ((i_8_) & (!g134) & (g135) & (g177) & (!sk[70]) & (g173)) + ((i_8_) & (!g134) & (g135) & (g177) & (sk[70]) & (!g173)) + ((i_8_) & (!g134) & (g135) & (g177) & (sk[70]) & (g173)) + ((i_8_) & (g134) & (!g135) & (!g177) & (!sk[70]) & (!g173)) + ((i_8_) & (g134) & (!g135) & (!g177) & (!sk[70]) & (g173)) + ((i_8_) & (g134) & (!g135) & (!g177) & (sk[70]) & (g173)) + ((i_8_) & (g134) & (!g135) & (g177) & (!sk[70]) & (!g173)) + ((i_8_) & (g134) & (!g135) & (g177) & (!sk[70]) & (g173)) + ((i_8_) & (g134) & (!g135) & (g177) & (sk[70]) & (g173)) + ((i_8_) & (g134) & (g135) & (!g177) & (!sk[70]) & (!g173)) + ((i_8_) & (g134) & (g135) & (!g177) & (!sk[70]) & (g173)) + ((i_8_) & (g134) & (g135) & (!g177) & (sk[70]) & (g173)) + ((i_8_) & (g134) & (g135) & (g177) & (!sk[70]) & (!g173)) + ((i_8_) & (g134) & (g135) & (g177) & (!sk[70]) & (g173)) + ((i_8_) & (g134) & (g135) & (g177) & (sk[70]) & (!g173)) + ((i_8_) & (g134) & (g135) & (g177) & (sk[70]) & (g173)));
	assign g437 = (((!i_8_) & (!sk[71]) & (!g100) & (g177) & (g172)) + ((!i_8_) & (!sk[71]) & (g100) & (!g177) & (!g172)) + ((!i_8_) & (!sk[71]) & (g100) & (!g177) & (g172)) + ((!i_8_) & (!sk[71]) & (g100) & (g177) & (!g172)) + ((!i_8_) & (!sk[71]) & (g100) & (g177) & (g172)) + ((i_8_) & (!sk[71]) & (!g100) & (g177) & (!g172)) + ((i_8_) & (!sk[71]) & (!g100) & (g177) & (g172)) + ((i_8_) & (!sk[71]) & (g100) & (!g177) & (!g172)) + ((i_8_) & (!sk[71]) & (g100) & (!g177) & (g172)) + ((i_8_) & (!sk[71]) & (g100) & (g177) & (!g172)) + ((i_8_) & (!sk[71]) & (g100) & (g177) & (g172)) + ((i_8_) & (sk[71]) & (g100) & (!g177) & (g172)) + ((i_8_) & (sk[71]) & (g100) & (g177) & (!g172)) + ((i_8_) & (sk[71]) & (g100) & (g177) & (g172)));
	assign g438 = (((!i_8_) & (!g108) & (!g226) & (!sk[72]) & (!g224) & (g231)) + ((!i_8_) & (!g108) & (!g226) & (!sk[72]) & (g224) & (g231)) + ((!i_8_) & (!g108) & (g226) & (!sk[72]) & (!g224) & (g231)) + ((!i_8_) & (!g108) & (g226) & (!sk[72]) & (g224) & (g231)) + ((!i_8_) & (g108) & (!g226) & (!sk[72]) & (!g224) & (g231)) + ((!i_8_) & (g108) & (!g226) & (!sk[72]) & (g224) & (g231)) + ((!i_8_) & (g108) & (!g226) & (sk[72]) & (!g224) & (!g231)) + ((!i_8_) & (g108) & (!g226) & (sk[72]) & (!g224) & (g231)) + ((!i_8_) & (g108) & (!g226) & (sk[72]) & (g224) & (!g231)) + ((!i_8_) & (g108) & (!g226) & (sk[72]) & (g224) & (g231)) + ((!i_8_) & (g108) & (g226) & (!sk[72]) & (!g224) & (g231)) + ((!i_8_) & (g108) & (g226) & (!sk[72]) & (g224) & (g231)) + ((!i_8_) & (g108) & (g226) & (sk[72]) & (!g224) & (!g231)) + ((!i_8_) & (g108) & (g226) & (sk[72]) & (g224) & (!g231)) + ((!i_8_) & (g108) & (g226) & (sk[72]) & (g224) & (g231)) + ((i_8_) & (!g108) & (!g226) & (!sk[72]) & (!g224) & (!g231)) + ((i_8_) & (!g108) & (!g226) & (!sk[72]) & (!g224) & (g231)) + ((i_8_) & (!g108) & (!g226) & (!sk[72]) & (g224) & (!g231)) + ((i_8_) & (!g108) & (!g226) & (!sk[72]) & (g224) & (g231)) + ((i_8_) & (!g108) & (g226) & (!sk[72]) & (!g224) & (!g231)) + ((i_8_) & (!g108) & (g226) & (!sk[72]) & (!g224) & (g231)) + ((i_8_) & (!g108) & (g226) & (!sk[72]) & (g224) & (!g231)) + ((i_8_) & (!g108) & (g226) & (!sk[72]) & (g224) & (g231)) + ((i_8_) & (g108) & (!g226) & (!sk[72]) & (!g224) & (!g231)) + ((i_8_) & (g108) & (!g226) & (!sk[72]) & (!g224) & (g231)) + ((i_8_) & (g108) & (!g226) & (!sk[72]) & (g224) & (!g231)) + ((i_8_) & (g108) & (!g226) & (!sk[72]) & (g224) & (g231)) + ((i_8_) & (g108) & (g226) & (!sk[72]) & (!g224) & (!g231)) + ((i_8_) & (g108) & (g226) & (!sk[72]) & (!g224) & (g231)) + ((i_8_) & (g108) & (g226) & (!sk[72]) & (g224) & (!g231)) + ((i_8_) & (g108) & (g226) & (!sk[72]) & (g224) & (g231)));
	assign g439 = (((!g434) & (!g435) & (!sk[73]) & (!g436) & (!g437) & (g438)) + ((!g434) & (!g435) & (!sk[73]) & (!g436) & (g437) & (g438)) + ((!g434) & (!g435) & (!sk[73]) & (g436) & (!g437) & (g438)) + ((!g434) & (!g435) & (!sk[73]) & (g436) & (g437) & (g438)) + ((!g434) & (!g435) & (sk[73]) & (!g436) & (!g437) & (!g438)) + ((!g434) & (g435) & (!sk[73]) & (!g436) & (!g437) & (g438)) + ((!g434) & (g435) & (!sk[73]) & (!g436) & (g437) & (g438)) + ((!g434) & (g435) & (!sk[73]) & (g436) & (!g437) & (g438)) + ((!g434) & (g435) & (!sk[73]) & (g436) & (g437) & (g438)) + ((g434) & (!g435) & (!sk[73]) & (!g436) & (!g437) & (!g438)) + ((g434) & (!g435) & (!sk[73]) & (!g436) & (!g437) & (g438)) + ((g434) & (!g435) & (!sk[73]) & (!g436) & (g437) & (!g438)) + ((g434) & (!g435) & (!sk[73]) & (!g436) & (g437) & (g438)) + ((g434) & (!g435) & (!sk[73]) & (g436) & (!g437) & (!g438)) + ((g434) & (!g435) & (!sk[73]) & (g436) & (!g437) & (g438)) + ((g434) & (!g435) & (!sk[73]) & (g436) & (g437) & (!g438)) + ((g434) & (!g435) & (!sk[73]) & (g436) & (g437) & (g438)) + ((g434) & (g435) & (!sk[73]) & (!g436) & (!g437) & (!g438)) + ((g434) & (g435) & (!sk[73]) & (!g436) & (!g437) & (g438)) + ((g434) & (g435) & (!sk[73]) & (!g436) & (g437) & (!g438)) + ((g434) & (g435) & (!sk[73]) & (!g436) & (g437) & (g438)) + ((g434) & (g435) & (!sk[73]) & (g436) & (!g437) & (!g438)) + ((g434) & (g435) & (!sk[73]) & (g436) & (!g437) & (g438)) + ((g434) & (g435) & (!sk[73]) & (g436) & (g437) & (!g438)) + ((g434) & (g435) & (!sk[73]) & (g436) & (g437) & (g438)));
	assign g440 = (((!i_8_) & (g4) & (g98) & (!g195) & (!g197) & (g173)) + ((!i_8_) & (g4) & (g98) & (!g195) & (g197) & (g173)) + ((!i_8_) & (g4) & (g98) & (g195) & (!g197) & (!g173)) + ((!i_8_) & (g4) & (g98) & (g195) & (!g197) & (g173)) + ((!i_8_) & (g4) & (g98) & (g195) & (g197) & (!g173)) + ((!i_8_) & (g4) & (g98) & (g195) & (g197) & (g173)) + ((i_8_) & (g4) & (g98) & (!g195) & (g197) & (!g173)) + ((i_8_) & (g4) & (g98) & (!g195) & (g197) & (g173)) + ((i_8_) & (g4) & (g98) & (g195) & (!g197) & (!g173)) + ((i_8_) & (g4) & (g98) & (g195) & (!g197) & (g173)) + ((i_8_) & (g4) & (g98) & (g195) & (g197) & (!g173)) + ((i_8_) & (g4) & (g98) & (g195) & (g197) & (g173)));
	assign g441 = (((!g109) & (!g146) & (!g195) & (!g232) & (!g173) & (!g440)) + ((!g109) & (!g146) & (!g195) & (!g232) & (g173) & (!g440)) + ((!g109) & (!g146) & (!g195) & (g232) & (!g173) & (!g440)) + ((!g109) & (!g146) & (!g195) & (g232) & (g173) & (!g440)) + ((!g109) & (g146) & (!g195) & (!g232) & (!g173) & (!g440)) + ((!g109) & (g146) & (!g195) & (!g232) & (g173) & (!g440)) + ((!g109) & (g146) & (!g195) & (g232) & (!g173) & (!g440)) + ((!g109) & (g146) & (!g195) & (g232) & (g173) & (!g440)) + ((!g109) & (g146) & (g195) & (!g232) & (!g173) & (!g440)) + ((!g109) & (g146) & (g195) & (!g232) & (g173) & (!g440)) + ((!g109) & (g146) & (g195) & (g232) & (!g173) & (!g440)) + ((!g109) & (g146) & (g195) & (g232) & (g173) & (!g440)) + ((g109) & (!g146) & (!g195) & (!g232) & (!g173) & (!g440)) + ((g109) & (g146) & (!g195) & (!g232) & (!g173) & (!g440)) + ((g109) & (g146) & (g195) & (!g232) & (!g173) & (!g440)));
	assign g442 = (((!i_8_) & (!g88) & (g224) & (!sk[76]) & (g197)) + ((!i_8_) & (g88) & (!g224) & (!sk[76]) & (!g197)) + ((!i_8_) & (g88) & (!g224) & (!sk[76]) & (g197)) + ((!i_8_) & (g88) & (!g224) & (sk[76]) & (g197)) + ((!i_8_) & (g88) & (g224) & (!sk[76]) & (!g197)) + ((!i_8_) & (g88) & (g224) & (!sk[76]) & (g197)) + ((!i_8_) & (g88) & (g224) & (sk[76]) & (!g197)) + ((!i_8_) & (g88) & (g224) & (sk[76]) & (g197)) + ((i_8_) & (!g88) & (g224) & (!sk[76]) & (!g197)) + ((i_8_) & (!g88) & (g224) & (!sk[76]) & (g197)) + ((i_8_) & (g88) & (!g224) & (!sk[76]) & (!g197)) + ((i_8_) & (g88) & (!g224) & (!sk[76]) & (g197)) + ((i_8_) & (g88) & (g224) & (!sk[76]) & (!g197)) + ((i_8_) & (g88) & (g224) & (!sk[76]) & (g197)));
	assign g443 = (((!g109) & (!g203) & (!g268) & (!g172) & (!g339) & (!g442)) + ((!g109) & (!g203) & (!g268) & (!g172) & (g339) & (!g442)) + ((!g109) & (!g203) & (!g268) & (g172) & (!g339) & (!g442)) + ((!g109) & (!g203) & (!g268) & (g172) & (g339) & (!g442)) + ((!g109) & (!g203) & (g268) & (!g172) & (!g339) & (!g442)) + ((!g109) & (!g203) & (g268) & (!g172) & (g339) & (!g442)) + ((!g109) & (!g203) & (g268) & (g172) & (!g339) & (!g442)) + ((!g109) & (!g203) & (g268) & (g172) & (g339) & (!g442)) + ((!g109) & (g203) & (!g268) & (!g172) & (!g339) & (!g442)) + ((!g109) & (g203) & (!g268) & (!g172) & (g339) & (!g442)) + ((!g109) & (g203) & (!g268) & (g172) & (!g339) & (!g442)) + ((!g109) & (g203) & (!g268) & (g172) & (g339) & (!g442)) + ((!g109) & (g203) & (g268) & (!g172) & (!g339) & (!g442)) + ((!g109) & (g203) & (g268) & (!g172) & (g339) & (!g442)) + ((!g109) & (g203) & (g268) & (g172) & (!g339) & (!g442)) + ((!g109) & (g203) & (g268) & (g172) & (g339) & (!g442)) + ((g109) & (!g203) & (!g268) & (!g172) & (!g339) & (!g442)));
	assign g444 = (((!i_8_) & (!sk[78]) & (!g88) & (g323) & (g231)) + ((!i_8_) & (!sk[78]) & (g88) & (!g323) & (!g231)) + ((!i_8_) & (!sk[78]) & (g88) & (!g323) & (g231)) + ((!i_8_) & (!sk[78]) & (g88) & (g323) & (!g231)) + ((!i_8_) & (!sk[78]) & (g88) & (g323) & (g231)) + ((!i_8_) & (sk[78]) & (!g88) & (g323) & (!g231)) + ((!i_8_) & (sk[78]) & (g88) & (!g323) & (!g231)) + ((!i_8_) & (sk[78]) & (g88) & (g323) & (!g231)) + ((i_8_) & (!sk[78]) & (!g88) & (g323) & (!g231)) + ((i_8_) & (!sk[78]) & (!g88) & (g323) & (g231)) + ((i_8_) & (!sk[78]) & (g88) & (!g323) & (!g231)) + ((i_8_) & (!sk[78]) & (g88) & (!g323) & (g231)) + ((i_8_) & (!sk[78]) & (g88) & (g323) & (!g231)) + ((i_8_) & (!sk[78]) & (g88) & (g323) & (g231)) + ((i_8_) & (sk[78]) & (!g88) & (g323) & (!g231)) + ((i_8_) & (sk[78]) & (g88) & (g323) & (!g231)));
	assign g445 = (((!i_8_) & (!g88) & (g232) & (!sk[79]) & (g339)) + ((!i_8_) & (g88) & (!g232) & (!sk[79]) & (!g339)) + ((!i_8_) & (g88) & (!g232) & (!sk[79]) & (g339)) + ((!i_8_) & (g88) & (!g232) & (sk[79]) & (g339)) + ((!i_8_) & (g88) & (g232) & (!sk[79]) & (!g339)) + ((!i_8_) & (g88) & (g232) & (!sk[79]) & (g339)) + ((!i_8_) & (g88) & (g232) & (sk[79]) & (!g339)) + ((!i_8_) & (g88) & (g232) & (sk[79]) & (g339)) + ((i_8_) & (!g88) & (g232) & (!sk[79]) & (!g339)) + ((i_8_) & (!g88) & (g232) & (!sk[79]) & (g339)) + ((i_8_) & (g88) & (!g232) & (!sk[79]) & (!g339)) + ((i_8_) & (g88) & (!g232) & (!sk[79]) & (g339)) + ((i_8_) & (g88) & (g232) & (!sk[79]) & (!g339)) + ((i_8_) & (g88) & (g232) & (!sk[79]) & (g339)));
	assign g446 = (((!i_8_) & (!g88) & (!sk[80]) & (g226) & (g349)) + ((!i_8_) & (g88) & (!sk[80]) & (!g226) & (!g349)) + ((!i_8_) & (g88) & (!sk[80]) & (!g226) & (g349)) + ((!i_8_) & (g88) & (!sk[80]) & (g226) & (!g349)) + ((!i_8_) & (g88) & (!sk[80]) & (g226) & (g349)) + ((!i_8_) & (g88) & (sk[80]) & (!g226) & (!g349)) + ((!i_8_) & (g88) & (sk[80]) & (!g226) & (g349)) + ((!i_8_) & (g88) & (sk[80]) & (g226) & (g349)) + ((i_8_) & (!g88) & (!sk[80]) & (g226) & (!g349)) + ((i_8_) & (!g88) & (!sk[80]) & (g226) & (g349)) + ((i_8_) & (g88) & (!sk[80]) & (!g226) & (!g349)) + ((i_8_) & (g88) & (!sk[80]) & (!g226) & (g349)) + ((i_8_) & (g88) & (!sk[80]) & (g226) & (!g349)) + ((i_8_) & (g88) & (!sk[80]) & (g226) & (g349)));
	assign g447 = (((!sk[81]) & (g134) & (!g226) & (!g349)) + ((!sk[81]) & (g134) & (!g226) & (g349)) + ((!sk[81]) & (g134) & (g226) & (!g349)) + ((!sk[81]) & (g134) & (g226) & (g349)) + ((sk[81]) & (g134) & (!g226) & (!g349)) + ((sk[81]) & (g134) & (!g226) & (g349)) + ((sk[81]) & (g134) & (g226) & (g349)));
	assign g448 = (((!sk[82]) & (!g224) & (!g232) & (g349) & (g423)) + ((!sk[82]) & (!g224) & (g232) & (!g349) & (!g423)) + ((!sk[82]) & (!g224) & (g232) & (!g349) & (g423)) + ((!sk[82]) & (!g224) & (g232) & (g349) & (!g423)) + ((!sk[82]) & (!g224) & (g232) & (g349) & (g423)) + ((!sk[82]) & (g224) & (!g232) & (g349) & (!g423)) + ((!sk[82]) & (g224) & (!g232) & (g349) & (g423)) + ((!sk[82]) & (g224) & (g232) & (!g349) & (!g423)) + ((!sk[82]) & (g224) & (g232) & (!g349) & (g423)) + ((!sk[82]) & (g224) & (g232) & (g349) & (!g423)) + ((!sk[82]) & (g224) & (g232) & (g349) & (g423)) + ((sk[82]) & (!g224) & (!g232) & (g349) & (g423)) + ((sk[82]) & (!g224) & (g232) & (!g349) & (g423)) + ((sk[82]) & (!g224) & (g232) & (g349) & (g423)) + ((sk[82]) & (g224) & (!g232) & (!g349) & (g423)) + ((sk[82]) & (g224) & (!g232) & (g349) & (g423)) + ((sk[82]) & (g224) & (g232) & (!g349) & (g423)) + ((sk[82]) & (g224) & (g232) & (g349) & (g423)));
	assign g449 = (((!g118) & (!g226) & (g203) & (!sk[83]) & (g349)) + ((!g118) & (g226) & (!g203) & (!sk[83]) & (!g349)) + ((!g118) & (g226) & (!g203) & (!sk[83]) & (g349)) + ((!g118) & (g226) & (g203) & (!sk[83]) & (!g349)) + ((!g118) & (g226) & (g203) & (!sk[83]) & (g349)) + ((g118) & (!g226) & (!g203) & (sk[83]) & (!g349)) + ((g118) & (!g226) & (!g203) & (sk[83]) & (g349)) + ((g118) & (!g226) & (g203) & (!sk[83]) & (!g349)) + ((g118) & (!g226) & (g203) & (!sk[83]) & (g349)) + ((g118) & (!g226) & (g203) & (sk[83]) & (!g349)) + ((g118) & (!g226) & (g203) & (sk[83]) & (g349)) + ((g118) & (g226) & (!g203) & (!sk[83]) & (!g349)) + ((g118) & (g226) & (!g203) & (!sk[83]) & (g349)) + ((g118) & (g226) & (!g203) & (sk[83]) & (g349)) + ((g118) & (g226) & (g203) & (!sk[83]) & (!g349)) + ((g118) & (g226) & (g203) & (!sk[83]) & (g349)) + ((g118) & (g226) & (g203) & (sk[83]) & (!g349)) + ((g118) & (g226) & (g203) & (sk[83]) & (g349)));
	assign g450 = (((!g444) & (!g445) & (!g446) & (!g447) & (!g448) & (!g449)));
	assign g451 = (((g99) & (!g226) & (!sk[85]) & (!g177)) + ((g99) & (!g226) & (!sk[85]) & (g177)) + ((g99) & (!g226) & (sk[85]) & (!g177)) + ((g99) & (!g226) & (sk[85]) & (g177)) + ((g99) & (g226) & (!sk[85]) & (!g177)) + ((g99) & (g226) & (!sk[85]) & (g177)) + ((g99) & (g226) & (sk[85]) & (g177)));
	assign g452 = (((!sk[86]) & (g149) & (!g226) & (!g177)) + ((!sk[86]) & (g149) & (!g226) & (g177)) + ((!sk[86]) & (g149) & (g226) & (!g177)) + ((!sk[86]) & (g149) & (g226) & (g177)) + ((sk[86]) & (!g149) & (!g226) & (!g177)) + ((sk[86]) & (!g149) & (!g226) & (g177)) + ((sk[86]) & (!g149) & (g226) & (!g177)) + ((sk[86]) & (!g149) & (g226) & (g177)) + ((sk[86]) & (g149) & (g226) & (!g177)));
	assign g453 = (((g59) & (!sk[87]) & (!g203) & (!g224)) + ((g59) & (!sk[87]) & (!g203) & (g224)) + ((g59) & (!sk[87]) & (g203) & (!g224)) + ((g59) & (!sk[87]) & (g203) & (g224)) + ((g59) & (sk[87]) & (!g203) & (g224)) + ((g59) & (sk[87]) & (g203) & (!g224)) + ((g59) & (sk[87]) & (g203) & (g224)));
	assign g454 = (((g149) & (!g199) & (!sk[88]) & (!g349)) + ((g149) & (!g199) & (!sk[88]) & (g349)) + ((g149) & (!g199) & (sk[88]) & (g349)) + ((g149) & (g199) & (!sk[88]) & (!g349)) + ((g149) & (g199) & (!sk[88]) & (g349)) + ((g149) & (g199) & (sk[88]) & (!g349)) + ((g149) & (g199) & (sk[88]) & (g349)));
	assign g455 = (((!g99) & (!sk[89]) & (!g199) & (!g197) & (!g268) & (g349)) + ((!g99) & (!sk[89]) & (!g199) & (!g197) & (g268) & (g349)) + ((!g99) & (!sk[89]) & (!g199) & (g197) & (!g268) & (g349)) + ((!g99) & (!sk[89]) & (!g199) & (g197) & (g268) & (g349)) + ((!g99) & (!sk[89]) & (g199) & (!g197) & (!g268) & (g349)) + ((!g99) & (!sk[89]) & (g199) & (!g197) & (g268) & (g349)) + ((!g99) & (!sk[89]) & (g199) & (g197) & (!g268) & (g349)) + ((!g99) & (!sk[89]) & (g199) & (g197) & (g268) & (g349)) + ((g99) & (!sk[89]) & (!g199) & (!g197) & (!g268) & (!g349)) + ((g99) & (!sk[89]) & (!g199) & (!g197) & (!g268) & (g349)) + ((g99) & (!sk[89]) & (!g199) & (!g197) & (g268) & (!g349)) + ((g99) & (!sk[89]) & (!g199) & (!g197) & (g268) & (g349)) + ((g99) & (!sk[89]) & (!g199) & (g197) & (!g268) & (!g349)) + ((g99) & (!sk[89]) & (!g199) & (g197) & (!g268) & (g349)) + ((g99) & (!sk[89]) & (!g199) & (g197) & (g268) & (!g349)) + ((g99) & (!sk[89]) & (!g199) & (g197) & (g268) & (g349)) + ((g99) & (!sk[89]) & (g199) & (!g197) & (!g268) & (!g349)) + ((g99) & (!sk[89]) & (g199) & (!g197) & (!g268) & (g349)) + ((g99) & (!sk[89]) & (g199) & (!g197) & (g268) & (!g349)) + ((g99) & (!sk[89]) & (g199) & (!g197) & (g268) & (g349)) + ((g99) & (!sk[89]) & (g199) & (g197) & (!g268) & (!g349)) + ((g99) & (!sk[89]) & (g199) & (g197) & (!g268) & (g349)) + ((g99) & (!sk[89]) & (g199) & (g197) & (g268) & (!g349)) + ((g99) & (!sk[89]) & (g199) & (g197) & (g268) & (g349)) + ((g99) & (sk[89]) & (!g199) & (!g197) & (!g268) & (g349)) + ((g99) & (sk[89]) & (!g199) & (!g197) & (g268) & (!g349)) + ((g99) & (sk[89]) & (!g199) & (!g197) & (g268) & (g349)) + ((g99) & (sk[89]) & (!g199) & (g197) & (!g268) & (!g349)) + ((g99) & (sk[89]) & (!g199) & (g197) & (!g268) & (g349)) + ((g99) & (sk[89]) & (!g199) & (g197) & (g268) & (!g349)) + ((g99) & (sk[89]) & (!g199) & (g197) & (g268) & (g349)) + ((g99) & (sk[89]) & (g199) & (!g197) & (!g268) & (!g349)) + ((g99) & (sk[89]) & (g199) & (!g197) & (!g268) & (g349)) + ((g99) & (sk[89]) & (g199) & (!g197) & (g268) & (!g349)) + ((g99) & (sk[89]) & (g199) & (!g197) & (g268) & (g349)) + ((g99) & (sk[89]) & (g199) & (g197) & (!g268) & (!g349)) + ((g99) & (sk[89]) & (g199) & (g197) & (!g268) & (g349)) + ((g99) & (sk[89]) & (g199) & (g197) & (g268) & (!g349)) + ((g99) & (sk[89]) & (g199) & (g197) & (g268) & (g349)));
	assign g456 = (((!g451) & (!g452) & (!g453) & (!sk[90]) & (!g454) & (g455)) + ((!g451) & (!g452) & (!g453) & (!sk[90]) & (g454) & (g455)) + ((!g451) & (!g452) & (g453) & (!sk[90]) & (!g454) & (g455)) + ((!g451) & (!g452) & (g453) & (!sk[90]) & (g454) & (g455)) + ((!g451) & (g452) & (!g453) & (!sk[90]) & (!g454) & (g455)) + ((!g451) & (g452) & (!g453) & (!sk[90]) & (g454) & (g455)) + ((!g451) & (g452) & (!g453) & (sk[90]) & (!g454) & (!g455)) + ((!g451) & (g452) & (g453) & (!sk[90]) & (!g454) & (g455)) + ((!g451) & (g452) & (g453) & (!sk[90]) & (g454) & (g455)) + ((g451) & (!g452) & (!g453) & (!sk[90]) & (!g454) & (!g455)) + ((g451) & (!g452) & (!g453) & (!sk[90]) & (!g454) & (g455)) + ((g451) & (!g452) & (!g453) & (!sk[90]) & (g454) & (!g455)) + ((g451) & (!g452) & (!g453) & (!sk[90]) & (g454) & (g455)) + ((g451) & (!g452) & (g453) & (!sk[90]) & (!g454) & (!g455)) + ((g451) & (!g452) & (g453) & (!sk[90]) & (!g454) & (g455)) + ((g451) & (!g452) & (g453) & (!sk[90]) & (g454) & (!g455)) + ((g451) & (!g452) & (g453) & (!sk[90]) & (g454) & (g455)) + ((g451) & (g452) & (!g453) & (!sk[90]) & (!g454) & (!g455)) + ((g451) & (g452) & (!g453) & (!sk[90]) & (!g454) & (g455)) + ((g451) & (g452) & (!g453) & (!sk[90]) & (g454) & (!g455)) + ((g451) & (g452) & (!g453) & (!sk[90]) & (g454) & (g455)) + ((g451) & (g452) & (g453) & (!sk[90]) & (!g454) & (!g455)) + ((g451) & (g452) & (g453) & (!sk[90]) & (!g454) & (g455)) + ((g451) & (g452) & (g453) & (!sk[90]) & (g454) & (!g455)) + ((g451) & (g452) & (g453) & (!sk[90]) & (g454) & (g455)));
	assign g457 = (((g433) & (g439) & (g441) & (g443) & (g450) & (g456)));
	assign g458 = (((!g136) & (!g195) & (g422) & (!g425) & (!g426) & (g457)) + ((!g136) & (g195) & (g422) & (!g425) & (!g426) & (g457)) + ((g136) & (!g195) & (g422) & (!g425) & (!g426) & (g457)));
	assign o_3_ = (((g73) & (!g169) & (!g275) & (!g336) & (!g420) & (!g458)) + ((g73) & (!g169) & (!g275) & (!g336) & (!g420) & (g458)) + ((g73) & (!g169) & (!g275) & (!g336) & (g420) & (!g458)) + ((g73) & (!g169) & (!g275) & (!g336) & (g420) & (g458)) + ((g73) & (!g169) & (!g275) & (g336) & (!g420) & (!g458)) + ((g73) & (!g169) & (!g275) & (g336) & (!g420) & (g458)) + ((g73) & (!g169) & (!g275) & (g336) & (g420) & (!g458)) + ((g73) & (!g169) & (!g275) & (g336) & (g420) & (g458)) + ((g73) & (!g169) & (g275) & (!g336) & (!g420) & (!g458)) + ((g73) & (!g169) & (g275) & (!g336) & (!g420) & (g458)) + ((g73) & (!g169) & (g275) & (!g336) & (g420) & (!g458)) + ((g73) & (!g169) & (g275) & (!g336) & (g420) & (g458)) + ((g73) & (!g169) & (g275) & (g336) & (!g420) & (!g458)) + ((g73) & (!g169) & (g275) & (g336) & (!g420) & (g458)) + ((g73) & (!g169) & (g275) & (g336) & (g420) & (!g458)) + ((g73) & (!g169) & (g275) & (g336) & (g420) & (g458)) + ((g73) & (g169) & (!g275) & (!g336) & (!g420) & (!g458)) + ((g73) & (g169) & (!g275) & (!g336) & (!g420) & (g458)) + ((g73) & (g169) & (!g275) & (!g336) & (g420) & (!g458)) + ((g73) & (g169) & (!g275) & (!g336) & (g420) & (g458)) + ((g73) & (g169) & (!g275) & (g336) & (!g420) & (!g458)) + ((g73) & (g169) & (!g275) & (g336) & (!g420) & (g458)) + ((g73) & (g169) & (!g275) & (g336) & (g420) & (!g458)) + ((g73) & (g169) & (!g275) & (g336) & (g420) & (g458)) + ((g73) & (g169) & (g275) & (!g336) & (!g420) & (!g458)) + ((g73) & (g169) & (g275) & (!g336) & (!g420) & (g458)) + ((g73) & (g169) & (g275) & (!g336) & (g420) & (!g458)) + ((g73) & (g169) & (g275) & (!g336) & (g420) & (g458)) + ((g73) & (g169) & (g275) & (g336) & (!g420) & (!g458)) + ((g73) & (g169) & (g275) & (g336) & (!g420) & (g458)) + ((g73) & (g169) & (g275) & (g336) & (g420) & (!g458)));
	assign g460 = (((!sk[94]) & (g48) & (!g158)) + ((!sk[94]) & (g48) & (g158)) + ((sk[94]) & (!g48) & (g158)));
	assign g461 = (((!i_14_) & (sk[95]) & (i_12_) & (i_13_)) + ((i_14_) & (!sk[95]) & (!i_12_) & (!i_13_)) + ((i_14_) & (!sk[95]) & (!i_12_) & (i_13_)) + ((i_14_) & (!sk[95]) & (i_12_) & (!i_13_)) + ((i_14_) & (!sk[95]) & (i_12_) & (i_13_)));
	assign g462 = (((!g18) & (sk[96]) & (!g461)) + ((g18) & (!sk[96]) & (!g461)) + ((g18) & (!sk[96]) & (g461)) + ((g18) & (sk[96]) & (!g461)) + ((g18) & (sk[96]) & (g461)));
	assign g463 = (((g151) & (!sk[97]) & (!g460) & (!g462)) + ((g151) & (!sk[97]) & (!g460) & (g462)) + ((g151) & (!sk[97]) & (g460) & (!g462)) + ((g151) & (!sk[97]) & (g460) & (g462)) + ((g151) & (sk[97]) & (!g460) & (!g462)) + ((g151) & (sk[97]) & (g460) & (!g462)) + ((g151) & (sk[97]) & (g460) & (g462)));
	assign g464 = (((!i_11_) & (!i_15_) & (!g113) & (sk[98]) & (!g48)) + ((!i_11_) & (!i_15_) & (!g113) & (sk[98]) & (g48)) + ((!i_11_) & (!i_15_) & (g113) & (!sk[98]) & (g48)) + ((!i_11_) & (!i_15_) & (g113) & (sk[98]) & (!g48)) + ((!i_11_) & (!i_15_) & (g113) & (sk[98]) & (g48)) + ((!i_11_) & (i_15_) & (!g113) & (!sk[98]) & (!g48)) + ((!i_11_) & (i_15_) & (!g113) & (!sk[98]) & (g48)) + ((!i_11_) & (i_15_) & (!g113) & (sk[98]) & (!g48)) + ((!i_11_) & (i_15_) & (!g113) & (sk[98]) & (g48)) + ((!i_11_) & (i_15_) & (g113) & (!sk[98]) & (!g48)) + ((!i_11_) & (i_15_) & (g113) & (!sk[98]) & (g48)) + ((!i_11_) & (i_15_) & (g113) & (sk[98]) & (g48)) + ((i_11_) & (!i_15_) & (!g113) & (sk[98]) & (!g48)) + ((i_11_) & (!i_15_) & (!g113) & (sk[98]) & (g48)) + ((i_11_) & (!i_15_) & (g113) & (!sk[98]) & (!g48)) + ((i_11_) & (!i_15_) & (g113) & (!sk[98]) & (g48)) + ((i_11_) & (!i_15_) & (g113) & (sk[98]) & (!g48)) + ((i_11_) & (!i_15_) & (g113) & (sk[98]) & (g48)) + ((i_11_) & (i_15_) & (!g113) & (!sk[98]) & (!g48)) + ((i_11_) & (i_15_) & (!g113) & (!sk[98]) & (g48)) + ((i_11_) & (i_15_) & (!g113) & (sk[98]) & (!g48)) + ((i_11_) & (i_15_) & (!g113) & (sk[98]) & (g48)) + ((i_11_) & (i_15_) & (g113) & (!sk[98]) & (!g48)) + ((i_11_) & (i_15_) & (g113) & (!sk[98]) & (g48)) + ((i_11_) & (i_15_) & (g113) & (sk[98]) & (!g48)) + ((i_11_) & (i_15_) & (g113) & (sk[98]) & (g48)));
	assign g465 = (((!i_11_) & (!sk[99]) & (!i_15_) & (g141) & (g48)) + ((!i_11_) & (!sk[99]) & (i_15_) & (!g141) & (!g48)) + ((!i_11_) & (!sk[99]) & (i_15_) & (!g141) & (g48)) + ((!i_11_) & (!sk[99]) & (i_15_) & (g141) & (!g48)) + ((!i_11_) & (!sk[99]) & (i_15_) & (g141) & (g48)) + ((!i_11_) & (sk[99]) & (!i_15_) & (!g141) & (!g48)) + ((!i_11_) & (sk[99]) & (!i_15_) & (!g141) & (g48)) + ((!i_11_) & (sk[99]) & (!i_15_) & (g141) & (!g48)) + ((!i_11_) & (sk[99]) & (!i_15_) & (g141) & (g48)) + ((!i_11_) & (sk[99]) & (i_15_) & (!g141) & (!g48)) + ((!i_11_) & (sk[99]) & (i_15_) & (!g141) & (g48)) + ((!i_11_) & (sk[99]) & (i_15_) & (g141) & (g48)) + ((i_11_) & (!sk[99]) & (!i_15_) & (g141) & (!g48)) + ((i_11_) & (!sk[99]) & (!i_15_) & (g141) & (g48)) + ((i_11_) & (!sk[99]) & (i_15_) & (!g141) & (!g48)) + ((i_11_) & (!sk[99]) & (i_15_) & (!g141) & (g48)) + ((i_11_) & (!sk[99]) & (i_15_) & (g141) & (!g48)) + ((i_11_) & (!sk[99]) & (i_15_) & (g141) & (g48)) + ((i_11_) & (sk[99]) & (!i_15_) & (!g141) & (!g48)) + ((i_11_) & (sk[99]) & (!i_15_) & (!g141) & (g48)) + ((i_11_) & (sk[99]) & (!i_15_) & (g141) & (!g48)) + ((i_11_) & (sk[99]) & (!i_15_) & (g141) & (g48)) + ((i_11_) & (sk[99]) & (i_15_) & (!g141) & (!g48)) + ((i_11_) & (sk[99]) & (i_15_) & (!g141) & (g48)) + ((i_11_) & (sk[99]) & (i_15_) & (g141) & (!g48)) + ((i_11_) & (sk[99]) & (i_15_) & (g141) & (g48)));
	assign g466 = (((!sk[100]) & (g284) & (!g460)) + ((!sk[100]) & (g284) & (g460)) + ((sk[100]) & (g284) & (g460)));
	assign g467 = (((!g6) & (sk[101]) & (!i_15_) & (!g48)) + ((!g6) & (sk[101]) & (!i_15_) & (g48)) + ((!g6) & (sk[101]) & (i_15_) & (!g48)) + ((!g6) & (sk[101]) & (i_15_) & (g48)) + ((g6) & (!sk[101]) & (!i_15_) & (!g48)) + ((g6) & (!sk[101]) & (!i_15_) & (g48)) + ((g6) & (!sk[101]) & (i_15_) & (!g48)) + ((g6) & (!sk[101]) & (i_15_) & (g48)) + ((g6) & (sk[101]) & (!i_15_) & (!g48)) + ((g6) & (sk[101]) & (!i_15_) & (g48)) + ((g6) & (sk[101]) & (i_15_) & (g48)));
	assign g468 = (((!g6) & (sk[102]) & (!i_15_) & (!g461)) + ((!g6) & (sk[102]) & (!i_15_) & (g461)) + ((!g6) & (sk[102]) & (i_15_) & (!g461)) + ((!g6) & (sk[102]) & (i_15_) & (g461)) + ((g6) & (!sk[102]) & (!i_15_) & (!g461)) + ((g6) & (!sk[102]) & (!i_15_) & (g461)) + ((g6) & (!sk[102]) & (i_15_) & (!g461)) + ((g6) & (!sk[102]) & (i_15_) & (g461)) + ((g6) & (sk[102]) & (!i_15_) & (!g461)) + ((g6) & (sk[102]) & (!i_15_) & (g461)) + ((g6) & (sk[102]) & (i_15_) & (!g461)));
	assign g469 = (((!sk[103]) & (g112) & (!g467) & (!g468)) + ((!sk[103]) & (g112) & (!g467) & (g468)) + ((!sk[103]) & (g112) & (g467) & (!g468)) + ((!sk[103]) & (g112) & (g467) & (g468)) + ((sk[103]) & (g112) & (!g467) & (!g468)) + ((sk[103]) & (g112) & (!g467) & (g468)) + ((sk[103]) & (g112) & (g467) & (!g468)));
	assign g470 = (((g158) & (!sk[104]) & (!g461)) + ((g158) & (!sk[104]) & (g461)) + ((g158) & (sk[104]) & (g461)));
	assign g471 = (((!g87) & (!g110) & (g111) & (!sk[105]) & (g465)) + ((!g87) & (g110) & (!g111) & (!sk[105]) & (!g465)) + ((!g87) & (g110) & (!g111) & (!sk[105]) & (g465)) + ((!g87) & (g110) & (g111) & (!sk[105]) & (!g465)) + ((!g87) & (g110) & (g111) & (!sk[105]) & (g465)) + ((!g87) & (g110) & (g111) & (sk[105]) & (!g465)) + ((g87) & (!g110) & (g111) & (!sk[105]) & (!g465)) + ((g87) & (!g110) & (g111) & (!sk[105]) & (g465)) + ((g87) & (!g110) & (g111) & (sk[105]) & (!g465)) + ((g87) & (g110) & (!g111) & (!sk[105]) & (!g465)) + ((g87) & (g110) & (!g111) & (!sk[105]) & (g465)) + ((g87) & (g110) & (g111) & (!sk[105]) & (!g465)) + ((g87) & (g110) & (g111) & (!sk[105]) & (g465)) + ((g87) & (g110) & (g111) & (sk[105]) & (!g465)));
	assign g472 = (((!i_8_) & (!g135) & (!g323) & (!g467) & (!g470) & (!g471)) + ((!i_8_) & (!g135) & (!g323) & (!g467) & (g470) & (!g471)) + ((!i_8_) & (!g135) & (!g323) & (g467) & (!g470) & (!g471)) + ((!i_8_) & (!g135) & (!g323) & (g467) & (g470) & (!g471)) + ((!i_8_) & (!g135) & (g323) & (g467) & (!g470) & (!g471)) + ((!i_8_) & (!g135) & (g323) & (g467) & (g470) & (!g471)) + ((!i_8_) & (g135) & (!g323) & (!g467) & (!g470) & (!g471)) + ((!i_8_) & (g135) & (!g323) & (!g467) & (g470) & (!g471)) + ((!i_8_) & (g135) & (!g323) & (g467) & (!g470) & (!g471)) + ((!i_8_) & (g135) & (!g323) & (g467) & (g470) & (!g471)) + ((!i_8_) & (g135) & (g323) & (g467) & (!g470) & (!g471)) + ((!i_8_) & (g135) & (g323) & (g467) & (g470) & (!g471)) + ((i_8_) & (!g135) & (!g323) & (!g467) & (!g470) & (!g471)) + ((i_8_) & (!g135) & (!g323) & (!g467) & (g470) & (!g471)) + ((i_8_) & (!g135) & (!g323) & (g467) & (!g470) & (!g471)) + ((i_8_) & (!g135) & (!g323) & (g467) & (g470) & (!g471)) + ((i_8_) & (!g135) & (g323) & (g467) & (!g470) & (!g471)) + ((i_8_) & (!g135) & (g323) & (g467) & (g470) & (!g471)) + ((i_8_) & (g135) & (!g323) & (!g467) & (!g470) & (!g471)) + ((i_8_) & (g135) & (!g323) & (g467) & (!g470) & (!g471)) + ((i_8_) & (g135) & (g323) & (g467) & (!g470) & (!g471)));
	assign g473 = (((!g101) & (!g464) & (!g465) & (!g466) & (!g469) & (g472)) + ((!g101) & (!g464) & (g465) & (!g466) & (!g469) & (g472)) + ((!g101) & (g464) & (!g465) & (!g466) & (!g469) & (g472)) + ((!g101) & (g464) & (g465) & (!g466) & (!g469) & (g472)) + ((g101) & (g464) & (g465) & (!g466) & (!g469) & (g472)));
	assign g474 = (((!g48) & (sk[108]) & (!g93)) + ((g48) & (!sk[108]) & (!g93)) + ((g48) & (!sk[108]) & (g93)));
	assign g475 = (((!g93) & (sk[109]) & (!g461)) + ((g93) & (!sk[109]) & (!g461)) + ((g93) & (!sk[109]) & (g461)) + ((g93) & (sk[109]) & (!g461)) + ((g93) & (sk[109]) & (g461)));
	assign g476 = (((!g338) & (sk[110]) & (!g474) & (!g475)) + ((!g338) & (sk[110]) & (g474) & (!g475)) + ((!g338) & (sk[110]) & (g474) & (g475)) + ((g338) & (!sk[110]) & (!g474) & (!g475)) + ((g338) & (!sk[110]) & (!g474) & (g475)) + ((g338) & (!sk[110]) & (g474) & (!g475)) + ((g338) & (!sk[110]) & (g474) & (g475)));
	assign g477 = (((!sk[111]) & (g48) & (!g115)) + ((!sk[111]) & (g48) & (g115)) + ((sk[111]) & (!g48) & (g115)) + ((sk[111]) & (g48) & (!g115)) + ((sk[111]) & (g48) & (g115)));
	assign g478 = (((!sk[112]) & (g48) & (!g124)) + ((!sk[112]) & (g48) & (g124)) + ((sk[112]) & (!g48) & (g124)));
	assign g479 = (((!sk[113]) & (!g112) & (!g323) & (g477) & (g478)) + ((!sk[113]) & (!g112) & (g323) & (!g477) & (!g478)) + ((!sk[113]) & (!g112) & (g323) & (!g477) & (g478)) + ((!sk[113]) & (!g112) & (g323) & (g477) & (!g478)) + ((!sk[113]) & (!g112) & (g323) & (g477) & (g478)) + ((!sk[113]) & (g112) & (!g323) & (g477) & (!g478)) + ((!sk[113]) & (g112) & (!g323) & (g477) & (g478)) + ((!sk[113]) & (g112) & (g323) & (!g477) & (!g478)) + ((!sk[113]) & (g112) & (g323) & (!g477) & (g478)) + ((!sk[113]) & (g112) & (g323) & (g477) & (!g478)) + ((!sk[113]) & (g112) & (g323) & (g477) & (g478)) + ((sk[113]) & (!g112) & (!g323) & (!g477) & (!g478)) + ((sk[113]) & (!g112) & (!g323) & (!g477) & (g478)) + ((sk[113]) & (!g112) & (!g323) & (g477) & (!g478)) + ((sk[113]) & (!g112) & (!g323) & (g477) & (g478)) + ((sk[113]) & (!g112) & (g323) & (g477) & (!g478)) + ((sk[113]) & (!g112) & (g323) & (g477) & (g478)) + ((sk[113]) & (g112) & (!g323) & (g477) & (!g478)) + ((sk[113]) & (g112) & (g323) & (g477) & (!g478)));
	assign g480 = (((!g112) & (sk[114]) & (g323) & (!g464)) + ((g112) & (!sk[114]) & (!g323) & (!g464)) + ((g112) & (!sk[114]) & (!g323) & (g464)) + ((g112) & (!sk[114]) & (g323) & (!g464)) + ((g112) & (!sk[114]) & (g323) & (g464)) + ((g112) & (sk[114]) & (!g323) & (!g464)) + ((g112) & (sk[114]) & (g323) & (!g464)));
	assign g481 = (((!sk[115]) & (g48) & (!g122)) + ((!sk[115]) & (g48) & (g122)) + ((sk[115]) & (!g48) & (g122)) + ((sk[115]) & (g48) & (!g122)) + ((sk[115]) & (g48) & (g122)));
	assign g482 = (((g323) & (!sk[116]) & (!g481) & (!g474)) + ((g323) & (!sk[116]) & (!g481) & (g474)) + ((g323) & (!sk[116]) & (g481) & (!g474)) + ((g323) & (!sk[116]) & (g481) & (g474)) + ((g323) & (sk[116]) & (!g481) & (!g474)) + ((g323) & (sk[116]) & (!g481) & (g474)) + ((g323) & (sk[116]) & (g481) & (g474)));
	assign g483 = (((!i_8_) & (!g88) & (!g112) & (!g460) & (!g470) & (!g475)) + ((!i_8_) & (!g88) & (!g112) & (!g460) & (!g470) & (g475)) + ((!i_8_) & (!g88) & (!g112) & (!g460) & (g470) & (!g475)) + ((!i_8_) & (!g88) & (!g112) & (!g460) & (g470) & (g475)) + ((!i_8_) & (!g88) & (!g112) & (g460) & (!g470) & (!g475)) + ((!i_8_) & (!g88) & (!g112) & (g460) & (!g470) & (g475)) + ((!i_8_) & (!g88) & (!g112) & (g460) & (g470) & (!g475)) + ((!i_8_) & (!g88) & (!g112) & (g460) & (g470) & (g475)) + ((!i_8_) & (!g88) & (g112) & (!g460) & (!g470) & (g475)) + ((!i_8_) & (g88) & (!g112) & (!g460) & (!g470) & (!g475)) + ((!i_8_) & (g88) & (!g112) & (!g460) & (!g470) & (g475)) + ((!i_8_) & (g88) & (!g112) & (!g460) & (g470) & (!g475)) + ((!i_8_) & (g88) & (!g112) & (!g460) & (g470) & (g475)) + ((!i_8_) & (g88) & (!g112) & (g460) & (!g470) & (!g475)) + ((!i_8_) & (g88) & (!g112) & (g460) & (!g470) & (g475)) + ((!i_8_) & (g88) & (!g112) & (g460) & (g470) & (!g475)) + ((!i_8_) & (g88) & (!g112) & (g460) & (g470) & (g475)) + ((!i_8_) & (g88) & (g112) & (!g460) & (!g470) & (g475)) + ((i_8_) & (!g88) & (!g112) & (!g460) & (!g470) & (!g475)) + ((i_8_) & (!g88) & (!g112) & (!g460) & (!g470) & (g475)) + ((i_8_) & (!g88) & (!g112) & (!g460) & (g470) & (!g475)) + ((i_8_) & (!g88) & (!g112) & (!g460) & (g470) & (g475)) + ((i_8_) & (!g88) & (!g112) & (g460) & (!g470) & (!g475)) + ((i_8_) & (!g88) & (!g112) & (g460) & (!g470) & (g475)) + ((i_8_) & (!g88) & (!g112) & (g460) & (g470) & (!g475)) + ((i_8_) & (!g88) & (!g112) & (g460) & (g470) & (g475)) + ((i_8_) & (!g88) & (g112) & (!g460) & (!g470) & (g475)) + ((i_8_) & (g88) & (!g112) & (!g460) & (!g470) & (!g475)) + ((i_8_) & (g88) & (!g112) & (!g460) & (!g470) & (g475)) + ((i_8_) & (g88) & (!g112) & (g460) & (!g470) & (!g475)) + ((i_8_) & (g88) & (!g112) & (g460) & (!g470) & (g475)) + ((i_8_) & (g88) & (g112) & (!g460) & (!g470) & (g475)));
	assign g484 = (((!sk[118]) & (!g476) & (!g479) & (!g480) & (!g482) & (g483)) + ((!sk[118]) & (!g476) & (!g479) & (!g480) & (g482) & (g483)) + ((!sk[118]) & (!g476) & (!g479) & (g480) & (!g482) & (g483)) + ((!sk[118]) & (!g476) & (!g479) & (g480) & (g482) & (g483)) + ((!sk[118]) & (!g476) & (g479) & (!g480) & (!g482) & (g483)) + ((!sk[118]) & (!g476) & (g479) & (!g480) & (g482) & (g483)) + ((!sk[118]) & (!g476) & (g479) & (g480) & (!g482) & (g483)) + ((!sk[118]) & (!g476) & (g479) & (g480) & (g482) & (g483)) + ((!sk[118]) & (g476) & (!g479) & (!g480) & (!g482) & (!g483)) + ((!sk[118]) & (g476) & (!g479) & (!g480) & (!g482) & (g483)) + ((!sk[118]) & (g476) & (!g479) & (!g480) & (g482) & (!g483)) + ((!sk[118]) & (g476) & (!g479) & (!g480) & (g482) & (g483)) + ((!sk[118]) & (g476) & (!g479) & (g480) & (!g482) & (!g483)) + ((!sk[118]) & (g476) & (!g479) & (g480) & (!g482) & (g483)) + ((!sk[118]) & (g476) & (!g479) & (g480) & (g482) & (!g483)) + ((!sk[118]) & (g476) & (!g479) & (g480) & (g482) & (g483)) + ((!sk[118]) & (g476) & (g479) & (!g480) & (!g482) & (!g483)) + ((!sk[118]) & (g476) & (g479) & (!g480) & (!g482) & (g483)) + ((!sk[118]) & (g476) & (g479) & (!g480) & (g482) & (!g483)) + ((!sk[118]) & (g476) & (g479) & (!g480) & (g482) & (g483)) + ((!sk[118]) & (g476) & (g479) & (g480) & (!g482) & (!g483)) + ((!sk[118]) & (g476) & (g479) & (g480) & (!g482) & (g483)) + ((!sk[118]) & (g476) & (g479) & (g480) & (g482) & (!g483)) + ((!sk[118]) & (g476) & (g479) & (g480) & (g482) & (g483)) + ((sk[118]) & (!g476) & (g479) & (!g480) & (!g482) & (g483)));
	assign g485 = (((!g122) & (sk[119]) & (g461)) + ((g122) & (!sk[119]) & (!g461)) + ((g122) & (!sk[119]) & (g461)));
	assign g486 = (((g145) & (!g485) & (!sk[120]) & (!g475)) + ((g145) & (!g485) & (!sk[120]) & (g475)) + ((g145) & (!g485) & (sk[120]) & (!g475)) + ((g145) & (g485) & (!sk[120]) & (!g475)) + ((g145) & (g485) & (!sk[120]) & (g475)) + ((g145) & (g485) & (sk[120]) & (!g475)) + ((g145) & (g485) & (sk[120]) & (g475)));
	assign g487 = (((!sk[121]) & (g115) & (!g461)) + ((!sk[121]) & (g115) & (g461)) + ((sk[121]) & (!g115) & (g461)));
	assign g488 = (((g145) & (!g487) & (!sk[122]) & (!g462)) + ((g145) & (!g487) & (!sk[122]) & (g462)) + ((g145) & (!g487) & (sk[122]) & (!g462)) + ((g145) & (g487) & (!sk[122]) & (!g462)) + ((g145) & (g487) & (!sk[122]) & (g462)) + ((g145) & (g487) & (sk[122]) & (!g462)) + ((g145) & (g487) & (sk[122]) & (g462)));
	assign g489 = (((!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!g48) & (g136)) + ((!i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!g48) & (g136)) + ((!i_11_) & (i_9_) & (i_10_) & (i_15_) & (!g48) & (g136)) + ((i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (!g48) & (g136)) + ((i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!g48) & (g136)) + ((i_11_) & (i_9_) & (i_10_) & (i_15_) & (!g48) & (g136)));
	assign g490 = (((!g463) & (g473) & (g484) & (!g486) & (!g488) & (!g489)));
	assign g491 = (((!sk[125]) & (g112) & (!g485)) + ((!sk[125]) & (g112) & (g485)) + ((sk[125]) & (!g112) & (!g485)) + ((sk[125]) & (!g112) & (g485)) + ((sk[125]) & (g112) & (!g485)));
	assign g492 = (((!sk[126]) & (!g59) & (!g135) & (g474) & (g460)) + ((!sk[126]) & (!g59) & (g135) & (!g474) & (!g460)) + ((!sk[126]) & (!g59) & (g135) & (!g474) & (g460)) + ((!sk[126]) & (!g59) & (g135) & (g474) & (!g460)) + ((!sk[126]) & (!g59) & (g135) & (g474) & (g460)) + ((!sk[126]) & (g59) & (!g135) & (g474) & (!g460)) + ((!sk[126]) & (g59) & (!g135) & (g474) & (g460)) + ((!sk[126]) & (g59) & (g135) & (!g474) & (!g460)) + ((!sk[126]) & (g59) & (g135) & (!g474) & (g460)) + ((!sk[126]) & (g59) & (g135) & (g474) & (!g460)) + ((!sk[126]) & (g59) & (g135) & (g474) & (g460)) + ((sk[126]) & (!g59) & (!g135) & (!g474) & (!g460)) + ((sk[126]) & (!g59) & (!g135) & (!g474) & (g460)) + ((sk[126]) & (!g59) & (!g135) & (g474) & (!g460)) + ((sk[126]) & (!g59) & (!g135) & (g474) & (g460)) + ((sk[126]) & (!g59) & (g135) & (!g474) & (!g460)) + ((sk[126]) & (!g59) & (g135) & (g474) & (!g460)) + ((sk[126]) & (g59) & (!g135) & (!g474) & (!g460)) + ((sk[126]) & (g59) & (!g135) & (!g474) & (g460)) + ((sk[126]) & (g59) & (g135) & (!g474) & (!g460)));
	assign g493 = (((!g99) & (!g118) & (!g464) & (!g467) & (!sk[127]) & (g468)) + ((!g99) & (!g118) & (!g464) & (!g467) & (sk[127]) & (!g468)) + ((!g99) & (!g118) & (!g464) & (!g467) & (sk[127]) & (g468)) + ((!g99) & (!g118) & (!g464) & (g467) & (!sk[127]) & (g468)) + ((!g99) & (!g118) & (!g464) & (g467) & (sk[127]) & (!g468)) + ((!g99) & (!g118) & (!g464) & (g467) & (sk[127]) & (g468)) + ((!g99) & (!g118) & (g464) & (!g467) & (!sk[127]) & (g468)) + ((!g99) & (!g118) & (g464) & (!g467) & (sk[127]) & (!g468)) + ((!g99) & (!g118) & (g464) & (!g467) & (sk[127]) & (g468)) + ((!g99) & (!g118) & (g464) & (g467) & (!sk[127]) & (g468)) + ((!g99) & (!g118) & (g464) & (g467) & (sk[127]) & (!g468)) + ((!g99) & (!g118) & (g464) & (g467) & (sk[127]) & (g468)) + ((!g99) & (g118) & (!g464) & (!g467) & (!sk[127]) & (g468)) + ((!g99) & (g118) & (!g464) & (g467) & (!sk[127]) & (g468)) + ((!g99) & (g118) & (g464) & (!g467) & (!sk[127]) & (g468)) + ((!g99) & (g118) & (g464) & (g467) & (!sk[127]) & (g468)) + ((!g99) & (g118) & (g464) & (g467) & (sk[127]) & (g468)) + ((g99) & (!g118) & (!g464) & (!g467) & (!sk[127]) & (!g468)) + ((g99) & (!g118) & (!g464) & (!g467) & (!sk[127]) & (g468)) + ((g99) & (!g118) & (!g464) & (g467) & (!sk[127]) & (!g468)) + ((g99) & (!g118) & (!g464) & (g467) & (!sk[127]) & (g468)) + ((g99) & (!g118) & (g464) & (!g467) & (!sk[127]) & (!g468)) + ((g99) & (!g118) & (g464) & (!g467) & (!sk[127]) & (g468)) + ((g99) & (!g118) & (g464) & (!g467) & (sk[127]) & (!g468)) + ((g99) & (!g118) & (g464) & (!g467) & (sk[127]) & (g468)) + ((g99) & (!g118) & (g464) & (g467) & (!sk[127]) & (!g468)) + ((g99) & (!g118) & (g464) & (g467) & (!sk[127]) & (g468)) + ((g99) & (!g118) & (g464) & (g467) & (sk[127]) & (!g468)) + ((g99) & (!g118) & (g464) & (g467) & (sk[127]) & (g468)) + ((g99) & (g118) & (!g464) & (!g467) & (!sk[127]) & (!g468)) + ((g99) & (g118) & (!g464) & (!g467) & (!sk[127]) & (g468)) + ((g99) & (g118) & (!g464) & (g467) & (!sk[127]) & (!g468)) + ((g99) & (g118) & (!g464) & (g467) & (!sk[127]) & (g468)) + ((g99) & (g118) & (g464) & (!g467) & (!sk[127]) & (!g468)) + ((g99) & (g118) & (g464) & (!g467) & (!sk[127]) & (g468)) + ((g99) & (g118) & (g464) & (g467) & (!sk[127]) & (!g468)) + ((g99) & (g118) & (g464) & (g467) & (!sk[127]) & (g468)) + ((g99) & (g118) & (g464) & (g467) & (sk[127]) & (g468)));
	assign g494 = (((!g59) & (!g429) & (!sk[0]) & (g465) & (g493)) + ((!g59) & (!g429) & (sk[0]) & (!g465) & (g493)) + ((!g59) & (!g429) & (sk[0]) & (g465) & (g493)) + ((!g59) & (g429) & (!sk[0]) & (!g465) & (!g493)) + ((!g59) & (g429) & (!sk[0]) & (!g465) & (g493)) + ((!g59) & (g429) & (!sk[0]) & (g465) & (!g493)) + ((!g59) & (g429) & (!sk[0]) & (g465) & (g493)) + ((!g59) & (g429) & (sk[0]) & (g465) & (g493)) + ((g59) & (!g429) & (!sk[0]) & (g465) & (!g493)) + ((g59) & (!g429) & (!sk[0]) & (g465) & (g493)) + ((g59) & (!g429) & (sk[0]) & (g465) & (g493)) + ((g59) & (g429) & (!sk[0]) & (!g465) & (!g493)) + ((g59) & (g429) & (!sk[0]) & (!g465) & (g493)) + ((g59) & (g429) & (!sk[0]) & (g465) & (!g493)) + ((g59) & (g429) & (!sk[0]) & (g465) & (g493)) + ((g59) & (g429) & (sk[0]) & (g465) & (g493)));
	assign g495 = (((!sk[1]) & (g30) & (!g110)) + ((!sk[1]) & (g30) & (g110)) + ((sk[1]) & (g30) & (g110)));
	assign g496 = (((!g124) & (!sk[2]) & (!g461) & (g474) & (g495)) + ((!g124) & (!sk[2]) & (g461) & (!g474) & (!g495)) + ((!g124) & (!sk[2]) & (g461) & (!g474) & (g495)) + ((!g124) & (!sk[2]) & (g461) & (g474) & (!g495)) + ((!g124) & (!sk[2]) & (g461) & (g474) & (g495)) + ((!g124) & (sk[2]) & (!g461) & (g474) & (g495)) + ((!g124) & (sk[2]) & (g461) & (g474) & (g495)) + ((g124) & (!sk[2]) & (!g461) & (g474) & (!g495)) + ((g124) & (!sk[2]) & (!g461) & (g474) & (g495)) + ((g124) & (!sk[2]) & (g461) & (!g474) & (!g495)) + ((g124) & (!sk[2]) & (g461) & (!g474) & (g495)) + ((g124) & (!sk[2]) & (g461) & (g474) & (!g495)) + ((g124) & (!sk[2]) & (g461) & (g474) & (g495)) + ((g124) & (sk[2]) & (!g461) & (g474) & (g495)) + ((g124) & (sk[2]) & (g461) & (!g474) & (g495)) + ((g124) & (sk[2]) & (g461) & (g474) & (g495)));
	assign g497 = (((g109) & (!sk[3]) & (!g465) & (!g462)) + ((g109) & (!sk[3]) & (!g465) & (g462)) + ((g109) & (!sk[3]) & (g465) & (!g462)) + ((g109) & (!sk[3]) & (g465) & (g462)) + ((g109) & (sk[3]) & (!g465) & (!g462)) + ((g109) & (sk[3]) & (!g465) & (g462)) + ((g109) & (sk[3]) & (g465) & (!g462)));
	assign g498 = (((!i_8_) & (!i_7_) & (!g400) & (!sk[4]) & (!g467) & (g487)) + ((!i_8_) & (!i_7_) & (!g400) & (!sk[4]) & (g467) & (g487)) + ((!i_8_) & (!i_7_) & (g400) & (!sk[4]) & (!g467) & (g487)) + ((!i_8_) & (!i_7_) & (g400) & (!sk[4]) & (g467) & (g487)) + ((!i_8_) & (!i_7_) & (g400) & (sk[4]) & (!g467) & (g487)) + ((!i_8_) & (!i_7_) & (g400) & (sk[4]) & (g467) & (g487)) + ((!i_8_) & (i_7_) & (!g400) & (!sk[4]) & (!g467) & (g487)) + ((!i_8_) & (i_7_) & (!g400) & (!sk[4]) & (g467) & (g487)) + ((!i_8_) & (i_7_) & (g400) & (!sk[4]) & (!g467) & (g487)) + ((!i_8_) & (i_7_) & (g400) & (!sk[4]) & (g467) & (g487)) + ((!i_8_) & (i_7_) & (g400) & (sk[4]) & (!g467) & (!g487)) + ((!i_8_) & (i_7_) & (g400) & (sk[4]) & (!g467) & (g487)) + ((i_8_) & (!i_7_) & (!g400) & (!sk[4]) & (!g467) & (!g487)) + ((i_8_) & (!i_7_) & (!g400) & (!sk[4]) & (!g467) & (g487)) + ((i_8_) & (!i_7_) & (!g400) & (!sk[4]) & (g467) & (!g487)) + ((i_8_) & (!i_7_) & (!g400) & (!sk[4]) & (g467) & (g487)) + ((i_8_) & (!i_7_) & (g400) & (!sk[4]) & (!g467) & (!g487)) + ((i_8_) & (!i_7_) & (g400) & (!sk[4]) & (!g467) & (g487)) + ((i_8_) & (!i_7_) & (g400) & (!sk[4]) & (g467) & (!g487)) + ((i_8_) & (!i_7_) & (g400) & (!sk[4]) & (g467) & (g487)) + ((i_8_) & (i_7_) & (!g400) & (!sk[4]) & (!g467) & (!g487)) + ((i_8_) & (i_7_) & (!g400) & (!sk[4]) & (!g467) & (g487)) + ((i_8_) & (i_7_) & (!g400) & (!sk[4]) & (g467) & (!g487)) + ((i_8_) & (i_7_) & (!g400) & (!sk[4]) & (g467) & (g487)) + ((i_8_) & (i_7_) & (g400) & (!sk[4]) & (!g467) & (!g487)) + ((i_8_) & (i_7_) & (g400) & (!sk[4]) & (!g467) & (g487)) + ((i_8_) & (i_7_) & (g400) & (!sk[4]) & (g467) & (!g487)) + ((i_8_) & (i_7_) & (g400) & (!sk[4]) & (g467) & (g487)));
	assign g499 = (((!g323) & (!sk[5]) & (!g478) & (!g496) & (!g497) & (g498)) + ((!g323) & (!sk[5]) & (!g478) & (!g496) & (g497) & (g498)) + ((!g323) & (!sk[5]) & (!g478) & (g496) & (!g497) & (g498)) + ((!g323) & (!sk[5]) & (!g478) & (g496) & (g497) & (g498)) + ((!g323) & (!sk[5]) & (g478) & (!g496) & (!g497) & (g498)) + ((!g323) & (!sk[5]) & (g478) & (!g496) & (g497) & (g498)) + ((!g323) & (!sk[5]) & (g478) & (g496) & (!g497) & (g498)) + ((!g323) & (!sk[5]) & (g478) & (g496) & (g497) & (g498)) + ((!g323) & (sk[5]) & (!g478) & (!g496) & (!g497) & (!g498)) + ((!g323) & (sk[5]) & (g478) & (!g496) & (!g497) & (!g498)) + ((g323) & (!sk[5]) & (!g478) & (!g496) & (!g497) & (!g498)) + ((g323) & (!sk[5]) & (!g478) & (!g496) & (!g497) & (g498)) + ((g323) & (!sk[5]) & (!g478) & (!g496) & (g497) & (!g498)) + ((g323) & (!sk[5]) & (!g478) & (!g496) & (g497) & (g498)) + ((g323) & (!sk[5]) & (!g478) & (g496) & (!g497) & (!g498)) + ((g323) & (!sk[5]) & (!g478) & (g496) & (!g497) & (g498)) + ((g323) & (!sk[5]) & (!g478) & (g496) & (g497) & (!g498)) + ((g323) & (!sk[5]) & (!g478) & (g496) & (g497) & (g498)) + ((g323) & (!sk[5]) & (g478) & (!g496) & (!g497) & (!g498)) + ((g323) & (!sk[5]) & (g478) & (!g496) & (!g497) & (g498)) + ((g323) & (!sk[5]) & (g478) & (!g496) & (g497) & (!g498)) + ((g323) & (!sk[5]) & (g478) & (!g496) & (g497) & (g498)) + ((g323) & (!sk[5]) & (g478) & (g496) & (!g497) & (!g498)) + ((g323) & (!sk[5]) & (g478) & (g496) & (!g497) & (g498)) + ((g323) & (!sk[5]) & (g478) & (g496) & (g497) & (!g498)) + ((g323) & (!sk[5]) & (g478) & (g496) & (g497) & (g498)) + ((g323) & (sk[5]) & (!g478) & (!g496) & (!g497) & (!g498)));
	assign g500 = (((g118) & (!g478) & (!sk[6]) & (!g487)) + ((g118) & (!g478) & (!sk[6]) & (g487)) + ((g118) & (!g478) & (sk[6]) & (g487)) + ((g118) & (g478) & (!sk[6]) & (!g487)) + ((g118) & (g478) & (!sk[6]) & (g487)) + ((g118) & (g478) & (sk[6]) & (!g487)) + ((g118) & (g478) & (sk[6]) & (g487)));
	assign g501 = (((!sk[7]) & (!g18) & (!g118) & (g228) & (g461)) + ((!sk[7]) & (!g18) & (g118) & (!g228) & (!g461)) + ((!sk[7]) & (!g18) & (g118) & (!g228) & (g461)) + ((!sk[7]) & (!g18) & (g118) & (g228) & (!g461)) + ((!sk[7]) & (!g18) & (g118) & (g228) & (g461)) + ((!sk[7]) & (g18) & (!g118) & (g228) & (!g461)) + ((!sk[7]) & (g18) & (!g118) & (g228) & (g461)) + ((!sk[7]) & (g18) & (g118) & (!g228) & (!g461)) + ((!sk[7]) & (g18) & (g118) & (!g228) & (g461)) + ((!sk[7]) & (g18) & (g118) & (g228) & (!g461)) + ((!sk[7]) & (g18) & (g118) & (g228) & (g461)) + ((sk[7]) & (!g18) & (g118) & (!g228) & (g461)) + ((sk[7]) & (!g18) & (g118) & (g228) & (g461)) + ((sk[7]) & (g18) & (g118) & (g228) & (g461)));
	assign g502 = (((!g22) & (!g88) & (!sk[8]) & (g124) & (g461)) + ((!g22) & (g88) & (!sk[8]) & (!g124) & (!g461)) + ((!g22) & (g88) & (!sk[8]) & (!g124) & (g461)) + ((!g22) & (g88) & (!sk[8]) & (g124) & (!g461)) + ((!g22) & (g88) & (!sk[8]) & (g124) & (g461)) + ((!g22) & (g88) & (sk[8]) & (g124) & (g461)) + ((g22) & (!g88) & (!sk[8]) & (g124) & (!g461)) + ((g22) & (!g88) & (!sk[8]) & (g124) & (g461)) + ((g22) & (g88) & (!sk[8]) & (!g124) & (!g461)) + ((g22) & (g88) & (!sk[8]) & (!g124) & (g461)) + ((g22) & (g88) & (!sk[8]) & (g124) & (!g461)) + ((g22) & (g88) & (!sk[8]) & (g124) & (g461)) + ((g22) & (g88) & (sk[8]) & (!g124) & (g461)) + ((g22) & (g88) & (sk[8]) & (g124) & (g461)));
	assign g503 = (((!sk[9]) & (!g22) & (!g134) & (!g93) & (!g124) & (g461)) + ((!sk[9]) & (!g22) & (!g134) & (!g93) & (g124) & (g461)) + ((!sk[9]) & (!g22) & (!g134) & (g93) & (!g124) & (g461)) + ((!sk[9]) & (!g22) & (!g134) & (g93) & (g124) & (g461)) + ((!sk[9]) & (!g22) & (g134) & (!g93) & (!g124) & (g461)) + ((!sk[9]) & (!g22) & (g134) & (!g93) & (g124) & (g461)) + ((!sk[9]) & (!g22) & (g134) & (g93) & (!g124) & (g461)) + ((!sk[9]) & (!g22) & (g134) & (g93) & (g124) & (g461)) + ((!sk[9]) & (g22) & (!g134) & (!g93) & (!g124) & (!g461)) + ((!sk[9]) & (g22) & (!g134) & (!g93) & (!g124) & (g461)) + ((!sk[9]) & (g22) & (!g134) & (!g93) & (g124) & (!g461)) + ((!sk[9]) & (g22) & (!g134) & (!g93) & (g124) & (g461)) + ((!sk[9]) & (g22) & (!g134) & (g93) & (!g124) & (!g461)) + ((!sk[9]) & (g22) & (!g134) & (g93) & (!g124) & (g461)) + ((!sk[9]) & (g22) & (!g134) & (g93) & (g124) & (!g461)) + ((!sk[9]) & (g22) & (!g134) & (g93) & (g124) & (g461)) + ((!sk[9]) & (g22) & (g134) & (!g93) & (!g124) & (!g461)) + ((!sk[9]) & (g22) & (g134) & (!g93) & (!g124) & (g461)) + ((!sk[9]) & (g22) & (g134) & (!g93) & (g124) & (!g461)) + ((!sk[9]) & (g22) & (g134) & (!g93) & (g124) & (g461)) + ((!sk[9]) & (g22) & (g134) & (g93) & (!g124) & (!g461)) + ((!sk[9]) & (g22) & (g134) & (g93) & (!g124) & (g461)) + ((!sk[9]) & (g22) & (g134) & (g93) & (g124) & (!g461)) + ((!sk[9]) & (g22) & (g134) & (g93) & (g124) & (g461)) + ((sk[9]) & (!g22) & (g134) & (!g93) & (!g124) & (g461)) + ((sk[9]) & (!g22) & (g134) & (!g93) & (g124) & (g461)) + ((sk[9]) & (!g22) & (g134) & (g93) & (g124) & (g461)) + ((sk[9]) & (g22) & (g134) & (!g93) & (!g124) & (g461)) + ((sk[9]) & (g22) & (g134) & (!g93) & (g124) & (g461)) + ((sk[9]) & (g22) & (g134) & (g93) & (!g124) & (g461)) + ((sk[9]) & (g22) & (g134) & (g93) & (g124) & (g461)));
	assign g504 = (((!g134) & (!g149) & (!g99) & (!g423) & (!g481) & (!g467)) + ((!g134) & (!g149) & (!g99) & (!g423) & (!g481) & (g467)) + ((!g134) & (!g149) & (!g99) & (!g423) & (g481) & (!g467)) + ((!g134) & (!g149) & (!g99) & (!g423) & (g481) & (g467)) + ((!g134) & (!g149) & (!g99) & (g423) & (g481) & (g467)) + ((!g134) & (!g149) & (g99) & (!g423) & (g481) & (!g467)) + ((!g134) & (!g149) & (g99) & (!g423) & (g481) & (g467)) + ((!g134) & (!g149) & (g99) & (g423) & (g481) & (g467)) + ((!g134) & (g149) & (!g99) & (!g423) & (g481) & (!g467)) + ((!g134) & (g149) & (!g99) & (!g423) & (g481) & (g467)) + ((!g134) & (g149) & (!g99) & (g423) & (g481) & (g467)) + ((!g134) & (g149) & (g99) & (!g423) & (g481) & (!g467)) + ((!g134) & (g149) & (g99) & (!g423) & (g481) & (g467)) + ((!g134) & (g149) & (g99) & (g423) & (g481) & (g467)) + ((g134) & (!g149) & (!g99) & (!g423) & (g481) & (!g467)) + ((g134) & (!g149) & (!g99) & (!g423) & (g481) & (g467)) + ((g134) & (!g149) & (!g99) & (g423) & (g481) & (g467)) + ((g134) & (!g149) & (g99) & (!g423) & (g481) & (!g467)) + ((g134) & (!g149) & (g99) & (!g423) & (g481) & (g467)) + ((g134) & (!g149) & (g99) & (g423) & (g481) & (g467)) + ((g134) & (g149) & (!g99) & (!g423) & (g481) & (!g467)) + ((g134) & (g149) & (!g99) & (!g423) & (g481) & (g467)) + ((g134) & (g149) & (!g99) & (g423) & (g481) & (g467)) + ((g134) & (g149) & (g99) & (!g423) & (g481) & (!g467)) + ((g134) & (g149) & (g99) & (!g423) & (g481) & (g467)) + ((g134) & (g149) & (g99) & (g423) & (g481) & (g467)));
	assign g505 = (((!g500) & (!g501) & (!g502) & (!g503) & (!sk[11]) & (g504)) + ((!g500) & (!g501) & (!g502) & (!g503) & (sk[11]) & (g504)) + ((!g500) & (!g501) & (!g502) & (g503) & (!sk[11]) & (g504)) + ((!g500) & (!g501) & (g502) & (!g503) & (!sk[11]) & (g504)) + ((!g500) & (!g501) & (g502) & (g503) & (!sk[11]) & (g504)) + ((!g500) & (g501) & (!g502) & (!g503) & (!sk[11]) & (g504)) + ((!g500) & (g501) & (!g502) & (g503) & (!sk[11]) & (g504)) + ((!g500) & (g501) & (g502) & (!g503) & (!sk[11]) & (g504)) + ((!g500) & (g501) & (g502) & (g503) & (!sk[11]) & (g504)) + ((g500) & (!g501) & (!g502) & (!g503) & (!sk[11]) & (!g504)) + ((g500) & (!g501) & (!g502) & (!g503) & (!sk[11]) & (g504)) + ((g500) & (!g501) & (!g502) & (g503) & (!sk[11]) & (!g504)) + ((g500) & (!g501) & (!g502) & (g503) & (!sk[11]) & (g504)) + ((g500) & (!g501) & (g502) & (!g503) & (!sk[11]) & (!g504)) + ((g500) & (!g501) & (g502) & (!g503) & (!sk[11]) & (g504)) + ((g500) & (!g501) & (g502) & (g503) & (!sk[11]) & (!g504)) + ((g500) & (!g501) & (g502) & (g503) & (!sk[11]) & (g504)) + ((g500) & (g501) & (!g502) & (!g503) & (!sk[11]) & (!g504)) + ((g500) & (g501) & (!g502) & (!g503) & (!sk[11]) & (g504)) + ((g500) & (g501) & (!g502) & (g503) & (!sk[11]) & (!g504)) + ((g500) & (g501) & (!g502) & (g503) & (!sk[11]) & (g504)) + ((g500) & (g501) & (g502) & (!g503) & (!sk[11]) & (!g504)) + ((g500) & (g501) & (g502) & (!g503) & (!sk[11]) & (g504)) + ((g500) & (g501) & (g502) & (g503) & (!sk[11]) & (!g504)) + ((g500) & (g501) & (g502) & (g503) & (!sk[11]) & (g504)));
	assign g506 = (((!sk[12]) & (g22) & (!g461)) + ((!sk[12]) & (g22) & (g461)) + ((sk[12]) & (g22) & (g461)));
	assign g507 = (((!sk[13]) & (!i_8_) & (!g108) & (g506) & (g470)) + ((!sk[13]) & (!i_8_) & (g108) & (!g506) & (!g470)) + ((!sk[13]) & (!i_8_) & (g108) & (!g506) & (g470)) + ((!sk[13]) & (!i_8_) & (g108) & (g506) & (!g470)) + ((!sk[13]) & (!i_8_) & (g108) & (g506) & (g470)) + ((!sk[13]) & (i_8_) & (!g108) & (g506) & (!g470)) + ((!sk[13]) & (i_8_) & (!g108) & (g506) & (g470)) + ((!sk[13]) & (i_8_) & (g108) & (!g506) & (!g470)) + ((!sk[13]) & (i_8_) & (g108) & (!g506) & (g470)) + ((!sk[13]) & (i_8_) & (g108) & (g506) & (!g470)) + ((!sk[13]) & (i_8_) & (g108) & (g506) & (g470)) + ((sk[13]) & (!i_8_) & (g108) & (!g506) & (g470)) + ((sk[13]) & (!i_8_) & (g108) & (g506) & (!g470)) + ((sk[13]) & (!i_8_) & (g108) & (g506) & (g470)) + ((sk[13]) & (i_8_) & (g108) & (g506) & (!g470)) + ((sk[13]) & (i_8_) & (g108) & (g506) & (g470)));
	assign g508 = (((!g136) & (!sk[14]) & (!g124) & (g115) & (g461)) + ((!g136) & (!sk[14]) & (g124) & (!g115) & (!g461)) + ((!g136) & (!sk[14]) & (g124) & (!g115) & (g461)) + ((!g136) & (!sk[14]) & (g124) & (g115) & (!g461)) + ((!g136) & (!sk[14]) & (g124) & (g115) & (g461)) + ((g136) & (!sk[14]) & (!g124) & (g115) & (!g461)) + ((g136) & (!sk[14]) & (!g124) & (g115) & (g461)) + ((g136) & (!sk[14]) & (g124) & (!g115) & (!g461)) + ((g136) & (!sk[14]) & (g124) & (!g115) & (g461)) + ((g136) & (!sk[14]) & (g124) & (g115) & (!g461)) + ((g136) & (!sk[14]) & (g124) & (g115) & (g461)) + ((g136) & (sk[14]) & (!g124) & (!g115) & (g461)) + ((g136) & (sk[14]) & (g124) & (!g115) & (g461)) + ((g136) & (sk[14]) & (g124) & (g115) & (g461)));
	assign g509 = (((!i_8_) & (!sk[15]) & (!g108) & (!g124) & (!g115) & (g461)) + ((!i_8_) & (!sk[15]) & (!g108) & (!g124) & (g115) & (g461)) + ((!i_8_) & (!sk[15]) & (!g108) & (g124) & (!g115) & (g461)) + ((!i_8_) & (!sk[15]) & (!g108) & (g124) & (g115) & (g461)) + ((!i_8_) & (!sk[15]) & (g108) & (!g124) & (!g115) & (g461)) + ((!i_8_) & (!sk[15]) & (g108) & (!g124) & (g115) & (g461)) + ((!i_8_) & (!sk[15]) & (g108) & (g124) & (!g115) & (g461)) + ((!i_8_) & (!sk[15]) & (g108) & (g124) & (g115) & (g461)) + ((!i_8_) & (sk[15]) & (g108) & (!g124) & (!g115) & (g461)) + ((!i_8_) & (sk[15]) & (g108) & (g124) & (!g115) & (g461)) + ((!i_8_) & (sk[15]) & (g108) & (g124) & (g115) & (g461)) + ((i_8_) & (!sk[15]) & (!g108) & (!g124) & (!g115) & (!g461)) + ((i_8_) & (!sk[15]) & (!g108) & (!g124) & (!g115) & (g461)) + ((i_8_) & (!sk[15]) & (!g108) & (!g124) & (g115) & (!g461)) + ((i_8_) & (!sk[15]) & (!g108) & (!g124) & (g115) & (g461)) + ((i_8_) & (!sk[15]) & (!g108) & (g124) & (!g115) & (!g461)) + ((i_8_) & (!sk[15]) & (!g108) & (g124) & (!g115) & (g461)) + ((i_8_) & (!sk[15]) & (!g108) & (g124) & (g115) & (!g461)) + ((i_8_) & (!sk[15]) & (!g108) & (g124) & (g115) & (g461)) + ((i_8_) & (!sk[15]) & (g108) & (!g124) & (!g115) & (!g461)) + ((i_8_) & (!sk[15]) & (g108) & (!g124) & (!g115) & (g461)) + ((i_8_) & (!sk[15]) & (g108) & (!g124) & (g115) & (!g461)) + ((i_8_) & (!sk[15]) & (g108) & (!g124) & (g115) & (g461)) + ((i_8_) & (!sk[15]) & (g108) & (g124) & (!g115) & (!g461)) + ((i_8_) & (!sk[15]) & (g108) & (g124) & (!g115) & (g461)) + ((i_8_) & (!sk[15]) & (g108) & (g124) & (g115) & (!g461)) + ((i_8_) & (!sk[15]) & (g108) & (g124) & (g115) & (g461)) + ((i_8_) & (sk[15]) & (g108) & (g124) & (!g115) & (g461)) + ((i_8_) & (sk[15]) & (g108) & (g124) & (g115) & (g461)));
	assign g510 = (((!sk[16]) & (!i_8_) & (!g108) & (g474) & (g475)) + ((!sk[16]) & (!i_8_) & (g108) & (!g474) & (!g475)) + ((!sk[16]) & (!i_8_) & (g108) & (!g474) & (g475)) + ((!sk[16]) & (!i_8_) & (g108) & (g474) & (!g475)) + ((!sk[16]) & (!i_8_) & (g108) & (g474) & (g475)) + ((!sk[16]) & (i_8_) & (!g108) & (g474) & (!g475)) + ((!sk[16]) & (i_8_) & (!g108) & (g474) & (g475)) + ((!sk[16]) & (i_8_) & (g108) & (!g474) & (!g475)) + ((!sk[16]) & (i_8_) & (g108) & (!g474) & (g475)) + ((!sk[16]) & (i_8_) & (g108) & (g474) & (!g475)) + ((!sk[16]) & (i_8_) & (g108) & (g474) & (g475)) + ((sk[16]) & (!i_8_) & (g108) & (!g474) & (!g475)) + ((sk[16]) & (!i_8_) & (g108) & (g474) & (!g475)) + ((sk[16]) & (!i_8_) & (g108) & (g474) & (g475)));
	assign g511 = (((!g149) & (!g109) & (!g477) & (!sk[17]) & (!g485) & (g510)) + ((!g149) & (!g109) & (!g477) & (!sk[17]) & (g485) & (g510)) + ((!g149) & (!g109) & (!g477) & (sk[17]) & (!g485) & (!g510)) + ((!g149) & (!g109) & (!g477) & (sk[17]) & (g485) & (!g510)) + ((!g149) & (!g109) & (g477) & (!sk[17]) & (!g485) & (g510)) + ((!g149) & (!g109) & (g477) & (!sk[17]) & (g485) & (g510)) + ((!g149) & (!g109) & (g477) & (sk[17]) & (!g485) & (!g510)) + ((!g149) & (!g109) & (g477) & (sk[17]) & (g485) & (!g510)) + ((!g149) & (g109) & (!g477) & (!sk[17]) & (!g485) & (g510)) + ((!g149) & (g109) & (!g477) & (!sk[17]) & (g485) & (g510)) + ((!g149) & (g109) & (g477) & (!sk[17]) & (!g485) & (g510)) + ((!g149) & (g109) & (g477) & (!sk[17]) & (g485) & (g510)) + ((!g149) & (g109) & (g477) & (sk[17]) & (!g485) & (!g510)) + ((g149) & (!g109) & (!g477) & (!sk[17]) & (!g485) & (!g510)) + ((g149) & (!g109) & (!g477) & (!sk[17]) & (!g485) & (g510)) + ((g149) & (!g109) & (!g477) & (!sk[17]) & (g485) & (!g510)) + ((g149) & (!g109) & (!g477) & (!sk[17]) & (g485) & (g510)) + ((g149) & (!g109) & (!g477) & (sk[17]) & (!g485) & (!g510)) + ((g149) & (!g109) & (g477) & (!sk[17]) & (!g485) & (!g510)) + ((g149) & (!g109) & (g477) & (!sk[17]) & (!g485) & (g510)) + ((g149) & (!g109) & (g477) & (!sk[17]) & (g485) & (!g510)) + ((g149) & (!g109) & (g477) & (!sk[17]) & (g485) & (g510)) + ((g149) & (!g109) & (g477) & (sk[17]) & (!g485) & (!g510)) + ((g149) & (g109) & (!g477) & (!sk[17]) & (!g485) & (!g510)) + ((g149) & (g109) & (!g477) & (!sk[17]) & (!g485) & (g510)) + ((g149) & (g109) & (!g477) & (!sk[17]) & (g485) & (!g510)) + ((g149) & (g109) & (!g477) & (!sk[17]) & (g485) & (g510)) + ((g149) & (g109) & (g477) & (!sk[17]) & (!g485) & (!g510)) + ((g149) & (g109) & (g477) & (!sk[17]) & (!g485) & (g510)) + ((g149) & (g109) & (g477) & (!sk[17]) & (g485) & (!g510)) + ((g149) & (g109) & (g477) & (!sk[17]) & (g485) & (g510)) + ((g149) & (g109) & (g477) & (sk[17]) & (!g485) & (!g510)));
	assign g512 = (((!g505) & (!g507) & (!sk[18]) & (!g508) & (!g509) & (g511)) + ((!g505) & (!g507) & (!sk[18]) & (!g508) & (g509) & (g511)) + ((!g505) & (!g507) & (!sk[18]) & (g508) & (!g509) & (g511)) + ((!g505) & (!g507) & (!sk[18]) & (g508) & (g509) & (g511)) + ((!g505) & (g507) & (!sk[18]) & (!g508) & (!g509) & (g511)) + ((!g505) & (g507) & (!sk[18]) & (!g508) & (g509) & (g511)) + ((!g505) & (g507) & (!sk[18]) & (g508) & (!g509) & (g511)) + ((!g505) & (g507) & (!sk[18]) & (g508) & (g509) & (g511)) + ((g505) & (!g507) & (!sk[18]) & (!g508) & (!g509) & (!g511)) + ((g505) & (!g507) & (!sk[18]) & (!g508) & (!g509) & (g511)) + ((g505) & (!g507) & (!sk[18]) & (!g508) & (g509) & (!g511)) + ((g505) & (!g507) & (!sk[18]) & (!g508) & (g509) & (g511)) + ((g505) & (!g507) & (!sk[18]) & (g508) & (!g509) & (!g511)) + ((g505) & (!g507) & (!sk[18]) & (g508) & (!g509) & (g511)) + ((g505) & (!g507) & (!sk[18]) & (g508) & (g509) & (!g511)) + ((g505) & (!g507) & (!sk[18]) & (g508) & (g509) & (g511)) + ((g505) & (!g507) & (sk[18]) & (!g508) & (!g509) & (g511)) + ((g505) & (g507) & (!sk[18]) & (!g508) & (!g509) & (!g511)) + ((g505) & (g507) & (!sk[18]) & (!g508) & (!g509) & (g511)) + ((g505) & (g507) & (!sk[18]) & (!g508) & (g509) & (!g511)) + ((g505) & (g507) & (!sk[18]) & (!g508) & (g509) & (g511)) + ((g505) & (g507) & (!sk[18]) & (g508) & (!g509) & (!g511)) + ((g505) & (g507) & (!sk[18]) & (g508) & (!g509) & (g511)) + ((g505) & (g507) & (!sk[18]) & (g508) & (g509) & (!g511)) + ((g505) & (g507) & (!sk[18]) & (g508) & (g509) & (g511)));
	assign g513 = (((!g110) & (!g111) & (!g428) & (!sk[19]) & (!g487) & (g506)) + ((!g110) & (!g111) & (!g428) & (!sk[19]) & (g487) & (g506)) + ((!g110) & (!g111) & (g428) & (!sk[19]) & (!g487) & (g506)) + ((!g110) & (!g111) & (g428) & (!sk[19]) & (g487) & (g506)) + ((!g110) & (g111) & (!g428) & (!sk[19]) & (!g487) & (g506)) + ((!g110) & (g111) & (!g428) & (!sk[19]) & (g487) & (g506)) + ((!g110) & (g111) & (g428) & (!sk[19]) & (!g487) & (g506)) + ((!g110) & (g111) & (g428) & (!sk[19]) & (g487) & (g506)) + ((!g110) & (g111) & (g428) & (sk[19]) & (g487) & (!g506)) + ((!g110) & (g111) & (g428) & (sk[19]) & (g487) & (g506)) + ((g110) & (!g111) & (!g428) & (!sk[19]) & (!g487) & (!g506)) + ((g110) & (!g111) & (!g428) & (!sk[19]) & (!g487) & (g506)) + ((g110) & (!g111) & (!g428) & (!sk[19]) & (g487) & (!g506)) + ((g110) & (!g111) & (!g428) & (!sk[19]) & (g487) & (g506)) + ((g110) & (!g111) & (g428) & (!sk[19]) & (!g487) & (!g506)) + ((g110) & (!g111) & (g428) & (!sk[19]) & (!g487) & (g506)) + ((g110) & (!g111) & (g428) & (!sk[19]) & (g487) & (!g506)) + ((g110) & (!g111) & (g428) & (!sk[19]) & (g487) & (g506)) + ((g110) & (g111) & (!g428) & (!sk[19]) & (!g487) & (!g506)) + ((g110) & (g111) & (!g428) & (!sk[19]) & (!g487) & (g506)) + ((g110) & (g111) & (!g428) & (!sk[19]) & (g487) & (!g506)) + ((g110) & (g111) & (!g428) & (!sk[19]) & (g487) & (g506)) + ((g110) & (g111) & (!g428) & (sk[19]) & (!g487) & (g506)) + ((g110) & (g111) & (!g428) & (sk[19]) & (g487) & (g506)) + ((g110) & (g111) & (g428) & (!sk[19]) & (!g487) & (!g506)) + ((g110) & (g111) & (g428) & (!sk[19]) & (!g487) & (g506)) + ((g110) & (g111) & (g428) & (!sk[19]) & (g487) & (!g506)) + ((g110) & (g111) & (g428) & (!sk[19]) & (g487) & (g506)) + ((g110) & (g111) & (g428) & (sk[19]) & (!g487) & (g506)) + ((g110) & (g111) & (g428) & (sk[19]) & (g487) & (!g506)) + ((g110) & (g111) & (g428) & (sk[19]) & (g487) & (g506)));
	assign g514 = (((!i_8_) & (!sk[20]) & (!g88) & (g108) & (g468)) + ((!i_8_) & (!sk[20]) & (g88) & (!g108) & (!g468)) + ((!i_8_) & (!sk[20]) & (g88) & (!g108) & (g468)) + ((!i_8_) & (!sk[20]) & (g88) & (g108) & (!g468)) + ((!i_8_) & (!sk[20]) & (g88) & (g108) & (g468)) + ((!i_8_) & (sk[20]) & (!g88) & (g108) & (!g468)) + ((!i_8_) & (sk[20]) & (g88) & (g108) & (!g468)) + ((i_8_) & (!sk[20]) & (!g88) & (g108) & (!g468)) + ((i_8_) & (!sk[20]) & (!g88) & (g108) & (g468)) + ((i_8_) & (!sk[20]) & (g88) & (!g108) & (!g468)) + ((i_8_) & (!sk[20]) & (g88) & (!g108) & (g468)) + ((i_8_) & (!sk[20]) & (g88) & (g108) & (!g468)) + ((i_8_) & (!sk[20]) & (g88) & (g108) & (g468)) + ((i_8_) & (sk[20]) & (!g88) & (g108) & (!g468)) + ((i_8_) & (sk[20]) & (g88) & (!g108) & (!g468)) + ((i_8_) & (sk[20]) & (g88) & (g108) & (!g468)));
	assign g515 = (((!i_8_) & (g135) & (!g485) & (!g506) & (!g468) & (!g475)) + ((!i_8_) & (g135) & (!g485) & (!g506) & (!g468) & (g475)) + ((!i_8_) & (g135) & (!g485) & (g506) & (!g468) & (!g475)) + ((!i_8_) & (g135) & (!g485) & (g506) & (!g468) & (g475)) + ((!i_8_) & (g135) & (g485) & (!g506) & (!g468) & (!g475)) + ((!i_8_) & (g135) & (g485) & (!g506) & (!g468) & (g475)) + ((!i_8_) & (g135) & (g485) & (g506) & (!g468) & (!g475)) + ((!i_8_) & (g135) & (g485) & (g506) & (!g468) & (g475)) + ((i_8_) & (g135) & (!g485) & (!g506) & (!g468) & (!g475)) + ((i_8_) & (g135) & (!g485) & (!g506) & (!g468) & (g475)) + ((i_8_) & (g135) & (!g485) & (!g506) & (g468) & (!g475)) + ((i_8_) & (g135) & (!g485) & (g506) & (!g468) & (!g475)) + ((i_8_) & (g135) & (!g485) & (g506) & (!g468) & (g475)) + ((i_8_) & (g135) & (!g485) & (g506) & (g468) & (!g475)) + ((i_8_) & (g135) & (!g485) & (g506) & (g468) & (g475)) + ((i_8_) & (g135) & (g485) & (!g506) & (!g468) & (!g475)) + ((i_8_) & (g135) & (g485) & (!g506) & (!g468) & (g475)) + ((i_8_) & (g135) & (g485) & (!g506) & (g468) & (!g475)) + ((i_8_) & (g135) & (g485) & (!g506) & (g468) & (g475)) + ((i_8_) & (g135) & (g485) & (g506) & (!g468) & (!g475)) + ((i_8_) & (g135) & (g485) & (g506) & (!g468) & (g475)) + ((i_8_) & (g135) & (g485) & (g506) & (g468) & (!g475)) + ((i_8_) & (g135) & (g485) & (g506) & (g468) & (g475)));
	assign g516 = (((!g100) & (!g506) & (!sk[22]) & (!g513) & (!g514) & (g515)) + ((!g100) & (!g506) & (!sk[22]) & (!g513) & (g514) & (g515)) + ((!g100) & (!g506) & (!sk[22]) & (g513) & (!g514) & (g515)) + ((!g100) & (!g506) & (!sk[22]) & (g513) & (g514) & (g515)) + ((!g100) & (!g506) & (sk[22]) & (!g513) & (!g514) & (!g515)) + ((!g100) & (g506) & (!sk[22]) & (!g513) & (!g514) & (g515)) + ((!g100) & (g506) & (!sk[22]) & (!g513) & (g514) & (g515)) + ((!g100) & (g506) & (!sk[22]) & (g513) & (!g514) & (g515)) + ((!g100) & (g506) & (!sk[22]) & (g513) & (g514) & (g515)) + ((!g100) & (g506) & (sk[22]) & (!g513) & (!g514) & (!g515)) + ((g100) & (!g506) & (!sk[22]) & (!g513) & (!g514) & (!g515)) + ((g100) & (!g506) & (!sk[22]) & (!g513) & (!g514) & (g515)) + ((g100) & (!g506) & (!sk[22]) & (!g513) & (g514) & (!g515)) + ((g100) & (!g506) & (!sk[22]) & (!g513) & (g514) & (g515)) + ((g100) & (!g506) & (!sk[22]) & (g513) & (!g514) & (!g515)) + ((g100) & (!g506) & (!sk[22]) & (g513) & (!g514) & (g515)) + ((g100) & (!g506) & (!sk[22]) & (g513) & (g514) & (!g515)) + ((g100) & (!g506) & (!sk[22]) & (g513) & (g514) & (g515)) + ((g100) & (!g506) & (sk[22]) & (!g513) & (!g514) & (!g515)) + ((g100) & (g506) & (!sk[22]) & (!g513) & (!g514) & (!g515)) + ((g100) & (g506) & (!sk[22]) & (!g513) & (!g514) & (g515)) + ((g100) & (g506) & (!sk[22]) & (!g513) & (g514) & (!g515)) + ((g100) & (g506) & (!sk[22]) & (!g513) & (g514) & (g515)) + ((g100) & (g506) & (!sk[22]) & (g513) & (!g514) & (!g515)) + ((g100) & (g506) & (!sk[22]) & (g513) & (!g514) & (g515)) + ((g100) & (g506) & (!sk[22]) & (g513) & (g514) & (!g515)) + ((g100) & (g506) & (!sk[22]) & (g513) & (g514) & (g515)));
	assign g517 = (((!g464) & (!g467) & (!sk[23]) & (!g474) & (!g465) & (g485)) + ((!g464) & (!g467) & (!sk[23]) & (!g474) & (g465) & (g485)) + ((!g464) & (!g467) & (!sk[23]) & (g474) & (!g465) & (g485)) + ((!g464) & (!g467) & (!sk[23]) & (g474) & (g465) & (g485)) + ((!g464) & (g467) & (!sk[23]) & (!g474) & (!g465) & (g485)) + ((!g464) & (g467) & (!sk[23]) & (!g474) & (g465) & (g485)) + ((!g464) & (g467) & (!sk[23]) & (g474) & (!g465) & (g485)) + ((!g464) & (g467) & (!sk[23]) & (g474) & (g465) & (g485)) + ((g464) & (!g467) & (!sk[23]) & (!g474) & (!g465) & (!g485)) + ((g464) & (!g467) & (!sk[23]) & (!g474) & (!g465) & (g485)) + ((g464) & (!g467) & (!sk[23]) & (!g474) & (g465) & (!g485)) + ((g464) & (!g467) & (!sk[23]) & (!g474) & (g465) & (g485)) + ((g464) & (!g467) & (!sk[23]) & (g474) & (!g465) & (!g485)) + ((g464) & (!g467) & (!sk[23]) & (g474) & (!g465) & (g485)) + ((g464) & (!g467) & (!sk[23]) & (g474) & (g465) & (!g485)) + ((g464) & (!g467) & (!sk[23]) & (g474) & (g465) & (g485)) + ((g464) & (g467) & (!sk[23]) & (!g474) & (!g465) & (!g485)) + ((g464) & (g467) & (!sk[23]) & (!g474) & (!g465) & (g485)) + ((g464) & (g467) & (!sk[23]) & (!g474) & (g465) & (!g485)) + ((g464) & (g467) & (!sk[23]) & (!g474) & (g465) & (g485)) + ((g464) & (g467) & (!sk[23]) & (g474) & (!g465) & (!g485)) + ((g464) & (g467) & (!sk[23]) & (g474) & (!g465) & (g485)) + ((g464) & (g467) & (!sk[23]) & (g474) & (g465) & (!g485)) + ((g464) & (g467) & (!sk[23]) & (g474) & (g465) & (g485)) + ((g464) & (g467) & (sk[23]) & (!g474) & (g465) & (!g485)));
	assign g518 = (((!i_11_) & (!sk[24]) & (!i_10_) & (i_15_) & (g461)) + ((!i_11_) & (!sk[24]) & (i_10_) & (!i_15_) & (!g461)) + ((!i_11_) & (!sk[24]) & (i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (!sk[24]) & (i_10_) & (i_15_) & (!g461)) + ((!i_11_) & (!sk[24]) & (i_10_) & (i_15_) & (g461)) + ((i_11_) & (!sk[24]) & (!i_10_) & (i_15_) & (!g461)) + ((i_11_) & (!sk[24]) & (!i_10_) & (i_15_) & (g461)) + ((i_11_) & (!sk[24]) & (i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (!sk[24]) & (i_10_) & (!i_15_) & (g461)) + ((i_11_) & (!sk[24]) & (i_10_) & (i_15_) & (!g461)) + ((i_11_) & (!sk[24]) & (i_10_) & (i_15_) & (g461)) + ((i_11_) & (sk[24]) & (!i_10_) & (i_15_) & (g461)));
	assign g519 = (((!g134) & (!g145) & (!g151) & (!g470) & (!g517) & (!g518)) + ((!g134) & (!g145) & (!g151) & (!g470) & (!g517) & (g518)) + ((!g134) & (!g145) & (!g151) & (!g470) & (g517) & (!g518)) + ((!g134) & (!g145) & (!g151) & (!g470) & (g517) & (g518)) + ((!g134) & (!g145) & (!g151) & (g470) & (!g517) & (!g518)) + ((!g134) & (!g145) & (!g151) & (g470) & (!g517) & (g518)) + ((!g134) & (!g145) & (!g151) & (g470) & (g517) & (!g518)) + ((!g134) & (!g145) & (!g151) & (g470) & (g517) & (g518)) + ((!g134) & (!g145) & (g151) & (!g470) & (!g517) & (!g518)) + ((!g134) & (!g145) & (g151) & (!g470) & (g517) & (!g518)) + ((!g134) & (!g145) & (g151) & (g470) & (!g517) & (!g518)) + ((!g134) & (!g145) & (g151) & (g470) & (g517) & (!g518)) + ((!g134) & (g145) & (!g151) & (!g470) & (!g517) & (!g518)) + ((!g134) & (g145) & (!g151) & (!g470) & (!g517) & (g518)) + ((!g134) & (g145) & (!g151) & (!g470) & (g517) & (!g518)) + ((!g134) & (g145) & (!g151) & (!g470) & (g517) & (g518)) + ((!g134) & (g145) & (g151) & (!g470) & (!g517) & (!g518)) + ((!g134) & (g145) & (g151) & (!g470) & (g517) & (!g518)) + ((g134) & (!g145) & (!g151) & (!g470) & (g517) & (!g518)) + ((g134) & (!g145) & (!g151) & (!g470) & (g517) & (g518)) + ((g134) & (!g145) & (g151) & (!g470) & (g517) & (!g518)) + ((g134) & (g145) & (!g151) & (!g470) & (g517) & (!g518)) + ((g134) & (g145) & (!g151) & (!g470) & (g517) & (g518)) + ((g134) & (g145) & (g151) & (!g470) & (g517) & (!g518)));
	assign g520 = (((!g109) & (!sk[26]) & (!g460) & (g516) & (g519)) + ((!g109) & (!sk[26]) & (g460) & (!g516) & (!g519)) + ((!g109) & (!sk[26]) & (g460) & (!g516) & (g519)) + ((!g109) & (!sk[26]) & (g460) & (g516) & (!g519)) + ((!g109) & (!sk[26]) & (g460) & (g516) & (g519)) + ((!g109) & (sk[26]) & (!g460) & (g516) & (g519)) + ((!g109) & (sk[26]) & (g460) & (g516) & (g519)) + ((g109) & (!sk[26]) & (!g460) & (g516) & (!g519)) + ((g109) & (!sk[26]) & (!g460) & (g516) & (g519)) + ((g109) & (!sk[26]) & (g460) & (!g516) & (!g519)) + ((g109) & (!sk[26]) & (g460) & (!g516) & (g519)) + ((g109) & (!sk[26]) & (g460) & (g516) & (!g519)) + ((g109) & (!sk[26]) & (g460) & (g516) & (g519)) + ((g109) & (sk[26]) & (!g460) & (g516) & (g519)));
	assign g521 = (((g490) & (g1737) & (g499) & (g1728) & (g512) & (g520)));
	assign g522 = (((!sk[28]) & (g93) & (!g171)) + ((!sk[28]) & (g93) & (g171)) + ((sk[28]) & (!g93) & (!g171)));
	assign g523 = (((!sk[29]) & (!g100) & (!g212) & (g251) & (g522)) + ((!sk[29]) & (!g100) & (g212) & (!g251) & (!g522)) + ((!sk[29]) & (!g100) & (g212) & (!g251) & (g522)) + ((!sk[29]) & (!g100) & (g212) & (g251) & (!g522)) + ((!sk[29]) & (!g100) & (g212) & (g251) & (g522)) + ((!sk[29]) & (g100) & (!g212) & (g251) & (!g522)) + ((!sk[29]) & (g100) & (!g212) & (g251) & (g522)) + ((!sk[29]) & (g100) & (g212) & (!g251) & (!g522)) + ((!sk[29]) & (g100) & (g212) & (!g251) & (g522)) + ((!sk[29]) & (g100) & (g212) & (g251) & (!g522)) + ((!sk[29]) & (g100) & (g212) & (g251) & (g522)) + ((sk[29]) & (!g100) & (!g212) & (!g251) & (g522)) + ((sk[29]) & (!g100) & (!g212) & (g251) & (g522)) + ((sk[29]) & (!g100) & (g212) & (g251) & (g522)) + ((sk[29]) & (g100) & (!g212) & (!g251) & (g522)) + ((sk[29]) & (g100) & (!g212) & (g251) & (g522)) + ((sk[29]) & (g100) & (g212) & (!g251) & (g522)) + ((sk[29]) & (g100) & (g212) & (g251) & (g522)));
	assign g524 = (((!i_11_) & (!sk[30]) & (!i_9_) & (i_15_) & (g375)) + ((!i_11_) & (!sk[30]) & (i_9_) & (!i_15_) & (!g375)) + ((!i_11_) & (!sk[30]) & (i_9_) & (!i_15_) & (g375)) + ((!i_11_) & (!sk[30]) & (i_9_) & (i_15_) & (!g375)) + ((!i_11_) & (!sk[30]) & (i_9_) & (i_15_) & (g375)) + ((i_11_) & (!sk[30]) & (!i_9_) & (i_15_) & (!g375)) + ((i_11_) & (!sk[30]) & (!i_9_) & (i_15_) & (g375)) + ((i_11_) & (!sk[30]) & (i_9_) & (!i_15_) & (!g375)) + ((i_11_) & (!sk[30]) & (i_9_) & (!i_15_) & (g375)) + ((i_11_) & (!sk[30]) & (i_9_) & (i_15_) & (!g375)) + ((i_11_) & (!sk[30]) & (i_9_) & (i_15_) & (g375)) + ((i_11_) & (sk[30]) & (!i_9_) & (i_15_) & (g375)));
	assign g525 = (((!i_11_) & (!i_9_) & (!g326) & (!g98) & (!sk[31]) & (g111)) + ((!i_11_) & (!i_9_) & (!g326) & (g98) & (!sk[31]) & (g111)) + ((!i_11_) & (!i_9_) & (g326) & (!g98) & (!sk[31]) & (g111)) + ((!i_11_) & (!i_9_) & (g326) & (g98) & (!sk[31]) & (g111)) + ((!i_11_) & (i_9_) & (!g326) & (!g98) & (!sk[31]) & (g111)) + ((!i_11_) & (i_9_) & (!g326) & (g98) & (!sk[31]) & (g111)) + ((!i_11_) & (i_9_) & (g326) & (!g98) & (!sk[31]) & (g111)) + ((!i_11_) & (i_9_) & (g326) & (g98) & (!sk[31]) & (g111)) + ((i_11_) & (!i_9_) & (!g326) & (!g98) & (!sk[31]) & (!g111)) + ((i_11_) & (!i_9_) & (!g326) & (!g98) & (!sk[31]) & (g111)) + ((i_11_) & (!i_9_) & (!g326) & (g98) & (!sk[31]) & (!g111)) + ((i_11_) & (!i_9_) & (!g326) & (g98) & (!sk[31]) & (g111)) + ((i_11_) & (!i_9_) & (g326) & (!g98) & (!sk[31]) & (!g111)) + ((i_11_) & (!i_9_) & (g326) & (!g98) & (!sk[31]) & (g111)) + ((i_11_) & (!i_9_) & (g326) & (g98) & (!sk[31]) & (!g111)) + ((i_11_) & (!i_9_) & (g326) & (g98) & (!sk[31]) & (g111)) + ((i_11_) & (!i_9_) & (g326) & (g98) & (sk[31]) & (g111)) + ((i_11_) & (i_9_) & (!g326) & (!g98) & (!sk[31]) & (!g111)) + ((i_11_) & (i_9_) & (!g326) & (!g98) & (!sk[31]) & (g111)) + ((i_11_) & (i_9_) & (!g326) & (g98) & (!sk[31]) & (!g111)) + ((i_11_) & (i_9_) & (!g326) & (g98) & (!sk[31]) & (g111)) + ((i_11_) & (i_9_) & (g326) & (!g98) & (!sk[31]) & (!g111)) + ((i_11_) & (i_9_) & (g326) & (!g98) & (!sk[31]) & (g111)) + ((i_11_) & (i_9_) & (g326) & (g98) & (!sk[31]) & (!g111)) + ((i_11_) & (i_9_) & (g326) & (g98) & (!sk[31]) & (g111)));
	assign g526 = (((!g297) & (!g216) & (!g227) & (!g231) & (!g238) & (!g349)) + ((!g297) & (!g216) & (!g227) & (!g231) & (!g238) & (g349)) + ((!g297) & (!g216) & (!g227) & (!g231) & (g238) & (!g349)) + ((!g297) & (!g216) & (!g227) & (!g231) & (g238) & (g349)) + ((!g297) & (!g216) & (!g227) & (g231) & (!g238) & (!g349)) + ((!g297) & (!g216) & (!g227) & (g231) & (!g238) & (g349)) + ((!g297) & (!g216) & (!g227) & (g231) & (g238) & (!g349)) + ((!g297) & (!g216) & (!g227) & (g231) & (g238) & (g349)) + ((!g297) & (!g216) & (g227) & (g231) & (!g238) & (!g349)) + ((!g297) & (!g216) & (g227) & (g231) & (g238) & (!g349)) + ((!g297) & (g216) & (!g227) & (!g231) & (!g238) & (!g349)) + ((!g297) & (g216) & (!g227) & (!g231) & (!g238) & (g349)) + ((!g297) & (g216) & (!g227) & (g231) & (!g238) & (!g349)) + ((!g297) & (g216) & (!g227) & (g231) & (!g238) & (g349)) + ((!g297) & (g216) & (g227) & (g231) & (!g238) & (!g349)) + ((g297) & (!g216) & (!g227) & (!g231) & (!g238) & (!g349)) + ((g297) & (!g216) & (!g227) & (!g231) & (!g238) & (g349)) + ((g297) & (!g216) & (!g227) & (g231) & (!g238) & (!g349)) + ((g297) & (!g216) & (!g227) & (g231) & (!g238) & (g349)) + ((g297) & (!g216) & (g227) & (g231) & (!g238) & (!g349)) + ((g297) & (g216) & (!g227) & (!g231) & (!g238) & (!g349)) + ((g297) & (g216) & (!g227) & (!g231) & (!g238) & (g349)) + ((g297) & (g216) & (!g227) & (g231) & (!g238) & (!g349)) + ((g297) & (g216) & (!g227) & (g231) & (!g238) & (g349)) + ((g297) & (g216) & (g227) & (g231) & (!g238) & (!g349)));
	assign g527 = (((!g261) & (!sk[33]) & (!g523) & (!g524) & (!g525) & (g526)) + ((!g261) & (!sk[33]) & (!g523) & (!g524) & (g525) & (g526)) + ((!g261) & (!sk[33]) & (!g523) & (g524) & (!g525) & (g526)) + ((!g261) & (!sk[33]) & (!g523) & (g524) & (g525) & (g526)) + ((!g261) & (!sk[33]) & (g523) & (!g524) & (!g525) & (g526)) + ((!g261) & (!sk[33]) & (g523) & (!g524) & (g525) & (g526)) + ((!g261) & (!sk[33]) & (g523) & (g524) & (!g525) & (g526)) + ((!g261) & (!sk[33]) & (g523) & (g524) & (g525) & (g526)) + ((!g261) & (sk[33]) & (!g523) & (!g524) & (!g525) & (g526)) + ((g261) & (!sk[33]) & (!g523) & (!g524) & (!g525) & (!g526)) + ((g261) & (!sk[33]) & (!g523) & (!g524) & (!g525) & (g526)) + ((g261) & (!sk[33]) & (!g523) & (!g524) & (g525) & (!g526)) + ((g261) & (!sk[33]) & (!g523) & (!g524) & (g525) & (g526)) + ((g261) & (!sk[33]) & (!g523) & (g524) & (!g525) & (!g526)) + ((g261) & (!sk[33]) & (!g523) & (g524) & (!g525) & (g526)) + ((g261) & (!sk[33]) & (!g523) & (g524) & (g525) & (!g526)) + ((g261) & (!sk[33]) & (!g523) & (g524) & (g525) & (g526)) + ((g261) & (!sk[33]) & (g523) & (!g524) & (!g525) & (!g526)) + ((g261) & (!sk[33]) & (g523) & (!g524) & (!g525) & (g526)) + ((g261) & (!sk[33]) & (g523) & (!g524) & (g525) & (!g526)) + ((g261) & (!sk[33]) & (g523) & (!g524) & (g525) & (g526)) + ((g261) & (!sk[33]) & (g523) & (g524) & (!g525) & (!g526)) + ((g261) & (!sk[33]) & (g523) & (g524) & (!g525) & (g526)) + ((g261) & (!sk[33]) & (g523) & (g524) & (g525) & (!g526)) + ((g261) & (!sk[33]) & (g523) & (g524) & (g525) & (g526)));
	assign g528 = (((!sk[34]) & (g45) & (!g197)) + ((!sk[34]) & (g45) & (g197)) + ((sk[34]) & (!g45) & (!g197)));
	assign g529 = (((!sk[35]) & (g467) & (!g528)) + ((!sk[35]) & (g467) & (g528)) + ((sk[35]) & (g467) & (g528)));
	assign g530 = (((!sk[36]) & (g22) & (!g171)) + ((!sk[36]) & (g22) & (g171)) + ((sk[36]) & (g22) & (!g171)));
	assign g531 = (((!sk[37]) & (g6) & (!i_15_) & (!g171)) + ((!sk[37]) & (g6) & (!i_15_) & (g171)) + ((!sk[37]) & (g6) & (i_15_) & (!g171)) + ((!sk[37]) & (g6) & (i_15_) & (g171)) + ((sk[37]) & (g6) & (i_15_) & (!g171)));
	assign g532 = (((!sk[38]) & (g13) & (!g124)) + ((!sk[38]) & (g13) & (g124)) + ((sk[38]) & (g13) & (g124)));
	assign g533 = (((!g134) & (!g195) & (g532) & (!sk[39]) & (g478)) + ((!g134) & (g195) & (!g532) & (!sk[39]) & (!g478)) + ((!g134) & (g195) & (!g532) & (!sk[39]) & (g478)) + ((!g134) & (g195) & (g532) & (!sk[39]) & (!g478)) + ((!g134) & (g195) & (g532) & (!sk[39]) & (g478)) + ((g134) & (!g195) & (!g532) & (sk[39]) & (g478)) + ((g134) & (!g195) & (g532) & (!sk[39]) & (!g478)) + ((g134) & (!g195) & (g532) & (!sk[39]) & (g478)) + ((g134) & (!g195) & (g532) & (sk[39]) & (!g478)) + ((g134) & (!g195) & (g532) & (sk[39]) & (g478)) + ((g134) & (g195) & (!g532) & (!sk[39]) & (!g478)) + ((g134) & (g195) & (!g532) & (!sk[39]) & (g478)) + ((g134) & (g195) & (!g532) & (sk[39]) & (!g478)) + ((g134) & (g195) & (!g532) & (sk[39]) & (g478)) + ((g134) & (g195) & (g532) & (!sk[39]) & (!g478)) + ((g134) & (g195) & (g532) & (!sk[39]) & (g478)) + ((g134) & (g195) & (g532) & (sk[39]) & (!g478)) + ((g134) & (g195) & (g532) & (sk[39]) & (g478)));
	assign g534 = (((!g171) & (sk[40]) & (g124)) + ((g171) & (!sk[40]) & (!g124)) + ((g171) & (!sk[40]) & (g124)));
	assign g535 = (((!sk[41]) & (g45) & (!g224) & (!g467)) + ((!sk[41]) & (g45) & (!g224) & (g467)) + ((!sk[41]) & (g45) & (g224) & (!g467)) + ((!sk[41]) & (g45) & (g224) & (g467)) + ((sk[41]) & (!g45) & (!g224) & (g467)));
	assign g536 = (((!g99) & (!sk[42]) & (!g534) & (!g530) & (!g531) & (g535)) + ((!g99) & (!sk[42]) & (!g534) & (!g530) & (g531) & (g535)) + ((!g99) & (!sk[42]) & (!g534) & (g530) & (!g531) & (g535)) + ((!g99) & (!sk[42]) & (!g534) & (g530) & (g531) & (g535)) + ((!g99) & (!sk[42]) & (g534) & (!g530) & (!g531) & (g535)) + ((!g99) & (!sk[42]) & (g534) & (!g530) & (g531) & (g535)) + ((!g99) & (!sk[42]) & (g534) & (g530) & (!g531) & (g535)) + ((!g99) & (!sk[42]) & (g534) & (g530) & (g531) & (g535)) + ((g99) & (!sk[42]) & (!g534) & (!g530) & (!g531) & (!g535)) + ((g99) & (!sk[42]) & (!g534) & (!g530) & (!g531) & (g535)) + ((g99) & (!sk[42]) & (!g534) & (!g530) & (g531) & (!g535)) + ((g99) & (!sk[42]) & (!g534) & (!g530) & (g531) & (g535)) + ((g99) & (!sk[42]) & (!g534) & (g530) & (!g531) & (!g535)) + ((g99) & (!sk[42]) & (!g534) & (g530) & (!g531) & (g535)) + ((g99) & (!sk[42]) & (!g534) & (g530) & (g531) & (!g535)) + ((g99) & (!sk[42]) & (!g534) & (g530) & (g531) & (g535)) + ((g99) & (!sk[42]) & (g534) & (!g530) & (!g531) & (!g535)) + ((g99) & (!sk[42]) & (g534) & (!g530) & (!g531) & (g535)) + ((g99) & (!sk[42]) & (g534) & (!g530) & (g531) & (!g535)) + ((g99) & (!sk[42]) & (g534) & (!g530) & (g531) & (g535)) + ((g99) & (!sk[42]) & (g534) & (g530) & (!g531) & (!g535)) + ((g99) & (!sk[42]) & (g534) & (g530) & (!g531) & (g535)) + ((g99) & (!sk[42]) & (g534) & (g530) & (g531) & (!g535)) + ((g99) & (!sk[42]) & (g534) & (g530) & (g531) & (g535)) + ((g99) & (sk[42]) & (!g534) & (!g530) & (!g531) & (!g535)) + ((g99) & (sk[42]) & (!g534) & (!g530) & (g531) & (!g535)) + ((g99) & (sk[42]) & (!g534) & (!g530) & (g531) & (g535)) + ((g99) & (sk[42]) & (!g534) & (g530) & (!g531) & (!g535)) + ((g99) & (sk[42]) & (!g534) & (g530) & (!g531) & (g535)) + ((g99) & (sk[42]) & (!g534) & (g530) & (g531) & (!g535)) + ((g99) & (sk[42]) & (!g534) & (g530) & (g531) & (g535)) + ((g99) & (sk[42]) & (g534) & (!g530) & (!g531) & (!g535)) + ((g99) & (sk[42]) & (g534) & (!g530) & (!g531) & (g535)) + ((g99) & (sk[42]) & (g534) & (!g530) & (g531) & (!g535)) + ((g99) & (sk[42]) & (g534) & (!g530) & (g531) & (g535)) + ((g99) & (sk[42]) & (g534) & (g530) & (!g531) & (!g535)) + ((g99) & (sk[42]) & (g534) & (g530) & (!g531) & (g535)) + ((g99) & (sk[42]) & (g534) & (g530) & (g531) & (!g535)) + ((g99) & (sk[42]) & (g534) & (g530) & (g531) & (g535)));
	assign g537 = (((!g423) & (!g464) & (!g478) & (!g533) & (!sk[43]) & (g536)) + ((!g423) & (!g464) & (!g478) & (!g533) & (sk[43]) & (!g536)) + ((!g423) & (!g464) & (!g478) & (g533) & (!sk[43]) & (g536)) + ((!g423) & (!g464) & (g478) & (!g533) & (!sk[43]) & (g536)) + ((!g423) & (!g464) & (g478) & (!g533) & (sk[43]) & (!g536)) + ((!g423) & (!g464) & (g478) & (g533) & (!sk[43]) & (g536)) + ((!g423) & (g464) & (!g478) & (!g533) & (!sk[43]) & (g536)) + ((!g423) & (g464) & (!g478) & (!g533) & (sk[43]) & (!g536)) + ((!g423) & (g464) & (!g478) & (g533) & (!sk[43]) & (g536)) + ((!g423) & (g464) & (g478) & (!g533) & (!sk[43]) & (g536)) + ((!g423) & (g464) & (g478) & (!g533) & (sk[43]) & (!g536)) + ((!g423) & (g464) & (g478) & (g533) & (!sk[43]) & (g536)) + ((g423) & (!g464) & (!g478) & (!g533) & (!sk[43]) & (!g536)) + ((g423) & (!g464) & (!g478) & (!g533) & (!sk[43]) & (g536)) + ((g423) & (!g464) & (!g478) & (g533) & (!sk[43]) & (!g536)) + ((g423) & (!g464) & (!g478) & (g533) & (!sk[43]) & (g536)) + ((g423) & (!g464) & (g478) & (!g533) & (!sk[43]) & (!g536)) + ((g423) & (!g464) & (g478) & (!g533) & (!sk[43]) & (g536)) + ((g423) & (!g464) & (g478) & (g533) & (!sk[43]) & (!g536)) + ((g423) & (!g464) & (g478) & (g533) & (!sk[43]) & (g536)) + ((g423) & (g464) & (!g478) & (!g533) & (!sk[43]) & (!g536)) + ((g423) & (g464) & (!g478) & (!g533) & (!sk[43]) & (g536)) + ((g423) & (g464) & (!g478) & (!g533) & (sk[43]) & (!g536)) + ((g423) & (g464) & (!g478) & (g533) & (!sk[43]) & (!g536)) + ((g423) & (g464) & (!g478) & (g533) & (!sk[43]) & (g536)) + ((g423) & (g464) & (g478) & (!g533) & (!sk[43]) & (!g536)) + ((g423) & (g464) & (g478) & (!g533) & (!sk[43]) & (g536)) + ((g423) & (g464) & (g478) & (g533) & (!sk[43]) & (!g536)) + ((g423) & (g464) & (g478) & (g533) & (!sk[43]) & (g536)));
	assign g538 = (((!sk[44]) & (!i_8_) & (!i_6_) & (!i_7_) & (!g98) & (g87)) + ((!sk[44]) & (!i_8_) & (!i_6_) & (!i_7_) & (g98) & (g87)) + ((!sk[44]) & (!i_8_) & (!i_6_) & (i_7_) & (!g98) & (g87)) + ((!sk[44]) & (!i_8_) & (!i_6_) & (i_7_) & (g98) & (g87)) + ((!sk[44]) & (!i_8_) & (i_6_) & (!i_7_) & (!g98) & (g87)) + ((!sk[44]) & (!i_8_) & (i_6_) & (!i_7_) & (g98) & (g87)) + ((!sk[44]) & (!i_8_) & (i_6_) & (i_7_) & (!g98) & (g87)) + ((!sk[44]) & (!i_8_) & (i_6_) & (i_7_) & (g98) & (g87)) + ((!sk[44]) & (i_8_) & (!i_6_) & (!i_7_) & (!g98) & (!g87)) + ((!sk[44]) & (i_8_) & (!i_6_) & (!i_7_) & (!g98) & (g87)) + ((!sk[44]) & (i_8_) & (!i_6_) & (!i_7_) & (g98) & (!g87)) + ((!sk[44]) & (i_8_) & (!i_6_) & (!i_7_) & (g98) & (g87)) + ((!sk[44]) & (i_8_) & (!i_6_) & (i_7_) & (!g98) & (!g87)) + ((!sk[44]) & (i_8_) & (!i_6_) & (i_7_) & (!g98) & (g87)) + ((!sk[44]) & (i_8_) & (!i_6_) & (i_7_) & (g98) & (!g87)) + ((!sk[44]) & (i_8_) & (!i_6_) & (i_7_) & (g98) & (g87)) + ((!sk[44]) & (i_8_) & (i_6_) & (!i_7_) & (!g98) & (!g87)) + ((!sk[44]) & (i_8_) & (i_6_) & (!i_7_) & (!g98) & (g87)) + ((!sk[44]) & (i_8_) & (i_6_) & (!i_7_) & (g98) & (!g87)) + ((!sk[44]) & (i_8_) & (i_6_) & (!i_7_) & (g98) & (g87)) + ((!sk[44]) & (i_8_) & (i_6_) & (i_7_) & (!g98) & (!g87)) + ((!sk[44]) & (i_8_) & (i_6_) & (i_7_) & (!g98) & (g87)) + ((!sk[44]) & (i_8_) & (i_6_) & (i_7_) & (g98) & (!g87)) + ((!sk[44]) & (i_8_) & (i_6_) & (i_7_) & (g98) & (g87)) + ((sk[44]) & (!i_8_) & (!i_6_) & (!i_7_) & (!g98) & (g87)) + ((sk[44]) & (!i_8_) & (!i_6_) & (!i_7_) & (g98) & (g87)) + ((sk[44]) & (!i_8_) & (!i_6_) & (i_7_) & (!g98) & (g87)) + ((sk[44]) & (!i_8_) & (!i_6_) & (i_7_) & (g98) & (!g87)) + ((sk[44]) & (!i_8_) & (!i_6_) & (i_7_) & (g98) & (g87)) + ((sk[44]) & (!i_8_) & (i_6_) & (!i_7_) & (g98) & (!g87)) + ((sk[44]) & (!i_8_) & (i_6_) & (!i_7_) & (g98) & (g87)) + ((sk[44]) & (!i_8_) & (i_6_) & (i_7_) & (g98) & (!g87)) + ((sk[44]) & (!i_8_) & (i_6_) & (i_7_) & (g98) & (g87)) + ((sk[44]) & (i_8_) & (!i_6_) & (i_7_) & (!g98) & (g87)) + ((sk[44]) & (i_8_) & (!i_6_) & (i_7_) & (g98) & (!g87)) + ((sk[44]) & (i_8_) & (!i_6_) & (i_7_) & (g98) & (g87)));
	assign g539 = (((!g99) & (!g251) & (g277) & (!g158) & (!g285) & (!g538)) + ((!g99) & (!g251) & (g277) & (!g158) & (g285) & (!g538)) + ((!g99) & (!g251) & (g277) & (g158) & (g285) & (!g538)) + ((!g99) & (g251) & (g277) & (!g158) & (!g285) & (!g538)) + ((!g99) & (g251) & (g277) & (!g158) & (g285) & (!g538)) + ((g99) & (!g251) & (g277) & (!g158) & (!g285) & (!g538)) + ((g99) & (!g251) & (g277) & (!g158) & (g285) & (!g538)) + ((g99) & (g251) & (g277) & (!g158) & (!g285) & (!g538)) + ((g99) & (g251) & (g277) & (!g158) & (g285) & (!g538)));
	assign g540 = (((!g171) & (sk[46]) & (!g122)) + ((g171) & (!sk[46]) & (!g122)) + ((g171) & (!sk[46]) & (g122)));
	assign g541 = (((!sk[47]) & (!i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (g171)) + ((!sk[47]) & (!i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (g171)) + ((!sk[47]) & (!i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (g171)) + ((!sk[47]) & (!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g171)) + ((!sk[47]) & (!i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (g171)) + ((!sk[47]) & (!i_11_) & (i_9_) & (!i_10_) & (i_15_) & (g171)) + ((!sk[47]) & (!i_11_) & (i_9_) & (i_10_) & (!i_15_) & (g171)) + ((!sk[47]) & (!i_11_) & (i_9_) & (i_10_) & (i_15_) & (g171)) + ((!sk[47]) & (i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (!g171)) + ((!sk[47]) & (i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (g171)) + ((!sk[47]) & (i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (!g171)) + ((!sk[47]) & (i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (g171)) + ((!sk[47]) & (i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (!g171)) + ((!sk[47]) & (i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (g171)) + ((!sk[47]) & (i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!g171)) + ((!sk[47]) & (i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g171)) + ((!sk[47]) & (i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (!g171)) + ((!sk[47]) & (i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (g171)) + ((!sk[47]) & (i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!g171)) + ((!sk[47]) & (i_11_) & (i_9_) & (!i_10_) & (i_15_) & (g171)) + ((!sk[47]) & (i_11_) & (i_9_) & (i_10_) & (!i_15_) & (!g171)) + ((!sk[47]) & (i_11_) & (i_9_) & (i_10_) & (!i_15_) & (g171)) + ((!sk[47]) & (i_11_) & (i_9_) & (i_10_) & (i_15_) & (!g171)) + ((!sk[47]) & (i_11_) & (i_9_) & (i_10_) & (i_15_) & (g171)) + ((sk[47]) & (!i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (!g171)) + ((sk[47]) & (i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!g171)));
	assign g542 = (((!g99) & (!g251) & (!g285) & (!g540) & (!sk[48]) & (g541)) + ((!g99) & (!g251) & (!g285) & (!g540) & (sk[48]) & (g541)) + ((!g99) & (!g251) & (!g285) & (g540) & (!sk[48]) & (g541)) + ((!g99) & (!g251) & (!g285) & (g540) & (sk[48]) & (g541)) + ((!g99) & (!g251) & (g285) & (!g540) & (!sk[48]) & (g541)) + ((!g99) & (!g251) & (g285) & (g540) & (!sk[48]) & (g541)) + ((!g99) & (!g251) & (g285) & (g540) & (sk[48]) & (g541)) + ((!g99) & (g251) & (!g285) & (!g540) & (!sk[48]) & (g541)) + ((!g99) & (g251) & (!g285) & (!g540) & (sk[48]) & (g541)) + ((!g99) & (g251) & (!g285) & (g540) & (!sk[48]) & (g541)) + ((!g99) & (g251) & (!g285) & (g540) & (sk[48]) & (g541)) + ((!g99) & (g251) & (g285) & (!g540) & (!sk[48]) & (g541)) + ((!g99) & (g251) & (g285) & (!g540) & (sk[48]) & (g541)) + ((!g99) & (g251) & (g285) & (g540) & (!sk[48]) & (g541)) + ((!g99) & (g251) & (g285) & (g540) & (sk[48]) & (g541)) + ((g99) & (!g251) & (!g285) & (!g540) & (!sk[48]) & (!g541)) + ((g99) & (!g251) & (!g285) & (!g540) & (!sk[48]) & (g541)) + ((g99) & (!g251) & (!g285) & (!g540) & (sk[48]) & (g541)) + ((g99) & (!g251) & (!g285) & (g540) & (!sk[48]) & (!g541)) + ((g99) & (!g251) & (!g285) & (g540) & (!sk[48]) & (g541)) + ((g99) & (!g251) & (!g285) & (g540) & (sk[48]) & (g541)) + ((g99) & (!g251) & (g285) & (!g540) & (!sk[48]) & (!g541)) + ((g99) & (!g251) & (g285) & (!g540) & (!sk[48]) & (g541)) + ((g99) & (!g251) & (g285) & (!g540) & (sk[48]) & (g541)) + ((g99) & (!g251) & (g285) & (g540) & (!sk[48]) & (!g541)) + ((g99) & (!g251) & (g285) & (g540) & (!sk[48]) & (g541)) + ((g99) & (!g251) & (g285) & (g540) & (sk[48]) & (g541)) + ((g99) & (g251) & (!g285) & (!g540) & (!sk[48]) & (!g541)) + ((g99) & (g251) & (!g285) & (!g540) & (!sk[48]) & (g541)) + ((g99) & (g251) & (!g285) & (!g540) & (sk[48]) & (g541)) + ((g99) & (g251) & (!g285) & (g540) & (!sk[48]) & (!g541)) + ((g99) & (g251) & (!g285) & (g540) & (!sk[48]) & (g541)) + ((g99) & (g251) & (!g285) & (g540) & (sk[48]) & (g541)) + ((g99) & (g251) & (g285) & (!g540) & (!sk[48]) & (!g541)) + ((g99) & (g251) & (g285) & (!g540) & (!sk[48]) & (g541)) + ((g99) & (g251) & (g285) & (!g540) & (sk[48]) & (g541)) + ((g99) & (g251) & (g285) & (g540) & (!sk[48]) & (!g541)) + ((g99) & (g251) & (g285) & (g540) & (!sk[48]) & (g541)) + ((g99) & (g251) & (g285) & (g540) & (sk[48]) & (g541)));
	assign g543 = (((!g109) & (!g529) & (g1721) & (g537) & (!g539) & (!g542)) + ((!g109) & (!g529) & (g1721) & (g537) & (g539) & (!g542)) + ((!g109) & (!g529) & (g1721) & (g537) & (g539) & (g542)) + ((!g109) & (g529) & (g1721) & (g537) & (!g539) & (!g542)) + ((!g109) & (g529) & (g1721) & (g537) & (g539) & (!g542)) + ((!g109) & (g529) & (g1721) & (g537) & (g539) & (g542)) + ((g109) & (g529) & (g1721) & (g537) & (!g539) & (!g542)) + ((g109) & (g529) & (g1721) & (g537) & (g539) & (!g542)) + ((g109) & (g529) & (g1721) & (g537) & (g539) & (g542)));
	assign g544 = (((!sk[50]) & (g6) & (!i_15_) & (!g461)) + ((!sk[50]) & (g6) & (!i_15_) & (g461)) + ((!sk[50]) & (g6) & (i_15_) & (!g461)) + ((!sk[50]) & (g6) & (i_15_) & (g461)) + ((sk[50]) & (!g6) & (!i_15_) & (!g461)) + ((sk[50]) & (!g6) & (!i_15_) & (g461)) + ((sk[50]) & (!g6) & (i_15_) & (!g461)) + ((sk[50]) & (!g6) & (i_15_) & (g461)) + ((sk[50]) & (g6) & (!i_15_) & (!g461)) + ((sk[50]) & (g6) & (i_15_) & (!g461)) + ((sk[50]) & (g6) & (i_15_) & (g461)));
	assign g545 = (((!g45) & (sk[51]) & (g118) & (!g544)) + ((g45) & (!sk[51]) & (!g118) & (!g544)) + ((g45) & (!sk[51]) & (!g118) & (g544)) + ((g45) & (!sk[51]) & (g118) & (!g544)) + ((g45) & (!sk[51]) & (g118) & (g544)) + ((g45) & (sk[51]) & (g118) & (!g544)) + ((g45) & (sk[51]) & (g118) & (g544)));
	assign g546 = (((g13) & (!sk[52]) & (!g115)) + ((g13) & (!sk[52]) & (g115)) + ((g13) & (sk[52]) & (!g115)));
	assign g547 = (((!sk[53]) & (g13) & (!g122)) + ((!sk[53]) & (g13) & (g122)) + ((sk[53]) & (!g13) & (!g122)) + ((sk[53]) & (!g13) & (g122)) + ((sk[53]) & (g13) & (g122)));
	assign g548 = (((g119) & (!sk[54]) & (!g461)) + ((g119) & (!sk[54]) & (g461)) + ((g119) & (sk[54]) & (g461)));
	assign g549 = (((!sk[55]) & (g547) & (!g548)) + ((!sk[55]) & (g547) & (g548)) + ((sk[55]) & (g547) & (!g548)));
	assign g550 = (((!sk[56]) & (g102) & (!g461)) + ((!sk[56]) & (g102) & (g461)) + ((sk[56]) & (!g102) & (g461)));
	assign g551 = (((g104) & (!sk[57]) & (!g461)) + ((g104) & (!sk[57]) & (g461)) + ((g104) & (sk[57]) & (g461)));
	assign g552 = (((!i_8_) & (g108) & (!g135) & (g550) & (!g546) & (!g551)) + ((!i_8_) & (g108) & (!g135) & (g550) & (!g546) & (g551)) + ((!i_8_) & (g108) & (!g135) & (g550) & (g546) & (!g551)) + ((!i_8_) & (g108) & (!g135) & (g550) & (g546) & (g551)) + ((!i_8_) & (g108) & (g135) & (g550) & (!g546) & (!g551)) + ((!i_8_) & (g108) & (g135) & (g550) & (!g546) & (g551)) + ((!i_8_) & (g108) & (g135) & (g550) & (g546) & (!g551)) + ((!i_8_) & (g108) & (g135) & (g550) & (g546) & (g551)) + ((i_8_) & (!g108) & (g135) & (!g550) & (!g546) & (g551)) + ((i_8_) & (!g108) & (g135) & (!g550) & (g546) & (!g551)) + ((i_8_) & (!g108) & (g135) & (!g550) & (g546) & (g551)) + ((i_8_) & (!g108) & (g135) & (g550) & (!g546) & (!g551)) + ((i_8_) & (!g108) & (g135) & (g550) & (!g546) & (g551)) + ((i_8_) & (!g108) & (g135) & (g550) & (g546) & (!g551)) + ((i_8_) & (!g108) & (g135) & (g550) & (g546) & (g551)) + ((i_8_) & (g108) & (!g135) & (!g550) & (!g546) & (g551)) + ((i_8_) & (g108) & (!g135) & (!g550) & (g546) & (g551)) + ((i_8_) & (g108) & (!g135) & (g550) & (!g546) & (g551)) + ((i_8_) & (g108) & (!g135) & (g550) & (g546) & (g551)) + ((i_8_) & (g108) & (g135) & (!g550) & (!g546) & (g551)) + ((i_8_) & (g108) & (g135) & (!g550) & (g546) & (!g551)) + ((i_8_) & (g108) & (g135) & (!g550) & (g546) & (g551)) + ((i_8_) & (g108) & (g135) & (g550) & (!g546) & (!g551)) + ((i_8_) & (g108) & (g135) & (g550) & (!g546) & (g551)) + ((i_8_) & (g108) & (g135) & (g550) & (g546) & (!g551)) + ((i_8_) & (g108) & (g135) & (g550) & (g546) & (g551)));
	assign g553 = (((!g149) & (!sk[59]) & (!g151) & (!g549) & (!g532) & (g552)) + ((!g149) & (!sk[59]) & (!g151) & (!g549) & (g532) & (g552)) + ((!g149) & (!sk[59]) & (!g151) & (g549) & (!g532) & (g552)) + ((!g149) & (!sk[59]) & (!g151) & (g549) & (g532) & (g552)) + ((!g149) & (!sk[59]) & (g151) & (!g549) & (!g532) & (g552)) + ((!g149) & (!sk[59]) & (g151) & (!g549) & (g532) & (g552)) + ((!g149) & (!sk[59]) & (g151) & (g549) & (!g532) & (g552)) + ((!g149) & (!sk[59]) & (g151) & (g549) & (g532) & (g552)) + ((!g149) & (sk[59]) & (!g151) & (!g549) & (!g532) & (!g552)) + ((!g149) & (sk[59]) & (!g151) & (!g549) & (g532) & (!g552)) + ((!g149) & (sk[59]) & (!g151) & (g549) & (!g532) & (!g552)) + ((!g149) & (sk[59]) & (!g151) & (g549) & (g532) & (!g552)) + ((!g149) & (sk[59]) & (g151) & (!g549) & (!g532) & (!g552)) + ((!g149) & (sk[59]) & (g151) & (g549) & (!g532) & (!g552)) + ((g149) & (!sk[59]) & (!g151) & (!g549) & (!g532) & (!g552)) + ((g149) & (!sk[59]) & (!g151) & (!g549) & (!g532) & (g552)) + ((g149) & (!sk[59]) & (!g151) & (!g549) & (g532) & (!g552)) + ((g149) & (!sk[59]) & (!g151) & (!g549) & (g532) & (g552)) + ((g149) & (!sk[59]) & (!g151) & (g549) & (!g532) & (!g552)) + ((g149) & (!sk[59]) & (!g151) & (g549) & (!g532) & (g552)) + ((g149) & (!sk[59]) & (!g151) & (g549) & (g532) & (!g552)) + ((g149) & (!sk[59]) & (!g151) & (g549) & (g532) & (g552)) + ((g149) & (!sk[59]) & (g151) & (!g549) & (!g532) & (!g552)) + ((g149) & (!sk[59]) & (g151) & (!g549) & (!g532) & (g552)) + ((g149) & (!sk[59]) & (g151) & (!g549) & (g532) & (!g552)) + ((g149) & (!sk[59]) & (g151) & (!g549) & (g532) & (g552)) + ((g149) & (!sk[59]) & (g151) & (g549) & (!g532) & (!g552)) + ((g149) & (!sk[59]) & (g151) & (g549) & (!g532) & (g552)) + ((g149) & (!sk[59]) & (g151) & (g549) & (g532) & (!g552)) + ((g149) & (!sk[59]) & (g151) & (g549) & (g532) & (g552)) + ((g149) & (sk[59]) & (!g151) & (g549) & (!g532) & (!g552)) + ((g149) & (sk[59]) & (!g151) & (g549) & (g532) & (!g552)) + ((g149) & (sk[59]) & (g151) & (g549) & (!g532) & (!g552)));
	assign g554 = (((!sk[60]) & (g95) & (!g461)) + ((!sk[60]) & (g95) & (g461)) + ((sk[60]) & (g95) & (g461)));
	assign g555 = (((g13) & (!sk[61]) & (!g93)) + ((g13) & (!sk[61]) & (g93)) + ((g13) & (sk[61]) & (!g93)));
	assign g556 = (((!g554) & (sk[62]) & (!g555)) + ((g554) & (!sk[62]) & (!g555)) + ((g554) & (!sk[62]) & (g555)));
	assign g557 = (((!sk[63]) & (!g18) & (!g15) & (g13) & (g461)) + ((!sk[63]) & (!g18) & (g15) & (!g13) & (!g461)) + ((!sk[63]) & (!g18) & (g15) & (!g13) & (g461)) + ((!sk[63]) & (!g18) & (g15) & (g13) & (!g461)) + ((!sk[63]) & (!g18) & (g15) & (g13) & (g461)) + ((!sk[63]) & (g18) & (!g15) & (g13) & (!g461)) + ((!sk[63]) & (g18) & (!g15) & (g13) & (g461)) + ((!sk[63]) & (g18) & (g15) & (!g13) & (!g461)) + ((!sk[63]) & (g18) & (g15) & (!g13) & (g461)) + ((!sk[63]) & (g18) & (g15) & (g13) & (!g461)) + ((!sk[63]) & (g18) & (g15) & (g13) & (g461)) + ((sk[63]) & (!g18) & (!g15) & (!g13) & (g461)) + ((sk[63]) & (!g18) & (!g15) & (g13) & (!g461)) + ((sk[63]) & (!g18) & (!g15) & (g13) & (g461)) + ((sk[63]) & (!g18) & (g15) & (g13) & (!g461)) + ((sk[63]) & (!g18) & (g15) & (g13) & (g461)) + ((sk[63]) & (g18) & (!g15) & (!g13) & (g461)) + ((sk[63]) & (g18) & (!g15) & (g13) & (g461)));
	assign g558 = (((!sk[64]) & (g45) & (!g556) & (!g557)) + ((!sk[64]) & (g45) & (!g556) & (g557)) + ((!sk[64]) & (g45) & (g556) & (!g557)) + ((!sk[64]) & (g45) & (g556) & (g557)) + ((sk[64]) & (!g45) & (g556) & (!g557)));
	assign g559 = (((!sk[65]) & (!g109) & (!g186) & (!g330) & (!g544) & (g558)) + ((!sk[65]) & (!g109) & (!g186) & (!g330) & (g544) & (g558)) + ((!sk[65]) & (!g109) & (!g186) & (g330) & (!g544) & (g558)) + ((!sk[65]) & (!g109) & (!g186) & (g330) & (g544) & (g558)) + ((!sk[65]) & (!g109) & (g186) & (!g330) & (!g544) & (g558)) + ((!sk[65]) & (!g109) & (g186) & (!g330) & (g544) & (g558)) + ((!sk[65]) & (!g109) & (g186) & (g330) & (!g544) & (g558)) + ((!sk[65]) & (!g109) & (g186) & (g330) & (g544) & (g558)) + ((!sk[65]) & (g109) & (!g186) & (!g330) & (!g544) & (!g558)) + ((!sk[65]) & (g109) & (!g186) & (!g330) & (!g544) & (g558)) + ((!sk[65]) & (g109) & (!g186) & (!g330) & (g544) & (!g558)) + ((!sk[65]) & (g109) & (!g186) & (!g330) & (g544) & (g558)) + ((!sk[65]) & (g109) & (!g186) & (g330) & (!g544) & (!g558)) + ((!sk[65]) & (g109) & (!g186) & (g330) & (!g544) & (g558)) + ((!sk[65]) & (g109) & (!g186) & (g330) & (g544) & (!g558)) + ((!sk[65]) & (g109) & (!g186) & (g330) & (g544) & (g558)) + ((!sk[65]) & (g109) & (g186) & (!g330) & (!g544) & (!g558)) + ((!sk[65]) & (g109) & (g186) & (!g330) & (!g544) & (g558)) + ((!sk[65]) & (g109) & (g186) & (!g330) & (g544) & (!g558)) + ((!sk[65]) & (g109) & (g186) & (!g330) & (g544) & (g558)) + ((!sk[65]) & (g109) & (g186) & (g330) & (!g544) & (!g558)) + ((!sk[65]) & (g109) & (g186) & (g330) & (!g544) & (g558)) + ((!sk[65]) & (g109) & (g186) & (g330) & (g544) & (!g558)) + ((!sk[65]) & (g109) & (g186) & (g330) & (g544) & (g558)) + ((sk[65]) & (!g109) & (!g186) & (!g330) & (g544) & (g558)) + ((sk[65]) & (!g109) & (!g186) & (g330) & (!g544) & (!g558)) + ((sk[65]) & (!g109) & (!g186) & (g330) & (!g544) & (g558)) + ((sk[65]) & (!g109) & (!g186) & (g330) & (g544) & (!g558)) + ((sk[65]) & (!g109) & (!g186) & (g330) & (g544) & (g558)) + ((sk[65]) & (!g109) & (g186) & (!g330) & (g544) & (g558)) + ((sk[65]) & (!g109) & (g186) & (g330) & (g544) & (!g558)) + ((sk[65]) & (!g109) & (g186) & (g330) & (g544) & (g558)) + ((sk[65]) & (g109) & (!g186) & (!g330) & (g544) & (g558)) + ((sk[65]) & (g109) & (!g186) & (g330) & (g544) & (!g558)) + ((sk[65]) & (g109) & (!g186) & (g330) & (g544) & (g558)) + ((sk[65]) & (g109) & (g186) & (!g330) & (g544) & (g558)) + ((sk[65]) & (g109) & (g186) & (g330) & (g544) & (!g558)) + ((sk[65]) & (g109) & (g186) & (g330) & (g544) & (g558)));
	assign g560 = (((!sk[66]) & (g13) & (!g22)) + ((!sk[66]) & (g13) & (g22)) + ((sk[66]) & (g13) & (g22)));
	assign g561 = (((g11) & (!sk[67]) & (!g461)) + ((g11) & (!sk[67]) & (g461)) + ((g11) & (sk[67]) & (g461)));
	assign g562 = (((!sk[68]) & (g112) & (!g560) & (!g561)) + ((!sk[68]) & (g112) & (!g560) & (g561)) + ((!sk[68]) & (g112) & (g560) & (!g561)) + ((!sk[68]) & (g112) & (g560) & (g561)) + ((sk[68]) & (g112) & (!g560) & (g561)) + ((sk[68]) & (g112) & (g560) & (!g561)) + ((sk[68]) & (g112) & (g560) & (g561)));
	assign g563 = (((!sk[69]) & (!i_8_) & (!g15) & (!g11) & (!g108) & (g461)) + ((!sk[69]) & (!i_8_) & (!g15) & (!g11) & (g108) & (g461)) + ((!sk[69]) & (!i_8_) & (!g15) & (g11) & (!g108) & (g461)) + ((!sk[69]) & (!i_8_) & (!g15) & (g11) & (g108) & (g461)) + ((!sk[69]) & (!i_8_) & (g15) & (!g11) & (!g108) & (g461)) + ((!sk[69]) & (!i_8_) & (g15) & (!g11) & (g108) & (g461)) + ((!sk[69]) & (!i_8_) & (g15) & (g11) & (!g108) & (g461)) + ((!sk[69]) & (!i_8_) & (g15) & (g11) & (g108) & (g461)) + ((!sk[69]) & (i_8_) & (!g15) & (!g11) & (!g108) & (!g461)) + ((!sk[69]) & (i_8_) & (!g15) & (!g11) & (!g108) & (g461)) + ((!sk[69]) & (i_8_) & (!g15) & (!g11) & (g108) & (!g461)) + ((!sk[69]) & (i_8_) & (!g15) & (!g11) & (g108) & (g461)) + ((!sk[69]) & (i_8_) & (!g15) & (g11) & (!g108) & (!g461)) + ((!sk[69]) & (i_8_) & (!g15) & (g11) & (!g108) & (g461)) + ((!sk[69]) & (i_8_) & (!g15) & (g11) & (g108) & (!g461)) + ((!sk[69]) & (i_8_) & (!g15) & (g11) & (g108) & (g461)) + ((!sk[69]) & (i_8_) & (g15) & (!g11) & (!g108) & (!g461)) + ((!sk[69]) & (i_8_) & (g15) & (!g11) & (!g108) & (g461)) + ((!sk[69]) & (i_8_) & (g15) & (!g11) & (g108) & (!g461)) + ((!sk[69]) & (i_8_) & (g15) & (!g11) & (g108) & (g461)) + ((!sk[69]) & (i_8_) & (g15) & (g11) & (!g108) & (!g461)) + ((!sk[69]) & (i_8_) & (g15) & (g11) & (!g108) & (g461)) + ((!sk[69]) & (i_8_) & (g15) & (g11) & (g108) & (!g461)) + ((!sk[69]) & (i_8_) & (g15) & (g11) & (g108) & (g461)) + ((sk[69]) & (!i_8_) & (!g15) & (!g11) & (g108) & (g461)) + ((sk[69]) & (!i_8_) & (!g15) & (g11) & (g108) & (g461)) + ((sk[69]) & (!i_8_) & (g15) & (g11) & (g108) & (g461)) + ((sk[69]) & (i_8_) & (!g15) & (g11) & (g108) & (g461)) + ((sk[69]) & (i_8_) & (g15) & (g11) & (g108) & (g461)));
	assign g564 = (((!i_8_) & (!g108) & (g548) & (!sk[70]) & (g554)) + ((!i_8_) & (g108) & (!g548) & (!sk[70]) & (!g554)) + ((!i_8_) & (g108) & (!g548) & (!sk[70]) & (g554)) + ((!i_8_) & (g108) & (!g548) & (sk[70]) & (g554)) + ((!i_8_) & (g108) & (g548) & (!sk[70]) & (!g554)) + ((!i_8_) & (g108) & (g548) & (!sk[70]) & (g554)) + ((!i_8_) & (g108) & (g548) & (sk[70]) & (!g554)) + ((!i_8_) & (g108) & (g548) & (sk[70]) & (g554)) + ((i_8_) & (!g108) & (g548) & (!sk[70]) & (!g554)) + ((i_8_) & (!g108) & (g548) & (!sk[70]) & (g554)) + ((i_8_) & (g108) & (!g548) & (!sk[70]) & (!g554)) + ((i_8_) & (g108) & (!g548) & (!sk[70]) & (g554)) + ((i_8_) & (g108) & (g548) & (!sk[70]) & (!g554)) + ((i_8_) & (g108) & (g548) & (!sk[70]) & (g554)));
	assign g565 = (((!g100) & (!g136) & (!g560) & (!g562) & (!g563) & (!g564)) + ((!g100) & (!g136) & (g560) & (!g562) & (!g563) & (!g564)) + ((!g100) & (g136) & (!g560) & (!g562) & (!g563) & (!g564)) + ((g100) & (!g136) & (!g560) & (!g562) & (!g563) & (!g564)) + ((g100) & (g136) & (!g560) & (!g562) & (!g563) & (!g564)));
	assign g566 = (((!sk[72]) & (g13) & (!g158)) + ((!sk[72]) & (g13) & (g158)) + ((sk[72]) & (g13) & (g158)));
	assign g567 = (((!g131) & (!g251) & (!g461) & (!sk[73]) & (!g566) & (g556)) + ((!g131) & (!g251) & (!g461) & (!sk[73]) & (g566) & (g556)) + ((!g131) & (!g251) & (g461) & (!sk[73]) & (!g566) & (g556)) + ((!g131) & (!g251) & (g461) & (!sk[73]) & (g566) & (g556)) + ((!g131) & (g251) & (!g461) & (!sk[73]) & (!g566) & (g556)) + ((!g131) & (g251) & (!g461) & (!sk[73]) & (g566) & (g556)) + ((!g131) & (g251) & (!g461) & (sk[73]) & (!g566) & (!g556)) + ((!g131) & (g251) & (!g461) & (sk[73]) & (g566) & (!g556)) + ((!g131) & (g251) & (!g461) & (sk[73]) & (g566) & (g556)) + ((!g131) & (g251) & (g461) & (!sk[73]) & (!g566) & (g556)) + ((!g131) & (g251) & (g461) & (!sk[73]) & (g566) & (g556)) + ((!g131) & (g251) & (g461) & (sk[73]) & (!g566) & (!g556)) + ((!g131) & (g251) & (g461) & (sk[73]) & (g566) & (!g556)) + ((!g131) & (g251) & (g461) & (sk[73]) & (g566) & (g556)) + ((g131) & (!g251) & (!g461) & (!sk[73]) & (!g566) & (!g556)) + ((g131) & (!g251) & (!g461) & (!sk[73]) & (!g566) & (g556)) + ((g131) & (!g251) & (!g461) & (!sk[73]) & (g566) & (!g556)) + ((g131) & (!g251) & (!g461) & (!sk[73]) & (g566) & (g556)) + ((g131) & (!g251) & (g461) & (!sk[73]) & (!g566) & (!g556)) + ((g131) & (!g251) & (g461) & (!sk[73]) & (!g566) & (g556)) + ((g131) & (!g251) & (g461) & (!sk[73]) & (g566) & (!g556)) + ((g131) & (!g251) & (g461) & (!sk[73]) & (g566) & (g556)) + ((g131) & (g251) & (!g461) & (!sk[73]) & (!g566) & (!g556)) + ((g131) & (g251) & (!g461) & (!sk[73]) & (!g566) & (g556)) + ((g131) & (g251) & (!g461) & (!sk[73]) & (g566) & (!g556)) + ((g131) & (g251) & (!g461) & (!sk[73]) & (g566) & (g556)) + ((g131) & (g251) & (!g461) & (sk[73]) & (!g566) & (!g556)) + ((g131) & (g251) & (!g461) & (sk[73]) & (g566) & (!g556)) + ((g131) & (g251) & (!g461) & (sk[73]) & (g566) & (g556)) + ((g131) & (g251) & (g461) & (!sk[73]) & (!g566) & (!g556)) + ((g131) & (g251) & (g461) & (!sk[73]) & (!g566) & (g556)) + ((g131) & (g251) & (g461) & (!sk[73]) & (g566) & (!g556)) + ((g131) & (g251) & (g461) & (!sk[73]) & (g566) & (g556)) + ((g131) & (g251) & (g461) & (sk[73]) & (!g566) & (!g556)) + ((g131) & (g251) & (g461) & (sk[73]) & (!g566) & (g556)) + ((g131) & (g251) & (g461) & (sk[73]) & (g566) & (!g556)) + ((g131) & (g251) & (g461) & (sk[73]) & (g566) & (g556)));
	assign g568 = (((!g545) & (g1708) & (g553) & (g559) & (g565) & (!g567)));
	assign g569 = (((g112) & (!sk[75]) & (!g566)) + ((g112) & (!sk[75]) & (g566)) + ((g112) & (sk[75]) & (g566)));
	assign g570 = (((i_14_) & (!i_12_) & (!i_13_) & (g99) & (!g101) & (!g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (g99) & (g101) & (!g115)) + ((i_14_) & (!i_12_) & (i_13_) & (!g99) & (g101) & (!g115)) + ((i_14_) & (!i_12_) & (i_13_) & (g99) & (!g101) & (!g115)) + ((i_14_) & (!i_12_) & (i_13_) & (g99) & (g101) & (!g115)) + ((i_14_) & (i_12_) & (!i_13_) & (!g99) & (g101) & (!g115)) + ((i_14_) & (i_12_) & (!i_13_) & (g99) & (!g101) & (!g115)) + ((i_14_) & (i_12_) & (!i_13_) & (g99) & (g101) & (!g115)));
	assign g571 = (((!sk[77]) & (!g45) & (!g547) & (g546) & (g532)) + ((!sk[77]) & (!g45) & (g547) & (!g546) & (!g532)) + ((!sk[77]) & (!g45) & (g547) & (!g546) & (g532)) + ((!sk[77]) & (!g45) & (g547) & (g546) & (!g532)) + ((!sk[77]) & (!g45) & (g547) & (g546) & (g532)) + ((!sk[77]) & (g45) & (!g547) & (g546) & (!g532)) + ((!sk[77]) & (g45) & (!g547) & (g546) & (g532)) + ((!sk[77]) & (g45) & (g547) & (!g546) & (!g532)) + ((!sk[77]) & (g45) & (g547) & (!g546) & (g532)) + ((!sk[77]) & (g45) & (g547) & (g546) & (!g532)) + ((!sk[77]) & (g45) & (g547) & (g546) & (g532)) + ((sk[77]) & (!g45) & (g547) & (!g546) & (!g532)));
	assign g572 = (((i_14_) & (!i_12_) & (!sk[78]) & (!i_13_)) + ((i_14_) & (!i_12_) & (!sk[78]) & (i_13_)) + ((i_14_) & (!i_12_) & (sk[78]) & (i_13_)) + ((i_14_) & (i_12_) & (!sk[78]) & (!i_13_)) + ((i_14_) & (i_12_) & (!sk[78]) & (i_13_)) + ((i_14_) & (i_12_) & (sk[78]) & (!i_13_)));
	assign g573 = (((!g13) & (!sk[79]) & (!g99) & (!g100) & (!g124) & (g572)) + ((!g13) & (!sk[79]) & (!g99) & (!g100) & (g124) & (g572)) + ((!g13) & (!sk[79]) & (!g99) & (g100) & (!g124) & (g572)) + ((!g13) & (!sk[79]) & (!g99) & (g100) & (g124) & (g572)) + ((!g13) & (!sk[79]) & (g99) & (!g100) & (!g124) & (g572)) + ((!g13) & (!sk[79]) & (g99) & (!g100) & (g124) & (g572)) + ((!g13) & (!sk[79]) & (g99) & (g100) & (!g124) & (g572)) + ((!g13) & (!sk[79]) & (g99) & (g100) & (g124) & (g572)) + ((!g13) & (sk[79]) & (!g99) & (g100) & (g124) & (g572)) + ((!g13) & (sk[79]) & (g99) & (g100) & (g124) & (g572)) + ((g13) & (!sk[79]) & (!g99) & (!g100) & (!g124) & (!g572)) + ((g13) & (!sk[79]) & (!g99) & (!g100) & (!g124) & (g572)) + ((g13) & (!sk[79]) & (!g99) & (!g100) & (g124) & (!g572)) + ((g13) & (!sk[79]) & (!g99) & (!g100) & (g124) & (g572)) + ((g13) & (!sk[79]) & (!g99) & (g100) & (!g124) & (!g572)) + ((g13) & (!sk[79]) & (!g99) & (g100) & (!g124) & (g572)) + ((g13) & (!sk[79]) & (!g99) & (g100) & (g124) & (!g572)) + ((g13) & (!sk[79]) & (!g99) & (g100) & (g124) & (g572)) + ((g13) & (!sk[79]) & (g99) & (!g100) & (!g124) & (!g572)) + ((g13) & (!sk[79]) & (g99) & (!g100) & (!g124) & (g572)) + ((g13) & (!sk[79]) & (g99) & (!g100) & (g124) & (!g572)) + ((g13) & (!sk[79]) & (g99) & (!g100) & (g124) & (g572)) + ((g13) & (!sk[79]) & (g99) & (g100) & (!g124) & (!g572)) + ((g13) & (!sk[79]) & (g99) & (g100) & (!g124) & (g572)) + ((g13) & (!sk[79]) & (g99) & (g100) & (g124) & (!g572)) + ((g13) & (!sk[79]) & (g99) & (g100) & (g124) & (g572)) + ((g13) & (sk[79]) & (!g99) & (g100) & (g124) & (g572)) + ((g13) & (sk[79]) & (g99) & (!g100) & (g124) & (!g572)) + ((g13) & (sk[79]) & (g99) & (!g100) & (g124) & (g572)) + ((g13) & (sk[79]) & (g99) & (g100) & (g124) & (!g572)) + ((g13) & (sk[79]) & (g99) & (g100) & (g124) & (g572)));
	assign g574 = (((!g122) & (sk[80]) & (g572)) + ((g122) & (!sk[80]) & (!g572)) + ((g122) & (!sk[80]) & (g572)));
	assign g575 = (((!g101) & (!g224) & (!g467) & (!g571) & (!g573) & (!g574)) + ((!g101) & (!g224) & (!g467) & (!g571) & (!g573) & (g574)) + ((!g101) & (!g224) & (!g467) & (g571) & (!g573) & (!g574)) + ((!g101) & (!g224) & (!g467) & (g571) & (!g573) & (g574)) + ((!g101) & (!g224) & (g467) & (!g571) & (!g573) & (!g574)) + ((!g101) & (!g224) & (g467) & (!g571) & (!g573) & (g574)) + ((!g101) & (!g224) & (g467) & (g571) & (!g573) & (!g574)) + ((!g101) & (!g224) & (g467) & (g571) & (!g573) & (g574)) + ((!g101) & (g224) & (!g467) & (!g571) & (!g573) & (!g574)) + ((!g101) & (g224) & (!g467) & (!g571) & (!g573) & (g574)) + ((!g101) & (g224) & (!g467) & (g571) & (!g573) & (!g574)) + ((!g101) & (g224) & (!g467) & (g571) & (!g573) & (g574)) + ((!g101) & (g224) & (g467) & (!g571) & (!g573) & (!g574)) + ((!g101) & (g224) & (g467) & (!g571) & (!g573) & (g574)) + ((!g101) & (g224) & (g467) & (g571) & (!g573) & (!g574)) + ((!g101) & (g224) & (g467) & (g571) & (!g573) & (g574)) + ((g101) & (!g224) & (g467) & (g571) & (!g573) & (!g574)));
	assign g576 = (((!sk[82]) & (g131) & (!g461) & (!g566)) + ((!sk[82]) & (g131) & (!g461) & (g566)) + ((!sk[82]) & (g131) & (g461) & (!g566)) + ((!sk[82]) & (g131) & (g461) & (g566)) + ((sk[82]) & (!g131) & (!g461) & (!g566)) + ((sk[82]) & (!g131) & (g461) & (!g566)) + ((sk[82]) & (g131) & (!g461) & (!g566)));
	assign g577 = (((!i_8_) & (!sk[83]) & (!g88) & (g284) & (g576)) + ((!i_8_) & (!sk[83]) & (g88) & (!g284) & (!g576)) + ((!i_8_) & (!sk[83]) & (g88) & (!g284) & (g576)) + ((!i_8_) & (!sk[83]) & (g88) & (g284) & (!g576)) + ((!i_8_) & (!sk[83]) & (g88) & (g284) & (g576)) + ((!i_8_) & (sk[83]) & (!g88) & (g284) & (!g576)) + ((!i_8_) & (sk[83]) & (g88) & (g284) & (!g576)) + ((i_8_) & (!sk[83]) & (!g88) & (g284) & (!g576)) + ((i_8_) & (!sk[83]) & (!g88) & (g284) & (g576)) + ((i_8_) & (!sk[83]) & (g88) & (!g284) & (!g576)) + ((i_8_) & (!sk[83]) & (g88) & (!g284) & (g576)) + ((i_8_) & (!sk[83]) & (g88) & (g284) & (!g576)) + ((i_8_) & (!sk[83]) & (g88) & (g284) & (g576)) + ((i_8_) & (sk[83]) & (!g88) & (g284) & (!g576)) + ((i_8_) & (sk[83]) & (g88) & (!g284) & (!g576)) + ((i_8_) & (sk[83]) & (g88) & (g284) & (!g576)));
	assign g578 = (((!i_8_) & (!g15) & (!sk[84]) & (!g119) & (!g108) & (g461)) + ((!i_8_) & (!g15) & (!sk[84]) & (!g119) & (g108) & (g461)) + ((!i_8_) & (!g15) & (!sk[84]) & (g119) & (!g108) & (g461)) + ((!i_8_) & (!g15) & (!sk[84]) & (g119) & (g108) & (g461)) + ((!i_8_) & (g15) & (!sk[84]) & (!g119) & (!g108) & (g461)) + ((!i_8_) & (g15) & (!sk[84]) & (!g119) & (g108) & (g461)) + ((!i_8_) & (g15) & (!sk[84]) & (g119) & (!g108) & (g461)) + ((!i_8_) & (g15) & (!sk[84]) & (g119) & (g108) & (g461)) + ((i_8_) & (!g15) & (!sk[84]) & (!g119) & (!g108) & (!g461)) + ((i_8_) & (!g15) & (!sk[84]) & (!g119) & (!g108) & (g461)) + ((i_8_) & (!g15) & (!sk[84]) & (!g119) & (g108) & (!g461)) + ((i_8_) & (!g15) & (!sk[84]) & (!g119) & (g108) & (g461)) + ((i_8_) & (!g15) & (!sk[84]) & (g119) & (!g108) & (!g461)) + ((i_8_) & (!g15) & (!sk[84]) & (g119) & (!g108) & (g461)) + ((i_8_) & (!g15) & (!sk[84]) & (g119) & (g108) & (!g461)) + ((i_8_) & (!g15) & (!sk[84]) & (g119) & (g108) & (g461)) + ((i_8_) & (!g15) & (sk[84]) & (!g119) & (g108) & (g461)) + ((i_8_) & (!g15) & (sk[84]) & (g119) & (g108) & (g461)) + ((i_8_) & (g15) & (!sk[84]) & (!g119) & (!g108) & (!g461)) + ((i_8_) & (g15) & (!sk[84]) & (!g119) & (!g108) & (g461)) + ((i_8_) & (g15) & (!sk[84]) & (!g119) & (g108) & (!g461)) + ((i_8_) & (g15) & (!sk[84]) & (!g119) & (g108) & (g461)) + ((i_8_) & (g15) & (!sk[84]) & (g119) & (!g108) & (!g461)) + ((i_8_) & (g15) & (!sk[84]) & (g119) & (!g108) & (g461)) + ((i_8_) & (g15) & (!sk[84]) & (g119) & (g108) & (!g461)) + ((i_8_) & (g15) & (!sk[84]) & (g119) & (g108) & (g461)) + ((i_8_) & (g15) & (sk[84]) & (g119) & (g108) & (g461)));
	assign g579 = (((!i_8_) & (!g108) & (!sk[85]) & (g554) & (g550)) + ((!i_8_) & (g108) & (!sk[85]) & (!g554) & (!g550)) + ((!i_8_) & (g108) & (!sk[85]) & (!g554) & (g550)) + ((!i_8_) & (g108) & (!sk[85]) & (g554) & (!g550)) + ((!i_8_) & (g108) & (!sk[85]) & (g554) & (g550)) + ((i_8_) & (!g108) & (!sk[85]) & (g554) & (!g550)) + ((i_8_) & (!g108) & (!sk[85]) & (g554) & (g550)) + ((i_8_) & (g108) & (!sk[85]) & (!g554) & (!g550)) + ((i_8_) & (g108) & (!sk[85]) & (!g554) & (g550)) + ((i_8_) & (g108) & (!sk[85]) & (g554) & (!g550)) + ((i_8_) & (g108) & (!sk[85]) & (g554) & (g550)) + ((i_8_) & (g108) & (sk[85]) & (!g554) & (g550)) + ((i_8_) & (g108) & (sk[85]) & (g554) & (!g550)) + ((i_8_) & (g108) & (sk[85]) & (g554) & (g550)));
	assign g580 = (((!g338) & (!g577) & (!sk[86]) & (!g556) & (!g578) & (g579)) + ((!g338) & (!g577) & (!sk[86]) & (!g556) & (g578) & (g579)) + ((!g338) & (!g577) & (!sk[86]) & (g556) & (!g578) & (g579)) + ((!g338) & (!g577) & (!sk[86]) & (g556) & (g578) & (g579)) + ((!g338) & (!g577) & (sk[86]) & (g556) & (!g578) & (!g579)) + ((!g338) & (g577) & (!sk[86]) & (!g556) & (!g578) & (g579)) + ((!g338) & (g577) & (!sk[86]) & (!g556) & (g578) & (g579)) + ((!g338) & (g577) & (!sk[86]) & (g556) & (!g578) & (g579)) + ((!g338) & (g577) & (!sk[86]) & (g556) & (g578) & (g579)) + ((g338) & (!g577) & (!sk[86]) & (!g556) & (!g578) & (!g579)) + ((g338) & (!g577) & (!sk[86]) & (!g556) & (!g578) & (g579)) + ((g338) & (!g577) & (!sk[86]) & (!g556) & (g578) & (!g579)) + ((g338) & (!g577) & (!sk[86]) & (!g556) & (g578) & (g579)) + ((g338) & (!g577) & (!sk[86]) & (g556) & (!g578) & (!g579)) + ((g338) & (!g577) & (!sk[86]) & (g556) & (!g578) & (g579)) + ((g338) & (!g577) & (!sk[86]) & (g556) & (g578) & (!g579)) + ((g338) & (!g577) & (!sk[86]) & (g556) & (g578) & (g579)) + ((g338) & (!g577) & (sk[86]) & (!g556) & (!g578) & (!g579)) + ((g338) & (!g577) & (sk[86]) & (g556) & (!g578) & (!g579)) + ((g338) & (g577) & (!sk[86]) & (!g556) & (!g578) & (!g579)) + ((g338) & (g577) & (!sk[86]) & (!g556) & (!g578) & (g579)) + ((g338) & (g577) & (!sk[86]) & (!g556) & (g578) & (!g579)) + ((g338) & (g577) & (!sk[86]) & (!g556) & (g578) & (g579)) + ((g338) & (g577) & (!sk[86]) & (g556) & (!g578) & (!g579)) + ((g338) & (g577) & (!sk[86]) & (g556) & (!g578) & (g579)) + ((g338) & (g577) & (!sk[86]) & (g556) & (g578) & (!g579)) + ((g338) & (g577) & (!sk[86]) & (g556) & (g578) & (g579)));
	assign g581 = (((!g102) & (!sk[87]) & (!g112) & (!g131) & (!g461) & (g546)) + ((!g102) & (!sk[87]) & (!g112) & (!g131) & (g461) & (g546)) + ((!g102) & (!sk[87]) & (!g112) & (g131) & (!g461) & (g546)) + ((!g102) & (!sk[87]) & (!g112) & (g131) & (g461) & (g546)) + ((!g102) & (!sk[87]) & (g112) & (!g131) & (!g461) & (g546)) + ((!g102) & (!sk[87]) & (g112) & (!g131) & (g461) & (g546)) + ((!g102) & (!sk[87]) & (g112) & (g131) & (!g461) & (g546)) + ((!g102) & (!sk[87]) & (g112) & (g131) & (g461) & (g546)) + ((!g102) & (sk[87]) & (g112) & (!g131) & (!g461) & (g546)) + ((!g102) & (sk[87]) & (g112) & (!g131) & (g461) & (!g546)) + ((!g102) & (sk[87]) & (g112) & (!g131) & (g461) & (g546)) + ((!g102) & (sk[87]) & (g112) & (g131) & (!g461) & (g546)) + ((!g102) & (sk[87]) & (g112) & (g131) & (g461) & (!g546)) + ((!g102) & (sk[87]) & (g112) & (g131) & (g461) & (g546)) + ((g102) & (!sk[87]) & (!g112) & (!g131) & (!g461) & (!g546)) + ((g102) & (!sk[87]) & (!g112) & (!g131) & (!g461) & (g546)) + ((g102) & (!sk[87]) & (!g112) & (!g131) & (g461) & (!g546)) + ((g102) & (!sk[87]) & (!g112) & (!g131) & (g461) & (g546)) + ((g102) & (!sk[87]) & (!g112) & (g131) & (!g461) & (!g546)) + ((g102) & (!sk[87]) & (!g112) & (g131) & (!g461) & (g546)) + ((g102) & (!sk[87]) & (!g112) & (g131) & (g461) & (!g546)) + ((g102) & (!sk[87]) & (!g112) & (g131) & (g461) & (g546)) + ((g102) & (!sk[87]) & (g112) & (!g131) & (!g461) & (!g546)) + ((g102) & (!sk[87]) & (g112) & (!g131) & (!g461) & (g546)) + ((g102) & (!sk[87]) & (g112) & (!g131) & (g461) & (!g546)) + ((g102) & (!sk[87]) & (g112) & (!g131) & (g461) & (g546)) + ((g102) & (!sk[87]) & (g112) & (g131) & (!g461) & (!g546)) + ((g102) & (!sk[87]) & (g112) & (g131) & (!g461) & (g546)) + ((g102) & (!sk[87]) & (g112) & (g131) & (g461) & (!g546)) + ((g102) & (!sk[87]) & (g112) & (g131) & (g461) & (g546)) + ((g102) & (sk[87]) & (g112) & (!g131) & (!g461) & (g546)) + ((g102) & (sk[87]) & (g112) & (!g131) & (g461) & (g546)) + ((g102) & (sk[87]) & (g112) & (g131) & (!g461) & (g546)) + ((g102) & (sk[87]) & (g112) & (g131) & (g461) & (!g546)) + ((g102) & (sk[87]) & (g112) & (g131) & (g461) & (g546)));
	assign g582 = (((!g151) & (sk[88]) & (!g554) & (!g581)) + ((!g151) & (sk[88]) & (g554) & (!g581)) + ((g151) & (!sk[88]) & (!g554) & (!g581)) + ((g151) & (!sk[88]) & (!g554) & (g581)) + ((g151) & (!sk[88]) & (g554) & (!g581)) + ((g151) & (!sk[88]) & (g554) & (g581)) + ((g151) & (sk[88]) & (!g554) & (!g581)));
	assign g583 = (((!g45) & (!sk[89]) & (!g195) & (g532) & (g478)) + ((!g45) & (!sk[89]) & (g195) & (!g532) & (!g478)) + ((!g45) & (!sk[89]) & (g195) & (!g532) & (g478)) + ((!g45) & (!sk[89]) & (g195) & (g532) & (!g478)) + ((!g45) & (!sk[89]) & (g195) & (g532) & (g478)) + ((!g45) & (sk[89]) & (!g195) & (!g532) & (!g478)) + ((g45) & (!sk[89]) & (!g195) & (g532) & (!g478)) + ((g45) & (!sk[89]) & (!g195) & (g532) & (g478)) + ((g45) & (!sk[89]) & (g195) & (!g532) & (!g478)) + ((g45) & (!sk[89]) & (g195) & (!g532) & (g478)) + ((g45) & (!sk[89]) & (g195) & (g532) & (!g478)) + ((g45) & (!sk[89]) & (g195) & (g532) & (g478)));
	assign g584 = (((!i_11_) & (!i_9_) & (!sk[90]) & (g48) & (g214)) + ((!i_11_) & (i_9_) & (!sk[90]) & (!g48) & (!g214)) + ((!i_11_) & (i_9_) & (!sk[90]) & (!g48) & (g214)) + ((!i_11_) & (i_9_) & (!sk[90]) & (g48) & (!g214)) + ((!i_11_) & (i_9_) & (!sk[90]) & (g48) & (g214)) + ((i_11_) & (!i_9_) & (!sk[90]) & (g48) & (!g214)) + ((i_11_) & (!i_9_) & (!sk[90]) & (g48) & (g214)) + ((i_11_) & (!i_9_) & (sk[90]) & (!g48) & (g214)) + ((i_11_) & (i_9_) & (!sk[90]) & (!g48) & (!g214)) + ((i_11_) & (i_9_) & (!sk[90]) & (!g48) & (g214)) + ((i_11_) & (i_9_) & (!sk[90]) & (g48) & (!g214)) + ((i_11_) & (i_9_) & (!sk[90]) & (g48) & (g214)));
	assign g585 = (((g141) & (!sk[91]) & (!g99) & (!g171)) + ((g141) & (!sk[91]) & (!g99) & (g171)) + ((g141) & (!sk[91]) & (g99) & (!g171)) + ((g141) & (!sk[91]) & (g99) & (g171)) + ((g141) & (sk[91]) & (g99) & (!g171)));
	assign g586 = (((!i_15_) & (!g89) & (!g583) & (!sk[92]) & (!g584) & (g585)) + ((!i_15_) & (!g89) & (!g583) & (!sk[92]) & (g584) & (g585)) + ((!i_15_) & (!g89) & (g583) & (!sk[92]) & (!g584) & (g585)) + ((!i_15_) & (!g89) & (g583) & (!sk[92]) & (g584) & (g585)) + ((!i_15_) & (!g89) & (g583) & (sk[92]) & (!g584) & (!g585)) + ((!i_15_) & (!g89) & (g583) & (sk[92]) & (!g584) & (g585)) + ((!i_15_) & (!g89) & (g583) & (sk[92]) & (g584) & (!g585)) + ((!i_15_) & (!g89) & (g583) & (sk[92]) & (g584) & (g585)) + ((!i_15_) & (g89) & (!g583) & (!sk[92]) & (!g584) & (g585)) + ((!i_15_) & (g89) & (!g583) & (!sk[92]) & (g584) & (g585)) + ((!i_15_) & (g89) & (!g583) & (sk[92]) & (!g584) & (!g585)) + ((!i_15_) & (g89) & (!g583) & (sk[92]) & (!g584) & (g585)) + ((!i_15_) & (g89) & (!g583) & (sk[92]) & (g584) & (!g585)) + ((!i_15_) & (g89) & (!g583) & (sk[92]) & (g584) & (g585)) + ((!i_15_) & (g89) & (g583) & (!sk[92]) & (!g584) & (g585)) + ((!i_15_) & (g89) & (g583) & (!sk[92]) & (g584) & (g585)) + ((!i_15_) & (g89) & (g583) & (sk[92]) & (!g584) & (!g585)) + ((!i_15_) & (g89) & (g583) & (sk[92]) & (!g584) & (g585)) + ((!i_15_) & (g89) & (g583) & (sk[92]) & (g584) & (!g585)) + ((!i_15_) & (g89) & (g583) & (sk[92]) & (g584) & (g585)) + ((i_15_) & (!g89) & (!g583) & (!sk[92]) & (!g584) & (!g585)) + ((i_15_) & (!g89) & (!g583) & (!sk[92]) & (!g584) & (g585)) + ((i_15_) & (!g89) & (!g583) & (!sk[92]) & (g584) & (!g585)) + ((i_15_) & (!g89) & (!g583) & (!sk[92]) & (g584) & (g585)) + ((i_15_) & (!g89) & (g583) & (!sk[92]) & (!g584) & (!g585)) + ((i_15_) & (!g89) & (g583) & (!sk[92]) & (!g584) & (g585)) + ((i_15_) & (!g89) & (g583) & (!sk[92]) & (g584) & (!g585)) + ((i_15_) & (!g89) & (g583) & (!sk[92]) & (g584) & (g585)) + ((i_15_) & (!g89) & (g583) & (sk[92]) & (!g584) & (!g585)) + ((i_15_) & (g89) & (!g583) & (!sk[92]) & (!g584) & (!g585)) + ((i_15_) & (g89) & (!g583) & (!sk[92]) & (!g584) & (g585)) + ((i_15_) & (g89) & (!g583) & (!sk[92]) & (g584) & (!g585)) + ((i_15_) & (g89) & (!g583) & (!sk[92]) & (g584) & (g585)) + ((i_15_) & (g89) & (!g583) & (sk[92]) & (!g584) & (!g585)) + ((i_15_) & (g89) & (g583) & (!sk[92]) & (!g584) & (!g585)) + ((i_15_) & (g89) & (g583) & (!sk[92]) & (!g584) & (g585)) + ((i_15_) & (g89) & (g583) & (!sk[92]) & (g584) & (!g585)) + ((i_15_) & (g89) & (g583) & (!sk[92]) & (g584) & (g585)) + ((i_15_) & (g89) & (g583) & (sk[92]) & (!g584) & (!g585)));
	assign g587 = (((!g569) & (!g570) & (g575) & (g580) & (g582) & (g586)));
	assign g588 = (((!i_12_) & (!sk[94]) & (!i_13_) & (g18) & (g179)) + ((!i_12_) & (!sk[94]) & (i_13_) & (!g18) & (!g179)) + ((!i_12_) & (!sk[94]) & (i_13_) & (!g18) & (g179)) + ((!i_12_) & (!sk[94]) & (i_13_) & (g18) & (!g179)) + ((!i_12_) & (!sk[94]) & (i_13_) & (g18) & (g179)) + ((!i_12_) & (sk[94]) & (!i_13_) & (!g18) & (!g179)) + ((!i_12_) & (sk[94]) & (!i_13_) & (g18) & (!g179)) + ((!i_12_) & (sk[94]) & (i_13_) & (!g18) & (!g179)) + ((!i_12_) & (sk[94]) & (i_13_) & (g18) & (!g179)) + ((i_12_) & (!sk[94]) & (!i_13_) & (g18) & (!g179)) + ((i_12_) & (!sk[94]) & (!i_13_) & (g18) & (g179)) + ((i_12_) & (!sk[94]) & (i_13_) & (!g18) & (!g179)) + ((i_12_) & (!sk[94]) & (i_13_) & (!g18) & (g179)) + ((i_12_) & (!sk[94]) & (i_13_) & (g18) & (!g179)) + ((i_12_) & (!sk[94]) & (i_13_) & (g18) & (g179)) + ((i_12_) & (sk[94]) & (!i_13_) & (!g18) & (!g179)) + ((i_12_) & (sk[94]) & (!i_13_) & (g18) & (!g179)) + ((i_12_) & (sk[94]) & (i_13_) & (g18) & (!g179)));
	assign g589 = (((!g109) & (!g330) & (!g413) & (!g414) & (!g531) & (g588)) + ((!g109) & (g330) & (!g413) & (!g414) & (!g531) & (!g588)) + ((!g109) & (g330) & (!g413) & (!g414) & (!g531) & (g588)) + ((!g109) & (g330) & (!g413) & (!g414) & (g531) & (!g588)) + ((!g109) & (g330) & (!g413) & (!g414) & (g531) & (g588)) + ((g109) & (!g330) & (!g413) & (!g414) & (!g531) & (g588)) + ((g109) & (g330) & (!g413) & (!g414) & (!g531) & (!g588)) + ((g109) & (g330) & (!g413) & (!g414) & (!g531) & (g588)));
	assign g590 = (((!i_11_) & (!i_9_) & (!sk[96]) & (!i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (!i_9_) & (!sk[96]) & (!i_10_) & (i_15_) & (g461)) + ((!i_11_) & (!i_9_) & (!sk[96]) & (i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (!i_9_) & (!sk[96]) & (i_10_) & (i_15_) & (g461)) + ((!i_11_) & (!i_9_) & (sk[96]) & (!i_10_) & (!i_15_) & (!g461)) + ((!i_11_) & (!i_9_) & (sk[96]) & (!i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (!i_9_) & (sk[96]) & (!i_10_) & (i_15_) & (!g461)) + ((!i_11_) & (!i_9_) & (sk[96]) & (!i_10_) & (i_15_) & (g461)) + ((!i_11_) & (!i_9_) & (sk[96]) & (i_10_) & (!i_15_) & (!g461)) + ((!i_11_) & (!i_9_) & (sk[96]) & (i_10_) & (i_15_) & (!g461)) + ((!i_11_) & (!i_9_) & (sk[96]) & (i_10_) & (i_15_) & (g461)) + ((!i_11_) & (i_9_) & (!sk[96]) & (!i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (i_9_) & (!sk[96]) & (!i_10_) & (i_15_) & (g461)) + ((!i_11_) & (i_9_) & (!sk[96]) & (i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (i_9_) & (!sk[96]) & (i_10_) & (i_15_) & (g461)) + ((!i_11_) & (i_9_) & (sk[96]) & (!i_10_) & (!i_15_) & (!g461)) + ((!i_11_) & (i_9_) & (sk[96]) & (!i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (i_9_) & (sk[96]) & (!i_10_) & (i_15_) & (!g461)) + ((!i_11_) & (i_9_) & (sk[96]) & (!i_10_) & (i_15_) & (g461)) + ((!i_11_) & (i_9_) & (sk[96]) & (i_10_) & (!i_15_) & (!g461)) + ((!i_11_) & (i_9_) & (sk[96]) & (i_10_) & (i_15_) & (!g461)) + ((!i_11_) & (i_9_) & (sk[96]) & (i_10_) & (i_15_) & (g461)) + ((i_11_) & (!i_9_) & (!sk[96]) & (!i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (!i_9_) & (!sk[96]) & (!i_10_) & (!i_15_) & (g461)) + ((i_11_) & (!i_9_) & (!sk[96]) & (!i_10_) & (i_15_) & (!g461)) + ((i_11_) & (!i_9_) & (!sk[96]) & (!i_10_) & (i_15_) & (g461)) + ((i_11_) & (!i_9_) & (!sk[96]) & (i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (!i_9_) & (!sk[96]) & (i_10_) & (!i_15_) & (g461)) + ((i_11_) & (!i_9_) & (!sk[96]) & (i_10_) & (i_15_) & (!g461)) + ((i_11_) & (!i_9_) & (!sk[96]) & (i_10_) & (i_15_) & (g461)) + ((i_11_) & (!i_9_) & (sk[96]) & (!i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (!i_9_) & (sk[96]) & (!i_10_) & (!i_15_) & (g461)) + ((i_11_) & (!i_9_) & (sk[96]) & (!i_10_) & (i_15_) & (!g461)) + ((i_11_) & (!i_9_) & (sk[96]) & (!i_10_) & (i_15_) & (g461)) + ((i_11_) & (!i_9_) & (sk[96]) & (i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (!i_9_) & (sk[96]) & (i_10_) & (i_15_) & (!g461)) + ((i_11_) & (!i_9_) & (sk[96]) & (i_10_) & (i_15_) & (g461)) + ((i_11_) & (i_9_) & (!sk[96]) & (!i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (i_9_) & (!sk[96]) & (!i_10_) & (!i_15_) & (g461)) + ((i_11_) & (i_9_) & (!sk[96]) & (!i_10_) & (i_15_) & (!g461)) + ((i_11_) & (i_9_) & (!sk[96]) & (!i_10_) & (i_15_) & (g461)) + ((i_11_) & (i_9_) & (!sk[96]) & (i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (i_9_) & (!sk[96]) & (i_10_) & (!i_15_) & (g461)) + ((i_11_) & (i_9_) & (!sk[96]) & (i_10_) & (i_15_) & (!g461)) + ((i_11_) & (i_9_) & (!sk[96]) & (i_10_) & (i_15_) & (g461)) + ((i_11_) & (i_9_) & (sk[96]) & (!i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (i_9_) & (sk[96]) & (!i_10_) & (i_15_) & (!g461)) + ((i_11_) & (i_9_) & (sk[96]) & (i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (i_9_) & (sk[96]) & (i_10_) & (i_15_) & (!g461)) + ((i_11_) & (i_9_) & (sk[96]) & (i_10_) & (i_15_) & (g461)));
	assign g591 = (((!i_11_) & (!i_9_) & (!i_10_) & (!sk[97]) & (!i_15_) & (g171)) + ((!i_11_) & (!i_9_) & (!i_10_) & (!sk[97]) & (i_15_) & (g171)) + ((!i_11_) & (!i_9_) & (i_10_) & (!sk[97]) & (!i_15_) & (g171)) + ((!i_11_) & (!i_9_) & (i_10_) & (!sk[97]) & (i_15_) & (g171)) + ((!i_11_) & (!i_9_) & (i_10_) & (sk[97]) & (!i_15_) & (!g171)) + ((!i_11_) & (!i_9_) & (i_10_) & (sk[97]) & (i_15_) & (!g171)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[97]) & (!i_15_) & (g171)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[97]) & (i_15_) & (g171)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[97]) & (!i_15_) & (g171)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[97]) & (i_15_) & (g171)) + ((!i_11_) & (i_9_) & (i_10_) & (sk[97]) & (i_15_) & (!g171)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[97]) & (!i_15_) & (!g171)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[97]) & (!i_15_) & (g171)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[97]) & (i_15_) & (!g171)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[97]) & (i_15_) & (g171)) + ((i_11_) & (!i_9_) & (!i_10_) & (sk[97]) & (!i_15_) & (!g171)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[97]) & (!i_15_) & (!g171)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[97]) & (!i_15_) & (g171)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[97]) & (i_15_) & (!g171)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[97]) & (i_15_) & (g171)) + ((i_11_) & (!i_9_) & (i_10_) & (sk[97]) & (!i_15_) & (!g171)) + ((i_11_) & (!i_9_) & (i_10_) & (sk[97]) & (i_15_) & (!g171)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[97]) & (!i_15_) & (!g171)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[97]) & (!i_15_) & (g171)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[97]) & (i_15_) & (!g171)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[97]) & (i_15_) & (g171)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[97]) & (!i_15_) & (!g171)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[97]) & (!i_15_) & (g171)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[97]) & (i_15_) & (!g171)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[97]) & (i_15_) & (g171)) + ((i_11_) & (i_9_) & (i_10_) & (sk[97]) & (i_15_) & (!g171)));
	assign g592 = (((!g204) & (!sk[98]) & (!g279) & (!g460) & (!g470) & (g591)) + ((!g204) & (!sk[98]) & (!g279) & (!g460) & (g470) & (g591)) + ((!g204) & (!sk[98]) & (!g279) & (g460) & (!g470) & (g591)) + ((!g204) & (!sk[98]) & (!g279) & (g460) & (g470) & (g591)) + ((!g204) & (!sk[98]) & (g279) & (!g460) & (!g470) & (g591)) + ((!g204) & (!sk[98]) & (g279) & (!g460) & (g470) & (g591)) + ((!g204) & (!sk[98]) & (g279) & (g460) & (!g470) & (g591)) + ((!g204) & (!sk[98]) & (g279) & (g460) & (g470) & (g591)) + ((!g204) & (sk[98]) & (!g279) & (!g460) & (!g470) & (!g591)) + ((!g204) & (sk[98]) & (!g279) & (!g460) & (!g470) & (g591)) + ((!g204) & (sk[98]) & (!g279) & (!g460) & (g470) & (!g591)) + ((!g204) & (sk[98]) & (!g279) & (!g460) & (g470) & (g591)) + ((!g204) & (sk[98]) & (!g279) & (g460) & (!g470) & (!g591)) + ((!g204) & (sk[98]) & (!g279) & (g460) & (!g470) & (g591)) + ((!g204) & (sk[98]) & (!g279) & (g460) & (g470) & (!g591)) + ((!g204) & (sk[98]) & (!g279) & (g460) & (g470) & (g591)) + ((!g204) & (sk[98]) & (g279) & (!g460) & (!g470) & (!g591)) + ((!g204) & (sk[98]) & (g279) & (!g460) & (!g470) & (g591)) + ((!g204) & (sk[98]) & (g279) & (!g460) & (g470) & (!g591)) + ((!g204) & (sk[98]) & (g279) & (!g460) & (g470) & (g591)) + ((!g204) & (sk[98]) & (g279) & (g460) & (!g470) & (!g591)) + ((!g204) & (sk[98]) & (g279) & (g460) & (!g470) & (g591)) + ((!g204) & (sk[98]) & (g279) & (g460) & (g470) & (!g591)) + ((!g204) & (sk[98]) & (g279) & (g460) & (g470) & (g591)) + ((g204) & (!sk[98]) & (!g279) & (!g460) & (!g470) & (!g591)) + ((g204) & (!sk[98]) & (!g279) & (!g460) & (!g470) & (g591)) + ((g204) & (!sk[98]) & (!g279) & (!g460) & (g470) & (!g591)) + ((g204) & (!sk[98]) & (!g279) & (!g460) & (g470) & (g591)) + ((g204) & (!sk[98]) & (!g279) & (g460) & (!g470) & (!g591)) + ((g204) & (!sk[98]) & (!g279) & (g460) & (!g470) & (g591)) + ((g204) & (!sk[98]) & (!g279) & (g460) & (g470) & (!g591)) + ((g204) & (!sk[98]) & (!g279) & (g460) & (g470) & (g591)) + ((g204) & (!sk[98]) & (g279) & (!g460) & (!g470) & (!g591)) + ((g204) & (!sk[98]) & (g279) & (!g460) & (!g470) & (g591)) + ((g204) & (!sk[98]) & (g279) & (!g460) & (g470) & (!g591)) + ((g204) & (!sk[98]) & (g279) & (!g460) & (g470) & (g591)) + ((g204) & (!sk[98]) & (g279) & (g460) & (!g470) & (!g591)) + ((g204) & (!sk[98]) & (g279) & (g460) & (!g470) & (g591)) + ((g204) & (!sk[98]) & (g279) & (g460) & (g470) & (!g591)) + ((g204) & (!sk[98]) & (g279) & (g460) & (g470) & (g591)) + ((g204) & (sk[98]) & (!g279) & (!g460) & (!g470) & (g591)) + ((g204) & (sk[98]) & (!g279) & (!g460) & (g470) & (!g591)) + ((g204) & (sk[98]) & (!g279) & (!g460) & (g470) & (g591)) + ((g204) & (sk[98]) & (!g279) & (g460) & (!g470) & (!g591)) + ((g204) & (sk[98]) & (!g279) & (g460) & (!g470) & (g591)) + ((g204) & (sk[98]) & (!g279) & (g460) & (g470) & (!g591)) + ((g204) & (sk[98]) & (!g279) & (g460) & (g470) & (g591)) + ((g204) & (sk[98]) & (g279) & (!g460) & (!g470) & (!g591)) + ((g204) & (sk[98]) & (g279) & (!g460) & (!g470) & (g591)) + ((g204) & (sk[98]) & (g279) & (!g460) & (g470) & (!g591)) + ((g204) & (sk[98]) & (g279) & (!g460) & (g470) & (g591)) + ((g204) & (sk[98]) & (g279) & (g460) & (!g470) & (!g591)) + ((g204) & (sk[98]) & (g279) & (g460) & (!g470) & (g591)) + ((g204) & (sk[98]) & (g279) & (g460) & (g470) & (!g591)) + ((g204) & (sk[98]) & (g279) & (g460) & (g470) & (g591)));
	assign g593 = (((!g177) & (!g560) & (sk[99]) & (!g561)) + ((g177) & (!g560) & (!sk[99]) & (!g561)) + ((g177) & (!g560) & (!sk[99]) & (g561)) + ((g177) & (g560) & (!sk[99]) & (!g561)) + ((g177) & (g560) & (!sk[99]) & (g561)));
	assign g594 = (((g464) & (!sk[100]) & (!g593)) + ((g464) & (!sk[100]) & (g593)) + ((g464) & (sk[100]) & (g593)));
	assign g595 = (((!g112) & (!g136) & (!g151) & (!g548) & (!g478) & (!g594)) + ((!g112) & (!g136) & (!g151) & (!g548) & (!g478) & (g594)) + ((!g112) & (!g136) & (!g151) & (!g548) & (g478) & (!g594)) + ((!g112) & (!g136) & (!g151) & (!g548) & (g478) & (g594)) + ((!g112) & (!g136) & (!g151) & (g548) & (!g478) & (!g594)) + ((!g112) & (!g136) & (!g151) & (g548) & (!g478) & (g594)) + ((!g112) & (!g136) & (!g151) & (g548) & (g478) & (!g594)) + ((!g112) & (!g136) & (!g151) & (g548) & (g478) & (g594)) + ((!g112) & (!g136) & (g151) & (!g548) & (!g478) & (g594)) + ((!g112) & (g136) & (!g151) & (!g548) & (!g478) & (!g594)) + ((!g112) & (g136) & (!g151) & (!g548) & (!g478) & (g594)) + ((!g112) & (g136) & (!g151) & (!g548) & (g478) & (!g594)) + ((!g112) & (g136) & (!g151) & (!g548) & (g478) & (g594)) + ((!g112) & (g136) & (g151) & (!g548) & (!g478) & (g594)) + ((g112) & (!g136) & (!g151) & (!g548) & (!g478) & (!g594)) + ((g112) & (!g136) & (!g151) & (!g548) & (!g478) & (g594)) + ((g112) & (!g136) & (!g151) & (!g548) & (g478) & (!g594)) + ((g112) & (!g136) & (!g151) & (!g548) & (g478) & (g594)) + ((g112) & (!g136) & (g151) & (!g548) & (!g478) & (g594)) + ((g112) & (g136) & (!g151) & (!g548) & (!g478) & (!g594)) + ((g112) & (g136) & (!g151) & (!g548) & (!g478) & (g594)) + ((g112) & (g136) & (!g151) & (!g548) & (g478) & (!g594)) + ((g112) & (g136) & (!g151) & (!g548) & (g478) & (g594)) + ((g112) & (g136) & (g151) & (!g548) & (!g478) & (g594)));
	assign g596 = (((!i_8_) & (!sk[102]) & (!g108) & (!g177) & (!g560) & (g464)) + ((!i_8_) & (!sk[102]) & (!g108) & (!g177) & (g560) & (g464)) + ((!i_8_) & (!sk[102]) & (!g108) & (g177) & (!g560) & (g464)) + ((!i_8_) & (!sk[102]) & (!g108) & (g177) & (g560) & (g464)) + ((!i_8_) & (!sk[102]) & (g108) & (!g177) & (!g560) & (g464)) + ((!i_8_) & (!sk[102]) & (g108) & (!g177) & (g560) & (g464)) + ((!i_8_) & (!sk[102]) & (g108) & (g177) & (!g560) & (g464)) + ((!i_8_) & (!sk[102]) & (g108) & (g177) & (g560) & (g464)) + ((i_8_) & (!sk[102]) & (!g108) & (!g177) & (!g560) & (!g464)) + ((i_8_) & (!sk[102]) & (!g108) & (!g177) & (!g560) & (g464)) + ((i_8_) & (!sk[102]) & (!g108) & (!g177) & (g560) & (!g464)) + ((i_8_) & (!sk[102]) & (!g108) & (!g177) & (g560) & (g464)) + ((i_8_) & (!sk[102]) & (!g108) & (g177) & (!g560) & (!g464)) + ((i_8_) & (!sk[102]) & (!g108) & (g177) & (!g560) & (g464)) + ((i_8_) & (!sk[102]) & (!g108) & (g177) & (g560) & (!g464)) + ((i_8_) & (!sk[102]) & (!g108) & (g177) & (g560) & (g464)) + ((i_8_) & (!sk[102]) & (g108) & (!g177) & (!g560) & (!g464)) + ((i_8_) & (!sk[102]) & (g108) & (!g177) & (!g560) & (g464)) + ((i_8_) & (!sk[102]) & (g108) & (!g177) & (g560) & (!g464)) + ((i_8_) & (!sk[102]) & (g108) & (!g177) & (g560) & (g464)) + ((i_8_) & (!sk[102]) & (g108) & (g177) & (!g560) & (!g464)) + ((i_8_) & (!sk[102]) & (g108) & (g177) & (!g560) & (g464)) + ((i_8_) & (!sk[102]) & (g108) & (g177) & (g560) & (!g464)) + ((i_8_) & (!sk[102]) & (g108) & (g177) & (g560) & (g464)) + ((i_8_) & (sk[102]) & (g108) & (!g177) & (!g560) & (!g464)) + ((i_8_) & (sk[102]) & (g108) & (!g177) & (g560) & (!g464)) + ((i_8_) & (sk[102]) & (g108) & (!g177) & (g560) & (g464)) + ((i_8_) & (sk[102]) & (g108) & (g177) & (!g560) & (!g464)) + ((i_8_) & (sk[102]) & (g108) & (g177) & (!g560) & (g464)) + ((i_8_) & (sk[102]) & (g108) & (g177) & (g560) & (!g464)) + ((i_8_) & (sk[102]) & (g108) & (g177) & (g560) & (g464)));
	assign g597 = (((!g145) & (!g195) & (!g532) & (!g596) & (!sk[103]) & (g478)) + ((!g145) & (!g195) & (!g532) & (!g596) & (sk[103]) & (!g478)) + ((!g145) & (!g195) & (!g532) & (!g596) & (sk[103]) & (g478)) + ((!g145) & (!g195) & (!g532) & (g596) & (!sk[103]) & (g478)) + ((!g145) & (!g195) & (g532) & (!g596) & (!sk[103]) & (g478)) + ((!g145) & (!g195) & (g532) & (!g596) & (sk[103]) & (!g478)) + ((!g145) & (!g195) & (g532) & (!g596) & (sk[103]) & (g478)) + ((!g145) & (!g195) & (g532) & (g596) & (!sk[103]) & (g478)) + ((!g145) & (g195) & (!g532) & (!g596) & (!sk[103]) & (g478)) + ((!g145) & (g195) & (!g532) & (!g596) & (sk[103]) & (!g478)) + ((!g145) & (g195) & (!g532) & (!g596) & (sk[103]) & (g478)) + ((!g145) & (g195) & (!g532) & (g596) & (!sk[103]) & (g478)) + ((!g145) & (g195) & (g532) & (!g596) & (!sk[103]) & (g478)) + ((!g145) & (g195) & (g532) & (!g596) & (sk[103]) & (!g478)) + ((!g145) & (g195) & (g532) & (!g596) & (sk[103]) & (g478)) + ((!g145) & (g195) & (g532) & (g596) & (!sk[103]) & (g478)) + ((g145) & (!g195) & (!g532) & (!g596) & (!sk[103]) & (!g478)) + ((g145) & (!g195) & (!g532) & (!g596) & (!sk[103]) & (g478)) + ((g145) & (!g195) & (!g532) & (!g596) & (sk[103]) & (!g478)) + ((g145) & (!g195) & (!g532) & (g596) & (!sk[103]) & (!g478)) + ((g145) & (!g195) & (!g532) & (g596) & (!sk[103]) & (g478)) + ((g145) & (!g195) & (g532) & (!g596) & (!sk[103]) & (!g478)) + ((g145) & (!g195) & (g532) & (!g596) & (!sk[103]) & (g478)) + ((g145) & (!g195) & (g532) & (g596) & (!sk[103]) & (!g478)) + ((g145) & (!g195) & (g532) & (g596) & (!sk[103]) & (g478)) + ((g145) & (g195) & (!g532) & (!g596) & (!sk[103]) & (!g478)) + ((g145) & (g195) & (!g532) & (!g596) & (!sk[103]) & (g478)) + ((g145) & (g195) & (!g532) & (g596) & (!sk[103]) & (!g478)) + ((g145) & (g195) & (!g532) & (g596) & (!sk[103]) & (g478)) + ((g145) & (g195) & (g532) & (!g596) & (!sk[103]) & (!g478)) + ((g145) & (g195) & (g532) & (!g596) & (!sk[103]) & (g478)) + ((g145) & (g195) & (g532) & (g596) & (!sk[103]) & (!g478)) + ((g145) & (g195) & (g532) & (g596) & (!sk[103]) & (g478)));
	assign g598 = (((!g99) & (!g203) & (g555) & (!sk[104]) & (g474)) + ((!g99) & (g203) & (!g555) & (!sk[104]) & (!g474)) + ((!g99) & (g203) & (!g555) & (!sk[104]) & (g474)) + ((!g99) & (g203) & (g555) & (!sk[104]) & (!g474)) + ((!g99) & (g203) & (g555) & (!sk[104]) & (g474)) + ((g99) & (!g203) & (!g555) & (sk[104]) & (g474)) + ((g99) & (!g203) & (g555) & (!sk[104]) & (!g474)) + ((g99) & (!g203) & (g555) & (!sk[104]) & (g474)) + ((g99) & (!g203) & (g555) & (sk[104]) & (!g474)) + ((g99) & (!g203) & (g555) & (sk[104]) & (g474)) + ((g99) & (g203) & (!g555) & (!sk[104]) & (!g474)) + ((g99) & (g203) & (!g555) & (!sk[104]) & (g474)) + ((g99) & (g203) & (!g555) & (sk[104]) & (!g474)) + ((g99) & (g203) & (!g555) & (sk[104]) & (g474)) + ((g99) & (g203) & (g555) & (!sk[104]) & (!g474)) + ((g99) & (g203) & (g555) & (!sk[104]) & (g474)) + ((g99) & (g203) & (g555) & (sk[104]) & (!g474)) + ((g99) & (g203) & (g555) & (sk[104]) & (g474)));
	assign g599 = (((!g100) & (sk[105]) & (g284) & (g470)) + ((g100) & (!sk[105]) & (!g284) & (!g470)) + ((g100) & (!sk[105]) & (!g284) & (g470)) + ((g100) & (!sk[105]) & (g284) & (!g470)) + ((g100) & (!sk[105]) & (g284) & (g470)) + ((g100) & (sk[105]) & (!g284) & (g470)) + ((g100) & (sk[105]) & (g284) & (g470)));
	assign g600 = (((!i_8_) & (!g4) & (!g98) & (!g279) & (!sk[106]) & (g173)) + ((!i_8_) & (!g4) & (!g98) & (g279) & (!sk[106]) & (g173)) + ((!i_8_) & (!g4) & (g98) & (!g279) & (!sk[106]) & (g173)) + ((!i_8_) & (!g4) & (g98) & (g279) & (!sk[106]) & (g173)) + ((!i_8_) & (g4) & (!g98) & (!g279) & (!sk[106]) & (g173)) + ((!i_8_) & (g4) & (!g98) & (g279) & (!sk[106]) & (g173)) + ((!i_8_) & (g4) & (g98) & (!g279) & (!sk[106]) & (g173)) + ((!i_8_) & (g4) & (g98) & (g279) & (!sk[106]) & (g173)) + ((!i_8_) & (g4) & (g98) & (g279) & (sk[106]) & (!g173)) + ((!i_8_) & (g4) & (g98) & (g279) & (sk[106]) & (g173)) + ((i_8_) & (!g4) & (!g98) & (!g279) & (!sk[106]) & (!g173)) + ((i_8_) & (!g4) & (!g98) & (!g279) & (!sk[106]) & (g173)) + ((i_8_) & (!g4) & (!g98) & (g279) & (!sk[106]) & (!g173)) + ((i_8_) & (!g4) & (!g98) & (g279) & (!sk[106]) & (g173)) + ((i_8_) & (!g4) & (g98) & (!g279) & (!sk[106]) & (!g173)) + ((i_8_) & (!g4) & (g98) & (!g279) & (!sk[106]) & (g173)) + ((i_8_) & (!g4) & (g98) & (g279) & (!sk[106]) & (!g173)) + ((i_8_) & (!g4) & (g98) & (g279) & (!sk[106]) & (g173)) + ((i_8_) & (g4) & (!g98) & (!g279) & (!sk[106]) & (!g173)) + ((i_8_) & (g4) & (!g98) & (!g279) & (!sk[106]) & (g173)) + ((i_8_) & (g4) & (!g98) & (g279) & (!sk[106]) & (!g173)) + ((i_8_) & (g4) & (!g98) & (g279) & (!sk[106]) & (g173)) + ((i_8_) & (g4) & (g98) & (!g279) & (!sk[106]) & (!g173)) + ((i_8_) & (g4) & (g98) & (!g279) & (!sk[106]) & (g173)) + ((i_8_) & (g4) & (g98) & (!g279) & (sk[106]) & (g173)) + ((i_8_) & (g4) & (g98) & (g279) & (!sk[106]) & (!g173)) + ((i_8_) & (g4) & (g98) & (g279) & (!sk[106]) & (g173)) + ((i_8_) & (g4) & (g98) & (g279) & (sk[106]) & (g173)));
	assign g601 = (((i_11_) & (!i_9_) & (!sk[107]) & (!g236)) + ((i_11_) & (!i_9_) & (!sk[107]) & (g236)) + ((i_11_) & (i_9_) & (!sk[107]) & (!g236)) + ((i_11_) & (i_9_) & (!sk[107]) & (g236)) + ((i_11_) & (i_9_) & (sk[107]) & (g236)));
	assign g602 = (((!sk[108]) & (!g134) & (!g149) & (g534) & (g522)) + ((!sk[108]) & (!g134) & (g149) & (!g534) & (!g522)) + ((!sk[108]) & (!g134) & (g149) & (!g534) & (g522)) + ((!sk[108]) & (!g134) & (g149) & (g534) & (!g522)) + ((!sk[108]) & (!g134) & (g149) & (g534) & (g522)) + ((!sk[108]) & (g134) & (!g149) & (g534) & (!g522)) + ((!sk[108]) & (g134) & (!g149) & (g534) & (g522)) + ((!sk[108]) & (g134) & (g149) & (!g534) & (!g522)) + ((!sk[108]) & (g134) & (g149) & (!g534) & (g522)) + ((!sk[108]) & (g134) & (g149) & (g534) & (!g522)) + ((!sk[108]) & (g134) & (g149) & (g534) & (g522)) + ((sk[108]) & (!g134) & (g149) & (!g534) & (g522)) + ((sk[108]) & (!g134) & (g149) & (g534) & (g522)) + ((sk[108]) & (g134) & (!g149) & (g534) & (!g522)) + ((sk[108]) & (g134) & (!g149) & (g534) & (g522)) + ((sk[108]) & (g134) & (g149) & (!g534) & (g522)) + ((sk[108]) & (g134) & (g149) & (g534) & (!g522)) + ((sk[108]) & (g134) & (g149) & (g534) & (g522)));
	assign g603 = (((!sk[109]) & (!i_8_) & (!g100) & (g199) & (g531)) + ((!sk[109]) & (!i_8_) & (g100) & (!g199) & (!g531)) + ((!sk[109]) & (!i_8_) & (g100) & (!g199) & (g531)) + ((!sk[109]) & (!i_8_) & (g100) & (g199) & (!g531)) + ((!sk[109]) & (!i_8_) & (g100) & (g199) & (g531)) + ((!sk[109]) & (i_8_) & (!g100) & (g199) & (!g531)) + ((!sk[109]) & (i_8_) & (!g100) & (g199) & (g531)) + ((!sk[109]) & (i_8_) & (g100) & (!g199) & (!g531)) + ((!sk[109]) & (i_8_) & (g100) & (!g199) & (g531)) + ((!sk[109]) & (i_8_) & (g100) & (g199) & (!g531)) + ((!sk[109]) & (i_8_) & (g100) & (g199) & (g531)) + ((sk[109]) & (i_8_) & (g100) & (!g199) & (g531)) + ((sk[109]) & (i_8_) & (g100) & (g199) & (!g531)) + ((sk[109]) & (i_8_) & (g100) & (g199) & (g531)));
	assign g604 = (((!g598) & (!g599) & (!g600) & (!g601) & (!g602) & (!g603)));
	assign g605 = (((!i_8_) & (!g108) & (!g177) & (!sk[111]) & (!g560) & (g464)) + ((!i_8_) & (!g108) & (!g177) & (!sk[111]) & (g560) & (g464)) + ((!i_8_) & (!g108) & (g177) & (!sk[111]) & (!g560) & (g464)) + ((!i_8_) & (!g108) & (g177) & (!sk[111]) & (g560) & (g464)) + ((!i_8_) & (g108) & (!g177) & (!sk[111]) & (!g560) & (g464)) + ((!i_8_) & (g108) & (!g177) & (!sk[111]) & (g560) & (g464)) + ((!i_8_) & (g108) & (!g177) & (sk[111]) & (!g560) & (!g464)) + ((!i_8_) & (g108) & (!g177) & (sk[111]) & (g560) & (!g464)) + ((!i_8_) & (g108) & (!g177) & (sk[111]) & (g560) & (g464)) + ((!i_8_) & (g108) & (g177) & (!sk[111]) & (!g560) & (g464)) + ((!i_8_) & (g108) & (g177) & (!sk[111]) & (g560) & (g464)) + ((!i_8_) & (g108) & (g177) & (sk[111]) & (!g560) & (!g464)) + ((!i_8_) & (g108) & (g177) & (sk[111]) & (!g560) & (g464)) + ((!i_8_) & (g108) & (g177) & (sk[111]) & (g560) & (!g464)) + ((!i_8_) & (g108) & (g177) & (sk[111]) & (g560) & (g464)) + ((i_8_) & (!g108) & (!g177) & (!sk[111]) & (!g560) & (!g464)) + ((i_8_) & (!g108) & (!g177) & (!sk[111]) & (!g560) & (g464)) + ((i_8_) & (!g108) & (!g177) & (!sk[111]) & (g560) & (!g464)) + ((i_8_) & (!g108) & (!g177) & (!sk[111]) & (g560) & (g464)) + ((i_8_) & (!g108) & (g177) & (!sk[111]) & (!g560) & (!g464)) + ((i_8_) & (!g108) & (g177) & (!sk[111]) & (!g560) & (g464)) + ((i_8_) & (!g108) & (g177) & (!sk[111]) & (g560) & (!g464)) + ((i_8_) & (!g108) & (g177) & (!sk[111]) & (g560) & (g464)) + ((i_8_) & (g108) & (!g177) & (!sk[111]) & (!g560) & (!g464)) + ((i_8_) & (g108) & (!g177) & (!sk[111]) & (!g560) & (g464)) + ((i_8_) & (g108) & (!g177) & (!sk[111]) & (g560) & (!g464)) + ((i_8_) & (g108) & (!g177) & (!sk[111]) & (g560) & (g464)) + ((i_8_) & (g108) & (g177) & (!sk[111]) & (!g560) & (!g464)) + ((i_8_) & (g108) & (g177) & (!sk[111]) & (!g560) & (g464)) + ((i_8_) & (g108) & (g177) & (!sk[111]) & (g560) & (!g464)) + ((i_8_) & (g108) & (g177) & (!sk[111]) & (g560) & (g464)));
	assign g606 = (((!g109) & (!sk[112]) & (!g195) & (!g605) & (!g532) & (g478)) + ((!g109) & (!sk[112]) & (!g195) & (!g605) & (g532) & (g478)) + ((!g109) & (!sk[112]) & (!g195) & (g605) & (!g532) & (g478)) + ((!g109) & (!sk[112]) & (!g195) & (g605) & (g532) & (g478)) + ((!g109) & (!sk[112]) & (g195) & (!g605) & (!g532) & (g478)) + ((!g109) & (!sk[112]) & (g195) & (!g605) & (g532) & (g478)) + ((!g109) & (!sk[112]) & (g195) & (g605) & (!g532) & (g478)) + ((!g109) & (!sk[112]) & (g195) & (g605) & (g532) & (g478)) + ((!g109) & (sk[112]) & (!g195) & (!g605) & (!g532) & (!g478)) + ((!g109) & (sk[112]) & (!g195) & (!g605) & (!g532) & (g478)) + ((!g109) & (sk[112]) & (!g195) & (!g605) & (g532) & (!g478)) + ((!g109) & (sk[112]) & (!g195) & (!g605) & (g532) & (g478)) + ((!g109) & (sk[112]) & (g195) & (!g605) & (!g532) & (!g478)) + ((!g109) & (sk[112]) & (g195) & (!g605) & (!g532) & (g478)) + ((!g109) & (sk[112]) & (g195) & (!g605) & (g532) & (!g478)) + ((!g109) & (sk[112]) & (g195) & (!g605) & (g532) & (g478)) + ((g109) & (!sk[112]) & (!g195) & (!g605) & (!g532) & (!g478)) + ((g109) & (!sk[112]) & (!g195) & (!g605) & (!g532) & (g478)) + ((g109) & (!sk[112]) & (!g195) & (!g605) & (g532) & (!g478)) + ((g109) & (!sk[112]) & (!g195) & (!g605) & (g532) & (g478)) + ((g109) & (!sk[112]) & (!g195) & (g605) & (!g532) & (!g478)) + ((g109) & (!sk[112]) & (!g195) & (g605) & (!g532) & (g478)) + ((g109) & (!sk[112]) & (!g195) & (g605) & (g532) & (!g478)) + ((g109) & (!sk[112]) & (!g195) & (g605) & (g532) & (g478)) + ((g109) & (!sk[112]) & (g195) & (!g605) & (!g532) & (!g478)) + ((g109) & (!sk[112]) & (g195) & (!g605) & (!g532) & (g478)) + ((g109) & (!sk[112]) & (g195) & (!g605) & (g532) & (!g478)) + ((g109) & (!sk[112]) & (g195) & (!g605) & (g532) & (g478)) + ((g109) & (!sk[112]) & (g195) & (g605) & (!g532) & (!g478)) + ((g109) & (!sk[112]) & (g195) & (g605) & (!g532) & (g478)) + ((g109) & (!sk[112]) & (g195) & (g605) & (g532) & (!g478)) + ((g109) & (!sk[112]) & (g195) & (g605) & (g532) & (g478)) + ((g109) & (sk[112]) & (!g195) & (!g605) & (!g532) & (!g478)));
	assign g607 = (((g589) & (!g1695) & (g595) & (g597) & (g604) & (g606)));
	assign g608 = (((!g136) & (!sk[114]) & (!g199) & (g547) & (g481)) + ((!g136) & (!sk[114]) & (g199) & (!g547) & (!g481)) + ((!g136) & (!sk[114]) & (g199) & (!g547) & (g481)) + ((!g136) & (!sk[114]) & (g199) & (g547) & (!g481)) + ((!g136) & (!sk[114]) & (g199) & (g547) & (g481)) + ((g136) & (!sk[114]) & (!g199) & (g547) & (!g481)) + ((g136) & (!sk[114]) & (!g199) & (g547) & (g481)) + ((g136) & (!sk[114]) & (g199) & (!g547) & (!g481)) + ((g136) & (!sk[114]) & (g199) & (!g547) & (g481)) + ((g136) & (!sk[114]) & (g199) & (g547) & (!g481)) + ((g136) & (!sk[114]) & (g199) & (g547) & (g481)) + ((g136) & (sk[114]) & (!g199) & (!g547) & (!g481)) + ((g136) & (sk[114]) & (!g199) & (!g547) & (g481)) + ((g136) & (sk[114]) & (!g199) & (g547) & (!g481)) + ((g136) & (sk[114]) & (g199) & (!g547) & (!g481)) + ((g136) & (sk[114]) & (g199) & (!g547) & (g481)) + ((g136) & (sk[114]) & (g199) & (g547) & (!g481)) + ((g136) & (sk[114]) & (g199) & (g547) & (g481)));
	assign g609 = (((!i_8_) & (!sk[115]) & (!g108) & (!g135) & (!g561) & (g544)) + ((!i_8_) & (!sk[115]) & (!g108) & (!g135) & (g561) & (g544)) + ((!i_8_) & (!sk[115]) & (!g108) & (g135) & (!g561) & (g544)) + ((!i_8_) & (!sk[115]) & (!g108) & (g135) & (g561) & (g544)) + ((!i_8_) & (!sk[115]) & (g108) & (!g135) & (!g561) & (g544)) + ((!i_8_) & (!sk[115]) & (g108) & (!g135) & (g561) & (g544)) + ((!i_8_) & (!sk[115]) & (g108) & (g135) & (!g561) & (g544)) + ((!i_8_) & (!sk[115]) & (g108) & (g135) & (g561) & (g544)) + ((i_8_) & (!sk[115]) & (!g108) & (!g135) & (!g561) & (!g544)) + ((i_8_) & (!sk[115]) & (!g108) & (!g135) & (!g561) & (g544)) + ((i_8_) & (!sk[115]) & (!g108) & (!g135) & (g561) & (!g544)) + ((i_8_) & (!sk[115]) & (!g108) & (!g135) & (g561) & (g544)) + ((i_8_) & (!sk[115]) & (!g108) & (g135) & (!g561) & (!g544)) + ((i_8_) & (!sk[115]) & (!g108) & (g135) & (!g561) & (g544)) + ((i_8_) & (!sk[115]) & (!g108) & (g135) & (g561) & (!g544)) + ((i_8_) & (!sk[115]) & (!g108) & (g135) & (g561) & (g544)) + ((i_8_) & (!sk[115]) & (g108) & (!g135) & (!g561) & (!g544)) + ((i_8_) & (!sk[115]) & (g108) & (!g135) & (!g561) & (g544)) + ((i_8_) & (!sk[115]) & (g108) & (!g135) & (g561) & (!g544)) + ((i_8_) & (!sk[115]) & (g108) & (!g135) & (g561) & (g544)) + ((i_8_) & (!sk[115]) & (g108) & (g135) & (!g561) & (!g544)) + ((i_8_) & (!sk[115]) & (g108) & (g135) & (!g561) & (g544)) + ((i_8_) & (!sk[115]) & (g108) & (g135) & (g561) & (!g544)) + ((i_8_) & (!sk[115]) & (g108) & (g135) & (g561) & (g544)) + ((i_8_) & (sk[115]) & (!g108) & (g135) & (g561) & (!g544)) + ((i_8_) & (sk[115]) & (!g108) & (g135) & (g561) & (g544)) + ((i_8_) & (sk[115]) & (g108) & (!g135) & (!g561) & (!g544)) + ((i_8_) & (sk[115]) & (g108) & (!g135) & (g561) & (!g544)) + ((i_8_) & (sk[115]) & (g108) & (g135) & (!g561) & (!g544)) + ((i_8_) & (sk[115]) & (g108) & (g135) & (g561) & (!g544)) + ((i_8_) & (sk[115]) & (g108) & (g135) & (g561) & (g544)));
	assign g610 = (((!i_11_) & (!i_15_) & (!g141) & (sk[116]) & (g461)) + ((!i_11_) & (!i_15_) & (g141) & (!sk[116]) & (g461)) + ((!i_11_) & (!i_15_) & (g141) & (sk[116]) & (g461)) + ((!i_11_) & (i_15_) & (!g141) & (!sk[116]) & (!g461)) + ((!i_11_) & (i_15_) & (!g141) & (!sk[116]) & (g461)) + ((!i_11_) & (i_15_) & (g141) & (!sk[116]) & (!g461)) + ((!i_11_) & (i_15_) & (g141) & (!sk[116]) & (g461)) + ((i_11_) & (!i_15_) & (!g141) & (sk[116]) & (g461)) + ((i_11_) & (!i_15_) & (g141) & (!sk[116]) & (!g461)) + ((i_11_) & (!i_15_) & (g141) & (!sk[116]) & (g461)) + ((i_11_) & (!i_15_) & (g141) & (sk[116]) & (g461)) + ((i_11_) & (i_15_) & (!g141) & (!sk[116]) & (!g461)) + ((i_11_) & (i_15_) & (!g141) & (!sk[116]) & (g461)) + ((i_11_) & (i_15_) & (g141) & (!sk[116]) & (!g461)) + ((i_11_) & (i_15_) & (g141) & (!sk[116]) & (g461)) + ((i_11_) & (i_15_) & (g141) & (sk[116]) & (g461)));
	assign g611 = (((!g6) & (!i_15_) & (!sk[117]) & (!g323) & (!g186) & (g610)) + ((!g6) & (!i_15_) & (!sk[117]) & (!g323) & (g186) & (g610)) + ((!g6) & (!i_15_) & (!sk[117]) & (g323) & (!g186) & (g610)) + ((!g6) & (!i_15_) & (!sk[117]) & (g323) & (g186) & (g610)) + ((!g6) & (i_15_) & (!sk[117]) & (!g323) & (!g186) & (g610)) + ((!g6) & (i_15_) & (!sk[117]) & (!g323) & (g186) & (g610)) + ((!g6) & (i_15_) & (!sk[117]) & (g323) & (!g186) & (g610)) + ((!g6) & (i_15_) & (!sk[117]) & (g323) & (g186) & (g610)) + ((!g6) & (i_15_) & (sk[117]) & (!g323) & (g186) & (g610)) + ((!g6) & (i_15_) & (sk[117]) & (g323) & (g186) & (g610)) + ((g6) & (!i_15_) & (!sk[117]) & (!g323) & (!g186) & (!g610)) + ((g6) & (!i_15_) & (!sk[117]) & (!g323) & (!g186) & (g610)) + ((g6) & (!i_15_) & (!sk[117]) & (!g323) & (g186) & (!g610)) + ((g6) & (!i_15_) & (!sk[117]) & (!g323) & (g186) & (g610)) + ((g6) & (!i_15_) & (!sk[117]) & (g323) & (!g186) & (!g610)) + ((g6) & (!i_15_) & (!sk[117]) & (g323) & (!g186) & (g610)) + ((g6) & (!i_15_) & (!sk[117]) & (g323) & (g186) & (!g610)) + ((g6) & (!i_15_) & (!sk[117]) & (g323) & (g186) & (g610)) + ((g6) & (!i_15_) & (sk[117]) & (g323) & (!g186) & (g610)) + ((g6) & (!i_15_) & (sk[117]) & (g323) & (g186) & (g610)) + ((g6) & (i_15_) & (!sk[117]) & (!g323) & (!g186) & (!g610)) + ((g6) & (i_15_) & (!sk[117]) & (!g323) & (!g186) & (g610)) + ((g6) & (i_15_) & (!sk[117]) & (!g323) & (g186) & (!g610)) + ((g6) & (i_15_) & (!sk[117]) & (!g323) & (g186) & (g610)) + ((g6) & (i_15_) & (!sk[117]) & (g323) & (!g186) & (!g610)) + ((g6) & (i_15_) & (!sk[117]) & (g323) & (!g186) & (g610)) + ((g6) & (i_15_) & (!sk[117]) & (g323) & (g186) & (!g610)) + ((g6) & (i_15_) & (!sk[117]) & (g323) & (g186) & (g610)) + ((g6) & (i_15_) & (sk[117]) & (!g323) & (g186) & (g610)) + ((g6) & (i_15_) & (sk[117]) & (g323) & (g186) & (g610)));
	assign g612 = (((!g136) & (!g532) & (!sk[118]) & (!g495) & (!g609) & (g611)) + ((!g136) & (!g532) & (!sk[118]) & (!g495) & (g609) & (g611)) + ((!g136) & (!g532) & (!sk[118]) & (g495) & (!g609) & (g611)) + ((!g136) & (!g532) & (!sk[118]) & (g495) & (g609) & (g611)) + ((!g136) & (!g532) & (sk[118]) & (!g495) & (!g609) & (!g611)) + ((!g136) & (!g532) & (sk[118]) & (g495) & (!g609) & (!g611)) + ((!g136) & (g532) & (!sk[118]) & (!g495) & (!g609) & (g611)) + ((!g136) & (g532) & (!sk[118]) & (!g495) & (g609) & (g611)) + ((!g136) & (g532) & (!sk[118]) & (g495) & (!g609) & (g611)) + ((!g136) & (g532) & (!sk[118]) & (g495) & (g609) & (g611)) + ((!g136) & (g532) & (sk[118]) & (!g495) & (!g609) & (!g611)) + ((g136) & (!g532) & (!sk[118]) & (!g495) & (!g609) & (!g611)) + ((g136) & (!g532) & (!sk[118]) & (!g495) & (!g609) & (g611)) + ((g136) & (!g532) & (!sk[118]) & (!g495) & (g609) & (!g611)) + ((g136) & (!g532) & (!sk[118]) & (!g495) & (g609) & (g611)) + ((g136) & (!g532) & (!sk[118]) & (g495) & (!g609) & (!g611)) + ((g136) & (!g532) & (!sk[118]) & (g495) & (!g609) & (g611)) + ((g136) & (!g532) & (!sk[118]) & (g495) & (g609) & (!g611)) + ((g136) & (!g532) & (!sk[118]) & (g495) & (g609) & (g611)) + ((g136) & (!g532) & (sk[118]) & (!g495) & (!g609) & (!g611)) + ((g136) & (!g532) & (sk[118]) & (g495) & (!g609) & (!g611)) + ((g136) & (g532) & (!sk[118]) & (!g495) & (!g609) & (!g611)) + ((g136) & (g532) & (!sk[118]) & (!g495) & (!g609) & (g611)) + ((g136) & (g532) & (!sk[118]) & (!g495) & (g609) & (!g611)) + ((g136) & (g532) & (!sk[118]) & (!g495) & (g609) & (g611)) + ((g136) & (g532) & (!sk[118]) & (g495) & (!g609) & (!g611)) + ((g136) & (g532) & (!sk[118]) & (g495) & (!g609) & (g611)) + ((g136) & (g532) & (!sk[118]) & (g495) & (g609) & (!g611)) + ((g136) & (g532) & (!sk[118]) & (g495) & (g609) & (g611)));
	assign g613 = (((!sk[119]) & (g199) & (!g547)) + ((!sk[119]) & (g199) & (g547)) + ((sk[119]) & (!g199) & (g547)));
	assign g614 = (((!g18) & (!g13) & (!g195) & (!sk[120]) & (!g124) & (g461)) + ((!g18) & (!g13) & (!g195) & (!sk[120]) & (g124) & (g461)) + ((!g18) & (!g13) & (!g195) & (sk[120]) & (!g124) & (!g461)) + ((!g18) & (!g13) & (!g195) & (sk[120]) & (g124) & (!g461)) + ((!g18) & (!g13) & (g195) & (!sk[120]) & (!g124) & (g461)) + ((!g18) & (!g13) & (g195) & (!sk[120]) & (g124) & (g461)) + ((!g18) & (g13) & (!g195) & (!sk[120]) & (!g124) & (g461)) + ((!g18) & (g13) & (!g195) & (!sk[120]) & (g124) & (g461)) + ((!g18) & (g13) & (!g195) & (sk[120]) & (!g124) & (!g461)) + ((!g18) & (g13) & (g195) & (!sk[120]) & (!g124) & (g461)) + ((!g18) & (g13) & (g195) & (!sk[120]) & (g124) & (g461)) + ((g18) & (!g13) & (!g195) & (!sk[120]) & (!g124) & (!g461)) + ((g18) & (!g13) & (!g195) & (!sk[120]) & (!g124) & (g461)) + ((g18) & (!g13) & (!g195) & (!sk[120]) & (g124) & (!g461)) + ((g18) & (!g13) & (!g195) & (!sk[120]) & (g124) & (g461)) + ((g18) & (!g13) & (!g195) & (sk[120]) & (!g124) & (!g461)) + ((g18) & (!g13) & (!g195) & (sk[120]) & (!g124) & (g461)) + ((g18) & (!g13) & (!g195) & (sk[120]) & (g124) & (!g461)) + ((g18) & (!g13) & (g195) & (!sk[120]) & (!g124) & (!g461)) + ((g18) & (!g13) & (g195) & (!sk[120]) & (!g124) & (g461)) + ((g18) & (!g13) & (g195) & (!sk[120]) & (g124) & (!g461)) + ((g18) & (!g13) & (g195) & (!sk[120]) & (g124) & (g461)) + ((g18) & (g13) & (!g195) & (!sk[120]) & (!g124) & (!g461)) + ((g18) & (g13) & (!g195) & (!sk[120]) & (!g124) & (g461)) + ((g18) & (g13) & (!g195) & (!sk[120]) & (g124) & (!g461)) + ((g18) & (g13) & (!g195) & (!sk[120]) & (g124) & (g461)) + ((g18) & (g13) & (!g195) & (sk[120]) & (!g124) & (!g461)) + ((g18) & (g13) & (!g195) & (sk[120]) & (!g124) & (g461)) + ((g18) & (g13) & (g195) & (!sk[120]) & (!g124) & (!g461)) + ((g18) & (g13) & (g195) & (!sk[120]) & (!g124) & (g461)) + ((g18) & (g13) & (g195) & (!sk[120]) & (g124) & (!g461)) + ((g18) & (g13) & (g195) & (!sk[120]) & (g124) & (g461)));
	assign g615 = (((!g177) & (!g560) & (!sk[121]) & (!g613) & (!g506) & (g614)) + ((!g177) & (!g560) & (!sk[121]) & (!g613) & (g506) & (g614)) + ((!g177) & (!g560) & (!sk[121]) & (g613) & (!g506) & (g614)) + ((!g177) & (!g560) & (!sk[121]) & (g613) & (g506) & (g614)) + ((!g177) & (!g560) & (sk[121]) & (g613) & (!g506) & (g614)) + ((!g177) & (g560) & (!sk[121]) & (!g613) & (!g506) & (g614)) + ((!g177) & (g560) & (!sk[121]) & (!g613) & (g506) & (g614)) + ((!g177) & (g560) & (!sk[121]) & (g613) & (!g506) & (g614)) + ((!g177) & (g560) & (!sk[121]) & (g613) & (g506) & (g614)) + ((g177) & (!g560) & (!sk[121]) & (!g613) & (!g506) & (!g614)) + ((g177) & (!g560) & (!sk[121]) & (!g613) & (!g506) & (g614)) + ((g177) & (!g560) & (!sk[121]) & (!g613) & (g506) & (!g614)) + ((g177) & (!g560) & (!sk[121]) & (!g613) & (g506) & (g614)) + ((g177) & (!g560) & (!sk[121]) & (g613) & (!g506) & (!g614)) + ((g177) & (!g560) & (!sk[121]) & (g613) & (!g506) & (g614)) + ((g177) & (!g560) & (!sk[121]) & (g613) & (g506) & (!g614)) + ((g177) & (!g560) & (!sk[121]) & (g613) & (g506) & (g614)) + ((g177) & (g560) & (!sk[121]) & (!g613) & (!g506) & (!g614)) + ((g177) & (g560) & (!sk[121]) & (!g613) & (!g506) & (g614)) + ((g177) & (g560) & (!sk[121]) & (!g613) & (g506) & (!g614)) + ((g177) & (g560) & (!sk[121]) & (!g613) & (g506) & (g614)) + ((g177) & (g560) & (!sk[121]) & (g613) & (!g506) & (!g614)) + ((g177) & (g560) & (!sk[121]) & (g613) & (!g506) & (g614)) + ((g177) & (g560) & (!sk[121]) & (g613) & (g506) & (!g614)) + ((g177) & (g560) & (!sk[121]) & (g613) & (g506) & (g614)));
	assign g616 = (((!i_11_) & (!sk[122]) & (!i_9_) & (!i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (!sk[122]) & (!i_9_) & (!i_10_) & (i_15_) & (g461)) + ((!i_11_) & (!sk[122]) & (!i_9_) & (i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (!sk[122]) & (!i_9_) & (i_10_) & (i_15_) & (g461)) + ((!i_11_) & (!sk[122]) & (i_9_) & (!i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (!sk[122]) & (i_9_) & (!i_10_) & (i_15_) & (g461)) + ((!i_11_) & (!sk[122]) & (i_9_) & (i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (!sk[122]) & (i_9_) & (i_10_) & (i_15_) & (g461)) + ((!i_11_) & (sk[122]) & (!i_9_) & (!i_10_) & (!i_15_) & (!g461)) + ((!i_11_) & (sk[122]) & (!i_9_) & (!i_10_) & (i_15_) & (!g461)) + ((!i_11_) & (sk[122]) & (!i_9_) & (!i_10_) & (i_15_) & (g461)) + ((!i_11_) & (sk[122]) & (!i_9_) & (i_10_) & (!i_15_) & (!g461)) + ((!i_11_) & (sk[122]) & (!i_9_) & (i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (sk[122]) & (!i_9_) & (i_10_) & (i_15_) & (!g461)) + ((!i_11_) & (sk[122]) & (!i_9_) & (i_10_) & (i_15_) & (g461)) + ((!i_11_) & (sk[122]) & (i_9_) & (!i_10_) & (!i_15_) & (!g461)) + ((!i_11_) & (sk[122]) & (i_9_) & (!i_10_) & (i_15_) & (!g461)) + ((!i_11_) & (sk[122]) & (i_9_) & (i_10_) & (!i_15_) & (!g461)) + ((!i_11_) & (sk[122]) & (i_9_) & (i_10_) & (!i_15_) & (g461)) + ((!i_11_) & (sk[122]) & (i_9_) & (i_10_) & (i_15_) & (!g461)) + ((!i_11_) & (sk[122]) & (i_9_) & (i_10_) & (i_15_) & (g461)) + ((i_11_) & (!sk[122]) & (!i_9_) & (!i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (!sk[122]) & (!i_9_) & (!i_10_) & (!i_15_) & (g461)) + ((i_11_) & (!sk[122]) & (!i_9_) & (!i_10_) & (i_15_) & (!g461)) + ((i_11_) & (!sk[122]) & (!i_9_) & (!i_10_) & (i_15_) & (g461)) + ((i_11_) & (!sk[122]) & (!i_9_) & (i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (!sk[122]) & (!i_9_) & (i_10_) & (!i_15_) & (g461)) + ((i_11_) & (!sk[122]) & (!i_9_) & (i_10_) & (i_15_) & (!g461)) + ((i_11_) & (!sk[122]) & (!i_9_) & (i_10_) & (i_15_) & (g461)) + ((i_11_) & (!sk[122]) & (i_9_) & (!i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (!sk[122]) & (i_9_) & (!i_10_) & (!i_15_) & (g461)) + ((i_11_) & (!sk[122]) & (i_9_) & (!i_10_) & (i_15_) & (!g461)) + ((i_11_) & (!sk[122]) & (i_9_) & (!i_10_) & (i_15_) & (g461)) + ((i_11_) & (!sk[122]) & (i_9_) & (i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (!sk[122]) & (i_9_) & (i_10_) & (!i_15_) & (g461)) + ((i_11_) & (!sk[122]) & (i_9_) & (i_10_) & (i_15_) & (!g461)) + ((i_11_) & (!sk[122]) & (i_9_) & (i_10_) & (i_15_) & (g461)) + ((i_11_) & (sk[122]) & (!i_9_) & (!i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (sk[122]) & (!i_9_) & (!i_10_) & (i_15_) & (!g461)) + ((i_11_) & (sk[122]) & (!i_9_) & (i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (sk[122]) & (!i_9_) & (i_10_) & (!i_15_) & (g461)) + ((i_11_) & (sk[122]) & (!i_9_) & (i_10_) & (i_15_) & (!g461)) + ((i_11_) & (sk[122]) & (i_9_) & (!i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (sk[122]) & (i_9_) & (!i_10_) & (!i_15_) & (g461)) + ((i_11_) & (sk[122]) & (i_9_) & (!i_10_) & (i_15_) & (!g461)) + ((i_11_) & (sk[122]) & (i_9_) & (!i_10_) & (i_15_) & (g461)) + ((i_11_) & (sk[122]) & (i_9_) & (i_10_) & (!i_15_) & (!g461)) + ((i_11_) & (sk[122]) & (i_9_) & (i_10_) & (!i_15_) & (g461)) + ((i_11_) & (sk[122]) & (i_9_) & (i_10_) & (i_15_) & (!g461)));
	assign g617 = (((!i_11_) & (!i_9_) & (!i_10_) & (!sk[123]) & (!i_15_) & (g13)) + ((!i_11_) & (!i_9_) & (!i_10_) & (!sk[123]) & (i_15_) & (g13)) + ((!i_11_) & (!i_9_) & (i_10_) & (!sk[123]) & (!i_15_) & (g13)) + ((!i_11_) & (!i_9_) & (i_10_) & (!sk[123]) & (i_15_) & (g13)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[123]) & (!i_15_) & (g13)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[123]) & (i_15_) & (g13)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[123]) & (!i_15_) & (g13)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[123]) & (i_15_) & (g13)) + ((!i_11_) & (i_9_) & (i_10_) & (sk[123]) & (i_15_) & (g13)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[123]) & (!i_15_) & (!g13)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[123]) & (!i_15_) & (g13)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[123]) & (i_15_) & (!g13)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[123]) & (i_15_) & (g13)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[123]) & (!i_15_) & (!g13)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[123]) & (!i_15_) & (g13)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[123]) & (i_15_) & (!g13)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[123]) & (i_15_) & (g13)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[123]) & (!i_15_) & (!g13)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[123]) & (!i_15_) & (g13)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[123]) & (i_15_) & (!g13)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[123]) & (i_15_) & (g13)) + ((i_11_) & (i_9_) & (!i_10_) & (sk[123]) & (i_15_) & (g13)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[123]) & (!i_15_) & (!g13)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[123]) & (!i_15_) & (g13)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[123]) & (i_15_) & (!g13)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[123]) & (i_15_) & (g13)));
	assign g618 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g99) & (!sk[124]) & (g158)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g99) & (!sk[124]) & (g158)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g99) & (!sk[124]) & (g158)) + ((!i_14_) & (!i_12_) & (i_13_) & (g99) & (!sk[124]) & (g158)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g99) & (!sk[124]) & (g158)) + ((!i_14_) & (i_12_) & (!i_13_) & (g99) & (!sk[124]) & (g158)) + ((!i_14_) & (i_12_) & (i_13_) & (!g99) & (!sk[124]) & (g158)) + ((!i_14_) & (i_12_) & (i_13_) & (g99) & (!sk[124]) & (g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g99) & (!sk[124]) & (!g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g99) & (!sk[124]) & (g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (g99) & (!sk[124]) & (!g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (g99) & (!sk[124]) & (g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (g99) & (sk[124]) & (g158)) + ((i_14_) & (!i_12_) & (i_13_) & (!g99) & (!sk[124]) & (!g158)) + ((i_14_) & (!i_12_) & (i_13_) & (!g99) & (!sk[124]) & (g158)) + ((i_14_) & (!i_12_) & (i_13_) & (g99) & (!sk[124]) & (!g158)) + ((i_14_) & (!i_12_) & (i_13_) & (g99) & (!sk[124]) & (g158)) + ((i_14_) & (!i_12_) & (i_13_) & (g99) & (sk[124]) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (!g99) & (!sk[124]) & (!g158)) + ((i_14_) & (i_12_) & (!i_13_) & (!g99) & (!sk[124]) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (g99) & (!sk[124]) & (!g158)) + ((i_14_) & (i_12_) & (!i_13_) & (g99) & (!sk[124]) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (g99) & (sk[124]) & (g158)) + ((i_14_) & (i_12_) & (i_13_) & (!g99) & (!sk[124]) & (!g158)) + ((i_14_) & (i_12_) & (i_13_) & (!g99) & (!sk[124]) & (g158)) + ((i_14_) & (i_12_) & (i_13_) & (g99) & (!sk[124]) & (!g158)) + ((i_14_) & (i_12_) & (i_13_) & (g99) & (!sk[124]) & (g158)));
	assign g619 = (((i_15_) & (!sk[125]) & (!g178) & (!g461)) + ((i_15_) & (!sk[125]) & (!g178) & (g461)) + ((i_15_) & (!sk[125]) & (g178) & (!g461)) + ((i_15_) & (!sk[125]) & (g178) & (g461)) + ((i_15_) & (sk[125]) & (g178) & (g461)));
	assign g620 = (((!sk[126]) & (g59) & (!g243) & (!g619)) + ((!sk[126]) & (g59) & (!g243) & (g619)) + ((!sk[126]) & (g59) & (g243) & (!g619)) + ((!sk[126]) & (g59) & (g243) & (g619)) + ((sk[126]) & (!g59) & (g243) & (g619)) + ((sk[126]) & (g59) & (!g243) & (g619)) + ((sk[126]) & (g59) & (g243) & (g619)));
	assign g621 = (((!sk[127]) & (g135) & (!g576)) + ((!sk[127]) & (g135) & (g576)) + ((sk[127]) & (g135) & (!g576)));
	assign g622 = (((!i_15_) & (!g113) & (!sk[0]) & (g118) & (g171)) + ((!i_15_) & (g113) & (!sk[0]) & (!g118) & (!g171)) + ((!i_15_) & (g113) & (!sk[0]) & (!g118) & (g171)) + ((!i_15_) & (g113) & (!sk[0]) & (g118) & (!g171)) + ((!i_15_) & (g113) & (!sk[0]) & (g118) & (g171)) + ((!i_15_) & (g113) & (sk[0]) & (g118) & (!g171)) + ((i_15_) & (!g113) & (!sk[0]) & (g118) & (!g171)) + ((i_15_) & (!g113) & (!sk[0]) & (g118) & (g171)) + ((i_15_) & (g113) & (!sk[0]) & (!g118) & (!g171)) + ((i_15_) & (g113) & (!sk[0]) & (!g118) & (g171)) + ((i_15_) & (g113) & (!sk[0]) & (g118) & (!g171)) + ((i_15_) & (g113) & (!sk[0]) & (g118) & (g171)));
	assign g623 = (((!g277) & (!g617) & (!g618) & (!g620) & (!g621) & (!g622)) + ((g277) & (!g617) & (!g618) & (!g620) & (!g621) & (!g622)) + ((g277) & (g617) & (!g618) & (!g620) & (!g621) & (!g622)));
	assign g624 = (((!g108) & (!g131) & (!sk[2]) & (!g171) & (!g164) & (g461)) + ((!g108) & (!g131) & (!sk[2]) & (!g171) & (g164) & (g461)) + ((!g108) & (!g131) & (!sk[2]) & (g171) & (!g164) & (g461)) + ((!g108) & (!g131) & (!sk[2]) & (g171) & (g164) & (g461)) + ((!g108) & (g131) & (!sk[2]) & (!g171) & (!g164) & (g461)) + ((!g108) & (g131) & (!sk[2]) & (!g171) & (g164) & (g461)) + ((!g108) & (g131) & (!sk[2]) & (g171) & (!g164) & (g461)) + ((!g108) & (g131) & (!sk[2]) & (g171) & (g164) & (g461)) + ((g108) & (!g131) & (!sk[2]) & (!g171) & (!g164) & (!g461)) + ((g108) & (!g131) & (!sk[2]) & (!g171) & (!g164) & (g461)) + ((g108) & (!g131) & (!sk[2]) & (!g171) & (g164) & (!g461)) + ((g108) & (!g131) & (!sk[2]) & (!g171) & (g164) & (g461)) + ((g108) & (!g131) & (!sk[2]) & (g171) & (!g164) & (!g461)) + ((g108) & (!g131) & (!sk[2]) & (g171) & (!g164) & (g461)) + ((g108) & (!g131) & (!sk[2]) & (g171) & (g164) & (!g461)) + ((g108) & (!g131) & (!sk[2]) & (g171) & (g164) & (g461)) + ((g108) & (!g131) & (sk[2]) & (!g171) & (g164) & (!g461)) + ((g108) & (!g131) & (sk[2]) & (!g171) & (g164) & (g461)) + ((g108) & (g131) & (!sk[2]) & (!g171) & (!g164) & (!g461)) + ((g108) & (g131) & (!sk[2]) & (!g171) & (!g164) & (g461)) + ((g108) & (g131) & (!sk[2]) & (!g171) & (g164) & (!g461)) + ((g108) & (g131) & (!sk[2]) & (!g171) & (g164) & (g461)) + ((g108) & (g131) & (!sk[2]) & (g171) & (!g164) & (!g461)) + ((g108) & (g131) & (!sk[2]) & (g171) & (!g164) & (g461)) + ((g108) & (g131) & (!sk[2]) & (g171) & (g164) & (!g461)) + ((g108) & (g131) & (!sk[2]) & (g171) & (g164) & (g461)) + ((g108) & (g131) & (sk[2]) & (!g171) & (!g164) & (g461)) + ((g108) & (g131) & (sk[2]) & (!g171) & (g164) & (!g461)) + ((g108) & (g131) & (sk[2]) & (!g171) & (g164) & (g461)) + ((g108) & (g131) & (sk[2]) & (g171) & (!g164) & (g461)) + ((g108) & (g131) & (sk[2]) & (g171) & (g164) & (g461)));
	assign g625 = (((!g47) & (!g566) & (!g546) & (sk[3]) & (!g555)) + ((!g47) & (!g566) & (g546) & (!sk[3]) & (g555)) + ((!g47) & (g566) & (!g546) & (!sk[3]) & (!g555)) + ((!g47) & (g566) & (!g546) & (!sk[3]) & (g555)) + ((!g47) & (g566) & (g546) & (!sk[3]) & (!g555)) + ((!g47) & (g566) & (g546) & (!sk[3]) & (g555)) + ((g47) & (!g566) & (g546) & (!sk[3]) & (!g555)) + ((g47) & (!g566) & (g546) & (!sk[3]) & (g555)) + ((g47) & (g566) & (!g546) & (!sk[3]) & (!g555)) + ((g47) & (g566) & (!g546) & (!sk[3]) & (g555)) + ((g47) & (g566) & (g546) & (!sk[3]) & (!g555)) + ((g47) & (g566) & (g546) & (!sk[3]) & (g555)));
	assign g626 = (((!sk[4]) & (g199) & (!g547) & (!g481)) + ((!sk[4]) & (g199) & (!g547) & (g481)) + ((!sk[4]) & (g199) & (g547) & (!g481)) + ((!sk[4]) & (g199) & (g547) & (g481)) + ((sk[4]) & (!g199) & (g547) & (g481)));
	assign g627 = (((!g177) & (sk[5]) & (!g560) & (g464)) + ((g177) & (!sk[5]) & (!g560) & (!g464)) + ((g177) & (!sk[5]) & (!g560) & (g464)) + ((g177) & (!sk[5]) & (g560) & (!g464)) + ((g177) & (!sk[5]) & (g560) & (g464)));
	assign g628 = (((!i_8_) & (!g88) & (!sk[6]) & (!g108) & (!g626) & (g627)) + ((!i_8_) & (!g88) & (!sk[6]) & (!g108) & (g626) & (g627)) + ((!i_8_) & (!g88) & (!sk[6]) & (g108) & (!g626) & (g627)) + ((!i_8_) & (!g88) & (!sk[6]) & (g108) & (g626) & (g627)) + ((!i_8_) & (!g88) & (sk[6]) & (g108) & (!g626) & (!g627)) + ((!i_8_) & (!g88) & (sk[6]) & (g108) & (!g626) & (g627)) + ((!i_8_) & (g88) & (!sk[6]) & (!g108) & (!g626) & (g627)) + ((!i_8_) & (g88) & (!sk[6]) & (!g108) & (g626) & (g627)) + ((!i_8_) & (g88) & (!sk[6]) & (g108) & (!g626) & (g627)) + ((!i_8_) & (g88) & (!sk[6]) & (g108) & (g626) & (g627)) + ((!i_8_) & (g88) & (sk[6]) & (!g108) & (!g626) & (!g627)) + ((!i_8_) & (g88) & (sk[6]) & (!g108) & (!g626) & (g627)) + ((!i_8_) & (g88) & (sk[6]) & (!g108) & (g626) & (!g627)) + ((!i_8_) & (g88) & (sk[6]) & (g108) & (!g626) & (!g627)) + ((!i_8_) & (g88) & (sk[6]) & (g108) & (!g626) & (g627)) + ((!i_8_) & (g88) & (sk[6]) & (g108) & (g626) & (!g627)) + ((i_8_) & (!g88) & (!sk[6]) & (!g108) & (!g626) & (!g627)) + ((i_8_) & (!g88) & (!sk[6]) & (!g108) & (!g626) & (g627)) + ((i_8_) & (!g88) & (!sk[6]) & (!g108) & (g626) & (!g627)) + ((i_8_) & (!g88) & (!sk[6]) & (!g108) & (g626) & (g627)) + ((i_8_) & (!g88) & (!sk[6]) & (g108) & (!g626) & (!g627)) + ((i_8_) & (!g88) & (!sk[6]) & (g108) & (!g626) & (g627)) + ((i_8_) & (!g88) & (!sk[6]) & (g108) & (g626) & (!g627)) + ((i_8_) & (!g88) & (!sk[6]) & (g108) & (g626) & (g627)) + ((i_8_) & (g88) & (!sk[6]) & (!g108) & (!g626) & (!g627)) + ((i_8_) & (g88) & (!sk[6]) & (!g108) & (!g626) & (g627)) + ((i_8_) & (g88) & (!sk[6]) & (!g108) & (g626) & (!g627)) + ((i_8_) & (g88) & (!sk[6]) & (!g108) & (g626) & (g627)) + ((i_8_) & (g88) & (!sk[6]) & (g108) & (!g626) & (!g627)) + ((i_8_) & (g88) & (!sk[6]) & (g108) & (!g626) & (g627)) + ((i_8_) & (g88) & (!sk[6]) & (g108) & (g626) & (!g627)) + ((i_8_) & (g88) & (!sk[6]) & (g108) & (g626) & (g627)));
	assign g629 = (((!sk[7]) & (!g109) & (!g534) & (!g624) & (!g625) & (g628)) + ((!sk[7]) & (!g109) & (!g534) & (!g624) & (g625) & (g628)) + ((!sk[7]) & (!g109) & (!g534) & (g624) & (!g625) & (g628)) + ((!sk[7]) & (!g109) & (!g534) & (g624) & (g625) & (g628)) + ((!sk[7]) & (!g109) & (g534) & (!g624) & (!g625) & (g628)) + ((!sk[7]) & (!g109) & (g534) & (!g624) & (g625) & (g628)) + ((!sk[7]) & (!g109) & (g534) & (g624) & (!g625) & (g628)) + ((!sk[7]) & (!g109) & (g534) & (g624) & (g625) & (g628)) + ((!sk[7]) & (g109) & (!g534) & (!g624) & (!g625) & (!g628)) + ((!sk[7]) & (g109) & (!g534) & (!g624) & (!g625) & (g628)) + ((!sk[7]) & (g109) & (!g534) & (!g624) & (g625) & (!g628)) + ((!sk[7]) & (g109) & (!g534) & (!g624) & (g625) & (g628)) + ((!sk[7]) & (g109) & (!g534) & (g624) & (!g625) & (!g628)) + ((!sk[7]) & (g109) & (!g534) & (g624) & (!g625) & (g628)) + ((!sk[7]) & (g109) & (!g534) & (g624) & (g625) & (!g628)) + ((!sk[7]) & (g109) & (!g534) & (g624) & (g625) & (g628)) + ((!sk[7]) & (g109) & (g534) & (!g624) & (!g625) & (!g628)) + ((!sk[7]) & (g109) & (g534) & (!g624) & (!g625) & (g628)) + ((!sk[7]) & (g109) & (g534) & (!g624) & (g625) & (!g628)) + ((!sk[7]) & (g109) & (g534) & (!g624) & (g625) & (g628)) + ((!sk[7]) & (g109) & (g534) & (g624) & (!g625) & (!g628)) + ((!sk[7]) & (g109) & (g534) & (g624) & (!g625) & (g628)) + ((!sk[7]) & (g109) & (g534) & (g624) & (g625) & (!g628)) + ((!sk[7]) & (g109) & (g534) & (g624) & (g625) & (g628)) + ((sk[7]) & (!g109) & (!g534) & (!g624) & (!g625) & (!g628)) + ((sk[7]) & (!g109) & (!g534) & (!g624) & (g625) & (!g628)) + ((sk[7]) & (!g109) & (g534) & (!g624) & (!g625) & (!g628)) + ((sk[7]) & (!g109) & (g534) & (!g624) & (g625) & (!g628)) + ((sk[7]) & (g109) & (!g534) & (!g624) & (g625) & (!g628)));
	assign g630 = (((!sk[8]) & (g171) & (!g115)) + ((!sk[8]) & (g171) & (g115)) + ((sk[8]) & (!g171) & (!g115)));
	assign g631 = (((!g548) & (!g550) & (!g561) & (sk[9]) & (!g630)) + ((!g548) & (!g550) & (g561) & (!sk[9]) & (g630)) + ((!g548) & (g550) & (!g561) & (!sk[9]) & (!g630)) + ((!g548) & (g550) & (!g561) & (!sk[9]) & (g630)) + ((!g548) & (g550) & (g561) & (!sk[9]) & (!g630)) + ((!g548) & (g550) & (g561) & (!sk[9]) & (g630)) + ((g548) & (!g550) & (g561) & (!sk[9]) & (!g630)) + ((g548) & (!g550) & (g561) & (!sk[9]) & (g630)) + ((g548) & (g550) & (!g561) & (!sk[9]) & (!g630)) + ((g548) & (g550) & (!g561) & (!sk[9]) & (g630)) + ((g548) & (g550) & (g561) & (!sk[9]) & (!g630)) + ((g548) & (g550) & (g561) & (!sk[9]) & (g630)));
	assign g632 = (((!g134) & (!g109) & (!g146) & (!g551) & (!sk[10]) & (g631)) + ((!g134) & (!g109) & (!g146) & (!g551) & (sk[10]) & (!g631)) + ((!g134) & (!g109) & (!g146) & (!g551) & (sk[10]) & (g631)) + ((!g134) & (!g109) & (!g146) & (g551) & (!sk[10]) & (g631)) + ((!g134) & (!g109) & (g146) & (!g551) & (!sk[10]) & (g631)) + ((!g134) & (!g109) & (g146) & (!g551) & (sk[10]) & (!g631)) + ((!g134) & (!g109) & (g146) & (!g551) & (sk[10]) & (g631)) + ((!g134) & (!g109) & (g146) & (g551) & (!sk[10]) & (g631)) + ((!g134) & (!g109) & (g146) & (g551) & (sk[10]) & (!g631)) + ((!g134) & (!g109) & (g146) & (g551) & (sk[10]) & (g631)) + ((!g134) & (g109) & (!g146) & (!g551) & (!sk[10]) & (g631)) + ((!g134) & (g109) & (!g146) & (!g551) & (sk[10]) & (!g631)) + ((!g134) & (g109) & (!g146) & (!g551) & (sk[10]) & (g631)) + ((!g134) & (g109) & (!g146) & (g551) & (!sk[10]) & (g631)) + ((!g134) & (g109) & (g146) & (!g551) & (!sk[10]) & (g631)) + ((!g134) & (g109) & (g146) & (!g551) & (sk[10]) & (!g631)) + ((!g134) & (g109) & (g146) & (!g551) & (sk[10]) & (g631)) + ((!g134) & (g109) & (g146) & (g551) & (!sk[10]) & (g631)) + ((g134) & (!g109) & (!g146) & (!g551) & (!sk[10]) & (!g631)) + ((g134) & (!g109) & (!g146) & (!g551) & (!sk[10]) & (g631)) + ((g134) & (!g109) & (!g146) & (!g551) & (sk[10]) & (g631)) + ((g134) & (!g109) & (!g146) & (g551) & (!sk[10]) & (!g631)) + ((g134) & (!g109) & (!g146) & (g551) & (!sk[10]) & (g631)) + ((g134) & (!g109) & (g146) & (!g551) & (!sk[10]) & (!g631)) + ((g134) & (!g109) & (g146) & (!g551) & (!sk[10]) & (g631)) + ((g134) & (!g109) & (g146) & (!g551) & (sk[10]) & (g631)) + ((g134) & (!g109) & (g146) & (g551) & (!sk[10]) & (!g631)) + ((g134) & (!g109) & (g146) & (g551) & (!sk[10]) & (g631)) + ((g134) & (g109) & (!g146) & (!g551) & (!sk[10]) & (!g631)) + ((g134) & (g109) & (!g146) & (!g551) & (!sk[10]) & (g631)) + ((g134) & (g109) & (!g146) & (!g551) & (sk[10]) & (g631)) + ((g134) & (g109) & (!g146) & (g551) & (!sk[10]) & (!g631)) + ((g134) & (g109) & (!g146) & (g551) & (!sk[10]) & (g631)) + ((g134) & (g109) & (g146) & (!g551) & (!sk[10]) & (!g631)) + ((g134) & (g109) & (g146) & (!g551) & (!sk[10]) & (g631)) + ((g134) & (g109) & (g146) & (!g551) & (sk[10]) & (g631)) + ((g134) & (g109) & (g146) & (g551) & (!sk[10]) & (!g631)) + ((g134) & (g109) & (g146) & (g551) & (!sk[10]) & (g631)));
	assign g633 = (((!g608) & (g612) & (g1686) & (g623) & (g629) & (g632)));
	assign g634 = (((g527) & (g543) & (g568) & (g587) & (g607) & (g633)));
	assign g635 = (((!g145) & (!g268) & (g555) & (!sk[13]) & (g474)) + ((!g145) & (g268) & (!g555) & (!sk[13]) & (!g474)) + ((!g145) & (g268) & (!g555) & (!sk[13]) & (g474)) + ((!g145) & (g268) & (g555) & (!sk[13]) & (!g474)) + ((!g145) & (g268) & (g555) & (!sk[13]) & (g474)) + ((g145) & (!g268) & (!g555) & (sk[13]) & (g474)) + ((g145) & (!g268) & (g555) & (!sk[13]) & (!g474)) + ((g145) & (!g268) & (g555) & (!sk[13]) & (g474)) + ((g145) & (!g268) & (g555) & (sk[13]) & (!g474)) + ((g145) & (!g268) & (g555) & (sk[13]) & (g474)) + ((g145) & (g268) & (!g555) & (!sk[13]) & (!g474)) + ((g145) & (g268) & (!g555) & (!sk[13]) & (g474)) + ((g145) & (g268) & (!g555) & (sk[13]) & (!g474)) + ((g145) & (g268) & (!g555) & (sk[13]) & (g474)) + ((g145) & (g268) & (g555) & (!sk[13]) & (!g474)) + ((g145) & (g268) & (g555) & (!sk[13]) & (g474)) + ((g145) & (g268) & (g555) & (sk[13]) & (!g474)) + ((g145) & (g268) & (g555) & (sk[13]) & (g474)));
	assign g636 = (((!g47) & (!g172) & (sk[14]) & (g465)) + ((g47) & (!g172) & (!sk[14]) & (!g465)) + ((g47) & (!g172) & (!sk[14]) & (g465)) + ((g47) & (g172) & (!sk[14]) & (!g465)) + ((g47) & (g172) & (!sk[14]) & (g465)));
	assign g637 = (((!g101) & (!sk[15]) & (!g151) & (g530) & (g636)) + ((!g101) & (!sk[15]) & (g151) & (!g530) & (!g636)) + ((!g101) & (!sk[15]) & (g151) & (!g530) & (g636)) + ((!g101) & (!sk[15]) & (g151) & (g530) & (!g636)) + ((!g101) & (!sk[15]) & (g151) & (g530) & (g636)) + ((!g101) & (sk[15]) & (g151) & (!g530) & (!g636)) + ((!g101) & (sk[15]) & (g151) & (g530) & (!g636)) + ((g101) & (!sk[15]) & (!g151) & (g530) & (!g636)) + ((g101) & (!sk[15]) & (!g151) & (g530) & (g636)) + ((g101) & (!sk[15]) & (g151) & (!g530) & (!g636)) + ((g101) & (!sk[15]) & (g151) & (!g530) & (g636)) + ((g101) & (!sk[15]) & (g151) & (g530) & (!g636)) + ((g101) & (!sk[15]) & (g151) & (g530) & (g636)) + ((g101) & (sk[15]) & (!g151) & (g530) & (!g636)) + ((g101) & (sk[15]) & (!g151) & (g530) & (g636)) + ((g101) & (sk[15]) & (g151) & (!g530) & (!g636)) + ((g101) & (sk[15]) & (g151) & (g530) & (!g636)) + ((g101) & (sk[15]) & (g151) & (g530) & (g636)));
	assign g638 = (((!sk[16]) & (g279) & (!g566) & (!g460)) + ((!sk[16]) & (g279) & (!g566) & (g460)) + ((!sk[16]) & (g279) & (g566) & (!g460)) + ((!sk[16]) & (g279) & (g566) & (g460)) + ((sk[16]) & (!g279) & (!g566) & (!g460)));
	assign g639 = (((!g101) & (!g145) & (!g203) & (!g555) & (!g474) & (!g638)) + ((!g101) & (!g145) & (!g203) & (!g555) & (!g474) & (g638)) + ((!g101) & (!g145) & (!g203) & (!g555) & (g474) & (!g638)) + ((!g101) & (!g145) & (!g203) & (!g555) & (g474) & (g638)) + ((!g101) & (!g145) & (!g203) & (g555) & (!g474) & (!g638)) + ((!g101) & (!g145) & (!g203) & (g555) & (!g474) & (g638)) + ((!g101) & (!g145) & (!g203) & (g555) & (g474) & (!g638)) + ((!g101) & (!g145) & (!g203) & (g555) & (g474) & (g638)) + ((!g101) & (!g145) & (g203) & (!g555) & (!g474) & (!g638)) + ((!g101) & (!g145) & (g203) & (!g555) & (!g474) & (g638)) + ((!g101) & (!g145) & (g203) & (!g555) & (g474) & (!g638)) + ((!g101) & (!g145) & (g203) & (!g555) & (g474) & (g638)) + ((!g101) & (!g145) & (g203) & (g555) & (!g474) & (!g638)) + ((!g101) & (!g145) & (g203) & (g555) & (!g474) & (g638)) + ((!g101) & (!g145) & (g203) & (g555) & (g474) & (!g638)) + ((!g101) & (!g145) & (g203) & (g555) & (g474) & (g638)) + ((!g101) & (g145) & (!g203) & (!g555) & (!g474) & (g638)) + ((!g101) & (g145) & (!g203) & (!g555) & (g474) & (g638)) + ((!g101) & (g145) & (!g203) & (g555) & (!g474) & (g638)) + ((!g101) & (g145) & (!g203) & (g555) & (g474) & (g638)) + ((!g101) & (g145) & (g203) & (!g555) & (!g474) & (g638)) + ((!g101) & (g145) & (g203) & (!g555) & (g474) & (g638)) + ((!g101) & (g145) & (g203) & (g555) & (!g474) & (g638)) + ((!g101) & (g145) & (g203) & (g555) & (g474) & (g638)) + ((g101) & (!g145) & (!g203) & (!g555) & (!g474) & (!g638)) + ((g101) & (!g145) & (!g203) & (!g555) & (!g474) & (g638)) + ((g101) & (g145) & (!g203) & (!g555) & (!g474) & (g638)));
	assign g640 = (((!sk[18]) & (g173) & (!g546) & (!g477)) + ((!sk[18]) & (g173) & (!g546) & (g477)) + ((!sk[18]) & (g173) & (g546) & (!g477)) + ((!sk[18]) & (g173) & (g546) & (g477)) + ((sk[18]) & (!g173) & (!g546) & (g477)));
	assign g641 = (((!g18) & (sk[19]) & (!g171)) + ((g18) & (!sk[19]) & (!g171)) + ((g18) & (!sk[19]) & (g171)));
	assign g642 = (((!g530) & (sk[20]) & (!g641) & (!g531)) + ((g530) & (!sk[20]) & (!g641) & (!g531)) + ((g530) & (!sk[20]) & (!g641) & (g531)) + ((g530) & (!sk[20]) & (g641) & (!g531)) + ((g530) & (!sk[20]) & (g641) & (g531)));
	assign g643 = (((!g15) & (!sk[21]) & (!g102) & (g461) & (g642)) + ((!g15) & (!sk[21]) & (g102) & (!g461) & (!g642)) + ((!g15) & (!sk[21]) & (g102) & (!g461) & (g642)) + ((!g15) & (!sk[21]) & (g102) & (g461) & (!g642)) + ((!g15) & (!sk[21]) & (g102) & (g461) & (g642)) + ((!g15) & (sk[21]) & (!g102) & (!g461) & (g642)) + ((!g15) & (sk[21]) & (g102) & (!g461) & (g642)) + ((g15) & (!sk[21]) & (!g102) & (g461) & (!g642)) + ((g15) & (!sk[21]) & (!g102) & (g461) & (g642)) + ((g15) & (!sk[21]) & (g102) & (!g461) & (!g642)) + ((g15) & (!sk[21]) & (g102) & (!g461) & (g642)) + ((g15) & (!sk[21]) & (g102) & (g461) & (!g642)) + ((g15) & (!sk[21]) & (g102) & (g461) & (g642)) + ((g15) & (sk[21]) & (!g102) & (!g461) & (g642)) + ((g15) & (sk[21]) & (g102) & (!g461) & (g642)) + ((g15) & (sk[21]) & (g102) & (g461) & (g642)));
	assign g644 = (((!g145) & (!g151) & (!g640) & (!g529) & (!sk[22]) & (g643)) + ((!g145) & (!g151) & (!g640) & (!g529) & (sk[22]) & (!g643)) + ((!g145) & (!g151) & (!g640) & (!g529) & (sk[22]) & (g643)) + ((!g145) & (!g151) & (!g640) & (g529) & (!sk[22]) & (g643)) + ((!g145) & (!g151) & (!g640) & (g529) & (sk[22]) & (!g643)) + ((!g145) & (!g151) & (!g640) & (g529) & (sk[22]) & (g643)) + ((!g145) & (!g151) & (g640) & (!g529) & (!sk[22]) & (g643)) + ((!g145) & (!g151) & (g640) & (!g529) & (sk[22]) & (!g643)) + ((!g145) & (!g151) & (g640) & (!g529) & (sk[22]) & (g643)) + ((!g145) & (!g151) & (g640) & (g529) & (!sk[22]) & (g643)) + ((!g145) & (!g151) & (g640) & (g529) & (sk[22]) & (!g643)) + ((!g145) & (!g151) & (g640) & (g529) & (sk[22]) & (g643)) + ((!g145) & (g151) & (!g640) & (!g529) & (!sk[22]) & (g643)) + ((!g145) & (g151) & (!g640) & (g529) & (!sk[22]) & (g643)) + ((!g145) & (g151) & (g640) & (!g529) & (!sk[22]) & (g643)) + ((!g145) & (g151) & (g640) & (g529) & (!sk[22]) & (g643)) + ((!g145) & (g151) & (g640) & (g529) & (sk[22]) & (g643)) + ((g145) & (!g151) & (!g640) & (!g529) & (!sk[22]) & (!g643)) + ((g145) & (!g151) & (!g640) & (!g529) & (!sk[22]) & (g643)) + ((g145) & (!g151) & (!g640) & (g529) & (!sk[22]) & (!g643)) + ((g145) & (!g151) & (!g640) & (g529) & (!sk[22]) & (g643)) + ((g145) & (!g151) & (g640) & (!g529) & (!sk[22]) & (!g643)) + ((g145) & (!g151) & (g640) & (!g529) & (!sk[22]) & (g643)) + ((g145) & (!g151) & (g640) & (!g529) & (sk[22]) & (!g643)) + ((g145) & (!g151) & (g640) & (!g529) & (sk[22]) & (g643)) + ((g145) & (!g151) & (g640) & (g529) & (!sk[22]) & (!g643)) + ((g145) & (!g151) & (g640) & (g529) & (!sk[22]) & (g643)) + ((g145) & (!g151) & (g640) & (g529) & (sk[22]) & (!g643)) + ((g145) & (!g151) & (g640) & (g529) & (sk[22]) & (g643)) + ((g145) & (g151) & (!g640) & (!g529) & (!sk[22]) & (!g643)) + ((g145) & (g151) & (!g640) & (!g529) & (!sk[22]) & (g643)) + ((g145) & (g151) & (!g640) & (g529) & (!sk[22]) & (!g643)) + ((g145) & (g151) & (!g640) & (g529) & (!sk[22]) & (g643)) + ((g145) & (g151) & (g640) & (!g529) & (!sk[22]) & (!g643)) + ((g145) & (g151) & (g640) & (!g529) & (!sk[22]) & (g643)) + ((g145) & (g151) & (g640) & (g529) & (!sk[22]) & (!g643)) + ((g145) & (g151) & (g640) & (g529) & (!sk[22]) & (g643)) + ((g145) & (g151) & (g640) & (g529) & (sk[22]) & (g643)));
	assign g645 = (((!g151) & (!g268) & (!g555) & (!g474) & (!sk[23]) & (g644)) + ((!g151) & (!g268) & (!g555) & (!g474) & (sk[23]) & (g644)) + ((!g151) & (!g268) & (!g555) & (g474) & (!sk[23]) & (g644)) + ((!g151) & (!g268) & (!g555) & (g474) & (sk[23]) & (g644)) + ((!g151) & (!g268) & (g555) & (!g474) & (!sk[23]) & (g644)) + ((!g151) & (!g268) & (g555) & (!g474) & (sk[23]) & (g644)) + ((!g151) & (!g268) & (g555) & (g474) & (!sk[23]) & (g644)) + ((!g151) & (!g268) & (g555) & (g474) & (sk[23]) & (g644)) + ((!g151) & (g268) & (!g555) & (!g474) & (!sk[23]) & (g644)) + ((!g151) & (g268) & (!g555) & (!g474) & (sk[23]) & (g644)) + ((!g151) & (g268) & (!g555) & (g474) & (!sk[23]) & (g644)) + ((!g151) & (g268) & (!g555) & (g474) & (sk[23]) & (g644)) + ((!g151) & (g268) & (g555) & (!g474) & (!sk[23]) & (g644)) + ((!g151) & (g268) & (g555) & (!g474) & (sk[23]) & (g644)) + ((!g151) & (g268) & (g555) & (g474) & (!sk[23]) & (g644)) + ((!g151) & (g268) & (g555) & (g474) & (sk[23]) & (g644)) + ((g151) & (!g268) & (!g555) & (!g474) & (!sk[23]) & (!g644)) + ((g151) & (!g268) & (!g555) & (!g474) & (!sk[23]) & (g644)) + ((g151) & (!g268) & (!g555) & (!g474) & (sk[23]) & (g644)) + ((g151) & (!g268) & (!g555) & (g474) & (!sk[23]) & (!g644)) + ((g151) & (!g268) & (!g555) & (g474) & (!sk[23]) & (g644)) + ((g151) & (!g268) & (g555) & (!g474) & (!sk[23]) & (!g644)) + ((g151) & (!g268) & (g555) & (!g474) & (!sk[23]) & (g644)) + ((g151) & (!g268) & (g555) & (g474) & (!sk[23]) & (!g644)) + ((g151) & (!g268) & (g555) & (g474) & (!sk[23]) & (g644)) + ((g151) & (g268) & (!g555) & (!g474) & (!sk[23]) & (!g644)) + ((g151) & (g268) & (!g555) & (!g474) & (!sk[23]) & (g644)) + ((g151) & (g268) & (!g555) & (g474) & (!sk[23]) & (!g644)) + ((g151) & (g268) & (!g555) & (g474) & (!sk[23]) & (g644)) + ((g151) & (g268) & (g555) & (!g474) & (!sk[23]) & (!g644)) + ((g151) & (g268) & (g555) & (!g474) & (!sk[23]) & (g644)) + ((g151) & (g268) & (g555) & (g474) & (!sk[23]) & (!g644)) + ((g151) & (g268) & (g555) & (g474) & (!sk[23]) & (g644)));
	assign g646 = (((!i_8_) & (!g88) & (!g108) & (!g112) & (!g135) & (!g284)) + ((!i_8_) & (!g88) & (!g108) & (!g112) & (g135) & (!g284)) + ((!i_8_) & (!g88) & (g108) & (!g112) & (!g135) & (!g284)) + ((!i_8_) & (!g88) & (g108) & (!g112) & (g135) & (!g284)) + ((!i_8_) & (g88) & (!g108) & (!g112) & (!g135) & (!g284)) + ((!i_8_) & (g88) & (!g108) & (!g112) & (g135) & (!g284)) + ((!i_8_) & (g88) & (g108) & (!g112) & (!g135) & (!g284)) + ((!i_8_) & (g88) & (g108) & (!g112) & (g135) & (!g284)) + ((i_8_) & (!g88) & (!g108) & (!g112) & (!g135) & (!g284)));
	assign g647 = (((!sk[25]) & (g171) & (!g158) & (!g646)) + ((!sk[25]) & (g171) & (!g158) & (g646)) + ((!sk[25]) & (g171) & (g158) & (!g646)) + ((!sk[25]) & (g171) & (g158) & (g646)) + ((sk[25]) & (!g171) & (g158) & (!g646)));
	assign g648 = (((!sk[26]) & (i_14_) & (!g101) & (!g158)) + ((!sk[26]) & (i_14_) & (!g101) & (g158)) + ((!sk[26]) & (i_14_) & (g101) & (!g158)) + ((!sk[26]) & (i_14_) & (g101) & (g158)) + ((sk[26]) & (i_14_) & (g101) & (g158)));
	assign g649 = (((g101) & (!g641) & (!sk[27]) & (!g630)) + ((g101) & (!g641) & (!sk[27]) & (g630)) + ((g101) & (!g641) & (sk[27]) & (g630)) + ((g101) & (g641) & (!sk[27]) & (!g630)) + ((g101) & (g641) & (!sk[27]) & (g630)) + ((g101) & (g641) & (sk[27]) & (!g630)) + ((g101) & (g641) & (sk[27]) & (g630)));
	assign g650 = (((!i_8_) & (!g88) & (g108) & (!sk[28]) & (g534)) + ((!i_8_) & (g88) & (!g108) & (!sk[28]) & (!g534)) + ((!i_8_) & (g88) & (!g108) & (!sk[28]) & (g534)) + ((!i_8_) & (g88) & (g108) & (!sk[28]) & (!g534)) + ((!i_8_) & (g88) & (g108) & (!sk[28]) & (g534)) + ((i_8_) & (!g88) & (g108) & (!sk[28]) & (!g534)) + ((i_8_) & (!g88) & (g108) & (!sk[28]) & (g534)) + ((i_8_) & (!g88) & (g108) & (sk[28]) & (g534)) + ((i_8_) & (g88) & (!g108) & (!sk[28]) & (!g534)) + ((i_8_) & (g88) & (!g108) & (!sk[28]) & (g534)) + ((i_8_) & (g88) & (!g108) & (sk[28]) & (g534)) + ((i_8_) & (g88) & (g108) & (!sk[28]) & (!g534)) + ((i_8_) & (g88) & (g108) & (!sk[28]) & (g534)) + ((i_8_) & (g88) & (g108) & (sk[28]) & (g534)));
	assign g651 = (((!sk[29]) & (!g112) & (!g534) & (g530) & (g540)) + ((!sk[29]) & (!g112) & (g534) & (!g530) & (!g540)) + ((!sk[29]) & (!g112) & (g534) & (!g530) & (g540)) + ((!sk[29]) & (!g112) & (g534) & (g530) & (!g540)) + ((!sk[29]) & (!g112) & (g534) & (g530) & (g540)) + ((!sk[29]) & (g112) & (!g534) & (g530) & (!g540)) + ((!sk[29]) & (g112) & (!g534) & (g530) & (g540)) + ((!sk[29]) & (g112) & (g534) & (!g530) & (!g540)) + ((!sk[29]) & (g112) & (g534) & (!g530) & (g540)) + ((!sk[29]) & (g112) & (g534) & (g530) & (!g540)) + ((!sk[29]) & (g112) & (g534) & (g530) & (g540)) + ((sk[29]) & (g112) & (!g534) & (!g530) & (g540)) + ((sk[29]) & (g112) & (!g534) & (g530) & (!g540)) + ((sk[29]) & (g112) & (!g534) & (g530) & (g540)) + ((sk[29]) & (g112) & (g534) & (!g530) & (!g540)) + ((sk[29]) & (g112) & (g534) & (!g530) & (g540)) + ((sk[29]) & (g112) & (g534) & (g530) & (!g540)) + ((sk[29]) & (g112) & (g534) & (g530) & (g540)));
	assign g652 = (((i_8_) & (g135) & (!g534) & (!g530) & (!g630) & (g540)) + ((i_8_) & (g135) & (!g534) & (!g530) & (g630) & (!g540)) + ((i_8_) & (g135) & (!g534) & (!g530) & (g630) & (g540)) + ((i_8_) & (g135) & (!g534) & (g530) & (!g630) & (!g540)) + ((i_8_) & (g135) & (!g534) & (g530) & (!g630) & (g540)) + ((i_8_) & (g135) & (!g534) & (g530) & (g630) & (!g540)) + ((i_8_) & (g135) & (!g534) & (g530) & (g630) & (g540)) + ((i_8_) & (g135) & (g534) & (!g530) & (!g630) & (!g540)) + ((i_8_) & (g135) & (g534) & (!g530) & (!g630) & (g540)) + ((i_8_) & (g135) & (g534) & (!g530) & (g630) & (!g540)) + ((i_8_) & (g135) & (g534) & (!g530) & (g630) & (g540)) + ((i_8_) & (g135) & (g534) & (g530) & (!g630) & (!g540)) + ((i_8_) & (g135) & (g534) & (g530) & (!g630) & (g540)) + ((i_8_) & (g135) & (g534) & (g530) & (g630) & (!g540)) + ((i_8_) & (g135) & (g534) & (g530) & (g630) & (g540)));
	assign g653 = (((!sk[31]) & (!g145) & (!g530) & (!g531) & (!g651) & (g652)) + ((!sk[31]) & (!g145) & (!g530) & (!g531) & (g651) & (g652)) + ((!sk[31]) & (!g145) & (!g530) & (g531) & (!g651) & (g652)) + ((!sk[31]) & (!g145) & (!g530) & (g531) & (g651) & (g652)) + ((!sk[31]) & (!g145) & (g530) & (!g531) & (!g651) & (g652)) + ((!sk[31]) & (!g145) & (g530) & (!g531) & (g651) & (g652)) + ((!sk[31]) & (!g145) & (g530) & (g531) & (!g651) & (g652)) + ((!sk[31]) & (!g145) & (g530) & (g531) & (g651) & (g652)) + ((!sk[31]) & (g145) & (!g530) & (!g531) & (!g651) & (!g652)) + ((!sk[31]) & (g145) & (!g530) & (!g531) & (!g651) & (g652)) + ((!sk[31]) & (g145) & (!g530) & (!g531) & (g651) & (!g652)) + ((!sk[31]) & (g145) & (!g530) & (!g531) & (g651) & (g652)) + ((!sk[31]) & (g145) & (!g530) & (g531) & (!g651) & (!g652)) + ((!sk[31]) & (g145) & (!g530) & (g531) & (!g651) & (g652)) + ((!sk[31]) & (g145) & (!g530) & (g531) & (g651) & (!g652)) + ((!sk[31]) & (g145) & (!g530) & (g531) & (g651) & (g652)) + ((!sk[31]) & (g145) & (g530) & (!g531) & (!g651) & (!g652)) + ((!sk[31]) & (g145) & (g530) & (!g531) & (!g651) & (g652)) + ((!sk[31]) & (g145) & (g530) & (!g531) & (g651) & (!g652)) + ((!sk[31]) & (g145) & (g530) & (!g531) & (g651) & (g652)) + ((!sk[31]) & (g145) & (g530) & (g531) & (!g651) & (!g652)) + ((!sk[31]) & (g145) & (g530) & (g531) & (!g651) & (g652)) + ((!sk[31]) & (g145) & (g530) & (g531) & (g651) & (!g652)) + ((!sk[31]) & (g145) & (g530) & (g531) & (g651) & (g652)) + ((sk[31]) & (!g145) & (!g530) & (!g531) & (!g651) & (!g652)) + ((sk[31]) & (!g145) & (!g530) & (g531) & (!g651) & (!g652)) + ((sk[31]) & (!g145) & (g530) & (!g531) & (!g651) & (!g652)) + ((sk[31]) & (!g145) & (g530) & (g531) & (!g651) & (!g652)) + ((sk[31]) & (g145) & (!g530) & (!g531) & (!g651) & (!g652)));
	assign g654 = (((!g45) & (g145) & (!g197) & (!g626) & (!g467) & (!g636)) + ((!g45) & (g145) & (!g197) & (!g626) & (!g467) & (g636)) + ((!g45) & (g145) & (!g197) & (!g626) & (g467) & (!g636)) + ((!g45) & (g145) & (!g197) & (!g626) & (g467) & (g636)) + ((!g45) & (g145) & (!g197) & (g626) & (!g467) & (!g636)) + ((!g45) & (g145) & (!g197) & (g626) & (!g467) & (g636)) + ((!g45) & (g145) & (!g197) & (g626) & (g467) & (!g636)) + ((!g45) & (g145) & (g197) & (!g626) & (!g467) & (!g636)) + ((!g45) & (g145) & (g197) & (!g626) & (!g467) & (g636)) + ((!g45) & (g145) & (g197) & (!g626) & (g467) & (!g636)) + ((!g45) & (g145) & (g197) & (!g626) & (g467) & (g636)) + ((!g45) & (g145) & (g197) & (g626) & (!g467) & (!g636)) + ((!g45) & (g145) & (g197) & (g626) & (!g467) & (g636)) + ((!g45) & (g145) & (g197) & (g626) & (g467) & (!g636)) + ((!g45) & (g145) & (g197) & (g626) & (g467) & (g636)) + ((g45) & (g145) & (!g197) & (!g626) & (!g467) & (!g636)) + ((g45) & (g145) & (!g197) & (!g626) & (!g467) & (g636)) + ((g45) & (g145) & (!g197) & (!g626) & (g467) & (!g636)) + ((g45) & (g145) & (!g197) & (!g626) & (g467) & (g636)) + ((g45) & (g145) & (!g197) & (g626) & (!g467) & (!g636)) + ((g45) & (g145) & (!g197) & (g626) & (!g467) & (g636)) + ((g45) & (g145) & (!g197) & (g626) & (g467) & (!g636)) + ((g45) & (g145) & (!g197) & (g626) & (g467) & (g636)) + ((g45) & (g145) & (g197) & (!g626) & (!g467) & (!g636)) + ((g45) & (g145) & (g197) & (!g626) & (!g467) & (g636)) + ((g45) & (g145) & (g197) & (!g626) & (g467) & (!g636)) + ((g45) & (g145) & (g197) & (!g626) & (g467) & (g636)) + ((g45) & (g145) & (g197) & (g626) & (!g467) & (!g636)) + ((g45) & (g145) & (g197) & (g626) & (!g467) & (g636)) + ((g45) & (g145) & (g197) & (g626) & (g467) & (!g636)) + ((g45) & (g145) & (g197) & (g626) & (g467) & (g636)));
	assign g655 = (((!g647) & (!g648) & (!g649) & (!g650) & (g653) & (!g654)));
	assign g656 = (((!i_8_) & (!g100) & (!g323) & (!g338) & (!sk[34]) & (g540)) + ((!i_8_) & (!g100) & (!g323) & (!g338) & (sk[34]) & (g540)) + ((!i_8_) & (!g100) & (!g323) & (g338) & (!sk[34]) & (g540)) + ((!i_8_) & (!g100) & (g323) & (!g338) & (!sk[34]) & (g540)) + ((!i_8_) & (!g100) & (g323) & (!g338) & (sk[34]) & (g540)) + ((!i_8_) & (!g100) & (g323) & (g338) & (!sk[34]) & (g540)) + ((!i_8_) & (!g100) & (g323) & (g338) & (sk[34]) & (g540)) + ((!i_8_) & (g100) & (!g323) & (!g338) & (!sk[34]) & (g540)) + ((!i_8_) & (g100) & (!g323) & (!g338) & (sk[34]) & (g540)) + ((!i_8_) & (g100) & (!g323) & (g338) & (!sk[34]) & (g540)) + ((!i_8_) & (g100) & (g323) & (!g338) & (!sk[34]) & (g540)) + ((!i_8_) & (g100) & (g323) & (!g338) & (sk[34]) & (g540)) + ((!i_8_) & (g100) & (g323) & (g338) & (!sk[34]) & (g540)) + ((!i_8_) & (g100) & (g323) & (g338) & (sk[34]) & (g540)) + ((i_8_) & (!g100) & (!g323) & (!g338) & (!sk[34]) & (!g540)) + ((i_8_) & (!g100) & (!g323) & (!g338) & (!sk[34]) & (g540)) + ((i_8_) & (!g100) & (!g323) & (!g338) & (sk[34]) & (g540)) + ((i_8_) & (!g100) & (!g323) & (g338) & (!sk[34]) & (!g540)) + ((i_8_) & (!g100) & (!g323) & (g338) & (!sk[34]) & (g540)) + ((i_8_) & (!g100) & (g323) & (!g338) & (!sk[34]) & (!g540)) + ((i_8_) & (!g100) & (g323) & (!g338) & (!sk[34]) & (g540)) + ((i_8_) & (!g100) & (g323) & (!g338) & (sk[34]) & (g540)) + ((i_8_) & (!g100) & (g323) & (g338) & (!sk[34]) & (!g540)) + ((i_8_) & (!g100) & (g323) & (g338) & (!sk[34]) & (g540)) + ((i_8_) & (!g100) & (g323) & (g338) & (sk[34]) & (g540)) + ((i_8_) & (g100) & (!g323) & (!g338) & (!sk[34]) & (!g540)) + ((i_8_) & (g100) & (!g323) & (!g338) & (!sk[34]) & (g540)) + ((i_8_) & (g100) & (!g323) & (!g338) & (sk[34]) & (g540)) + ((i_8_) & (g100) & (!g323) & (g338) & (!sk[34]) & (!g540)) + ((i_8_) & (g100) & (!g323) & (g338) & (!sk[34]) & (g540)) + ((i_8_) & (g100) & (!g323) & (g338) & (sk[34]) & (g540)) + ((i_8_) & (g100) & (g323) & (!g338) & (!sk[34]) & (!g540)) + ((i_8_) & (g100) & (g323) & (!g338) & (!sk[34]) & (g540)) + ((i_8_) & (g100) & (g323) & (!g338) & (sk[34]) & (g540)) + ((i_8_) & (g100) & (g323) & (g338) & (!sk[34]) & (!g540)) + ((i_8_) & (g100) & (g323) & (g338) & (!sk[34]) & (g540)) + ((i_8_) & (g100) & (g323) & (g338) & (sk[34]) & (g540)));
	assign g657 = (((!g101) & (!sk[35]) & (!g151) & (!g534) & (!g626) & (g656)) + ((!g101) & (!sk[35]) & (!g151) & (!g534) & (g626) & (g656)) + ((!g101) & (!sk[35]) & (!g151) & (g534) & (!g626) & (g656)) + ((!g101) & (!sk[35]) & (!g151) & (g534) & (g626) & (g656)) + ((!g101) & (!sk[35]) & (g151) & (!g534) & (!g626) & (g656)) + ((!g101) & (!sk[35]) & (g151) & (!g534) & (g626) & (g656)) + ((!g101) & (!sk[35]) & (g151) & (g534) & (!g626) & (g656)) + ((!g101) & (!sk[35]) & (g151) & (g534) & (g626) & (g656)) + ((!g101) & (sk[35]) & (!g151) & (!g534) & (!g626) & (!g656)) + ((!g101) & (sk[35]) & (!g151) & (!g534) & (g626) & (!g656)) + ((!g101) & (sk[35]) & (!g151) & (g534) & (!g626) & (!g656)) + ((!g101) & (sk[35]) & (!g151) & (g534) & (g626) & (!g656)) + ((!g101) & (sk[35]) & (g151) & (!g534) & (g626) & (!g656)) + ((!g101) & (sk[35]) & (g151) & (g534) & (g626) & (!g656)) + ((g101) & (!sk[35]) & (!g151) & (!g534) & (!g626) & (!g656)) + ((g101) & (!sk[35]) & (!g151) & (!g534) & (!g626) & (g656)) + ((g101) & (!sk[35]) & (!g151) & (!g534) & (g626) & (!g656)) + ((g101) & (!sk[35]) & (!g151) & (!g534) & (g626) & (g656)) + ((g101) & (!sk[35]) & (!g151) & (g534) & (!g626) & (!g656)) + ((g101) & (!sk[35]) & (!g151) & (g534) & (!g626) & (g656)) + ((g101) & (!sk[35]) & (!g151) & (g534) & (g626) & (!g656)) + ((g101) & (!sk[35]) & (!g151) & (g534) & (g626) & (g656)) + ((g101) & (!sk[35]) & (g151) & (!g534) & (!g626) & (!g656)) + ((g101) & (!sk[35]) & (g151) & (!g534) & (!g626) & (g656)) + ((g101) & (!sk[35]) & (g151) & (!g534) & (g626) & (!g656)) + ((g101) & (!sk[35]) & (g151) & (!g534) & (g626) & (g656)) + ((g101) & (!sk[35]) & (g151) & (g534) & (!g626) & (!g656)) + ((g101) & (!sk[35]) & (g151) & (g534) & (!g626) & (g656)) + ((g101) & (!sk[35]) & (g151) & (g534) & (g626) & (!g656)) + ((g101) & (!sk[35]) & (g151) & (g534) & (g626) & (g656)) + ((g101) & (sk[35]) & (!g151) & (!g534) & (!g626) & (!g656)) + ((g101) & (sk[35]) & (!g151) & (!g534) & (g626) & (!g656)) + ((g101) & (sk[35]) & (g151) & (!g534) & (g626) & (!g656)));
	assign g658 = (((!sk[36]) & (i_11_) & (!g141) & (!g377)) + ((!sk[36]) & (i_11_) & (!g141) & (g377)) + ((!sk[36]) & (i_11_) & (g141) & (!g377)) + ((!sk[36]) & (i_11_) & (g141) & (g377)) + ((sk[36]) & (i_11_) & (g141) & (g377)));
	assign g659 = (((i_11_) & (!sk[37]) & (!g5) & (!g377)) + ((i_11_) & (!sk[37]) & (!g5) & (g377)) + ((i_11_) & (!sk[37]) & (g5) & (!g377)) + ((i_11_) & (!sk[37]) & (g5) & (g377)) + ((i_11_) & (sk[37]) & (g5) & (g377)));
	assign g660 = (((!i_3_) & (!i_4_) & (!i_8_) & (!g34) & (!sk[38]) & (g57)) + ((!i_3_) & (!i_4_) & (!i_8_) & (g34) & (!sk[38]) & (g57)) + ((!i_3_) & (!i_4_) & (i_8_) & (!g34) & (!sk[38]) & (g57)) + ((!i_3_) & (!i_4_) & (i_8_) & (g34) & (!sk[38]) & (g57)) + ((!i_3_) & (i_4_) & (!i_8_) & (!g34) & (!sk[38]) & (g57)) + ((!i_3_) & (i_4_) & (!i_8_) & (g34) & (!sk[38]) & (g57)) + ((!i_3_) & (i_4_) & (i_8_) & (!g34) & (!sk[38]) & (g57)) + ((!i_3_) & (i_4_) & (i_8_) & (g34) & (!sk[38]) & (g57)) + ((!i_3_) & (i_4_) & (i_8_) & (g34) & (sk[38]) & (g57)) + ((i_3_) & (!i_4_) & (!i_8_) & (!g34) & (!sk[38]) & (!g57)) + ((i_3_) & (!i_4_) & (!i_8_) & (!g34) & (!sk[38]) & (g57)) + ((i_3_) & (!i_4_) & (!i_8_) & (g34) & (!sk[38]) & (!g57)) + ((i_3_) & (!i_4_) & (!i_8_) & (g34) & (!sk[38]) & (g57)) + ((i_3_) & (!i_4_) & (i_8_) & (!g34) & (!sk[38]) & (!g57)) + ((i_3_) & (!i_4_) & (i_8_) & (!g34) & (!sk[38]) & (g57)) + ((i_3_) & (!i_4_) & (i_8_) & (g34) & (!sk[38]) & (!g57)) + ((i_3_) & (!i_4_) & (i_8_) & (g34) & (!sk[38]) & (g57)) + ((i_3_) & (i_4_) & (!i_8_) & (!g34) & (!sk[38]) & (!g57)) + ((i_3_) & (i_4_) & (!i_8_) & (!g34) & (!sk[38]) & (g57)) + ((i_3_) & (i_4_) & (!i_8_) & (g34) & (!sk[38]) & (!g57)) + ((i_3_) & (i_4_) & (!i_8_) & (g34) & (!sk[38]) & (g57)) + ((i_3_) & (i_4_) & (i_8_) & (!g34) & (!sk[38]) & (!g57)) + ((i_3_) & (i_4_) & (i_8_) & (!g34) & (!sk[38]) & (g57)) + ((i_3_) & (i_4_) & (i_8_) & (g34) & (!sk[38]) & (!g57)) + ((i_3_) & (i_4_) & (i_8_) & (g34) & (!sk[38]) & (g57)));
	assign g661 = (((!i_14_) & (!i_12_) & (!g112) & (!sk[39]) & (!g199) & (g122)) + ((!i_14_) & (!i_12_) & (!g112) & (!sk[39]) & (g199) & (g122)) + ((!i_14_) & (!i_12_) & (g112) & (!sk[39]) & (!g199) & (g122)) + ((!i_14_) & (!i_12_) & (g112) & (!sk[39]) & (g199) & (g122)) + ((!i_14_) & (!i_12_) & (g112) & (sk[39]) & (g199) & (!g122)) + ((!i_14_) & (!i_12_) & (g112) & (sk[39]) & (g199) & (g122)) + ((!i_14_) & (i_12_) & (!g112) & (!sk[39]) & (!g199) & (g122)) + ((!i_14_) & (i_12_) & (!g112) & (!sk[39]) & (g199) & (g122)) + ((!i_14_) & (i_12_) & (g112) & (!sk[39]) & (!g199) & (g122)) + ((!i_14_) & (i_12_) & (g112) & (!sk[39]) & (g199) & (g122)) + ((!i_14_) & (i_12_) & (g112) & (sk[39]) & (g199) & (!g122)) + ((!i_14_) & (i_12_) & (g112) & (sk[39]) & (g199) & (g122)) + ((i_14_) & (!i_12_) & (!g112) & (!sk[39]) & (!g199) & (!g122)) + ((i_14_) & (!i_12_) & (!g112) & (!sk[39]) & (!g199) & (g122)) + ((i_14_) & (!i_12_) & (!g112) & (!sk[39]) & (g199) & (!g122)) + ((i_14_) & (!i_12_) & (!g112) & (!sk[39]) & (g199) & (g122)) + ((i_14_) & (!i_12_) & (g112) & (!sk[39]) & (!g199) & (!g122)) + ((i_14_) & (!i_12_) & (g112) & (!sk[39]) & (!g199) & (g122)) + ((i_14_) & (!i_12_) & (g112) & (!sk[39]) & (g199) & (!g122)) + ((i_14_) & (!i_12_) & (g112) & (!sk[39]) & (g199) & (g122)) + ((i_14_) & (!i_12_) & (g112) & (sk[39]) & (!g199) & (!g122)) + ((i_14_) & (!i_12_) & (g112) & (sk[39]) & (g199) & (!g122)) + ((i_14_) & (!i_12_) & (g112) & (sk[39]) & (g199) & (g122)) + ((i_14_) & (i_12_) & (!g112) & (!sk[39]) & (!g199) & (!g122)) + ((i_14_) & (i_12_) & (!g112) & (!sk[39]) & (!g199) & (g122)) + ((i_14_) & (i_12_) & (!g112) & (!sk[39]) & (g199) & (!g122)) + ((i_14_) & (i_12_) & (!g112) & (!sk[39]) & (g199) & (g122)) + ((i_14_) & (i_12_) & (g112) & (!sk[39]) & (!g199) & (!g122)) + ((i_14_) & (i_12_) & (g112) & (!sk[39]) & (!g199) & (g122)) + ((i_14_) & (i_12_) & (g112) & (!sk[39]) & (g199) & (!g122)) + ((i_14_) & (i_12_) & (g112) & (!sk[39]) & (g199) & (g122)) + ((i_14_) & (i_12_) & (g112) & (sk[39]) & (g199) & (!g122)) + ((i_14_) & (i_12_) & (g112) & (sk[39]) & (g199) & (g122)));
	assign g662 = (((!g338) & (!g658) & (!g659) & (!g522) & (!g660) & (!g661)) + ((!g338) & (!g658) & (!g659) & (!g522) & (g660) & (!g661)) + ((g338) & (!g658) & (!g659) & (!g522) & (!g660) & (!g661)) + ((g338) & (!g658) & (!g659) & (!g522) & (g660) & (!g661)) + ((g338) & (!g658) & (!g659) & (g522) & (!g660) & (!g661)));
	assign g663 = (((!g146) & (!g630) & (!sk[41]) & (g657) & (g662)) + ((!g146) & (!g630) & (sk[41]) & (g657) & (g662)) + ((!g146) & (g630) & (!sk[41]) & (!g657) & (!g662)) + ((!g146) & (g630) & (!sk[41]) & (!g657) & (g662)) + ((!g146) & (g630) & (!sk[41]) & (g657) & (!g662)) + ((!g146) & (g630) & (!sk[41]) & (g657) & (g662)) + ((g146) & (!g630) & (!sk[41]) & (g657) & (!g662)) + ((g146) & (!g630) & (!sk[41]) & (g657) & (g662)) + ((g146) & (!g630) & (sk[41]) & (g657) & (g662)) + ((g146) & (g630) & (!sk[41]) & (!g657) & (!g662)) + ((g146) & (g630) & (!sk[41]) & (!g657) & (g662)) + ((g146) & (g630) & (!sk[41]) & (g657) & (!g662)) + ((g146) & (g630) & (!sk[41]) & (g657) & (g662)) + ((g146) & (g630) & (sk[41]) & (g657) & (g662)));
	assign g664 = (((!g635) & (!g637) & (g639) & (g645) & (g655) & (g663)));
	assign o_4_ = (((g73) & (!g358) & (!g458) & (!g521) & (!g634) & (!g664)) + ((g73) & (!g358) & (!g458) & (!g521) & (!g634) & (g664)) + ((g73) & (!g358) & (!g458) & (!g521) & (g634) & (!g664)) + ((g73) & (!g358) & (!g458) & (!g521) & (g634) & (g664)) + ((g73) & (!g358) & (!g458) & (g521) & (!g634) & (!g664)) + ((g73) & (!g358) & (!g458) & (g521) & (!g634) & (g664)) + ((g73) & (!g358) & (!g458) & (g521) & (g634) & (!g664)) + ((g73) & (!g358) & (!g458) & (g521) & (g634) & (g664)) + ((g73) & (!g358) & (g458) & (!g521) & (!g634) & (!g664)) + ((g73) & (!g358) & (g458) & (!g521) & (!g634) & (g664)) + ((g73) & (!g358) & (g458) & (!g521) & (g634) & (!g664)) + ((g73) & (!g358) & (g458) & (!g521) & (g634) & (g664)) + ((g73) & (!g358) & (g458) & (g521) & (!g634) & (!g664)) + ((g73) & (!g358) & (g458) & (g521) & (!g634) & (g664)) + ((g73) & (!g358) & (g458) & (g521) & (g634) & (!g664)) + ((g73) & (!g358) & (g458) & (g521) & (g634) & (g664)) + ((g73) & (g358) & (!g458) & (!g521) & (!g634) & (!g664)) + ((g73) & (g358) & (!g458) & (!g521) & (!g634) & (g664)) + ((g73) & (g358) & (!g458) & (!g521) & (g634) & (!g664)) + ((g73) & (g358) & (!g458) & (!g521) & (g634) & (g664)) + ((g73) & (g358) & (!g458) & (g521) & (!g634) & (!g664)) + ((g73) & (g358) & (!g458) & (g521) & (!g634) & (g664)) + ((g73) & (g358) & (!g458) & (g521) & (g634) & (!g664)) + ((g73) & (g358) & (!g458) & (g521) & (g634) & (g664)) + ((g73) & (g358) & (g458) & (!g521) & (!g634) & (!g664)) + ((g73) & (g358) & (g458) & (!g521) & (!g634) & (g664)) + ((g73) & (g358) & (g458) & (!g521) & (g634) & (!g664)) + ((g73) & (g358) & (g458) & (!g521) & (g634) & (g664)) + ((g73) & (g358) & (g458) & (g521) & (!g634) & (!g664)) + ((g73) & (g358) & (g458) & (g521) & (!g634) & (g664)) + ((g73) & (g358) & (g458) & (g521) & (g634) & (!g664)));
	assign g666 = (((!g107) & (!g130) & (!sk[44]) & (!g1782) & (!g148) & (g157)) + ((!g107) & (!g130) & (!sk[44]) & (!g1782) & (g148) & (g157)) + ((!g107) & (!g130) & (!sk[44]) & (g1782) & (!g148) & (g157)) + ((!g107) & (!g130) & (!sk[44]) & (g1782) & (g148) & (g157)) + ((!g107) & (g130) & (!sk[44]) & (!g1782) & (!g148) & (g157)) + ((!g107) & (g130) & (!sk[44]) & (!g1782) & (g148) & (g157)) + ((!g107) & (g130) & (!sk[44]) & (g1782) & (!g148) & (g157)) + ((!g107) & (g130) & (!sk[44]) & (g1782) & (g148) & (g157)) + ((g107) & (!g130) & (!sk[44]) & (!g1782) & (!g148) & (!g157)) + ((g107) & (!g130) & (!sk[44]) & (!g1782) & (!g148) & (g157)) + ((g107) & (!g130) & (!sk[44]) & (!g1782) & (g148) & (!g157)) + ((g107) & (!g130) & (!sk[44]) & (!g1782) & (g148) & (g157)) + ((g107) & (!g130) & (!sk[44]) & (g1782) & (!g148) & (!g157)) + ((g107) & (!g130) & (!sk[44]) & (g1782) & (!g148) & (g157)) + ((g107) & (!g130) & (!sk[44]) & (g1782) & (g148) & (!g157)) + ((g107) & (!g130) & (!sk[44]) & (g1782) & (g148) & (g157)) + ((g107) & (g130) & (!sk[44]) & (!g1782) & (!g148) & (!g157)) + ((g107) & (g130) & (!sk[44]) & (!g1782) & (!g148) & (g157)) + ((g107) & (g130) & (!sk[44]) & (!g1782) & (g148) & (!g157)) + ((g107) & (g130) & (!sk[44]) & (!g1782) & (g148) & (g157)) + ((g107) & (g130) & (!sk[44]) & (g1782) & (!g148) & (!g157)) + ((g107) & (g130) & (!sk[44]) & (g1782) & (!g148) & (g157)) + ((g107) & (g130) & (!sk[44]) & (g1782) & (g148) & (!g157)) + ((g107) & (g130) & (!sk[44]) & (g1782) & (g148) & (g157)) + ((g107) & (g130) & (sk[44]) & (g1782) & (g148) & (g157)));
	assign g667 = (((!g490) & (!g1737) & (!g499) & (!g1728) & (!sk[45]) & (g512)) + ((!g490) & (!g1737) & (!g499) & (g1728) & (!sk[45]) & (g512)) + ((!g490) & (!g1737) & (g499) & (!g1728) & (!sk[45]) & (g512)) + ((!g490) & (!g1737) & (g499) & (g1728) & (!sk[45]) & (g512)) + ((!g490) & (g1737) & (!g499) & (!g1728) & (!sk[45]) & (g512)) + ((!g490) & (g1737) & (!g499) & (g1728) & (!sk[45]) & (g512)) + ((!g490) & (g1737) & (g499) & (!g1728) & (!sk[45]) & (g512)) + ((!g490) & (g1737) & (g499) & (g1728) & (!sk[45]) & (g512)) + ((g490) & (!g1737) & (!g499) & (!g1728) & (!sk[45]) & (!g512)) + ((g490) & (!g1737) & (!g499) & (!g1728) & (!sk[45]) & (g512)) + ((g490) & (!g1737) & (!g499) & (g1728) & (!sk[45]) & (!g512)) + ((g490) & (!g1737) & (!g499) & (g1728) & (!sk[45]) & (g512)) + ((g490) & (!g1737) & (g499) & (!g1728) & (!sk[45]) & (!g512)) + ((g490) & (!g1737) & (g499) & (!g1728) & (!sk[45]) & (g512)) + ((g490) & (!g1737) & (g499) & (g1728) & (!sk[45]) & (!g512)) + ((g490) & (!g1737) & (g499) & (g1728) & (!sk[45]) & (g512)) + ((g490) & (g1737) & (!g499) & (!g1728) & (!sk[45]) & (!g512)) + ((g490) & (g1737) & (!g499) & (!g1728) & (!sk[45]) & (g512)) + ((g490) & (g1737) & (!g499) & (g1728) & (!sk[45]) & (!g512)) + ((g490) & (g1737) & (!g499) & (g1728) & (!sk[45]) & (g512)) + ((g490) & (g1737) & (g499) & (!g1728) & (!sk[45]) & (!g512)) + ((g490) & (g1737) & (g499) & (!g1728) & (!sk[45]) & (g512)) + ((g490) & (g1737) & (g499) & (g1728) & (!sk[45]) & (!g512)) + ((g490) & (g1737) & (g499) & (g1728) & (!sk[45]) & (g512)) + ((g490) & (g1737) & (g499) & (g1728) & (sk[45]) & (g512)));
	assign g668 = (((!g19) & (sk[46]) & (!g16) & (g145)) + ((g19) & (!sk[46]) & (!g16) & (!g145)) + ((g19) & (!sk[46]) & (!g16) & (g145)) + ((g19) & (!sk[46]) & (g16) & (!g145)) + ((g19) & (!sk[46]) & (g16) & (g145)) + ((g19) & (sk[46]) & (!g16) & (g145)) + ((g19) & (sk[46]) & (g16) & (g145)));
	assign g669 = (((!g7) & (sk[47]) & (!g93)) + ((!g7) & (sk[47]) & (g93)) + ((g7) & (!sk[47]) & (!g93)) + ((g7) & (!sk[47]) & (g93)) + ((g7) & (sk[47]) & (g93)));
	assign g670 = (((!sk[48]) & (g9) & (!g119)) + ((!sk[48]) & (g9) & (g119)) + ((sk[48]) & (g9) & (g119)));
	assign g671 = (((g7) & (!sk[49]) & (!g122)) + ((g7) & (!sk[49]) & (g122)) + ((g7) & (sk[49]) & (!g122)));
	assign g672 = (((!sk[50]) & (g9) & (!g102)) + ((!sk[50]) & (g9) & (g102)) + ((sk[50]) & (g9) & (!g102)));
	assign g673 = (((!i_8_) & (!sk[51]) & (!g16) & (g100) & (g672)) + ((!i_8_) & (!sk[51]) & (g16) & (!g100) & (!g672)) + ((!i_8_) & (!sk[51]) & (g16) & (!g100) & (g672)) + ((!i_8_) & (!sk[51]) & (g16) & (g100) & (!g672)) + ((!i_8_) & (!sk[51]) & (g16) & (g100) & (g672)) + ((i_8_) & (!sk[51]) & (!g16) & (g100) & (!g672)) + ((i_8_) & (!sk[51]) & (!g16) & (g100) & (g672)) + ((i_8_) & (!sk[51]) & (g16) & (!g100) & (!g672)) + ((i_8_) & (!sk[51]) & (g16) & (!g100) & (g672)) + ((i_8_) & (!sk[51]) & (g16) & (g100) & (!g672)) + ((i_8_) & (!sk[51]) & (g16) & (g100) & (g672)) + ((i_8_) & (sk[51]) & (!g16) & (g100) & (!g672)) + ((i_8_) & (sk[51]) & (!g16) & (g100) & (g672)) + ((i_8_) & (sk[51]) & (g16) & (g100) & (g672)));
	assign g674 = (((!g101) & (!g145) & (!g669) & (!g670) & (!g671) & (!g673)) + ((!g101) & (!g145) & (!g669) & (!g670) & (g671) & (!g673)) + ((!g101) & (!g145) & (!g669) & (g670) & (!g671) & (!g673)) + ((!g101) & (!g145) & (!g669) & (g670) & (g671) & (!g673)) + ((!g101) & (!g145) & (g669) & (!g670) & (!g671) & (!g673)) + ((!g101) & (!g145) & (g669) & (!g670) & (g671) & (!g673)) + ((!g101) & (!g145) & (g669) & (g670) & (!g671) & (!g673)) + ((!g101) & (!g145) & (g669) & (g670) & (g671) & (!g673)) + ((!g101) & (g145) & (g669) & (!g670) & (!g671) & (!g673)) + ((g101) & (!g145) & (!g669) & (!g670) & (!g671) & (!g673)) + ((g101) & (!g145) & (!g669) & (!g670) & (g671) & (!g673)) + ((g101) & (!g145) & (g669) & (!g670) & (!g671) & (!g673)) + ((g101) & (!g145) & (g669) & (!g670) & (g671) & (!g673)) + ((g101) & (g145) & (g669) & (!g670) & (!g671) & (!g673)));
	assign g675 = (((!sk[53]) & (g7) & (!g115)) + ((!sk[53]) & (g7) & (g115)) + ((sk[53]) & (g7) & (!g115)));
	assign g676 = (((g7) & (!sk[54]) & (!g158)) + ((g7) & (!sk[54]) & (g158)) + ((g7) & (sk[54]) & (g158)));
	assign g677 = (((g9) & (!sk[55]) & (!g131)) + ((g9) & (!sk[55]) & (g131)) + ((g9) & (sk[55]) & (g131)));
	assign g678 = (((!g9) & (sk[56]) & (!g95)) + ((!g9) & (sk[56]) & (g95)) + ((g9) & (!sk[56]) & (!g95)) + ((g9) & (!sk[56]) & (g95)) + ((g9) & (sk[56]) & (!g95)));
	assign g679 = (((!g323) & (!g284) & (!sk[57]) & (g678) & (g677)) + ((!g323) & (!g284) & (sk[57]) & (!g678) & (!g677)) + ((!g323) & (!g284) & (sk[57]) & (!g678) & (g677)) + ((!g323) & (!g284) & (sk[57]) & (g678) & (!g677)) + ((!g323) & (!g284) & (sk[57]) & (g678) & (g677)) + ((!g323) & (g284) & (!sk[57]) & (!g678) & (!g677)) + ((!g323) & (g284) & (!sk[57]) & (!g678) & (g677)) + ((!g323) & (g284) & (!sk[57]) & (g678) & (!g677)) + ((!g323) & (g284) & (!sk[57]) & (g678) & (g677)) + ((!g323) & (g284) & (sk[57]) & (!g678) & (!g677)) + ((!g323) & (g284) & (sk[57]) & (g678) & (!g677)) + ((g323) & (!g284) & (!sk[57]) & (g678) & (!g677)) + ((g323) & (!g284) & (!sk[57]) & (g678) & (g677)) + ((g323) & (!g284) & (sk[57]) & (g678) & (!g677)) + ((g323) & (g284) & (!sk[57]) & (!g678) & (!g677)) + ((g323) & (g284) & (!sk[57]) & (!g678) & (g677)) + ((g323) & (g284) & (!sk[57]) & (g678) & (!g677)) + ((g323) & (g284) & (!sk[57]) & (g678) & (g677)) + ((g323) & (g284) & (sk[57]) & (g678) & (!g677)));
	assign g680 = (((!g145) & (!g675) & (!g672) & (!g676) & (!g677) & (g679)) + ((!g145) & (!g675) & (!g672) & (!g676) & (g677) & (g679)) + ((!g145) & (!g675) & (!g672) & (g676) & (!g677) & (g679)) + ((!g145) & (!g675) & (!g672) & (g676) & (g677) & (g679)) + ((!g145) & (!g675) & (g672) & (!g676) & (!g677) & (g679)) + ((!g145) & (!g675) & (g672) & (!g676) & (g677) & (g679)) + ((!g145) & (!g675) & (g672) & (g676) & (!g677) & (g679)) + ((!g145) & (!g675) & (g672) & (g676) & (g677) & (g679)) + ((!g145) & (g675) & (!g672) & (!g676) & (!g677) & (g679)) + ((!g145) & (g675) & (!g672) & (!g676) & (g677) & (g679)) + ((!g145) & (g675) & (!g672) & (g676) & (!g677) & (g679)) + ((!g145) & (g675) & (!g672) & (g676) & (g677) & (g679)) + ((!g145) & (g675) & (g672) & (!g676) & (!g677) & (g679)) + ((!g145) & (g675) & (g672) & (!g676) & (g677) & (g679)) + ((!g145) & (g675) & (g672) & (g676) & (!g677) & (g679)) + ((!g145) & (g675) & (g672) & (g676) & (g677) & (g679)) + ((g145) & (!g675) & (!g672) & (!g676) & (!g677) & (g679)));
	assign g681 = (((!sk[59]) & (g19) & (!g16) & (!g112)) + ((!sk[59]) & (g19) & (!g16) & (g112)) + ((!sk[59]) & (g19) & (g16) & (!g112)) + ((!sk[59]) & (g19) & (g16) & (g112)) + ((sk[59]) & (!g19) & (!g16) & (g112)) + ((sk[59]) & (g19) & (!g16) & (g112)) + ((sk[59]) & (g19) & (g16) & (g112)));
	assign g682 = (((g112) & (!sk[60]) & (!g678) & (!g669)) + ((g112) & (!sk[60]) & (!g678) & (g669)) + ((g112) & (!sk[60]) & (g678) & (!g669)) + ((g112) & (!sk[60]) & (g678) & (g669)) + ((g112) & (sk[60]) & (!g678) & (!g669)) + ((g112) & (sk[60]) & (!g678) & (g669)) + ((g112) & (sk[60]) & (g678) & (!g669)));
	assign g683 = (((g112) & (!sk[61]) & (!g676) & (!g677)) + ((g112) & (!sk[61]) & (!g676) & (g677)) + ((g112) & (!sk[61]) & (g676) & (!g677)) + ((g112) & (!sk[61]) & (g676) & (g677)) + ((g112) & (sk[61]) & (!g676) & (g677)) + ((g112) & (sk[61]) & (g676) & (!g677)) + ((g112) & (sk[61]) & (g676) & (g677)));
	assign g684 = (((g112) & (!g675) & (!sk[62]) & (!g672)) + ((g112) & (!g675) & (!sk[62]) & (g672)) + ((g112) & (!g675) & (sk[62]) & (g672)) + ((g112) & (g675) & (!sk[62]) & (!g672)) + ((g112) & (g675) & (!sk[62]) & (g672)) + ((g112) & (g675) & (sk[62]) & (!g672)) + ((g112) & (g675) & (sk[62]) & (g672)));
	assign g685 = (((!i_8_) & (!sk[63]) & (!g100) & (g678) & (g677)) + ((!i_8_) & (!sk[63]) & (g100) & (!g678) & (!g677)) + ((!i_8_) & (!sk[63]) & (g100) & (!g678) & (g677)) + ((!i_8_) & (!sk[63]) & (g100) & (g678) & (!g677)) + ((!i_8_) & (!sk[63]) & (g100) & (g678) & (g677)) + ((i_8_) & (!sk[63]) & (!g100) & (g678) & (!g677)) + ((i_8_) & (!sk[63]) & (!g100) & (g678) & (g677)) + ((i_8_) & (!sk[63]) & (g100) & (!g678) & (!g677)) + ((i_8_) & (!sk[63]) & (g100) & (!g678) & (g677)) + ((i_8_) & (!sk[63]) & (g100) & (g678) & (!g677)) + ((i_8_) & (!sk[63]) & (g100) & (g678) & (g677)) + ((i_8_) & (sk[63]) & (g100) & (!g678) & (!g677)) + ((i_8_) & (sk[63]) & (g100) & (!g678) & (g677)) + ((i_8_) & (sk[63]) & (g100) & (g678) & (g677)));
	assign g686 = (((!g12) & (!sk[64]) & (!g112) & (g323) & (g670)) + ((!g12) & (!sk[64]) & (g112) & (!g323) & (!g670)) + ((!g12) & (!sk[64]) & (g112) & (!g323) & (g670)) + ((!g12) & (!sk[64]) & (g112) & (g323) & (!g670)) + ((!g12) & (!sk[64]) & (g112) & (g323) & (g670)) + ((!g12) & (sk[64]) & (!g112) & (!g323) & (!g670)) + ((!g12) & (sk[64]) & (!g112) & (!g323) & (g670)) + ((!g12) & (sk[64]) & (!g112) & (g323) & (!g670)) + ((!g12) & (sk[64]) & (!g112) & (g323) & (g670)) + ((!g12) & (sk[64]) & (g112) & (!g323) & (!g670)) + ((!g12) & (sk[64]) & (g112) & (g323) & (!g670)) + ((g12) & (!sk[64]) & (!g112) & (g323) & (!g670)) + ((g12) & (!sk[64]) & (!g112) & (g323) & (g670)) + ((g12) & (!sk[64]) & (g112) & (!g323) & (!g670)) + ((g12) & (!sk[64]) & (g112) & (!g323) & (g670)) + ((g12) & (!sk[64]) & (g112) & (g323) & (!g670)) + ((g12) & (!sk[64]) & (g112) & (g323) & (g670)) + ((g12) & (sk[64]) & (!g112) & (!g323) & (!g670)) + ((g12) & (sk[64]) & (!g112) & (!g323) & (g670)));
	assign g687 = (((!g681) & (!g682) & (!g683) & (!g684) & (!g685) & (g686)));
	assign g688 = (((!g19) & (!g16) & (!g136) & (!g151) & (!g678) & (!g669)) + ((!g19) & (!g16) & (!g136) & (!g151) & (!g678) & (g669)) + ((!g19) & (!g16) & (!g136) & (!g151) & (g678) & (!g669)) + ((!g19) & (!g16) & (!g136) & (!g151) & (g678) & (g669)) + ((!g19) & (g16) & (!g136) & (!g151) & (!g678) & (!g669)) + ((!g19) & (g16) & (!g136) & (!g151) & (!g678) & (g669)) + ((!g19) & (g16) & (!g136) & (!g151) & (g678) & (!g669)) + ((!g19) & (g16) & (!g136) & (!g151) & (g678) & (g669)) + ((!g19) & (g16) & (!g136) & (g151) & (g678) & (g669)) + ((!g19) & (g16) & (g136) & (!g151) & (!g678) & (!g669)) + ((!g19) & (g16) & (g136) & (!g151) & (!g678) & (g669)) + ((!g19) & (g16) & (g136) & (!g151) & (g678) & (!g669)) + ((!g19) & (g16) & (g136) & (!g151) & (g678) & (g669)) + ((!g19) & (g16) & (g136) & (g151) & (g678) & (g669)) + ((g19) & (!g16) & (!g136) & (!g151) & (!g678) & (!g669)) + ((g19) & (!g16) & (!g136) & (!g151) & (!g678) & (g669)) + ((g19) & (!g16) & (!g136) & (!g151) & (g678) & (!g669)) + ((g19) & (!g16) & (!g136) & (!g151) & (g678) & (g669)) + ((g19) & (g16) & (!g136) & (!g151) & (!g678) & (!g669)) + ((g19) & (g16) & (!g136) & (!g151) & (!g678) & (g669)) + ((g19) & (g16) & (!g136) & (!g151) & (g678) & (!g669)) + ((g19) & (g16) & (!g136) & (!g151) & (g678) & (g669)));
	assign g689 = (((!i_8_) & (!g12) & (!sk[67]) & (g135) & (g672)) + ((!i_8_) & (g12) & (!sk[67]) & (!g135) & (!g672)) + ((!i_8_) & (g12) & (!sk[67]) & (!g135) & (g672)) + ((!i_8_) & (g12) & (!sk[67]) & (g135) & (!g672)) + ((!i_8_) & (g12) & (!sk[67]) & (g135) & (g672)) + ((i_8_) & (!g12) & (!sk[67]) & (g135) & (!g672)) + ((i_8_) & (!g12) & (!sk[67]) & (g135) & (g672)) + ((i_8_) & (!g12) & (sk[67]) & (g135) & (g672)) + ((i_8_) & (g12) & (!sk[67]) & (!g135) & (!g672)) + ((i_8_) & (g12) & (!sk[67]) & (!g135) & (g672)) + ((i_8_) & (g12) & (!sk[67]) & (g135) & (!g672)) + ((i_8_) & (g12) & (!sk[67]) & (g135) & (g672)) + ((i_8_) & (g12) & (sk[67]) & (g135) & (!g672)) + ((i_8_) & (g12) & (sk[67]) & (g135) & (g672)));
	assign g690 = (((!i_8_) & (!sk[68]) & (!g135) & (g669) & (g676)) + ((!i_8_) & (!sk[68]) & (g135) & (!g669) & (!g676)) + ((!i_8_) & (!sk[68]) & (g135) & (!g669) & (g676)) + ((!i_8_) & (!sk[68]) & (g135) & (g669) & (!g676)) + ((!i_8_) & (!sk[68]) & (g135) & (g669) & (g676)) + ((i_8_) & (!sk[68]) & (!g135) & (g669) & (!g676)) + ((i_8_) & (!sk[68]) & (!g135) & (g669) & (g676)) + ((i_8_) & (!sk[68]) & (g135) & (!g669) & (!g676)) + ((i_8_) & (!sk[68]) & (g135) & (!g669) & (g676)) + ((i_8_) & (!sk[68]) & (g135) & (g669) & (!g676)) + ((i_8_) & (!sk[68]) & (g135) & (g669) & (g676)) + ((i_8_) & (sk[68]) & (g135) & (!g669) & (!g676)) + ((i_8_) & (sk[68]) & (g135) & (!g669) & (g676)) + ((i_8_) & (sk[68]) & (g135) & (g669) & (g676)));
	assign g691 = (((!sk[69]) & (!i_8_) & (!g135) & (g678) & (g670)) + ((!sk[69]) & (!i_8_) & (g135) & (!g678) & (!g670)) + ((!sk[69]) & (!i_8_) & (g135) & (!g678) & (g670)) + ((!sk[69]) & (!i_8_) & (g135) & (g678) & (!g670)) + ((!sk[69]) & (!i_8_) & (g135) & (g678) & (g670)) + ((!sk[69]) & (i_8_) & (!g135) & (g678) & (!g670)) + ((!sk[69]) & (i_8_) & (!g135) & (g678) & (g670)) + ((!sk[69]) & (i_8_) & (g135) & (!g678) & (!g670)) + ((!sk[69]) & (i_8_) & (g135) & (!g678) & (g670)) + ((!sk[69]) & (i_8_) & (g135) & (g678) & (!g670)) + ((!sk[69]) & (i_8_) & (g135) & (g678) & (g670)) + ((sk[69]) & (i_8_) & (g135) & (!g678) & (!g670)) + ((sk[69]) & (i_8_) & (g135) & (!g678) & (g670)) + ((sk[69]) & (i_8_) & (g135) & (g678) & (g670)));
	assign g692 = (((i_8_) & (!g12) & (g88) & (!g108) & (!g675) & (g676)) + ((i_8_) & (!g12) & (g88) & (!g108) & (g675) & (!g676)) + ((i_8_) & (!g12) & (g88) & (!g108) & (g675) & (g676)) + ((i_8_) & (!g12) & (g88) & (g108) & (!g675) & (g676)) + ((i_8_) & (!g12) & (g88) & (g108) & (g675) & (!g676)) + ((i_8_) & (!g12) & (g88) & (g108) & (g675) & (g676)) + ((i_8_) & (g12) & (!g88) & (g108) & (!g675) & (!g676)) + ((i_8_) & (g12) & (!g88) & (g108) & (!g675) & (g676)) + ((i_8_) & (g12) & (!g88) & (g108) & (g675) & (!g676)) + ((i_8_) & (g12) & (!g88) & (g108) & (g675) & (g676)) + ((i_8_) & (g12) & (g88) & (!g108) & (!g675) & (!g676)) + ((i_8_) & (g12) & (g88) & (!g108) & (!g675) & (g676)) + ((i_8_) & (g12) & (g88) & (!g108) & (g675) & (!g676)) + ((i_8_) & (g12) & (g88) & (!g108) & (g675) & (g676)) + ((i_8_) & (g12) & (g88) & (g108) & (!g675) & (!g676)) + ((i_8_) & (g12) & (g88) & (g108) & (!g675) & (g676)) + ((i_8_) & (g12) & (g88) & (g108) & (g675) & (!g676)) + ((i_8_) & (g12) & (g88) & (g108) & (g675) & (g676)));
	assign g693 = (((!g151) & (!g670) & (!g689) & (!g690) & (!g691) & (!g692)) + ((!g151) & (g670) & (!g689) & (!g690) & (!g691) & (!g692)) + ((g151) & (!g670) & (!g689) & (!g690) & (!g691) & (!g692)));
	assign g694 = (((!g668) & (g674) & (g680) & (g687) & (g688) & (g693)));
	assign g695 = (((!sk[73]) & (g8) & (!g145)) + ((!sk[73]) & (g8) & (g145)) + ((sk[73]) & (!g8) & (g145)));
	assign g696 = (((!g9) & (sk[74]) & (!g104)) + ((!g9) & (sk[74]) & (g104)) + ((g9) & (!sk[74]) & (!g104)) + ((g9) & (!sk[74]) & (g104)) + ((g9) & (sk[74]) & (!g104)));
	assign g697 = (((!sk[75]) & (!g112) & (!g136) & (g151) & (g696)) + ((!sk[75]) & (!g112) & (g136) & (!g151) & (!g696)) + ((!sk[75]) & (!g112) & (g136) & (!g151) & (g696)) + ((!sk[75]) & (!g112) & (g136) & (g151) & (!g696)) + ((!sk[75]) & (!g112) & (g136) & (g151) & (g696)) + ((!sk[75]) & (g112) & (!g136) & (g151) & (!g696)) + ((!sk[75]) & (g112) & (!g136) & (g151) & (g696)) + ((!sk[75]) & (g112) & (g136) & (!g151) & (!g696)) + ((!sk[75]) & (g112) & (g136) & (!g151) & (g696)) + ((!sk[75]) & (g112) & (g136) & (g151) & (!g696)) + ((!sk[75]) & (g112) & (g136) & (g151) & (g696)) + ((sk[75]) & (!g112) & (!g136) & (g151) & (!g696)) + ((sk[75]) & (!g112) & (g136) & (!g151) & (!g696)) + ((sk[75]) & (!g112) & (g136) & (g151) & (!g696)) + ((sk[75]) & (g112) & (!g136) & (!g151) & (!g696)) + ((sk[75]) & (g112) & (!g136) & (g151) & (!g696)) + ((sk[75]) & (g112) & (g136) & (!g151) & (!g696)) + ((sk[75]) & (g112) & (g136) & (g151) & (!g696)));
	assign g698 = (((!g8) & (!g10) & (!g112) & (!g323) & (!g696) & (!g670)) + ((!g8) & (!g10) & (!g112) & (!g323) & (!g696) & (g670)) + ((!g8) & (!g10) & (!g112) & (!g323) & (g696) & (!g670)) + ((!g8) & (!g10) & (!g112) & (!g323) & (g696) & (g670)) + ((!g8) & (!g10) & (!g112) & (g323) & (g696) & (!g670)) + ((!g8) & (g10) & (!g112) & (!g323) & (!g696) & (!g670)) + ((!g8) & (g10) & (!g112) & (!g323) & (!g696) & (g670)) + ((!g8) & (g10) & (!g112) & (!g323) & (g696) & (!g670)) + ((!g8) & (g10) & (!g112) & (!g323) & (g696) & (g670)) + ((g8) & (!g10) & (!g112) & (!g323) & (!g696) & (!g670)) + ((g8) & (!g10) & (!g112) & (!g323) & (!g696) & (g670)) + ((g8) & (!g10) & (!g112) & (!g323) & (g696) & (!g670)) + ((g8) & (!g10) & (!g112) & (!g323) & (g696) & (g670)) + ((g8) & (!g10) & (!g112) & (g323) & (g696) & (!g670)) + ((g8) & (!g10) & (g112) & (!g323) & (!g696) & (!g670)) + ((g8) & (!g10) & (g112) & (!g323) & (!g696) & (g670)) + ((g8) & (!g10) & (g112) & (!g323) & (g696) & (!g670)) + ((g8) & (!g10) & (g112) & (!g323) & (g696) & (g670)) + ((g8) & (!g10) & (g112) & (g323) & (g696) & (!g670)) + ((g8) & (g10) & (!g112) & (!g323) & (!g696) & (!g670)) + ((g8) & (g10) & (!g112) & (!g323) & (!g696) & (g670)) + ((g8) & (g10) & (!g112) & (!g323) & (g696) & (!g670)) + ((g8) & (g10) & (!g112) & (!g323) & (g696) & (g670)));
	assign g699 = (((!g10) & (!g12) & (!g101) & (!g145) & (!g696) & (g698)) + ((!g10) & (!g12) & (!g101) & (!g145) & (g696) & (g698)) + ((!g10) & (!g12) & (!g101) & (g145) & (g696) & (g698)) + ((!g10) & (!g12) & (g101) & (!g145) & (g696) & (g698)) + ((!g10) & (!g12) & (g101) & (g145) & (g696) & (g698)) + ((!g10) & (g12) & (!g101) & (!g145) & (!g696) & (g698)) + ((!g10) & (g12) & (!g101) & (!g145) & (g696) & (g698)) + ((!g10) & (g12) & (!g101) & (g145) & (g696) & (g698)) + ((g10) & (!g12) & (!g101) & (!g145) & (!g696) & (g698)) + ((g10) & (!g12) & (!g101) & (!g145) & (g696) & (g698)) + ((g10) & (!g12) & (!g101) & (g145) & (g696) & (g698)) + ((g10) & (g12) & (!g101) & (!g145) & (!g696) & (g698)) + ((g10) & (g12) & (!g101) & (!g145) & (g696) & (g698)) + ((g10) & (g12) & (!g101) & (g145) & (g696) & (g698)));
	assign g700 = (((!g8) & (!g10) & (!g23) & (!g136) & (!sk[78]) & (g151)) + ((!g8) & (!g10) & (!g23) & (!g136) & (sk[78]) & (!g151)) + ((!g8) & (!g10) & (!g23) & (g136) & (!sk[78]) & (g151)) + ((!g8) & (!g10) & (g23) & (!g136) & (!sk[78]) & (g151)) + ((!g8) & (!g10) & (g23) & (!g136) & (sk[78]) & (!g151)) + ((!g8) & (!g10) & (g23) & (g136) & (!sk[78]) & (g151)) + ((!g8) & (g10) & (!g23) & (!g136) & (!sk[78]) & (g151)) + ((!g8) & (g10) & (!g23) & (!g136) & (sk[78]) & (!g151)) + ((!g8) & (g10) & (!g23) & (g136) & (!sk[78]) & (g151)) + ((!g8) & (g10) & (g23) & (!g136) & (!sk[78]) & (g151)) + ((!g8) & (g10) & (g23) & (!g136) & (sk[78]) & (!g151)) + ((!g8) & (g10) & (g23) & (g136) & (!sk[78]) & (g151)) + ((g8) & (!g10) & (!g23) & (!g136) & (!sk[78]) & (!g151)) + ((g8) & (!g10) & (!g23) & (!g136) & (!sk[78]) & (g151)) + ((g8) & (!g10) & (!g23) & (!g136) & (sk[78]) & (!g151)) + ((g8) & (!g10) & (!g23) & (!g136) & (sk[78]) & (g151)) + ((g8) & (!g10) & (!g23) & (g136) & (!sk[78]) & (!g151)) + ((g8) & (!g10) & (!g23) & (g136) & (!sk[78]) & (g151)) + ((g8) & (!g10) & (!g23) & (g136) & (sk[78]) & (!g151)) + ((g8) & (!g10) & (!g23) & (g136) & (sk[78]) & (g151)) + ((g8) & (!g10) & (g23) & (!g136) & (!sk[78]) & (!g151)) + ((g8) & (!g10) & (g23) & (!g136) & (!sk[78]) & (g151)) + ((g8) & (!g10) & (g23) & (!g136) & (sk[78]) & (!g151)) + ((g8) & (!g10) & (g23) & (!g136) & (sk[78]) & (g151)) + ((g8) & (!g10) & (g23) & (g136) & (!sk[78]) & (!g151)) + ((g8) & (!g10) & (g23) & (g136) & (!sk[78]) & (g151)) + ((g8) & (g10) & (!g23) & (!g136) & (!sk[78]) & (!g151)) + ((g8) & (g10) & (!g23) & (!g136) & (!sk[78]) & (g151)) + ((g8) & (g10) & (!g23) & (!g136) & (sk[78]) & (!g151)) + ((g8) & (g10) & (!g23) & (g136) & (!sk[78]) & (!g151)) + ((g8) & (g10) & (!g23) & (g136) & (!sk[78]) & (g151)) + ((g8) & (g10) & (g23) & (!g136) & (!sk[78]) & (!g151)) + ((g8) & (g10) & (g23) & (!g136) & (!sk[78]) & (g151)) + ((g8) & (g10) & (g23) & (!g136) & (sk[78]) & (!g151)) + ((g8) & (g10) & (g23) & (g136) & (!sk[78]) & (!g151)) + ((g8) & (g10) & (g23) & (g136) & (!sk[78]) & (g151)));
	assign g701 = (((!g695) & (!sk[79]) & (!g697) & (g699) & (g700)) + ((!g695) & (!sk[79]) & (g697) & (!g699) & (!g700)) + ((!g695) & (!sk[79]) & (g697) & (!g699) & (g700)) + ((!g695) & (!sk[79]) & (g697) & (g699) & (!g700)) + ((!g695) & (!sk[79]) & (g697) & (g699) & (g700)) + ((!g695) & (sk[79]) & (!g697) & (g699) & (g700)) + ((g695) & (!sk[79]) & (!g697) & (g699) & (!g700)) + ((g695) & (!sk[79]) & (!g697) & (g699) & (g700)) + ((g695) & (!sk[79]) & (g697) & (!g699) & (!g700)) + ((g695) & (!sk[79]) & (g697) & (!g699) & (g700)) + ((g695) & (!sk[79]) & (g697) & (g699) & (!g700)) + ((g695) & (!sk[79]) & (g697) & (g699) & (g700)));
	assign g702 = (((g9) & (!sk[80]) & (!g124)) + ((g9) & (!sk[80]) & (g124)) + ((g9) & (sk[80]) & (g124)));
	assign g703 = (((g9) & (!sk[81]) & (!g22)) + ((g9) & (!sk[81]) & (g22)) + ((g9) & (sk[81]) & (g22)));
	assign g704 = (((!sk[82]) & (g9) & (!g122)) + ((!sk[82]) & (g9) & (g122)) + ((sk[82]) & (g9) & (!g122)));
	assign g705 = (((!g46) & (!sk[83]) & (!g118) & (g702) & (g704)) + ((!g46) & (!sk[83]) & (g118) & (!g702) & (!g704)) + ((!g46) & (!sk[83]) & (g118) & (!g702) & (g704)) + ((!g46) & (!sk[83]) & (g118) & (g702) & (!g704)) + ((!g46) & (!sk[83]) & (g118) & (g702) & (g704)) + ((!g46) & (sk[83]) & (g118) & (!g702) & (g704)) + ((!g46) & (sk[83]) & (g118) & (g702) & (!g704)) + ((!g46) & (sk[83]) & (g118) & (g702) & (g704)) + ((g46) & (!sk[83]) & (!g118) & (g702) & (!g704)) + ((g46) & (!sk[83]) & (!g118) & (g702) & (g704)) + ((g46) & (!sk[83]) & (g118) & (!g702) & (!g704)) + ((g46) & (!sk[83]) & (g118) & (!g702) & (g704)) + ((g46) & (!sk[83]) & (g118) & (g702) & (!g704)) + ((g46) & (!sk[83]) & (g118) & (g702) & (g704)) + ((g46) & (sk[83]) & (g118) & (!g702) & (!g704)) + ((g46) & (sk[83]) & (g118) & (!g702) & (g704)) + ((g46) & (sk[83]) & (g118) & (g702) & (!g704)) + ((g46) & (sk[83]) & (g118) & (g702) & (g704)));
	assign g706 = (((g9) & (!sk[84]) & (!g115)) + ((g9) & (!sk[84]) & (g115)) + ((g9) & (sk[84]) & (!g115)));
	assign g707 = (((!sk[85]) & (g477) & (!g703)) + ((!sk[85]) & (g477) & (g703)) + ((sk[85]) & (g477) & (!g703)));
	assign g708 = (((!i_8_) & (g108) & (!g464) & (!g696) & (!g706) & (!g707)) + ((!i_8_) & (g108) & (!g464) & (!g696) & (!g706) & (g707)) + ((!i_8_) & (g108) & (!g464) & (!g696) & (g706) & (!g707)) + ((!i_8_) & (g108) & (!g464) & (!g696) & (g706) & (g707)) + ((!i_8_) & (g108) & (!g464) & (g696) & (!g706) & (!g707)) + ((!i_8_) & (g108) & (!g464) & (g696) & (!g706) & (g707)) + ((!i_8_) & (g108) & (!g464) & (g696) & (g706) & (!g707)) + ((!i_8_) & (g108) & (!g464) & (g696) & (g706) & (g707)) + ((!i_8_) & (g108) & (g464) & (!g696) & (!g706) & (!g707)) + ((!i_8_) & (g108) & (g464) & (!g696) & (!g706) & (g707)) + ((!i_8_) & (g108) & (g464) & (!g696) & (g706) & (!g707)) + ((!i_8_) & (g108) & (g464) & (!g696) & (g706) & (g707)) + ((!i_8_) & (g108) & (g464) & (g696) & (g706) & (!g707)) + ((!i_8_) & (g108) & (g464) & (g696) & (g706) & (g707)) + ((i_8_) & (g108) & (!g464) & (!g696) & (!g706) & (!g707)) + ((i_8_) & (g108) & (!g464) & (!g696) & (!g706) & (g707)) + ((i_8_) & (g108) & (!g464) & (!g696) & (g706) & (!g707)) + ((i_8_) & (g108) & (!g464) & (!g696) & (g706) & (g707)) + ((i_8_) & (g108) & (!g464) & (g696) & (!g706) & (!g707)) + ((i_8_) & (g108) & (!g464) & (g696) & (!g706) & (g707)) + ((i_8_) & (g108) & (!g464) & (g696) & (g706) & (!g707)) + ((i_8_) & (g108) & (!g464) & (g696) & (g706) & (g707)) + ((i_8_) & (g108) & (g464) & (!g696) & (!g706) & (!g707)) + ((i_8_) & (g108) & (g464) & (!g696) & (g706) & (!g707)) + ((i_8_) & (g108) & (g464) & (!g696) & (g706) & (g707)) + ((i_8_) & (g108) & (g464) & (g696) & (!g706) & (!g707)) + ((i_8_) & (g108) & (g464) & (g696) & (g706) & (!g707)) + ((i_8_) & (g108) & (g464) & (g696) & (g706) & (g707)));
	assign g709 = (((!g109) & (!g702) & (!sk[87]) & (!g703) & (!g705) & (g708)) + ((!g109) & (!g702) & (!sk[87]) & (!g703) & (g705) & (g708)) + ((!g109) & (!g702) & (!sk[87]) & (g703) & (!g705) & (g708)) + ((!g109) & (!g702) & (!sk[87]) & (g703) & (g705) & (g708)) + ((!g109) & (!g702) & (sk[87]) & (!g703) & (!g705) & (!g708)) + ((!g109) & (!g702) & (sk[87]) & (g703) & (!g705) & (!g708)) + ((!g109) & (g702) & (!sk[87]) & (!g703) & (!g705) & (g708)) + ((!g109) & (g702) & (!sk[87]) & (!g703) & (g705) & (g708)) + ((!g109) & (g702) & (!sk[87]) & (g703) & (!g705) & (g708)) + ((!g109) & (g702) & (!sk[87]) & (g703) & (g705) & (g708)) + ((!g109) & (g702) & (sk[87]) & (!g703) & (!g705) & (!g708)) + ((!g109) & (g702) & (sk[87]) & (g703) & (!g705) & (!g708)) + ((g109) & (!g702) & (!sk[87]) & (!g703) & (!g705) & (!g708)) + ((g109) & (!g702) & (!sk[87]) & (!g703) & (!g705) & (g708)) + ((g109) & (!g702) & (!sk[87]) & (!g703) & (g705) & (!g708)) + ((g109) & (!g702) & (!sk[87]) & (!g703) & (g705) & (g708)) + ((g109) & (!g702) & (!sk[87]) & (g703) & (!g705) & (!g708)) + ((g109) & (!g702) & (!sk[87]) & (g703) & (!g705) & (g708)) + ((g109) & (!g702) & (!sk[87]) & (g703) & (g705) & (!g708)) + ((g109) & (!g702) & (!sk[87]) & (g703) & (g705) & (g708)) + ((g109) & (!g702) & (sk[87]) & (!g703) & (!g705) & (!g708)) + ((g109) & (g702) & (!sk[87]) & (!g703) & (!g705) & (!g708)) + ((g109) & (g702) & (!sk[87]) & (!g703) & (!g705) & (g708)) + ((g109) & (g702) & (!sk[87]) & (!g703) & (g705) & (!g708)) + ((g109) & (g702) & (!sk[87]) & (!g703) & (g705) & (g708)) + ((g109) & (g702) & (!sk[87]) & (g703) & (!g705) & (!g708)) + ((g109) & (g702) & (!sk[87]) & (g703) & (!g705) & (g708)) + ((g109) & (g702) & (!sk[87]) & (g703) & (g705) & (!g708)) + ((g109) & (g702) & (!sk[87]) & (g703) & (g705) & (g708)));
	assign g710 = (((g9) & (!sk[88]) & (!g158)) + ((g9) & (!sk[88]) & (g158)) + ((g9) & (sk[88]) & (g158)));
	assign g711 = (((!sk[89]) & (i_14_) & (!i_12_)) + ((!sk[89]) & (i_14_) & (i_12_)) + ((sk[89]) & (!i_14_) & (i_12_)));
	assign g712 = (((!g7) & (!i_8_) & (!sk[90]) & (!g115) & (!g122) & (g711)) + ((!g7) & (!i_8_) & (!sk[90]) & (!g115) & (g122) & (g711)) + ((!g7) & (!i_8_) & (!sk[90]) & (g115) & (!g122) & (g711)) + ((!g7) & (!i_8_) & (!sk[90]) & (g115) & (g122) & (g711)) + ((!g7) & (i_8_) & (!sk[90]) & (!g115) & (!g122) & (g711)) + ((!g7) & (i_8_) & (!sk[90]) & (!g115) & (g122) & (g711)) + ((!g7) & (i_8_) & (!sk[90]) & (g115) & (!g122) & (g711)) + ((!g7) & (i_8_) & (!sk[90]) & (g115) & (g122) & (g711)) + ((!g7) & (i_8_) & (sk[90]) & (!g115) & (!g122) & (g711)) + ((!g7) & (i_8_) & (sk[90]) & (!g115) & (g122) & (g711)) + ((!g7) & (i_8_) & (sk[90]) & (g115) & (!g122) & (g711)) + ((g7) & (!i_8_) & (!sk[90]) & (!g115) & (!g122) & (!g711)) + ((g7) & (!i_8_) & (!sk[90]) & (!g115) & (!g122) & (g711)) + ((g7) & (!i_8_) & (!sk[90]) & (!g115) & (g122) & (!g711)) + ((g7) & (!i_8_) & (!sk[90]) & (!g115) & (g122) & (g711)) + ((g7) & (!i_8_) & (!sk[90]) & (g115) & (!g122) & (!g711)) + ((g7) & (!i_8_) & (!sk[90]) & (g115) & (!g122) & (g711)) + ((g7) & (!i_8_) & (!sk[90]) & (g115) & (g122) & (!g711)) + ((g7) & (!i_8_) & (!sk[90]) & (g115) & (g122) & (g711)) + ((g7) & (!i_8_) & (sk[90]) & (!g115) & (!g122) & (!g711)) + ((g7) & (!i_8_) & (sk[90]) & (!g115) & (!g122) & (g711)) + ((g7) & (!i_8_) & (sk[90]) & (!g115) & (g122) & (!g711)) + ((g7) & (!i_8_) & (sk[90]) & (!g115) & (g122) & (g711)) + ((g7) & (i_8_) & (!sk[90]) & (!g115) & (!g122) & (!g711)) + ((g7) & (i_8_) & (!sk[90]) & (!g115) & (!g122) & (g711)) + ((g7) & (i_8_) & (!sk[90]) & (!g115) & (g122) & (!g711)) + ((g7) & (i_8_) & (!sk[90]) & (!g115) & (g122) & (g711)) + ((g7) & (i_8_) & (!sk[90]) & (g115) & (!g122) & (!g711)) + ((g7) & (i_8_) & (!sk[90]) & (g115) & (!g122) & (g711)) + ((g7) & (i_8_) & (!sk[90]) & (g115) & (g122) & (!g711)) + ((g7) & (i_8_) & (!sk[90]) & (g115) & (g122) & (g711)) + ((g7) & (i_8_) & (sk[90]) & (!g115) & (!g122) & (!g711)) + ((g7) & (i_8_) & (sk[90]) & (!g115) & (!g122) & (g711)) + ((g7) & (i_8_) & (sk[90]) & (!g115) & (g122) & (!g711)) + ((g7) & (i_8_) & (sk[90]) & (!g115) & (g122) & (g711)) + ((g7) & (i_8_) & (sk[90]) & (g115) & (!g122) & (!g711)) + ((g7) & (i_8_) & (sk[90]) & (g115) & (!g122) & (g711)));
	assign g713 = (((!g6) & (!i_15_) & (!sk[91]) & (g7) & (g461)) + ((!g6) & (i_15_) & (!sk[91]) & (!g7) & (!g461)) + ((!g6) & (i_15_) & (!sk[91]) & (!g7) & (g461)) + ((!g6) & (i_15_) & (!sk[91]) & (g7) & (!g461)) + ((!g6) & (i_15_) & (!sk[91]) & (g7) & (g461)) + ((g6) & (!i_15_) & (!sk[91]) & (g7) & (!g461)) + ((g6) & (!i_15_) & (!sk[91]) & (g7) & (g461)) + ((g6) & (i_15_) & (!sk[91]) & (!g7) & (!g461)) + ((g6) & (i_15_) & (!sk[91]) & (!g7) & (g461)) + ((g6) & (i_15_) & (!sk[91]) & (g7) & (!g461)) + ((g6) & (i_15_) & (!sk[91]) & (g7) & (g461)) + ((g6) & (i_15_) & (sk[91]) & (!g7) & (g461)) + ((g6) & (i_15_) & (sk[91]) & (g7) & (!g461)) + ((g6) & (i_15_) & (sk[91]) & (g7) & (g461)));
	assign g714 = (((!g4) & (!sk[92]) & (!g98) & (!g92) & (!g712) & (g713)) + ((!g4) & (!sk[92]) & (!g98) & (!g92) & (g712) & (g713)) + ((!g4) & (!sk[92]) & (!g98) & (g92) & (!g712) & (g713)) + ((!g4) & (!sk[92]) & (!g98) & (g92) & (g712) & (g713)) + ((!g4) & (!sk[92]) & (g98) & (!g92) & (!g712) & (g713)) + ((!g4) & (!sk[92]) & (g98) & (!g92) & (g712) & (g713)) + ((!g4) & (!sk[92]) & (g98) & (g92) & (!g712) & (g713)) + ((!g4) & (!sk[92]) & (g98) & (g92) & (g712) & (g713)) + ((g4) & (!sk[92]) & (!g98) & (!g92) & (!g712) & (!g713)) + ((g4) & (!sk[92]) & (!g98) & (!g92) & (!g712) & (g713)) + ((g4) & (!sk[92]) & (!g98) & (!g92) & (g712) & (!g713)) + ((g4) & (!sk[92]) & (!g98) & (!g92) & (g712) & (g713)) + ((g4) & (!sk[92]) & (!g98) & (g92) & (!g712) & (!g713)) + ((g4) & (!sk[92]) & (!g98) & (g92) & (!g712) & (g713)) + ((g4) & (!sk[92]) & (!g98) & (g92) & (g712) & (!g713)) + ((g4) & (!sk[92]) & (!g98) & (g92) & (g712) & (g713)) + ((g4) & (!sk[92]) & (g98) & (!g92) & (!g712) & (!g713)) + ((g4) & (!sk[92]) & (g98) & (!g92) & (!g712) & (g713)) + ((g4) & (!sk[92]) & (g98) & (!g92) & (g712) & (!g713)) + ((g4) & (!sk[92]) & (g98) & (!g92) & (g712) & (g713)) + ((g4) & (!sk[92]) & (g98) & (g92) & (!g712) & (!g713)) + ((g4) & (!sk[92]) & (g98) & (g92) & (!g712) & (g713)) + ((g4) & (!sk[92]) & (g98) & (g92) & (g712) & (!g713)) + ((g4) & (!sk[92]) & (g98) & (g92) & (g712) & (g713)) + ((g4) & (sk[92]) & (g98) & (!g92) & (!g712) & (!g713)) + ((g4) & (sk[92]) & (g98) & (!g92) & (!g712) & (g713)) + ((g4) & (sk[92]) & (g98) & (!g92) & (g712) & (!g713)) + ((g4) & (sk[92]) & (g98) & (!g92) & (g712) & (g713)) + ((g4) & (sk[92]) & (g98) & (g92) & (!g712) & (g713)) + ((g4) & (sk[92]) & (g98) & (g92) & (g712) & (!g713)) + ((g4) & (sk[92]) & (g98) & (g92) & (g712) & (g713)));
	assign g715 = (((!g251) & (!g281) & (!g710) & (sk[93]) & (!g714)) + ((!g251) & (!g281) & (g710) & (!sk[93]) & (g714)) + ((!g251) & (!g281) & (g710) & (sk[93]) & (!g714)) + ((!g251) & (g281) & (!g710) & (!sk[93]) & (!g714)) + ((!g251) & (g281) & (!g710) & (!sk[93]) & (g714)) + ((!g251) & (g281) & (!g710) & (sk[93]) & (!g714)) + ((!g251) & (g281) & (g710) & (!sk[93]) & (!g714)) + ((!g251) & (g281) & (g710) & (!sk[93]) & (g714)) + ((!g251) & (g281) & (g710) & (sk[93]) & (!g714)) + ((g251) & (!g281) & (g710) & (!sk[93]) & (!g714)) + ((g251) & (!g281) & (g710) & (!sk[93]) & (g714)) + ((g251) & (g281) & (!g710) & (!sk[93]) & (!g714)) + ((g251) & (g281) & (!g710) & (!sk[93]) & (g714)) + ((g251) & (g281) & (!g710) & (sk[93]) & (!g714)) + ((g251) & (g281) & (g710) & (!sk[93]) & (!g714)) + ((g251) & (g281) & (g710) & (!sk[93]) & (g714)));
	assign g716 = (((!i_8_) & (!g99) & (!sk[94]) & (g108) & (g467)) + ((!i_8_) & (g99) & (!sk[94]) & (!g108) & (!g467)) + ((!i_8_) & (g99) & (!sk[94]) & (!g108) & (g467)) + ((!i_8_) & (g99) & (!sk[94]) & (g108) & (!g467)) + ((!i_8_) & (g99) & (!sk[94]) & (g108) & (g467)) + ((!i_8_) & (g99) & (sk[94]) & (!g108) & (!g467)) + ((!i_8_) & (g99) & (sk[94]) & (g108) & (!g467)) + ((i_8_) & (!g99) & (!sk[94]) & (g108) & (!g467)) + ((i_8_) & (!g99) & (!sk[94]) & (g108) & (g467)) + ((i_8_) & (!g99) & (sk[94]) & (g108) & (!g467)) + ((i_8_) & (g99) & (!sk[94]) & (!g108) & (!g467)) + ((i_8_) & (g99) & (!sk[94]) & (!g108) & (g467)) + ((i_8_) & (g99) & (!sk[94]) & (g108) & (!g467)) + ((i_8_) & (g99) & (!sk[94]) & (g108) & (g467)) + ((i_8_) & (g99) & (sk[94]) & (!g108) & (!g467)) + ((i_8_) & (g99) & (sk[94]) & (g108) & (!g467)));
	assign g717 = (((!g19) & (!g99) & (!sk[95]) & (g115) & (g711)) + ((!g19) & (g99) & (!sk[95]) & (!g115) & (!g711)) + ((!g19) & (g99) & (!sk[95]) & (!g115) & (g711)) + ((!g19) & (g99) & (!sk[95]) & (g115) & (!g711)) + ((!g19) & (g99) & (!sk[95]) & (g115) & (g711)) + ((!g19) & (g99) & (sk[95]) & (!g115) & (g711)) + ((g19) & (!g99) & (!sk[95]) & (g115) & (!g711)) + ((g19) & (!g99) & (!sk[95]) & (g115) & (g711)) + ((g19) & (g99) & (!sk[95]) & (!g115) & (!g711)) + ((g19) & (g99) & (!sk[95]) & (!g115) & (g711)) + ((g19) & (g99) & (!sk[95]) & (g115) & (!g711)) + ((g19) & (g99) & (!sk[95]) & (g115) & (g711)) + ((g19) & (g99) & (sk[95]) & (!g115) & (!g711)) + ((g19) & (g99) & (sk[95]) & (!g115) & (g711)) + ((g19) & (g99) & (sk[95]) & (g115) & (!g711)) + ((g19) & (g99) & (sk[95]) & (g115) & (g711)));
	assign g718 = (((!i_8_) & (!g46) & (g88) & (!sk[96]) & (g704)) + ((!i_8_) & (!g46) & (g88) & (sk[96]) & (g704)) + ((!i_8_) & (g46) & (!g88) & (!sk[96]) & (!g704)) + ((!i_8_) & (g46) & (!g88) & (!sk[96]) & (g704)) + ((!i_8_) & (g46) & (g88) & (!sk[96]) & (!g704)) + ((!i_8_) & (g46) & (g88) & (!sk[96]) & (g704)) + ((!i_8_) & (g46) & (g88) & (sk[96]) & (!g704)) + ((!i_8_) & (g46) & (g88) & (sk[96]) & (g704)) + ((i_8_) & (!g46) & (g88) & (!sk[96]) & (!g704)) + ((i_8_) & (!g46) & (g88) & (!sk[96]) & (g704)) + ((i_8_) & (g46) & (!g88) & (!sk[96]) & (!g704)) + ((i_8_) & (g46) & (!g88) & (!sk[96]) & (g704)) + ((i_8_) & (g46) & (g88) & (!sk[96]) & (!g704)) + ((i_8_) & (g46) & (g88) & (!sk[96]) & (g704)));
	assign g719 = (((!i_8_) & (!g100) & (!sk[97]) & (g474) & (g460)) + ((!i_8_) & (g100) & (!sk[97]) & (!g474) & (!g460)) + ((!i_8_) & (g100) & (!sk[97]) & (!g474) & (g460)) + ((!i_8_) & (g100) & (!sk[97]) & (g474) & (!g460)) + ((!i_8_) & (g100) & (!sk[97]) & (g474) & (g460)) + ((i_8_) & (!g100) & (!sk[97]) & (g474) & (!g460)) + ((i_8_) & (!g100) & (!sk[97]) & (g474) & (g460)) + ((i_8_) & (g100) & (!sk[97]) & (!g474) & (!g460)) + ((i_8_) & (g100) & (!sk[97]) & (!g474) & (g460)) + ((i_8_) & (g100) & (!sk[97]) & (g474) & (!g460)) + ((i_8_) & (g100) & (!sk[97]) & (g474) & (g460)) + ((i_8_) & (g100) & (sk[97]) & (!g474) & (g460)) + ((i_8_) & (g100) & (sk[97]) & (g474) & (!g460)) + ((i_8_) & (g100) & (sk[97]) & (g474) & (g460)));
	assign g720 = (((!g112) & (!g186) & (!g120) & (!g477) & (!g474) & (!g671)) + ((!g112) & (!g186) & (!g120) & (!g477) & (!g474) & (g671)) + ((!g112) & (!g186) & (!g120) & (!g477) & (g474) & (!g671)) + ((!g112) & (!g186) & (!g120) & (!g477) & (g474) & (g671)) + ((!g112) & (!g186) & (!g120) & (g477) & (!g474) & (!g671)) + ((!g112) & (!g186) & (!g120) & (g477) & (!g474) & (g671)) + ((!g112) & (!g186) & (!g120) & (g477) & (g474) & (!g671)) + ((!g112) & (!g186) & (!g120) & (g477) & (g474) & (g671)) + ((!g112) & (!g186) & (g120) & (!g477) & (!g474) & (!g671)) + ((!g112) & (!g186) & (g120) & (!g477) & (!g474) & (g671)) + ((!g112) & (!g186) & (g120) & (!g477) & (g474) & (!g671)) + ((!g112) & (!g186) & (g120) & (!g477) & (g474) & (g671)) + ((!g112) & (!g186) & (g120) & (g477) & (!g474) & (!g671)) + ((!g112) & (!g186) & (g120) & (g477) & (!g474) & (g671)) + ((!g112) & (!g186) & (g120) & (g477) & (g474) & (!g671)) + ((!g112) & (!g186) & (g120) & (g477) & (g474) & (g671)) + ((!g112) & (g186) & (!g120) & (g477) & (!g474) & (!g671)) + ((!g112) & (g186) & (!g120) & (g477) & (!g474) & (g671)) + ((!g112) & (g186) & (g120) & (g477) & (!g474) & (!g671)) + ((!g112) & (g186) & (g120) & (g477) & (!g474) & (g671)) + ((g112) & (!g186) & (g120) & (!g477) & (!g474) & (!g671)) + ((g112) & (!g186) & (g120) & (!g477) & (g474) & (!g671)) + ((g112) & (!g186) & (g120) & (g477) & (!g474) & (!g671)) + ((g112) & (!g186) & (g120) & (g477) & (g474) & (!g671)) + ((g112) & (g186) & (g120) & (g477) & (!g474) & (!g671)));
	assign g721 = (((!sk[99]) & (!g716) & (!g717) & (!g718) & (!g719) & (g720)) + ((!sk[99]) & (!g716) & (!g717) & (!g718) & (g719) & (g720)) + ((!sk[99]) & (!g716) & (!g717) & (g718) & (!g719) & (g720)) + ((!sk[99]) & (!g716) & (!g717) & (g718) & (g719) & (g720)) + ((!sk[99]) & (!g716) & (g717) & (!g718) & (!g719) & (g720)) + ((!sk[99]) & (!g716) & (g717) & (!g718) & (g719) & (g720)) + ((!sk[99]) & (!g716) & (g717) & (g718) & (!g719) & (g720)) + ((!sk[99]) & (!g716) & (g717) & (g718) & (g719) & (g720)) + ((!sk[99]) & (g716) & (!g717) & (!g718) & (!g719) & (!g720)) + ((!sk[99]) & (g716) & (!g717) & (!g718) & (!g719) & (g720)) + ((!sk[99]) & (g716) & (!g717) & (!g718) & (g719) & (!g720)) + ((!sk[99]) & (g716) & (!g717) & (!g718) & (g719) & (g720)) + ((!sk[99]) & (g716) & (!g717) & (g718) & (!g719) & (!g720)) + ((!sk[99]) & (g716) & (!g717) & (g718) & (!g719) & (g720)) + ((!sk[99]) & (g716) & (!g717) & (g718) & (g719) & (!g720)) + ((!sk[99]) & (g716) & (!g717) & (g718) & (g719) & (g720)) + ((!sk[99]) & (g716) & (g717) & (!g718) & (!g719) & (!g720)) + ((!sk[99]) & (g716) & (g717) & (!g718) & (!g719) & (g720)) + ((!sk[99]) & (g716) & (g717) & (!g718) & (g719) & (!g720)) + ((!sk[99]) & (g716) & (g717) & (!g718) & (g719) & (g720)) + ((!sk[99]) & (g716) & (g717) & (g718) & (!g719) & (!g720)) + ((!sk[99]) & (g716) & (g717) & (g718) & (!g719) & (g720)) + ((!sk[99]) & (g716) & (g717) & (g718) & (g719) & (!g720)) + ((!sk[99]) & (g716) & (g717) & (g718) & (g719) & (g720)) + ((sk[99]) & (!g716) & (!g717) & (!g718) & (!g719) & (g720)));
	assign g722 = (((g44) & (!sk[100]) & (!g118) & (!g186)) + ((g44) & (!sk[100]) & (!g118) & (g186)) + ((g44) & (!sk[100]) & (g118) & (!g186)) + ((g44) & (!sk[100]) & (g118) & (g186)) + ((g44) & (sk[100]) & (!g118) & (g186)) + ((g44) & (sk[100]) & (g118) & (!g186)) + ((g44) & (sk[100]) & (g118) & (g186)));
	assign g723 = (((!g44) & (sk[101]) & (g108) & (g710)) + ((g44) & (!sk[101]) & (!g108) & (!g710)) + ((g44) & (!sk[101]) & (!g108) & (g710)) + ((g44) & (!sk[101]) & (g108) & (!g710)) + ((g44) & (!sk[101]) & (g108) & (g710)) + ((g44) & (sk[101]) & (g108) & (!g710)) + ((g44) & (sk[101]) & (g108) & (g710)));
	assign g724 = (((!g7) & (g158) & (sk[102]) & (g711)) + ((g7) & (!g158) & (!sk[102]) & (!g711)) + ((g7) & (!g158) & (!sk[102]) & (g711)) + ((g7) & (g158) & (!sk[102]) & (!g711)) + ((g7) & (g158) & (!sk[102]) & (g711)) + ((g7) & (g158) & (sk[102]) & (!g711)) + ((g7) & (g158) & (sk[102]) & (g711)));
	assign g725 = (((!g99) & (!g724) & (!sk[103]) & (g677) & (g710)) + ((!g99) & (g724) & (!sk[103]) & (!g677) & (!g710)) + ((!g99) & (g724) & (!sk[103]) & (!g677) & (g710)) + ((!g99) & (g724) & (!sk[103]) & (g677) & (!g710)) + ((!g99) & (g724) & (!sk[103]) & (g677) & (g710)) + ((g99) & (!g724) & (!sk[103]) & (g677) & (!g710)) + ((g99) & (!g724) & (!sk[103]) & (g677) & (g710)) + ((g99) & (!g724) & (sk[103]) & (!g677) & (g710)) + ((g99) & (!g724) & (sk[103]) & (g677) & (!g710)) + ((g99) & (!g724) & (sk[103]) & (g677) & (g710)) + ((g99) & (g724) & (!sk[103]) & (!g677) & (!g710)) + ((g99) & (g724) & (!sk[103]) & (!g677) & (g710)) + ((g99) & (g724) & (!sk[103]) & (g677) & (!g710)) + ((g99) & (g724) & (!sk[103]) & (g677) & (g710)) + ((g99) & (g724) & (sk[103]) & (!g677) & (!g710)) + ((g99) & (g724) & (sk[103]) & (!g677) & (g710)) + ((g99) & (g724) & (sk[103]) & (g677) & (!g710)) + ((g99) & (g724) & (sk[103]) & (g677) & (g710)));
	assign g726 = (((!g7) & (sk[104]) & (!g711)) + ((g7) & (!sk[104]) & (!g711)) + ((g7) & (!sk[104]) & (g711)));
	assign g727 = (((!g6) & (!sk[105]) & (!i_15_) & (!i_14_) & (!i_12_) & (i_13_)) + ((!g6) & (!sk[105]) & (!i_15_) & (!i_14_) & (i_12_) & (i_13_)) + ((!g6) & (!sk[105]) & (!i_15_) & (i_14_) & (!i_12_) & (i_13_)) + ((!g6) & (!sk[105]) & (!i_15_) & (i_14_) & (i_12_) & (i_13_)) + ((!g6) & (!sk[105]) & (i_15_) & (!i_14_) & (!i_12_) & (i_13_)) + ((!g6) & (!sk[105]) & (i_15_) & (!i_14_) & (i_12_) & (i_13_)) + ((!g6) & (!sk[105]) & (i_15_) & (i_14_) & (!i_12_) & (i_13_)) + ((!g6) & (!sk[105]) & (i_15_) & (i_14_) & (i_12_) & (i_13_)) + ((g6) & (!sk[105]) & (!i_15_) & (!i_14_) & (!i_12_) & (!i_13_)) + ((g6) & (!sk[105]) & (!i_15_) & (!i_14_) & (!i_12_) & (i_13_)) + ((g6) & (!sk[105]) & (!i_15_) & (!i_14_) & (i_12_) & (!i_13_)) + ((g6) & (!sk[105]) & (!i_15_) & (!i_14_) & (i_12_) & (i_13_)) + ((g6) & (!sk[105]) & (!i_15_) & (i_14_) & (!i_12_) & (!i_13_)) + ((g6) & (!sk[105]) & (!i_15_) & (i_14_) & (!i_12_) & (i_13_)) + ((g6) & (!sk[105]) & (!i_15_) & (i_14_) & (i_12_) & (!i_13_)) + ((g6) & (!sk[105]) & (!i_15_) & (i_14_) & (i_12_) & (i_13_)) + ((g6) & (!sk[105]) & (i_15_) & (!i_14_) & (!i_12_) & (!i_13_)) + ((g6) & (!sk[105]) & (i_15_) & (!i_14_) & (!i_12_) & (i_13_)) + ((g6) & (!sk[105]) & (i_15_) & (!i_14_) & (i_12_) & (!i_13_)) + ((g6) & (!sk[105]) & (i_15_) & (!i_14_) & (i_12_) & (i_13_)) + ((g6) & (!sk[105]) & (i_15_) & (i_14_) & (!i_12_) & (!i_13_)) + ((g6) & (!sk[105]) & (i_15_) & (i_14_) & (!i_12_) & (i_13_)) + ((g6) & (!sk[105]) & (i_15_) & (i_14_) & (i_12_) & (!i_13_)) + ((g6) & (!sk[105]) & (i_15_) & (i_14_) & (i_12_) & (i_13_)) + ((g6) & (sk[105]) & (i_15_) & (!i_14_) & (!i_12_) & (!i_13_)) + ((g6) & (sk[105]) & (i_15_) & (!i_14_) & (i_12_) & (!i_13_)) + ((g6) & (sk[105]) & (i_15_) & (!i_14_) & (i_12_) & (i_13_)));
	assign g728 = (((!sk[106]) & (!g18) & (!g59) & (g726) & (g727)) + ((!sk[106]) & (!g18) & (g59) & (!g726) & (!g727)) + ((!sk[106]) & (!g18) & (g59) & (!g726) & (g727)) + ((!sk[106]) & (!g18) & (g59) & (g726) & (!g727)) + ((!sk[106]) & (!g18) & (g59) & (g726) & (g727)) + ((!sk[106]) & (g18) & (!g59) & (g726) & (!g727)) + ((!sk[106]) & (g18) & (!g59) & (g726) & (g727)) + ((!sk[106]) & (g18) & (g59) & (!g726) & (!g727)) + ((!sk[106]) & (g18) & (g59) & (!g726) & (g727)) + ((!sk[106]) & (g18) & (g59) & (g726) & (!g727)) + ((!sk[106]) & (g18) & (g59) & (g726) & (g727)) + ((sk[106]) & (!g18) & (g59) & (!g726) & (!g727)) + ((sk[106]) & (!g18) & (g59) & (!g726) & (g727)) + ((sk[106]) & (!g18) & (g59) & (g726) & (g727)) + ((sk[106]) & (g18) & (g59) & (!g726) & (g727)) + ((sk[106]) & (g18) & (g59) & (g726) & (g727)));
	assign g729 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g59) & (g99) & (!g93)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g59) & (!g99) & (!g93)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g59) & (g99) & (!g93)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g59) & (g99) & (!g93)) + ((!i_14_) & (!i_12_) & (i_13_) & (g59) & (g99) & (!g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g59) & (g99) & (!g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (g59) & (!g99) & (!g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (g59) & (g99) & (!g93)) + ((!i_14_) & (i_12_) & (i_13_) & (!g59) & (g99) & (!g93)) + ((!i_14_) & (i_12_) & (i_13_) & (g59) & (!g99) & (!g93)) + ((!i_14_) & (i_12_) & (i_13_) & (g59) & (g99) & (!g93)));
	assign g730 = (((!g722) & (!g723) & (!g725) & (!sk[108]) & (!g728) & (g729)) + ((!g722) & (!g723) & (!g725) & (!sk[108]) & (g728) & (g729)) + ((!g722) & (!g723) & (!g725) & (sk[108]) & (!g728) & (!g729)) + ((!g722) & (!g723) & (g725) & (!sk[108]) & (!g728) & (g729)) + ((!g722) & (!g723) & (g725) & (!sk[108]) & (g728) & (g729)) + ((!g722) & (g723) & (!g725) & (!sk[108]) & (!g728) & (g729)) + ((!g722) & (g723) & (!g725) & (!sk[108]) & (g728) & (g729)) + ((!g722) & (g723) & (g725) & (!sk[108]) & (!g728) & (g729)) + ((!g722) & (g723) & (g725) & (!sk[108]) & (g728) & (g729)) + ((g722) & (!g723) & (!g725) & (!sk[108]) & (!g728) & (!g729)) + ((g722) & (!g723) & (!g725) & (!sk[108]) & (!g728) & (g729)) + ((g722) & (!g723) & (!g725) & (!sk[108]) & (g728) & (!g729)) + ((g722) & (!g723) & (!g725) & (!sk[108]) & (g728) & (g729)) + ((g722) & (!g723) & (g725) & (!sk[108]) & (!g728) & (!g729)) + ((g722) & (!g723) & (g725) & (!sk[108]) & (!g728) & (g729)) + ((g722) & (!g723) & (g725) & (!sk[108]) & (g728) & (!g729)) + ((g722) & (!g723) & (g725) & (!sk[108]) & (g728) & (g729)) + ((g722) & (g723) & (!g725) & (!sk[108]) & (!g728) & (!g729)) + ((g722) & (g723) & (!g725) & (!sk[108]) & (!g728) & (g729)) + ((g722) & (g723) & (!g725) & (!sk[108]) & (g728) & (!g729)) + ((g722) & (g723) & (!g725) & (!sk[108]) & (g728) & (g729)) + ((g722) & (g723) & (g725) & (!sk[108]) & (!g728) & (!g729)) + ((g722) & (g723) & (g725) & (!sk[108]) & (!g728) & (g729)) + ((g722) & (g723) & (g725) & (!sk[108]) & (g728) & (!g729)) + ((g722) & (g723) & (g725) & (!sk[108]) & (g728) & (g729)));
	assign g731 = (((!sk[109]) & (!g44) & (!g46) & (g99) & (g678)) + ((!sk[109]) & (!g44) & (g46) & (!g99) & (!g678)) + ((!sk[109]) & (!g44) & (g46) & (!g99) & (g678)) + ((!sk[109]) & (!g44) & (g46) & (g99) & (!g678)) + ((!sk[109]) & (!g44) & (g46) & (g99) & (g678)) + ((!sk[109]) & (g44) & (!g46) & (g99) & (!g678)) + ((!sk[109]) & (g44) & (!g46) & (g99) & (g678)) + ((!sk[109]) & (g44) & (g46) & (!g99) & (!g678)) + ((!sk[109]) & (g44) & (g46) & (!g99) & (g678)) + ((!sk[109]) & (g44) & (g46) & (g99) & (!g678)) + ((!sk[109]) & (g44) & (g46) & (g99) & (g678)) + ((sk[109]) & (!g44) & (!g46) & (g99) & (!g678)) + ((sk[109]) & (!g44) & (g46) & (g99) & (!g678)) + ((sk[109]) & (!g44) & (g46) & (g99) & (g678)) + ((sk[109]) & (g44) & (!g46) & (g99) & (!g678)) + ((sk[109]) & (g44) & (!g46) & (g99) & (g678)) + ((sk[109]) & (g44) & (g46) & (g99) & (!g678)) + ((sk[109]) & (g44) & (g46) & (g99) & (g678)));
	assign g732 = (((!sk[110]) & (!g99) & (!g477) & (g474) & (g460)) + ((!sk[110]) & (!g99) & (g477) & (!g474) & (!g460)) + ((!sk[110]) & (!g99) & (g477) & (!g474) & (g460)) + ((!sk[110]) & (!g99) & (g477) & (g474) & (!g460)) + ((!sk[110]) & (!g99) & (g477) & (g474) & (g460)) + ((!sk[110]) & (g99) & (!g477) & (g474) & (!g460)) + ((!sk[110]) & (g99) & (!g477) & (g474) & (g460)) + ((!sk[110]) & (g99) & (g477) & (!g474) & (!g460)) + ((!sk[110]) & (g99) & (g477) & (!g474) & (g460)) + ((!sk[110]) & (g99) & (g477) & (g474) & (!g460)) + ((!sk[110]) & (g99) & (g477) & (g474) & (g460)) + ((sk[110]) & (g99) & (!g477) & (!g474) & (!g460)) + ((sk[110]) & (g99) & (!g477) & (!g474) & (g460)) + ((sk[110]) & (g99) & (!g477) & (g474) & (!g460)) + ((sk[110]) & (g99) & (!g477) & (g474) & (g460)) + ((sk[110]) & (g99) & (g477) & (!g474) & (g460)) + ((sk[110]) & (g99) & (g477) & (g474) & (!g460)) + ((sk[110]) & (g99) & (g477) & (g474) & (g460)));
	assign g733 = (((!g99) & (!sk[111]) & (!g702) & (g706) & (g703)) + ((!g99) & (!sk[111]) & (g702) & (!g706) & (!g703)) + ((!g99) & (!sk[111]) & (g702) & (!g706) & (g703)) + ((!g99) & (!sk[111]) & (g702) & (g706) & (!g703)) + ((!g99) & (!sk[111]) & (g702) & (g706) & (g703)) + ((g99) & (!sk[111]) & (!g702) & (g706) & (!g703)) + ((g99) & (!sk[111]) & (!g702) & (g706) & (g703)) + ((g99) & (!sk[111]) & (g702) & (!g706) & (!g703)) + ((g99) & (!sk[111]) & (g702) & (!g706) & (g703)) + ((g99) & (!sk[111]) & (g702) & (g706) & (!g703)) + ((g99) & (!sk[111]) & (g702) & (g706) & (g703)) + ((g99) & (sk[111]) & (!g702) & (!g706) & (g703)) + ((g99) & (sk[111]) & (!g702) & (g706) & (!g703)) + ((g99) & (sk[111]) & (!g702) & (g706) & (g703)) + ((g99) & (sk[111]) & (g702) & (!g706) & (!g703)) + ((g99) & (sk[111]) & (g702) & (!g706) & (g703)) + ((g99) & (sk[111]) & (g702) & (g706) & (!g703)) + ((g99) & (sk[111]) & (g702) & (g706) & (g703)));
	assign g734 = (((g7) & (!sk[112]) & (!g124)) + ((g7) & (!sk[112]) & (g124)) + ((g7) & (sk[112]) & (g124)));
	assign g735 = (((!g134) & (!g478) & (g734) & (!sk[113]) & (g702)) + ((!g134) & (g478) & (!g734) & (!sk[113]) & (!g702)) + ((!g134) & (g478) & (!g734) & (!sk[113]) & (g702)) + ((!g134) & (g478) & (g734) & (!sk[113]) & (!g702)) + ((!g134) & (g478) & (g734) & (!sk[113]) & (g702)) + ((g134) & (!g478) & (!g734) & (sk[113]) & (g702)) + ((g134) & (!g478) & (g734) & (!sk[113]) & (!g702)) + ((g134) & (!g478) & (g734) & (!sk[113]) & (g702)) + ((g134) & (!g478) & (g734) & (sk[113]) & (!g702)) + ((g134) & (!g478) & (g734) & (sk[113]) & (g702)) + ((g134) & (g478) & (!g734) & (!sk[113]) & (!g702)) + ((g134) & (g478) & (!g734) & (!sk[113]) & (g702)) + ((g134) & (g478) & (!g734) & (sk[113]) & (!g702)) + ((g134) & (g478) & (!g734) & (sk[113]) & (g702)) + ((g134) & (g478) & (g734) & (!sk[113]) & (!g702)) + ((g134) & (g478) & (g734) & (!sk[113]) & (g702)) + ((g134) & (g478) & (g734) & (sk[113]) & (!g702)) + ((g134) & (g478) & (g734) & (sk[113]) & (g702)));
	assign g736 = (((!i_8_) & (!i_6_) & (i_7_) & (g98) & (!g478) & (g704)) + ((!i_8_) & (!i_6_) & (i_7_) & (g98) & (g478) & (!g704)) + ((!i_8_) & (!i_6_) & (i_7_) & (g98) & (g478) & (g704)) + ((!i_8_) & (i_6_) & (i_7_) & (g98) & (!g478) & (g704)) + ((!i_8_) & (i_6_) & (i_7_) & (g98) & (g478) & (!g704)) + ((!i_8_) & (i_6_) & (i_7_) & (g98) & (g478) & (g704)) + ((i_8_) & (!i_6_) & (i_7_) & (g98) & (g478) & (!g704)) + ((i_8_) & (!i_6_) & (i_7_) & (g98) & (g478) & (g704)) + ((i_8_) & (i_6_) & (i_7_) & (g98) & (!g478) & (g704)) + ((i_8_) & (i_6_) & (i_7_) & (g98) & (g478) & (g704)));
	assign g737 = (((!g731) & (!g732) & (!g733) & (!g735) & (!sk[115]) & (g736)) + ((!g731) & (!g732) & (!g733) & (!g735) & (sk[115]) & (!g736)) + ((!g731) & (!g732) & (!g733) & (g735) & (!sk[115]) & (g736)) + ((!g731) & (!g732) & (g733) & (!g735) & (!sk[115]) & (g736)) + ((!g731) & (!g732) & (g733) & (g735) & (!sk[115]) & (g736)) + ((!g731) & (g732) & (!g733) & (!g735) & (!sk[115]) & (g736)) + ((!g731) & (g732) & (!g733) & (g735) & (!sk[115]) & (g736)) + ((!g731) & (g732) & (g733) & (!g735) & (!sk[115]) & (g736)) + ((!g731) & (g732) & (g733) & (g735) & (!sk[115]) & (g736)) + ((g731) & (!g732) & (!g733) & (!g735) & (!sk[115]) & (!g736)) + ((g731) & (!g732) & (!g733) & (!g735) & (!sk[115]) & (g736)) + ((g731) & (!g732) & (!g733) & (g735) & (!sk[115]) & (!g736)) + ((g731) & (!g732) & (!g733) & (g735) & (!sk[115]) & (g736)) + ((g731) & (!g732) & (g733) & (!g735) & (!sk[115]) & (!g736)) + ((g731) & (!g732) & (g733) & (!g735) & (!sk[115]) & (g736)) + ((g731) & (!g732) & (g733) & (g735) & (!sk[115]) & (!g736)) + ((g731) & (!g732) & (g733) & (g735) & (!sk[115]) & (g736)) + ((g731) & (g732) & (!g733) & (!g735) & (!sk[115]) & (!g736)) + ((g731) & (g732) & (!g733) & (!g735) & (!sk[115]) & (g736)) + ((g731) & (g732) & (!g733) & (g735) & (!sk[115]) & (!g736)) + ((g731) & (g732) & (!g733) & (g735) & (!sk[115]) & (g736)) + ((g731) & (g732) & (g733) & (!g735) & (!sk[115]) & (!g736)) + ((g731) & (g732) & (g733) & (!g735) & (!sk[115]) & (g736)) + ((g731) & (g732) & (g733) & (g735) & (!sk[115]) & (!g736)) + ((g731) & (g732) & (g733) & (g735) & (!sk[115]) & (g736)));
	assign g738 = (((!sk[116]) & (!i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (g7)) + ((!sk[116]) & (!i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (g7)) + ((!sk[116]) & (!i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (g7)) + ((!sk[116]) & (!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g7)) + ((!sk[116]) & (!i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (g7)) + ((!sk[116]) & (!i_11_) & (i_9_) & (!i_10_) & (i_15_) & (g7)) + ((!sk[116]) & (!i_11_) & (i_9_) & (i_10_) & (!i_15_) & (g7)) + ((!sk[116]) & (!i_11_) & (i_9_) & (i_10_) & (i_15_) & (g7)) + ((!sk[116]) & (i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (!g7)) + ((!sk[116]) & (i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (g7)) + ((!sk[116]) & (i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (!g7)) + ((!sk[116]) & (i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (g7)) + ((!sk[116]) & (i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (!g7)) + ((!sk[116]) & (i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (g7)) + ((!sk[116]) & (i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!g7)) + ((!sk[116]) & (i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g7)) + ((!sk[116]) & (i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (!g7)) + ((!sk[116]) & (i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (g7)) + ((!sk[116]) & (i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!g7)) + ((!sk[116]) & (i_11_) & (i_9_) & (!i_10_) & (i_15_) & (g7)) + ((!sk[116]) & (i_11_) & (i_9_) & (i_10_) & (!i_15_) & (!g7)) + ((!sk[116]) & (i_11_) & (i_9_) & (i_10_) & (!i_15_) & (g7)) + ((!sk[116]) & (i_11_) & (i_9_) & (i_10_) & (i_15_) & (!g7)) + ((!sk[116]) & (i_11_) & (i_9_) & (i_10_) & (i_15_) & (g7)) + ((sk[116]) & (!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g7)) + ((sk[116]) & (!i_11_) & (i_9_) & (!i_10_) & (i_15_) & (g7)) + ((sk[116]) & (i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g7)));
	assign g739 = (((!sk[117]) & (!g23) & (!g96) & (!g734) & (!g669) & (g738)) + ((!sk[117]) & (!g23) & (!g96) & (!g734) & (g669) & (g738)) + ((!sk[117]) & (!g23) & (!g96) & (g734) & (!g669) & (g738)) + ((!sk[117]) & (!g23) & (!g96) & (g734) & (g669) & (g738)) + ((!sk[117]) & (!g23) & (g96) & (!g734) & (!g669) & (g738)) + ((!sk[117]) & (!g23) & (g96) & (!g734) & (g669) & (g738)) + ((!sk[117]) & (!g23) & (g96) & (g734) & (!g669) & (g738)) + ((!sk[117]) & (!g23) & (g96) & (g734) & (g669) & (g738)) + ((!sk[117]) & (g23) & (!g96) & (!g734) & (!g669) & (!g738)) + ((!sk[117]) & (g23) & (!g96) & (!g734) & (!g669) & (g738)) + ((!sk[117]) & (g23) & (!g96) & (!g734) & (g669) & (!g738)) + ((!sk[117]) & (g23) & (!g96) & (!g734) & (g669) & (g738)) + ((!sk[117]) & (g23) & (!g96) & (g734) & (!g669) & (!g738)) + ((!sk[117]) & (g23) & (!g96) & (g734) & (!g669) & (g738)) + ((!sk[117]) & (g23) & (!g96) & (g734) & (g669) & (!g738)) + ((!sk[117]) & (g23) & (!g96) & (g734) & (g669) & (g738)) + ((!sk[117]) & (g23) & (g96) & (!g734) & (!g669) & (!g738)) + ((!sk[117]) & (g23) & (g96) & (!g734) & (!g669) & (g738)) + ((!sk[117]) & (g23) & (g96) & (!g734) & (g669) & (!g738)) + ((!sk[117]) & (g23) & (g96) & (!g734) & (g669) & (g738)) + ((!sk[117]) & (g23) & (g96) & (g734) & (!g669) & (!g738)) + ((!sk[117]) & (g23) & (g96) & (g734) & (!g669) & (g738)) + ((!sk[117]) & (g23) & (g96) & (g734) & (g669) & (!g738)) + ((!sk[117]) & (g23) & (g96) & (g734) & (g669) & (g738)) + ((sk[117]) & (!g23) & (g96) & (!g734) & (g669) & (!g738)));
	assign g740 = (((!g46) & (!g90) & (!sk[118]) & (g704) & (g739)) + ((!g46) & (g90) & (!sk[118]) & (!g704) & (!g739)) + ((!g46) & (g90) & (!sk[118]) & (!g704) & (g739)) + ((!g46) & (g90) & (!sk[118]) & (g704) & (!g739)) + ((!g46) & (g90) & (!sk[118]) & (g704) & (g739)) + ((!g46) & (g90) & (sk[118]) & (!g704) & (g739)) + ((g46) & (!g90) & (!sk[118]) & (g704) & (!g739)) + ((g46) & (!g90) & (!sk[118]) & (g704) & (g739)) + ((g46) & (g90) & (!sk[118]) & (!g704) & (!g739)) + ((g46) & (g90) & (!sk[118]) & (!g704) & (g739)) + ((g46) & (g90) & (!sk[118]) & (g704) & (!g739)) + ((g46) & (g90) & (!sk[118]) & (g704) & (g739)));
	assign g741 = (((!g243) & (!g251) & (!g460) & (!sk[119]) & (!g724) & (g740)) + ((!g243) & (!g251) & (!g460) & (!sk[119]) & (g724) & (g740)) + ((!g243) & (!g251) & (!g460) & (sk[119]) & (!g724) & (!g740)) + ((!g243) & (!g251) & (!g460) & (sk[119]) & (!g724) & (g740)) + ((!g243) & (!g251) & (!g460) & (sk[119]) & (g724) & (!g740)) + ((!g243) & (!g251) & (!g460) & (sk[119]) & (g724) & (g740)) + ((!g243) & (!g251) & (g460) & (!sk[119]) & (!g724) & (g740)) + ((!g243) & (!g251) & (g460) & (!sk[119]) & (g724) & (g740)) + ((!g243) & (!g251) & (g460) & (sk[119]) & (!g724) & (!g740)) + ((!g243) & (!g251) & (g460) & (sk[119]) & (!g724) & (g740)) + ((!g243) & (!g251) & (g460) & (sk[119]) & (g724) & (!g740)) + ((!g243) & (!g251) & (g460) & (sk[119]) & (g724) & (g740)) + ((!g243) & (g251) & (!g460) & (!sk[119]) & (!g724) & (g740)) + ((!g243) & (g251) & (!g460) & (!sk[119]) & (g724) & (g740)) + ((!g243) & (g251) & (!g460) & (sk[119]) & (!g724) & (!g740)) + ((!g243) & (g251) & (!g460) & (sk[119]) & (!g724) & (g740)) + ((!g243) & (g251) & (g460) & (!sk[119]) & (!g724) & (g740)) + ((!g243) & (g251) & (g460) & (!sk[119]) & (g724) & (g740)) + ((g243) & (!g251) & (!g460) & (!sk[119]) & (!g724) & (!g740)) + ((g243) & (!g251) & (!g460) & (!sk[119]) & (!g724) & (g740)) + ((g243) & (!g251) & (!g460) & (!sk[119]) & (g724) & (!g740)) + ((g243) & (!g251) & (!g460) & (!sk[119]) & (g724) & (g740)) + ((g243) & (!g251) & (!g460) & (sk[119]) & (!g724) & (g740)) + ((g243) & (!g251) & (!g460) & (sk[119]) & (g724) & (g740)) + ((g243) & (!g251) & (g460) & (!sk[119]) & (!g724) & (!g740)) + ((g243) & (!g251) & (g460) & (!sk[119]) & (!g724) & (g740)) + ((g243) & (!g251) & (g460) & (!sk[119]) & (g724) & (!g740)) + ((g243) & (!g251) & (g460) & (!sk[119]) & (g724) & (g740)) + ((g243) & (!g251) & (g460) & (sk[119]) & (!g724) & (g740)) + ((g243) & (!g251) & (g460) & (sk[119]) & (g724) & (g740)) + ((g243) & (g251) & (!g460) & (!sk[119]) & (!g724) & (!g740)) + ((g243) & (g251) & (!g460) & (!sk[119]) & (!g724) & (g740)) + ((g243) & (g251) & (!g460) & (!sk[119]) & (g724) & (!g740)) + ((g243) & (g251) & (!g460) & (!sk[119]) & (g724) & (g740)) + ((g243) & (g251) & (!g460) & (sk[119]) & (!g724) & (g740)) + ((g243) & (g251) & (g460) & (!sk[119]) & (!g724) & (!g740)) + ((g243) & (g251) & (g460) & (!sk[119]) & (!g724) & (g740)) + ((g243) & (g251) & (g460) & (!sk[119]) & (g724) & (!g740)) + ((g243) & (g251) & (g460) & (!sk[119]) & (g724) & (g740)));
	assign g742 = (((!sk[120]) & (!g715) & (!g721) & (!g730) & (!g737) & (g741)) + ((!sk[120]) & (!g715) & (!g721) & (!g730) & (g737) & (g741)) + ((!sk[120]) & (!g715) & (!g721) & (g730) & (!g737) & (g741)) + ((!sk[120]) & (!g715) & (!g721) & (g730) & (g737) & (g741)) + ((!sk[120]) & (!g715) & (g721) & (!g730) & (!g737) & (g741)) + ((!sk[120]) & (!g715) & (g721) & (!g730) & (g737) & (g741)) + ((!sk[120]) & (!g715) & (g721) & (g730) & (!g737) & (g741)) + ((!sk[120]) & (!g715) & (g721) & (g730) & (g737) & (g741)) + ((!sk[120]) & (g715) & (!g721) & (!g730) & (!g737) & (!g741)) + ((!sk[120]) & (g715) & (!g721) & (!g730) & (!g737) & (g741)) + ((!sk[120]) & (g715) & (!g721) & (!g730) & (g737) & (!g741)) + ((!sk[120]) & (g715) & (!g721) & (!g730) & (g737) & (g741)) + ((!sk[120]) & (g715) & (!g721) & (g730) & (!g737) & (!g741)) + ((!sk[120]) & (g715) & (!g721) & (g730) & (!g737) & (g741)) + ((!sk[120]) & (g715) & (!g721) & (g730) & (g737) & (!g741)) + ((!sk[120]) & (g715) & (!g721) & (g730) & (g737) & (g741)) + ((!sk[120]) & (g715) & (g721) & (!g730) & (!g737) & (!g741)) + ((!sk[120]) & (g715) & (g721) & (!g730) & (!g737) & (g741)) + ((!sk[120]) & (g715) & (g721) & (!g730) & (g737) & (!g741)) + ((!sk[120]) & (g715) & (g721) & (!g730) & (g737) & (g741)) + ((!sk[120]) & (g715) & (g721) & (g730) & (!g737) & (!g741)) + ((!sk[120]) & (g715) & (g721) & (g730) & (!g737) & (g741)) + ((!sk[120]) & (g715) & (g721) & (g730) & (g737) & (!g741)) + ((!sk[120]) & (g715) & (g721) & (g730) & (g737) & (g741)) + ((sk[120]) & (g715) & (g721) & (g730) & (g737) & (g741)));
	assign g743 = (((!sk[121]) & (!g7) & (!g9) & (!g22) & (!g100) & (g277)) + ((!sk[121]) & (!g7) & (!g9) & (!g22) & (g100) & (g277)) + ((!sk[121]) & (!g7) & (!g9) & (g22) & (!g100) & (g277)) + ((!sk[121]) & (!g7) & (!g9) & (g22) & (g100) & (g277)) + ((!sk[121]) & (!g7) & (g9) & (!g22) & (!g100) & (g277)) + ((!sk[121]) & (!g7) & (g9) & (!g22) & (g100) & (g277)) + ((!sk[121]) & (!g7) & (g9) & (g22) & (!g100) & (g277)) + ((!sk[121]) & (!g7) & (g9) & (g22) & (g100) & (g277)) + ((!sk[121]) & (g7) & (!g9) & (!g22) & (!g100) & (!g277)) + ((!sk[121]) & (g7) & (!g9) & (!g22) & (!g100) & (g277)) + ((!sk[121]) & (g7) & (!g9) & (!g22) & (g100) & (!g277)) + ((!sk[121]) & (g7) & (!g9) & (!g22) & (g100) & (g277)) + ((!sk[121]) & (g7) & (!g9) & (g22) & (!g100) & (!g277)) + ((!sk[121]) & (g7) & (!g9) & (g22) & (!g100) & (g277)) + ((!sk[121]) & (g7) & (!g9) & (g22) & (g100) & (!g277)) + ((!sk[121]) & (g7) & (!g9) & (g22) & (g100) & (g277)) + ((!sk[121]) & (g7) & (g9) & (!g22) & (!g100) & (!g277)) + ((!sk[121]) & (g7) & (g9) & (!g22) & (!g100) & (g277)) + ((!sk[121]) & (g7) & (g9) & (!g22) & (g100) & (!g277)) + ((!sk[121]) & (g7) & (g9) & (!g22) & (g100) & (g277)) + ((!sk[121]) & (g7) & (g9) & (g22) & (!g100) & (!g277)) + ((!sk[121]) & (g7) & (g9) & (g22) & (!g100) & (g277)) + ((!sk[121]) & (g7) & (g9) & (g22) & (g100) & (!g277)) + ((!sk[121]) & (g7) & (g9) & (g22) & (g100) & (g277)) + ((sk[121]) & (!g7) & (g9) & (g22) & (!g100) & (!g277)) + ((sk[121]) & (!g7) & (g9) & (g22) & (g100) & (!g277)) + ((sk[121]) & (g7) & (!g9) & (g22) & (g100) & (!g277)) + ((sk[121]) & (g7) & (!g9) & (g22) & (g100) & (g277)) + ((sk[121]) & (g7) & (g9) & (g22) & (!g100) & (!g277)) + ((sk[121]) & (g7) & (g9) & (g22) & (g100) & (!g277)) + ((sk[121]) & (g7) & (g9) & (g22) & (g100) & (g277)));
	assign g744 = (((!i_14_) & (!i_12_) & (!i_13_) & (g101) & (!g145) & (!g93)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g101) & (g145) & (!g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (g101) & (!g145) & (!g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (g101) & (g145) & (!g93)) + ((!i_14_) & (i_12_) & (i_13_) & (g101) & (!g145) & (!g93)) + ((!i_14_) & (i_12_) & (i_13_) & (g101) & (g145) & (!g93)) + ((i_14_) & (!i_12_) & (i_13_) & (!g101) & (g145) & (!g93)) + ((i_14_) & (!i_12_) & (i_13_) & (g101) & (g145) & (!g93)));
	assign g745 = (((!i_8_) & (!g18) & (g4) & (g98) & (!g122) & (!g726)) + ((!i_8_) & (g18) & (g4) & (g98) & (!g122) & (!g726)) + ((i_8_) & (!g18) & (g4) & (g98) & (!g122) & (!g726)) + ((i_8_) & (!g18) & (g4) & (g98) & (g122) & (!g726)));
	assign g746 = (((!i_6_) & (sk[124]) & (g87)) + ((i_6_) & (!sk[124]) & (!g87)) + ((i_6_) & (!sk[124]) & (g87)));
	assign g747 = (((!i_8_) & (!g134) & (!g135) & (g746) & (g671) & (!g704)) + ((!i_8_) & (!g134) & (!g135) & (g746) & (g671) & (g704)) + ((!i_8_) & (!g134) & (g135) & (g746) & (g671) & (!g704)) + ((!i_8_) & (!g134) & (g135) & (g746) & (g671) & (g704)) + ((!i_8_) & (g134) & (!g135) & (!g746) & (!g671) & (g704)) + ((!i_8_) & (g134) & (!g135) & (!g746) & (g671) & (g704)) + ((!i_8_) & (g134) & (!g135) & (g746) & (!g671) & (g704)) + ((!i_8_) & (g134) & (!g135) & (g746) & (g671) & (!g704)) + ((!i_8_) & (g134) & (!g135) & (g746) & (g671) & (g704)) + ((!i_8_) & (g134) & (g135) & (!g746) & (!g671) & (g704)) + ((!i_8_) & (g134) & (g135) & (!g746) & (g671) & (g704)) + ((!i_8_) & (g134) & (g135) & (g746) & (!g671) & (g704)) + ((!i_8_) & (g134) & (g135) & (g746) & (g671) & (!g704)) + ((!i_8_) & (g134) & (g135) & (g746) & (g671) & (g704)) + ((i_8_) & (!g134) & (!g135) & (g746) & (g671) & (!g704)) + ((i_8_) & (!g134) & (!g135) & (g746) & (g671) & (g704)) + ((i_8_) & (!g134) & (g135) & (!g746) & (g671) & (!g704)) + ((i_8_) & (!g134) & (g135) & (!g746) & (g671) & (g704)) + ((i_8_) & (!g134) & (g135) & (g746) & (g671) & (!g704)) + ((i_8_) & (!g134) & (g135) & (g746) & (g671) & (g704)) + ((i_8_) & (g134) & (!g135) & (!g746) & (!g671) & (g704)) + ((i_8_) & (g134) & (!g135) & (!g746) & (g671) & (g704)) + ((i_8_) & (g134) & (!g135) & (g746) & (!g671) & (g704)) + ((i_8_) & (g134) & (!g135) & (g746) & (g671) & (!g704)) + ((i_8_) & (g134) & (!g135) & (g746) & (g671) & (g704)) + ((i_8_) & (g134) & (g135) & (!g746) & (!g671) & (g704)) + ((i_8_) & (g134) & (g135) & (!g746) & (g671) & (!g704)) + ((i_8_) & (g134) & (g135) & (!g746) & (g671) & (g704)) + ((i_8_) & (g134) & (g135) & (g746) & (!g671) & (g704)) + ((i_8_) & (g134) & (g135) & (g746) & (g671) & (!g704)) + ((i_8_) & (g134) & (g135) & (g746) & (g671) & (g704)));
	assign g748 = (((!g145) & (!g135) & (!g460) & (!g710) & (!g745) & (!g747)) + ((!g145) & (!g135) & (!g460) & (g710) & (!g745) & (!g747)) + ((!g145) & (!g135) & (g460) & (!g710) & (!g745) & (!g747)) + ((!g145) & (!g135) & (g460) & (g710) & (!g745) & (!g747)) + ((!g145) & (g135) & (!g460) & (!g710) & (!g745) & (!g747)) + ((!g145) & (g135) & (g460) & (!g710) & (!g745) & (!g747)) + ((g145) & (!g135) & (!g460) & (!g710) & (!g745) & (!g747)) + ((g145) & (!g135) & (!g460) & (g710) & (!g745) & (!g747)) + ((g145) & (g135) & (!g460) & (!g710) & (!g745) & (!g747)));
	assign g749 = (((i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g9) & (!g660)) + ((i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g9) & (g660)) + ((i_11_) & (i_9_) & (!i_10_) & (i_15_) & (g9) & (g660)));
	assign g750 = (((!g134) & (!g251) & (!sk[0]) & (!g660) & (!g704) & (g749)) + ((!g134) & (!g251) & (!sk[0]) & (!g660) & (g704) & (g749)) + ((!g134) & (!g251) & (!sk[0]) & (g660) & (!g704) & (g749)) + ((!g134) & (!g251) & (!sk[0]) & (g660) & (g704) & (g749)) + ((!g134) & (!g251) & (sk[0]) & (g660) & (g704) & (g749)) + ((!g134) & (g251) & (!sk[0]) & (!g660) & (!g704) & (g749)) + ((!g134) & (g251) & (!sk[0]) & (!g660) & (g704) & (g749)) + ((!g134) & (g251) & (!sk[0]) & (g660) & (!g704) & (g749)) + ((!g134) & (g251) & (!sk[0]) & (g660) & (g704) & (g749)) + ((!g134) & (g251) & (sk[0]) & (!g660) & (!g704) & (g749)) + ((!g134) & (g251) & (sk[0]) & (!g660) & (g704) & (g749)) + ((!g134) & (g251) & (sk[0]) & (g660) & (!g704) & (g749)) + ((!g134) & (g251) & (sk[0]) & (g660) & (g704) & (g749)) + ((g134) & (!g251) & (!sk[0]) & (!g660) & (!g704) & (!g749)) + ((g134) & (!g251) & (!sk[0]) & (!g660) & (!g704) & (g749)) + ((g134) & (!g251) & (!sk[0]) & (!g660) & (g704) & (!g749)) + ((g134) & (!g251) & (!sk[0]) & (!g660) & (g704) & (g749)) + ((g134) & (!g251) & (!sk[0]) & (g660) & (!g704) & (!g749)) + ((g134) & (!g251) & (!sk[0]) & (g660) & (!g704) & (g749)) + ((g134) & (!g251) & (!sk[0]) & (g660) & (g704) & (!g749)) + ((g134) & (!g251) & (!sk[0]) & (g660) & (g704) & (g749)) + ((g134) & (!g251) & (sk[0]) & (!g660) & (!g704) & (g749)) + ((g134) & (!g251) & (sk[0]) & (!g660) & (g704) & (g749)) + ((g134) & (!g251) & (sk[0]) & (g660) & (!g704) & (g749)) + ((g134) & (!g251) & (sk[0]) & (g660) & (g704) & (g749)) + ((g134) & (g251) & (!sk[0]) & (!g660) & (!g704) & (!g749)) + ((g134) & (g251) & (!sk[0]) & (!g660) & (!g704) & (g749)) + ((g134) & (g251) & (!sk[0]) & (!g660) & (g704) & (!g749)) + ((g134) & (g251) & (!sk[0]) & (!g660) & (g704) & (g749)) + ((g134) & (g251) & (!sk[0]) & (g660) & (!g704) & (!g749)) + ((g134) & (g251) & (!sk[0]) & (g660) & (!g704) & (g749)) + ((g134) & (g251) & (!sk[0]) & (g660) & (g704) & (!g749)) + ((g134) & (g251) & (!sk[0]) & (g660) & (g704) & (g749)) + ((g134) & (g251) & (sk[0]) & (!g660) & (!g704) & (g749)) + ((g134) & (g251) & (sk[0]) & (!g660) & (g704) & (g749)) + ((g134) & (g251) & (sk[0]) & (g660) & (!g704) & (g749)) + ((g134) & (g251) & (sk[0]) & (g660) & (g704) & (g749)));
	assign g751 = (((!sk[1]) & (!i_8_) & (!g10) & (!g4) & (!g46) & (g98)) + ((!sk[1]) & (!i_8_) & (!g10) & (!g4) & (g46) & (g98)) + ((!sk[1]) & (!i_8_) & (!g10) & (g4) & (!g46) & (g98)) + ((!sk[1]) & (!i_8_) & (!g10) & (g4) & (g46) & (g98)) + ((!sk[1]) & (!i_8_) & (g10) & (!g4) & (!g46) & (g98)) + ((!sk[1]) & (!i_8_) & (g10) & (!g4) & (g46) & (g98)) + ((!sk[1]) & (!i_8_) & (g10) & (g4) & (!g46) & (g98)) + ((!sk[1]) & (!i_8_) & (g10) & (g4) & (g46) & (g98)) + ((!sk[1]) & (i_8_) & (!g10) & (!g4) & (!g46) & (!g98)) + ((!sk[1]) & (i_8_) & (!g10) & (!g4) & (!g46) & (g98)) + ((!sk[1]) & (i_8_) & (!g10) & (!g4) & (g46) & (!g98)) + ((!sk[1]) & (i_8_) & (!g10) & (!g4) & (g46) & (g98)) + ((!sk[1]) & (i_8_) & (!g10) & (g4) & (!g46) & (!g98)) + ((!sk[1]) & (i_8_) & (!g10) & (g4) & (!g46) & (g98)) + ((!sk[1]) & (i_8_) & (!g10) & (g4) & (g46) & (!g98)) + ((!sk[1]) & (i_8_) & (!g10) & (g4) & (g46) & (g98)) + ((!sk[1]) & (i_8_) & (g10) & (!g4) & (!g46) & (!g98)) + ((!sk[1]) & (i_8_) & (g10) & (!g4) & (!g46) & (g98)) + ((!sk[1]) & (i_8_) & (g10) & (!g4) & (g46) & (!g98)) + ((!sk[1]) & (i_8_) & (g10) & (!g4) & (g46) & (g98)) + ((!sk[1]) & (i_8_) & (g10) & (g4) & (!g46) & (!g98)) + ((!sk[1]) & (i_8_) & (g10) & (g4) & (!g46) & (g98)) + ((!sk[1]) & (i_8_) & (g10) & (g4) & (g46) & (!g98)) + ((!sk[1]) & (i_8_) & (g10) & (g4) & (g46) & (g98)) + ((sk[1]) & (!i_8_) & (g10) & (g4) & (!g46) & (g98)) + ((sk[1]) & (!i_8_) & (g10) & (g4) & (g46) & (g98)) + ((sk[1]) & (i_8_) & (!g10) & (g4) & (g46) & (g98)) + ((sk[1]) & (i_8_) & (g10) & (g4) & (g46) & (g98)));
	assign g752 = (((!g186) & (!sk[2]) & (!g423) & (g702) & (g703)) + ((!g186) & (!sk[2]) & (g423) & (!g702) & (!g703)) + ((!g186) & (!sk[2]) & (g423) & (!g702) & (g703)) + ((!g186) & (!sk[2]) & (g423) & (g702) & (!g703)) + ((!g186) & (!sk[2]) & (g423) & (g702) & (g703)) + ((!g186) & (sk[2]) & (g423) & (g702) & (!g703)) + ((!g186) & (sk[2]) & (g423) & (g702) & (g703)) + ((g186) & (!sk[2]) & (!g423) & (g702) & (!g703)) + ((g186) & (!sk[2]) & (!g423) & (g702) & (g703)) + ((g186) & (!sk[2]) & (g423) & (!g702) & (!g703)) + ((g186) & (!sk[2]) & (g423) & (!g702) & (g703)) + ((g186) & (!sk[2]) & (g423) & (g702) & (!g703)) + ((g186) & (!sk[2]) & (g423) & (g702) & (g703)) + ((g186) & (sk[2]) & (!g423) & (!g702) & (g703)) + ((g186) & (sk[2]) & (!g423) & (g702) & (g703)) + ((g186) & (sk[2]) & (g423) & (!g702) & (g703)) + ((g186) & (sk[2]) & (g423) & (g702) & (!g703)) + ((g186) & (sk[2]) & (g423) & (g702) & (g703)));
	assign g753 = (((!sk[3]) & (g481) & (!g702)) + ((!sk[3]) & (g481) & (g702)) + ((sk[3]) & (g481) & (!g702)));
	assign g754 = (((!i_8_) & (!g88) & (g108) & (!g467) & (!g465) & (!g753)) + ((!i_8_) & (!g88) & (g108) & (!g467) & (!g465) & (g753)) + ((!i_8_) & (!g88) & (g108) & (!g467) & (g465) & (!g753)) + ((!i_8_) & (!g88) & (g108) & (!g467) & (g465) & (g753)) + ((!i_8_) & (g88) & (!g108) & (!g467) & (!g465) & (!g753)) + ((!i_8_) & (g88) & (!g108) & (!g467) & (g465) & (!g753)) + ((!i_8_) & (g88) & (!g108) & (g467) & (!g465) & (!g753)) + ((!i_8_) & (g88) & (!g108) & (g467) & (g465) & (!g753)) + ((!i_8_) & (g88) & (g108) & (!g467) & (!g465) & (!g753)) + ((!i_8_) & (g88) & (g108) & (!g467) & (!g465) & (g753)) + ((!i_8_) & (g88) & (g108) & (!g467) & (g465) & (!g753)) + ((!i_8_) & (g88) & (g108) & (!g467) & (g465) & (g753)) + ((!i_8_) & (g88) & (g108) & (g467) & (!g465) & (!g753)) + ((!i_8_) & (g88) & (g108) & (g467) & (g465) & (!g753)) + ((i_8_) & (g88) & (!g108) & (!g467) & (!g465) & (!g753)) + ((i_8_) & (g88) & (!g108) & (!g467) & (!g465) & (g753)) + ((i_8_) & (g88) & (!g108) & (!g467) & (g465) & (!g753)) + ((i_8_) & (g88) & (!g108) & (!g467) & (g465) & (g753)) + ((i_8_) & (g88) & (!g108) & (g467) & (!g465) & (!g753)) + ((i_8_) & (g88) & (!g108) & (g467) & (!g465) & (g753)) + ((i_8_) & (g88) & (!g108) & (g467) & (g465) & (!g753)) + ((i_8_) & (g88) & (g108) & (!g467) & (!g465) & (!g753)) + ((i_8_) & (g88) & (g108) & (!g467) & (!g465) & (g753)) + ((i_8_) & (g88) & (g108) & (!g467) & (g465) & (!g753)) + ((i_8_) & (g88) & (g108) & (!g467) & (g465) & (g753)) + ((i_8_) & (g88) & (g108) & (g467) & (!g465) & (!g753)) + ((i_8_) & (g88) & (g108) & (g467) & (!g465) & (g753)) + ((i_8_) & (g88) & (g108) & (g467) & (g465) & (!g753)));
	assign g755 = (((!g186) & (!g677) & (!g751) & (!g752) & (!sk[5]) & (g754)) + ((!g186) & (!g677) & (!g751) & (!g752) & (sk[5]) & (!g754)) + ((!g186) & (!g677) & (!g751) & (g752) & (!sk[5]) & (g754)) + ((!g186) & (!g677) & (g751) & (!g752) & (!sk[5]) & (g754)) + ((!g186) & (!g677) & (g751) & (g752) & (!sk[5]) & (g754)) + ((!g186) & (g677) & (!g751) & (!g752) & (!sk[5]) & (g754)) + ((!g186) & (g677) & (!g751) & (!g752) & (sk[5]) & (!g754)) + ((!g186) & (g677) & (!g751) & (g752) & (!sk[5]) & (g754)) + ((!g186) & (g677) & (g751) & (!g752) & (!sk[5]) & (g754)) + ((!g186) & (g677) & (g751) & (g752) & (!sk[5]) & (g754)) + ((g186) & (!g677) & (!g751) & (!g752) & (!sk[5]) & (!g754)) + ((g186) & (!g677) & (!g751) & (!g752) & (!sk[5]) & (g754)) + ((g186) & (!g677) & (!g751) & (!g752) & (sk[5]) & (!g754)) + ((g186) & (!g677) & (!g751) & (g752) & (!sk[5]) & (!g754)) + ((g186) & (!g677) & (!g751) & (g752) & (!sk[5]) & (g754)) + ((g186) & (!g677) & (g751) & (!g752) & (!sk[5]) & (!g754)) + ((g186) & (!g677) & (g751) & (!g752) & (!sk[5]) & (g754)) + ((g186) & (!g677) & (g751) & (g752) & (!sk[5]) & (!g754)) + ((g186) & (!g677) & (g751) & (g752) & (!sk[5]) & (g754)) + ((g186) & (g677) & (!g751) & (!g752) & (!sk[5]) & (!g754)) + ((g186) & (g677) & (!g751) & (!g752) & (!sk[5]) & (g754)) + ((g186) & (g677) & (!g751) & (g752) & (!sk[5]) & (!g754)) + ((g186) & (g677) & (!g751) & (g752) & (!sk[5]) & (g754)) + ((g186) & (g677) & (g751) & (!g752) & (!sk[5]) & (!g754)) + ((g186) & (g677) & (g751) & (!g752) & (!sk[5]) & (g754)) + ((g186) & (g677) & (g751) & (g752) & (!sk[5]) & (!g754)) + ((g186) & (g677) & (g751) & (g752) & (!sk[5]) & (g754)));
	assign g756 = (((!sk[6]) & (g9) & (!g93)) + ((!sk[6]) & (g9) & (g93)) + ((sk[6]) & (g9) & (!g93)));
	assign g757 = (((!g44) & (!g46) & (!g109) & (!g330) & (!g215) & (!g756)) + ((!g44) & (!g46) & (!g109) & (!g330) & (g215) & (!g756)) + ((!g44) & (!g46) & (!g109) & (g330) & (!g215) & (!g756)) + ((!g44) & (!g46) & (!g109) & (g330) & (g215) & (!g756)) + ((!g44) & (!g46) & (!g109) & (g330) & (g215) & (g756)) + ((!g44) & (!g46) & (g109) & (!g330) & (!g215) & (!g756)) + ((!g44) & (!g46) & (g109) & (!g330) & (g215) & (!g756)) + ((!g44) & (!g46) & (g109) & (g330) & (!g215) & (!g756)) + ((!g44) & (!g46) & (g109) & (g330) & (g215) & (!g756)) + ((!g44) & (g46) & (!g109) & (g330) & (!g215) & (!g756)) + ((!g44) & (g46) & (!g109) & (g330) & (g215) & (!g756)) + ((!g44) & (g46) & (!g109) & (g330) & (g215) & (g756)) + ((g44) & (!g46) & (!g109) & (g330) & (!g215) & (!g756)) + ((g44) & (!g46) & (!g109) & (g330) & (g215) & (!g756)) + ((g44) & (!g46) & (!g109) & (g330) & (g215) & (g756)) + ((g44) & (!g46) & (g109) & (g330) & (!g215) & (!g756)) + ((g44) & (!g46) & (g109) & (g330) & (g215) & (!g756)) + ((g44) & (g46) & (!g109) & (g330) & (!g215) & (!g756)) + ((g44) & (g46) & (!g109) & (g330) & (g215) & (!g756)) + ((g44) & (g46) & (!g109) & (g330) & (g215) & (g756)));
	assign g758 = (((!g743) & (!g744) & (g748) & (!g750) & (g755) & (g757)));
	assign g759 = (((g411) & (g694) & (g701) & (g709) & (g742) & (g758)));
	assign g760 = (((!i_8_) & (!g135) & (g481) & (!sk[10]) & (g704)) + ((!i_8_) & (g135) & (!g481) & (!sk[10]) & (!g704)) + ((!i_8_) & (g135) & (!g481) & (!sk[10]) & (g704)) + ((!i_8_) & (g135) & (g481) & (!sk[10]) & (!g704)) + ((!i_8_) & (g135) & (g481) & (!sk[10]) & (g704)) + ((i_8_) & (!g135) & (g481) & (!sk[10]) & (!g704)) + ((i_8_) & (!g135) & (g481) & (!sk[10]) & (g704)) + ((i_8_) & (g135) & (!g481) & (!sk[10]) & (!g704)) + ((i_8_) & (g135) & (!g481) & (!sk[10]) & (g704)) + ((i_8_) & (g135) & (!g481) & (sk[10]) & (!g704)) + ((i_8_) & (g135) & (!g481) & (sk[10]) & (g704)) + ((i_8_) & (g135) & (g481) & (!sk[10]) & (!g704)) + ((i_8_) & (g135) & (g481) & (!sk[10]) & (g704)) + ((i_8_) & (g135) & (g481) & (sk[10]) & (g704)));
	assign g761 = (((!i_8_) & (!g108) & (!sk[11]) & (g702) & (g756)) + ((!i_8_) & (g108) & (!sk[11]) & (!g702) & (!g756)) + ((!i_8_) & (g108) & (!sk[11]) & (!g702) & (g756)) + ((!i_8_) & (g108) & (!sk[11]) & (g702) & (!g756)) + ((!i_8_) & (g108) & (!sk[11]) & (g702) & (g756)) + ((i_8_) & (!g108) & (!sk[11]) & (g702) & (!g756)) + ((i_8_) & (!g108) & (!sk[11]) & (g702) & (g756)) + ((i_8_) & (g108) & (!sk[11]) & (!g702) & (!g756)) + ((i_8_) & (g108) & (!sk[11]) & (!g702) & (g756)) + ((i_8_) & (g108) & (!sk[11]) & (g702) & (!g756)) + ((i_8_) & (g108) & (!sk[11]) & (g702) & (g756)) + ((i_8_) & (g108) & (sk[11]) & (!g702) & (g756)) + ((i_8_) & (g108) & (sk[11]) & (g702) & (!g756)) + ((i_8_) & (g108) & (sk[11]) & (g702) & (g756)));
	assign g762 = (((!i_8_) & (!g135) & (g706) & (!sk[12]) & (g703)) + ((!i_8_) & (g135) & (!g706) & (!sk[12]) & (!g703)) + ((!i_8_) & (g135) & (!g706) & (!sk[12]) & (g703)) + ((!i_8_) & (g135) & (g706) & (!sk[12]) & (!g703)) + ((!i_8_) & (g135) & (g706) & (!sk[12]) & (g703)) + ((i_8_) & (!g135) & (g706) & (!sk[12]) & (!g703)) + ((i_8_) & (!g135) & (g706) & (!sk[12]) & (g703)) + ((i_8_) & (g135) & (!g706) & (!sk[12]) & (!g703)) + ((i_8_) & (g135) & (!g706) & (!sk[12]) & (g703)) + ((i_8_) & (g135) & (!g706) & (sk[12]) & (g703)) + ((i_8_) & (g135) & (g706) & (!sk[12]) & (!g703)) + ((i_8_) & (g135) & (g706) & (!sk[12]) & (g703)) + ((i_8_) & (g135) & (g706) & (sk[12]) & (!g703)) + ((i_8_) & (g135) & (g706) & (sk[12]) & (g703)));
	assign g763 = (((!i_8_) & (!g100) & (!g481) & (!g467) & (!sk[13]) & (g478)) + ((!i_8_) & (!g100) & (!g481) & (g467) & (!sk[13]) & (g478)) + ((!i_8_) & (!g100) & (g481) & (!g467) & (!sk[13]) & (g478)) + ((!i_8_) & (!g100) & (g481) & (g467) & (!sk[13]) & (g478)) + ((!i_8_) & (g100) & (!g481) & (!g467) & (!sk[13]) & (g478)) + ((!i_8_) & (g100) & (!g481) & (g467) & (!sk[13]) & (g478)) + ((!i_8_) & (g100) & (g481) & (!g467) & (!sk[13]) & (g478)) + ((!i_8_) & (g100) & (g481) & (g467) & (!sk[13]) & (g478)) + ((i_8_) & (!g100) & (!g481) & (!g467) & (!sk[13]) & (!g478)) + ((i_8_) & (!g100) & (!g481) & (!g467) & (!sk[13]) & (g478)) + ((i_8_) & (!g100) & (!g481) & (g467) & (!sk[13]) & (!g478)) + ((i_8_) & (!g100) & (!g481) & (g467) & (!sk[13]) & (g478)) + ((i_8_) & (!g100) & (g481) & (!g467) & (!sk[13]) & (!g478)) + ((i_8_) & (!g100) & (g481) & (!g467) & (!sk[13]) & (g478)) + ((i_8_) & (!g100) & (g481) & (g467) & (!sk[13]) & (!g478)) + ((i_8_) & (!g100) & (g481) & (g467) & (!sk[13]) & (g478)) + ((i_8_) & (g100) & (!g481) & (!g467) & (!sk[13]) & (!g478)) + ((i_8_) & (g100) & (!g481) & (!g467) & (!sk[13]) & (g478)) + ((i_8_) & (g100) & (!g481) & (!g467) & (sk[13]) & (!g478)) + ((i_8_) & (g100) & (!g481) & (!g467) & (sk[13]) & (g478)) + ((i_8_) & (g100) & (!g481) & (g467) & (!sk[13]) & (!g478)) + ((i_8_) & (g100) & (!g481) & (g467) & (!sk[13]) & (g478)) + ((i_8_) & (g100) & (!g481) & (g467) & (sk[13]) & (!g478)) + ((i_8_) & (g100) & (!g481) & (g467) & (sk[13]) & (g478)) + ((i_8_) & (g100) & (g481) & (!g467) & (!sk[13]) & (!g478)) + ((i_8_) & (g100) & (g481) & (!g467) & (!sk[13]) & (g478)) + ((i_8_) & (g100) & (g481) & (!g467) & (sk[13]) & (!g478)) + ((i_8_) & (g100) & (g481) & (!g467) & (sk[13]) & (g478)) + ((i_8_) & (g100) & (g481) & (g467) & (!sk[13]) & (!g478)) + ((i_8_) & (g100) & (g481) & (g467) & (!sk[13]) & (g478)) + ((i_8_) & (g100) & (g481) & (g467) & (sk[13]) & (g478)));
	assign g764 = (((!g284) & (!g724) & (!g760) & (!g761) & (!g762) & (!g763)) + ((!g284) & (g724) & (!g760) & (!g761) & (!g762) & (!g763)) + ((g284) & (!g724) & (!g760) & (!g761) & (!g762) & (!g763)));
	assign g765 = (((!g46) & (!g151) & (!g284) & (!g706) & (!g756) & (!g710)) + ((!g46) & (!g151) & (!g284) & (!g706) & (!g756) & (g710)) + ((!g46) & (!g151) & (!g284) & (!g706) & (g756) & (!g710)) + ((!g46) & (!g151) & (!g284) & (!g706) & (g756) & (g710)) + ((!g46) & (!g151) & (!g284) & (g706) & (!g756) & (!g710)) + ((!g46) & (!g151) & (!g284) & (g706) & (!g756) & (g710)) + ((!g46) & (!g151) & (!g284) & (g706) & (g756) & (!g710)) + ((!g46) & (!g151) & (!g284) & (g706) & (g756) & (g710)) + ((!g46) & (!g151) & (g284) & (!g706) & (!g756) & (!g710)) + ((!g46) & (!g151) & (g284) & (!g706) & (g756) & (!g710)) + ((!g46) & (!g151) & (g284) & (g706) & (!g756) & (!g710)) + ((!g46) & (!g151) & (g284) & (g706) & (g756) & (!g710)) + ((!g46) & (g151) & (!g284) & (!g706) & (!g756) & (!g710)) + ((!g46) & (g151) & (g284) & (!g706) & (!g756) & (!g710)) + ((g46) & (!g151) & (!g284) & (!g706) & (!g756) & (!g710)) + ((g46) & (!g151) & (!g284) & (!g706) & (!g756) & (g710)) + ((g46) & (!g151) & (!g284) & (!g706) & (g756) & (!g710)) + ((g46) & (!g151) & (!g284) & (!g706) & (g756) & (g710)) + ((g46) & (!g151) & (!g284) & (g706) & (!g756) & (!g710)) + ((g46) & (!g151) & (!g284) & (g706) & (!g756) & (g710)) + ((g46) & (!g151) & (!g284) & (g706) & (g756) & (!g710)) + ((g46) & (!g151) & (!g284) & (g706) & (g756) & (g710)) + ((g46) & (!g151) & (g284) & (!g706) & (!g756) & (!g710)) + ((g46) & (!g151) & (g284) & (!g706) & (g756) & (!g710)) + ((g46) & (!g151) & (g284) & (g706) & (!g756) & (!g710)) + ((g46) & (!g151) & (g284) & (g706) & (g756) & (!g710)));
	assign g766 = (((!g46) & (!g101) & (!g145) & (!g136) & (!g323) & (!g702)) + ((!g46) & (!g101) & (!g145) & (!g136) & (!g323) & (g702)) + ((!g46) & (!g101) & (!g145) & (!g136) & (g323) & (!g702)) + ((!g46) & (!g101) & (!g145) & (g136) & (!g323) & (!g702)) + ((!g46) & (!g101) & (!g145) & (g136) & (g323) & (!g702)) + ((!g46) & (!g101) & (g145) & (!g136) & (!g323) & (!g702)) + ((!g46) & (!g101) & (g145) & (!g136) & (!g323) & (g702)) + ((!g46) & (!g101) & (g145) & (!g136) & (g323) & (!g702)) + ((!g46) & (!g101) & (g145) & (g136) & (!g323) & (!g702)) + ((!g46) & (!g101) & (g145) & (g136) & (g323) & (!g702)) + ((!g46) & (g101) & (!g145) & (!g136) & (!g323) & (!g702)) + ((!g46) & (g101) & (!g145) & (!g136) & (g323) & (!g702)) + ((!g46) & (g101) & (!g145) & (g136) & (!g323) & (!g702)) + ((!g46) & (g101) & (!g145) & (g136) & (g323) & (!g702)) + ((!g46) & (g101) & (g145) & (!g136) & (!g323) & (!g702)) + ((!g46) & (g101) & (g145) & (!g136) & (g323) & (!g702)) + ((!g46) & (g101) & (g145) & (g136) & (!g323) & (!g702)) + ((!g46) & (g101) & (g145) & (g136) & (g323) & (!g702)) + ((g46) & (!g101) & (!g145) & (!g136) & (!g323) & (!g702)) + ((g46) & (!g101) & (!g145) & (!g136) & (!g323) & (g702)) + ((g46) & (!g101) & (!g145) & (!g136) & (g323) & (!g702)) + ((g46) & (!g101) & (!g145) & (g136) & (!g323) & (!g702)) + ((g46) & (!g101) & (!g145) & (g136) & (g323) & (!g702)) + ((g46) & (g101) & (!g145) & (!g136) & (!g323) & (!g702)) + ((g46) & (g101) & (!g145) & (!g136) & (g323) & (!g702)) + ((g46) & (g101) & (!g145) & (g136) & (!g323) & (!g702)) + ((g46) & (g101) & (!g145) & (g136) & (g323) & (!g702)));
	assign g767 = (((!i_8_) & (!sk[17]) & (!g100) & (g477) & (g706)) + ((!i_8_) & (!sk[17]) & (g100) & (!g477) & (!g706)) + ((!i_8_) & (!sk[17]) & (g100) & (!g477) & (g706)) + ((!i_8_) & (!sk[17]) & (g100) & (g477) & (!g706)) + ((!i_8_) & (!sk[17]) & (g100) & (g477) & (g706)) + ((i_8_) & (!sk[17]) & (!g100) & (g477) & (!g706)) + ((i_8_) & (!sk[17]) & (!g100) & (g477) & (g706)) + ((i_8_) & (!sk[17]) & (g100) & (!g477) & (!g706)) + ((i_8_) & (!sk[17]) & (g100) & (!g477) & (g706)) + ((i_8_) & (!sk[17]) & (g100) & (g477) & (!g706)) + ((i_8_) & (!sk[17]) & (g100) & (g477) & (g706)) + ((i_8_) & (sk[17]) & (g100) & (!g477) & (!g706)) + ((i_8_) & (sk[17]) & (g100) & (!g477) & (g706)) + ((i_8_) & (sk[17]) & (g100) & (g477) & (g706)));
	assign g768 = (((!g112) & (!g702) & (!sk[18]) & (g706) & (g703)) + ((!g112) & (g702) & (!sk[18]) & (!g706) & (!g703)) + ((!g112) & (g702) & (!sk[18]) & (!g706) & (g703)) + ((!g112) & (g702) & (!sk[18]) & (g706) & (!g703)) + ((!g112) & (g702) & (!sk[18]) & (g706) & (g703)) + ((g112) & (!g702) & (!sk[18]) & (g706) & (!g703)) + ((g112) & (!g702) & (!sk[18]) & (g706) & (g703)) + ((g112) & (!g702) & (sk[18]) & (!g706) & (g703)) + ((g112) & (!g702) & (sk[18]) & (g706) & (!g703)) + ((g112) & (!g702) & (sk[18]) & (g706) & (g703)) + ((g112) & (g702) & (!sk[18]) & (!g706) & (!g703)) + ((g112) & (g702) & (!sk[18]) & (!g706) & (g703)) + ((g112) & (g702) & (!sk[18]) & (g706) & (!g703)) + ((g112) & (g702) & (!sk[18]) & (g706) & (g703)) + ((g112) & (g702) & (sk[18]) & (!g706) & (!g703)) + ((g112) & (g702) & (sk[18]) & (!g706) & (g703)) + ((g112) & (g702) & (sk[18]) & (g706) & (!g703)) + ((g112) & (g702) & (sk[18]) & (g706) & (g703)));
	assign g769 = (((!g112) & (!g481) & (!sk[19]) & (g704) & (g710)) + ((!g112) & (g481) & (!sk[19]) & (!g704) & (!g710)) + ((!g112) & (g481) & (!sk[19]) & (!g704) & (g710)) + ((!g112) & (g481) & (!sk[19]) & (g704) & (!g710)) + ((!g112) & (g481) & (!sk[19]) & (g704) & (g710)) + ((g112) & (!g481) & (!sk[19]) & (g704) & (!g710)) + ((g112) & (!g481) & (!sk[19]) & (g704) & (g710)) + ((g112) & (!g481) & (sk[19]) & (!g704) & (!g710)) + ((g112) & (!g481) & (sk[19]) & (!g704) & (g710)) + ((g112) & (!g481) & (sk[19]) & (g704) & (!g710)) + ((g112) & (!g481) & (sk[19]) & (g704) & (g710)) + ((g112) & (g481) & (!sk[19]) & (!g704) & (!g710)) + ((g112) & (g481) & (!sk[19]) & (!g704) & (g710)) + ((g112) & (g481) & (!sk[19]) & (g704) & (!g710)) + ((g112) & (g481) & (!sk[19]) & (g704) & (g710)) + ((g112) & (g481) & (sk[19]) & (!g704) & (g710)) + ((g112) & (g481) & (sk[19]) & (g704) & (!g710)) + ((g112) & (g481) & (sk[19]) & (g704) & (g710)));
	assign g770 = (((!i_8_) & (!g100) & (!sk[20]) & (g703) & (g710)) + ((!i_8_) & (g100) & (!sk[20]) & (!g703) & (!g710)) + ((!i_8_) & (g100) & (!sk[20]) & (!g703) & (g710)) + ((!i_8_) & (g100) & (!sk[20]) & (g703) & (!g710)) + ((!i_8_) & (g100) & (!sk[20]) & (g703) & (g710)) + ((i_8_) & (!g100) & (!sk[20]) & (g703) & (!g710)) + ((i_8_) & (!g100) & (!sk[20]) & (g703) & (g710)) + ((i_8_) & (g100) & (!sk[20]) & (!g703) & (!g710)) + ((i_8_) & (g100) & (!sk[20]) & (!g703) & (g710)) + ((i_8_) & (g100) & (!sk[20]) & (g703) & (!g710)) + ((i_8_) & (g100) & (!sk[20]) & (g703) & (g710)) + ((i_8_) & (g100) & (sk[20]) & (!g703) & (g710)) + ((i_8_) & (g100) & (sk[20]) & (g703) & (!g710)) + ((i_8_) & (g100) & (sk[20]) & (g703) & (g710)));
	assign g771 = (((!i_8_) & (!g44) & (!g100) & (!g323) & (!g703) & (!g756)) + ((!i_8_) & (!g44) & (!g100) & (!g323) & (!g703) & (g756)) + ((!i_8_) & (!g44) & (!g100) & (!g323) & (g703) & (!g756)) + ((!i_8_) & (!g44) & (!g100) & (!g323) & (g703) & (g756)) + ((!i_8_) & (!g44) & (!g100) & (g323) & (!g703) & (!g756)) + ((!i_8_) & (!g44) & (g100) & (!g323) & (!g703) & (!g756)) + ((!i_8_) & (!g44) & (g100) & (!g323) & (!g703) & (g756)) + ((!i_8_) & (!g44) & (g100) & (!g323) & (g703) & (!g756)) + ((!i_8_) & (!g44) & (g100) & (!g323) & (g703) & (g756)) + ((!i_8_) & (!g44) & (g100) & (g323) & (!g703) & (!g756)) + ((!i_8_) & (g44) & (!g100) & (!g323) & (!g703) & (!g756)) + ((!i_8_) & (g44) & (!g100) & (!g323) & (!g703) & (g756)) + ((!i_8_) & (g44) & (!g100) & (!g323) & (g703) & (!g756)) + ((!i_8_) & (g44) & (!g100) & (!g323) & (g703) & (g756)) + ((!i_8_) & (g44) & (g100) & (!g323) & (!g703) & (!g756)) + ((!i_8_) & (g44) & (g100) & (!g323) & (!g703) & (g756)) + ((!i_8_) & (g44) & (g100) & (!g323) & (g703) & (!g756)) + ((!i_8_) & (g44) & (g100) & (!g323) & (g703) & (g756)) + ((i_8_) & (!g44) & (!g100) & (!g323) & (!g703) & (!g756)) + ((i_8_) & (!g44) & (!g100) & (!g323) & (!g703) & (g756)) + ((i_8_) & (!g44) & (!g100) & (!g323) & (g703) & (!g756)) + ((i_8_) & (!g44) & (!g100) & (!g323) & (g703) & (g756)) + ((i_8_) & (!g44) & (!g100) & (g323) & (!g703) & (!g756)) + ((i_8_) & (!g44) & (g100) & (!g323) & (!g703) & (!g756)) + ((i_8_) & (!g44) & (g100) & (!g323) & (g703) & (!g756)) + ((i_8_) & (!g44) & (g100) & (g323) & (!g703) & (!g756)) + ((i_8_) & (g44) & (!g100) & (!g323) & (!g703) & (!g756)) + ((i_8_) & (g44) & (!g100) & (!g323) & (!g703) & (g756)) + ((i_8_) & (g44) & (!g100) & (!g323) & (g703) & (!g756)) + ((i_8_) & (g44) & (!g100) & (!g323) & (g703) & (g756)));
	assign g772 = (((!g767) & (!g768) & (!sk[22]) & (!g769) & (!g770) & (g771)) + ((!g767) & (!g768) & (!sk[22]) & (!g769) & (g770) & (g771)) + ((!g767) & (!g768) & (!sk[22]) & (g769) & (!g770) & (g771)) + ((!g767) & (!g768) & (!sk[22]) & (g769) & (g770) & (g771)) + ((!g767) & (!g768) & (sk[22]) & (!g769) & (!g770) & (g771)) + ((!g767) & (g768) & (!sk[22]) & (!g769) & (!g770) & (g771)) + ((!g767) & (g768) & (!sk[22]) & (!g769) & (g770) & (g771)) + ((!g767) & (g768) & (!sk[22]) & (g769) & (!g770) & (g771)) + ((!g767) & (g768) & (!sk[22]) & (g769) & (g770) & (g771)) + ((g767) & (!g768) & (!sk[22]) & (!g769) & (!g770) & (!g771)) + ((g767) & (!g768) & (!sk[22]) & (!g769) & (!g770) & (g771)) + ((g767) & (!g768) & (!sk[22]) & (!g769) & (g770) & (!g771)) + ((g767) & (!g768) & (!sk[22]) & (!g769) & (g770) & (g771)) + ((g767) & (!g768) & (!sk[22]) & (g769) & (!g770) & (!g771)) + ((g767) & (!g768) & (!sk[22]) & (g769) & (!g770) & (g771)) + ((g767) & (!g768) & (!sk[22]) & (g769) & (g770) & (!g771)) + ((g767) & (!g768) & (!sk[22]) & (g769) & (g770) & (g771)) + ((g767) & (g768) & (!sk[22]) & (!g769) & (!g770) & (!g771)) + ((g767) & (g768) & (!sk[22]) & (!g769) & (!g770) & (g771)) + ((g767) & (g768) & (!sk[22]) & (!g769) & (g770) & (!g771)) + ((g767) & (g768) & (!sk[22]) & (!g769) & (g770) & (g771)) + ((g767) & (g768) & (!sk[22]) & (g769) & (!g770) & (!g771)) + ((g767) & (g768) & (!sk[22]) & (g769) & (!g770) & (g771)) + ((g767) & (g768) & (!sk[22]) & (g769) & (g770) & (!g771)) + ((g767) & (g768) & (!sk[22]) & (g769) & (g770) & (g771)));
	assign g773 = (((!g764) & (!g765) & (!sk[23]) & (g766) & (g772)) + ((!g764) & (g765) & (!sk[23]) & (!g766) & (!g772)) + ((!g764) & (g765) & (!sk[23]) & (!g766) & (g772)) + ((!g764) & (g765) & (!sk[23]) & (g766) & (!g772)) + ((!g764) & (g765) & (!sk[23]) & (g766) & (g772)) + ((g764) & (!g765) & (!sk[23]) & (g766) & (!g772)) + ((g764) & (!g765) & (!sk[23]) & (g766) & (g772)) + ((g764) & (g765) & (!sk[23]) & (!g766) & (!g772)) + ((g764) & (g765) & (!sk[23]) & (!g766) & (g772)) + ((g764) & (g765) & (!sk[23]) & (g766) & (!g772)) + ((g764) & (g765) & (!sk[23]) & (g766) & (g772)) + ((g764) & (g765) & (sk[23]) & (g766) & (g772)));
	assign g774 = (((!g8) & (!g10) & (sk[24]) & (g118)) + ((!g8) & (g10) & (sk[24]) & (g118)) + ((g8) & (!g10) & (!sk[24]) & (!g118)) + ((g8) & (!g10) & (!sk[24]) & (g118)) + ((g8) & (g10) & (!sk[24]) & (!g118)) + ((g8) & (g10) & (!sk[24]) & (g118)) + ((g8) & (g10) & (sk[24]) & (g118)));
	assign g775 = (((!i_8_) & (!g19) & (g23) & (!sk[25]) & (g108)) + ((!i_8_) & (g19) & (!g23) & (!sk[25]) & (!g108)) + ((!i_8_) & (g19) & (!g23) & (!sk[25]) & (g108)) + ((!i_8_) & (g19) & (!g23) & (sk[25]) & (g108)) + ((!i_8_) & (g19) & (g23) & (!sk[25]) & (!g108)) + ((!i_8_) & (g19) & (g23) & (!sk[25]) & (g108)) + ((!i_8_) & (g19) & (g23) & (sk[25]) & (g108)) + ((i_8_) & (!g19) & (g23) & (!sk[25]) & (!g108)) + ((i_8_) & (!g19) & (g23) & (!sk[25]) & (g108)) + ((i_8_) & (!g19) & (g23) & (sk[25]) & (g108)) + ((i_8_) & (g19) & (!g23) & (!sk[25]) & (!g108)) + ((i_8_) & (g19) & (!g23) & (!sk[25]) & (g108)) + ((i_8_) & (g19) & (g23) & (!sk[25]) & (!g108)) + ((i_8_) & (g19) & (g23) & (!sk[25]) & (g108)) + ((i_8_) & (g19) & (g23) & (sk[25]) & (g108)));
	assign g776 = (((!i_9_) & (!g53) & (!g9) & (!g119) & (!sk[26]) & (g214)) + ((!i_9_) & (!g53) & (!g9) & (g119) & (!sk[26]) & (g214)) + ((!i_9_) & (!g53) & (g9) & (!g119) & (!sk[26]) & (g214)) + ((!i_9_) & (!g53) & (g9) & (g119) & (!sk[26]) & (g214)) + ((!i_9_) & (!g53) & (g9) & (g119) & (sk[26]) & (g214)) + ((!i_9_) & (g53) & (!g9) & (!g119) & (!sk[26]) & (g214)) + ((!i_9_) & (g53) & (!g9) & (g119) & (!sk[26]) & (g214)) + ((!i_9_) & (g53) & (g9) & (!g119) & (!sk[26]) & (g214)) + ((!i_9_) & (g53) & (g9) & (g119) & (!sk[26]) & (g214)) + ((!i_9_) & (g53) & (g9) & (g119) & (sk[26]) & (g214)) + ((i_9_) & (!g53) & (!g9) & (!g119) & (!sk[26]) & (!g214)) + ((i_9_) & (!g53) & (!g9) & (!g119) & (!sk[26]) & (g214)) + ((i_9_) & (!g53) & (!g9) & (g119) & (!sk[26]) & (!g214)) + ((i_9_) & (!g53) & (!g9) & (g119) & (!sk[26]) & (g214)) + ((i_9_) & (!g53) & (g9) & (!g119) & (!sk[26]) & (!g214)) + ((i_9_) & (!g53) & (g9) & (!g119) & (!sk[26]) & (g214)) + ((i_9_) & (!g53) & (g9) & (g119) & (!sk[26]) & (!g214)) + ((i_9_) & (!g53) & (g9) & (g119) & (!sk[26]) & (g214)) + ((i_9_) & (!g53) & (g9) & (g119) & (sk[26]) & (g214)) + ((i_9_) & (g53) & (!g9) & (!g119) & (!sk[26]) & (!g214)) + ((i_9_) & (g53) & (!g9) & (!g119) & (!sk[26]) & (g214)) + ((i_9_) & (g53) & (!g9) & (g119) & (!sk[26]) & (!g214)) + ((i_9_) & (g53) & (!g9) & (g119) & (!sk[26]) & (g214)) + ((i_9_) & (g53) & (g9) & (!g119) & (!sk[26]) & (!g214)) + ((i_9_) & (g53) & (g9) & (!g119) & (!sk[26]) & (g214)) + ((i_9_) & (g53) & (g9) & (!g119) & (sk[26]) & (g214)) + ((i_9_) & (g53) & (g9) & (g119) & (!sk[26]) & (!g214)) + ((i_9_) & (g53) & (g9) & (g119) & (!sk[26]) & (g214)) + ((i_9_) & (g53) & (g9) & (g119) & (sk[26]) & (g214)));
	assign g777 = (((!i_8_) & (!sk[27]) & (!g88) & (g423) & (g696)) + ((!i_8_) & (!sk[27]) & (g88) & (!g423) & (!g696)) + ((!i_8_) & (!sk[27]) & (g88) & (!g423) & (g696)) + ((!i_8_) & (!sk[27]) & (g88) & (g423) & (!g696)) + ((!i_8_) & (!sk[27]) & (g88) & (g423) & (g696)) + ((!i_8_) & (sk[27]) & (!g88) & (g423) & (!g696)) + ((!i_8_) & (sk[27]) & (g88) & (!g423) & (!g696)) + ((!i_8_) & (sk[27]) & (g88) & (g423) & (!g696)) + ((i_8_) & (!sk[27]) & (!g88) & (g423) & (!g696)) + ((i_8_) & (!sk[27]) & (!g88) & (g423) & (g696)) + ((i_8_) & (!sk[27]) & (g88) & (!g423) & (!g696)) + ((i_8_) & (!sk[27]) & (g88) & (!g423) & (g696)) + ((i_8_) & (!sk[27]) & (g88) & (g423) & (!g696)) + ((i_8_) & (!sk[27]) & (g88) & (g423) & (g696)) + ((i_8_) & (sk[27]) & (!g88) & (g423) & (!g696)) + ((i_8_) & (sk[27]) & (g88) & (g423) & (!g696)));
	assign g778 = (((!g429) & (!g678) & (!g774) & (!g775) & (!g776) & (!g777)) + ((!g429) & (g678) & (!g774) & (!g775) & (!g776) & (!g777)) + ((g429) & (g678) & (!g774) & (!g775) & (!g776) & (!g777)));
	assign g779 = (((!g134) & (!sk[29]) & (!g696) & (g675) & (g672)) + ((!g134) & (!sk[29]) & (g696) & (!g675) & (!g672)) + ((!g134) & (!sk[29]) & (g696) & (!g675) & (g672)) + ((!g134) & (!sk[29]) & (g696) & (g675) & (!g672)) + ((!g134) & (!sk[29]) & (g696) & (g675) & (g672)) + ((g134) & (!sk[29]) & (!g696) & (g675) & (!g672)) + ((g134) & (!sk[29]) & (!g696) & (g675) & (g672)) + ((g134) & (!sk[29]) & (g696) & (!g675) & (!g672)) + ((g134) & (!sk[29]) & (g696) & (!g675) & (g672)) + ((g134) & (!sk[29]) & (g696) & (g675) & (!g672)) + ((g134) & (!sk[29]) & (g696) & (g675) & (g672)) + ((g134) & (sk[29]) & (!g696) & (!g675) & (!g672)) + ((g134) & (sk[29]) & (!g696) & (!g675) & (g672)) + ((g134) & (sk[29]) & (!g696) & (g675) & (!g672)) + ((g134) & (sk[29]) & (!g696) & (g675) & (g672)) + ((g134) & (sk[29]) & (g696) & (!g675) & (g672)) + ((g134) & (sk[29]) & (g696) & (g675) & (!g672)) + ((g134) & (sk[29]) & (g696) & (g675) & (g672)));
	assign g780 = (((!g19) & (!g16) & (g89) & (!g678) & (!g669) & (!g779)) + ((!g19) & (!g16) & (g89) & (!g678) & (g669) & (!g779)) + ((!g19) & (!g16) & (g89) & (g678) & (!g669) & (!g779)) + ((!g19) & (!g16) & (g89) & (g678) & (g669) & (!g779)) + ((!g19) & (g16) & (!g89) & (g678) & (g669) & (!g779)) + ((!g19) & (g16) & (g89) & (!g678) & (!g669) & (!g779)) + ((!g19) & (g16) & (g89) & (!g678) & (g669) & (!g779)) + ((!g19) & (g16) & (g89) & (g678) & (!g669) & (!g779)) + ((!g19) & (g16) & (g89) & (g678) & (g669) & (!g779)) + ((g19) & (!g16) & (g89) & (!g678) & (!g669) & (!g779)) + ((g19) & (!g16) & (g89) & (!g678) & (g669) & (!g779)) + ((g19) & (!g16) & (g89) & (g678) & (!g669) & (!g779)) + ((g19) & (!g16) & (g89) & (g678) & (g669) & (!g779)) + ((g19) & (g16) & (g89) & (!g678) & (!g669) & (!g779)) + ((g19) & (g16) & (g89) & (!g678) & (g669) & (!g779)) + ((g19) & (g16) & (g89) & (g678) & (!g669) & (!g779)) + ((g19) & (g16) & (g89) & (g678) & (g669) & (!g779)));
	assign g781 = (((!g19) & (!g16) & (sk[31]) & (g134)) + ((g19) & (!g16) & (!sk[31]) & (!g134)) + ((g19) & (!g16) & (!sk[31]) & (g134)) + ((g19) & (!g16) & (sk[31]) & (g134)) + ((g19) & (g16) & (!sk[31]) & (!g134)) + ((g19) & (g16) & (!sk[31]) & (g134)) + ((g19) & (g16) & (sk[31]) & (g134)));
	assign g782 = (((g118) & (!sk[32]) & (!g670) & (!g671)) + ((g118) & (!sk[32]) & (!g670) & (g671)) + ((g118) & (!sk[32]) & (g670) & (!g671)) + ((g118) & (!sk[32]) & (g670) & (g671)) + ((g118) & (sk[32]) & (!g670) & (g671)) + ((g118) & (sk[32]) & (g670) & (!g671)) + ((g118) & (sk[32]) & (g670) & (g671)));
	assign g783 = (((g134) & (!sk[33]) & (!g670) & (!g671)) + ((g134) & (!sk[33]) & (!g670) & (g671)) + ((g134) & (!sk[33]) & (g670) & (!g671)) + ((g134) & (!sk[33]) & (g670) & (g671)) + ((g134) & (sk[33]) & (!g670) & (g671)) + ((g134) & (sk[33]) & (g670) & (!g671)) + ((g134) & (sk[33]) & (g670) & (g671)));
	assign g784 = (((!g8) & (!i_8_) & (!sk[34]) & (g88) & (g675)) + ((!g8) & (!i_8_) & (sk[34]) & (g88) & (!g675)) + ((!g8) & (!i_8_) & (sk[34]) & (g88) & (g675)) + ((!g8) & (i_8_) & (!sk[34]) & (!g88) & (!g675)) + ((!g8) & (i_8_) & (!sk[34]) & (!g88) & (g675)) + ((!g8) & (i_8_) & (!sk[34]) & (g88) & (!g675)) + ((!g8) & (i_8_) & (!sk[34]) & (g88) & (g675)) + ((g8) & (!i_8_) & (!sk[34]) & (g88) & (!g675)) + ((g8) & (!i_8_) & (!sk[34]) & (g88) & (g675)) + ((g8) & (!i_8_) & (sk[34]) & (g88) & (g675)) + ((g8) & (i_8_) & (!sk[34]) & (!g88) & (!g675)) + ((g8) & (i_8_) & (!sk[34]) & (!g88) & (g675)) + ((g8) & (i_8_) & (!sk[34]) & (g88) & (!g675)) + ((g8) & (i_8_) & (!sk[34]) & (g88) & (g675)));
	assign g785 = (((!g8) & (!i_8_) & (g108) & (!g678) & (!g670) & (!g671)) + ((!g8) & (!i_8_) & (g108) & (!g678) & (!g670) & (g671)) + ((!g8) & (!i_8_) & (g108) & (!g678) & (g670) & (!g671)) + ((!g8) & (!i_8_) & (g108) & (!g678) & (g670) & (g671)) + ((!g8) & (!i_8_) & (g108) & (g678) & (!g670) & (!g671)) + ((!g8) & (!i_8_) & (g108) & (g678) & (!g670) & (g671)) + ((!g8) & (!i_8_) & (g108) & (g678) & (g670) & (!g671)) + ((!g8) & (!i_8_) & (g108) & (g678) & (g670) & (g671)) + ((g8) & (!i_8_) & (g108) & (!g678) & (!g670) & (!g671)) + ((g8) & (!i_8_) & (g108) & (!g678) & (!g670) & (g671)) + ((g8) & (!i_8_) & (g108) & (!g678) & (g670) & (!g671)) + ((g8) & (!i_8_) & (g108) & (!g678) & (g670) & (g671)) + ((g8) & (!i_8_) & (g108) & (g678) & (!g670) & (g671)) + ((g8) & (!i_8_) & (g108) & (g678) & (g670) & (!g671)) + ((g8) & (!i_8_) & (g108) & (g678) & (g670) & (g671)));
	assign g786 = (((!g781) & (!g782) & (!sk[36]) & (!g783) & (!g784) & (g785)) + ((!g781) & (!g782) & (!sk[36]) & (!g783) & (g784) & (g785)) + ((!g781) & (!g782) & (!sk[36]) & (g783) & (!g784) & (g785)) + ((!g781) & (!g782) & (!sk[36]) & (g783) & (g784) & (g785)) + ((!g781) & (!g782) & (sk[36]) & (!g783) & (!g784) & (!g785)) + ((!g781) & (g782) & (!sk[36]) & (!g783) & (!g784) & (g785)) + ((!g781) & (g782) & (!sk[36]) & (!g783) & (g784) & (g785)) + ((!g781) & (g782) & (!sk[36]) & (g783) & (!g784) & (g785)) + ((!g781) & (g782) & (!sk[36]) & (g783) & (g784) & (g785)) + ((g781) & (!g782) & (!sk[36]) & (!g783) & (!g784) & (!g785)) + ((g781) & (!g782) & (!sk[36]) & (!g783) & (!g784) & (g785)) + ((g781) & (!g782) & (!sk[36]) & (!g783) & (g784) & (!g785)) + ((g781) & (!g782) & (!sk[36]) & (!g783) & (g784) & (g785)) + ((g781) & (!g782) & (!sk[36]) & (g783) & (!g784) & (!g785)) + ((g781) & (!g782) & (!sk[36]) & (g783) & (!g784) & (g785)) + ((g781) & (!g782) & (!sk[36]) & (g783) & (g784) & (!g785)) + ((g781) & (!g782) & (!sk[36]) & (g783) & (g784) & (g785)) + ((g781) & (g782) & (!sk[36]) & (!g783) & (!g784) & (!g785)) + ((g781) & (g782) & (!sk[36]) & (!g783) & (!g784) & (g785)) + ((g781) & (g782) & (!sk[36]) & (!g783) & (g784) & (!g785)) + ((g781) & (g782) & (!sk[36]) & (!g783) & (g784) & (g785)) + ((g781) & (g782) & (!sk[36]) & (g783) & (!g784) & (!g785)) + ((g781) & (g782) & (!sk[36]) & (g783) & (!g784) & (g785)) + ((g781) & (g782) & (!sk[36]) & (g783) & (g784) & (!g785)) + ((g781) & (g782) & (!sk[36]) & (g783) & (g784) & (g785)));
	assign g787 = (((!g10) & (sk[37]) & (g12) & (g134)) + ((g10) & (!sk[37]) & (!g12) & (!g134)) + ((g10) & (!sk[37]) & (!g12) & (g134)) + ((g10) & (!sk[37]) & (g12) & (!g134)) + ((g10) & (!sk[37]) & (g12) & (g134)) + ((g10) & (sk[37]) & (!g12) & (g134)) + ((g10) & (sk[37]) & (g12) & (g134)));
	assign g788 = (((!sk[38]) & (g12) & (!g16) & (!g99)) + ((!sk[38]) & (g12) & (!g16) & (g99)) + ((!sk[38]) & (g12) & (g16) & (!g99)) + ((!sk[38]) & (g12) & (g16) & (g99)) + ((sk[38]) & (!g12) & (!g16) & (g99)) + ((sk[38]) & (g12) & (!g16) & (g99)) + ((sk[38]) & (g12) & (g16) & (g99)));
	assign g789 = (((!g23) & (g88) & (sk[39]) & (g734)) + ((g23) & (!g88) & (!sk[39]) & (!g734)) + ((g23) & (!g88) & (!sk[39]) & (g734)) + ((g23) & (g88) & (!sk[39]) & (!g734)) + ((g23) & (g88) & (!sk[39]) & (g734)) + ((g23) & (g88) & (sk[39]) & (!g734)) + ((g23) & (g88) & (sk[39]) & (g734)));
	assign g790 = (((!g23) & (g112) & (sk[40]) & (g734)) + ((g23) & (!g112) & (!sk[40]) & (!g734)) + ((g23) & (!g112) & (!sk[40]) & (g734)) + ((g23) & (g112) & (!sk[40]) & (!g734)) + ((g23) & (g112) & (!sk[40]) & (g734)) + ((g23) & (g112) & (sk[40]) & (!g734)) + ((g23) & (g112) & (sk[40]) & (g734)));
	assign g791 = (((!i_8_) & (!g108) & (g734) & (!sk[41]) & (g669)) + ((!i_8_) & (g108) & (!g734) & (!sk[41]) & (!g669)) + ((!i_8_) & (g108) & (!g734) & (!sk[41]) & (g669)) + ((!i_8_) & (g108) & (!g734) & (sk[41]) & (!g669)) + ((!i_8_) & (g108) & (g734) & (!sk[41]) & (!g669)) + ((!i_8_) & (g108) & (g734) & (!sk[41]) & (g669)) + ((!i_8_) & (g108) & (g734) & (sk[41]) & (!g669)) + ((!i_8_) & (g108) & (g734) & (sk[41]) & (g669)) + ((i_8_) & (!g108) & (g734) & (!sk[41]) & (!g669)) + ((i_8_) & (!g108) & (g734) & (!sk[41]) & (g669)) + ((i_8_) & (g108) & (!g734) & (!sk[41]) & (!g669)) + ((i_8_) & (g108) & (!g734) & (!sk[41]) & (g669)) + ((i_8_) & (g108) & (g734) & (!sk[41]) & (!g669)) + ((i_8_) & (g108) & (g734) & (!sk[41]) & (g669)) + ((i_8_) & (g108) & (g734) & (sk[41]) & (!g669)) + ((i_8_) & (g108) & (g734) & (sk[41]) & (g669)));
	assign g792 = (((!i_8_) & (!g135) & (!sk[42]) & (g734) & (g675)) + ((!i_8_) & (g135) & (!sk[42]) & (!g734) & (!g675)) + ((!i_8_) & (g135) & (!sk[42]) & (!g734) & (g675)) + ((!i_8_) & (g135) & (!sk[42]) & (g734) & (!g675)) + ((!i_8_) & (g135) & (!sk[42]) & (g734) & (g675)) + ((i_8_) & (!g135) & (!sk[42]) & (g734) & (!g675)) + ((i_8_) & (!g135) & (!sk[42]) & (g734) & (g675)) + ((i_8_) & (g135) & (!sk[42]) & (!g734) & (!g675)) + ((i_8_) & (g135) & (!sk[42]) & (!g734) & (g675)) + ((i_8_) & (g135) & (!sk[42]) & (g734) & (!g675)) + ((i_8_) & (g135) & (!sk[42]) & (g734) & (g675)) + ((i_8_) & (g135) & (sk[42]) & (!g734) & (g675)) + ((i_8_) & (g135) & (sk[42]) & (g734) & (!g675)) + ((i_8_) & (g135) & (sk[42]) & (g734) & (g675)));
	assign g793 = (((!g787) & (!g788) & (!g789) & (!g790) & (!g791) & (!g792)));
	assign g794 = (((!g99) & (!g696) & (!sk[44]) & (g670) & (g672)) + ((!g99) & (g696) & (!sk[44]) & (!g670) & (!g672)) + ((!g99) & (g696) & (!sk[44]) & (!g670) & (g672)) + ((!g99) & (g696) & (!sk[44]) & (g670) & (!g672)) + ((!g99) & (g696) & (!sk[44]) & (g670) & (g672)) + ((g99) & (!g696) & (!sk[44]) & (g670) & (!g672)) + ((g99) & (!g696) & (!sk[44]) & (g670) & (g672)) + ((g99) & (!g696) & (sk[44]) & (!g670) & (!g672)) + ((g99) & (!g696) & (sk[44]) & (!g670) & (g672)) + ((g99) & (!g696) & (sk[44]) & (g670) & (!g672)) + ((g99) & (!g696) & (sk[44]) & (g670) & (g672)) + ((g99) & (g696) & (!sk[44]) & (!g670) & (!g672)) + ((g99) & (g696) & (!sk[44]) & (!g670) & (g672)) + ((g99) & (g696) & (!sk[44]) & (g670) & (!g672)) + ((g99) & (g696) & (!sk[44]) & (g670) & (g672)) + ((g99) & (g696) & (sk[44]) & (!g670) & (g672)) + ((g99) & (g696) & (sk[44]) & (g670) & (!g672)) + ((g99) & (g696) & (sk[44]) & (g670) & (g672)));
	assign g795 = (((!sk[45]) & (!g10) & (!g16) & (g59) & (g678)) + ((!sk[45]) & (!g10) & (g16) & (!g59) & (!g678)) + ((!sk[45]) & (!g10) & (g16) & (!g59) & (g678)) + ((!sk[45]) & (!g10) & (g16) & (g59) & (!g678)) + ((!sk[45]) & (!g10) & (g16) & (g59) & (g678)) + ((!sk[45]) & (g10) & (!g16) & (g59) & (!g678)) + ((!sk[45]) & (g10) & (!g16) & (g59) & (g678)) + ((!sk[45]) & (g10) & (g16) & (!g59) & (!g678)) + ((!sk[45]) & (g10) & (g16) & (!g59) & (g678)) + ((!sk[45]) & (g10) & (g16) & (g59) & (!g678)) + ((!sk[45]) & (g10) & (g16) & (g59) & (g678)) + ((sk[45]) & (!g10) & (!g16) & (g59) & (!g678)) + ((sk[45]) & (!g10) & (!g16) & (g59) & (g678)) + ((sk[45]) & (!g10) & (g16) & (g59) & (!g678)) + ((sk[45]) & (g10) & (!g16) & (g59) & (!g678)) + ((sk[45]) & (g10) & (!g16) & (g59) & (g678)) + ((sk[45]) & (g10) & (g16) & (g59) & (!g678)) + ((sk[45]) & (g10) & (g16) & (g59) & (g678)));
	assign g796 = (((!g8) & (!g23) & (g134) & (!sk[46]) & (g669)) + ((!g8) & (!g23) & (g134) & (sk[46]) & (!g669)) + ((!g8) & (!g23) & (g134) & (sk[46]) & (g669)) + ((!g8) & (g23) & (!g134) & (!sk[46]) & (!g669)) + ((!g8) & (g23) & (!g134) & (!sk[46]) & (g669)) + ((!g8) & (g23) & (g134) & (!sk[46]) & (!g669)) + ((!g8) & (g23) & (g134) & (!sk[46]) & (g669)) + ((!g8) & (g23) & (g134) & (sk[46]) & (!g669)) + ((!g8) & (g23) & (g134) & (sk[46]) & (g669)) + ((g8) & (!g23) & (g134) & (!sk[46]) & (!g669)) + ((g8) & (!g23) & (g134) & (!sk[46]) & (g669)) + ((g8) & (!g23) & (g134) & (sk[46]) & (!g669)) + ((g8) & (g23) & (!g134) & (!sk[46]) & (!g669)) + ((g8) & (g23) & (!g134) & (!sk[46]) & (g669)) + ((g8) & (g23) & (g134) & (!sk[46]) & (!g669)) + ((g8) & (g23) & (g134) & (!sk[46]) & (g669)) + ((g8) & (g23) & (g134) & (sk[46]) & (!g669)) + ((g8) & (g23) & (g134) & (sk[46]) & (g669)));
	assign g797 = (((!sk[47]) & (i_9_) & (!g53) & (!g9)) + ((!sk[47]) & (i_9_) & (!g53) & (g9)) + ((!sk[47]) & (i_9_) & (g53) & (!g9)) + ((!sk[47]) & (i_9_) & (g53) & (g9)) + ((sk[47]) & (!i_9_) & (g53) & (g9)));
	assign g798 = (((!g12) & (!g118) & (!sk[48]) & (g696) & (g797)) + ((!g12) & (g118) & (!sk[48]) & (!g696) & (!g797)) + ((!g12) & (g118) & (!sk[48]) & (!g696) & (g797)) + ((!g12) & (g118) & (!sk[48]) & (g696) & (!g797)) + ((!g12) & (g118) & (!sk[48]) & (g696) & (g797)) + ((!g12) & (g118) & (sk[48]) & (!g696) & (!g797)) + ((!g12) & (g118) & (sk[48]) & (!g696) & (g797)) + ((!g12) & (g118) & (sk[48]) & (g696) & (g797)) + ((g12) & (!g118) & (!sk[48]) & (g696) & (!g797)) + ((g12) & (!g118) & (!sk[48]) & (g696) & (g797)) + ((g12) & (g118) & (!sk[48]) & (!g696) & (!g797)) + ((g12) & (g118) & (!sk[48]) & (!g696) & (g797)) + ((g12) & (g118) & (!sk[48]) & (g696) & (!g797)) + ((g12) & (g118) & (!sk[48]) & (g696) & (g797)) + ((g12) & (g118) & (sk[48]) & (!g696) & (!g797)) + ((g12) & (g118) & (sk[48]) & (!g696) & (g797)) + ((g12) & (g118) & (sk[48]) & (g696) & (!g797)) + ((g12) & (g118) & (sk[48]) & (g696) & (g797)));
	assign g799 = (((!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g7) & (g118)) + ((!i_11_) & (i_9_) & (i_10_) & (i_15_) & (g7) & (g118)) + ((i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (g7) & (g118)) + ((i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g7) & (g118)) + ((i_11_) & (i_9_) & (i_10_) & (i_15_) & (g7) & (g118)));
	assign g800 = (((!g794) & (!sk[50]) & (!g795) & (!g796) & (!g798) & (g799)) + ((!g794) & (!sk[50]) & (!g795) & (!g796) & (g798) & (g799)) + ((!g794) & (!sk[50]) & (!g795) & (g796) & (!g798) & (g799)) + ((!g794) & (!sk[50]) & (!g795) & (g796) & (g798) & (g799)) + ((!g794) & (!sk[50]) & (g795) & (!g796) & (!g798) & (g799)) + ((!g794) & (!sk[50]) & (g795) & (!g796) & (g798) & (g799)) + ((!g794) & (!sk[50]) & (g795) & (g796) & (!g798) & (g799)) + ((!g794) & (!sk[50]) & (g795) & (g796) & (g798) & (g799)) + ((!g794) & (sk[50]) & (!g795) & (!g796) & (!g798) & (!g799)) + ((g794) & (!sk[50]) & (!g795) & (!g796) & (!g798) & (!g799)) + ((g794) & (!sk[50]) & (!g795) & (!g796) & (!g798) & (g799)) + ((g794) & (!sk[50]) & (!g795) & (!g796) & (g798) & (!g799)) + ((g794) & (!sk[50]) & (!g795) & (!g796) & (g798) & (g799)) + ((g794) & (!sk[50]) & (!g795) & (g796) & (!g798) & (!g799)) + ((g794) & (!sk[50]) & (!g795) & (g796) & (!g798) & (g799)) + ((g794) & (!sk[50]) & (!g795) & (g796) & (g798) & (!g799)) + ((g794) & (!sk[50]) & (!g795) & (g796) & (g798) & (g799)) + ((g794) & (!sk[50]) & (g795) & (!g796) & (!g798) & (!g799)) + ((g794) & (!sk[50]) & (g795) & (!g796) & (!g798) & (g799)) + ((g794) & (!sk[50]) & (g795) & (!g796) & (g798) & (!g799)) + ((g794) & (!sk[50]) & (g795) & (!g796) & (g798) & (g799)) + ((g794) & (!sk[50]) & (g795) & (g796) & (!g798) & (!g799)) + ((g794) & (!sk[50]) & (g795) & (g796) & (!g798) & (g799)) + ((g794) & (!sk[50]) & (g795) & (g796) & (g798) & (!g799)) + ((g794) & (!sk[50]) & (g795) & (g796) & (g798) & (g799)));
	assign g801 = (((!sk[51]) & (g676) & (!g677)) + ((!sk[51]) & (g676) & (g677)) + ((sk[51]) & (!g676) & (!g677)));
	assign g802 = (((!g23) & (!g12) & (g109) & (!g675) & (!g672) & (!g801)) + ((!g23) & (!g12) & (g109) & (!g675) & (g672) & (!g801)) + ((!g23) & (!g12) & (g109) & (!g675) & (g672) & (g801)) + ((!g23) & (!g12) & (g109) & (g675) & (!g672) & (!g801)) + ((!g23) & (!g12) & (g109) & (g675) & (!g672) & (g801)) + ((!g23) & (!g12) & (g109) & (g675) & (g672) & (!g801)) + ((!g23) & (!g12) & (g109) & (g675) & (g672) & (g801)) + ((!g23) & (g12) & (g109) & (!g675) & (!g672) & (!g801)) + ((!g23) & (g12) & (g109) & (!g675) & (!g672) & (g801)) + ((!g23) & (g12) & (g109) & (!g675) & (g672) & (!g801)) + ((!g23) & (g12) & (g109) & (!g675) & (g672) & (g801)) + ((!g23) & (g12) & (g109) & (g675) & (!g672) & (!g801)) + ((!g23) & (g12) & (g109) & (g675) & (!g672) & (g801)) + ((!g23) & (g12) & (g109) & (g675) & (g672) & (!g801)) + ((!g23) & (g12) & (g109) & (g675) & (g672) & (g801)) + ((g23) & (!g12) & (g109) & (!g675) & (!g672) & (!g801)) + ((g23) & (!g12) & (g109) & (!g675) & (!g672) & (g801)) + ((g23) & (!g12) & (g109) & (!g675) & (g672) & (!g801)) + ((g23) & (!g12) & (g109) & (!g675) & (g672) & (g801)) + ((g23) & (!g12) & (g109) & (g675) & (!g672) & (!g801)) + ((g23) & (!g12) & (g109) & (g675) & (!g672) & (g801)) + ((g23) & (!g12) & (g109) & (g675) & (g672) & (!g801)) + ((g23) & (!g12) & (g109) & (g675) & (g672) & (g801)) + ((g23) & (g12) & (g109) & (!g675) & (!g672) & (!g801)) + ((g23) & (g12) & (g109) & (!g675) & (!g672) & (g801)) + ((g23) & (g12) & (g109) & (!g675) & (g672) & (!g801)) + ((g23) & (g12) & (g109) & (!g675) & (g672) & (g801)) + ((g23) & (g12) & (g109) & (g675) & (!g672) & (!g801)) + ((g23) & (g12) & (g109) & (g675) & (!g672) & (g801)) + ((g23) & (g12) & (g109) & (g675) & (g672) & (!g801)) + ((g23) & (g12) & (g109) & (g675) & (g672) & (g801)));
	assign g803 = (((g778) & (g780) & (g786) & (g793) & (g800) & (!g802)));
	assign g804 = (((!g21) & (!g112) & (g127) & (!sk[54]) & (g506)) + ((!g21) & (g112) & (!g127) & (!sk[54]) & (!g506)) + ((!g21) & (g112) & (!g127) & (!sk[54]) & (g506)) + ((!g21) & (g112) & (!g127) & (sk[54]) & (!g506)) + ((!g21) & (g112) & (!g127) & (sk[54]) & (g506)) + ((!g21) & (g112) & (g127) & (!sk[54]) & (!g506)) + ((!g21) & (g112) & (g127) & (!sk[54]) & (g506)) + ((!g21) & (g112) & (g127) & (sk[54]) & (g506)) + ((g21) & (!g112) & (g127) & (!sk[54]) & (!g506)) + ((g21) & (!g112) & (g127) & (!sk[54]) & (g506)) + ((g21) & (g112) & (!g127) & (!sk[54]) & (!g506)) + ((g21) & (g112) & (!g127) & (!sk[54]) & (g506)) + ((g21) & (g112) & (!g127) & (sk[54]) & (!g506)) + ((g21) & (g112) & (!g127) & (sk[54]) & (g506)) + ((g21) & (g112) & (g127) & (!sk[54]) & (!g506)) + ((g21) & (g112) & (g127) & (!sk[54]) & (g506)) + ((g21) & (g112) & (g127) & (sk[54]) & (!g506)) + ((g21) & (g112) & (g127) & (sk[54]) & (g506)));
	assign g805 = (((!sk[55]) & (g20) & (!g59)) + ((!sk[55]) & (g20) & (g59)) + ((sk[55]) & (!g20) & (g59)));
	assign g806 = (((!sk[56]) & (g18) & (!g711)) + ((!sk[56]) & (g18) & (g711)) + ((sk[56]) & (!g18) & (g711)));
	assign g807 = (((!sk[57]) & (g20) & (!g806)) + ((!sk[57]) & (g20) & (g806)) + ((sk[57]) & (g20) & (!g806)));
	assign g808 = (((!sk[58]) & (!i_8_) & (!g20) & (g21) & (g135)) + ((!sk[58]) & (!i_8_) & (g20) & (!g21) & (!g135)) + ((!sk[58]) & (!i_8_) & (g20) & (!g21) & (g135)) + ((!sk[58]) & (!i_8_) & (g20) & (g21) & (!g135)) + ((!sk[58]) & (!i_8_) & (g20) & (g21) & (g135)) + ((!sk[58]) & (i_8_) & (!g20) & (g21) & (!g135)) + ((!sk[58]) & (i_8_) & (!g20) & (g21) & (g135)) + ((!sk[58]) & (i_8_) & (g20) & (!g21) & (!g135)) + ((!sk[58]) & (i_8_) & (g20) & (!g21) & (g135)) + ((!sk[58]) & (i_8_) & (g20) & (g21) & (!g135)) + ((!sk[58]) & (i_8_) & (g20) & (g21) & (g135)) + ((sk[58]) & (!i_8_) & (!g20) & (!g21) & (g135)) + ((sk[58]) & (!i_8_) & (!g20) & (g21) & (g135)) + ((sk[58]) & (i_8_) & (!g20) & (!g21) & (g135)) + ((sk[58]) & (i_8_) & (!g20) & (g21) & (g135)) + ((sk[58]) & (i_8_) & (g20) & (g21) & (g135)));
	assign g809 = (((!g20) & (!g16) & (!g118) & (sk[59]) & (g423)) + ((!g20) & (!g16) & (g118) & (!sk[59]) & (g423)) + ((!g20) & (!g16) & (g118) & (sk[59]) & (!g423)) + ((!g20) & (!g16) & (g118) & (sk[59]) & (g423)) + ((!g20) & (g16) & (!g118) & (!sk[59]) & (!g423)) + ((!g20) & (g16) & (!g118) & (!sk[59]) & (g423)) + ((!g20) & (g16) & (g118) & (!sk[59]) & (!g423)) + ((!g20) & (g16) & (g118) & (!sk[59]) & (g423)) + ((!g20) & (g16) & (g118) & (sk[59]) & (!g423)) + ((!g20) & (g16) & (g118) & (sk[59]) & (g423)) + ((g20) & (!g16) & (!g118) & (sk[59]) & (g423)) + ((g20) & (!g16) & (g118) & (!sk[59]) & (!g423)) + ((g20) & (!g16) & (g118) & (!sk[59]) & (g423)) + ((g20) & (!g16) & (g118) & (sk[59]) & (g423)) + ((g20) & (g16) & (!g118) & (!sk[59]) & (!g423)) + ((g20) & (g16) & (!g118) & (!sk[59]) & (g423)) + ((g20) & (g16) & (g118) & (!sk[59]) & (!g423)) + ((g20) & (g16) & (g118) & (!sk[59]) & (g423)));
	assign g810 = (((!g136) & (!g127) & (!g506) & (!g808) & (!sk[60]) & (g809)) + ((!g136) & (!g127) & (!g506) & (!g808) & (sk[60]) & (!g809)) + ((!g136) & (!g127) & (!g506) & (g808) & (!sk[60]) & (g809)) + ((!g136) & (!g127) & (g506) & (!g808) & (!sk[60]) & (g809)) + ((!g136) & (!g127) & (g506) & (!g808) & (sk[60]) & (!g809)) + ((!g136) & (!g127) & (g506) & (g808) & (!sk[60]) & (g809)) + ((!g136) & (g127) & (!g506) & (!g808) & (!sk[60]) & (g809)) + ((!g136) & (g127) & (!g506) & (!g808) & (sk[60]) & (!g809)) + ((!g136) & (g127) & (!g506) & (g808) & (!sk[60]) & (g809)) + ((!g136) & (g127) & (g506) & (!g808) & (!sk[60]) & (g809)) + ((!g136) & (g127) & (g506) & (!g808) & (sk[60]) & (!g809)) + ((!g136) & (g127) & (g506) & (g808) & (!sk[60]) & (g809)) + ((g136) & (!g127) & (!g506) & (!g808) & (!sk[60]) & (!g809)) + ((g136) & (!g127) & (!g506) & (!g808) & (!sk[60]) & (g809)) + ((g136) & (!g127) & (!g506) & (g808) & (!sk[60]) & (!g809)) + ((g136) & (!g127) & (!g506) & (g808) & (!sk[60]) & (g809)) + ((g136) & (!g127) & (g506) & (!g808) & (!sk[60]) & (!g809)) + ((g136) & (!g127) & (g506) & (!g808) & (!sk[60]) & (g809)) + ((g136) & (!g127) & (g506) & (g808) & (!sk[60]) & (!g809)) + ((g136) & (!g127) & (g506) & (g808) & (!sk[60]) & (g809)) + ((g136) & (g127) & (!g506) & (!g808) & (!sk[60]) & (!g809)) + ((g136) & (g127) & (!g506) & (!g808) & (!sk[60]) & (g809)) + ((g136) & (g127) & (!g506) & (!g808) & (sk[60]) & (!g809)) + ((g136) & (g127) & (!g506) & (g808) & (!sk[60]) & (!g809)) + ((g136) & (g127) & (!g506) & (g808) & (!sk[60]) & (g809)) + ((g136) & (g127) & (g506) & (!g808) & (!sk[60]) & (!g809)) + ((g136) & (g127) & (g506) & (!g808) & (!sk[60]) & (g809)) + ((g136) & (g127) & (g506) & (g808) & (!sk[60]) & (!g809)) + ((g136) & (g127) & (g506) & (g808) & (!sk[60]) & (g809)));
	assign g811 = (((!g6) & (!i_15_) & (!sk[61]) & (!i_14_) & (!i_12_) & (i_13_)) + ((!g6) & (!i_15_) & (!sk[61]) & (!i_14_) & (i_12_) & (i_13_)) + ((!g6) & (!i_15_) & (!sk[61]) & (i_14_) & (!i_12_) & (i_13_)) + ((!g6) & (!i_15_) & (!sk[61]) & (i_14_) & (i_12_) & (i_13_)) + ((!g6) & (i_15_) & (!sk[61]) & (!i_14_) & (!i_12_) & (i_13_)) + ((!g6) & (i_15_) & (!sk[61]) & (!i_14_) & (i_12_) & (i_13_)) + ((!g6) & (i_15_) & (!sk[61]) & (i_14_) & (!i_12_) & (i_13_)) + ((!g6) & (i_15_) & (!sk[61]) & (i_14_) & (i_12_) & (i_13_)) + ((g6) & (!i_15_) & (!sk[61]) & (!i_14_) & (!i_12_) & (!i_13_)) + ((g6) & (!i_15_) & (!sk[61]) & (!i_14_) & (!i_12_) & (i_13_)) + ((g6) & (!i_15_) & (!sk[61]) & (!i_14_) & (i_12_) & (!i_13_)) + ((g6) & (!i_15_) & (!sk[61]) & (!i_14_) & (i_12_) & (i_13_)) + ((g6) & (!i_15_) & (!sk[61]) & (i_14_) & (!i_12_) & (!i_13_)) + ((g6) & (!i_15_) & (!sk[61]) & (i_14_) & (!i_12_) & (i_13_)) + ((g6) & (!i_15_) & (!sk[61]) & (i_14_) & (i_12_) & (!i_13_)) + ((g6) & (!i_15_) & (!sk[61]) & (i_14_) & (i_12_) & (i_13_)) + ((g6) & (!i_15_) & (sk[61]) & (i_14_) & (!i_12_) & (!i_13_)) + ((g6) & (!i_15_) & (sk[61]) & (i_14_) & (!i_12_) & (i_13_)) + ((g6) & (i_15_) & (!sk[61]) & (!i_14_) & (!i_12_) & (!i_13_)) + ((g6) & (i_15_) & (!sk[61]) & (!i_14_) & (!i_12_) & (i_13_)) + ((g6) & (i_15_) & (!sk[61]) & (!i_14_) & (i_12_) & (!i_13_)) + ((g6) & (i_15_) & (!sk[61]) & (!i_14_) & (i_12_) & (i_13_)) + ((g6) & (i_15_) & (!sk[61]) & (i_14_) & (!i_12_) & (!i_13_)) + ((g6) & (i_15_) & (!sk[61]) & (i_14_) & (!i_12_) & (i_13_)) + ((g6) & (i_15_) & (!sk[61]) & (i_14_) & (i_12_) & (!i_13_)) + ((g6) & (i_15_) & (!sk[61]) & (i_14_) & (i_12_) & (i_13_)) + ((g6) & (i_15_) & (sk[61]) & (!i_14_) & (i_12_) & (i_13_)));
	assign g812 = (((!g186) & (!sk[62]) & (!g122) & (g280) & (g711)) + ((!g186) & (!sk[62]) & (g122) & (!g280) & (!g711)) + ((!g186) & (!sk[62]) & (g122) & (!g280) & (g711)) + ((!g186) & (!sk[62]) & (g122) & (g280) & (!g711)) + ((!g186) & (!sk[62]) & (g122) & (g280) & (g711)) + ((g186) & (!sk[62]) & (!g122) & (g280) & (!g711)) + ((g186) & (!sk[62]) & (!g122) & (g280) & (g711)) + ((g186) & (!sk[62]) & (g122) & (!g280) & (!g711)) + ((g186) & (!sk[62]) & (g122) & (!g280) & (g711)) + ((g186) & (!sk[62]) & (g122) & (g280) & (!g711)) + ((g186) & (!sk[62]) & (g122) & (g280) & (g711)) + ((g186) & (sk[62]) & (!g122) & (!g280) & (g711)) + ((g186) & (sk[62]) & (!g122) & (g280) & (!g711)) + ((g186) & (sk[62]) & (!g122) & (g280) & (g711)) + ((g186) & (sk[62]) & (g122) & (g280) & (!g711)) + ((g186) & (sk[62]) & (g122) & (g280) & (g711)));
	assign g813 = (((i_14_) & (!sk[63]) & (!i_12_) & (!g95)) + ((i_14_) & (!sk[63]) & (!i_12_) & (g95)) + ((i_14_) & (!sk[63]) & (i_12_) & (!g95)) + ((i_14_) & (!sk[63]) & (i_12_) & (g95)) + ((i_14_) & (sk[63]) & (!i_12_) & (g95)));
	assign g814 = (((!g297) & (!g270) & (!sk[64]) & (!g243) & (!g813) & (g495)) + ((!g297) & (!g270) & (!sk[64]) & (!g243) & (g813) & (g495)) + ((!g297) & (!g270) & (!sk[64]) & (g243) & (!g813) & (g495)) + ((!g297) & (!g270) & (!sk[64]) & (g243) & (g813) & (g495)) + ((!g297) & (!g270) & (sk[64]) & (!g243) & (!g813) & (!g495)) + ((!g297) & (!g270) & (sk[64]) & (!g243) & (!g813) & (g495)) + ((!g297) & (!g270) & (sk[64]) & (!g243) & (g813) & (!g495)) + ((!g297) & (g270) & (!sk[64]) & (!g243) & (!g813) & (g495)) + ((!g297) & (g270) & (!sk[64]) & (!g243) & (g813) & (g495)) + ((!g297) & (g270) & (!sk[64]) & (g243) & (!g813) & (g495)) + ((!g297) & (g270) & (!sk[64]) & (g243) & (g813) & (g495)) + ((!g297) & (g270) & (sk[64]) & (!g243) & (!g813) & (!g495)) + ((!g297) & (g270) & (sk[64]) & (!g243) & (!g813) & (g495)) + ((!g297) & (g270) & (sk[64]) & (!g243) & (g813) & (!g495)) + ((!g297) & (g270) & (sk[64]) & (g243) & (!g813) & (!g495)) + ((!g297) & (g270) & (sk[64]) & (g243) & (!g813) & (g495)) + ((!g297) & (g270) & (sk[64]) & (g243) & (g813) & (!g495)) + ((g297) & (!g270) & (!sk[64]) & (!g243) & (!g813) & (!g495)) + ((g297) & (!g270) & (!sk[64]) & (!g243) & (!g813) & (g495)) + ((g297) & (!g270) & (!sk[64]) & (!g243) & (g813) & (!g495)) + ((g297) & (!g270) & (!sk[64]) & (!g243) & (g813) & (g495)) + ((g297) & (!g270) & (!sk[64]) & (g243) & (!g813) & (!g495)) + ((g297) & (!g270) & (!sk[64]) & (g243) & (!g813) & (g495)) + ((g297) & (!g270) & (!sk[64]) & (g243) & (g813) & (!g495)) + ((g297) & (!g270) & (!sk[64]) & (g243) & (g813) & (g495)) + ((g297) & (!g270) & (sk[64]) & (!g243) & (!g813) & (!g495)) + ((g297) & (!g270) & (sk[64]) & (!g243) & (g813) & (!g495)) + ((g297) & (g270) & (!sk[64]) & (!g243) & (!g813) & (!g495)) + ((g297) & (g270) & (!sk[64]) & (!g243) & (!g813) & (g495)) + ((g297) & (g270) & (!sk[64]) & (!g243) & (g813) & (!g495)) + ((g297) & (g270) & (!sk[64]) & (!g243) & (g813) & (g495)) + ((g297) & (g270) & (!sk[64]) & (g243) & (!g813) & (!g495)) + ((g297) & (g270) & (!sk[64]) & (g243) & (!g813) & (g495)) + ((g297) & (g270) & (!sk[64]) & (g243) & (g813) & (!g495)) + ((g297) & (g270) & (!sk[64]) & (g243) & (g813) & (g495)) + ((g297) & (g270) & (sk[64]) & (!g243) & (!g813) & (!g495)) + ((g297) & (g270) & (sk[64]) & (!g243) & (g813) & (!g495)) + ((g297) & (g270) & (sk[64]) & (g243) & (!g813) & (!g495)) + ((g297) & (g270) & (sk[64]) & (g243) & (g813) & (!g495)));
	assign g815 = (((!g101) & (!g109) & (!g811) & (!g676) & (!g812) & (g814)) + ((!g101) & (!g109) & (!g811) & (g676) & (!g812) & (g814)) + ((!g101) & (!g109) & (g811) & (!g676) & (!g812) & (g814)) + ((!g101) & (!g109) & (g811) & (g676) & (!g812) & (g814)) + ((!g101) & (g109) & (!g811) & (!g676) & (!g812) & (g814)) + ((!g101) & (g109) & (!g811) & (g676) & (!g812) & (g814)) + ((g101) & (!g109) & (!g811) & (!g676) & (!g812) & (g814)) + ((g101) & (!g109) & (g811) & (!g676) & (!g812) & (g814)) + ((g101) & (g109) & (!g811) & (!g676) & (!g812) & (g814)));
	assign g816 = (((!g804) & (!g805) & (g1673) & (g810) & (g1666) & (g815)));
	assign g817 = (((!g6) & (!i_15_) & (!i_14_) & (!sk[67]) & (!i_12_) & (i_13_)) + ((!g6) & (!i_15_) & (!i_14_) & (!sk[67]) & (i_12_) & (i_13_)) + ((!g6) & (!i_15_) & (i_14_) & (!sk[67]) & (!i_12_) & (i_13_)) + ((!g6) & (!i_15_) & (i_14_) & (!sk[67]) & (i_12_) & (i_13_)) + ((!g6) & (i_15_) & (!i_14_) & (!sk[67]) & (!i_12_) & (i_13_)) + ((!g6) & (i_15_) & (!i_14_) & (!sk[67]) & (i_12_) & (i_13_)) + ((!g6) & (i_15_) & (i_14_) & (!sk[67]) & (!i_12_) & (i_13_)) + ((!g6) & (i_15_) & (i_14_) & (!sk[67]) & (i_12_) & (i_13_)) + ((g6) & (!i_15_) & (!i_14_) & (!sk[67]) & (!i_12_) & (!i_13_)) + ((g6) & (!i_15_) & (!i_14_) & (!sk[67]) & (!i_12_) & (i_13_)) + ((g6) & (!i_15_) & (!i_14_) & (!sk[67]) & (i_12_) & (!i_13_)) + ((g6) & (!i_15_) & (!i_14_) & (!sk[67]) & (i_12_) & (i_13_)) + ((g6) & (!i_15_) & (i_14_) & (!sk[67]) & (!i_12_) & (!i_13_)) + ((g6) & (!i_15_) & (i_14_) & (!sk[67]) & (!i_12_) & (i_13_)) + ((g6) & (!i_15_) & (i_14_) & (!sk[67]) & (i_12_) & (!i_13_)) + ((g6) & (!i_15_) & (i_14_) & (!sk[67]) & (i_12_) & (i_13_)) + ((g6) & (!i_15_) & (i_14_) & (sk[67]) & (!i_12_) & (!i_13_)) + ((g6) & (i_15_) & (!i_14_) & (!sk[67]) & (!i_12_) & (!i_13_)) + ((g6) & (i_15_) & (!i_14_) & (!sk[67]) & (!i_12_) & (i_13_)) + ((g6) & (i_15_) & (!i_14_) & (!sk[67]) & (i_12_) & (!i_13_)) + ((g6) & (i_15_) & (!i_14_) & (!sk[67]) & (i_12_) & (i_13_)) + ((g6) & (i_15_) & (!i_14_) & (sk[67]) & (i_12_) & (!i_13_)) + ((g6) & (i_15_) & (!i_14_) & (sk[67]) & (i_12_) & (i_13_)) + ((g6) & (i_15_) & (i_14_) & (!sk[67]) & (!i_12_) & (!i_13_)) + ((g6) & (i_15_) & (i_14_) & (!sk[67]) & (!i_12_) & (i_13_)) + ((g6) & (i_15_) & (i_14_) & (!sk[67]) & (i_12_) & (!i_13_)) + ((g6) & (i_15_) & (i_14_) & (!sk[67]) & (i_12_) & (i_13_)));
	assign g818 = (((!g304) & (!g94) & (sk[68]) & (g475)) + ((g304) & (!g94) & (!sk[68]) & (!g475)) + ((g304) & (!g94) & (!sk[68]) & (g475)) + ((g304) & (g94) & (!sk[68]) & (!g475)) + ((g304) & (g94) & (!sk[68]) & (g475)));
	assign g819 = (((!i_8_) & (!sk[69]) & (!g10) & (!g108) & (!g158) & (g572)) + ((!i_8_) & (!sk[69]) & (!g10) & (!g108) & (g158) & (g572)) + ((!i_8_) & (!sk[69]) & (!g10) & (g108) & (!g158) & (g572)) + ((!i_8_) & (!sk[69]) & (!g10) & (g108) & (g158) & (g572)) + ((!i_8_) & (!sk[69]) & (g10) & (!g108) & (!g158) & (g572)) + ((!i_8_) & (!sk[69]) & (g10) & (!g108) & (g158) & (g572)) + ((!i_8_) & (!sk[69]) & (g10) & (g108) & (!g158) & (g572)) + ((!i_8_) & (!sk[69]) & (g10) & (g108) & (g158) & (g572)) + ((!i_8_) & (sk[69]) & (!g10) & (g108) & (g158) & (g572)) + ((!i_8_) & (sk[69]) & (g10) & (g108) & (g158) & (g572)) + ((i_8_) & (!sk[69]) & (!g10) & (!g108) & (!g158) & (!g572)) + ((i_8_) & (!sk[69]) & (!g10) & (!g108) & (!g158) & (g572)) + ((i_8_) & (!sk[69]) & (!g10) & (!g108) & (g158) & (!g572)) + ((i_8_) & (!sk[69]) & (!g10) & (!g108) & (g158) & (g572)) + ((i_8_) & (!sk[69]) & (!g10) & (g108) & (!g158) & (!g572)) + ((i_8_) & (!sk[69]) & (!g10) & (g108) & (!g158) & (g572)) + ((i_8_) & (!sk[69]) & (!g10) & (g108) & (g158) & (!g572)) + ((i_8_) & (!sk[69]) & (!g10) & (g108) & (g158) & (g572)) + ((i_8_) & (!sk[69]) & (g10) & (!g108) & (!g158) & (!g572)) + ((i_8_) & (!sk[69]) & (g10) & (!g108) & (!g158) & (g572)) + ((i_8_) & (!sk[69]) & (g10) & (!g108) & (g158) & (!g572)) + ((i_8_) & (!sk[69]) & (g10) & (!g108) & (g158) & (g572)) + ((i_8_) & (!sk[69]) & (g10) & (g108) & (!g158) & (!g572)) + ((i_8_) & (!sk[69]) & (g10) & (g108) & (!g158) & (g572)) + ((i_8_) & (!sk[69]) & (g10) & (g108) & (g158) & (!g572)) + ((i_8_) & (!sk[69]) & (g10) & (g108) & (g158) & (g572)) + ((i_8_) & (sk[69]) & (g10) & (g108) & (!g158) & (!g572)) + ((i_8_) & (sk[69]) & (g10) & (g108) & (!g158) & (g572)) + ((i_8_) & (sk[69]) & (g10) & (g108) & (g158) & (!g572)) + ((i_8_) & (sk[69]) & (g10) & (g108) & (g158) & (g572)));
	assign g820 = (((!g216) & (!g423) & (!g817) & (!sk[70]) & (!g818) & (g819)) + ((!g216) & (!g423) & (!g817) & (!sk[70]) & (g818) & (g819)) + ((!g216) & (!g423) & (!g817) & (sk[70]) & (!g818) & (!g819)) + ((!g216) & (!g423) & (!g817) & (sk[70]) & (g818) & (!g819)) + ((!g216) & (!g423) & (g817) & (!sk[70]) & (!g818) & (g819)) + ((!g216) & (!g423) & (g817) & (!sk[70]) & (g818) & (g819)) + ((!g216) & (!g423) & (g817) & (sk[70]) & (!g818) & (!g819)) + ((!g216) & (!g423) & (g817) & (sk[70]) & (g818) & (!g819)) + ((!g216) & (g423) & (!g817) & (!sk[70]) & (!g818) & (g819)) + ((!g216) & (g423) & (!g817) & (!sk[70]) & (g818) & (g819)) + ((!g216) & (g423) & (!g817) & (sk[70]) & (g818) & (!g819)) + ((!g216) & (g423) & (g817) & (!sk[70]) & (!g818) & (g819)) + ((!g216) & (g423) & (g817) & (!sk[70]) & (g818) & (g819)) + ((g216) & (!g423) & (!g817) & (!sk[70]) & (!g818) & (!g819)) + ((g216) & (!g423) & (!g817) & (!sk[70]) & (!g818) & (g819)) + ((g216) & (!g423) & (!g817) & (!sk[70]) & (g818) & (!g819)) + ((g216) & (!g423) & (!g817) & (!sk[70]) & (g818) & (g819)) + ((g216) & (!g423) & (!g817) & (sk[70]) & (!g818) & (!g819)) + ((g216) & (!g423) & (!g817) & (sk[70]) & (g818) & (!g819)) + ((g216) & (!g423) & (g817) & (!sk[70]) & (!g818) & (!g819)) + ((g216) & (!g423) & (g817) & (!sk[70]) & (!g818) & (g819)) + ((g216) & (!g423) & (g817) & (!sk[70]) & (g818) & (!g819)) + ((g216) & (!g423) & (g817) & (!sk[70]) & (g818) & (g819)) + ((g216) & (!g423) & (g817) & (sk[70]) & (!g818) & (!g819)) + ((g216) & (!g423) & (g817) & (sk[70]) & (g818) & (!g819)) + ((g216) & (g423) & (!g817) & (!sk[70]) & (!g818) & (!g819)) + ((g216) & (g423) & (!g817) & (!sk[70]) & (!g818) & (g819)) + ((g216) & (g423) & (!g817) & (!sk[70]) & (g818) & (!g819)) + ((g216) & (g423) & (!g817) & (!sk[70]) & (g818) & (g819)) + ((g216) & (g423) & (g817) & (!sk[70]) & (!g818) & (!g819)) + ((g216) & (g423) & (g817) & (!sk[70]) & (!g818) & (g819)) + ((g216) & (g423) & (g817) & (!sk[70]) & (g818) & (!g819)) + ((g216) & (g423) & (g817) & (!sk[70]) & (g818) & (g819)));
	assign g821 = (((g301) & (g1768) & (g306) & (g313) & (g321) & (g820)));
	assign g822 = (((!i_14_) & (!i_12_) & (!sk[72]) & (g18) & (g119)) + ((!i_14_) & (i_12_) & (!sk[72]) & (!g18) & (!g119)) + ((!i_14_) & (i_12_) & (!sk[72]) & (!g18) & (g119)) + ((!i_14_) & (i_12_) & (!sk[72]) & (g18) & (!g119)) + ((!i_14_) & (i_12_) & (!sk[72]) & (g18) & (g119)) + ((!i_14_) & (i_12_) & (sk[72]) & (!g18) & (!g119)) + ((!i_14_) & (i_12_) & (sk[72]) & (!g18) & (g119)) + ((i_14_) & (!i_12_) & (!sk[72]) & (g18) & (!g119)) + ((i_14_) & (!i_12_) & (!sk[72]) & (g18) & (g119)) + ((i_14_) & (!i_12_) & (sk[72]) & (!g18) & (g119)) + ((i_14_) & (!i_12_) & (sk[72]) & (g18) & (g119)) + ((i_14_) & (i_12_) & (!sk[72]) & (!g18) & (!g119)) + ((i_14_) & (i_12_) & (!sk[72]) & (!g18) & (g119)) + ((i_14_) & (i_12_) & (!sk[72]) & (g18) & (!g119)) + ((i_14_) & (i_12_) & (!sk[72]) & (g18) & (g119)));
	assign g823 = (((!g270) & (!g204) & (!sk[73]) & (!g817) & (!g724) & (g822)) + ((!g270) & (!g204) & (!sk[73]) & (!g817) & (g724) & (g822)) + ((!g270) & (!g204) & (!sk[73]) & (g817) & (!g724) & (g822)) + ((!g270) & (!g204) & (!sk[73]) & (g817) & (g724) & (g822)) + ((!g270) & (g204) & (!sk[73]) & (!g817) & (!g724) & (g822)) + ((!g270) & (g204) & (!sk[73]) & (!g817) & (g724) & (g822)) + ((!g270) & (g204) & (!sk[73]) & (g817) & (!g724) & (g822)) + ((!g270) & (g204) & (!sk[73]) & (g817) & (g724) & (g822)) + ((g270) & (!g204) & (!sk[73]) & (!g817) & (!g724) & (!g822)) + ((g270) & (!g204) & (!sk[73]) & (!g817) & (!g724) & (g822)) + ((g270) & (!g204) & (!sk[73]) & (!g817) & (g724) & (!g822)) + ((g270) & (!g204) & (!sk[73]) & (!g817) & (g724) & (g822)) + ((g270) & (!g204) & (!sk[73]) & (g817) & (!g724) & (!g822)) + ((g270) & (!g204) & (!sk[73]) & (g817) & (!g724) & (g822)) + ((g270) & (!g204) & (!sk[73]) & (g817) & (g724) & (!g822)) + ((g270) & (!g204) & (!sk[73]) & (g817) & (g724) & (g822)) + ((g270) & (g204) & (!sk[73]) & (!g817) & (!g724) & (!g822)) + ((g270) & (g204) & (!sk[73]) & (!g817) & (!g724) & (g822)) + ((g270) & (g204) & (!sk[73]) & (!g817) & (g724) & (!g822)) + ((g270) & (g204) & (!sk[73]) & (!g817) & (g724) & (g822)) + ((g270) & (g204) & (!sk[73]) & (g817) & (!g724) & (!g822)) + ((g270) & (g204) & (!sk[73]) & (g817) & (!g724) & (g822)) + ((g270) & (g204) & (!sk[73]) & (g817) & (g724) & (!g822)) + ((g270) & (g204) & (!sk[73]) & (g817) & (g724) & (g822)) + ((g270) & (g204) & (sk[73]) & (!g817) & (!g724) & (!g822)));
	assign g824 = (((!g246) & (!g421) & (!g517) & (!g678) & (!sk[74]) & (g823)) + ((!g246) & (!g421) & (!g517) & (g678) & (!sk[74]) & (g823)) + ((!g246) & (!g421) & (g517) & (!g678) & (!sk[74]) & (g823)) + ((!g246) & (!g421) & (g517) & (g678) & (!sk[74]) & (g823)) + ((!g246) & (g421) & (!g517) & (!g678) & (!sk[74]) & (g823)) + ((!g246) & (g421) & (!g517) & (g678) & (!sk[74]) & (g823)) + ((!g246) & (g421) & (g517) & (!g678) & (!sk[74]) & (g823)) + ((!g246) & (g421) & (g517) & (g678) & (!sk[74]) & (g823)) + ((!g246) & (g421) & (g517) & (g678) & (sk[74]) & (g823)) + ((g246) & (!g421) & (!g517) & (!g678) & (!sk[74]) & (!g823)) + ((g246) & (!g421) & (!g517) & (!g678) & (!sk[74]) & (g823)) + ((g246) & (!g421) & (!g517) & (g678) & (!sk[74]) & (!g823)) + ((g246) & (!g421) & (!g517) & (g678) & (!sk[74]) & (g823)) + ((g246) & (!g421) & (g517) & (!g678) & (!sk[74]) & (!g823)) + ((g246) & (!g421) & (g517) & (!g678) & (!sk[74]) & (g823)) + ((g246) & (!g421) & (g517) & (g678) & (!sk[74]) & (!g823)) + ((g246) & (!g421) & (g517) & (g678) & (!sk[74]) & (g823)) + ((g246) & (g421) & (!g517) & (!g678) & (!sk[74]) & (!g823)) + ((g246) & (g421) & (!g517) & (!g678) & (!sk[74]) & (g823)) + ((g246) & (g421) & (!g517) & (g678) & (!sk[74]) & (!g823)) + ((g246) & (g421) & (!g517) & (g678) & (!sk[74]) & (g823)) + ((g246) & (g421) & (g517) & (!g678) & (!sk[74]) & (!g823)) + ((g246) & (g421) & (g517) & (!g678) & (!sk[74]) & (g823)) + ((g246) & (g421) & (g517) & (g678) & (!sk[74]) & (!g823)) + ((g246) & (g421) & (g517) & (g678) & (!sk[74]) & (g823)));
	assign g825 = (((g134) & (!sk[75]) & (!g824)) + ((g134) & (!sk[75]) & (g824)) + ((g134) & (sk[75]) & (!g824)));
	assign g826 = (((g464) & (!sk[76]) & (!g478) & (!g487)) + ((g464) & (!sk[76]) & (!g478) & (g487)) + ((g464) & (!sk[76]) & (g478) & (!g487)) + ((g464) & (!sk[76]) & (g478) & (g487)) + ((g464) & (sk[76]) & (!g478) & (!g487)));
	assign g827 = (((!g264) & (sk[77]) & (!g115) & (!g711)) + ((!g264) & (sk[77]) & (g115) & (!g711)) + ((!g264) & (sk[77]) & (g115) & (g711)) + ((g264) & (!sk[77]) & (!g115) & (!g711)) + ((g264) & (!sk[77]) & (!g115) & (g711)) + ((g264) & (!sk[77]) & (g115) & (!g711)) + ((g264) & (!sk[77]) & (g115) & (g711)));
	assign g828 = (((!i_8_) & (!g124) & (!sk[78]) & (g572) & (g672)) + ((!i_8_) & (g124) & (!sk[78]) & (!g572) & (!g672)) + ((!i_8_) & (g124) & (!sk[78]) & (!g572) & (g672)) + ((!i_8_) & (g124) & (!sk[78]) & (g572) & (!g672)) + ((!i_8_) & (g124) & (!sk[78]) & (g572) & (g672)) + ((!i_8_) & (g124) & (sk[78]) & (g572) & (!g672)) + ((!i_8_) & (g124) & (sk[78]) & (g572) & (g672)) + ((i_8_) & (!g124) & (!sk[78]) & (g572) & (!g672)) + ((i_8_) & (!g124) & (!sk[78]) & (g572) & (g672)) + ((i_8_) & (!g124) & (sk[78]) & (!g572) & (g672)) + ((i_8_) & (!g124) & (sk[78]) & (g572) & (g672)) + ((i_8_) & (g124) & (!sk[78]) & (!g572) & (!g672)) + ((i_8_) & (g124) & (!sk[78]) & (!g572) & (g672)) + ((i_8_) & (g124) & (!sk[78]) & (g572) & (!g672)) + ((i_8_) & (g124) & (!sk[78]) & (g572) & (g672)) + ((i_8_) & (g124) & (sk[78]) & (!g572) & (g672)) + ((i_8_) & (g124) & (sk[78]) & (g572) & (g672)));
	assign g829 = (((!g243) & (!g423) & (g827) & (!sk[79]) & (g828)) + ((!g243) & (g423) & (!g827) & (!sk[79]) & (!g828)) + ((!g243) & (g423) & (!g827) & (!sk[79]) & (g828)) + ((!g243) & (g423) & (!g827) & (sk[79]) & (!g828)) + ((!g243) & (g423) & (!g827) & (sk[79]) & (g828)) + ((!g243) & (g423) & (g827) & (!sk[79]) & (!g828)) + ((!g243) & (g423) & (g827) & (!sk[79]) & (g828)) + ((g243) & (!g423) & (!g827) & (sk[79]) & (g828)) + ((g243) & (!g423) & (g827) & (!sk[79]) & (!g828)) + ((g243) & (!g423) & (g827) & (!sk[79]) & (g828)) + ((g243) & (!g423) & (g827) & (sk[79]) & (g828)) + ((g243) & (g423) & (!g827) & (!sk[79]) & (!g828)) + ((g243) & (g423) & (!g827) & (!sk[79]) & (g828)) + ((g243) & (g423) & (!g827) & (sk[79]) & (!g828)) + ((g243) & (g423) & (!g827) & (sk[79]) & (g828)) + ((g243) & (g423) & (g827) & (!sk[79]) & (!g828)) + ((g243) & (g423) & (g827) & (!sk[79]) & (g828)) + ((g243) & (g423) & (g827) & (sk[79]) & (g828)));
	assign g830 = (((!g113) & (!g326) & (!g88) & (!g826) & (!sk[80]) & (g829)) + ((!g113) & (!g326) & (!g88) & (!g826) & (sk[80]) & (!g829)) + ((!g113) & (!g326) & (!g88) & (g826) & (!sk[80]) & (g829)) + ((!g113) & (!g326) & (!g88) & (g826) & (sk[80]) & (!g829)) + ((!g113) & (!g326) & (g88) & (!g826) & (!sk[80]) & (g829)) + ((!g113) & (!g326) & (g88) & (g826) & (!sk[80]) & (g829)) + ((!g113) & (!g326) & (g88) & (g826) & (sk[80]) & (!g829)) + ((!g113) & (g326) & (!g88) & (!g826) & (!sk[80]) & (g829)) + ((!g113) & (g326) & (!g88) & (!g826) & (sk[80]) & (!g829)) + ((!g113) & (g326) & (!g88) & (g826) & (!sk[80]) & (g829)) + ((!g113) & (g326) & (!g88) & (g826) & (sk[80]) & (!g829)) + ((!g113) & (g326) & (g88) & (!g826) & (!sk[80]) & (g829)) + ((!g113) & (g326) & (g88) & (g826) & (!sk[80]) & (g829)) + ((!g113) & (g326) & (g88) & (g826) & (sk[80]) & (!g829)) + ((g113) & (!g326) & (!g88) & (!g826) & (!sk[80]) & (!g829)) + ((g113) & (!g326) & (!g88) & (!g826) & (!sk[80]) & (g829)) + ((g113) & (!g326) & (!g88) & (!g826) & (sk[80]) & (!g829)) + ((g113) & (!g326) & (!g88) & (g826) & (!sk[80]) & (!g829)) + ((g113) & (!g326) & (!g88) & (g826) & (!sk[80]) & (g829)) + ((g113) & (!g326) & (!g88) & (g826) & (sk[80]) & (!g829)) + ((g113) & (!g326) & (g88) & (!g826) & (!sk[80]) & (!g829)) + ((g113) & (!g326) & (g88) & (!g826) & (!sk[80]) & (g829)) + ((g113) & (!g326) & (g88) & (g826) & (!sk[80]) & (!g829)) + ((g113) & (!g326) & (g88) & (g826) & (!sk[80]) & (g829)) + ((g113) & (!g326) & (g88) & (g826) & (sk[80]) & (!g829)) + ((g113) & (g326) & (!g88) & (!g826) & (!sk[80]) & (!g829)) + ((g113) & (g326) & (!g88) & (!g826) & (!sk[80]) & (g829)) + ((g113) & (g326) & (!g88) & (!g826) & (sk[80]) & (!g829)) + ((g113) & (g326) & (!g88) & (g826) & (!sk[80]) & (!g829)) + ((g113) & (g326) & (!g88) & (g826) & (!sk[80]) & (g829)) + ((g113) & (g326) & (!g88) & (g826) & (sk[80]) & (!g829)) + ((g113) & (g326) & (g88) & (!g826) & (!sk[80]) & (!g829)) + ((g113) & (g326) & (g88) & (!g826) & (!sk[80]) & (g829)) + ((g113) & (g326) & (g88) & (g826) & (!sk[80]) & (!g829)) + ((g113) & (g326) & (g88) & (g826) & (!sk[80]) & (g829)));
	assign g831 = (((!sk[81]) & (!g135) & (!g195) & (g412) & (g677)) + ((!sk[81]) & (!g135) & (g195) & (!g412) & (!g677)) + ((!sk[81]) & (!g135) & (g195) & (!g412) & (g677)) + ((!sk[81]) & (!g135) & (g195) & (g412) & (!g677)) + ((!sk[81]) & (!g135) & (g195) & (g412) & (g677)) + ((!sk[81]) & (g135) & (!g195) & (g412) & (!g677)) + ((!sk[81]) & (g135) & (!g195) & (g412) & (g677)) + ((!sk[81]) & (g135) & (g195) & (!g412) & (!g677)) + ((!sk[81]) & (g135) & (g195) & (!g412) & (g677)) + ((!sk[81]) & (g135) & (g195) & (g412) & (!g677)) + ((!sk[81]) & (g135) & (g195) & (g412) & (g677)) + ((sk[81]) & (g135) & (!g195) & (!g412) & (!g677)) + ((sk[81]) & (g135) & (!g195) & (!g412) & (g677)) + ((sk[81]) & (g135) & (!g195) & (g412) & (g677)) + ((sk[81]) & (g135) & (g195) & (!g412) & (!g677)) + ((sk[81]) & (g135) & (g195) & (!g412) & (g677)) + ((sk[81]) & (g135) & (g195) & (g412) & (!g677)) + ((sk[81]) & (g135) & (g195) & (g412) & (g677)));
	assign g832 = (((!g6) & (!g141) & (!g326) & (!g59) & (!g89) & (!g831)) + ((!g6) & (!g141) & (!g326) & (!g59) & (g89) & (!g831)) + ((!g6) & (!g141) & (!g326) & (g59) & (!g89) & (!g831)) + ((!g6) & (!g141) & (!g326) & (g59) & (g89) & (!g831)) + ((!g6) & (!g141) & (g326) & (!g59) & (!g89) & (!g831)) + ((!g6) & (!g141) & (g326) & (!g59) & (g89) & (!g831)) + ((!g6) & (!g141) & (g326) & (g59) & (!g89) & (!g831)) + ((!g6) & (!g141) & (g326) & (g59) & (g89) & (!g831)) + ((!g6) & (g141) & (!g326) & (!g59) & (!g89) & (!g831)) + ((!g6) & (g141) & (!g326) & (!g59) & (g89) & (!g831)) + ((!g6) & (g141) & (!g326) & (g59) & (!g89) & (!g831)) + ((!g6) & (g141) & (!g326) & (g59) & (g89) & (!g831)) + ((!g6) & (g141) & (g326) & (!g59) & (g89) & (!g831)) + ((!g6) & (g141) & (g326) & (g59) & (g89) & (!g831)) + ((g6) & (!g141) & (!g326) & (!g59) & (!g89) & (!g831)) + ((g6) & (!g141) & (!g326) & (!g59) & (g89) & (!g831)) + ((g6) & (!g141) & (!g326) & (g59) & (!g89) & (!g831)) + ((g6) & (!g141) & (!g326) & (g59) & (g89) & (!g831)) + ((g6) & (!g141) & (g326) & (!g59) & (g89) & (!g831)) + ((g6) & (g141) & (!g326) & (!g59) & (!g89) & (!g831)) + ((g6) & (g141) & (!g326) & (!g59) & (g89) & (!g831)) + ((g6) & (g141) & (!g326) & (g59) & (!g89) & (!g831)) + ((g6) & (g141) & (!g326) & (g59) & (g89) & (!g831)) + ((g6) & (g141) & (g326) & (!g59) & (g89) & (!g831)));
	assign g833 = (((!i_8_) & (!g10) & (!g16) & (g108) & (!g574) & (!g678)) + ((!i_8_) & (!g10) & (!g16) & (g108) & (!g574) & (g678)) + ((!i_8_) & (!g10) & (!g16) & (g108) & (g574) & (!g678)) + ((!i_8_) & (!g10) & (!g16) & (g108) & (g574) & (g678)) + ((!i_8_) & (!g10) & (g16) & (g108) & (g574) & (!g678)) + ((!i_8_) & (!g10) & (g16) & (g108) & (g574) & (g678)) + ((!i_8_) & (g10) & (!g16) & (g108) & (!g574) & (!g678)) + ((!i_8_) & (g10) & (!g16) & (g108) & (!g574) & (g678)) + ((!i_8_) & (g10) & (!g16) & (g108) & (g574) & (!g678)) + ((!i_8_) & (g10) & (!g16) & (g108) & (g574) & (g678)) + ((!i_8_) & (g10) & (g16) & (g108) & (!g574) & (!g678)) + ((!i_8_) & (g10) & (g16) & (g108) & (!g574) & (g678)) + ((!i_8_) & (g10) & (g16) & (g108) & (g574) & (!g678)) + ((!i_8_) & (g10) & (g16) & (g108) & (g574) & (g678)) + ((i_8_) & (!g10) & (!g16) & (g108) & (!g574) & (!g678)) + ((i_8_) & (!g10) & (!g16) & (g108) & (g574) & (!g678)) + ((i_8_) & (!g10) & (!g16) & (g108) & (g574) & (g678)) + ((i_8_) & (!g10) & (g16) & (g108) & (!g574) & (!g678)) + ((i_8_) & (!g10) & (g16) & (g108) & (g574) & (!g678)) + ((i_8_) & (!g10) & (g16) & (g108) & (g574) & (g678)) + ((i_8_) & (g10) & (!g16) & (g108) & (!g574) & (!g678)) + ((i_8_) & (g10) & (!g16) & (g108) & (g574) & (!g678)) + ((i_8_) & (g10) & (!g16) & (g108) & (g574) & (g678)) + ((i_8_) & (g10) & (g16) & (g108) & (!g574) & (!g678)) + ((i_8_) & (g10) & (g16) & (g108) & (g574) & (!g678)) + ((i_8_) & (g10) & (g16) & (g108) & (g574) & (g678)));
	assign g834 = (((!sk[84]) & (!g145) & (!g339) & (g465) & (g833)) + ((!sk[84]) & (!g145) & (g339) & (!g465) & (!g833)) + ((!sk[84]) & (!g145) & (g339) & (!g465) & (g833)) + ((!sk[84]) & (!g145) & (g339) & (g465) & (!g833)) + ((!sk[84]) & (!g145) & (g339) & (g465) & (g833)) + ((!sk[84]) & (g145) & (!g339) & (g465) & (!g833)) + ((!sk[84]) & (g145) & (!g339) & (g465) & (g833)) + ((!sk[84]) & (g145) & (g339) & (!g465) & (!g833)) + ((!sk[84]) & (g145) & (g339) & (!g465) & (g833)) + ((!sk[84]) & (g145) & (g339) & (g465) & (!g833)) + ((!sk[84]) & (g145) & (g339) & (g465) & (g833)) + ((sk[84]) & (!g145) & (!g339) & (!g465) & (!g833)) + ((sk[84]) & (!g145) & (!g339) & (g465) & (!g833)) + ((sk[84]) & (!g145) & (g339) & (!g465) & (!g833)) + ((sk[84]) & (!g145) & (g339) & (g465) & (!g833)) + ((sk[84]) & (g145) & (!g339) & (g465) & (!g833)));
	assign g835 = (((!g216) & (!g122) & (sk[85]) & (!g711)) + ((!g216) & (g122) & (sk[85]) & (!g711)) + ((!g216) & (g122) & (sk[85]) & (g711)) + ((g216) & (!g122) & (!sk[85]) & (!g711)) + ((g216) & (!g122) & (!sk[85]) & (g711)) + ((g216) & (g122) & (!sk[85]) & (!g711)) + ((g216) & (g122) & (!sk[85]) & (g711)));
	assign g836 = (((!i_14_) & (!i_12_) & (g100) & (!g108) & (!g131) & (g734)) + ((!i_14_) & (!i_12_) & (g100) & (!g108) & (g131) & (g734)) + ((!i_14_) & (!i_12_) & (g100) & (g108) & (!g131) & (g734)) + ((!i_14_) & (!i_12_) & (g100) & (g108) & (g131) & (g734)) + ((!i_14_) & (i_12_) & (g100) & (!g108) & (!g131) & (g734)) + ((!i_14_) & (i_12_) & (g100) & (!g108) & (g131) & (g734)) + ((!i_14_) & (i_12_) & (g100) & (g108) & (!g131) & (g734)) + ((!i_14_) & (i_12_) & (g100) & (g108) & (g131) & (g734)) + ((i_14_) & (!i_12_) & (g100) & (!g108) & (!g131) & (g734)) + ((i_14_) & (!i_12_) & (g100) & (!g108) & (g131) & (g734)) + ((i_14_) & (!i_12_) & (g100) & (g108) & (!g131) & (g734)) + ((i_14_) & (!i_12_) & (g100) & (g108) & (g131) & (g734)) + ((i_14_) & (i_12_) & (!g100) & (g108) & (g131) & (!g734)) + ((i_14_) & (i_12_) & (!g100) & (g108) & (g131) & (g734)) + ((i_14_) & (i_12_) & (g100) & (!g108) & (!g131) & (g734)) + ((i_14_) & (i_12_) & (g100) & (!g108) & (g131) & (g734)) + ((i_14_) & (i_12_) & (g100) & (g108) & (!g131) & (g734)) + ((i_14_) & (i_12_) & (g100) & (g108) & (g131) & (!g734)) + ((i_14_) & (i_12_) & (g100) & (g108) & (g131) & (g734)));
	assign g837 = (((!sk[87]) & (g297) & (!g124) & (!g711)) + ((!sk[87]) & (g297) & (!g124) & (g711)) + ((!sk[87]) & (g297) & (g124) & (!g711)) + ((!sk[87]) & (g297) & (g124) & (g711)) + ((sk[87]) & (!g297) & (!g124) & (!g711)) + ((sk[87]) & (!g297) & (!g124) & (g711)) + ((sk[87]) & (!g297) & (g124) & (!g711)));
	assign g838 = (((!sk[88]) & (g21) & (!g22) & (!g711)) + ((!sk[88]) & (g21) & (!g22) & (g711)) + ((!sk[88]) & (g21) & (g22) & (!g711)) + ((!sk[88]) & (g21) & (g22) & (g711)) + ((sk[88]) & (!g21) & (!g22) & (!g711)) + ((sk[88]) & (!g21) & (!g22) & (g711)) + ((sk[88]) & (!g21) & (g22) & (!g711)));
	assign g839 = (((!g99) & (!g323) & (!g423) & (!sk[89]) & (!g837) & (g838)) + ((!g99) & (!g323) & (!g423) & (!sk[89]) & (g837) & (g838)) + ((!g99) & (!g323) & (!g423) & (sk[89]) & (!g837) & (!g838)) + ((!g99) & (!g323) & (!g423) & (sk[89]) & (!g837) & (g838)) + ((!g99) & (!g323) & (!g423) & (sk[89]) & (g837) & (!g838)) + ((!g99) & (!g323) & (!g423) & (sk[89]) & (g837) & (g838)) + ((!g99) & (!g323) & (g423) & (!sk[89]) & (!g837) & (g838)) + ((!g99) & (!g323) & (g423) & (!sk[89]) & (g837) & (g838)) + ((!g99) & (!g323) & (g423) & (sk[89]) & (g837) & (g838)) + ((!g99) & (g323) & (!g423) & (!sk[89]) & (!g837) & (g838)) + ((!g99) & (g323) & (!g423) & (!sk[89]) & (g837) & (g838)) + ((!g99) & (g323) & (!g423) & (sk[89]) & (g837) & (g838)) + ((!g99) & (g323) & (g423) & (!sk[89]) & (!g837) & (g838)) + ((!g99) & (g323) & (g423) & (!sk[89]) & (g837) & (g838)) + ((!g99) & (g323) & (g423) & (sk[89]) & (g837) & (g838)) + ((g99) & (!g323) & (!g423) & (!sk[89]) & (!g837) & (!g838)) + ((g99) & (!g323) & (!g423) & (!sk[89]) & (!g837) & (g838)) + ((g99) & (!g323) & (!g423) & (!sk[89]) & (g837) & (!g838)) + ((g99) & (!g323) & (!g423) & (!sk[89]) & (g837) & (g838)) + ((g99) & (!g323) & (!g423) & (sk[89]) & (g837) & (g838)) + ((g99) & (!g323) & (g423) & (!sk[89]) & (!g837) & (!g838)) + ((g99) & (!g323) & (g423) & (!sk[89]) & (!g837) & (g838)) + ((g99) & (!g323) & (g423) & (!sk[89]) & (g837) & (!g838)) + ((g99) & (!g323) & (g423) & (!sk[89]) & (g837) & (g838)) + ((g99) & (!g323) & (g423) & (sk[89]) & (g837) & (g838)) + ((g99) & (g323) & (!g423) & (!sk[89]) & (!g837) & (!g838)) + ((g99) & (g323) & (!g423) & (!sk[89]) & (!g837) & (g838)) + ((g99) & (g323) & (!g423) & (!sk[89]) & (g837) & (!g838)) + ((g99) & (g323) & (!g423) & (!sk[89]) & (g837) & (g838)) + ((g99) & (g323) & (!g423) & (sk[89]) & (g837) & (g838)) + ((g99) & (g323) & (g423) & (!sk[89]) & (!g837) & (!g838)) + ((g99) & (g323) & (g423) & (!sk[89]) & (!g837) & (g838)) + ((g99) & (g323) & (g423) & (!sk[89]) & (g837) & (!g838)) + ((g99) & (g323) & (g423) & (!sk[89]) & (g837) & (g838)) + ((g99) & (g323) & (g423) & (sk[89]) & (g837) & (g838)));
	assign g840 = (((!sk[90]) & (!g21) & (!g118) & (!g835) & (!g836) & (g839)) + ((!sk[90]) & (!g21) & (!g118) & (!g835) & (g836) & (g839)) + ((!sk[90]) & (!g21) & (!g118) & (g835) & (!g836) & (g839)) + ((!sk[90]) & (!g21) & (!g118) & (g835) & (g836) & (g839)) + ((!sk[90]) & (!g21) & (g118) & (!g835) & (!g836) & (g839)) + ((!sk[90]) & (!g21) & (g118) & (!g835) & (g836) & (g839)) + ((!sk[90]) & (!g21) & (g118) & (g835) & (!g836) & (g839)) + ((!sk[90]) & (!g21) & (g118) & (g835) & (g836) & (g839)) + ((!sk[90]) & (g21) & (!g118) & (!g835) & (!g836) & (!g839)) + ((!sk[90]) & (g21) & (!g118) & (!g835) & (!g836) & (g839)) + ((!sk[90]) & (g21) & (!g118) & (!g835) & (g836) & (!g839)) + ((!sk[90]) & (g21) & (!g118) & (!g835) & (g836) & (g839)) + ((!sk[90]) & (g21) & (!g118) & (g835) & (!g836) & (!g839)) + ((!sk[90]) & (g21) & (!g118) & (g835) & (!g836) & (g839)) + ((!sk[90]) & (g21) & (!g118) & (g835) & (g836) & (!g839)) + ((!sk[90]) & (g21) & (!g118) & (g835) & (g836) & (g839)) + ((!sk[90]) & (g21) & (g118) & (!g835) & (!g836) & (!g839)) + ((!sk[90]) & (g21) & (g118) & (!g835) & (!g836) & (g839)) + ((!sk[90]) & (g21) & (g118) & (!g835) & (g836) & (!g839)) + ((!sk[90]) & (g21) & (g118) & (!g835) & (g836) & (g839)) + ((!sk[90]) & (g21) & (g118) & (g835) & (!g836) & (!g839)) + ((!sk[90]) & (g21) & (g118) & (g835) & (!g836) & (g839)) + ((!sk[90]) & (g21) & (g118) & (g835) & (g836) & (!g839)) + ((!sk[90]) & (g21) & (g118) & (g835) & (g836) & (g839)) + ((sk[90]) & (!g21) & (!g118) & (!g835) & (!g836) & (g839)) + ((sk[90]) & (!g21) & (!g118) & (g835) & (!g836) & (g839)) + ((sk[90]) & (!g21) & (g118) & (g835) & (!g836) & (g839)) + ((sk[90]) & (g21) & (!g118) & (!g835) & (!g836) & (g839)) + ((sk[90]) & (g21) & (!g118) & (g835) & (!g836) & (g839)));
	assign g841 = (((!g825) & (g1653) & (g830) & (g832) & (g834) & (g840)));
	assign g842 = (((g457) & (g773) & (g803) & (g816) & (g821) & (g841)));
	assign g843 = (((!g136) & (!g462) & (g817) & (!sk[93]) & (g818)) + ((!g136) & (g462) & (!g817) & (!sk[93]) & (!g818)) + ((!g136) & (g462) & (!g817) & (!sk[93]) & (g818)) + ((!g136) & (g462) & (g817) & (!sk[93]) & (!g818)) + ((!g136) & (g462) & (g817) & (!sk[93]) & (g818)) + ((g136) & (!g462) & (!g817) & (sk[93]) & (!g818)) + ((g136) & (!g462) & (!g817) & (sk[93]) & (g818)) + ((g136) & (!g462) & (g817) & (!sk[93]) & (!g818)) + ((g136) & (!g462) & (g817) & (!sk[93]) & (g818)) + ((g136) & (!g462) & (g817) & (sk[93]) & (!g818)) + ((g136) & (!g462) & (g817) & (sk[93]) & (g818)) + ((g136) & (g462) & (!g817) & (!sk[93]) & (!g818)) + ((g136) & (g462) & (!g817) & (!sk[93]) & (g818)) + ((g136) & (g462) & (!g817) & (sk[93]) & (!g818)) + ((g136) & (g462) & (g817) & (!sk[93]) & (!g818)) + ((g136) & (g462) & (g817) & (!sk[93]) & (g818)) + ((g136) & (g462) & (g817) & (sk[93]) & (!g818)) + ((g136) & (g462) & (g817) & (sk[93]) & (g818)));
	assign g844 = (((!i_8_) & (!g21) & (!g22) & (!g100) & (!g711) & (g837)) + ((!i_8_) & (!g21) & (!g22) & (!g100) & (g711) & (g837)) + ((!i_8_) & (!g21) & (!g22) & (g100) & (!g711) & (g837)) + ((!i_8_) & (!g21) & (!g22) & (g100) & (g711) & (g837)) + ((!i_8_) & (!g21) & (g22) & (!g100) & (!g711) & (g837)) + ((!i_8_) & (!g21) & (g22) & (g100) & (!g711) & (g837)) + ((!i_8_) & (g21) & (!g22) & (!g100) & (!g711) & (g837)) + ((!i_8_) & (g21) & (!g22) & (!g100) & (g711) & (g837)) + ((!i_8_) & (g21) & (!g22) & (g100) & (!g711) & (g837)) + ((!i_8_) & (g21) & (!g22) & (g100) & (g711) & (g837)) + ((!i_8_) & (g21) & (g22) & (!g100) & (!g711) & (g837)) + ((!i_8_) & (g21) & (g22) & (g100) & (!g711) & (g837)) + ((i_8_) & (!g21) & (!g22) & (!g100) & (!g711) & (g837)) + ((i_8_) & (!g21) & (!g22) & (!g100) & (g711) & (g837)) + ((i_8_) & (!g21) & (!g22) & (g100) & (!g711) & (g837)) + ((i_8_) & (!g21) & (!g22) & (g100) & (g711) & (g837)) + ((i_8_) & (!g21) & (g22) & (!g100) & (!g711) & (g837)) + ((i_8_) & (!g21) & (g22) & (g100) & (!g711) & (g837)) + ((i_8_) & (g21) & (!g22) & (!g100) & (!g711) & (g837)) + ((i_8_) & (g21) & (!g22) & (!g100) & (g711) & (g837)) + ((i_8_) & (g21) & (g22) & (!g100) & (!g711) & (g837)));
	assign g845 = (((!g101) & (!g136) & (!g216) & (!g123) & (!g485) & (!g844)) + ((!g101) & (!g136) & (!g216) & (!g123) & (!g485) & (g844)) + ((!g101) & (!g136) & (!g216) & (!g123) & (g485) & (!g844)) + ((!g101) & (!g136) & (!g216) & (!g123) & (g485) & (g844)) + ((!g101) & (!g136) & (!g216) & (g123) & (!g485) & (!g844)) + ((!g101) & (!g136) & (!g216) & (g123) & (!g485) & (g844)) + ((!g101) & (!g136) & (!g216) & (g123) & (g485) & (!g844)) + ((!g101) & (!g136) & (!g216) & (g123) & (g485) & (g844)) + ((!g101) & (!g136) & (g216) & (!g123) & (!g485) & (!g844)) + ((!g101) & (!g136) & (g216) & (!g123) & (!g485) & (g844)) + ((!g101) & (!g136) & (g216) & (!g123) & (g485) & (!g844)) + ((!g101) & (!g136) & (g216) & (!g123) & (g485) & (g844)) + ((!g101) & (!g136) & (g216) & (g123) & (!g485) & (!g844)) + ((!g101) & (!g136) & (g216) & (g123) & (!g485) & (g844)) + ((!g101) & (!g136) & (g216) & (g123) & (g485) & (!g844)) + ((!g101) & (!g136) & (g216) & (g123) & (g485) & (g844)) + ((!g101) & (g136) & (!g216) & (!g123) & (!g485) & (!g844)) + ((!g101) & (g136) & (!g216) & (!g123) & (!g485) & (g844)) + ((g101) & (!g136) & (!g216) & (!g123) & (!g485) & (g844)) + ((g101) & (!g136) & (!g216) & (!g123) & (g485) & (g844)) + ((g101) & (!g136) & (!g216) & (g123) & (!g485) & (g844)) + ((g101) & (!g136) & (!g216) & (g123) & (g485) & (g844)) + ((g101) & (!g136) & (g216) & (!g123) & (!g485) & (g844)) + ((g101) & (!g136) & (g216) & (!g123) & (g485) & (g844)) + ((g101) & (!g136) & (g216) & (g123) & (!g485) & (g844)) + ((g101) & (!g136) & (g216) & (g123) & (g485) & (g844)) + ((g101) & (g136) & (!g216) & (!g123) & (!g485) & (g844)));
	assign g846 = (((!g14) & (!g112) & (!g323) & (!g835) & (!g807) & (!g827)) + ((!g14) & (!g112) & (!g323) & (!g835) & (!g807) & (g827)) + ((!g14) & (!g112) & (!g323) & (!g835) & (g807) & (!g827)) + ((!g14) & (!g112) & (!g323) & (!g835) & (g807) & (g827)) + ((!g14) & (!g112) & (!g323) & (g835) & (!g807) & (!g827)) + ((!g14) & (!g112) & (!g323) & (g835) & (!g807) & (g827)) + ((!g14) & (!g112) & (!g323) & (g835) & (g807) & (!g827)) + ((!g14) & (!g112) & (!g323) & (g835) & (g807) & (g827)) + ((!g14) & (!g112) & (g323) & (g835) & (g807) & (g827)) + ((!g14) & (g112) & (!g323) & (!g835) & (g807) & (g827)) + ((!g14) & (g112) & (!g323) & (g835) & (g807) & (g827)) + ((!g14) & (g112) & (g323) & (g835) & (g807) & (g827)) + ((g14) & (!g112) & (!g323) & (!g835) & (!g807) & (!g827)) + ((g14) & (!g112) & (!g323) & (!g835) & (!g807) & (g827)) + ((g14) & (!g112) & (!g323) & (!g835) & (g807) & (!g827)) + ((g14) & (!g112) & (!g323) & (!g835) & (g807) & (g827)) + ((g14) & (!g112) & (!g323) & (g835) & (!g807) & (!g827)) + ((g14) & (!g112) & (!g323) & (g835) & (!g807) & (g827)) + ((g14) & (!g112) & (!g323) & (g835) & (g807) & (!g827)) + ((g14) & (!g112) & (!g323) & (g835) & (g807) & (g827)) + ((g14) & (!g112) & (g323) & (g835) & (g807) & (g827)));
	assign g847 = (((!g145) & (!g151) & (!sk[97]) & (g811) & (g846)) + ((!g145) & (!g151) & (sk[97]) & (!g811) & (g846)) + ((!g145) & (!g151) & (sk[97]) & (g811) & (g846)) + ((!g145) & (g151) & (!sk[97]) & (!g811) & (!g846)) + ((!g145) & (g151) & (!sk[97]) & (!g811) & (g846)) + ((!g145) & (g151) & (!sk[97]) & (g811) & (!g846)) + ((!g145) & (g151) & (!sk[97]) & (g811) & (g846)) + ((!g145) & (g151) & (sk[97]) & (!g811) & (g846)) + ((g145) & (!g151) & (!sk[97]) & (g811) & (!g846)) + ((g145) & (!g151) & (!sk[97]) & (g811) & (g846)) + ((g145) & (!g151) & (sk[97]) & (!g811) & (g846)) + ((g145) & (g151) & (!sk[97]) & (!g811) & (!g846)) + ((g145) & (g151) & (!sk[97]) & (!g811) & (g846)) + ((g145) & (g151) & (!sk[97]) & (g811) & (!g846)) + ((g145) & (g151) & (!sk[97]) & (g811) & (g846)) + ((g145) & (g151) & (sk[97]) & (!g811) & (g846)));
	assign g848 = (((!g316) & (!g158) & (sk[98]) & (!g711)) + ((!g316) & (!g158) & (sk[98]) & (g711)) + ((!g316) & (g158) & (sk[98]) & (!g711)) + ((g316) & (!g158) & (!sk[98]) & (!g711)) + ((g316) & (!g158) & (!sk[98]) & (g711)) + ((g316) & (g158) & (!sk[98]) & (!g711)) + ((g316) & (g158) & (!sk[98]) & (g711)));
	assign g849 = (((!i_8_) & (!g88) & (g813) & (!sk[99]) & (g475)) + ((!i_8_) & (g88) & (!g813) & (!sk[99]) & (!g475)) + ((!i_8_) & (g88) & (!g813) & (!sk[99]) & (g475)) + ((!i_8_) & (g88) & (g813) & (!sk[99]) & (!g475)) + ((!i_8_) & (g88) & (g813) & (!sk[99]) & (g475)) + ((i_8_) & (!g88) & (g813) & (!sk[99]) & (!g475)) + ((i_8_) & (!g88) & (g813) & (!sk[99]) & (g475)) + ((i_8_) & (g88) & (!g813) & (!sk[99]) & (!g475)) + ((i_8_) & (g88) & (!g813) & (!sk[99]) & (g475)) + ((i_8_) & (g88) & (!g813) & (sk[99]) & (!g475)) + ((i_8_) & (g88) & (g813) & (!sk[99]) & (!g475)) + ((i_8_) & (g88) & (g813) & (!sk[99]) & (g475)) + ((i_8_) & (g88) & (g813) & (sk[99]) & (!g475)) + ((i_8_) & (g88) & (g813) & (sk[99]) & (g475)));
	assign g850 = (((!sk[100]) & (g323) & (!g817) & (!g818)) + ((!sk[100]) & (g323) & (!g817) & (g818)) + ((!sk[100]) & (g323) & (g817) & (!g818)) + ((!sk[100]) & (g323) & (g817) & (g818)) + ((sk[100]) & (g323) & (!g817) & (!g818)) + ((sk[100]) & (g323) & (g817) & (!g818)) + ((sk[100]) & (g323) & (g817) & (g818)));
	assign g851 = (((!g101) & (!sk[101]) & (!g145) & (!g848) & (!g849) & (g850)) + ((!g101) & (!sk[101]) & (!g145) & (!g848) & (g849) & (g850)) + ((!g101) & (!sk[101]) & (!g145) & (g848) & (!g849) & (g850)) + ((!g101) & (!sk[101]) & (!g145) & (g848) & (g849) & (g850)) + ((!g101) & (!sk[101]) & (g145) & (!g848) & (!g849) & (g850)) + ((!g101) & (!sk[101]) & (g145) & (!g848) & (g849) & (g850)) + ((!g101) & (!sk[101]) & (g145) & (g848) & (!g849) & (g850)) + ((!g101) & (!sk[101]) & (g145) & (g848) & (g849) & (g850)) + ((!g101) & (sk[101]) & (!g145) & (!g848) & (!g849) & (!g850)) + ((!g101) & (sk[101]) & (!g145) & (g848) & (!g849) & (!g850)) + ((!g101) & (sk[101]) & (g145) & (g848) & (!g849) & (!g850)) + ((g101) & (!sk[101]) & (!g145) & (!g848) & (!g849) & (!g850)) + ((g101) & (!sk[101]) & (!g145) & (!g848) & (!g849) & (g850)) + ((g101) & (!sk[101]) & (!g145) & (!g848) & (g849) & (!g850)) + ((g101) & (!sk[101]) & (!g145) & (!g848) & (g849) & (g850)) + ((g101) & (!sk[101]) & (!g145) & (g848) & (!g849) & (!g850)) + ((g101) & (!sk[101]) & (!g145) & (g848) & (!g849) & (g850)) + ((g101) & (!sk[101]) & (!g145) & (g848) & (g849) & (!g850)) + ((g101) & (!sk[101]) & (!g145) & (g848) & (g849) & (g850)) + ((g101) & (!sk[101]) & (g145) & (!g848) & (!g849) & (!g850)) + ((g101) & (!sk[101]) & (g145) & (!g848) & (!g849) & (g850)) + ((g101) & (!sk[101]) & (g145) & (!g848) & (g849) & (!g850)) + ((g101) & (!sk[101]) & (g145) & (!g848) & (g849) & (g850)) + ((g101) & (!sk[101]) & (g145) & (g848) & (!g849) & (!g850)) + ((g101) & (!sk[101]) & (g145) & (g848) & (!g849) & (g850)) + ((g101) & (!sk[101]) & (g145) & (g848) & (g849) & (!g850)) + ((g101) & (!sk[101]) & (g145) & (g848) & (g849) & (g850)) + ((g101) & (sk[101]) & (!g145) & (g848) & (!g849) & (!g850)) + ((g101) & (sk[101]) & (g145) & (g848) & (!g849) & (!g850)));
	assign g852 = (((!g843) & (!g845) & (!sk[102]) & (g847) & (g851)) + ((!g843) & (g845) & (!sk[102]) & (!g847) & (!g851)) + ((!g843) & (g845) & (!sk[102]) & (!g847) & (g851)) + ((!g843) & (g845) & (!sk[102]) & (g847) & (!g851)) + ((!g843) & (g845) & (!sk[102]) & (g847) & (g851)) + ((!g843) & (g845) & (sk[102]) & (g847) & (g851)) + ((g843) & (!g845) & (!sk[102]) & (g847) & (!g851)) + ((g843) & (!g845) & (!sk[102]) & (g847) & (g851)) + ((g843) & (g845) & (!sk[102]) & (!g847) & (!g851)) + ((g843) & (g845) & (!sk[102]) & (!g847) & (g851)) + ((g843) & (g845) & (!sk[102]) & (g847) & (!g851)) + ((g843) & (g845) & (!sk[102]) & (g847) & (g851)));
	assign g853 = (((g235) & (g274) & (g358) & (g374) & (g398) & (g852)));
	assign g854 = (((!g73) & (!g666) & (!g667) & (!g759) & (!g842) & (!g853)) + ((!g73) & (!g666) & (!g667) & (!g759) & (!g842) & (g853)) + ((!g73) & (!g666) & (!g667) & (!g759) & (g842) & (!g853)) + ((!g73) & (!g666) & (!g667) & (!g759) & (g842) & (g853)) + ((!g73) & (!g666) & (!g667) & (g759) & (!g842) & (!g853)) + ((!g73) & (!g666) & (!g667) & (g759) & (!g842) & (g853)) + ((!g73) & (!g666) & (!g667) & (g759) & (g842) & (!g853)) + ((!g73) & (!g666) & (!g667) & (g759) & (g842) & (g853)) + ((!g73) & (!g666) & (g667) & (!g759) & (!g842) & (!g853)) + ((!g73) & (!g666) & (g667) & (!g759) & (!g842) & (g853)) + ((!g73) & (!g666) & (g667) & (!g759) & (g842) & (!g853)) + ((!g73) & (!g666) & (g667) & (!g759) & (g842) & (g853)) + ((!g73) & (!g666) & (g667) & (g759) & (!g842) & (!g853)) + ((!g73) & (!g666) & (g667) & (g759) & (!g842) & (g853)) + ((!g73) & (!g666) & (g667) & (g759) & (g842) & (!g853)) + ((!g73) & (!g666) & (g667) & (g759) & (g842) & (g853)) + ((!g73) & (g666) & (!g667) & (!g759) & (!g842) & (!g853)) + ((!g73) & (g666) & (!g667) & (!g759) & (!g842) & (g853)) + ((!g73) & (g666) & (!g667) & (!g759) & (g842) & (!g853)) + ((!g73) & (g666) & (!g667) & (!g759) & (g842) & (g853)) + ((!g73) & (g666) & (!g667) & (g759) & (!g842) & (!g853)) + ((!g73) & (g666) & (!g667) & (g759) & (!g842) & (g853)) + ((!g73) & (g666) & (!g667) & (g759) & (g842) & (!g853)) + ((!g73) & (g666) & (!g667) & (g759) & (g842) & (g853)) + ((!g73) & (g666) & (g667) & (!g759) & (!g842) & (!g853)) + ((!g73) & (g666) & (g667) & (!g759) & (!g842) & (g853)) + ((!g73) & (g666) & (g667) & (!g759) & (g842) & (!g853)) + ((!g73) & (g666) & (g667) & (!g759) & (g842) & (g853)) + ((!g73) & (g666) & (g667) & (g759) & (!g842) & (!g853)) + ((!g73) & (g666) & (g667) & (g759) & (!g842) & (g853)) + ((!g73) & (g666) & (g667) & (g759) & (g842) & (!g853)) + ((!g73) & (g666) & (g667) & (g759) & (g842) & (g853)) + ((g73) & (g666) & (g667) & (g759) & (g842) & (g853)));
	assign g855 = (((!sk[105]) & (!i_5_) & (!i_3_) & (i_4_) & (g29)) + ((!sk[105]) & (!i_5_) & (i_3_) & (!i_4_) & (!g29)) + ((!sk[105]) & (!i_5_) & (i_3_) & (!i_4_) & (g29)) + ((!sk[105]) & (!i_5_) & (i_3_) & (i_4_) & (!g29)) + ((!sk[105]) & (!i_5_) & (i_3_) & (i_4_) & (g29)) + ((!sk[105]) & (i_5_) & (!i_3_) & (i_4_) & (!g29)) + ((!sk[105]) & (i_5_) & (!i_3_) & (i_4_) & (g29)) + ((!sk[105]) & (i_5_) & (i_3_) & (!i_4_) & (!g29)) + ((!sk[105]) & (i_5_) & (i_3_) & (!i_4_) & (g29)) + ((!sk[105]) & (i_5_) & (i_3_) & (i_4_) & (!g29)) + ((!sk[105]) & (i_5_) & (i_3_) & (i_4_) & (g29)) + ((sk[105]) & (!i_5_) & (!i_3_) & (!i_4_) & (g29)));
	assign o_7_ = (((!g2) & (!g36) & (!sk[106]) & (!g73) & (!g111) & (g855)) + ((!g2) & (!g36) & (!sk[106]) & (!g73) & (g111) & (g855)) + ((!g2) & (!g36) & (!sk[106]) & (g73) & (!g111) & (g855)) + ((!g2) & (!g36) & (!sk[106]) & (g73) & (g111) & (g855)) + ((!g2) & (!g36) & (sk[106]) & (g73) & (!g111) & (!g855)) + ((!g2) & (!g36) & (sk[106]) & (g73) & (!g111) & (g855)) + ((!g2) & (!g36) & (sk[106]) & (g73) & (g111) & (!g855)) + ((!g2) & (!g36) & (sk[106]) & (g73) & (g111) & (g855)) + ((!g2) & (g36) & (!sk[106]) & (!g73) & (!g111) & (g855)) + ((!g2) & (g36) & (!sk[106]) & (!g73) & (g111) & (g855)) + ((!g2) & (g36) & (!sk[106]) & (g73) & (!g111) & (g855)) + ((!g2) & (g36) & (!sk[106]) & (g73) & (g111) & (g855)) + ((!g2) & (g36) & (sk[106]) & (g73) & (!g111) & (g855)) + ((!g2) & (g36) & (sk[106]) & (g73) & (g111) & (g855)) + ((g2) & (!g36) & (!sk[106]) & (!g73) & (!g111) & (!g855)) + ((g2) & (!g36) & (!sk[106]) & (!g73) & (!g111) & (g855)) + ((g2) & (!g36) & (!sk[106]) & (!g73) & (g111) & (!g855)) + ((g2) & (!g36) & (!sk[106]) & (!g73) & (g111) & (g855)) + ((g2) & (!g36) & (!sk[106]) & (g73) & (!g111) & (!g855)) + ((g2) & (!g36) & (!sk[106]) & (g73) & (!g111) & (g855)) + ((g2) & (!g36) & (!sk[106]) & (g73) & (g111) & (!g855)) + ((g2) & (!g36) & (!sk[106]) & (g73) & (g111) & (g855)) + ((g2) & (!g36) & (sk[106]) & (g73) & (!g111) & (!g855)) + ((g2) & (!g36) & (sk[106]) & (g73) & (!g111) & (g855)) + ((g2) & (!g36) & (sk[106]) & (g73) & (g111) & (!g855)) + ((g2) & (!g36) & (sk[106]) & (g73) & (g111) & (g855)) + ((g2) & (g36) & (!sk[106]) & (!g73) & (!g111) & (!g855)) + ((g2) & (g36) & (!sk[106]) & (!g73) & (!g111) & (g855)) + ((g2) & (g36) & (!sk[106]) & (!g73) & (g111) & (!g855)) + ((g2) & (g36) & (!sk[106]) & (!g73) & (g111) & (g855)) + ((g2) & (g36) & (!sk[106]) & (g73) & (!g111) & (!g855)) + ((g2) & (g36) & (!sk[106]) & (g73) & (!g111) & (g855)) + ((g2) & (g36) & (!sk[106]) & (g73) & (g111) & (!g855)) + ((g2) & (g36) & (!sk[106]) & (g73) & (g111) & (g855)) + ((g2) & (g36) & (sk[106]) & (g73) & (!g111) & (g855)) + ((g2) & (g36) & (sk[106]) & (g73) & (g111) & (!g855)) + ((g2) & (g36) & (sk[106]) & (g73) & (g111) & (g855)));
	assign g857 = (((!g10) & (!g16) & (!g134) & (!g109) & (!g678) & (!g801)) + ((!g10) & (!g16) & (!g134) & (!g109) & (!g678) & (g801)) + ((!g10) & (!g16) & (!g134) & (!g109) & (g678) & (!g801)) + ((!g10) & (!g16) & (!g134) & (!g109) & (g678) & (g801)) + ((!g10) & (!g16) & (g134) & (!g109) & (g678) & (g801)) + ((!g10) & (g16) & (!g134) & (!g109) & (!g678) & (!g801)) + ((!g10) & (g16) & (!g134) & (!g109) & (!g678) & (g801)) + ((!g10) & (g16) & (!g134) & (!g109) & (g678) & (!g801)) + ((!g10) & (g16) & (!g134) & (!g109) & (g678) & (g801)) + ((!g10) & (g16) & (!g134) & (g109) & (!g678) & (!g801)) + ((!g10) & (g16) & (!g134) & (g109) & (!g678) & (g801)) + ((!g10) & (g16) & (!g134) & (g109) & (g678) & (!g801)) + ((!g10) & (g16) & (!g134) & (g109) & (g678) & (g801)) + ((!g10) & (g16) & (g134) & (!g109) & (g678) & (g801)) + ((!g10) & (g16) & (g134) & (g109) & (g678) & (g801)) + ((g10) & (!g16) & (!g134) & (!g109) & (!g678) & (!g801)) + ((g10) & (!g16) & (!g134) & (!g109) & (!g678) & (g801)) + ((g10) & (!g16) & (!g134) & (!g109) & (g678) & (!g801)) + ((g10) & (!g16) & (!g134) & (!g109) & (g678) & (g801)) + ((g10) & (!g16) & (g134) & (!g109) & (g678) & (g801)) + ((g10) & (g16) & (!g134) & (!g109) & (!g678) & (!g801)) + ((g10) & (g16) & (!g134) & (!g109) & (!g678) & (g801)) + ((g10) & (g16) & (!g134) & (!g109) & (g678) & (!g801)) + ((g10) & (g16) & (!g134) & (!g109) & (g678) & (g801)) + ((g10) & (g16) & (g134) & (!g109) & (g678) & (g801)));
	assign g858 = (((!g251) & (!g672) & (!sk[108]) & (g803) & (g857)) + ((!g251) & (!g672) & (sk[108]) & (g803) & (g857)) + ((!g251) & (g672) & (!sk[108]) & (!g803) & (!g857)) + ((!g251) & (g672) & (!sk[108]) & (!g803) & (g857)) + ((!g251) & (g672) & (!sk[108]) & (g803) & (!g857)) + ((!g251) & (g672) & (!sk[108]) & (g803) & (g857)) + ((!g251) & (g672) & (sk[108]) & (g803) & (g857)) + ((g251) & (!g672) & (!sk[108]) & (g803) & (!g857)) + ((g251) & (!g672) & (!sk[108]) & (g803) & (g857)) + ((g251) & (!g672) & (sk[108]) & (g803) & (g857)) + ((g251) & (g672) & (!sk[108]) & (!g803) & (!g857)) + ((g251) & (g672) & (!sk[108]) & (!g803) & (g857)) + ((g251) & (g672) & (!sk[108]) & (g803) & (!g857)) + ((g251) & (g672) & (!sk[108]) & (g803) & (g857)));
	assign g859 = (((!sk[109]) & (!g145) & (!g151) & (g142) & (g103)) + ((!sk[109]) & (!g145) & (g151) & (!g142) & (!g103)) + ((!sk[109]) & (!g145) & (g151) & (!g142) & (g103)) + ((!sk[109]) & (!g145) & (g151) & (g142) & (!g103)) + ((!sk[109]) & (!g145) & (g151) & (g142) & (g103)) + ((!sk[109]) & (g145) & (!g151) & (g142) & (!g103)) + ((!sk[109]) & (g145) & (!g151) & (g142) & (g103)) + ((!sk[109]) & (g145) & (g151) & (!g142) & (!g103)) + ((!sk[109]) & (g145) & (g151) & (!g142) & (g103)) + ((!sk[109]) & (g145) & (g151) & (g142) & (!g103)) + ((!sk[109]) & (g145) & (g151) & (g142) & (g103)) + ((sk[109]) & (!g145) & (!g151) & (!g142) & (!g103)) + ((sk[109]) & (!g145) & (!g151) & (!g142) & (g103)) + ((sk[109]) & (!g145) & (!g151) & (g142) & (!g103)) + ((sk[109]) & (!g145) & (!g151) & (g142) & (g103)) + ((sk[109]) & (!g145) & (g151) & (!g142) & (g103)) + ((sk[109]) & (g145) & (!g151) & (!g142) & (g103)) + ((sk[109]) & (g145) & (!g151) & (g142) & (g103)) + ((sk[109]) & (g145) & (g151) & (!g142) & (g103)));
	assign g860 = (((!g764) & (!sk[110]) & (!g765) & (!g766) & (!g772) & (g859)) + ((!g764) & (!sk[110]) & (!g765) & (!g766) & (g772) & (g859)) + ((!g764) & (!sk[110]) & (!g765) & (g766) & (!g772) & (g859)) + ((!g764) & (!sk[110]) & (!g765) & (g766) & (g772) & (g859)) + ((!g764) & (!sk[110]) & (g765) & (!g766) & (!g772) & (g859)) + ((!g764) & (!sk[110]) & (g765) & (!g766) & (g772) & (g859)) + ((!g764) & (!sk[110]) & (g765) & (g766) & (!g772) & (g859)) + ((!g764) & (!sk[110]) & (g765) & (g766) & (g772) & (g859)) + ((g764) & (!sk[110]) & (!g765) & (!g766) & (!g772) & (!g859)) + ((g764) & (!sk[110]) & (!g765) & (!g766) & (!g772) & (g859)) + ((g764) & (!sk[110]) & (!g765) & (!g766) & (g772) & (!g859)) + ((g764) & (!sk[110]) & (!g765) & (!g766) & (g772) & (g859)) + ((g764) & (!sk[110]) & (!g765) & (g766) & (!g772) & (!g859)) + ((g764) & (!sk[110]) & (!g765) & (g766) & (!g772) & (g859)) + ((g764) & (!sk[110]) & (!g765) & (g766) & (g772) & (!g859)) + ((g764) & (!sk[110]) & (!g765) & (g766) & (g772) & (g859)) + ((g764) & (!sk[110]) & (g765) & (!g766) & (!g772) & (!g859)) + ((g764) & (!sk[110]) & (g765) & (!g766) & (!g772) & (g859)) + ((g764) & (!sk[110]) & (g765) & (!g766) & (g772) & (!g859)) + ((g764) & (!sk[110]) & (g765) & (!g766) & (g772) & (g859)) + ((g764) & (!sk[110]) & (g765) & (g766) & (!g772) & (!g859)) + ((g764) & (!sk[110]) & (g765) & (g766) & (!g772) & (g859)) + ((g764) & (!sk[110]) & (g765) & (g766) & (g772) & (!g859)) + ((g764) & (!sk[110]) & (g765) & (g766) & (g772) & (g859)) + ((g764) & (sk[110]) & (g765) & (g766) & (g772) & (g859)));
	assign g861 = (((!i_8_) & (!g88) & (!sk[111]) & (!g108) & (!g678) & (g672)) + ((!i_8_) & (!g88) & (!sk[111]) & (!g108) & (g678) & (g672)) + ((!i_8_) & (!g88) & (!sk[111]) & (g108) & (!g678) & (g672)) + ((!i_8_) & (!g88) & (!sk[111]) & (g108) & (g678) & (g672)) + ((!i_8_) & (g88) & (!sk[111]) & (!g108) & (!g678) & (g672)) + ((!i_8_) & (g88) & (!sk[111]) & (!g108) & (g678) & (g672)) + ((!i_8_) & (g88) & (!sk[111]) & (g108) & (!g678) & (g672)) + ((!i_8_) & (g88) & (!sk[111]) & (g108) & (g678) & (g672)) + ((i_8_) & (!g88) & (!sk[111]) & (!g108) & (!g678) & (!g672)) + ((i_8_) & (!g88) & (!sk[111]) & (!g108) & (!g678) & (g672)) + ((i_8_) & (!g88) & (!sk[111]) & (!g108) & (g678) & (!g672)) + ((i_8_) & (!g88) & (!sk[111]) & (!g108) & (g678) & (g672)) + ((i_8_) & (!g88) & (!sk[111]) & (g108) & (!g678) & (!g672)) + ((i_8_) & (!g88) & (!sk[111]) & (g108) & (!g678) & (g672)) + ((i_8_) & (!g88) & (!sk[111]) & (g108) & (g678) & (!g672)) + ((i_8_) & (!g88) & (!sk[111]) & (g108) & (g678) & (g672)) + ((i_8_) & (!g88) & (sk[111]) & (g108) & (!g678) & (!g672)) + ((i_8_) & (!g88) & (sk[111]) & (g108) & (!g678) & (g672)) + ((i_8_) & (g88) & (!sk[111]) & (!g108) & (!g678) & (!g672)) + ((i_8_) & (g88) & (!sk[111]) & (!g108) & (!g678) & (g672)) + ((i_8_) & (g88) & (!sk[111]) & (!g108) & (g678) & (!g672)) + ((i_8_) & (g88) & (!sk[111]) & (!g108) & (g678) & (g672)) + ((i_8_) & (g88) & (!sk[111]) & (g108) & (!g678) & (!g672)) + ((i_8_) & (g88) & (!sk[111]) & (g108) & (!g678) & (g672)) + ((i_8_) & (g88) & (!sk[111]) & (g108) & (g678) & (!g672)) + ((i_8_) & (g88) & (!sk[111]) & (g108) & (g678) & (g672)) + ((i_8_) & (g88) & (sk[111]) & (!g108) & (!g678) & (g672)) + ((i_8_) & (g88) & (sk[111]) & (!g108) & (g678) & (g672)) + ((i_8_) & (g88) & (sk[111]) & (g108) & (!g678) & (!g672)) + ((i_8_) & (g88) & (sk[111]) & (g108) & (!g678) & (g672)) + ((i_8_) & (g88) & (sk[111]) & (g108) & (g678) & (g672)));
	assign g862 = (((!sk[112]) & (!g136) & (!g186) & (!g677) & (!g826) & (g861)) + ((!sk[112]) & (!g136) & (!g186) & (!g677) & (g826) & (g861)) + ((!sk[112]) & (!g136) & (!g186) & (g677) & (!g826) & (g861)) + ((!sk[112]) & (!g136) & (!g186) & (g677) & (g826) & (g861)) + ((!sk[112]) & (!g136) & (g186) & (!g677) & (!g826) & (g861)) + ((!sk[112]) & (!g136) & (g186) & (!g677) & (g826) & (g861)) + ((!sk[112]) & (!g136) & (g186) & (g677) & (!g826) & (g861)) + ((!sk[112]) & (!g136) & (g186) & (g677) & (g826) & (g861)) + ((!sk[112]) & (g136) & (!g186) & (!g677) & (!g826) & (!g861)) + ((!sk[112]) & (g136) & (!g186) & (!g677) & (!g826) & (g861)) + ((!sk[112]) & (g136) & (!g186) & (!g677) & (g826) & (!g861)) + ((!sk[112]) & (g136) & (!g186) & (!g677) & (g826) & (g861)) + ((!sk[112]) & (g136) & (!g186) & (g677) & (!g826) & (!g861)) + ((!sk[112]) & (g136) & (!g186) & (g677) & (!g826) & (g861)) + ((!sk[112]) & (g136) & (!g186) & (g677) & (g826) & (!g861)) + ((!sk[112]) & (g136) & (!g186) & (g677) & (g826) & (g861)) + ((!sk[112]) & (g136) & (g186) & (!g677) & (!g826) & (!g861)) + ((!sk[112]) & (g136) & (g186) & (!g677) & (!g826) & (g861)) + ((!sk[112]) & (g136) & (g186) & (!g677) & (g826) & (!g861)) + ((!sk[112]) & (g136) & (g186) & (!g677) & (g826) & (g861)) + ((!sk[112]) & (g136) & (g186) & (g677) & (!g826) & (!g861)) + ((!sk[112]) & (g136) & (g186) & (g677) & (!g826) & (g861)) + ((!sk[112]) & (g136) & (g186) & (g677) & (g826) & (!g861)) + ((!sk[112]) & (g136) & (g186) & (g677) & (g826) & (g861)) + ((sk[112]) & (!g136) & (!g186) & (!g677) & (!g826) & (!g861)) + ((sk[112]) & (!g136) & (!g186) & (!g677) & (g826) & (!g861)) + ((sk[112]) & (!g136) & (!g186) & (g677) & (!g826) & (!g861)) + ((sk[112]) & (!g136) & (!g186) & (g677) & (g826) & (!g861)) + ((sk[112]) & (!g136) & (g186) & (!g677) & (g826) & (!g861)) + ((sk[112]) & (!g136) & (g186) & (g677) & (g826) & (!g861)) + ((sk[112]) & (g136) & (!g186) & (!g677) & (!g826) & (!g861)) + ((sk[112]) & (g136) & (!g186) & (!g677) & (g826) & (!g861)) + ((sk[112]) & (g136) & (g186) & (!g677) & (g826) & (!g861)));
	assign g863 = (((!sk[113]) & (!i_8_) & (!g108) & (g481) & (g465)) + ((!sk[113]) & (!i_8_) & (g108) & (!g481) & (!g465)) + ((!sk[113]) & (!i_8_) & (g108) & (!g481) & (g465)) + ((!sk[113]) & (!i_8_) & (g108) & (g481) & (!g465)) + ((!sk[113]) & (!i_8_) & (g108) & (g481) & (g465)) + ((!sk[113]) & (i_8_) & (!g108) & (g481) & (!g465)) + ((!sk[113]) & (i_8_) & (!g108) & (g481) & (g465)) + ((!sk[113]) & (i_8_) & (g108) & (!g481) & (!g465)) + ((!sk[113]) & (i_8_) & (g108) & (!g481) & (g465)) + ((!sk[113]) & (i_8_) & (g108) & (g481) & (!g465)) + ((!sk[113]) & (i_8_) & (g108) & (g481) & (g465)) + ((sk[113]) & (!i_8_) & (g108) & (!g481) & (!g465)) + ((sk[113]) & (!i_8_) & (g108) & (!g481) & (g465)) + ((sk[113]) & (i_8_) & (g108) & (!g481) & (!g465)) + ((sk[113]) & (i_8_) & (g108) & (!g481) & (g465)) + ((sk[113]) & (i_8_) & (g108) & (g481) & (!g465)));
	assign g864 = (((!i_8_) & (!g100) & (!g124) & (!g158) & (!sk[114]) & (g726)) + ((!i_8_) & (!g100) & (!g124) & (g158) & (!sk[114]) & (g726)) + ((!i_8_) & (!g100) & (g124) & (!g158) & (!sk[114]) & (g726)) + ((!i_8_) & (!g100) & (g124) & (g158) & (!sk[114]) & (g726)) + ((!i_8_) & (g100) & (!g124) & (!g158) & (!sk[114]) & (g726)) + ((!i_8_) & (g100) & (!g124) & (g158) & (!sk[114]) & (g726)) + ((!i_8_) & (g100) & (g124) & (!g158) & (!sk[114]) & (g726)) + ((!i_8_) & (g100) & (g124) & (!g158) & (sk[114]) & (!g726)) + ((!i_8_) & (g100) & (g124) & (g158) & (!sk[114]) & (g726)) + ((!i_8_) & (g100) & (g124) & (g158) & (sk[114]) & (!g726)) + ((i_8_) & (!g100) & (!g124) & (!g158) & (!sk[114]) & (!g726)) + ((i_8_) & (!g100) & (!g124) & (!g158) & (!sk[114]) & (g726)) + ((i_8_) & (!g100) & (!g124) & (g158) & (!sk[114]) & (!g726)) + ((i_8_) & (!g100) & (!g124) & (g158) & (!sk[114]) & (g726)) + ((i_8_) & (!g100) & (g124) & (!g158) & (!sk[114]) & (!g726)) + ((i_8_) & (!g100) & (g124) & (!g158) & (!sk[114]) & (g726)) + ((i_8_) & (!g100) & (g124) & (g158) & (!sk[114]) & (!g726)) + ((i_8_) & (!g100) & (g124) & (g158) & (!sk[114]) & (g726)) + ((i_8_) & (g100) & (!g124) & (!g158) & (!sk[114]) & (!g726)) + ((i_8_) & (g100) & (!g124) & (!g158) & (!sk[114]) & (g726)) + ((i_8_) & (g100) & (!g124) & (g158) & (!sk[114]) & (!g726)) + ((i_8_) & (g100) & (!g124) & (g158) & (!sk[114]) & (g726)) + ((i_8_) & (g100) & (!g124) & (g158) & (sk[114]) & (!g726)) + ((i_8_) & (g100) & (g124) & (!g158) & (!sk[114]) & (!g726)) + ((i_8_) & (g100) & (g124) & (!g158) & (!sk[114]) & (g726)) + ((i_8_) & (g100) & (g124) & (!g158) & (sk[114]) & (!g726)) + ((i_8_) & (g100) & (g124) & (g158) & (!sk[114]) & (!g726)) + ((i_8_) & (g100) & (g124) & (g158) & (!sk[114]) & (g726)) + ((i_8_) & (g100) & (g124) & (g158) & (sk[114]) & (!g726)));
	assign g865 = (((!g10) & (!sk[115]) & (!g145) & (!g136) & (!g127) & (g864)) + ((!g10) & (!sk[115]) & (!g145) & (!g136) & (g127) & (g864)) + ((!g10) & (!sk[115]) & (!g145) & (g136) & (!g127) & (g864)) + ((!g10) & (!sk[115]) & (!g145) & (g136) & (g127) & (g864)) + ((!g10) & (!sk[115]) & (g145) & (!g136) & (!g127) & (g864)) + ((!g10) & (!sk[115]) & (g145) & (!g136) & (g127) & (g864)) + ((!g10) & (!sk[115]) & (g145) & (g136) & (!g127) & (g864)) + ((!g10) & (!sk[115]) & (g145) & (g136) & (g127) & (g864)) + ((!g10) & (sk[115]) & (!g145) & (!g136) & (!g127) & (!g864)) + ((!g10) & (sk[115]) & (!g145) & (!g136) & (g127) & (!g864)) + ((!g10) & (sk[115]) & (!g145) & (g136) & (g127) & (!g864)) + ((!g10) & (sk[115]) & (g145) & (!g136) & (!g127) & (!g864)) + ((!g10) & (sk[115]) & (g145) & (!g136) & (g127) & (!g864)) + ((!g10) & (sk[115]) & (g145) & (g136) & (g127) & (!g864)) + ((g10) & (!sk[115]) & (!g145) & (!g136) & (!g127) & (!g864)) + ((g10) & (!sk[115]) & (!g145) & (!g136) & (!g127) & (g864)) + ((g10) & (!sk[115]) & (!g145) & (!g136) & (g127) & (!g864)) + ((g10) & (!sk[115]) & (!g145) & (!g136) & (g127) & (g864)) + ((g10) & (!sk[115]) & (!g145) & (g136) & (!g127) & (!g864)) + ((g10) & (!sk[115]) & (!g145) & (g136) & (!g127) & (g864)) + ((g10) & (!sk[115]) & (!g145) & (g136) & (g127) & (!g864)) + ((g10) & (!sk[115]) & (!g145) & (g136) & (g127) & (g864)) + ((g10) & (!sk[115]) & (g145) & (!g136) & (!g127) & (!g864)) + ((g10) & (!sk[115]) & (g145) & (!g136) & (!g127) & (g864)) + ((g10) & (!sk[115]) & (g145) & (!g136) & (g127) & (!g864)) + ((g10) & (!sk[115]) & (g145) & (!g136) & (g127) & (g864)) + ((g10) & (!sk[115]) & (g145) & (g136) & (!g127) & (!g864)) + ((g10) & (!sk[115]) & (g145) & (g136) & (!g127) & (g864)) + ((g10) & (!sk[115]) & (g145) & (g136) & (g127) & (!g864)) + ((g10) & (!sk[115]) & (g145) & (g136) & (g127) & (g864)) + ((g10) & (sk[115]) & (!g145) & (!g136) & (!g127) & (!g864)) + ((g10) & (sk[115]) & (!g145) & (!g136) & (g127) & (!g864)) + ((g10) & (sk[115]) & (!g145) & (g136) & (g127) & (!g864)));
	assign g866 = (((!i_8_) & (!g30) & (g5) & (!sk[116]) & (g40)) + ((!i_8_) & (g30) & (!g5) & (!sk[116]) & (!g40)) + ((!i_8_) & (g30) & (!g5) & (!sk[116]) & (g40)) + ((!i_8_) & (g30) & (g5) & (!sk[116]) & (!g40)) + ((!i_8_) & (g30) & (g5) & (!sk[116]) & (g40)) + ((!i_8_) & (g30) & (g5) & (sk[116]) & (g40)) + ((i_8_) & (!g30) & (g5) & (!sk[116]) & (!g40)) + ((i_8_) & (!g30) & (g5) & (!sk[116]) & (g40)) + ((i_8_) & (g30) & (!g5) & (!sk[116]) & (!g40)) + ((i_8_) & (g30) & (!g5) & (!sk[116]) & (g40)) + ((i_8_) & (g30) & (!g5) & (sk[116]) & (g40)) + ((i_8_) & (g30) & (g5) & (!sk[116]) & (!g40)) + ((i_8_) & (g30) & (g5) & (!sk[116]) & (g40)) + ((i_8_) & (g30) & (g5) & (sk[116]) & (g40)));
	assign g867 = (((!i_8_) & (!g100) & (!g120) & (!g746) & (!g103) & (!g866)) + ((!i_8_) & (!g100) & (!g120) & (!g746) & (g103) & (!g866)) + ((!i_8_) & (!g100) & (g120) & (!g746) & (!g103) & (!g866)) + ((!i_8_) & (!g100) & (g120) & (!g746) & (g103) & (!g866)) + ((!i_8_) & (!g100) & (g120) & (g746) & (!g103) & (!g866)) + ((!i_8_) & (!g100) & (g120) & (g746) & (g103) & (!g866)) + ((!i_8_) & (g100) & (!g120) & (!g746) & (!g103) & (!g866)) + ((!i_8_) & (g100) & (!g120) & (!g746) & (g103) & (!g866)) + ((!i_8_) & (g100) & (g120) & (!g746) & (!g103) & (!g866)) + ((!i_8_) & (g100) & (g120) & (!g746) & (g103) & (!g866)) + ((!i_8_) & (g100) & (g120) & (g746) & (!g103) & (!g866)) + ((!i_8_) & (g100) & (g120) & (g746) & (g103) & (!g866)) + ((i_8_) & (!g100) & (!g120) & (!g746) & (!g103) & (!g866)) + ((i_8_) & (!g100) & (!g120) & (!g746) & (g103) & (!g866)) + ((i_8_) & (!g100) & (g120) & (!g746) & (!g103) & (!g866)) + ((i_8_) & (!g100) & (g120) & (!g746) & (g103) & (!g866)) + ((i_8_) & (!g100) & (g120) & (g746) & (!g103) & (!g866)) + ((i_8_) & (!g100) & (g120) & (g746) & (g103) & (!g866)) + ((i_8_) & (g100) & (g120) & (!g746) & (g103) & (!g866)) + ((i_8_) & (g100) & (g120) & (g746) & (g103) & (!g866)));
	assign g868 = (((!g59) & (!g112) & (!g135) & (!g96) & (!g462) & (g867)) + ((!g59) & (!g112) & (!g135) & (!g96) & (g462) & (g867)) + ((!g59) & (!g112) & (!g135) & (g96) & (!g462) & (g867)) + ((!g59) & (!g112) & (!g135) & (g96) & (g462) & (g867)) + ((!g59) & (!g112) & (g135) & (!g96) & (g462) & (g867)) + ((!g59) & (!g112) & (g135) & (g96) & (g462) & (g867)) + ((!g59) & (g112) & (!g135) & (g96) & (g462) & (g867)) + ((!g59) & (g112) & (g135) & (g96) & (g462) & (g867)) + ((g59) & (!g112) & (!g135) & (g96) & (!g462) & (g867)) + ((g59) & (!g112) & (!g135) & (g96) & (g462) & (g867)) + ((g59) & (!g112) & (g135) & (g96) & (g462) & (g867)) + ((g59) & (g112) & (!g135) & (g96) & (g462) & (g867)) + ((g59) & (g112) & (g135) & (g96) & (g462) & (g867)));
	assign g869 = (((!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!g91) & (g711)) + ((!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g91) & (g711)) + ((!i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!g91) & (!g711)) + ((!i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!g91) & (g711)) + ((!i_11_) & (i_9_) & (i_10_) & (i_15_) & (!g91) & (g711)) + ((!i_11_) & (i_9_) & (i_10_) & (i_15_) & (g91) & (g711)) + ((i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (!g91) & (!g711)) + ((i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (!g91) & (g711)) + ((i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!g91) & (!g711)) + ((i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!g91) & (g711)) + ((i_11_) & (i_9_) & (i_10_) & (i_15_) & (!g91) & (g711)) + ((i_11_) & (i_9_) & (i_10_) & (i_15_) & (g91) & (g711)));
	assign g870 = (((!g16) & (!g243) & (!sk[120]) & (g619) & (g869)) + ((!g16) & (g243) & (!sk[120]) & (!g619) & (!g869)) + ((!g16) & (g243) & (!sk[120]) & (!g619) & (g869)) + ((!g16) & (g243) & (!sk[120]) & (g619) & (!g869)) + ((!g16) & (g243) & (!sk[120]) & (g619) & (g869)) + ((!g16) & (g243) & (sk[120]) & (!g619) & (!g869)) + ((!g16) & (g243) & (sk[120]) & (!g619) & (g869)) + ((!g16) & (g243) & (sk[120]) & (g619) & (!g869)) + ((!g16) & (g243) & (sk[120]) & (g619) & (g869)) + ((g16) & (!g243) & (!sk[120]) & (g619) & (!g869)) + ((g16) & (!g243) & (!sk[120]) & (g619) & (g869)) + ((g16) & (g243) & (!sk[120]) & (!g619) & (!g869)) + ((g16) & (g243) & (!sk[120]) & (!g619) & (g869)) + ((g16) & (g243) & (!sk[120]) & (g619) & (!g869)) + ((g16) & (g243) & (!sk[120]) & (g619) & (g869)) + ((g16) & (g243) & (sk[120]) & (!g619) & (g869)) + ((g16) & (g243) & (sk[120]) & (g619) & (!g869)) + ((g16) & (g243) & (sk[120]) & (g619) & (g869)));
	assign g871 = (((!g251) & (!g132) & (!sk[121]) & (!g122) & (!g711) & (g870)) + ((!g251) & (!g132) & (!sk[121]) & (!g122) & (g711) & (g870)) + ((!g251) & (!g132) & (!sk[121]) & (g122) & (!g711) & (g870)) + ((!g251) & (!g132) & (!sk[121]) & (g122) & (g711) & (g870)) + ((!g251) & (!g132) & (sk[121]) & (!g122) & (!g711) & (!g870)) + ((!g251) & (!g132) & (sk[121]) & (!g122) & (g711) & (!g870)) + ((!g251) & (!g132) & (sk[121]) & (g122) & (!g711) & (!g870)) + ((!g251) & (!g132) & (sk[121]) & (g122) & (g711) & (!g870)) + ((!g251) & (g132) & (!sk[121]) & (!g122) & (!g711) & (g870)) + ((!g251) & (g132) & (!sk[121]) & (!g122) & (g711) & (g870)) + ((!g251) & (g132) & (!sk[121]) & (g122) & (!g711) & (g870)) + ((!g251) & (g132) & (!sk[121]) & (g122) & (g711) & (g870)) + ((!g251) & (g132) & (sk[121]) & (!g122) & (!g711) & (!g870)) + ((!g251) & (g132) & (sk[121]) & (!g122) & (g711) & (!g870)) + ((!g251) & (g132) & (sk[121]) & (g122) & (!g711) & (!g870)) + ((!g251) & (g132) & (sk[121]) & (g122) & (g711) & (!g870)) + ((g251) & (!g132) & (!sk[121]) & (!g122) & (!g711) & (!g870)) + ((g251) & (!g132) & (!sk[121]) & (!g122) & (!g711) & (g870)) + ((g251) & (!g132) & (!sk[121]) & (!g122) & (g711) & (!g870)) + ((g251) & (!g132) & (!sk[121]) & (!g122) & (g711) & (g870)) + ((g251) & (!g132) & (!sk[121]) & (g122) & (!g711) & (!g870)) + ((g251) & (!g132) & (!sk[121]) & (g122) & (!g711) & (g870)) + ((g251) & (!g132) & (!sk[121]) & (g122) & (g711) & (!g870)) + ((g251) & (!g132) & (!sk[121]) & (g122) & (g711) & (g870)) + ((g251) & (g132) & (!sk[121]) & (!g122) & (!g711) & (!g870)) + ((g251) & (g132) & (!sk[121]) & (!g122) & (!g711) & (g870)) + ((g251) & (g132) & (!sk[121]) & (!g122) & (g711) & (!g870)) + ((g251) & (g132) & (!sk[121]) & (!g122) & (g711) & (g870)) + ((g251) & (g132) & (!sk[121]) & (g122) & (!g711) & (!g870)) + ((g251) & (g132) & (!sk[121]) & (g122) & (!g711) & (g870)) + ((g251) & (g132) & (!sk[121]) & (g122) & (g711) & (!g870)) + ((g251) & (g132) & (!sk[121]) & (g122) & (g711) & (g870)) + ((g251) & (g132) & (sk[121]) & (!g122) & (!g711) & (!g870)) + ((g251) & (g132) & (sk[121]) & (g122) & (!g711) & (!g870)) + ((g251) & (g132) & (sk[121]) & (g122) & (g711) & (!g870)));
	assign g872 = (((!g99) & (!g132) & (!g863) & (g865) & (g868) & (g871)) + ((!g99) & (g132) & (!g863) & (g865) & (g868) & (g871)) + ((g99) & (g132) & (!g863) & (g865) & (g868) & (g871)));
	assign g873 = (((!g82) & (!sk[123]) & (!g860) & (g862) & (g872)) + ((!g82) & (!sk[123]) & (g860) & (!g862) & (!g872)) + ((!g82) & (!sk[123]) & (g860) & (!g862) & (g872)) + ((!g82) & (!sk[123]) & (g860) & (g862) & (!g872)) + ((!g82) & (!sk[123]) & (g860) & (g862) & (g872)) + ((g82) & (!sk[123]) & (!g860) & (g862) & (!g872)) + ((g82) & (!sk[123]) & (!g860) & (g862) & (g872)) + ((g82) & (!sk[123]) & (g860) & (!g862) & (!g872)) + ((g82) & (!sk[123]) & (g860) & (!g862) & (g872)) + ((g82) & (!sk[123]) & (g860) & (g862) & (!g872)) + ((g82) & (!sk[123]) & (g860) & (g862) & (g872)) + ((g82) & (sk[123]) & (g860) & (g862) & (g872)));
	assign g874 = (((!g73) & (!g169) & (!g521) & (!g759) & (!g858) & (!g873)) + ((!g73) & (!g169) & (!g521) & (!g759) & (!g858) & (g873)) + ((!g73) & (!g169) & (!g521) & (!g759) & (g858) & (!g873)) + ((!g73) & (!g169) & (!g521) & (!g759) & (g858) & (g873)) + ((!g73) & (!g169) & (!g521) & (g759) & (!g858) & (!g873)) + ((!g73) & (!g169) & (!g521) & (g759) & (!g858) & (g873)) + ((!g73) & (!g169) & (!g521) & (g759) & (g858) & (!g873)) + ((!g73) & (!g169) & (!g521) & (g759) & (g858) & (g873)) + ((!g73) & (!g169) & (g521) & (!g759) & (!g858) & (!g873)) + ((!g73) & (!g169) & (g521) & (!g759) & (!g858) & (g873)) + ((!g73) & (!g169) & (g521) & (!g759) & (g858) & (!g873)) + ((!g73) & (!g169) & (g521) & (!g759) & (g858) & (g873)) + ((!g73) & (!g169) & (g521) & (g759) & (!g858) & (!g873)) + ((!g73) & (!g169) & (g521) & (g759) & (!g858) & (g873)) + ((!g73) & (!g169) & (g521) & (g759) & (g858) & (!g873)) + ((!g73) & (!g169) & (g521) & (g759) & (g858) & (g873)) + ((!g73) & (g169) & (!g521) & (!g759) & (!g858) & (!g873)) + ((!g73) & (g169) & (!g521) & (!g759) & (!g858) & (g873)) + ((!g73) & (g169) & (!g521) & (!g759) & (g858) & (!g873)) + ((!g73) & (g169) & (!g521) & (!g759) & (g858) & (g873)) + ((!g73) & (g169) & (!g521) & (g759) & (!g858) & (!g873)) + ((!g73) & (g169) & (!g521) & (g759) & (!g858) & (g873)) + ((!g73) & (g169) & (!g521) & (g759) & (g858) & (!g873)) + ((!g73) & (g169) & (!g521) & (g759) & (g858) & (g873)) + ((!g73) & (g169) & (g521) & (!g759) & (!g858) & (!g873)) + ((!g73) & (g169) & (g521) & (!g759) & (!g858) & (g873)) + ((!g73) & (g169) & (g521) & (!g759) & (g858) & (!g873)) + ((!g73) & (g169) & (g521) & (!g759) & (g858) & (g873)) + ((!g73) & (g169) & (g521) & (g759) & (!g858) & (!g873)) + ((!g73) & (g169) & (g521) & (g759) & (!g858) & (g873)) + ((!g73) & (g169) & (g521) & (g759) & (g858) & (!g873)) + ((!g73) & (g169) & (g521) & (g759) & (g858) & (g873)) + ((g73) & (g169) & (g521) & (g759) & (g858) & (g873)));
	assign g875 = (((!i_15_) & (sk[125]) & (g7)) + ((i_15_) & (!sk[125]) & (!g7)) + ((i_15_) & (!sk[125]) & (g7)));
	assign g876 = (((!i_11_) & (!i_9_) & (i_10_) & (!sk[126]) & (g875)) + ((!i_11_) & (!i_9_) & (i_10_) & (sk[126]) & (g875)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[126]) & (!g875)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[126]) & (g875)) + ((!i_11_) & (i_9_) & (!i_10_) & (sk[126]) & (g875)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[126]) & (!g875)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[126]) & (g875)) + ((i_11_) & (!i_9_) & (!i_10_) & (sk[126]) & (g875)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[126]) & (!g875)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[126]) & (g875)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[126]) & (!g875)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[126]) & (g875)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[126]) & (!g875)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[126]) & (g875)));
	assign g877 = (((!i_11_) & (!i_9_) & (!sk[127]) & (i_10_) & (g875)) + ((!i_11_) & (!i_9_) & (sk[127]) & (!i_10_) & (g875)) + ((!i_11_) & (i_9_) & (!sk[127]) & (!i_10_) & (!g875)) + ((!i_11_) & (i_9_) & (!sk[127]) & (!i_10_) & (g875)) + ((!i_11_) & (i_9_) & (!sk[127]) & (i_10_) & (!g875)) + ((!i_11_) & (i_9_) & (!sk[127]) & (i_10_) & (g875)) + ((i_11_) & (!i_9_) & (!sk[127]) & (i_10_) & (!g875)) + ((i_11_) & (!i_9_) & (!sk[127]) & (i_10_) & (g875)) + ((i_11_) & (!i_9_) & (sk[127]) & (i_10_) & (g875)) + ((i_11_) & (i_9_) & (!sk[127]) & (!i_10_) & (!g875)) + ((i_11_) & (i_9_) & (!sk[127]) & (!i_10_) & (g875)) + ((i_11_) & (i_9_) & (!sk[127]) & (i_10_) & (!g875)) + ((i_11_) & (i_9_) & (!sk[127]) & (i_10_) & (g875)));
	assign g878 = (((!g99) & (!sk[0]) & (!g251) & (g285) & (g877)) + ((!g99) & (!sk[0]) & (g251) & (!g285) & (!g877)) + ((!g99) & (!sk[0]) & (g251) & (!g285) & (g877)) + ((!g99) & (!sk[0]) & (g251) & (g285) & (!g877)) + ((!g99) & (!sk[0]) & (g251) & (g285) & (g877)) + ((!g99) & (sk[0]) & (!g251) & (!g285) & (g877)) + ((!g99) & (sk[0]) & (g251) & (!g285) & (g877)) + ((!g99) & (sk[0]) & (g251) & (g285) & (g877)) + ((g99) & (!sk[0]) & (!g251) & (g285) & (!g877)) + ((g99) & (!sk[0]) & (!g251) & (g285) & (g877)) + ((g99) & (!sk[0]) & (g251) & (!g285) & (!g877)) + ((g99) & (!sk[0]) & (g251) & (!g285) & (g877)) + ((g99) & (!sk[0]) & (g251) & (g285) & (!g877)) + ((g99) & (!sk[0]) & (g251) & (g285) & (g877)) + ((g99) & (sk[0]) & (!g251) & (!g285) & (g877)) + ((g99) & (sk[0]) & (!g251) & (g285) & (g877)) + ((g99) & (sk[0]) & (g251) & (!g285) & (g877)) + ((g99) & (sk[0]) & (g251) & (g285) & (g877)));
	assign g879 = (((!g212) & (!sk[1]) & (!g568) & (g876) & (g878)) + ((!g212) & (!sk[1]) & (g568) & (!g876) & (!g878)) + ((!g212) & (!sk[1]) & (g568) & (!g876) & (g878)) + ((!g212) & (!sk[1]) & (g568) & (g876) & (!g878)) + ((!g212) & (!sk[1]) & (g568) & (g876) & (g878)) + ((!g212) & (sk[1]) & (g568) & (!g876) & (!g878)) + ((g212) & (!sk[1]) & (!g568) & (g876) & (!g878)) + ((g212) & (!sk[1]) & (!g568) & (g876) & (g878)) + ((g212) & (!sk[1]) & (g568) & (!g876) & (!g878)) + ((g212) & (!sk[1]) & (g568) & (!g876) & (g878)) + ((g212) & (!sk[1]) & (g568) & (g876) & (!g878)) + ((g212) & (!sk[1]) & (g568) & (g876) & (g878)) + ((g212) & (sk[1]) & (g568) & (!g876) & (!g878)) + ((g212) & (sk[1]) & (g568) & (g876) & (!g878)));
	assign g880 = (((!sk[2]) & (g569) & (!g580) & (!g582)) + ((!sk[2]) & (g569) & (!g580) & (g582)) + ((!sk[2]) & (g569) & (g580) & (!g582)) + ((!sk[2]) & (g569) & (g580) & (g582)) + ((sk[2]) & (!g569) & (g580) & (g582)));
	assign g881 = (((!sk[3]) & (g7) & (!g104)) + ((!sk[3]) & (g7) & (g104)) + ((sk[3]) & (g7) & (g104)));
	assign g882 = (((!sk[4]) & (g551) & (!g734)) + ((!sk[4]) & (g551) & (g734)) + ((sk[4]) & (!g551) & (!g734)));
	assign g883 = (((!sk[5]) & (!i_8_) & (!g23) & (!g206) & (!g100) & (g561)) + ((!sk[5]) & (!i_8_) & (!g23) & (!g206) & (g100) & (g561)) + ((!sk[5]) & (!i_8_) & (!g23) & (g206) & (!g100) & (g561)) + ((!sk[5]) & (!i_8_) & (!g23) & (g206) & (g100) & (g561)) + ((!sk[5]) & (!i_8_) & (g23) & (!g206) & (!g100) & (g561)) + ((!sk[5]) & (!i_8_) & (g23) & (!g206) & (g100) & (g561)) + ((!sk[5]) & (!i_8_) & (g23) & (g206) & (!g100) & (g561)) + ((!sk[5]) & (!i_8_) & (g23) & (g206) & (g100) & (g561)) + ((!sk[5]) & (i_8_) & (!g23) & (!g206) & (!g100) & (!g561)) + ((!sk[5]) & (i_8_) & (!g23) & (!g206) & (!g100) & (g561)) + ((!sk[5]) & (i_8_) & (!g23) & (!g206) & (g100) & (!g561)) + ((!sk[5]) & (i_8_) & (!g23) & (!g206) & (g100) & (g561)) + ((!sk[5]) & (i_8_) & (!g23) & (g206) & (!g100) & (!g561)) + ((!sk[5]) & (i_8_) & (!g23) & (g206) & (!g100) & (g561)) + ((!sk[5]) & (i_8_) & (!g23) & (g206) & (g100) & (!g561)) + ((!sk[5]) & (i_8_) & (!g23) & (g206) & (g100) & (g561)) + ((!sk[5]) & (i_8_) & (g23) & (!g206) & (!g100) & (!g561)) + ((!sk[5]) & (i_8_) & (g23) & (!g206) & (!g100) & (g561)) + ((!sk[5]) & (i_8_) & (g23) & (!g206) & (g100) & (!g561)) + ((!sk[5]) & (i_8_) & (g23) & (!g206) & (g100) & (g561)) + ((!sk[5]) & (i_8_) & (g23) & (g206) & (!g100) & (!g561)) + ((!sk[5]) & (i_8_) & (g23) & (g206) & (!g100) & (g561)) + ((!sk[5]) & (i_8_) & (g23) & (g206) & (g100) & (!g561)) + ((!sk[5]) & (i_8_) & (g23) & (g206) & (g100) & (g561)) + ((sk[5]) & (!i_8_) & (!g23) & (!g206) & (!g100) & (!g561)) + ((sk[5]) & (!i_8_) & (!g23) & (!g206) & (g100) & (!g561)) + ((sk[5]) & (!i_8_) & (!g23) & (g206) & (!g100) & (!g561)) + ((sk[5]) & (!i_8_) & (!g23) & (g206) & (g100) & (!g561)) + ((sk[5]) & (i_8_) & (!g23) & (!g206) & (!g100) & (!g561)) + ((sk[5]) & (i_8_) & (!g23) & (g206) & (!g100) & (!g561)) + ((sk[5]) & (i_8_) & (!g23) & (g206) & (g100) & (!g561)));
	assign g884 = (((!g101) & (!g185) & (!g881) & (!sk[6]) & (!g882) & (g883)) + ((!g101) & (!g185) & (!g881) & (!sk[6]) & (g882) & (g883)) + ((!g101) & (!g185) & (g881) & (!sk[6]) & (!g882) & (g883)) + ((!g101) & (!g185) & (g881) & (!sk[6]) & (g882) & (g883)) + ((!g101) & (g185) & (!g881) & (!sk[6]) & (!g882) & (g883)) + ((!g101) & (g185) & (!g881) & (!sk[6]) & (g882) & (g883)) + ((!g101) & (g185) & (g881) & (!sk[6]) & (!g882) & (g883)) + ((!g101) & (g185) & (g881) & (!sk[6]) & (g882) & (g883)) + ((g101) & (!g185) & (!g881) & (!sk[6]) & (!g882) & (!g883)) + ((g101) & (!g185) & (!g881) & (!sk[6]) & (!g882) & (g883)) + ((g101) & (!g185) & (!g881) & (!sk[6]) & (g882) & (!g883)) + ((g101) & (!g185) & (!g881) & (!sk[6]) & (g882) & (g883)) + ((g101) & (!g185) & (!g881) & (sk[6]) & (!g882) & (!g883)) + ((g101) & (!g185) & (!g881) & (sk[6]) & (!g882) & (g883)) + ((g101) & (!g185) & (!g881) & (sk[6]) & (g882) & (!g883)) + ((g101) & (!g185) & (!g881) & (sk[6]) & (g882) & (g883)) + ((g101) & (!g185) & (g881) & (!sk[6]) & (!g882) & (!g883)) + ((g101) & (!g185) & (g881) & (!sk[6]) & (!g882) & (g883)) + ((g101) & (!g185) & (g881) & (!sk[6]) & (g882) & (!g883)) + ((g101) & (!g185) & (g881) & (!sk[6]) & (g882) & (g883)) + ((g101) & (!g185) & (g881) & (sk[6]) & (!g882) & (!g883)) + ((g101) & (!g185) & (g881) & (sk[6]) & (!g882) & (g883)) + ((g101) & (!g185) & (g881) & (sk[6]) & (g882) & (!g883)) + ((g101) & (!g185) & (g881) & (sk[6]) & (g882) & (g883)) + ((g101) & (g185) & (!g881) & (!sk[6]) & (!g882) & (!g883)) + ((g101) & (g185) & (!g881) & (!sk[6]) & (!g882) & (g883)) + ((g101) & (g185) & (!g881) & (!sk[6]) & (g882) & (!g883)) + ((g101) & (g185) & (!g881) & (!sk[6]) & (g882) & (g883)) + ((g101) & (g185) & (!g881) & (sk[6]) & (!g882) & (!g883)) + ((g101) & (g185) & (!g881) & (sk[6]) & (!g882) & (g883)) + ((g101) & (g185) & (!g881) & (sk[6]) & (g882) & (!g883)) + ((g101) & (g185) & (g881) & (!sk[6]) & (!g882) & (!g883)) + ((g101) & (g185) & (g881) & (!sk[6]) & (!g882) & (g883)) + ((g101) & (g185) & (g881) & (!sk[6]) & (g882) & (!g883)) + ((g101) & (g185) & (g881) & (!sk[6]) & (g882) & (g883)) + ((g101) & (g185) & (g881) & (sk[6]) & (!g882) & (!g883)) + ((g101) & (g185) & (g881) & (sk[6]) & (!g882) & (g883)) + ((g101) & (g185) & (g881) & (sk[6]) & (g882) & (!g883)) + ((g101) & (g185) & (g881) & (sk[6]) & (g882) & (g883)));
	assign g885 = (((!sk[7]) & (!i_11_) & (!i_9_) & (!i_10_) & (!g323) & (g875)) + ((!sk[7]) & (!i_11_) & (!i_9_) & (!i_10_) & (g323) & (g875)) + ((!sk[7]) & (!i_11_) & (!i_9_) & (i_10_) & (!g323) & (g875)) + ((!sk[7]) & (!i_11_) & (!i_9_) & (i_10_) & (g323) & (g875)) + ((!sk[7]) & (!i_11_) & (i_9_) & (!i_10_) & (!g323) & (g875)) + ((!sk[7]) & (!i_11_) & (i_9_) & (!i_10_) & (g323) & (g875)) + ((!sk[7]) & (!i_11_) & (i_9_) & (i_10_) & (!g323) & (g875)) + ((!sk[7]) & (!i_11_) & (i_9_) & (i_10_) & (g323) & (g875)) + ((!sk[7]) & (i_11_) & (!i_9_) & (!i_10_) & (!g323) & (!g875)) + ((!sk[7]) & (i_11_) & (!i_9_) & (!i_10_) & (!g323) & (g875)) + ((!sk[7]) & (i_11_) & (!i_9_) & (!i_10_) & (g323) & (!g875)) + ((!sk[7]) & (i_11_) & (!i_9_) & (!i_10_) & (g323) & (g875)) + ((!sk[7]) & (i_11_) & (!i_9_) & (i_10_) & (!g323) & (!g875)) + ((!sk[7]) & (i_11_) & (!i_9_) & (i_10_) & (!g323) & (g875)) + ((!sk[7]) & (i_11_) & (!i_9_) & (i_10_) & (g323) & (!g875)) + ((!sk[7]) & (i_11_) & (!i_9_) & (i_10_) & (g323) & (g875)) + ((!sk[7]) & (i_11_) & (i_9_) & (!i_10_) & (!g323) & (!g875)) + ((!sk[7]) & (i_11_) & (i_9_) & (!i_10_) & (!g323) & (g875)) + ((!sk[7]) & (i_11_) & (i_9_) & (!i_10_) & (g323) & (!g875)) + ((!sk[7]) & (i_11_) & (i_9_) & (!i_10_) & (g323) & (g875)) + ((!sk[7]) & (i_11_) & (i_9_) & (i_10_) & (!g323) & (!g875)) + ((!sk[7]) & (i_11_) & (i_9_) & (i_10_) & (!g323) & (g875)) + ((!sk[7]) & (i_11_) & (i_9_) & (i_10_) & (g323) & (!g875)) + ((!sk[7]) & (i_11_) & (i_9_) & (i_10_) & (g323) & (g875)) + ((sk[7]) & (!i_11_) & (i_9_) & (!i_10_) & (g323) & (g875)) + ((sk[7]) & (i_11_) & (i_9_) & (i_10_) & (g323) & (g875)));
	assign g886 = (((!i_8_) & (!g10) & (!sk[8]) & (!g66) & (!g100) & (g108)) + ((!i_8_) & (!g10) & (!sk[8]) & (!g66) & (g100) & (g108)) + ((!i_8_) & (!g10) & (!sk[8]) & (g66) & (!g100) & (g108)) + ((!i_8_) & (!g10) & (!sk[8]) & (g66) & (g100) & (g108)) + ((!i_8_) & (g10) & (!sk[8]) & (!g66) & (!g100) & (g108)) + ((!i_8_) & (g10) & (!sk[8]) & (!g66) & (g100) & (g108)) + ((!i_8_) & (g10) & (!sk[8]) & (g66) & (!g100) & (g108)) + ((!i_8_) & (g10) & (!sk[8]) & (g66) & (g100) & (g108)) + ((i_8_) & (!g10) & (!sk[8]) & (!g66) & (!g100) & (!g108)) + ((i_8_) & (!g10) & (!sk[8]) & (!g66) & (!g100) & (g108)) + ((i_8_) & (!g10) & (!sk[8]) & (!g66) & (g100) & (!g108)) + ((i_8_) & (!g10) & (!sk[8]) & (!g66) & (g100) & (g108)) + ((i_8_) & (!g10) & (!sk[8]) & (g66) & (!g100) & (!g108)) + ((i_8_) & (!g10) & (!sk[8]) & (g66) & (!g100) & (g108)) + ((i_8_) & (!g10) & (!sk[8]) & (g66) & (g100) & (!g108)) + ((i_8_) & (!g10) & (!sk[8]) & (g66) & (g100) & (g108)) + ((i_8_) & (!g10) & (sk[8]) & (g66) & (!g100) & (g108)) + ((i_8_) & (!g10) & (sk[8]) & (g66) & (g100) & (!g108)) + ((i_8_) & (!g10) & (sk[8]) & (g66) & (g100) & (g108)) + ((i_8_) & (g10) & (!sk[8]) & (!g66) & (!g100) & (!g108)) + ((i_8_) & (g10) & (!sk[8]) & (!g66) & (!g100) & (g108)) + ((i_8_) & (g10) & (!sk[8]) & (!g66) & (g100) & (!g108)) + ((i_8_) & (g10) & (!sk[8]) & (!g66) & (g100) & (g108)) + ((i_8_) & (g10) & (!sk[8]) & (g66) & (!g100) & (!g108)) + ((i_8_) & (g10) & (!sk[8]) & (g66) & (!g100) & (g108)) + ((i_8_) & (g10) & (!sk[8]) & (g66) & (g100) & (!g108)) + ((i_8_) & (g10) & (!sk[8]) & (g66) & (g100) & (g108)) + ((i_8_) & (g10) & (sk[8]) & (!g66) & (!g100) & (g108)) + ((i_8_) & (g10) & (sk[8]) & (!g66) & (g100) & (g108)) + ((i_8_) & (g10) & (sk[8]) & (g66) & (!g100) & (g108)) + ((i_8_) & (g10) & (sk[8]) & (g66) & (g100) & (!g108)) + ((i_8_) & (g10) & (sk[8]) & (g66) & (g100) & (g108)));
	assign g887 = (((!g181) & (sk[9]) & (!g548) & (!g671)) + ((g181) & (!sk[9]) & (!g548) & (!g671)) + ((g181) & (!sk[9]) & (!g548) & (g671)) + ((g181) & (!sk[9]) & (g548) & (!g671)) + ((g181) & (!sk[9]) & (g548) & (g671)));
	assign g888 = (((!g8) & (!g221) & (!g323) & (!sk[10]) & (!g544) & (g887)) + ((!g8) & (!g221) & (!g323) & (!sk[10]) & (g544) & (g887)) + ((!g8) & (!g221) & (g323) & (!sk[10]) & (!g544) & (g887)) + ((!g8) & (!g221) & (g323) & (!sk[10]) & (g544) & (g887)) + ((!g8) & (!g221) & (g323) & (sk[10]) & (!g544) & (!g887)) + ((!g8) & (!g221) & (g323) & (sk[10]) & (!g544) & (g887)) + ((!g8) & (!g221) & (g323) & (sk[10]) & (g544) & (!g887)) + ((!g8) & (!g221) & (g323) & (sk[10]) & (g544) & (g887)) + ((!g8) & (g221) & (!g323) & (!sk[10]) & (!g544) & (g887)) + ((!g8) & (g221) & (!g323) & (!sk[10]) & (g544) & (g887)) + ((!g8) & (g221) & (g323) & (!sk[10]) & (!g544) & (g887)) + ((!g8) & (g221) & (g323) & (!sk[10]) & (g544) & (g887)) + ((!g8) & (g221) & (g323) & (sk[10]) & (!g544) & (!g887)) + ((!g8) & (g221) & (g323) & (sk[10]) & (!g544) & (g887)) + ((!g8) & (g221) & (g323) & (sk[10]) & (g544) & (!g887)) + ((!g8) & (g221) & (g323) & (sk[10]) & (g544) & (g887)) + ((g8) & (!g221) & (!g323) & (!sk[10]) & (!g544) & (!g887)) + ((g8) & (!g221) & (!g323) & (!sk[10]) & (!g544) & (g887)) + ((g8) & (!g221) & (!g323) & (!sk[10]) & (g544) & (!g887)) + ((g8) & (!g221) & (!g323) & (!sk[10]) & (g544) & (g887)) + ((g8) & (!g221) & (g323) & (!sk[10]) & (!g544) & (!g887)) + ((g8) & (!g221) & (g323) & (!sk[10]) & (!g544) & (g887)) + ((g8) & (!g221) & (g323) & (!sk[10]) & (g544) & (!g887)) + ((g8) & (!g221) & (g323) & (!sk[10]) & (g544) & (g887)) + ((g8) & (!g221) & (g323) & (sk[10]) & (!g544) & (!g887)) + ((g8) & (!g221) & (g323) & (sk[10]) & (!g544) & (g887)) + ((g8) & (!g221) & (g323) & (sk[10]) & (g544) & (!g887)) + ((g8) & (!g221) & (g323) & (sk[10]) & (g544) & (g887)) + ((g8) & (g221) & (!g323) & (!sk[10]) & (!g544) & (!g887)) + ((g8) & (g221) & (!g323) & (!sk[10]) & (!g544) & (g887)) + ((g8) & (g221) & (!g323) & (!sk[10]) & (g544) & (!g887)) + ((g8) & (g221) & (!g323) & (!sk[10]) & (g544) & (g887)) + ((g8) & (g221) & (g323) & (!sk[10]) & (!g544) & (!g887)) + ((g8) & (g221) & (g323) & (!sk[10]) & (!g544) & (g887)) + ((g8) & (g221) & (g323) & (!sk[10]) & (g544) & (!g887)) + ((g8) & (g221) & (g323) & (!sk[10]) & (g544) & (g887)) + ((g8) & (g221) & (g323) & (sk[10]) & (!g544) & (!g887)) + ((g8) & (g221) & (g323) & (sk[10]) & (!g544) & (g887)) + ((g8) & (g221) & (g323) & (sk[10]) & (g544) & (!g887)));
	assign g889 = (((!g136) & (!g609) & (!g881) & (!g885) & (!g886) & (!g888)) + ((!g136) & (!g609) & (g881) & (!g885) & (!g886) & (!g888)) + ((g136) & (!g609) & (!g881) & (!g885) & (!g886) & (!g888)));
	assign g890 = (((!g695) & (!g697) & (g699) & (g700) & (!g884) & (g889)));
	assign g891 = (((!sk[13]) & (g270) & (!g554) & (!g669)) + ((!sk[13]) & (g270) & (!g554) & (g669)) + ((!sk[13]) & (g270) & (g554) & (!g669)) + ((!sk[13]) & (g270) & (g554) & (g669)) + ((sk[13]) & (g270) & (!g554) & (g669)));
	assign g892 = (((!sk[14]) & (i_8_) & (!i_7_) & (!g98)) + ((!sk[14]) & (i_8_) & (!i_7_) & (g98)) + ((!sk[14]) & (i_8_) & (i_7_) & (!g98)) + ((!sk[14]) & (i_8_) & (i_7_) & (g98)) + ((sk[14]) & (i_8_) & (i_7_) & (g98)));
	assign g893 = (((!i_6_) & (!sk[15]) & (!g43) & (!g131) & (!g461) & (g892)) + ((!i_6_) & (!sk[15]) & (!g43) & (!g131) & (g461) & (g892)) + ((!i_6_) & (!sk[15]) & (!g43) & (g131) & (!g461) & (g892)) + ((!i_6_) & (!sk[15]) & (!g43) & (g131) & (g461) & (g892)) + ((!i_6_) & (!sk[15]) & (g43) & (!g131) & (!g461) & (g892)) + ((!i_6_) & (!sk[15]) & (g43) & (!g131) & (g461) & (g892)) + ((!i_6_) & (!sk[15]) & (g43) & (g131) & (!g461) & (g892)) + ((!i_6_) & (!sk[15]) & (g43) & (g131) & (g461) & (g892)) + ((!i_6_) & (sk[15]) & (!g43) & (g131) & (g461) & (g892)) + ((!i_6_) & (sk[15]) & (g43) & (g131) & (g461) & (g892)) + ((i_6_) & (!sk[15]) & (!g43) & (!g131) & (!g461) & (!g892)) + ((i_6_) & (!sk[15]) & (!g43) & (!g131) & (!g461) & (g892)) + ((i_6_) & (!sk[15]) & (!g43) & (!g131) & (g461) & (!g892)) + ((i_6_) & (!sk[15]) & (!g43) & (!g131) & (g461) & (g892)) + ((i_6_) & (!sk[15]) & (!g43) & (g131) & (!g461) & (!g892)) + ((i_6_) & (!sk[15]) & (!g43) & (g131) & (!g461) & (g892)) + ((i_6_) & (!sk[15]) & (!g43) & (g131) & (g461) & (!g892)) + ((i_6_) & (!sk[15]) & (!g43) & (g131) & (g461) & (g892)) + ((i_6_) & (!sk[15]) & (g43) & (!g131) & (!g461) & (!g892)) + ((i_6_) & (!sk[15]) & (g43) & (!g131) & (!g461) & (g892)) + ((i_6_) & (!sk[15]) & (g43) & (!g131) & (g461) & (!g892)) + ((i_6_) & (!sk[15]) & (g43) & (!g131) & (g461) & (g892)) + ((i_6_) & (!sk[15]) & (g43) & (g131) & (!g461) & (!g892)) + ((i_6_) & (!sk[15]) & (g43) & (g131) & (!g461) & (g892)) + ((i_6_) & (!sk[15]) & (g43) & (g131) & (g461) & (!g892)) + ((i_6_) & (!sk[15]) & (g43) & (g131) & (g461) & (g892)) + ((i_6_) & (sk[15]) & (g43) & (!g131) & (!g461) & (g892)) + ((i_6_) & (sk[15]) & (g43) & (!g131) & (g461) & (g892)) + ((i_6_) & (sk[15]) & (g43) & (g131) & (!g461) & (g892)) + ((i_6_) & (sk[15]) & (g43) & (g131) & (g461) & (g892)));
	assign g894 = (((!g101) & (!g136) & (!sk[16]) & (!g576) & (!g891) & (g893)) + ((!g101) & (!g136) & (!sk[16]) & (!g576) & (g891) & (g893)) + ((!g101) & (!g136) & (!sk[16]) & (g576) & (!g891) & (g893)) + ((!g101) & (!g136) & (!sk[16]) & (g576) & (g891) & (g893)) + ((!g101) & (!g136) & (sk[16]) & (!g576) & (!g891) & (!g893)) + ((!g101) & (!g136) & (sk[16]) & (!g576) & (g891) & (!g893)) + ((!g101) & (!g136) & (sk[16]) & (g576) & (!g891) & (!g893)) + ((!g101) & (!g136) & (sk[16]) & (g576) & (g891) & (!g893)) + ((!g101) & (g136) & (!sk[16]) & (!g576) & (!g891) & (g893)) + ((!g101) & (g136) & (!sk[16]) & (!g576) & (g891) & (g893)) + ((!g101) & (g136) & (!sk[16]) & (g576) & (!g891) & (g893)) + ((!g101) & (g136) & (!sk[16]) & (g576) & (g891) & (g893)) + ((!g101) & (g136) & (sk[16]) & (g576) & (!g891) & (!g893)) + ((!g101) & (g136) & (sk[16]) & (g576) & (g891) & (!g893)) + ((g101) & (!g136) & (!sk[16]) & (!g576) & (!g891) & (!g893)) + ((g101) & (!g136) & (!sk[16]) & (!g576) & (!g891) & (g893)) + ((g101) & (!g136) & (!sk[16]) & (!g576) & (g891) & (!g893)) + ((g101) & (!g136) & (!sk[16]) & (!g576) & (g891) & (g893)) + ((g101) & (!g136) & (!sk[16]) & (g576) & (!g891) & (!g893)) + ((g101) & (!g136) & (!sk[16]) & (g576) & (!g891) & (g893)) + ((g101) & (!g136) & (!sk[16]) & (g576) & (g891) & (!g893)) + ((g101) & (!g136) & (!sk[16]) & (g576) & (g891) & (g893)) + ((g101) & (!g136) & (sk[16]) & (!g576) & (g891) & (!g893)) + ((g101) & (!g136) & (sk[16]) & (g576) & (g891) & (!g893)) + ((g101) & (g136) & (!sk[16]) & (!g576) & (!g891) & (!g893)) + ((g101) & (g136) & (!sk[16]) & (!g576) & (!g891) & (g893)) + ((g101) & (g136) & (!sk[16]) & (!g576) & (g891) & (!g893)) + ((g101) & (g136) & (!sk[16]) & (!g576) & (g891) & (g893)) + ((g101) & (g136) & (!sk[16]) & (g576) & (!g891) & (!g893)) + ((g101) & (g136) & (!sk[16]) & (g576) & (!g891) & (g893)) + ((g101) & (g136) & (!sk[16]) & (g576) & (g891) & (!g893)) + ((g101) & (g136) & (!sk[16]) & (g576) & (g891) & (g893)) + ((g101) & (g136) & (sk[16]) & (g576) & (g891) & (!g893)));
	assign g895 = (((!sk[17]) & (g7) & (!g119)) + ((!sk[17]) & (g7) & (g119)) + ((sk[17]) & (g7) & (g119)));
	assign g896 = (((!i_11_) & (!i_9_) & (i_10_) & (!sk[18]) & (g875)) + ((!i_11_) & (!i_9_) & (i_10_) & (sk[18]) & (g875)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[18]) & (!g875)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[18]) & (g875)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[18]) & (!g875)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[18]) & (g875)) + ((i_11_) & (!i_9_) & (!i_10_) & (sk[18]) & (g875)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[18]) & (!g875)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[18]) & (g875)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[18]) & (!g875)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[18]) & (g875)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[18]) & (!g875)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[18]) & (g875)));
	assign g897 = (((!i_5_) & (!g141) & (!g326) & (!sk[19]) & (!g660) & (g896)) + ((!i_5_) & (!g141) & (!g326) & (!sk[19]) & (g660) & (g896)) + ((!i_5_) & (!g141) & (!g326) & (sk[19]) & (g660) & (g896)) + ((!i_5_) & (!g141) & (g326) & (!sk[19]) & (!g660) & (g896)) + ((!i_5_) & (!g141) & (g326) & (!sk[19]) & (g660) & (g896)) + ((!i_5_) & (!g141) & (g326) & (sk[19]) & (g660) & (g896)) + ((!i_5_) & (g141) & (!g326) & (!sk[19]) & (!g660) & (g896)) + ((!i_5_) & (g141) & (!g326) & (!sk[19]) & (g660) & (g896)) + ((!i_5_) & (g141) & (!g326) & (sk[19]) & (g660) & (g896)) + ((!i_5_) & (g141) & (g326) & (!sk[19]) & (!g660) & (g896)) + ((!i_5_) & (g141) & (g326) & (!sk[19]) & (g660) & (g896)) + ((!i_5_) & (g141) & (g326) & (sk[19]) & (g660) & (!g896)) + ((!i_5_) & (g141) & (g326) & (sk[19]) & (g660) & (g896)) + ((i_5_) & (!g141) & (!g326) & (!sk[19]) & (!g660) & (!g896)) + ((i_5_) & (!g141) & (!g326) & (!sk[19]) & (!g660) & (g896)) + ((i_5_) & (!g141) & (!g326) & (!sk[19]) & (g660) & (!g896)) + ((i_5_) & (!g141) & (!g326) & (!sk[19]) & (g660) & (g896)) + ((i_5_) & (!g141) & (!g326) & (sk[19]) & (g660) & (g896)) + ((i_5_) & (!g141) & (g326) & (!sk[19]) & (!g660) & (!g896)) + ((i_5_) & (!g141) & (g326) & (!sk[19]) & (!g660) & (g896)) + ((i_5_) & (!g141) & (g326) & (!sk[19]) & (g660) & (!g896)) + ((i_5_) & (!g141) & (g326) & (!sk[19]) & (g660) & (g896)) + ((i_5_) & (!g141) & (g326) & (sk[19]) & (g660) & (g896)) + ((i_5_) & (g141) & (!g326) & (!sk[19]) & (!g660) & (!g896)) + ((i_5_) & (g141) & (!g326) & (!sk[19]) & (!g660) & (g896)) + ((i_5_) & (g141) & (!g326) & (!sk[19]) & (g660) & (!g896)) + ((i_5_) & (g141) & (!g326) & (!sk[19]) & (g660) & (g896)) + ((i_5_) & (g141) & (!g326) & (sk[19]) & (g660) & (g896)) + ((i_5_) & (g141) & (g326) & (!sk[19]) & (!g660) & (!g896)) + ((i_5_) & (g141) & (g326) & (!sk[19]) & (!g660) & (g896)) + ((i_5_) & (g141) & (g326) & (!sk[19]) & (g660) & (!g896)) + ((i_5_) & (g141) & (g326) & (!sk[19]) & (g660) & (g896)) + ((i_5_) & (g141) & (g326) & (sk[19]) & (g660) & (g896)));
	assign g898 = (((!sk[20]) & (g15) & (!g711)) + ((!sk[20]) & (g15) & (g711)) + ((sk[20]) & (!g15) & (g711)));
	assign g899 = (((!g19) & (sk[21]) & (!g898)) + ((g19) & (!sk[21]) & (!g898)) + ((g19) & (!sk[21]) & (g898)));
	assign g900 = (((!sk[22]) & (i_8_) & (!g100) & (!g899)) + ((!sk[22]) & (i_8_) & (!g100) & (g899)) + ((!sk[22]) & (i_8_) & (g100) & (!g899)) + ((!sk[22]) & (i_8_) & (g100) & (g899)) + ((sk[22]) & (i_8_) & (g100) & (!g899)));
	assign g901 = (((i_8_) & (!g181) & (g135) & (!g548) & (!g671) & (g895)) + ((i_8_) & (!g181) & (g135) & (!g548) & (g671) & (!g895)) + ((i_8_) & (!g181) & (g135) & (!g548) & (g671) & (g895)) + ((i_8_) & (!g181) & (g135) & (g548) & (!g671) & (!g895)) + ((i_8_) & (!g181) & (g135) & (g548) & (!g671) & (g895)) + ((i_8_) & (!g181) & (g135) & (g548) & (g671) & (!g895)) + ((i_8_) & (!g181) & (g135) & (g548) & (g671) & (g895)) + ((i_8_) & (g181) & (g135) & (!g548) & (!g671) & (!g895)) + ((i_8_) & (g181) & (g135) & (!g548) & (!g671) & (g895)) + ((i_8_) & (g181) & (g135) & (!g548) & (g671) & (!g895)) + ((i_8_) & (g181) & (g135) & (!g548) & (g671) & (g895)) + ((i_8_) & (g181) & (g135) & (g548) & (!g671) & (!g895)) + ((i_8_) & (g181) & (g135) & (g548) & (!g671) & (g895)) + ((i_8_) & (g181) & (g135) & (g548) & (g671) & (!g895)) + ((i_8_) & (g181) & (g135) & (g548) & (g671) & (g895)));
	assign g902 = (((!g151) & (!g895) & (!sk[24]) & (!g897) & (!g900) & (g901)) + ((!g151) & (!g895) & (!sk[24]) & (!g897) & (g900) & (g901)) + ((!g151) & (!g895) & (!sk[24]) & (g897) & (!g900) & (g901)) + ((!g151) & (!g895) & (!sk[24]) & (g897) & (g900) & (g901)) + ((!g151) & (!g895) & (sk[24]) & (!g897) & (!g900) & (!g901)) + ((!g151) & (g895) & (!sk[24]) & (!g897) & (!g900) & (g901)) + ((!g151) & (g895) & (!sk[24]) & (!g897) & (g900) & (g901)) + ((!g151) & (g895) & (!sk[24]) & (g897) & (!g900) & (g901)) + ((!g151) & (g895) & (!sk[24]) & (g897) & (g900) & (g901)) + ((!g151) & (g895) & (sk[24]) & (!g897) & (!g900) & (!g901)) + ((g151) & (!g895) & (!sk[24]) & (!g897) & (!g900) & (!g901)) + ((g151) & (!g895) & (!sk[24]) & (!g897) & (!g900) & (g901)) + ((g151) & (!g895) & (!sk[24]) & (!g897) & (g900) & (!g901)) + ((g151) & (!g895) & (!sk[24]) & (!g897) & (g900) & (g901)) + ((g151) & (!g895) & (!sk[24]) & (g897) & (!g900) & (!g901)) + ((g151) & (!g895) & (!sk[24]) & (g897) & (!g900) & (g901)) + ((g151) & (!g895) & (!sk[24]) & (g897) & (g900) & (!g901)) + ((g151) & (!g895) & (!sk[24]) & (g897) & (g900) & (g901)) + ((g151) & (!g895) & (sk[24]) & (!g897) & (!g900) & (!g901)) + ((g151) & (g895) & (!sk[24]) & (!g897) & (!g900) & (!g901)) + ((g151) & (g895) & (!sk[24]) & (!g897) & (!g900) & (g901)) + ((g151) & (g895) & (!sk[24]) & (!g897) & (g900) & (!g901)) + ((g151) & (g895) & (!sk[24]) & (!g897) & (g900) & (g901)) + ((g151) & (g895) & (!sk[24]) & (g897) & (!g900) & (!g901)) + ((g151) & (g895) & (!sk[24]) & (g897) & (!g900) & (g901)) + ((g151) & (g895) & (!sk[24]) & (g897) & (g900) & (!g901)) + ((g151) & (g895) & (!sk[24]) & (g897) & (g900) & (g901)));
	assign g903 = (((!i_8_) & (!sk[25]) & (!g91) & (!g100) & (!g131) & (g461)) + ((!i_8_) & (!sk[25]) & (!g91) & (!g100) & (g131) & (g461)) + ((!i_8_) & (!sk[25]) & (!g91) & (g100) & (!g131) & (g461)) + ((!i_8_) & (!sk[25]) & (!g91) & (g100) & (g131) & (g461)) + ((!i_8_) & (!sk[25]) & (g91) & (!g100) & (!g131) & (g461)) + ((!i_8_) & (!sk[25]) & (g91) & (!g100) & (g131) & (g461)) + ((!i_8_) & (!sk[25]) & (g91) & (g100) & (!g131) & (g461)) + ((!i_8_) & (!sk[25]) & (g91) & (g100) & (g131) & (g461)) + ((!i_8_) & (sk[25]) & (!g91) & (!g100) & (g131) & (g461)) + ((!i_8_) & (sk[25]) & (!g91) & (g100) & (g131) & (g461)) + ((!i_8_) & (sk[25]) & (g91) & (!g100) & (g131) & (g461)) + ((!i_8_) & (sk[25]) & (g91) & (g100) & (g131) & (g461)) + ((i_8_) & (!sk[25]) & (!g91) & (!g100) & (!g131) & (!g461)) + ((i_8_) & (!sk[25]) & (!g91) & (!g100) & (!g131) & (g461)) + ((i_8_) & (!sk[25]) & (!g91) & (!g100) & (g131) & (!g461)) + ((i_8_) & (!sk[25]) & (!g91) & (!g100) & (g131) & (g461)) + ((i_8_) & (!sk[25]) & (!g91) & (g100) & (!g131) & (!g461)) + ((i_8_) & (!sk[25]) & (!g91) & (g100) & (!g131) & (g461)) + ((i_8_) & (!sk[25]) & (!g91) & (g100) & (g131) & (!g461)) + ((i_8_) & (!sk[25]) & (!g91) & (g100) & (g131) & (g461)) + ((i_8_) & (!sk[25]) & (g91) & (!g100) & (!g131) & (!g461)) + ((i_8_) & (!sk[25]) & (g91) & (!g100) & (!g131) & (g461)) + ((i_8_) & (!sk[25]) & (g91) & (!g100) & (g131) & (!g461)) + ((i_8_) & (!sk[25]) & (g91) & (!g100) & (g131) & (g461)) + ((i_8_) & (!sk[25]) & (g91) & (g100) & (!g131) & (!g461)) + ((i_8_) & (!sk[25]) & (g91) & (g100) & (!g131) & (g461)) + ((i_8_) & (!sk[25]) & (g91) & (g100) & (g131) & (!g461)) + ((i_8_) & (!sk[25]) & (g91) & (g100) & (g131) & (g461)) + ((i_8_) & (sk[25]) & (!g91) & (!g100) & (g131) & (g461)) + ((i_8_) & (sk[25]) & (!g91) & (g100) & (g131) & (!g461)) + ((i_8_) & (sk[25]) & (!g91) & (g100) & (g131) & (g461)) + ((i_8_) & (sk[25]) & (g91) & (!g100) & (g131) & (g461)) + ((i_8_) & (sk[25]) & (g91) & (g100) & (g131) & (g461)));
	assign g904 = (((!g101) & (!g136) & (!g676) & (!g677) & (!g861) & (!g903)) + ((!g101) & (!g136) & (!g676) & (!g677) & (!g861) & (g903)) + ((!g101) & (!g136) & (!g676) & (g677) & (!g861) & (!g903)) + ((!g101) & (!g136) & (!g676) & (g677) & (!g861) & (g903)) + ((!g101) & (!g136) & (g676) & (!g677) & (!g861) & (!g903)) + ((!g101) & (!g136) & (g676) & (!g677) & (!g861) & (g903)) + ((!g101) & (!g136) & (g676) & (g677) & (!g861) & (!g903)) + ((!g101) & (!g136) & (g676) & (g677) & (!g861) & (g903)) + ((!g101) & (g136) & (!g676) & (!g677) & (!g861) & (!g903)) + ((!g101) & (g136) & (!g676) & (!g677) & (!g861) & (g903)) + ((!g101) & (g136) & (g676) & (!g677) & (!g861) & (!g903)) + ((!g101) & (g136) & (g676) & (!g677) & (!g861) & (g903)) + ((g101) & (!g136) & (!g676) & (!g677) & (!g861) & (!g903)) + ((g101) & (!g136) & (!g676) & (g677) & (!g861) & (!g903)) + ((g101) & (g136) & (!g676) & (!g677) & (!g861) & (!g903)));
	assign g905 = (((!g7) & (!g102) & (!g131) & (!sk[27]) & (!g146) & (g646)) + ((!g7) & (!g102) & (!g131) & (!sk[27]) & (g146) & (g646)) + ((!g7) & (!g102) & (g131) & (!sk[27]) & (!g146) & (g646)) + ((!g7) & (!g102) & (g131) & (!sk[27]) & (g146) & (g646)) + ((!g7) & (g102) & (!g131) & (!sk[27]) & (!g146) & (g646)) + ((!g7) & (g102) & (!g131) & (!sk[27]) & (g146) & (g646)) + ((!g7) & (g102) & (g131) & (!sk[27]) & (!g146) & (g646)) + ((!g7) & (g102) & (g131) & (!sk[27]) & (g146) & (g646)) + ((g7) & (!g102) & (!g131) & (!sk[27]) & (!g146) & (!g646)) + ((g7) & (!g102) & (!g131) & (!sk[27]) & (!g146) & (g646)) + ((g7) & (!g102) & (!g131) & (!sk[27]) & (g146) & (!g646)) + ((g7) & (!g102) & (!g131) & (!sk[27]) & (g146) & (g646)) + ((g7) & (!g102) & (!g131) & (sk[27]) & (!g146) & (!g646)) + ((g7) & (!g102) & (!g131) & (sk[27]) & (!g146) & (g646)) + ((g7) & (!g102) & (g131) & (!sk[27]) & (!g146) & (!g646)) + ((g7) & (!g102) & (g131) & (!sk[27]) & (!g146) & (g646)) + ((g7) & (!g102) & (g131) & (!sk[27]) & (g146) & (!g646)) + ((g7) & (!g102) & (g131) & (!sk[27]) & (g146) & (g646)) + ((g7) & (!g102) & (g131) & (sk[27]) & (!g146) & (!g646)) + ((g7) & (!g102) & (g131) & (sk[27]) & (!g146) & (g646)) + ((g7) & (!g102) & (g131) & (sk[27]) & (g146) & (!g646)) + ((g7) & (g102) & (!g131) & (!sk[27]) & (!g146) & (!g646)) + ((g7) & (g102) & (!g131) & (!sk[27]) & (!g146) & (g646)) + ((g7) & (g102) & (!g131) & (!sk[27]) & (g146) & (!g646)) + ((g7) & (g102) & (!g131) & (!sk[27]) & (g146) & (g646)) + ((g7) & (g102) & (g131) & (!sk[27]) & (!g146) & (!g646)) + ((g7) & (g102) & (g131) & (!sk[27]) & (!g146) & (g646)) + ((g7) & (g102) & (g131) & (!sk[27]) & (g146) & (!g646)) + ((g7) & (g102) & (g131) & (!sk[27]) & (g146) & (g646)) + ((g7) & (g102) & (g131) & (sk[27]) & (!g146) & (!g646)) + ((g7) & (g102) & (g131) & (sk[27]) & (g146) & (!g646)));
	assign g906 = (((!sk[28]) & (!g7) & (!i_8_) & (!g95) & (!g100) & (g131)) + ((!sk[28]) & (!g7) & (!i_8_) & (!g95) & (g100) & (g131)) + ((!sk[28]) & (!g7) & (!i_8_) & (g95) & (!g100) & (g131)) + ((!sk[28]) & (!g7) & (!i_8_) & (g95) & (g100) & (g131)) + ((!sk[28]) & (!g7) & (i_8_) & (!g95) & (!g100) & (g131)) + ((!sk[28]) & (!g7) & (i_8_) & (!g95) & (g100) & (g131)) + ((!sk[28]) & (!g7) & (i_8_) & (g95) & (!g100) & (g131)) + ((!sk[28]) & (!g7) & (i_8_) & (g95) & (g100) & (g131)) + ((!sk[28]) & (g7) & (!i_8_) & (!g95) & (!g100) & (!g131)) + ((!sk[28]) & (g7) & (!i_8_) & (!g95) & (!g100) & (g131)) + ((!sk[28]) & (g7) & (!i_8_) & (!g95) & (g100) & (!g131)) + ((!sk[28]) & (g7) & (!i_8_) & (!g95) & (g100) & (g131)) + ((!sk[28]) & (g7) & (!i_8_) & (g95) & (!g100) & (!g131)) + ((!sk[28]) & (g7) & (!i_8_) & (g95) & (!g100) & (g131)) + ((!sk[28]) & (g7) & (!i_8_) & (g95) & (g100) & (!g131)) + ((!sk[28]) & (g7) & (!i_8_) & (g95) & (g100) & (g131)) + ((!sk[28]) & (g7) & (i_8_) & (!g95) & (!g100) & (!g131)) + ((!sk[28]) & (g7) & (i_8_) & (!g95) & (!g100) & (g131)) + ((!sk[28]) & (g7) & (i_8_) & (!g95) & (g100) & (!g131)) + ((!sk[28]) & (g7) & (i_8_) & (!g95) & (g100) & (g131)) + ((!sk[28]) & (g7) & (i_8_) & (g95) & (!g100) & (!g131)) + ((!sk[28]) & (g7) & (i_8_) & (g95) & (!g100) & (g131)) + ((!sk[28]) & (g7) & (i_8_) & (g95) & (g100) & (!g131)) + ((!sk[28]) & (g7) & (i_8_) & (g95) & (g100) & (g131)) + ((sk[28]) & (g7) & (i_8_) & (!g95) & (g100) & (g131)) + ((sk[28]) & (g7) & (i_8_) & (g95) & (g100) & (!g131)) + ((sk[28]) & (g7) & (i_8_) & (g95) & (g100) & (g131)));
	assign g907 = (((!sk[29]) & (g7) & (!g102)) + ((!sk[29]) & (g7) & (g102)) + ((sk[29]) & (g7) & (!g102)));
	assign g908 = (((!sk[30]) & (g7) & (!g11)) + ((!sk[30]) & (g7) & (g11)) + ((sk[30]) & (g7) & (g11)));
	assign g909 = (((!i_8_) & (!sk[31]) & (!g100) & (g907) & (g908)) + ((!i_8_) & (!sk[31]) & (g100) & (!g907) & (!g908)) + ((!i_8_) & (!sk[31]) & (g100) & (!g907) & (g908)) + ((!i_8_) & (!sk[31]) & (g100) & (g907) & (!g908)) + ((!i_8_) & (!sk[31]) & (g100) & (g907) & (g908)) + ((i_8_) & (!sk[31]) & (!g100) & (g907) & (!g908)) + ((i_8_) & (!sk[31]) & (!g100) & (g907) & (g908)) + ((i_8_) & (!sk[31]) & (g100) & (!g907) & (!g908)) + ((i_8_) & (!sk[31]) & (g100) & (!g907) & (g908)) + ((i_8_) & (!sk[31]) & (g100) & (g907) & (!g908)) + ((i_8_) & (!sk[31]) & (g100) & (g907) & (g908)) + ((i_8_) & (sk[31]) & (g100) & (!g907) & (g908)) + ((i_8_) & (sk[31]) & (g100) & (g907) & (!g908)) + ((i_8_) & (sk[31]) & (g100) & (g907) & (g908)));
	assign g910 = (((!i_8_) & (!g135) & (!sk[32]) & (g907) & (g908)) + ((!i_8_) & (g135) & (!sk[32]) & (!g907) & (!g908)) + ((!i_8_) & (g135) & (!sk[32]) & (!g907) & (g908)) + ((!i_8_) & (g135) & (!sk[32]) & (g907) & (!g908)) + ((!i_8_) & (g135) & (!sk[32]) & (g907) & (g908)) + ((i_8_) & (!g135) & (!sk[32]) & (g907) & (!g908)) + ((i_8_) & (!g135) & (!sk[32]) & (g907) & (g908)) + ((i_8_) & (g135) & (!sk[32]) & (!g907) & (!g908)) + ((i_8_) & (g135) & (!sk[32]) & (!g907) & (g908)) + ((i_8_) & (g135) & (!sk[32]) & (g907) & (!g908)) + ((i_8_) & (g135) & (!sk[32]) & (g907) & (g908)) + ((i_8_) & (g135) & (sk[32]) & (!g907) & (g908)) + ((i_8_) & (g135) & (sk[32]) & (g907) & (!g908)) + ((i_8_) & (g135) & (sk[32]) & (g907) & (g908)));
	assign g911 = (((!sk[33]) & (!g112) & (!g895) & (g908) & (g881)) + ((!sk[33]) & (!g112) & (g895) & (!g908) & (!g881)) + ((!sk[33]) & (!g112) & (g895) & (!g908) & (g881)) + ((!sk[33]) & (!g112) & (g895) & (g908) & (!g881)) + ((!sk[33]) & (!g112) & (g895) & (g908) & (g881)) + ((!sk[33]) & (g112) & (!g895) & (g908) & (!g881)) + ((!sk[33]) & (g112) & (!g895) & (g908) & (g881)) + ((!sk[33]) & (g112) & (g895) & (!g908) & (!g881)) + ((!sk[33]) & (g112) & (g895) & (!g908) & (g881)) + ((!sk[33]) & (g112) & (g895) & (g908) & (!g881)) + ((!sk[33]) & (g112) & (g895) & (g908) & (g881)) + ((sk[33]) & (g112) & (!g895) & (!g908) & (g881)) + ((sk[33]) & (g112) & (!g895) & (g908) & (!g881)) + ((sk[33]) & (g112) & (!g895) & (g908) & (g881)) + ((sk[33]) & (g112) & (g895) & (!g908) & (!g881)) + ((sk[33]) & (g112) & (g895) & (!g908) & (g881)) + ((sk[33]) & (g112) & (g895) & (g908) & (!g881)) + ((sk[33]) & (g112) & (g895) & (g908) & (g881)));
	assign g912 = (((i_8_) & (!g264) & (g108) & (!g895) & (!g907) & (g881)) + ((i_8_) & (!g264) & (g108) & (!g895) & (g907) & (!g881)) + ((i_8_) & (!g264) & (g108) & (!g895) & (g907) & (g881)) + ((i_8_) & (!g264) & (g108) & (g895) & (!g907) & (!g881)) + ((i_8_) & (!g264) & (g108) & (g895) & (!g907) & (g881)) + ((i_8_) & (!g264) & (g108) & (g895) & (g907) & (!g881)) + ((i_8_) & (!g264) & (g108) & (g895) & (g907) & (g881)) + ((i_8_) & (g264) & (g108) & (!g895) & (!g907) & (!g881)) + ((i_8_) & (g264) & (g108) & (!g895) & (!g907) & (g881)) + ((i_8_) & (g264) & (g108) & (!g895) & (g907) & (!g881)) + ((i_8_) & (g264) & (g108) & (!g895) & (g907) & (g881)) + ((i_8_) & (g264) & (g108) & (g895) & (!g907) & (!g881)) + ((i_8_) & (g264) & (g108) & (g895) & (!g907) & (g881)) + ((i_8_) & (g264) & (g108) & (g895) & (g907) & (!g881)) + ((i_8_) & (g264) & (g108) & (g895) & (g907) & (g881)));
	assign g913 = (((!g906) & (!g909) & (!g910) & (!sk[35]) & (!g911) & (g912)) + ((!g906) & (!g909) & (!g910) & (!sk[35]) & (g911) & (g912)) + ((!g906) & (!g909) & (!g910) & (sk[35]) & (!g911) & (!g912)) + ((!g906) & (!g909) & (g910) & (!sk[35]) & (!g911) & (g912)) + ((!g906) & (!g909) & (g910) & (!sk[35]) & (g911) & (g912)) + ((!g906) & (g909) & (!g910) & (!sk[35]) & (!g911) & (g912)) + ((!g906) & (g909) & (!g910) & (!sk[35]) & (g911) & (g912)) + ((!g906) & (g909) & (g910) & (!sk[35]) & (!g911) & (g912)) + ((!g906) & (g909) & (g910) & (!sk[35]) & (g911) & (g912)) + ((g906) & (!g909) & (!g910) & (!sk[35]) & (!g911) & (!g912)) + ((g906) & (!g909) & (!g910) & (!sk[35]) & (!g911) & (g912)) + ((g906) & (!g909) & (!g910) & (!sk[35]) & (g911) & (!g912)) + ((g906) & (!g909) & (!g910) & (!sk[35]) & (g911) & (g912)) + ((g906) & (!g909) & (g910) & (!sk[35]) & (!g911) & (!g912)) + ((g906) & (!g909) & (g910) & (!sk[35]) & (!g911) & (g912)) + ((g906) & (!g909) & (g910) & (!sk[35]) & (g911) & (!g912)) + ((g906) & (!g909) & (g910) & (!sk[35]) & (g911) & (g912)) + ((g906) & (g909) & (!g910) & (!sk[35]) & (!g911) & (!g912)) + ((g906) & (g909) & (!g910) & (!sk[35]) & (!g911) & (g912)) + ((g906) & (g909) & (!g910) & (!sk[35]) & (g911) & (!g912)) + ((g906) & (g909) & (!g910) & (!sk[35]) & (g911) & (g912)) + ((g906) & (g909) & (g910) & (!sk[35]) & (!g911) & (!g912)) + ((g906) & (g909) & (g910) & (!sk[35]) & (!g911) & (g912)) + ((g906) & (g909) & (g910) & (!sk[35]) & (g911) & (!g912)) + ((g906) & (g909) & (g910) & (!sk[35]) & (g911) & (g912)));
	assign g914 = (((!sk[36]) & (g102) & (!g711) & (!g675)) + ((!sk[36]) & (g102) & (!g711) & (g675)) + ((!sk[36]) & (g102) & (g711) & (!g675)) + ((!sk[36]) & (g102) & (g711) & (g675)) + ((sk[36]) & (!g102) & (!g711) & (!g675)) + ((sk[36]) & (g102) & (!g711) & (!g675)) + ((sk[36]) & (g102) & (g711) & (!g675)));
	assign g915 = (((!i_8_) & (!g100) & (!g112) & (!g887) & (!sk[37]) & (g914)) + ((!i_8_) & (!g100) & (!g112) & (g887) & (!sk[37]) & (g914)) + ((!i_8_) & (!g100) & (g112) & (!g887) & (!sk[37]) & (g914)) + ((!i_8_) & (!g100) & (g112) & (!g887) & (sk[37]) & (!g914)) + ((!i_8_) & (!g100) & (g112) & (!g887) & (sk[37]) & (g914)) + ((!i_8_) & (!g100) & (g112) & (g887) & (!sk[37]) & (g914)) + ((!i_8_) & (g100) & (!g112) & (!g887) & (!sk[37]) & (g914)) + ((!i_8_) & (g100) & (!g112) & (g887) & (!sk[37]) & (g914)) + ((!i_8_) & (g100) & (g112) & (!g887) & (!sk[37]) & (g914)) + ((!i_8_) & (g100) & (g112) & (!g887) & (sk[37]) & (!g914)) + ((!i_8_) & (g100) & (g112) & (!g887) & (sk[37]) & (g914)) + ((!i_8_) & (g100) & (g112) & (g887) & (!sk[37]) & (g914)) + ((i_8_) & (!g100) & (!g112) & (!g887) & (!sk[37]) & (!g914)) + ((i_8_) & (!g100) & (!g112) & (!g887) & (!sk[37]) & (g914)) + ((i_8_) & (!g100) & (!g112) & (g887) & (!sk[37]) & (!g914)) + ((i_8_) & (!g100) & (!g112) & (g887) & (!sk[37]) & (g914)) + ((i_8_) & (!g100) & (g112) & (!g887) & (!sk[37]) & (!g914)) + ((i_8_) & (!g100) & (g112) & (!g887) & (!sk[37]) & (g914)) + ((i_8_) & (!g100) & (g112) & (!g887) & (sk[37]) & (!g914)) + ((i_8_) & (!g100) & (g112) & (!g887) & (sk[37]) & (g914)) + ((i_8_) & (!g100) & (g112) & (g887) & (!sk[37]) & (!g914)) + ((i_8_) & (!g100) & (g112) & (g887) & (!sk[37]) & (g914)) + ((i_8_) & (g100) & (!g112) & (!g887) & (!sk[37]) & (!g914)) + ((i_8_) & (g100) & (!g112) & (!g887) & (!sk[37]) & (g914)) + ((i_8_) & (g100) & (!g112) & (!g887) & (sk[37]) & (!g914)) + ((i_8_) & (g100) & (!g112) & (!g887) & (sk[37]) & (g914)) + ((i_8_) & (g100) & (!g112) & (g887) & (!sk[37]) & (!g914)) + ((i_8_) & (g100) & (!g112) & (g887) & (!sk[37]) & (g914)) + ((i_8_) & (g100) & (!g112) & (g887) & (sk[37]) & (!g914)) + ((i_8_) & (g100) & (g112) & (!g887) & (!sk[37]) & (!g914)) + ((i_8_) & (g100) & (g112) & (!g887) & (!sk[37]) & (g914)) + ((i_8_) & (g100) & (g112) & (!g887) & (sk[37]) & (!g914)) + ((i_8_) & (g100) & (g112) & (!g887) & (sk[37]) & (g914)) + ((i_8_) & (g100) & (g112) & (g887) & (!sk[37]) & (!g914)) + ((i_8_) & (g100) & (g112) & (g887) & (!sk[37]) & (g914)) + ((i_8_) & (g100) & (g112) & (g887) & (sk[37]) & (!g914)));
	assign g916 = (((!sk[38]) & (!g323) & (!g914) & (!g908) & (!g899) & (g915)) + ((!sk[38]) & (!g323) & (!g914) & (!g908) & (g899) & (g915)) + ((!sk[38]) & (!g323) & (!g914) & (g908) & (!g899) & (g915)) + ((!sk[38]) & (!g323) & (!g914) & (g908) & (g899) & (g915)) + ((!sk[38]) & (!g323) & (g914) & (!g908) & (!g899) & (g915)) + ((!sk[38]) & (!g323) & (g914) & (!g908) & (g899) & (g915)) + ((!sk[38]) & (!g323) & (g914) & (g908) & (!g899) & (g915)) + ((!sk[38]) & (!g323) & (g914) & (g908) & (g899) & (g915)) + ((!sk[38]) & (g323) & (!g914) & (!g908) & (!g899) & (!g915)) + ((!sk[38]) & (g323) & (!g914) & (!g908) & (!g899) & (g915)) + ((!sk[38]) & (g323) & (!g914) & (!g908) & (g899) & (!g915)) + ((!sk[38]) & (g323) & (!g914) & (!g908) & (g899) & (g915)) + ((!sk[38]) & (g323) & (!g914) & (g908) & (!g899) & (!g915)) + ((!sk[38]) & (g323) & (!g914) & (g908) & (!g899) & (g915)) + ((!sk[38]) & (g323) & (!g914) & (g908) & (g899) & (!g915)) + ((!sk[38]) & (g323) & (!g914) & (g908) & (g899) & (g915)) + ((!sk[38]) & (g323) & (g914) & (!g908) & (!g899) & (!g915)) + ((!sk[38]) & (g323) & (g914) & (!g908) & (!g899) & (g915)) + ((!sk[38]) & (g323) & (g914) & (!g908) & (g899) & (!g915)) + ((!sk[38]) & (g323) & (g914) & (!g908) & (g899) & (g915)) + ((!sk[38]) & (g323) & (g914) & (g908) & (!g899) & (!g915)) + ((!sk[38]) & (g323) & (g914) & (g908) & (!g899) & (g915)) + ((!sk[38]) & (g323) & (g914) & (g908) & (g899) & (!g915)) + ((!sk[38]) & (g323) & (g914) & (g908) & (g899) & (g915)) + ((sk[38]) & (!g323) & (!g914) & (!g908) & (!g899) & (!g915)) + ((sk[38]) & (!g323) & (!g914) & (!g908) & (g899) & (!g915)) + ((sk[38]) & (!g323) & (!g914) & (g908) & (!g899) & (!g915)) + ((sk[38]) & (!g323) & (!g914) & (g908) & (g899) & (!g915)) + ((sk[38]) & (!g323) & (g914) & (!g908) & (!g899) & (!g915)) + ((sk[38]) & (!g323) & (g914) & (!g908) & (g899) & (!g915)) + ((sk[38]) & (!g323) & (g914) & (g908) & (!g899) & (!g915)) + ((sk[38]) & (!g323) & (g914) & (g908) & (g899) & (!g915)) + ((sk[38]) & (g323) & (g914) & (!g908) & (g899) & (!g915)));
	assign g917 = (((g894) & (g902) & (g904) & (!g905) & (g913) & (g916)));
	assign g918 = (((!g880) & (!g694) & (!sk[40]) & (g890) & (g917)) + ((!g880) & (g694) & (!sk[40]) & (!g890) & (!g917)) + ((!g880) & (g694) & (!sk[40]) & (!g890) & (g917)) + ((!g880) & (g694) & (!sk[40]) & (g890) & (!g917)) + ((!g880) & (g694) & (!sk[40]) & (g890) & (g917)) + ((g880) & (!g694) & (!sk[40]) & (g890) & (!g917)) + ((g880) & (!g694) & (!sk[40]) & (g890) & (g917)) + ((g880) & (g694) & (!sk[40]) & (!g890) & (!g917)) + ((g880) & (g694) & (!sk[40]) & (!g890) & (g917)) + ((g880) & (g694) & (!sk[40]) & (g890) & (!g917)) + ((g880) & (g694) & (!sk[40]) & (g890) & (g917)) + ((g880) & (g694) & (sk[40]) & (g890) & (g917)));
	assign g919 = (((!g316) & (!g216) & (!g207) & (sk[41]) & (!g895)) + ((!g316) & (!g216) & (g207) & (!sk[41]) & (g895)) + ((!g316) & (g216) & (!g207) & (!sk[41]) & (!g895)) + ((!g316) & (g216) & (!g207) & (!sk[41]) & (g895)) + ((!g316) & (g216) & (g207) & (!sk[41]) & (!g895)) + ((!g316) & (g216) & (g207) & (!sk[41]) & (g895)) + ((g316) & (!g216) & (g207) & (!sk[41]) & (!g895)) + ((g316) & (!g216) & (g207) & (!sk[41]) & (g895)) + ((g316) & (g216) & (!g207) & (!sk[41]) & (!g895)) + ((g316) & (g216) & (!g207) & (!sk[41]) & (g895)) + ((g316) & (g216) & (g207) & (!sk[41]) & (!g895)) + ((g316) & (g216) & (g207) & (!sk[41]) & (g895)));
	assign g920 = (((!sk[42]) & (!g547) & (!g532) & (g676) & (g896)) + ((!sk[42]) & (!g547) & (g532) & (!g676) & (!g896)) + ((!sk[42]) & (!g547) & (g532) & (!g676) & (g896)) + ((!sk[42]) & (!g547) & (g532) & (g676) & (!g896)) + ((!sk[42]) & (!g547) & (g532) & (g676) & (g896)) + ((!sk[42]) & (g547) & (!g532) & (g676) & (!g896)) + ((!sk[42]) & (g547) & (!g532) & (g676) & (g896)) + ((!sk[42]) & (g547) & (g532) & (!g676) & (!g896)) + ((!sk[42]) & (g547) & (g532) & (!g676) & (g896)) + ((!sk[42]) & (g547) & (g532) & (g676) & (!g896)) + ((!sk[42]) & (g547) & (g532) & (g676) & (g896)) + ((sk[42]) & (g547) & (!g532) & (!g676) & (!g896)));
	assign g921 = (((g185) & (!sk[43]) & (!g551) & (!g734)) + ((g185) & (!sk[43]) & (!g551) & (g734)) + ((g185) & (!sk[43]) & (g551) & (!g734)) + ((g185) & (!sk[43]) & (g551) & (g734)) + ((g185) & (sk[43]) & (!g551) & (!g734)));
	assign g922 = (((!sk[44]) & (g134) & (!g881) & (!g921)) + ((!sk[44]) & (g134) & (!g881) & (g921)) + ((!sk[44]) & (g134) & (g881) & (!g921)) + ((!sk[44]) & (g134) & (g881) & (g921)) + ((sk[44]) & (g134) & (!g881) & (!g921)) + ((sk[44]) & (g134) & (g881) & (!g921)) + ((sk[44]) & (g134) & (g881) & (g921)));
	assign g923 = (((!g251) & (!sk[45]) & (!g919) & (g920) & (g922)) + ((!g251) & (!sk[45]) & (g919) & (!g920) & (!g922)) + ((!g251) & (!sk[45]) & (g919) & (!g920) & (g922)) + ((!g251) & (!sk[45]) & (g919) & (g920) & (!g922)) + ((!g251) & (!sk[45]) & (g919) & (g920) & (g922)) + ((!g251) & (sk[45]) & (!g919) & (!g920) & (!g922)) + ((!g251) & (sk[45]) & (!g919) & (g920) & (!g922)) + ((!g251) & (sk[45]) & (g919) & (!g920) & (!g922)) + ((!g251) & (sk[45]) & (g919) & (g920) & (!g922)) + ((g251) & (!sk[45]) & (!g919) & (g920) & (!g922)) + ((g251) & (!sk[45]) & (!g919) & (g920) & (g922)) + ((g251) & (!sk[45]) & (g919) & (!g920) & (!g922)) + ((g251) & (!sk[45]) & (g919) & (!g920) & (g922)) + ((g251) & (!sk[45]) & (g919) & (g920) & (!g922)) + ((g251) & (!sk[45]) & (g919) & (g920) & (g922)) + ((g251) & (sk[45]) & (g919) & (g920) & (!g922)));
	assign g924 = (((!g19) & (!g15) & (!g91) & (!g99) & (!sk[46]) & (g461)) + ((!g19) & (!g15) & (!g91) & (g99) & (!sk[46]) & (g461)) + ((!g19) & (!g15) & (!g91) & (g99) & (sk[46]) & (!g461)) + ((!g19) & (!g15) & (!g91) & (g99) & (sk[46]) & (g461)) + ((!g19) & (!g15) & (g91) & (!g99) & (!sk[46]) & (g461)) + ((!g19) & (!g15) & (g91) & (g99) & (!sk[46]) & (g461)) + ((!g19) & (!g15) & (g91) & (g99) & (sk[46]) & (g461)) + ((!g19) & (g15) & (!g91) & (!g99) & (!sk[46]) & (g461)) + ((!g19) & (g15) & (!g91) & (g99) & (!sk[46]) & (g461)) + ((!g19) & (g15) & (g91) & (!g99) & (!sk[46]) & (g461)) + ((!g19) & (g15) & (g91) & (g99) & (!sk[46]) & (g461)) + ((g19) & (!g15) & (!g91) & (!g99) & (!sk[46]) & (!g461)) + ((g19) & (!g15) & (!g91) & (!g99) & (!sk[46]) & (g461)) + ((g19) & (!g15) & (!g91) & (g99) & (!sk[46]) & (!g461)) + ((g19) & (!g15) & (!g91) & (g99) & (!sk[46]) & (g461)) + ((g19) & (!g15) & (!g91) & (g99) & (sk[46]) & (!g461)) + ((g19) & (!g15) & (!g91) & (g99) & (sk[46]) & (g461)) + ((g19) & (!g15) & (g91) & (!g99) & (!sk[46]) & (!g461)) + ((g19) & (!g15) & (g91) & (!g99) & (!sk[46]) & (g461)) + ((g19) & (!g15) & (g91) & (g99) & (!sk[46]) & (!g461)) + ((g19) & (!g15) & (g91) & (g99) & (!sk[46]) & (g461)) + ((g19) & (!g15) & (g91) & (g99) & (sk[46]) & (!g461)) + ((g19) & (!g15) & (g91) & (g99) & (sk[46]) & (g461)) + ((g19) & (g15) & (!g91) & (!g99) & (!sk[46]) & (!g461)) + ((g19) & (g15) & (!g91) & (!g99) & (!sk[46]) & (g461)) + ((g19) & (g15) & (!g91) & (g99) & (!sk[46]) & (!g461)) + ((g19) & (g15) & (!g91) & (g99) & (!sk[46]) & (g461)) + ((g19) & (g15) & (!g91) & (g99) & (sk[46]) & (!g461)) + ((g19) & (g15) & (!g91) & (g99) & (sk[46]) & (g461)) + ((g19) & (g15) & (g91) & (!g99) & (!sk[46]) & (!g461)) + ((g19) & (g15) & (g91) & (!g99) & (!sk[46]) & (g461)) + ((g19) & (g15) & (g91) & (g99) & (!sk[46]) & (!g461)) + ((g19) & (g15) & (g91) & (g99) & (!sk[46]) & (g461)) + ((g19) & (g15) & (g91) & (g99) & (sk[46]) & (!g461)) + ((g19) & (g15) & (g91) & (g99) & (sk[46]) & (g461)));
	assign g925 = (((!g316) & (!g669) & (g676) & (!sk[47]) & (g896)) + ((!g316) & (g669) & (!g676) & (!sk[47]) & (!g896)) + ((!g316) & (g669) & (!g676) & (!sk[47]) & (g896)) + ((!g316) & (g669) & (!g676) & (sk[47]) & (!g896)) + ((!g316) & (g669) & (g676) & (!sk[47]) & (!g896)) + ((!g316) & (g669) & (g676) & (!sk[47]) & (g896)) + ((g316) & (!g669) & (g676) & (!sk[47]) & (!g896)) + ((g316) & (!g669) & (g676) & (!sk[47]) & (g896)) + ((g316) & (g669) & (!g676) & (!sk[47]) & (!g896)) + ((g316) & (g669) & (!g676) & (!sk[47]) & (g896)) + ((g316) & (g669) & (g676) & (!sk[47]) & (!g896)) + ((g316) & (g669) & (g676) & (!sk[47]) & (g896)));
	assign g926 = (((!g99) & (!g887) & (!sk[48]) & (g924) & (g925)) + ((!g99) & (!g887) & (sk[48]) & (!g924) & (!g925)) + ((!g99) & (!g887) & (sk[48]) & (!g924) & (g925)) + ((!g99) & (g887) & (!sk[48]) & (!g924) & (!g925)) + ((!g99) & (g887) & (!sk[48]) & (!g924) & (g925)) + ((!g99) & (g887) & (!sk[48]) & (g924) & (!g925)) + ((!g99) & (g887) & (!sk[48]) & (g924) & (g925)) + ((!g99) & (g887) & (sk[48]) & (!g924) & (!g925)) + ((!g99) & (g887) & (sk[48]) & (!g924) & (g925)) + ((g99) & (!g887) & (!sk[48]) & (g924) & (!g925)) + ((g99) & (!g887) & (!sk[48]) & (g924) & (g925)) + ((g99) & (g887) & (!sk[48]) & (!g924) & (!g925)) + ((g99) & (g887) & (!sk[48]) & (!g924) & (g925)) + ((g99) & (g887) & (!sk[48]) & (g924) & (!g925)) + ((g99) & (g887) & (!sk[48]) & (g924) & (g925)) + ((g99) & (g887) & (sk[48]) & (!g924) & (g925)));
	assign g927 = (((!sk[49]) & (!g47) & (!g108) & (g560) & (g926)) + ((!sk[49]) & (!g47) & (g108) & (!g560) & (!g926)) + ((!sk[49]) & (!g47) & (g108) & (!g560) & (g926)) + ((!sk[49]) & (!g47) & (g108) & (g560) & (!g926)) + ((!sk[49]) & (!g47) & (g108) & (g560) & (g926)) + ((!sk[49]) & (g47) & (!g108) & (g560) & (!g926)) + ((!sk[49]) & (g47) & (!g108) & (g560) & (g926)) + ((!sk[49]) & (g47) & (g108) & (!g560) & (!g926)) + ((!sk[49]) & (g47) & (g108) & (!g560) & (g926)) + ((!sk[49]) & (g47) & (g108) & (g560) & (!g926)) + ((!sk[49]) & (g47) & (g108) & (g560) & (g926)) + ((sk[49]) & (!g47) & (!g108) & (!g560) & (g926)) + ((sk[49]) & (!g47) & (!g108) & (g560) & (g926)) + ((sk[49]) & (!g47) & (g108) & (!g560) & (g926)) + ((sk[49]) & (g47) & (!g108) & (!g560) & (g926)) + ((sk[49]) & (g47) & (!g108) & (g560) & (g926)));
	assign g928 = (((!g23) & (!g206) & (!sk[50]) & (g99) & (g561)) + ((!g23) & (!g206) & (sk[50]) & (g99) & (!g561)) + ((!g23) & (!g206) & (sk[50]) & (g99) & (g561)) + ((!g23) & (g206) & (!sk[50]) & (!g99) & (!g561)) + ((!g23) & (g206) & (!sk[50]) & (!g99) & (g561)) + ((!g23) & (g206) & (!sk[50]) & (g99) & (!g561)) + ((!g23) & (g206) & (!sk[50]) & (g99) & (g561)) + ((!g23) & (g206) & (sk[50]) & (g99) & (g561)) + ((g23) & (!g206) & (!sk[50]) & (g99) & (!g561)) + ((g23) & (!g206) & (!sk[50]) & (g99) & (g561)) + ((g23) & (!g206) & (sk[50]) & (g99) & (!g561)) + ((g23) & (!g206) & (sk[50]) & (g99) & (g561)) + ((g23) & (g206) & (!sk[50]) & (!g99) & (!g561)) + ((g23) & (g206) & (!sk[50]) & (!g99) & (g561)) + ((g23) & (g206) & (!sk[50]) & (g99) & (!g561)) + ((g23) & (g206) & (!sk[50]) & (g99) & (g561)) + ((g23) & (g206) & (sk[50]) & (g99) & (!g561)) + ((g23) & (g206) & (sk[50]) & (g99) & (g561)));
	assign g929 = (((!g99) & (!g220) & (g550) & (!sk[51]) & (g675)) + ((!g99) & (g220) & (!g550) & (!sk[51]) & (!g675)) + ((!g99) & (g220) & (!g550) & (!sk[51]) & (g675)) + ((!g99) & (g220) & (g550) & (!sk[51]) & (!g675)) + ((!g99) & (g220) & (g550) & (!sk[51]) & (g675)) + ((g99) & (!g220) & (!g550) & (sk[51]) & (g675)) + ((g99) & (!g220) & (g550) & (!sk[51]) & (!g675)) + ((g99) & (!g220) & (g550) & (!sk[51]) & (g675)) + ((g99) & (!g220) & (g550) & (sk[51]) & (!g675)) + ((g99) & (!g220) & (g550) & (sk[51]) & (g675)) + ((g99) & (g220) & (!g550) & (!sk[51]) & (!g675)) + ((g99) & (g220) & (!g550) & (!sk[51]) & (g675)) + ((g99) & (g220) & (!g550) & (sk[51]) & (!g675)) + ((g99) & (g220) & (!g550) & (sk[51]) & (g675)) + ((g99) & (g220) & (g550) & (!sk[51]) & (!g675)) + ((g99) & (g220) & (g550) & (!sk[51]) & (g675)) + ((g99) & (g220) & (g550) & (sk[51]) & (!g675)) + ((g99) & (g220) & (g550) & (sk[51]) & (g675)));
	assign g930 = (((!g45) & (!g746) & (!sk[52]) & (g928) & (g929)) + ((!g45) & (!g746) & (sk[52]) & (!g928) & (!g929)) + ((!g45) & (g746) & (!sk[52]) & (!g928) & (!g929)) + ((!g45) & (g746) & (!sk[52]) & (!g928) & (g929)) + ((!g45) & (g746) & (!sk[52]) & (g928) & (!g929)) + ((!g45) & (g746) & (!sk[52]) & (g928) & (g929)) + ((!g45) & (g746) & (sk[52]) & (!g928) & (!g929)) + ((g45) & (!g746) & (!sk[52]) & (g928) & (!g929)) + ((g45) & (!g746) & (!sk[52]) & (g928) & (g929)) + ((g45) & (!g746) & (sk[52]) & (!g928) & (!g929)) + ((g45) & (g746) & (!sk[52]) & (!g928) & (!g929)) + ((g45) & (g746) & (!sk[52]) & (!g928) & (g929)) + ((g45) & (g746) & (!sk[52]) & (g928) & (!g929)) + ((g45) & (g746) & (!sk[52]) & (g928) & (g929)));
	assign g931 = (((!sk[53]) & (g99) & (!g185) & (!g882)) + ((!sk[53]) & (g99) & (!g185) & (g882)) + ((!sk[53]) & (g99) & (g185) & (!g882)) + ((!sk[53]) & (g99) & (g185) & (g882)) + ((sk[53]) & (g99) & (!g185) & (!g882)) + ((sk[53]) & (g99) & (!g185) & (g882)) + ((sk[53]) & (g99) & (g185) & (!g882)));
	assign g932 = (((!g8) & (!sk[54]) & (!g10) & (!g99) & (!g221) & (g544)) + ((!g8) & (!sk[54]) & (!g10) & (!g99) & (g221) & (g544)) + ((!g8) & (!sk[54]) & (!g10) & (g99) & (!g221) & (g544)) + ((!g8) & (!sk[54]) & (!g10) & (g99) & (g221) & (g544)) + ((!g8) & (!sk[54]) & (g10) & (!g99) & (!g221) & (g544)) + ((!g8) & (!sk[54]) & (g10) & (!g99) & (g221) & (g544)) + ((!g8) & (!sk[54]) & (g10) & (g99) & (!g221) & (g544)) + ((!g8) & (!sk[54]) & (g10) & (g99) & (g221) & (g544)) + ((!g8) & (sk[54]) & (!g10) & (g99) & (!g221) & (!g544)) + ((!g8) & (sk[54]) & (!g10) & (g99) & (!g221) & (g544)) + ((!g8) & (sk[54]) & (!g10) & (g99) & (g221) & (!g544)) + ((!g8) & (sk[54]) & (!g10) & (g99) & (g221) & (g544)) + ((!g8) & (sk[54]) & (g10) & (g99) & (!g221) & (!g544)) + ((!g8) & (sk[54]) & (g10) & (g99) & (!g221) & (g544)) + ((!g8) & (sk[54]) & (g10) & (g99) & (g221) & (!g544)) + ((!g8) & (sk[54]) & (g10) & (g99) & (g221) & (g544)) + ((g8) & (!sk[54]) & (!g10) & (!g99) & (!g221) & (!g544)) + ((g8) & (!sk[54]) & (!g10) & (!g99) & (!g221) & (g544)) + ((g8) & (!sk[54]) & (!g10) & (!g99) & (g221) & (!g544)) + ((g8) & (!sk[54]) & (!g10) & (!g99) & (g221) & (g544)) + ((g8) & (!sk[54]) & (!g10) & (g99) & (!g221) & (!g544)) + ((g8) & (!sk[54]) & (!g10) & (g99) & (!g221) & (g544)) + ((g8) & (!sk[54]) & (!g10) & (g99) & (g221) & (!g544)) + ((g8) & (!sk[54]) & (!g10) & (g99) & (g221) & (g544)) + ((g8) & (!sk[54]) & (g10) & (!g99) & (!g221) & (!g544)) + ((g8) & (!sk[54]) & (g10) & (!g99) & (!g221) & (g544)) + ((g8) & (!sk[54]) & (g10) & (!g99) & (g221) & (!g544)) + ((g8) & (!sk[54]) & (g10) & (!g99) & (g221) & (g544)) + ((g8) & (!sk[54]) & (g10) & (g99) & (!g221) & (!g544)) + ((g8) & (!sk[54]) & (g10) & (g99) & (!g221) & (g544)) + ((g8) & (!sk[54]) & (g10) & (g99) & (g221) & (!g544)) + ((g8) & (!sk[54]) & (g10) & (g99) & (g221) & (g544)) + ((g8) & (sk[54]) & (!g10) & (g99) & (!g221) & (!g544)) + ((g8) & (sk[54]) & (!g10) & (g99) & (!g221) & (g544)) + ((g8) & (sk[54]) & (!g10) & (g99) & (g221) & (!g544)) + ((g8) & (sk[54]) & (g10) & (g99) & (!g221) & (!g544)) + ((g8) & (sk[54]) & (g10) & (g99) & (!g221) & (g544)) + ((g8) & (sk[54]) & (g10) & (g99) & (g221) & (!g544)) + ((g8) & (sk[54]) & (g10) & (g99) & (g221) & (g544)));
	assign g933 = (((!g264) & (!g101) & (!sk[55]) & (g931) & (g932)) + ((!g264) & (!g101) & (sk[55]) & (!g931) & (!g932)) + ((!g264) & (g101) & (!sk[55]) & (!g931) & (!g932)) + ((!g264) & (g101) & (!sk[55]) & (!g931) & (g932)) + ((!g264) & (g101) & (!sk[55]) & (g931) & (!g932)) + ((!g264) & (g101) & (!sk[55]) & (g931) & (g932)) + ((!g264) & (g101) & (sk[55]) & (!g931) & (!g932)) + ((g264) & (!g101) & (!sk[55]) & (g931) & (!g932)) + ((g264) & (!g101) & (!sk[55]) & (g931) & (g932)) + ((g264) & (!g101) & (sk[55]) & (!g931) & (!g932)) + ((g264) & (g101) & (!sk[55]) & (!g931) & (!g932)) + ((g264) & (g101) & (!sk[55]) & (!g931) & (g932)) + ((g264) & (g101) & (!sk[55]) & (g931) & (!g932)) + ((g264) & (g101) & (!sk[55]) & (g931) & (g932)));
	assign g934 = (((g108) & (!sk[56]) & (!g908)) + ((g108) & (!sk[56]) & (g908)) + ((g108) & (sk[56]) & (g908)));
	assign g935 = (((!g23) & (!g206) & (g423) & (!sk[57]) & (g561)) + ((!g23) & (!g206) & (g423) & (sk[57]) & (!g561)) + ((!g23) & (!g206) & (g423) & (sk[57]) & (g561)) + ((!g23) & (g206) & (!g423) & (!sk[57]) & (!g561)) + ((!g23) & (g206) & (!g423) & (!sk[57]) & (g561)) + ((!g23) & (g206) & (g423) & (!sk[57]) & (!g561)) + ((!g23) & (g206) & (g423) & (!sk[57]) & (g561)) + ((!g23) & (g206) & (g423) & (sk[57]) & (g561)) + ((g23) & (!g206) & (g423) & (!sk[57]) & (!g561)) + ((g23) & (!g206) & (g423) & (!sk[57]) & (g561)) + ((g23) & (!g206) & (g423) & (sk[57]) & (!g561)) + ((g23) & (!g206) & (g423) & (sk[57]) & (g561)) + ((g23) & (g206) & (!g423) & (!sk[57]) & (!g561)) + ((g23) & (g206) & (!g423) & (!sk[57]) & (g561)) + ((g23) & (g206) & (g423) & (!sk[57]) & (!g561)) + ((g23) & (g206) & (g423) & (!sk[57]) & (g561)) + ((g23) & (g206) & (g423) & (sk[57]) & (!g561)) + ((g23) & (g206) & (g423) & (sk[57]) & (g561)));
	assign g936 = (((!i_14_) & (!i_12_) & (!sk[58]) & (!i_13_) & (!g99) & (g131)) + ((!i_14_) & (!i_12_) & (!sk[58]) & (!i_13_) & (g99) & (g131)) + ((!i_14_) & (!i_12_) & (!sk[58]) & (i_13_) & (!g99) & (g131)) + ((!i_14_) & (!i_12_) & (!sk[58]) & (i_13_) & (g99) & (g131)) + ((!i_14_) & (!i_12_) & (sk[58]) & (i_13_) & (g99) & (g131)) + ((!i_14_) & (i_12_) & (!sk[58]) & (!i_13_) & (!g99) & (g131)) + ((!i_14_) & (i_12_) & (!sk[58]) & (!i_13_) & (g99) & (g131)) + ((!i_14_) & (i_12_) & (!sk[58]) & (i_13_) & (!g99) & (g131)) + ((!i_14_) & (i_12_) & (!sk[58]) & (i_13_) & (g99) & (g131)) + ((!i_14_) & (i_12_) & (sk[58]) & (!i_13_) & (g99) & (g131)) + ((!i_14_) & (i_12_) & (sk[58]) & (i_13_) & (g99) & (g131)) + ((i_14_) & (!i_12_) & (!sk[58]) & (!i_13_) & (!g99) & (!g131)) + ((i_14_) & (!i_12_) & (!sk[58]) & (!i_13_) & (!g99) & (g131)) + ((i_14_) & (!i_12_) & (!sk[58]) & (!i_13_) & (g99) & (!g131)) + ((i_14_) & (!i_12_) & (!sk[58]) & (!i_13_) & (g99) & (g131)) + ((i_14_) & (!i_12_) & (!sk[58]) & (i_13_) & (!g99) & (!g131)) + ((i_14_) & (!i_12_) & (!sk[58]) & (i_13_) & (!g99) & (g131)) + ((i_14_) & (!i_12_) & (!sk[58]) & (i_13_) & (g99) & (!g131)) + ((i_14_) & (!i_12_) & (!sk[58]) & (i_13_) & (g99) & (g131)) + ((i_14_) & (i_12_) & (!sk[58]) & (!i_13_) & (!g99) & (!g131)) + ((i_14_) & (i_12_) & (!sk[58]) & (!i_13_) & (!g99) & (g131)) + ((i_14_) & (i_12_) & (!sk[58]) & (!i_13_) & (g99) & (!g131)) + ((i_14_) & (i_12_) & (!sk[58]) & (!i_13_) & (g99) & (g131)) + ((i_14_) & (i_12_) & (!sk[58]) & (i_13_) & (!g99) & (!g131)) + ((i_14_) & (i_12_) & (!sk[58]) & (i_13_) & (!g99) & (g131)) + ((i_14_) & (i_12_) & (!sk[58]) & (i_13_) & (g99) & (!g131)) + ((i_14_) & (i_12_) & (!sk[58]) & (i_13_) & (g99) & (g131)));
	assign g937 = (((!sk[59]) & (!i_14_) & (!i_12_) & (!i_13_) & (!g99) & (g95)) + ((!sk[59]) & (!i_14_) & (!i_12_) & (!i_13_) & (g99) & (g95)) + ((!sk[59]) & (!i_14_) & (!i_12_) & (i_13_) & (!g99) & (g95)) + ((!sk[59]) & (!i_14_) & (!i_12_) & (i_13_) & (g99) & (g95)) + ((!sk[59]) & (!i_14_) & (i_12_) & (!i_13_) & (!g99) & (g95)) + ((!sk[59]) & (!i_14_) & (i_12_) & (!i_13_) & (g99) & (g95)) + ((!sk[59]) & (!i_14_) & (i_12_) & (i_13_) & (!g99) & (g95)) + ((!sk[59]) & (!i_14_) & (i_12_) & (i_13_) & (g99) & (g95)) + ((!sk[59]) & (i_14_) & (!i_12_) & (!i_13_) & (!g99) & (!g95)) + ((!sk[59]) & (i_14_) & (!i_12_) & (!i_13_) & (!g99) & (g95)) + ((!sk[59]) & (i_14_) & (!i_12_) & (!i_13_) & (g99) & (!g95)) + ((!sk[59]) & (i_14_) & (!i_12_) & (!i_13_) & (g99) & (g95)) + ((!sk[59]) & (i_14_) & (!i_12_) & (i_13_) & (!g99) & (!g95)) + ((!sk[59]) & (i_14_) & (!i_12_) & (i_13_) & (!g99) & (g95)) + ((!sk[59]) & (i_14_) & (!i_12_) & (i_13_) & (g99) & (!g95)) + ((!sk[59]) & (i_14_) & (!i_12_) & (i_13_) & (g99) & (g95)) + ((!sk[59]) & (i_14_) & (i_12_) & (!i_13_) & (!g99) & (!g95)) + ((!sk[59]) & (i_14_) & (i_12_) & (!i_13_) & (!g99) & (g95)) + ((!sk[59]) & (i_14_) & (i_12_) & (!i_13_) & (g99) & (!g95)) + ((!sk[59]) & (i_14_) & (i_12_) & (!i_13_) & (g99) & (g95)) + ((!sk[59]) & (i_14_) & (i_12_) & (i_13_) & (!g99) & (!g95)) + ((!sk[59]) & (i_14_) & (i_12_) & (i_13_) & (!g99) & (g95)) + ((!sk[59]) & (i_14_) & (i_12_) & (i_13_) & (g99) & (!g95)) + ((!sk[59]) & (i_14_) & (i_12_) & (i_13_) & (g99) & (g95)) + ((sk[59]) & (!i_14_) & (!i_12_) & (i_13_) & (g99) & (g95)) + ((sk[59]) & (!i_14_) & (i_12_) & (!i_13_) & (g99) & (g95)) + ((sk[59]) & (!i_14_) & (i_12_) & (i_13_) & (g99) & (g95)));
	assign g938 = (((!g99) & (!g908) & (!sk[60]) & (!g935) & (!g936) & (g937)) + ((!g99) & (!g908) & (!sk[60]) & (!g935) & (g936) & (g937)) + ((!g99) & (!g908) & (!sk[60]) & (g935) & (!g936) & (g937)) + ((!g99) & (!g908) & (!sk[60]) & (g935) & (g936) & (g937)) + ((!g99) & (!g908) & (sk[60]) & (!g935) & (!g936) & (!g937)) + ((!g99) & (g908) & (!sk[60]) & (!g935) & (!g936) & (g937)) + ((!g99) & (g908) & (!sk[60]) & (!g935) & (g936) & (g937)) + ((!g99) & (g908) & (!sk[60]) & (g935) & (!g936) & (g937)) + ((!g99) & (g908) & (!sk[60]) & (g935) & (g936) & (g937)) + ((!g99) & (g908) & (sk[60]) & (!g935) & (!g936) & (!g937)) + ((g99) & (!g908) & (!sk[60]) & (!g935) & (!g936) & (!g937)) + ((g99) & (!g908) & (!sk[60]) & (!g935) & (!g936) & (g937)) + ((g99) & (!g908) & (!sk[60]) & (!g935) & (g936) & (!g937)) + ((g99) & (!g908) & (!sk[60]) & (!g935) & (g936) & (g937)) + ((g99) & (!g908) & (!sk[60]) & (g935) & (!g936) & (!g937)) + ((g99) & (!g908) & (!sk[60]) & (g935) & (!g936) & (g937)) + ((g99) & (!g908) & (!sk[60]) & (g935) & (g936) & (!g937)) + ((g99) & (!g908) & (!sk[60]) & (g935) & (g936) & (g937)) + ((g99) & (!g908) & (sk[60]) & (!g935) & (!g936) & (!g937)) + ((g99) & (g908) & (!sk[60]) & (!g935) & (!g936) & (!g937)) + ((g99) & (g908) & (!sk[60]) & (!g935) & (!g936) & (g937)) + ((g99) & (g908) & (!sk[60]) & (!g935) & (g936) & (!g937)) + ((g99) & (g908) & (!sk[60]) & (!g935) & (g936) & (g937)) + ((g99) & (g908) & (!sk[60]) & (g935) & (!g936) & (!g937)) + ((g99) & (g908) & (!sk[60]) & (g935) & (!g936) & (g937)) + ((g99) & (g908) & (!sk[60]) & (g935) & (g936) & (!g937)) + ((g99) & (g908) & (!sk[60]) & (g935) & (g936) & (g937)));
	assign g939 = (((!g112) & (!g135) & (!g547) & (!g934) & (!sk[61]) & (g938)) + ((!g112) & (!g135) & (!g547) & (!g934) & (sk[61]) & (g938)) + ((!g112) & (!g135) & (!g547) & (g934) & (!sk[61]) & (g938)) + ((!g112) & (!g135) & (g547) & (!g934) & (!sk[61]) & (g938)) + ((!g112) & (!g135) & (g547) & (!g934) & (sk[61]) & (g938)) + ((!g112) & (!g135) & (g547) & (g934) & (!sk[61]) & (g938)) + ((!g112) & (g135) & (!g547) & (!g934) & (!sk[61]) & (g938)) + ((!g112) & (g135) & (!g547) & (g934) & (!sk[61]) & (g938)) + ((!g112) & (g135) & (g547) & (!g934) & (!sk[61]) & (g938)) + ((!g112) & (g135) & (g547) & (!g934) & (sk[61]) & (g938)) + ((!g112) & (g135) & (g547) & (g934) & (!sk[61]) & (g938)) + ((g112) & (!g135) & (!g547) & (!g934) & (!sk[61]) & (!g938)) + ((g112) & (!g135) & (!g547) & (!g934) & (!sk[61]) & (g938)) + ((g112) & (!g135) & (!g547) & (g934) & (!sk[61]) & (!g938)) + ((g112) & (!g135) & (!g547) & (g934) & (!sk[61]) & (g938)) + ((g112) & (!g135) & (g547) & (!g934) & (!sk[61]) & (!g938)) + ((g112) & (!g135) & (g547) & (!g934) & (!sk[61]) & (g938)) + ((g112) & (!g135) & (g547) & (!g934) & (sk[61]) & (g938)) + ((g112) & (!g135) & (g547) & (g934) & (!sk[61]) & (!g938)) + ((g112) & (!g135) & (g547) & (g934) & (!sk[61]) & (g938)) + ((g112) & (g135) & (!g547) & (!g934) & (!sk[61]) & (!g938)) + ((g112) & (g135) & (!g547) & (!g934) & (!sk[61]) & (g938)) + ((g112) & (g135) & (!g547) & (g934) & (!sk[61]) & (!g938)) + ((g112) & (g135) & (!g547) & (g934) & (!sk[61]) & (g938)) + ((g112) & (g135) & (g547) & (!g934) & (!sk[61]) & (!g938)) + ((g112) & (g135) & (g547) & (!g934) & (!sk[61]) & (g938)) + ((g112) & (g135) & (g547) & (!g934) & (sk[61]) & (g938)) + ((g112) & (g135) & (g547) & (g934) & (!sk[61]) & (!g938)) + ((g112) & (g135) & (g547) & (g934) & (!sk[61]) & (g938)));
	assign g940 = (((!g100) & (!g108) & (!g566) & (!g555) & (!sk[62]) & (g571)) + ((!g100) & (!g108) & (!g566) & (!g555) & (sk[62]) & (!g571)) + ((!g100) & (!g108) & (!g566) & (!g555) & (sk[62]) & (g571)) + ((!g100) & (!g108) & (!g566) & (g555) & (!sk[62]) & (g571)) + ((!g100) & (!g108) & (!g566) & (g555) & (sk[62]) & (!g571)) + ((!g100) & (!g108) & (!g566) & (g555) & (sk[62]) & (g571)) + ((!g100) & (!g108) & (g566) & (!g555) & (!sk[62]) & (g571)) + ((!g100) & (!g108) & (g566) & (!g555) & (sk[62]) & (!g571)) + ((!g100) & (!g108) & (g566) & (!g555) & (sk[62]) & (g571)) + ((!g100) & (!g108) & (g566) & (g555) & (!sk[62]) & (g571)) + ((!g100) & (!g108) & (g566) & (g555) & (sk[62]) & (!g571)) + ((!g100) & (!g108) & (g566) & (g555) & (sk[62]) & (g571)) + ((!g100) & (g108) & (!g566) & (!g555) & (!sk[62]) & (g571)) + ((!g100) & (g108) & (!g566) & (!g555) & (sk[62]) & (g571)) + ((!g100) & (g108) & (!g566) & (g555) & (!sk[62]) & (g571)) + ((!g100) & (g108) & (g566) & (!g555) & (!sk[62]) & (g571)) + ((!g100) & (g108) & (g566) & (g555) & (!sk[62]) & (g571)) + ((g100) & (!g108) & (!g566) & (!g555) & (!sk[62]) & (!g571)) + ((g100) & (!g108) & (!g566) & (!g555) & (!sk[62]) & (g571)) + ((g100) & (!g108) & (!g566) & (!g555) & (sk[62]) & (g571)) + ((g100) & (!g108) & (!g566) & (g555) & (!sk[62]) & (!g571)) + ((g100) & (!g108) & (!g566) & (g555) & (!sk[62]) & (g571)) + ((g100) & (!g108) & (g566) & (!g555) & (!sk[62]) & (!g571)) + ((g100) & (!g108) & (g566) & (!g555) & (!sk[62]) & (g571)) + ((g100) & (!g108) & (g566) & (g555) & (!sk[62]) & (!g571)) + ((g100) & (!g108) & (g566) & (g555) & (!sk[62]) & (g571)) + ((g100) & (g108) & (!g566) & (!g555) & (!sk[62]) & (!g571)) + ((g100) & (g108) & (!g566) & (!g555) & (!sk[62]) & (g571)) + ((g100) & (g108) & (!g566) & (!g555) & (sk[62]) & (g571)) + ((g100) & (g108) & (!g566) & (g555) & (!sk[62]) & (!g571)) + ((g100) & (g108) & (!g566) & (g555) & (!sk[62]) & (g571)) + ((g100) & (g108) & (g566) & (!g555) & (!sk[62]) & (!g571)) + ((g100) & (g108) & (g566) & (!g555) & (!sk[62]) & (g571)) + ((g100) & (g108) & (g566) & (g555) & (!sk[62]) & (!g571)) + ((g100) & (g108) & (g566) & (g555) & (!sk[62]) & (g571)));
	assign g941 = (((!g8) & (!g221) & (!sk[63]) & (!g101) & (!g544) & (g940)) + ((!g8) & (!g221) & (!sk[63]) & (!g101) & (g544) & (g940)) + ((!g8) & (!g221) & (!sk[63]) & (g101) & (!g544) & (g940)) + ((!g8) & (!g221) & (!sk[63]) & (g101) & (g544) & (g940)) + ((!g8) & (!g221) & (sk[63]) & (!g101) & (!g544) & (g940)) + ((!g8) & (!g221) & (sk[63]) & (!g101) & (g544) & (g940)) + ((!g8) & (g221) & (!sk[63]) & (!g101) & (!g544) & (g940)) + ((!g8) & (g221) & (!sk[63]) & (!g101) & (g544) & (g940)) + ((!g8) & (g221) & (!sk[63]) & (g101) & (!g544) & (g940)) + ((!g8) & (g221) & (!sk[63]) & (g101) & (g544) & (g940)) + ((!g8) & (g221) & (sk[63]) & (!g101) & (!g544) & (g940)) + ((!g8) & (g221) & (sk[63]) & (!g101) & (g544) & (g940)) + ((g8) & (!g221) & (!sk[63]) & (!g101) & (!g544) & (!g940)) + ((g8) & (!g221) & (!sk[63]) & (!g101) & (!g544) & (g940)) + ((g8) & (!g221) & (!sk[63]) & (!g101) & (g544) & (!g940)) + ((g8) & (!g221) & (!sk[63]) & (!g101) & (g544) & (g940)) + ((g8) & (!g221) & (!sk[63]) & (g101) & (!g544) & (!g940)) + ((g8) & (!g221) & (!sk[63]) & (g101) & (!g544) & (g940)) + ((g8) & (!g221) & (!sk[63]) & (g101) & (g544) & (!g940)) + ((g8) & (!g221) & (!sk[63]) & (g101) & (g544) & (g940)) + ((g8) & (!g221) & (sk[63]) & (!g101) & (!g544) & (g940)) + ((g8) & (!g221) & (sk[63]) & (!g101) & (g544) & (g940)) + ((g8) & (g221) & (!sk[63]) & (!g101) & (!g544) & (!g940)) + ((g8) & (g221) & (!sk[63]) & (!g101) & (!g544) & (g940)) + ((g8) & (g221) & (!sk[63]) & (!g101) & (g544) & (!g940)) + ((g8) & (g221) & (!sk[63]) & (!g101) & (g544) & (g940)) + ((g8) & (g221) & (!sk[63]) & (g101) & (!g544) & (!g940)) + ((g8) & (g221) & (!sk[63]) & (g101) & (!g544) & (g940)) + ((g8) & (g221) & (!sk[63]) & (g101) & (g544) & (!g940)) + ((g8) & (g221) & (!sk[63]) & (g101) & (g544) & (g940)) + ((g8) & (g221) & (sk[63]) & (!g101) & (!g544) & (g940)) + ((g8) & (g221) & (sk[63]) & (!g101) & (g544) & (g940)) + ((g8) & (g221) & (sk[63]) & (g101) & (g544) & (g940)));
	assign g942 = (((g923) & (g927) & (g930) & (g933) & (g939) & (g941)));
	assign g943 = (((!sk[65]) & (g220) & (!g898)) + ((!sk[65]) & (g220) & (g898)) + ((sk[65]) & (!g220) & (!g898)));
	assign g944 = (((g186) & (!g548) & (!g550) & (!g671) & (!g677) & (!g943)) + ((g186) & (!g548) & (!g550) & (!g671) & (g677) & (!g943)) + ((g186) & (!g548) & (!g550) & (!g671) & (g677) & (g943)) + ((g186) & (!g548) & (!g550) & (g671) & (!g677) & (!g943)) + ((g186) & (!g548) & (!g550) & (g671) & (!g677) & (g943)) + ((g186) & (!g548) & (!g550) & (g671) & (g677) & (!g943)) + ((g186) & (!g548) & (!g550) & (g671) & (g677) & (g943)) + ((g186) & (!g548) & (g550) & (!g671) & (!g677) & (!g943)) + ((g186) & (!g548) & (g550) & (!g671) & (!g677) & (g943)) + ((g186) & (!g548) & (g550) & (!g671) & (g677) & (!g943)) + ((g186) & (!g548) & (g550) & (!g671) & (g677) & (g943)) + ((g186) & (!g548) & (g550) & (g671) & (!g677) & (!g943)) + ((g186) & (!g548) & (g550) & (g671) & (!g677) & (g943)) + ((g186) & (!g548) & (g550) & (g671) & (g677) & (!g943)) + ((g186) & (!g548) & (g550) & (g671) & (g677) & (g943)) + ((g186) & (g548) & (!g550) & (!g671) & (!g677) & (!g943)) + ((g186) & (g548) & (!g550) & (!g671) & (!g677) & (g943)) + ((g186) & (g548) & (!g550) & (!g671) & (g677) & (!g943)) + ((g186) & (g548) & (!g550) & (!g671) & (g677) & (g943)) + ((g186) & (g548) & (!g550) & (g671) & (!g677) & (!g943)) + ((g186) & (g548) & (!g550) & (g671) & (!g677) & (g943)) + ((g186) & (g548) & (!g550) & (g671) & (g677) & (!g943)) + ((g186) & (g548) & (!g550) & (g671) & (g677) & (g943)) + ((g186) & (g548) & (g550) & (!g671) & (!g677) & (!g943)) + ((g186) & (g548) & (g550) & (!g671) & (!g677) & (g943)) + ((g186) & (g548) & (g550) & (!g671) & (g677) & (!g943)) + ((g186) & (g548) & (g550) & (!g671) & (g677) & (g943)) + ((g186) & (g548) & (g550) & (g671) & (!g677) & (!g943)) + ((g186) & (g548) & (g550) & (g671) & (!g677) & (g943)) + ((g186) & (g548) & (g550) & (g671) & (g677) & (!g943)) + ((g186) & (g548) & (g550) & (g671) & (g677) & (g943)));
	assign g945 = (((!g99) & (!g109) & (!g423) & (!g429) & (!g881) & (!g921)) + ((!g99) & (!g109) & (!g423) & (!g429) & (!g881) & (g921)) + ((!g99) & (!g109) & (!g423) & (!g429) & (g881) & (!g921)) + ((!g99) & (!g109) & (!g423) & (!g429) & (g881) & (g921)) + ((!g99) & (!g109) & (!g423) & (g429) & (!g881) & (!g921)) + ((!g99) & (!g109) & (!g423) & (g429) & (!g881) & (g921)) + ((!g99) & (!g109) & (g423) & (!g429) & (!g881) & (g921)) + ((!g99) & (!g109) & (g423) & (!g429) & (g881) & (g921)) + ((!g99) & (!g109) & (g423) & (g429) & (!g881) & (g921)) + ((!g99) & (g109) & (!g423) & (!g429) & (!g881) & (!g921)) + ((!g99) & (g109) & (!g423) & (!g429) & (!g881) & (g921)) + ((!g99) & (g109) & (!g423) & (g429) & (!g881) & (!g921)) + ((!g99) & (g109) & (!g423) & (g429) & (!g881) & (g921)) + ((!g99) & (g109) & (g423) & (!g429) & (!g881) & (g921)) + ((!g99) & (g109) & (g423) & (g429) & (!g881) & (g921)) + ((g99) & (!g109) & (!g423) & (!g429) & (!g881) & (!g921)) + ((g99) & (!g109) & (!g423) & (!g429) & (!g881) & (g921)) + ((g99) & (!g109) & (!g423) & (g429) & (!g881) & (!g921)) + ((g99) & (!g109) & (!g423) & (g429) & (!g881) & (g921)) + ((g99) & (!g109) & (g423) & (!g429) & (!g881) & (g921)) + ((g99) & (!g109) & (g423) & (g429) & (!g881) & (g921)) + ((g99) & (g109) & (!g423) & (!g429) & (!g881) & (!g921)) + ((g99) & (g109) & (!g423) & (!g429) & (!g881) & (g921)) + ((g99) & (g109) & (!g423) & (g429) & (!g881) & (!g921)) + ((g99) & (g109) & (!g423) & (g429) & (!g881) & (g921)) + ((g99) & (g109) & (g423) & (!g429) & (!g881) & (g921)) + ((g99) & (g109) & (g423) & (g429) & (!g881) & (g921)));
	assign g946 = (((!i_11_) & (i_9_) & (!i_10_) & (!g99) & (g186) & (g875)) + ((!i_11_) & (i_9_) & (!i_10_) & (g99) & (!g186) & (g875)) + ((!i_11_) & (i_9_) & (!i_10_) & (g99) & (g186) & (g875)) + ((!i_11_) & (i_9_) & (i_10_) & (!g99) & (g186) & (g875)) + ((!i_11_) & (i_9_) & (i_10_) & (g99) & (g186) & (g875)));
	assign g947 = (((!g16) & (!g270) & (g243) & (!sk[69]) & (g669)) + ((!g16) & (!g270) & (g243) & (sk[69]) & (!g669)) + ((!g16) & (!g270) & (g243) & (sk[69]) & (g669)) + ((!g16) & (g270) & (!g243) & (!sk[69]) & (!g669)) + ((!g16) & (g270) & (!g243) & (!sk[69]) & (g669)) + ((!g16) & (g270) & (g243) & (!sk[69]) & (!g669)) + ((!g16) & (g270) & (g243) & (!sk[69]) & (g669)) + ((!g16) & (g270) & (g243) & (sk[69]) & (!g669)) + ((!g16) & (g270) & (g243) & (sk[69]) & (g669)) + ((g16) & (!g270) & (g243) & (!sk[69]) & (!g669)) + ((g16) & (!g270) & (g243) & (!sk[69]) & (g669)) + ((g16) & (!g270) & (g243) & (sk[69]) & (!g669)) + ((g16) & (!g270) & (g243) & (sk[69]) & (g669)) + ((g16) & (g270) & (!g243) & (!sk[69]) & (!g669)) + ((g16) & (g270) & (!g243) & (!sk[69]) & (g669)) + ((g16) & (g270) & (g243) & (!sk[69]) & (!g669)) + ((g16) & (g270) & (g243) & (!sk[69]) & (g669)) + ((g16) & (g270) & (g243) & (sk[69]) & (!g669)));
	assign g948 = (((!g101) & (!g216) & (!g146) & (!sk[70]) & (!g946) & (g947)) + ((!g101) & (!g216) & (!g146) & (!sk[70]) & (g946) & (g947)) + ((!g101) & (!g216) & (!g146) & (sk[70]) & (!g946) & (!g947)) + ((!g101) & (!g216) & (g146) & (!sk[70]) & (!g946) & (g947)) + ((!g101) & (!g216) & (g146) & (!sk[70]) & (g946) & (g947)) + ((!g101) & (!g216) & (g146) & (sk[70]) & (!g946) & (!g947)) + ((!g101) & (g216) & (!g146) & (!sk[70]) & (!g946) & (g947)) + ((!g101) & (g216) & (!g146) & (!sk[70]) & (g946) & (g947)) + ((!g101) & (g216) & (g146) & (!sk[70]) & (!g946) & (g947)) + ((!g101) & (g216) & (g146) & (!sk[70]) & (g946) & (g947)) + ((!g101) & (g216) & (g146) & (sk[70]) & (!g946) & (!g947)) + ((g101) & (!g216) & (!g146) & (!sk[70]) & (!g946) & (!g947)) + ((g101) & (!g216) & (!g146) & (!sk[70]) & (!g946) & (g947)) + ((g101) & (!g216) & (!g146) & (!sk[70]) & (g946) & (!g947)) + ((g101) & (!g216) & (!g146) & (!sk[70]) & (g946) & (g947)) + ((g101) & (!g216) & (!g146) & (sk[70]) & (!g946) & (!g947)) + ((g101) & (!g216) & (g146) & (!sk[70]) & (!g946) & (!g947)) + ((g101) & (!g216) & (g146) & (!sk[70]) & (!g946) & (g947)) + ((g101) & (!g216) & (g146) & (!sk[70]) & (g946) & (!g947)) + ((g101) & (!g216) & (g146) & (!sk[70]) & (g946) & (g947)) + ((g101) & (!g216) & (g146) & (sk[70]) & (!g946) & (!g947)) + ((g101) & (g216) & (!g146) & (!sk[70]) & (!g946) & (!g947)) + ((g101) & (g216) & (!g146) & (!sk[70]) & (!g946) & (g947)) + ((g101) & (g216) & (!g146) & (!sk[70]) & (g946) & (!g947)) + ((g101) & (g216) & (!g146) & (!sk[70]) & (g946) & (g947)) + ((g101) & (g216) & (g146) & (!sk[70]) & (!g946) & (!g947)) + ((g101) & (g216) & (g146) & (!sk[70]) & (!g946) & (g947)) + ((g101) & (g216) & (g146) & (!sk[70]) & (g946) & (!g947)) + ((g101) & (g216) & (g146) & (!sk[70]) & (g946) & (g947)));
	assign g949 = (((!g47) & (!g546) & (!sk[71]) & (g555) & (g617)) + ((!g47) & (!g546) & (sk[71]) & (!g555) & (!g617)) + ((!g47) & (g546) & (!sk[71]) & (!g555) & (!g617)) + ((!g47) & (g546) & (!sk[71]) & (!g555) & (g617)) + ((!g47) & (g546) & (!sk[71]) & (g555) & (!g617)) + ((!g47) & (g546) & (!sk[71]) & (g555) & (g617)) + ((g47) & (!g546) & (!sk[71]) & (g555) & (!g617)) + ((g47) & (!g546) & (!sk[71]) & (g555) & (g617)) + ((g47) & (g546) & (!sk[71]) & (!g555) & (!g617)) + ((g47) & (g546) & (!sk[71]) & (!g555) & (g617)) + ((g47) & (g546) & (!sk[71]) & (g555) & (!g617)) + ((g47) & (g546) & (!sk[71]) & (g555) & (g617)));
	assign g950 = (((g221) & (!sk[72]) & (!g181) & (!g738)) + ((g221) & (!sk[72]) & (!g181) & (g738)) + ((g221) & (!sk[72]) & (g181) & (!g738)) + ((g221) & (!sk[72]) & (g181) & (g738)) + ((g221) & (sk[72]) & (!g181) & (!g738)));
	assign g951 = (((!i_8_) & (!i_6_) & (!i_7_) & (g87) & (!g949) & (!g950)) + ((!i_8_) & (!i_6_) & (!i_7_) & (g87) & (g949) & (!g950)) + ((i_8_) & (!i_6_) & (i_7_) & (g87) & (!g949) & (!g950)) + ((i_8_) & (!i_6_) & (i_7_) & (g87) & (!g949) & (g950)));
	assign g952 = (((!g88) & (!sk[74]) & (!g551) & (g561) & (g881)) + ((!g88) & (!sk[74]) & (g551) & (!g561) & (!g881)) + ((!g88) & (!sk[74]) & (g551) & (!g561) & (g881)) + ((!g88) & (!sk[74]) & (g551) & (g561) & (!g881)) + ((!g88) & (!sk[74]) & (g551) & (g561) & (g881)) + ((g88) & (!sk[74]) & (!g551) & (g561) & (!g881)) + ((g88) & (!sk[74]) & (!g551) & (g561) & (g881)) + ((g88) & (!sk[74]) & (g551) & (!g561) & (!g881)) + ((g88) & (!sk[74]) & (g551) & (!g561) & (g881)) + ((g88) & (!sk[74]) & (g551) & (g561) & (!g881)) + ((g88) & (!sk[74]) & (g551) & (g561) & (g881)) + ((g88) & (sk[74]) & (!g551) & (!g561) & (g881)) + ((g88) & (sk[74]) & (!g551) & (g561) & (!g881)) + ((g88) & (sk[74]) & (!g551) & (g561) & (g881)) + ((g88) & (sk[74]) & (g551) & (!g561) & (!g881)) + ((g88) & (sk[74]) & (g551) & (!g561) & (g881)) + ((g88) & (sk[74]) & (g551) & (g561) & (!g881)) + ((g88) & (sk[74]) & (g551) & (g561) & (g881)));
	assign g953 = (((!i_8_) & (!g100) & (!sk[75]) & (g108) & (g895)) + ((!i_8_) & (!g100) & (sk[75]) & (g108) & (g895)) + ((!i_8_) & (g100) & (!sk[75]) & (!g108) & (!g895)) + ((!i_8_) & (g100) & (!sk[75]) & (!g108) & (g895)) + ((!i_8_) & (g100) & (!sk[75]) & (g108) & (!g895)) + ((!i_8_) & (g100) & (!sk[75]) & (g108) & (g895)) + ((!i_8_) & (g100) & (sk[75]) & (!g108) & (g895)) + ((!i_8_) & (g100) & (sk[75]) & (g108) & (g895)) + ((i_8_) & (!g100) & (!sk[75]) & (g108) & (!g895)) + ((i_8_) & (!g100) & (!sk[75]) & (g108) & (g895)) + ((i_8_) & (g100) & (!sk[75]) & (!g108) & (!g895)) + ((i_8_) & (g100) & (!sk[75]) & (!g108) & (g895)) + ((i_8_) & (g100) & (!sk[75]) & (g108) & (!g895)) + ((i_8_) & (g100) & (!sk[75]) & (g108) & (g895)) + ((i_8_) & (g100) & (sk[75]) & (!g108) & (g895)) + ((i_8_) & (g100) & (sk[75]) & (g108) & (g895)));
	assign g954 = (((!i_11_) & (!i_9_) & (!i_10_) & (!sk[76]) & (!i_15_) & (g7)) + ((!i_11_) & (!i_9_) & (!i_10_) & (!sk[76]) & (i_15_) & (g7)) + ((!i_11_) & (!i_9_) & (i_10_) & (!sk[76]) & (!i_15_) & (g7)) + ((!i_11_) & (!i_9_) & (i_10_) & (!sk[76]) & (i_15_) & (g7)) + ((!i_11_) & (!i_9_) & (i_10_) & (sk[76]) & (i_15_) & (g7)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[76]) & (!i_15_) & (g7)) + ((!i_11_) & (i_9_) & (!i_10_) & (!sk[76]) & (i_15_) & (g7)) + ((!i_11_) & (i_9_) & (!i_10_) & (sk[76]) & (i_15_) & (g7)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[76]) & (!i_15_) & (g7)) + ((!i_11_) & (i_9_) & (i_10_) & (!sk[76]) & (i_15_) & (g7)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[76]) & (!i_15_) & (!g7)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[76]) & (!i_15_) & (g7)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[76]) & (i_15_) & (!g7)) + ((i_11_) & (!i_9_) & (!i_10_) & (!sk[76]) & (i_15_) & (g7)) + ((i_11_) & (!i_9_) & (!i_10_) & (sk[76]) & (i_15_) & (g7)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[76]) & (!i_15_) & (!g7)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[76]) & (!i_15_) & (g7)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[76]) & (i_15_) & (!g7)) + ((i_11_) & (!i_9_) & (i_10_) & (!sk[76]) & (i_15_) & (g7)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[76]) & (!i_15_) & (!g7)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[76]) & (!i_15_) & (g7)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[76]) & (i_15_) & (!g7)) + ((i_11_) & (i_9_) & (!i_10_) & (!sk[76]) & (i_15_) & (g7)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[76]) & (!i_15_) & (!g7)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[76]) & (!i_15_) & (g7)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[76]) & (i_15_) & (!g7)) + ((i_11_) & (i_9_) & (i_10_) & (!sk[76]) & (i_15_) & (g7)));
	assign g955 = (((!g59) & (!sk[77]) & (!g66) & (!g118) & (!g943) & (g954)) + ((!g59) & (!sk[77]) & (!g66) & (!g118) & (g943) & (g954)) + ((!g59) & (!sk[77]) & (!g66) & (g118) & (!g943) & (g954)) + ((!g59) & (!sk[77]) & (!g66) & (g118) & (g943) & (g954)) + ((!g59) & (!sk[77]) & (g66) & (!g118) & (!g943) & (g954)) + ((!g59) & (!sk[77]) & (g66) & (!g118) & (g943) & (g954)) + ((!g59) & (!sk[77]) & (g66) & (g118) & (!g943) & (g954)) + ((!g59) & (!sk[77]) & (g66) & (g118) & (g943) & (g954)) + ((!g59) & (sk[77]) & (!g66) & (!g118) & (!g943) & (!g954)) + ((!g59) & (sk[77]) & (!g66) & (!g118) & (!g943) & (g954)) + ((!g59) & (sk[77]) & (!g66) & (!g118) & (g943) & (!g954)) + ((!g59) & (sk[77]) & (!g66) & (!g118) & (g943) & (g954)) + ((!g59) & (sk[77]) & (!g66) & (g118) & (g943) & (!g954)) + ((!g59) & (sk[77]) & (!g66) & (g118) & (g943) & (g954)) + ((!g59) & (sk[77]) & (g66) & (!g118) & (!g943) & (!g954)) + ((!g59) & (sk[77]) & (g66) & (!g118) & (!g943) & (g954)) + ((!g59) & (sk[77]) & (g66) & (!g118) & (g943) & (!g954)) + ((!g59) & (sk[77]) & (g66) & (!g118) & (g943) & (g954)) + ((g59) & (!sk[77]) & (!g66) & (!g118) & (!g943) & (!g954)) + ((g59) & (!sk[77]) & (!g66) & (!g118) & (!g943) & (g954)) + ((g59) & (!sk[77]) & (!g66) & (!g118) & (g943) & (!g954)) + ((g59) & (!sk[77]) & (!g66) & (!g118) & (g943) & (g954)) + ((g59) & (!sk[77]) & (!g66) & (g118) & (!g943) & (!g954)) + ((g59) & (!sk[77]) & (!g66) & (g118) & (!g943) & (g954)) + ((g59) & (!sk[77]) & (!g66) & (g118) & (g943) & (!g954)) + ((g59) & (!sk[77]) & (!g66) & (g118) & (g943) & (g954)) + ((g59) & (!sk[77]) & (g66) & (!g118) & (!g943) & (!g954)) + ((g59) & (!sk[77]) & (g66) & (!g118) & (!g943) & (g954)) + ((g59) & (!sk[77]) & (g66) & (!g118) & (g943) & (!g954)) + ((g59) & (!sk[77]) & (g66) & (!g118) & (g943) & (g954)) + ((g59) & (!sk[77]) & (g66) & (g118) & (!g943) & (!g954)) + ((g59) & (!sk[77]) & (g66) & (g118) & (!g943) & (g954)) + ((g59) & (!sk[77]) & (g66) & (g118) & (g943) & (!g954)) + ((g59) & (!sk[77]) & (g66) & (g118) & (g943) & (g954)) + ((g59) & (sk[77]) & (!g66) & (!g118) & (!g943) & (!g954)) + ((g59) & (sk[77]) & (!g66) & (!g118) & (g943) & (!g954)) + ((g59) & (sk[77]) & (!g66) & (g118) & (g943) & (!g954)) + ((g59) & (sk[77]) & (g66) & (!g118) & (!g943) & (!g954)) + ((g59) & (sk[77]) & (g66) & (!g118) & (g943) & (!g954)));
	assign g956 = (((!sk[78]) & (!g284) & (!g676) & (!g952) & (!g953) & (g955)) + ((!sk[78]) & (!g284) & (!g676) & (!g952) & (g953) & (g955)) + ((!sk[78]) & (!g284) & (!g676) & (g952) & (!g953) & (g955)) + ((!sk[78]) & (!g284) & (!g676) & (g952) & (g953) & (g955)) + ((!sk[78]) & (!g284) & (g676) & (!g952) & (!g953) & (g955)) + ((!sk[78]) & (!g284) & (g676) & (!g952) & (g953) & (g955)) + ((!sk[78]) & (!g284) & (g676) & (g952) & (!g953) & (g955)) + ((!sk[78]) & (!g284) & (g676) & (g952) & (g953) & (g955)) + ((!sk[78]) & (g284) & (!g676) & (!g952) & (!g953) & (!g955)) + ((!sk[78]) & (g284) & (!g676) & (!g952) & (!g953) & (g955)) + ((!sk[78]) & (g284) & (!g676) & (!g952) & (g953) & (!g955)) + ((!sk[78]) & (g284) & (!g676) & (!g952) & (g953) & (g955)) + ((!sk[78]) & (g284) & (!g676) & (g952) & (!g953) & (!g955)) + ((!sk[78]) & (g284) & (!g676) & (g952) & (!g953) & (g955)) + ((!sk[78]) & (g284) & (!g676) & (g952) & (g953) & (!g955)) + ((!sk[78]) & (g284) & (!g676) & (g952) & (g953) & (g955)) + ((!sk[78]) & (g284) & (g676) & (!g952) & (!g953) & (!g955)) + ((!sk[78]) & (g284) & (g676) & (!g952) & (!g953) & (g955)) + ((!sk[78]) & (g284) & (g676) & (!g952) & (g953) & (!g955)) + ((!sk[78]) & (g284) & (g676) & (!g952) & (g953) & (g955)) + ((!sk[78]) & (g284) & (g676) & (g952) & (!g953) & (!g955)) + ((!sk[78]) & (g284) & (g676) & (g952) & (!g953) & (g955)) + ((!sk[78]) & (g284) & (g676) & (g952) & (g953) & (!g955)) + ((!sk[78]) & (g284) & (g676) & (g952) & (g953) & (g955)) + ((sk[78]) & (!g284) & (!g676) & (!g952) & (!g953) & (g955)) + ((sk[78]) & (!g284) & (g676) & (!g952) & (!g953) & (g955)) + ((sk[78]) & (g284) & (!g676) & (!g952) & (!g953) & (g955)));
	assign g957 = (((!i_11_) & (!i_9_) & (!sk[79]) & (i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (!sk[79]) & (!i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (!sk[79]) & (!i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (!sk[79]) & (i_10_) & (!i_15_)) + ((!i_11_) & (i_9_) & (!sk[79]) & (i_10_) & (i_15_)) + ((!i_11_) & (i_9_) & (sk[79]) & (i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (!sk[79]) & (i_10_) & (!i_15_)) + ((i_11_) & (!i_9_) & (!sk[79]) & (i_10_) & (i_15_)) + ((i_11_) & (!i_9_) & (sk[79]) & (!i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (!sk[79]) & (!i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (!sk[79]) & (!i_10_) & (i_15_)) + ((i_11_) & (i_9_) & (!sk[79]) & (i_10_) & (!i_15_)) + ((i_11_) & (i_9_) & (!sk[79]) & (i_10_) & (i_15_)));
	assign g958 = (((!i_15_) & (!g13) & (!sk[80]) & (!g59) & (!g112) & (g957)) + ((!i_15_) & (!g13) & (!sk[80]) & (!g59) & (g112) & (g957)) + ((!i_15_) & (!g13) & (!sk[80]) & (g59) & (!g112) & (g957)) + ((!i_15_) & (!g13) & (!sk[80]) & (g59) & (g112) & (g957)) + ((!i_15_) & (g13) & (!sk[80]) & (!g59) & (!g112) & (g957)) + ((!i_15_) & (g13) & (!sk[80]) & (!g59) & (g112) & (g957)) + ((!i_15_) & (g13) & (!sk[80]) & (g59) & (!g112) & (g957)) + ((!i_15_) & (g13) & (!sk[80]) & (g59) & (g112) & (g957)) + ((!i_15_) & (g13) & (sk[80]) & (!g59) & (g112) & (g957)) + ((!i_15_) & (g13) & (sk[80]) & (g59) & (!g112) & (g957)) + ((!i_15_) & (g13) & (sk[80]) & (g59) & (g112) & (g957)) + ((i_15_) & (!g13) & (!sk[80]) & (!g59) & (!g112) & (!g957)) + ((i_15_) & (!g13) & (!sk[80]) & (!g59) & (!g112) & (g957)) + ((i_15_) & (!g13) & (!sk[80]) & (!g59) & (g112) & (!g957)) + ((i_15_) & (!g13) & (!sk[80]) & (!g59) & (g112) & (g957)) + ((i_15_) & (!g13) & (!sk[80]) & (g59) & (!g112) & (!g957)) + ((i_15_) & (!g13) & (!sk[80]) & (g59) & (!g112) & (g957)) + ((i_15_) & (!g13) & (!sk[80]) & (g59) & (g112) & (!g957)) + ((i_15_) & (!g13) & (!sk[80]) & (g59) & (g112) & (g957)) + ((i_15_) & (g13) & (!sk[80]) & (!g59) & (!g112) & (!g957)) + ((i_15_) & (g13) & (!sk[80]) & (!g59) & (!g112) & (g957)) + ((i_15_) & (g13) & (!sk[80]) & (!g59) & (g112) & (!g957)) + ((i_15_) & (g13) & (!sk[80]) & (!g59) & (g112) & (g957)) + ((i_15_) & (g13) & (!sk[80]) & (g59) & (!g112) & (!g957)) + ((i_15_) & (g13) & (!sk[80]) & (g59) & (!g112) & (g957)) + ((i_15_) & (g13) & (!sk[80]) & (g59) & (g112) & (!g957)) + ((i_15_) & (g13) & (!sk[80]) & (g59) & (g112) & (g957)) + ((i_15_) & (g13) & (sk[80]) & (!g59) & (!g112) & (g957)) + ((i_15_) & (g13) & (sk[80]) & (!g59) & (g112) & (g957)) + ((i_15_) & (g13) & (sk[80]) & (g59) & (!g112) & (g957)) + ((i_15_) & (g13) & (sk[80]) & (g59) & (g112) & (g957)));
	assign g959 = (((!i_15_) & (!g134) & (!g251) & (!g576) & (!g895) & (!g958)) + ((!i_15_) & (!g134) & (!g251) & (!g576) & (g895) & (!g958)) + ((!i_15_) & (!g134) & (!g251) & (g576) & (!g895) & (!g958)) + ((!i_15_) & (!g134) & (!g251) & (g576) & (g895) & (!g958)) + ((!i_15_) & (!g134) & (g251) & (!g576) & (!g895) & (!g958)) + ((!i_15_) & (!g134) & (g251) & (!g576) & (g895) & (!g958)) + ((!i_15_) & (!g134) & (g251) & (g576) & (!g895) & (!g958)) + ((!i_15_) & (!g134) & (g251) & (g576) & (g895) & (!g958)) + ((!i_15_) & (g134) & (!g251) & (g576) & (!g895) & (!g958)) + ((!i_15_) & (g134) & (g251) & (g576) & (!g895) & (!g958)) + ((i_15_) & (!g134) & (!g251) & (!g576) & (!g895) & (!g958)) + ((i_15_) & (!g134) & (!g251) & (!g576) & (!g895) & (g958)) + ((i_15_) & (!g134) & (!g251) & (!g576) & (g895) & (!g958)) + ((i_15_) & (!g134) & (!g251) & (!g576) & (g895) & (g958)) + ((i_15_) & (!g134) & (!g251) & (g576) & (!g895) & (!g958)) + ((i_15_) & (!g134) & (!g251) & (g576) & (!g895) & (g958)) + ((i_15_) & (!g134) & (!g251) & (g576) & (g895) & (!g958)) + ((i_15_) & (!g134) & (!g251) & (g576) & (g895) & (g958)) + ((i_15_) & (!g134) & (g251) & (!g576) & (!g895) & (!g958)) + ((i_15_) & (!g134) & (g251) & (!g576) & (g895) & (!g958)) + ((i_15_) & (!g134) & (g251) & (g576) & (!g895) & (!g958)) + ((i_15_) & (!g134) & (g251) & (g576) & (g895) & (!g958)) + ((i_15_) & (g134) & (!g251) & (g576) & (!g895) & (!g958)) + ((i_15_) & (g134) & (g251) & (g576) & (!g895) & (!g958)));
	assign g960 = (((!g944) & (g945) & (g948) & (!g951) & (g956) & (g959)));
	assign g961 = (((!sk[83]) & (!i_14_) & (!i_12_) & (i_13_) & (g104)) + ((!sk[83]) & (!i_14_) & (i_12_) & (!i_13_) & (!g104)) + ((!sk[83]) & (!i_14_) & (i_12_) & (!i_13_) & (g104)) + ((!sk[83]) & (!i_14_) & (i_12_) & (i_13_) & (!g104)) + ((!sk[83]) & (!i_14_) & (i_12_) & (i_13_) & (g104)) + ((!sk[83]) & (i_14_) & (!i_12_) & (i_13_) & (!g104)) + ((!sk[83]) & (i_14_) & (!i_12_) & (i_13_) & (g104)) + ((!sk[83]) & (i_14_) & (i_12_) & (!i_13_) & (!g104)) + ((!sk[83]) & (i_14_) & (i_12_) & (!i_13_) & (g104)) + ((!sk[83]) & (i_14_) & (i_12_) & (i_13_) & (!g104)) + ((!sk[83]) & (i_14_) & (i_12_) & (i_13_) & (g104)) + ((sk[83]) & (!i_14_) & (!i_12_) & (i_13_) & (g104)) + ((sk[83]) & (!i_14_) & (i_12_) & (!i_13_) & (g104)) + ((sk[83]) & (!i_14_) & (i_12_) & (i_13_) & (g104)));
	assign g962 = (((!g23) & (!sk[84]) & (!g206) & (!g323) & (!g561) & (g921)) + ((!g23) & (!sk[84]) & (!g206) & (!g323) & (g561) & (g921)) + ((!g23) & (!sk[84]) & (!g206) & (g323) & (!g561) & (g921)) + ((!g23) & (!sk[84]) & (!g206) & (g323) & (g561) & (g921)) + ((!g23) & (!sk[84]) & (g206) & (!g323) & (!g561) & (g921)) + ((!g23) & (!sk[84]) & (g206) & (!g323) & (g561) & (g921)) + ((!g23) & (!sk[84]) & (g206) & (g323) & (!g561) & (g921)) + ((!g23) & (!sk[84]) & (g206) & (g323) & (g561) & (g921)) + ((!g23) & (sk[84]) & (!g206) & (g323) & (!g561) & (!g921)) + ((!g23) & (sk[84]) & (!g206) & (g323) & (!g561) & (g921)) + ((!g23) & (sk[84]) & (!g206) & (g323) & (g561) & (!g921)) + ((!g23) & (sk[84]) & (!g206) & (g323) & (g561) & (g921)) + ((!g23) & (sk[84]) & (g206) & (g323) & (!g561) & (!g921)) + ((!g23) & (sk[84]) & (g206) & (g323) & (g561) & (!g921)) + ((!g23) & (sk[84]) & (g206) & (g323) & (g561) & (g921)) + ((g23) & (!sk[84]) & (!g206) & (!g323) & (!g561) & (!g921)) + ((g23) & (!sk[84]) & (!g206) & (!g323) & (!g561) & (g921)) + ((g23) & (!sk[84]) & (!g206) & (!g323) & (g561) & (!g921)) + ((g23) & (!sk[84]) & (!g206) & (!g323) & (g561) & (g921)) + ((g23) & (!sk[84]) & (!g206) & (g323) & (!g561) & (!g921)) + ((g23) & (!sk[84]) & (!g206) & (g323) & (!g561) & (g921)) + ((g23) & (!sk[84]) & (!g206) & (g323) & (g561) & (!g921)) + ((g23) & (!sk[84]) & (!g206) & (g323) & (g561) & (g921)) + ((g23) & (!sk[84]) & (g206) & (!g323) & (!g561) & (!g921)) + ((g23) & (!sk[84]) & (g206) & (!g323) & (!g561) & (g921)) + ((g23) & (!sk[84]) & (g206) & (!g323) & (g561) & (!g921)) + ((g23) & (!sk[84]) & (g206) & (!g323) & (g561) & (g921)) + ((g23) & (!sk[84]) & (g206) & (g323) & (!g561) & (!g921)) + ((g23) & (!sk[84]) & (g206) & (g323) & (!g561) & (g921)) + ((g23) & (!sk[84]) & (g206) & (g323) & (g561) & (!g921)) + ((g23) & (!sk[84]) & (g206) & (g323) & (g561) & (g921)) + ((g23) & (sk[84]) & (!g206) & (g323) & (!g561) & (!g921)) + ((g23) & (sk[84]) & (!g206) & (g323) & (!g561) & (g921)) + ((g23) & (sk[84]) & (!g206) & (g323) & (g561) & (!g921)) + ((g23) & (sk[84]) & (!g206) & (g323) & (g561) & (g921)) + ((g23) & (sk[84]) & (g206) & (g323) & (!g561) & (!g921)) + ((g23) & (sk[84]) & (g206) & (g323) & (!g561) & (g921)) + ((g23) & (sk[84]) & (g206) & (g323) & (g561) & (!g921)) + ((g23) & (sk[84]) & (g206) & (g323) & (g561) & (g921)));
	assign g963 = (((!g112) & (!g135) & (!sk[85]) & (g532) & (g962)) + ((!g112) & (!g135) & (sk[85]) & (!g532) & (!g962)) + ((!g112) & (!g135) & (sk[85]) & (g532) & (!g962)) + ((!g112) & (g135) & (!sk[85]) & (!g532) & (!g962)) + ((!g112) & (g135) & (!sk[85]) & (!g532) & (g962)) + ((!g112) & (g135) & (!sk[85]) & (g532) & (!g962)) + ((!g112) & (g135) & (!sk[85]) & (g532) & (g962)) + ((!g112) & (g135) & (sk[85]) & (!g532) & (!g962)) + ((g112) & (!g135) & (!sk[85]) & (g532) & (!g962)) + ((g112) & (!g135) & (!sk[85]) & (g532) & (g962)) + ((g112) & (!g135) & (sk[85]) & (!g532) & (!g962)) + ((g112) & (g135) & (!sk[85]) & (!g532) & (!g962)) + ((g112) & (g135) & (!sk[85]) & (!g532) & (g962)) + ((g112) & (g135) & (!sk[85]) & (g532) & (!g962)) + ((g112) & (g135) & (!sk[85]) & (g532) & (g962)) + ((g112) & (g135) & (sk[85]) & (!g532) & (!g962)));
	assign g964 = (((!i_12_) & (!i_13_) & (!i_8_) & (!g108) & (!sk[86]) & (g135)) + ((!i_12_) & (!i_13_) & (!i_8_) & (g108) & (!sk[86]) & (g135)) + ((!i_12_) & (!i_13_) & (i_8_) & (!g108) & (!sk[86]) & (g135)) + ((!i_12_) & (!i_13_) & (i_8_) & (g108) & (!sk[86]) & (g135)) + ((!i_12_) & (i_13_) & (!i_8_) & (!g108) & (!sk[86]) & (g135)) + ((!i_12_) & (i_13_) & (!i_8_) & (g108) & (!sk[86]) & (g135)) + ((!i_12_) & (i_13_) & (i_8_) & (!g108) & (!sk[86]) & (g135)) + ((!i_12_) & (i_13_) & (i_8_) & (g108) & (!sk[86]) & (g135)) + ((i_12_) & (!i_13_) & (!i_8_) & (!g108) & (!sk[86]) & (!g135)) + ((i_12_) & (!i_13_) & (!i_8_) & (!g108) & (!sk[86]) & (g135)) + ((i_12_) & (!i_13_) & (!i_8_) & (g108) & (!sk[86]) & (!g135)) + ((i_12_) & (!i_13_) & (!i_8_) & (g108) & (!sk[86]) & (g135)) + ((i_12_) & (!i_13_) & (i_8_) & (!g108) & (!sk[86]) & (!g135)) + ((i_12_) & (!i_13_) & (i_8_) & (!g108) & (!sk[86]) & (g135)) + ((i_12_) & (!i_13_) & (i_8_) & (!g108) & (sk[86]) & (g135)) + ((i_12_) & (!i_13_) & (i_8_) & (g108) & (!sk[86]) & (!g135)) + ((i_12_) & (!i_13_) & (i_8_) & (g108) & (!sk[86]) & (g135)) + ((i_12_) & (!i_13_) & (i_8_) & (g108) & (sk[86]) & (g135)) + ((i_12_) & (i_13_) & (!i_8_) & (!g108) & (!sk[86]) & (!g135)) + ((i_12_) & (i_13_) & (!i_8_) & (!g108) & (!sk[86]) & (g135)) + ((i_12_) & (i_13_) & (!i_8_) & (g108) & (!sk[86]) & (!g135)) + ((i_12_) & (i_13_) & (!i_8_) & (g108) & (!sk[86]) & (g135)) + ((i_12_) & (i_13_) & (!i_8_) & (g108) & (sk[86]) & (!g135)) + ((i_12_) & (i_13_) & (!i_8_) & (g108) & (sk[86]) & (g135)) + ((i_12_) & (i_13_) & (i_8_) & (!g108) & (!sk[86]) & (!g135)) + ((i_12_) & (i_13_) & (i_8_) & (!g108) & (!sk[86]) & (g135)) + ((i_12_) & (i_13_) & (i_8_) & (g108) & (!sk[86]) & (!g135)) + ((i_12_) & (i_13_) & (i_8_) & (g108) & (!sk[86]) & (g135)));
	assign g965 = (((!g548) & (!g550) & (!g561) & (sk[87]) & (!g908)) + ((!g548) & (!g550) & (g561) & (!sk[87]) & (g908)) + ((!g548) & (g550) & (!g561) & (!sk[87]) & (!g908)) + ((!g548) & (g550) & (!g561) & (!sk[87]) & (g908)) + ((!g548) & (g550) & (g561) & (!sk[87]) & (!g908)) + ((!g548) & (g550) & (g561) & (!sk[87]) & (g908)) + ((g548) & (!g550) & (g561) & (!sk[87]) & (!g908)) + ((g548) & (!g550) & (g561) & (!sk[87]) & (g908)) + ((g548) & (g550) & (!g561) & (!sk[87]) & (!g908)) + ((g548) & (g550) & (!g561) & (!sk[87]) & (g908)) + ((g548) & (g550) & (g561) & (!sk[87]) & (!g908)) + ((g548) & (g550) & (g561) & (!sk[87]) & (g908)));
	assign g966 = (((!i_14_) & (!sk[88]) & (!g131) & (!g277) & (!g964) & (g965)) + ((!i_14_) & (!sk[88]) & (!g131) & (!g277) & (g964) & (g965)) + ((!i_14_) & (!sk[88]) & (!g131) & (g277) & (!g964) & (g965)) + ((!i_14_) & (!sk[88]) & (!g131) & (g277) & (g964) & (g965)) + ((!i_14_) & (!sk[88]) & (g131) & (!g277) & (!g964) & (g965)) + ((!i_14_) & (!sk[88]) & (g131) & (!g277) & (g964) & (g965)) + ((!i_14_) & (!sk[88]) & (g131) & (g277) & (!g964) & (g965)) + ((!i_14_) & (!sk[88]) & (g131) & (g277) & (g964) & (g965)) + ((!i_14_) & (sk[88]) & (!g131) & (!g277) & (!g964) & (!g965)) + ((!i_14_) & (sk[88]) & (!g131) & (!g277) & (g964) & (!g965)) + ((!i_14_) & (sk[88]) & (g131) & (!g277) & (!g964) & (!g965)) + ((!i_14_) & (sk[88]) & (g131) & (!g277) & (g964) & (!g965)) + ((!i_14_) & (sk[88]) & (g131) & (!g277) & (g964) & (g965)) + ((!i_14_) & (sk[88]) & (g131) & (g277) & (g964) & (!g965)) + ((!i_14_) & (sk[88]) & (g131) & (g277) & (g964) & (g965)) + ((i_14_) & (!sk[88]) & (!g131) & (!g277) & (!g964) & (!g965)) + ((i_14_) & (!sk[88]) & (!g131) & (!g277) & (!g964) & (g965)) + ((i_14_) & (!sk[88]) & (!g131) & (!g277) & (g964) & (!g965)) + ((i_14_) & (!sk[88]) & (!g131) & (!g277) & (g964) & (g965)) + ((i_14_) & (!sk[88]) & (!g131) & (g277) & (!g964) & (!g965)) + ((i_14_) & (!sk[88]) & (!g131) & (g277) & (!g964) & (g965)) + ((i_14_) & (!sk[88]) & (!g131) & (g277) & (g964) & (!g965)) + ((i_14_) & (!sk[88]) & (!g131) & (g277) & (g964) & (g965)) + ((i_14_) & (!sk[88]) & (g131) & (!g277) & (!g964) & (!g965)) + ((i_14_) & (!sk[88]) & (g131) & (!g277) & (!g964) & (g965)) + ((i_14_) & (!sk[88]) & (g131) & (!g277) & (g964) & (!g965)) + ((i_14_) & (!sk[88]) & (g131) & (!g277) & (g964) & (g965)) + ((i_14_) & (!sk[88]) & (g131) & (g277) & (!g964) & (!g965)) + ((i_14_) & (!sk[88]) & (g131) & (g277) & (!g964) & (g965)) + ((i_14_) & (!sk[88]) & (g131) & (g277) & (g964) & (!g965)) + ((i_14_) & (!sk[88]) & (g131) & (g277) & (g964) & (g965)) + ((i_14_) & (sk[88]) & (!g131) & (!g277) & (!g964) & (!g965)) + ((i_14_) & (sk[88]) & (!g131) & (!g277) & (g964) & (!g965)) + ((i_14_) & (sk[88]) & (g131) & (!g277) & (!g964) & (!g965)) + ((i_14_) & (sk[88]) & (g131) & (!g277) & (g964) & (!g965)));
	assign g967 = (((!g109) & (!g551) & (!g495) & (!g961) & (g963) & (!g966)) + ((!g109) & (!g551) & (!g495) & (g961) & (g963) & (!g966)) + ((!g109) & (!g551) & (g495) & (!g961) & (g963) & (!g966)) + ((!g109) & (!g551) & (g495) & (g961) & (g963) & (!g966)) + ((!g109) & (g551) & (!g495) & (!g961) & (g963) & (!g966)) + ((!g109) & (g551) & (!g495) & (g961) & (g963) & (!g966)) + ((g109) & (!g551) & (!g495) & (!g961) & (g963) & (!g966)) + ((g109) & (!g551) & (g495) & (!g961) & (g963) & (!g966)) + ((g109) & (g551) & (!g495) & (!g961) & (g963) & (!g966)));
	assign g968 = (((g322) & (g325) & (g335) & (g374) & (g960) & (g967)));
	assign o_9_ = (((g73) & (!g858) & (!g879) & (!g918) & (!g942) & (!g968)) + ((g73) & (!g858) & (!g879) & (!g918) & (!g942) & (g968)) + ((g73) & (!g858) & (!g879) & (!g918) & (g942) & (!g968)) + ((g73) & (!g858) & (!g879) & (!g918) & (g942) & (g968)) + ((g73) & (!g858) & (!g879) & (g918) & (!g942) & (!g968)) + ((g73) & (!g858) & (!g879) & (g918) & (!g942) & (g968)) + ((g73) & (!g858) & (!g879) & (g918) & (g942) & (!g968)) + ((g73) & (!g858) & (!g879) & (g918) & (g942) & (g968)) + ((g73) & (!g858) & (g879) & (!g918) & (!g942) & (!g968)) + ((g73) & (!g858) & (g879) & (!g918) & (!g942) & (g968)) + ((g73) & (!g858) & (g879) & (!g918) & (g942) & (!g968)) + ((g73) & (!g858) & (g879) & (!g918) & (g942) & (g968)) + ((g73) & (!g858) & (g879) & (g918) & (!g942) & (!g968)) + ((g73) & (!g858) & (g879) & (g918) & (!g942) & (g968)) + ((g73) & (!g858) & (g879) & (g918) & (g942) & (!g968)) + ((g73) & (!g858) & (g879) & (g918) & (g942) & (g968)) + ((g73) & (g858) & (!g879) & (!g918) & (!g942) & (!g968)) + ((g73) & (g858) & (!g879) & (!g918) & (!g942) & (g968)) + ((g73) & (g858) & (!g879) & (!g918) & (g942) & (!g968)) + ((g73) & (g858) & (!g879) & (!g918) & (g942) & (g968)) + ((g73) & (g858) & (!g879) & (g918) & (!g942) & (!g968)) + ((g73) & (g858) & (!g879) & (g918) & (!g942) & (g968)) + ((g73) & (g858) & (!g879) & (g918) & (g942) & (!g968)) + ((g73) & (g858) & (!g879) & (g918) & (g942) & (g968)) + ((g73) & (g858) & (g879) & (!g918) & (!g942) & (!g968)) + ((g73) & (g858) & (g879) & (!g918) & (!g942) & (g968)) + ((g73) & (g858) & (g879) & (!g918) & (g942) & (!g968)) + ((g73) & (g858) & (g879) & (!g918) & (g942) & (g968)) + ((g73) & (g858) & (g879) & (g918) & (!g942) & (!g968)) + ((g73) & (g858) & (g879) & (g918) & (!g942) & (g968)) + ((g73) & (g858) & (g879) & (g918) & (g942) & (!g968)));
	assign g970 = (((!g20) & (g101) & (sk[92]) & (!g806)) + ((!g20) & (g101) & (sk[92]) & (g806)) + ((g20) & (!g101) & (!sk[92]) & (!g806)) + ((g20) & (!g101) & (!sk[92]) & (g806)) + ((g20) & (g101) & (!sk[92]) & (!g806)) + ((g20) & (g101) & (!sk[92]) & (g806)) + ((g20) & (g101) & (sk[92]) & (g806)));
	assign g971 = (((!g101) & (!sk[93]) & (!g339) & (g465) & (g924)) + ((!g101) & (!sk[93]) & (g339) & (!g465) & (!g924)) + ((!g101) & (!sk[93]) & (g339) & (!g465) & (g924)) + ((!g101) & (!sk[93]) & (g339) & (g465) & (!g924)) + ((!g101) & (!sk[93]) & (g339) & (g465) & (g924)) + ((!g101) & (sk[93]) & (!g339) & (!g465) & (!g924)) + ((!g101) & (sk[93]) & (!g339) & (g465) & (!g924)) + ((!g101) & (sk[93]) & (g339) & (!g465) & (!g924)) + ((!g101) & (sk[93]) & (g339) & (g465) & (!g924)) + ((g101) & (!sk[93]) & (!g339) & (g465) & (!g924)) + ((g101) & (!sk[93]) & (!g339) & (g465) & (g924)) + ((g101) & (!sk[93]) & (g339) & (!g465) & (!g924)) + ((g101) & (!sk[93]) & (g339) & (!g465) & (g924)) + ((g101) & (!sk[93]) & (g339) & (g465) & (!g924)) + ((g101) & (!sk[93]) & (g339) & (g465) & (g924)) + ((g101) & (sk[93]) & (!g339) & (g465) & (!g924)));
	assign g972 = (((!sk[94]) & (!i_8_) & (!g21) & (!g22) & (!g100) & (g711)) + ((!sk[94]) & (!i_8_) & (!g21) & (!g22) & (g100) & (g711)) + ((!sk[94]) & (!i_8_) & (!g21) & (g22) & (!g100) & (g711)) + ((!sk[94]) & (!i_8_) & (!g21) & (g22) & (g100) & (g711)) + ((!sk[94]) & (!i_8_) & (g21) & (!g22) & (!g100) & (g711)) + ((!sk[94]) & (!i_8_) & (g21) & (!g22) & (g100) & (g711)) + ((!sk[94]) & (!i_8_) & (g21) & (g22) & (!g100) & (g711)) + ((!sk[94]) & (!i_8_) & (g21) & (g22) & (g100) & (g711)) + ((!sk[94]) & (i_8_) & (!g21) & (!g22) & (!g100) & (!g711)) + ((!sk[94]) & (i_8_) & (!g21) & (!g22) & (!g100) & (g711)) + ((!sk[94]) & (i_8_) & (!g21) & (!g22) & (g100) & (!g711)) + ((!sk[94]) & (i_8_) & (!g21) & (!g22) & (g100) & (g711)) + ((!sk[94]) & (i_8_) & (!g21) & (g22) & (!g100) & (!g711)) + ((!sk[94]) & (i_8_) & (!g21) & (g22) & (!g100) & (g711)) + ((!sk[94]) & (i_8_) & (!g21) & (g22) & (g100) & (!g711)) + ((!sk[94]) & (i_8_) & (!g21) & (g22) & (g100) & (g711)) + ((!sk[94]) & (i_8_) & (g21) & (!g22) & (!g100) & (!g711)) + ((!sk[94]) & (i_8_) & (g21) & (!g22) & (!g100) & (g711)) + ((!sk[94]) & (i_8_) & (g21) & (!g22) & (g100) & (!g711)) + ((!sk[94]) & (i_8_) & (g21) & (!g22) & (g100) & (g711)) + ((!sk[94]) & (i_8_) & (g21) & (g22) & (!g100) & (!g711)) + ((!sk[94]) & (i_8_) & (g21) & (g22) & (!g100) & (g711)) + ((!sk[94]) & (i_8_) & (g21) & (g22) & (g100) & (!g711)) + ((!sk[94]) & (i_8_) & (g21) & (g22) & (g100) & (g711)) + ((sk[94]) & (i_8_) & (!g21) & (g22) & (g100) & (g711)) + ((sk[94]) & (i_8_) & (g21) & (!g22) & (g100) & (!g711)) + ((sk[94]) & (i_8_) & (g21) & (!g22) & (g100) & (g711)) + ((sk[94]) & (i_8_) & (g21) & (g22) & (g100) & (!g711)) + ((sk[94]) & (i_8_) & (g21) & (g22) & (g100) & (g711)));
	assign g973 = (((!i_14_) & (!i_12_) & (i_13_) & (!g18) & (!g15) & (g99)) + ((!i_14_) & (!i_12_) & (i_13_) & (g18) & (!g15) & (g99)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g18) & (!g15) & (g99)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g18) & (g15) & (g99)) + ((i_14_) & (!i_12_) & (!i_13_) & (g18) & (!g15) & (g99)) + ((i_14_) & (i_12_) & (!i_13_) & (!g18) & (!g15) & (g99)) + ((i_14_) & (i_12_) & (!i_13_) & (!g18) & (g15) & (g99)) + ((i_14_) & (i_12_) & (i_13_) & (!g18) & (!g15) & (g99)) + ((i_14_) & (i_12_) & (i_13_) & (g18) & (!g15) & (g99)));
	assign g974 = (((!g99) & (!g152) & (!g465) & (!g462) & (!g972) & (!g973)) + ((!g99) & (!g152) & (!g465) & (g462) & (!g972) & (!g973)) + ((!g99) & (!g152) & (g465) & (!g462) & (!g972) & (!g973)) + ((!g99) & (!g152) & (g465) & (g462) & (!g972) & (!g973)) + ((g99) & (!g152) & (g465) & (g462) & (!g972) & (!g973)));
	assign g975 = (((!sk[97]) & (!g47) & (!g101) & (!g172) & (!g142) & (g883)) + ((!sk[97]) & (!g47) & (!g101) & (!g172) & (g142) & (g883)) + ((!sk[97]) & (!g47) & (!g101) & (g172) & (!g142) & (g883)) + ((!sk[97]) & (!g47) & (!g101) & (g172) & (g142) & (g883)) + ((!sk[97]) & (!g47) & (g101) & (!g172) & (!g142) & (g883)) + ((!sk[97]) & (!g47) & (g101) & (!g172) & (g142) & (g883)) + ((!sk[97]) & (!g47) & (g101) & (g172) & (!g142) & (g883)) + ((!sk[97]) & (!g47) & (g101) & (g172) & (g142) & (g883)) + ((!sk[97]) & (g47) & (!g101) & (!g172) & (!g142) & (!g883)) + ((!sk[97]) & (g47) & (!g101) & (!g172) & (!g142) & (g883)) + ((!sk[97]) & (g47) & (!g101) & (!g172) & (g142) & (!g883)) + ((!sk[97]) & (g47) & (!g101) & (!g172) & (g142) & (g883)) + ((!sk[97]) & (g47) & (!g101) & (g172) & (!g142) & (!g883)) + ((!sk[97]) & (g47) & (!g101) & (g172) & (!g142) & (g883)) + ((!sk[97]) & (g47) & (!g101) & (g172) & (g142) & (!g883)) + ((!sk[97]) & (g47) & (!g101) & (g172) & (g142) & (g883)) + ((!sk[97]) & (g47) & (g101) & (!g172) & (!g142) & (!g883)) + ((!sk[97]) & (g47) & (g101) & (!g172) & (!g142) & (g883)) + ((!sk[97]) & (g47) & (g101) & (!g172) & (g142) & (!g883)) + ((!sk[97]) & (g47) & (g101) & (!g172) & (g142) & (g883)) + ((!sk[97]) & (g47) & (g101) & (g172) & (!g142) & (!g883)) + ((!sk[97]) & (g47) & (g101) & (g172) & (!g142) & (g883)) + ((!sk[97]) & (g47) & (g101) & (g172) & (g142) & (!g883)) + ((!sk[97]) & (g47) & (g101) & (g172) & (g142) & (g883)) + ((sk[97]) & (!g47) & (g101) & (!g172) & (!g142) & (!g883)) + ((sk[97]) & (!g47) & (g101) & (!g172) & (g142) & (!g883)) + ((sk[97]) & (!g47) & (g101) & (!g172) & (g142) & (g883)) + ((sk[97]) & (!g47) & (g101) & (g172) & (!g142) & (!g883)) + ((sk[97]) & (!g47) & (g101) & (g172) & (!g142) & (g883)) + ((sk[97]) & (!g47) & (g101) & (g172) & (g142) & (!g883)) + ((sk[97]) & (!g47) & (g101) & (g172) & (g142) & (g883)) + ((sk[97]) & (g47) & (g101) & (!g172) & (!g142) & (!g883)) + ((sk[97]) & (g47) & (g101) & (!g172) & (!g142) & (g883)) + ((sk[97]) & (g47) & (g101) & (!g172) & (g142) & (!g883)) + ((sk[97]) & (g47) & (g101) & (!g172) & (g142) & (g883)) + ((sk[97]) & (g47) & (g101) & (g172) & (!g142) & (!g883)) + ((sk[97]) & (g47) & (g101) & (g172) & (!g142) & (g883)) + ((sk[97]) & (g47) & (g101) & (g172) & (g142) & (!g883)) + ((sk[97]) & (g47) & (g101) & (g172) & (g142) & (g883)));
	assign g976 = (((!g12) & (!g101) & (!g970) & (g971) & (g974) & (!g975)) + ((!g12) & (g101) & (!g970) & (g971) & (g974) & (!g975)) + ((g12) & (!g101) & (!g970) & (g971) & (g974) & (!g975)));
	assign g977 = (((!g99) & (!g114) & (!sk[99]) & (!g560) & (!g464) & (g838)) + ((!g99) & (!g114) & (!sk[99]) & (!g560) & (g464) & (g838)) + ((!g99) & (!g114) & (!sk[99]) & (g560) & (!g464) & (g838)) + ((!g99) & (!g114) & (!sk[99]) & (g560) & (g464) & (g838)) + ((!g99) & (g114) & (!sk[99]) & (!g560) & (!g464) & (g838)) + ((!g99) & (g114) & (!sk[99]) & (!g560) & (g464) & (g838)) + ((!g99) & (g114) & (!sk[99]) & (g560) & (!g464) & (g838)) + ((!g99) & (g114) & (!sk[99]) & (g560) & (g464) & (g838)) + ((g99) & (!g114) & (!sk[99]) & (!g560) & (!g464) & (!g838)) + ((g99) & (!g114) & (!sk[99]) & (!g560) & (!g464) & (g838)) + ((g99) & (!g114) & (!sk[99]) & (!g560) & (g464) & (!g838)) + ((g99) & (!g114) & (!sk[99]) & (!g560) & (g464) & (g838)) + ((g99) & (!g114) & (!sk[99]) & (g560) & (!g464) & (!g838)) + ((g99) & (!g114) & (!sk[99]) & (g560) & (!g464) & (g838)) + ((g99) & (!g114) & (!sk[99]) & (g560) & (g464) & (!g838)) + ((g99) & (!g114) & (!sk[99]) & (g560) & (g464) & (g838)) + ((g99) & (!g114) & (sk[99]) & (!g560) & (!g464) & (!g838)) + ((g99) & (!g114) & (sk[99]) & (!g560) & (!g464) & (g838)) + ((g99) & (!g114) & (sk[99]) & (!g560) & (g464) & (!g838)) + ((g99) & (!g114) & (sk[99]) & (g560) & (!g464) & (!g838)) + ((g99) & (!g114) & (sk[99]) & (g560) & (!g464) & (g838)) + ((g99) & (!g114) & (sk[99]) & (g560) & (g464) & (!g838)) + ((g99) & (!g114) & (sk[99]) & (g560) & (g464) & (g838)) + ((g99) & (g114) & (!sk[99]) & (!g560) & (!g464) & (!g838)) + ((g99) & (g114) & (!sk[99]) & (!g560) & (!g464) & (g838)) + ((g99) & (g114) & (!sk[99]) & (!g560) & (g464) & (!g838)) + ((g99) & (g114) & (!sk[99]) & (!g560) & (g464) & (g838)) + ((g99) & (g114) & (!sk[99]) & (g560) & (!g464) & (!g838)) + ((g99) & (g114) & (!sk[99]) & (g560) & (!g464) & (g838)) + ((g99) & (g114) & (!sk[99]) & (g560) & (g464) & (!g838)) + ((g99) & (g114) & (!sk[99]) & (g560) & (g464) & (g838)) + ((g99) & (g114) & (sk[99]) & (!g560) & (!g464) & (!g838)) + ((g99) & (g114) & (sk[99]) & (!g560) & (!g464) & (g838)) + ((g99) & (g114) & (sk[99]) & (!g560) & (g464) & (!g838)) + ((g99) & (g114) & (sk[99]) & (!g560) & (g464) & (g838)) + ((g99) & (g114) & (sk[99]) & (g560) & (!g464) & (!g838)) + ((g99) & (g114) & (sk[99]) & (g560) & (!g464) & (g838)) + ((g99) & (g114) & (sk[99]) & (g560) & (g464) & (!g838)) + ((g99) & (g114) & (sk[99]) & (g560) & (g464) & (g838)));
	assign g978 = (((!g451) & (sk[100]) & (!g928) & (!g977)) + ((g451) & (!sk[100]) & (!g928) & (!g977)) + ((g451) & (!sk[100]) & (!g928) & (g977)) + ((g451) & (!sk[100]) & (g928) & (!g977)) + ((g451) & (!sk[100]) & (g928) & (g977)));
	assign g979 = (((!g630) & (sk[101]) & (!g907)) + ((g630) & (!sk[101]) & (!g907)) + ((g630) & (!sk[101]) & (g907)));
	assign g980 = (((!sk[102]) & (g193) & (!g706)) + ((!sk[102]) & (g193) & (g706)) + ((sk[102]) & (!g193) & (!g706)));
	assign g981 = (((g99) & (!sk[103]) & (!g979) & (!g980)) + ((g99) & (!sk[103]) & (!g979) & (g980)) + ((g99) & (!sk[103]) & (g979) & (!g980)) + ((g99) & (!sk[103]) & (g979) & (g980)) + ((g99) & (sk[103]) & (!g979) & (!g980)) + ((g99) & (sk[103]) & (!g979) & (g980)) + ((g99) & (sk[103]) & (g979) & (!g980)));
	assign g982 = (((!g702) & (sk[104]) & (!g881)) + ((g702) & (!sk[104]) & (!g881)) + ((g702) & (!sk[104]) & (g881)));
	assign g983 = (((!g101) & (!g193) & (!g630) & (!g706) & (!g981) & (!g982)) + ((!g101) & (!g193) & (!g630) & (!g706) & (!g981) & (g982)) + ((!g101) & (!g193) & (!g630) & (g706) & (!g981) & (!g982)) + ((!g101) & (!g193) & (!g630) & (g706) & (!g981) & (g982)) + ((!g101) & (!g193) & (g630) & (!g706) & (!g981) & (!g982)) + ((!g101) & (!g193) & (g630) & (!g706) & (!g981) & (g982)) + ((!g101) & (!g193) & (g630) & (g706) & (!g981) & (!g982)) + ((!g101) & (!g193) & (g630) & (g706) & (!g981) & (g982)) + ((!g101) & (g193) & (!g630) & (!g706) & (!g981) & (!g982)) + ((!g101) & (g193) & (!g630) & (!g706) & (!g981) & (g982)) + ((!g101) & (g193) & (!g630) & (g706) & (!g981) & (!g982)) + ((!g101) & (g193) & (!g630) & (g706) & (!g981) & (g982)) + ((!g101) & (g193) & (g630) & (!g706) & (!g981) & (!g982)) + ((!g101) & (g193) & (g630) & (!g706) & (!g981) & (g982)) + ((!g101) & (g193) & (g630) & (g706) & (!g981) & (!g982)) + ((!g101) & (g193) & (g630) & (g706) & (!g981) & (g982)) + ((g101) & (!g193) & (!g630) & (!g706) & (!g981) & (g982)));
	assign g984 = (((!g12) & (!g16) & (!sk[106]) & (!g99) & (!g101) & (g187)) + ((!g12) & (!g16) & (!sk[106]) & (!g99) & (g101) & (g187)) + ((!g12) & (!g16) & (!sk[106]) & (g99) & (!g101) & (g187)) + ((!g12) & (!g16) & (!sk[106]) & (g99) & (g101) & (g187)) + ((!g12) & (!g16) & (sk[106]) & (!g99) & (!g101) & (!g187)) + ((!g12) & (!g16) & (sk[106]) & (!g99) & (!g101) & (g187)) + ((!g12) & (!g16) & (sk[106]) & (g99) & (!g101) & (!g187)) + ((!g12) & (!g16) & (sk[106]) & (g99) & (!g101) & (g187)) + ((!g12) & (g16) & (!sk[106]) & (!g99) & (!g101) & (g187)) + ((!g12) & (g16) & (!sk[106]) & (!g99) & (g101) & (g187)) + ((!g12) & (g16) & (!sk[106]) & (g99) & (!g101) & (g187)) + ((!g12) & (g16) & (!sk[106]) & (g99) & (g101) & (g187)) + ((!g12) & (g16) & (sk[106]) & (!g99) & (!g101) & (!g187)) + ((!g12) & (g16) & (sk[106]) & (!g99) & (!g101) & (g187)) + ((!g12) & (g16) & (sk[106]) & (!g99) & (g101) & (!g187)) + ((!g12) & (g16) & (sk[106]) & (g99) & (!g101) & (!g187)) + ((!g12) & (g16) & (sk[106]) & (g99) & (!g101) & (g187)) + ((!g12) & (g16) & (sk[106]) & (g99) & (g101) & (!g187)) + ((g12) & (!g16) & (!sk[106]) & (!g99) & (!g101) & (!g187)) + ((g12) & (!g16) & (!sk[106]) & (!g99) & (!g101) & (g187)) + ((g12) & (!g16) & (!sk[106]) & (!g99) & (g101) & (!g187)) + ((g12) & (!g16) & (!sk[106]) & (!g99) & (g101) & (g187)) + ((g12) & (!g16) & (!sk[106]) & (g99) & (!g101) & (!g187)) + ((g12) & (!g16) & (!sk[106]) & (g99) & (!g101) & (g187)) + ((g12) & (!g16) & (!sk[106]) & (g99) & (g101) & (!g187)) + ((g12) & (!g16) & (!sk[106]) & (g99) & (g101) & (g187)) + ((g12) & (!g16) & (sk[106]) & (!g99) & (!g101) & (!g187)) + ((g12) & (!g16) & (sk[106]) & (!g99) & (!g101) & (g187)) + ((g12) & (g16) & (!sk[106]) & (!g99) & (!g101) & (!g187)) + ((g12) & (g16) & (!sk[106]) & (!g99) & (!g101) & (g187)) + ((g12) & (g16) & (!sk[106]) & (!g99) & (g101) & (!g187)) + ((g12) & (g16) & (!sk[106]) & (!g99) & (g101) & (g187)) + ((g12) & (g16) & (!sk[106]) & (g99) & (!g101) & (!g187)) + ((g12) & (g16) & (!sk[106]) & (g99) & (!g101) & (g187)) + ((g12) & (g16) & (!sk[106]) & (g99) & (g101) & (!g187)) + ((g12) & (g16) & (!sk[106]) & (g99) & (g101) & (g187)) + ((g12) & (g16) & (sk[106]) & (!g99) & (!g101) & (!g187)) + ((g12) & (g16) & (sk[106]) & (!g99) & (!g101) & (g187)) + ((g12) & (g16) & (sk[106]) & (!g99) & (g101) & (!g187)));
	assign g985 = (((!g101) & (!g534) & (!g899) & (g978) & (g983) & (g984)) + ((!g101) & (!g534) & (g899) & (g978) & (g983) & (g984)) + ((!g101) & (g534) & (!g899) & (g978) & (g983) & (g984)) + ((!g101) & (g534) & (g899) & (g978) & (g983) & (g984)) + ((g101) & (!g534) & (g899) & (g978) & (g983) & (g984)));
	assign g986 = (((g7) & (!sk[108]) & (!g95)) + ((g7) & (!sk[108]) & (g95)) + ((g7) & (sk[108]) & (g95)));
	assign g987 = (((!i_8_) & (!g100) & (!sk[109]) & (g522) & (g986)) + ((!i_8_) & (g100) & (!sk[109]) & (!g522) & (!g986)) + ((!i_8_) & (g100) & (!sk[109]) & (!g522) & (g986)) + ((!i_8_) & (g100) & (!sk[109]) & (g522) & (!g986)) + ((!i_8_) & (g100) & (!sk[109]) & (g522) & (g986)) + ((!i_8_) & (g100) & (sk[109]) & (!g522) & (g986)) + ((!i_8_) & (g100) & (sk[109]) & (g522) & (!g986)) + ((!i_8_) & (g100) & (sk[109]) & (g522) & (g986)) + ((i_8_) & (!g100) & (!sk[109]) & (g522) & (!g986)) + ((i_8_) & (!g100) & (!sk[109]) & (g522) & (g986)) + ((i_8_) & (g100) & (!sk[109]) & (!g522) & (!g986)) + ((i_8_) & (g100) & (!sk[109]) & (!g522) & (g986)) + ((i_8_) & (g100) & (!sk[109]) & (g522) & (!g986)) + ((i_8_) & (g100) & (!sk[109]) & (g522) & (g986)) + ((i_8_) & (g100) & (sk[109]) & (g522) & (!g986)) + ((i_8_) & (g100) & (sk[109]) & (g522) & (g986)));
	assign g988 = (((g99) & (!g835) & (!sk[110]) & (!g887)) + ((g99) & (!g835) & (!sk[110]) & (g887)) + ((g99) & (!g835) & (sk[110]) & (!g887)) + ((g99) & (!g835) & (sk[110]) & (g887)) + ((g99) & (g835) & (!sk[110]) & (!g887)) + ((g99) & (g835) & (!sk[110]) & (g887)) + ((g99) & (g835) & (sk[110]) & (!g887)));
	assign g989 = (((!sk[111]) & (!g46) & (!g66) & (!g99) & (!g209) & (g531)) + ((!sk[111]) & (!g46) & (!g66) & (!g99) & (g209) & (g531)) + ((!sk[111]) & (!g46) & (!g66) & (g99) & (!g209) & (g531)) + ((!sk[111]) & (!g46) & (!g66) & (g99) & (g209) & (g531)) + ((!sk[111]) & (!g46) & (g66) & (!g99) & (!g209) & (g531)) + ((!sk[111]) & (!g46) & (g66) & (!g99) & (g209) & (g531)) + ((!sk[111]) & (!g46) & (g66) & (g99) & (!g209) & (g531)) + ((!sk[111]) & (!g46) & (g66) & (g99) & (g209) & (g531)) + ((!sk[111]) & (g46) & (!g66) & (!g99) & (!g209) & (!g531)) + ((!sk[111]) & (g46) & (!g66) & (!g99) & (!g209) & (g531)) + ((!sk[111]) & (g46) & (!g66) & (!g99) & (g209) & (!g531)) + ((!sk[111]) & (g46) & (!g66) & (!g99) & (g209) & (g531)) + ((!sk[111]) & (g46) & (!g66) & (g99) & (!g209) & (!g531)) + ((!sk[111]) & (g46) & (!g66) & (g99) & (!g209) & (g531)) + ((!sk[111]) & (g46) & (!g66) & (g99) & (g209) & (!g531)) + ((!sk[111]) & (g46) & (!g66) & (g99) & (g209) & (g531)) + ((!sk[111]) & (g46) & (g66) & (!g99) & (!g209) & (!g531)) + ((!sk[111]) & (g46) & (g66) & (!g99) & (!g209) & (g531)) + ((!sk[111]) & (g46) & (g66) & (!g99) & (g209) & (!g531)) + ((!sk[111]) & (g46) & (g66) & (!g99) & (g209) & (g531)) + ((!sk[111]) & (g46) & (g66) & (g99) & (!g209) & (!g531)) + ((!sk[111]) & (g46) & (g66) & (g99) & (!g209) & (g531)) + ((!sk[111]) & (g46) & (g66) & (g99) & (g209) & (!g531)) + ((!sk[111]) & (g46) & (g66) & (g99) & (g209) & (g531)) + ((sk[111]) & (!g46) & (!g66) & (g99) & (!g209) & (g531)) + ((sk[111]) & (!g46) & (!g66) & (g99) & (g209) & (!g531)) + ((sk[111]) & (!g46) & (!g66) & (g99) & (g209) & (g531)) + ((sk[111]) & (!g46) & (g66) & (g99) & (!g209) & (!g531)) + ((sk[111]) & (!g46) & (g66) & (g99) & (!g209) & (g531)) + ((sk[111]) & (!g46) & (g66) & (g99) & (g209) & (!g531)) + ((sk[111]) & (!g46) & (g66) & (g99) & (g209) & (g531)) + ((sk[111]) & (g46) & (!g66) & (g99) & (!g209) & (!g531)) + ((sk[111]) & (g46) & (!g66) & (g99) & (!g209) & (g531)) + ((sk[111]) & (g46) & (!g66) & (g99) & (g209) & (!g531)) + ((sk[111]) & (g46) & (!g66) & (g99) & (g209) & (g531)) + ((sk[111]) & (g46) & (g66) & (g99) & (!g209) & (!g531)) + ((sk[111]) & (g46) & (g66) & (g99) & (!g209) & (g531)) + ((sk[111]) & (g46) & (g66) & (g99) & (g209) & (!g531)) + ((sk[111]) & (g46) & (g66) & (g99) & (g209) & (g531)));
	assign g990 = (((!g7) & (!g101) & (!g131) & (!g540) & (!g710) & (!g989)) + ((!g7) & (!g101) & (!g131) & (!g540) & (g710) & (!g989)) + ((!g7) & (!g101) & (!g131) & (g540) & (!g710) & (!g989)) + ((!g7) & (!g101) & (!g131) & (g540) & (g710) & (!g989)) + ((!g7) & (!g101) & (g131) & (!g540) & (!g710) & (!g989)) + ((!g7) & (!g101) & (g131) & (!g540) & (g710) & (!g989)) + ((!g7) & (!g101) & (g131) & (g540) & (!g710) & (!g989)) + ((!g7) & (!g101) & (g131) & (g540) & (g710) & (!g989)) + ((!g7) & (g101) & (!g131) & (!g540) & (!g710) & (!g989)) + ((!g7) & (g101) & (g131) & (!g540) & (!g710) & (!g989)) + ((g7) & (!g101) & (!g131) & (!g540) & (!g710) & (!g989)) + ((g7) & (!g101) & (!g131) & (!g540) & (g710) & (!g989)) + ((g7) & (!g101) & (!g131) & (g540) & (!g710) & (!g989)) + ((g7) & (!g101) & (!g131) & (g540) & (g710) & (!g989)) + ((g7) & (!g101) & (g131) & (!g540) & (!g710) & (!g989)) + ((g7) & (!g101) & (g131) & (!g540) & (g710) & (!g989)) + ((g7) & (!g101) & (g131) & (g540) & (!g710) & (!g989)) + ((g7) & (!g101) & (g131) & (g540) & (g710) & (!g989)) + ((g7) & (g101) & (!g131) & (!g540) & (!g710) & (!g989)));
	assign g991 = (((!i_8_) & (!g4) & (!sk[113]) & (!g98) & (!g213) & (g986)) + ((!i_8_) & (!g4) & (!sk[113]) & (!g98) & (g213) & (g986)) + ((!i_8_) & (!g4) & (!sk[113]) & (g98) & (!g213) & (g986)) + ((!i_8_) & (!g4) & (!sk[113]) & (g98) & (g213) & (g986)) + ((!i_8_) & (g4) & (!sk[113]) & (!g98) & (!g213) & (g986)) + ((!i_8_) & (g4) & (!sk[113]) & (!g98) & (g213) & (g986)) + ((!i_8_) & (g4) & (!sk[113]) & (g98) & (!g213) & (g986)) + ((!i_8_) & (g4) & (!sk[113]) & (g98) & (g213) & (g986)) + ((!i_8_) & (g4) & (sk[113]) & (g98) & (g213) & (!g986)) + ((!i_8_) & (g4) & (sk[113]) & (g98) & (g213) & (g986)) + ((i_8_) & (!g4) & (!sk[113]) & (!g98) & (!g213) & (!g986)) + ((i_8_) & (!g4) & (!sk[113]) & (!g98) & (!g213) & (g986)) + ((i_8_) & (!g4) & (!sk[113]) & (!g98) & (g213) & (!g986)) + ((i_8_) & (!g4) & (!sk[113]) & (!g98) & (g213) & (g986)) + ((i_8_) & (!g4) & (!sk[113]) & (g98) & (!g213) & (!g986)) + ((i_8_) & (!g4) & (!sk[113]) & (g98) & (!g213) & (g986)) + ((i_8_) & (!g4) & (!sk[113]) & (g98) & (g213) & (!g986)) + ((i_8_) & (!g4) & (!sk[113]) & (g98) & (g213) & (g986)) + ((i_8_) & (g4) & (!sk[113]) & (!g98) & (!g213) & (!g986)) + ((i_8_) & (g4) & (!sk[113]) & (!g98) & (!g213) & (g986)) + ((i_8_) & (g4) & (!sk[113]) & (!g98) & (g213) & (!g986)) + ((i_8_) & (g4) & (!sk[113]) & (!g98) & (g213) & (g986)) + ((i_8_) & (g4) & (!sk[113]) & (g98) & (!g213) & (!g986)) + ((i_8_) & (g4) & (!sk[113]) & (g98) & (!g213) & (g986)) + ((i_8_) & (g4) & (!sk[113]) & (g98) & (g213) & (!g986)) + ((i_8_) & (g4) & (!sk[113]) & (g98) & (g213) & (g986)) + ((i_8_) & (g4) & (sk[113]) & (g98) & (!g213) & (g986)) + ((i_8_) & (g4) & (sk[113]) & (g98) & (g213) & (!g986)) + ((i_8_) & (g4) & (sk[113]) & (g98) & (g213) & (g986)));
	assign g992 = (((!g99) & (!sk[114]) & (!g101) & (g756) & (g991)) + ((!g99) & (!sk[114]) & (g101) & (!g756) & (!g991)) + ((!g99) & (!sk[114]) & (g101) & (!g756) & (g991)) + ((!g99) & (!sk[114]) & (g101) & (g756) & (!g991)) + ((!g99) & (!sk[114]) & (g101) & (g756) & (g991)) + ((!g99) & (sk[114]) & (!g101) & (!g756) & (!g991)) + ((!g99) & (sk[114]) & (!g101) & (g756) & (!g991)) + ((!g99) & (sk[114]) & (g101) & (!g756) & (!g991)) + ((g99) & (!sk[114]) & (!g101) & (g756) & (!g991)) + ((g99) & (!sk[114]) & (!g101) & (g756) & (g991)) + ((g99) & (!sk[114]) & (g101) & (!g756) & (!g991)) + ((g99) & (!sk[114]) & (g101) & (!g756) & (g991)) + ((g99) & (!sk[114]) & (g101) & (g756) & (!g991)) + ((g99) & (!sk[114]) & (g101) & (g756) & (g991)) + ((g99) & (sk[114]) & (!g101) & (!g756) & (!g991)) + ((g99) & (sk[114]) & (g101) & (!g756) & (!g991)));
	assign g993 = (((!sk[115]) & (!g101) & (!g183) & (g704) & (g895)) + ((!sk[115]) & (!g101) & (g183) & (!g704) & (!g895)) + ((!sk[115]) & (!g101) & (g183) & (!g704) & (g895)) + ((!sk[115]) & (!g101) & (g183) & (g704) & (!g895)) + ((!sk[115]) & (!g101) & (g183) & (g704) & (g895)) + ((!sk[115]) & (g101) & (!g183) & (g704) & (!g895)) + ((!sk[115]) & (g101) & (!g183) & (g704) & (g895)) + ((!sk[115]) & (g101) & (g183) & (!g704) & (!g895)) + ((!sk[115]) & (g101) & (g183) & (!g704) & (g895)) + ((!sk[115]) & (g101) & (g183) & (g704) & (!g895)) + ((!sk[115]) & (g101) & (g183) & (g704) & (g895)) + ((sk[115]) & (g101) & (!g183) & (!g704) & (g895)) + ((sk[115]) & (g101) & (!g183) & (g704) & (!g895)) + ((sk[115]) & (g101) & (!g183) & (g704) & (g895)) + ((sk[115]) & (g101) & (g183) & (!g704) & (!g895)) + ((sk[115]) & (g101) & (g183) & (!g704) & (g895)) + ((sk[115]) & (g101) & (g183) & (g704) & (!g895)) + ((sk[115]) & (g101) & (g183) & (g704) & (g895)));
	assign g994 = (((!g987) & (!g988) & (!g990) & (!sk[116]) & (!g992) & (g993)) + ((!g987) & (!g988) & (!g990) & (!sk[116]) & (g992) & (g993)) + ((!g987) & (!g988) & (g990) & (!sk[116]) & (!g992) & (g993)) + ((!g987) & (!g988) & (g990) & (!sk[116]) & (g992) & (g993)) + ((!g987) & (!g988) & (g990) & (sk[116]) & (g992) & (!g993)) + ((!g987) & (g988) & (!g990) & (!sk[116]) & (!g992) & (g993)) + ((!g987) & (g988) & (!g990) & (!sk[116]) & (g992) & (g993)) + ((!g987) & (g988) & (g990) & (!sk[116]) & (!g992) & (g993)) + ((!g987) & (g988) & (g990) & (!sk[116]) & (g992) & (g993)) + ((g987) & (!g988) & (!g990) & (!sk[116]) & (!g992) & (!g993)) + ((g987) & (!g988) & (!g990) & (!sk[116]) & (!g992) & (g993)) + ((g987) & (!g988) & (!g990) & (!sk[116]) & (g992) & (!g993)) + ((g987) & (!g988) & (!g990) & (!sk[116]) & (g992) & (g993)) + ((g987) & (!g988) & (g990) & (!sk[116]) & (!g992) & (!g993)) + ((g987) & (!g988) & (g990) & (!sk[116]) & (!g992) & (g993)) + ((g987) & (!g988) & (g990) & (!sk[116]) & (g992) & (!g993)) + ((g987) & (!g988) & (g990) & (!sk[116]) & (g992) & (g993)) + ((g987) & (g988) & (!g990) & (!sk[116]) & (!g992) & (!g993)) + ((g987) & (g988) & (!g990) & (!sk[116]) & (!g992) & (g993)) + ((g987) & (g988) & (!g990) & (!sk[116]) & (g992) & (!g993)) + ((g987) & (g988) & (!g990) & (!sk[116]) & (g992) & (g993)) + ((g987) & (g988) & (g990) & (!sk[116]) & (!g992) & (!g993)) + ((g987) & (g988) & (g990) & (!sk[116]) & (!g992) & (g993)) + ((g987) & (g988) & (g990) & (!sk[116]) & (g992) & (!g993)) + ((g987) & (g988) & (g990) & (!sk[116]) & (g992) & (g993)));
	assign g995 = (((!i_8_) & (g4) & (!g44) & (g98) & (!g530) & (g641)) + ((!i_8_) & (g4) & (!g44) & (g98) & (g530) & (!g641)) + ((!i_8_) & (g4) & (!g44) & (g98) & (g530) & (g641)) + ((!i_8_) & (g4) & (g44) & (g98) & (!g530) & (!g641)) + ((!i_8_) & (g4) & (g44) & (g98) & (!g530) & (g641)) + ((!i_8_) & (g4) & (g44) & (g98) & (g530) & (!g641)) + ((!i_8_) & (g4) & (g44) & (g98) & (g530) & (g641)) + ((i_8_) & (g4) & (!g44) & (g98) & (!g530) & (g641)) + ((i_8_) & (g4) & (!g44) & (g98) & (g530) & (g641)) + ((i_8_) & (g4) & (g44) & (g98) & (!g530) & (!g641)) + ((i_8_) & (g4) & (g44) & (g98) & (!g530) & (g641)) + ((i_8_) & (g4) & (g44) & (g98) & (g530) & (!g641)) + ((i_8_) & (g4) & (g44) & (g98) & (g530) & (g641)));
	assign g996 = (((!g4) & (!g43) & (!sk[118]) & (!g98) & (!g191) & (g995)) + ((!g4) & (!g43) & (!sk[118]) & (!g98) & (g191) & (g995)) + ((!g4) & (!g43) & (!sk[118]) & (g98) & (!g191) & (g995)) + ((!g4) & (!g43) & (!sk[118]) & (g98) & (g191) & (g995)) + ((!g4) & (!g43) & (sk[118]) & (!g98) & (!g191) & (!g995)) + ((!g4) & (!g43) & (sk[118]) & (!g98) & (g191) & (!g995)) + ((!g4) & (!g43) & (sk[118]) & (g98) & (!g191) & (!g995)) + ((!g4) & (!g43) & (sk[118]) & (g98) & (g191) & (!g995)) + ((!g4) & (g43) & (!sk[118]) & (!g98) & (!g191) & (g995)) + ((!g4) & (g43) & (!sk[118]) & (!g98) & (g191) & (g995)) + ((!g4) & (g43) & (!sk[118]) & (g98) & (!g191) & (g995)) + ((!g4) & (g43) & (!sk[118]) & (g98) & (g191) & (g995)) + ((!g4) & (g43) & (sk[118]) & (!g98) & (!g191) & (!g995)) + ((!g4) & (g43) & (sk[118]) & (!g98) & (g191) & (!g995)) + ((!g4) & (g43) & (sk[118]) & (g98) & (!g191) & (!g995)) + ((!g4) & (g43) & (sk[118]) & (g98) & (g191) & (!g995)) + ((g4) & (!g43) & (!sk[118]) & (!g98) & (!g191) & (!g995)) + ((g4) & (!g43) & (!sk[118]) & (!g98) & (!g191) & (g995)) + ((g4) & (!g43) & (!sk[118]) & (!g98) & (g191) & (!g995)) + ((g4) & (!g43) & (!sk[118]) & (!g98) & (g191) & (g995)) + ((g4) & (!g43) & (!sk[118]) & (g98) & (!g191) & (!g995)) + ((g4) & (!g43) & (!sk[118]) & (g98) & (!g191) & (g995)) + ((g4) & (!g43) & (!sk[118]) & (g98) & (g191) & (!g995)) + ((g4) & (!g43) & (!sk[118]) & (g98) & (g191) & (g995)) + ((g4) & (!g43) & (sk[118]) & (!g98) & (!g191) & (!g995)) + ((g4) & (!g43) & (sk[118]) & (!g98) & (g191) & (!g995)) + ((g4) & (!g43) & (sk[118]) & (g98) & (!g191) & (!g995)) + ((g4) & (g43) & (!sk[118]) & (!g98) & (!g191) & (!g995)) + ((g4) & (g43) & (!sk[118]) & (!g98) & (!g191) & (g995)) + ((g4) & (g43) & (!sk[118]) & (!g98) & (g191) & (!g995)) + ((g4) & (g43) & (!sk[118]) & (!g98) & (g191) & (g995)) + ((g4) & (g43) & (!sk[118]) & (g98) & (!g191) & (!g995)) + ((g4) & (g43) & (!sk[118]) & (g98) & (!g191) & (g995)) + ((g4) & (g43) & (!sk[118]) & (g98) & (g191) & (!g995)) + ((g4) & (g43) & (!sk[118]) & (g98) & (g191) & (g995)) + ((g4) & (g43) & (sk[118]) & (!g98) & (!g191) & (!g995)) + ((g4) & (g43) & (sk[118]) & (!g98) & (g191) & (!g995)));
	assign g997 = (((!g99) & (!g101) & (!sk[119]) & (!g187) & (!g534) & (g907)) + ((!g99) & (!g101) & (!sk[119]) & (!g187) & (g534) & (g907)) + ((!g99) & (!g101) & (!sk[119]) & (g187) & (!g534) & (g907)) + ((!g99) & (!g101) & (!sk[119]) & (g187) & (g534) & (g907)) + ((!g99) & (!g101) & (sk[119]) & (!g187) & (!g534) & (!g907)) + ((!g99) & (!g101) & (sk[119]) & (!g187) & (!g534) & (g907)) + ((!g99) & (!g101) & (sk[119]) & (!g187) & (g534) & (!g907)) + ((!g99) & (!g101) & (sk[119]) & (!g187) & (g534) & (g907)) + ((!g99) & (!g101) & (sk[119]) & (g187) & (!g534) & (!g907)) + ((!g99) & (!g101) & (sk[119]) & (g187) & (!g534) & (g907)) + ((!g99) & (!g101) & (sk[119]) & (g187) & (g534) & (!g907)) + ((!g99) & (!g101) & (sk[119]) & (g187) & (g534) & (g907)) + ((!g99) & (g101) & (!sk[119]) & (!g187) & (!g534) & (g907)) + ((!g99) & (g101) & (!sk[119]) & (!g187) & (g534) & (g907)) + ((!g99) & (g101) & (!sk[119]) & (g187) & (!g534) & (g907)) + ((!g99) & (g101) & (!sk[119]) & (g187) & (g534) & (g907)) + ((!g99) & (g101) & (sk[119]) & (!g187) & (!g534) & (!g907)) + ((!g99) & (g101) & (sk[119]) & (!g187) & (g534) & (!g907)) + ((!g99) & (g101) & (sk[119]) & (g187) & (!g534) & (!g907)) + ((!g99) & (g101) & (sk[119]) & (g187) & (g534) & (!g907)) + ((g99) & (!g101) & (!sk[119]) & (!g187) & (!g534) & (!g907)) + ((g99) & (!g101) & (!sk[119]) & (!g187) & (!g534) & (g907)) + ((g99) & (!g101) & (!sk[119]) & (!g187) & (g534) & (!g907)) + ((g99) & (!g101) & (!sk[119]) & (!g187) & (g534) & (g907)) + ((g99) & (!g101) & (!sk[119]) & (g187) & (!g534) & (!g907)) + ((g99) & (!g101) & (!sk[119]) & (g187) & (!g534) & (g907)) + ((g99) & (!g101) & (!sk[119]) & (g187) & (g534) & (!g907)) + ((g99) & (!g101) & (!sk[119]) & (g187) & (g534) & (g907)) + ((g99) & (!g101) & (sk[119]) & (!g187) & (!g534) & (!g907)) + ((g99) & (!g101) & (sk[119]) & (!g187) & (!g534) & (g907)) + ((g99) & (g101) & (!sk[119]) & (!g187) & (!g534) & (!g907)) + ((g99) & (g101) & (!sk[119]) & (!g187) & (!g534) & (g907)) + ((g99) & (g101) & (!sk[119]) & (!g187) & (g534) & (!g907)) + ((g99) & (g101) & (!sk[119]) & (!g187) & (g534) & (g907)) + ((g99) & (g101) & (!sk[119]) & (g187) & (!g534) & (!g907)) + ((g99) & (g101) & (!sk[119]) & (g187) & (!g534) & (g907)) + ((g99) & (g101) & (!sk[119]) & (g187) & (g534) & (!g907)) + ((g99) & (g101) & (!sk[119]) & (g187) & (g534) & (g907)) + ((g99) & (g101) & (sk[119]) & (!g187) & (!g534) & (!g907)));
	assign g998 = (((!g99) & (!sk[120]) & (!g201) & (g702) & (g881)) + ((!g99) & (!sk[120]) & (g201) & (!g702) & (!g881)) + ((!g99) & (!sk[120]) & (g201) & (!g702) & (g881)) + ((!g99) & (!sk[120]) & (g201) & (g702) & (!g881)) + ((!g99) & (!sk[120]) & (g201) & (g702) & (g881)) + ((g99) & (!sk[120]) & (!g201) & (g702) & (!g881)) + ((g99) & (!sk[120]) & (!g201) & (g702) & (g881)) + ((g99) & (!sk[120]) & (g201) & (!g702) & (!g881)) + ((g99) & (!sk[120]) & (g201) & (!g702) & (g881)) + ((g99) & (!sk[120]) & (g201) & (g702) & (!g881)) + ((g99) & (!sk[120]) & (g201) & (g702) & (g881)) + ((g99) & (sk[120]) & (!g201) & (!g702) & (!g881)) + ((g99) & (sk[120]) & (!g201) & (!g702) & (g881)) + ((g99) & (sk[120]) & (!g201) & (g702) & (!g881)) + ((g99) & (sk[120]) & (!g201) & (g702) & (g881)) + ((g99) & (sk[120]) & (g201) & (!g702) & (g881)) + ((g99) & (sk[120]) & (g201) & (g702) & (!g881)) + ((g99) & (sk[120]) & (g201) & (g702) & (g881)));
	assign g999 = (((!sk[121]) & (g996) & (!g997) & (!g998)) + ((!sk[121]) & (g996) & (!g997) & (g998)) + ((!sk[121]) & (g996) & (g997) & (!g998)) + ((!sk[121]) & (g996) & (g997) & (g998)) + ((sk[121]) & (g996) & (g997) & (!g998)));
	assign g1000 = (((!g976) & (!g985) & (g994) & (!sk[122]) & (g999)) + ((!g976) & (g985) & (!g994) & (!sk[122]) & (!g999)) + ((!g976) & (g985) & (!g994) & (!sk[122]) & (g999)) + ((!g976) & (g985) & (g994) & (!sk[122]) & (!g999)) + ((!g976) & (g985) & (g994) & (!sk[122]) & (g999)) + ((g976) & (!g985) & (g994) & (!sk[122]) & (!g999)) + ((g976) & (!g985) & (g994) & (!sk[122]) & (g999)) + ((g976) & (g985) & (!g994) & (!sk[122]) & (!g999)) + ((g976) & (g985) & (!g994) & (!sk[122]) & (g999)) + ((g976) & (g985) & (g994) & (!sk[122]) & (!g999)) + ((g976) & (g985) & (g994) & (!sk[122]) & (g999)) + ((g976) & (g985) & (g994) & (sk[122]) & (g999)));
	assign g1001 = (((!g46) & (sk[123]) & (!g209) & (!g531)) + ((g46) & (!sk[123]) & (!g209) & (!g531)) + ((g46) & (!sk[123]) & (!g209) & (g531)) + ((g46) & (!sk[123]) & (g209) & (!g531)) + ((g46) & (!sk[123]) & (g209) & (g531)));
	assign g1002 = (((!i_14_) & (!i_12_) & (i_13_) & (g99) & (g95) & (!g93)) + ((!i_14_) & (!i_12_) & (i_13_) & (g99) & (g95) & (g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (g99) & (g95) & (!g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (g99) & (g95) & (g93)) + ((!i_14_) & (i_12_) & (i_13_) & (g99) & (g95) & (!g93)) + ((!i_14_) & (i_12_) & (i_13_) & (g99) & (g95) & (g93)) + ((i_14_) & (!i_12_) & (!i_13_) & (g99) & (!g95) & (!g93)) + ((i_14_) & (!i_12_) & (!i_13_) & (g99) & (g95) & (!g93)) + ((i_14_) & (!i_12_) & (i_13_) & (g99) & (!g95) & (!g93)) + ((i_14_) & (!i_12_) & (i_13_) & (g99) & (g95) & (!g93)) + ((i_14_) & (i_12_) & (!i_13_) & (g99) & (!g95) & (!g93)) + ((i_14_) & (i_12_) & (!i_13_) & (g99) & (g95) & (!g93)));
	assign g1003 = (((!g99) & (!g268) & (!sk[125]) & (!g96) & (!g669) & (g818)) + ((!g99) & (!g268) & (!sk[125]) & (!g96) & (g669) & (g818)) + ((!g99) & (!g268) & (!sk[125]) & (g96) & (!g669) & (g818)) + ((!g99) & (!g268) & (!sk[125]) & (g96) & (g669) & (g818)) + ((!g99) & (g268) & (!sk[125]) & (!g96) & (!g669) & (g818)) + ((!g99) & (g268) & (!sk[125]) & (!g96) & (g669) & (g818)) + ((!g99) & (g268) & (!sk[125]) & (g96) & (!g669) & (g818)) + ((!g99) & (g268) & (!sk[125]) & (g96) & (g669) & (g818)) + ((g99) & (!g268) & (!sk[125]) & (!g96) & (!g669) & (!g818)) + ((g99) & (!g268) & (!sk[125]) & (!g96) & (!g669) & (g818)) + ((g99) & (!g268) & (!sk[125]) & (!g96) & (g669) & (!g818)) + ((g99) & (!g268) & (!sk[125]) & (!g96) & (g669) & (g818)) + ((g99) & (!g268) & (!sk[125]) & (g96) & (!g669) & (!g818)) + ((g99) & (!g268) & (!sk[125]) & (g96) & (!g669) & (g818)) + ((g99) & (!g268) & (!sk[125]) & (g96) & (g669) & (!g818)) + ((g99) & (!g268) & (!sk[125]) & (g96) & (g669) & (g818)) + ((g99) & (!g268) & (sk[125]) & (!g96) & (!g669) & (!g818)) + ((g99) & (!g268) & (sk[125]) & (!g96) & (!g669) & (g818)) + ((g99) & (!g268) & (sk[125]) & (!g96) & (g669) & (!g818)) + ((g99) & (!g268) & (sk[125]) & (!g96) & (g669) & (g818)) + ((g99) & (!g268) & (sk[125]) & (g96) & (!g669) & (!g818)) + ((g99) & (!g268) & (sk[125]) & (g96) & (!g669) & (g818)) + ((g99) & (!g268) & (sk[125]) & (g96) & (g669) & (!g818)) + ((g99) & (g268) & (!sk[125]) & (!g96) & (!g669) & (!g818)) + ((g99) & (g268) & (!sk[125]) & (!g96) & (!g669) & (g818)) + ((g99) & (g268) & (!sk[125]) & (!g96) & (g669) & (!g818)) + ((g99) & (g268) & (!sk[125]) & (!g96) & (g669) & (g818)) + ((g99) & (g268) & (!sk[125]) & (g96) & (!g669) & (!g818)) + ((g99) & (g268) & (!sk[125]) & (g96) & (!g669) & (g818)) + ((g99) & (g268) & (!sk[125]) & (g96) & (g669) & (!g818)) + ((g99) & (g268) & (!sk[125]) & (g96) & (g669) & (g818)) + ((g99) & (g268) & (sk[125]) & (!g96) & (!g669) & (!g818)) + ((g99) & (g268) & (sk[125]) & (!g96) & (!g669) & (g818)) + ((g99) & (g268) & (sk[125]) & (!g96) & (g669) & (!g818)) + ((g99) & (g268) & (sk[125]) & (!g96) & (g669) & (g818)) + ((g99) & (g268) & (sk[125]) & (g96) & (!g669) & (!g818)) + ((g99) & (g268) & (sk[125]) & (g96) & (!g669) & (g818)) + ((g99) & (g268) & (sk[125]) & (g96) & (g669) & (!g818)) + ((g99) & (g268) & (sk[125]) & (g96) & (g669) & (g818)));
	assign g1004 = (((i_14_) & (!i_12_) & (!i_13_) & (!g95) & (g101) & (!g93)) + ((i_14_) & (!i_12_) & (!i_13_) & (g95) & (g101) & (!g93)) + ((i_14_) & (!i_12_) & (!i_13_) & (g95) & (g101) & (g93)) + ((i_14_) & (!i_12_) & (i_13_) & (!g95) & (g101) & (!g93)) + ((i_14_) & (!i_12_) & (i_13_) & (g95) & (g101) & (!g93)) + ((i_14_) & (!i_12_) & (i_13_) & (g95) & (g101) & (g93)) + ((i_14_) & (i_12_) & (!i_13_) & (!g95) & (g101) & (!g93)) + ((i_14_) & (i_12_) & (!i_13_) & (g95) & (g101) & (!g93)) + ((i_14_) & (i_12_) & (i_13_) & (g95) & (g101) & (!g93)) + ((i_14_) & (i_12_) & (i_13_) & (g95) & (g101) & (g93)));
	assign g1005 = (((!g101) & (!sk[127]) & (!g94) & (!g475) & (!g678) & (g891)) + ((!g101) & (!sk[127]) & (!g94) & (!g475) & (g678) & (g891)) + ((!g101) & (!sk[127]) & (!g94) & (g475) & (!g678) & (g891)) + ((!g101) & (!sk[127]) & (!g94) & (g475) & (g678) & (g891)) + ((!g101) & (!sk[127]) & (g94) & (!g475) & (!g678) & (g891)) + ((!g101) & (!sk[127]) & (g94) & (!g475) & (g678) & (g891)) + ((!g101) & (!sk[127]) & (g94) & (g475) & (!g678) & (g891)) + ((!g101) & (!sk[127]) & (g94) & (g475) & (g678) & (g891)) + ((g101) & (!sk[127]) & (!g94) & (!g475) & (!g678) & (!g891)) + ((g101) & (!sk[127]) & (!g94) & (!g475) & (!g678) & (g891)) + ((g101) & (!sk[127]) & (!g94) & (!g475) & (g678) & (!g891)) + ((g101) & (!sk[127]) & (!g94) & (!g475) & (g678) & (g891)) + ((g101) & (!sk[127]) & (!g94) & (g475) & (!g678) & (!g891)) + ((g101) & (!sk[127]) & (!g94) & (g475) & (!g678) & (g891)) + ((g101) & (!sk[127]) & (!g94) & (g475) & (g678) & (!g891)) + ((g101) & (!sk[127]) & (!g94) & (g475) & (g678) & (g891)) + ((g101) & (!sk[127]) & (g94) & (!g475) & (!g678) & (!g891)) + ((g101) & (!sk[127]) & (g94) & (!g475) & (!g678) & (g891)) + ((g101) & (!sk[127]) & (g94) & (!g475) & (g678) & (!g891)) + ((g101) & (!sk[127]) & (g94) & (!g475) & (g678) & (g891)) + ((g101) & (!sk[127]) & (g94) & (g475) & (!g678) & (!g891)) + ((g101) & (!sk[127]) & (g94) & (g475) & (!g678) & (g891)) + ((g101) & (!sk[127]) & (g94) & (g475) & (g678) & (!g891)) + ((g101) & (!sk[127]) & (g94) & (g475) & (g678) & (g891)) + ((g101) & (sk[127]) & (!g94) & (!g475) & (!g678) & (!g891)) + ((g101) & (sk[127]) & (!g94) & (!g475) & (!g678) & (g891)) + ((g101) & (sk[127]) & (!g94) & (!g475) & (g678) & (!g891)) + ((g101) & (sk[127]) & (!g94) & (!g475) & (g678) & (g891)) + ((g101) & (sk[127]) & (!g94) & (g475) & (!g678) & (!g891)) + ((g101) & (sk[127]) & (!g94) & (g475) & (!g678) & (g891)) + ((g101) & (sk[127]) & (!g94) & (g475) & (g678) & (!g891)) + ((g101) & (sk[127]) & (g94) & (!g475) & (!g678) & (!g891)) + ((g101) & (sk[127]) & (g94) & (!g475) & (!g678) & (g891)) + ((g101) & (sk[127]) & (g94) & (!g475) & (g678) & (!g891)) + ((g101) & (sk[127]) & (g94) & (!g475) & (g678) & (g891)) + ((g101) & (sk[127]) & (g94) & (g475) & (!g678) & (!g891)) + ((g101) & (sk[127]) & (g94) & (g475) & (!g678) & (g891)) + ((g101) & (sk[127]) & (g94) & (g475) & (g678) & (!g891)) + ((g101) & (sk[127]) & (g94) & (g475) & (g678) & (g891)));
	assign g1006 = (((!g1002) & (!g1003) & (!sk[0]) & (g1004) & (g1005)) + ((!g1002) & (!g1003) & (sk[0]) & (!g1004) & (!g1005)) + ((!g1002) & (g1003) & (!sk[0]) & (!g1004) & (!g1005)) + ((!g1002) & (g1003) & (!sk[0]) & (!g1004) & (g1005)) + ((!g1002) & (g1003) & (!sk[0]) & (g1004) & (!g1005)) + ((!g1002) & (g1003) & (!sk[0]) & (g1004) & (g1005)) + ((g1002) & (!g1003) & (!sk[0]) & (g1004) & (!g1005)) + ((g1002) & (!g1003) & (!sk[0]) & (g1004) & (g1005)) + ((g1002) & (g1003) & (!sk[0]) & (!g1004) & (!g1005)) + ((g1002) & (g1003) & (!sk[0]) & (!g1004) & (g1005)) + ((g1002) & (g1003) & (!sk[0]) & (g1004) & (!g1005)) + ((g1002) & (g1003) & (!sk[0]) & (g1004) & (g1005)));
	assign g1007 = (((!i_9_) & (!i_8_) & (!sk[1]) & (!g30) & (!g326) & (g98)) + ((!i_9_) & (!i_8_) & (!sk[1]) & (!g30) & (g326) & (g98)) + ((!i_9_) & (!i_8_) & (!sk[1]) & (g30) & (!g326) & (g98)) + ((!i_9_) & (!i_8_) & (!sk[1]) & (g30) & (g326) & (g98)) + ((!i_9_) & (i_8_) & (!sk[1]) & (!g30) & (!g326) & (g98)) + ((!i_9_) & (i_8_) & (!sk[1]) & (!g30) & (g326) & (g98)) + ((!i_9_) & (i_8_) & (!sk[1]) & (g30) & (!g326) & (g98)) + ((!i_9_) & (i_8_) & (!sk[1]) & (g30) & (g326) & (g98)) + ((!i_9_) & (i_8_) & (sk[1]) & (g30) & (g326) & (g98)) + ((i_9_) & (!i_8_) & (!sk[1]) & (!g30) & (!g326) & (!g98)) + ((i_9_) & (!i_8_) & (!sk[1]) & (!g30) & (!g326) & (g98)) + ((i_9_) & (!i_8_) & (!sk[1]) & (!g30) & (g326) & (!g98)) + ((i_9_) & (!i_8_) & (!sk[1]) & (!g30) & (g326) & (g98)) + ((i_9_) & (!i_8_) & (!sk[1]) & (g30) & (!g326) & (!g98)) + ((i_9_) & (!i_8_) & (!sk[1]) & (g30) & (!g326) & (g98)) + ((i_9_) & (!i_8_) & (!sk[1]) & (g30) & (g326) & (!g98)) + ((i_9_) & (!i_8_) & (!sk[1]) & (g30) & (g326) & (g98)) + ((i_9_) & (!i_8_) & (sk[1]) & (g30) & (g326) & (g98)) + ((i_9_) & (i_8_) & (!sk[1]) & (!g30) & (!g326) & (!g98)) + ((i_9_) & (i_8_) & (!sk[1]) & (!g30) & (!g326) & (g98)) + ((i_9_) & (i_8_) & (!sk[1]) & (!g30) & (g326) & (!g98)) + ((i_9_) & (i_8_) & (!sk[1]) & (!g30) & (g326) & (g98)) + ((i_9_) & (i_8_) & (!sk[1]) & (g30) & (!g326) & (!g98)) + ((i_9_) & (i_8_) & (!sk[1]) & (g30) & (!g326) & (g98)) + ((i_9_) & (i_8_) & (!sk[1]) & (g30) & (g326) & (!g98)) + ((i_9_) & (i_8_) & (!sk[1]) & (g30) & (g326) & (g98)));
	assign g1008 = (((!g101) & (!sk[2]) & (!g1001) & (g1006) & (g1007)) + ((!g101) & (!sk[2]) & (g1001) & (!g1006) & (!g1007)) + ((!g101) & (!sk[2]) & (g1001) & (!g1006) & (g1007)) + ((!g101) & (!sk[2]) & (g1001) & (g1006) & (!g1007)) + ((!g101) & (!sk[2]) & (g1001) & (g1006) & (g1007)) + ((!g101) & (sk[2]) & (!g1001) & (g1006) & (!g1007)) + ((!g101) & (sk[2]) & (g1001) & (g1006) & (!g1007)) + ((g101) & (!sk[2]) & (!g1001) & (g1006) & (!g1007)) + ((g101) & (!sk[2]) & (!g1001) & (g1006) & (g1007)) + ((g101) & (!sk[2]) & (g1001) & (!g1006) & (!g1007)) + ((g101) & (!sk[2]) & (g1001) & (!g1006) & (g1007)) + ((g101) & (!sk[2]) & (g1001) & (g1006) & (!g1007)) + ((g101) & (!sk[2]) & (g1001) & (g1006) & (g1007)) + ((g101) & (sk[2]) & (g1001) & (g1006) & (!g1007)));
	assign g1009 = (((!sk[3]) & (!g99) & (!g264) & (!g115) & (!g711) & (g672)) + ((!sk[3]) & (!g99) & (!g264) & (!g115) & (g711) & (g672)) + ((!sk[3]) & (!g99) & (!g264) & (g115) & (!g711) & (g672)) + ((!sk[3]) & (!g99) & (!g264) & (g115) & (g711) & (g672)) + ((!sk[3]) & (!g99) & (g264) & (!g115) & (!g711) & (g672)) + ((!sk[3]) & (!g99) & (g264) & (!g115) & (g711) & (g672)) + ((!sk[3]) & (!g99) & (g264) & (g115) & (!g711) & (g672)) + ((!sk[3]) & (!g99) & (g264) & (g115) & (g711) & (g672)) + ((!sk[3]) & (g99) & (!g264) & (!g115) & (!g711) & (!g672)) + ((!sk[3]) & (g99) & (!g264) & (!g115) & (!g711) & (g672)) + ((!sk[3]) & (g99) & (!g264) & (!g115) & (g711) & (!g672)) + ((!sk[3]) & (g99) & (!g264) & (!g115) & (g711) & (g672)) + ((!sk[3]) & (g99) & (!g264) & (g115) & (!g711) & (!g672)) + ((!sk[3]) & (g99) & (!g264) & (g115) & (!g711) & (g672)) + ((!sk[3]) & (g99) & (!g264) & (g115) & (g711) & (!g672)) + ((!sk[3]) & (g99) & (!g264) & (g115) & (g711) & (g672)) + ((!sk[3]) & (g99) & (g264) & (!g115) & (!g711) & (!g672)) + ((!sk[3]) & (g99) & (g264) & (!g115) & (!g711) & (g672)) + ((!sk[3]) & (g99) & (g264) & (!g115) & (g711) & (!g672)) + ((!sk[3]) & (g99) & (g264) & (!g115) & (g711) & (g672)) + ((!sk[3]) & (g99) & (g264) & (g115) & (!g711) & (!g672)) + ((!sk[3]) & (g99) & (g264) & (g115) & (!g711) & (g672)) + ((!sk[3]) & (g99) & (g264) & (g115) & (g711) & (!g672)) + ((!sk[3]) & (g99) & (g264) & (g115) & (g711) & (g672)) + ((sk[3]) & (g99) & (!g264) & (!g115) & (!g711) & (g672)) + ((sk[3]) & (g99) & (!g264) & (!g115) & (g711) & (!g672)) + ((sk[3]) & (g99) & (!g264) & (!g115) & (g711) & (g672)) + ((sk[3]) & (g99) & (!g264) & (g115) & (!g711) & (g672)) + ((sk[3]) & (g99) & (!g264) & (g115) & (g711) & (g672)) + ((sk[3]) & (g99) & (g264) & (!g115) & (!g711) & (!g672)) + ((sk[3]) & (g99) & (g264) & (!g115) & (!g711) & (g672)) + ((sk[3]) & (g99) & (g264) & (!g115) & (g711) & (!g672)) + ((sk[3]) & (g99) & (g264) & (!g115) & (g711) & (g672)) + ((sk[3]) & (g99) & (g264) & (g115) & (!g711) & (!g672)) + ((sk[3]) & (g99) & (g264) & (g115) & (!g711) & (g672)) + ((sk[3]) & (g99) & (g264) & (g115) & (g711) & (!g672)) + ((sk[3]) & (g99) & (g264) & (g115) & (g711) & (g672)));
	assign g1010 = (((!g101) & (!g696) & (!sk[4]) & (g672) & (g1009)) + ((!g101) & (!g696) & (sk[4]) & (!g672) & (!g1009)) + ((!g101) & (!g696) & (sk[4]) & (g672) & (!g1009)) + ((!g101) & (g696) & (!sk[4]) & (!g672) & (!g1009)) + ((!g101) & (g696) & (!sk[4]) & (!g672) & (g1009)) + ((!g101) & (g696) & (!sk[4]) & (g672) & (!g1009)) + ((!g101) & (g696) & (!sk[4]) & (g672) & (g1009)) + ((!g101) & (g696) & (sk[4]) & (!g672) & (!g1009)) + ((!g101) & (g696) & (sk[4]) & (g672) & (!g1009)) + ((g101) & (!g696) & (!sk[4]) & (g672) & (!g1009)) + ((g101) & (!g696) & (!sk[4]) & (g672) & (g1009)) + ((g101) & (g696) & (!sk[4]) & (!g672) & (!g1009)) + ((g101) & (g696) & (!sk[4]) & (!g672) & (g1009)) + ((g101) & (g696) & (!sk[4]) & (g672) & (!g1009)) + ((g101) & (g696) & (!sk[4]) & (g672) & (g1009)) + ((g101) & (g696) & (sk[4]) & (!g672) & (!g1009)));
	assign g1011 = (((!sk[5]) & (!g99) & (!g101) & (g696) & (g670)) + ((!sk[5]) & (!g99) & (g101) & (!g696) & (!g670)) + ((!sk[5]) & (!g99) & (g101) & (!g696) & (g670)) + ((!sk[5]) & (!g99) & (g101) & (g696) & (!g670)) + ((!sk[5]) & (!g99) & (g101) & (g696) & (g670)) + ((!sk[5]) & (g99) & (!g101) & (g696) & (!g670)) + ((!sk[5]) & (g99) & (!g101) & (g696) & (g670)) + ((!sk[5]) & (g99) & (g101) & (!g696) & (!g670)) + ((!sk[5]) & (g99) & (g101) & (!g696) & (g670)) + ((!sk[5]) & (g99) & (g101) & (g696) & (!g670)) + ((!sk[5]) & (g99) & (g101) & (g696) & (g670)) + ((sk[5]) & (!g99) & (g101) & (!g696) & (g670)) + ((sk[5]) & (!g99) & (g101) & (g696) & (g670)) + ((sk[5]) & (g99) & (!g101) & (!g696) & (!g670)) + ((sk[5]) & (g99) & (!g101) & (!g696) & (g670)) + ((sk[5]) & (g99) & (g101) & (!g696) & (!g670)) + ((sk[5]) & (g99) & (g101) & (!g696) & (g670)) + ((sk[5]) & (g99) & (g101) & (g696) & (g670)));
	assign g1012 = (((!g10) & (g99) & (!g220) & (!g221) & (!g550) & (!g544)) + ((!g10) & (g99) & (!g220) & (!g221) & (!g550) & (g544)) + ((!g10) & (g99) & (!g220) & (!g221) & (g550) & (!g544)) + ((!g10) & (g99) & (!g220) & (!g221) & (g550) & (g544)) + ((!g10) & (g99) & (!g220) & (g221) & (!g550) & (!g544)) + ((!g10) & (g99) & (!g220) & (g221) & (g550) & (!g544)) + ((!g10) & (g99) & (!g220) & (g221) & (g550) & (g544)) + ((!g10) & (g99) & (g220) & (!g221) & (!g550) & (!g544)) + ((!g10) & (g99) & (g220) & (!g221) & (!g550) & (g544)) + ((!g10) & (g99) & (g220) & (!g221) & (g550) & (!g544)) + ((!g10) & (g99) & (g220) & (!g221) & (g550) & (g544)) + ((!g10) & (g99) & (g220) & (g221) & (!g550) & (!g544)) + ((!g10) & (g99) & (g220) & (g221) & (!g550) & (g544)) + ((!g10) & (g99) & (g220) & (g221) & (g550) & (!g544)) + ((!g10) & (g99) & (g220) & (g221) & (g550) & (g544)) + ((g10) & (g99) & (!g220) & (!g221) & (!g550) & (!g544)) + ((g10) & (g99) & (!g220) & (!g221) & (!g550) & (g544)) + ((g10) & (g99) & (!g220) & (!g221) & (g550) & (!g544)) + ((g10) & (g99) & (!g220) & (!g221) & (g550) & (g544)) + ((g10) & (g99) & (!g220) & (g221) & (!g550) & (!g544)) + ((g10) & (g99) & (!g220) & (g221) & (!g550) & (g544)) + ((g10) & (g99) & (!g220) & (g221) & (g550) & (!g544)) + ((g10) & (g99) & (!g220) & (g221) & (g550) & (g544)) + ((g10) & (g99) & (g220) & (!g221) & (!g550) & (!g544)) + ((g10) & (g99) & (g220) & (!g221) & (!g550) & (g544)) + ((g10) & (g99) & (g220) & (!g221) & (g550) & (!g544)) + ((g10) & (g99) & (g220) & (!g221) & (g550) & (g544)) + ((g10) & (g99) & (g220) & (g221) & (!g550) & (!g544)) + ((g10) & (g99) & (g220) & (g221) & (!g550) & (g544)) + ((g10) & (g99) & (g220) & (g221) & (g550) & (!g544)) + ((g10) & (g99) & (g220) & (g221) & (g550) & (g544)));
	assign g1013 = (((!g10) & (!g14) & (!g101) & (!g677) & (!g903) & (!g1012)) + ((!g10) & (!g14) & (!g101) & (!g677) & (g903) & (!g1012)) + ((!g10) & (!g14) & (!g101) & (g677) & (!g903) & (!g1012)) + ((!g10) & (!g14) & (!g101) & (g677) & (g903) & (!g1012)) + ((!g10) & (!g14) & (g101) & (!g677) & (!g903) & (!g1012)) + ((!g10) & (g14) & (!g101) & (!g677) & (!g903) & (!g1012)) + ((!g10) & (g14) & (!g101) & (!g677) & (g903) & (!g1012)) + ((!g10) & (g14) & (!g101) & (g677) & (!g903) & (!g1012)) + ((!g10) & (g14) & (!g101) & (g677) & (g903) & (!g1012)) + ((g10) & (!g14) & (!g101) & (!g677) & (!g903) & (!g1012)) + ((g10) & (!g14) & (!g101) & (!g677) & (g903) & (!g1012)) + ((g10) & (!g14) & (!g101) & (g677) & (!g903) & (!g1012)) + ((g10) & (!g14) & (!g101) & (g677) & (g903) & (!g1012)) + ((g10) & (g14) & (!g101) & (!g677) & (!g903) & (!g1012)) + ((g10) & (g14) & (!g101) & (!g677) & (g903) & (!g1012)) + ((g10) & (g14) & (!g101) & (g677) & (!g903) & (!g1012)) + ((g10) & (g14) & (!g101) & (g677) & (g903) & (!g1012)));
	assign g1014 = (((!g102) & (!sk[8]) & (!g119) & (g544) & (g711)) + ((!g102) & (!sk[8]) & (g119) & (!g544) & (!g711)) + ((!g102) & (!sk[8]) & (g119) & (!g544) & (g711)) + ((!g102) & (!sk[8]) & (g119) & (g544) & (!g711)) + ((!g102) & (!sk[8]) & (g119) & (g544) & (g711)) + ((!g102) & (sk[8]) & (!g119) & (g544) & (!g711)) + ((!g102) & (sk[8]) & (g119) & (g544) & (!g711)) + ((g102) & (!sk[8]) & (!g119) & (g544) & (!g711)) + ((g102) & (!sk[8]) & (!g119) & (g544) & (g711)) + ((g102) & (!sk[8]) & (g119) & (!g544) & (!g711)) + ((g102) & (!sk[8]) & (g119) & (!g544) & (g711)) + ((g102) & (!sk[8]) & (g119) & (g544) & (!g711)) + ((g102) & (!sk[8]) & (g119) & (g544) & (g711)) + ((g102) & (sk[8]) & (!g119) & (g544) & (!g711)) + ((g102) & (sk[8]) & (!g119) & (g544) & (g711)) + ((g102) & (sk[8]) & (g119) & (g544) & (!g711)));
	assign g1015 = (((!i_8_) & (!g100) & (g551) & (!sk[9]) & (g1014)) + ((!i_8_) & (g100) & (!g551) & (!sk[9]) & (!g1014)) + ((!i_8_) & (g100) & (!g551) & (!sk[9]) & (g1014)) + ((!i_8_) & (g100) & (g551) & (!sk[9]) & (!g1014)) + ((!i_8_) & (g100) & (g551) & (!sk[9]) & (g1014)) + ((!i_8_) & (g100) & (g551) & (sk[9]) & (!g1014)) + ((!i_8_) & (g100) & (g551) & (sk[9]) & (g1014)) + ((i_8_) & (!g100) & (g551) & (!sk[9]) & (!g1014)) + ((i_8_) & (!g100) & (g551) & (!sk[9]) & (g1014)) + ((i_8_) & (g100) & (!g551) & (!sk[9]) & (!g1014)) + ((i_8_) & (g100) & (!g551) & (!sk[9]) & (g1014)) + ((i_8_) & (g100) & (!g551) & (sk[9]) & (!g1014)) + ((i_8_) & (g100) & (g551) & (!sk[9]) & (!g1014)) + ((i_8_) & (g100) & (g551) & (!sk[9]) & (g1014)) + ((i_8_) & (g100) & (g551) & (sk[9]) & (!g1014)) + ((i_8_) & (g100) & (g551) & (sk[9]) & (g1014)));
	assign g1016 = (((!g324) & (!g440) & (!sk[10]) & (g864) & (g1015)) + ((!g324) & (!g440) & (sk[10]) & (!g864) & (!g1015)) + ((!g324) & (g440) & (!sk[10]) & (!g864) & (!g1015)) + ((!g324) & (g440) & (!sk[10]) & (!g864) & (g1015)) + ((!g324) & (g440) & (!sk[10]) & (g864) & (!g1015)) + ((!g324) & (g440) & (!sk[10]) & (g864) & (g1015)) + ((g324) & (!g440) & (!sk[10]) & (g864) & (!g1015)) + ((g324) & (!g440) & (!sk[10]) & (g864) & (g1015)) + ((g324) & (g440) & (!sk[10]) & (!g864) & (!g1015)) + ((g324) & (g440) & (!sk[10]) & (!g864) & (g1015)) + ((g324) & (g440) & (!sk[10]) & (g864) & (!g1015)) + ((g324) & (g440) & (!sk[10]) & (g864) & (g1015)));
	assign g1017 = (((!g267) & (!sk[11]) & (!g714) & (!g1011) & (!g1013) & (g1016)) + ((!g267) & (!sk[11]) & (!g714) & (!g1011) & (g1013) & (g1016)) + ((!g267) & (!sk[11]) & (!g714) & (g1011) & (!g1013) & (g1016)) + ((!g267) & (!sk[11]) & (!g714) & (g1011) & (g1013) & (g1016)) + ((!g267) & (!sk[11]) & (g714) & (!g1011) & (!g1013) & (g1016)) + ((!g267) & (!sk[11]) & (g714) & (!g1011) & (g1013) & (g1016)) + ((!g267) & (!sk[11]) & (g714) & (g1011) & (!g1013) & (g1016)) + ((!g267) & (!sk[11]) & (g714) & (g1011) & (g1013) & (g1016)) + ((g267) & (!sk[11]) & (!g714) & (!g1011) & (!g1013) & (!g1016)) + ((g267) & (!sk[11]) & (!g714) & (!g1011) & (!g1013) & (g1016)) + ((g267) & (!sk[11]) & (!g714) & (!g1011) & (g1013) & (!g1016)) + ((g267) & (!sk[11]) & (!g714) & (!g1011) & (g1013) & (g1016)) + ((g267) & (!sk[11]) & (!g714) & (g1011) & (!g1013) & (!g1016)) + ((g267) & (!sk[11]) & (!g714) & (g1011) & (!g1013) & (g1016)) + ((g267) & (!sk[11]) & (!g714) & (g1011) & (g1013) & (!g1016)) + ((g267) & (!sk[11]) & (!g714) & (g1011) & (g1013) & (g1016)) + ((g267) & (!sk[11]) & (g714) & (!g1011) & (!g1013) & (!g1016)) + ((g267) & (!sk[11]) & (g714) & (!g1011) & (!g1013) & (g1016)) + ((g267) & (!sk[11]) & (g714) & (!g1011) & (g1013) & (!g1016)) + ((g267) & (!sk[11]) & (g714) & (!g1011) & (g1013) & (g1016)) + ((g267) & (!sk[11]) & (g714) & (g1011) & (!g1013) & (!g1016)) + ((g267) & (!sk[11]) & (g714) & (g1011) & (!g1013) & (g1016)) + ((g267) & (!sk[11]) & (g714) & (g1011) & (g1013) & (!g1016)) + ((g267) & (!sk[11]) & (g714) & (g1011) & (g1013) & (g1016)) + ((g267) & (sk[11]) & (!g714) & (!g1011) & (g1013) & (g1016)));
	assign g1018 = (((!g106) & (!g570) & (!g575) & (!g1010) & (!sk[12]) & (g1017)) + ((!g106) & (!g570) & (!g575) & (g1010) & (!sk[12]) & (g1017)) + ((!g106) & (!g570) & (g575) & (!g1010) & (!sk[12]) & (g1017)) + ((!g106) & (!g570) & (g575) & (g1010) & (!sk[12]) & (g1017)) + ((!g106) & (g570) & (!g575) & (!g1010) & (!sk[12]) & (g1017)) + ((!g106) & (g570) & (!g575) & (g1010) & (!sk[12]) & (g1017)) + ((!g106) & (g570) & (g575) & (!g1010) & (!sk[12]) & (g1017)) + ((!g106) & (g570) & (g575) & (g1010) & (!sk[12]) & (g1017)) + ((g106) & (!g570) & (!g575) & (!g1010) & (!sk[12]) & (!g1017)) + ((g106) & (!g570) & (!g575) & (!g1010) & (!sk[12]) & (g1017)) + ((g106) & (!g570) & (!g575) & (g1010) & (!sk[12]) & (!g1017)) + ((g106) & (!g570) & (!g575) & (g1010) & (!sk[12]) & (g1017)) + ((g106) & (!g570) & (g575) & (!g1010) & (!sk[12]) & (!g1017)) + ((g106) & (!g570) & (g575) & (!g1010) & (!sk[12]) & (g1017)) + ((g106) & (!g570) & (g575) & (g1010) & (!sk[12]) & (!g1017)) + ((g106) & (!g570) & (g575) & (g1010) & (!sk[12]) & (g1017)) + ((g106) & (!g570) & (g575) & (g1010) & (sk[12]) & (g1017)) + ((g106) & (g570) & (!g575) & (!g1010) & (!sk[12]) & (!g1017)) + ((g106) & (g570) & (!g575) & (!g1010) & (!sk[12]) & (g1017)) + ((g106) & (g570) & (!g575) & (g1010) & (!sk[12]) & (!g1017)) + ((g106) & (g570) & (!g575) & (g1010) & (!sk[12]) & (g1017)) + ((g106) & (g570) & (g575) & (!g1010) & (!sk[12]) & (!g1017)) + ((g106) & (g570) & (g575) & (!g1010) & (!sk[12]) & (g1017)) + ((g106) & (g570) & (g575) & (g1010) & (!sk[12]) & (!g1017)) + ((g106) & (g570) & (g575) & (g1010) & (!sk[12]) & (g1017)));
	assign g1019 = (((!i_8_) & (!g100) & (!sk[13]) & (!g177) & (!g114) & (g560)) + ((!i_8_) & (!g100) & (!sk[13]) & (!g177) & (g114) & (g560)) + ((!i_8_) & (!g100) & (!sk[13]) & (g177) & (!g114) & (g560)) + ((!i_8_) & (!g100) & (!sk[13]) & (g177) & (g114) & (g560)) + ((!i_8_) & (!g100) & (sk[13]) & (!g177) & (!g114) & (!g560)) + ((!i_8_) & (!g100) & (sk[13]) & (!g177) & (g114) & (!g560)) + ((!i_8_) & (!g100) & (sk[13]) & (g177) & (!g114) & (!g560)) + ((!i_8_) & (!g100) & (sk[13]) & (g177) & (g114) & (!g560)) + ((!i_8_) & (g100) & (!sk[13]) & (!g177) & (!g114) & (g560)) + ((!i_8_) & (g100) & (!sk[13]) & (!g177) & (g114) & (g560)) + ((!i_8_) & (g100) & (!sk[13]) & (g177) & (!g114) & (g560)) + ((!i_8_) & (g100) & (!sk[13]) & (g177) & (g114) & (g560)) + ((!i_8_) & (g100) & (sk[13]) & (!g177) & (!g114) & (!g560)) + ((!i_8_) & (g100) & (sk[13]) & (!g177) & (g114) & (!g560)) + ((!i_8_) & (g100) & (sk[13]) & (g177) & (!g114) & (!g560)) + ((!i_8_) & (g100) & (sk[13]) & (g177) & (g114) & (!g560)) + ((i_8_) & (!g100) & (!sk[13]) & (!g177) & (!g114) & (!g560)) + ((i_8_) & (!g100) & (!sk[13]) & (!g177) & (!g114) & (g560)) + ((i_8_) & (!g100) & (!sk[13]) & (!g177) & (g114) & (!g560)) + ((i_8_) & (!g100) & (!sk[13]) & (!g177) & (g114) & (g560)) + ((i_8_) & (!g100) & (!sk[13]) & (g177) & (!g114) & (!g560)) + ((i_8_) & (!g100) & (!sk[13]) & (g177) & (!g114) & (g560)) + ((i_8_) & (!g100) & (!sk[13]) & (g177) & (g114) & (!g560)) + ((i_8_) & (!g100) & (!sk[13]) & (g177) & (g114) & (g560)) + ((i_8_) & (!g100) & (sk[13]) & (!g177) & (!g114) & (!g560)) + ((i_8_) & (!g100) & (sk[13]) & (!g177) & (g114) & (!g560)) + ((i_8_) & (!g100) & (sk[13]) & (g177) & (!g114) & (!g560)) + ((i_8_) & (!g100) & (sk[13]) & (g177) & (g114) & (!g560)) + ((i_8_) & (g100) & (!sk[13]) & (!g177) & (!g114) & (!g560)) + ((i_8_) & (g100) & (!sk[13]) & (!g177) & (!g114) & (g560)) + ((i_8_) & (g100) & (!sk[13]) & (!g177) & (g114) & (!g560)) + ((i_8_) & (g100) & (!sk[13]) & (!g177) & (g114) & (g560)) + ((i_8_) & (g100) & (!sk[13]) & (g177) & (!g114) & (!g560)) + ((i_8_) & (g100) & (!sk[13]) & (g177) & (!g114) & (g560)) + ((i_8_) & (g100) & (!sk[13]) & (g177) & (g114) & (!g560)) + ((i_8_) & (g100) & (!sk[13]) & (g177) & (g114) & (g560)) + ((i_8_) & (g100) & (sk[13]) & (!g177) & (!g114) & (!g560)));
	assign g1020 = (((!sk[14]) & (g101) & (!g1019)) + ((!sk[14]) & (g101) & (g1019)) + ((sk[14]) & (g101) & (!g1019)));
	assign g1021 = (((!g99) & (!g101) & (!g226) & (!g464) & (!g703) & (!g908)) + ((!g99) & (!g101) & (!g226) & (!g464) & (!g703) & (g908)) + ((!g99) & (!g101) & (!g226) & (!g464) & (g703) & (!g908)) + ((!g99) & (!g101) & (!g226) & (!g464) & (g703) & (g908)) + ((!g99) & (!g101) & (!g226) & (g464) & (!g703) & (!g908)) + ((!g99) & (!g101) & (!g226) & (g464) & (!g703) & (g908)) + ((!g99) & (!g101) & (!g226) & (g464) & (g703) & (!g908)) + ((!g99) & (!g101) & (!g226) & (g464) & (g703) & (g908)) + ((!g99) & (!g101) & (g226) & (!g464) & (!g703) & (!g908)) + ((!g99) & (!g101) & (g226) & (!g464) & (!g703) & (g908)) + ((!g99) & (!g101) & (g226) & (!g464) & (g703) & (!g908)) + ((!g99) & (!g101) & (g226) & (!g464) & (g703) & (g908)) + ((!g99) & (!g101) & (g226) & (g464) & (!g703) & (!g908)) + ((!g99) & (!g101) & (g226) & (g464) & (!g703) & (g908)) + ((!g99) & (!g101) & (g226) & (g464) & (g703) & (!g908)) + ((!g99) & (!g101) & (g226) & (g464) & (g703) & (g908)) + ((!g99) & (g101) & (g226) & (g464) & (!g703) & (!g908)) + ((g99) & (!g101) & (!g226) & (!g464) & (!g703) & (!g908)) + ((g99) & (!g101) & (!g226) & (g464) & (!g703) & (!g908)) + ((g99) & (!g101) & (g226) & (!g464) & (!g703) & (!g908)) + ((g99) & (!g101) & (g226) & (g464) & (!g703) & (!g908)) + ((g99) & (g101) & (g226) & (g464) & (!g703) & (!g908)));
	assign g1022 = (((!i_14_) & (!i_12_) & (i_13_) & (g99) & (!g119) & (!g122)) + ((!i_14_) & (!i_12_) & (i_13_) & (g99) & (g119) & (!g122)) + ((!i_14_) & (!i_12_) & (i_13_) & (g99) & (g119) & (g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (g99) & (!g119) & (!g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (g99) & (g119) & (!g122)) + ((i_14_) & (!i_12_) & (i_13_) & (g99) & (!g119) & (!g122)) + ((i_14_) & (!i_12_) & (i_13_) & (g99) & (g119) & (!g122)) + ((i_14_) & (!i_12_) & (i_13_) & (g99) & (g119) & (g122)) + ((i_14_) & (i_12_) & (!i_13_) & (g99) & (!g119) & (!g122)) + ((i_14_) & (i_12_) & (!i_13_) & (g99) & (g119) & (!g122)) + ((i_14_) & (i_12_) & (!i_13_) & (g99) & (g119) & (g122)) + ((i_14_) & (i_12_) & (i_13_) & (g99) & (!g119) & (!g122)) + ((i_14_) & (i_12_) & (i_13_) & (g99) & (g119) & (!g122)) + ((i_14_) & (i_12_) & (i_13_) & (g99) & (g119) & (g122)));
	assign g1023 = (((!g99) & (sk[17]) & (!g535) & (!g1022)) + ((!g99) & (sk[17]) & (g535) & (!g1022)) + ((g99) & (!sk[17]) & (!g535) & (!g1022)) + ((g99) & (!sk[17]) & (!g535) & (g1022)) + ((g99) & (!sk[17]) & (g535) & (!g1022)) + ((g99) & (!sk[17]) & (g535) & (g1022)) + ((g99) & (sk[17]) & (g535) & (!g1022)));
	assign g1024 = (((!g14) & (!g99) & (!sk[18]) & (!g197) & (!g90) & (g895)) + ((!g14) & (!g99) & (!sk[18]) & (!g197) & (g90) & (g895)) + ((!g14) & (!g99) & (!sk[18]) & (g197) & (!g90) & (g895)) + ((!g14) & (!g99) & (!sk[18]) & (g197) & (g90) & (g895)) + ((!g14) & (g99) & (!sk[18]) & (!g197) & (!g90) & (g895)) + ((!g14) & (g99) & (!sk[18]) & (!g197) & (g90) & (g895)) + ((!g14) & (g99) & (!sk[18]) & (g197) & (!g90) & (g895)) + ((!g14) & (g99) & (!sk[18]) & (g197) & (g90) & (g895)) + ((!g14) & (g99) & (sk[18]) & (!g197) & (!g90) & (!g895)) + ((!g14) & (g99) & (sk[18]) & (!g197) & (!g90) & (g895)) + ((!g14) & (g99) & (sk[18]) & (!g197) & (g90) & (g895)) + ((!g14) & (g99) & (sk[18]) & (g197) & (!g90) & (!g895)) + ((!g14) & (g99) & (sk[18]) & (g197) & (!g90) & (g895)) + ((!g14) & (g99) & (sk[18]) & (g197) & (g90) & (!g895)) + ((!g14) & (g99) & (sk[18]) & (g197) & (g90) & (g895)) + ((g14) & (!g99) & (!sk[18]) & (!g197) & (!g90) & (!g895)) + ((g14) & (!g99) & (!sk[18]) & (!g197) & (!g90) & (g895)) + ((g14) & (!g99) & (!sk[18]) & (!g197) & (g90) & (!g895)) + ((g14) & (!g99) & (!sk[18]) & (!g197) & (g90) & (g895)) + ((g14) & (!g99) & (!sk[18]) & (g197) & (!g90) & (!g895)) + ((g14) & (!g99) & (!sk[18]) & (g197) & (!g90) & (g895)) + ((g14) & (!g99) & (!sk[18]) & (g197) & (g90) & (!g895)) + ((g14) & (!g99) & (!sk[18]) & (g197) & (g90) & (g895)) + ((g14) & (g99) & (!sk[18]) & (!g197) & (!g90) & (!g895)) + ((g14) & (g99) & (!sk[18]) & (!g197) & (!g90) & (g895)) + ((g14) & (g99) & (!sk[18]) & (!g197) & (g90) & (!g895)) + ((g14) & (g99) & (!sk[18]) & (!g197) & (g90) & (g895)) + ((g14) & (g99) & (!sk[18]) & (g197) & (!g90) & (!g895)) + ((g14) & (g99) & (!sk[18]) & (g197) & (!g90) & (g895)) + ((g14) & (g99) & (!sk[18]) & (g197) & (g90) & (!g895)) + ((g14) & (g99) & (!sk[18]) & (g197) & (g90) & (g895)) + ((g14) & (g99) & (sk[18]) & (!g197) & (!g90) & (!g895)) + ((g14) & (g99) & (sk[18]) & (!g197) & (!g90) & (g895)) + ((g14) & (g99) & (sk[18]) & (!g197) & (g90) & (!g895)) + ((g14) & (g99) & (sk[18]) & (!g197) & (g90) & (g895)) + ((g14) & (g99) & (sk[18]) & (g197) & (!g90) & (!g895)) + ((g14) & (g99) & (sk[18]) & (g197) & (!g90) & (g895)) + ((g14) & (g99) & (sk[18]) & (g197) & (g90) & (!g895)) + ((g14) & (g99) & (sk[18]) & (g197) & (g90) & (g895)));
	assign g1025 = (((!g101) & (!g201) & (!g530) & (sk[19]) & (!g1024)) + ((!g101) & (!g201) & (g530) & (!sk[19]) & (g1024)) + ((!g101) & (!g201) & (g530) & (sk[19]) & (!g1024)) + ((!g101) & (g201) & (!g530) & (!sk[19]) & (!g1024)) + ((!g101) & (g201) & (!g530) & (!sk[19]) & (g1024)) + ((!g101) & (g201) & (!g530) & (sk[19]) & (!g1024)) + ((!g101) & (g201) & (g530) & (!sk[19]) & (!g1024)) + ((!g101) & (g201) & (g530) & (!sk[19]) & (g1024)) + ((!g101) & (g201) & (g530) & (sk[19]) & (!g1024)) + ((g101) & (!g201) & (g530) & (!sk[19]) & (!g1024)) + ((g101) & (!g201) & (g530) & (!sk[19]) & (g1024)) + ((g101) & (g201) & (!g530) & (!sk[19]) & (!g1024)) + ((g101) & (g201) & (!g530) & (!sk[19]) & (g1024)) + ((g101) & (g201) & (!g530) & (sk[19]) & (!g1024)) + ((g101) & (g201) & (g530) & (!sk[19]) & (!g1024)) + ((g101) & (g201) & (g530) & (!sk[19]) & (g1024)));
	assign g1026 = (((!g7) & (!g131) & (!g171) & (sk[20]) & (g158)) + ((!g7) & (!g131) & (g171) & (!sk[20]) & (g158)) + ((!g7) & (g131) & (!g171) & (!sk[20]) & (!g158)) + ((!g7) & (g131) & (!g171) & (!sk[20]) & (g158)) + ((!g7) & (g131) & (!g171) & (sk[20]) & (g158)) + ((!g7) & (g131) & (g171) & (!sk[20]) & (!g158)) + ((!g7) & (g131) & (g171) & (!sk[20]) & (g158)) + ((g7) & (!g131) & (!g171) & (sk[20]) & (g158)) + ((g7) & (!g131) & (g171) & (!sk[20]) & (!g158)) + ((g7) & (!g131) & (g171) & (!sk[20]) & (g158)) + ((g7) & (g131) & (!g171) & (!sk[20]) & (!g158)) + ((g7) & (g131) & (!g171) & (!sk[20]) & (g158)) + ((g7) & (g131) & (!g171) & (sk[20]) & (!g158)) + ((g7) & (g131) & (!g171) & (sk[20]) & (g158)) + ((g7) & (g131) & (g171) & (!sk[20]) & (!g158)) + ((g7) & (g131) & (g171) & (!sk[20]) & (g158)) + ((g7) & (g131) & (g171) & (sk[20]) & (!g158)) + ((g7) & (g131) & (g171) & (sk[20]) & (g158)));
	assign g1027 = (((i_8_) & (!g66) & (g100) & (!g253) & (!g132) & (!g279)) + ((i_8_) & (!g66) & (g100) & (!g253) & (!g132) & (g279)) + ((i_8_) & (!g66) & (g100) & (!g253) & (g132) & (g279)) + ((i_8_) & (!g66) & (g100) & (g253) & (!g132) & (!g279)) + ((i_8_) & (!g66) & (g100) & (g253) & (!g132) & (g279)) + ((i_8_) & (!g66) & (g100) & (g253) & (g132) & (!g279)) + ((i_8_) & (!g66) & (g100) & (g253) & (g132) & (g279)) + ((i_8_) & (g66) & (g100) & (!g253) & (!g132) & (!g279)) + ((i_8_) & (g66) & (g100) & (!g253) & (!g132) & (g279)) + ((i_8_) & (g66) & (g100) & (!g253) & (g132) & (!g279)) + ((i_8_) & (g66) & (g100) & (!g253) & (g132) & (g279)) + ((i_8_) & (g66) & (g100) & (g253) & (!g132) & (!g279)) + ((i_8_) & (g66) & (g100) & (g253) & (!g132) & (g279)) + ((i_8_) & (g66) & (g100) & (g253) & (g132) & (!g279)) + ((i_8_) & (g66) & (g100) & (g253) & (g132) & (g279)));
	assign g1028 = (((!g648) & (!g1020) & (g1021) & (g1023) & (g1025) & (g1542)));
	assign g1029 = (((!sk[23]) & (!g73) & (!g1000) & (!g1008) & (!g1018) & (g1028)) + ((!sk[23]) & (!g73) & (!g1000) & (!g1008) & (g1018) & (g1028)) + ((!sk[23]) & (!g73) & (!g1000) & (g1008) & (!g1018) & (g1028)) + ((!sk[23]) & (!g73) & (!g1000) & (g1008) & (g1018) & (g1028)) + ((!sk[23]) & (!g73) & (g1000) & (!g1008) & (!g1018) & (g1028)) + ((!sk[23]) & (!g73) & (g1000) & (!g1008) & (g1018) & (g1028)) + ((!sk[23]) & (!g73) & (g1000) & (g1008) & (!g1018) & (g1028)) + ((!sk[23]) & (!g73) & (g1000) & (g1008) & (g1018) & (g1028)) + ((!sk[23]) & (g73) & (!g1000) & (!g1008) & (!g1018) & (!g1028)) + ((!sk[23]) & (g73) & (!g1000) & (!g1008) & (!g1018) & (g1028)) + ((!sk[23]) & (g73) & (!g1000) & (!g1008) & (g1018) & (!g1028)) + ((!sk[23]) & (g73) & (!g1000) & (!g1008) & (g1018) & (g1028)) + ((!sk[23]) & (g73) & (!g1000) & (g1008) & (!g1018) & (!g1028)) + ((!sk[23]) & (g73) & (!g1000) & (g1008) & (!g1018) & (g1028)) + ((!sk[23]) & (g73) & (!g1000) & (g1008) & (g1018) & (!g1028)) + ((!sk[23]) & (g73) & (!g1000) & (g1008) & (g1018) & (g1028)) + ((!sk[23]) & (g73) & (g1000) & (!g1008) & (!g1018) & (!g1028)) + ((!sk[23]) & (g73) & (g1000) & (!g1008) & (!g1018) & (g1028)) + ((!sk[23]) & (g73) & (g1000) & (!g1008) & (g1018) & (!g1028)) + ((!sk[23]) & (g73) & (g1000) & (!g1008) & (g1018) & (g1028)) + ((!sk[23]) & (g73) & (g1000) & (g1008) & (!g1018) & (!g1028)) + ((!sk[23]) & (g73) & (g1000) & (g1008) & (!g1018) & (g1028)) + ((!sk[23]) & (g73) & (g1000) & (g1008) & (g1018) & (!g1028)) + ((!sk[23]) & (g73) & (g1000) & (g1008) & (g1018) & (g1028)) + ((sk[23]) & (!g73) & (!g1000) & (!g1008) & (!g1018) & (!g1028)) + ((sk[23]) & (!g73) & (!g1000) & (!g1008) & (!g1018) & (g1028)) + ((sk[23]) & (!g73) & (!g1000) & (!g1008) & (g1018) & (!g1028)) + ((sk[23]) & (!g73) & (!g1000) & (!g1008) & (g1018) & (g1028)) + ((sk[23]) & (!g73) & (!g1000) & (g1008) & (!g1018) & (!g1028)) + ((sk[23]) & (!g73) & (!g1000) & (g1008) & (!g1018) & (g1028)) + ((sk[23]) & (!g73) & (!g1000) & (g1008) & (g1018) & (!g1028)) + ((sk[23]) & (!g73) & (!g1000) & (g1008) & (g1018) & (g1028)) + ((sk[23]) & (!g73) & (g1000) & (!g1008) & (!g1018) & (!g1028)) + ((sk[23]) & (!g73) & (g1000) & (!g1008) & (!g1018) & (g1028)) + ((sk[23]) & (!g73) & (g1000) & (!g1008) & (g1018) & (!g1028)) + ((sk[23]) & (!g73) & (g1000) & (!g1008) & (g1018) & (g1028)) + ((sk[23]) & (!g73) & (g1000) & (g1008) & (!g1018) & (!g1028)) + ((sk[23]) & (!g73) & (g1000) & (g1008) & (!g1018) & (g1028)) + ((sk[23]) & (!g73) & (g1000) & (g1008) & (g1018) & (!g1028)) + ((sk[23]) & (!g73) & (g1000) & (g1008) & (g1018) & (g1028)) + ((sk[23]) & (g73) & (g1000) & (g1008) & (g1018) & (g1028)));
	assign g1030 = (((!g213) & (!g557) & (!sk[24]) & (g522) & (g756)) + ((!g213) & (!g557) & (sk[24]) & (!g522) & (!g756)) + ((!g213) & (g557) & (!sk[24]) & (!g522) & (!g756)) + ((!g213) & (g557) & (!sk[24]) & (!g522) & (g756)) + ((!g213) & (g557) & (!sk[24]) & (g522) & (!g756)) + ((!g213) & (g557) & (!sk[24]) & (g522) & (g756)) + ((g213) & (!g557) & (!sk[24]) & (g522) & (!g756)) + ((g213) & (!g557) & (!sk[24]) & (g522) & (g756)) + ((g213) & (g557) & (!sk[24]) & (!g522) & (!g756)) + ((g213) & (g557) & (!sk[24]) & (!g522) & (g756)) + ((g213) & (g557) & (!sk[24]) & (g522) & (!g756)) + ((g213) & (g557) & (!sk[24]) & (g522) & (g756)));
	assign g1031 = (((!g44) & (g556) & (g544) & (!g641) & (!g876) & (g1030)));
	assign g1032 = (((!i_14_) & (!i_12_) & (!sk[26]) & (!i_13_) & (!g131) & (g158)) + ((!i_14_) & (!i_12_) & (!sk[26]) & (!i_13_) & (g131) & (g158)) + ((!i_14_) & (!i_12_) & (!sk[26]) & (i_13_) & (!g131) & (g158)) + ((!i_14_) & (!i_12_) & (!sk[26]) & (i_13_) & (g131) & (g158)) + ((!i_14_) & (!i_12_) & (sk[26]) & (!i_13_) & (!g131) & (!g158)) + ((!i_14_) & (!i_12_) & (sk[26]) & (!i_13_) & (!g131) & (g158)) + ((!i_14_) & (!i_12_) & (sk[26]) & (i_13_) & (!g131) & (!g158)) + ((!i_14_) & (i_12_) & (!sk[26]) & (!i_13_) & (!g131) & (g158)) + ((!i_14_) & (i_12_) & (!sk[26]) & (!i_13_) & (g131) & (g158)) + ((!i_14_) & (i_12_) & (!sk[26]) & (i_13_) & (!g131) & (g158)) + ((!i_14_) & (i_12_) & (!sk[26]) & (i_13_) & (g131) & (g158)) + ((!i_14_) & (i_12_) & (sk[26]) & (!i_13_) & (!g131) & (!g158)) + ((!i_14_) & (i_12_) & (sk[26]) & (!i_13_) & (!g131) & (g158)) + ((!i_14_) & (i_12_) & (sk[26]) & (i_13_) & (!g131) & (!g158)) + ((!i_14_) & (i_12_) & (sk[26]) & (i_13_) & (!g131) & (g158)) + ((i_14_) & (!i_12_) & (!sk[26]) & (!i_13_) & (!g131) & (!g158)) + ((i_14_) & (!i_12_) & (!sk[26]) & (!i_13_) & (!g131) & (g158)) + ((i_14_) & (!i_12_) & (!sk[26]) & (!i_13_) & (g131) & (!g158)) + ((i_14_) & (!i_12_) & (!sk[26]) & (!i_13_) & (g131) & (g158)) + ((i_14_) & (!i_12_) & (!sk[26]) & (i_13_) & (!g131) & (!g158)) + ((i_14_) & (!i_12_) & (!sk[26]) & (i_13_) & (!g131) & (g158)) + ((i_14_) & (!i_12_) & (!sk[26]) & (i_13_) & (g131) & (!g158)) + ((i_14_) & (!i_12_) & (!sk[26]) & (i_13_) & (g131) & (g158)) + ((i_14_) & (!i_12_) & (sk[26]) & (!i_13_) & (!g131) & (!g158)) + ((i_14_) & (!i_12_) & (sk[26]) & (!i_13_) & (g131) & (!g158)) + ((i_14_) & (!i_12_) & (sk[26]) & (i_13_) & (!g131) & (!g158)) + ((i_14_) & (!i_12_) & (sk[26]) & (i_13_) & (!g131) & (g158)) + ((i_14_) & (!i_12_) & (sk[26]) & (i_13_) & (g131) & (!g158)) + ((i_14_) & (!i_12_) & (sk[26]) & (i_13_) & (g131) & (g158)) + ((i_14_) & (i_12_) & (!sk[26]) & (!i_13_) & (!g131) & (!g158)) + ((i_14_) & (i_12_) & (!sk[26]) & (!i_13_) & (!g131) & (g158)) + ((i_14_) & (i_12_) & (!sk[26]) & (!i_13_) & (g131) & (!g158)) + ((i_14_) & (i_12_) & (!sk[26]) & (!i_13_) & (g131) & (g158)) + ((i_14_) & (i_12_) & (!sk[26]) & (i_13_) & (!g131) & (!g158)) + ((i_14_) & (i_12_) & (!sk[26]) & (i_13_) & (!g131) & (g158)) + ((i_14_) & (i_12_) & (!sk[26]) & (i_13_) & (g131) & (!g158)) + ((i_14_) & (i_12_) & (!sk[26]) & (i_13_) & (g131) & (g158)) + ((i_14_) & (i_12_) & (sk[26]) & (!i_13_) & (!g131) & (!g158)) + ((i_14_) & (i_12_) & (sk[26]) & (!i_13_) & (!g131) & (g158)) + ((i_14_) & (i_12_) & (sk[26]) & (i_13_) & (!g131) & (!g158)) + ((i_14_) & (i_12_) & (sk[26]) & (i_13_) & (g131) & (!g158)));
	assign g1033 = (((g6) & (!i_15_) & (!i_14_) & (!i_12_) & (i_13_) & (g59)) + ((g6) & (!i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g59)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g59)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (i_13_) & (g59)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (!i_13_) & (g59)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (i_13_) & (g59)) + ((g6) & (i_15_) & (!i_14_) & (!i_12_) & (!i_13_) & (g59)) + ((g6) & (i_15_) & (!i_14_) & (!i_12_) & (i_13_) & (g59)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g59)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (i_13_) & (g59)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g59)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (i_13_) & (g59)) + ((g6) & (i_15_) & (i_14_) & (i_12_) & (!i_13_) & (g59)) + ((g6) & (i_15_) & (i_14_) & (i_12_) & (i_13_) & (g59)));
	assign g1034 = (((!g18) & (!g59) & (!g142) & (!g465) & (!sk[28]) & (g726)) + ((!g18) & (!g59) & (!g142) & (g465) & (!sk[28]) & (g726)) + ((!g18) & (!g59) & (g142) & (!g465) & (!sk[28]) & (g726)) + ((!g18) & (!g59) & (g142) & (g465) & (!sk[28]) & (g726)) + ((!g18) & (g59) & (!g142) & (!g465) & (!sk[28]) & (g726)) + ((!g18) & (g59) & (!g142) & (!g465) & (sk[28]) & (!g726)) + ((!g18) & (g59) & (!g142) & (!g465) & (sk[28]) & (g726)) + ((!g18) & (g59) & (!g142) & (g465) & (!sk[28]) & (g726)) + ((!g18) & (g59) & (!g142) & (g465) & (sk[28]) & (!g726)) + ((!g18) & (g59) & (g142) & (!g465) & (!sk[28]) & (g726)) + ((!g18) & (g59) & (g142) & (!g465) & (sk[28]) & (!g726)) + ((!g18) & (g59) & (g142) & (!g465) & (sk[28]) & (g726)) + ((!g18) & (g59) & (g142) & (g465) & (!sk[28]) & (g726)) + ((!g18) & (g59) & (g142) & (g465) & (sk[28]) & (!g726)) + ((!g18) & (g59) & (g142) & (g465) & (sk[28]) & (g726)) + ((g18) & (!g59) & (!g142) & (!g465) & (!sk[28]) & (!g726)) + ((g18) & (!g59) & (!g142) & (!g465) & (!sk[28]) & (g726)) + ((g18) & (!g59) & (!g142) & (g465) & (!sk[28]) & (!g726)) + ((g18) & (!g59) & (!g142) & (g465) & (!sk[28]) & (g726)) + ((g18) & (!g59) & (g142) & (!g465) & (!sk[28]) & (!g726)) + ((g18) & (!g59) & (g142) & (!g465) & (!sk[28]) & (g726)) + ((g18) & (!g59) & (g142) & (g465) & (!sk[28]) & (!g726)) + ((g18) & (!g59) & (g142) & (g465) & (!sk[28]) & (g726)) + ((g18) & (g59) & (!g142) & (!g465) & (!sk[28]) & (!g726)) + ((g18) & (g59) & (!g142) & (!g465) & (!sk[28]) & (g726)) + ((g18) & (g59) & (!g142) & (!g465) & (sk[28]) & (!g726)) + ((g18) & (g59) & (!g142) & (!g465) & (sk[28]) & (g726)) + ((g18) & (g59) & (!g142) & (g465) & (!sk[28]) & (!g726)) + ((g18) & (g59) & (!g142) & (g465) & (!sk[28]) & (g726)) + ((g18) & (g59) & (g142) & (!g465) & (!sk[28]) & (!g726)) + ((g18) & (g59) & (g142) & (!g465) & (!sk[28]) & (g726)) + ((g18) & (g59) & (g142) & (!g465) & (sk[28]) & (!g726)) + ((g18) & (g59) & (g142) & (!g465) & (sk[28]) & (g726)) + ((g18) & (g59) & (g142) & (g465) & (!sk[28]) & (!g726)) + ((g18) & (g59) & (g142) & (g465) & (!sk[28]) & (g726)) + ((g18) & (g59) & (g142) & (g465) & (sk[28]) & (!g726)) + ((g18) & (g59) & (g142) & (g465) & (sk[28]) & (g726)));
	assign g1035 = (((!i_14_) & (!i_12_) & (i_13_) & (!g18) & (!g15) & (g59)) + ((!i_14_) & (!i_12_) & (i_13_) & (g18) & (!g15) & (g59)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g18) & (!g15) & (g59)) + ((!i_14_) & (i_12_) & (!i_13_) & (g18) & (!g15) & (g59)) + ((i_14_) & (i_12_) & (!i_13_) & (!g18) & (!g15) & (g59)) + ((i_14_) & (i_12_) & (!i_13_) & (!g18) & (g15) & (g59)) + ((i_14_) & (i_12_) & (!i_13_) & (g18) & (!g15) & (g59)) + ((i_14_) & (i_12_) & (i_13_) & (!g18) & (!g15) & (g59)) + ((i_14_) & (i_12_) & (i_13_) & (g18) & (!g15) & (g59)));
	assign g1036 = (((!i_14_) & (!i_12_) & (!i_13_) & (g59) & (!g95) & (!g93)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g59) & (g95) & (!g93)) + ((!i_14_) & (!i_12_) & (i_13_) & (g59) & (g95) & (!g93)) + ((!i_14_) & (!i_12_) & (i_13_) & (g59) & (g95) & (g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (g59) & (!g95) & (!g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (g59) & (g95) & (!g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (g59) & (g95) & (g93)) + ((!i_14_) & (i_12_) & (i_13_) & (g59) & (!g95) & (!g93)) + ((!i_14_) & (i_12_) & (i_13_) & (g59) & (g95) & (!g93)) + ((i_14_) & (!i_12_) & (!i_13_) & (g59) & (g95) & (!g93)) + ((i_14_) & (!i_12_) & (!i_13_) & (g59) & (g95) & (g93)) + ((i_14_) & (!i_12_) & (i_13_) & (g59) & (!g95) & (!g93)) + ((i_14_) & (!i_12_) & (i_13_) & (g59) & (g95) & (!g93)) + ((i_14_) & (!i_12_) & (i_13_) & (g59) & (g95) & (g93)) + ((i_14_) & (i_12_) & (!i_13_) & (g59) & (!g95) & (!g93)) + ((i_14_) & (i_12_) & (!i_13_) & (g59) & (g95) & (!g93)) + ((i_14_) & (i_12_) & (i_13_) & (g59) & (g95) & (!g93)) + ((i_14_) & (i_12_) & (i_13_) & (g59) & (g95) & (g93)));
	assign g1037 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g131) & (g158) & (g284)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g131) & (g158) & (g284)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g131) & (g158) & (g284)) + ((!i_14_) & (i_12_) & (!i_13_) & (g131) & (g158) & (g284)) + ((!i_14_) & (i_12_) & (i_13_) & (!g131) & (g158) & (g284)) + ((!i_14_) & (i_12_) & (i_13_) & (g131) & (g158) & (g284)) + ((i_14_) & (!i_12_) & (!i_13_) & (g131) & (!g158) & (g284)) + ((i_14_) & (!i_12_) & (!i_13_) & (g131) & (g158) & (g284)) + ((i_14_) & (!i_12_) & (i_13_) & (!g131) & (g158) & (g284)) + ((i_14_) & (!i_12_) & (i_13_) & (g131) & (!g158) & (g284)) + ((i_14_) & (!i_12_) & (i_13_) & (g131) & (g158) & (g284)) + ((i_14_) & (i_12_) & (!i_13_) & (!g131) & (g158) & (g284)) + ((i_14_) & (i_12_) & (!i_13_) & (g131) & (g158) & (g284)) + ((i_14_) & (i_12_) & (i_13_) & (g131) & (!g158) & (g284)) + ((i_14_) & (i_12_) & (i_13_) & (g131) & (g158) & (g284)));
	assign g1038 = (((!g1033) & (!g1034) & (!sk[32]) & (!g1035) & (!g1036) & (g1037)) + ((!g1033) & (!g1034) & (!sk[32]) & (!g1035) & (g1036) & (g1037)) + ((!g1033) & (!g1034) & (!sk[32]) & (g1035) & (!g1036) & (g1037)) + ((!g1033) & (!g1034) & (!sk[32]) & (g1035) & (g1036) & (g1037)) + ((!g1033) & (!g1034) & (sk[32]) & (!g1035) & (!g1036) & (!g1037)) + ((!g1033) & (g1034) & (!sk[32]) & (!g1035) & (!g1036) & (g1037)) + ((!g1033) & (g1034) & (!sk[32]) & (!g1035) & (g1036) & (g1037)) + ((!g1033) & (g1034) & (!sk[32]) & (g1035) & (!g1036) & (g1037)) + ((!g1033) & (g1034) & (!sk[32]) & (g1035) & (g1036) & (g1037)) + ((g1033) & (!g1034) & (!sk[32]) & (!g1035) & (!g1036) & (!g1037)) + ((g1033) & (!g1034) & (!sk[32]) & (!g1035) & (!g1036) & (g1037)) + ((g1033) & (!g1034) & (!sk[32]) & (!g1035) & (g1036) & (!g1037)) + ((g1033) & (!g1034) & (!sk[32]) & (!g1035) & (g1036) & (g1037)) + ((g1033) & (!g1034) & (!sk[32]) & (g1035) & (!g1036) & (!g1037)) + ((g1033) & (!g1034) & (!sk[32]) & (g1035) & (!g1036) & (g1037)) + ((g1033) & (!g1034) & (!sk[32]) & (g1035) & (g1036) & (!g1037)) + ((g1033) & (!g1034) & (!sk[32]) & (g1035) & (g1036) & (g1037)) + ((g1033) & (g1034) & (!sk[32]) & (!g1035) & (!g1036) & (!g1037)) + ((g1033) & (g1034) & (!sk[32]) & (!g1035) & (!g1036) & (g1037)) + ((g1033) & (g1034) & (!sk[32]) & (!g1035) & (g1036) & (!g1037)) + ((g1033) & (g1034) & (!sk[32]) & (!g1035) & (g1036) & (g1037)) + ((g1033) & (g1034) & (!sk[32]) & (g1035) & (!g1036) & (!g1037)) + ((g1033) & (g1034) & (!sk[32]) & (g1035) & (!g1036) & (g1037)) + ((g1033) & (g1034) & (!sk[32]) & (g1035) & (g1036) & (!g1037)) + ((g1033) & (g1034) & (!sk[32]) & (g1035) & (g1036) & (g1037)));
	assign g1039 = (((!i_11_) & (!i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g113)) + ((!i_11_) & (!i_15_) & (!i_14_) & (i_12_) & (i_13_) & (g113)) + ((!i_11_) & (!i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g113)) + ((!i_11_) & (!i_15_) & (i_14_) & (!i_12_) & (i_13_) & (g113)) + ((!i_11_) & (!i_15_) & (i_14_) & (i_12_) & (i_13_) & (g113)) + ((!i_11_) & (i_15_) & (!i_14_) & (!i_12_) & (!i_13_) & (g113)) + ((!i_11_) & (i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g113)) + ((!i_11_) & (i_15_) & (!i_14_) & (i_12_) & (i_13_) & (g113)) + ((!i_11_) & (i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g113)));
	assign g1040 = (((g323) & (!sk[34]) & (!g1039)) + ((g323) & (!sk[34]) & (g1039)) + ((g323) & (sk[34]) & (g1039)));
	assign g1041 = (((!g12) & (!g177) & (!g114) & (sk[35]) & (!g560)) + ((!g12) & (!g177) & (g114) & (!sk[35]) & (g560)) + ((!g12) & (g177) & (!g114) & (!sk[35]) & (!g560)) + ((!g12) & (g177) & (!g114) & (!sk[35]) & (g560)) + ((!g12) & (g177) & (g114) & (!sk[35]) & (!g560)) + ((!g12) & (g177) & (g114) & (!sk[35]) & (g560)) + ((g12) & (!g177) & (g114) & (!sk[35]) & (!g560)) + ((g12) & (!g177) & (g114) & (!sk[35]) & (g560)) + ((g12) & (g177) & (!g114) & (!sk[35]) & (!g560)) + ((g12) & (g177) & (!g114) & (!sk[35]) & (g560)) + ((g12) & (g177) & (g114) & (!sk[35]) & (!g560)) + ((g12) & (g177) & (g114) & (!sk[35]) & (g560)));
	assign g1042 = (((g323) & (!sk[36]) & (!g187) & (!g534)) + ((g323) & (!sk[36]) & (!g187) & (g534)) + ((g323) & (!sk[36]) & (g187) & (!g534)) + ((g323) & (!sk[36]) & (g187) & (g534)) + ((g323) & (sk[36]) & (!g187) & (g534)) + ((g323) & (sk[36]) & (g187) & (!g534)) + ((g323) & (sk[36]) & (g187) & (g534)));
	assign g1043 = (((!sk[37]) & (!g12) & (!g323) & (!g201) & (!g703) & (g908)) + ((!sk[37]) & (!g12) & (!g323) & (!g201) & (g703) & (g908)) + ((!sk[37]) & (!g12) & (!g323) & (g201) & (!g703) & (g908)) + ((!sk[37]) & (!g12) & (!g323) & (g201) & (g703) & (g908)) + ((!sk[37]) & (!g12) & (g323) & (!g201) & (!g703) & (g908)) + ((!sk[37]) & (!g12) & (g323) & (!g201) & (g703) & (g908)) + ((!sk[37]) & (!g12) & (g323) & (g201) & (!g703) & (g908)) + ((!sk[37]) & (!g12) & (g323) & (g201) & (g703) & (g908)) + ((!sk[37]) & (g12) & (!g323) & (!g201) & (!g703) & (!g908)) + ((!sk[37]) & (g12) & (!g323) & (!g201) & (!g703) & (g908)) + ((!sk[37]) & (g12) & (!g323) & (!g201) & (g703) & (!g908)) + ((!sk[37]) & (g12) & (!g323) & (!g201) & (g703) & (g908)) + ((!sk[37]) & (g12) & (!g323) & (g201) & (!g703) & (!g908)) + ((!sk[37]) & (g12) & (!g323) & (g201) & (!g703) & (g908)) + ((!sk[37]) & (g12) & (!g323) & (g201) & (g703) & (!g908)) + ((!sk[37]) & (g12) & (!g323) & (g201) & (g703) & (g908)) + ((!sk[37]) & (g12) & (g323) & (!g201) & (!g703) & (!g908)) + ((!sk[37]) & (g12) & (g323) & (!g201) & (!g703) & (g908)) + ((!sk[37]) & (g12) & (g323) & (!g201) & (g703) & (!g908)) + ((!sk[37]) & (g12) & (g323) & (!g201) & (g703) & (g908)) + ((!sk[37]) & (g12) & (g323) & (g201) & (!g703) & (!g908)) + ((!sk[37]) & (g12) & (g323) & (g201) & (!g703) & (g908)) + ((!sk[37]) & (g12) & (g323) & (g201) & (g703) & (!g908)) + ((!sk[37]) & (g12) & (g323) & (g201) & (g703) & (g908)) + ((sk[37]) & (!g12) & (g323) & (!g201) & (!g703) & (!g908)) + ((sk[37]) & (!g12) & (g323) & (!g201) & (!g703) & (g908)) + ((sk[37]) & (!g12) & (g323) & (!g201) & (g703) & (!g908)) + ((sk[37]) & (!g12) & (g323) & (!g201) & (g703) & (g908)) + ((sk[37]) & (!g12) & (g323) & (g201) & (!g703) & (g908)) + ((sk[37]) & (!g12) & (g323) & (g201) & (g703) & (!g908)) + ((sk[37]) & (!g12) & (g323) & (g201) & (g703) & (g908)) + ((sk[37]) & (g12) & (g323) & (!g201) & (!g703) & (!g908)) + ((sk[37]) & (g12) & (g323) & (!g201) & (!g703) & (g908)) + ((sk[37]) & (g12) & (g323) & (!g201) & (g703) & (!g908)) + ((sk[37]) & (g12) & (g323) & (!g201) & (g703) & (g908)) + ((sk[37]) & (g12) & (g323) & (g201) & (!g703) & (!g908)) + ((sk[37]) & (g12) & (g323) & (g201) & (!g703) & (g908)) + ((sk[37]) & (g12) & (g323) & (g201) & (g703) & (!g908)) + ((sk[37]) & (g12) & (g323) & (g201) & (g703) & (g908)));
	assign g1044 = (((!g423) & (!g838) & (!sk[38]) & (!g935) & (!g1042) & (g1043)) + ((!g423) & (!g838) & (!sk[38]) & (!g935) & (g1042) & (g1043)) + ((!g423) & (!g838) & (!sk[38]) & (g935) & (!g1042) & (g1043)) + ((!g423) & (!g838) & (!sk[38]) & (g935) & (g1042) & (g1043)) + ((!g423) & (!g838) & (sk[38]) & (!g935) & (!g1042) & (!g1043)) + ((!g423) & (g838) & (!sk[38]) & (!g935) & (!g1042) & (g1043)) + ((!g423) & (g838) & (!sk[38]) & (!g935) & (g1042) & (g1043)) + ((!g423) & (g838) & (!sk[38]) & (g935) & (!g1042) & (g1043)) + ((!g423) & (g838) & (!sk[38]) & (g935) & (g1042) & (g1043)) + ((!g423) & (g838) & (sk[38]) & (!g935) & (!g1042) & (!g1043)) + ((g423) & (!g838) & (!sk[38]) & (!g935) & (!g1042) & (!g1043)) + ((g423) & (!g838) & (!sk[38]) & (!g935) & (!g1042) & (g1043)) + ((g423) & (!g838) & (!sk[38]) & (!g935) & (g1042) & (!g1043)) + ((g423) & (!g838) & (!sk[38]) & (!g935) & (g1042) & (g1043)) + ((g423) & (!g838) & (!sk[38]) & (g935) & (!g1042) & (!g1043)) + ((g423) & (!g838) & (!sk[38]) & (g935) & (!g1042) & (g1043)) + ((g423) & (!g838) & (!sk[38]) & (g935) & (g1042) & (!g1043)) + ((g423) & (!g838) & (!sk[38]) & (g935) & (g1042) & (g1043)) + ((g423) & (g838) & (!sk[38]) & (!g935) & (!g1042) & (!g1043)) + ((g423) & (g838) & (!sk[38]) & (!g935) & (!g1042) & (g1043)) + ((g423) & (g838) & (!sk[38]) & (!g935) & (g1042) & (!g1043)) + ((g423) & (g838) & (!sk[38]) & (!g935) & (g1042) & (g1043)) + ((g423) & (g838) & (!sk[38]) & (g935) & (!g1042) & (!g1043)) + ((g423) & (g838) & (!sk[38]) & (g935) & (!g1042) & (g1043)) + ((g423) & (g838) & (!sk[38]) & (g935) & (g1042) & (!g1043)) + ((g423) & (g838) & (!sk[38]) & (g935) & (g1042) & (g1043)) + ((g423) & (g838) & (sk[38]) & (!g935) & (!g1042) & (!g1043)));
	assign g1045 = (((!g423) & (!g1040) & (!g1041) & (sk[39]) & (g1044)) + ((!g423) & (!g1040) & (g1041) & (!sk[39]) & (g1044)) + ((!g423) & (!g1040) & (g1041) & (sk[39]) & (g1044)) + ((!g423) & (g1040) & (!g1041) & (!sk[39]) & (!g1044)) + ((!g423) & (g1040) & (!g1041) & (!sk[39]) & (g1044)) + ((!g423) & (g1040) & (g1041) & (!sk[39]) & (!g1044)) + ((!g423) & (g1040) & (g1041) & (!sk[39]) & (g1044)) + ((g423) & (!g1040) & (g1041) & (!sk[39]) & (!g1044)) + ((g423) & (!g1040) & (g1041) & (!sk[39]) & (g1044)) + ((g423) & (!g1040) & (g1041) & (sk[39]) & (g1044)) + ((g423) & (g1040) & (!g1041) & (!sk[39]) & (!g1044)) + ((g423) & (g1040) & (!g1041) & (!sk[39]) & (g1044)) + ((g423) & (g1040) & (g1041) & (!sk[39]) & (!g1044)) + ((g423) & (g1040) & (g1041) & (!sk[39]) & (g1044)));
	assign g1046 = (((g323) & (!sk[40]) & (!g226) & (!g464)) + ((g323) & (!sk[40]) & (!g226) & (g464)) + ((g323) & (!sk[40]) & (g226) & (!g464)) + ((g323) & (!sk[40]) & (g226) & (g464)) + ((g323) & (sk[40]) & (!g226) & (!g464)) + ((g323) & (sk[40]) & (!g226) & (g464)) + ((g323) & (sk[40]) & (g226) & (!g464)));
	assign g1047 = (((!g323) & (!g224) & (!g423) & (!g467) & (!g817) & (!g1046)) + ((!g323) & (!g224) & (!g423) & (!g467) & (g817) & (!g1046)) + ((!g323) & (!g224) & (!g423) & (g467) & (!g817) & (!g1046)) + ((!g323) & (!g224) & (!g423) & (g467) & (g817) & (!g1046)) + ((!g323) & (!g224) & (g423) & (g467) & (!g817) & (!g1046)) + ((!g323) & (g224) & (!g423) & (!g467) & (!g817) & (!g1046)) + ((!g323) & (g224) & (!g423) & (!g467) & (g817) & (!g1046)) + ((!g323) & (g224) & (!g423) & (g467) & (!g817) & (!g1046)) + ((!g323) & (g224) & (!g423) & (g467) & (g817) & (!g1046)) + ((g323) & (!g224) & (!g423) & (g467) & (!g817) & (!g1046)) + ((g323) & (!g224) & (g423) & (g467) & (!g817) & (!g1046)));
	assign g1048 = (((!sk[42]) & (!i_14_) & (!i_12_) & (!i_13_) & (!g119) & (g122)) + ((!sk[42]) & (!i_14_) & (!i_12_) & (!i_13_) & (g119) & (g122)) + ((!sk[42]) & (!i_14_) & (!i_12_) & (i_13_) & (!g119) & (g122)) + ((!sk[42]) & (!i_14_) & (!i_12_) & (i_13_) & (g119) & (g122)) + ((!sk[42]) & (!i_14_) & (i_12_) & (!i_13_) & (!g119) & (g122)) + ((!sk[42]) & (!i_14_) & (i_12_) & (!i_13_) & (g119) & (g122)) + ((!sk[42]) & (!i_14_) & (i_12_) & (i_13_) & (!g119) & (g122)) + ((!sk[42]) & (!i_14_) & (i_12_) & (i_13_) & (g119) & (g122)) + ((!sk[42]) & (i_14_) & (!i_12_) & (!i_13_) & (!g119) & (!g122)) + ((!sk[42]) & (i_14_) & (!i_12_) & (!i_13_) & (!g119) & (g122)) + ((!sk[42]) & (i_14_) & (!i_12_) & (!i_13_) & (g119) & (!g122)) + ((!sk[42]) & (i_14_) & (!i_12_) & (!i_13_) & (g119) & (g122)) + ((!sk[42]) & (i_14_) & (!i_12_) & (i_13_) & (!g119) & (!g122)) + ((!sk[42]) & (i_14_) & (!i_12_) & (i_13_) & (!g119) & (g122)) + ((!sk[42]) & (i_14_) & (!i_12_) & (i_13_) & (g119) & (!g122)) + ((!sk[42]) & (i_14_) & (!i_12_) & (i_13_) & (g119) & (g122)) + ((!sk[42]) & (i_14_) & (i_12_) & (!i_13_) & (!g119) & (!g122)) + ((!sk[42]) & (i_14_) & (i_12_) & (!i_13_) & (!g119) & (g122)) + ((!sk[42]) & (i_14_) & (i_12_) & (!i_13_) & (g119) & (!g122)) + ((!sk[42]) & (i_14_) & (i_12_) & (!i_13_) & (g119) & (g122)) + ((!sk[42]) & (i_14_) & (i_12_) & (i_13_) & (!g119) & (!g122)) + ((!sk[42]) & (i_14_) & (i_12_) & (i_13_) & (!g119) & (g122)) + ((!sk[42]) & (i_14_) & (i_12_) & (i_13_) & (g119) & (!g122)) + ((!sk[42]) & (i_14_) & (i_12_) & (i_13_) & (g119) & (g122)) + ((sk[42]) & (!i_14_) & (!i_12_) & (!i_13_) & (!g119) & (!g122)) + ((sk[42]) & (!i_14_) & (!i_12_) & (!i_13_) & (g119) & (!g122)) + ((sk[42]) & (!i_14_) & (!i_12_) & (i_13_) & (g119) & (!g122)) + ((sk[42]) & (!i_14_) & (!i_12_) & (i_13_) & (g119) & (g122)) + ((sk[42]) & (!i_14_) & (i_12_) & (!i_13_) & (!g119) & (!g122)) + ((sk[42]) & (!i_14_) & (i_12_) & (!i_13_) & (g119) & (!g122)) + ((sk[42]) & (!i_14_) & (i_12_) & (!i_13_) & (g119) & (g122)) + ((sk[42]) & (!i_14_) & (i_12_) & (i_13_) & (!g119) & (!g122)) + ((sk[42]) & (!i_14_) & (i_12_) & (i_13_) & (g119) & (!g122)) + ((sk[42]) & (!i_14_) & (i_12_) & (i_13_) & (g119) & (g122)) + ((sk[42]) & (i_14_) & (!i_12_) & (!i_13_) & (g119) & (!g122)) + ((sk[42]) & (i_14_) & (!i_12_) & (!i_13_) & (g119) & (g122)));
	assign g1049 = (((!i_14_) & (!sk[43]) & (!i_12_) & (!i_13_) & (!g104) & (g124)) + ((!i_14_) & (!sk[43]) & (!i_12_) & (!i_13_) & (g104) & (g124)) + ((!i_14_) & (!sk[43]) & (!i_12_) & (i_13_) & (!g104) & (g124)) + ((!i_14_) & (!sk[43]) & (!i_12_) & (i_13_) & (g104) & (g124)) + ((!i_14_) & (!sk[43]) & (i_12_) & (!i_13_) & (!g104) & (g124)) + ((!i_14_) & (!sk[43]) & (i_12_) & (!i_13_) & (g104) & (g124)) + ((!i_14_) & (!sk[43]) & (i_12_) & (i_13_) & (!g104) & (g124)) + ((!i_14_) & (!sk[43]) & (i_12_) & (i_13_) & (g104) & (g124)) + ((!i_14_) & (sk[43]) & (i_12_) & (!i_13_) & (!g104) & (g124)) + ((!i_14_) & (sk[43]) & (i_12_) & (!i_13_) & (g104) & (g124)) + ((!i_14_) & (sk[43]) & (i_12_) & (i_13_) & (!g104) & (g124)) + ((!i_14_) & (sk[43]) & (i_12_) & (i_13_) & (g104) & (g124)) + ((i_14_) & (!sk[43]) & (!i_12_) & (!i_13_) & (!g104) & (!g124)) + ((i_14_) & (!sk[43]) & (!i_12_) & (!i_13_) & (!g104) & (g124)) + ((i_14_) & (!sk[43]) & (!i_12_) & (!i_13_) & (g104) & (!g124)) + ((i_14_) & (!sk[43]) & (!i_12_) & (!i_13_) & (g104) & (g124)) + ((i_14_) & (!sk[43]) & (!i_12_) & (i_13_) & (!g104) & (!g124)) + ((i_14_) & (!sk[43]) & (!i_12_) & (i_13_) & (!g104) & (g124)) + ((i_14_) & (!sk[43]) & (!i_12_) & (i_13_) & (g104) & (!g124)) + ((i_14_) & (!sk[43]) & (!i_12_) & (i_13_) & (g104) & (g124)) + ((i_14_) & (!sk[43]) & (i_12_) & (!i_13_) & (!g104) & (!g124)) + ((i_14_) & (!sk[43]) & (i_12_) & (!i_13_) & (!g104) & (g124)) + ((i_14_) & (!sk[43]) & (i_12_) & (!i_13_) & (g104) & (!g124)) + ((i_14_) & (!sk[43]) & (i_12_) & (!i_13_) & (g104) & (g124)) + ((i_14_) & (!sk[43]) & (i_12_) & (i_13_) & (!g104) & (!g124)) + ((i_14_) & (!sk[43]) & (i_12_) & (i_13_) & (!g104) & (g124)) + ((i_14_) & (!sk[43]) & (i_12_) & (i_13_) & (g104) & (!g124)) + ((i_14_) & (!sk[43]) & (i_12_) & (i_13_) & (g104) & (g124)) + ((i_14_) & (sk[43]) & (!i_12_) & (!i_13_) & (!g104) & (g124)) + ((i_14_) & (sk[43]) & (!i_12_) & (!i_13_) & (g104) & (!g124)) + ((i_14_) & (sk[43]) & (!i_12_) & (!i_13_) & (g104) & (g124)) + ((i_14_) & (sk[43]) & (!i_12_) & (i_13_) & (g104) & (!g124)) + ((i_14_) & (sk[43]) & (!i_12_) & (i_13_) & (g104) & (g124)) + ((i_14_) & (sk[43]) & (i_12_) & (i_13_) & (g104) & (!g124)) + ((i_14_) & (sk[43]) & (i_12_) & (i_13_) & (g104) & (g124)));
	assign g1050 = (((!g323) & (!g90) & (!sk[44]) & (!g528) & (!g921) & (g1049)) + ((!g323) & (!g90) & (!sk[44]) & (!g528) & (g921) & (g1049)) + ((!g323) & (!g90) & (!sk[44]) & (g528) & (!g921) & (g1049)) + ((!g323) & (!g90) & (!sk[44]) & (g528) & (g921) & (g1049)) + ((!g323) & (g90) & (!sk[44]) & (!g528) & (!g921) & (g1049)) + ((!g323) & (g90) & (!sk[44]) & (!g528) & (g921) & (g1049)) + ((!g323) & (g90) & (!sk[44]) & (g528) & (!g921) & (g1049)) + ((!g323) & (g90) & (!sk[44]) & (g528) & (g921) & (g1049)) + ((g323) & (!g90) & (!sk[44]) & (!g528) & (!g921) & (!g1049)) + ((g323) & (!g90) & (!sk[44]) & (!g528) & (!g921) & (g1049)) + ((g323) & (!g90) & (!sk[44]) & (!g528) & (g921) & (!g1049)) + ((g323) & (!g90) & (!sk[44]) & (!g528) & (g921) & (g1049)) + ((g323) & (!g90) & (!sk[44]) & (g528) & (!g921) & (!g1049)) + ((g323) & (!g90) & (!sk[44]) & (g528) & (!g921) & (g1049)) + ((g323) & (!g90) & (!sk[44]) & (g528) & (g921) & (!g1049)) + ((g323) & (!g90) & (!sk[44]) & (g528) & (g921) & (g1049)) + ((g323) & (!g90) & (sk[44]) & (!g528) & (!g921) & (!g1049)) + ((g323) & (!g90) & (sk[44]) & (!g528) & (!g921) & (g1049)) + ((g323) & (!g90) & (sk[44]) & (!g528) & (g921) & (!g1049)) + ((g323) & (!g90) & (sk[44]) & (!g528) & (g921) & (g1049)) + ((g323) & (!g90) & (sk[44]) & (g528) & (!g921) & (!g1049)) + ((g323) & (!g90) & (sk[44]) & (g528) & (!g921) & (g1049)) + ((g323) & (!g90) & (sk[44]) & (g528) & (g921) & (!g1049)) + ((g323) & (!g90) & (sk[44]) & (g528) & (g921) & (g1049)) + ((g323) & (g90) & (!sk[44]) & (!g528) & (!g921) & (!g1049)) + ((g323) & (g90) & (!sk[44]) & (!g528) & (!g921) & (g1049)) + ((g323) & (g90) & (!sk[44]) & (!g528) & (g921) & (!g1049)) + ((g323) & (g90) & (!sk[44]) & (!g528) & (g921) & (g1049)) + ((g323) & (g90) & (!sk[44]) & (g528) & (!g921) & (!g1049)) + ((g323) & (g90) & (!sk[44]) & (g528) & (!g921) & (g1049)) + ((g323) & (g90) & (!sk[44]) & (g528) & (g921) & (!g1049)) + ((g323) & (g90) & (!sk[44]) & (g528) & (g921) & (g1049)) + ((g323) & (g90) & (sk[44]) & (!g528) & (!g921) & (!g1049)) + ((g323) & (g90) & (sk[44]) & (!g528) & (!g921) & (g1049)) + ((g323) & (g90) & (sk[44]) & (!g528) & (g921) & (!g1049)) + ((g323) & (g90) & (sk[44]) & (!g528) & (g921) & (g1049)) + ((g323) & (g90) & (sk[44]) & (g528) & (!g921) & (!g1049)) + ((g323) & (g90) & (sk[44]) & (g528) & (!g921) & (g1049)) + ((g323) & (g90) & (sk[44]) & (g528) & (g921) & (g1049)));
	assign g1051 = (((!g423) & (!g1048) & (sk[45]) & (!g1050)) + ((!g423) & (g1048) & (sk[45]) & (!g1050)) + ((g423) & (!g1048) & (!sk[45]) & (!g1050)) + ((g423) & (!g1048) & (!sk[45]) & (g1050)) + ((g423) & (!g1048) & (sk[45]) & (!g1050)) + ((g423) & (g1048) & (!sk[45]) & (!g1050)) + ((g423) & (g1048) & (!sk[45]) & (g1050)));
	assign g1052 = (((!sk[46]) & (!i_14_) & (!i_12_) & (!i_13_) & (!g95) & (g93)) + ((!sk[46]) & (!i_14_) & (!i_12_) & (!i_13_) & (g95) & (g93)) + ((!sk[46]) & (!i_14_) & (!i_12_) & (i_13_) & (!g95) & (g93)) + ((!sk[46]) & (!i_14_) & (!i_12_) & (i_13_) & (g95) & (g93)) + ((!sk[46]) & (!i_14_) & (i_12_) & (!i_13_) & (!g95) & (g93)) + ((!sk[46]) & (!i_14_) & (i_12_) & (!i_13_) & (g95) & (g93)) + ((!sk[46]) & (!i_14_) & (i_12_) & (i_13_) & (!g95) & (g93)) + ((!sk[46]) & (!i_14_) & (i_12_) & (i_13_) & (g95) & (g93)) + ((!sk[46]) & (i_14_) & (!i_12_) & (!i_13_) & (!g95) & (!g93)) + ((!sk[46]) & (i_14_) & (!i_12_) & (!i_13_) & (!g95) & (g93)) + ((!sk[46]) & (i_14_) & (!i_12_) & (!i_13_) & (g95) & (!g93)) + ((!sk[46]) & (i_14_) & (!i_12_) & (!i_13_) & (g95) & (g93)) + ((!sk[46]) & (i_14_) & (!i_12_) & (i_13_) & (!g95) & (!g93)) + ((!sk[46]) & (i_14_) & (!i_12_) & (i_13_) & (!g95) & (g93)) + ((!sk[46]) & (i_14_) & (!i_12_) & (i_13_) & (g95) & (!g93)) + ((!sk[46]) & (i_14_) & (!i_12_) & (i_13_) & (g95) & (g93)) + ((!sk[46]) & (i_14_) & (i_12_) & (!i_13_) & (!g95) & (!g93)) + ((!sk[46]) & (i_14_) & (i_12_) & (!i_13_) & (!g95) & (g93)) + ((!sk[46]) & (i_14_) & (i_12_) & (!i_13_) & (g95) & (!g93)) + ((!sk[46]) & (i_14_) & (i_12_) & (!i_13_) & (g95) & (g93)) + ((!sk[46]) & (i_14_) & (i_12_) & (i_13_) & (!g95) & (!g93)) + ((!sk[46]) & (i_14_) & (i_12_) & (i_13_) & (!g95) & (g93)) + ((!sk[46]) & (i_14_) & (i_12_) & (i_13_) & (g95) & (!g93)) + ((!sk[46]) & (i_14_) & (i_12_) & (i_13_) & (g95) & (g93)) + ((sk[46]) & (!i_14_) & (!i_12_) & (!i_13_) & (!g95) & (g93)) + ((sk[46]) & (!i_14_) & (!i_12_) & (!i_13_) & (g95) & (g93)) + ((sk[46]) & (!i_14_) & (!i_12_) & (i_13_) & (!g95) & (!g93)) + ((sk[46]) & (!i_14_) & (!i_12_) & (i_13_) & (!g95) & (g93)) + ((sk[46]) & (!i_14_) & (i_12_) & (!i_13_) & (!g95) & (g93)) + ((sk[46]) & (!i_14_) & (i_12_) & (i_13_) & (!g95) & (g93)) + ((sk[46]) & (i_14_) & (!i_12_) & (!i_13_) & (!g95) & (g93)) + ((sk[46]) & (i_14_) & (!i_12_) & (i_13_) & (!g95) & (g93)) + ((sk[46]) & (i_14_) & (i_12_) & (!i_13_) & (!g95) & (g93)) + ((sk[46]) & (i_14_) & (i_12_) & (!i_13_) & (g95) & (g93)) + ((sk[46]) & (i_14_) & (i_12_) & (i_13_) & (!g95) & (!g93)) + ((sk[46]) & (i_14_) & (i_12_) & (i_13_) & (!g95) & (g93)));
	assign g1053 = (((!g120) & (!sk[47]) & (!g349) & (!g423) & (!g613) & (g481)) + ((!g120) & (!sk[47]) & (!g349) & (!g423) & (g613) & (g481)) + ((!g120) & (!sk[47]) & (!g349) & (g423) & (!g613) & (g481)) + ((!g120) & (!sk[47]) & (!g349) & (g423) & (g613) & (g481)) + ((!g120) & (!sk[47]) & (g349) & (!g423) & (!g613) & (g481)) + ((!g120) & (!sk[47]) & (g349) & (!g423) & (g613) & (g481)) + ((!g120) & (!sk[47]) & (g349) & (g423) & (!g613) & (g481)) + ((!g120) & (!sk[47]) & (g349) & (g423) & (g613) & (g481)) + ((!g120) & (sk[47]) & (!g349) & (g423) & (!g613) & (!g481)) + ((!g120) & (sk[47]) & (!g349) & (g423) & (!g613) & (g481)) + ((!g120) & (sk[47]) & (!g349) & (g423) & (g613) & (!g481)) + ((!g120) & (sk[47]) & (!g349) & (g423) & (g613) & (g481)) + ((!g120) & (sk[47]) & (g349) & (g423) & (!g613) & (!g481)) + ((!g120) & (sk[47]) & (g349) & (g423) & (!g613) & (g481)) + ((!g120) & (sk[47]) & (g349) & (g423) & (g613) & (!g481)) + ((!g120) & (sk[47]) & (g349) & (g423) & (g613) & (g481)) + ((g120) & (!sk[47]) & (!g349) & (!g423) & (!g613) & (!g481)) + ((g120) & (!sk[47]) & (!g349) & (!g423) & (!g613) & (g481)) + ((g120) & (!sk[47]) & (!g349) & (!g423) & (g613) & (!g481)) + ((g120) & (!sk[47]) & (!g349) & (!g423) & (g613) & (g481)) + ((g120) & (!sk[47]) & (!g349) & (g423) & (!g613) & (!g481)) + ((g120) & (!sk[47]) & (!g349) & (g423) & (!g613) & (g481)) + ((g120) & (!sk[47]) & (!g349) & (g423) & (g613) & (!g481)) + ((g120) & (!sk[47]) & (!g349) & (g423) & (g613) & (g481)) + ((g120) & (!sk[47]) & (g349) & (!g423) & (!g613) & (!g481)) + ((g120) & (!sk[47]) & (g349) & (!g423) & (!g613) & (g481)) + ((g120) & (!sk[47]) & (g349) & (!g423) & (g613) & (!g481)) + ((g120) & (!sk[47]) & (g349) & (!g423) & (g613) & (g481)) + ((g120) & (!sk[47]) & (g349) & (g423) & (!g613) & (!g481)) + ((g120) & (!sk[47]) & (g349) & (g423) & (!g613) & (g481)) + ((g120) & (!sk[47]) & (g349) & (g423) & (g613) & (!g481)) + ((g120) & (!sk[47]) & (g349) & (g423) & (g613) & (g481)) + ((g120) & (sk[47]) & (!g349) & (g423) & (!g613) & (!g481)) + ((g120) & (sk[47]) & (!g349) & (g423) & (!g613) & (g481)) + ((g120) & (sk[47]) & (!g349) & (g423) & (g613) & (!g481)) + ((g120) & (sk[47]) & (g349) & (g423) & (!g613) & (!g481)) + ((g120) & (sk[47]) & (g349) & (g423) & (!g613) & (g481)) + ((g120) & (sk[47]) & (g349) & (g423) & (g613) & (!g481)) + ((g120) & (sk[47]) & (g349) & (g423) & (g613) & (g481)));
	assign g1054 = (((!g323) & (!g835) & (sk[48]) & (!g1053)) + ((!g323) & (g835) & (sk[48]) & (!g1053)) + ((g323) & (!g835) & (!sk[48]) & (!g1053)) + ((g323) & (!g835) & (!sk[48]) & (g1053)) + ((g323) & (g835) & (!sk[48]) & (!g1053)) + ((g323) & (g835) & (!sk[48]) & (g1053)) + ((g323) & (g835) & (sk[48]) & (!g1053)));
	assign g1055 = (((!sk[49]) & (!i_14_) & (!i_12_) & (!i_13_) & (!g95) & (g93)) + ((!sk[49]) & (!i_14_) & (!i_12_) & (!i_13_) & (g95) & (g93)) + ((!sk[49]) & (!i_14_) & (!i_12_) & (i_13_) & (!g95) & (g93)) + ((!sk[49]) & (!i_14_) & (!i_12_) & (i_13_) & (g95) & (g93)) + ((!sk[49]) & (!i_14_) & (i_12_) & (!i_13_) & (!g95) & (g93)) + ((!sk[49]) & (!i_14_) & (i_12_) & (!i_13_) & (g95) & (g93)) + ((!sk[49]) & (!i_14_) & (i_12_) & (i_13_) & (!g95) & (g93)) + ((!sk[49]) & (!i_14_) & (i_12_) & (i_13_) & (g95) & (g93)) + ((!sk[49]) & (i_14_) & (!i_12_) & (!i_13_) & (!g95) & (!g93)) + ((!sk[49]) & (i_14_) & (!i_12_) & (!i_13_) & (!g95) & (g93)) + ((!sk[49]) & (i_14_) & (!i_12_) & (!i_13_) & (g95) & (!g93)) + ((!sk[49]) & (i_14_) & (!i_12_) & (!i_13_) & (g95) & (g93)) + ((!sk[49]) & (i_14_) & (!i_12_) & (i_13_) & (!g95) & (!g93)) + ((!sk[49]) & (i_14_) & (!i_12_) & (i_13_) & (!g95) & (g93)) + ((!sk[49]) & (i_14_) & (!i_12_) & (i_13_) & (g95) & (!g93)) + ((!sk[49]) & (i_14_) & (!i_12_) & (i_13_) & (g95) & (g93)) + ((!sk[49]) & (i_14_) & (i_12_) & (!i_13_) & (!g95) & (!g93)) + ((!sk[49]) & (i_14_) & (i_12_) & (!i_13_) & (!g95) & (g93)) + ((!sk[49]) & (i_14_) & (i_12_) & (!i_13_) & (g95) & (!g93)) + ((!sk[49]) & (i_14_) & (i_12_) & (!i_13_) & (g95) & (g93)) + ((!sk[49]) & (i_14_) & (i_12_) & (i_13_) & (!g95) & (!g93)) + ((!sk[49]) & (i_14_) & (i_12_) & (i_13_) & (!g95) & (g93)) + ((!sk[49]) & (i_14_) & (i_12_) & (i_13_) & (g95) & (!g93)) + ((!sk[49]) & (i_14_) & (i_12_) & (i_13_) & (g95) & (g93)) + ((sk[49]) & (!i_14_) & (!i_12_) & (!i_13_) & (!g95) & (!g93)) + ((sk[49]) & (!i_14_) & (!i_12_) & (!i_13_) & (g95) & (!g93)) + ((sk[49]) & (!i_14_) & (i_12_) & (!i_13_) & (g95) & (!g93)) + ((sk[49]) & (!i_14_) & (i_12_) & (!i_13_) & (g95) & (g93)) + ((sk[49]) & (!i_14_) & (i_12_) & (i_13_) & (g95) & (!g93)) + ((sk[49]) & (!i_14_) & (i_12_) & (i_13_) & (g95) & (g93)) + ((sk[49]) & (i_14_) & (!i_12_) & (!i_13_) & (!g95) & (!g93)) + ((sk[49]) & (i_14_) & (!i_12_) & (!i_13_) & (g95) & (!g93)) + ((sk[49]) & (i_14_) & (!i_12_) & (i_13_) & (g95) & (!g93)) + ((sk[49]) & (i_14_) & (!i_12_) & (i_13_) & (g95) & (g93)) + ((sk[49]) & (i_14_) & (i_12_) & (i_13_) & (g95) & (!g93)) + ((sk[49]) & (i_14_) & (i_12_) & (i_13_) & (g95) & (g93)));
	assign g1056 = (((!g323) & (!g678) & (!sk[50]) & (g670) & (g756)) + ((!g323) & (g678) & (!sk[50]) & (!g670) & (!g756)) + ((!g323) & (g678) & (!sk[50]) & (!g670) & (g756)) + ((!g323) & (g678) & (!sk[50]) & (g670) & (!g756)) + ((!g323) & (g678) & (!sk[50]) & (g670) & (g756)) + ((g323) & (!g678) & (!sk[50]) & (g670) & (!g756)) + ((g323) & (!g678) & (!sk[50]) & (g670) & (g756)) + ((g323) & (!g678) & (sk[50]) & (!g670) & (!g756)) + ((g323) & (!g678) & (sk[50]) & (!g670) & (g756)) + ((g323) & (!g678) & (sk[50]) & (g670) & (!g756)) + ((g323) & (!g678) & (sk[50]) & (g670) & (g756)) + ((g323) & (g678) & (!sk[50]) & (!g670) & (!g756)) + ((g323) & (g678) & (!sk[50]) & (!g670) & (g756)) + ((g323) & (g678) & (!sk[50]) & (g670) & (!g756)) + ((g323) & (g678) & (!sk[50]) & (g670) & (g756)) + ((g323) & (g678) & (sk[50]) & (!g670) & (g756)) + ((g323) & (g678) & (sk[50]) & (g670) & (!g756)) + ((g323) & (g678) & (sk[50]) & (g670) & (g756)));
	assign g1057 = (((!g323) & (!g203) & (!sk[51]) & (g213) & (g474)) + ((!g323) & (g203) & (!sk[51]) & (!g213) & (!g474)) + ((!g323) & (g203) & (!sk[51]) & (!g213) & (g474)) + ((!g323) & (g203) & (!sk[51]) & (g213) & (!g474)) + ((!g323) & (g203) & (!sk[51]) & (g213) & (g474)) + ((g323) & (!g203) & (!sk[51]) & (g213) & (!g474)) + ((g323) & (!g203) & (!sk[51]) & (g213) & (g474)) + ((g323) & (!g203) & (sk[51]) & (!g213) & (g474)) + ((g323) & (!g203) & (sk[51]) & (g213) & (!g474)) + ((g323) & (!g203) & (sk[51]) & (g213) & (g474)) + ((g323) & (g203) & (!sk[51]) & (!g213) & (!g474)) + ((g323) & (g203) & (!sk[51]) & (!g213) & (g474)) + ((g323) & (g203) & (!sk[51]) & (g213) & (!g474)) + ((g323) & (g203) & (!sk[51]) & (g213) & (g474)) + ((g323) & (g203) & (sk[51]) & (!g213) & (!g474)) + ((g323) & (g203) & (sk[51]) & (!g213) & (g474)) + ((g323) & (g203) & (sk[51]) & (g213) & (!g474)) + ((g323) & (g203) & (sk[51]) & (g213) & (g474)));
	assign g1058 = (((!g323) & (!g818) & (!g887) & (!g1055) & (!g1056) & (!g1057)) + ((!g323) & (!g818) & (!g887) & (g1055) & (!g1056) & (!g1057)) + ((!g323) & (!g818) & (g887) & (!g1055) & (!g1056) & (!g1057)) + ((!g323) & (!g818) & (g887) & (g1055) & (!g1056) & (!g1057)) + ((!g323) & (g818) & (!g887) & (!g1055) & (!g1056) & (!g1057)) + ((!g323) & (g818) & (!g887) & (g1055) & (!g1056) & (!g1057)) + ((!g323) & (g818) & (g887) & (!g1055) & (!g1056) & (!g1057)) + ((!g323) & (g818) & (g887) & (g1055) & (!g1056) & (!g1057)) + ((g323) & (g818) & (g887) & (!g1055) & (!g1056) & (!g1057)));
	assign g1059 = (((!g423) & (!g1052) & (!sk[53]) & (g1054) & (g1058)) + ((!g423) & (!g1052) & (sk[53]) & (g1054) & (g1058)) + ((!g423) & (g1052) & (!sk[53]) & (!g1054) & (!g1058)) + ((!g423) & (g1052) & (!sk[53]) & (!g1054) & (g1058)) + ((!g423) & (g1052) & (!sk[53]) & (g1054) & (!g1058)) + ((!g423) & (g1052) & (!sk[53]) & (g1054) & (g1058)) + ((!g423) & (g1052) & (sk[53]) & (g1054) & (g1058)) + ((g423) & (!g1052) & (!sk[53]) & (g1054) & (!g1058)) + ((g423) & (!g1052) & (!sk[53]) & (g1054) & (g1058)) + ((g423) & (g1052) & (!sk[53]) & (!g1054) & (!g1058)) + ((g423) & (g1052) & (!sk[53]) & (!g1054) & (g1058)) + ((g423) & (g1052) & (!sk[53]) & (g1054) & (!g1058)) + ((g423) & (g1052) & (!sk[53]) & (g1054) & (g1058)) + ((g423) & (g1052) & (sk[53]) & (g1054) & (g1058)));
	assign g1060 = (((!g6) & (!sk[54]) & (!i_15_) & (g7) & (g182)) + ((!g6) & (!sk[54]) & (i_15_) & (!g7) & (!g182)) + ((!g6) & (!sk[54]) & (i_15_) & (!g7) & (g182)) + ((!g6) & (!sk[54]) & (i_15_) & (g7) & (!g182)) + ((!g6) & (!sk[54]) & (i_15_) & (g7) & (g182)) + ((g6) & (!sk[54]) & (!i_15_) & (g7) & (!g182)) + ((g6) & (!sk[54]) & (!i_15_) & (g7) & (g182)) + ((g6) & (!sk[54]) & (i_15_) & (!g7) & (!g182)) + ((g6) & (!sk[54]) & (i_15_) & (!g7) & (g182)) + ((g6) & (!sk[54]) & (i_15_) & (g7) & (!g182)) + ((g6) & (!sk[54]) & (i_15_) & (g7) & (g182)) + ((g6) & (sk[54]) & (!i_15_) & (!g7) & (g182)) + ((g6) & (sk[54]) & (!i_15_) & (g7) & (!g182)) + ((g6) & (sk[54]) & (!i_15_) & (g7) & (g182)));
	assign g1061 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g131) & (!sk[55]) & (g158)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g131) & (!sk[55]) & (g158)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g131) & (sk[55]) & (!g158)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g131) & (sk[55]) & (g158)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g131) & (!sk[55]) & (g158)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g131) & (sk[55]) & (g158)) + ((!i_14_) & (!i_12_) & (i_13_) & (g131) & (!sk[55]) & (g158)) + ((!i_14_) & (!i_12_) & (i_13_) & (g131) & (sk[55]) & (g158)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g131) & (!sk[55]) & (g158)) + ((!i_14_) & (i_12_) & (!i_13_) & (g131) & (!sk[55]) & (g158)) + ((!i_14_) & (i_12_) & (i_13_) & (!g131) & (!sk[55]) & (g158)) + ((!i_14_) & (i_12_) & (i_13_) & (g131) & (!sk[55]) & (g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g131) & (!sk[55]) & (!g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g131) & (!sk[55]) & (g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (g131) & (!sk[55]) & (!g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (g131) & (!sk[55]) & (g158)) + ((i_14_) & (!i_12_) & (i_13_) & (!g131) & (!sk[55]) & (!g158)) + ((i_14_) & (!i_12_) & (i_13_) & (!g131) & (!sk[55]) & (g158)) + ((i_14_) & (!i_12_) & (i_13_) & (!g131) & (sk[55]) & (g158)) + ((i_14_) & (!i_12_) & (i_13_) & (g131) & (!sk[55]) & (!g158)) + ((i_14_) & (!i_12_) & (i_13_) & (g131) & (!sk[55]) & (g158)) + ((i_14_) & (!i_12_) & (i_13_) & (g131) & (sk[55]) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (!g131) & (!sk[55]) & (!g158)) + ((i_14_) & (i_12_) & (!i_13_) & (!g131) & (!sk[55]) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (!g131) & (sk[55]) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (g131) & (!sk[55]) & (!g158)) + ((i_14_) & (i_12_) & (!i_13_) & (g131) & (!sk[55]) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (g131) & (sk[55]) & (!g158)) + ((i_14_) & (i_12_) & (!i_13_) & (g131) & (sk[55]) & (g158)) + ((i_14_) & (i_12_) & (i_13_) & (!g131) & (!sk[55]) & (!g158)) + ((i_14_) & (i_12_) & (i_13_) & (!g131) & (!sk[55]) & (g158)) + ((i_14_) & (i_12_) & (i_13_) & (!g131) & (sk[55]) & (g158)) + ((i_14_) & (i_12_) & (i_13_) & (g131) & (!sk[55]) & (!g158)) + ((i_14_) & (i_12_) & (i_13_) & (g131) & (!sk[55]) & (g158)) + ((i_14_) & (i_12_) & (i_13_) & (g131) & (sk[55]) & (g158)));
	assign g1062 = (((!g46) & (!sk[56]) & (!g642) & (!g522) & (!g896) & (g1061)) + ((!g46) & (!sk[56]) & (!g642) & (!g522) & (g896) & (g1061)) + ((!g46) & (!sk[56]) & (!g642) & (g522) & (!g896) & (g1061)) + ((!g46) & (!sk[56]) & (!g642) & (g522) & (g896) & (g1061)) + ((!g46) & (!sk[56]) & (g642) & (!g522) & (!g896) & (g1061)) + ((!g46) & (!sk[56]) & (g642) & (!g522) & (g896) & (g1061)) + ((!g46) & (!sk[56]) & (g642) & (g522) & (!g896) & (g1061)) + ((!g46) & (!sk[56]) & (g642) & (g522) & (g896) & (g1061)) + ((!g46) & (sk[56]) & (g642) & (!g522) & (!g896) & (!g1061)) + ((g46) & (!sk[56]) & (!g642) & (!g522) & (!g896) & (!g1061)) + ((g46) & (!sk[56]) & (!g642) & (!g522) & (!g896) & (g1061)) + ((g46) & (!sk[56]) & (!g642) & (!g522) & (g896) & (!g1061)) + ((g46) & (!sk[56]) & (!g642) & (!g522) & (g896) & (g1061)) + ((g46) & (!sk[56]) & (!g642) & (g522) & (!g896) & (!g1061)) + ((g46) & (!sk[56]) & (!g642) & (g522) & (!g896) & (g1061)) + ((g46) & (!sk[56]) & (!g642) & (g522) & (g896) & (!g1061)) + ((g46) & (!sk[56]) & (!g642) & (g522) & (g896) & (g1061)) + ((g46) & (!sk[56]) & (g642) & (!g522) & (!g896) & (!g1061)) + ((g46) & (!sk[56]) & (g642) & (!g522) & (!g896) & (g1061)) + ((g46) & (!sk[56]) & (g642) & (!g522) & (g896) & (!g1061)) + ((g46) & (!sk[56]) & (g642) & (!g522) & (g896) & (g1061)) + ((g46) & (!sk[56]) & (g642) & (g522) & (!g896) & (!g1061)) + ((g46) & (!sk[56]) & (g642) & (g522) & (!g896) & (g1061)) + ((g46) & (!sk[56]) & (g642) & (g522) & (g896) & (!g1061)) + ((g46) & (!sk[56]) & (g642) & (g522) & (g896) & (g1061)));
	assign g1063 = (((!i_11_) & (!sk[57]) & (!g113) & (!g9) & (!g423) & (g1049)) + ((!i_11_) & (!sk[57]) & (!g113) & (!g9) & (g423) & (g1049)) + ((!i_11_) & (!sk[57]) & (!g113) & (g9) & (!g423) & (g1049)) + ((!i_11_) & (!sk[57]) & (!g113) & (g9) & (g423) & (g1049)) + ((!i_11_) & (!sk[57]) & (g113) & (!g9) & (!g423) & (g1049)) + ((!i_11_) & (!sk[57]) & (g113) & (!g9) & (g423) & (g1049)) + ((!i_11_) & (!sk[57]) & (g113) & (g9) & (!g423) & (g1049)) + ((!i_11_) & (!sk[57]) & (g113) & (g9) & (g423) & (g1049)) + ((!i_11_) & (sk[57]) & (!g113) & (!g9) & (g423) & (g1049)) + ((!i_11_) & (sk[57]) & (!g113) & (g9) & (g423) & (g1049)) + ((!i_11_) & (sk[57]) & (g113) & (!g9) & (g423) & (g1049)) + ((!i_11_) & (sk[57]) & (g113) & (g9) & (g423) & (g1049)) + ((i_11_) & (!sk[57]) & (!g113) & (!g9) & (!g423) & (!g1049)) + ((i_11_) & (!sk[57]) & (!g113) & (!g9) & (!g423) & (g1049)) + ((i_11_) & (!sk[57]) & (!g113) & (!g9) & (g423) & (!g1049)) + ((i_11_) & (!sk[57]) & (!g113) & (!g9) & (g423) & (g1049)) + ((i_11_) & (!sk[57]) & (!g113) & (g9) & (!g423) & (!g1049)) + ((i_11_) & (!sk[57]) & (!g113) & (g9) & (!g423) & (g1049)) + ((i_11_) & (!sk[57]) & (!g113) & (g9) & (g423) & (!g1049)) + ((i_11_) & (!sk[57]) & (!g113) & (g9) & (g423) & (g1049)) + ((i_11_) & (!sk[57]) & (g113) & (!g9) & (!g423) & (!g1049)) + ((i_11_) & (!sk[57]) & (g113) & (!g9) & (!g423) & (g1049)) + ((i_11_) & (!sk[57]) & (g113) & (!g9) & (g423) & (!g1049)) + ((i_11_) & (!sk[57]) & (g113) & (!g9) & (g423) & (g1049)) + ((i_11_) & (!sk[57]) & (g113) & (g9) & (!g423) & (!g1049)) + ((i_11_) & (!sk[57]) & (g113) & (g9) & (!g423) & (g1049)) + ((i_11_) & (!sk[57]) & (g113) & (g9) & (g423) & (!g1049)) + ((i_11_) & (!sk[57]) & (g113) & (g9) & (g423) & (g1049)) + ((i_11_) & (sk[57]) & (!g113) & (!g9) & (g423) & (g1049)) + ((i_11_) & (sk[57]) & (!g113) & (g9) & (g423) & (g1049)) + ((i_11_) & (sk[57]) & (g113) & (!g9) & (g423) & (g1049)) + ((i_11_) & (sk[57]) & (g113) & (g9) & (g423) & (!g1049)) + ((i_11_) & (sk[57]) & (g113) & (g9) & (g423) & (g1049)));
	assign g1064 = (((!g183) & (sk[58]) & (!g704) & (!g895)) + ((g183) & (!sk[58]) & (!g704) & (!g895)) + ((g183) & (!sk[58]) & (!g704) & (g895)) + ((g183) & (!sk[58]) & (g704) & (!g895)) + ((g183) & (!sk[58]) & (g704) & (g895)));
	assign g1065 = (((!g323) & (!g120) & (!sk[59]) & (g613) & (g1064)) + ((!g323) & (g120) & (!sk[59]) & (!g613) & (!g1064)) + ((!g323) & (g120) & (!sk[59]) & (!g613) & (g1064)) + ((!g323) & (g120) & (!sk[59]) & (g613) & (!g1064)) + ((!g323) & (g120) & (!sk[59]) & (g613) & (g1064)) + ((g323) & (!g120) & (!sk[59]) & (g613) & (!g1064)) + ((g323) & (!g120) & (!sk[59]) & (g613) & (g1064)) + ((g323) & (!g120) & (sk[59]) & (!g613) & (!g1064)) + ((g323) & (!g120) & (sk[59]) & (!g613) & (g1064)) + ((g323) & (!g120) & (sk[59]) & (g613) & (!g1064)) + ((g323) & (!g120) & (sk[59]) & (g613) & (g1064)) + ((g323) & (g120) & (!sk[59]) & (!g613) & (!g1064)) + ((g323) & (g120) & (!sk[59]) & (!g613) & (g1064)) + ((g323) & (g120) & (!sk[59]) & (g613) & (!g1064)) + ((g323) & (g120) & (!sk[59]) & (g613) & (g1064)) + ((g323) & (g120) & (sk[59]) & (!g613) & (!g1064)) + ((g323) & (g120) & (sk[59]) & (!g613) & (g1064)) + ((g323) & (g120) & (sk[59]) & (g613) & (!g1064)));
	assign g1066 = (((!g47) & (!sk[60]) & (!g323) & (g172) & (g142)) + ((!g47) & (!sk[60]) & (g323) & (!g172) & (!g142)) + ((!g47) & (!sk[60]) & (g323) & (!g172) & (g142)) + ((!g47) & (!sk[60]) & (g323) & (g172) & (!g142)) + ((!g47) & (!sk[60]) & (g323) & (g172) & (g142)) + ((!g47) & (sk[60]) & (g323) & (!g172) & (g142)) + ((!g47) & (sk[60]) & (g323) & (g172) & (!g142)) + ((!g47) & (sk[60]) & (g323) & (g172) & (g142)) + ((g47) & (!sk[60]) & (!g323) & (g172) & (!g142)) + ((g47) & (!sk[60]) & (!g323) & (g172) & (g142)) + ((g47) & (!sk[60]) & (g323) & (!g172) & (!g142)) + ((g47) & (!sk[60]) & (g323) & (!g172) & (g142)) + ((g47) & (!sk[60]) & (g323) & (g172) & (!g142)) + ((g47) & (!sk[60]) & (g323) & (g172) & (g142)) + ((g47) & (sk[60]) & (g323) & (!g172) & (!g142)) + ((g47) & (sk[60]) & (g323) & (!g172) & (g142)) + ((g47) & (sk[60]) & (g323) & (g172) & (!g142)) + ((g47) & (sk[60]) & (g323) & (g172) & (g142)));
	assign g1067 = (((!g44) & (!g323) & (!g191) & (!g339) & (!sk[61]) & (g807)) + ((!g44) & (!g323) & (!g191) & (g339) & (!sk[61]) & (g807)) + ((!g44) & (!g323) & (g191) & (!g339) & (!sk[61]) & (g807)) + ((!g44) & (!g323) & (g191) & (g339) & (!sk[61]) & (g807)) + ((!g44) & (g323) & (!g191) & (!g339) & (!sk[61]) & (g807)) + ((!g44) & (g323) & (!g191) & (!g339) & (sk[61]) & (!g807)) + ((!g44) & (g323) & (!g191) & (g339) & (!sk[61]) & (g807)) + ((!g44) & (g323) & (!g191) & (g339) & (sk[61]) & (!g807)) + ((!g44) & (g323) & (!g191) & (g339) & (sk[61]) & (g807)) + ((!g44) & (g323) & (g191) & (!g339) & (!sk[61]) & (g807)) + ((!g44) & (g323) & (g191) & (!g339) & (sk[61]) & (!g807)) + ((!g44) & (g323) & (g191) & (!g339) & (sk[61]) & (g807)) + ((!g44) & (g323) & (g191) & (g339) & (!sk[61]) & (g807)) + ((!g44) & (g323) & (g191) & (g339) & (sk[61]) & (!g807)) + ((!g44) & (g323) & (g191) & (g339) & (sk[61]) & (g807)) + ((g44) & (!g323) & (!g191) & (!g339) & (!sk[61]) & (!g807)) + ((g44) & (!g323) & (!g191) & (!g339) & (!sk[61]) & (g807)) + ((g44) & (!g323) & (!g191) & (g339) & (!sk[61]) & (!g807)) + ((g44) & (!g323) & (!g191) & (g339) & (!sk[61]) & (g807)) + ((g44) & (!g323) & (g191) & (!g339) & (!sk[61]) & (!g807)) + ((g44) & (!g323) & (g191) & (!g339) & (!sk[61]) & (g807)) + ((g44) & (!g323) & (g191) & (g339) & (!sk[61]) & (!g807)) + ((g44) & (!g323) & (g191) & (g339) & (!sk[61]) & (g807)) + ((g44) & (g323) & (!g191) & (!g339) & (!sk[61]) & (!g807)) + ((g44) & (g323) & (!g191) & (!g339) & (!sk[61]) & (g807)) + ((g44) & (g323) & (!g191) & (!g339) & (sk[61]) & (!g807)) + ((g44) & (g323) & (!g191) & (!g339) & (sk[61]) & (g807)) + ((g44) & (g323) & (!g191) & (g339) & (!sk[61]) & (!g807)) + ((g44) & (g323) & (!g191) & (g339) & (!sk[61]) & (g807)) + ((g44) & (g323) & (!g191) & (g339) & (sk[61]) & (!g807)) + ((g44) & (g323) & (!g191) & (g339) & (sk[61]) & (g807)) + ((g44) & (g323) & (g191) & (!g339) & (!sk[61]) & (!g807)) + ((g44) & (g323) & (g191) & (!g339) & (!sk[61]) & (g807)) + ((g44) & (g323) & (g191) & (!g339) & (sk[61]) & (!g807)) + ((g44) & (g323) & (g191) & (!g339) & (sk[61]) & (g807)) + ((g44) & (g323) & (g191) & (g339) & (!sk[61]) & (!g807)) + ((g44) & (g323) & (g191) & (g339) & (!sk[61]) & (g807)) + ((g44) & (g323) & (g191) & (g339) & (sk[61]) & (!g807)) + ((g44) & (g323) & (g191) & (g339) & (sk[61]) & (g807)));
	assign g1068 = (((!g323) & (!g465) & (!g899) & (!g1066) & (!sk[62]) & (g1067)) + ((!g323) & (!g465) & (!g899) & (!g1066) & (sk[62]) & (!g1067)) + ((!g323) & (!g465) & (!g899) & (g1066) & (!sk[62]) & (g1067)) + ((!g323) & (!g465) & (g899) & (!g1066) & (!sk[62]) & (g1067)) + ((!g323) & (!g465) & (g899) & (!g1066) & (sk[62]) & (!g1067)) + ((!g323) & (!g465) & (g899) & (g1066) & (!sk[62]) & (g1067)) + ((!g323) & (g465) & (!g899) & (!g1066) & (!sk[62]) & (g1067)) + ((!g323) & (g465) & (!g899) & (!g1066) & (sk[62]) & (!g1067)) + ((!g323) & (g465) & (!g899) & (g1066) & (!sk[62]) & (g1067)) + ((!g323) & (g465) & (g899) & (!g1066) & (!sk[62]) & (g1067)) + ((!g323) & (g465) & (g899) & (!g1066) & (sk[62]) & (!g1067)) + ((!g323) & (g465) & (g899) & (g1066) & (!sk[62]) & (g1067)) + ((g323) & (!g465) & (!g899) & (!g1066) & (!sk[62]) & (!g1067)) + ((g323) & (!g465) & (!g899) & (!g1066) & (!sk[62]) & (g1067)) + ((g323) & (!g465) & (!g899) & (g1066) & (!sk[62]) & (!g1067)) + ((g323) & (!g465) & (!g899) & (g1066) & (!sk[62]) & (g1067)) + ((g323) & (!g465) & (g899) & (!g1066) & (!sk[62]) & (!g1067)) + ((g323) & (!g465) & (g899) & (!g1066) & (!sk[62]) & (g1067)) + ((g323) & (!g465) & (g899) & (g1066) & (!sk[62]) & (!g1067)) + ((g323) & (!g465) & (g899) & (g1066) & (!sk[62]) & (g1067)) + ((g323) & (g465) & (!g899) & (!g1066) & (!sk[62]) & (!g1067)) + ((g323) & (g465) & (!g899) & (!g1066) & (!sk[62]) & (g1067)) + ((g323) & (g465) & (!g899) & (g1066) & (!sk[62]) & (!g1067)) + ((g323) & (g465) & (!g899) & (g1066) & (!sk[62]) & (g1067)) + ((g323) & (g465) & (g899) & (!g1066) & (!sk[62]) & (!g1067)) + ((g323) & (g465) & (g899) & (!g1066) & (!sk[62]) & (g1067)) + ((g323) & (g465) & (g899) & (!g1066) & (sk[62]) & (!g1067)) + ((g323) & (g465) & (g899) & (g1066) & (!sk[62]) & (!g1067)) + ((g323) & (g465) & (g899) & (g1066) & (!sk[62]) & (g1067)));
	assign g1069 = (((!g323) & (!g349) & (!sk[63]) & (g481) & (g540)) + ((!g323) & (g349) & (!sk[63]) & (!g481) & (!g540)) + ((!g323) & (g349) & (!sk[63]) & (!g481) & (g540)) + ((!g323) & (g349) & (!sk[63]) & (g481) & (!g540)) + ((!g323) & (g349) & (!sk[63]) & (g481) & (g540)) + ((g323) & (!g349) & (!sk[63]) & (g481) & (!g540)) + ((g323) & (!g349) & (!sk[63]) & (g481) & (g540)) + ((g323) & (!g349) & (sk[63]) & (!g481) & (!g540)) + ((g323) & (!g349) & (sk[63]) & (!g481) & (g540)) + ((g323) & (!g349) & (sk[63]) & (g481) & (g540)) + ((g323) & (g349) & (!sk[63]) & (!g481) & (!g540)) + ((g323) & (g349) & (!sk[63]) & (!g481) & (g540)) + ((g323) & (g349) & (!sk[63]) & (g481) & (!g540)) + ((g323) & (g349) & (!sk[63]) & (g481) & (g540)) + ((g323) & (g349) & (sk[63]) & (!g481) & (!g540)) + ((g323) & (g349) & (sk[63]) & (!g481) & (g540)) + ((g323) & (g349) & (sk[63]) & (g481) & (!g540)) + ((g323) & (g349) & (sk[63]) & (g481) & (g540)));
	assign g1070 = (((!g10) & (!g323) & (!g423) & (!g677) & (!g921) & (!g1069)) + ((!g10) & (!g323) & (!g423) & (!g677) & (g921) & (!g1069)) + ((!g10) & (!g323) & (!g423) & (g677) & (!g921) & (!g1069)) + ((!g10) & (!g323) & (!g423) & (g677) & (g921) & (!g1069)) + ((!g10) & (!g323) & (g423) & (!g677) & (g921) & (!g1069)) + ((!g10) & (!g323) & (g423) & (g677) & (g921) & (!g1069)) + ((!g10) & (g323) & (!g423) & (!g677) & (!g921) & (!g1069)) + ((!g10) & (g323) & (!g423) & (!g677) & (g921) & (!g1069)) + ((!g10) & (g323) & (g423) & (!g677) & (g921) & (!g1069)) + ((g10) & (!g323) & (!g423) & (!g677) & (!g921) & (!g1069)) + ((g10) & (!g323) & (!g423) & (!g677) & (g921) & (!g1069)) + ((g10) & (!g323) & (!g423) & (g677) & (!g921) & (!g1069)) + ((g10) & (!g323) & (!g423) & (g677) & (g921) & (!g1069)) + ((g10) & (!g323) & (g423) & (!g677) & (g921) & (!g1069)) + ((g10) & (!g323) & (g423) & (g677) & (g921) & (!g1069)));
	assign g1071 = (((!g207) & (!g323) & (!sk[65]) & (!g246) & (!g576) & (g724)) + ((!g207) & (!g323) & (!sk[65]) & (!g246) & (g576) & (g724)) + ((!g207) & (!g323) & (!sk[65]) & (g246) & (!g576) & (g724)) + ((!g207) & (!g323) & (!sk[65]) & (g246) & (g576) & (g724)) + ((!g207) & (g323) & (!sk[65]) & (!g246) & (!g576) & (g724)) + ((!g207) & (g323) & (!sk[65]) & (!g246) & (g576) & (g724)) + ((!g207) & (g323) & (!sk[65]) & (g246) & (!g576) & (g724)) + ((!g207) & (g323) & (!sk[65]) & (g246) & (g576) & (g724)) + ((!g207) & (g323) & (sk[65]) & (!g246) & (!g576) & (!g724)) + ((!g207) & (g323) & (sk[65]) & (!g246) & (!g576) & (g724)) + ((!g207) & (g323) & (sk[65]) & (!g246) & (g576) & (g724)) + ((!g207) & (g323) & (sk[65]) & (g246) & (!g576) & (!g724)) + ((!g207) & (g323) & (sk[65]) & (g246) & (!g576) & (g724)) + ((!g207) & (g323) & (sk[65]) & (g246) & (g576) & (!g724)) + ((!g207) & (g323) & (sk[65]) & (g246) & (g576) & (g724)) + ((g207) & (!g323) & (!sk[65]) & (!g246) & (!g576) & (!g724)) + ((g207) & (!g323) & (!sk[65]) & (!g246) & (!g576) & (g724)) + ((g207) & (!g323) & (!sk[65]) & (!g246) & (g576) & (!g724)) + ((g207) & (!g323) & (!sk[65]) & (!g246) & (g576) & (g724)) + ((g207) & (!g323) & (!sk[65]) & (g246) & (!g576) & (!g724)) + ((g207) & (!g323) & (!sk[65]) & (g246) & (!g576) & (g724)) + ((g207) & (!g323) & (!sk[65]) & (g246) & (g576) & (!g724)) + ((g207) & (!g323) & (!sk[65]) & (g246) & (g576) & (g724)) + ((g207) & (g323) & (!sk[65]) & (!g246) & (!g576) & (!g724)) + ((g207) & (g323) & (!sk[65]) & (!g246) & (!g576) & (g724)) + ((g207) & (g323) & (!sk[65]) & (!g246) & (g576) & (!g724)) + ((g207) & (g323) & (!sk[65]) & (!g246) & (g576) & (g724)) + ((g207) & (g323) & (!sk[65]) & (g246) & (!g576) & (!g724)) + ((g207) & (g323) & (!sk[65]) & (g246) & (!g576) & (g724)) + ((g207) & (g323) & (!sk[65]) & (g246) & (g576) & (!g724)) + ((g207) & (g323) & (!sk[65]) & (g246) & (g576) & (g724)) + ((g207) & (g323) & (sk[65]) & (!g246) & (!g576) & (!g724)) + ((g207) & (g323) & (sk[65]) & (!g246) & (!g576) & (g724)) + ((g207) & (g323) & (sk[65]) & (!g246) & (g576) & (!g724)) + ((g207) & (g323) & (sk[65]) & (!g246) & (g576) & (g724)) + ((g207) & (g323) & (sk[65]) & (g246) & (!g576) & (!g724)) + ((g207) & (g323) & (sk[65]) & (g246) & (!g576) & (g724)) + ((g207) & (g323) & (sk[65]) & (g246) & (g576) & (!g724)) + ((g207) & (g323) & (sk[65]) & (g246) & (g576) & (g724)));
	assign g1072 = (((!g8) & (!g221) & (!g323) & (!sk[66]) & (!g544) & (g1071)) + ((!g8) & (!g221) & (!g323) & (!sk[66]) & (g544) & (g1071)) + ((!g8) & (!g221) & (!g323) & (sk[66]) & (!g544) & (!g1071)) + ((!g8) & (!g221) & (!g323) & (sk[66]) & (g544) & (!g1071)) + ((!g8) & (!g221) & (g323) & (!sk[66]) & (!g544) & (g1071)) + ((!g8) & (!g221) & (g323) & (!sk[66]) & (g544) & (g1071)) + ((!g8) & (g221) & (!g323) & (!sk[66]) & (!g544) & (g1071)) + ((!g8) & (g221) & (!g323) & (!sk[66]) & (g544) & (g1071)) + ((!g8) & (g221) & (!g323) & (sk[66]) & (!g544) & (!g1071)) + ((!g8) & (g221) & (!g323) & (sk[66]) & (g544) & (!g1071)) + ((!g8) & (g221) & (g323) & (!sk[66]) & (!g544) & (g1071)) + ((!g8) & (g221) & (g323) & (!sk[66]) & (g544) & (g1071)) + ((g8) & (!g221) & (!g323) & (!sk[66]) & (!g544) & (!g1071)) + ((g8) & (!g221) & (!g323) & (!sk[66]) & (!g544) & (g1071)) + ((g8) & (!g221) & (!g323) & (!sk[66]) & (g544) & (!g1071)) + ((g8) & (!g221) & (!g323) & (!sk[66]) & (g544) & (g1071)) + ((g8) & (!g221) & (!g323) & (sk[66]) & (!g544) & (!g1071)) + ((g8) & (!g221) & (!g323) & (sk[66]) & (g544) & (!g1071)) + ((g8) & (!g221) & (g323) & (!sk[66]) & (!g544) & (!g1071)) + ((g8) & (!g221) & (g323) & (!sk[66]) & (!g544) & (g1071)) + ((g8) & (!g221) & (g323) & (!sk[66]) & (g544) & (!g1071)) + ((g8) & (!g221) & (g323) & (!sk[66]) & (g544) & (g1071)) + ((g8) & (g221) & (!g323) & (!sk[66]) & (!g544) & (!g1071)) + ((g8) & (g221) & (!g323) & (!sk[66]) & (!g544) & (g1071)) + ((g8) & (g221) & (!g323) & (!sk[66]) & (g544) & (!g1071)) + ((g8) & (g221) & (!g323) & (!sk[66]) & (g544) & (g1071)) + ((g8) & (g221) & (!g323) & (sk[66]) & (!g544) & (!g1071)) + ((g8) & (g221) & (!g323) & (sk[66]) & (g544) & (!g1071)) + ((g8) & (g221) & (g323) & (!sk[66]) & (!g544) & (!g1071)) + ((g8) & (g221) & (g323) & (!sk[66]) & (!g544) & (g1071)) + ((g8) & (g221) & (g323) & (!sk[66]) & (g544) & (!g1071)) + ((g8) & (g221) & (g323) & (!sk[66]) & (g544) & (g1071)) + ((g8) & (g221) & (g323) & (sk[66]) & (g544) & (!g1071)));
	assign g1073 = (((!sk[67]) & (!g1063) & (!g1065) & (!g1068) & (!g1070) & (g1072)) + ((!sk[67]) & (!g1063) & (!g1065) & (!g1068) & (g1070) & (g1072)) + ((!sk[67]) & (!g1063) & (!g1065) & (g1068) & (!g1070) & (g1072)) + ((!sk[67]) & (!g1063) & (!g1065) & (g1068) & (g1070) & (g1072)) + ((!sk[67]) & (!g1063) & (g1065) & (!g1068) & (!g1070) & (g1072)) + ((!sk[67]) & (!g1063) & (g1065) & (!g1068) & (g1070) & (g1072)) + ((!sk[67]) & (!g1063) & (g1065) & (g1068) & (!g1070) & (g1072)) + ((!sk[67]) & (!g1063) & (g1065) & (g1068) & (g1070) & (g1072)) + ((!sk[67]) & (g1063) & (!g1065) & (!g1068) & (!g1070) & (!g1072)) + ((!sk[67]) & (g1063) & (!g1065) & (!g1068) & (!g1070) & (g1072)) + ((!sk[67]) & (g1063) & (!g1065) & (!g1068) & (g1070) & (!g1072)) + ((!sk[67]) & (g1063) & (!g1065) & (!g1068) & (g1070) & (g1072)) + ((!sk[67]) & (g1063) & (!g1065) & (g1068) & (!g1070) & (!g1072)) + ((!sk[67]) & (g1063) & (!g1065) & (g1068) & (!g1070) & (g1072)) + ((!sk[67]) & (g1063) & (!g1065) & (g1068) & (g1070) & (!g1072)) + ((!sk[67]) & (g1063) & (!g1065) & (g1068) & (g1070) & (g1072)) + ((!sk[67]) & (g1063) & (g1065) & (!g1068) & (!g1070) & (!g1072)) + ((!sk[67]) & (g1063) & (g1065) & (!g1068) & (!g1070) & (g1072)) + ((!sk[67]) & (g1063) & (g1065) & (!g1068) & (g1070) & (!g1072)) + ((!sk[67]) & (g1063) & (g1065) & (!g1068) & (g1070) & (g1072)) + ((!sk[67]) & (g1063) & (g1065) & (g1068) & (!g1070) & (!g1072)) + ((!sk[67]) & (g1063) & (g1065) & (g1068) & (!g1070) & (g1072)) + ((!sk[67]) & (g1063) & (g1065) & (g1068) & (g1070) & (!g1072)) + ((!sk[67]) & (g1063) & (g1065) & (g1068) & (g1070) & (g1072)) + ((sk[67]) & (!g1063) & (!g1065) & (g1068) & (g1070) & (g1072)));
	assign g1074 = (((!sk[68]) & (!g243) & (!g1673) & (!g1060) & (!g1062) & (g1073)) + ((!sk[68]) & (!g243) & (!g1673) & (!g1060) & (g1062) & (g1073)) + ((!sk[68]) & (!g243) & (!g1673) & (g1060) & (!g1062) & (g1073)) + ((!sk[68]) & (!g243) & (!g1673) & (g1060) & (g1062) & (g1073)) + ((!sk[68]) & (!g243) & (g1673) & (!g1060) & (!g1062) & (g1073)) + ((!sk[68]) & (!g243) & (g1673) & (!g1060) & (g1062) & (g1073)) + ((!sk[68]) & (!g243) & (g1673) & (g1060) & (!g1062) & (g1073)) + ((!sk[68]) & (!g243) & (g1673) & (g1060) & (g1062) & (g1073)) + ((!sk[68]) & (g243) & (!g1673) & (!g1060) & (!g1062) & (!g1073)) + ((!sk[68]) & (g243) & (!g1673) & (!g1060) & (!g1062) & (g1073)) + ((!sk[68]) & (g243) & (!g1673) & (!g1060) & (g1062) & (!g1073)) + ((!sk[68]) & (g243) & (!g1673) & (!g1060) & (g1062) & (g1073)) + ((!sk[68]) & (g243) & (!g1673) & (g1060) & (!g1062) & (!g1073)) + ((!sk[68]) & (g243) & (!g1673) & (g1060) & (!g1062) & (g1073)) + ((!sk[68]) & (g243) & (!g1673) & (g1060) & (g1062) & (!g1073)) + ((!sk[68]) & (g243) & (!g1673) & (g1060) & (g1062) & (g1073)) + ((!sk[68]) & (g243) & (g1673) & (!g1060) & (!g1062) & (!g1073)) + ((!sk[68]) & (g243) & (g1673) & (!g1060) & (!g1062) & (g1073)) + ((!sk[68]) & (g243) & (g1673) & (!g1060) & (g1062) & (!g1073)) + ((!sk[68]) & (g243) & (g1673) & (!g1060) & (g1062) & (g1073)) + ((!sk[68]) & (g243) & (g1673) & (g1060) & (!g1062) & (!g1073)) + ((!sk[68]) & (g243) & (g1673) & (g1060) & (!g1062) & (g1073)) + ((!sk[68]) & (g243) & (g1673) & (g1060) & (g1062) & (!g1073)) + ((!sk[68]) & (g243) & (g1673) & (g1060) & (g1062) & (g1073)) + ((sk[68]) & (!g243) & (g1673) & (!g1060) & (!g1062) & (g1073)) + ((sk[68]) & (!g243) & (g1673) & (!g1060) & (g1062) & (g1073)) + ((sk[68]) & (!g243) & (g1673) & (g1060) & (!g1062) & (g1073)) + ((sk[68]) & (!g243) & (g1673) & (g1060) & (g1062) & (g1073)) + ((sk[68]) & (g243) & (g1673) & (!g1060) & (g1062) & (g1073)));
	assign g1075 = (((!g142) & (!sk[69]) & (!g540) & (g724) & (g895)) + ((!g142) & (!sk[69]) & (g540) & (!g724) & (!g895)) + ((!g142) & (!sk[69]) & (g540) & (!g724) & (g895)) + ((!g142) & (!sk[69]) & (g540) & (g724) & (!g895)) + ((!g142) & (!sk[69]) & (g540) & (g724) & (g895)) + ((!g142) & (sk[69]) & (!g540) & (!g724) & (!g895)) + ((g142) & (!sk[69]) & (!g540) & (g724) & (!g895)) + ((g142) & (!sk[69]) & (!g540) & (g724) & (g895)) + ((g142) & (!sk[69]) & (g540) & (!g724) & (!g895)) + ((g142) & (!sk[69]) & (g540) & (!g724) & (g895)) + ((g142) & (!sk[69]) & (g540) & (g724) & (!g895)) + ((g142) & (!sk[69]) & (g540) & (g724) & (g895)));
	assign g1076 = (((!sk[70]) & (!i_14_) & (!i_12_) & (i_13_) & (g102)) + ((!sk[70]) & (!i_14_) & (i_12_) & (!i_13_) & (!g102)) + ((!sk[70]) & (!i_14_) & (i_12_) & (!i_13_) & (g102)) + ((!sk[70]) & (!i_14_) & (i_12_) & (i_13_) & (!g102)) + ((!sk[70]) & (!i_14_) & (i_12_) & (i_13_) & (g102)) + ((!sk[70]) & (i_14_) & (!i_12_) & (i_13_) & (!g102)) + ((!sk[70]) & (i_14_) & (!i_12_) & (i_13_) & (g102)) + ((!sk[70]) & (i_14_) & (i_12_) & (!i_13_) & (!g102)) + ((!sk[70]) & (i_14_) & (i_12_) & (!i_13_) & (g102)) + ((!sk[70]) & (i_14_) & (i_12_) & (i_13_) & (!g102)) + ((!sk[70]) & (i_14_) & (i_12_) & (i_13_) & (g102)) + ((sk[70]) & (!i_14_) & (!i_12_) & (i_13_) & (!g102)) + ((sk[70]) & (!i_14_) & (i_12_) & (!i_13_) & (!g102)) + ((sk[70]) & (!i_14_) & (i_12_) & (i_13_) & (!g102)));
	assign g1077 = (((!g6) & (!i_15_) & (!i_14_) & (!i_12_) & (!sk[71]) & (i_13_)) + ((!g6) & (!i_15_) & (!i_14_) & (i_12_) & (!sk[71]) & (i_13_)) + ((!g6) & (!i_15_) & (i_14_) & (!i_12_) & (!sk[71]) & (i_13_)) + ((!g6) & (!i_15_) & (i_14_) & (i_12_) & (!sk[71]) & (i_13_)) + ((!g6) & (i_15_) & (!i_14_) & (!i_12_) & (!sk[71]) & (i_13_)) + ((!g6) & (i_15_) & (!i_14_) & (i_12_) & (!sk[71]) & (i_13_)) + ((!g6) & (i_15_) & (i_14_) & (!i_12_) & (!sk[71]) & (i_13_)) + ((!g6) & (i_15_) & (i_14_) & (i_12_) & (!sk[71]) & (i_13_)) + ((g6) & (!i_15_) & (!i_14_) & (!i_12_) & (!sk[71]) & (!i_13_)) + ((g6) & (!i_15_) & (!i_14_) & (!i_12_) & (!sk[71]) & (i_13_)) + ((g6) & (!i_15_) & (!i_14_) & (!i_12_) & (sk[71]) & (i_13_)) + ((g6) & (!i_15_) & (!i_14_) & (i_12_) & (!sk[71]) & (!i_13_)) + ((g6) & (!i_15_) & (!i_14_) & (i_12_) & (!sk[71]) & (i_13_)) + ((g6) & (!i_15_) & (!i_14_) & (i_12_) & (sk[71]) & (!i_13_)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (!sk[71]) & (!i_13_)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (!sk[71]) & (i_13_)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (sk[71]) & (i_13_)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (!sk[71]) & (!i_13_)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (!sk[71]) & (i_13_)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (sk[71]) & (i_13_)) + ((g6) & (i_15_) & (!i_14_) & (!i_12_) & (!sk[71]) & (!i_13_)) + ((g6) & (i_15_) & (!i_14_) & (!i_12_) & (!sk[71]) & (i_13_)) + ((g6) & (i_15_) & (!i_14_) & (!i_12_) & (sk[71]) & (!i_13_)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (!sk[71]) & (!i_13_)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (!sk[71]) & (i_13_)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (!sk[71]) & (!i_13_)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (!sk[71]) & (i_13_)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (sk[71]) & (!i_13_)) + ((g6) & (i_15_) & (i_14_) & (i_12_) & (!sk[71]) & (!i_13_)) + ((g6) & (i_15_) & (i_14_) & (i_12_) & (!sk[71]) & (i_13_)));
	assign g1078 = (((!g232) & (!g103) & (!sk[72]) & (g1076) & (g1077)) + ((!g232) & (g103) & (!sk[72]) & (!g1076) & (!g1077)) + ((!g232) & (g103) & (!sk[72]) & (!g1076) & (g1077)) + ((!g232) & (g103) & (!sk[72]) & (g1076) & (!g1077)) + ((!g232) & (g103) & (!sk[72]) & (g1076) & (g1077)) + ((!g232) & (g103) & (sk[72]) & (!g1076) & (!g1077)) + ((g232) & (!g103) & (!sk[72]) & (g1076) & (!g1077)) + ((g232) & (!g103) & (!sk[72]) & (g1076) & (g1077)) + ((g232) & (g103) & (!sk[72]) & (!g1076) & (!g1077)) + ((g232) & (g103) & (!sk[72]) & (!g1076) & (g1077)) + ((g232) & (g103) & (!sk[72]) & (g1076) & (!g1077)) + ((g232) & (g103) & (!sk[72]) & (g1076) & (g1077)));
	assign g1079 = (((!g44) & (!g183) & (!g191) & (!sk[73]) & (!g704) & (g756)) + ((!g44) & (!g183) & (!g191) & (!sk[73]) & (g704) & (g756)) + ((!g44) & (!g183) & (!g191) & (sk[73]) & (!g704) & (!g756)) + ((!g44) & (!g183) & (g191) & (!sk[73]) & (!g704) & (g756)) + ((!g44) & (!g183) & (g191) & (!sk[73]) & (g704) & (g756)) + ((!g44) & (g183) & (!g191) & (!sk[73]) & (!g704) & (g756)) + ((!g44) & (g183) & (!g191) & (!sk[73]) & (g704) & (g756)) + ((!g44) & (g183) & (g191) & (!sk[73]) & (!g704) & (g756)) + ((!g44) & (g183) & (g191) & (!sk[73]) & (g704) & (g756)) + ((g44) & (!g183) & (!g191) & (!sk[73]) & (!g704) & (!g756)) + ((g44) & (!g183) & (!g191) & (!sk[73]) & (!g704) & (g756)) + ((g44) & (!g183) & (!g191) & (!sk[73]) & (g704) & (!g756)) + ((g44) & (!g183) & (!g191) & (!sk[73]) & (g704) & (g756)) + ((g44) & (!g183) & (g191) & (!sk[73]) & (!g704) & (!g756)) + ((g44) & (!g183) & (g191) & (!sk[73]) & (!g704) & (g756)) + ((g44) & (!g183) & (g191) & (!sk[73]) & (g704) & (!g756)) + ((g44) & (!g183) & (g191) & (!sk[73]) & (g704) & (g756)) + ((g44) & (g183) & (!g191) & (!sk[73]) & (!g704) & (!g756)) + ((g44) & (g183) & (!g191) & (!sk[73]) & (!g704) & (g756)) + ((g44) & (g183) & (!g191) & (!sk[73]) & (g704) & (!g756)) + ((g44) & (g183) & (!g191) & (!sk[73]) & (g704) & (g756)) + ((g44) & (g183) & (g191) & (!sk[73]) & (!g704) & (!g756)) + ((g44) & (g183) & (g191) & (!sk[73]) & (!g704) & (g756)) + ((g44) & (g183) & (g191) & (!sk[73]) & (g704) & (!g756)) + ((g44) & (g183) & (g191) & (!sk[73]) & (g704) & (g756)));
	assign g1080 = (((!g316) & (!g172) & (!sk[74]) & (!g173) & (!g339) & (g1079)) + ((!g316) & (!g172) & (!sk[74]) & (!g173) & (g339) & (g1079)) + ((!g316) & (!g172) & (!sk[74]) & (g173) & (!g339) & (g1079)) + ((!g316) & (!g172) & (!sk[74]) & (g173) & (g339) & (g1079)) + ((!g316) & (!g172) & (sk[74]) & (!g173) & (!g339) & (g1079)) + ((!g316) & (g172) & (!sk[74]) & (!g173) & (!g339) & (g1079)) + ((!g316) & (g172) & (!sk[74]) & (!g173) & (g339) & (g1079)) + ((!g316) & (g172) & (!sk[74]) & (g173) & (!g339) & (g1079)) + ((!g316) & (g172) & (!sk[74]) & (g173) & (g339) & (g1079)) + ((g316) & (!g172) & (!sk[74]) & (!g173) & (!g339) & (!g1079)) + ((g316) & (!g172) & (!sk[74]) & (!g173) & (!g339) & (g1079)) + ((g316) & (!g172) & (!sk[74]) & (!g173) & (g339) & (!g1079)) + ((g316) & (!g172) & (!sk[74]) & (!g173) & (g339) & (g1079)) + ((g316) & (!g172) & (!sk[74]) & (g173) & (!g339) & (!g1079)) + ((g316) & (!g172) & (!sk[74]) & (g173) & (!g339) & (g1079)) + ((g316) & (!g172) & (!sk[74]) & (g173) & (g339) & (!g1079)) + ((g316) & (!g172) & (!sk[74]) & (g173) & (g339) & (g1079)) + ((g316) & (g172) & (!sk[74]) & (!g173) & (!g339) & (!g1079)) + ((g316) & (g172) & (!sk[74]) & (!g173) & (!g339) & (g1079)) + ((g316) & (g172) & (!sk[74]) & (!g173) & (g339) & (!g1079)) + ((g316) & (g172) & (!sk[74]) & (!g173) & (g339) & (g1079)) + ((g316) & (g172) & (!sk[74]) & (g173) & (!g339) & (!g1079)) + ((g316) & (g172) & (!sk[74]) & (g173) & (!g339) & (g1079)) + ((g316) & (g172) & (!sk[74]) & (g173) & (g339) & (!g1079)) + ((g316) & (g172) & (!sk[74]) & (g173) & (g339) & (g1079)));
	assign g1081 = (((!g222) & (!g908) & (!g1075) & (!sk[75]) & (!g1078) & (g1080)) + ((!g222) & (!g908) & (!g1075) & (!sk[75]) & (g1078) & (g1080)) + ((!g222) & (!g908) & (g1075) & (!sk[75]) & (!g1078) & (g1080)) + ((!g222) & (!g908) & (g1075) & (!sk[75]) & (g1078) & (g1080)) + ((!g222) & (!g908) & (g1075) & (sk[75]) & (g1078) & (g1080)) + ((!g222) & (g908) & (!g1075) & (!sk[75]) & (!g1078) & (g1080)) + ((!g222) & (g908) & (!g1075) & (!sk[75]) & (g1078) & (g1080)) + ((!g222) & (g908) & (g1075) & (!sk[75]) & (!g1078) & (g1080)) + ((!g222) & (g908) & (g1075) & (!sk[75]) & (g1078) & (g1080)) + ((g222) & (!g908) & (!g1075) & (!sk[75]) & (!g1078) & (!g1080)) + ((g222) & (!g908) & (!g1075) & (!sk[75]) & (!g1078) & (g1080)) + ((g222) & (!g908) & (!g1075) & (!sk[75]) & (g1078) & (!g1080)) + ((g222) & (!g908) & (!g1075) & (!sk[75]) & (g1078) & (g1080)) + ((g222) & (!g908) & (g1075) & (!sk[75]) & (!g1078) & (!g1080)) + ((g222) & (!g908) & (g1075) & (!sk[75]) & (!g1078) & (g1080)) + ((g222) & (!g908) & (g1075) & (!sk[75]) & (g1078) & (!g1080)) + ((g222) & (!g908) & (g1075) & (!sk[75]) & (g1078) & (g1080)) + ((g222) & (g908) & (!g1075) & (!sk[75]) & (!g1078) & (!g1080)) + ((g222) & (g908) & (!g1075) & (!sk[75]) & (!g1078) & (g1080)) + ((g222) & (g908) & (!g1075) & (!sk[75]) & (g1078) & (!g1080)) + ((g222) & (g908) & (!g1075) & (!sk[75]) & (g1078) & (g1080)) + ((g222) & (g908) & (g1075) & (!sk[75]) & (!g1078) & (!g1080)) + ((g222) & (g908) & (g1075) & (!sk[75]) & (!g1078) & (g1080)) + ((g222) & (g908) & (g1075) & (!sk[75]) & (g1078) & (!g1080)) + ((g222) & (g908) & (g1075) & (!sk[75]) & (g1078) & (g1080)));
	assign g1082 = (((i_14_) & (!sk[76]) & (!i_12_) & (!g115)) + ((i_14_) & (!sk[76]) & (!i_12_) & (g115)) + ((i_14_) & (!sk[76]) & (i_12_) & (!g115)) + ((i_14_) & (!sk[76]) & (i_12_) & (g115)) + ((i_14_) & (sk[76]) & (!i_12_) & (!g115)));
	assign g1083 = (((!g19) & (g201) & (!g675) & (!g797) & (!g703) & (!g1082)));
	assign g1084 = (((!g132) & (!g576) & (!sk[78]) & (!g557) & (!g465) & (g1083)) + ((!g132) & (!g576) & (!sk[78]) & (!g557) & (g465) & (g1083)) + ((!g132) & (!g576) & (!sk[78]) & (g557) & (!g465) & (g1083)) + ((!g132) & (!g576) & (!sk[78]) & (g557) & (g465) & (g1083)) + ((!g132) & (g576) & (!sk[78]) & (!g557) & (!g465) & (g1083)) + ((!g132) & (g576) & (!sk[78]) & (!g557) & (g465) & (g1083)) + ((!g132) & (g576) & (!sk[78]) & (g557) & (!g465) & (g1083)) + ((!g132) & (g576) & (!sk[78]) & (g557) & (g465) & (g1083)) + ((g132) & (!g576) & (!sk[78]) & (!g557) & (!g465) & (!g1083)) + ((g132) & (!g576) & (!sk[78]) & (!g557) & (!g465) & (g1083)) + ((g132) & (!g576) & (!sk[78]) & (!g557) & (g465) & (!g1083)) + ((g132) & (!g576) & (!sk[78]) & (!g557) & (g465) & (g1083)) + ((g132) & (!g576) & (!sk[78]) & (g557) & (!g465) & (!g1083)) + ((g132) & (!g576) & (!sk[78]) & (g557) & (!g465) & (g1083)) + ((g132) & (!g576) & (!sk[78]) & (g557) & (g465) & (!g1083)) + ((g132) & (!g576) & (!sk[78]) & (g557) & (g465) & (g1083)) + ((g132) & (g576) & (!sk[78]) & (!g557) & (!g465) & (!g1083)) + ((g132) & (g576) & (!sk[78]) & (!g557) & (!g465) & (g1083)) + ((g132) & (g576) & (!sk[78]) & (!g557) & (g465) & (!g1083)) + ((g132) & (g576) & (!sk[78]) & (!g557) & (g465) & (g1083)) + ((g132) & (g576) & (!sk[78]) & (g557) & (!g465) & (!g1083)) + ((g132) & (g576) & (!sk[78]) & (g557) & (!g465) & (g1083)) + ((g132) & (g576) & (!sk[78]) & (g557) & (g465) & (!g1083)) + ((g132) & (g576) & (!sk[78]) & (g557) & (g465) & (g1083)) + ((g132) & (g576) & (sk[78]) & (!g557) & (g465) & (g1083)));
	assign g1085 = (((!g207) & (!g213) & (!g279) & (!sk[79]) & (!g544) & (g881)) + ((!g207) & (!g213) & (!g279) & (!sk[79]) & (g544) & (g881)) + ((!g207) & (!g213) & (!g279) & (sk[79]) & (g544) & (!g881)) + ((!g207) & (!g213) & (g279) & (!sk[79]) & (!g544) & (g881)) + ((!g207) & (!g213) & (g279) & (!sk[79]) & (g544) & (g881)) + ((!g207) & (g213) & (!g279) & (!sk[79]) & (!g544) & (g881)) + ((!g207) & (g213) & (!g279) & (!sk[79]) & (g544) & (g881)) + ((!g207) & (g213) & (g279) & (!sk[79]) & (!g544) & (g881)) + ((!g207) & (g213) & (g279) & (!sk[79]) & (g544) & (g881)) + ((g207) & (!g213) & (!g279) & (!sk[79]) & (!g544) & (!g881)) + ((g207) & (!g213) & (!g279) & (!sk[79]) & (!g544) & (g881)) + ((g207) & (!g213) & (!g279) & (!sk[79]) & (g544) & (!g881)) + ((g207) & (!g213) & (!g279) & (!sk[79]) & (g544) & (g881)) + ((g207) & (!g213) & (g279) & (!sk[79]) & (!g544) & (!g881)) + ((g207) & (!g213) & (g279) & (!sk[79]) & (!g544) & (g881)) + ((g207) & (!g213) & (g279) & (!sk[79]) & (g544) & (!g881)) + ((g207) & (!g213) & (g279) & (!sk[79]) & (g544) & (g881)) + ((g207) & (g213) & (!g279) & (!sk[79]) & (!g544) & (!g881)) + ((g207) & (g213) & (!g279) & (!sk[79]) & (!g544) & (g881)) + ((g207) & (g213) & (!g279) & (!sk[79]) & (g544) & (!g881)) + ((g207) & (g213) & (!g279) & (!sk[79]) & (g544) & (g881)) + ((g207) & (g213) & (g279) & (!sk[79]) & (!g544) & (!g881)) + ((g207) & (g213) & (g279) & (!sk[79]) & (!g544) & (g881)) + ((g207) & (g213) & (g279) & (!sk[79]) & (g544) & (!g881)) + ((g207) & (g213) & (g279) & (!sk[79]) & (g544) & (g881)));
	assign g1086 = (((!sk[80]) & (g243) & (!g630) & (!g980)) + ((!sk[80]) & (g243) & (!g630) & (g980)) + ((!sk[80]) & (g243) & (g630) & (!g980)) + ((!sk[80]) & (g243) & (g630) & (g980)) + ((sk[80]) & (g243) & (!g630) & (!g980)) + ((sk[80]) & (g243) & (g630) & (!g980)) + ((sk[80]) & (g243) & (g630) & (g980)));
	assign g1087 = (((!g323) & (!sk[81]) & (!g173) & (g103) & (g546)) + ((!g323) & (!sk[81]) & (g173) & (!g103) & (!g546)) + ((!g323) & (!sk[81]) & (g173) & (!g103) & (g546)) + ((!g323) & (!sk[81]) & (g173) & (g103) & (!g546)) + ((!g323) & (!sk[81]) & (g173) & (g103) & (g546)) + ((g323) & (!sk[81]) & (!g173) & (g103) & (!g546)) + ((g323) & (!sk[81]) & (!g173) & (g103) & (g546)) + ((g323) & (!sk[81]) & (g173) & (!g103) & (!g546)) + ((g323) & (!sk[81]) & (g173) & (!g103) & (g546)) + ((g323) & (!sk[81]) & (g173) & (g103) & (!g546)) + ((g323) & (!sk[81]) & (g173) & (g103) & (g546)) + ((g323) & (sk[81]) & (!g173) & (!g103) & (!g546)) + ((g323) & (sk[81]) & (!g173) & (!g103) & (g546)) + ((g323) & (sk[81]) & (!g173) & (g103) & (g546)) + ((g323) & (sk[81]) & (g173) & (!g103) & (!g546)) + ((g323) & (sk[81]) & (g173) & (!g103) & (g546)) + ((g323) & (sk[81]) & (g173) & (g103) & (!g546)) + ((g323) & (sk[81]) & (g173) & (g103) & (g546)));
	assign g1088 = (((!g187) & (!g423) & (!g534) & (!sk[82]) & (!g907) & (g1087)) + ((!g187) & (!g423) & (!g534) & (!sk[82]) & (g907) & (g1087)) + ((!g187) & (!g423) & (!g534) & (sk[82]) & (!g907) & (!g1087)) + ((!g187) & (!g423) & (!g534) & (sk[82]) & (g907) & (!g1087)) + ((!g187) & (!g423) & (g534) & (!sk[82]) & (!g907) & (g1087)) + ((!g187) & (!g423) & (g534) & (!sk[82]) & (g907) & (g1087)) + ((!g187) & (!g423) & (g534) & (sk[82]) & (!g907) & (!g1087)) + ((!g187) & (!g423) & (g534) & (sk[82]) & (g907) & (!g1087)) + ((!g187) & (g423) & (!g534) & (!sk[82]) & (!g907) & (g1087)) + ((!g187) & (g423) & (!g534) & (!sk[82]) & (g907) & (g1087)) + ((!g187) & (g423) & (!g534) & (sk[82]) & (!g907) & (!g1087)) + ((!g187) & (g423) & (g534) & (!sk[82]) & (!g907) & (g1087)) + ((!g187) & (g423) & (g534) & (!sk[82]) & (g907) & (g1087)) + ((g187) & (!g423) & (!g534) & (!sk[82]) & (!g907) & (!g1087)) + ((g187) & (!g423) & (!g534) & (!sk[82]) & (!g907) & (g1087)) + ((g187) & (!g423) & (!g534) & (!sk[82]) & (g907) & (!g1087)) + ((g187) & (!g423) & (!g534) & (!sk[82]) & (g907) & (g1087)) + ((g187) & (!g423) & (!g534) & (sk[82]) & (!g907) & (!g1087)) + ((g187) & (!g423) & (!g534) & (sk[82]) & (g907) & (!g1087)) + ((g187) & (!g423) & (g534) & (!sk[82]) & (!g907) & (!g1087)) + ((g187) & (!g423) & (g534) & (!sk[82]) & (!g907) & (g1087)) + ((g187) & (!g423) & (g534) & (!sk[82]) & (g907) & (!g1087)) + ((g187) & (!g423) & (g534) & (!sk[82]) & (g907) & (g1087)) + ((g187) & (!g423) & (g534) & (sk[82]) & (!g907) & (!g1087)) + ((g187) & (!g423) & (g534) & (sk[82]) & (g907) & (!g1087)) + ((g187) & (g423) & (!g534) & (!sk[82]) & (!g907) & (!g1087)) + ((g187) & (g423) & (!g534) & (!sk[82]) & (!g907) & (g1087)) + ((g187) & (g423) & (!g534) & (!sk[82]) & (g907) & (!g1087)) + ((g187) & (g423) & (!g534) & (!sk[82]) & (g907) & (g1087)) + ((g187) & (g423) & (g534) & (!sk[82]) & (!g907) & (!g1087)) + ((g187) & (g423) & (g534) & (!sk[82]) & (!g907) & (g1087)) + ((g187) & (g423) & (g534) & (!sk[82]) & (g907) & (!g1087)) + ((g187) & (g423) & (g534) & (!sk[82]) & (g907) & (g1087)));
	assign g1089 = (((!sk[83]) & (!i_11_) & (!i_10_) & (g323) & (g875)) + ((!sk[83]) & (!i_11_) & (i_10_) & (!g323) & (!g875)) + ((!sk[83]) & (!i_11_) & (i_10_) & (!g323) & (g875)) + ((!sk[83]) & (!i_11_) & (i_10_) & (g323) & (!g875)) + ((!sk[83]) & (!i_11_) & (i_10_) & (g323) & (g875)) + ((!sk[83]) & (i_11_) & (!i_10_) & (g323) & (!g875)) + ((!sk[83]) & (i_11_) & (!i_10_) & (g323) & (g875)) + ((!sk[83]) & (i_11_) & (i_10_) & (!g323) & (!g875)) + ((!sk[83]) & (i_11_) & (i_10_) & (!g323) & (g875)) + ((!sk[83]) & (i_11_) & (i_10_) & (g323) & (!g875)) + ((!sk[83]) & (i_11_) & (i_10_) & (g323) & (g875)) + ((sk[83]) & (i_11_) & (i_10_) & (g323) & (g875)));
	assign g1090 = (((!g48) & (!sk[84]) & (!g323) & (!g182) & (!g124) & (g115)) + ((!g48) & (!sk[84]) & (!g323) & (!g182) & (g124) & (g115)) + ((!g48) & (!sk[84]) & (!g323) & (g182) & (!g124) & (g115)) + ((!g48) & (!sk[84]) & (!g323) & (g182) & (g124) & (g115)) + ((!g48) & (!sk[84]) & (g323) & (!g182) & (!g124) & (g115)) + ((!g48) & (!sk[84]) & (g323) & (!g182) & (g124) & (g115)) + ((!g48) & (!sk[84]) & (g323) & (g182) & (!g124) & (g115)) + ((!g48) & (!sk[84]) & (g323) & (g182) & (g124) & (g115)) + ((!g48) & (sk[84]) & (g323) & (!g182) & (!g124) & (!g115)) + ((!g48) & (sk[84]) & (g323) & (!g182) & (g124) & (!g115)) + ((!g48) & (sk[84]) & (g323) & (!g182) & (g124) & (g115)) + ((!g48) & (sk[84]) & (g323) & (g182) & (!g124) & (!g115)) + ((!g48) & (sk[84]) & (g323) & (g182) & (g124) & (!g115)) + ((!g48) & (sk[84]) & (g323) & (g182) & (g124) & (g115)) + ((g48) & (!sk[84]) & (!g323) & (!g182) & (!g124) & (!g115)) + ((g48) & (!sk[84]) & (!g323) & (!g182) & (!g124) & (g115)) + ((g48) & (!sk[84]) & (!g323) & (!g182) & (g124) & (!g115)) + ((g48) & (!sk[84]) & (!g323) & (!g182) & (g124) & (g115)) + ((g48) & (!sk[84]) & (!g323) & (g182) & (!g124) & (!g115)) + ((g48) & (!sk[84]) & (!g323) & (g182) & (!g124) & (g115)) + ((g48) & (!sk[84]) & (!g323) & (g182) & (g124) & (!g115)) + ((g48) & (!sk[84]) & (!g323) & (g182) & (g124) & (g115)) + ((g48) & (!sk[84]) & (g323) & (!g182) & (!g124) & (!g115)) + ((g48) & (!sk[84]) & (g323) & (!g182) & (!g124) & (g115)) + ((g48) & (!sk[84]) & (g323) & (!g182) & (g124) & (!g115)) + ((g48) & (!sk[84]) & (g323) & (!g182) & (g124) & (g115)) + ((g48) & (!sk[84]) & (g323) & (g182) & (!g124) & (!g115)) + ((g48) & (!sk[84]) & (g323) & (g182) & (!g124) & (g115)) + ((g48) & (!sk[84]) & (g323) & (g182) & (g124) & (!g115)) + ((g48) & (!sk[84]) & (g323) & (g182) & (g124) & (g115)) + ((g48) & (sk[84]) & (g323) & (g182) & (!g124) & (!g115)) + ((g48) & (sk[84]) & (g323) & (g182) & (g124) & (!g115)) + ((g48) & (sk[84]) & (g323) & (g182) & (g124) & (g115)));
	assign g1091 = (((!g323) & (!g696) & (!g702) & (!g827) & (!g914) & (!g1090)) + ((!g323) & (!g696) & (!g702) & (!g827) & (g914) & (!g1090)) + ((!g323) & (!g696) & (!g702) & (g827) & (!g914) & (!g1090)) + ((!g323) & (!g696) & (!g702) & (g827) & (g914) & (!g1090)) + ((!g323) & (!g696) & (g702) & (!g827) & (!g914) & (!g1090)) + ((!g323) & (!g696) & (g702) & (!g827) & (g914) & (!g1090)) + ((!g323) & (!g696) & (g702) & (g827) & (!g914) & (!g1090)) + ((!g323) & (!g696) & (g702) & (g827) & (g914) & (!g1090)) + ((!g323) & (g696) & (!g702) & (!g827) & (!g914) & (!g1090)) + ((!g323) & (g696) & (!g702) & (!g827) & (g914) & (!g1090)) + ((!g323) & (g696) & (!g702) & (g827) & (!g914) & (!g1090)) + ((!g323) & (g696) & (!g702) & (g827) & (g914) & (!g1090)) + ((!g323) & (g696) & (g702) & (!g827) & (!g914) & (!g1090)) + ((!g323) & (g696) & (g702) & (!g827) & (g914) & (!g1090)) + ((!g323) & (g696) & (g702) & (g827) & (!g914) & (!g1090)) + ((!g323) & (g696) & (g702) & (g827) & (g914) & (!g1090)) + ((g323) & (g696) & (!g702) & (g827) & (g914) & (!g1090)));
	assign g1092 = (((!g829) & (!g1086) & (!g1088) & (!sk[86]) & (!g1089) & (g1091)) + ((!g829) & (!g1086) & (!g1088) & (!sk[86]) & (g1089) & (g1091)) + ((!g829) & (!g1086) & (g1088) & (!sk[86]) & (!g1089) & (g1091)) + ((!g829) & (!g1086) & (g1088) & (!sk[86]) & (g1089) & (g1091)) + ((!g829) & (!g1086) & (g1088) & (sk[86]) & (!g1089) & (g1091)) + ((!g829) & (g1086) & (!g1088) & (!sk[86]) & (!g1089) & (g1091)) + ((!g829) & (g1086) & (!g1088) & (!sk[86]) & (g1089) & (g1091)) + ((!g829) & (g1086) & (g1088) & (!sk[86]) & (!g1089) & (g1091)) + ((!g829) & (g1086) & (g1088) & (!sk[86]) & (g1089) & (g1091)) + ((g829) & (!g1086) & (!g1088) & (!sk[86]) & (!g1089) & (!g1091)) + ((g829) & (!g1086) & (!g1088) & (!sk[86]) & (!g1089) & (g1091)) + ((g829) & (!g1086) & (!g1088) & (!sk[86]) & (g1089) & (!g1091)) + ((g829) & (!g1086) & (!g1088) & (!sk[86]) & (g1089) & (g1091)) + ((g829) & (!g1086) & (g1088) & (!sk[86]) & (!g1089) & (!g1091)) + ((g829) & (!g1086) & (g1088) & (!sk[86]) & (!g1089) & (g1091)) + ((g829) & (!g1086) & (g1088) & (!sk[86]) & (g1089) & (!g1091)) + ((g829) & (!g1086) & (g1088) & (!sk[86]) & (g1089) & (g1091)) + ((g829) & (g1086) & (!g1088) & (!sk[86]) & (!g1089) & (!g1091)) + ((g829) & (g1086) & (!g1088) & (!sk[86]) & (!g1089) & (g1091)) + ((g829) & (g1086) & (!g1088) & (!sk[86]) & (g1089) & (!g1091)) + ((g829) & (g1086) & (!g1088) & (!sk[86]) & (g1089) & (g1091)) + ((g829) & (g1086) & (g1088) & (!sk[86]) & (!g1089) & (!g1091)) + ((g829) & (g1086) & (g1088) & (!sk[86]) & (!g1089) & (g1091)) + ((g829) & (g1086) & (g1088) & (!sk[86]) & (g1089) & (!g1091)) + ((g829) & (g1086) & (g1088) & (!sk[86]) & (g1089) & (g1091)));
	assign g1093 = (((!g423) & (!g1081) & (!sk[87]) & (!g1084) & (!g1085) & (g1092)) + ((!g423) & (!g1081) & (!sk[87]) & (!g1084) & (g1085) & (g1092)) + ((!g423) & (!g1081) & (!sk[87]) & (g1084) & (!g1085) & (g1092)) + ((!g423) & (!g1081) & (!sk[87]) & (g1084) & (g1085) & (g1092)) + ((!g423) & (!g1081) & (sk[87]) & (!g1084) & (!g1085) & (g1092)) + ((!g423) & (!g1081) & (sk[87]) & (!g1084) & (g1085) & (g1092)) + ((!g423) & (!g1081) & (sk[87]) & (g1084) & (!g1085) & (g1092)) + ((!g423) & (!g1081) & (sk[87]) & (g1084) & (g1085) & (g1092)) + ((!g423) & (g1081) & (!sk[87]) & (!g1084) & (!g1085) & (g1092)) + ((!g423) & (g1081) & (!sk[87]) & (!g1084) & (g1085) & (g1092)) + ((!g423) & (g1081) & (!sk[87]) & (g1084) & (!g1085) & (g1092)) + ((!g423) & (g1081) & (!sk[87]) & (g1084) & (g1085) & (g1092)) + ((!g423) & (g1081) & (sk[87]) & (!g1084) & (!g1085) & (g1092)) + ((!g423) & (g1081) & (sk[87]) & (!g1084) & (g1085) & (g1092)) + ((!g423) & (g1081) & (sk[87]) & (g1084) & (!g1085) & (g1092)) + ((!g423) & (g1081) & (sk[87]) & (g1084) & (g1085) & (g1092)) + ((g423) & (!g1081) & (!sk[87]) & (!g1084) & (!g1085) & (!g1092)) + ((g423) & (!g1081) & (!sk[87]) & (!g1084) & (!g1085) & (g1092)) + ((g423) & (!g1081) & (!sk[87]) & (!g1084) & (g1085) & (!g1092)) + ((g423) & (!g1081) & (!sk[87]) & (!g1084) & (g1085) & (g1092)) + ((g423) & (!g1081) & (!sk[87]) & (g1084) & (!g1085) & (!g1092)) + ((g423) & (!g1081) & (!sk[87]) & (g1084) & (!g1085) & (g1092)) + ((g423) & (!g1081) & (!sk[87]) & (g1084) & (g1085) & (!g1092)) + ((g423) & (!g1081) & (!sk[87]) & (g1084) & (g1085) & (g1092)) + ((g423) & (g1081) & (!sk[87]) & (!g1084) & (!g1085) & (!g1092)) + ((g423) & (g1081) & (!sk[87]) & (!g1084) & (!g1085) & (g1092)) + ((g423) & (g1081) & (!sk[87]) & (!g1084) & (g1085) & (!g1092)) + ((g423) & (g1081) & (!sk[87]) & (!g1084) & (g1085) & (g1092)) + ((g423) & (g1081) & (!sk[87]) & (g1084) & (!g1085) & (!g1092)) + ((g423) & (g1081) & (!sk[87]) & (g1084) & (!g1085) & (g1092)) + ((g423) & (g1081) & (!sk[87]) & (g1084) & (g1085) & (!g1092)) + ((g423) & (g1081) & (!sk[87]) & (g1084) & (g1085) & (g1092)) + ((g423) & (g1081) & (sk[87]) & (g1084) & (g1085) & (g1092)));
	assign g1094 = (((g1045) & (g1047) & (g1051) & (g1059) & (g1074) & (g1093)));
	assign g1095 = (((!sk[89]) & (g89) & (!g627)) + ((!sk[89]) & (g89) & (g627)) + ((sk[89]) & (!g89) & (!g627)));
	assign g1096 = (((!sk[90]) & (g21) & (!g114)) + ((!sk[90]) & (g21) & (g114)) + ((sk[90]) & (!g21) & (!g114)));
	assign g1097 = (((!i_14_) & (!i_13_) & (sk[91]) & (g22)) + ((i_14_) & (!i_13_) & (!sk[91]) & (!g22)) + ((i_14_) & (!i_13_) & (!sk[91]) & (g22)) + ((i_14_) & (i_13_) & (!sk[91]) & (!g22)) + ((i_14_) & (i_13_) & (!sk[91]) & (g22)));
	assign g1098 = (((!g151) & (!sk[92]) & (!g506) & (!g594) & (!g1096) & (g1097)) + ((!g151) & (!sk[92]) & (!g506) & (!g594) & (g1096) & (g1097)) + ((!g151) & (!sk[92]) & (!g506) & (g594) & (!g1096) & (g1097)) + ((!g151) & (!sk[92]) & (!g506) & (g594) & (g1096) & (g1097)) + ((!g151) & (!sk[92]) & (g506) & (!g594) & (!g1096) & (g1097)) + ((!g151) & (!sk[92]) & (g506) & (!g594) & (g1096) & (g1097)) + ((!g151) & (!sk[92]) & (g506) & (g594) & (!g1096) & (g1097)) + ((!g151) & (!sk[92]) & (g506) & (g594) & (g1096) & (g1097)) + ((g151) & (!sk[92]) & (!g506) & (!g594) & (!g1096) & (!g1097)) + ((g151) & (!sk[92]) & (!g506) & (!g594) & (!g1096) & (g1097)) + ((g151) & (!sk[92]) & (!g506) & (!g594) & (g1096) & (!g1097)) + ((g151) & (!sk[92]) & (!g506) & (!g594) & (g1096) & (g1097)) + ((g151) & (!sk[92]) & (!g506) & (g594) & (!g1096) & (!g1097)) + ((g151) & (!sk[92]) & (!g506) & (g594) & (!g1096) & (g1097)) + ((g151) & (!sk[92]) & (!g506) & (g594) & (g1096) & (!g1097)) + ((g151) & (!sk[92]) & (!g506) & (g594) & (g1096) & (g1097)) + ((g151) & (!sk[92]) & (g506) & (!g594) & (!g1096) & (!g1097)) + ((g151) & (!sk[92]) & (g506) & (!g594) & (!g1096) & (g1097)) + ((g151) & (!sk[92]) & (g506) & (!g594) & (g1096) & (!g1097)) + ((g151) & (!sk[92]) & (g506) & (!g594) & (g1096) & (g1097)) + ((g151) & (!sk[92]) & (g506) & (g594) & (!g1096) & (!g1097)) + ((g151) & (!sk[92]) & (g506) & (g594) & (!g1096) & (g1097)) + ((g151) & (!sk[92]) & (g506) & (g594) & (g1096) & (!g1097)) + ((g151) & (!sk[92]) & (g506) & (g594) & (g1096) & (g1097)) + ((g151) & (sk[92]) & (!g506) & (!g594) & (!g1096) & (!g1097)) + ((g151) & (sk[92]) & (!g506) & (!g594) & (!g1096) & (g1097)) + ((g151) & (sk[92]) & (!g506) & (!g594) & (g1096) & (!g1097)) + ((g151) & (sk[92]) & (!g506) & (!g594) & (g1096) & (g1097)) + ((g151) & (sk[92]) & (!g506) & (g594) & (!g1096) & (!g1097)) + ((g151) & (sk[92]) & (!g506) & (g594) & (!g1096) & (g1097)) + ((g151) & (sk[92]) & (!g506) & (g594) & (g1096) & (g1097)) + ((g151) & (sk[92]) & (g506) & (!g594) & (!g1096) & (!g1097)) + ((g151) & (sk[92]) & (g506) & (!g594) & (!g1096) & (g1097)) + ((g151) & (sk[92]) & (g506) & (!g594) & (g1096) & (!g1097)) + ((g151) & (sk[92]) & (g506) & (!g594) & (g1096) & (g1097)) + ((g151) & (sk[92]) & (g506) & (g594) & (!g1096) & (!g1097)) + ((g151) & (sk[92]) & (g506) & (g594) & (!g1096) & (g1097)) + ((g151) & (sk[92]) & (g506) & (g594) & (g1096) & (!g1097)) + ((g151) & (sk[92]) & (g506) & (g594) & (g1096) & (g1097)));
	assign g1099 = (((!sk[93]) & (g187) & (!g982)) + ((!sk[93]) & (g187) & (g982)) + ((sk[93]) & (!g187) & (g982)));
	assign g1100 = (((!sk[94]) & (g151) & (!g534) & (!g1099)) + ((!sk[94]) & (g151) & (!g534) & (g1099)) + ((!sk[94]) & (g151) & (g534) & (!g1099)) + ((!sk[94]) & (g151) & (g534) & (g1099)) + ((sk[94]) & (g151) & (!g534) & (!g1099)) + ((sk[94]) & (g151) & (g534) & (!g1099)) + ((sk[94]) & (g151) & (g534) & (g1099)));
	assign g1101 = (((!g1095) & (!sk[95]) & (!g1098) & (g1100) & (g1541)) + ((!g1095) & (!sk[95]) & (g1098) & (!g1100) & (!g1541)) + ((!g1095) & (!sk[95]) & (g1098) & (!g1100) & (g1541)) + ((!g1095) & (!sk[95]) & (g1098) & (g1100) & (!g1541)) + ((!g1095) & (!sk[95]) & (g1098) & (g1100) & (g1541)) + ((!g1095) & (sk[95]) & (!g1098) & (!g1100) & (g1541)) + ((g1095) & (!sk[95]) & (!g1098) & (g1100) & (!g1541)) + ((g1095) & (!sk[95]) & (!g1098) & (g1100) & (g1541)) + ((g1095) & (!sk[95]) & (g1098) & (!g1100) & (!g1541)) + ((g1095) & (!sk[95]) & (g1098) & (!g1100) & (g1541)) + ((g1095) & (!sk[95]) & (g1098) & (g1100) & (!g1541)) + ((g1095) & (!sk[95]) & (g1098) & (g1100) & (g1541)));
	assign g1102 = (((!i_8_) & (!g46) & (!sk[96]) & (!g88) & (!g224) & (g811)) + ((!i_8_) & (!g46) & (!sk[96]) & (!g88) & (g224) & (g811)) + ((!i_8_) & (!g46) & (!sk[96]) & (g88) & (!g224) & (g811)) + ((!i_8_) & (!g46) & (!sk[96]) & (g88) & (g224) & (g811)) + ((!i_8_) & (!g46) & (sk[96]) & (!g88) & (!g224) & (!g811)) + ((!i_8_) & (!g46) & (sk[96]) & (!g88) & (!g224) & (g811)) + ((!i_8_) & (!g46) & (sk[96]) & (!g88) & (g224) & (!g811)) + ((!i_8_) & (!g46) & (sk[96]) & (!g88) & (g224) & (g811)) + ((!i_8_) & (!g46) & (sk[96]) & (g88) & (!g224) & (!g811)) + ((!i_8_) & (!g46) & (sk[96]) & (g88) & (!g224) & (g811)) + ((!i_8_) & (!g46) & (sk[96]) & (g88) & (g224) & (!g811)) + ((!i_8_) & (!g46) & (sk[96]) & (g88) & (g224) & (g811)) + ((!i_8_) & (g46) & (!sk[96]) & (!g88) & (!g224) & (g811)) + ((!i_8_) & (g46) & (!sk[96]) & (!g88) & (g224) & (g811)) + ((!i_8_) & (g46) & (!sk[96]) & (g88) & (!g224) & (g811)) + ((!i_8_) & (g46) & (!sk[96]) & (g88) & (g224) & (g811)) + ((!i_8_) & (g46) & (sk[96]) & (!g88) & (!g224) & (!g811)) + ((!i_8_) & (g46) & (sk[96]) & (!g88) & (!g224) & (g811)) + ((!i_8_) & (g46) & (sk[96]) & (!g88) & (g224) & (!g811)) + ((!i_8_) & (g46) & (sk[96]) & (!g88) & (g224) & (g811)) + ((!i_8_) & (g46) & (sk[96]) & (g88) & (!g224) & (!g811)) + ((!i_8_) & (g46) & (sk[96]) & (g88) & (!g224) & (g811)) + ((!i_8_) & (g46) & (sk[96]) & (g88) & (g224) & (!g811)) + ((!i_8_) & (g46) & (sk[96]) & (g88) & (g224) & (g811)) + ((i_8_) & (!g46) & (!sk[96]) & (!g88) & (!g224) & (!g811)) + ((i_8_) & (!g46) & (!sk[96]) & (!g88) & (!g224) & (g811)) + ((i_8_) & (!g46) & (!sk[96]) & (!g88) & (g224) & (!g811)) + ((i_8_) & (!g46) & (!sk[96]) & (!g88) & (g224) & (g811)) + ((i_8_) & (!g46) & (!sk[96]) & (g88) & (!g224) & (!g811)) + ((i_8_) & (!g46) & (!sk[96]) & (g88) & (!g224) & (g811)) + ((i_8_) & (!g46) & (!sk[96]) & (g88) & (g224) & (!g811)) + ((i_8_) & (!g46) & (!sk[96]) & (g88) & (g224) & (g811)) + ((i_8_) & (!g46) & (sk[96]) & (!g88) & (!g224) & (!g811)) + ((i_8_) & (!g46) & (sk[96]) & (!g88) & (!g224) & (g811)) + ((i_8_) & (!g46) & (sk[96]) & (!g88) & (g224) & (!g811)) + ((i_8_) & (!g46) & (sk[96]) & (!g88) & (g224) & (g811)) + ((i_8_) & (!g46) & (sk[96]) & (g88) & (!g224) & (!g811)) + ((i_8_) & (g46) & (!sk[96]) & (!g88) & (!g224) & (!g811)) + ((i_8_) & (g46) & (!sk[96]) & (!g88) & (!g224) & (g811)) + ((i_8_) & (g46) & (!sk[96]) & (!g88) & (g224) & (!g811)) + ((i_8_) & (g46) & (!sk[96]) & (!g88) & (g224) & (g811)) + ((i_8_) & (g46) & (!sk[96]) & (g88) & (!g224) & (!g811)) + ((i_8_) & (g46) & (!sk[96]) & (g88) & (!g224) & (g811)) + ((i_8_) & (g46) & (!sk[96]) & (g88) & (g224) & (!g811)) + ((i_8_) & (g46) & (!sk[96]) & (g88) & (g224) & (g811)) + ((i_8_) & (g46) & (sk[96]) & (!g88) & (!g224) & (!g811)) + ((i_8_) & (g46) & (sk[96]) & (!g88) & (!g224) & (g811)) + ((i_8_) & (g46) & (sk[96]) & (!g88) & (g224) & (!g811)) + ((i_8_) & (g46) & (sk[96]) & (!g88) & (g224) & (g811)));
	assign g1103 = (((!sk[97]) & (!i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g124)) + ((!sk[97]) & (!i_14_) & (!i_12_) & (!i_13_) & (g104) & (g124)) + ((!sk[97]) & (!i_14_) & (!i_12_) & (i_13_) & (!g104) & (g124)) + ((!sk[97]) & (!i_14_) & (!i_12_) & (i_13_) & (g104) & (g124)) + ((!sk[97]) & (!i_14_) & (i_12_) & (!i_13_) & (!g104) & (g124)) + ((!sk[97]) & (!i_14_) & (i_12_) & (!i_13_) & (g104) & (g124)) + ((!sk[97]) & (!i_14_) & (i_12_) & (i_13_) & (!g104) & (g124)) + ((!sk[97]) & (!i_14_) & (i_12_) & (i_13_) & (g104) & (g124)) + ((!sk[97]) & (i_14_) & (!i_12_) & (!i_13_) & (!g104) & (!g124)) + ((!sk[97]) & (i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g124)) + ((!sk[97]) & (i_14_) & (!i_12_) & (!i_13_) & (g104) & (!g124)) + ((!sk[97]) & (i_14_) & (!i_12_) & (!i_13_) & (g104) & (g124)) + ((!sk[97]) & (i_14_) & (!i_12_) & (i_13_) & (!g104) & (!g124)) + ((!sk[97]) & (i_14_) & (!i_12_) & (i_13_) & (!g104) & (g124)) + ((!sk[97]) & (i_14_) & (!i_12_) & (i_13_) & (g104) & (!g124)) + ((!sk[97]) & (i_14_) & (!i_12_) & (i_13_) & (g104) & (g124)) + ((!sk[97]) & (i_14_) & (i_12_) & (!i_13_) & (!g104) & (!g124)) + ((!sk[97]) & (i_14_) & (i_12_) & (!i_13_) & (!g104) & (g124)) + ((!sk[97]) & (i_14_) & (i_12_) & (!i_13_) & (g104) & (!g124)) + ((!sk[97]) & (i_14_) & (i_12_) & (!i_13_) & (g104) & (g124)) + ((!sk[97]) & (i_14_) & (i_12_) & (i_13_) & (!g104) & (!g124)) + ((!sk[97]) & (i_14_) & (i_12_) & (i_13_) & (!g104) & (g124)) + ((!sk[97]) & (i_14_) & (i_12_) & (i_13_) & (g104) & (!g124)) + ((!sk[97]) & (i_14_) & (i_12_) & (i_13_) & (g104) & (g124)) + ((sk[97]) & (!i_14_) & (!i_12_) & (!i_13_) & (!g104) & (!g124)) + ((sk[97]) & (!i_14_) & (!i_12_) & (!i_13_) & (g104) & (!g124)) + ((sk[97]) & (!i_14_) & (!i_12_) & (i_13_) & (!g104) & (!g124)) + ((sk[97]) & (!i_14_) & (!i_12_) & (i_13_) & (!g104) & (g124)) + ((sk[97]) & (!i_14_) & (!i_12_) & (i_13_) & (g104) & (!g124)) + ((sk[97]) & (!i_14_) & (!i_12_) & (i_13_) & (g104) & (g124)) + ((sk[97]) & (!i_14_) & (i_12_) & (!i_13_) & (!g104) & (!g124)) + ((sk[97]) & (!i_14_) & (i_12_) & (!i_13_) & (g104) & (!g124)) + ((sk[97]) & (!i_14_) & (i_12_) & (i_13_) & (!g104) & (!g124)) + ((sk[97]) & (i_14_) & (!i_12_) & (!i_13_) & (!g104) & (!g124)) + ((sk[97]) & (i_14_) & (!i_12_) & (i_13_) & (!g104) & (!g124)) + ((sk[97]) & (i_14_) & (i_12_) & (!i_13_) & (!g104) & (!g124)) + ((sk[97]) & (i_14_) & (i_12_) & (!i_13_) & (g104) & (!g124)) + ((sk[97]) & (i_14_) & (i_12_) & (i_13_) & (!g104) & (!g124)) + ((sk[97]) & (i_14_) & (i_12_) & (i_13_) & (!g104) & (g124)));
	assign g1104 = (((!g14) & (!g46) & (!g89) & (!g442) & (!sk[98]) & (g1103)) + ((!g14) & (!g46) & (!g89) & (!g442) & (sk[98]) & (g1103)) + ((!g14) & (!g46) & (!g89) & (g442) & (!sk[98]) & (g1103)) + ((!g14) & (!g46) & (g89) & (!g442) & (!sk[98]) & (g1103)) + ((!g14) & (!g46) & (g89) & (!g442) & (sk[98]) & (!g1103)) + ((!g14) & (!g46) & (g89) & (!g442) & (sk[98]) & (g1103)) + ((!g14) & (!g46) & (g89) & (g442) & (!sk[98]) & (g1103)) + ((!g14) & (g46) & (!g89) & (!g442) & (!sk[98]) & (g1103)) + ((!g14) & (g46) & (!g89) & (g442) & (!sk[98]) & (g1103)) + ((!g14) & (g46) & (g89) & (!g442) & (!sk[98]) & (g1103)) + ((!g14) & (g46) & (g89) & (!g442) & (sk[98]) & (!g1103)) + ((!g14) & (g46) & (g89) & (!g442) & (sk[98]) & (g1103)) + ((!g14) & (g46) & (g89) & (g442) & (!sk[98]) & (g1103)) + ((g14) & (!g46) & (!g89) & (!g442) & (!sk[98]) & (!g1103)) + ((g14) & (!g46) & (!g89) & (!g442) & (!sk[98]) & (g1103)) + ((g14) & (!g46) & (!g89) & (g442) & (!sk[98]) & (!g1103)) + ((g14) & (!g46) & (!g89) & (g442) & (!sk[98]) & (g1103)) + ((g14) & (!g46) & (g89) & (!g442) & (!sk[98]) & (!g1103)) + ((g14) & (!g46) & (g89) & (!g442) & (!sk[98]) & (g1103)) + ((g14) & (!g46) & (g89) & (!g442) & (sk[98]) & (!g1103)) + ((g14) & (!g46) & (g89) & (!g442) & (sk[98]) & (g1103)) + ((g14) & (!g46) & (g89) & (g442) & (!sk[98]) & (!g1103)) + ((g14) & (!g46) & (g89) & (g442) & (!sk[98]) & (g1103)) + ((g14) & (g46) & (!g89) & (!g442) & (!sk[98]) & (!g1103)) + ((g14) & (g46) & (!g89) & (!g442) & (!sk[98]) & (g1103)) + ((g14) & (g46) & (!g89) & (g442) & (!sk[98]) & (!g1103)) + ((g14) & (g46) & (!g89) & (g442) & (!sk[98]) & (g1103)) + ((g14) & (g46) & (g89) & (!g442) & (!sk[98]) & (!g1103)) + ((g14) & (g46) & (g89) & (!g442) & (!sk[98]) & (g1103)) + ((g14) & (g46) & (g89) & (!g442) & (sk[98]) & (!g1103)) + ((g14) & (g46) & (g89) & (!g442) & (sk[98]) & (g1103)) + ((g14) & (g46) & (g89) & (g442) & (!sk[98]) & (!g1103)) + ((g14) & (g46) & (g89) & (g442) & (!sk[98]) & (g1103)));
	assign g1105 = (((g1628) & (!sk[99]) & (!g1622) & (!g1104)) + ((g1628) & (!sk[99]) & (!g1622) & (g1104)) + ((g1628) & (!sk[99]) & (g1622) & (!g1104)) + ((g1628) & (!sk[99]) & (g1622) & (g1104)) + ((g1628) & (sk[99]) & (g1622) & (g1104)));
	assign g1106 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g95) & (g151) & (!g93)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g95) & (g151) & (!g93)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g95) & (g151) & (g93)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g95) & (g151) & (!g93)) + ((!i_14_) & (!i_12_) & (i_13_) & (g95) & (g151) & (!g93)) + ((!i_14_) & (!i_12_) & (i_13_) & (g95) & (g151) & (g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g95) & (g151) & (!g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (g95) & (g151) & (!g93)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g95) & (g151) & (!g93)) + ((i_14_) & (!i_12_) & (!i_13_) & (g95) & (g151) & (!g93)) + ((i_14_) & (!i_12_) & (i_13_) & (!g95) & (g151) & (!g93)) + ((i_14_) & (!i_12_) & (i_13_) & (g95) & (g151) & (!g93)) + ((i_14_) & (i_12_) & (i_13_) & (!g95) & (g151) & (!g93)) + ((i_14_) & (i_12_) & (i_13_) & (g95) & (g151) & (!g93)) + ((i_14_) & (i_12_) & (i_13_) & (g95) & (g151) & (g93)));
	assign g1107 = (((!i_8_) & (!g88) & (g203) & (!sk[101]) & (g475)) + ((!i_8_) & (g88) & (!g203) & (!sk[101]) & (!g475)) + ((!i_8_) & (g88) & (!g203) & (!sk[101]) & (g475)) + ((!i_8_) & (g88) & (!g203) & (sk[101]) & (!g475)) + ((!i_8_) & (g88) & (g203) & (!sk[101]) & (!g475)) + ((!i_8_) & (g88) & (g203) & (!sk[101]) & (g475)) + ((!i_8_) & (g88) & (g203) & (sk[101]) & (!g475)) + ((i_8_) & (!g88) & (g203) & (!sk[101]) & (!g475)) + ((i_8_) & (!g88) & (g203) & (!sk[101]) & (g475)) + ((i_8_) & (g88) & (!g203) & (!sk[101]) & (!g475)) + ((i_8_) & (g88) & (!g203) & (!sk[101]) & (g475)) + ((i_8_) & (g88) & (g203) & (!sk[101]) & (!g475)) + ((i_8_) & (g88) & (g203) & (!sk[101]) & (g475)) + ((i_8_) & (g88) & (g203) & (sk[101]) & (!g475)) + ((i_8_) & (g88) & (g203) & (sk[101]) & (g475)));
	assign g1108 = (((!sk[102]) & (!i_8_) & (!g88) & (!g304) & (!g270) & (g213)) + ((!sk[102]) & (!i_8_) & (!g88) & (!g304) & (g270) & (g213)) + ((!sk[102]) & (!i_8_) & (!g88) & (g304) & (!g270) & (g213)) + ((!sk[102]) & (!i_8_) & (!g88) & (g304) & (g270) & (g213)) + ((!sk[102]) & (!i_8_) & (g88) & (!g304) & (!g270) & (g213)) + ((!sk[102]) & (!i_8_) & (g88) & (!g304) & (g270) & (g213)) + ((!sk[102]) & (!i_8_) & (g88) & (g304) & (!g270) & (g213)) + ((!sk[102]) & (!i_8_) & (g88) & (g304) & (g270) & (g213)) + ((!sk[102]) & (i_8_) & (!g88) & (!g304) & (!g270) & (!g213)) + ((!sk[102]) & (i_8_) & (!g88) & (!g304) & (!g270) & (g213)) + ((!sk[102]) & (i_8_) & (!g88) & (!g304) & (g270) & (!g213)) + ((!sk[102]) & (i_8_) & (!g88) & (!g304) & (g270) & (g213)) + ((!sk[102]) & (i_8_) & (!g88) & (g304) & (!g270) & (!g213)) + ((!sk[102]) & (i_8_) & (!g88) & (g304) & (!g270) & (g213)) + ((!sk[102]) & (i_8_) & (!g88) & (g304) & (g270) & (!g213)) + ((!sk[102]) & (i_8_) & (!g88) & (g304) & (g270) & (g213)) + ((!sk[102]) & (i_8_) & (g88) & (!g304) & (!g270) & (!g213)) + ((!sk[102]) & (i_8_) & (g88) & (!g304) & (!g270) & (g213)) + ((!sk[102]) & (i_8_) & (g88) & (!g304) & (g270) & (!g213)) + ((!sk[102]) & (i_8_) & (g88) & (!g304) & (g270) & (g213)) + ((!sk[102]) & (i_8_) & (g88) & (g304) & (!g270) & (!g213)) + ((!sk[102]) & (i_8_) & (g88) & (g304) & (!g270) & (g213)) + ((!sk[102]) & (i_8_) & (g88) & (g304) & (g270) & (!g213)) + ((!sk[102]) & (i_8_) & (g88) & (g304) & (g270) & (g213)) + ((sk[102]) & (!i_8_) & (g88) & (!g304) & (!g270) & (!g213)) + ((sk[102]) & (!i_8_) & (g88) & (!g304) & (!g270) & (g213)) + ((sk[102]) & (!i_8_) & (g88) & (g304) & (!g270) & (!g213)) + ((sk[102]) & (!i_8_) & (g88) & (g304) & (!g270) & (g213)) + ((sk[102]) & (!i_8_) & (g88) & (g304) & (g270) & (!g213)) + ((sk[102]) & (!i_8_) & (g88) & (g304) & (g270) & (g213)) + ((sk[102]) & (i_8_) & (g88) & (!g304) & (!g270) & (!g213)) + ((sk[102]) & (i_8_) & (g88) & (!g304) & (!g270) & (g213)) + ((sk[102]) & (i_8_) & (g88) & (!g304) & (g270) & (g213)) + ((sk[102]) & (i_8_) & (g88) & (g304) & (!g270) & (!g213)) + ((sk[102]) & (i_8_) & (g88) & (g304) & (!g270) & (g213)) + ((sk[102]) & (i_8_) & (g88) & (g304) & (g270) & (g213)));
	assign g1109 = (((!g89) & (!g93) & (!g572) & (!g849) & (!g1107) & (!g1108)) + ((!g89) & (g93) & (!g572) & (!g849) & (!g1107) & (!g1108)) + ((!g89) & (g93) & (g572) & (!g849) & (!g1107) & (!g1108)) + ((g89) & (!g93) & (!g572) & (!g849) & (!g1107) & (!g1108)) + ((g89) & (!g93) & (g572) & (!g849) & (!g1107) & (!g1108)) + ((g89) & (g93) & (!g572) & (!g849) & (!g1107) & (!g1108)) + ((g89) & (g93) & (g572) & (!g849) & (!g1107) & (!g1108)));
	assign g1110 = (((!g89) & (!g97) & (g678) & (g669) & (!g1106) & (g1109)) + ((g89) & (!g97) & (!g678) & (!g669) & (!g1106) & (g1109)) + ((g89) & (!g97) & (!g678) & (g669) & (!g1106) & (g1109)) + ((g89) & (!g97) & (g678) & (!g669) & (!g1106) & (g1109)) + ((g89) & (!g97) & (g678) & (g669) & (!g1106) & (g1109)));
	assign g1111 = (((!g268) & (!g172) & (!sk[105]) & (!g556) & (!g986) & (g1030)) + ((!g268) & (!g172) & (!sk[105]) & (!g556) & (g986) & (g1030)) + ((!g268) & (!g172) & (!sk[105]) & (g556) & (!g986) & (g1030)) + ((!g268) & (!g172) & (!sk[105]) & (g556) & (g986) & (g1030)) + ((!g268) & (!g172) & (sk[105]) & (g556) & (!g986) & (g1030)) + ((!g268) & (g172) & (!sk[105]) & (!g556) & (!g986) & (g1030)) + ((!g268) & (g172) & (!sk[105]) & (!g556) & (g986) & (g1030)) + ((!g268) & (g172) & (!sk[105]) & (g556) & (!g986) & (g1030)) + ((!g268) & (g172) & (!sk[105]) & (g556) & (g986) & (g1030)) + ((g268) & (!g172) & (!sk[105]) & (!g556) & (!g986) & (!g1030)) + ((g268) & (!g172) & (!sk[105]) & (!g556) & (!g986) & (g1030)) + ((g268) & (!g172) & (!sk[105]) & (!g556) & (g986) & (!g1030)) + ((g268) & (!g172) & (!sk[105]) & (!g556) & (g986) & (g1030)) + ((g268) & (!g172) & (!sk[105]) & (g556) & (!g986) & (!g1030)) + ((g268) & (!g172) & (!sk[105]) & (g556) & (!g986) & (g1030)) + ((g268) & (!g172) & (!sk[105]) & (g556) & (g986) & (!g1030)) + ((g268) & (!g172) & (!sk[105]) & (g556) & (g986) & (g1030)) + ((g268) & (g172) & (!sk[105]) & (!g556) & (!g986) & (!g1030)) + ((g268) & (g172) & (!sk[105]) & (!g556) & (!g986) & (g1030)) + ((g268) & (g172) & (!sk[105]) & (!g556) & (g986) & (!g1030)) + ((g268) & (g172) & (!sk[105]) & (!g556) & (g986) & (g1030)) + ((g268) & (g172) & (!sk[105]) & (g556) & (!g986) & (!g1030)) + ((g268) & (g172) & (!sk[105]) & (g556) & (!g986) & (g1030)) + ((g268) & (g172) & (!sk[105]) & (g556) & (g986) & (!g1030)) + ((g268) & (g172) & (!sk[105]) & (g556) & (g986) & (g1030)));
	assign g1112 = (((!g20) & (!g460) & (!sk[106]) & (g1032) & (g1111)) + ((!g20) & (g460) & (!sk[106]) & (!g1032) & (!g1111)) + ((!g20) & (g460) & (!sk[106]) & (!g1032) & (g1111)) + ((!g20) & (g460) & (!sk[106]) & (g1032) & (!g1111)) + ((!g20) & (g460) & (!sk[106]) & (g1032) & (g1111)) + ((g20) & (!g460) & (!sk[106]) & (g1032) & (!g1111)) + ((g20) & (!g460) & (!sk[106]) & (g1032) & (g1111)) + ((g20) & (!g460) & (sk[106]) & (g1032) & (g1111)) + ((g20) & (g460) & (!sk[106]) & (!g1032) & (!g1111)) + ((g20) & (g460) & (!sk[106]) & (!g1032) & (g1111)) + ((g20) & (g460) & (!sk[106]) & (g1032) & (!g1111)) + ((g20) & (g460) & (!sk[106]) & (g1032) & (g1111)));
	assign g1113 = (((!g204) & (!g548) & (!sk[107]) & (!g881) & (!g1096) & (g1075)) + ((!g204) & (!g548) & (!sk[107]) & (!g881) & (g1096) & (g1075)) + ((!g204) & (!g548) & (!sk[107]) & (g881) & (!g1096) & (g1075)) + ((!g204) & (!g548) & (!sk[107]) & (g881) & (g1096) & (g1075)) + ((!g204) & (g548) & (!sk[107]) & (!g881) & (!g1096) & (g1075)) + ((!g204) & (g548) & (!sk[107]) & (!g881) & (g1096) & (g1075)) + ((!g204) & (g548) & (!sk[107]) & (g881) & (!g1096) & (g1075)) + ((!g204) & (g548) & (!sk[107]) & (g881) & (g1096) & (g1075)) + ((g204) & (!g548) & (!sk[107]) & (!g881) & (!g1096) & (!g1075)) + ((g204) & (!g548) & (!sk[107]) & (!g881) & (!g1096) & (g1075)) + ((g204) & (!g548) & (!sk[107]) & (!g881) & (g1096) & (!g1075)) + ((g204) & (!g548) & (!sk[107]) & (!g881) & (g1096) & (g1075)) + ((g204) & (!g548) & (!sk[107]) & (g881) & (!g1096) & (!g1075)) + ((g204) & (!g548) & (!sk[107]) & (g881) & (!g1096) & (g1075)) + ((g204) & (!g548) & (!sk[107]) & (g881) & (g1096) & (!g1075)) + ((g204) & (!g548) & (!sk[107]) & (g881) & (g1096) & (g1075)) + ((g204) & (!g548) & (sk[107]) & (!g881) & (g1096) & (g1075)) + ((g204) & (g548) & (!sk[107]) & (!g881) & (!g1096) & (!g1075)) + ((g204) & (g548) & (!sk[107]) & (!g881) & (!g1096) & (g1075)) + ((g204) & (g548) & (!sk[107]) & (!g881) & (g1096) & (!g1075)) + ((g204) & (g548) & (!sk[107]) & (!g881) & (g1096) & (g1075)) + ((g204) & (g548) & (!sk[107]) & (g881) & (!g1096) & (!g1075)) + ((g204) & (g548) & (!sk[107]) & (g881) & (!g1096) & (g1075)) + ((g204) & (g548) & (!sk[107]) & (g881) & (g1096) & (!g1075)) + ((g204) & (g548) & (!sk[107]) & (g881) & (g1096) & (g1075)));
	assign g1114 = (((!g181) & (!g123) & (!g670) & (!g671) & (!sk[108]) & (g702)) + ((!g181) & (!g123) & (!g670) & (!g671) & (sk[108]) & (!g702)) + ((!g181) & (!g123) & (!g670) & (g671) & (!sk[108]) & (g702)) + ((!g181) & (!g123) & (g670) & (!g671) & (!sk[108]) & (g702)) + ((!g181) & (!g123) & (g670) & (g671) & (!sk[108]) & (g702)) + ((!g181) & (g123) & (!g670) & (!g671) & (!sk[108]) & (g702)) + ((!g181) & (g123) & (!g670) & (g671) & (!sk[108]) & (g702)) + ((!g181) & (g123) & (g670) & (!g671) & (!sk[108]) & (g702)) + ((!g181) & (g123) & (g670) & (g671) & (!sk[108]) & (g702)) + ((g181) & (!g123) & (!g670) & (!g671) & (!sk[108]) & (!g702)) + ((g181) & (!g123) & (!g670) & (!g671) & (!sk[108]) & (g702)) + ((g181) & (!g123) & (!g670) & (g671) & (!sk[108]) & (!g702)) + ((g181) & (!g123) & (!g670) & (g671) & (!sk[108]) & (g702)) + ((g181) & (!g123) & (g670) & (!g671) & (!sk[108]) & (!g702)) + ((g181) & (!g123) & (g670) & (!g671) & (!sk[108]) & (g702)) + ((g181) & (!g123) & (g670) & (g671) & (!sk[108]) & (!g702)) + ((g181) & (!g123) & (g670) & (g671) & (!sk[108]) & (g702)) + ((g181) & (g123) & (!g670) & (!g671) & (!sk[108]) & (!g702)) + ((g181) & (g123) & (!g670) & (!g671) & (!sk[108]) & (g702)) + ((g181) & (g123) & (!g670) & (g671) & (!sk[108]) & (!g702)) + ((g181) & (g123) & (!g670) & (g671) & (!sk[108]) & (g702)) + ((g181) & (g123) & (g670) & (!g671) & (!sk[108]) & (!g702)) + ((g181) & (g123) & (g670) & (!g671) & (!sk[108]) & (g702)) + ((g181) & (g123) & (g670) & (g671) & (!sk[108]) & (!g702)) + ((g181) & (g123) & (g670) & (g671) & (!sk[108]) & (g702)));
	assign g1115 = (((!g10) & (!g45) & (!g221) & (!sk[109]) & (!g187) & (g1114)) + ((!g10) & (!g45) & (!g221) & (!sk[109]) & (g187) & (g1114)) + ((!g10) & (!g45) & (g221) & (!sk[109]) & (!g187) & (g1114)) + ((!g10) & (!g45) & (g221) & (!sk[109]) & (g187) & (g1114)) + ((!g10) & (!g45) & (g221) & (sk[109]) & (!g187) & (g1114)) + ((!g10) & (g45) & (!g221) & (!sk[109]) & (!g187) & (g1114)) + ((!g10) & (g45) & (!g221) & (!sk[109]) & (g187) & (g1114)) + ((!g10) & (g45) & (g221) & (!sk[109]) & (!g187) & (g1114)) + ((!g10) & (g45) & (g221) & (!sk[109]) & (g187) & (g1114)) + ((g10) & (!g45) & (!g221) & (!sk[109]) & (!g187) & (!g1114)) + ((g10) & (!g45) & (!g221) & (!sk[109]) & (!g187) & (g1114)) + ((g10) & (!g45) & (!g221) & (!sk[109]) & (g187) & (!g1114)) + ((g10) & (!g45) & (!g221) & (!sk[109]) & (g187) & (g1114)) + ((g10) & (!g45) & (g221) & (!sk[109]) & (!g187) & (!g1114)) + ((g10) & (!g45) & (g221) & (!sk[109]) & (!g187) & (g1114)) + ((g10) & (!g45) & (g221) & (!sk[109]) & (g187) & (!g1114)) + ((g10) & (!g45) & (g221) & (!sk[109]) & (g187) & (g1114)) + ((g10) & (g45) & (!g221) & (!sk[109]) & (!g187) & (!g1114)) + ((g10) & (g45) & (!g221) & (!sk[109]) & (!g187) & (g1114)) + ((g10) & (g45) & (!g221) & (!sk[109]) & (g187) & (!g1114)) + ((g10) & (g45) & (!g221) & (!sk[109]) & (g187) & (g1114)) + ((g10) & (g45) & (g221) & (!sk[109]) & (!g187) & (!g1114)) + ((g10) & (g45) & (g221) & (!sk[109]) & (!g187) & (g1114)) + ((g10) & (g45) & (g221) & (!sk[109]) & (g187) & (!g1114)) + ((g10) & (g45) & (g221) & (!sk[109]) & (g187) & (g1114)));
	assign g1116 = (((!sk[110]) & (!i_8_) & (!g88) & (!g534) & (!g979) & (g980)) + ((!sk[110]) & (!i_8_) & (!g88) & (!g534) & (g979) & (g980)) + ((!sk[110]) & (!i_8_) & (!g88) & (g534) & (!g979) & (g980)) + ((!sk[110]) & (!i_8_) & (!g88) & (g534) & (g979) & (g980)) + ((!sk[110]) & (!i_8_) & (g88) & (!g534) & (!g979) & (g980)) + ((!sk[110]) & (!i_8_) & (g88) & (!g534) & (g979) & (g980)) + ((!sk[110]) & (!i_8_) & (g88) & (g534) & (!g979) & (g980)) + ((!sk[110]) & (!i_8_) & (g88) & (g534) & (g979) & (g980)) + ((!sk[110]) & (i_8_) & (!g88) & (!g534) & (!g979) & (!g980)) + ((!sk[110]) & (i_8_) & (!g88) & (!g534) & (!g979) & (g980)) + ((!sk[110]) & (i_8_) & (!g88) & (!g534) & (g979) & (!g980)) + ((!sk[110]) & (i_8_) & (!g88) & (!g534) & (g979) & (g980)) + ((!sk[110]) & (i_8_) & (!g88) & (g534) & (!g979) & (!g980)) + ((!sk[110]) & (i_8_) & (!g88) & (g534) & (!g979) & (g980)) + ((!sk[110]) & (i_8_) & (!g88) & (g534) & (g979) & (!g980)) + ((!sk[110]) & (i_8_) & (!g88) & (g534) & (g979) & (g980)) + ((!sk[110]) & (i_8_) & (g88) & (!g534) & (!g979) & (!g980)) + ((!sk[110]) & (i_8_) & (g88) & (!g534) & (!g979) & (g980)) + ((!sk[110]) & (i_8_) & (g88) & (!g534) & (g979) & (!g980)) + ((!sk[110]) & (i_8_) & (g88) & (!g534) & (g979) & (g980)) + ((!sk[110]) & (i_8_) & (g88) & (g534) & (!g979) & (!g980)) + ((!sk[110]) & (i_8_) & (g88) & (g534) & (!g979) & (g980)) + ((!sk[110]) & (i_8_) & (g88) & (g534) & (g979) & (!g980)) + ((!sk[110]) & (i_8_) & (g88) & (g534) & (g979) & (g980)) + ((sk[110]) & (!i_8_) & (!g88) & (!g534) & (!g979) & (!g980)) + ((sk[110]) & (!i_8_) & (!g88) & (!g534) & (!g979) & (g980)) + ((sk[110]) & (!i_8_) & (!g88) & (!g534) & (g979) & (!g980)) + ((sk[110]) & (!i_8_) & (!g88) & (!g534) & (g979) & (g980)) + ((sk[110]) & (!i_8_) & (!g88) & (g534) & (!g979) & (!g980)) + ((sk[110]) & (!i_8_) & (!g88) & (g534) & (!g979) & (g980)) + ((sk[110]) & (!i_8_) & (!g88) & (g534) & (g979) & (!g980)) + ((sk[110]) & (!i_8_) & (!g88) & (g534) & (g979) & (g980)) + ((sk[110]) & (!i_8_) & (g88) & (!g534) & (g979) & (g980)) + ((sk[110]) & (i_8_) & (!g88) & (!g534) & (!g979) & (!g980)) + ((sk[110]) & (i_8_) & (!g88) & (!g534) & (!g979) & (g980)) + ((sk[110]) & (i_8_) & (!g88) & (!g534) & (g979) & (!g980)) + ((sk[110]) & (i_8_) & (!g88) & (!g534) & (g979) & (g980)) + ((sk[110]) & (i_8_) & (!g88) & (g534) & (!g979) & (!g980)) + ((sk[110]) & (i_8_) & (!g88) & (g534) & (!g979) & (g980)) + ((sk[110]) & (i_8_) & (!g88) & (g534) & (g979) & (!g980)) + ((sk[110]) & (i_8_) & (!g88) & (g534) & (g979) & (g980)) + ((sk[110]) & (i_8_) & (g88) & (!g534) & (g979) & (g980)) + ((sk[110]) & (i_8_) & (g88) & (g534) & (g979) & (g980)));
	assign g1117 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g102) & (!sk[111]) & (g115)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g102) & (!sk[111]) & (g115)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g102) & (!sk[111]) & (g115)) + ((!i_14_) & (!i_12_) & (i_13_) & (g102) & (!sk[111]) & (g115)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g102) & (!sk[111]) & (g115)) + ((!i_14_) & (i_12_) & (!i_13_) & (g102) & (!sk[111]) & (g115)) + ((!i_14_) & (i_12_) & (i_13_) & (!g102) & (!sk[111]) & (g115)) + ((!i_14_) & (i_12_) & (i_13_) & (!g102) & (sk[111]) & (!g115)) + ((!i_14_) & (i_12_) & (i_13_) & (g102) & (!sk[111]) & (g115)) + ((!i_14_) & (i_12_) & (i_13_) & (g102) & (sk[111]) & (!g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g102) & (!sk[111]) & (!g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g102) & (!sk[111]) & (g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g102) & (sk[111]) & (!g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g102) & (sk[111]) & (g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (g102) & (!sk[111]) & (!g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (g102) & (!sk[111]) & (g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (g102) & (sk[111]) & (!g115)) + ((i_14_) & (!i_12_) & (i_13_) & (!g102) & (!sk[111]) & (!g115)) + ((i_14_) & (!i_12_) & (i_13_) & (!g102) & (!sk[111]) & (g115)) + ((i_14_) & (!i_12_) & (i_13_) & (!g102) & (sk[111]) & (!g115)) + ((i_14_) & (!i_12_) & (i_13_) & (!g102) & (sk[111]) & (g115)) + ((i_14_) & (!i_12_) & (i_13_) & (g102) & (!sk[111]) & (!g115)) + ((i_14_) & (!i_12_) & (i_13_) & (g102) & (!sk[111]) & (g115)) + ((i_14_) & (!i_12_) & (i_13_) & (g102) & (sk[111]) & (!g115)) + ((i_14_) & (i_12_) & (!i_13_) & (!g102) & (!sk[111]) & (!g115)) + ((i_14_) & (i_12_) & (!i_13_) & (!g102) & (!sk[111]) & (g115)) + ((i_14_) & (i_12_) & (!i_13_) & (g102) & (!sk[111]) & (!g115)) + ((i_14_) & (i_12_) & (!i_13_) & (g102) & (!sk[111]) & (g115)) + ((i_14_) & (i_12_) & (i_13_) & (!g102) & (!sk[111]) & (!g115)) + ((i_14_) & (i_12_) & (i_13_) & (!g102) & (!sk[111]) & (g115)) + ((i_14_) & (i_12_) & (i_13_) & (!g102) & (sk[111]) & (!g115)) + ((i_14_) & (i_12_) & (i_13_) & (!g102) & (sk[111]) & (g115)) + ((i_14_) & (i_12_) & (i_13_) & (g102) & (!sk[111]) & (!g115)) + ((i_14_) & (i_12_) & (i_13_) & (g102) & (!sk[111]) & (g115)));
	assign g1118 = (((!i_8_) & (!g88) & (!g232) & (!sk[112]) & (!g116) & (g675)) + ((!i_8_) & (!g88) & (!g232) & (!sk[112]) & (g116) & (g675)) + ((!i_8_) & (!g88) & (!g232) & (sk[112]) & (!g116) & (!g675)) + ((!i_8_) & (!g88) & (!g232) & (sk[112]) & (!g116) & (g675)) + ((!i_8_) & (!g88) & (!g232) & (sk[112]) & (g116) & (!g675)) + ((!i_8_) & (!g88) & (!g232) & (sk[112]) & (g116) & (g675)) + ((!i_8_) & (!g88) & (g232) & (!sk[112]) & (!g116) & (g675)) + ((!i_8_) & (!g88) & (g232) & (!sk[112]) & (g116) & (g675)) + ((!i_8_) & (!g88) & (g232) & (sk[112]) & (!g116) & (!g675)) + ((!i_8_) & (!g88) & (g232) & (sk[112]) & (!g116) & (g675)) + ((!i_8_) & (!g88) & (g232) & (sk[112]) & (g116) & (!g675)) + ((!i_8_) & (!g88) & (g232) & (sk[112]) & (g116) & (g675)) + ((!i_8_) & (g88) & (!g232) & (!sk[112]) & (!g116) & (g675)) + ((!i_8_) & (g88) & (!g232) & (!sk[112]) & (g116) & (g675)) + ((!i_8_) & (g88) & (!g232) & (sk[112]) & (!g116) & (!g675)) + ((!i_8_) & (g88) & (g232) & (!sk[112]) & (!g116) & (g675)) + ((!i_8_) & (g88) & (g232) & (!sk[112]) & (g116) & (g675)) + ((i_8_) & (!g88) & (!g232) & (!sk[112]) & (!g116) & (!g675)) + ((i_8_) & (!g88) & (!g232) & (!sk[112]) & (!g116) & (g675)) + ((i_8_) & (!g88) & (!g232) & (!sk[112]) & (g116) & (!g675)) + ((i_8_) & (!g88) & (!g232) & (!sk[112]) & (g116) & (g675)) + ((i_8_) & (!g88) & (!g232) & (sk[112]) & (!g116) & (!g675)) + ((i_8_) & (!g88) & (!g232) & (sk[112]) & (!g116) & (g675)) + ((i_8_) & (!g88) & (!g232) & (sk[112]) & (g116) & (!g675)) + ((i_8_) & (!g88) & (!g232) & (sk[112]) & (g116) & (g675)) + ((i_8_) & (!g88) & (g232) & (!sk[112]) & (!g116) & (!g675)) + ((i_8_) & (!g88) & (g232) & (!sk[112]) & (!g116) & (g675)) + ((i_8_) & (!g88) & (g232) & (!sk[112]) & (g116) & (!g675)) + ((i_8_) & (!g88) & (g232) & (!sk[112]) & (g116) & (g675)) + ((i_8_) & (!g88) & (g232) & (sk[112]) & (!g116) & (!g675)) + ((i_8_) & (!g88) & (g232) & (sk[112]) & (!g116) & (g675)) + ((i_8_) & (!g88) & (g232) & (sk[112]) & (g116) & (!g675)) + ((i_8_) & (!g88) & (g232) & (sk[112]) & (g116) & (g675)) + ((i_8_) & (g88) & (!g232) & (!sk[112]) & (!g116) & (!g675)) + ((i_8_) & (g88) & (!g232) & (!sk[112]) & (!g116) & (g675)) + ((i_8_) & (g88) & (!g232) & (!sk[112]) & (g116) & (!g675)) + ((i_8_) & (g88) & (!g232) & (!sk[112]) & (g116) & (g675)) + ((i_8_) & (g88) & (!g232) & (sk[112]) & (!g116) & (!g675)) + ((i_8_) & (g88) & (!g232) & (sk[112]) & (!g116) & (g675)) + ((i_8_) & (g88) & (!g232) & (sk[112]) & (g116) & (!g675)) + ((i_8_) & (g88) & (!g232) & (sk[112]) & (g116) & (g675)) + ((i_8_) & (g88) & (g232) & (!sk[112]) & (!g116) & (!g675)) + ((i_8_) & (g88) & (g232) & (!sk[112]) & (!g116) & (g675)) + ((i_8_) & (g88) & (g232) & (!sk[112]) & (g116) & (!g675)) + ((i_8_) & (g88) & (g232) & (!sk[112]) & (g116) & (g675)));
	assign g1119 = (((!sk[113]) & (!g89) & (!g1112) & (!g1113) & (!g1115) & (g1616)) + ((!sk[113]) & (!g89) & (!g1112) & (!g1113) & (g1115) & (g1616)) + ((!sk[113]) & (!g89) & (!g1112) & (g1113) & (!g1115) & (g1616)) + ((!sk[113]) & (!g89) & (!g1112) & (g1113) & (g1115) & (g1616)) + ((!sk[113]) & (!g89) & (g1112) & (!g1113) & (!g1115) & (g1616)) + ((!sk[113]) & (!g89) & (g1112) & (!g1113) & (g1115) & (g1616)) + ((!sk[113]) & (!g89) & (g1112) & (g1113) & (!g1115) & (g1616)) + ((!sk[113]) & (!g89) & (g1112) & (g1113) & (g1115) & (g1616)) + ((!sk[113]) & (g89) & (!g1112) & (!g1113) & (!g1115) & (!g1616)) + ((!sk[113]) & (g89) & (!g1112) & (!g1113) & (!g1115) & (g1616)) + ((!sk[113]) & (g89) & (!g1112) & (!g1113) & (g1115) & (!g1616)) + ((!sk[113]) & (g89) & (!g1112) & (!g1113) & (g1115) & (g1616)) + ((!sk[113]) & (g89) & (!g1112) & (g1113) & (!g1115) & (!g1616)) + ((!sk[113]) & (g89) & (!g1112) & (g1113) & (!g1115) & (g1616)) + ((!sk[113]) & (g89) & (!g1112) & (g1113) & (g1115) & (!g1616)) + ((!sk[113]) & (g89) & (!g1112) & (g1113) & (g1115) & (g1616)) + ((!sk[113]) & (g89) & (g1112) & (!g1113) & (!g1115) & (!g1616)) + ((!sk[113]) & (g89) & (g1112) & (!g1113) & (!g1115) & (g1616)) + ((!sk[113]) & (g89) & (g1112) & (!g1113) & (g1115) & (!g1616)) + ((!sk[113]) & (g89) & (g1112) & (!g1113) & (g1115) & (g1616)) + ((!sk[113]) & (g89) & (g1112) & (g1113) & (!g1115) & (!g1616)) + ((!sk[113]) & (g89) & (g1112) & (g1113) & (!g1115) & (g1616)) + ((!sk[113]) & (g89) & (g1112) & (g1113) & (g1115) & (!g1616)) + ((!sk[113]) & (g89) & (g1112) & (g1113) & (g1115) & (g1616)) + ((sk[113]) & (!g89) & (g1112) & (g1113) & (g1115) & (g1616)) + ((sk[113]) & (g89) & (!g1112) & (!g1113) & (!g1115) & (g1616)) + ((sk[113]) & (g89) & (!g1112) & (!g1113) & (g1115) & (g1616)) + ((sk[113]) & (g89) & (!g1112) & (g1113) & (!g1115) & (g1616)) + ((sk[113]) & (g89) & (!g1112) & (g1113) & (g1115) & (g1616)) + ((sk[113]) & (g89) & (g1112) & (!g1113) & (!g1115) & (g1616)) + ((sk[113]) & (g89) & (g1112) & (!g1113) & (g1115) & (g1616)) + ((sk[113]) & (g89) & (g1112) & (g1113) & (!g1115) & (g1616)) + ((sk[113]) & (g89) & (g1112) & (g1113) & (g1115) & (g1616)));
	assign g1120 = (((!sk[114]) & (!g115) & (!g554) & (g460) & (g711)) + ((!sk[114]) & (!g115) & (g554) & (!g460) & (!g711)) + ((!sk[114]) & (!g115) & (g554) & (!g460) & (g711)) + ((!sk[114]) & (!g115) & (g554) & (g460) & (!g711)) + ((!sk[114]) & (!g115) & (g554) & (g460) & (g711)) + ((!sk[114]) & (g115) & (!g554) & (g460) & (!g711)) + ((!sk[114]) & (g115) & (!g554) & (g460) & (g711)) + ((!sk[114]) & (g115) & (g554) & (!g460) & (!g711)) + ((!sk[114]) & (g115) & (g554) & (!g460) & (g711)) + ((!sk[114]) & (g115) & (g554) & (g460) & (!g711)) + ((!sk[114]) & (g115) & (g554) & (g460) & (g711)) + ((sk[114]) & (!g115) & (!g554) & (!g460) & (!g711)) + ((sk[114]) & (g115) & (!g554) & (!g460) & (!g711)) + ((sk[114]) & (g115) & (!g554) & (!g460) & (g711)));
	assign g1121 = (((!g253) & (!g710) & (!g1026) & (sk[115]) & (g1120)) + ((!g253) & (!g710) & (g1026) & (!sk[115]) & (g1120)) + ((!g253) & (g710) & (!g1026) & (!sk[115]) & (!g1120)) + ((!g253) & (g710) & (!g1026) & (!sk[115]) & (g1120)) + ((!g253) & (g710) & (g1026) & (!sk[115]) & (!g1120)) + ((!g253) & (g710) & (g1026) & (!sk[115]) & (g1120)) + ((g253) & (!g710) & (g1026) & (!sk[115]) & (!g1120)) + ((g253) & (!g710) & (g1026) & (!sk[115]) & (g1120)) + ((g253) & (g710) & (!g1026) & (!sk[115]) & (!g1120)) + ((g253) & (g710) & (!g1026) & (!sk[115]) & (g1120)) + ((g253) & (g710) & (g1026) & (!sk[115]) & (!g1120)) + ((g253) & (g710) & (g1026) & (!sk[115]) & (g1120)));
	assign g1122 = (((!g44) & (!g191) & (sk[116]) & (!g641)) + ((g44) & (!g191) & (!sk[116]) & (!g641)) + ((g44) & (!g191) & (!sk[116]) & (g641)) + ((g44) & (g191) & (!sk[116]) & (!g641)) + ((g44) & (g191) & (!sk[116]) & (g641)));
	assign g1123 = (((!g6) & (!i_15_) & (!i_14_) & (i_12_) & (i_13_) & (!g122)) + ((!g6) & (!i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (!g122)) + ((!g6) & (!i_15_) & (i_14_) & (!i_12_) & (i_13_) & (!g122)) + ((!g6) & (i_15_) & (!i_14_) & (i_12_) & (i_13_) & (!g122)) + ((!g6) & (i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (!g122)) + ((!g6) & (i_15_) & (i_14_) & (!i_12_) & (i_13_) & (!g122)) + ((g6) & (!i_15_) & (!i_14_) & (i_12_) & (i_13_) & (!g122)) + ((g6) & (!i_15_) & (!i_14_) & (i_12_) & (i_13_) & (g122)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (!g122)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (i_13_) & (!g122)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (!i_13_) & (!g122)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (!i_13_) & (g122)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (i_13_) & (!g122)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (!g122)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (i_13_) & (!g122)) + ((g6) & (i_15_) & (i_14_) & (i_12_) & (i_13_) & (!g122)) + ((g6) & (i_15_) & (i_14_) & (i_12_) & (i_13_) & (g122)));
	assign g1124 = (((!i_9_) & (!i_10_) & (!sk[118]) & (!g7) & (!g53) & (g91)) + ((!i_9_) & (!i_10_) & (!sk[118]) & (!g7) & (g53) & (g91)) + ((!i_9_) & (!i_10_) & (!sk[118]) & (g7) & (!g53) & (g91)) + ((!i_9_) & (!i_10_) & (!sk[118]) & (g7) & (g53) & (g91)) + ((!i_9_) & (i_10_) & (!sk[118]) & (!g7) & (!g53) & (g91)) + ((!i_9_) & (i_10_) & (!sk[118]) & (!g7) & (g53) & (g91)) + ((!i_9_) & (i_10_) & (!sk[118]) & (g7) & (!g53) & (g91)) + ((!i_9_) & (i_10_) & (!sk[118]) & (g7) & (g53) & (g91)) + ((!i_9_) & (i_10_) & (sk[118]) & (!g7) & (g53) & (!g91)) + ((!i_9_) & (i_10_) & (sk[118]) & (g7) & (g53) & (!g91)) + ((!i_9_) & (i_10_) & (sk[118]) & (g7) & (g53) & (g91)) + ((i_9_) & (!i_10_) & (!sk[118]) & (!g7) & (!g53) & (!g91)) + ((i_9_) & (!i_10_) & (!sk[118]) & (!g7) & (!g53) & (g91)) + ((i_9_) & (!i_10_) & (!sk[118]) & (!g7) & (g53) & (!g91)) + ((i_9_) & (!i_10_) & (!sk[118]) & (!g7) & (g53) & (g91)) + ((i_9_) & (!i_10_) & (!sk[118]) & (g7) & (!g53) & (!g91)) + ((i_9_) & (!i_10_) & (!sk[118]) & (g7) & (!g53) & (g91)) + ((i_9_) & (!i_10_) & (!sk[118]) & (g7) & (g53) & (!g91)) + ((i_9_) & (!i_10_) & (!sk[118]) & (g7) & (g53) & (g91)) + ((i_9_) & (!i_10_) & (sk[118]) & (g7) & (g53) & (!g91)) + ((i_9_) & (!i_10_) & (sk[118]) & (g7) & (g53) & (g91)) + ((i_9_) & (i_10_) & (!sk[118]) & (!g7) & (!g53) & (!g91)) + ((i_9_) & (i_10_) & (!sk[118]) & (!g7) & (!g53) & (g91)) + ((i_9_) & (i_10_) & (!sk[118]) & (!g7) & (g53) & (!g91)) + ((i_9_) & (i_10_) & (!sk[118]) & (!g7) & (g53) & (g91)) + ((i_9_) & (i_10_) & (!sk[118]) & (g7) & (!g53) & (!g91)) + ((i_9_) & (i_10_) & (!sk[118]) & (g7) & (!g53) & (g91)) + ((i_9_) & (i_10_) & (!sk[118]) & (g7) & (g53) & (!g91)) + ((i_9_) & (i_10_) & (!sk[118]) & (g7) & (g53) & (g91)) + ((i_9_) & (i_10_) & (sk[118]) & (g7) & (g53) & (!g91)) + ((i_9_) & (i_10_) & (sk[118]) & (g7) & (g53) & (g91)));
	assign g1125 = (((!g1076) & (!g1122) & (g1123) & (!sk[119]) & (g1124)) + ((!g1076) & (g1122) & (!g1123) & (!sk[119]) & (!g1124)) + ((!g1076) & (g1122) & (!g1123) & (!sk[119]) & (g1124)) + ((!g1076) & (g1122) & (!g1123) & (sk[119]) & (!g1124)) + ((!g1076) & (g1122) & (g1123) & (!sk[119]) & (!g1124)) + ((!g1076) & (g1122) & (g1123) & (!sk[119]) & (g1124)) + ((g1076) & (!g1122) & (g1123) & (!sk[119]) & (!g1124)) + ((g1076) & (!g1122) & (g1123) & (!sk[119]) & (g1124)) + ((g1076) & (g1122) & (!g1123) & (!sk[119]) & (!g1124)) + ((g1076) & (g1122) & (!g1123) & (!sk[119]) & (g1124)) + ((g1076) & (g1122) & (g1123) & (!sk[119]) & (!g1124)) + ((g1076) & (g1122) & (g1123) & (!sk[119]) & (g1124)));
	assign g1126 = (((!sk[120]) & (!i_8_) & (!g88) & (!g1084) & (!g1121) & (g1125)) + ((!sk[120]) & (!i_8_) & (!g88) & (!g1084) & (g1121) & (g1125)) + ((!sk[120]) & (!i_8_) & (!g88) & (g1084) & (!g1121) & (g1125)) + ((!sk[120]) & (!i_8_) & (!g88) & (g1084) & (g1121) & (g1125)) + ((!sk[120]) & (!i_8_) & (g88) & (!g1084) & (!g1121) & (g1125)) + ((!sk[120]) & (!i_8_) & (g88) & (!g1084) & (g1121) & (g1125)) + ((!sk[120]) & (!i_8_) & (g88) & (g1084) & (!g1121) & (g1125)) + ((!sk[120]) & (!i_8_) & (g88) & (g1084) & (g1121) & (g1125)) + ((!sk[120]) & (i_8_) & (!g88) & (!g1084) & (!g1121) & (!g1125)) + ((!sk[120]) & (i_8_) & (!g88) & (!g1084) & (!g1121) & (g1125)) + ((!sk[120]) & (i_8_) & (!g88) & (!g1084) & (g1121) & (!g1125)) + ((!sk[120]) & (i_8_) & (!g88) & (!g1084) & (g1121) & (g1125)) + ((!sk[120]) & (i_8_) & (!g88) & (g1084) & (!g1121) & (!g1125)) + ((!sk[120]) & (i_8_) & (!g88) & (g1084) & (!g1121) & (g1125)) + ((!sk[120]) & (i_8_) & (!g88) & (g1084) & (g1121) & (!g1125)) + ((!sk[120]) & (i_8_) & (!g88) & (g1084) & (g1121) & (g1125)) + ((!sk[120]) & (i_8_) & (g88) & (!g1084) & (!g1121) & (!g1125)) + ((!sk[120]) & (i_8_) & (g88) & (!g1084) & (!g1121) & (g1125)) + ((!sk[120]) & (i_8_) & (g88) & (!g1084) & (g1121) & (!g1125)) + ((!sk[120]) & (i_8_) & (g88) & (!g1084) & (g1121) & (g1125)) + ((!sk[120]) & (i_8_) & (g88) & (g1084) & (!g1121) & (!g1125)) + ((!sk[120]) & (i_8_) & (g88) & (g1084) & (!g1121) & (g1125)) + ((!sk[120]) & (i_8_) & (g88) & (g1084) & (g1121) & (!g1125)) + ((!sk[120]) & (i_8_) & (g88) & (g1084) & (g1121) & (g1125)) + ((sk[120]) & (!i_8_) & (g88) & (!g1084) & (!g1121) & (!g1125)) + ((sk[120]) & (!i_8_) & (g88) & (!g1084) & (g1121) & (!g1125)) + ((sk[120]) & (!i_8_) & (g88) & (g1084) & (!g1121) & (!g1125)) + ((sk[120]) & (!i_8_) & (g88) & (g1084) & (g1121) & (!g1125)) + ((sk[120]) & (i_8_) & (g88) & (!g1084) & (!g1121) & (!g1125)) + ((sk[120]) & (i_8_) & (g88) & (!g1084) & (!g1121) & (g1125)) + ((sk[120]) & (i_8_) & (g88) & (!g1084) & (g1121) & (!g1125)) + ((sk[120]) & (i_8_) & (g88) & (!g1084) & (g1121) & (g1125)) + ((sk[120]) & (i_8_) & (g88) & (g1084) & (!g1121) & (!g1125)) + ((sk[120]) & (i_8_) & (g88) & (g1084) & (!g1121) & (g1125)) + ((sk[120]) & (i_8_) & (g88) & (g1084) & (g1121) & (!g1125)));
	assign g1127 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g119) & (!sk[121]) & (g122)) + ((!i_14_) & (!i_12_) & (!i_13_) & (!g119) & (sk[121]) & (!g122)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g119) & (!sk[121]) & (g122)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g119) & (sk[121]) & (!g122)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g119) & (!sk[121]) & (g122)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g119) & (sk[121]) & (!g122)) + ((!i_14_) & (!i_12_) & (i_13_) & (g119) & (!sk[121]) & (g122)) + ((!i_14_) & (!i_12_) & (i_13_) & (g119) & (sk[121]) & (!g122)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g119) & (!sk[121]) & (g122)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g119) & (sk[121]) & (!g122)) + ((!i_14_) & (i_12_) & (!i_13_) & (g119) & (!sk[121]) & (g122)) + ((!i_14_) & (i_12_) & (!i_13_) & (g119) & (sk[121]) & (!g122)) + ((!i_14_) & (i_12_) & (i_13_) & (!g119) & (!sk[121]) & (g122)) + ((!i_14_) & (i_12_) & (i_13_) & (g119) & (!sk[121]) & (g122)) + ((!i_14_) & (i_12_) & (i_13_) & (g119) & (sk[121]) & (!g122)) + ((!i_14_) & (i_12_) & (i_13_) & (g119) & (sk[121]) & (g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g119) & (!sk[121]) & (!g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g119) & (!sk[121]) & (g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (g119) & (!sk[121]) & (!g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (g119) & (!sk[121]) & (g122)) + ((i_14_) & (!i_12_) & (i_13_) & (!g119) & (!sk[121]) & (!g122)) + ((i_14_) & (!i_12_) & (i_13_) & (!g119) & (!sk[121]) & (g122)) + ((i_14_) & (!i_12_) & (i_13_) & (g119) & (!sk[121]) & (!g122)) + ((i_14_) & (!i_12_) & (i_13_) & (g119) & (!sk[121]) & (g122)) + ((i_14_) & (i_12_) & (!i_13_) & (!g119) & (!sk[121]) & (!g122)) + ((i_14_) & (i_12_) & (!i_13_) & (!g119) & (!sk[121]) & (g122)) + ((i_14_) & (i_12_) & (!i_13_) & (g119) & (!sk[121]) & (!g122)) + ((i_14_) & (i_12_) & (!i_13_) & (g119) & (!sk[121]) & (g122)) + ((i_14_) & (i_12_) & (!i_13_) & (g119) & (sk[121]) & (!g122)) + ((i_14_) & (i_12_) & (!i_13_) & (g119) & (sk[121]) & (g122)) + ((i_14_) & (i_12_) & (i_13_) & (!g119) & (!sk[121]) & (!g122)) + ((i_14_) & (i_12_) & (i_13_) & (!g119) & (!sk[121]) & (g122)) + ((i_14_) & (i_12_) & (i_13_) & (!g119) & (sk[121]) & (!g122)) + ((i_14_) & (i_12_) & (i_13_) & (g119) & (!sk[121]) & (!g122)) + ((i_14_) & (i_12_) & (i_13_) & (g119) & (!sk[121]) & (g122)) + ((i_14_) & (i_12_) & (i_13_) & (g119) & (sk[121]) & (!g122)));
	assign g1128 = (((!i_8_) & (g88) & (!g349) & (!g670) & (g704) & (!g895)) + ((!i_8_) & (g88) & (!g349) & (!g670) & (g704) & (g895)) + ((!i_8_) & (g88) & (!g349) & (g670) & (g704) & (!g895)) + ((!i_8_) & (g88) & (!g349) & (g670) & (g704) & (g895)) + ((!i_8_) & (g88) & (g349) & (!g670) & (!g704) & (!g895)) + ((!i_8_) & (g88) & (g349) & (!g670) & (!g704) & (g895)) + ((!i_8_) & (g88) & (g349) & (!g670) & (g704) & (!g895)) + ((!i_8_) & (g88) & (g349) & (!g670) & (g704) & (g895)) + ((!i_8_) & (g88) & (g349) & (g670) & (!g704) & (!g895)) + ((!i_8_) & (g88) & (g349) & (g670) & (!g704) & (g895)) + ((!i_8_) & (g88) & (g349) & (g670) & (g704) & (!g895)) + ((!i_8_) & (g88) & (g349) & (g670) & (g704) & (g895)) + ((i_8_) & (g88) & (!g349) & (!g670) & (!g704) & (g895)) + ((i_8_) & (g88) & (!g349) & (!g670) & (g704) & (g895)) + ((i_8_) & (g88) & (!g349) & (g670) & (!g704) & (!g895)) + ((i_8_) & (g88) & (!g349) & (g670) & (!g704) & (g895)) + ((i_8_) & (g88) & (!g349) & (g670) & (g704) & (!g895)) + ((i_8_) & (g88) & (!g349) & (g670) & (g704) & (g895)) + ((i_8_) & (g88) & (g349) & (!g670) & (!g704) & (!g895)) + ((i_8_) & (g88) & (g349) & (!g670) & (!g704) & (g895)) + ((i_8_) & (g88) & (g349) & (!g670) & (g704) & (!g895)) + ((i_8_) & (g88) & (g349) & (!g670) & (g704) & (g895)) + ((i_8_) & (g88) & (g349) & (g670) & (!g704) & (!g895)) + ((i_8_) & (g88) & (g349) & (g670) & (!g704) & (g895)) + ((i_8_) & (g88) & (g349) & (g670) & (g704) & (!g895)) + ((i_8_) & (g88) & (g349) & (g670) & (g704) & (g895)));
	assign g1129 = (((!i_8_) & (!g88) & (!g181) & (!g183) & (!g1127) & (!g1128)) + ((!i_8_) & (!g88) & (!g181) & (!g183) & (g1127) & (!g1128)) + ((!i_8_) & (!g88) & (!g181) & (g183) & (!g1127) & (!g1128)) + ((!i_8_) & (!g88) & (!g181) & (g183) & (g1127) & (!g1128)) + ((!i_8_) & (!g88) & (g181) & (!g183) & (!g1127) & (!g1128)) + ((!i_8_) & (!g88) & (g181) & (!g183) & (g1127) & (!g1128)) + ((!i_8_) & (!g88) & (g181) & (g183) & (!g1127) & (!g1128)) + ((!i_8_) & (!g88) & (g181) & (g183) & (g1127) & (!g1128)) + ((!i_8_) & (g88) & (!g181) & (!g183) & (!g1127) & (!g1128)) + ((!i_8_) & (g88) & (!g181) & (!g183) & (g1127) & (!g1128)) + ((!i_8_) & (g88) & (g181) & (!g183) & (!g1127) & (!g1128)) + ((!i_8_) & (g88) & (g181) & (!g183) & (g1127) & (!g1128)) + ((i_8_) & (!g88) & (!g181) & (!g183) & (!g1127) & (!g1128)) + ((i_8_) & (!g88) & (!g181) & (!g183) & (g1127) & (!g1128)) + ((i_8_) & (!g88) & (!g181) & (g183) & (!g1127) & (!g1128)) + ((i_8_) & (!g88) & (!g181) & (g183) & (g1127) & (!g1128)) + ((i_8_) & (!g88) & (g181) & (!g183) & (!g1127) & (!g1128)) + ((i_8_) & (!g88) & (g181) & (!g183) & (g1127) & (!g1128)) + ((i_8_) & (!g88) & (g181) & (g183) & (!g1127) & (!g1128)) + ((i_8_) & (!g88) & (g181) & (g183) & (g1127) & (!g1128)) + ((i_8_) & (g88) & (!g181) & (!g183) & (!g1127) & (!g1128)) + ((i_8_) & (g88) & (!g181) & (g183) & (!g1127) & (!g1128)));
	assign g1130 = (((!i_8_) & (!g88) & (!g339) & (!g117) & (!sk[124]) & (g806)) + ((!i_8_) & (!g88) & (!g339) & (g117) & (!sk[124]) & (g806)) + ((!i_8_) & (!g88) & (g339) & (!g117) & (!sk[124]) & (g806)) + ((!i_8_) & (!g88) & (g339) & (g117) & (!sk[124]) & (g806)) + ((!i_8_) & (g88) & (!g339) & (!g117) & (!sk[124]) & (g806)) + ((!i_8_) & (g88) & (!g339) & (g117) & (!sk[124]) & (g806)) + ((!i_8_) & (g88) & (!g339) & (g117) & (sk[124]) & (!g806)) + ((!i_8_) & (g88) & (!g339) & (g117) & (sk[124]) & (g806)) + ((!i_8_) & (g88) & (g339) & (!g117) & (!sk[124]) & (g806)) + ((!i_8_) & (g88) & (g339) & (!g117) & (sk[124]) & (!g806)) + ((!i_8_) & (g88) & (g339) & (!g117) & (sk[124]) & (g806)) + ((!i_8_) & (g88) & (g339) & (g117) & (!sk[124]) & (g806)) + ((!i_8_) & (g88) & (g339) & (g117) & (sk[124]) & (!g806)) + ((!i_8_) & (g88) & (g339) & (g117) & (sk[124]) & (g806)) + ((i_8_) & (!g88) & (!g339) & (!g117) & (!sk[124]) & (!g806)) + ((i_8_) & (!g88) & (!g339) & (!g117) & (!sk[124]) & (g806)) + ((i_8_) & (!g88) & (!g339) & (g117) & (!sk[124]) & (!g806)) + ((i_8_) & (!g88) & (!g339) & (g117) & (!sk[124]) & (g806)) + ((i_8_) & (!g88) & (g339) & (!g117) & (!sk[124]) & (!g806)) + ((i_8_) & (!g88) & (g339) & (!g117) & (!sk[124]) & (g806)) + ((i_8_) & (!g88) & (g339) & (g117) & (!sk[124]) & (!g806)) + ((i_8_) & (!g88) & (g339) & (g117) & (!sk[124]) & (g806)) + ((i_8_) & (g88) & (!g339) & (!g117) & (!sk[124]) & (!g806)) + ((i_8_) & (g88) & (!g339) & (!g117) & (!sk[124]) & (g806)) + ((i_8_) & (g88) & (!g339) & (!g117) & (sk[124]) & (g806)) + ((i_8_) & (g88) & (!g339) & (g117) & (!sk[124]) & (!g806)) + ((i_8_) & (g88) & (!g339) & (g117) & (!sk[124]) & (g806)) + ((i_8_) & (g88) & (!g339) & (g117) & (sk[124]) & (g806)) + ((i_8_) & (g88) & (g339) & (!g117) & (!sk[124]) & (!g806)) + ((i_8_) & (g88) & (g339) & (!g117) & (!sk[124]) & (g806)) + ((i_8_) & (g88) & (g339) & (!g117) & (sk[124]) & (!g806)) + ((i_8_) & (g88) & (g339) & (!g117) & (sk[124]) & (g806)) + ((i_8_) & (g88) & (g339) & (g117) & (!sk[124]) & (!g806)) + ((i_8_) & (g88) & (g339) & (g117) & (!sk[124]) & (g806)) + ((i_8_) & (g88) & (g339) & (g117) & (sk[124]) & (!g806)) + ((i_8_) & (g88) & (g339) & (g117) & (sk[124]) & (g806)));
	assign g1131 = (((!g19) & (!g16) & (g89) & (!g465) & (!g462) & (!g1130)) + ((!g19) & (!g16) & (g89) & (!g465) & (g462) & (!g1130)) + ((!g19) & (!g16) & (g89) & (g465) & (!g462) & (!g1130)) + ((!g19) & (!g16) & (g89) & (g465) & (g462) & (!g1130)) + ((!g19) & (g16) & (!g89) & (g465) & (g462) & (!g1130)) + ((!g19) & (g16) & (g89) & (!g465) & (!g462) & (!g1130)) + ((!g19) & (g16) & (g89) & (!g465) & (g462) & (!g1130)) + ((!g19) & (g16) & (g89) & (g465) & (!g462) & (!g1130)) + ((!g19) & (g16) & (g89) & (g465) & (g462) & (!g1130)) + ((g19) & (!g16) & (g89) & (!g465) & (!g462) & (!g1130)) + ((g19) & (!g16) & (g89) & (!g465) & (g462) & (!g1130)) + ((g19) & (!g16) & (g89) & (g465) & (!g462) & (!g1130)) + ((g19) & (!g16) & (g89) & (g465) & (g462) & (!g1130)) + ((g19) & (g16) & (g89) & (!g465) & (!g462) & (!g1130)) + ((g19) & (g16) & (g89) & (!g465) & (g462) & (!g1130)) + ((g19) & (g16) & (g89) & (g465) & (!g462) & (!g1130)) + ((g19) & (g16) & (g89) & (g465) & (g462) & (!g1130)));
	assign g1132 = (((!sk[126]) & (!i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g124)) + ((!sk[126]) & (!i_14_) & (!i_12_) & (!i_13_) & (g104) & (g124)) + ((!sk[126]) & (!i_14_) & (!i_12_) & (i_13_) & (!g104) & (g124)) + ((!sk[126]) & (!i_14_) & (!i_12_) & (i_13_) & (g104) & (g124)) + ((!sk[126]) & (!i_14_) & (i_12_) & (!i_13_) & (!g104) & (g124)) + ((!sk[126]) & (!i_14_) & (i_12_) & (!i_13_) & (g104) & (g124)) + ((!sk[126]) & (!i_14_) & (i_12_) & (i_13_) & (!g104) & (g124)) + ((!sk[126]) & (!i_14_) & (i_12_) & (i_13_) & (g104) & (g124)) + ((!sk[126]) & (i_14_) & (!i_12_) & (!i_13_) & (!g104) & (!g124)) + ((!sk[126]) & (i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g124)) + ((!sk[126]) & (i_14_) & (!i_12_) & (!i_13_) & (g104) & (!g124)) + ((!sk[126]) & (i_14_) & (!i_12_) & (!i_13_) & (g104) & (g124)) + ((!sk[126]) & (i_14_) & (!i_12_) & (i_13_) & (!g104) & (!g124)) + ((!sk[126]) & (i_14_) & (!i_12_) & (i_13_) & (!g104) & (g124)) + ((!sk[126]) & (i_14_) & (!i_12_) & (i_13_) & (g104) & (!g124)) + ((!sk[126]) & (i_14_) & (!i_12_) & (i_13_) & (g104) & (g124)) + ((!sk[126]) & (i_14_) & (i_12_) & (!i_13_) & (!g104) & (!g124)) + ((!sk[126]) & (i_14_) & (i_12_) & (!i_13_) & (!g104) & (g124)) + ((!sk[126]) & (i_14_) & (i_12_) & (!i_13_) & (g104) & (!g124)) + ((!sk[126]) & (i_14_) & (i_12_) & (!i_13_) & (g104) & (g124)) + ((!sk[126]) & (i_14_) & (i_12_) & (i_13_) & (!g104) & (!g124)) + ((!sk[126]) & (i_14_) & (i_12_) & (i_13_) & (!g104) & (g124)) + ((!sk[126]) & (i_14_) & (i_12_) & (i_13_) & (g104) & (!g124)) + ((!sk[126]) & (i_14_) & (i_12_) & (i_13_) & (g104) & (g124)) + ((sk[126]) & (!i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g124)) + ((sk[126]) & (!i_14_) & (!i_12_) & (!i_13_) & (g104) & (g124)) + ((sk[126]) & (!i_14_) & (i_12_) & (!i_13_) & (!g104) & (g124)) + ((sk[126]) & (!i_14_) & (i_12_) & (!i_13_) & (g104) & (g124)) + ((sk[126]) & (!i_14_) & (i_12_) & (i_13_) & (!g104) & (g124)) + ((sk[126]) & (!i_14_) & (i_12_) & (i_13_) & (g104) & (!g124)) + ((sk[126]) & (!i_14_) & (i_12_) & (i_13_) & (g104) & (g124)) + ((sk[126]) & (i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g124)) + ((sk[126]) & (i_14_) & (!i_12_) & (!i_13_) & (g104) & (!g124)) + ((sk[126]) & (i_14_) & (!i_12_) & (!i_13_) & (g104) & (g124)) + ((sk[126]) & (i_14_) & (!i_12_) & (i_13_) & (!g104) & (g124)) + ((sk[126]) & (i_14_) & (!i_12_) & (i_13_) & (g104) & (!g124)) + ((sk[126]) & (i_14_) & (!i_12_) & (i_13_) & (g104) & (g124)) + ((sk[126]) & (i_14_) & (i_12_) & (i_13_) & (g104) & (!g124)) + ((sk[126]) & (i_14_) & (i_12_) & (i_13_) & (g104) & (g124)));
	assign g1133 = (((!i_8_) & (!g88) & (!sk[127]) & (!g185) & (!g696) & (g1132)) + ((!i_8_) & (!g88) & (!sk[127]) & (!g185) & (g696) & (g1132)) + ((!i_8_) & (!g88) & (!sk[127]) & (g185) & (!g696) & (g1132)) + ((!i_8_) & (!g88) & (!sk[127]) & (g185) & (g696) & (g1132)) + ((!i_8_) & (g88) & (!sk[127]) & (!g185) & (!g696) & (g1132)) + ((!i_8_) & (g88) & (!sk[127]) & (!g185) & (g696) & (g1132)) + ((!i_8_) & (g88) & (!sk[127]) & (g185) & (!g696) & (g1132)) + ((!i_8_) & (g88) & (!sk[127]) & (g185) & (g696) & (g1132)) + ((!i_8_) & (g88) & (sk[127]) & (!g185) & (!g696) & (!g1132)) + ((!i_8_) & (g88) & (sk[127]) & (!g185) & (!g696) & (g1132)) + ((!i_8_) & (g88) & (sk[127]) & (!g185) & (g696) & (!g1132)) + ((!i_8_) & (g88) & (sk[127]) & (!g185) & (g696) & (g1132)) + ((!i_8_) & (g88) & (sk[127]) & (g185) & (!g696) & (!g1132)) + ((!i_8_) & (g88) & (sk[127]) & (g185) & (!g696) & (g1132)) + ((i_8_) & (!g88) & (!sk[127]) & (!g185) & (!g696) & (!g1132)) + ((i_8_) & (!g88) & (!sk[127]) & (!g185) & (!g696) & (g1132)) + ((i_8_) & (!g88) & (!sk[127]) & (!g185) & (g696) & (!g1132)) + ((i_8_) & (!g88) & (!sk[127]) & (!g185) & (g696) & (g1132)) + ((i_8_) & (!g88) & (!sk[127]) & (g185) & (!g696) & (!g1132)) + ((i_8_) & (!g88) & (!sk[127]) & (g185) & (!g696) & (g1132)) + ((i_8_) & (!g88) & (!sk[127]) & (g185) & (g696) & (!g1132)) + ((i_8_) & (!g88) & (!sk[127]) & (g185) & (g696) & (g1132)) + ((i_8_) & (g88) & (!sk[127]) & (!g185) & (!g696) & (!g1132)) + ((i_8_) & (g88) & (!sk[127]) & (!g185) & (!g696) & (g1132)) + ((i_8_) & (g88) & (!sk[127]) & (!g185) & (g696) & (!g1132)) + ((i_8_) & (g88) & (!sk[127]) & (!g185) & (g696) & (g1132)) + ((i_8_) & (g88) & (!sk[127]) & (g185) & (!g696) & (!g1132)) + ((i_8_) & (g88) & (!sk[127]) & (g185) & (!g696) & (g1132)) + ((i_8_) & (g88) & (!sk[127]) & (g185) & (g696) & (!g1132)) + ((i_8_) & (g88) & (!sk[127]) & (g185) & (g696) & (g1132)) + ((i_8_) & (g88) & (sk[127]) & (!g185) & (!g696) & (g1132)) + ((i_8_) & (g88) & (sk[127]) & (!g185) & (g696) & (g1132)) + ((i_8_) & (g88) & (sk[127]) & (g185) & (!g696) & (g1132)) + ((i_8_) & (g88) & (sk[127]) & (g185) & (g696) & (g1132)));
	assign g1134 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g131) & (g151) & (g158)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g131) & (g151) & (g158)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g131) & (g151) & (g158)) + ((!i_14_) & (i_12_) & (!i_13_) & (g131) & (g151) & (!g158)) + ((!i_14_) & (i_12_) & (!i_13_) & (g131) & (g151) & (g158)) + ((!i_14_) & (i_12_) & (i_13_) & (!g131) & (g151) & (g158)) + ((!i_14_) & (i_12_) & (i_13_) & (g131) & (g151) & (g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (g131) & (g151) & (!g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (g131) & (g151) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (!g131) & (g151) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (g131) & (g151) & (g158)) + ((i_14_) & (i_12_) & (i_13_) & (g131) & (g151) & (!g158)) + ((i_14_) & (i_12_) & (i_13_) & (g131) & (g151) & (g158)));
	assign g1135 = (((!g8) & (!sk[1]) & (!g10) & (!g151) & (!g1133) & (g1134)) + ((!g8) & (!sk[1]) & (!g10) & (!g151) & (g1133) & (g1134)) + ((!g8) & (!sk[1]) & (!g10) & (g151) & (!g1133) & (g1134)) + ((!g8) & (!sk[1]) & (!g10) & (g151) & (g1133) & (g1134)) + ((!g8) & (!sk[1]) & (g10) & (!g151) & (!g1133) & (g1134)) + ((!g8) & (!sk[1]) & (g10) & (!g151) & (g1133) & (g1134)) + ((!g8) & (!sk[1]) & (g10) & (g151) & (!g1133) & (g1134)) + ((!g8) & (!sk[1]) & (g10) & (g151) & (g1133) & (g1134)) + ((!g8) & (sk[1]) & (!g10) & (!g151) & (!g1133) & (!g1134)) + ((!g8) & (sk[1]) & (g10) & (!g151) & (!g1133) & (!g1134)) + ((g8) & (!sk[1]) & (!g10) & (!g151) & (!g1133) & (!g1134)) + ((g8) & (!sk[1]) & (!g10) & (!g151) & (!g1133) & (g1134)) + ((g8) & (!sk[1]) & (!g10) & (!g151) & (g1133) & (!g1134)) + ((g8) & (!sk[1]) & (!g10) & (!g151) & (g1133) & (g1134)) + ((g8) & (!sk[1]) & (!g10) & (g151) & (!g1133) & (!g1134)) + ((g8) & (!sk[1]) & (!g10) & (g151) & (!g1133) & (g1134)) + ((g8) & (!sk[1]) & (!g10) & (g151) & (g1133) & (!g1134)) + ((g8) & (!sk[1]) & (!g10) & (g151) & (g1133) & (g1134)) + ((g8) & (!sk[1]) & (g10) & (!g151) & (!g1133) & (!g1134)) + ((g8) & (!sk[1]) & (g10) & (!g151) & (!g1133) & (g1134)) + ((g8) & (!sk[1]) & (g10) & (!g151) & (g1133) & (!g1134)) + ((g8) & (!sk[1]) & (g10) & (!g151) & (g1133) & (g1134)) + ((g8) & (!sk[1]) & (g10) & (g151) & (!g1133) & (!g1134)) + ((g8) & (!sk[1]) & (g10) & (g151) & (!g1133) & (g1134)) + ((g8) & (!sk[1]) & (g10) & (g151) & (g1133) & (!g1134)) + ((g8) & (!sk[1]) & (g10) & (g151) & (g1133) & (g1134)) + ((g8) & (sk[1]) & (!g10) & (!g151) & (!g1133) & (!g1134)) + ((g8) & (sk[1]) & (!g10) & (g151) & (!g1133) & (!g1134)) + ((g8) & (sk[1]) & (g10) & (!g151) & (!g1133) & (!g1134)));
	assign g1136 = (((!g176) & (!g1126) & (!g1129) & (!g1131) & (!sk[2]) & (g1135)) + ((!g176) & (!g1126) & (!g1129) & (g1131) & (!sk[2]) & (g1135)) + ((!g176) & (!g1126) & (g1129) & (!g1131) & (!sk[2]) & (g1135)) + ((!g176) & (!g1126) & (g1129) & (g1131) & (!sk[2]) & (g1135)) + ((!g176) & (!g1126) & (g1129) & (g1131) & (sk[2]) & (g1135)) + ((!g176) & (g1126) & (!g1129) & (!g1131) & (!sk[2]) & (g1135)) + ((!g176) & (g1126) & (!g1129) & (g1131) & (!sk[2]) & (g1135)) + ((!g176) & (g1126) & (g1129) & (!g1131) & (!sk[2]) & (g1135)) + ((!g176) & (g1126) & (g1129) & (g1131) & (!sk[2]) & (g1135)) + ((g176) & (!g1126) & (!g1129) & (!g1131) & (!sk[2]) & (!g1135)) + ((g176) & (!g1126) & (!g1129) & (!g1131) & (!sk[2]) & (g1135)) + ((g176) & (!g1126) & (!g1129) & (g1131) & (!sk[2]) & (!g1135)) + ((g176) & (!g1126) & (!g1129) & (g1131) & (!sk[2]) & (g1135)) + ((g176) & (!g1126) & (g1129) & (!g1131) & (!sk[2]) & (!g1135)) + ((g176) & (!g1126) & (g1129) & (!g1131) & (!sk[2]) & (g1135)) + ((g176) & (!g1126) & (g1129) & (g1131) & (!sk[2]) & (!g1135)) + ((g176) & (!g1126) & (g1129) & (g1131) & (!sk[2]) & (g1135)) + ((g176) & (g1126) & (!g1129) & (!g1131) & (!sk[2]) & (!g1135)) + ((g176) & (g1126) & (!g1129) & (!g1131) & (!sk[2]) & (g1135)) + ((g176) & (g1126) & (!g1129) & (g1131) & (!sk[2]) & (!g1135)) + ((g176) & (g1126) & (!g1129) & (g1131) & (!sk[2]) & (g1135)) + ((g176) & (g1126) & (g1129) & (!g1131) & (!sk[2]) & (!g1135)) + ((g176) & (g1126) & (g1129) & (!g1131) & (!sk[2]) & (g1135)) + ((g176) & (g1126) & (g1129) & (g1131) & (!sk[2]) & (!g1135)) + ((g176) & (g1126) & (g1129) & (g1131) & (!sk[2]) & (g1135)));
	assign g1137 = (((!g1101) & (!sk[3]) & (!g1105) & (!g1110) & (!g1119) & (g1136)) + ((!g1101) & (!sk[3]) & (!g1105) & (!g1110) & (g1119) & (g1136)) + ((!g1101) & (!sk[3]) & (!g1105) & (g1110) & (!g1119) & (g1136)) + ((!g1101) & (!sk[3]) & (!g1105) & (g1110) & (g1119) & (g1136)) + ((!g1101) & (!sk[3]) & (g1105) & (!g1110) & (!g1119) & (g1136)) + ((!g1101) & (!sk[3]) & (g1105) & (!g1110) & (g1119) & (g1136)) + ((!g1101) & (!sk[3]) & (g1105) & (g1110) & (!g1119) & (g1136)) + ((!g1101) & (!sk[3]) & (g1105) & (g1110) & (g1119) & (g1136)) + ((g1101) & (!sk[3]) & (!g1105) & (!g1110) & (!g1119) & (!g1136)) + ((g1101) & (!sk[3]) & (!g1105) & (!g1110) & (!g1119) & (g1136)) + ((g1101) & (!sk[3]) & (!g1105) & (!g1110) & (g1119) & (!g1136)) + ((g1101) & (!sk[3]) & (!g1105) & (!g1110) & (g1119) & (g1136)) + ((g1101) & (!sk[3]) & (!g1105) & (g1110) & (!g1119) & (!g1136)) + ((g1101) & (!sk[3]) & (!g1105) & (g1110) & (!g1119) & (g1136)) + ((g1101) & (!sk[3]) & (!g1105) & (g1110) & (g1119) & (!g1136)) + ((g1101) & (!sk[3]) & (!g1105) & (g1110) & (g1119) & (g1136)) + ((g1101) & (!sk[3]) & (g1105) & (!g1110) & (!g1119) & (!g1136)) + ((g1101) & (!sk[3]) & (g1105) & (!g1110) & (!g1119) & (g1136)) + ((g1101) & (!sk[3]) & (g1105) & (!g1110) & (g1119) & (!g1136)) + ((g1101) & (!sk[3]) & (g1105) & (!g1110) & (g1119) & (g1136)) + ((g1101) & (!sk[3]) & (g1105) & (g1110) & (!g1119) & (!g1136)) + ((g1101) & (!sk[3]) & (g1105) & (g1110) & (!g1119) & (g1136)) + ((g1101) & (!sk[3]) & (g1105) & (g1110) & (g1119) & (!g1136)) + ((g1101) & (!sk[3]) & (g1105) & (g1110) & (g1119) & (g1136)) + ((g1101) & (sk[3]) & (g1105) & (g1110) & (g1119) & (g1136)));
	assign g1138 = (((!i_1_) & (sk[4]) & (!i_0_) & (!i_2_)) + ((!i_1_) & (sk[4]) & (i_0_) & (i_2_)) + ((i_1_) & (!sk[4]) & (!i_0_) & (!i_2_)) + ((i_1_) & (!sk[4]) & (!i_0_) & (i_2_)) + ((i_1_) & (!sk[4]) & (i_0_) & (!i_2_)) + ((i_1_) & (!sk[4]) & (i_0_) & (i_2_)) + ((i_1_) & (sk[4]) & (!i_0_) & (!i_2_)) + ((i_1_) & (sk[4]) & (i_0_) & (!i_2_)) + ((i_1_) & (sk[4]) & (i_0_) & (i_2_)));
	assign g1139 = (((!sk[5]) & (g20) & (!g460) & (!g710)) + ((!sk[5]) & (g20) & (!g460) & (g710)) + ((!sk[5]) & (g20) & (g460) & (!g710)) + ((!sk[5]) & (g20) & (g460) & (g710)) + ((sk[5]) & (g20) & (!g460) & (!g710)));
	assign g1140 = (((g528) & (!sk[6]) & (!g1031)) + ((g528) & (!sk[6]) & (g1031)) + ((g528) & (sk[6]) & (g1031)));
	assign g1141 = (((!i_8_) & (!sk[7]) & (!g23) & (g108) & (g506)) + ((!i_8_) & (!sk[7]) & (g23) & (!g108) & (!g506)) + ((!i_8_) & (!sk[7]) & (g23) & (!g108) & (g506)) + ((!i_8_) & (!sk[7]) & (g23) & (g108) & (!g506)) + ((!i_8_) & (!sk[7]) & (g23) & (g108) & (g506)) + ((i_8_) & (!sk[7]) & (!g23) & (g108) & (!g506)) + ((i_8_) & (!sk[7]) & (!g23) & (g108) & (g506)) + ((i_8_) & (!sk[7]) & (g23) & (!g108) & (!g506)) + ((i_8_) & (!sk[7]) & (g23) & (!g108) & (g506)) + ((i_8_) & (!sk[7]) & (g23) & (g108) & (!g506)) + ((i_8_) & (!sk[7]) & (g23) & (g108) & (g506)) + ((i_8_) & (sk[7]) & (!g23) & (g108) & (g506)) + ((i_8_) & (sk[7]) & (g23) & (g108) & (!g506)) + ((i_8_) & (sk[7]) & (g23) & (g108) & (g506)));
	assign g1142 = (((!sk[8]) & (!i_8_) & (!g21) & (g108) & (g561)) + ((!sk[8]) & (!i_8_) & (g21) & (!g108) & (!g561)) + ((!sk[8]) & (!i_8_) & (g21) & (!g108) & (g561)) + ((!sk[8]) & (!i_8_) & (g21) & (g108) & (!g561)) + ((!sk[8]) & (!i_8_) & (g21) & (g108) & (g561)) + ((!sk[8]) & (i_8_) & (!g21) & (g108) & (!g561)) + ((!sk[8]) & (i_8_) & (!g21) & (g108) & (g561)) + ((!sk[8]) & (i_8_) & (g21) & (!g108) & (!g561)) + ((!sk[8]) & (i_8_) & (g21) & (!g108) & (g561)) + ((!sk[8]) & (i_8_) & (g21) & (g108) & (!g561)) + ((!sk[8]) & (i_8_) & (g21) & (g108) & (g561)) + ((sk[8]) & (i_8_) & (!g21) & (g108) & (g561)) + ((sk[8]) & (i_8_) & (g21) & (g108) & (!g561)) + ((sk[8]) & (i_8_) & (g21) & (g108) & (g561)));
	assign g1143 = (((!g145) & (!g127) & (!g114) & (!g596) & (!g1141) & (!g1142)) + ((!g145) & (!g127) & (g114) & (!g596) & (!g1141) & (!g1142)) + ((!g145) & (g127) & (!g114) & (!g596) & (!g1141) & (!g1142)) + ((!g145) & (g127) & (g114) & (!g596) & (!g1141) & (!g1142)) + ((g145) & (g127) & (!g114) & (!g596) & (!g1141) & (!g1142)));
	assign g1144 = (((!g112) & (!g136) & (!g474) & (!g1139) & (!g1140) & (g1143)) + ((!g112) & (!g136) & (!g474) & (!g1139) & (g1140) & (g1143)) + ((!g112) & (!g136) & (!g474) & (g1139) & (!g1140) & (g1143)) + ((!g112) & (!g136) & (!g474) & (g1139) & (g1140) & (g1143)) + ((!g112) & (!g136) & (g474) & (!g1139) & (!g1140) & (g1143)) + ((!g112) & (!g136) & (g474) & (!g1139) & (g1140) & (g1143)) + ((!g112) & (!g136) & (g474) & (g1139) & (!g1140) & (g1143)) + ((!g112) & (!g136) & (g474) & (g1139) & (g1140) & (g1143)) + ((!g112) & (g136) & (!g474) & (g1139) & (g1140) & (g1143)) + ((!g112) & (g136) & (g474) & (g1139) & (g1140) & (g1143)) + ((g112) & (!g136) & (!g474) & (!g1139) & (g1140) & (g1143)) + ((g112) & (!g136) & (!g474) & (g1139) & (g1140) & (g1143)) + ((g112) & (g136) & (!g474) & (g1139) & (g1140) & (g1143)));
	assign g1145 = (((g880) & (g694) & (g860) & (g890) & (g917) & (g1144)));
	assign g1146 = (((!i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (!g7) & (g9)) + ((!i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (g7) & (g9)) + ((!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!g7) & (g9)) + ((!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (g7) & (g9)) + ((!i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (g7) & (!g9)) + ((!i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (g7) & (g9)) + ((!i_11_) & (i_9_) & (i_10_) & (!i_15_) & (g7) & (!g9)) + ((!i_11_) & (i_9_) & (i_10_) & (!i_15_) & (g7) & (g9)) + ((!i_11_) & (i_9_) & (i_10_) & (i_15_) & (!g7) & (g9)) + ((!i_11_) & (i_9_) & (i_10_) & (i_15_) & (g7) & (g9)));
	assign g1147 = (((!g151) & (!g544) & (!sk[13]) & (g487) & (g1146)) + ((!g151) & (g544) & (!sk[13]) & (!g487) & (!g1146)) + ((!g151) & (g544) & (!sk[13]) & (!g487) & (g1146)) + ((!g151) & (g544) & (!sk[13]) & (g487) & (!g1146)) + ((!g151) & (g544) & (!sk[13]) & (g487) & (g1146)) + ((g151) & (!g544) & (!sk[13]) & (g487) & (!g1146)) + ((g151) & (!g544) & (!sk[13]) & (g487) & (g1146)) + ((g151) & (!g544) & (sk[13]) & (!g487) & (!g1146)) + ((g151) & (!g544) & (sk[13]) & (!g487) & (g1146)) + ((g151) & (!g544) & (sk[13]) & (g487) & (!g1146)) + ((g151) & (!g544) & (sk[13]) & (g487) & (g1146)) + ((g151) & (g544) & (!sk[13]) & (!g487) & (!g1146)) + ((g151) & (g544) & (!sk[13]) & (!g487) & (g1146)) + ((g151) & (g544) & (!sk[13]) & (g487) & (!g1146)) + ((g151) & (g544) & (!sk[13]) & (g487) & (g1146)) + ((g151) & (g544) & (sk[13]) & (!g487) & (g1146)) + ((g151) & (g544) & (sk[13]) & (g487) & (!g1146)) + ((g151) & (g544) & (sk[13]) & (g487) & (g1146)));
	assign g1148 = (((!sk[14]) & (g112) & (!g114) & (!g464)) + ((!sk[14]) & (g112) & (!g114) & (g464)) + ((!sk[14]) & (g112) & (g114) & (!g464)) + ((!sk[14]) & (g112) & (g114) & (g464)) + ((sk[14]) & (g112) & (!g114) & (!g464)) + ((sk[14]) & (g112) & (g114) & (!g464)) + ((sk[14]) & (g112) & (g114) & (g464)));
	assign g1149 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g11) & (g22) & (g112)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g11) & (g22) & (g112)) + ((!i_14_) & (!i_12_) & (i_13_) & (g11) & (!g22) & (g112)) + ((!i_14_) & (!i_12_) & (i_13_) & (g11) & (g22) & (g112)) + ((!i_14_) & (i_12_) & (!i_13_) & (g11) & (!g22) & (g112)) + ((!i_14_) & (i_12_) & (!i_13_) & (g11) & (g22) & (g112)) + ((i_14_) & (i_12_) & (!i_13_) & (!g11) & (g22) & (g112)) + ((i_14_) & (i_12_) & (!i_13_) & (g11) & (g22) & (g112)) + ((i_14_) & (i_12_) & (i_13_) & (g11) & (!g22) & (g112)) + ((i_14_) & (i_12_) & (i_13_) & (g11) & (g22) & (g112)));
	assign g1150 = (((!g112) & (!g183) & (!sk[16]) & (!g123) & (!g670) & (g887)) + ((!g112) & (!g183) & (!sk[16]) & (!g123) & (g670) & (g887)) + ((!g112) & (!g183) & (!sk[16]) & (g123) & (!g670) & (g887)) + ((!g112) & (!g183) & (!sk[16]) & (g123) & (g670) & (g887)) + ((!g112) & (g183) & (!sk[16]) & (!g123) & (!g670) & (g887)) + ((!g112) & (g183) & (!sk[16]) & (!g123) & (g670) & (g887)) + ((!g112) & (g183) & (!sk[16]) & (g123) & (!g670) & (g887)) + ((!g112) & (g183) & (!sk[16]) & (g123) & (g670) & (g887)) + ((g112) & (!g183) & (!sk[16]) & (!g123) & (!g670) & (!g887)) + ((g112) & (!g183) & (!sk[16]) & (!g123) & (!g670) & (g887)) + ((g112) & (!g183) & (!sk[16]) & (!g123) & (g670) & (!g887)) + ((g112) & (!g183) & (!sk[16]) & (!g123) & (g670) & (g887)) + ((g112) & (!g183) & (!sk[16]) & (g123) & (!g670) & (!g887)) + ((g112) & (!g183) & (!sk[16]) & (g123) & (!g670) & (g887)) + ((g112) & (!g183) & (!sk[16]) & (g123) & (g670) & (!g887)) + ((g112) & (!g183) & (!sk[16]) & (g123) & (g670) & (g887)) + ((g112) & (!g183) & (sk[16]) & (!g123) & (!g670) & (!g887)) + ((g112) & (!g183) & (sk[16]) & (!g123) & (g670) & (!g887)) + ((g112) & (!g183) & (sk[16]) & (!g123) & (g670) & (g887)) + ((g112) & (!g183) & (sk[16]) & (g123) & (!g670) & (!g887)) + ((g112) & (!g183) & (sk[16]) & (g123) & (!g670) & (g887)) + ((g112) & (!g183) & (sk[16]) & (g123) & (g670) & (!g887)) + ((g112) & (!g183) & (sk[16]) & (g123) & (g670) & (g887)) + ((g112) & (g183) & (!sk[16]) & (!g123) & (!g670) & (!g887)) + ((g112) & (g183) & (!sk[16]) & (!g123) & (!g670) & (g887)) + ((g112) & (g183) & (!sk[16]) & (!g123) & (g670) & (!g887)) + ((g112) & (g183) & (!sk[16]) & (!g123) & (g670) & (g887)) + ((g112) & (g183) & (!sk[16]) & (g123) & (!g670) & (!g887)) + ((g112) & (g183) & (!sk[16]) & (g123) & (!g670) & (g887)) + ((g112) & (g183) & (!sk[16]) & (g123) & (g670) & (!g887)) + ((g112) & (g183) & (!sk[16]) & (g123) & (g670) & (g887)) + ((g112) & (g183) & (sk[16]) & (!g123) & (!g670) & (!g887)) + ((g112) & (g183) & (sk[16]) & (!g123) & (!g670) & (g887)) + ((g112) & (g183) & (sk[16]) & (!g123) & (g670) & (!g887)) + ((g112) & (g183) & (sk[16]) & (!g123) & (g670) & (g887)) + ((g112) & (g183) & (sk[16]) & (g123) & (!g670) & (!g887)) + ((g112) & (g183) & (sk[16]) & (g123) & (!g670) & (g887)) + ((g112) & (g183) & (sk[16]) & (g123) & (g670) & (!g887)) + ((g112) & (g183) & (sk[16]) & (g123) & (g670) & (g887)));
	assign g1151 = (((!g562) & (!g804) & (!g1148) & (!sk[17]) & (!g1149) & (g1150)) + ((!g562) & (!g804) & (!g1148) & (!sk[17]) & (g1149) & (g1150)) + ((!g562) & (!g804) & (!g1148) & (sk[17]) & (!g1149) & (!g1150)) + ((!g562) & (!g804) & (g1148) & (!sk[17]) & (!g1149) & (g1150)) + ((!g562) & (!g804) & (g1148) & (!sk[17]) & (g1149) & (g1150)) + ((!g562) & (g804) & (!g1148) & (!sk[17]) & (!g1149) & (g1150)) + ((!g562) & (g804) & (!g1148) & (!sk[17]) & (g1149) & (g1150)) + ((!g562) & (g804) & (g1148) & (!sk[17]) & (!g1149) & (g1150)) + ((!g562) & (g804) & (g1148) & (!sk[17]) & (g1149) & (g1150)) + ((g562) & (!g804) & (!g1148) & (!sk[17]) & (!g1149) & (!g1150)) + ((g562) & (!g804) & (!g1148) & (!sk[17]) & (!g1149) & (g1150)) + ((g562) & (!g804) & (!g1148) & (!sk[17]) & (g1149) & (!g1150)) + ((g562) & (!g804) & (!g1148) & (!sk[17]) & (g1149) & (g1150)) + ((g562) & (!g804) & (g1148) & (!sk[17]) & (!g1149) & (!g1150)) + ((g562) & (!g804) & (g1148) & (!sk[17]) & (!g1149) & (g1150)) + ((g562) & (!g804) & (g1148) & (!sk[17]) & (g1149) & (!g1150)) + ((g562) & (!g804) & (g1148) & (!sk[17]) & (g1149) & (g1150)) + ((g562) & (g804) & (!g1148) & (!sk[17]) & (!g1149) & (!g1150)) + ((g562) & (g804) & (!g1148) & (!sk[17]) & (!g1149) & (g1150)) + ((g562) & (g804) & (!g1148) & (!sk[17]) & (g1149) & (!g1150)) + ((g562) & (g804) & (!g1148) & (!sk[17]) & (g1149) & (g1150)) + ((g562) & (g804) & (g1148) & (!sk[17]) & (!g1149) & (!g1150)) + ((g562) & (g804) & (g1148) & (!sk[17]) & (!g1149) & (g1150)) + ((g562) & (g804) & (g1148) & (!sk[17]) & (g1149) & (!g1150)) + ((g562) & (g804) & (g1148) & (!sk[17]) & (g1149) & (g1150)));
	assign g1152 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g136) & (g124)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g104) & (g136) & (g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g104) & (g136) & (g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (g104) & (g136) & (!g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (g104) & (g136) & (g124)) + ((!i_14_) & (i_12_) & (i_13_) & (!g104) & (g136) & (g124)) + ((!i_14_) & (i_12_) & (i_13_) & (g104) & (g136) & (!g124)) + ((!i_14_) & (i_12_) & (i_13_) & (g104) & (g136) & (g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g136) & (g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (g104) & (g136) & (!g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (g104) & (g136) & (g124)) + ((i_14_) & (!i_12_) & (i_13_) & (g104) & (g136) & (!g124)) + ((i_14_) & (!i_12_) & (i_13_) & (g104) & (g136) & (g124)) + ((i_14_) & (i_12_) & (i_13_) & (g104) & (g136) & (!g124)) + ((i_14_) & (i_12_) & (i_13_) & (g104) & (g136) & (g124)));
	assign g1153 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g112) & (g124)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g104) & (g112) & (g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g104) & (g112) & (g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (g104) & (g112) & (!g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (g104) & (g112) & (g124)) + ((!i_14_) & (i_12_) & (i_13_) & (!g104) & (g112) & (g124)) + ((!i_14_) & (i_12_) & (i_13_) & (g104) & (g112) & (!g124)) + ((!i_14_) & (i_12_) & (i_13_) & (g104) & (g112) & (g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g112) & (g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (g104) & (g112) & (!g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (g104) & (g112) & (g124)) + ((i_14_) & (!i_12_) & (i_13_) & (g104) & (g112) & (!g124)) + ((i_14_) & (!i_12_) & (i_13_) & (g104) & (g112) & (g124)) + ((i_14_) & (i_12_) & (i_13_) & (g104) & (g112) & (!g124)) + ((i_14_) & (i_12_) & (i_13_) & (g104) & (g112) & (g124)));
	assign g1154 = (((!sk[20]) & (!g101) & (!g323) & (!g231) & (!g478) & (g1001)) + ((!sk[20]) & (!g101) & (!g323) & (!g231) & (g478) & (g1001)) + ((!sk[20]) & (!g101) & (!g323) & (g231) & (!g478) & (g1001)) + ((!sk[20]) & (!g101) & (!g323) & (g231) & (g478) & (g1001)) + ((!sk[20]) & (!g101) & (g323) & (!g231) & (!g478) & (g1001)) + ((!sk[20]) & (!g101) & (g323) & (!g231) & (g478) & (g1001)) + ((!sk[20]) & (!g101) & (g323) & (g231) & (!g478) & (g1001)) + ((!sk[20]) & (!g101) & (g323) & (g231) & (g478) & (g1001)) + ((!sk[20]) & (g101) & (!g323) & (!g231) & (!g478) & (!g1001)) + ((!sk[20]) & (g101) & (!g323) & (!g231) & (!g478) & (g1001)) + ((!sk[20]) & (g101) & (!g323) & (!g231) & (g478) & (!g1001)) + ((!sk[20]) & (g101) & (!g323) & (!g231) & (g478) & (g1001)) + ((!sk[20]) & (g101) & (!g323) & (g231) & (!g478) & (!g1001)) + ((!sk[20]) & (g101) & (!g323) & (g231) & (!g478) & (g1001)) + ((!sk[20]) & (g101) & (!g323) & (g231) & (g478) & (!g1001)) + ((!sk[20]) & (g101) & (!g323) & (g231) & (g478) & (g1001)) + ((!sk[20]) & (g101) & (g323) & (!g231) & (!g478) & (!g1001)) + ((!sk[20]) & (g101) & (g323) & (!g231) & (!g478) & (g1001)) + ((!sk[20]) & (g101) & (g323) & (!g231) & (g478) & (!g1001)) + ((!sk[20]) & (g101) & (g323) & (!g231) & (g478) & (g1001)) + ((!sk[20]) & (g101) & (g323) & (g231) & (!g478) & (!g1001)) + ((!sk[20]) & (g101) & (g323) & (g231) & (!g478) & (g1001)) + ((!sk[20]) & (g101) & (g323) & (g231) & (g478) & (!g1001)) + ((!sk[20]) & (g101) & (g323) & (g231) & (g478) & (g1001)) + ((sk[20]) & (!g101) & (!g323) & (!g231) & (!g478) & (!g1001)) + ((sk[20]) & (!g101) & (!g323) & (!g231) & (!g478) & (g1001)) + ((sk[20]) & (!g101) & (!g323) & (!g231) & (g478) & (!g1001)) + ((sk[20]) & (!g101) & (!g323) & (!g231) & (g478) & (g1001)) + ((sk[20]) & (!g101) & (!g323) & (g231) & (!g478) & (!g1001)) + ((sk[20]) & (!g101) & (!g323) & (g231) & (!g478) & (g1001)) + ((sk[20]) & (!g101) & (!g323) & (g231) & (g478) & (!g1001)) + ((sk[20]) & (!g101) & (!g323) & (g231) & (g478) & (g1001)) + ((sk[20]) & (!g101) & (g323) & (g231) & (!g478) & (!g1001)) + ((sk[20]) & (!g101) & (g323) & (g231) & (!g478) & (g1001)) + ((sk[20]) & (g101) & (!g323) & (!g231) & (!g478) & (g1001)) + ((sk[20]) & (g101) & (!g323) & (!g231) & (g478) & (g1001)) + ((sk[20]) & (g101) & (!g323) & (g231) & (!g478) & (g1001)) + ((sk[20]) & (g101) & (!g323) & (g231) & (g478) & (g1001)) + ((sk[20]) & (g101) & (g323) & (g231) & (!g478) & (g1001)));
	assign g1155 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g145) & (g124)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g104) & (g145) & (g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g104) & (g145) & (g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (g104) & (g145) & (g124)) + ((!i_14_) & (i_12_) & (i_13_) & (!g104) & (g145) & (g124)) + ((!i_14_) & (i_12_) & (i_13_) & (g104) & (g145) & (!g124)) + ((!i_14_) & (i_12_) & (i_13_) & (g104) & (g145) & (g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g145) & (g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (g104) & (g145) & (!g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (g104) & (g145) & (g124)) + ((i_14_) & (!i_12_) & (i_13_) & (!g104) & (g145) & (g124)) + ((i_14_) & (!i_12_) & (i_13_) & (g104) & (g145) & (!g124)) + ((i_14_) & (!i_12_) & (i_13_) & (g104) & (g145) & (g124)) + ((i_14_) & (i_12_) & (i_13_) & (g104) & (g145) & (!g124)) + ((i_14_) & (i_12_) & (i_13_) & (g104) & (g145) & (g124)));
	assign g1156 = (((!g1151) & (!g1152) & (!g1153) & (!sk[22]) & (!g1154) & (g1155)) + ((!g1151) & (!g1152) & (!g1153) & (!sk[22]) & (g1154) & (g1155)) + ((!g1151) & (!g1152) & (g1153) & (!sk[22]) & (!g1154) & (g1155)) + ((!g1151) & (!g1152) & (g1153) & (!sk[22]) & (g1154) & (g1155)) + ((!g1151) & (g1152) & (!g1153) & (!sk[22]) & (!g1154) & (g1155)) + ((!g1151) & (g1152) & (!g1153) & (!sk[22]) & (g1154) & (g1155)) + ((!g1151) & (g1152) & (g1153) & (!sk[22]) & (!g1154) & (g1155)) + ((!g1151) & (g1152) & (g1153) & (!sk[22]) & (g1154) & (g1155)) + ((g1151) & (!g1152) & (!g1153) & (!sk[22]) & (!g1154) & (!g1155)) + ((g1151) & (!g1152) & (!g1153) & (!sk[22]) & (!g1154) & (g1155)) + ((g1151) & (!g1152) & (!g1153) & (!sk[22]) & (g1154) & (!g1155)) + ((g1151) & (!g1152) & (!g1153) & (!sk[22]) & (g1154) & (g1155)) + ((g1151) & (!g1152) & (!g1153) & (sk[22]) & (g1154) & (!g1155)) + ((g1151) & (!g1152) & (g1153) & (!sk[22]) & (!g1154) & (!g1155)) + ((g1151) & (!g1152) & (g1153) & (!sk[22]) & (!g1154) & (g1155)) + ((g1151) & (!g1152) & (g1153) & (!sk[22]) & (g1154) & (!g1155)) + ((g1151) & (!g1152) & (g1153) & (!sk[22]) & (g1154) & (g1155)) + ((g1151) & (g1152) & (!g1153) & (!sk[22]) & (!g1154) & (!g1155)) + ((g1151) & (g1152) & (!g1153) & (!sk[22]) & (!g1154) & (g1155)) + ((g1151) & (g1152) & (!g1153) & (!sk[22]) & (g1154) & (!g1155)) + ((g1151) & (g1152) & (!g1153) & (!sk[22]) & (g1154) & (g1155)) + ((g1151) & (g1152) & (g1153) & (!sk[22]) & (!g1154) & (!g1155)) + ((g1151) & (g1152) & (g1153) & (!sk[22]) & (!g1154) & (g1155)) + ((g1151) & (g1152) & (g1153) & (!sk[22]) & (g1154) & (!g1155)) + ((g1151) & (g1152) & (g1153) & (!sk[22]) & (g1154) & (g1155)));
	assign g1157 = (((!i_8_) & (!g108) & (!sk[23]) & (!g183) & (!g540) & (g704)) + ((!i_8_) & (!g108) & (!sk[23]) & (!g183) & (g540) & (g704)) + ((!i_8_) & (!g108) & (!sk[23]) & (g183) & (!g540) & (g704)) + ((!i_8_) & (!g108) & (!sk[23]) & (g183) & (g540) & (g704)) + ((!i_8_) & (!g108) & (sk[23]) & (!g183) & (!g540) & (!g704)) + ((!i_8_) & (!g108) & (sk[23]) & (g183) & (!g540) & (!g704)) + ((!i_8_) & (g108) & (!sk[23]) & (!g183) & (!g540) & (g704)) + ((!i_8_) & (g108) & (!sk[23]) & (!g183) & (g540) & (g704)) + ((!i_8_) & (g108) & (!sk[23]) & (g183) & (!g540) & (g704)) + ((!i_8_) & (g108) & (!sk[23]) & (g183) & (g540) & (g704)) + ((!i_8_) & (g108) & (sk[23]) & (!g183) & (!g540) & (!g704)) + ((!i_8_) & (g108) & (sk[23]) & (g183) & (!g540) & (!g704)) + ((i_8_) & (!g108) & (!sk[23]) & (!g183) & (!g540) & (!g704)) + ((i_8_) & (!g108) & (!sk[23]) & (!g183) & (!g540) & (g704)) + ((i_8_) & (!g108) & (!sk[23]) & (!g183) & (g540) & (!g704)) + ((i_8_) & (!g108) & (!sk[23]) & (!g183) & (g540) & (g704)) + ((i_8_) & (!g108) & (!sk[23]) & (g183) & (!g540) & (!g704)) + ((i_8_) & (!g108) & (!sk[23]) & (g183) & (!g540) & (g704)) + ((i_8_) & (!g108) & (!sk[23]) & (g183) & (g540) & (!g704)) + ((i_8_) & (!g108) & (!sk[23]) & (g183) & (g540) & (g704)) + ((i_8_) & (!g108) & (sk[23]) & (!g183) & (!g540) & (!g704)) + ((i_8_) & (!g108) & (sk[23]) & (g183) & (!g540) & (!g704)) + ((i_8_) & (g108) & (!sk[23]) & (!g183) & (!g540) & (!g704)) + ((i_8_) & (g108) & (!sk[23]) & (!g183) & (!g540) & (g704)) + ((i_8_) & (g108) & (!sk[23]) & (!g183) & (g540) & (!g704)) + ((i_8_) & (g108) & (!sk[23]) & (!g183) & (g540) & (g704)) + ((i_8_) & (g108) & (!sk[23]) & (g183) & (!g540) & (!g704)) + ((i_8_) & (g108) & (!sk[23]) & (g183) & (!g540) & (g704)) + ((i_8_) & (g108) & (!sk[23]) & (g183) & (g540) & (!g704)) + ((i_8_) & (g108) & (!sk[23]) & (g183) & (g540) & (g704)) + ((i_8_) & (g108) & (sk[23]) & (!g183) & (!g540) & (!g704)));
	assign g1158 = (((!sk[24]) & (g145) & (!g1157)) + ((!sk[24]) & (g145) & (g1157)) + ((sk[24]) & (g145) & (!g1157)));
	assign g1159 = (((!g268) & (!g556) & (!sk[25]) & (!g669) & (!g672) & (g979)) + ((!g268) & (!g556) & (!sk[25]) & (!g669) & (g672) & (g979)) + ((!g268) & (!g556) & (!sk[25]) & (g669) & (!g672) & (g979)) + ((!g268) & (!g556) & (!sk[25]) & (g669) & (g672) & (g979)) + ((!g268) & (g556) & (!sk[25]) & (!g669) & (!g672) & (g979)) + ((!g268) & (g556) & (!sk[25]) & (!g669) & (g672) & (g979)) + ((!g268) & (g556) & (!sk[25]) & (g669) & (!g672) & (g979)) + ((!g268) & (g556) & (!sk[25]) & (g669) & (g672) & (g979)) + ((!g268) & (g556) & (sk[25]) & (g669) & (!g672) & (g979)) + ((g268) & (!g556) & (!sk[25]) & (!g669) & (!g672) & (!g979)) + ((g268) & (!g556) & (!sk[25]) & (!g669) & (!g672) & (g979)) + ((g268) & (!g556) & (!sk[25]) & (!g669) & (g672) & (!g979)) + ((g268) & (!g556) & (!sk[25]) & (!g669) & (g672) & (g979)) + ((g268) & (!g556) & (!sk[25]) & (g669) & (!g672) & (!g979)) + ((g268) & (!g556) & (!sk[25]) & (g669) & (!g672) & (g979)) + ((g268) & (!g556) & (!sk[25]) & (g669) & (g672) & (!g979)) + ((g268) & (!g556) & (!sk[25]) & (g669) & (g672) & (g979)) + ((g268) & (g556) & (!sk[25]) & (!g669) & (!g672) & (!g979)) + ((g268) & (g556) & (!sk[25]) & (!g669) & (!g672) & (g979)) + ((g268) & (g556) & (!sk[25]) & (!g669) & (g672) & (!g979)) + ((g268) & (g556) & (!sk[25]) & (!g669) & (g672) & (g979)) + ((g268) & (g556) & (!sk[25]) & (g669) & (!g672) & (!g979)) + ((g268) & (g556) & (!sk[25]) & (g669) & (!g672) & (g979)) + ((g268) & (g556) & (!sk[25]) & (g669) & (g672) & (!g979)) + ((g268) & (g556) & (!sk[25]) & (g669) & (g672) & (g979)));
	assign g1160 = (((!g16) & (g323) & (!g534) & (!g980) & (!g1062) & (!g1159)) + ((!g16) & (g323) & (!g534) & (!g980) & (!g1062) & (g1159)) + ((!g16) & (g323) & (!g534) & (!g980) & (g1062) & (!g1159)) + ((!g16) & (g323) & (!g534) & (!g980) & (g1062) & (g1159)) + ((!g16) & (g323) & (!g534) & (g980) & (!g1062) & (!g1159)) + ((!g16) & (g323) & (!g534) & (g980) & (!g1062) & (g1159)) + ((!g16) & (g323) & (!g534) & (g980) & (g1062) & (!g1159)) + ((!g16) & (g323) & (!g534) & (g980) & (g1062) & (g1159)) + ((!g16) & (g323) & (g534) & (!g980) & (!g1062) & (!g1159)) + ((!g16) & (g323) & (g534) & (!g980) & (!g1062) & (g1159)) + ((!g16) & (g323) & (g534) & (!g980) & (g1062) & (!g1159)) + ((!g16) & (g323) & (g534) & (!g980) & (g1062) & (g1159)) + ((!g16) & (g323) & (g534) & (g980) & (!g1062) & (!g1159)) + ((!g16) & (g323) & (g534) & (g980) & (!g1062) & (g1159)) + ((!g16) & (g323) & (g534) & (g980) & (g1062) & (!g1159)) + ((!g16) & (g323) & (g534) & (g980) & (g1062) & (g1159)) + ((g16) & (g323) & (!g534) & (!g980) & (!g1062) & (!g1159)) + ((g16) & (g323) & (!g534) & (!g980) & (!g1062) & (g1159)) + ((g16) & (g323) & (!g534) & (!g980) & (g1062) & (!g1159)) + ((g16) & (g323) & (!g534) & (!g980) & (g1062) & (g1159)) + ((g16) & (g323) & (!g534) & (g980) & (!g1062) & (!g1159)) + ((g16) & (g323) & (!g534) & (g980) & (!g1062) & (g1159)) + ((g16) & (g323) & (!g534) & (g980) & (g1062) & (!g1159)) + ((g16) & (g323) & (g534) & (!g980) & (!g1062) & (!g1159)) + ((g16) & (g323) & (g534) & (!g980) & (!g1062) & (g1159)) + ((g16) & (g323) & (g534) & (!g980) & (g1062) & (!g1159)) + ((g16) & (g323) & (g534) & (!g980) & (g1062) & (g1159)) + ((g16) & (g323) & (g534) & (g980) & (!g1062) & (!g1159)) + ((g16) & (g323) & (g534) & (g980) & (!g1062) & (g1159)) + ((g16) & (g323) & (g534) & (g980) & (g1062) & (!g1159)) + ((g16) & (g323) & (g534) & (g980) & (g1062) & (g1159)));
	assign g1161 = (((!sk[27]) & (!i_14_) & (!i_12_) & (g119) & (g485)) + ((!sk[27]) & (!i_14_) & (i_12_) & (!g119) & (!g485)) + ((!sk[27]) & (!i_14_) & (i_12_) & (!g119) & (g485)) + ((!sk[27]) & (!i_14_) & (i_12_) & (g119) & (!g485)) + ((!sk[27]) & (!i_14_) & (i_12_) & (g119) & (g485)) + ((!sk[27]) & (i_14_) & (!i_12_) & (g119) & (!g485)) + ((!sk[27]) & (i_14_) & (!i_12_) & (g119) & (g485)) + ((!sk[27]) & (i_14_) & (i_12_) & (!g119) & (!g485)) + ((!sk[27]) & (i_14_) & (i_12_) & (!g119) & (g485)) + ((!sk[27]) & (i_14_) & (i_12_) & (g119) & (!g485)) + ((!sk[27]) & (i_14_) & (i_12_) & (g119) & (g485)) + ((sk[27]) & (!i_14_) & (!i_12_) & (!g119) & (!g485)) + ((sk[27]) & (!i_14_) & (!i_12_) & (g119) & (!g485)) + ((sk[27]) & (!i_14_) & (i_12_) & (!g119) & (!g485)) + ((sk[27]) & (!i_14_) & (i_12_) & (g119) & (!g485)) + ((sk[27]) & (i_14_) & (!i_12_) & (!g119) & (!g485)) + ((sk[27]) & (i_14_) & (i_12_) & (!g119) & (!g485)) + ((sk[27]) & (i_14_) & (i_12_) & (g119) & (!g485)));
	assign g1162 = (((g112) & (!g199) & (!sk[28]) & (!g547)) + ((g112) & (!g199) & (!sk[28]) & (g547)) + ((g112) & (!g199) & (sk[28]) & (!g547)) + ((g112) & (g199) & (!sk[28]) & (!g547)) + ((g112) & (g199) & (!sk[28]) & (g547)) + ((g112) & (g199) & (sk[28]) & (!g547)) + ((g112) & (g199) & (sk[28]) & (g547)));
	assign g1163 = (((!g101) & (!g151) & (!sk[29]) & (!g1064) & (!g1161) & (g1162)) + ((!g101) & (!g151) & (!sk[29]) & (!g1064) & (g1161) & (g1162)) + ((!g101) & (!g151) & (!sk[29]) & (g1064) & (!g1161) & (g1162)) + ((!g101) & (!g151) & (!sk[29]) & (g1064) & (g1161) & (g1162)) + ((!g101) & (!g151) & (sk[29]) & (!g1064) & (!g1161) & (!g1162)) + ((!g101) & (!g151) & (sk[29]) & (!g1064) & (g1161) & (!g1162)) + ((!g101) & (!g151) & (sk[29]) & (g1064) & (!g1161) & (!g1162)) + ((!g101) & (!g151) & (sk[29]) & (g1064) & (g1161) & (!g1162)) + ((!g101) & (g151) & (!sk[29]) & (!g1064) & (!g1161) & (g1162)) + ((!g101) & (g151) & (!sk[29]) & (!g1064) & (g1161) & (g1162)) + ((!g101) & (g151) & (!sk[29]) & (g1064) & (!g1161) & (g1162)) + ((!g101) & (g151) & (!sk[29]) & (g1064) & (g1161) & (g1162)) + ((!g101) & (g151) & (sk[29]) & (!g1064) & (g1161) & (!g1162)) + ((!g101) & (g151) & (sk[29]) & (g1064) & (g1161) & (!g1162)) + ((g101) & (!g151) & (!sk[29]) & (!g1064) & (!g1161) & (!g1162)) + ((g101) & (!g151) & (!sk[29]) & (!g1064) & (!g1161) & (g1162)) + ((g101) & (!g151) & (!sk[29]) & (!g1064) & (g1161) & (!g1162)) + ((g101) & (!g151) & (!sk[29]) & (!g1064) & (g1161) & (g1162)) + ((g101) & (!g151) & (!sk[29]) & (g1064) & (!g1161) & (!g1162)) + ((g101) & (!g151) & (!sk[29]) & (g1064) & (!g1161) & (g1162)) + ((g101) & (!g151) & (!sk[29]) & (g1064) & (g1161) & (!g1162)) + ((g101) & (!g151) & (!sk[29]) & (g1064) & (g1161) & (g1162)) + ((g101) & (!g151) & (sk[29]) & (g1064) & (!g1161) & (!g1162)) + ((g101) & (!g151) & (sk[29]) & (g1064) & (g1161) & (!g1162)) + ((g101) & (g151) & (!sk[29]) & (!g1064) & (!g1161) & (!g1162)) + ((g101) & (g151) & (!sk[29]) & (!g1064) & (!g1161) & (g1162)) + ((g101) & (g151) & (!sk[29]) & (!g1064) & (g1161) & (!g1162)) + ((g101) & (g151) & (!sk[29]) & (!g1064) & (g1161) & (g1162)) + ((g101) & (g151) & (!sk[29]) & (g1064) & (!g1161) & (!g1162)) + ((g101) & (g151) & (!sk[29]) & (g1064) & (!g1161) & (g1162)) + ((g101) & (g151) & (!sk[29]) & (g1064) & (g1161) & (!g1162)) + ((g101) & (g151) & (!sk[29]) & (g1064) & (g1161) & (g1162)) + ((g101) & (g151) & (sk[29]) & (g1064) & (g1161) & (!g1162)));
	assign g1164 = (((g6) & (!i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g101)) + ((g6) & (!i_15_) & (!i_14_) & (i_12_) & (i_13_) & (g101)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g101)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (i_13_) & (g101)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (i_13_) & (g101)) + ((g6) & (i_15_) & (!i_14_) & (!i_12_) & (!i_13_) & (g101)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g101)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (i_13_) & (g101)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g101)));
	assign g1165 = (((!i_8_) & (!sk[31]) & (!g108) & (!g201) & (!g703) & (g908)) + ((!i_8_) & (!sk[31]) & (!g108) & (!g201) & (g703) & (g908)) + ((!i_8_) & (!sk[31]) & (!g108) & (g201) & (!g703) & (g908)) + ((!i_8_) & (!sk[31]) & (!g108) & (g201) & (g703) & (g908)) + ((!i_8_) & (!sk[31]) & (g108) & (!g201) & (!g703) & (g908)) + ((!i_8_) & (!sk[31]) & (g108) & (!g201) & (g703) & (g908)) + ((!i_8_) & (!sk[31]) & (g108) & (g201) & (!g703) & (g908)) + ((!i_8_) & (!sk[31]) & (g108) & (g201) & (g703) & (g908)) + ((i_8_) & (!sk[31]) & (!g108) & (!g201) & (!g703) & (!g908)) + ((i_8_) & (!sk[31]) & (!g108) & (!g201) & (!g703) & (g908)) + ((i_8_) & (!sk[31]) & (!g108) & (!g201) & (g703) & (!g908)) + ((i_8_) & (!sk[31]) & (!g108) & (!g201) & (g703) & (g908)) + ((i_8_) & (!sk[31]) & (!g108) & (g201) & (!g703) & (!g908)) + ((i_8_) & (!sk[31]) & (!g108) & (g201) & (!g703) & (g908)) + ((i_8_) & (!sk[31]) & (!g108) & (g201) & (g703) & (!g908)) + ((i_8_) & (!sk[31]) & (!g108) & (g201) & (g703) & (g908)) + ((i_8_) & (!sk[31]) & (g108) & (!g201) & (!g703) & (!g908)) + ((i_8_) & (!sk[31]) & (g108) & (!g201) & (!g703) & (g908)) + ((i_8_) & (!sk[31]) & (g108) & (!g201) & (g703) & (!g908)) + ((i_8_) & (!sk[31]) & (g108) & (!g201) & (g703) & (g908)) + ((i_8_) & (!sk[31]) & (g108) & (g201) & (!g703) & (!g908)) + ((i_8_) & (!sk[31]) & (g108) & (g201) & (!g703) & (g908)) + ((i_8_) & (!sk[31]) & (g108) & (g201) & (g703) & (!g908)) + ((i_8_) & (!sk[31]) & (g108) & (g201) & (g703) & (g908)) + ((i_8_) & (sk[31]) & (g108) & (!g201) & (!g703) & (!g908)) + ((i_8_) & (sk[31]) & (g108) & (!g201) & (!g703) & (g908)) + ((i_8_) & (sk[31]) & (g108) & (!g201) & (g703) & (!g908)) + ((i_8_) & (sk[31]) & (g108) & (!g201) & (g703) & (g908)) + ((i_8_) & (sk[31]) & (g108) & (g201) & (!g703) & (g908)) + ((i_8_) & (sk[31]) & (g108) & (g201) & (g703) & (!g908)) + ((i_8_) & (sk[31]) & (g108) & (g201) & (g703) & (g908)));
	assign g1166 = (((!g101) & (!g199) & (!g120) & (!g547) & (!sk[32]) & (g1165)) + ((!g101) & (!g199) & (!g120) & (!g547) & (sk[32]) & (!g1165)) + ((!g101) & (!g199) & (!g120) & (g547) & (!sk[32]) & (g1165)) + ((!g101) & (!g199) & (!g120) & (g547) & (sk[32]) & (!g1165)) + ((!g101) & (!g199) & (g120) & (!g547) & (!sk[32]) & (g1165)) + ((!g101) & (!g199) & (g120) & (!g547) & (sk[32]) & (!g1165)) + ((!g101) & (!g199) & (g120) & (g547) & (!sk[32]) & (g1165)) + ((!g101) & (!g199) & (g120) & (g547) & (sk[32]) & (!g1165)) + ((!g101) & (g199) & (!g120) & (!g547) & (!sk[32]) & (g1165)) + ((!g101) & (g199) & (!g120) & (!g547) & (sk[32]) & (!g1165)) + ((!g101) & (g199) & (!g120) & (g547) & (!sk[32]) & (g1165)) + ((!g101) & (g199) & (!g120) & (g547) & (sk[32]) & (!g1165)) + ((!g101) & (g199) & (g120) & (!g547) & (!sk[32]) & (g1165)) + ((!g101) & (g199) & (g120) & (!g547) & (sk[32]) & (!g1165)) + ((!g101) & (g199) & (g120) & (g547) & (!sk[32]) & (g1165)) + ((!g101) & (g199) & (g120) & (g547) & (sk[32]) & (!g1165)) + ((g101) & (!g199) & (!g120) & (!g547) & (!sk[32]) & (!g1165)) + ((g101) & (!g199) & (!g120) & (!g547) & (!sk[32]) & (g1165)) + ((g101) & (!g199) & (!g120) & (g547) & (!sk[32]) & (!g1165)) + ((g101) & (!g199) & (!g120) & (g547) & (!sk[32]) & (g1165)) + ((g101) & (!g199) & (g120) & (!g547) & (!sk[32]) & (!g1165)) + ((g101) & (!g199) & (g120) & (!g547) & (!sk[32]) & (g1165)) + ((g101) & (!g199) & (g120) & (g547) & (!sk[32]) & (!g1165)) + ((g101) & (!g199) & (g120) & (g547) & (!sk[32]) & (g1165)) + ((g101) & (!g199) & (g120) & (g547) & (sk[32]) & (!g1165)) + ((g101) & (g199) & (!g120) & (!g547) & (!sk[32]) & (!g1165)) + ((g101) & (g199) & (!g120) & (!g547) & (!sk[32]) & (g1165)) + ((g101) & (g199) & (!g120) & (g547) & (!sk[32]) & (!g1165)) + ((g101) & (g199) & (!g120) & (g547) & (!sk[32]) & (g1165)) + ((g101) & (g199) & (g120) & (!g547) & (!sk[32]) & (!g1165)) + ((g101) & (g199) & (g120) & (!g547) & (!sk[32]) & (g1165)) + ((g101) & (g199) & (g120) & (g547) & (!sk[32]) & (!g1165)) + ((g101) & (g199) & (g120) & (g547) & (!sk[32]) & (g1165)));
	assign g1167 = (((!g1065) & (!g1158) & (!g1160) & (g1163) & (!g1164) & (g1166)));
	assign g1168 = (((i_12_) & (!i_13_) & (!sk[34]) & (!g93)) + ((i_12_) & (!i_13_) & (!sk[34]) & (g93)) + ((i_12_) & (i_13_) & (!sk[34]) & (!g93)) + ((i_12_) & (i_13_) & (!sk[34]) & (g93)) + ((i_12_) & (i_13_) & (sk[34]) & (!g93)));
	assign g1169 = (((!sk[35]) & (g13) & (!g115) & (!g711)) + ((!sk[35]) & (g13) & (!g115) & (g711)) + ((!sk[35]) & (g13) & (g115) & (!g711)) + ((!sk[35]) & (g13) & (g115) & (g711)) + ((sk[35]) & (!g13) & (!g115) & (g711)) + ((sk[35]) & (g13) & (!g115) & (!g711)) + ((sk[35]) & (g13) & (!g115) & (g711)));
	assign g1170 = (((!i_8_) & (!sk[36]) & (!g264) & (!g100) & (!g103) & (g1169)) + ((!i_8_) & (!sk[36]) & (!g264) & (!g100) & (g103) & (g1169)) + ((!i_8_) & (!sk[36]) & (!g264) & (g100) & (!g103) & (g1169)) + ((!i_8_) & (!sk[36]) & (!g264) & (g100) & (g103) & (g1169)) + ((!i_8_) & (!sk[36]) & (g264) & (!g100) & (!g103) & (g1169)) + ((!i_8_) & (!sk[36]) & (g264) & (!g100) & (g103) & (g1169)) + ((!i_8_) & (!sk[36]) & (g264) & (g100) & (!g103) & (g1169)) + ((!i_8_) & (!sk[36]) & (g264) & (g100) & (g103) & (g1169)) + ((!i_8_) & (sk[36]) & (!g264) & (!g100) & (!g103) & (!g1169)) + ((!i_8_) & (sk[36]) & (!g264) & (!g100) & (g103) & (!g1169)) + ((!i_8_) & (sk[36]) & (!g264) & (g100) & (!g103) & (!g1169)) + ((!i_8_) & (sk[36]) & (!g264) & (g100) & (g103) & (!g1169)) + ((!i_8_) & (sk[36]) & (g264) & (!g100) & (!g103) & (!g1169)) + ((!i_8_) & (sk[36]) & (g264) & (!g100) & (g103) & (!g1169)) + ((!i_8_) & (sk[36]) & (g264) & (g100) & (!g103) & (!g1169)) + ((!i_8_) & (sk[36]) & (g264) & (g100) & (g103) & (!g1169)) + ((i_8_) & (!sk[36]) & (!g264) & (!g100) & (!g103) & (!g1169)) + ((i_8_) & (!sk[36]) & (!g264) & (!g100) & (!g103) & (g1169)) + ((i_8_) & (!sk[36]) & (!g264) & (!g100) & (g103) & (!g1169)) + ((i_8_) & (!sk[36]) & (!g264) & (!g100) & (g103) & (g1169)) + ((i_8_) & (!sk[36]) & (!g264) & (g100) & (!g103) & (!g1169)) + ((i_8_) & (!sk[36]) & (!g264) & (g100) & (!g103) & (g1169)) + ((i_8_) & (!sk[36]) & (!g264) & (g100) & (g103) & (!g1169)) + ((i_8_) & (!sk[36]) & (!g264) & (g100) & (g103) & (g1169)) + ((i_8_) & (!sk[36]) & (g264) & (!g100) & (!g103) & (!g1169)) + ((i_8_) & (!sk[36]) & (g264) & (!g100) & (!g103) & (g1169)) + ((i_8_) & (!sk[36]) & (g264) & (!g100) & (g103) & (!g1169)) + ((i_8_) & (!sk[36]) & (g264) & (!g100) & (g103) & (g1169)) + ((i_8_) & (!sk[36]) & (g264) & (g100) & (!g103) & (!g1169)) + ((i_8_) & (!sk[36]) & (g264) & (g100) & (!g103) & (g1169)) + ((i_8_) & (!sk[36]) & (g264) & (g100) & (g103) & (!g1169)) + ((i_8_) & (!sk[36]) & (g264) & (g100) & (g103) & (g1169)) + ((i_8_) & (sk[36]) & (!g264) & (!g100) & (!g103) & (!g1169)) + ((i_8_) & (sk[36]) & (!g264) & (!g100) & (g103) & (!g1169)) + ((i_8_) & (sk[36]) & (!g264) & (g100) & (g103) & (!g1169)) + ((i_8_) & (sk[36]) & (g264) & (!g100) & (!g103) & (!g1169)) + ((i_8_) & (sk[36]) & (g264) & (!g100) & (g103) & (!g1169)));
	assign g1171 = (((!g20) & (g101) & (!g173) & (!g806) & (!g1168) & (!g1170)) + ((!g20) & (g101) & (!g173) & (!g806) & (!g1168) & (g1170)) + ((!g20) & (g101) & (!g173) & (!g806) & (g1168) & (!g1170)) + ((!g20) & (g101) & (!g173) & (!g806) & (g1168) & (g1170)) + ((!g20) & (g101) & (!g173) & (g806) & (!g1168) & (!g1170)) + ((!g20) & (g101) & (!g173) & (g806) & (!g1168) & (g1170)) + ((!g20) & (g101) & (!g173) & (g806) & (g1168) & (!g1170)) + ((!g20) & (g101) & (!g173) & (g806) & (g1168) & (g1170)) + ((!g20) & (g101) & (g173) & (!g806) & (!g1168) & (!g1170)) + ((!g20) & (g101) & (g173) & (!g806) & (!g1168) & (g1170)) + ((!g20) & (g101) & (g173) & (!g806) & (g1168) & (!g1170)) + ((!g20) & (g101) & (g173) & (!g806) & (g1168) & (g1170)) + ((!g20) & (g101) & (g173) & (g806) & (!g1168) & (!g1170)) + ((!g20) & (g101) & (g173) & (g806) & (!g1168) & (g1170)) + ((!g20) & (g101) & (g173) & (g806) & (g1168) & (!g1170)) + ((!g20) & (g101) & (g173) & (g806) & (g1168) & (g1170)) + ((g20) & (g101) & (!g173) & (!g806) & (!g1168) & (!g1170)) + ((g20) & (g101) & (!g173) & (!g806) & (g1168) & (!g1170)) + ((g20) & (g101) & (!g173) & (!g806) & (g1168) & (g1170)) + ((g20) & (g101) & (!g173) & (g806) & (!g1168) & (!g1170)) + ((g20) & (g101) & (!g173) & (g806) & (!g1168) & (g1170)) + ((g20) & (g101) & (!g173) & (g806) & (g1168) & (!g1170)) + ((g20) & (g101) & (!g173) & (g806) & (g1168) & (g1170)) + ((g20) & (g101) & (g173) & (!g806) & (!g1168) & (!g1170)) + ((g20) & (g101) & (g173) & (!g806) & (!g1168) & (g1170)) + ((g20) & (g101) & (g173) & (!g806) & (g1168) & (!g1170)) + ((g20) & (g101) & (g173) & (!g806) & (g1168) & (g1170)) + ((g20) & (g101) & (g173) & (g806) & (!g1168) & (!g1170)) + ((g20) & (g101) & (g173) & (g806) & (!g1168) & (g1170)) + ((g20) & (g101) & (g173) & (g806) & (g1168) & (!g1170)) + ((g20) & (g101) & (g173) & (g806) & (g1168) & (g1170)));
	assign g1172 = (((!g145) & (!g261) & (!g524) & (!g525) & (!g710) & (!g1122)) + ((!g145) & (!g261) & (!g524) & (!g525) & (!g710) & (g1122)) + ((!g145) & (!g261) & (!g524) & (!g525) & (g710) & (!g1122)) + ((!g145) & (!g261) & (!g524) & (!g525) & (g710) & (g1122)) + ((g145) & (!g261) & (!g524) & (!g525) & (!g710) & (g1122)));
	assign g1173 = (((!g843) & (g845) & (g847) & (g851) & (!g1171) & (g1172)));
	assign g1174 = (((!g112) & (!g216) & (g120) & (!sk[40]) & (g485)) + ((!g112) & (g216) & (!g120) & (!sk[40]) & (!g485)) + ((!g112) & (g216) & (!g120) & (!sk[40]) & (g485)) + ((!g112) & (g216) & (g120) & (!sk[40]) & (!g485)) + ((!g112) & (g216) & (g120) & (!sk[40]) & (g485)) + ((g112) & (!g216) & (!g120) & (sk[40]) & (!g485)) + ((g112) & (!g216) & (!g120) & (sk[40]) & (g485)) + ((g112) & (!g216) & (g120) & (!sk[40]) & (!g485)) + ((g112) & (!g216) & (g120) & (!sk[40]) & (g485)) + ((g112) & (!g216) & (g120) & (sk[40]) & (g485)) + ((g112) & (g216) & (!g120) & (!sk[40]) & (!g485)) + ((g112) & (g216) & (!g120) & (!sk[40]) & (g485)) + ((g112) & (g216) & (!g120) & (sk[40]) & (!g485)) + ((g112) & (g216) & (!g120) & (sk[40]) & (g485)) + ((g112) & (g216) & (g120) & (!sk[40]) & (!g485)) + ((g112) & (g216) & (g120) & (!sk[40]) & (g485)) + ((g112) & (g216) & (g120) & (sk[40]) & (!g485)) + ((g112) & (g216) & (g120) & (sk[40]) & (g485)));
	assign g1175 = (((!g136) & (!sk[41]) & (!g226) & (!g506) & (!g670) & (g1001)) + ((!g136) & (!sk[41]) & (!g226) & (!g506) & (g670) & (g1001)) + ((!g136) & (!sk[41]) & (!g226) & (g506) & (!g670) & (g1001)) + ((!g136) & (!sk[41]) & (!g226) & (g506) & (g670) & (g1001)) + ((!g136) & (!sk[41]) & (g226) & (!g506) & (!g670) & (g1001)) + ((!g136) & (!sk[41]) & (g226) & (!g506) & (g670) & (g1001)) + ((!g136) & (!sk[41]) & (g226) & (g506) & (!g670) & (g1001)) + ((!g136) & (!sk[41]) & (g226) & (g506) & (g670) & (g1001)) + ((g136) & (!sk[41]) & (!g226) & (!g506) & (!g670) & (!g1001)) + ((g136) & (!sk[41]) & (!g226) & (!g506) & (!g670) & (g1001)) + ((g136) & (!sk[41]) & (!g226) & (!g506) & (g670) & (!g1001)) + ((g136) & (!sk[41]) & (!g226) & (!g506) & (g670) & (g1001)) + ((g136) & (!sk[41]) & (!g226) & (g506) & (!g670) & (!g1001)) + ((g136) & (!sk[41]) & (!g226) & (g506) & (!g670) & (g1001)) + ((g136) & (!sk[41]) & (!g226) & (g506) & (g670) & (!g1001)) + ((g136) & (!sk[41]) & (!g226) & (g506) & (g670) & (g1001)) + ((g136) & (!sk[41]) & (g226) & (!g506) & (!g670) & (!g1001)) + ((g136) & (!sk[41]) & (g226) & (!g506) & (!g670) & (g1001)) + ((g136) & (!sk[41]) & (g226) & (!g506) & (g670) & (!g1001)) + ((g136) & (!sk[41]) & (g226) & (!g506) & (g670) & (g1001)) + ((g136) & (!sk[41]) & (g226) & (g506) & (!g670) & (!g1001)) + ((g136) & (!sk[41]) & (g226) & (g506) & (!g670) & (g1001)) + ((g136) & (!sk[41]) & (g226) & (g506) & (g670) & (!g1001)) + ((g136) & (!sk[41]) & (g226) & (g506) & (g670) & (g1001)) + ((g136) & (sk[41]) & (!g226) & (!g506) & (!g670) & (!g1001)) + ((g136) & (sk[41]) & (!g226) & (!g506) & (!g670) & (g1001)) + ((g136) & (sk[41]) & (!g226) & (!g506) & (g670) & (!g1001)) + ((g136) & (sk[41]) & (!g226) & (!g506) & (g670) & (g1001)) + ((g136) & (sk[41]) & (!g226) & (g506) & (!g670) & (!g1001)) + ((g136) & (sk[41]) & (!g226) & (g506) & (!g670) & (g1001)) + ((g136) & (sk[41]) & (!g226) & (g506) & (g670) & (!g1001)) + ((g136) & (sk[41]) & (!g226) & (g506) & (g670) & (g1001)) + ((g136) & (sk[41]) & (g226) & (!g506) & (!g670) & (!g1001)) + ((g136) & (sk[41]) & (g226) & (!g506) & (g670) & (!g1001)) + ((g136) & (sk[41]) & (g226) & (!g506) & (g670) & (g1001)) + ((g136) & (sk[41]) & (g226) & (g506) & (!g670) & (!g1001)) + ((g136) & (sk[41]) & (g226) & (g506) & (!g670) & (g1001)) + ((g136) & (sk[41]) & (g226) & (g506) & (g670) & (!g1001)) + ((g136) & (sk[41]) & (g226) & (g506) & (g670) & (g1001)));
	assign g1176 = (((!i_8_) & (!g135) & (!g114) & (!sk[42]) & (!g560) & (g464)) + ((!i_8_) & (!g135) & (!g114) & (!sk[42]) & (g560) & (g464)) + ((!i_8_) & (!g135) & (g114) & (!sk[42]) & (!g560) & (g464)) + ((!i_8_) & (!g135) & (g114) & (!sk[42]) & (g560) & (g464)) + ((!i_8_) & (g135) & (!g114) & (!sk[42]) & (!g560) & (g464)) + ((!i_8_) & (g135) & (!g114) & (!sk[42]) & (g560) & (g464)) + ((!i_8_) & (g135) & (g114) & (!sk[42]) & (!g560) & (g464)) + ((!i_8_) & (g135) & (g114) & (!sk[42]) & (g560) & (g464)) + ((i_8_) & (!g135) & (!g114) & (!sk[42]) & (!g560) & (!g464)) + ((i_8_) & (!g135) & (!g114) & (!sk[42]) & (!g560) & (g464)) + ((i_8_) & (!g135) & (!g114) & (!sk[42]) & (g560) & (!g464)) + ((i_8_) & (!g135) & (!g114) & (!sk[42]) & (g560) & (g464)) + ((i_8_) & (!g135) & (g114) & (!sk[42]) & (!g560) & (!g464)) + ((i_8_) & (!g135) & (g114) & (!sk[42]) & (!g560) & (g464)) + ((i_8_) & (!g135) & (g114) & (!sk[42]) & (g560) & (!g464)) + ((i_8_) & (!g135) & (g114) & (!sk[42]) & (g560) & (g464)) + ((i_8_) & (g135) & (!g114) & (!sk[42]) & (!g560) & (!g464)) + ((i_8_) & (g135) & (!g114) & (!sk[42]) & (!g560) & (g464)) + ((i_8_) & (g135) & (!g114) & (!sk[42]) & (g560) & (!g464)) + ((i_8_) & (g135) & (!g114) & (!sk[42]) & (g560) & (g464)) + ((i_8_) & (g135) & (!g114) & (sk[42]) & (!g560) & (!g464)) + ((i_8_) & (g135) & (!g114) & (sk[42]) & (g560) & (!g464)) + ((i_8_) & (g135) & (!g114) & (sk[42]) & (g560) & (g464)) + ((i_8_) & (g135) & (g114) & (!sk[42]) & (!g560) & (!g464)) + ((i_8_) & (g135) & (g114) & (!sk[42]) & (!g560) & (g464)) + ((i_8_) & (g135) & (g114) & (!sk[42]) & (g560) & (!g464)) + ((i_8_) & (g135) & (g114) & (!sk[42]) & (g560) & (g464)) + ((i_8_) & (g135) & (g114) & (sk[42]) & (!g560) & (!g464)) + ((i_8_) & (g135) & (g114) & (sk[42]) & (!g560) & (g464)) + ((i_8_) & (g135) & (g114) & (sk[42]) & (g560) & (!g464)) + ((i_8_) & (g135) & (g114) & (sk[42]) & (g560) & (g464)));
	assign g1177 = (((!g21) & (!sk[43]) & (!g136) & (!g177) & (!g120) & (g1176)) + ((!g21) & (!sk[43]) & (!g136) & (!g177) & (g120) & (g1176)) + ((!g21) & (!sk[43]) & (!g136) & (g177) & (!g120) & (g1176)) + ((!g21) & (!sk[43]) & (!g136) & (g177) & (g120) & (g1176)) + ((!g21) & (!sk[43]) & (g136) & (!g177) & (!g120) & (g1176)) + ((!g21) & (!sk[43]) & (g136) & (!g177) & (g120) & (g1176)) + ((!g21) & (!sk[43]) & (g136) & (g177) & (!g120) & (g1176)) + ((!g21) & (!sk[43]) & (g136) & (g177) & (g120) & (g1176)) + ((!g21) & (sk[43]) & (!g136) & (!g177) & (!g120) & (!g1176)) + ((!g21) & (sk[43]) & (!g136) & (!g177) & (g120) & (!g1176)) + ((!g21) & (sk[43]) & (!g136) & (g177) & (!g120) & (!g1176)) + ((!g21) & (sk[43]) & (!g136) & (g177) & (g120) & (!g1176)) + ((!g21) & (sk[43]) & (g136) & (!g177) & (g120) & (!g1176)) + ((g21) & (!sk[43]) & (!g136) & (!g177) & (!g120) & (!g1176)) + ((g21) & (!sk[43]) & (!g136) & (!g177) & (!g120) & (g1176)) + ((g21) & (!sk[43]) & (!g136) & (!g177) & (g120) & (!g1176)) + ((g21) & (!sk[43]) & (!g136) & (!g177) & (g120) & (g1176)) + ((g21) & (!sk[43]) & (!g136) & (g177) & (!g120) & (!g1176)) + ((g21) & (!sk[43]) & (!g136) & (g177) & (!g120) & (g1176)) + ((g21) & (!sk[43]) & (!g136) & (g177) & (g120) & (!g1176)) + ((g21) & (!sk[43]) & (!g136) & (g177) & (g120) & (g1176)) + ((g21) & (!sk[43]) & (g136) & (!g177) & (!g120) & (!g1176)) + ((g21) & (!sk[43]) & (g136) & (!g177) & (!g120) & (g1176)) + ((g21) & (!sk[43]) & (g136) & (!g177) & (g120) & (!g1176)) + ((g21) & (!sk[43]) & (g136) & (!g177) & (g120) & (g1176)) + ((g21) & (!sk[43]) & (g136) & (g177) & (!g120) & (!g1176)) + ((g21) & (!sk[43]) & (g136) & (g177) & (!g120) & (g1176)) + ((g21) & (!sk[43]) & (g136) & (g177) & (g120) & (!g1176)) + ((g21) & (!sk[43]) & (g136) & (g177) & (g120) & (g1176)) + ((g21) & (sk[43]) & (!g136) & (!g177) & (!g120) & (!g1176)) + ((g21) & (sk[43]) & (!g136) & (!g177) & (g120) & (!g1176)) + ((g21) & (sk[43]) & (!g136) & (g177) & (!g120) & (!g1176)) + ((g21) & (sk[43]) & (!g136) & (g177) & (g120) & (!g1176)));
	assign g1178 = (((!sk[44]) & (!g608) & (!g1174) & (g1175) & (g1177)) + ((!sk[44]) & (!g608) & (g1174) & (!g1175) & (!g1177)) + ((!sk[44]) & (!g608) & (g1174) & (!g1175) & (g1177)) + ((!sk[44]) & (!g608) & (g1174) & (g1175) & (!g1177)) + ((!sk[44]) & (!g608) & (g1174) & (g1175) & (g1177)) + ((!sk[44]) & (g608) & (!g1174) & (g1175) & (!g1177)) + ((!sk[44]) & (g608) & (!g1174) & (g1175) & (g1177)) + ((!sk[44]) & (g608) & (g1174) & (!g1175) & (!g1177)) + ((!sk[44]) & (g608) & (g1174) & (!g1175) & (g1177)) + ((!sk[44]) & (g608) & (g1174) & (g1175) & (!g1177)) + ((!sk[44]) & (g608) & (g1174) & (g1175) & (g1177)) + ((sk[44]) & (!g608) & (!g1174) & (!g1175) & (g1177)));
	assign g1179 = (((!i_8_) & (!g108) & (!sk[45]) & (g630) & (g980)) + ((!i_8_) & (g108) & (!sk[45]) & (!g630) & (!g980)) + ((!i_8_) & (g108) & (!sk[45]) & (!g630) & (g980)) + ((!i_8_) & (g108) & (!sk[45]) & (g630) & (!g980)) + ((!i_8_) & (g108) & (!sk[45]) & (g630) & (g980)) + ((i_8_) & (!g108) & (!sk[45]) & (g630) & (!g980)) + ((i_8_) & (!g108) & (!sk[45]) & (g630) & (g980)) + ((i_8_) & (g108) & (!sk[45]) & (!g630) & (!g980)) + ((i_8_) & (g108) & (!sk[45]) & (!g630) & (g980)) + ((i_8_) & (g108) & (!sk[45]) & (g630) & (!g980)) + ((i_8_) & (g108) & (!sk[45]) & (g630) & (g980)) + ((i_8_) & (g108) & (sk[45]) & (!g630) & (!g980)) + ((i_8_) & (g108) & (sk[45]) & (g630) & (!g980)) + ((i_8_) & (g108) & (sk[45]) & (g630) & (g980)));
	assign g1180 = (((!g47) & (!sk[46]) & (!g101) & (!g172) & (!g142) & (g1179)) + ((!g47) & (!sk[46]) & (!g101) & (!g172) & (g142) & (g1179)) + ((!g47) & (!sk[46]) & (!g101) & (g172) & (!g142) & (g1179)) + ((!g47) & (!sk[46]) & (!g101) & (g172) & (g142) & (g1179)) + ((!g47) & (!sk[46]) & (g101) & (!g172) & (!g142) & (g1179)) + ((!g47) & (!sk[46]) & (g101) & (!g172) & (g142) & (g1179)) + ((!g47) & (!sk[46]) & (g101) & (g172) & (!g142) & (g1179)) + ((!g47) & (!sk[46]) & (g101) & (g172) & (g142) & (g1179)) + ((!g47) & (sk[46]) & (!g101) & (!g172) & (!g142) & (!g1179)) + ((!g47) & (sk[46]) & (!g101) & (!g172) & (g142) & (!g1179)) + ((!g47) & (sk[46]) & (!g101) & (g172) & (!g142) & (!g1179)) + ((!g47) & (sk[46]) & (!g101) & (g172) & (g142) & (!g1179)) + ((!g47) & (sk[46]) & (g101) & (!g172) & (!g142) & (!g1179)) + ((g47) & (!sk[46]) & (!g101) & (!g172) & (!g142) & (!g1179)) + ((g47) & (!sk[46]) & (!g101) & (!g172) & (!g142) & (g1179)) + ((g47) & (!sk[46]) & (!g101) & (!g172) & (g142) & (!g1179)) + ((g47) & (!sk[46]) & (!g101) & (!g172) & (g142) & (g1179)) + ((g47) & (!sk[46]) & (!g101) & (g172) & (!g142) & (!g1179)) + ((g47) & (!sk[46]) & (!g101) & (g172) & (!g142) & (g1179)) + ((g47) & (!sk[46]) & (!g101) & (g172) & (g142) & (!g1179)) + ((g47) & (!sk[46]) & (!g101) & (g172) & (g142) & (g1179)) + ((g47) & (!sk[46]) & (g101) & (!g172) & (!g142) & (!g1179)) + ((g47) & (!sk[46]) & (g101) & (!g172) & (!g142) & (g1179)) + ((g47) & (!sk[46]) & (g101) & (!g172) & (g142) & (!g1179)) + ((g47) & (!sk[46]) & (g101) & (!g172) & (g142) & (g1179)) + ((g47) & (!sk[46]) & (g101) & (g172) & (!g142) & (!g1179)) + ((g47) & (!sk[46]) & (g101) & (g172) & (!g142) & (g1179)) + ((g47) & (!sk[46]) & (g101) & (g172) & (g142) & (!g1179)) + ((g47) & (!sk[46]) & (g101) & (g172) & (g142) & (g1179)) + ((g47) & (sk[46]) & (!g101) & (!g172) & (!g142) & (!g1179)) + ((g47) & (sk[46]) & (!g101) & (!g172) & (g142) & (!g1179)) + ((g47) & (sk[46]) & (!g101) & (g172) & (!g142) & (!g1179)) + ((g47) & (sk[46]) & (!g101) & (g172) & (g142) & (!g1179)));
	assign g1181 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g102) & (g136) & (!g115)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g102) & (g136) & (!g115)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g102) & (g136) & (!g115)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g102) & (g136) & (g115)) + ((!i_14_) & (i_12_) & (!i_13_) & (g102) & (g136) & (!g115)) + ((!i_14_) & (i_12_) & (i_13_) & (!g102) & (g136) & (!g115)) + ((!i_14_) & (i_12_) & (i_13_) & (!g102) & (g136) & (g115)) + ((!i_14_) & (i_12_) & (i_13_) & (g102) & (g136) & (!g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g102) & (g136) & (!g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g102) & (g136) & (g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (g102) & (g136) & (!g115)) + ((i_14_) & (!i_12_) & (i_13_) & (!g102) & (g136) & (!g115)) + ((i_14_) & (!i_12_) & (i_13_) & (!g102) & (g136) & (g115)) + ((i_14_) & (i_12_) & (i_13_) & (!g102) & (g136) & (!g115)) + ((i_14_) & (i_12_) & (i_13_) & (!g102) & (g136) & (g115)));
	assign g1182 = (((!g1050) & (!g1071) & (!g1040) & (sk[48]) & (!g1066)) + ((!g1050) & (!g1071) & (g1040) & (!sk[48]) & (g1066)) + ((!g1050) & (g1071) & (!g1040) & (!sk[48]) & (!g1066)) + ((!g1050) & (g1071) & (!g1040) & (!sk[48]) & (g1066)) + ((!g1050) & (g1071) & (g1040) & (!sk[48]) & (!g1066)) + ((!g1050) & (g1071) & (g1040) & (!sk[48]) & (g1066)) + ((g1050) & (!g1071) & (g1040) & (!sk[48]) & (!g1066)) + ((g1050) & (!g1071) & (g1040) & (!sk[48]) & (g1066)) + ((g1050) & (g1071) & (!g1040) & (!sk[48]) & (!g1066)) + ((g1050) & (g1071) & (!g1040) & (!sk[48]) & (g1066)) + ((g1050) & (g1071) & (g1040) & (!sk[48]) & (!g1066)) + ((g1050) & (g1071) & (g1040) & (!sk[48]) & (g1066)));
	assign g1183 = (((!sk[49]) & (!g151) & (!g1127) & (g1099) & (g1132)) + ((!sk[49]) & (!g151) & (g1127) & (!g1099) & (!g1132)) + ((!sk[49]) & (!g151) & (g1127) & (!g1099) & (g1132)) + ((!sk[49]) & (!g151) & (g1127) & (g1099) & (!g1132)) + ((!sk[49]) & (!g151) & (g1127) & (g1099) & (g1132)) + ((!sk[49]) & (g151) & (!g1127) & (g1099) & (!g1132)) + ((!sk[49]) & (g151) & (!g1127) & (g1099) & (g1132)) + ((!sk[49]) & (g151) & (g1127) & (!g1099) & (!g1132)) + ((!sk[49]) & (g151) & (g1127) & (!g1099) & (g1132)) + ((!sk[49]) & (g151) & (g1127) & (g1099) & (!g1132)) + ((!sk[49]) & (g151) & (g1127) & (g1099) & (g1132)) + ((sk[49]) & (g151) & (!g1127) & (!g1099) & (!g1132)) + ((sk[49]) & (g151) & (!g1127) & (!g1099) & (g1132)) + ((sk[49]) & (g151) & (!g1127) & (g1099) & (g1132)) + ((sk[49]) & (g151) & (g1127) & (!g1099) & (!g1132)) + ((sk[49]) & (g151) & (g1127) & (!g1099) & (g1132)) + ((sk[49]) & (g151) & (g1127) & (g1099) & (!g1132)) + ((sk[49]) & (g151) & (g1127) & (g1099) & (g1132)));
	assign g1184 = (((!i_8_) & (!g100) & (!sk[50]) & (!g195) & (!g105) & (g532)) + ((!i_8_) & (!g100) & (!sk[50]) & (!g195) & (g105) & (g532)) + ((!i_8_) & (!g100) & (!sk[50]) & (g195) & (!g105) & (g532)) + ((!i_8_) & (!g100) & (!sk[50]) & (g195) & (g105) & (g532)) + ((!i_8_) & (!g100) & (sk[50]) & (!g195) & (!g105) & (!g532)) + ((!i_8_) & (!g100) & (sk[50]) & (!g195) & (g105) & (!g532)) + ((!i_8_) & (g100) & (!sk[50]) & (!g195) & (!g105) & (g532)) + ((!i_8_) & (g100) & (!sk[50]) & (!g195) & (g105) & (g532)) + ((!i_8_) & (g100) & (!sk[50]) & (g195) & (!g105) & (g532)) + ((!i_8_) & (g100) & (!sk[50]) & (g195) & (g105) & (g532)) + ((!i_8_) & (g100) & (sk[50]) & (!g195) & (!g105) & (!g532)) + ((!i_8_) & (g100) & (sk[50]) & (!g195) & (g105) & (!g532)) + ((i_8_) & (!g100) & (!sk[50]) & (!g195) & (!g105) & (!g532)) + ((i_8_) & (!g100) & (!sk[50]) & (!g195) & (!g105) & (g532)) + ((i_8_) & (!g100) & (!sk[50]) & (!g195) & (g105) & (!g532)) + ((i_8_) & (!g100) & (!sk[50]) & (!g195) & (g105) & (g532)) + ((i_8_) & (!g100) & (!sk[50]) & (g195) & (!g105) & (!g532)) + ((i_8_) & (!g100) & (!sk[50]) & (g195) & (!g105) & (g532)) + ((i_8_) & (!g100) & (!sk[50]) & (g195) & (g105) & (!g532)) + ((i_8_) & (!g100) & (!sk[50]) & (g195) & (g105) & (g532)) + ((i_8_) & (!g100) & (sk[50]) & (!g195) & (!g105) & (!g532)) + ((i_8_) & (!g100) & (sk[50]) & (!g195) & (g105) & (!g532)) + ((i_8_) & (g100) & (!sk[50]) & (!g195) & (!g105) & (!g532)) + ((i_8_) & (g100) & (!sk[50]) & (!g195) & (!g105) & (g532)) + ((i_8_) & (g100) & (!sk[50]) & (!g195) & (g105) & (!g532)) + ((i_8_) & (g100) & (!sk[50]) & (!g195) & (g105) & (g532)) + ((i_8_) & (g100) & (!sk[50]) & (g195) & (!g105) & (!g532)) + ((i_8_) & (g100) & (!sk[50]) & (g195) & (!g105) & (g532)) + ((i_8_) & (g100) & (!sk[50]) & (g195) & (g105) & (!g532)) + ((i_8_) & (g100) & (!sk[50]) & (g195) & (g105) & (g532)) + ((i_8_) & (g100) & (sk[50]) & (!g195) & (!g105) & (!g532)));
	assign g1185 = (((!sk[51]) & (g20) & (!g98) & (!g111)) + ((!sk[51]) & (g20) & (!g98) & (g111)) + ((!sk[51]) & (g20) & (g98) & (!g111)) + ((!sk[51]) & (g20) & (g98) & (g111)) + ((sk[51]) & (!g20) & (g98) & (g111)));
	assign g1186 = (((!i_8_) & (!g100) & (!g112) & (!g1185) & (!g835) & (!g1001)) + ((!i_8_) & (!g100) & (!g112) & (!g1185) & (!g835) & (g1001)) + ((!i_8_) & (!g100) & (!g112) & (!g1185) & (g835) & (!g1001)) + ((!i_8_) & (!g100) & (!g112) & (!g1185) & (g835) & (g1001)) + ((!i_8_) & (!g100) & (g112) & (!g1185) & (!g835) & (g1001)) + ((!i_8_) & (!g100) & (g112) & (!g1185) & (g835) & (g1001)) + ((!i_8_) & (g100) & (!g112) & (!g1185) & (!g835) & (!g1001)) + ((!i_8_) & (g100) & (!g112) & (!g1185) & (!g835) & (g1001)) + ((!i_8_) & (g100) & (!g112) & (!g1185) & (g835) & (!g1001)) + ((!i_8_) & (g100) & (!g112) & (!g1185) & (g835) & (g1001)) + ((!i_8_) & (g100) & (g112) & (!g1185) & (!g835) & (g1001)) + ((!i_8_) & (g100) & (g112) & (!g1185) & (g835) & (g1001)) + ((i_8_) & (!g100) & (!g112) & (!g1185) & (!g835) & (!g1001)) + ((i_8_) & (!g100) & (!g112) & (!g1185) & (!g835) & (g1001)) + ((i_8_) & (!g100) & (!g112) & (!g1185) & (g835) & (!g1001)) + ((i_8_) & (!g100) & (!g112) & (!g1185) & (g835) & (g1001)) + ((i_8_) & (!g100) & (g112) & (!g1185) & (!g835) & (g1001)) + ((i_8_) & (!g100) & (g112) & (!g1185) & (g835) & (g1001)) + ((i_8_) & (g100) & (!g112) & (!g1185) & (g835) & (!g1001)) + ((i_8_) & (g100) & (!g112) & (!g1185) & (g835) & (g1001)) + ((i_8_) & (g100) & (g112) & (!g1185) & (g835) & (g1001)));
	assign g1187 = (((!g101) & (!sk[53]) & (!g1019) & (!g1087) & (!g1184) & (g1186)) + ((!g101) & (!sk[53]) & (!g1019) & (!g1087) & (g1184) & (g1186)) + ((!g101) & (!sk[53]) & (!g1019) & (g1087) & (!g1184) & (g1186)) + ((!g101) & (!sk[53]) & (!g1019) & (g1087) & (g1184) & (g1186)) + ((!g101) & (!sk[53]) & (g1019) & (!g1087) & (!g1184) & (g1186)) + ((!g101) & (!sk[53]) & (g1019) & (!g1087) & (g1184) & (g1186)) + ((!g101) & (!sk[53]) & (g1019) & (g1087) & (!g1184) & (g1186)) + ((!g101) & (!sk[53]) & (g1019) & (g1087) & (g1184) & (g1186)) + ((!g101) & (sk[53]) & (!g1019) & (!g1087) & (!g1184) & (g1186)) + ((!g101) & (sk[53]) & (!g1019) & (!g1087) & (g1184) & (g1186)) + ((!g101) & (sk[53]) & (g1019) & (!g1087) & (!g1184) & (g1186)) + ((!g101) & (sk[53]) & (g1019) & (!g1087) & (g1184) & (g1186)) + ((g101) & (!sk[53]) & (!g1019) & (!g1087) & (!g1184) & (!g1186)) + ((g101) & (!sk[53]) & (!g1019) & (!g1087) & (!g1184) & (g1186)) + ((g101) & (!sk[53]) & (!g1019) & (!g1087) & (g1184) & (!g1186)) + ((g101) & (!sk[53]) & (!g1019) & (!g1087) & (g1184) & (g1186)) + ((g101) & (!sk[53]) & (!g1019) & (g1087) & (!g1184) & (!g1186)) + ((g101) & (!sk[53]) & (!g1019) & (g1087) & (!g1184) & (g1186)) + ((g101) & (!sk[53]) & (!g1019) & (g1087) & (g1184) & (!g1186)) + ((g101) & (!sk[53]) & (!g1019) & (g1087) & (g1184) & (g1186)) + ((g101) & (!sk[53]) & (g1019) & (!g1087) & (!g1184) & (!g1186)) + ((g101) & (!sk[53]) & (g1019) & (!g1087) & (!g1184) & (g1186)) + ((g101) & (!sk[53]) & (g1019) & (!g1087) & (g1184) & (!g1186)) + ((g101) & (!sk[53]) & (g1019) & (!g1087) & (g1184) & (g1186)) + ((g101) & (!sk[53]) & (g1019) & (g1087) & (!g1184) & (!g1186)) + ((g101) & (!sk[53]) & (g1019) & (g1087) & (!g1184) & (g1186)) + ((g101) & (!sk[53]) & (g1019) & (g1087) & (g1184) & (!g1186)) + ((g101) & (!sk[53]) & (g1019) & (g1087) & (g1184) & (g1186)) + ((g101) & (sk[53]) & (g1019) & (!g1087) & (g1184) & (g1186)));
	assign g1188 = (((!g1098) & (g1180) & (!g1181) & (g1182) & (!g1183) & (g1187)));
	assign g1189 = (((!g1147) & (g1156) & (g1167) & (g1173) & (g1178) & (g1188)));
	assign o_16_ = (((g73) & (!g420) & (!g490) & (!g664) & (!g1145) & (!g1189)) + ((g73) & (!g420) & (!g490) & (!g664) & (!g1145) & (g1189)) + ((g73) & (!g420) & (!g490) & (!g664) & (g1145) & (!g1189)) + ((g73) & (!g420) & (!g490) & (!g664) & (g1145) & (g1189)) + ((g73) & (!g420) & (!g490) & (g664) & (!g1145) & (!g1189)) + ((g73) & (!g420) & (!g490) & (g664) & (!g1145) & (g1189)) + ((g73) & (!g420) & (!g490) & (g664) & (g1145) & (!g1189)) + ((g73) & (!g420) & (!g490) & (g664) & (g1145) & (g1189)) + ((g73) & (!g420) & (g490) & (!g664) & (!g1145) & (!g1189)) + ((g73) & (!g420) & (g490) & (!g664) & (!g1145) & (g1189)) + ((g73) & (!g420) & (g490) & (!g664) & (g1145) & (!g1189)) + ((g73) & (!g420) & (g490) & (!g664) & (g1145) & (g1189)) + ((g73) & (!g420) & (g490) & (g664) & (!g1145) & (!g1189)) + ((g73) & (!g420) & (g490) & (g664) & (!g1145) & (g1189)) + ((g73) & (!g420) & (g490) & (g664) & (g1145) & (!g1189)) + ((g73) & (!g420) & (g490) & (g664) & (g1145) & (g1189)) + ((g73) & (g420) & (!g490) & (!g664) & (!g1145) & (!g1189)) + ((g73) & (g420) & (!g490) & (!g664) & (!g1145) & (g1189)) + ((g73) & (g420) & (!g490) & (!g664) & (g1145) & (!g1189)) + ((g73) & (g420) & (!g490) & (!g664) & (g1145) & (g1189)) + ((g73) & (g420) & (!g490) & (g664) & (!g1145) & (!g1189)) + ((g73) & (g420) & (!g490) & (g664) & (!g1145) & (g1189)) + ((g73) & (g420) & (!g490) & (g664) & (g1145) & (!g1189)) + ((g73) & (g420) & (!g490) & (g664) & (g1145) & (g1189)) + ((g73) & (g420) & (g490) & (!g664) & (!g1145) & (!g1189)) + ((g73) & (g420) & (g490) & (!g664) & (!g1145) & (g1189)) + ((g73) & (g420) & (g490) & (!g664) & (g1145) & (!g1189)) + ((g73) & (g420) & (g490) & (!g664) & (g1145) & (g1189)) + ((g73) & (g420) & (g490) & (g664) & (!g1145) & (!g1189)) + ((g73) & (g420) & (g490) & (g664) & (!g1145) & (g1189)) + ((g73) & (g420) & (g490) & (g664) & (g1145) & (!g1189)));
	assign g1191 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g109) & (g124)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g104) & (g109) & (g124)) + ((!i_14_) & (!i_12_) & (i_13_) & (g104) & (g109) & (!g124)) + ((!i_14_) & (!i_12_) & (i_13_) & (g104) & (g109) & (g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g104) & (g109) & (g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (g104) & (g109) & (!g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (g104) & (g109) & (g124)) + ((!i_14_) & (i_12_) & (i_13_) & (!g104) & (g109) & (g124)) + ((!i_14_) & (i_12_) & (i_13_) & (g104) & (g109) & (!g124)) + ((!i_14_) & (i_12_) & (i_13_) & (g104) & (g109) & (g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g109) & (g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (g104) & (g109) & (!g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (g104) & (g109) & (g124)) + ((i_14_) & (!i_12_) & (i_13_) & (!g104) & (g109) & (g124)) + ((i_14_) & (!i_12_) & (i_13_) & (g104) & (g109) & (!g124)) + ((i_14_) & (!i_12_) & (i_13_) & (g104) & (g109) & (g124)) + ((i_14_) & (i_12_) & (!i_13_) & (!g104) & (g109) & (g124)) + ((i_14_) & (i_12_) & (!i_13_) & (g104) & (g109) & (g124)) + ((i_14_) & (i_12_) & (i_13_) & (g104) & (g109) & (!g124)) + ((i_14_) & (i_12_) & (i_13_) & (g104) & (g109) & (g124)));
	assign g1192 = (((g6) & (!i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g145)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g145)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (i_13_) & (g145)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (i_13_) & (g145)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g145)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (i_13_) & (g145)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g145)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (i_13_) & (g145)) + ((g6) & (i_15_) & (i_14_) & (i_12_) & (!i_13_) & (g145)));
	assign g1193 = (((!g10) & (!sk[59]) & (!g99) & (!g109) & (!g92) & (g468)) + ((!g10) & (!sk[59]) & (!g99) & (!g109) & (g92) & (g468)) + ((!g10) & (!sk[59]) & (!g99) & (g109) & (!g92) & (g468)) + ((!g10) & (!sk[59]) & (!g99) & (g109) & (g92) & (g468)) + ((!g10) & (!sk[59]) & (g99) & (!g109) & (!g92) & (g468)) + ((!g10) & (!sk[59]) & (g99) & (!g109) & (g92) & (g468)) + ((!g10) & (!sk[59]) & (g99) & (g109) & (!g92) & (g468)) + ((!g10) & (!sk[59]) & (g99) & (g109) & (g92) & (g468)) + ((!g10) & (sk[59]) & (!g99) & (!g109) & (!g92) & (!g468)) + ((!g10) & (sk[59]) & (!g99) & (!g109) & (!g92) & (g468)) + ((!g10) & (sk[59]) & (!g99) & (!g109) & (g92) & (!g468)) + ((!g10) & (sk[59]) & (!g99) & (!g109) & (g92) & (g468)) + ((!g10) & (sk[59]) & (!g99) & (g109) & (!g92) & (!g468)) + ((!g10) & (sk[59]) & (!g99) & (g109) & (!g92) & (g468)) + ((!g10) & (sk[59]) & (!g99) & (g109) & (g92) & (!g468)) + ((!g10) & (sk[59]) & (!g99) & (g109) & (g92) & (g468)) + ((!g10) & (sk[59]) & (g99) & (!g109) & (g92) & (g468)) + ((!g10) & (sk[59]) & (g99) & (g109) & (g92) & (g468)) + ((g10) & (!sk[59]) & (!g99) & (!g109) & (!g92) & (!g468)) + ((g10) & (!sk[59]) & (!g99) & (!g109) & (!g92) & (g468)) + ((g10) & (!sk[59]) & (!g99) & (!g109) & (g92) & (!g468)) + ((g10) & (!sk[59]) & (!g99) & (!g109) & (g92) & (g468)) + ((g10) & (!sk[59]) & (!g99) & (g109) & (!g92) & (!g468)) + ((g10) & (!sk[59]) & (!g99) & (g109) & (!g92) & (g468)) + ((g10) & (!sk[59]) & (!g99) & (g109) & (g92) & (!g468)) + ((g10) & (!sk[59]) & (!g99) & (g109) & (g92) & (g468)) + ((g10) & (!sk[59]) & (g99) & (!g109) & (!g92) & (!g468)) + ((g10) & (!sk[59]) & (g99) & (!g109) & (!g92) & (g468)) + ((g10) & (!sk[59]) & (g99) & (!g109) & (g92) & (!g468)) + ((g10) & (!sk[59]) & (g99) & (!g109) & (g92) & (g468)) + ((g10) & (!sk[59]) & (g99) & (g109) & (!g92) & (!g468)) + ((g10) & (!sk[59]) & (g99) & (g109) & (!g92) & (g468)) + ((g10) & (!sk[59]) & (g99) & (g109) & (g92) & (!g468)) + ((g10) & (!sk[59]) & (g99) & (g109) & (g92) & (g468)) + ((g10) & (sk[59]) & (!g99) & (!g109) & (!g92) & (!g468)) + ((g10) & (sk[59]) & (!g99) & (!g109) & (!g92) & (g468)) + ((g10) & (sk[59]) & (!g99) & (!g109) & (g92) & (!g468)) + ((g10) & (sk[59]) & (!g99) & (!g109) & (g92) & (g468)) + ((g10) & (sk[59]) & (g99) & (!g109) & (g92) & (g468)));
	assign g1194 = (((!g101) & (!g224) & (!g467) & (!g574) & (!g1192) & (g1193)) + ((!g101) & (!g224) & (!g467) & (g574) & (!g1192) & (g1193)) + ((!g101) & (!g224) & (g467) & (!g574) & (!g1192) & (g1193)) + ((!g101) & (!g224) & (g467) & (g574) & (!g1192) & (g1193)) + ((!g101) & (g224) & (!g467) & (!g574) & (!g1192) & (g1193)) + ((!g101) & (g224) & (!g467) & (g574) & (!g1192) & (g1193)) + ((!g101) & (g224) & (g467) & (!g574) & (!g1192) & (g1193)) + ((!g101) & (g224) & (g467) & (g574) & (!g1192) & (g1193)) + ((g101) & (!g224) & (g467) & (!g574) & (!g1192) & (g1193)));
	assign g1195 = (((!g932) & (g978) & (!g1164) & (g1166) & (!g1191) & (g1194)));
	assign g1196 = (((!sk[62]) & (g1020) & (!g1021)) + ((!sk[62]) & (g1020) & (g1021)) + ((sk[62]) & (!g1020) & (g1021)));
	assign g1197 = (((!sk[63]) & (!g21) & (!g12) & (g134) & (g136)) + ((!sk[63]) & (!g21) & (g12) & (!g134) & (!g136)) + ((!sk[63]) & (!g21) & (g12) & (!g134) & (g136)) + ((!sk[63]) & (!g21) & (g12) & (g134) & (!g136)) + ((!sk[63]) & (!g21) & (g12) & (g134) & (g136)) + ((!sk[63]) & (g21) & (!g12) & (g134) & (!g136)) + ((!sk[63]) & (g21) & (!g12) & (g134) & (g136)) + ((!sk[63]) & (g21) & (g12) & (!g134) & (!g136)) + ((!sk[63]) & (g21) & (g12) & (!g134) & (g136)) + ((!sk[63]) & (g21) & (g12) & (g134) & (!g136)) + ((!sk[63]) & (g21) & (g12) & (g134) & (g136)) + ((sk[63]) & (!g21) & (!g12) & (!g134) & (!g136)) + ((sk[63]) & (!g21) & (!g12) & (!g134) & (g136)) + ((sk[63]) & (!g21) & (!g12) & (g134) & (!g136)) + ((sk[63]) & (!g21) & (!g12) & (g134) & (g136)) + ((sk[63]) & (!g21) & (g12) & (!g134) & (!g136)) + ((sk[63]) & (g21) & (!g12) & (!g134) & (!g136)) + ((sk[63]) & (g21) & (!g12) & (!g134) & (g136)) + ((sk[63]) & (g21) & (g12) & (!g134) & (!g136)));
	assign g1198 = (((!i_14_) & (!i_12_) & (!i_13_) & (g11) & (!g22) & (g136)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g11) & (g22) & (g136)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g11) & (g22) & (g136)) + ((!i_14_) & (!i_12_) & (i_13_) & (g11) & (g22) & (g136)) + ((!i_14_) & (i_12_) & (i_13_) & (g11) & (!g22) & (g136)) + ((!i_14_) & (i_12_) & (i_13_) & (g11) & (g22) & (g136)) + ((i_14_) & (i_12_) & (!i_13_) & (g11) & (!g22) & (g136)) + ((i_14_) & (i_12_) & (!i_13_) & (g11) & (g22) & (g136)) + ((i_14_) & (i_12_) & (i_13_) & (!g11) & (g22) & (g136)) + ((i_14_) & (i_12_) & (i_13_) & (g11) & (g22) & (g136)));
	assign g1199 = (((!i_14_) & (!sk[65]) & (!i_12_) & (!i_13_) & (!g11) & (g22)) + ((!i_14_) & (!sk[65]) & (!i_12_) & (!i_13_) & (g11) & (g22)) + ((!i_14_) & (!sk[65]) & (!i_12_) & (i_13_) & (!g11) & (g22)) + ((!i_14_) & (!sk[65]) & (!i_12_) & (i_13_) & (g11) & (g22)) + ((!i_14_) & (!sk[65]) & (i_12_) & (!i_13_) & (!g11) & (g22)) + ((!i_14_) & (!sk[65]) & (i_12_) & (!i_13_) & (g11) & (g22)) + ((!i_14_) & (!sk[65]) & (i_12_) & (i_13_) & (!g11) & (g22)) + ((!i_14_) & (!sk[65]) & (i_12_) & (i_13_) & (g11) & (g22)) + ((!i_14_) & (sk[65]) & (!i_12_) & (!i_13_) & (!g11) & (g22)) + ((!i_14_) & (sk[65]) & (!i_12_) & (!i_13_) & (g11) & (!g22)) + ((!i_14_) & (sk[65]) & (!i_12_) & (!i_13_) & (g11) & (g22)) + ((!i_14_) & (sk[65]) & (!i_12_) & (i_13_) & (!g11) & (g22)) + ((!i_14_) & (sk[65]) & (!i_12_) & (i_13_) & (g11) & (g22)) + ((!i_14_) & (sk[65]) & (i_12_) & (!i_13_) & (g11) & (!g22)) + ((!i_14_) & (sk[65]) & (i_12_) & (!i_13_) & (g11) & (g22)) + ((i_14_) & (!sk[65]) & (!i_12_) & (!i_13_) & (!g11) & (!g22)) + ((i_14_) & (!sk[65]) & (!i_12_) & (!i_13_) & (!g11) & (g22)) + ((i_14_) & (!sk[65]) & (!i_12_) & (!i_13_) & (g11) & (!g22)) + ((i_14_) & (!sk[65]) & (!i_12_) & (!i_13_) & (g11) & (g22)) + ((i_14_) & (!sk[65]) & (!i_12_) & (i_13_) & (!g11) & (!g22)) + ((i_14_) & (!sk[65]) & (!i_12_) & (i_13_) & (!g11) & (g22)) + ((i_14_) & (!sk[65]) & (!i_12_) & (i_13_) & (g11) & (!g22)) + ((i_14_) & (!sk[65]) & (!i_12_) & (i_13_) & (g11) & (g22)) + ((i_14_) & (!sk[65]) & (i_12_) & (!i_13_) & (!g11) & (!g22)) + ((i_14_) & (!sk[65]) & (i_12_) & (!i_13_) & (!g11) & (g22)) + ((i_14_) & (!sk[65]) & (i_12_) & (!i_13_) & (g11) & (!g22)) + ((i_14_) & (!sk[65]) & (i_12_) & (!i_13_) & (g11) & (g22)) + ((i_14_) & (!sk[65]) & (i_12_) & (i_13_) & (!g11) & (!g22)) + ((i_14_) & (!sk[65]) & (i_12_) & (i_13_) & (!g11) & (g22)) + ((i_14_) & (!sk[65]) & (i_12_) & (i_13_) & (g11) & (!g22)) + ((i_14_) & (!sk[65]) & (i_12_) & (i_13_) & (g11) & (g22)) + ((i_14_) & (sk[65]) & (i_12_) & (!i_13_) & (!g11) & (g22)) + ((i_14_) & (sk[65]) & (i_12_) & (!i_13_) & (g11) & (!g22)) + ((i_14_) & (sk[65]) & (i_12_) & (!i_13_) & (g11) & (g22)));
	assign g1200 = (((!sk[66]) & (!g112) & (!g201) & (!g530) & (!g703) & (g908)) + ((!sk[66]) & (!g112) & (!g201) & (!g530) & (g703) & (g908)) + ((!sk[66]) & (!g112) & (!g201) & (g530) & (!g703) & (g908)) + ((!sk[66]) & (!g112) & (!g201) & (g530) & (g703) & (g908)) + ((!sk[66]) & (!g112) & (g201) & (!g530) & (!g703) & (g908)) + ((!sk[66]) & (!g112) & (g201) & (!g530) & (g703) & (g908)) + ((!sk[66]) & (!g112) & (g201) & (g530) & (!g703) & (g908)) + ((!sk[66]) & (!g112) & (g201) & (g530) & (g703) & (g908)) + ((!sk[66]) & (g112) & (!g201) & (!g530) & (!g703) & (!g908)) + ((!sk[66]) & (g112) & (!g201) & (!g530) & (!g703) & (g908)) + ((!sk[66]) & (g112) & (!g201) & (!g530) & (g703) & (!g908)) + ((!sk[66]) & (g112) & (!g201) & (!g530) & (g703) & (g908)) + ((!sk[66]) & (g112) & (!g201) & (g530) & (!g703) & (!g908)) + ((!sk[66]) & (g112) & (!g201) & (g530) & (!g703) & (g908)) + ((!sk[66]) & (g112) & (!g201) & (g530) & (g703) & (!g908)) + ((!sk[66]) & (g112) & (!g201) & (g530) & (g703) & (g908)) + ((!sk[66]) & (g112) & (g201) & (!g530) & (!g703) & (!g908)) + ((!sk[66]) & (g112) & (g201) & (!g530) & (!g703) & (g908)) + ((!sk[66]) & (g112) & (g201) & (!g530) & (g703) & (!g908)) + ((!sk[66]) & (g112) & (g201) & (!g530) & (g703) & (g908)) + ((!sk[66]) & (g112) & (g201) & (g530) & (!g703) & (!g908)) + ((!sk[66]) & (g112) & (g201) & (g530) & (!g703) & (g908)) + ((!sk[66]) & (g112) & (g201) & (g530) & (g703) & (!g908)) + ((!sk[66]) & (g112) & (g201) & (g530) & (g703) & (g908)) + ((sk[66]) & (g112) & (!g201) & (!g530) & (!g703) & (!g908)) + ((sk[66]) & (g112) & (!g201) & (!g530) & (!g703) & (g908)) + ((sk[66]) & (g112) & (!g201) & (!g530) & (g703) & (!g908)) + ((sk[66]) & (g112) & (!g201) & (!g530) & (g703) & (g908)) + ((sk[66]) & (g112) & (!g201) & (g530) & (!g703) & (!g908)) + ((sk[66]) & (g112) & (!g201) & (g530) & (!g703) & (g908)) + ((sk[66]) & (g112) & (!g201) & (g530) & (g703) & (!g908)) + ((sk[66]) & (g112) & (!g201) & (g530) & (g703) & (g908)) + ((sk[66]) & (g112) & (g201) & (!g530) & (!g703) & (g908)) + ((sk[66]) & (g112) & (g201) & (!g530) & (g703) & (!g908)) + ((sk[66]) & (g112) & (g201) & (!g530) & (g703) & (g908)) + ((sk[66]) & (g112) & (g201) & (g530) & (!g703) & (!g908)) + ((sk[66]) & (g112) & (g201) & (g530) & (!g703) & (g908)) + ((sk[66]) & (g112) & (g201) & (g530) & (g703) & (!g908)) + ((sk[66]) & (g112) & (g201) & (g530) & (g703) & (g908)));
	assign g1201 = (((!sk[67]) & (g134) & (!g1199) & (!g1200)) + ((!sk[67]) & (g134) & (!g1199) & (g1200)) + ((!sk[67]) & (g134) & (g1199) & (!g1200)) + ((!sk[67]) & (g134) & (g1199) & (g1200)) + ((sk[67]) & (!g134) & (!g1199) & (!g1200)) + ((sk[67]) & (!g134) & (g1199) & (!g1200)) + ((sk[67]) & (g134) & (!g1199) & (!g1200)));
	assign g1202 = (((!g134) & (!g153) & (!g506) & (g1197) & (!g1198) & (g1201)) + ((!g134) & (!g153) & (g506) & (g1197) & (!g1198) & (g1201)) + ((g134) & (!g153) & (!g506) & (g1197) & (!g1198) & (g1201)));
	assign g1203 = (((!g21) & (!g109) & (!g114) & (!sk[69]) & (!g605) & (g908)) + ((!g21) & (!g109) & (!g114) & (!sk[69]) & (g605) & (g908)) + ((!g21) & (!g109) & (!g114) & (sk[69]) & (!g605) & (!g908)) + ((!g21) & (!g109) & (!g114) & (sk[69]) & (!g605) & (g908)) + ((!g21) & (!g109) & (g114) & (!sk[69]) & (!g605) & (g908)) + ((!g21) & (!g109) & (g114) & (!sk[69]) & (g605) & (g908)) + ((!g21) & (!g109) & (g114) & (sk[69]) & (!g605) & (!g908)) + ((!g21) & (!g109) & (g114) & (sk[69]) & (!g605) & (g908)) + ((!g21) & (g109) & (!g114) & (!sk[69]) & (!g605) & (g908)) + ((!g21) & (g109) & (!g114) & (!sk[69]) & (g605) & (g908)) + ((!g21) & (g109) & (!g114) & (sk[69]) & (!g605) & (!g908)) + ((!g21) & (g109) & (g114) & (!sk[69]) & (!g605) & (g908)) + ((!g21) & (g109) & (g114) & (!sk[69]) & (g605) & (g908)) + ((g21) & (!g109) & (!g114) & (!sk[69]) & (!g605) & (!g908)) + ((g21) & (!g109) & (!g114) & (!sk[69]) & (!g605) & (g908)) + ((g21) & (!g109) & (!g114) & (!sk[69]) & (g605) & (!g908)) + ((g21) & (!g109) & (!g114) & (!sk[69]) & (g605) & (g908)) + ((g21) & (!g109) & (!g114) & (sk[69]) & (!g605) & (!g908)) + ((g21) & (!g109) & (!g114) & (sk[69]) & (!g605) & (g908)) + ((g21) & (!g109) & (g114) & (!sk[69]) & (!g605) & (!g908)) + ((g21) & (!g109) & (g114) & (!sk[69]) & (!g605) & (g908)) + ((g21) & (!g109) & (g114) & (!sk[69]) & (g605) & (!g908)) + ((g21) & (!g109) & (g114) & (!sk[69]) & (g605) & (g908)) + ((g21) & (!g109) & (g114) & (sk[69]) & (!g605) & (!g908)) + ((g21) & (!g109) & (g114) & (sk[69]) & (!g605) & (g908)) + ((g21) & (g109) & (!g114) & (!sk[69]) & (!g605) & (!g908)) + ((g21) & (g109) & (!g114) & (!sk[69]) & (!g605) & (g908)) + ((g21) & (g109) & (!g114) & (!sk[69]) & (g605) & (!g908)) + ((g21) & (g109) & (!g114) & (!sk[69]) & (g605) & (g908)) + ((g21) & (g109) & (g114) & (!sk[69]) & (!g605) & (!g908)) + ((g21) & (g109) & (g114) & (!sk[69]) & (!g605) & (g908)) + ((g21) & (g109) & (g114) & (!sk[69]) & (g605) & (!g908)) + ((g21) & (g109) & (g114) & (!sk[69]) & (g605) & (g908)));
	assign g1204 = (((!i_8_) & (!g108) & (!sk[70]) & (g530) & (g703)) + ((!i_8_) & (g108) & (!sk[70]) & (!g530) & (!g703)) + ((!i_8_) & (g108) & (!sk[70]) & (!g530) & (g703)) + ((!i_8_) & (g108) & (!sk[70]) & (g530) & (!g703)) + ((!i_8_) & (g108) & (!sk[70]) & (g530) & (g703)) + ((!i_8_) & (g108) & (sk[70]) & (!g530) & (g703)) + ((!i_8_) & (g108) & (sk[70]) & (g530) & (g703)) + ((i_8_) & (!g108) & (!sk[70]) & (g530) & (!g703)) + ((i_8_) & (!g108) & (!sk[70]) & (g530) & (g703)) + ((i_8_) & (g108) & (!sk[70]) & (!g530) & (!g703)) + ((i_8_) & (g108) & (!sk[70]) & (!g530) & (g703)) + ((i_8_) & (g108) & (!sk[70]) & (g530) & (!g703)) + ((i_8_) & (g108) & (!sk[70]) & (g530) & (g703)) + ((i_8_) & (g108) & (sk[70]) & (g530) & (!g703)) + ((i_8_) & (g108) & (sk[70]) & (g530) & (g703)));
	assign g1205 = (((!i_8_) & (!g12) & (!g206) & (g108) & (!g226) & (!g506)) + ((!i_8_) & (!g12) & (!g206) & (g108) & (!g226) & (g506)) + ((!i_8_) & (!g12) & (!g206) & (g108) & (g226) & (g506)) + ((!i_8_) & (!g12) & (g206) & (g108) & (!g226) & (!g506)) + ((!i_8_) & (!g12) & (g206) & (g108) & (!g226) & (g506)) + ((!i_8_) & (!g12) & (g206) & (g108) & (g226) & (g506)) + ((!i_8_) & (g12) & (!g206) & (g108) & (!g226) & (!g506)) + ((!i_8_) & (g12) & (!g206) & (g108) & (!g226) & (g506)) + ((!i_8_) & (g12) & (!g206) & (g108) & (g226) & (g506)) + ((!i_8_) & (g12) & (g206) & (g108) & (!g226) & (!g506)) + ((!i_8_) & (g12) & (g206) & (g108) & (!g226) & (g506)) + ((!i_8_) & (g12) & (g206) & (g108) & (g226) & (g506)) + ((i_8_) & (!g12) & (!g206) & (g108) & (!g226) & (!g506)) + ((i_8_) & (!g12) & (!g206) & (g108) & (!g226) & (g506)) + ((i_8_) & (!g12) & (!g206) & (g108) & (g226) & (!g506)) + ((i_8_) & (!g12) & (!g206) & (g108) & (g226) & (g506)) + ((i_8_) & (!g12) & (g206) & (g108) & (!g226) & (!g506)) + ((i_8_) & (!g12) & (g206) & (g108) & (!g226) & (g506)) + ((i_8_) & (g12) & (!g206) & (g108) & (!g226) & (!g506)) + ((i_8_) & (g12) & (!g206) & (g108) & (!g226) & (g506)) + ((i_8_) & (g12) & (!g206) & (g108) & (g226) & (!g506)) + ((i_8_) & (g12) & (!g206) & (g108) & (g226) & (g506)) + ((i_8_) & (g12) & (g206) & (g108) & (!g226) & (!g506)) + ((i_8_) & (g12) & (g206) & (g108) & (!g226) & (g506)) + ((i_8_) & (g12) & (g206) & (g108) & (g226) & (!g506)) + ((i_8_) & (g12) & (g206) & (g108) & (g226) & (g506)));
	assign g1206 = (((!g1143) & (!sk[72]) & (!g1203) & (g1204) & (g1205)) + ((!g1143) & (!sk[72]) & (g1203) & (!g1204) & (!g1205)) + ((!g1143) & (!sk[72]) & (g1203) & (!g1204) & (g1205)) + ((!g1143) & (!sk[72]) & (g1203) & (g1204) & (!g1205)) + ((!g1143) & (!sk[72]) & (g1203) & (g1204) & (g1205)) + ((g1143) & (!sk[72]) & (!g1203) & (g1204) & (!g1205)) + ((g1143) & (!sk[72]) & (!g1203) & (g1204) & (g1205)) + ((g1143) & (!sk[72]) & (g1203) & (!g1204) & (!g1205)) + ((g1143) & (!sk[72]) & (g1203) & (!g1204) & (g1205)) + ((g1143) & (!sk[72]) & (g1203) & (g1204) & (!g1205)) + ((g1143) & (!sk[72]) & (g1203) & (g1204) & (g1205)) + ((g1143) & (sk[72]) & (g1203) & (!g1204) & (!g1205)));
	assign g1207 = (((!g562) & (!g804) & (!g1148) & (sk[73]) & (!g1149)) + ((!g562) & (!g804) & (g1148) & (!sk[73]) & (g1149)) + ((!g562) & (g804) & (!g1148) & (!sk[73]) & (!g1149)) + ((!g562) & (g804) & (!g1148) & (!sk[73]) & (g1149)) + ((!g562) & (g804) & (g1148) & (!sk[73]) & (!g1149)) + ((!g562) & (g804) & (g1148) & (!sk[73]) & (g1149)) + ((g562) & (!g804) & (g1148) & (!sk[73]) & (!g1149)) + ((g562) & (!g804) & (g1148) & (!sk[73]) & (g1149)) + ((g562) & (g804) & (!g1148) & (!sk[73]) & (!g1149)) + ((g562) & (g804) & (!g1148) & (!sk[73]) & (g1149)) + ((g562) & (g804) & (g1148) & (!sk[73]) & (!g1149)) + ((g562) & (g804) & (g1148) & (!sk[73]) & (g1149)));
	assign g1208 = (((!sk[74]) & (g136) & (!g177) & (!g1176)) + ((!sk[74]) & (g136) & (!g177) & (g1176)) + ((!sk[74]) & (g136) & (g177) & (!g1176)) + ((!sk[74]) & (g136) & (g177) & (g1176)) + ((sk[74]) & (!g136) & (!g177) & (!g1176)) + ((sk[74]) & (!g136) & (g177) & (!g1176)) + ((sk[74]) & (g136) & (!g177) & (!g1176)));
	assign g1209 = (((!i_8_) & (!i_6_) & (!i_7_) & (g87) & (!g424) & (g530)) + ((!i_8_) & (!i_6_) & (!i_7_) & (g87) & (g424) & (g530)) + ((!i_8_) & (i_6_) & (i_7_) & (g87) & (g424) & (!g530)) + ((!i_8_) & (i_6_) & (i_7_) & (g87) & (g424) & (g530)) + ((i_8_) & (!i_6_) & (!i_7_) & (g87) & (!g424) & (g530)) + ((i_8_) & (!i_6_) & (!i_7_) & (g87) & (g424) & (g530)));
	assign g1210 = (((!g151) & (!g201) & (!g423) & (!g703) & (!sk[76]) & (g1209)) + ((!g151) & (!g201) & (!g423) & (!g703) & (sk[76]) & (!g1209)) + ((!g151) & (!g201) & (!g423) & (g703) & (!sk[76]) & (g1209)) + ((!g151) & (!g201) & (!g423) & (g703) & (sk[76]) & (!g1209)) + ((!g151) & (!g201) & (g423) & (!g703) & (!sk[76]) & (g1209)) + ((!g151) & (!g201) & (g423) & (g703) & (!sk[76]) & (g1209)) + ((!g151) & (g201) & (!g423) & (!g703) & (!sk[76]) & (g1209)) + ((!g151) & (g201) & (!g423) & (!g703) & (sk[76]) & (!g1209)) + ((!g151) & (g201) & (!g423) & (g703) & (!sk[76]) & (g1209)) + ((!g151) & (g201) & (!g423) & (g703) & (sk[76]) & (!g1209)) + ((!g151) & (g201) & (g423) & (!g703) & (!sk[76]) & (g1209)) + ((!g151) & (g201) & (g423) & (!g703) & (sk[76]) & (!g1209)) + ((!g151) & (g201) & (g423) & (g703) & (!sk[76]) & (g1209)) + ((g151) & (!g201) & (!g423) & (!g703) & (!sk[76]) & (!g1209)) + ((g151) & (!g201) & (!g423) & (!g703) & (!sk[76]) & (g1209)) + ((g151) & (!g201) & (!g423) & (g703) & (!sk[76]) & (!g1209)) + ((g151) & (!g201) & (!g423) & (g703) & (!sk[76]) & (g1209)) + ((g151) & (!g201) & (g423) & (!g703) & (!sk[76]) & (!g1209)) + ((g151) & (!g201) & (g423) & (!g703) & (!sk[76]) & (g1209)) + ((g151) & (!g201) & (g423) & (g703) & (!sk[76]) & (!g1209)) + ((g151) & (!g201) & (g423) & (g703) & (!sk[76]) & (g1209)) + ((g151) & (g201) & (!g423) & (!g703) & (!sk[76]) & (!g1209)) + ((g151) & (g201) & (!g423) & (!g703) & (!sk[76]) & (g1209)) + ((g151) & (g201) & (!g423) & (!g703) & (sk[76]) & (!g1209)) + ((g151) & (g201) & (!g423) & (g703) & (!sk[76]) & (!g1209)) + ((g151) & (g201) & (!g423) & (g703) & (!sk[76]) & (g1209)) + ((g151) & (g201) & (g423) & (!g703) & (!sk[76]) & (!g1209)) + ((g151) & (g201) & (g423) & (!g703) & (!sk[76]) & (g1209)) + ((g151) & (g201) & (g423) & (!g703) & (sk[76]) & (!g1209)) + ((g151) & (g201) & (g423) & (g703) & (!sk[76]) & (!g1209)) + ((g151) & (g201) & (g423) & (g703) & (!sk[76]) & (g1209)));
	assign g1211 = (((!g134) & (!g89) & (!g118) & (!sk[77]) & (!g593) & (g1096)) + ((!g134) & (!g89) & (!g118) & (!sk[77]) & (g593) & (g1096)) + ((!g134) & (!g89) & (!g118) & (sk[77]) & (!g593) & (g1096)) + ((!g134) & (!g89) & (!g118) & (sk[77]) & (g593) & (g1096)) + ((!g134) & (!g89) & (g118) & (!sk[77]) & (!g593) & (g1096)) + ((!g134) & (!g89) & (g118) & (!sk[77]) & (g593) & (g1096)) + ((!g134) & (!g89) & (g118) & (sk[77]) & (g593) & (g1096)) + ((!g134) & (g89) & (!g118) & (!sk[77]) & (!g593) & (g1096)) + ((!g134) & (g89) & (!g118) & (!sk[77]) & (g593) & (g1096)) + ((!g134) & (g89) & (!g118) & (sk[77]) & (!g593) & (!g1096)) + ((!g134) & (g89) & (!g118) & (sk[77]) & (!g593) & (g1096)) + ((!g134) & (g89) & (!g118) & (sk[77]) & (g593) & (!g1096)) + ((!g134) & (g89) & (!g118) & (sk[77]) & (g593) & (g1096)) + ((!g134) & (g89) & (g118) & (!sk[77]) & (!g593) & (g1096)) + ((!g134) & (g89) & (g118) & (!sk[77]) & (g593) & (g1096)) + ((!g134) & (g89) & (g118) & (sk[77]) & (g593) & (g1096)) + ((g134) & (!g89) & (!g118) & (!sk[77]) & (!g593) & (!g1096)) + ((g134) & (!g89) & (!g118) & (!sk[77]) & (!g593) & (g1096)) + ((g134) & (!g89) & (!g118) & (!sk[77]) & (g593) & (!g1096)) + ((g134) & (!g89) & (!g118) & (!sk[77]) & (g593) & (g1096)) + ((g134) & (!g89) & (!g118) & (sk[77]) & (g593) & (g1096)) + ((g134) & (!g89) & (g118) & (!sk[77]) & (!g593) & (!g1096)) + ((g134) & (!g89) & (g118) & (!sk[77]) & (!g593) & (g1096)) + ((g134) & (!g89) & (g118) & (!sk[77]) & (g593) & (!g1096)) + ((g134) & (!g89) & (g118) & (!sk[77]) & (g593) & (g1096)) + ((g134) & (!g89) & (g118) & (sk[77]) & (g593) & (g1096)) + ((g134) & (g89) & (!g118) & (!sk[77]) & (!g593) & (!g1096)) + ((g134) & (g89) & (!g118) & (!sk[77]) & (!g593) & (g1096)) + ((g134) & (g89) & (!g118) & (!sk[77]) & (g593) & (!g1096)) + ((g134) & (g89) & (!g118) & (!sk[77]) & (g593) & (g1096)) + ((g134) & (g89) & (!g118) & (sk[77]) & (g593) & (!g1096)) + ((g134) & (g89) & (!g118) & (sk[77]) & (g593) & (g1096)) + ((g134) & (g89) & (g118) & (!sk[77]) & (!g593) & (!g1096)) + ((g134) & (g89) & (g118) & (!sk[77]) & (!g593) & (g1096)) + ((g134) & (g89) & (g118) & (!sk[77]) & (g593) & (!g1096)) + ((g134) & (g89) & (g118) & (!sk[77]) & (g593) & (g1096)) + ((g134) & (g89) & (g118) & (sk[77]) & (g593) & (g1096)));
	assign g1212 = (((g99) & (!sk[78]) & (!g201)) + ((g99) & (!sk[78]) & (g201)) + ((g99) & (sk[78]) & (!g201)));
	assign g1213 = (((g118) & (!sk[79]) & (!g506)) + ((g118) & (!sk[79]) & (g506)) + ((g118) & (sk[79]) & (g506)));
	assign g1214 = (((g134) & (!sk[80]) & (!g464)) + ((g134) & (!sk[80]) & (g464)) + ((g134) & (sk[80]) & (!g464)));
	assign g1215 = (((!i_8_) & (!g23) & (!g206) & (!sk[81]) & (!g135) & (g226)) + ((!i_8_) & (!g23) & (!g206) & (!sk[81]) & (g135) & (g226)) + ((!i_8_) & (!g23) & (g206) & (!sk[81]) & (!g135) & (g226)) + ((!i_8_) & (!g23) & (g206) & (!sk[81]) & (g135) & (g226)) + ((!i_8_) & (g23) & (!g206) & (!sk[81]) & (!g135) & (g226)) + ((!i_8_) & (g23) & (!g206) & (!sk[81]) & (g135) & (g226)) + ((!i_8_) & (g23) & (g206) & (!sk[81]) & (!g135) & (g226)) + ((!i_8_) & (g23) & (g206) & (!sk[81]) & (g135) & (g226)) + ((i_8_) & (!g23) & (!g206) & (!sk[81]) & (!g135) & (!g226)) + ((i_8_) & (!g23) & (!g206) & (!sk[81]) & (!g135) & (g226)) + ((i_8_) & (!g23) & (!g206) & (!sk[81]) & (g135) & (!g226)) + ((i_8_) & (!g23) & (!g206) & (!sk[81]) & (g135) & (g226)) + ((i_8_) & (!g23) & (!g206) & (sk[81]) & (g135) & (!g226)) + ((i_8_) & (!g23) & (!g206) & (sk[81]) & (g135) & (g226)) + ((i_8_) & (!g23) & (g206) & (!sk[81]) & (!g135) & (!g226)) + ((i_8_) & (!g23) & (g206) & (!sk[81]) & (!g135) & (g226)) + ((i_8_) & (!g23) & (g206) & (!sk[81]) & (g135) & (!g226)) + ((i_8_) & (!g23) & (g206) & (!sk[81]) & (g135) & (g226)) + ((i_8_) & (!g23) & (g206) & (sk[81]) & (g135) & (!g226)) + ((i_8_) & (g23) & (!g206) & (!sk[81]) & (!g135) & (!g226)) + ((i_8_) & (g23) & (!g206) & (!sk[81]) & (!g135) & (g226)) + ((i_8_) & (g23) & (!g206) & (!sk[81]) & (g135) & (!g226)) + ((i_8_) & (g23) & (!g206) & (!sk[81]) & (g135) & (g226)) + ((i_8_) & (g23) & (!g206) & (sk[81]) & (g135) & (!g226)) + ((i_8_) & (g23) & (!g206) & (sk[81]) & (g135) & (g226)) + ((i_8_) & (g23) & (g206) & (!sk[81]) & (!g135) & (!g226)) + ((i_8_) & (g23) & (g206) & (!sk[81]) & (!g135) & (g226)) + ((i_8_) & (g23) & (g206) & (!sk[81]) & (g135) & (!g226)) + ((i_8_) & (g23) & (g206) & (!sk[81]) & (g135) & (g226)) + ((i_8_) & (g23) & (g206) & (sk[81]) & (g135) & (!g226)) + ((i_8_) & (g23) & (g206) & (sk[81]) & (g135) & (g226)));
	assign g1216 = (((!g297) & (!g1212) & (!g238) & (!g1213) & (!g1214) & (!g1215)) + ((!g297) & (!g1212) & (g238) & (!g1213) & (!g1214) & (!g1215)) + ((g297) & (!g1212) & (!g238) & (!g1213) & (!g1214) & (!g1215)));
	assign g1217 = (((g1207) & (g1208) & (g1210) & (g1607) & (g1211) & (g1216)));
	assign g1218 = (((!i_14_) & (!i_12_) & (!i_13_) & (g11) & (!g22) & (g118)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g11) & (g22) & (g118)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g11) & (g22) & (g118)) + ((!i_14_) & (!i_12_) & (i_13_) & (g11) & (!g22) & (g118)) + ((!i_14_) & (!i_12_) & (i_13_) & (g11) & (g22) & (g118)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g11) & (g22) & (g118)) + ((!i_14_) & (i_12_) & (!i_13_) & (g11) & (g22) & (g118)) + ((i_14_) & (i_12_) & (!i_13_) & (!g11) & (g22) & (g118)) + ((i_14_) & (i_12_) & (!i_13_) & (g11) & (!g22) & (g118)) + ((i_14_) & (i_12_) & (!i_13_) & (g11) & (g22) & (g118)) + ((i_14_) & (i_12_) & (i_13_) & (!g11) & (g22) & (g118)) + ((i_14_) & (i_12_) & (i_13_) & (g11) & (g22) & (g118)));
	assign g1219 = (((!g23) & (!g206) & (!g118) & (!g260) & (!g464) & (!g1218)) + ((!g23) & (!g206) & (!g118) & (!g260) & (g464) & (!g1218)) + ((!g23) & (g206) & (!g118) & (!g260) & (!g464) & (!g1218)) + ((!g23) & (g206) & (!g118) & (!g260) & (g464) & (!g1218)) + ((!g23) & (g206) & (g118) & (!g260) & (g464) & (!g1218)) + ((g23) & (!g206) & (!g118) & (!g260) & (!g464) & (!g1218)) + ((g23) & (!g206) & (!g118) & (!g260) & (g464) & (!g1218)) + ((g23) & (g206) & (!g118) & (!g260) & (!g464) & (!g1218)) + ((g23) & (g206) & (!g118) & (!g260) & (g464) & (!g1218)));
	assign g1220 = (((!g1095) & (!sk[86]) & (!g1098) & (!g1100) & (!g1541) & (g1219)) + ((!g1095) & (!sk[86]) & (!g1098) & (!g1100) & (g1541) & (g1219)) + ((!g1095) & (!sk[86]) & (!g1098) & (g1100) & (!g1541) & (g1219)) + ((!g1095) & (!sk[86]) & (!g1098) & (g1100) & (g1541) & (g1219)) + ((!g1095) & (!sk[86]) & (g1098) & (!g1100) & (!g1541) & (g1219)) + ((!g1095) & (!sk[86]) & (g1098) & (!g1100) & (g1541) & (g1219)) + ((!g1095) & (!sk[86]) & (g1098) & (g1100) & (!g1541) & (g1219)) + ((!g1095) & (!sk[86]) & (g1098) & (g1100) & (g1541) & (g1219)) + ((!g1095) & (sk[86]) & (!g1098) & (!g1100) & (g1541) & (g1219)) + ((g1095) & (!sk[86]) & (!g1098) & (!g1100) & (!g1541) & (!g1219)) + ((g1095) & (!sk[86]) & (!g1098) & (!g1100) & (!g1541) & (g1219)) + ((g1095) & (!sk[86]) & (!g1098) & (!g1100) & (g1541) & (!g1219)) + ((g1095) & (!sk[86]) & (!g1098) & (!g1100) & (g1541) & (g1219)) + ((g1095) & (!sk[86]) & (!g1098) & (g1100) & (!g1541) & (!g1219)) + ((g1095) & (!sk[86]) & (!g1098) & (g1100) & (!g1541) & (g1219)) + ((g1095) & (!sk[86]) & (!g1098) & (g1100) & (g1541) & (!g1219)) + ((g1095) & (!sk[86]) & (!g1098) & (g1100) & (g1541) & (g1219)) + ((g1095) & (!sk[86]) & (g1098) & (!g1100) & (!g1541) & (!g1219)) + ((g1095) & (!sk[86]) & (g1098) & (!g1100) & (!g1541) & (g1219)) + ((g1095) & (!sk[86]) & (g1098) & (!g1100) & (g1541) & (!g1219)) + ((g1095) & (!sk[86]) & (g1098) & (!g1100) & (g1541) & (g1219)) + ((g1095) & (!sk[86]) & (g1098) & (g1100) & (!g1541) & (!g1219)) + ((g1095) & (!sk[86]) & (g1098) & (g1100) & (!g1541) & (g1219)) + ((g1095) & (!sk[86]) & (g1098) & (g1100) & (g1541) & (!g1219)) + ((g1095) & (!sk[86]) & (g1098) & (g1100) & (g1541) & (g1219)));
	assign g1221 = (((g1196) & (g1045) & (g1202) & (g1206) & (g1217) & (g1220)));
	assign g1222 = (((!sk[88]) & (i_8_) & (!g135) & (!g224)) + ((!sk[88]) & (i_8_) & (!g135) & (g224)) + ((!sk[88]) & (i_8_) & (g135) & (!g224)) + ((!sk[88]) & (i_8_) & (g135) & (g224)) + ((sk[88]) & (i_8_) & (g135) & (g224)));
	assign g1223 = (((!sk[89]) & (g10) & (!g134)) + ((!sk[89]) & (g10) & (g134)) + ((sk[89]) & (g10) & (g134)));
	assign g1224 = (((!sk[90]) & (g66) & (!g118)) + ((!sk[90]) & (g66) & (g118)) + ((sk[90]) & (g66) & (g118)));
	assign g1225 = (((!sk[91]) & (!i_8_) & (!g134) & (!g221) & (!g135) & (g127)) + ((!sk[91]) & (!i_8_) & (!g134) & (!g221) & (g135) & (g127)) + ((!sk[91]) & (!i_8_) & (!g134) & (g221) & (!g135) & (g127)) + ((!sk[91]) & (!i_8_) & (!g134) & (g221) & (g135) & (g127)) + ((!sk[91]) & (!i_8_) & (g134) & (!g221) & (!g135) & (g127)) + ((!sk[91]) & (!i_8_) & (g134) & (!g221) & (g135) & (g127)) + ((!sk[91]) & (!i_8_) & (g134) & (g221) & (!g135) & (g127)) + ((!sk[91]) & (!i_8_) & (g134) & (g221) & (g135) & (g127)) + ((!sk[91]) & (i_8_) & (!g134) & (!g221) & (!g135) & (!g127)) + ((!sk[91]) & (i_8_) & (!g134) & (!g221) & (!g135) & (g127)) + ((!sk[91]) & (i_8_) & (!g134) & (!g221) & (g135) & (!g127)) + ((!sk[91]) & (i_8_) & (!g134) & (!g221) & (g135) & (g127)) + ((!sk[91]) & (i_8_) & (!g134) & (g221) & (!g135) & (!g127)) + ((!sk[91]) & (i_8_) & (!g134) & (g221) & (!g135) & (g127)) + ((!sk[91]) & (i_8_) & (!g134) & (g221) & (g135) & (!g127)) + ((!sk[91]) & (i_8_) & (!g134) & (g221) & (g135) & (g127)) + ((!sk[91]) & (i_8_) & (g134) & (!g221) & (!g135) & (!g127)) + ((!sk[91]) & (i_8_) & (g134) & (!g221) & (!g135) & (g127)) + ((!sk[91]) & (i_8_) & (g134) & (!g221) & (g135) & (!g127)) + ((!sk[91]) & (i_8_) & (g134) & (!g221) & (g135) & (g127)) + ((!sk[91]) & (i_8_) & (g134) & (g221) & (!g135) & (!g127)) + ((!sk[91]) & (i_8_) & (g134) & (g221) & (!g135) & (g127)) + ((!sk[91]) & (i_8_) & (g134) & (g221) & (g135) & (!g127)) + ((!sk[91]) & (i_8_) & (g134) & (g221) & (g135) & (g127)) + ((sk[91]) & (!i_8_) & (g134) & (!g221) & (!g135) & (!g127)) + ((sk[91]) & (!i_8_) & (g134) & (!g221) & (!g135) & (g127)) + ((sk[91]) & (!i_8_) & (g134) & (!g221) & (g135) & (!g127)) + ((sk[91]) & (!i_8_) & (g134) & (!g221) & (g135) & (g127)) + ((sk[91]) & (i_8_) & (!g134) & (!g221) & (g135) & (!g127)) + ((sk[91]) & (i_8_) & (!g134) & (g221) & (g135) & (!g127)) + ((sk[91]) & (i_8_) & (g134) & (!g221) & (!g135) & (!g127)) + ((sk[91]) & (i_8_) & (g134) & (!g221) & (!g135) & (g127)) + ((sk[91]) & (i_8_) & (g134) & (!g221) & (g135) & (!g127)) + ((sk[91]) & (i_8_) & (g134) & (!g221) & (g135) & (g127)) + ((sk[91]) & (i_8_) & (g134) & (g221) & (g135) & (!g127)));
	assign g1226 = (((!i_8_) & (!sk[92]) & (!g134) & (!g135) & (!g90) & (g467)) + ((!i_8_) & (!sk[92]) & (!g134) & (!g135) & (g90) & (g467)) + ((!i_8_) & (!sk[92]) & (!g134) & (g135) & (!g90) & (g467)) + ((!i_8_) & (!sk[92]) & (!g134) & (g135) & (g90) & (g467)) + ((!i_8_) & (!sk[92]) & (g134) & (!g135) & (!g90) & (g467)) + ((!i_8_) & (!sk[92]) & (g134) & (!g135) & (g90) & (g467)) + ((!i_8_) & (!sk[92]) & (g134) & (g135) & (!g90) & (g467)) + ((!i_8_) & (!sk[92]) & (g134) & (g135) & (g90) & (g467)) + ((!i_8_) & (sk[92]) & (g134) & (!g135) & (!g90) & (!g467)) + ((!i_8_) & (sk[92]) & (g134) & (!g135) & (!g90) & (g467)) + ((!i_8_) & (sk[92]) & (g134) & (g135) & (!g90) & (!g467)) + ((!i_8_) & (sk[92]) & (g134) & (g135) & (!g90) & (g467)) + ((i_8_) & (!sk[92]) & (!g134) & (!g135) & (!g90) & (!g467)) + ((i_8_) & (!sk[92]) & (!g134) & (!g135) & (!g90) & (g467)) + ((i_8_) & (!sk[92]) & (!g134) & (!g135) & (g90) & (!g467)) + ((i_8_) & (!sk[92]) & (!g134) & (!g135) & (g90) & (g467)) + ((i_8_) & (!sk[92]) & (!g134) & (g135) & (!g90) & (!g467)) + ((i_8_) & (!sk[92]) & (!g134) & (g135) & (!g90) & (g467)) + ((i_8_) & (!sk[92]) & (!g134) & (g135) & (g90) & (!g467)) + ((i_8_) & (!sk[92]) & (!g134) & (g135) & (g90) & (g467)) + ((i_8_) & (!sk[92]) & (g134) & (!g135) & (!g90) & (!g467)) + ((i_8_) & (!sk[92]) & (g134) & (!g135) & (!g90) & (g467)) + ((i_8_) & (!sk[92]) & (g134) & (!g135) & (g90) & (!g467)) + ((i_8_) & (!sk[92]) & (g134) & (!g135) & (g90) & (g467)) + ((i_8_) & (!sk[92]) & (g134) & (g135) & (!g90) & (!g467)) + ((i_8_) & (!sk[92]) & (g134) & (g135) & (!g90) & (g467)) + ((i_8_) & (!sk[92]) & (g134) & (g135) & (g90) & (!g467)) + ((i_8_) & (!sk[92]) & (g134) & (g135) & (g90) & (g467)) + ((i_8_) & (sk[92]) & (!g134) & (g135) & (!g90) & (!g467)) + ((i_8_) & (sk[92]) & (!g134) & (g135) & (!g90) & (g467)) + ((i_8_) & (sk[92]) & (!g134) & (g135) & (g90) & (!g467)) + ((i_8_) & (sk[92]) & (g134) & (!g135) & (!g90) & (!g467)) + ((i_8_) & (sk[92]) & (g134) & (!g135) & (!g90) & (g467)) + ((i_8_) & (sk[92]) & (g134) & (g135) & (!g90) & (!g467)) + ((i_8_) & (sk[92]) & (g134) & (g135) & (!g90) & (g467)) + ((i_8_) & (sk[92]) & (g134) & (g135) & (g90) & (!g467)));
	assign g1227 = (((!g370) & (!g1222) & (!g1223) & (!g1224) & (!g1225) & (!g1226)));
	assign g1228 = (((!g8) & (!i_8_) & (g135) & (!g528) & (!g817) & (!g1001)) + ((!g8) & (!i_8_) & (g135) & (!g528) & (!g817) & (g1001)) + ((!g8) & (!i_8_) & (g135) & (!g528) & (g817) & (!g1001)) + ((!g8) & (!i_8_) & (g135) & (!g528) & (g817) & (g1001)) + ((!g8) & (!i_8_) & (g135) & (g528) & (!g817) & (!g1001)) + ((!g8) & (!i_8_) & (g135) & (g528) & (!g817) & (g1001)) + ((!g8) & (!i_8_) & (g135) & (g528) & (g817) & (!g1001)) + ((!g8) & (!i_8_) & (g135) & (g528) & (g817) & (g1001)) + ((!g8) & (i_8_) & (g135) & (!g528) & (!g817) & (!g1001)) + ((!g8) & (i_8_) & (g135) & (!g528) & (!g817) & (g1001)) + ((!g8) & (i_8_) & (g135) & (!g528) & (g817) & (!g1001)) + ((!g8) & (i_8_) & (g135) & (!g528) & (g817) & (g1001)) + ((!g8) & (i_8_) & (g135) & (g528) & (g817) & (!g1001)) + ((!g8) & (i_8_) & (g135) & (g528) & (g817) & (g1001)) + ((g8) & (!i_8_) & (g135) & (!g528) & (!g817) & (!g1001)) + ((g8) & (!i_8_) & (g135) & (!g528) & (!g817) & (g1001)) + ((g8) & (!i_8_) & (g135) & (!g528) & (g817) & (!g1001)) + ((g8) & (!i_8_) & (g135) & (!g528) & (g817) & (g1001)) + ((g8) & (!i_8_) & (g135) & (g528) & (!g817) & (!g1001)) + ((g8) & (!i_8_) & (g135) & (g528) & (g817) & (!g1001)) + ((g8) & (i_8_) & (g135) & (!g528) & (!g817) & (!g1001)) + ((g8) & (i_8_) & (g135) & (!g528) & (!g817) & (g1001)) + ((g8) & (i_8_) & (g135) & (!g528) & (g817) & (!g1001)) + ((g8) & (i_8_) & (g135) & (!g528) & (g817) & (g1001)) + ((g8) & (i_8_) & (g135) & (g528) & (g817) & (!g1001)) + ((g8) & (i_8_) & (g135) & (g528) & (g817) & (g1001)));
	assign g1229 = (((!g608) & (!g1174) & (!g1175) & (g1177) & (g1227) & (!g1228)));
	assign g1230 = (((!g145) & (!g187) & (!sk[96]) & (!g534) & (!g702) & (g881)) + ((!g145) & (!g187) & (!sk[96]) & (!g534) & (g702) & (g881)) + ((!g145) & (!g187) & (!sk[96]) & (g534) & (!g702) & (g881)) + ((!g145) & (!g187) & (!sk[96]) & (g534) & (g702) & (g881)) + ((!g145) & (g187) & (!sk[96]) & (!g534) & (!g702) & (g881)) + ((!g145) & (g187) & (!sk[96]) & (!g534) & (g702) & (g881)) + ((!g145) & (g187) & (!sk[96]) & (g534) & (!g702) & (g881)) + ((!g145) & (g187) & (!sk[96]) & (g534) & (g702) & (g881)) + ((g145) & (!g187) & (!sk[96]) & (!g534) & (!g702) & (!g881)) + ((g145) & (!g187) & (!sk[96]) & (!g534) & (!g702) & (g881)) + ((g145) & (!g187) & (!sk[96]) & (!g534) & (g702) & (!g881)) + ((g145) & (!g187) & (!sk[96]) & (!g534) & (g702) & (g881)) + ((g145) & (!g187) & (!sk[96]) & (g534) & (!g702) & (!g881)) + ((g145) & (!g187) & (!sk[96]) & (g534) & (!g702) & (g881)) + ((g145) & (!g187) & (!sk[96]) & (g534) & (g702) & (!g881)) + ((g145) & (!g187) & (!sk[96]) & (g534) & (g702) & (g881)) + ((g145) & (!g187) & (sk[96]) & (!g534) & (!g702) & (g881)) + ((g145) & (!g187) & (sk[96]) & (!g534) & (g702) & (!g881)) + ((g145) & (!g187) & (sk[96]) & (!g534) & (g702) & (g881)) + ((g145) & (!g187) & (sk[96]) & (g534) & (!g702) & (!g881)) + ((g145) & (!g187) & (sk[96]) & (g534) & (!g702) & (g881)) + ((g145) & (!g187) & (sk[96]) & (g534) & (g702) & (!g881)) + ((g145) & (!g187) & (sk[96]) & (g534) & (g702) & (g881)) + ((g145) & (g187) & (!sk[96]) & (!g534) & (!g702) & (!g881)) + ((g145) & (g187) & (!sk[96]) & (!g534) & (!g702) & (g881)) + ((g145) & (g187) & (!sk[96]) & (!g534) & (g702) & (!g881)) + ((g145) & (g187) & (!sk[96]) & (!g534) & (g702) & (g881)) + ((g145) & (g187) & (!sk[96]) & (g534) & (!g702) & (!g881)) + ((g145) & (g187) & (!sk[96]) & (g534) & (!g702) & (g881)) + ((g145) & (g187) & (!sk[96]) & (g534) & (g702) & (!g881)) + ((g145) & (g187) & (!sk[96]) & (g534) & (g702) & (g881)) + ((g145) & (g187) & (sk[96]) & (!g534) & (!g702) & (!g881)) + ((g145) & (g187) & (sk[96]) & (!g534) & (!g702) & (g881)) + ((g145) & (g187) & (sk[96]) & (!g534) & (g702) & (!g881)) + ((g145) & (g187) & (sk[96]) & (!g534) & (g702) & (g881)) + ((g145) & (g187) & (sk[96]) & (g534) & (!g702) & (!g881)) + ((g145) & (g187) & (sk[96]) & (g534) & (!g702) & (g881)) + ((g145) & (g187) & (sk[96]) & (g534) & (g702) & (!g881)) + ((g145) & (g187) & (sk[96]) & (g534) & (g702) & (g881)));
	assign g1231 = (((g6) & (!i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g109)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g109)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (i_13_) & (g109)) + ((g6) & (i_15_) & (!i_14_) & (!i_12_) & (!i_13_) & (g109)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g109)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (i_13_) & (g109)) + ((g6) & (i_15_) & (i_14_) & (i_12_) & (!i_13_) & (g109)));
	assign g1232 = (((!i_8_) & (!g46) & (!g209) & (!sk[98]) & (!g531) & (g1060)) + ((!i_8_) & (!g46) & (!g209) & (!sk[98]) & (g531) & (g1060)) + ((!i_8_) & (!g46) & (!g209) & (sk[98]) & (!g531) & (!g1060)) + ((!i_8_) & (!g46) & (!g209) & (sk[98]) & (g531) & (!g1060)) + ((!i_8_) & (!g46) & (g209) & (!sk[98]) & (!g531) & (g1060)) + ((!i_8_) & (!g46) & (g209) & (!sk[98]) & (g531) & (g1060)) + ((!i_8_) & (!g46) & (g209) & (sk[98]) & (!g531) & (!g1060)) + ((!i_8_) & (!g46) & (g209) & (sk[98]) & (g531) & (!g1060)) + ((!i_8_) & (g46) & (!g209) & (!sk[98]) & (!g531) & (g1060)) + ((!i_8_) & (g46) & (!g209) & (!sk[98]) & (g531) & (g1060)) + ((!i_8_) & (g46) & (g209) & (!sk[98]) & (!g531) & (g1060)) + ((!i_8_) & (g46) & (g209) & (!sk[98]) & (g531) & (g1060)) + ((i_8_) & (!g46) & (!g209) & (!sk[98]) & (!g531) & (!g1060)) + ((i_8_) & (!g46) & (!g209) & (!sk[98]) & (!g531) & (g1060)) + ((i_8_) & (!g46) & (!g209) & (!sk[98]) & (g531) & (!g1060)) + ((i_8_) & (!g46) & (!g209) & (!sk[98]) & (g531) & (g1060)) + ((i_8_) & (!g46) & (!g209) & (sk[98]) & (!g531) & (!g1060)) + ((i_8_) & (!g46) & (!g209) & (sk[98]) & (!g531) & (g1060)) + ((i_8_) & (!g46) & (g209) & (!sk[98]) & (!g531) & (!g1060)) + ((i_8_) & (!g46) & (g209) & (!sk[98]) & (!g531) & (g1060)) + ((i_8_) & (!g46) & (g209) & (!sk[98]) & (g531) & (!g1060)) + ((i_8_) & (!g46) & (g209) & (!sk[98]) & (g531) & (g1060)) + ((i_8_) & (g46) & (!g209) & (!sk[98]) & (!g531) & (!g1060)) + ((i_8_) & (g46) & (!g209) & (!sk[98]) & (!g531) & (g1060)) + ((i_8_) & (g46) & (!g209) & (!sk[98]) & (g531) & (!g1060)) + ((i_8_) & (g46) & (!g209) & (!sk[98]) & (g531) & (g1060)) + ((i_8_) & (g46) & (!g209) & (sk[98]) & (!g531) & (!g1060)) + ((i_8_) & (g46) & (!g209) & (sk[98]) & (!g531) & (g1060)) + ((i_8_) & (g46) & (g209) & (!sk[98]) & (!g531) & (!g1060)) + ((i_8_) & (g46) & (g209) & (!sk[98]) & (!g531) & (g1060)) + ((i_8_) & (g46) & (g209) & (!sk[98]) & (g531) & (!g1060)) + ((i_8_) & (g46) & (g209) & (!sk[98]) & (g531) & (g1060)));
	assign g1233 = (((!i_8_) & (!g206) & (!g108) & (!sk[99]) & (!g127) & (g561)) + ((!i_8_) & (!g206) & (!g108) & (!sk[99]) & (g127) & (g561)) + ((!i_8_) & (!g206) & (g108) & (!sk[99]) & (!g127) & (g561)) + ((!i_8_) & (!g206) & (g108) & (!sk[99]) & (g127) & (g561)) + ((!i_8_) & (!g206) & (g108) & (sk[99]) & (!g127) & (!g561)) + ((!i_8_) & (!g206) & (g108) & (sk[99]) & (!g127) & (g561)) + ((!i_8_) & (!g206) & (g108) & (sk[99]) & (g127) & (!g561)) + ((!i_8_) & (!g206) & (g108) & (sk[99]) & (g127) & (g561)) + ((!i_8_) & (g206) & (!g108) & (!sk[99]) & (!g127) & (g561)) + ((!i_8_) & (g206) & (!g108) & (!sk[99]) & (g127) & (g561)) + ((!i_8_) & (g206) & (g108) & (!sk[99]) & (!g127) & (g561)) + ((!i_8_) & (g206) & (g108) & (!sk[99]) & (g127) & (g561)) + ((!i_8_) & (g206) & (g108) & (sk[99]) & (!g127) & (!g561)) + ((!i_8_) & (g206) & (g108) & (sk[99]) & (!g127) & (g561)) + ((!i_8_) & (g206) & (g108) & (sk[99]) & (g127) & (g561)) + ((i_8_) & (!g206) & (!g108) & (!sk[99]) & (!g127) & (!g561)) + ((i_8_) & (!g206) & (!g108) & (!sk[99]) & (!g127) & (g561)) + ((i_8_) & (!g206) & (!g108) & (!sk[99]) & (g127) & (!g561)) + ((i_8_) & (!g206) & (!g108) & (!sk[99]) & (g127) & (g561)) + ((i_8_) & (!g206) & (g108) & (!sk[99]) & (!g127) & (!g561)) + ((i_8_) & (!g206) & (g108) & (!sk[99]) & (!g127) & (g561)) + ((i_8_) & (!g206) & (g108) & (!sk[99]) & (g127) & (!g561)) + ((i_8_) & (!g206) & (g108) & (!sk[99]) & (g127) & (g561)) + ((i_8_) & (g206) & (!g108) & (!sk[99]) & (!g127) & (!g561)) + ((i_8_) & (g206) & (!g108) & (!sk[99]) & (!g127) & (g561)) + ((i_8_) & (g206) & (!g108) & (!sk[99]) & (g127) & (!g561)) + ((i_8_) & (g206) & (!g108) & (!sk[99]) & (g127) & (g561)) + ((i_8_) & (g206) & (g108) & (!sk[99]) & (!g127) & (!g561)) + ((i_8_) & (g206) & (g108) & (!sk[99]) & (!g127) & (g561)) + ((i_8_) & (g206) & (g108) & (!sk[99]) & (g127) & (!g561)) + ((i_8_) & (g206) & (g108) & (!sk[99]) & (g127) & (g561)));
	assign g1234 = (((!i_8_) & (!g23) & (!g12) & (!g108) & (!g1232) & (!g1233)) + ((!i_8_) & (!g23) & (!g12) & (!g108) & (g1232) & (!g1233)) + ((!i_8_) & (!g23) & (!g12) & (g108) & (g1232) & (!g1233)) + ((!i_8_) & (!g23) & (g12) & (!g108) & (!g1232) & (!g1233)) + ((!i_8_) & (!g23) & (g12) & (!g108) & (g1232) & (!g1233)) + ((!i_8_) & (g23) & (!g12) & (!g108) & (!g1232) & (!g1233)) + ((!i_8_) & (g23) & (!g12) & (!g108) & (g1232) & (!g1233)) + ((!i_8_) & (g23) & (g12) & (!g108) & (!g1232) & (!g1233)) + ((!i_8_) & (g23) & (g12) & (!g108) & (g1232) & (!g1233)) + ((i_8_) & (!g23) & (!g12) & (!g108) & (!g1232) & (!g1233)) + ((i_8_) & (!g23) & (!g12) & (!g108) & (g1232) & (!g1233)) + ((i_8_) & (!g23) & (!g12) & (g108) & (g1232) & (!g1233)) + ((i_8_) & (!g23) & (g12) & (!g108) & (!g1232) & (!g1233)) + ((i_8_) & (!g23) & (g12) & (!g108) & (g1232) & (!g1233)) + ((i_8_) & (!g23) & (g12) & (g108) & (g1232) & (!g1233)) + ((i_8_) & (g23) & (!g12) & (!g108) & (!g1232) & (!g1233)) + ((i_8_) & (g23) & (!g12) & (!g108) & (g1232) & (!g1233)) + ((i_8_) & (g23) & (!g12) & (g108) & (g1232) & (!g1233)) + ((i_8_) & (g23) & (g12) & (!g108) & (!g1232) & (!g1233)) + ((i_8_) & (g23) & (g12) & (!g108) & (g1232) & (!g1233)) + ((i_8_) & (g23) & (g12) & (g108) & (g1232) & (!g1233)));
	assign g1235 = (((g1628) & (g1622) & (g1104) & (!g1230) & (!g1231) & (g1234)));
	assign g1236 = (((g6) & (!i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g112)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g112)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (i_13_) & (g112)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (!i_13_) & (g112)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (i_13_) & (g112)) + ((g6) & (i_15_) & (!i_14_) & (!i_12_) & (i_13_) & (g112)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g112)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (i_13_) & (g112)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g112)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (i_13_) & (g112)) + ((g6) & (i_15_) & (i_14_) & (i_12_) & (!i_13_) & (g112)) + ((g6) & (i_15_) & (i_14_) & (i_12_) & (i_13_) & (g112)));
	assign g1237 = (((g6) & (!i_15_) & (!i_14_) & (!i_12_) & (i_13_) & (g118)) + ((g6) & (!i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g118)) + ((g6) & (!i_15_) & (!i_14_) & (i_12_) & (i_13_) & (g118)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g118)) + ((g6) & (!i_15_) & (i_14_) & (!i_12_) & (i_13_) & (g118)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (!i_13_) & (g118)) + ((g6) & (!i_15_) & (i_14_) & (i_12_) & (i_13_) & (g118)) + ((g6) & (i_15_) & (!i_14_) & (!i_12_) & (!i_13_) & (g118)) + ((g6) & (i_15_) & (!i_14_) & (!i_12_) & (i_13_) & (g118)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (!i_13_) & (g118)) + ((g6) & (i_15_) & (!i_14_) & (i_12_) & (i_13_) & (g118)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (!i_13_) & (g118)) + ((g6) & (i_15_) & (i_14_) & (!i_12_) & (i_13_) & (g118)) + ((g6) & (i_15_) & (i_14_) & (i_12_) & (!i_13_) & (g118)));
	assign g1238 = (((!sk[104]) & (g1236) & (!g1237)) + ((!sk[104]) & (g1236) & (g1237)) + ((sk[104]) & (!g1236) & (!g1237)));
	assign g1239 = (((!g109) & (!g529) & (!sk[105]) & (!g1721) & (!g537) & (g1238)) + ((!g109) & (!g529) & (!sk[105]) & (!g1721) & (g537) & (g1238)) + ((!g109) & (!g529) & (!sk[105]) & (g1721) & (!g537) & (g1238)) + ((!g109) & (!g529) & (!sk[105]) & (g1721) & (g537) & (g1238)) + ((!g109) & (!g529) & (sk[105]) & (g1721) & (g537) & (g1238)) + ((!g109) & (g529) & (!sk[105]) & (!g1721) & (!g537) & (g1238)) + ((!g109) & (g529) & (!sk[105]) & (!g1721) & (g537) & (g1238)) + ((!g109) & (g529) & (!sk[105]) & (g1721) & (!g537) & (g1238)) + ((!g109) & (g529) & (!sk[105]) & (g1721) & (g537) & (g1238)) + ((!g109) & (g529) & (sk[105]) & (g1721) & (g537) & (g1238)) + ((g109) & (!g529) & (!sk[105]) & (!g1721) & (!g537) & (!g1238)) + ((g109) & (!g529) & (!sk[105]) & (!g1721) & (!g537) & (g1238)) + ((g109) & (!g529) & (!sk[105]) & (!g1721) & (g537) & (!g1238)) + ((g109) & (!g529) & (!sk[105]) & (!g1721) & (g537) & (g1238)) + ((g109) & (!g529) & (!sk[105]) & (g1721) & (!g537) & (!g1238)) + ((g109) & (!g529) & (!sk[105]) & (g1721) & (!g537) & (g1238)) + ((g109) & (!g529) & (!sk[105]) & (g1721) & (g537) & (!g1238)) + ((g109) & (!g529) & (!sk[105]) & (g1721) & (g537) & (g1238)) + ((g109) & (g529) & (!sk[105]) & (!g1721) & (!g537) & (!g1238)) + ((g109) & (g529) & (!sk[105]) & (!g1721) & (!g537) & (g1238)) + ((g109) & (g529) & (!sk[105]) & (!g1721) & (g537) & (!g1238)) + ((g109) & (g529) & (!sk[105]) & (!g1721) & (g537) & (g1238)) + ((g109) & (g529) & (!sk[105]) & (g1721) & (!g537) & (!g1238)) + ((g109) & (g529) & (!sk[105]) & (g1721) & (!g537) & (g1238)) + ((g109) & (g529) & (!sk[105]) & (g1721) & (g537) & (!g1238)) + ((g109) & (g529) & (!sk[105]) & (g1721) & (g537) & (g1238)) + ((g109) & (g529) & (sk[105]) & (g1721) & (g537) & (g1238)));
	assign g1240 = (((!sk[106]) & (g46) & (!g243)) + ((!sk[106]) & (g46) & (g243)) + ((sk[106]) & (g46) & (g243)));
	assign g1241 = (((!g185) & (!g151) & (!g187) & (!g429) & (!g1033) & (!g1240)) + ((!g185) & (!g151) & (!g187) & (g429) & (!g1033) & (!g1240)) + ((!g185) & (!g151) & (g187) & (!g429) & (!g1033) & (!g1240)) + ((g185) & (!g151) & (!g187) & (!g429) & (!g1033) & (!g1240)) + ((g185) & (!g151) & (!g187) & (g429) & (!g1033) & (!g1240)) + ((g185) & (!g151) & (g187) & (!g429) & (!g1033) & (!g1240)) + ((g185) & (g151) & (!g187) & (!g429) & (!g1033) & (!g1240)) + ((g185) & (g151) & (!g187) & (g429) & (!g1033) & (!g1240)) + ((g185) & (g151) & (g187) & (!g429) & (!g1033) & (!g1240)));
	assign g1242 = (((!g8) & (!g197) & (g90) & (!sk[108]) & (g424)) + ((!g8) & (g197) & (!g90) & (!sk[108]) & (!g424)) + ((!g8) & (g197) & (!g90) & (!sk[108]) & (g424)) + ((!g8) & (g197) & (g90) & (!sk[108]) & (!g424)) + ((!g8) & (g197) & (g90) & (!sk[108]) & (g424)) + ((g8) & (!g197) & (g90) & (!sk[108]) & (!g424)) + ((g8) & (!g197) & (g90) & (!sk[108]) & (g424)) + ((g8) & (!g197) & (g90) & (sk[108]) & (!g424)) + ((g8) & (g197) & (!g90) & (!sk[108]) & (!g424)) + ((g8) & (g197) & (!g90) & (!sk[108]) & (g424)) + ((g8) & (g197) & (g90) & (!sk[108]) & (!g424)) + ((g8) & (g197) & (g90) & (!sk[108]) & (g424)));
	assign g1243 = (((!i_8_) & (!g108) & (g185) & (!sk[109]) & (g231)) + ((!i_8_) & (g108) & (!g185) & (!sk[109]) & (!g231)) + ((!i_8_) & (g108) & (!g185) & (!sk[109]) & (g231)) + ((!i_8_) & (g108) & (g185) & (!sk[109]) & (!g231)) + ((!i_8_) & (g108) & (g185) & (!sk[109]) & (g231)) + ((i_8_) & (!g108) & (g185) & (!sk[109]) & (!g231)) + ((i_8_) & (!g108) & (g185) & (!sk[109]) & (g231)) + ((i_8_) & (g108) & (!g185) & (!sk[109]) & (!g231)) + ((i_8_) & (g108) & (!g185) & (!sk[109]) & (g231)) + ((i_8_) & (g108) & (!g185) & (sk[109]) & (!g231)) + ((i_8_) & (g108) & (!g185) & (sk[109]) & (g231)) + ((i_8_) & (g108) & (g185) & (!sk[109]) & (!g231)) + ((i_8_) & (g108) & (g185) & (!sk[109]) & (g231)) + ((i_8_) & (g108) & (g185) & (sk[109]) & (!g231)));
	assign g1244 = (((!sk[110]) & (!g66) & (!g330) & (!g423) & (!g1242) & (g1243)) + ((!sk[110]) & (!g66) & (!g330) & (!g423) & (g1242) & (g1243)) + ((!sk[110]) & (!g66) & (!g330) & (g423) & (!g1242) & (g1243)) + ((!sk[110]) & (!g66) & (!g330) & (g423) & (g1242) & (g1243)) + ((!sk[110]) & (!g66) & (g330) & (!g423) & (!g1242) & (g1243)) + ((!sk[110]) & (!g66) & (g330) & (!g423) & (g1242) & (g1243)) + ((!sk[110]) & (!g66) & (g330) & (g423) & (!g1242) & (g1243)) + ((!sk[110]) & (!g66) & (g330) & (g423) & (g1242) & (g1243)) + ((!sk[110]) & (g66) & (!g330) & (!g423) & (!g1242) & (!g1243)) + ((!sk[110]) & (g66) & (!g330) & (!g423) & (!g1242) & (g1243)) + ((!sk[110]) & (g66) & (!g330) & (!g423) & (g1242) & (!g1243)) + ((!sk[110]) & (g66) & (!g330) & (!g423) & (g1242) & (g1243)) + ((!sk[110]) & (g66) & (!g330) & (g423) & (!g1242) & (!g1243)) + ((!sk[110]) & (g66) & (!g330) & (g423) & (!g1242) & (g1243)) + ((!sk[110]) & (g66) & (!g330) & (g423) & (g1242) & (!g1243)) + ((!sk[110]) & (g66) & (!g330) & (g423) & (g1242) & (g1243)) + ((!sk[110]) & (g66) & (g330) & (!g423) & (!g1242) & (!g1243)) + ((!sk[110]) & (g66) & (g330) & (!g423) & (!g1242) & (g1243)) + ((!sk[110]) & (g66) & (g330) & (!g423) & (g1242) & (!g1243)) + ((!sk[110]) & (g66) & (g330) & (!g423) & (g1242) & (g1243)) + ((!sk[110]) & (g66) & (g330) & (g423) & (!g1242) & (!g1243)) + ((!sk[110]) & (g66) & (g330) & (g423) & (!g1242) & (g1243)) + ((!sk[110]) & (g66) & (g330) & (g423) & (g1242) & (!g1243)) + ((!sk[110]) & (g66) & (g330) & (g423) & (g1242) & (g1243)) + ((sk[110]) & (!g66) & (!g330) & (!g423) & (!g1242) & (!g1243)) + ((sk[110]) & (!g66) & (!g330) & (!g423) & (g1242) & (!g1243)) + ((sk[110]) & (!g66) & (!g330) & (g423) & (g1242) & (!g1243)) + ((sk[110]) & (!g66) & (g330) & (!g423) & (!g1242) & (!g1243)) + ((sk[110]) & (!g66) & (g330) & (!g423) & (g1242) & (!g1243)) + ((sk[110]) & (!g66) & (g330) & (g423) & (g1242) & (!g1243)) + ((sk[110]) & (g66) & (g330) & (!g423) & (!g1242) & (!g1243)) + ((sk[110]) & (g66) & (g330) & (!g423) & (g1242) & (!g1243)) + ((sk[110]) & (g66) & (g330) & (g423) & (g1242) & (!g1243)));
	assign g1245 = (((!i_8_) & (!sk[111]) & (!g88) & (g108) & (g531)) + ((!i_8_) & (!sk[111]) & (g88) & (!g108) & (!g531)) + ((!i_8_) & (!sk[111]) & (g88) & (!g108) & (g531)) + ((!i_8_) & (!sk[111]) & (g88) & (g108) & (!g531)) + ((!i_8_) & (!sk[111]) & (g88) & (g108) & (g531)) + ((!i_8_) & (sk[111]) & (!g88) & (g108) & (g531)) + ((!i_8_) & (sk[111]) & (g88) & (g108) & (g531)) + ((i_8_) & (!sk[111]) & (!g88) & (g108) & (!g531)) + ((i_8_) & (!sk[111]) & (!g88) & (g108) & (g531)) + ((i_8_) & (!sk[111]) & (g88) & (!g108) & (!g531)) + ((i_8_) & (!sk[111]) & (g88) & (!g108) & (g531)) + ((i_8_) & (!sk[111]) & (g88) & (g108) & (!g531)) + ((i_8_) & (!sk[111]) & (g88) & (g108) & (g531)) + ((i_8_) & (sk[111]) & (g88) & (!g108) & (g531)) + ((i_8_) & (sk[111]) & (g88) & (g108) & (g531)));
	assign g1246 = (((!g227) & (!g209) & (!sk[112]) & (g746) & (g349)) + ((!g227) & (g209) & (!sk[112]) & (!g746) & (!g349)) + ((!g227) & (g209) & (!sk[112]) & (!g746) & (g349)) + ((!g227) & (g209) & (!sk[112]) & (g746) & (!g349)) + ((!g227) & (g209) & (!sk[112]) & (g746) & (g349)) + ((!g227) & (g209) & (sk[112]) & (g746) & (!g349)) + ((!g227) & (g209) & (sk[112]) & (g746) & (g349)) + ((g227) & (!g209) & (!sk[112]) & (g746) & (!g349)) + ((g227) & (!g209) & (!sk[112]) & (g746) & (g349)) + ((g227) & (!g209) & (sk[112]) & (!g746) & (g349)) + ((g227) & (!g209) & (sk[112]) & (g746) & (g349)) + ((g227) & (g209) & (!sk[112]) & (!g746) & (!g349)) + ((g227) & (g209) & (!sk[112]) & (!g746) & (g349)) + ((g227) & (g209) & (!sk[112]) & (g746) & (!g349)) + ((g227) & (g209) & (!sk[112]) & (g746) & (g349)) + ((g227) & (g209) & (sk[112]) & (!g746) & (g349)) + ((g227) & (g209) & (sk[112]) & (g746) & (!g349)) + ((g227) & (g209) & (sk[112]) & (g746) & (g349)));
	assign g1247 = (((!sk[113]) & (g12) & (!g46) & (!g99)) + ((!sk[113]) & (g12) & (!g46) & (g99)) + ((!sk[113]) & (g12) & (g46) & (!g99)) + ((!sk[113]) & (g12) & (g46) & (g99)) + ((sk[113]) & (!g12) & (g46) & (g99)) + ((sk[113]) & (g12) & (!g46) & (g99)) + ((sk[113]) & (g12) & (g46) & (g99)));
	assign g1248 = (((!g134) & (!g118) & (!g231) & (!sk[114]) & (!g534) & (g478)) + ((!g134) & (!g118) & (!g231) & (!sk[114]) & (g534) & (g478)) + ((!g134) & (!g118) & (!g231) & (sk[114]) & (!g534) & (!g478)) + ((!g134) & (!g118) & (!g231) & (sk[114]) & (!g534) & (g478)) + ((!g134) & (!g118) & (!g231) & (sk[114]) & (g534) & (!g478)) + ((!g134) & (!g118) & (!g231) & (sk[114]) & (g534) & (g478)) + ((!g134) & (!g118) & (g231) & (!sk[114]) & (!g534) & (g478)) + ((!g134) & (!g118) & (g231) & (!sk[114]) & (g534) & (g478)) + ((!g134) & (!g118) & (g231) & (sk[114]) & (!g534) & (!g478)) + ((!g134) & (!g118) & (g231) & (sk[114]) & (!g534) & (g478)) + ((!g134) & (!g118) & (g231) & (sk[114]) & (g534) & (!g478)) + ((!g134) & (!g118) & (g231) & (sk[114]) & (g534) & (g478)) + ((!g134) & (g118) & (!g231) & (!sk[114]) & (!g534) & (g478)) + ((!g134) & (g118) & (!g231) & (!sk[114]) & (g534) & (g478)) + ((!g134) & (g118) & (g231) & (!sk[114]) & (!g534) & (g478)) + ((!g134) & (g118) & (g231) & (!sk[114]) & (g534) & (g478)) + ((!g134) & (g118) & (g231) & (sk[114]) & (!g534) & (!g478)) + ((g134) & (!g118) & (!g231) & (!sk[114]) & (!g534) & (!g478)) + ((g134) & (!g118) & (!g231) & (!sk[114]) & (!g534) & (g478)) + ((g134) & (!g118) & (!g231) & (!sk[114]) & (g534) & (!g478)) + ((g134) & (!g118) & (!g231) & (!sk[114]) & (g534) & (g478)) + ((g134) & (!g118) & (g231) & (!sk[114]) & (!g534) & (!g478)) + ((g134) & (!g118) & (g231) & (!sk[114]) & (!g534) & (g478)) + ((g134) & (!g118) & (g231) & (!sk[114]) & (g534) & (!g478)) + ((g134) & (!g118) & (g231) & (!sk[114]) & (g534) & (g478)) + ((g134) & (!g118) & (g231) & (sk[114]) & (!g534) & (!g478)) + ((g134) & (!g118) & (g231) & (sk[114]) & (!g534) & (g478)) + ((g134) & (!g118) & (g231) & (sk[114]) & (g534) & (!g478)) + ((g134) & (!g118) & (g231) & (sk[114]) & (g534) & (g478)) + ((g134) & (g118) & (!g231) & (!sk[114]) & (!g534) & (!g478)) + ((g134) & (g118) & (!g231) & (!sk[114]) & (!g534) & (g478)) + ((g134) & (g118) & (!g231) & (!sk[114]) & (g534) & (!g478)) + ((g134) & (g118) & (!g231) & (!sk[114]) & (g534) & (g478)) + ((g134) & (g118) & (g231) & (!sk[114]) & (!g534) & (!g478)) + ((g134) & (g118) & (g231) & (!sk[114]) & (!g534) & (g478)) + ((g134) & (g118) & (g231) & (!sk[114]) & (g534) & (!g478)) + ((g134) & (g118) & (g231) & (!sk[114]) & (g534) & (g478)) + ((g134) & (g118) & (g231) & (sk[114]) & (!g534) & (!g478)));
	assign g1249 = (((!g972) & (!g1245) & (!g1246) & (!g1247) & (!sk[115]) & (g1248)) + ((!g972) & (!g1245) & (!g1246) & (!g1247) & (sk[115]) & (g1248)) + ((!g972) & (!g1245) & (!g1246) & (g1247) & (!sk[115]) & (g1248)) + ((!g972) & (!g1245) & (g1246) & (!g1247) & (!sk[115]) & (g1248)) + ((!g972) & (!g1245) & (g1246) & (g1247) & (!sk[115]) & (g1248)) + ((!g972) & (g1245) & (!g1246) & (!g1247) & (!sk[115]) & (g1248)) + ((!g972) & (g1245) & (!g1246) & (g1247) & (!sk[115]) & (g1248)) + ((!g972) & (g1245) & (g1246) & (!g1247) & (!sk[115]) & (g1248)) + ((!g972) & (g1245) & (g1246) & (g1247) & (!sk[115]) & (g1248)) + ((g972) & (!g1245) & (!g1246) & (!g1247) & (!sk[115]) & (!g1248)) + ((g972) & (!g1245) & (!g1246) & (!g1247) & (!sk[115]) & (g1248)) + ((g972) & (!g1245) & (!g1246) & (g1247) & (!sk[115]) & (!g1248)) + ((g972) & (!g1245) & (!g1246) & (g1247) & (!sk[115]) & (g1248)) + ((g972) & (!g1245) & (g1246) & (!g1247) & (!sk[115]) & (!g1248)) + ((g972) & (!g1245) & (g1246) & (!g1247) & (!sk[115]) & (g1248)) + ((g972) & (!g1245) & (g1246) & (g1247) & (!sk[115]) & (!g1248)) + ((g972) & (!g1245) & (g1246) & (g1247) & (!sk[115]) & (g1248)) + ((g972) & (g1245) & (!g1246) & (!g1247) & (!sk[115]) & (!g1248)) + ((g972) & (g1245) & (!g1246) & (!g1247) & (!sk[115]) & (g1248)) + ((g972) & (g1245) & (!g1246) & (g1247) & (!sk[115]) & (!g1248)) + ((g972) & (g1245) & (!g1246) & (g1247) & (!sk[115]) & (g1248)) + ((g972) & (g1245) & (g1246) & (!g1247) & (!sk[115]) & (!g1248)) + ((g972) & (g1245) & (g1246) & (!g1247) & (!sk[115]) & (g1248)) + ((g972) & (g1245) & (g1246) & (g1247) & (!sk[115]) & (!g1248)) + ((g972) & (g1245) & (g1246) & (g1247) & (!sk[115]) & (g1248)));
	assign g1250 = (((g766) & (g1025) & (g1054) & (g1241) & (g1244) & (g1249)));
	assign g1251 = (((!sk[117]) & (!g10) & (!g45) & (g221) & (g534)) + ((!sk[117]) & (!g10) & (g45) & (!g221) & (!g534)) + ((!sk[117]) & (!g10) & (g45) & (!g221) & (g534)) + ((!sk[117]) & (!g10) & (g45) & (g221) & (!g534)) + ((!sk[117]) & (!g10) & (g45) & (g221) & (g534)) + ((!sk[117]) & (g10) & (!g45) & (g221) & (!g534)) + ((!sk[117]) & (g10) & (!g45) & (g221) & (g534)) + ((!sk[117]) & (g10) & (g45) & (!g221) & (!g534)) + ((!sk[117]) & (g10) & (g45) & (!g221) & (g534)) + ((!sk[117]) & (g10) & (g45) & (g221) & (!g534)) + ((!sk[117]) & (g10) & (g45) & (g221) & (g534)) + ((sk[117]) & (!g10) & (!g45) & (g221) & (!g534)));
	assign g1252 = (((!sk[118]) & (!g134) & (!g224) & (g467) & (g817)) + ((!sk[118]) & (!g134) & (g224) & (!g467) & (!g817)) + ((!sk[118]) & (!g134) & (g224) & (!g467) & (g817)) + ((!sk[118]) & (!g134) & (g224) & (g467) & (!g817)) + ((!sk[118]) & (!g134) & (g224) & (g467) & (g817)) + ((!sk[118]) & (g134) & (!g224) & (g467) & (!g817)) + ((!sk[118]) & (g134) & (!g224) & (g467) & (g817)) + ((!sk[118]) & (g134) & (g224) & (!g467) & (!g817)) + ((!sk[118]) & (g134) & (g224) & (!g467) & (g817)) + ((!sk[118]) & (g134) & (g224) & (g467) & (!g817)) + ((!sk[118]) & (g134) & (g224) & (g467) & (g817)) + ((sk[118]) & (g134) & (!g224) & (!g467) & (!g817)) + ((sk[118]) & (g134) & (!g224) & (!g467) & (g817)) + ((sk[118]) & (g134) & (!g224) & (g467) & (g817)) + ((sk[118]) & (g134) & (g224) & (!g467) & (!g817)) + ((sk[118]) & (g134) & (g224) & (!g467) & (g817)) + ((sk[118]) & (g134) & (g224) & (g467) & (!g817)) + ((sk[118]) & (g134) & (g224) & (g467) & (g817)));
	assign g1253 = (((!g214) & (!g946) & (!sk[119]) & (g1251) & (g1252)) + ((!g214) & (!g946) & (sk[119]) & (!g1251) & (!g1252)) + ((!g214) & (!g946) & (sk[119]) & (g1251) & (!g1252)) + ((!g214) & (g946) & (!sk[119]) & (!g1251) & (!g1252)) + ((!g214) & (g946) & (!sk[119]) & (!g1251) & (g1252)) + ((!g214) & (g946) & (!sk[119]) & (g1251) & (!g1252)) + ((!g214) & (g946) & (!sk[119]) & (g1251) & (g1252)) + ((g214) & (!g946) & (!sk[119]) & (g1251) & (!g1252)) + ((g214) & (!g946) & (!sk[119]) & (g1251) & (g1252)) + ((g214) & (!g946) & (sk[119]) & (g1251) & (!g1252)) + ((g214) & (g946) & (!sk[119]) & (!g1251) & (!g1252)) + ((g214) & (g946) & (!sk[119]) & (!g1251) & (g1252)) + ((g214) & (g946) & (!sk[119]) & (g1251) & (!g1252)) + ((g214) & (g946) & (!sk[119]) & (g1251) & (g1252)));
	assign g1254 = (((!i_11_) & (!sk[120]) & (!i_9_) & (!i_10_) & (!g326) & (g238)) + ((!i_11_) & (!sk[120]) & (!i_9_) & (!i_10_) & (g326) & (g238)) + ((!i_11_) & (!sk[120]) & (!i_9_) & (i_10_) & (!g326) & (g238)) + ((!i_11_) & (!sk[120]) & (!i_9_) & (i_10_) & (g326) & (g238)) + ((!i_11_) & (!sk[120]) & (i_9_) & (!i_10_) & (!g326) & (g238)) + ((!i_11_) & (!sk[120]) & (i_9_) & (!i_10_) & (g326) & (g238)) + ((!i_11_) & (!sk[120]) & (i_9_) & (i_10_) & (!g326) & (g238)) + ((!i_11_) & (!sk[120]) & (i_9_) & (i_10_) & (g326) & (g238)) + ((!i_11_) & (sk[120]) & (i_9_) & (i_10_) & (g326) & (g238)) + ((i_11_) & (!sk[120]) & (!i_9_) & (!i_10_) & (!g326) & (!g238)) + ((i_11_) & (!sk[120]) & (!i_9_) & (!i_10_) & (!g326) & (g238)) + ((i_11_) & (!sk[120]) & (!i_9_) & (!i_10_) & (g326) & (!g238)) + ((i_11_) & (!sk[120]) & (!i_9_) & (!i_10_) & (g326) & (g238)) + ((i_11_) & (!sk[120]) & (!i_9_) & (i_10_) & (!g326) & (!g238)) + ((i_11_) & (!sk[120]) & (!i_9_) & (i_10_) & (!g326) & (g238)) + ((i_11_) & (!sk[120]) & (!i_9_) & (i_10_) & (g326) & (!g238)) + ((i_11_) & (!sk[120]) & (!i_9_) & (i_10_) & (g326) & (g238)) + ((i_11_) & (!sk[120]) & (i_9_) & (!i_10_) & (!g326) & (!g238)) + ((i_11_) & (!sk[120]) & (i_9_) & (!i_10_) & (!g326) & (g238)) + ((i_11_) & (!sk[120]) & (i_9_) & (!i_10_) & (g326) & (!g238)) + ((i_11_) & (!sk[120]) & (i_9_) & (!i_10_) & (g326) & (g238)) + ((i_11_) & (!sk[120]) & (i_9_) & (i_10_) & (!g326) & (!g238)) + ((i_11_) & (!sk[120]) & (i_9_) & (i_10_) & (!g326) & (g238)) + ((i_11_) & (!sk[120]) & (i_9_) & (i_10_) & (g326) & (!g238)) + ((i_11_) & (!sk[120]) & (i_9_) & (i_10_) & (g326) & (g238)) + ((i_11_) & (sk[120]) & (i_9_) & (!i_10_) & (g326) & (g238)));
	assign g1255 = (((!i_14_) & (!i_12_) & (!sk[121]) & (i_13_) & (g122)) + ((!i_14_) & (!i_12_) & (sk[121]) & (i_13_) & (!g122)) + ((!i_14_) & (i_12_) & (!sk[121]) & (!i_13_) & (!g122)) + ((!i_14_) & (i_12_) & (!sk[121]) & (!i_13_) & (g122)) + ((!i_14_) & (i_12_) & (!sk[121]) & (i_13_) & (!g122)) + ((!i_14_) & (i_12_) & (!sk[121]) & (i_13_) & (g122)) + ((i_14_) & (!i_12_) & (!sk[121]) & (i_13_) & (!g122)) + ((i_14_) & (!i_12_) & (!sk[121]) & (i_13_) & (g122)) + ((i_14_) & (i_12_) & (!sk[121]) & (!i_13_) & (!g122)) + ((i_14_) & (i_12_) & (!sk[121]) & (!i_13_) & (g122)) + ((i_14_) & (i_12_) & (!sk[121]) & (i_13_) & (!g122)) + ((i_14_) & (i_12_) & (!sk[121]) & (i_13_) & (g122)) + ((i_14_) & (i_12_) & (sk[121]) & (i_13_) & (!g122)));
	assign g1256 = (((!g109) & (!g186) & (!g330) & (!sk[122]) & (!g544) & (g1255)) + ((!g109) & (!g186) & (!g330) & (!sk[122]) & (g544) & (g1255)) + ((!g109) & (!g186) & (!g330) & (sk[122]) & (g544) & (!g1255)) + ((!g109) & (!g186) & (!g330) & (sk[122]) & (g544) & (g1255)) + ((!g109) & (!g186) & (g330) & (!sk[122]) & (!g544) & (g1255)) + ((!g109) & (!g186) & (g330) & (!sk[122]) & (g544) & (g1255)) + ((!g109) & (!g186) & (g330) & (sk[122]) & (!g544) & (!g1255)) + ((!g109) & (!g186) & (g330) & (sk[122]) & (!g544) & (g1255)) + ((!g109) & (!g186) & (g330) & (sk[122]) & (g544) & (!g1255)) + ((!g109) & (!g186) & (g330) & (sk[122]) & (g544) & (g1255)) + ((!g109) & (g186) & (!g330) & (!sk[122]) & (!g544) & (g1255)) + ((!g109) & (g186) & (!g330) & (!sk[122]) & (g544) & (g1255)) + ((!g109) & (g186) & (!g330) & (sk[122]) & (g544) & (!g1255)) + ((!g109) & (g186) & (!g330) & (sk[122]) & (g544) & (g1255)) + ((!g109) & (g186) & (g330) & (!sk[122]) & (!g544) & (g1255)) + ((!g109) & (g186) & (g330) & (!sk[122]) & (g544) & (g1255)) + ((!g109) & (g186) & (g330) & (sk[122]) & (g544) & (!g1255)) + ((!g109) & (g186) & (g330) & (sk[122]) & (g544) & (g1255)) + ((g109) & (!g186) & (!g330) & (!sk[122]) & (!g544) & (!g1255)) + ((g109) & (!g186) & (!g330) & (!sk[122]) & (!g544) & (g1255)) + ((g109) & (!g186) & (!g330) & (!sk[122]) & (g544) & (!g1255)) + ((g109) & (!g186) & (!g330) & (!sk[122]) & (g544) & (g1255)) + ((g109) & (!g186) & (!g330) & (sk[122]) & (g544) & (!g1255)) + ((g109) & (!g186) & (g330) & (!sk[122]) & (!g544) & (!g1255)) + ((g109) & (!g186) & (g330) & (!sk[122]) & (!g544) & (g1255)) + ((g109) & (!g186) & (g330) & (!sk[122]) & (g544) & (!g1255)) + ((g109) & (!g186) & (g330) & (!sk[122]) & (g544) & (g1255)) + ((g109) & (!g186) & (g330) & (sk[122]) & (g544) & (!g1255)) + ((g109) & (g186) & (!g330) & (!sk[122]) & (!g544) & (!g1255)) + ((g109) & (g186) & (!g330) & (!sk[122]) & (!g544) & (g1255)) + ((g109) & (g186) & (!g330) & (!sk[122]) & (g544) & (!g1255)) + ((g109) & (g186) & (!g330) & (!sk[122]) & (g544) & (g1255)) + ((g109) & (g186) & (!g330) & (sk[122]) & (g544) & (!g1255)) + ((g109) & (g186) & (g330) & (!sk[122]) & (!g544) & (!g1255)) + ((g109) & (g186) & (g330) & (!sk[122]) & (!g544) & (g1255)) + ((g109) & (g186) & (g330) & (!sk[122]) & (g544) & (!g1255)) + ((g109) & (g186) & (g330) & (!sk[122]) & (g544) & (g1255)) + ((g109) & (g186) & (g330) & (sk[122]) & (g544) & (!g1255)));
	assign g1257 = (((g242) & (g1253) & (g1047) & (g1051) & (!g1254) & (g1256)));
	assign g1258 = (((g890) & (g1229) & (g1235) & (g1239) & (g1250) & (g1257)));
	assign g1259 = (((!g1065) & (!g1158) & (sk[125]) & (g1163)) + ((g1065) & (!g1158) & (!sk[125]) & (!g1163)) + ((g1065) & (!g1158) & (!sk[125]) & (g1163)) + ((g1065) & (g1158) & (!sk[125]) & (!g1163)) + ((g1065) & (g1158) & (!sk[125]) & (g1163)));
	assign g1260 = (((!sk[126]) & (g187) & (!g534) & (!g702)) + ((!sk[126]) & (g187) & (!g534) & (g702)) + ((!sk[126]) & (g187) & (g534) & (!g702)) + ((!sk[126]) & (g187) & (g534) & (g702)) + ((sk[126]) & (!g187) & (!g534) & (!g702)));
	assign g1261 = (((!g89) & (!g109) & (!sk[127]) & (g1099) & (g1260)) + ((!g89) & (!g109) & (sk[127]) & (!g1099) & (!g1260)) + ((!g89) & (!g109) & (sk[127]) & (!g1099) & (g1260)) + ((!g89) & (g109) & (!sk[127]) & (!g1099) & (!g1260)) + ((!g89) & (g109) & (!sk[127]) & (!g1099) & (g1260)) + ((!g89) & (g109) & (!sk[127]) & (g1099) & (!g1260)) + ((!g89) & (g109) & (!sk[127]) & (g1099) & (g1260)) + ((!g89) & (g109) & (sk[127]) & (!g1099) & (!g1260)) + ((!g89) & (g109) & (sk[127]) & (!g1099) & (g1260)) + ((!g89) & (g109) & (sk[127]) & (g1099) & (!g1260)) + ((g89) & (!g109) & (!sk[127]) & (g1099) & (!g1260)) + ((g89) & (!g109) & (!sk[127]) & (g1099) & (g1260)) + ((g89) & (g109) & (!sk[127]) & (!g1099) & (!g1260)) + ((g89) & (g109) & (!sk[127]) & (!g1099) & (g1260)) + ((g89) & (g109) & (!sk[127]) & (g1099) & (!g1260)) + ((g89) & (g109) & (!sk[127]) & (g1099) & (g1260)) + ((g89) & (g109) & (sk[127]) & (!g1099) & (!g1260)) + ((g89) & (g109) & (sk[127]) & (g1099) & (!g1260)));
	assign g1262 = (((!i_8_) & (!g134) & (!g135) & (!g187) & (!g534) & (!g702)) + ((!i_8_) & (!g134) & (!g135) & (!g187) & (!g534) & (g702)) + ((!i_8_) & (!g134) & (!g135) & (!g187) & (g534) & (!g702)) + ((!i_8_) & (!g134) & (!g135) & (!g187) & (g534) & (g702)) + ((!i_8_) & (!g134) & (!g135) & (g187) & (!g534) & (!g702)) + ((!i_8_) & (!g134) & (!g135) & (g187) & (!g534) & (g702)) + ((!i_8_) & (!g134) & (!g135) & (g187) & (g534) & (!g702)) + ((!i_8_) & (!g134) & (!g135) & (g187) & (g534) & (g702)) + ((!i_8_) & (!g134) & (g135) & (!g187) & (!g534) & (!g702)) + ((!i_8_) & (!g134) & (g135) & (!g187) & (!g534) & (g702)) + ((!i_8_) & (!g134) & (g135) & (!g187) & (g534) & (!g702)) + ((!i_8_) & (!g134) & (g135) & (!g187) & (g534) & (g702)) + ((!i_8_) & (!g134) & (g135) & (g187) & (!g534) & (!g702)) + ((!i_8_) & (!g134) & (g135) & (g187) & (!g534) & (g702)) + ((!i_8_) & (!g134) & (g135) & (g187) & (g534) & (!g702)) + ((!i_8_) & (!g134) & (g135) & (g187) & (g534) & (g702)) + ((!i_8_) & (g134) & (!g135) & (!g187) & (!g534) & (!g702)) + ((!i_8_) & (g134) & (g135) & (!g187) & (!g534) & (!g702)) + ((i_8_) & (!g134) & (!g135) & (!g187) & (!g534) & (!g702)) + ((i_8_) & (!g134) & (!g135) & (!g187) & (!g534) & (g702)) + ((i_8_) & (!g134) & (!g135) & (!g187) & (g534) & (!g702)) + ((i_8_) & (!g134) & (!g135) & (!g187) & (g534) & (g702)) + ((i_8_) & (!g134) & (!g135) & (g187) & (!g534) & (!g702)) + ((i_8_) & (!g134) & (!g135) & (g187) & (!g534) & (g702)) + ((i_8_) & (!g134) & (!g135) & (g187) & (g534) & (!g702)) + ((i_8_) & (!g134) & (!g135) & (g187) & (g534) & (g702)) + ((i_8_) & (!g134) & (g135) & (!g187) & (!g534) & (!g702)) + ((i_8_) & (!g134) & (g135) & (!g187) & (!g534) & (g702)) + ((i_8_) & (g134) & (!g135) & (!g187) & (!g534) & (!g702)) + ((i_8_) & (g134) & (g135) & (!g187) & (!g534) & (!g702)));
	assign g1263 = (((!g136) & (!g231) & (!g478) & (!sk[1]) & (!g922) & (g1262)) + ((!g136) & (!g231) & (!g478) & (!sk[1]) & (g922) & (g1262)) + ((!g136) & (!g231) & (!g478) & (sk[1]) & (!g922) & (g1262)) + ((!g136) & (!g231) & (g478) & (!sk[1]) & (!g922) & (g1262)) + ((!g136) & (!g231) & (g478) & (!sk[1]) & (g922) & (g1262)) + ((!g136) & (!g231) & (g478) & (sk[1]) & (!g922) & (g1262)) + ((!g136) & (g231) & (!g478) & (!sk[1]) & (!g922) & (g1262)) + ((!g136) & (g231) & (!g478) & (!sk[1]) & (g922) & (g1262)) + ((!g136) & (g231) & (!g478) & (sk[1]) & (!g922) & (g1262)) + ((!g136) & (g231) & (g478) & (!sk[1]) & (!g922) & (g1262)) + ((!g136) & (g231) & (g478) & (!sk[1]) & (g922) & (g1262)) + ((!g136) & (g231) & (g478) & (sk[1]) & (!g922) & (g1262)) + ((g136) & (!g231) & (!g478) & (!sk[1]) & (!g922) & (!g1262)) + ((g136) & (!g231) & (!g478) & (!sk[1]) & (!g922) & (g1262)) + ((g136) & (!g231) & (!g478) & (!sk[1]) & (g922) & (!g1262)) + ((g136) & (!g231) & (!g478) & (!sk[1]) & (g922) & (g1262)) + ((g136) & (!g231) & (g478) & (!sk[1]) & (!g922) & (!g1262)) + ((g136) & (!g231) & (g478) & (!sk[1]) & (!g922) & (g1262)) + ((g136) & (!g231) & (g478) & (!sk[1]) & (g922) & (!g1262)) + ((g136) & (!g231) & (g478) & (!sk[1]) & (g922) & (g1262)) + ((g136) & (g231) & (!g478) & (!sk[1]) & (!g922) & (!g1262)) + ((g136) & (g231) & (!g478) & (!sk[1]) & (!g922) & (g1262)) + ((g136) & (g231) & (!g478) & (!sk[1]) & (g922) & (!g1262)) + ((g136) & (g231) & (!g478) & (!sk[1]) & (g922) & (g1262)) + ((g136) & (g231) & (!g478) & (sk[1]) & (!g922) & (g1262)) + ((g136) & (g231) & (g478) & (!sk[1]) & (!g922) & (!g1262)) + ((g136) & (g231) & (g478) & (!sk[1]) & (!g922) & (g1262)) + ((g136) & (g231) & (g478) & (!sk[1]) & (g922) & (!g1262)) + ((g136) & (g231) & (g478) & (!sk[1]) & (g922) & (g1262)));
	assign g1264 = (((!g134) & (!g99) & (!g105) & (!g837) & (!g696) & (!g702)) + ((!g134) & (!g99) & (!g105) & (!g837) & (!g696) & (g702)) + ((!g134) & (!g99) & (!g105) & (!g837) & (g696) & (!g702)) + ((!g134) & (!g99) & (!g105) & (!g837) & (g696) & (g702)) + ((!g134) & (!g99) & (!g105) & (g837) & (!g696) & (!g702)) + ((!g134) & (!g99) & (!g105) & (g837) & (!g696) & (g702)) + ((!g134) & (!g99) & (!g105) & (g837) & (g696) & (!g702)) + ((!g134) & (!g99) & (!g105) & (g837) & (g696) & (g702)) + ((!g134) & (!g99) & (g105) & (!g837) & (!g696) & (!g702)) + ((!g134) & (!g99) & (g105) & (!g837) & (!g696) & (g702)) + ((!g134) & (!g99) & (g105) & (!g837) & (g696) & (!g702)) + ((!g134) & (!g99) & (g105) & (!g837) & (g696) & (g702)) + ((!g134) & (!g99) & (g105) & (g837) & (!g696) & (!g702)) + ((!g134) & (!g99) & (g105) & (g837) & (!g696) & (g702)) + ((!g134) & (!g99) & (g105) & (g837) & (g696) & (!g702)) + ((!g134) & (!g99) & (g105) & (g837) & (g696) & (g702)) + ((!g134) & (g99) & (!g105) & (!g837) & (!g696) & (!g702)) + ((!g134) & (g99) & (!g105) & (!g837) & (g696) & (!g702)) + ((!g134) & (g99) & (!g105) & (g837) & (!g696) & (!g702)) + ((!g134) & (g99) & (!g105) & (g837) & (g696) & (!g702)) + ((!g134) & (g99) & (g105) & (!g837) & (!g696) & (!g702)) + ((!g134) & (g99) & (g105) & (!g837) & (g696) & (!g702)) + ((!g134) & (g99) & (g105) & (g837) & (!g696) & (!g702)) + ((!g134) & (g99) & (g105) & (g837) & (g696) & (!g702)) + ((g134) & (!g99) & (!g105) & (g837) & (g696) & (!g702)) + ((g134) & (!g99) & (!g105) & (g837) & (g696) & (g702)) + ((g134) & (g99) & (!g105) & (g837) & (g696) & (!g702)));
	assign g1265 = (((g945) & (!g1063) & (!g1261) & (g1263) & (!g1133) & (g1264)));
	assign g1266 = (((!sk[4]) & (g101) & (!g1184)) + ((!sk[4]) & (g101) & (g1184)) + ((sk[4]) & (g101) & (!g1184)));
	assign g1267 = (((!g99) & (!g195) & (!sk[5]) & (g105) & (g696)) + ((!g99) & (g195) & (!sk[5]) & (!g105) & (!g696)) + ((!g99) & (g195) & (!sk[5]) & (!g105) & (g696)) + ((!g99) & (g195) & (!sk[5]) & (g105) & (!g696)) + ((!g99) & (g195) & (!sk[5]) & (g105) & (g696)) + ((g99) & (!g195) & (!sk[5]) & (g105) & (!g696)) + ((g99) & (!g195) & (!sk[5]) & (g105) & (g696)) + ((g99) & (!g195) & (sk[5]) & (!g105) & (!g696)) + ((g99) & (!g195) & (sk[5]) & (g105) & (!g696)) + ((g99) & (!g195) & (sk[5]) & (g105) & (g696)) + ((g99) & (g195) & (!sk[5]) & (!g105) & (!g696)) + ((g99) & (g195) & (!sk[5]) & (!g105) & (g696)) + ((g99) & (g195) & (!sk[5]) & (g105) & (!g696)) + ((g99) & (g195) & (!sk[5]) & (g105) & (g696)) + ((g99) & (g195) & (sk[5]) & (!g105) & (!g696)) + ((g99) & (g195) & (sk[5]) & (!g105) & (g696)) + ((g99) & (g195) & (sk[5]) & (g105) & (!g696)) + ((g99) & (g195) & (sk[5]) & (g105) & (g696)));
	assign g1268 = (((!g99) & (!sk[6]) & (!g101) & (!g573) & (!g837) & (g1267)) + ((!g99) & (!sk[6]) & (!g101) & (!g573) & (g837) & (g1267)) + ((!g99) & (!sk[6]) & (!g101) & (g573) & (!g837) & (g1267)) + ((!g99) & (!sk[6]) & (!g101) & (g573) & (g837) & (g1267)) + ((!g99) & (!sk[6]) & (g101) & (!g573) & (!g837) & (g1267)) + ((!g99) & (!sk[6]) & (g101) & (!g573) & (g837) & (g1267)) + ((!g99) & (!sk[6]) & (g101) & (g573) & (!g837) & (g1267)) + ((!g99) & (!sk[6]) & (g101) & (g573) & (g837) & (g1267)) + ((!g99) & (sk[6]) & (!g101) & (!g573) & (!g837) & (!g1267)) + ((!g99) & (sk[6]) & (!g101) & (!g573) & (g837) & (!g1267)) + ((!g99) & (sk[6]) & (g101) & (!g573) & (g837) & (!g1267)) + ((g99) & (!sk[6]) & (!g101) & (!g573) & (!g837) & (!g1267)) + ((g99) & (!sk[6]) & (!g101) & (!g573) & (!g837) & (g1267)) + ((g99) & (!sk[6]) & (!g101) & (!g573) & (g837) & (!g1267)) + ((g99) & (!sk[6]) & (!g101) & (!g573) & (g837) & (g1267)) + ((g99) & (!sk[6]) & (!g101) & (g573) & (!g837) & (!g1267)) + ((g99) & (!sk[6]) & (!g101) & (g573) & (!g837) & (g1267)) + ((g99) & (!sk[6]) & (!g101) & (g573) & (g837) & (!g1267)) + ((g99) & (!sk[6]) & (!g101) & (g573) & (g837) & (g1267)) + ((g99) & (!sk[6]) & (g101) & (!g573) & (!g837) & (!g1267)) + ((g99) & (!sk[6]) & (g101) & (!g573) & (!g837) & (g1267)) + ((g99) & (!sk[6]) & (g101) & (!g573) & (g837) & (!g1267)) + ((g99) & (!sk[6]) & (g101) & (!g573) & (g837) & (g1267)) + ((g99) & (!sk[6]) & (g101) & (g573) & (!g837) & (!g1267)) + ((g99) & (!sk[6]) & (g101) & (g573) & (!g837) & (g1267)) + ((g99) & (!sk[6]) & (g101) & (g573) & (g837) & (!g1267)) + ((g99) & (!sk[6]) & (g101) & (g573) & (g837) & (g1267)) + ((g99) & (sk[6]) & (!g101) & (!g573) & (g837) & (!g1267)) + ((g99) & (sk[6]) & (g101) & (!g573) & (g837) & (!g1267)));
	assign g1269 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g104) & (!g112) & (!g124)) + ((!i_14_) & (!i_12_) & (!i_13_) & (!g104) & (!g112) & (g124)) + ((!i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g112) & (!g124)) + ((!i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g112) & (g124)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g104) & (!g112) & (!g124)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g104) & (!g112) & (g124)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g104) & (!g112) & (!g124)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g104) & (g112) & (!g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g104) & (!g112) & (!g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g104) & (!g112) & (g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g104) & (g112) & (!g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g104) & (g112) & (g124)) + ((!i_14_) & (i_12_) & (i_13_) & (!g104) & (!g112) & (!g124)) + ((!i_14_) & (i_12_) & (i_13_) & (!g104) & (g112) & (!g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g104) & (!g112) & (!g124)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g104) & (g112) & (!g124)) + ((i_14_) & (!i_12_) & (i_13_) & (!g104) & (!g112) & (!g124)) + ((i_14_) & (!i_12_) & (i_13_) & (!g104) & (!g112) & (g124)) + ((i_14_) & (!i_12_) & (i_13_) & (!g104) & (g112) & (!g124)) + ((i_14_) & (!i_12_) & (i_13_) & (!g104) & (g112) & (g124)) + ((i_14_) & (i_12_) & (!i_13_) & (!g104) & (!g112) & (!g124)) + ((i_14_) & (i_12_) & (!i_13_) & (!g104) & (!g112) & (g124)) + ((i_14_) & (i_12_) & (!i_13_) & (!g104) & (g112) & (!g124)) + ((i_14_) & (i_12_) & (!i_13_) & (!g104) & (g112) & (g124)) + ((i_14_) & (i_12_) & (!i_13_) & (g104) & (!g112) & (!g124)) + ((i_14_) & (i_12_) & (!i_13_) & (g104) & (!g112) & (g124)) + ((i_14_) & (i_12_) & (!i_13_) & (g104) & (g112) & (!g124)) + ((i_14_) & (i_12_) & (!i_13_) & (g104) & (g112) & (g124)) + ((i_14_) & (i_12_) & (i_13_) & (!g104) & (!g112) & (!g124)) + ((i_14_) & (i_12_) & (i_13_) & (!g104) & (!g112) & (g124)) + ((i_14_) & (i_12_) & (i_13_) & (!g104) & (g112) & (!g124)) + ((i_14_) & (i_12_) & (i_13_) & (!g104) & (g112) & (g124)));
	assign g1270 = (((!sk[8]) & (!i_8_) & (!g495) & (g982) & (g1269)) + ((!sk[8]) & (!i_8_) & (g495) & (!g982) & (!g1269)) + ((!sk[8]) & (!i_8_) & (g495) & (!g982) & (g1269)) + ((!sk[8]) & (!i_8_) & (g495) & (g982) & (!g1269)) + ((!sk[8]) & (!i_8_) & (g495) & (g982) & (g1269)) + ((!sk[8]) & (i_8_) & (!g495) & (g982) & (!g1269)) + ((!sk[8]) & (i_8_) & (!g495) & (g982) & (g1269)) + ((!sk[8]) & (i_8_) & (g495) & (!g982) & (!g1269)) + ((!sk[8]) & (i_8_) & (g495) & (!g982) & (g1269)) + ((!sk[8]) & (i_8_) & (g495) & (g982) & (!g1269)) + ((!sk[8]) & (i_8_) & (g495) & (g982) & (g1269)) + ((sk[8]) & (!i_8_) & (g495) & (!g982) & (!g1269)) + ((sk[8]) & (!i_8_) & (g495) & (g982) & (!g1269)) + ((sk[8]) & (i_8_) & (g495) & (!g982) & (!g1269)));
	assign g1271 = (((!i_14_) & (!i_12_) & (!i_13_) & (g118) & (!g112) & (g124)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g118) & (g112) & (g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (g118) & (!g112) & (g124)) + ((!i_14_) & (i_12_) & (!i_13_) & (g118) & (g112) & (g124)) + ((i_14_) & (!i_12_) & (i_13_) & (!g118) & (g112) & (g124)) + ((i_14_) & (!i_12_) & (i_13_) & (g118) & (g112) & (g124)) + ((i_14_) & (i_12_) & (!i_13_) & (!g118) & (g112) & (g124)) + ((i_14_) & (i_12_) & (!i_13_) & (g118) & (g112) & (g124)) + ((i_14_) & (i_12_) & (i_13_) & (!g118) & (g112) & (g124)) + ((i_14_) & (i_12_) & (i_13_) & (g118) & (g112) & (g124)));
	assign g1272 = (((!i_11_) & (!g113) & (!g112) & (!g187) & (!g236) & (!g1271)) + ((!i_11_) & (!g113) & (!g112) & (!g187) & (g236) & (!g1271)) + ((!i_11_) & (!g113) & (!g112) & (g187) & (!g236) & (!g1271)) + ((!i_11_) & (!g113) & (!g112) & (g187) & (g236) & (!g1271)) + ((!i_11_) & (!g113) & (g112) & (!g187) & (!g236) & (!g1271)) + ((!i_11_) & (!g113) & (g112) & (!g187) & (g236) & (!g1271)) + ((!i_11_) & (g113) & (!g112) & (!g187) & (!g236) & (!g1271)) + ((!i_11_) & (g113) & (!g112) & (!g187) & (g236) & (!g1271)) + ((!i_11_) & (g113) & (!g112) & (g187) & (!g236) & (!g1271)) + ((!i_11_) & (g113) & (!g112) & (g187) & (g236) & (!g1271)) + ((!i_11_) & (g113) & (g112) & (!g187) & (!g236) & (!g1271)) + ((!i_11_) & (g113) & (g112) & (!g187) & (g236) & (!g1271)) + ((i_11_) & (!g113) & (!g112) & (!g187) & (!g236) & (!g1271)) + ((i_11_) & (!g113) & (!g112) & (!g187) & (g236) & (!g1271)) + ((i_11_) & (!g113) & (!g112) & (g187) & (!g236) & (!g1271)) + ((i_11_) & (!g113) & (!g112) & (g187) & (g236) & (!g1271)) + ((i_11_) & (!g113) & (g112) & (!g187) & (!g236) & (!g1271)) + ((i_11_) & (!g113) & (g112) & (!g187) & (g236) & (!g1271)) + ((i_11_) & (g113) & (!g112) & (!g187) & (!g236) & (!g1271)) + ((i_11_) & (g113) & (!g112) & (g187) & (!g236) & (!g1271)) + ((i_11_) & (g113) & (g112) & (!g187) & (!g236) & (!g1271)));
	assign g1273 = (((!g931) & (!g1266) & (!g1268) & (!g1270) & (!sk[11]) & (g1272)) + ((!g931) & (!g1266) & (!g1268) & (g1270) & (!sk[11]) & (g1272)) + ((!g931) & (!g1266) & (g1268) & (!g1270) & (!sk[11]) & (g1272)) + ((!g931) & (!g1266) & (g1268) & (!g1270) & (sk[11]) & (g1272)) + ((!g931) & (!g1266) & (g1268) & (g1270) & (!sk[11]) & (g1272)) + ((!g931) & (g1266) & (!g1268) & (!g1270) & (!sk[11]) & (g1272)) + ((!g931) & (g1266) & (!g1268) & (g1270) & (!sk[11]) & (g1272)) + ((!g931) & (g1266) & (g1268) & (!g1270) & (!sk[11]) & (g1272)) + ((!g931) & (g1266) & (g1268) & (g1270) & (!sk[11]) & (g1272)) + ((g931) & (!g1266) & (!g1268) & (!g1270) & (!sk[11]) & (!g1272)) + ((g931) & (!g1266) & (!g1268) & (!g1270) & (!sk[11]) & (g1272)) + ((g931) & (!g1266) & (!g1268) & (g1270) & (!sk[11]) & (!g1272)) + ((g931) & (!g1266) & (!g1268) & (g1270) & (!sk[11]) & (g1272)) + ((g931) & (!g1266) & (g1268) & (!g1270) & (!sk[11]) & (!g1272)) + ((g931) & (!g1266) & (g1268) & (!g1270) & (!sk[11]) & (g1272)) + ((g931) & (!g1266) & (g1268) & (g1270) & (!sk[11]) & (!g1272)) + ((g931) & (!g1266) & (g1268) & (g1270) & (!sk[11]) & (g1272)) + ((g931) & (g1266) & (!g1268) & (!g1270) & (!sk[11]) & (!g1272)) + ((g931) & (g1266) & (!g1268) & (!g1270) & (!sk[11]) & (g1272)) + ((g931) & (g1266) & (!g1268) & (g1270) & (!sk[11]) & (!g1272)) + ((g931) & (g1266) & (!g1268) & (g1270) & (!sk[11]) & (g1272)) + ((g931) & (g1266) & (g1268) & (!g1270) & (!sk[11]) & (!g1272)) + ((g931) & (g1266) & (g1268) & (!g1270) & (!sk[11]) & (g1272)) + ((g931) & (g1266) & (g1268) & (g1270) & (!sk[11]) & (!g1272)) + ((g931) & (g1266) & (g1268) & (g1270) & (!sk[11]) & (g1272)));
	assign g1274 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g119) & (g118) & (!g122)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g119) & (g118) & (!g122)) + ((!i_14_) & (!i_12_) & (i_13_) & (!g119) & (g118) & (!g122)) + ((!i_14_) & (!i_12_) & (i_13_) & (g119) & (g118) & (!g122)) + ((!i_14_) & (!i_12_) & (i_13_) & (g119) & (g118) & (g122)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g119) & (g118) & (!g122)) + ((!i_14_) & (i_12_) & (!i_13_) & (g119) & (g118) & (!g122)) + ((!i_14_) & (i_12_) & (!i_13_) & (g119) & (g118) & (g122)) + ((!i_14_) & (i_12_) & (i_13_) & (!g119) & (g118) & (!g122)) + ((!i_14_) & (i_12_) & (i_13_) & (g119) & (g118) & (!g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (g119) & (g118) & (!g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (g119) & (g118) & (g122)) + ((i_14_) & (!i_12_) & (i_13_) & (!g119) & (g118) & (!g122)) + ((i_14_) & (!i_12_) & (i_13_) & (g119) & (g118) & (!g122)) + ((i_14_) & (!i_12_) & (i_13_) & (g119) & (g118) & (g122)) + ((i_14_) & (i_12_) & (!i_13_) & (!g119) & (g118) & (!g122)) + ((i_14_) & (i_12_) & (!i_13_) & (g119) & (g118) & (!g122)) + ((i_14_) & (i_12_) & (!i_13_) & (g119) & (g118) & (g122)));
	assign g1275 = (((!i_11_) & (!sk[13]) & (!i_9_) & (!i_10_) & (!g236) & (g1274)) + ((!i_11_) & (!sk[13]) & (!i_9_) & (!i_10_) & (g236) & (g1274)) + ((!i_11_) & (!sk[13]) & (!i_9_) & (i_10_) & (!g236) & (g1274)) + ((!i_11_) & (!sk[13]) & (!i_9_) & (i_10_) & (g236) & (g1274)) + ((!i_11_) & (!sk[13]) & (i_9_) & (!i_10_) & (!g236) & (g1274)) + ((!i_11_) & (!sk[13]) & (i_9_) & (!i_10_) & (g236) & (g1274)) + ((!i_11_) & (!sk[13]) & (i_9_) & (i_10_) & (!g236) & (g1274)) + ((!i_11_) & (!sk[13]) & (i_9_) & (i_10_) & (g236) & (g1274)) + ((!i_11_) & (sk[13]) & (!i_9_) & (!i_10_) & (!g236) & (!g1274)) + ((!i_11_) & (sk[13]) & (!i_9_) & (!i_10_) & (g236) & (!g1274)) + ((!i_11_) & (sk[13]) & (!i_9_) & (i_10_) & (!g236) & (!g1274)) + ((!i_11_) & (sk[13]) & (!i_9_) & (i_10_) & (g236) & (!g1274)) + ((!i_11_) & (sk[13]) & (i_9_) & (!i_10_) & (!g236) & (!g1274)) + ((!i_11_) & (sk[13]) & (i_9_) & (!i_10_) & (g236) & (!g1274)) + ((!i_11_) & (sk[13]) & (i_9_) & (i_10_) & (!g236) & (!g1274)) + ((!i_11_) & (sk[13]) & (i_9_) & (i_10_) & (g236) & (!g1274)) + ((i_11_) & (!sk[13]) & (!i_9_) & (!i_10_) & (!g236) & (!g1274)) + ((i_11_) & (!sk[13]) & (!i_9_) & (!i_10_) & (!g236) & (g1274)) + ((i_11_) & (!sk[13]) & (!i_9_) & (!i_10_) & (g236) & (!g1274)) + ((i_11_) & (!sk[13]) & (!i_9_) & (!i_10_) & (g236) & (g1274)) + ((i_11_) & (!sk[13]) & (!i_9_) & (i_10_) & (!g236) & (!g1274)) + ((i_11_) & (!sk[13]) & (!i_9_) & (i_10_) & (!g236) & (g1274)) + ((i_11_) & (!sk[13]) & (!i_9_) & (i_10_) & (g236) & (!g1274)) + ((i_11_) & (!sk[13]) & (!i_9_) & (i_10_) & (g236) & (g1274)) + ((i_11_) & (!sk[13]) & (i_9_) & (!i_10_) & (!g236) & (!g1274)) + ((i_11_) & (!sk[13]) & (i_9_) & (!i_10_) & (!g236) & (g1274)) + ((i_11_) & (!sk[13]) & (i_9_) & (!i_10_) & (g236) & (!g1274)) + ((i_11_) & (!sk[13]) & (i_9_) & (!i_10_) & (g236) & (g1274)) + ((i_11_) & (!sk[13]) & (i_9_) & (i_10_) & (!g236) & (!g1274)) + ((i_11_) & (!sk[13]) & (i_9_) & (i_10_) & (!g236) & (g1274)) + ((i_11_) & (!sk[13]) & (i_9_) & (i_10_) & (g236) & (!g1274)) + ((i_11_) & (!sk[13]) & (i_9_) & (i_10_) & (g236) & (g1274)) + ((i_11_) & (sk[13]) & (!i_9_) & (!i_10_) & (!g236) & (!g1274)) + ((i_11_) & (sk[13]) & (!i_9_) & (!i_10_) & (g236) & (!g1274)) + ((i_11_) & (sk[13]) & (!i_9_) & (i_10_) & (!g236) & (!g1274)) + ((i_11_) & (sk[13]) & (!i_9_) & (i_10_) & (g236) & (!g1274)) + ((i_11_) & (sk[13]) & (i_9_) & (!i_10_) & (!g236) & (!g1274)) + ((i_11_) & (sk[13]) & (i_9_) & (i_10_) & (!g236) & (!g1274)) + ((i_11_) & (sk[13]) & (i_9_) & (i_10_) & (g236) & (!g1274)));
	assign g1276 = (((!sk[14]) & (!i_8_) & (!g108) & (g216) & (g548)) + ((!sk[14]) & (!i_8_) & (g108) & (!g216) & (!g548)) + ((!sk[14]) & (!i_8_) & (g108) & (!g216) & (g548)) + ((!sk[14]) & (!i_8_) & (g108) & (g216) & (!g548)) + ((!sk[14]) & (!i_8_) & (g108) & (g216) & (g548)) + ((!sk[14]) & (i_8_) & (!g108) & (g216) & (!g548)) + ((!sk[14]) & (i_8_) & (!g108) & (g216) & (g548)) + ((!sk[14]) & (i_8_) & (g108) & (!g216) & (!g548)) + ((!sk[14]) & (i_8_) & (g108) & (!g216) & (g548)) + ((!sk[14]) & (i_8_) & (g108) & (g216) & (!g548)) + ((!sk[14]) & (i_8_) & (g108) & (g216) & (g548)) + ((sk[14]) & (!i_8_) & (g108) & (!g216) & (g548)) + ((sk[14]) & (!i_8_) & (g108) & (g216) & (g548)) + ((sk[14]) & (i_8_) & (g108) & (!g216) & (g548)) + ((sk[14]) & (i_8_) & (g108) & (g216) & (!g548)) + ((sk[14]) & (i_8_) & (g108) & (g216) & (g548)));
	assign g1277 = (((!i_8_) & (!sk[15]) & (!g181) & (!g108) & (!g123) & (g485)) + ((!i_8_) & (!sk[15]) & (!g181) & (!g108) & (g123) & (g485)) + ((!i_8_) & (!sk[15]) & (!g181) & (g108) & (!g123) & (g485)) + ((!i_8_) & (!sk[15]) & (!g181) & (g108) & (g123) & (g485)) + ((!i_8_) & (!sk[15]) & (g181) & (!g108) & (!g123) & (g485)) + ((!i_8_) & (!sk[15]) & (g181) & (!g108) & (g123) & (g485)) + ((!i_8_) & (!sk[15]) & (g181) & (g108) & (!g123) & (g485)) + ((!i_8_) & (!sk[15]) & (g181) & (g108) & (g123) & (g485)) + ((!i_8_) & (sk[15]) & (!g181) & (g108) & (!g123) & (g485)) + ((!i_8_) & (sk[15]) & (!g181) & (g108) & (g123) & (!g485)) + ((!i_8_) & (sk[15]) & (!g181) & (g108) & (g123) & (g485)) + ((!i_8_) & (sk[15]) & (g181) & (g108) & (!g123) & (!g485)) + ((!i_8_) & (sk[15]) & (g181) & (g108) & (!g123) & (g485)) + ((!i_8_) & (sk[15]) & (g181) & (g108) & (g123) & (!g485)) + ((!i_8_) & (sk[15]) & (g181) & (g108) & (g123) & (g485)) + ((i_8_) & (!sk[15]) & (!g181) & (!g108) & (!g123) & (!g485)) + ((i_8_) & (!sk[15]) & (!g181) & (!g108) & (!g123) & (g485)) + ((i_8_) & (!sk[15]) & (!g181) & (!g108) & (g123) & (!g485)) + ((i_8_) & (!sk[15]) & (!g181) & (!g108) & (g123) & (g485)) + ((i_8_) & (!sk[15]) & (!g181) & (g108) & (!g123) & (!g485)) + ((i_8_) & (!sk[15]) & (!g181) & (g108) & (!g123) & (g485)) + ((i_8_) & (!sk[15]) & (!g181) & (g108) & (g123) & (!g485)) + ((i_8_) & (!sk[15]) & (!g181) & (g108) & (g123) & (g485)) + ((i_8_) & (!sk[15]) & (g181) & (!g108) & (!g123) & (!g485)) + ((i_8_) & (!sk[15]) & (g181) & (!g108) & (!g123) & (g485)) + ((i_8_) & (!sk[15]) & (g181) & (!g108) & (g123) & (!g485)) + ((i_8_) & (!sk[15]) & (g181) & (!g108) & (g123) & (g485)) + ((i_8_) & (!sk[15]) & (g181) & (g108) & (!g123) & (!g485)) + ((i_8_) & (!sk[15]) & (g181) & (g108) & (!g123) & (g485)) + ((i_8_) & (!sk[15]) & (g181) & (g108) & (g123) & (!g485)) + ((i_8_) & (!sk[15]) & (g181) & (g108) & (g123) & (g485)) + ((i_8_) & (sk[15]) & (!g181) & (g108) & (!g123) & (g485)) + ((i_8_) & (sk[15]) & (!g181) & (g108) & (g123) & (g485)) + ((i_8_) & (sk[15]) & (g181) & (g108) & (!g123) & (!g485)) + ((i_8_) & (sk[15]) & (g181) & (g108) & (!g123) & (g485)) + ((i_8_) & (sk[15]) & (g181) & (g108) & (g123) & (!g485)) + ((i_8_) & (sk[15]) & (g181) & (g108) & (g123) & (g485)));
	assign g1278 = (((!i_8_) & (!g108) & (!g670) & (!g671) & (!g1276) & (!g1277)) + ((!i_8_) & (!g108) & (!g670) & (g671) & (!g1276) & (!g1277)) + ((!i_8_) & (!g108) & (g670) & (!g671) & (!g1276) & (!g1277)) + ((!i_8_) & (!g108) & (g670) & (g671) & (!g1276) & (!g1277)) + ((!i_8_) & (g108) & (!g670) & (!g671) & (!g1276) & (!g1277)) + ((!i_8_) & (g108) & (g670) & (!g671) & (!g1276) & (!g1277)) + ((i_8_) & (!g108) & (!g670) & (!g671) & (!g1276) & (!g1277)) + ((i_8_) & (!g108) & (!g670) & (g671) & (!g1276) & (!g1277)) + ((i_8_) & (!g108) & (g670) & (!g671) & (!g1276) & (!g1277)) + ((i_8_) & (!g108) & (g670) & (g671) & (!g1276) & (!g1277)) + ((i_8_) & (g108) & (!g670) & (!g671) & (!g1276) & (!g1277)));
	assign g1279 = (((!i_8_) & (g108) & (!g216) & (!g120) & (!g123) & (!g670)) + ((!i_8_) & (g108) & (!g216) & (!g120) & (!g123) & (g670)) + ((!i_8_) & (g108) & (!g216) & (!g120) & (g123) & (!g670)) + ((!i_8_) & (g108) & (!g216) & (!g120) & (g123) & (g670)) + ((!i_8_) & (g108) & (!g216) & (g120) & (!g123) & (g670)) + ((!i_8_) & (g108) & (!g216) & (g120) & (g123) & (g670)) + ((!i_8_) & (g108) & (g216) & (!g120) & (!g123) & (!g670)) + ((!i_8_) & (g108) & (g216) & (!g120) & (!g123) & (g670)) + ((!i_8_) & (g108) & (g216) & (!g120) & (g123) & (!g670)) + ((!i_8_) & (g108) & (g216) & (!g120) & (g123) & (g670)) + ((!i_8_) & (g108) & (g216) & (g120) & (!g123) & (!g670)) + ((!i_8_) & (g108) & (g216) & (g120) & (!g123) & (g670)) + ((!i_8_) & (g108) & (g216) & (g120) & (g123) & (!g670)) + ((!i_8_) & (g108) & (g216) & (g120) & (g123) & (g670)) + ((i_8_) & (g108) & (!g216) & (!g120) & (!g123) & (!g670)) + ((i_8_) & (g108) & (!g216) & (!g120) & (!g123) & (g670)) + ((i_8_) & (g108) & (!g216) & (!g120) & (g123) & (!g670)) + ((i_8_) & (g108) & (!g216) & (!g120) & (g123) & (g670)) + ((i_8_) & (g108) & (!g216) & (g120) & (g123) & (!g670)) + ((i_8_) & (g108) & (!g216) & (g120) & (g123) & (g670)) + ((i_8_) & (g108) & (g216) & (!g120) & (!g123) & (!g670)) + ((i_8_) & (g108) & (g216) & (!g120) & (!g123) & (g670)) + ((i_8_) & (g108) & (g216) & (!g120) & (g123) & (!g670)) + ((i_8_) & (g108) & (g216) & (!g120) & (g123) & (g670)) + ((i_8_) & (g108) & (g216) & (g120) & (g123) & (!g670)) + ((i_8_) & (g108) & (g216) & (g120) & (g123) & (g670)));
	assign g1280 = (((!sk[18]) & (g108) & (!g349)) + ((!sk[18]) & (g108) & (g349)) + ((sk[18]) & (g108) & (g349)));
	assign g1281 = (((!g101) & (!g835) & (!g670) & (!g887) & (!sk[19]) & (g1280)) + ((!g101) & (!g835) & (!g670) & (!g887) & (sk[19]) & (!g1280)) + ((!g101) & (!g835) & (!g670) & (g887) & (!sk[19]) & (g1280)) + ((!g101) & (!g835) & (!g670) & (g887) & (sk[19]) & (!g1280)) + ((!g101) & (!g835) & (g670) & (!g887) & (!sk[19]) & (g1280)) + ((!g101) & (!g835) & (g670) & (!g887) & (sk[19]) & (!g1280)) + ((!g101) & (!g835) & (g670) & (g887) & (!sk[19]) & (g1280)) + ((!g101) & (!g835) & (g670) & (g887) & (sk[19]) & (!g1280)) + ((!g101) & (g835) & (!g670) & (!g887) & (!sk[19]) & (g1280)) + ((!g101) & (g835) & (!g670) & (!g887) & (sk[19]) & (!g1280)) + ((!g101) & (g835) & (!g670) & (g887) & (!sk[19]) & (g1280)) + ((!g101) & (g835) & (!g670) & (g887) & (sk[19]) & (!g1280)) + ((!g101) & (g835) & (g670) & (!g887) & (!sk[19]) & (g1280)) + ((!g101) & (g835) & (g670) & (!g887) & (sk[19]) & (!g1280)) + ((!g101) & (g835) & (g670) & (g887) & (!sk[19]) & (g1280)) + ((!g101) & (g835) & (g670) & (g887) & (sk[19]) & (!g1280)) + ((g101) & (!g835) & (!g670) & (!g887) & (!sk[19]) & (!g1280)) + ((g101) & (!g835) & (!g670) & (!g887) & (!sk[19]) & (g1280)) + ((g101) & (!g835) & (!g670) & (g887) & (!sk[19]) & (!g1280)) + ((g101) & (!g835) & (!g670) & (g887) & (!sk[19]) & (g1280)) + ((g101) & (!g835) & (g670) & (!g887) & (!sk[19]) & (!g1280)) + ((g101) & (!g835) & (g670) & (!g887) & (!sk[19]) & (g1280)) + ((g101) & (!g835) & (g670) & (g887) & (!sk[19]) & (!g1280)) + ((g101) & (!g835) & (g670) & (g887) & (!sk[19]) & (g1280)) + ((g101) & (g835) & (!g670) & (!g887) & (!sk[19]) & (!g1280)) + ((g101) & (g835) & (!g670) & (!g887) & (!sk[19]) & (g1280)) + ((g101) & (g835) & (!g670) & (g887) & (!sk[19]) & (!g1280)) + ((g101) & (g835) & (!g670) & (g887) & (!sk[19]) & (g1280)) + ((g101) & (g835) & (!g670) & (g887) & (sk[19]) & (!g1280)) + ((g101) & (g835) & (g670) & (!g887) & (!sk[19]) & (!g1280)) + ((g101) & (g835) & (g670) & (!g887) & (!sk[19]) & (g1280)) + ((g101) & (g835) & (g670) & (g887) & (!sk[19]) & (!g1280)) + ((g101) & (g835) & (g670) & (g887) & (!sk[19]) & (g1280)));
	assign g1282 = (((!i_8_) & (!g108) & (!sk[20]) & (g626) & (g895)) + ((!i_8_) & (g108) & (!sk[20]) & (!g626) & (!g895)) + ((!i_8_) & (g108) & (!sk[20]) & (!g626) & (g895)) + ((!i_8_) & (g108) & (!sk[20]) & (g626) & (!g895)) + ((!i_8_) & (g108) & (!sk[20]) & (g626) & (g895)) + ((!i_8_) & (g108) & (sk[20]) & (!g626) & (!g895)) + ((!i_8_) & (g108) & (sk[20]) & (!g626) & (g895)) + ((!i_8_) & (g108) & (sk[20]) & (g626) & (g895)) + ((i_8_) & (!g108) & (!sk[20]) & (g626) & (!g895)) + ((i_8_) & (!g108) & (!sk[20]) & (g626) & (g895)) + ((i_8_) & (g108) & (!sk[20]) & (!g626) & (!g895)) + ((i_8_) & (g108) & (!sk[20]) & (!g626) & (g895)) + ((i_8_) & (g108) & (!sk[20]) & (g626) & (!g895)) + ((i_8_) & (g108) & (!sk[20]) & (g626) & (g895)) + ((i_8_) & (g108) & (sk[20]) & (!g626) & (!g895)) + ((i_8_) & (g108) & (sk[20]) & (!g626) & (g895)));
	assign g1283 = (((g657) & (g1275) & (g1278) & (!g1279) & (g1281) & (!g1282)));
	assign g1284 = (((!i_8_) & (!g88) & (!g120) & (!sk[22]) & (!g626) & (g1048)) + ((!i_8_) & (!g88) & (!g120) & (!sk[22]) & (g626) & (g1048)) + ((!i_8_) & (!g88) & (g120) & (!sk[22]) & (!g626) & (g1048)) + ((!i_8_) & (!g88) & (g120) & (!sk[22]) & (g626) & (g1048)) + ((!i_8_) & (g88) & (!g120) & (!sk[22]) & (!g626) & (g1048)) + ((!i_8_) & (g88) & (!g120) & (!sk[22]) & (g626) & (g1048)) + ((!i_8_) & (g88) & (!g120) & (sk[22]) & (!g626) & (!g1048)) + ((!i_8_) & (g88) & (!g120) & (sk[22]) & (!g626) & (g1048)) + ((!i_8_) & (g88) & (!g120) & (sk[22]) & (g626) & (!g1048)) + ((!i_8_) & (g88) & (!g120) & (sk[22]) & (g626) & (g1048)) + ((!i_8_) & (g88) & (g120) & (!sk[22]) & (!g626) & (g1048)) + ((!i_8_) & (g88) & (g120) & (!sk[22]) & (g626) & (g1048)) + ((!i_8_) & (g88) & (g120) & (sk[22]) & (!g626) & (!g1048)) + ((!i_8_) & (g88) & (g120) & (sk[22]) & (!g626) & (g1048)) + ((!i_8_) & (g88) & (g120) & (sk[22]) & (g626) & (g1048)) + ((i_8_) & (!g88) & (!g120) & (!sk[22]) & (!g626) & (!g1048)) + ((i_8_) & (!g88) & (!g120) & (!sk[22]) & (!g626) & (g1048)) + ((i_8_) & (!g88) & (!g120) & (!sk[22]) & (g626) & (!g1048)) + ((i_8_) & (!g88) & (!g120) & (!sk[22]) & (g626) & (g1048)) + ((i_8_) & (!g88) & (g120) & (!sk[22]) & (!g626) & (!g1048)) + ((i_8_) & (!g88) & (g120) & (!sk[22]) & (!g626) & (g1048)) + ((i_8_) & (!g88) & (g120) & (!sk[22]) & (g626) & (!g1048)) + ((i_8_) & (!g88) & (g120) & (!sk[22]) & (g626) & (g1048)) + ((i_8_) & (g88) & (!g120) & (!sk[22]) & (!g626) & (!g1048)) + ((i_8_) & (g88) & (!g120) & (!sk[22]) & (!g626) & (g1048)) + ((i_8_) & (g88) & (!g120) & (!sk[22]) & (g626) & (!g1048)) + ((i_8_) & (g88) & (!g120) & (!sk[22]) & (g626) & (g1048)) + ((i_8_) & (g88) & (g120) & (!sk[22]) & (!g626) & (!g1048)) + ((i_8_) & (g88) & (g120) & (!sk[22]) & (!g626) & (g1048)) + ((i_8_) & (g88) & (g120) & (!sk[22]) & (g626) & (!g1048)) + ((i_8_) & (g88) & (g120) & (!sk[22]) & (g626) & (g1048)));
	assign g1285 = (((!g101) & (!g136) & (!sk[23]) & (!g187) & (!g670) & (g1284)) + ((!g101) & (!g136) & (!sk[23]) & (!g187) & (g670) & (g1284)) + ((!g101) & (!g136) & (!sk[23]) & (g187) & (!g670) & (g1284)) + ((!g101) & (!g136) & (!sk[23]) & (g187) & (g670) & (g1284)) + ((!g101) & (!g136) & (sk[23]) & (!g187) & (!g670) & (!g1284)) + ((!g101) & (!g136) & (sk[23]) & (!g187) & (g670) & (!g1284)) + ((!g101) & (!g136) & (sk[23]) & (g187) & (!g670) & (!g1284)) + ((!g101) & (!g136) & (sk[23]) & (g187) & (g670) & (!g1284)) + ((!g101) & (g136) & (!sk[23]) & (!g187) & (!g670) & (g1284)) + ((!g101) & (g136) & (!sk[23]) & (!g187) & (g670) & (g1284)) + ((!g101) & (g136) & (!sk[23]) & (g187) & (!g670) & (g1284)) + ((!g101) & (g136) & (!sk[23]) & (g187) & (g670) & (g1284)) + ((!g101) & (g136) & (sk[23]) & (!g187) & (!g670) & (!g1284)) + ((!g101) & (g136) & (sk[23]) & (g187) & (!g670) & (!g1284)) + ((g101) & (!g136) & (!sk[23]) & (!g187) & (!g670) & (!g1284)) + ((g101) & (!g136) & (!sk[23]) & (!g187) & (!g670) & (g1284)) + ((g101) & (!g136) & (!sk[23]) & (!g187) & (g670) & (!g1284)) + ((g101) & (!g136) & (!sk[23]) & (!g187) & (g670) & (g1284)) + ((g101) & (!g136) & (!sk[23]) & (g187) & (!g670) & (!g1284)) + ((g101) & (!g136) & (!sk[23]) & (g187) & (!g670) & (g1284)) + ((g101) & (!g136) & (!sk[23]) & (g187) & (g670) & (!g1284)) + ((g101) & (!g136) & (!sk[23]) & (g187) & (g670) & (g1284)) + ((g101) & (!g136) & (sk[23]) & (!g187) & (!g670) & (!g1284)) + ((g101) & (!g136) & (sk[23]) & (!g187) & (g670) & (!g1284)) + ((g101) & (g136) & (!sk[23]) & (!g187) & (!g670) & (!g1284)) + ((g101) & (g136) & (!sk[23]) & (!g187) & (!g670) & (g1284)) + ((g101) & (g136) & (!sk[23]) & (!g187) & (g670) & (!g1284)) + ((g101) & (g136) & (!sk[23]) & (!g187) & (g670) & (g1284)) + ((g101) & (g136) & (!sk[23]) & (g187) & (!g670) & (!g1284)) + ((g101) & (g136) & (!sk[23]) & (g187) & (!g670) & (g1284)) + ((g101) & (g136) & (!sk[23]) & (g187) & (g670) & (!g1284)) + ((g101) & (g136) & (!sk[23]) & (g187) & (g670) & (g1284)) + ((g101) & (g136) & (sk[23]) & (!g187) & (!g670) & (!g1284)));
	assign g1286 = (((!i_14_) & (i_12_) & (i_13_) & (g149) & (!g119) & (!g122)) + ((!i_14_) & (i_12_) & (i_13_) & (g149) & (g119) & (!g122)) + ((!i_14_) & (i_12_) & (i_13_) & (g149) & (g119) & (g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (g149) & (!g119) & (!g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (g149) & (g119) & (!g122)) + ((i_14_) & (!i_12_) & (i_13_) & (g149) & (!g119) & (!g122)) + ((i_14_) & (!i_12_) & (i_13_) & (g149) & (g119) & (!g122)) + ((i_14_) & (i_12_) & (!i_13_) & (g149) & (!g119) & (!g122)) + ((i_14_) & (i_12_) & (!i_13_) & (g149) & (g119) & (!g122)) + ((i_14_) & (i_12_) & (i_13_) & (g149) & (!g119) & (!g122)) + ((i_14_) & (i_12_) & (i_13_) & (g149) & (g119) & (!g122)) + ((i_14_) & (i_12_) & (i_13_) & (g149) & (g119) & (g122)));
	assign g1287 = (((!g277) & (!g214) & (g613) & (!g540) & (!g895) & (!g1286)) + ((!g277) & (g214) & (g613) & (!g540) & (!g895) & (!g1286)) + ((g277) & (!g214) & (!g613) & (!g540) & (!g895) & (!g1286)) + ((g277) & (!g214) & (!g613) & (!g540) & (g895) & (!g1286)) + ((g277) & (!g214) & (!g613) & (g540) & (!g895) & (!g1286)) + ((g277) & (!g214) & (!g613) & (g540) & (g895) & (!g1286)) + ((g277) & (!g214) & (g613) & (!g540) & (!g895) & (!g1286)) + ((g277) & (!g214) & (g613) & (!g540) & (g895) & (!g1286)) + ((g277) & (!g214) & (g613) & (g540) & (!g895) & (!g1286)) + ((g277) & (!g214) & (g613) & (g540) & (g895) & (!g1286)) + ((g277) & (g214) & (!g613) & (!g540) & (!g895) & (!g1286)) + ((g277) & (g214) & (g613) & (!g540) & (!g895) & (!g1286)));
	assign g1288 = (((!g988) & (sk[26]) & (!g1022)) + ((g988) & (!sk[26]) & (!g1022)) + ((g988) & (!sk[26]) & (g1022)));
	assign g1289 = (((!sk[27]) & (i_8_) & (!g108) & (!g895)) + ((!sk[27]) & (i_8_) & (!g108) & (g895)) + ((!sk[27]) & (i_8_) & (g108) & (!g895)) + ((!sk[27]) & (i_8_) & (g108) & (g895)) + ((sk[27]) & (i_8_) & (g108) & (g895)));
	assign g1290 = (((!sk[28]) & (g134) & (!g1161)) + ((!sk[28]) & (g134) & (g1161)) + ((sk[28]) & (g134) & (!g1161)));
	assign g1291 = (((!g183) & (sk[29]) & (g423) & (g704)) + ((g183) & (!sk[29]) & (!g423) & (!g704)) + ((g183) & (!sk[29]) & (!g423) & (g704)) + ((g183) & (!sk[29]) & (g423) & (!g704)) + ((g183) & (!sk[29]) & (g423) & (g704)) + ((g183) & (sk[29]) & (g423) & (!g704)) + ((g183) & (sk[29]) & (g423) & (g704)));
	assign g1292 = (((!g134) & (g118) & (sk[30]) & (g548)) + ((g134) & (!g118) & (!sk[30]) & (!g548)) + ((g134) & (!g118) & (!sk[30]) & (g548)) + ((g134) & (!g118) & (sk[30]) & (g548)) + ((g134) & (g118) & (!sk[30]) & (!g548)) + ((g134) & (g118) & (!sk[30]) & (g548)) + ((g134) & (g118) & (sk[30]) & (g548)));
	assign g1293 = (((!sk[31]) & (!g112) & (!g323) & (g349) & (g481)) + ((!sk[31]) & (!g112) & (g323) & (!g349) & (!g481)) + ((!sk[31]) & (!g112) & (g323) & (!g349) & (g481)) + ((!sk[31]) & (!g112) & (g323) & (g349) & (!g481)) + ((!sk[31]) & (!g112) & (g323) & (g349) & (g481)) + ((!sk[31]) & (g112) & (!g323) & (g349) & (!g481)) + ((!sk[31]) & (g112) & (!g323) & (g349) & (g481)) + ((!sk[31]) & (g112) & (g323) & (!g349) & (!g481)) + ((!sk[31]) & (g112) & (g323) & (!g349) & (g481)) + ((!sk[31]) & (g112) & (g323) & (g349) & (!g481)) + ((!sk[31]) & (g112) & (g323) & (g349) & (g481)) + ((sk[31]) & (!g112) & (!g323) & (!g349) & (!g481)) + ((sk[31]) & (!g112) & (!g323) & (!g349) & (g481)) + ((sk[31]) & (!g112) & (!g323) & (g349) & (!g481)) + ((sk[31]) & (!g112) & (!g323) & (g349) & (g481)) + ((sk[31]) & (!g112) & (g323) & (!g349) & (g481)) + ((sk[31]) & (g112) & (!g323) & (!g349) & (g481)) + ((sk[31]) & (g112) & (!g323) & (g349) & (g481)) + ((sk[31]) & (g112) & (g323) & (!g349) & (g481)));
	assign g1294 = (((g491) & (!g1289) & (!g1290) & (!g1291) & (!g1292) & (g1293)));
	assign g1295 = (((!g1150) & (g1129) & (g1285) & (g1287) & (g1288) & (g1294)));
	assign g1296 = (((!g112) & (!g349) & (!g540) & (!sk[34]) & (!g704) & (g895)) + ((!g112) & (!g349) & (!g540) & (!sk[34]) & (g704) & (g895)) + ((!g112) & (!g349) & (g540) & (!sk[34]) & (!g704) & (g895)) + ((!g112) & (!g349) & (g540) & (!sk[34]) & (g704) & (g895)) + ((!g112) & (g349) & (!g540) & (!sk[34]) & (!g704) & (g895)) + ((!g112) & (g349) & (!g540) & (!sk[34]) & (g704) & (g895)) + ((!g112) & (g349) & (g540) & (!sk[34]) & (!g704) & (g895)) + ((!g112) & (g349) & (g540) & (!sk[34]) & (g704) & (g895)) + ((g112) & (!g349) & (!g540) & (!sk[34]) & (!g704) & (!g895)) + ((g112) & (!g349) & (!g540) & (!sk[34]) & (!g704) & (g895)) + ((g112) & (!g349) & (!g540) & (!sk[34]) & (g704) & (!g895)) + ((g112) & (!g349) & (!g540) & (!sk[34]) & (g704) & (g895)) + ((g112) & (!g349) & (!g540) & (sk[34]) & (!g704) & (g895)) + ((g112) & (!g349) & (!g540) & (sk[34]) & (g704) & (!g895)) + ((g112) & (!g349) & (!g540) & (sk[34]) & (g704) & (g895)) + ((g112) & (!g349) & (g540) & (!sk[34]) & (!g704) & (!g895)) + ((g112) & (!g349) & (g540) & (!sk[34]) & (!g704) & (g895)) + ((g112) & (!g349) & (g540) & (!sk[34]) & (g704) & (!g895)) + ((g112) & (!g349) & (g540) & (!sk[34]) & (g704) & (g895)) + ((g112) & (!g349) & (g540) & (sk[34]) & (!g704) & (!g895)) + ((g112) & (!g349) & (g540) & (sk[34]) & (!g704) & (g895)) + ((g112) & (!g349) & (g540) & (sk[34]) & (g704) & (!g895)) + ((g112) & (!g349) & (g540) & (sk[34]) & (g704) & (g895)) + ((g112) & (g349) & (!g540) & (!sk[34]) & (!g704) & (!g895)) + ((g112) & (g349) & (!g540) & (!sk[34]) & (!g704) & (g895)) + ((g112) & (g349) & (!g540) & (!sk[34]) & (g704) & (!g895)) + ((g112) & (g349) & (!g540) & (!sk[34]) & (g704) & (g895)) + ((g112) & (g349) & (!g540) & (sk[34]) & (!g704) & (!g895)) + ((g112) & (g349) & (!g540) & (sk[34]) & (!g704) & (g895)) + ((g112) & (g349) & (!g540) & (sk[34]) & (g704) & (!g895)) + ((g112) & (g349) & (!g540) & (sk[34]) & (g704) & (g895)) + ((g112) & (g349) & (g540) & (!sk[34]) & (!g704) & (!g895)) + ((g112) & (g349) & (g540) & (!sk[34]) & (!g704) & (g895)) + ((g112) & (g349) & (g540) & (!sk[34]) & (g704) & (!g895)) + ((g112) & (g349) & (g540) & (!sk[34]) & (g704) & (g895)) + ((g112) & (g349) & (g540) & (sk[34]) & (!g704) & (!g895)) + ((g112) & (g349) & (g540) & (sk[34]) & (!g704) & (g895)) + ((g112) & (g349) & (g540) & (sk[34]) & (g704) & (!g895)) + ((g112) & (g349) & (g540) & (sk[34]) & (g704) & (g895)));
	assign g1297 = (((!sk[35]) & (!g134) & (!g136) & (!g120) & (!g123) & (g1296)) + ((!sk[35]) & (!g134) & (!g136) & (!g120) & (g123) & (g1296)) + ((!sk[35]) & (!g134) & (!g136) & (g120) & (!g123) & (g1296)) + ((!sk[35]) & (!g134) & (!g136) & (g120) & (g123) & (g1296)) + ((!sk[35]) & (!g134) & (g136) & (!g120) & (!g123) & (g1296)) + ((!sk[35]) & (!g134) & (g136) & (!g120) & (g123) & (g1296)) + ((!sk[35]) & (!g134) & (g136) & (g120) & (!g123) & (g1296)) + ((!sk[35]) & (!g134) & (g136) & (g120) & (g123) & (g1296)) + ((!sk[35]) & (g134) & (!g136) & (!g120) & (!g123) & (!g1296)) + ((!sk[35]) & (g134) & (!g136) & (!g120) & (!g123) & (g1296)) + ((!sk[35]) & (g134) & (!g136) & (!g120) & (g123) & (!g1296)) + ((!sk[35]) & (g134) & (!g136) & (!g120) & (g123) & (g1296)) + ((!sk[35]) & (g134) & (!g136) & (g120) & (!g123) & (!g1296)) + ((!sk[35]) & (g134) & (!g136) & (g120) & (!g123) & (g1296)) + ((!sk[35]) & (g134) & (!g136) & (g120) & (g123) & (!g1296)) + ((!sk[35]) & (g134) & (!g136) & (g120) & (g123) & (g1296)) + ((!sk[35]) & (g134) & (g136) & (!g120) & (!g123) & (!g1296)) + ((!sk[35]) & (g134) & (g136) & (!g120) & (!g123) & (g1296)) + ((!sk[35]) & (g134) & (g136) & (!g120) & (g123) & (!g1296)) + ((!sk[35]) & (g134) & (g136) & (!g120) & (g123) & (g1296)) + ((!sk[35]) & (g134) & (g136) & (g120) & (!g123) & (!g1296)) + ((!sk[35]) & (g134) & (g136) & (g120) & (!g123) & (g1296)) + ((!sk[35]) & (g134) & (g136) & (g120) & (g123) & (!g1296)) + ((!sk[35]) & (g134) & (g136) & (g120) & (g123) & (g1296)) + ((sk[35]) & (!g134) & (!g136) & (!g120) & (!g123) & (!g1296)) + ((sk[35]) & (!g134) & (!g136) & (!g120) & (g123) & (!g1296)) + ((sk[35]) & (!g134) & (!g136) & (g120) & (!g123) & (!g1296)) + ((sk[35]) & (!g134) & (!g136) & (g120) & (g123) & (!g1296)) + ((sk[35]) & (!g134) & (g136) & (g120) & (!g123) & (!g1296)) + ((sk[35]) & (!g134) & (g136) & (g120) & (g123) & (!g1296)) + ((sk[35]) & (g134) & (!g136) & (!g120) & (!g123) & (!g1296)) + ((sk[35]) & (g134) & (!g136) & (g120) & (!g123) & (!g1296)) + ((sk[35]) & (g134) & (g136) & (g120) & (!g123) & (!g1296)));
	assign g1298 = (((g136) & (!sk[36]) & (!g349) & (!g540)) + ((g136) & (!sk[36]) & (!g349) & (g540)) + ((g136) & (!sk[36]) & (g349) & (!g540)) + ((g136) & (!sk[36]) & (g349) & (g540)) + ((g136) & (sk[36]) & (!g349) & (g540)) + ((g136) & (sk[36]) & (g349) & (!g540)) + ((g136) & (sk[36]) & (g349) & (g540)));
	assign g1299 = (((!i_14_) & (!i_12_) & (!i_13_) & (!g119) & (g136) & (!g122)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g119) & (g136) & (!g122)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g119) & (g136) & (g122)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g119) & (g136) & (!g122)) + ((!i_14_) & (i_12_) & (!i_13_) & (g119) & (g136) & (!g122)) + ((!i_14_) & (i_12_) & (!i_13_) & (g119) & (g136) & (g122)) + ((!i_14_) & (i_12_) & (i_13_) & (!g119) & (g136) & (!g122)) + ((!i_14_) & (i_12_) & (i_13_) & (g119) & (g136) & (!g122)) + ((!i_14_) & (i_12_) & (i_13_) & (g119) & (g136) & (g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (!g119) & (g136) & (!g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (g119) & (g136) & (!g122)) + ((i_14_) & (!i_12_) & (!i_13_) & (g119) & (g136) & (g122)) + ((i_14_) & (i_12_) & (i_13_) & (g119) & (g136) & (!g122)) + ((i_14_) & (i_12_) & (i_13_) & (g119) & (g136) & (g122)));
	assign g1300 = (((!sk[38]) & (!g760) & (!g1297) & (!g1298) & (!g1596) & (g1299)) + ((!sk[38]) & (!g760) & (!g1297) & (!g1298) & (g1596) & (g1299)) + ((!sk[38]) & (!g760) & (!g1297) & (g1298) & (!g1596) & (g1299)) + ((!sk[38]) & (!g760) & (!g1297) & (g1298) & (g1596) & (g1299)) + ((!sk[38]) & (!g760) & (g1297) & (!g1298) & (!g1596) & (g1299)) + ((!sk[38]) & (!g760) & (g1297) & (!g1298) & (g1596) & (g1299)) + ((!sk[38]) & (!g760) & (g1297) & (g1298) & (!g1596) & (g1299)) + ((!sk[38]) & (!g760) & (g1297) & (g1298) & (g1596) & (g1299)) + ((!sk[38]) & (g760) & (!g1297) & (!g1298) & (!g1596) & (!g1299)) + ((!sk[38]) & (g760) & (!g1297) & (!g1298) & (!g1596) & (g1299)) + ((!sk[38]) & (g760) & (!g1297) & (!g1298) & (g1596) & (!g1299)) + ((!sk[38]) & (g760) & (!g1297) & (!g1298) & (g1596) & (g1299)) + ((!sk[38]) & (g760) & (!g1297) & (g1298) & (!g1596) & (!g1299)) + ((!sk[38]) & (g760) & (!g1297) & (g1298) & (!g1596) & (g1299)) + ((!sk[38]) & (g760) & (!g1297) & (g1298) & (g1596) & (!g1299)) + ((!sk[38]) & (g760) & (!g1297) & (g1298) & (g1596) & (g1299)) + ((!sk[38]) & (g760) & (g1297) & (!g1298) & (!g1596) & (!g1299)) + ((!sk[38]) & (g760) & (g1297) & (!g1298) & (!g1596) & (g1299)) + ((!sk[38]) & (g760) & (g1297) & (!g1298) & (g1596) & (!g1299)) + ((!sk[38]) & (g760) & (g1297) & (!g1298) & (g1596) & (g1299)) + ((!sk[38]) & (g760) & (g1297) & (g1298) & (!g1596) & (!g1299)) + ((!sk[38]) & (g760) & (g1297) & (g1298) & (!g1596) & (g1299)) + ((!sk[38]) & (g760) & (g1297) & (g1298) & (g1596) & (!g1299)) + ((!sk[38]) & (g760) & (g1297) & (g1298) & (g1596) & (g1299)) + ((sk[38]) & (!g760) & (g1297) & (!g1298) & (g1596) & (!g1299)));
	assign g1301 = (((g1259) & (g1265) & (g1273) & (g1283) & (g1295) & (g1300)));
	assign o_17_ = (((g73) & (!g1156) & (!g1195) & (!g1221) & (!g1258) & (!g1301)) + ((g73) & (!g1156) & (!g1195) & (!g1221) & (!g1258) & (g1301)) + ((g73) & (!g1156) & (!g1195) & (!g1221) & (g1258) & (!g1301)) + ((g73) & (!g1156) & (!g1195) & (!g1221) & (g1258) & (g1301)) + ((g73) & (!g1156) & (!g1195) & (g1221) & (!g1258) & (!g1301)) + ((g73) & (!g1156) & (!g1195) & (g1221) & (!g1258) & (g1301)) + ((g73) & (!g1156) & (!g1195) & (g1221) & (g1258) & (!g1301)) + ((g73) & (!g1156) & (!g1195) & (g1221) & (g1258) & (g1301)) + ((g73) & (!g1156) & (g1195) & (!g1221) & (!g1258) & (!g1301)) + ((g73) & (!g1156) & (g1195) & (!g1221) & (!g1258) & (g1301)) + ((g73) & (!g1156) & (g1195) & (!g1221) & (g1258) & (!g1301)) + ((g73) & (!g1156) & (g1195) & (!g1221) & (g1258) & (g1301)) + ((g73) & (!g1156) & (g1195) & (g1221) & (!g1258) & (!g1301)) + ((g73) & (!g1156) & (g1195) & (g1221) & (!g1258) & (g1301)) + ((g73) & (!g1156) & (g1195) & (g1221) & (g1258) & (!g1301)) + ((g73) & (!g1156) & (g1195) & (g1221) & (g1258) & (g1301)) + ((g73) & (g1156) & (!g1195) & (!g1221) & (!g1258) & (!g1301)) + ((g73) & (g1156) & (!g1195) & (!g1221) & (!g1258) & (g1301)) + ((g73) & (g1156) & (!g1195) & (!g1221) & (g1258) & (!g1301)) + ((g73) & (g1156) & (!g1195) & (!g1221) & (g1258) & (g1301)) + ((g73) & (g1156) & (!g1195) & (g1221) & (!g1258) & (!g1301)) + ((g73) & (g1156) & (!g1195) & (g1221) & (!g1258) & (g1301)) + ((g73) & (g1156) & (!g1195) & (g1221) & (g1258) & (!g1301)) + ((g73) & (g1156) & (!g1195) & (g1221) & (g1258) & (g1301)) + ((g73) & (g1156) & (g1195) & (!g1221) & (!g1258) & (!g1301)) + ((g73) & (g1156) & (g1195) & (!g1221) & (!g1258) & (g1301)) + ((g73) & (g1156) & (g1195) & (!g1221) & (g1258) & (!g1301)) + ((g73) & (g1156) & (g1195) & (!g1221) & (g1258) & (g1301)) + ((g73) & (g1156) & (g1195) & (g1221) & (!g1258) & (!g1301)) + ((g73) & (g1156) & (g1195) & (g1221) & (!g1258) & (g1301)) + ((g73) & (g1156) & (g1195) & (g1221) & (g1258) & (!g1301)));
	assign g1303 = (((g1265) & (!sk[41]) & (!g1273)) + ((g1265) & (!sk[41]) & (g1273)) + ((g1265) & (sk[41]) & (g1273)));
	assign g1304 = (((!i_14_) & (!i_12_) & (!sk[42]) & (!i_13_) & (!g102) & (g115)) + ((!i_14_) & (!i_12_) & (!sk[42]) & (!i_13_) & (g102) & (g115)) + ((!i_14_) & (!i_12_) & (!sk[42]) & (i_13_) & (!g102) & (g115)) + ((!i_14_) & (!i_12_) & (!sk[42]) & (i_13_) & (g102) & (g115)) + ((!i_14_) & (!i_12_) & (sk[42]) & (i_13_) & (!g102) & (!g115)) + ((!i_14_) & (!i_12_) & (sk[42]) & (i_13_) & (!g102) & (g115)) + ((!i_14_) & (i_12_) & (!sk[42]) & (!i_13_) & (!g102) & (g115)) + ((!i_14_) & (i_12_) & (!sk[42]) & (!i_13_) & (g102) & (g115)) + ((!i_14_) & (i_12_) & (!sk[42]) & (i_13_) & (!g102) & (g115)) + ((!i_14_) & (i_12_) & (!sk[42]) & (i_13_) & (g102) & (g115)) + ((!i_14_) & (i_12_) & (sk[42]) & (!i_13_) & (!g102) & (!g115)) + ((!i_14_) & (i_12_) & (sk[42]) & (!i_13_) & (!g102) & (g115)) + ((!i_14_) & (i_12_) & (sk[42]) & (!i_13_) & (g102) & (!g115)) + ((!i_14_) & (i_12_) & (sk[42]) & (i_13_) & (!g102) & (!g115)) + ((!i_14_) & (i_12_) & (sk[42]) & (i_13_) & (!g102) & (g115)) + ((i_14_) & (!i_12_) & (!sk[42]) & (!i_13_) & (!g102) & (!g115)) + ((i_14_) & (!i_12_) & (!sk[42]) & (!i_13_) & (!g102) & (g115)) + ((i_14_) & (!i_12_) & (!sk[42]) & (!i_13_) & (g102) & (!g115)) + ((i_14_) & (!i_12_) & (!sk[42]) & (!i_13_) & (g102) & (g115)) + ((i_14_) & (!i_12_) & (!sk[42]) & (i_13_) & (!g102) & (!g115)) + ((i_14_) & (!i_12_) & (!sk[42]) & (i_13_) & (!g102) & (g115)) + ((i_14_) & (!i_12_) & (!sk[42]) & (i_13_) & (g102) & (!g115)) + ((i_14_) & (!i_12_) & (!sk[42]) & (i_13_) & (g102) & (g115)) + ((i_14_) & (!i_12_) & (sk[42]) & (!i_13_) & (!g102) & (!g115)) + ((i_14_) & (!i_12_) & (sk[42]) & (!i_13_) & (!g102) & (g115)) + ((i_14_) & (!i_12_) & (sk[42]) & (i_13_) & (!g102) & (!g115)) + ((i_14_) & (!i_12_) & (sk[42]) & (i_13_) & (!g102) & (g115)) + ((i_14_) & (!i_12_) & (sk[42]) & (i_13_) & (g102) & (!g115)) + ((i_14_) & (i_12_) & (!sk[42]) & (!i_13_) & (!g102) & (!g115)) + ((i_14_) & (i_12_) & (!sk[42]) & (!i_13_) & (!g102) & (g115)) + ((i_14_) & (i_12_) & (!sk[42]) & (!i_13_) & (g102) & (!g115)) + ((i_14_) & (i_12_) & (!sk[42]) & (!i_13_) & (g102) & (g115)) + ((i_14_) & (i_12_) & (!sk[42]) & (i_13_) & (!g102) & (!g115)) + ((i_14_) & (i_12_) & (!sk[42]) & (i_13_) & (!g102) & (g115)) + ((i_14_) & (i_12_) & (!sk[42]) & (i_13_) & (g102) & (!g115)) + ((i_14_) & (i_12_) & (!sk[42]) & (i_13_) & (g102) & (g115)) + ((i_14_) & (i_12_) & (sk[42]) & (!i_13_) & (!g102) & (!g115)) + ((i_14_) & (i_12_) & (sk[42]) & (!i_13_) & (g102) & (!g115)));
	assign g1305 = (((!g118) & (!g187) & (!g534) & (!g980) & (!sk[43]) & (g1304)) + ((!g118) & (!g187) & (!g534) & (g980) & (!sk[43]) & (g1304)) + ((!g118) & (!g187) & (g534) & (!g980) & (!sk[43]) & (g1304)) + ((!g118) & (!g187) & (g534) & (g980) & (!sk[43]) & (g1304)) + ((!g118) & (g187) & (!g534) & (!g980) & (!sk[43]) & (g1304)) + ((!g118) & (g187) & (!g534) & (g980) & (!sk[43]) & (g1304)) + ((!g118) & (g187) & (g534) & (!g980) & (!sk[43]) & (g1304)) + ((!g118) & (g187) & (g534) & (g980) & (!sk[43]) & (g1304)) + ((g118) & (!g187) & (!g534) & (!g980) & (!sk[43]) & (!g1304)) + ((g118) & (!g187) & (!g534) & (!g980) & (!sk[43]) & (g1304)) + ((g118) & (!g187) & (!g534) & (!g980) & (sk[43]) & (!g1304)) + ((g118) & (!g187) & (!g534) & (!g980) & (sk[43]) & (g1304)) + ((g118) & (!g187) & (!g534) & (g980) & (!sk[43]) & (!g1304)) + ((g118) & (!g187) & (!g534) & (g980) & (!sk[43]) & (g1304)) + ((g118) & (!g187) & (!g534) & (g980) & (sk[43]) & (g1304)) + ((g118) & (!g187) & (g534) & (!g980) & (!sk[43]) & (!g1304)) + ((g118) & (!g187) & (g534) & (!g980) & (!sk[43]) & (g1304)) + ((g118) & (!g187) & (g534) & (!g980) & (sk[43]) & (!g1304)) + ((g118) & (!g187) & (g534) & (!g980) & (sk[43]) & (g1304)) + ((g118) & (!g187) & (g534) & (g980) & (!sk[43]) & (!g1304)) + ((g118) & (!g187) & (g534) & (g980) & (!sk[43]) & (g1304)) + ((g118) & (!g187) & (g534) & (g980) & (sk[43]) & (!g1304)) + ((g118) & (!g187) & (g534) & (g980) & (sk[43]) & (g1304)) + ((g118) & (g187) & (!g534) & (!g980) & (!sk[43]) & (!g1304)) + ((g118) & (g187) & (!g534) & (!g980) & (!sk[43]) & (g1304)) + ((g118) & (g187) & (!g534) & (!g980) & (sk[43]) & (!g1304)) + ((g118) & (g187) & (!g534) & (!g980) & (sk[43]) & (g1304)) + ((g118) & (g187) & (!g534) & (g980) & (!sk[43]) & (!g1304)) + ((g118) & (g187) & (!g534) & (g980) & (!sk[43]) & (g1304)) + ((g118) & (g187) & (!g534) & (g980) & (sk[43]) & (!g1304)) + ((g118) & (g187) & (!g534) & (g980) & (sk[43]) & (g1304)) + ((g118) & (g187) & (g534) & (!g980) & (!sk[43]) & (!g1304)) + ((g118) & (g187) & (g534) & (!g980) & (!sk[43]) & (g1304)) + ((g118) & (g187) & (g534) & (!g980) & (sk[43]) & (!g1304)) + ((g118) & (g187) & (g534) & (!g980) & (sk[43]) & (g1304)) + ((g118) & (g187) & (g534) & (g980) & (!sk[43]) & (!g1304)) + ((g118) & (g187) & (g534) & (g980) & (!sk[43]) & (g1304)) + ((g118) & (g187) & (g534) & (g980) & (sk[43]) & (!g1304)) + ((g118) & (g187) & (g534) & (g980) & (sk[43]) & (g1304)));
	assign g1306 = (((!g546) & (!g477) & (!sk[44]) & (g706) & (g979)) + ((!g546) & (g477) & (!sk[44]) & (!g706) & (!g979)) + ((!g546) & (g477) & (!sk[44]) & (!g706) & (g979)) + ((!g546) & (g477) & (!sk[44]) & (g706) & (!g979)) + ((!g546) & (g477) & (!sk[44]) & (g706) & (g979)) + ((!g546) & (g477) & (sk[44]) & (!g706) & (g979)) + ((g546) & (!g477) & (!sk[44]) & (g706) & (!g979)) + ((g546) & (!g477) & (!sk[44]) & (g706) & (g979)) + ((g546) & (g477) & (!sk[44]) & (!g706) & (!g979)) + ((g546) & (g477) & (!sk[44]) & (!g706) & (g979)) + ((g546) & (g477) & (!sk[44]) & (g706) & (!g979)) + ((g546) & (g477) & (!sk[44]) & (g706) & (g979)));
	assign g1307 = (((!g109) & (!g1179) & (!sk[45]) & (g1243) & (g1306)) + ((!g109) & (!g1179) & (sk[45]) & (!g1243) & (!g1306)) + ((!g109) & (!g1179) & (sk[45]) & (!g1243) & (g1306)) + ((!g109) & (g1179) & (!sk[45]) & (!g1243) & (!g1306)) + ((!g109) & (g1179) & (!sk[45]) & (!g1243) & (g1306)) + ((!g109) & (g1179) & (!sk[45]) & (g1243) & (!g1306)) + ((!g109) & (g1179) & (!sk[45]) & (g1243) & (g1306)) + ((g109) & (!g1179) & (!sk[45]) & (g1243) & (!g1306)) + ((g109) & (!g1179) & (!sk[45]) & (g1243) & (g1306)) + ((g109) & (!g1179) & (sk[45]) & (!g1243) & (g1306)) + ((g109) & (g1179) & (!sk[45]) & (!g1243) & (!g1306)) + ((g109) & (g1179) & (!sk[45]) & (!g1243) & (g1306)) + ((g109) & (g1179) & (!sk[45]) & (g1243) & (!g1306)) + ((g109) & (g1179) & (!sk[45]) & (g1243) & (g1306)));
	assign g1308 = (((!i_8_) & (g108) & (!g193) & (!g232) & (!g173) & (!g103)) + ((!i_8_) & (g108) & (!g193) & (!g232) & (g173) & (!g103)) + ((!i_8_) & (g108) & (!g193) & (!g232) & (g173) & (g103)) + ((!i_8_) & (g108) & (!g193) & (g232) & (!g173) & (!g103)) + ((!i_8_) & (g108) & (!g193) & (g232) & (!g173) & (g103)) + ((!i_8_) & (g108) & (!g193) & (g232) & (g173) & (!g103)) + ((!i_8_) & (g108) & (!g193) & (g232) & (g173) & (g103)) + ((!i_8_) & (g108) & (g193) & (!g232) & (!g173) & (!g103)) + ((!i_8_) & (g108) & (g193) & (!g232) & (!g173) & (g103)) + ((!i_8_) & (g108) & (g193) & (!g232) & (g173) & (!g103)) + ((!i_8_) & (g108) & (g193) & (!g232) & (g173) & (g103)) + ((!i_8_) & (g108) & (g193) & (g232) & (!g173) & (!g103)) + ((!i_8_) & (g108) & (g193) & (g232) & (!g173) & (g103)) + ((!i_8_) & (g108) & (g193) & (g232) & (g173) & (!g103)) + ((!i_8_) & (g108) & (g193) & (g232) & (g173) & (g103)));
	assign g1309 = (((!i_8_) & (!g264) & (!g108) & (!g696) & (!g907) & (!g1308)) + ((!i_8_) & (!g264) & (!g108) & (!g696) & (g907) & (!g1308)) + ((!i_8_) & (!g264) & (!g108) & (g696) & (!g907) & (!g1308)) + ((!i_8_) & (!g264) & (!g108) & (g696) & (g907) & (!g1308)) + ((!i_8_) & (!g264) & (g108) & (!g696) & (!g907) & (!g1308)) + ((!i_8_) & (!g264) & (g108) & (!g696) & (g907) & (!g1308)) + ((!i_8_) & (!g264) & (g108) & (g696) & (!g907) & (!g1308)) + ((!i_8_) & (!g264) & (g108) & (g696) & (g907) & (!g1308)) + ((!i_8_) & (g264) & (!g108) & (!g696) & (!g907) & (!g1308)) + ((!i_8_) & (g264) & (!g108) & (!g696) & (g907) & (!g1308)) + ((!i_8_) & (g264) & (!g108) & (g696) & (!g907) & (!g1308)) + ((!i_8_) & (g264) & (!g108) & (g696) & (g907) & (!g1308)) + ((i_8_) & (!g264) & (!g108) & (!g696) & (!g907) & (!g1308)) + ((i_8_) & (!g264) & (!g108) & (!g696) & (g907) & (!g1308)) + ((i_8_) & (!g264) & (!g108) & (g696) & (!g907) & (!g1308)) + ((i_8_) & (!g264) & (!g108) & (g696) & (g907) & (!g1308)) + ((i_8_) & (!g264) & (g108) & (g696) & (!g907) & (!g1308)) + ((i_8_) & (g264) & (!g108) & (!g696) & (!g907) & (!g1308)) + ((i_8_) & (g264) & (!g108) & (!g696) & (g907) & (!g1308)) + ((i_8_) & (g264) & (!g108) & (g696) & (!g907) & (!g1308)) + ((i_8_) & (g264) & (!g108) & (g696) & (g907) & (!g1308)) + ((i_8_) & (g264) & (g108) & (g696) & (!g907) & (!g1308)));
	assign g1310 = (((!g220) & (sk[48]) & (g112) & (!g827)) + ((g220) & (!sk[48]) & (!g112) & (!g827)) + ((g220) & (!sk[48]) & (!g112) & (g827)) + ((g220) & (!sk[48]) & (g112) & (!g827)) + ((g220) & (!sk[48]) & (g112) & (g827)) + ((g220) & (sk[48]) & (g112) & (!g827)) + ((g220) & (sk[48]) & (g112) & (g827)));
	assign g1311 = (((!g48) & (!sk[49]) & (!g102) & (!g112) & (!g182) & (g115)) + ((!g48) & (!sk[49]) & (!g102) & (!g112) & (g182) & (g115)) + ((!g48) & (!sk[49]) & (!g102) & (g112) & (!g182) & (g115)) + ((!g48) & (!sk[49]) & (!g102) & (g112) & (g182) & (g115)) + ((!g48) & (!sk[49]) & (g102) & (!g112) & (!g182) & (g115)) + ((!g48) & (!sk[49]) & (g102) & (!g112) & (g182) & (g115)) + ((!g48) & (!sk[49]) & (g102) & (g112) & (!g182) & (g115)) + ((!g48) & (!sk[49]) & (g102) & (g112) & (g182) & (g115)) + ((!g48) & (sk[49]) & (!g102) & (g112) & (!g182) & (!g115)) + ((!g48) & (sk[49]) & (!g102) & (g112) & (!g182) & (g115)) + ((!g48) & (sk[49]) & (!g102) & (g112) & (g182) & (!g115)) + ((!g48) & (sk[49]) & (!g102) & (g112) & (g182) & (g115)) + ((!g48) & (sk[49]) & (g102) & (g112) & (!g182) & (!g115)) + ((!g48) & (sk[49]) & (g102) & (g112) & (g182) & (!g115)) + ((g48) & (!sk[49]) & (!g102) & (!g112) & (!g182) & (!g115)) + ((g48) & (!sk[49]) & (!g102) & (!g112) & (!g182) & (g115)) + ((g48) & (!sk[49]) & (!g102) & (!g112) & (g182) & (!g115)) + ((g48) & (!sk[49]) & (!g102) & (!g112) & (g182) & (g115)) + ((g48) & (!sk[49]) & (!g102) & (g112) & (!g182) & (!g115)) + ((g48) & (!sk[49]) & (!g102) & (g112) & (!g182) & (g115)) + ((g48) & (!sk[49]) & (!g102) & (g112) & (g182) & (!g115)) + ((g48) & (!sk[49]) & (!g102) & (g112) & (g182) & (g115)) + ((g48) & (!sk[49]) & (g102) & (!g112) & (!g182) & (!g115)) + ((g48) & (!sk[49]) & (g102) & (!g112) & (!g182) & (g115)) + ((g48) & (!sk[49]) & (g102) & (!g112) & (g182) & (!g115)) + ((g48) & (!sk[49]) & (g102) & (!g112) & (g182) & (g115)) + ((g48) & (!sk[49]) & (g102) & (g112) & (!g182) & (!g115)) + ((g48) & (!sk[49]) & (g102) & (g112) & (!g182) & (g115)) + ((g48) & (!sk[49]) & (g102) & (g112) & (g182) & (!g115)) + ((g48) & (!sk[49]) & (g102) & (g112) & (g182) & (g115)) + ((g48) & (sk[49]) & (!g102) & (g112) & (g182) & (!g115)) + ((g48) & (sk[49]) & (!g102) & (g112) & (g182) & (g115)) + ((g48) & (sk[49]) & (g102) & (g112) & (g182) & (!g115)));
	assign g1312 = (((!g112) & (!sk[50]) & (!g675) & (g672) & (g706)) + ((!g112) & (!sk[50]) & (g675) & (!g672) & (!g706)) + ((!g112) & (!sk[50]) & (g675) & (!g672) & (g706)) + ((!g112) & (!sk[50]) & (g675) & (g672) & (!g706)) + ((!g112) & (!sk[50]) & (g675) & (g672) & (g706)) + ((g112) & (!sk[50]) & (!g675) & (g672) & (!g706)) + ((g112) & (!sk[50]) & (!g675) & (g672) & (g706)) + ((g112) & (!sk[50]) & (g675) & (!g672) & (!g706)) + ((g112) & (!sk[50]) & (g675) & (!g672) & (g706)) + ((g112) & (!sk[50]) & (g675) & (g672) & (!g706)) + ((g112) & (!sk[50]) & (g675) & (g672) & (g706)) + ((g112) & (sk[50]) & (!g675) & (!g672) & (g706)) + ((g112) & (sk[50]) & (!g675) & (g672) & (!g706)) + ((g112) & (sk[50]) & (!g675) & (g672) & (g706)) + ((g112) & (sk[50]) & (g675) & (!g672) & (!g706)) + ((g112) & (sk[50]) & (g675) & (!g672) & (g706)) + ((g112) & (sk[50]) & (g675) & (g672) & (!g706)) + ((g112) & (sk[50]) & (g675) & (g672) & (g706)));
	assign g1313 = (((!sk[51]) & (!g118) & (!g231) & (!g478) & (!g487) & (g675)) + ((!sk[51]) & (!g118) & (!g231) & (!g478) & (g487) & (g675)) + ((!sk[51]) & (!g118) & (!g231) & (g478) & (!g487) & (g675)) + ((!sk[51]) & (!g118) & (!g231) & (g478) & (g487) & (g675)) + ((!sk[51]) & (!g118) & (g231) & (!g478) & (!g487) & (g675)) + ((!sk[51]) & (!g118) & (g231) & (!g478) & (g487) & (g675)) + ((!sk[51]) & (!g118) & (g231) & (g478) & (!g487) & (g675)) + ((!sk[51]) & (!g118) & (g231) & (g478) & (g487) & (g675)) + ((!sk[51]) & (g118) & (!g231) & (!g478) & (!g487) & (!g675)) + ((!sk[51]) & (g118) & (!g231) & (!g478) & (!g487) & (g675)) + ((!sk[51]) & (g118) & (!g231) & (!g478) & (g487) & (!g675)) + ((!sk[51]) & (g118) & (!g231) & (!g478) & (g487) & (g675)) + ((!sk[51]) & (g118) & (!g231) & (g478) & (!g487) & (!g675)) + ((!sk[51]) & (g118) & (!g231) & (g478) & (!g487) & (g675)) + ((!sk[51]) & (g118) & (!g231) & (g478) & (g487) & (!g675)) + ((!sk[51]) & (g118) & (!g231) & (g478) & (g487) & (g675)) + ((!sk[51]) & (g118) & (g231) & (!g478) & (!g487) & (!g675)) + ((!sk[51]) & (g118) & (g231) & (!g478) & (!g487) & (g675)) + ((!sk[51]) & (g118) & (g231) & (!g478) & (g487) & (!g675)) + ((!sk[51]) & (g118) & (g231) & (!g478) & (g487) & (g675)) + ((!sk[51]) & (g118) & (g231) & (g478) & (!g487) & (!g675)) + ((!sk[51]) & (g118) & (g231) & (g478) & (!g487) & (g675)) + ((!sk[51]) & (g118) & (g231) & (g478) & (g487) & (!g675)) + ((!sk[51]) & (g118) & (g231) & (g478) & (g487) & (g675)) + ((sk[51]) & (g118) & (!g231) & (!g478) & (!g487) & (!g675)) + ((sk[51]) & (g118) & (!g231) & (!g478) & (!g487) & (g675)) + ((sk[51]) & (g118) & (!g231) & (!g478) & (g487) & (!g675)) + ((sk[51]) & (g118) & (!g231) & (!g478) & (g487) & (g675)) + ((sk[51]) & (g118) & (!g231) & (g478) & (!g487) & (!g675)) + ((sk[51]) & (g118) & (!g231) & (g478) & (!g487) & (g675)) + ((sk[51]) & (g118) & (!g231) & (g478) & (g487) & (!g675)) + ((sk[51]) & (g118) & (!g231) & (g478) & (g487) & (g675)) + ((sk[51]) & (g118) & (g231) & (!g478) & (!g487) & (g675)) + ((sk[51]) & (g118) & (g231) & (!g478) & (g487) & (!g675)) + ((sk[51]) & (g118) & (g231) & (!g478) & (g487) & (g675)) + ((sk[51]) & (g118) & (g231) & (g478) & (!g487) & (!g675)) + ((sk[51]) & (g118) & (g231) & (g478) & (!g487) & (g675)) + ((sk[51]) & (g118) & (g231) & (g478) & (g487) & (!g675)) + ((sk[51]) & (g118) & (g231) & (g478) & (g487) & (g675)));
	assign g1314 = (((!sk[52]) & (!g658) & (!g1310) & (!g1311) & (!g1312) & (g1313)) + ((!sk[52]) & (!g658) & (!g1310) & (!g1311) & (g1312) & (g1313)) + ((!sk[52]) & (!g658) & (!g1310) & (g1311) & (!g1312) & (g1313)) + ((!sk[52]) & (!g658) & (!g1310) & (g1311) & (g1312) & (g1313)) + ((!sk[52]) & (!g658) & (g1310) & (!g1311) & (!g1312) & (g1313)) + ((!sk[52]) & (!g658) & (g1310) & (!g1311) & (g1312) & (g1313)) + ((!sk[52]) & (!g658) & (g1310) & (g1311) & (!g1312) & (g1313)) + ((!sk[52]) & (!g658) & (g1310) & (g1311) & (g1312) & (g1313)) + ((!sk[52]) & (g658) & (!g1310) & (!g1311) & (!g1312) & (!g1313)) + ((!sk[52]) & (g658) & (!g1310) & (!g1311) & (!g1312) & (g1313)) + ((!sk[52]) & (g658) & (!g1310) & (!g1311) & (g1312) & (!g1313)) + ((!sk[52]) & (g658) & (!g1310) & (!g1311) & (g1312) & (g1313)) + ((!sk[52]) & (g658) & (!g1310) & (g1311) & (!g1312) & (!g1313)) + ((!sk[52]) & (g658) & (!g1310) & (g1311) & (!g1312) & (g1313)) + ((!sk[52]) & (g658) & (!g1310) & (g1311) & (g1312) & (!g1313)) + ((!sk[52]) & (g658) & (!g1310) & (g1311) & (g1312) & (g1313)) + ((!sk[52]) & (g658) & (g1310) & (!g1311) & (!g1312) & (!g1313)) + ((!sk[52]) & (g658) & (g1310) & (!g1311) & (!g1312) & (g1313)) + ((!sk[52]) & (g658) & (g1310) & (!g1311) & (g1312) & (!g1313)) + ((!sk[52]) & (g658) & (g1310) & (!g1311) & (g1312) & (g1313)) + ((!sk[52]) & (g658) & (g1310) & (g1311) & (!g1312) & (!g1313)) + ((!sk[52]) & (g658) & (g1310) & (g1311) & (!g1312) & (g1313)) + ((!sk[52]) & (g658) & (g1310) & (g1311) & (g1312) & (!g1313)) + ((!sk[52]) & (g658) & (g1310) & (g1311) & (g1312) & (g1313)) + ((sk[52]) & (!g658) & (!g1310) & (!g1311) & (!g1312) & (!g1313)));
	assign g1315 = (((!sk[53]) & (g173) & (!g546) & (!g907)) + ((!sk[53]) & (g173) & (!g546) & (g907)) + ((!sk[53]) & (g173) & (g546) & (!g907)) + ((!sk[53]) & (g173) & (g546) & (g907)) + ((sk[53]) & (!g173) & (!g546) & (!g907)));
	assign g1316 = (((!g550) & (!g630) & (sk[54]) & (g696)) + ((g550) & (!g630) & (!sk[54]) & (!g696)) + ((g550) & (!g630) & (!sk[54]) & (g696)) + ((g550) & (g630) & (!sk[54]) & (!g696)) + ((g550) & (g630) & (!sk[54]) & (g696)));
	assign g1317 = (((!g112) & (!g495) & (!g1153) & (!g1315) & (!sk[55]) & (g1316)) + ((!g112) & (!g495) & (!g1153) & (!g1315) & (sk[55]) & (!g1316)) + ((!g112) & (!g495) & (!g1153) & (!g1315) & (sk[55]) & (g1316)) + ((!g112) & (!g495) & (!g1153) & (g1315) & (!sk[55]) & (g1316)) + ((!g112) & (!g495) & (!g1153) & (g1315) & (sk[55]) & (!g1316)) + ((!g112) & (!g495) & (!g1153) & (g1315) & (sk[55]) & (g1316)) + ((!g112) & (!g495) & (g1153) & (!g1315) & (!sk[55]) & (g1316)) + ((!g112) & (!g495) & (g1153) & (g1315) & (!sk[55]) & (g1316)) + ((!g112) & (g495) & (!g1153) & (!g1315) & (!sk[55]) & (g1316)) + ((!g112) & (g495) & (!g1153) & (g1315) & (!sk[55]) & (g1316)) + ((!g112) & (g495) & (!g1153) & (g1315) & (sk[55]) & (!g1316)) + ((!g112) & (g495) & (!g1153) & (g1315) & (sk[55]) & (g1316)) + ((!g112) & (g495) & (g1153) & (!g1315) & (!sk[55]) & (g1316)) + ((!g112) & (g495) & (g1153) & (g1315) & (!sk[55]) & (g1316)) + ((g112) & (!g495) & (!g1153) & (!g1315) & (!sk[55]) & (!g1316)) + ((g112) & (!g495) & (!g1153) & (!g1315) & (!sk[55]) & (g1316)) + ((g112) & (!g495) & (!g1153) & (!g1315) & (sk[55]) & (g1316)) + ((g112) & (!g495) & (!g1153) & (g1315) & (!sk[55]) & (!g1316)) + ((g112) & (!g495) & (!g1153) & (g1315) & (!sk[55]) & (g1316)) + ((g112) & (!g495) & (!g1153) & (g1315) & (sk[55]) & (g1316)) + ((g112) & (!g495) & (g1153) & (!g1315) & (!sk[55]) & (!g1316)) + ((g112) & (!g495) & (g1153) & (!g1315) & (!sk[55]) & (g1316)) + ((g112) & (!g495) & (g1153) & (g1315) & (!sk[55]) & (!g1316)) + ((g112) & (!g495) & (g1153) & (g1315) & (!sk[55]) & (g1316)) + ((g112) & (g495) & (!g1153) & (!g1315) & (!sk[55]) & (!g1316)) + ((g112) & (g495) & (!g1153) & (!g1315) & (!sk[55]) & (g1316)) + ((g112) & (g495) & (!g1153) & (g1315) & (!sk[55]) & (!g1316)) + ((g112) & (g495) & (!g1153) & (g1315) & (!sk[55]) & (g1316)) + ((g112) & (g495) & (!g1153) & (g1315) & (sk[55]) & (g1316)) + ((g112) & (g495) & (g1153) & (!g1315) & (!sk[55]) & (!g1316)) + ((g112) & (g495) & (g1153) & (!g1315) & (!sk[55]) & (g1316)) + ((g112) & (g495) & (g1153) & (g1315) & (!sk[55]) & (!g1316)) + ((g112) & (g495) & (g1153) & (g1315) & (!sk[55]) & (g1316)));
	assign g1318 = (((!g1155) & (!g1305) & (g1307) & (g1309) & (g1314) & (g1317)));
	assign g1319 = (((g101) & (!g185) & (!g173) & (!g914) & (!g882) & (!g1170)) + ((g101) & (!g185) & (!g173) & (!g914) & (!g882) & (g1170)) + ((g101) & (!g185) & (!g173) & (!g914) & (g882) & (!g1170)) + ((g101) & (!g185) & (!g173) & (!g914) & (g882) & (g1170)) + ((g101) & (!g185) & (!g173) & (g914) & (!g882) & (!g1170)) + ((g101) & (!g185) & (!g173) & (g914) & (!g882) & (g1170)) + ((g101) & (!g185) & (!g173) & (g914) & (g882) & (!g1170)) + ((g101) & (!g185) & (!g173) & (g914) & (g882) & (g1170)) + ((g101) & (!g185) & (g173) & (!g914) & (!g882) & (!g1170)) + ((g101) & (!g185) & (g173) & (!g914) & (!g882) & (g1170)) + ((g101) & (!g185) & (g173) & (!g914) & (g882) & (!g1170)) + ((g101) & (!g185) & (g173) & (!g914) & (g882) & (g1170)) + ((g101) & (!g185) & (g173) & (g914) & (!g882) & (!g1170)) + ((g101) & (!g185) & (g173) & (g914) & (!g882) & (g1170)) + ((g101) & (!g185) & (g173) & (g914) & (g882) & (!g1170)) + ((g101) & (!g185) & (g173) & (g914) & (g882) & (g1170)) + ((g101) & (g185) & (!g173) & (!g914) & (!g882) & (!g1170)) + ((g101) & (g185) & (!g173) & (!g914) & (!g882) & (g1170)) + ((g101) & (g185) & (!g173) & (!g914) & (g882) & (!g1170)) + ((g101) & (g185) & (!g173) & (!g914) & (g882) & (g1170)) + ((g101) & (g185) & (!g173) & (g914) & (!g882) & (!g1170)) + ((g101) & (g185) & (!g173) & (g914) & (!g882) & (g1170)) + ((g101) & (g185) & (!g173) & (g914) & (g882) & (!g1170)) + ((g101) & (g185) & (g173) & (!g914) & (!g882) & (!g1170)) + ((g101) & (g185) & (g173) & (!g914) & (!g882) & (g1170)) + ((g101) & (g185) & (g173) & (!g914) & (g882) & (!g1170)) + ((g101) & (g185) & (g173) & (!g914) & (g882) & (g1170)) + ((g101) & (g185) & (g173) & (g914) & (!g882) & (!g1170)) + ((g101) & (g185) & (g173) & (g914) & (!g882) & (g1170)) + ((g101) & (g185) & (g173) & (g914) & (g882) & (!g1170)) + ((g101) & (g185) & (g173) & (g914) & (g882) & (g1170)));
	assign g1320 = (((!g99) & (!g173) & (!g103) & (sk[58]) & (!g929)) + ((!g99) & (!g173) & (g103) & (!sk[58]) & (g929)) + ((!g99) & (!g173) & (g103) & (sk[58]) & (!g929)) + ((!g99) & (g173) & (!g103) & (!sk[58]) & (!g929)) + ((!g99) & (g173) & (!g103) & (!sk[58]) & (g929)) + ((!g99) & (g173) & (!g103) & (sk[58]) & (!g929)) + ((!g99) & (g173) & (g103) & (!sk[58]) & (!g929)) + ((!g99) & (g173) & (g103) & (!sk[58]) & (g929)) + ((!g99) & (g173) & (g103) & (sk[58]) & (!g929)) + ((g99) & (!g173) & (g103) & (!sk[58]) & (!g929)) + ((g99) & (!g173) & (g103) & (!sk[58]) & (g929)) + ((g99) & (!g173) & (g103) & (sk[58]) & (!g929)) + ((g99) & (g173) & (!g103) & (!sk[58]) & (!g929)) + ((g99) & (g173) & (!g103) & (!sk[58]) & (g929)) + ((g99) & (g173) & (g103) & (!sk[58]) & (!g929)) + ((g99) & (g173) & (g103) & (!sk[58]) & (g929)));
	assign g1321 = (((!g570) & (!g1010) & (g1319) & (!sk[59]) & (g1320)) + ((!g570) & (g1010) & (!g1319) & (!sk[59]) & (!g1320)) + ((!g570) & (g1010) & (!g1319) & (!sk[59]) & (g1320)) + ((!g570) & (g1010) & (!g1319) & (sk[59]) & (g1320)) + ((!g570) & (g1010) & (g1319) & (!sk[59]) & (!g1320)) + ((!g570) & (g1010) & (g1319) & (!sk[59]) & (g1320)) + ((g570) & (!g1010) & (g1319) & (!sk[59]) & (!g1320)) + ((g570) & (!g1010) & (g1319) & (!sk[59]) & (g1320)) + ((g570) & (g1010) & (!g1319) & (!sk[59]) & (!g1320)) + ((g570) & (g1010) & (!g1319) & (!sk[59]) & (g1320)) + ((g570) & (g1010) & (g1319) & (!sk[59]) & (!g1320)) + ((g570) & (g1010) & (g1319) & (!sk[59]) & (g1320)));
	assign g1322 = (((!sk[60]) & (!g136) & (!g193) & (!g696) & (!g672) & (g702)) + ((!sk[60]) & (!g136) & (!g193) & (!g696) & (g672) & (g702)) + ((!sk[60]) & (!g136) & (!g193) & (g696) & (!g672) & (g702)) + ((!sk[60]) & (!g136) & (!g193) & (g696) & (g672) & (g702)) + ((!sk[60]) & (!g136) & (g193) & (!g696) & (!g672) & (g702)) + ((!sk[60]) & (!g136) & (g193) & (!g696) & (g672) & (g702)) + ((!sk[60]) & (!g136) & (g193) & (g696) & (!g672) & (g702)) + ((!sk[60]) & (!g136) & (g193) & (g696) & (g672) & (g702)) + ((!sk[60]) & (g136) & (!g193) & (!g696) & (!g672) & (!g702)) + ((!sk[60]) & (g136) & (!g193) & (!g696) & (!g672) & (g702)) + ((!sk[60]) & (g136) & (!g193) & (!g696) & (g672) & (!g702)) + ((!sk[60]) & (g136) & (!g193) & (!g696) & (g672) & (g702)) + ((!sk[60]) & (g136) & (!g193) & (g696) & (!g672) & (!g702)) + ((!sk[60]) & (g136) & (!g193) & (g696) & (!g672) & (g702)) + ((!sk[60]) & (g136) & (!g193) & (g696) & (g672) & (!g702)) + ((!sk[60]) & (g136) & (!g193) & (g696) & (g672) & (g702)) + ((!sk[60]) & (g136) & (g193) & (!g696) & (!g672) & (!g702)) + ((!sk[60]) & (g136) & (g193) & (!g696) & (!g672) & (g702)) + ((!sk[60]) & (g136) & (g193) & (!g696) & (g672) & (!g702)) + ((!sk[60]) & (g136) & (g193) & (!g696) & (g672) & (g702)) + ((!sk[60]) & (g136) & (g193) & (g696) & (!g672) & (!g702)) + ((!sk[60]) & (g136) & (g193) & (g696) & (!g672) & (g702)) + ((!sk[60]) & (g136) & (g193) & (g696) & (g672) & (!g702)) + ((!sk[60]) & (g136) & (g193) & (g696) & (g672) & (g702)) + ((sk[60]) & (g136) & (!g193) & (!g696) & (!g672) & (!g702)) + ((sk[60]) & (g136) & (!g193) & (!g696) & (!g672) & (g702)) + ((sk[60]) & (g136) & (!g193) & (!g696) & (g672) & (!g702)) + ((sk[60]) & (g136) & (!g193) & (!g696) & (g672) & (g702)) + ((sk[60]) & (g136) & (!g193) & (g696) & (!g672) & (g702)) + ((sk[60]) & (g136) & (!g193) & (g696) & (g672) & (!g702)) + ((sk[60]) & (g136) & (!g193) & (g696) & (g672) & (g702)) + ((sk[60]) & (g136) & (g193) & (!g696) & (!g672) & (!g702)) + ((sk[60]) & (g136) & (g193) & (!g696) & (!g672) & (g702)) + ((sk[60]) & (g136) & (g193) & (!g696) & (g672) & (!g702)) + ((sk[60]) & (g136) & (g193) & (!g696) & (g672) & (g702)) + ((sk[60]) & (g136) & (g193) & (g696) & (!g672) & (!g702)) + ((sk[60]) & (g136) & (g193) & (g696) & (!g672) & (g702)) + ((sk[60]) & (g136) & (g193) & (g696) & (g672) & (!g702)) + ((sk[60]) & (g136) & (g193) & (g696) & (g672) & (g702)));
	assign g1323 = (((!i_14_) & (!i_12_) & (!i_13_) & (!sk[61]) & (!g102) & (g115)) + ((!i_14_) & (!i_12_) & (!i_13_) & (!sk[61]) & (g102) & (g115)) + ((!i_14_) & (!i_12_) & (!i_13_) & (sk[61]) & (g102) & (!g115)) + ((!i_14_) & (!i_12_) & (!i_13_) & (sk[61]) & (g102) & (g115)) + ((!i_14_) & (!i_12_) & (i_13_) & (!sk[61]) & (!g102) & (g115)) + ((!i_14_) & (!i_12_) & (i_13_) & (!sk[61]) & (g102) & (g115)) + ((!i_14_) & (!i_12_) & (i_13_) & (sk[61]) & (!g102) & (g115)) + ((!i_14_) & (!i_12_) & (i_13_) & (sk[61]) & (g102) & (g115)) + ((!i_14_) & (i_12_) & (!i_13_) & (!sk[61]) & (!g102) & (g115)) + ((!i_14_) & (i_12_) & (!i_13_) & (!sk[61]) & (g102) & (g115)) + ((!i_14_) & (i_12_) & (!i_13_) & (sk[61]) & (!g102) & (g115)) + ((!i_14_) & (i_12_) & (!i_13_) & (sk[61]) & (g102) & (g115)) + ((!i_14_) & (i_12_) & (i_13_) & (!sk[61]) & (!g102) & (g115)) + ((!i_14_) & (i_12_) & (i_13_) & (!sk[61]) & (g102) & (g115)) + ((!i_14_) & (i_12_) & (i_13_) & (sk[61]) & (g102) & (g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (!sk[61]) & (!g102) & (!g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (!sk[61]) & (!g102) & (g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (!sk[61]) & (g102) & (!g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (!sk[61]) & (g102) & (g115)) + ((i_14_) & (!i_12_) & (!i_13_) & (sk[61]) & (g102) & (g115)) + ((i_14_) & (!i_12_) & (i_13_) & (!sk[61]) & (!g102) & (!g115)) + ((i_14_) & (!i_12_) & (i_13_) & (!sk[61]) & (!g102) & (g115)) + ((i_14_) & (!i_12_) & (i_13_) & (!sk[61]) & (g102) & (!g115)) + ((i_14_) & (!i_12_) & (i_13_) & (!sk[61]) & (g102) & (g115)) + ((i_14_) & (!i_12_) & (i_13_) & (sk[61]) & (!g102) & (g115)) + ((i_14_) & (!i_12_) & (i_13_) & (sk[61]) & (g102) & (g115)) + ((i_14_) & (i_12_) & (!i_13_) & (!sk[61]) & (!g102) & (!g115)) + ((i_14_) & (i_12_) & (!i_13_) & (!sk[61]) & (!g102) & (g115)) + ((i_14_) & (i_12_) & (!i_13_) & (!sk[61]) & (g102) & (!g115)) + ((i_14_) & (i_12_) & (!i_13_) & (!sk[61]) & (g102) & (g115)) + ((i_14_) & (i_12_) & (!i_13_) & (sk[61]) & (g102) & (g115)) + ((i_14_) & (i_12_) & (i_13_) & (!sk[61]) & (!g102) & (!g115)) + ((i_14_) & (i_12_) & (i_13_) & (!sk[61]) & (!g102) & (g115)) + ((i_14_) & (i_12_) & (i_13_) & (!sk[61]) & (g102) & (!g115)) + ((i_14_) & (i_12_) & (i_13_) & (!sk[61]) & (g102) & (g115)) + ((i_14_) & (i_12_) & (i_13_) & (sk[61]) & (g102) & (g115)));
	assign g1324 = (((!g134) & (!sk[62]) & (!g533) & (g779) & (g1323)) + ((!g134) & (!sk[62]) & (g533) & (!g779) & (!g1323)) + ((!g134) & (!sk[62]) & (g533) & (!g779) & (g1323)) + ((!g134) & (!sk[62]) & (g533) & (g779) & (!g1323)) + ((!g134) & (!sk[62]) & (g533) & (g779) & (g1323)) + ((!g134) & (sk[62]) & (!g533) & (!g779) & (!g1323)) + ((!g134) & (sk[62]) & (!g533) & (!g779) & (g1323)) + ((g134) & (!sk[62]) & (!g533) & (g779) & (!g1323)) + ((g134) & (!sk[62]) & (!g533) & (g779) & (g1323)) + ((g134) & (!sk[62]) & (g533) & (!g779) & (!g1323)) + ((g134) & (!sk[62]) & (g533) & (!g779) & (g1323)) + ((g134) & (!sk[62]) & (g533) & (g779) & (!g1323)) + ((g134) & (!sk[62]) & (g533) & (g779) & (g1323)) + ((g134) & (sk[62]) & (!g533) & (!g779) & (g1323)));
	assign g1325 = (((!g134) & (!sk[63]) & (!g136) & (g231) & (g232)) + ((!g134) & (!sk[63]) & (g136) & (!g231) & (!g232)) + ((!g134) & (!sk[63]) & (g136) & (!g231) & (g232)) + ((!g134) & (!sk[63]) & (g136) & (g231) & (!g232)) + ((!g134) & (!sk[63]) & (g136) & (g231) & (g232)) + ((!g134) & (sk[63]) & (g136) & (!g231) & (g232)) + ((!g134) & (sk[63]) & (g136) & (g231) & (g232)) + ((g134) & (!sk[63]) & (!g136) & (g231) & (!g232)) + ((g134) & (!sk[63]) & (!g136) & (g231) & (g232)) + ((g134) & (!sk[63]) & (g136) & (!g231) & (!g232)) + ((g134) & (!sk[63]) & (g136) & (!g231) & (g232)) + ((g134) & (!sk[63]) & (g136) & (g231) & (!g232)) + ((g134) & (!sk[63]) & (g136) & (g231) & (g232)) + ((g134) & (sk[63]) & (!g136) & (!g231) & (!g232)) + ((g134) & (sk[63]) & (!g136) & (!g231) & (g232)) + ((g134) & (sk[63]) & (g136) & (!g231) & (!g232)) + ((g134) & (sk[63]) & (g136) & (!g231) & (g232)) + ((g134) & (sk[63]) & (g136) & (g231) & (g232)));
	assign g1326 = (((!sk[64]) & (!i_8_) & (!g135) & (g907) & (g881)) + ((!sk[64]) & (!i_8_) & (g135) & (!g907) & (!g881)) + ((!sk[64]) & (!i_8_) & (g135) & (!g907) & (g881)) + ((!sk[64]) & (!i_8_) & (g135) & (g907) & (!g881)) + ((!sk[64]) & (!i_8_) & (g135) & (g907) & (g881)) + ((!sk[64]) & (i_8_) & (!g135) & (g907) & (!g881)) + ((!sk[64]) & (i_8_) & (!g135) & (g907) & (g881)) + ((!sk[64]) & (i_8_) & (g135) & (!g907) & (!g881)) + ((!sk[64]) & (i_8_) & (g135) & (!g907) & (g881)) + ((!sk[64]) & (i_8_) & (g135) & (g907) & (!g881)) + ((!sk[64]) & (i_8_) & (g135) & (g907) & (g881)) + ((sk[64]) & (i_8_) & (g135) & (!g907) & (g881)) + ((sk[64]) & (i_8_) & (g135) & (g907) & (!g881)) + ((sk[64]) & (i_8_) & (g135) & (g907) & (g881)));
	assign g1327 = (((!g134) & (!g220) & (!g103) & (!g105) & (!sk[65]) & (g837)) + ((!g134) & (!g220) & (!g103) & (g105) & (!sk[65]) & (g837)) + ((!g134) & (!g220) & (g103) & (!g105) & (!sk[65]) & (g837)) + ((!g134) & (!g220) & (g103) & (g105) & (!sk[65]) & (g837)) + ((!g134) & (g220) & (!g103) & (!g105) & (!sk[65]) & (g837)) + ((!g134) & (g220) & (!g103) & (g105) & (!sk[65]) & (g837)) + ((!g134) & (g220) & (g103) & (!g105) & (!sk[65]) & (g837)) + ((!g134) & (g220) & (g103) & (g105) & (!sk[65]) & (g837)) + ((g134) & (!g220) & (!g103) & (!g105) & (!sk[65]) & (!g837)) + ((g134) & (!g220) & (!g103) & (!g105) & (!sk[65]) & (g837)) + ((g134) & (!g220) & (!g103) & (!g105) & (sk[65]) & (!g837)) + ((g134) & (!g220) & (!g103) & (!g105) & (sk[65]) & (g837)) + ((g134) & (!g220) & (!g103) & (g105) & (!sk[65]) & (!g837)) + ((g134) & (!g220) & (!g103) & (g105) & (!sk[65]) & (g837)) + ((g134) & (!g220) & (!g103) & (g105) & (sk[65]) & (!g837)) + ((g134) & (!g220) & (!g103) & (g105) & (sk[65]) & (g837)) + ((g134) & (!g220) & (g103) & (!g105) & (!sk[65]) & (!g837)) + ((g134) & (!g220) & (g103) & (!g105) & (!sk[65]) & (g837)) + ((g134) & (!g220) & (g103) & (!g105) & (sk[65]) & (!g837)) + ((g134) & (!g220) & (g103) & (g105) & (!sk[65]) & (!g837)) + ((g134) & (!g220) & (g103) & (g105) & (!sk[65]) & (g837)) + ((g134) & (!g220) & (g103) & (g105) & (sk[65]) & (!g837)) + ((g134) & (!g220) & (g103) & (g105) & (sk[65]) & (g837)) + ((g134) & (g220) & (!g103) & (!g105) & (!sk[65]) & (!g837)) + ((g134) & (g220) & (!g103) & (!g105) & (!sk[65]) & (g837)) + ((g134) & (g220) & (!g103) & (!g105) & (sk[65]) & (!g837)) + ((g134) & (g220) & (!g103) & (!g105) & (sk[65]) & (g837)) + ((g134) & (g220) & (!g103) & (g105) & (!sk[65]) & (!g837)) + ((g134) & (g220) & (!g103) & (g105) & (!sk[65]) & (g837)) + ((g134) & (g220) & (!g103) & (g105) & (sk[65]) & (!g837)) + ((g134) & (g220) & (!g103) & (g105) & (sk[65]) & (g837)) + ((g134) & (g220) & (g103) & (!g105) & (!sk[65]) & (!g837)) + ((g134) & (g220) & (g103) & (!g105) & (!sk[65]) & (g837)) + ((g134) & (g220) & (g103) & (!g105) & (sk[65]) & (!g837)) + ((g134) & (g220) & (g103) & (!g105) & (sk[65]) & (g837)) + ((g134) & (g220) & (g103) & (g105) & (!sk[65]) & (!g837)) + ((g134) & (g220) & (g103) & (g105) & (!sk[65]) & (g837)) + ((g134) & (g220) & (g103) & (g105) & (sk[65]) & (!g837)) + ((g134) & (g220) & (g103) & (g105) & (sk[65]) & (g837)));
	assign g1328 = (((!g136) & (!g477) & (!g630) & (!g706) & (!g1326) & (!g1327)) + ((!g136) & (!g477) & (!g630) & (g706) & (!g1326) & (!g1327)) + ((!g136) & (!g477) & (g630) & (!g706) & (!g1326) & (!g1327)) + ((!g136) & (!g477) & (g630) & (g706) & (!g1326) & (!g1327)) + ((!g136) & (g477) & (!g630) & (!g706) & (!g1326) & (!g1327)) + ((!g136) & (g477) & (!g630) & (g706) & (!g1326) & (!g1327)) + ((!g136) & (g477) & (g630) & (!g706) & (!g1326) & (!g1327)) + ((!g136) & (g477) & (g630) & (g706) & (!g1326) & (!g1327)) + ((g136) & (g477) & (!g630) & (!g706) & (!g1326) & (!g1327)));
	assign g1329 = (((!g1152) & (!g1181) & (!g1322) & (g1324) & (!g1325) & (g1328)));
	assign g1330 = (((!g145) & (!sk[68]) & (!g269) & (!g1082) & (!g1191) & (g1589)) + ((!g145) & (!sk[68]) & (!g269) & (!g1082) & (g1191) & (g1589)) + ((!g145) & (!sk[68]) & (!g269) & (g1082) & (!g1191) & (g1589)) + ((!g145) & (!sk[68]) & (!g269) & (g1082) & (g1191) & (g1589)) + ((!g145) & (!sk[68]) & (g269) & (!g1082) & (!g1191) & (g1589)) + ((!g145) & (!sk[68]) & (g269) & (!g1082) & (g1191) & (g1589)) + ((!g145) & (!sk[68]) & (g269) & (g1082) & (!g1191) & (g1589)) + ((!g145) & (!sk[68]) & (g269) & (g1082) & (g1191) & (g1589)) + ((!g145) & (sk[68]) & (!g269) & (!g1082) & (!g1191) & (g1589)) + ((!g145) & (sk[68]) & (!g269) & (g1082) & (!g1191) & (g1589)) + ((!g145) & (sk[68]) & (g269) & (!g1082) & (!g1191) & (g1589)) + ((!g145) & (sk[68]) & (g269) & (g1082) & (!g1191) & (g1589)) + ((g145) & (!sk[68]) & (!g269) & (!g1082) & (!g1191) & (!g1589)) + ((g145) & (!sk[68]) & (!g269) & (!g1082) & (!g1191) & (g1589)) + ((g145) & (!sk[68]) & (!g269) & (!g1082) & (g1191) & (!g1589)) + ((g145) & (!sk[68]) & (!g269) & (!g1082) & (g1191) & (g1589)) + ((g145) & (!sk[68]) & (!g269) & (g1082) & (!g1191) & (!g1589)) + ((g145) & (!sk[68]) & (!g269) & (g1082) & (!g1191) & (g1589)) + ((g145) & (!sk[68]) & (!g269) & (g1082) & (g1191) & (!g1589)) + ((g145) & (!sk[68]) & (!g269) & (g1082) & (g1191) & (g1589)) + ((g145) & (!sk[68]) & (g269) & (!g1082) & (!g1191) & (!g1589)) + ((g145) & (!sk[68]) & (g269) & (!g1082) & (!g1191) & (g1589)) + ((g145) & (!sk[68]) & (g269) & (!g1082) & (g1191) & (!g1589)) + ((g145) & (!sk[68]) & (g269) & (!g1082) & (g1191) & (g1589)) + ((g145) & (!sk[68]) & (g269) & (g1082) & (!g1191) & (!g1589)) + ((g145) & (!sk[68]) & (g269) & (g1082) & (!g1191) & (g1589)) + ((g145) & (!sk[68]) & (g269) & (g1082) & (g1191) & (!g1589)) + ((g145) & (!sk[68]) & (g269) & (g1082) & (g1191) & (g1589)) + ((g145) & (sk[68]) & (!g269) & (!g1082) & (!g1191) & (g1589)));
	assign g1331 = (((!sk[69]) & (g89) & (!g1103)) + ((!sk[69]) & (g89) & (g1103)) + ((sk[69]) & (!g89) & (!g1103)));
	assign g1332 = (((!g323) & (!g195) & (!g105) & (!sk[70]) & (!g532) & (g921)) + ((!g323) & (!g195) & (!g105) & (!sk[70]) & (g532) & (g921)) + ((!g323) & (!g195) & (g105) & (!sk[70]) & (!g532) & (g921)) + ((!g323) & (!g195) & (g105) & (!sk[70]) & (g532) & (g921)) + ((!g323) & (g195) & (!g105) & (!sk[70]) & (!g532) & (g921)) + ((!g323) & (g195) & (!g105) & (!sk[70]) & (g532) & (g921)) + ((!g323) & (g195) & (g105) & (!sk[70]) & (!g532) & (g921)) + ((!g323) & (g195) & (g105) & (!sk[70]) & (g532) & (g921)) + ((g323) & (!g195) & (!g105) & (!sk[70]) & (!g532) & (!g921)) + ((g323) & (!g195) & (!g105) & (!sk[70]) & (!g532) & (g921)) + ((g323) & (!g195) & (!g105) & (!sk[70]) & (g532) & (!g921)) + ((g323) & (!g195) & (!g105) & (!sk[70]) & (g532) & (g921)) + ((g323) & (!g195) & (!g105) & (sk[70]) & (!g532) & (!g921)) + ((g323) & (!g195) & (!g105) & (sk[70]) & (g532) & (!g921)) + ((g323) & (!g195) & (!g105) & (sk[70]) & (g532) & (g921)) + ((g323) & (!g195) & (g105) & (!sk[70]) & (!g532) & (!g921)) + ((g323) & (!g195) & (g105) & (!sk[70]) & (!g532) & (g921)) + ((g323) & (!g195) & (g105) & (!sk[70]) & (g532) & (!g921)) + ((g323) & (!g195) & (g105) & (!sk[70]) & (g532) & (g921)) + ((g323) & (!g195) & (g105) & (sk[70]) & (!g532) & (!g921)) + ((g323) & (!g195) & (g105) & (sk[70]) & (!g532) & (g921)) + ((g323) & (!g195) & (g105) & (sk[70]) & (g532) & (!g921)) + ((g323) & (!g195) & (g105) & (sk[70]) & (g532) & (g921)) + ((g323) & (g195) & (!g105) & (!sk[70]) & (!g532) & (!g921)) + ((g323) & (g195) & (!g105) & (!sk[70]) & (!g532) & (g921)) + ((g323) & (g195) & (!g105) & (!sk[70]) & (g532) & (!g921)) + ((g323) & (g195) & (!g105) & (!sk[70]) & (g532) & (g921)) + ((g323) & (g195) & (!g105) & (sk[70]) & (!g532) & (!g921)) + ((g323) & (g195) & (!g105) & (sk[70]) & (!g532) & (g921)) + ((g323) & (g195) & (!g105) & (sk[70]) & (g532) & (!g921)) + ((g323) & (g195) & (!g105) & (sk[70]) & (g532) & (g921)) + ((g323) & (g195) & (g105) & (!sk[70]) & (!g532) & (!g921)) + ((g323) & (g195) & (g105) & (!sk[70]) & (!g532) & (g921)) + ((g323) & (g195) & (g105) & (!sk[70]) & (g532) & (!g921)) + ((g323) & (g195) & (g105) & (!sk[70]) & (g532) & (g921)) + ((g323) & (g195) & (g105) & (sk[70]) & (!g532) & (!g921)) + ((g323) & (g195) & (g105) & (sk[70]) & (!g532) & (g921)) + ((g323) & (g195) & (g105) & (sk[70]) & (g532) & (!g921)) + ((g323) & (g195) & (g105) & (sk[70]) & (g532) & (g921)));
	assign g1333 = (((!i_8_) & (!g88) & (g115) & (!sk[71]) & (g711)) + ((!i_8_) & (g88) & (!g115) & (!sk[71]) & (!g711)) + ((!i_8_) & (g88) & (!g115) & (!sk[71]) & (g711)) + ((!i_8_) & (g88) & (g115) & (!sk[71]) & (!g711)) + ((!i_8_) & (g88) & (g115) & (!sk[71]) & (g711)) + ((i_8_) & (!g88) & (g115) & (!sk[71]) & (!g711)) + ((i_8_) & (!g88) & (g115) & (!sk[71]) & (g711)) + ((i_8_) & (g88) & (!g115) & (!sk[71]) & (!g711)) + ((i_8_) & (g88) & (!g115) & (!sk[71]) & (g711)) + ((i_8_) & (g88) & (!g115) & (sk[71]) & (g711)) + ((i_8_) & (g88) & (g115) & (!sk[71]) & (!g711)) + ((i_8_) & (g88) & (g115) & (!sk[71]) & (g711)));
	assign g1334 = (((!sk[72]) & (!g118) & (!g232) & (g423) & (g630)) + ((!sk[72]) & (!g118) & (g232) & (!g423) & (!g630)) + ((!sk[72]) & (!g118) & (g232) & (!g423) & (g630)) + ((!sk[72]) & (!g118) & (g232) & (g423) & (!g630)) + ((!sk[72]) & (!g118) & (g232) & (g423) & (g630)) + ((!sk[72]) & (g118) & (!g232) & (g423) & (!g630)) + ((!sk[72]) & (g118) & (!g232) & (g423) & (g630)) + ((!sk[72]) & (g118) & (g232) & (!g423) & (!g630)) + ((!sk[72]) & (g118) & (g232) & (!g423) & (g630)) + ((!sk[72]) & (g118) & (g232) & (g423) & (!g630)) + ((!sk[72]) & (g118) & (g232) & (g423) & (g630)) + ((sk[72]) & (!g118) & (g232) & (g423) & (!g630)) + ((sk[72]) & (!g118) & (g232) & (g423) & (g630)) + ((sk[72]) & (g118) & (!g232) & (!g423) & (g630)) + ((sk[72]) & (g118) & (!g232) & (g423) & (g630)) + ((sk[72]) & (g118) & (g232) & (!g423) & (g630)) + ((sk[72]) & (g118) & (g232) & (g423) & (!g630)) + ((sk[72]) & (g118) & (g232) & (g423) & (g630)));
	assign g1335 = (((!g88) & (!sk[73]) & (!g103) & (g423) & (g1076)) + ((!g88) & (!sk[73]) & (g103) & (!g423) & (!g1076)) + ((!g88) & (!sk[73]) & (g103) & (!g423) & (g1076)) + ((!g88) & (!sk[73]) & (g103) & (g423) & (!g1076)) + ((!g88) & (!sk[73]) & (g103) & (g423) & (g1076)) + ((!g88) & (sk[73]) & (!g103) & (!g423) & (!g1076)) + ((!g88) & (sk[73]) & (!g103) & (!g423) & (g1076)) + ((!g88) & (sk[73]) & (g103) & (!g423) & (!g1076)) + ((!g88) & (sk[73]) & (g103) & (!g423) & (g1076)) + ((!g88) & (sk[73]) & (g103) & (g423) & (!g1076)) + ((g88) & (!sk[73]) & (!g103) & (g423) & (!g1076)) + ((g88) & (!sk[73]) & (!g103) & (g423) & (g1076)) + ((g88) & (!sk[73]) & (g103) & (!g423) & (!g1076)) + ((g88) & (!sk[73]) & (g103) & (!g423) & (g1076)) + ((g88) & (!sk[73]) & (g103) & (g423) & (!g1076)) + ((g88) & (!sk[73]) & (g103) & (g423) & (g1076)) + ((g88) & (sk[73]) & (!g103) & (!g423) & (!g1076)) + ((g88) & (sk[73]) & (g103) & (!g423) & (!g1076)) + ((g88) & (sk[73]) & (g103) & (g423) & (!g1076)));
	assign g1336 = (((!i_8_) & (!g88) & (!g264) & (!g103) & (g423) & (g675)) + ((!i_8_) & (!g88) & (!g264) & (g103) & (g423) & (g675)) + ((!i_8_) & (!g88) & (g264) & (!g103) & (g423) & (g675)) + ((!i_8_) & (!g88) & (g264) & (g103) & (g423) & (g675)) + ((!i_8_) & (g88) & (!g264) & (!g103) & (g423) & (g675)) + ((!i_8_) & (g88) & (!g264) & (g103) & (g423) & (g675)) + ((!i_8_) & (g88) & (g264) & (!g103) & (g423) & (g675)) + ((!i_8_) & (g88) & (g264) & (g103) & (g423) & (g675)) + ((i_8_) & (!g88) & (!g264) & (!g103) & (g423) & (g675)) + ((i_8_) & (!g88) & (!g264) & (g103) & (g423) & (g675)) + ((i_8_) & (!g88) & (g264) & (!g103) & (g423) & (g675)) + ((i_8_) & (!g88) & (g264) & (g103) & (g423) & (g675)) + ((i_8_) & (g88) & (!g264) & (!g103) & (!g423) & (!g675)) + ((i_8_) & (g88) & (!g264) & (!g103) & (!g423) & (g675)) + ((i_8_) & (g88) & (!g264) & (!g103) & (g423) & (!g675)) + ((i_8_) & (g88) & (!g264) & (!g103) & (g423) & (g675)) + ((i_8_) & (g88) & (!g264) & (g103) & (!g423) & (g675)) + ((i_8_) & (g88) & (!g264) & (g103) & (g423) & (g675)) + ((i_8_) & (g88) & (g264) & (!g103) & (!g423) & (!g675)) + ((i_8_) & (g88) & (g264) & (!g103) & (!g423) & (g675)) + ((i_8_) & (g88) & (g264) & (!g103) & (g423) & (!g675)) + ((i_8_) & (g88) & (g264) & (!g103) & (g423) & (g675)) + ((i_8_) & (g88) & (g264) & (g103) & (!g423) & (!g675)) + ((i_8_) & (g88) & (g264) & (g103) & (!g423) & (g675)) + ((i_8_) & (g88) & (g264) & (g103) & (g423) & (!g675)) + ((i_8_) & (g88) & (g264) & (g103) & (g423) & (g675)));
	assign g1337 = (((!g323) & (!g837) & (!g1333) & (!g1334) & (g1335) & (!g1336)) + ((!g323) & (g837) & (!g1333) & (!g1334) & (g1335) & (!g1336)) + ((g323) & (g837) & (!g1333) & (!g1334) & (g1335) & (!g1336)));
	assign g1338 = (((!sk[76]) & (!i_8_) & (!g88) & (g423) & (g640)) + ((!sk[76]) & (!i_8_) & (g88) & (!g423) & (!g640)) + ((!sk[76]) & (!i_8_) & (g88) & (!g423) & (g640)) + ((!sk[76]) & (!i_8_) & (g88) & (g423) & (!g640)) + ((!sk[76]) & (!i_8_) & (g88) & (g423) & (g640)) + ((!sk[76]) & (i_8_) & (!g88) & (g423) & (!g640)) + ((!sk[76]) & (i_8_) & (!g88) & (g423) & (g640)) + ((!sk[76]) & (i_8_) & (g88) & (!g423) & (!g640)) + ((!sk[76]) & (i_8_) & (g88) & (!g423) & (g640)) + ((!sk[76]) & (i_8_) & (g88) & (g423) & (!g640)) + ((!sk[76]) & (i_8_) & (g88) & (g423) & (g640)) + ((sk[76]) & (!i_8_) & (!g88) & (g423) & (!g640)) + ((sk[76]) & (!i_8_) & (g88) & (g423) & (!g640)) + ((sk[76]) & (i_8_) & (!g88) & (g423) & (!g640)) + ((sk[76]) & (i_8_) & (g88) & (!g423) & (!g640)) + ((sk[76]) & (i_8_) & (g88) & (g423) & (!g640)));
	assign g1339 = (((!g145) & (!g187) & (!g534) & (!g702) & (!g881) & (!g1338)) + ((!g145) & (!g187) & (!g534) & (!g702) & (g881) & (!g1338)) + ((!g145) & (!g187) & (!g534) & (g702) & (!g881) & (!g1338)) + ((!g145) & (!g187) & (!g534) & (g702) & (g881) & (!g1338)) + ((!g145) & (!g187) & (g534) & (!g702) & (!g881) & (!g1338)) + ((!g145) & (!g187) & (g534) & (!g702) & (g881) & (!g1338)) + ((!g145) & (!g187) & (g534) & (g702) & (!g881) & (!g1338)) + ((!g145) & (!g187) & (g534) & (g702) & (g881) & (!g1338)) + ((!g145) & (g187) & (!g534) & (!g702) & (!g881) & (!g1338)) + ((!g145) & (g187) & (!g534) & (!g702) & (g881) & (!g1338)) + ((!g145) & (g187) & (!g534) & (g702) & (!g881) & (!g1338)) + ((!g145) & (g187) & (!g534) & (g702) & (g881) & (!g1338)) + ((!g145) & (g187) & (g534) & (!g702) & (!g881) & (!g1338)) + ((!g145) & (g187) & (g534) & (!g702) & (g881) & (!g1338)) + ((!g145) & (g187) & (g534) & (g702) & (!g881) & (!g1338)) + ((!g145) & (g187) & (g534) & (g702) & (g881) & (!g1338)) + ((g145) & (!g187) & (!g534) & (!g702) & (!g881) & (!g1338)));
	assign g1340 = (((g997) & (!g1331) & (g1616) & (!g1332) & (g1337) & (g1339)));
	assign g1341 = (((g1092) & (g1318) & (g1321) & (g1329) & (g1330) & (g1340)));
	assign g1342 = (((!sk[80]) & (!g44) & (!g43) & (g191) & (g530)) + ((!sk[80]) & (!g44) & (g43) & (!g191) & (!g530)) + ((!sk[80]) & (!g44) & (g43) & (!g191) & (g530)) + ((!sk[80]) & (!g44) & (g43) & (g191) & (!g530)) + ((!sk[80]) & (!g44) & (g43) & (g191) & (g530)) + ((!sk[80]) & (g44) & (!g43) & (g191) & (!g530)) + ((!sk[80]) & (g44) & (!g43) & (g191) & (g530)) + ((!sk[80]) & (g44) & (g43) & (!g191) & (!g530)) + ((!sk[80]) & (g44) & (g43) & (!g191) & (g530)) + ((!sk[80]) & (g44) & (g43) & (g191) & (!g530)) + ((!sk[80]) & (g44) & (g43) & (g191) & (g530)) + ((sk[80]) & (!g44) & (!g43) & (!g191) & (!g530)));
	assign g1343 = (((!i_8_) & (!sk[81]) & (!g108) & (!g142) & (!g117) & (g1342)) + ((!i_8_) & (!sk[81]) & (!g108) & (!g142) & (g117) & (g1342)) + ((!i_8_) & (!sk[81]) & (!g108) & (g142) & (!g117) & (g1342)) + ((!i_8_) & (!sk[81]) & (!g108) & (g142) & (g117) & (g1342)) + ((!i_8_) & (!sk[81]) & (g108) & (!g142) & (!g117) & (g1342)) + ((!i_8_) & (!sk[81]) & (g108) & (!g142) & (g117) & (g1342)) + ((!i_8_) & (!sk[81]) & (g108) & (g142) & (!g117) & (g1342)) + ((!i_8_) & (!sk[81]) & (g108) & (g142) & (g117) & (g1342)) + ((!i_8_) & (sk[81]) & (g108) & (!g142) & (!g117) & (!g1342)) + ((!i_8_) & (sk[81]) & (g108) & (!g142) & (g117) & (!g1342)) + ((!i_8_) & (sk[81]) & (g108) & (!g142) & (g117) & (g1342)) + ((!i_8_) & (sk[81]) & (g108) & (g142) & (!g117) & (!g1342)) + ((!i_8_) & (sk[81]) & (g108) & (g142) & (!g117) & (g1342)) + ((!i_8_) & (sk[81]) & (g108) & (g142) & (g117) & (!g1342)) + ((!i_8_) & (sk[81]) & (g108) & (g142) & (g117) & (g1342)) + ((i_8_) & (!sk[81]) & (!g108) & (!g142) & (!g117) & (!g1342)) + ((i_8_) & (!sk[81]) & (!g108) & (!g142) & (!g117) & (g1342)) + ((i_8_) & (!sk[81]) & (!g108) & (!g142) & (g117) & (!g1342)) + ((i_8_) & (!sk[81]) & (!g108) & (!g142) & (g117) & (g1342)) + ((i_8_) & (!sk[81]) & (!g108) & (g142) & (!g117) & (!g1342)) + ((i_8_) & (!sk[81]) & (!g108) & (g142) & (!g117) & (g1342)) + ((i_8_) & (!sk[81]) & (!g108) & (g142) & (g117) & (!g1342)) + ((i_8_) & (!sk[81]) & (!g108) & (g142) & (g117) & (g1342)) + ((i_8_) & (!sk[81]) & (g108) & (!g142) & (!g117) & (!g1342)) + ((i_8_) & (!sk[81]) & (g108) & (!g142) & (!g117) & (g1342)) + ((i_8_) & (!sk[81]) & (g108) & (!g142) & (g117) & (!g1342)) + ((i_8_) & (!sk[81]) & (g108) & (!g142) & (g117) & (g1342)) + ((i_8_) & (!sk[81]) & (g108) & (g142) & (!g117) & (!g1342)) + ((i_8_) & (!sk[81]) & (g108) & (g142) & (!g117) & (g1342)) + ((i_8_) & (!sk[81]) & (g108) & (g142) & (g117) & (!g1342)) + ((i_8_) & (!sk[81]) & (g108) & (g142) & (g117) & (g1342)) + ((i_8_) & (sk[81]) & (g108) & (!g142) & (g117) & (!g1342)) + ((i_8_) & (sk[81]) & (g108) & (!g142) & (g117) & (g1342)) + ((i_8_) & (sk[81]) & (g108) & (g142) & (!g117) & (!g1342)) + ((i_8_) & (sk[81]) & (g108) & (g142) & (!g117) & (g1342)) + ((i_8_) & (sk[81]) & (g108) & (g142) & (g117) & (!g1342)) + ((i_8_) & (sk[81]) & (g108) & (g142) & (g117) & (g1342)));
	assign g1344 = (((!i_8_) & (!g19) & (g108) & (!sk[82]) & (g462)) + ((!i_8_) & (g19) & (!g108) & (!sk[82]) & (!g462)) + ((!i_8_) & (g19) & (!g108) & (!sk[82]) & (g462)) + ((!i_8_) & (g19) & (g108) & (!sk[82]) & (!g462)) + ((!i_8_) & (g19) & (g108) & (!sk[82]) & (g462)) + ((!i_8_) & (g19) & (g108) & (sk[82]) & (!g462)) + ((!i_8_) & (g19) & (g108) & (sk[82]) & (g462)) + ((i_8_) & (!g19) & (g108) & (!sk[82]) & (!g462)) + ((i_8_) & (!g19) & (g108) & (!sk[82]) & (g462)) + ((i_8_) & (!g19) & (g108) & (sk[82]) & (!g462)) + ((i_8_) & (g19) & (!g108) & (!sk[82]) & (!g462)) + ((i_8_) & (g19) & (!g108) & (!sk[82]) & (g462)) + ((i_8_) & (g19) & (g108) & (!sk[82]) & (!g462)) + ((i_8_) & (g19) & (g108) & (!sk[82]) & (g462)) + ((i_8_) & (g19) & (g108) & (sk[82]) & (!g462)));
	assign g1345 = (((!i_14_) & (!i_12_) & (!i_13_) & (i_8_) & (!g15) & (g108)) + ((!i_14_) & (i_12_) & (!i_13_) & (!i_8_) & (!g15) & (g108)) + ((!i_14_) & (i_12_) & (!i_13_) & (i_8_) & (!g15) & (g108)) + ((!i_14_) & (i_12_) & (i_13_) & (!i_8_) & (!g15) & (g108)) + ((!i_14_) & (i_12_) & (i_13_) & (i_8_) & (!g15) & (g108)) + ((i_14_) & (!i_12_) & (!i_13_) & (!i_8_) & (!g15) & (g108)) + ((i_14_) & (!i_12_) & (!i_13_) & (i_8_) & (!g15) & (g108)));
	assign g1346 = (((!g109) & (!g201) & (!g172) & (!g339) & (!g1344) & (!g1345)) + ((!g109) & (!g201) & (!g172) & (g339) & (!g1344) & (!g1345)) + ((!g109) & (!g201) & (g172) & (!g339) & (!g1344) & (!g1345)) + ((!g109) & (!g201) & (g172) & (g339) & (!g1344) & (!g1345)) + ((!g109) & (g201) & (!g172) & (!g339) & (!g1344) & (!g1345)) + ((!g109) & (g201) & (!g172) & (g339) & (!g1344) & (!g1345)) + ((!g109) & (g201) & (g172) & (!g339) & (!g1344) & (!g1345)) + ((!g109) & (g201) & (g172) & (g339) & (!g1344) & (!g1345)) + ((g109) & (g201) & (!g172) & (!g339) & (!g1344) & (!g1345)));
	assign g1347 = (((!g145) & (!g497) & (!g668) & (!g1122) & (!g1343) & (g1346)) + ((!g145) & (!g497) & (!g668) & (g1122) & (!g1343) & (g1346)) + ((g145) & (!g497) & (!g668) & (g1122) & (!g1343) & (g1346)));
	assign g1348 = (((!g134) & (!sk[86]) & (!g136) & (g142) & (g465)) + ((!g134) & (!sk[86]) & (g136) & (!g142) & (!g465)) + ((!g134) & (!sk[86]) & (g136) & (!g142) & (g465)) + ((!g134) & (!sk[86]) & (g136) & (g142) & (!g465)) + ((!g134) & (!sk[86]) & (g136) & (g142) & (g465)) + ((!g134) & (sk[86]) & (g136) & (!g142) & (!g465)) + ((!g134) & (sk[86]) & (g136) & (g142) & (!g465)) + ((g134) & (!sk[86]) & (!g136) & (g142) & (!g465)) + ((g134) & (!sk[86]) & (!g136) & (g142) & (g465)) + ((g134) & (!sk[86]) & (g136) & (!g142) & (!g465)) + ((g134) & (!sk[86]) & (g136) & (!g142) & (g465)) + ((g134) & (!sk[86]) & (g136) & (g142) & (!g465)) + ((g134) & (!sk[86]) & (g136) & (g142) & (g465)) + ((g134) & (sk[86]) & (!g136) & (g142) & (!g465)) + ((g134) & (sk[86]) & (!g136) & (g142) & (g465)) + ((g134) & (sk[86]) & (g136) & (!g142) & (!g465)) + ((g134) & (sk[86]) & (g136) & (g142) & (!g465)) + ((g134) & (sk[86]) & (g136) & (g142) & (g465)));
	assign g1349 = (((!sk[87]) & (g134) & (!g222) & (!g530)) + ((!sk[87]) & (g134) & (!g222) & (g530)) + ((!sk[87]) & (g134) & (g222) & (!g530)) + ((!sk[87]) & (g134) & (g222) & (g530)) + ((sk[87]) & (g134) & (!g222) & (g530)) + ((sk[87]) & (g134) & (g222) & (!g530)) + ((sk[87]) & (g134) & (g222) & (g530)));
	assign g1350 = (((!g43) & (!g135) & (!sk[88]) & (!g781) & (!g1122) & (g1349)) + ((!g43) & (!g135) & (!sk[88]) & (!g781) & (g1122) & (g1349)) + ((!g43) & (!g135) & (!sk[88]) & (g781) & (!g1122) & (g1349)) + ((!g43) & (!g135) & (!sk[88]) & (g781) & (g1122) & (g1349)) + ((!g43) & (!g135) & (sk[88]) & (!g781) & (!g1122) & (!g1349)) + ((!g43) & (!g135) & (sk[88]) & (!g781) & (g1122) & (!g1349)) + ((!g43) & (g135) & (!sk[88]) & (!g781) & (!g1122) & (g1349)) + ((!g43) & (g135) & (!sk[88]) & (!g781) & (g1122) & (g1349)) + ((!g43) & (g135) & (!sk[88]) & (g781) & (!g1122) & (g1349)) + ((!g43) & (g135) & (!sk[88]) & (g781) & (g1122) & (g1349)) + ((!g43) & (g135) & (sk[88]) & (!g781) & (g1122) & (!g1349)) + ((g43) & (!g135) & (!sk[88]) & (!g781) & (!g1122) & (!g1349)) + ((g43) & (!g135) & (!sk[88]) & (!g781) & (!g1122) & (g1349)) + ((g43) & (!g135) & (!sk[88]) & (!g781) & (g1122) & (!g1349)) + ((g43) & (!g135) & (!sk[88]) & (!g781) & (g1122) & (g1349)) + ((g43) & (!g135) & (!sk[88]) & (g781) & (!g1122) & (!g1349)) + ((g43) & (!g135) & (!sk[88]) & (g781) & (!g1122) & (g1349)) + ((g43) & (!g135) & (!sk[88]) & (g781) & (g1122) & (!g1349)) + ((g43) & (!g135) & (!sk[88]) & (g781) & (g1122) & (g1349)) + ((g43) & (!g135) & (sk[88]) & (!g781) & (!g1122) & (!g1349)) + ((g43) & (!g135) & (sk[88]) & (!g781) & (g1122) & (!g1349)) + ((g43) & (g135) & (!sk[88]) & (!g781) & (!g1122) & (!g1349)) + ((g43) & (g135) & (!sk[88]) & (!g781) & (!g1122) & (g1349)) + ((g43) & (g135) & (!sk[88]) & (!g781) & (g1122) & (!g1349)) + ((g43) & (g135) & (!sk[88]) & (!g781) & (g1122) & (g1349)) + ((g43) & (g135) & (!sk[88]) & (g781) & (!g1122) & (!g1349)) + ((g43) & (g135) & (!sk[88]) & (g781) & (!g1122) & (g1349)) + ((g43) & (g135) & (!sk[88]) & (g781) & (g1122) & (!g1349)) + ((g43) & (g135) & (!sk[88]) & (g781) & (g1122) & (g1349)));
	assign g1351 = (((!g19) & (!sk[89]) & (!g16) & (!g136) & (!g222) & (g399)) + ((!g19) & (!sk[89]) & (!g16) & (!g136) & (g222) & (g399)) + ((!g19) & (!sk[89]) & (!g16) & (g136) & (!g222) & (g399)) + ((!g19) & (!sk[89]) & (!g16) & (g136) & (g222) & (g399)) + ((!g19) & (!sk[89]) & (g16) & (!g136) & (!g222) & (g399)) + ((!g19) & (!sk[89]) & (g16) & (!g136) & (g222) & (g399)) + ((!g19) & (!sk[89]) & (g16) & (g136) & (!g222) & (g399)) + ((!g19) & (!sk[89]) & (g16) & (g136) & (g222) & (g399)) + ((!g19) & (sk[89]) & (!g16) & (g136) & (!g222) & (!g399)) + ((!g19) & (sk[89]) & (!g16) & (g136) & (!g222) & (g399)) + ((!g19) & (sk[89]) & (!g16) & (g136) & (g222) & (!g399)) + ((!g19) & (sk[89]) & (!g16) & (g136) & (g222) & (g399)) + ((!g19) & (sk[89]) & (g16) & (g136) & (!g222) & (!g399)) + ((!g19) & (sk[89]) & (g16) & (g136) & (g222) & (!g399)) + ((!g19) & (sk[89]) & (g16) & (g136) & (g222) & (g399)) + ((g19) & (!sk[89]) & (!g16) & (!g136) & (!g222) & (!g399)) + ((g19) & (!sk[89]) & (!g16) & (!g136) & (!g222) & (g399)) + ((g19) & (!sk[89]) & (!g16) & (!g136) & (g222) & (!g399)) + ((g19) & (!sk[89]) & (!g16) & (!g136) & (g222) & (g399)) + ((g19) & (!sk[89]) & (!g16) & (g136) & (!g222) & (!g399)) + ((g19) & (!sk[89]) & (!g16) & (g136) & (!g222) & (g399)) + ((g19) & (!sk[89]) & (!g16) & (g136) & (g222) & (!g399)) + ((g19) & (!sk[89]) & (!g16) & (g136) & (g222) & (g399)) + ((g19) & (!sk[89]) & (g16) & (!g136) & (!g222) & (!g399)) + ((g19) & (!sk[89]) & (g16) & (!g136) & (!g222) & (g399)) + ((g19) & (!sk[89]) & (g16) & (!g136) & (g222) & (!g399)) + ((g19) & (!sk[89]) & (g16) & (!g136) & (g222) & (g399)) + ((g19) & (!sk[89]) & (g16) & (g136) & (!g222) & (!g399)) + ((g19) & (!sk[89]) & (g16) & (g136) & (!g222) & (g399)) + ((g19) & (!sk[89]) & (g16) & (g136) & (g222) & (!g399)) + ((g19) & (!sk[89]) & (g16) & (g136) & (g222) & (g399)) + ((g19) & (sk[89]) & (!g16) & (g136) & (!g222) & (!g399)) + ((g19) & (sk[89]) & (!g16) & (g136) & (!g222) & (g399)) + ((g19) & (sk[89]) & (!g16) & (g136) & (g222) & (!g399)) + ((g19) & (sk[89]) & (!g16) & (g136) & (g222) & (g399)) + ((g19) & (sk[89]) & (g16) & (g136) & (!g222) & (!g399)) + ((g19) & (sk[89]) & (g16) & (g136) & (!g222) & (g399)) + ((g19) & (sk[89]) & (g16) & (g136) & (g222) & (!g399)) + ((g19) & (sk[89]) & (g16) & (g136) & (g222) & (g399)));
	assign g1352 = (((!g136) & (!g339) & (!g1348) & (!sk[90]) & (!g1350) & (g1351)) + ((!g136) & (!g339) & (!g1348) & (!sk[90]) & (g1350) & (g1351)) + ((!g136) & (!g339) & (!g1348) & (sk[90]) & (g1350) & (!g1351)) + ((!g136) & (!g339) & (g1348) & (!sk[90]) & (!g1350) & (g1351)) + ((!g136) & (!g339) & (g1348) & (!sk[90]) & (g1350) & (g1351)) + ((!g136) & (g339) & (!g1348) & (!sk[90]) & (!g1350) & (g1351)) + ((!g136) & (g339) & (!g1348) & (!sk[90]) & (g1350) & (g1351)) + ((!g136) & (g339) & (!g1348) & (sk[90]) & (g1350) & (!g1351)) + ((!g136) & (g339) & (g1348) & (!sk[90]) & (!g1350) & (g1351)) + ((!g136) & (g339) & (g1348) & (!sk[90]) & (g1350) & (g1351)) + ((g136) & (!g339) & (!g1348) & (!sk[90]) & (!g1350) & (!g1351)) + ((g136) & (!g339) & (!g1348) & (!sk[90]) & (!g1350) & (g1351)) + ((g136) & (!g339) & (!g1348) & (!sk[90]) & (g1350) & (!g1351)) + ((g136) & (!g339) & (!g1348) & (!sk[90]) & (g1350) & (g1351)) + ((g136) & (!g339) & (!g1348) & (sk[90]) & (g1350) & (!g1351)) + ((g136) & (!g339) & (g1348) & (!sk[90]) & (!g1350) & (!g1351)) + ((g136) & (!g339) & (g1348) & (!sk[90]) & (!g1350) & (g1351)) + ((g136) & (!g339) & (g1348) & (!sk[90]) & (g1350) & (!g1351)) + ((g136) & (!g339) & (g1348) & (!sk[90]) & (g1350) & (g1351)) + ((g136) & (g339) & (!g1348) & (!sk[90]) & (!g1350) & (!g1351)) + ((g136) & (g339) & (!g1348) & (!sk[90]) & (!g1350) & (g1351)) + ((g136) & (g339) & (!g1348) & (!sk[90]) & (g1350) & (!g1351)) + ((g136) & (g339) & (!g1348) & (!sk[90]) & (g1350) & (g1351)) + ((g136) & (g339) & (g1348) & (!sk[90]) & (!g1350) & (!g1351)) + ((g136) & (g339) & (g1348) & (!sk[90]) & (!g1350) & (g1351)) + ((g136) & (g339) & (g1348) & (!sk[90]) & (g1350) & (!g1351)) + ((g136) & (g339) & (g1348) & (!sk[90]) & (g1350) & (g1351)));
	assign g1353 = (((!g149) & (!g191) & (!g338) & (!g340) & (g399) & (!g361)) + ((!g149) & (!g191) & (g338) & (!g340) & (!g399) & (!g361)) + ((!g149) & (!g191) & (g338) & (!g340) & (g399) & (!g361)) + ((!g149) & (g191) & (g338) & (!g340) & (!g399) & (!g361)) + ((!g149) & (g191) & (g338) & (!g340) & (g399) & (!g361)) + ((g149) & (!g191) & (!g338) & (!g340) & (g399) & (!g361)) + ((g149) & (!g191) & (g338) & (!g340) & (!g399) & (!g361)) + ((g149) & (!g191) & (g338) & (!g340) & (g399) & (!g361)));
	assign g1354 = (((!g804) & (!g805) & (g1673) & (g810) & (g1666) & (g1353)));
	assign g1355 = (((!g19) & (!g118) & (g117) & (!sk[93]) & (g462)) + ((!g19) & (g118) & (!g117) & (!sk[93]) & (!g462)) + ((!g19) & (g118) & (!g117) & (!sk[93]) & (g462)) + ((!g19) & (g118) & (!g117) & (sk[93]) & (!g462)) + ((!g19) & (g118) & (g117) & (!sk[93]) & (!g462)) + ((!g19) & (g118) & (g117) & (!sk[93]) & (g462)) + ((!g19) & (g118) & (g117) & (sk[93]) & (!g462)) + ((!g19) & (g118) & (g117) & (sk[93]) & (g462)) + ((g19) & (!g118) & (g117) & (!sk[93]) & (!g462)) + ((g19) & (!g118) & (g117) & (!sk[93]) & (g462)) + ((g19) & (g118) & (!g117) & (!sk[93]) & (!g462)) + ((g19) & (g118) & (!g117) & (!sk[93]) & (g462)) + ((g19) & (g118) & (!g117) & (sk[93]) & (!g462)) + ((g19) & (g118) & (!g117) & (sk[93]) & (g462)) + ((g19) & (g118) & (g117) & (!sk[93]) & (!g462)) + ((g19) & (g118) & (g117) & (!sk[93]) & (g462)) + ((g19) & (g118) & (g117) & (sk[93]) & (!g462)) + ((g19) & (g118) & (g117) & (sk[93]) & (g462)));
	assign g1356 = (((g112) & (!g222) & (!sk[94]) & (!g807)) + ((g112) & (!g222) & (!sk[94]) & (g807)) + ((g112) & (!g222) & (sk[94]) & (!g807)) + ((g112) & (g222) & (!sk[94]) & (!g807)) + ((g112) & (g222) & (!sk[94]) & (g807)) + ((g112) & (g222) & (sk[94]) & (!g807)) + ((g112) & (g222) & (sk[94]) & (g807)));
	assign g1357 = (((!g19) & (!g16) & (g112) & (!g142) & (!g339) & (!g465)) + ((!g19) & (!g16) & (g112) & (!g142) & (!g339) & (g465)) + ((!g19) & (!g16) & (g112) & (!g142) & (g339) & (!g465)) + ((!g19) & (!g16) & (g112) & (!g142) & (g339) & (g465)) + ((!g19) & (!g16) & (g112) & (g142) & (!g339) & (!g465)) + ((!g19) & (!g16) & (g112) & (g142) & (!g339) & (g465)) + ((!g19) & (!g16) & (g112) & (g142) & (g339) & (!g465)) + ((!g19) & (!g16) & (g112) & (g142) & (g339) & (g465)) + ((!g19) & (g16) & (g112) & (!g142) & (!g339) & (!g465)) + ((!g19) & (g16) & (g112) & (!g142) & (g339) & (!g465)) + ((!g19) & (g16) & (g112) & (!g142) & (g339) & (g465)) + ((!g19) & (g16) & (g112) & (g142) & (!g339) & (!g465)) + ((!g19) & (g16) & (g112) & (g142) & (!g339) & (g465)) + ((!g19) & (g16) & (g112) & (g142) & (g339) & (!g465)) + ((!g19) & (g16) & (g112) & (g142) & (g339) & (g465)) + ((g19) & (!g16) & (g112) & (!g142) & (!g339) & (!g465)) + ((g19) & (!g16) & (g112) & (!g142) & (!g339) & (g465)) + ((g19) & (!g16) & (g112) & (!g142) & (g339) & (!g465)) + ((g19) & (!g16) & (g112) & (!g142) & (g339) & (g465)) + ((g19) & (!g16) & (g112) & (g142) & (!g339) & (!g465)) + ((g19) & (!g16) & (g112) & (g142) & (!g339) & (g465)) + ((g19) & (!g16) & (g112) & (g142) & (g339) & (!g465)) + ((g19) & (!g16) & (g112) & (g142) & (g339) & (g465)) + ((g19) & (g16) & (g112) & (!g142) & (!g339) & (!g465)) + ((g19) & (g16) & (g112) & (!g142) & (!g339) & (g465)) + ((g19) & (g16) & (g112) & (!g142) & (g339) & (!g465)) + ((g19) & (g16) & (g112) & (!g142) & (g339) & (g465)) + ((g19) & (g16) & (g112) & (g142) & (!g339) & (!g465)) + ((g19) & (g16) & (g112) & (g142) & (!g339) & (g465)) + ((g19) & (g16) & (g112) & (g142) & (g339) & (!g465)) + ((g19) & (g16) & (g112) & (g142) & (g339) & (g465)));
	assign g1358 = (((!g16) & (!g118) & (!g378) & (!g1355) & (!g1356) & (!g1357)) + ((g16) & (!g118) & (!g378) & (!g1355) & (!g1356) & (!g1357)) + ((g16) & (g118) & (!g378) & (!g1355) & (!g1356) & (!g1357)));
	assign g1359 = (((!i_8_) & (g108) & (!g201) & (g641) & (!g703) & (!g908)) + ((!i_8_) & (g108) & (!g201) & (g641) & (!g703) & (g908)) + ((!i_8_) & (g108) & (!g201) & (g641) & (g703) & (!g908)) + ((!i_8_) & (g108) & (!g201) & (g641) & (g703) & (g908)) + ((!i_8_) & (g108) & (g201) & (g641) & (!g703) & (!g908)) + ((!i_8_) & (g108) & (g201) & (g641) & (!g703) & (g908)) + ((!i_8_) & (g108) & (g201) & (g641) & (g703) & (!g908)) + ((!i_8_) & (g108) & (g201) & (g641) & (g703) & (g908)) + ((i_8_) & (g108) & (!g201) & (!g641) & (!g703) & (!g908)) + ((i_8_) & (g108) & (!g201) & (!g641) & (!g703) & (g908)) + ((i_8_) & (g108) & (!g201) & (!g641) & (g703) & (!g908)) + ((i_8_) & (g108) & (!g201) & (!g641) & (g703) & (g908)) + ((i_8_) & (g108) & (!g201) & (g641) & (!g703) & (!g908)) + ((i_8_) & (g108) & (!g201) & (g641) & (!g703) & (g908)) + ((i_8_) & (g108) & (!g201) & (g641) & (g703) & (!g908)) + ((i_8_) & (g108) & (!g201) & (g641) & (g703) & (g908)) + ((i_8_) & (g108) & (g201) & (!g641) & (!g703) & (g908)) + ((i_8_) & (g108) & (g201) & (!g641) & (g703) & (!g908)) + ((i_8_) & (g108) & (g201) & (!g641) & (g703) & (g908)) + ((i_8_) & (g108) & (g201) & (g641) & (!g703) & (g908)) + ((i_8_) & (g108) & (g201) & (g641) & (g703) & (!g908)) + ((i_8_) & (g108) & (g201) & (g641) & (g703) & (g908)));
	assign g1360 = (((!sk[98]) & (g996) & (!g1359)) + ((!sk[98]) & (g996) & (g1359)) + ((sk[98]) & (g996) & (!g1359)));
	assign g1361 = (((!g43) & (sk[99]) & (!g641)) + ((g43) & (!sk[99]) & (!g641)) + ((g43) & (!sk[99]) & (g641)));
	assign g1362 = (((!g118) & (!g186) & (!sk[100]) & (g142) & (g898)) + ((!g118) & (!g186) & (sk[100]) & (!g142) & (!g898)) + ((!g118) & (!g186) & (sk[100]) & (!g142) & (g898)) + ((!g118) & (!g186) & (sk[100]) & (g142) & (!g898)) + ((!g118) & (!g186) & (sk[100]) & (g142) & (g898)) + ((!g118) & (g186) & (!sk[100]) & (!g142) & (!g898)) + ((!g118) & (g186) & (!sk[100]) & (!g142) & (g898)) + ((!g118) & (g186) & (!sk[100]) & (g142) & (!g898)) + ((!g118) & (g186) & (!sk[100]) & (g142) & (g898)) + ((!g118) & (g186) & (sk[100]) & (!g142) & (!g898)) + ((g118) & (!g186) & (!sk[100]) & (g142) & (!g898)) + ((g118) & (!g186) & (!sk[100]) & (g142) & (g898)) + ((g118) & (!g186) & (sk[100]) & (!g142) & (!g898)) + ((g118) & (g186) & (!sk[100]) & (!g142) & (!g898)) + ((g118) & (g186) & (!sk[100]) & (!g142) & (g898)) + ((g118) & (g186) & (!sk[100]) & (g142) & (!g898)) + ((g118) & (g186) & (!sk[100]) & (g142) & (g898)) + ((g118) & (g186) & (sk[100]) & (!g142) & (!g898)));
	assign g1363 = (((!g59) & (!g44) & (!sk[101]) & (g186) & (g495)) + ((!g59) & (g44) & (!sk[101]) & (!g186) & (!g495)) + ((!g59) & (g44) & (!sk[101]) & (!g186) & (g495)) + ((!g59) & (g44) & (!sk[101]) & (g186) & (!g495)) + ((!g59) & (g44) & (!sk[101]) & (g186) & (g495)) + ((!g59) & (g44) & (sk[101]) & (!g186) & (g495)) + ((!g59) & (g44) & (sk[101]) & (g186) & (!g495)) + ((!g59) & (g44) & (sk[101]) & (g186) & (g495)) + ((g59) & (!g44) & (!sk[101]) & (g186) & (!g495)) + ((g59) & (!g44) & (!sk[101]) & (g186) & (g495)) + ((g59) & (g44) & (!sk[101]) & (!g186) & (!g495)) + ((g59) & (g44) & (!sk[101]) & (!g186) & (g495)) + ((g59) & (g44) & (!sk[101]) & (g186) & (!g495)) + ((g59) & (g44) & (!sk[101]) & (g186) & (g495)) + ((g59) & (g44) & (sk[101]) & (!g186) & (!g495)) + ((g59) & (g44) & (sk[101]) & (!g186) & (g495)) + ((g59) & (g44) & (sk[101]) & (g186) & (!g495)) + ((g59) & (g44) & (sk[101]) & (g186) & (g495)));
	assign g1364 = (((!g59) & (!g146) & (!g251) & (g1361) & (g1362) & (!g1363)) + ((!g59) & (!g146) & (g251) & (g1361) & (g1362) & (!g1363)) + ((!g59) & (g146) & (!g251) & (!g1361) & (g1362) & (!g1363)) + ((!g59) & (g146) & (!g251) & (g1361) & (g1362) & (!g1363)) + ((!g59) & (g146) & (g251) & (g1361) & (g1362) & (!g1363)) + ((g59) & (!g146) & (!g251) & (g1361) & (g1362) & (!g1363)) + ((g59) & (!g146) & (g251) & (g1361) & (g1362) & (!g1363)) + ((g59) & (g146) & (!g251) & (g1361) & (g1362) & (!g1363)) + ((g59) & (g146) & (g251) & (g1361) & (g1362) & (!g1363)));
	assign g1365 = (((i_8_) & (!sk[103]) & (!g100) & (!g201)) + ((i_8_) & (!sk[103]) & (!g100) & (g201)) + ((i_8_) & (!sk[103]) & (g100) & (!g201)) + ((i_8_) & (!sk[103]) & (g100) & (g201)) + ((i_8_) & (sk[103]) & (g100) & (!g201)));
	assign g1366 = (((g134) & (!sk[104]) & (!g117)) + ((g134) & (!sk[104]) & (g117)) + ((g134) & (sk[104]) & (g117)));
	assign g1367 = (((!sk[105]) & (g20) & (!g88)) + ((!sk[105]) & (g20) & (g88)) + ((sk[105]) & (!g20) & (g88)));
	assign g1368 = (((g186) & (!sk[106]) & (!g908)) + ((g186) & (!sk[106]) & (g908)) + ((g186) & (sk[106]) & (g908)));
	assign g1369 = (((!sk[107]) & (g98) & (!g264) & (!g111)) + ((!sk[107]) & (g98) & (!g264) & (g111)) + ((!sk[107]) & (g98) & (g264) & (!g111)) + ((!sk[107]) & (g98) & (g264) & (g111)) + ((sk[107]) & (g98) & (g264) & (g111)));
	assign g1370 = (((!g1365) & (!g1366) & (!g1046) & (!g1367) & (!g1368) & (!g1369)));
	assign g1371 = (((!g15) & (!sk[109]) & (!g59) & (!g112) & (!g135) & (g461)) + ((!g15) & (!sk[109]) & (!g59) & (!g112) & (g135) & (g461)) + ((!g15) & (!sk[109]) & (!g59) & (g112) & (!g135) & (g461)) + ((!g15) & (!sk[109]) & (!g59) & (g112) & (g135) & (g461)) + ((!g15) & (!sk[109]) & (g59) & (!g112) & (!g135) & (g461)) + ((!g15) & (!sk[109]) & (g59) & (!g112) & (g135) & (g461)) + ((!g15) & (!sk[109]) & (g59) & (g112) & (!g135) & (g461)) + ((!g15) & (!sk[109]) & (g59) & (g112) & (g135) & (g461)) + ((!g15) & (sk[109]) & (!g59) & (!g112) & (g135) & (g461)) + ((!g15) & (sk[109]) & (!g59) & (g112) & (!g135) & (g461)) + ((!g15) & (sk[109]) & (!g59) & (g112) & (g135) & (g461)) + ((!g15) & (sk[109]) & (g59) & (!g112) & (!g135) & (g461)) + ((!g15) & (sk[109]) & (g59) & (!g112) & (g135) & (g461)) + ((!g15) & (sk[109]) & (g59) & (g112) & (!g135) & (g461)) + ((!g15) & (sk[109]) & (g59) & (g112) & (g135) & (g461)) + ((g15) & (!sk[109]) & (!g59) & (!g112) & (!g135) & (!g461)) + ((g15) & (!sk[109]) & (!g59) & (!g112) & (!g135) & (g461)) + ((g15) & (!sk[109]) & (!g59) & (!g112) & (g135) & (!g461)) + ((g15) & (!sk[109]) & (!g59) & (!g112) & (g135) & (g461)) + ((g15) & (!sk[109]) & (!g59) & (g112) & (!g135) & (!g461)) + ((g15) & (!sk[109]) & (!g59) & (g112) & (!g135) & (g461)) + ((g15) & (!sk[109]) & (!g59) & (g112) & (g135) & (!g461)) + ((g15) & (!sk[109]) & (!g59) & (g112) & (g135) & (g461)) + ((g15) & (!sk[109]) & (g59) & (!g112) & (!g135) & (!g461)) + ((g15) & (!sk[109]) & (g59) & (!g112) & (!g135) & (g461)) + ((g15) & (!sk[109]) & (g59) & (!g112) & (g135) & (!g461)) + ((g15) & (!sk[109]) & (g59) & (!g112) & (g135) & (g461)) + ((g15) & (!sk[109]) & (g59) & (g112) & (!g135) & (!g461)) + ((g15) & (!sk[109]) & (g59) & (g112) & (!g135) & (g461)) + ((g15) & (!sk[109]) & (g59) & (g112) & (g135) & (!g461)) + ((g15) & (!sk[109]) & (g59) & (g112) & (g135) & (g461)));
	assign g1372 = (((!g375) & (!g164) & (!g1371) & (!sk[110]) & (!g1034) & (g1035)) + ((!g375) & (!g164) & (!g1371) & (!sk[110]) & (g1034) & (g1035)) + ((!g375) & (!g164) & (!g1371) & (sk[110]) & (!g1034) & (!g1035)) + ((!g375) & (!g164) & (g1371) & (!sk[110]) & (!g1034) & (g1035)) + ((!g375) & (!g164) & (g1371) & (!sk[110]) & (g1034) & (g1035)) + ((!g375) & (g164) & (!g1371) & (!sk[110]) & (!g1034) & (g1035)) + ((!g375) & (g164) & (!g1371) & (!sk[110]) & (g1034) & (g1035)) + ((!g375) & (g164) & (!g1371) & (sk[110]) & (!g1034) & (!g1035)) + ((!g375) & (g164) & (g1371) & (!sk[110]) & (!g1034) & (g1035)) + ((!g375) & (g164) & (g1371) & (!sk[110]) & (g1034) & (g1035)) + ((g375) & (!g164) & (!g1371) & (!sk[110]) & (!g1034) & (!g1035)) + ((g375) & (!g164) & (!g1371) & (!sk[110]) & (!g1034) & (g1035)) + ((g375) & (!g164) & (!g1371) & (!sk[110]) & (g1034) & (!g1035)) + ((g375) & (!g164) & (!g1371) & (!sk[110]) & (g1034) & (g1035)) + ((g375) & (!g164) & (!g1371) & (sk[110]) & (!g1034) & (!g1035)) + ((g375) & (!g164) & (g1371) & (!sk[110]) & (!g1034) & (!g1035)) + ((g375) & (!g164) & (g1371) & (!sk[110]) & (!g1034) & (g1035)) + ((g375) & (!g164) & (g1371) & (!sk[110]) & (g1034) & (!g1035)) + ((g375) & (!g164) & (g1371) & (!sk[110]) & (g1034) & (g1035)) + ((g375) & (g164) & (!g1371) & (!sk[110]) & (!g1034) & (!g1035)) + ((g375) & (g164) & (!g1371) & (!sk[110]) & (!g1034) & (g1035)) + ((g375) & (g164) & (!g1371) & (!sk[110]) & (g1034) & (!g1035)) + ((g375) & (g164) & (!g1371) & (!sk[110]) & (g1034) & (g1035)) + ((g375) & (g164) & (g1371) & (!sk[110]) & (!g1034) & (!g1035)) + ((g375) & (g164) & (g1371) & (!sk[110]) & (!g1034) & (g1035)) + ((g375) & (g164) & (g1371) & (!sk[110]) & (g1034) & (!g1035)) + ((g375) & (g164) & (g1371) & (!sk[110]) & (g1034) & (g1035)));
	assign g1373 = (((g1358) & (g1360) & (g1580) & (g1364) & (g1370) & (g1372)));
	assign g1374 = (((!g23) & (!g12) & (!g109) & (sk[112]) & (!g1233)) + ((!g23) & (!g12) & (g109) & (!sk[112]) & (g1233)) + ((!g23) & (!g12) & (g109) & (sk[112]) & (!g1233)) + ((!g23) & (g12) & (!g109) & (!sk[112]) & (!g1233)) + ((!g23) & (g12) & (!g109) & (!sk[112]) & (g1233)) + ((!g23) & (g12) & (!g109) & (sk[112]) & (!g1233)) + ((!g23) & (g12) & (g109) & (!sk[112]) & (!g1233)) + ((!g23) & (g12) & (g109) & (!sk[112]) & (g1233)) + ((g23) & (!g12) & (!g109) & (sk[112]) & (!g1233)) + ((g23) & (!g12) & (g109) & (!sk[112]) & (!g1233)) + ((g23) & (!g12) & (g109) & (!sk[112]) & (g1233)) + ((g23) & (g12) & (!g109) & (!sk[112]) & (!g1233)) + ((g23) & (g12) & (!g109) & (!sk[112]) & (g1233)) + ((g23) & (g12) & (!g109) & (sk[112]) & (!g1233)) + ((g23) & (g12) & (g109) & (!sk[112]) & (!g1233)) + ((g23) & (g12) & (g109) & (!sk[112]) & (g1233)));
	assign g1375 = (((!g31) & (!sk[113]) & (!g19) & (!g87) & (!g339) & (g465)) + ((!g31) & (!sk[113]) & (!g19) & (!g87) & (g339) & (g465)) + ((!g31) & (!sk[113]) & (!g19) & (g87) & (!g339) & (g465)) + ((!g31) & (!sk[113]) & (!g19) & (g87) & (g339) & (g465)) + ((!g31) & (!sk[113]) & (g19) & (!g87) & (!g339) & (g465)) + ((!g31) & (!sk[113]) & (g19) & (!g87) & (g339) & (g465)) + ((!g31) & (!sk[113]) & (g19) & (g87) & (!g339) & (g465)) + ((!g31) & (!sk[113]) & (g19) & (g87) & (g339) & (g465)) + ((g31) & (!sk[113]) & (!g19) & (!g87) & (!g339) & (!g465)) + ((g31) & (!sk[113]) & (!g19) & (!g87) & (!g339) & (g465)) + ((g31) & (!sk[113]) & (!g19) & (!g87) & (g339) & (!g465)) + ((g31) & (!sk[113]) & (!g19) & (!g87) & (g339) & (g465)) + ((g31) & (!sk[113]) & (!g19) & (g87) & (!g339) & (!g465)) + ((g31) & (!sk[113]) & (!g19) & (g87) & (!g339) & (g465)) + ((g31) & (!sk[113]) & (!g19) & (g87) & (g339) & (!g465)) + ((g31) & (!sk[113]) & (!g19) & (g87) & (g339) & (g465)) + ((g31) & (!sk[113]) & (g19) & (!g87) & (!g339) & (!g465)) + ((g31) & (!sk[113]) & (g19) & (!g87) & (!g339) & (g465)) + ((g31) & (!sk[113]) & (g19) & (!g87) & (g339) & (!g465)) + ((g31) & (!sk[113]) & (g19) & (!g87) & (g339) & (g465)) + ((g31) & (!sk[113]) & (g19) & (g87) & (!g339) & (!g465)) + ((g31) & (!sk[113]) & (g19) & (g87) & (!g339) & (g465)) + ((g31) & (!sk[113]) & (g19) & (g87) & (g339) & (!g465)) + ((g31) & (!sk[113]) & (g19) & (g87) & (g339) & (g465)) + ((g31) & (sk[113]) & (!g19) & (g87) & (!g339) & (!g465)) + ((g31) & (sk[113]) & (!g19) & (g87) & (g339) & (!g465)) + ((g31) & (sk[113]) & (!g19) & (g87) & (g339) & (g465)) + ((g31) & (sk[113]) & (g19) & (g87) & (!g339) & (!g465)) + ((g31) & (sk[113]) & (g19) & (g87) & (!g339) & (g465)) + ((g31) & (sk[113]) & (g19) & (g87) & (g339) & (!g465)) + ((g31) & (sk[113]) & (g19) & (g87) & (g339) & (g465)));
	assign g1376 = (((!g172) & (!sk[114]) & (!g214) & (g495) & (g1375)) + ((!g172) & (!sk[114]) & (g214) & (!g495) & (!g1375)) + ((!g172) & (!sk[114]) & (g214) & (!g495) & (g1375)) + ((!g172) & (!sk[114]) & (g214) & (g495) & (!g1375)) + ((!g172) & (!sk[114]) & (g214) & (g495) & (g1375)) + ((!g172) & (sk[114]) & (!g214) & (!g495) & (!g1375)) + ((!g172) & (sk[114]) & (!g214) & (g495) & (!g1375)) + ((!g172) & (sk[114]) & (g214) & (!g495) & (!g1375)) + ((!g172) & (sk[114]) & (g214) & (g495) & (!g1375)) + ((g172) & (!sk[114]) & (!g214) & (g495) & (!g1375)) + ((g172) & (!sk[114]) & (!g214) & (g495) & (g1375)) + ((g172) & (!sk[114]) & (g214) & (!g495) & (!g1375)) + ((g172) & (!sk[114]) & (g214) & (!g495) & (g1375)) + ((g172) & (!sk[114]) & (g214) & (g495) & (!g1375)) + ((g172) & (!sk[114]) & (g214) & (g495) & (g1375)) + ((g172) & (sk[114]) & (!g214) & (!g495) & (!g1375)));
	assign g1377 = (((!g277) & (!g339) & (!sk[115]) & (g465) & (g1376)) + ((!g277) & (!g339) & (sk[115]) & (g465) & (g1376)) + ((!g277) & (g339) & (!sk[115]) & (!g465) & (!g1376)) + ((!g277) & (g339) & (!sk[115]) & (!g465) & (g1376)) + ((!g277) & (g339) & (!sk[115]) & (g465) & (!g1376)) + ((!g277) & (g339) & (!sk[115]) & (g465) & (g1376)) + ((g277) & (!g339) & (!sk[115]) & (g465) & (!g1376)) + ((g277) & (!g339) & (!sk[115]) & (g465) & (g1376)) + ((g277) & (!g339) & (sk[115]) & (!g465) & (g1376)) + ((g277) & (!g339) & (sk[115]) & (g465) & (g1376)) + ((g277) & (g339) & (!sk[115]) & (!g465) & (!g1376)) + ((g277) & (g339) & (!sk[115]) & (!g465) & (g1376)) + ((g277) & (g339) & (!sk[115]) & (g465) & (!g1376)) + ((g277) & (g339) & (!sk[115]) & (g465) & (g1376)) + ((g277) & (g339) & (sk[115]) & (!g465) & (g1376)) + ((g277) & (g339) & (sk[115]) & (g465) & (g1376)));
	assign g1378 = (((!i_8_) & (!g19) & (!g16) & (!g88) & (!g231) & (!g262)) + ((!i_8_) & (!g19) & (!g16) & (!g88) & (g231) & (!g262)) + ((!i_8_) & (!g19) & (!g16) & (g88) & (!g231) & (!g262)) + ((!i_8_) & (!g19) & (!g16) & (g88) & (g231) & (!g262)) + ((!i_8_) & (!g19) & (g16) & (!g88) & (!g231) & (!g262)) + ((!i_8_) & (!g19) & (g16) & (!g88) & (g231) & (!g262)) + ((!i_8_) & (!g19) & (g16) & (g88) & (!g231) & (!g262)) + ((!i_8_) & (!g19) & (g16) & (g88) & (g231) & (!g262)) + ((!i_8_) & (g19) & (!g16) & (!g88) & (!g231) & (!g262)) + ((!i_8_) & (g19) & (!g16) & (!g88) & (g231) & (!g262)) + ((!i_8_) & (g19) & (!g16) & (g88) & (!g231) & (!g262)) + ((!i_8_) & (g19) & (!g16) & (g88) & (g231) & (!g262)) + ((!i_8_) & (g19) & (g16) & (!g88) & (!g231) & (!g262)) + ((!i_8_) & (g19) & (g16) & (!g88) & (g231) & (!g262)) + ((!i_8_) & (g19) & (g16) & (g88) & (!g231) & (!g262)) + ((!i_8_) & (g19) & (g16) & (g88) & (g231) & (!g262)) + ((i_8_) & (!g19) & (!g16) & (!g88) & (!g231) & (!g262)) + ((i_8_) & (!g19) & (!g16) & (!g88) & (g231) & (!g262)) + ((i_8_) & (!g19) & (g16) & (!g88) & (!g231) & (!g262)) + ((i_8_) & (!g19) & (g16) & (!g88) & (g231) & (!g262)) + ((i_8_) & (!g19) & (g16) & (g88) & (g231) & (!g262)) + ((i_8_) & (g19) & (!g16) & (!g88) & (!g231) & (!g262)) + ((i_8_) & (g19) & (!g16) & (!g88) & (g231) & (!g262)) + ((i_8_) & (g19) & (g16) & (!g88) & (!g231) & (!g262)) + ((i_8_) & (g19) & (g16) & (!g88) & (g231) & (!g262)));
	assign g1379 = (((!sk[117]) & (!g101) & (!g151) & (!g530) & (!g636) & (g1378)) + ((!sk[117]) & (!g101) & (!g151) & (!g530) & (g636) & (g1378)) + ((!sk[117]) & (!g101) & (!g151) & (g530) & (!g636) & (g1378)) + ((!sk[117]) & (!g101) & (!g151) & (g530) & (g636) & (g1378)) + ((!sk[117]) & (!g101) & (g151) & (!g530) & (!g636) & (g1378)) + ((!sk[117]) & (!g101) & (g151) & (!g530) & (g636) & (g1378)) + ((!sk[117]) & (!g101) & (g151) & (g530) & (!g636) & (g1378)) + ((!sk[117]) & (!g101) & (g151) & (g530) & (g636) & (g1378)) + ((!sk[117]) & (g101) & (!g151) & (!g530) & (!g636) & (!g1378)) + ((!sk[117]) & (g101) & (!g151) & (!g530) & (!g636) & (g1378)) + ((!sk[117]) & (g101) & (!g151) & (!g530) & (g636) & (!g1378)) + ((!sk[117]) & (g101) & (!g151) & (!g530) & (g636) & (g1378)) + ((!sk[117]) & (g101) & (!g151) & (g530) & (!g636) & (!g1378)) + ((!sk[117]) & (g101) & (!g151) & (g530) & (!g636) & (g1378)) + ((!sk[117]) & (g101) & (!g151) & (g530) & (g636) & (!g1378)) + ((!sk[117]) & (g101) & (!g151) & (g530) & (g636) & (g1378)) + ((!sk[117]) & (g101) & (g151) & (!g530) & (!g636) & (!g1378)) + ((!sk[117]) & (g101) & (g151) & (!g530) & (!g636) & (g1378)) + ((!sk[117]) & (g101) & (g151) & (!g530) & (g636) & (!g1378)) + ((!sk[117]) & (g101) & (g151) & (!g530) & (g636) & (g1378)) + ((!sk[117]) & (g101) & (g151) & (g530) & (!g636) & (!g1378)) + ((!sk[117]) & (g101) & (g151) & (g530) & (!g636) & (g1378)) + ((!sk[117]) & (g101) & (g151) & (g530) & (g636) & (!g1378)) + ((!sk[117]) & (g101) & (g151) & (g530) & (g636) & (g1378)) + ((sk[117]) & (!g101) & (!g151) & (!g530) & (!g636) & (g1378)) + ((sk[117]) & (!g101) & (!g151) & (!g530) & (g636) & (g1378)) + ((sk[117]) & (!g101) & (!g151) & (g530) & (!g636) & (g1378)) + ((sk[117]) & (!g101) & (!g151) & (g530) & (g636) & (g1378)) + ((sk[117]) & (!g101) & (g151) & (!g530) & (g636) & (g1378)) + ((sk[117]) & (!g101) & (g151) & (g530) & (g636) & (g1378)) + ((sk[117]) & (g101) & (!g151) & (!g530) & (!g636) & (g1378)) + ((sk[117]) & (g101) & (!g151) & (!g530) & (g636) & (g1378)) + ((sk[117]) & (g101) & (g151) & (!g530) & (g636) & (g1378)));
	assign g1380 = (((!i_8_) & (!sk[118]) & (!g16) & (!g108) & (!g339) & (g636)) + ((!i_8_) & (!sk[118]) & (!g16) & (!g108) & (g339) & (g636)) + ((!i_8_) & (!sk[118]) & (!g16) & (g108) & (!g339) & (g636)) + ((!i_8_) & (!sk[118]) & (!g16) & (g108) & (g339) & (g636)) + ((!i_8_) & (!sk[118]) & (g16) & (!g108) & (!g339) & (g636)) + ((!i_8_) & (!sk[118]) & (g16) & (!g108) & (g339) & (g636)) + ((!i_8_) & (!sk[118]) & (g16) & (g108) & (!g339) & (g636)) + ((!i_8_) & (!sk[118]) & (g16) & (g108) & (g339) & (g636)) + ((!i_8_) & (sk[118]) & (!g16) & (g108) & (!g339) & (!g636)) + ((!i_8_) & (sk[118]) & (!g16) & (g108) & (!g339) & (g636)) + ((!i_8_) & (sk[118]) & (!g16) & (g108) & (g339) & (!g636)) + ((!i_8_) & (sk[118]) & (!g16) & (g108) & (g339) & (g636)) + ((i_8_) & (!sk[118]) & (!g16) & (!g108) & (!g339) & (!g636)) + ((i_8_) & (!sk[118]) & (!g16) & (!g108) & (!g339) & (g636)) + ((i_8_) & (!sk[118]) & (!g16) & (!g108) & (g339) & (!g636)) + ((i_8_) & (!sk[118]) & (!g16) & (!g108) & (g339) & (g636)) + ((i_8_) & (!sk[118]) & (!g16) & (g108) & (!g339) & (!g636)) + ((i_8_) & (!sk[118]) & (!g16) & (g108) & (!g339) & (g636)) + ((i_8_) & (!sk[118]) & (!g16) & (g108) & (g339) & (!g636)) + ((i_8_) & (!sk[118]) & (!g16) & (g108) & (g339) & (g636)) + ((i_8_) & (!sk[118]) & (g16) & (!g108) & (!g339) & (!g636)) + ((i_8_) & (!sk[118]) & (g16) & (!g108) & (!g339) & (g636)) + ((i_8_) & (!sk[118]) & (g16) & (!g108) & (g339) & (!g636)) + ((i_8_) & (!sk[118]) & (g16) & (!g108) & (g339) & (g636)) + ((i_8_) & (!sk[118]) & (g16) & (g108) & (!g339) & (!g636)) + ((i_8_) & (!sk[118]) & (g16) & (g108) & (!g339) & (g636)) + ((i_8_) & (!sk[118]) & (g16) & (g108) & (g339) & (!g636)) + ((i_8_) & (!sk[118]) & (g16) & (g108) & (g339) & (g636)) + ((i_8_) & (sk[118]) & (!g16) & (g108) & (!g339) & (!g636)) + ((i_8_) & (sk[118]) & (!g16) & (g108) & (g339) & (!g636)) + ((i_8_) & (sk[118]) & (!g16) & (g108) & (g339) & (g636)) + ((i_8_) & (sk[118]) & (g16) & (g108) & (!g339) & (!g636)) + ((i_8_) & (sk[118]) & (g16) & (g108) & (g339) & (!g636)) + ((i_8_) & (sk[118]) & (g16) & (g108) & (g339) & (g636)));
	assign g1381 = (((g1374) & (g1377) & (g1379) & (!g1380) & (g1068) & (g1131)));
	assign g1382 = (((g976) & (g1347) & (g1352) & (g1354) & (g1373) & (g1381)));
	assign o_18_ = (((g73) & (!g985) & (!g1221) & (!g1303) & (!g1341) & (!g1382)) + ((g73) & (!g985) & (!g1221) & (!g1303) & (!g1341) & (g1382)) + ((g73) & (!g985) & (!g1221) & (!g1303) & (g1341) & (!g1382)) + ((g73) & (!g985) & (!g1221) & (!g1303) & (g1341) & (g1382)) + ((g73) & (!g985) & (!g1221) & (g1303) & (!g1341) & (!g1382)) + ((g73) & (!g985) & (!g1221) & (g1303) & (!g1341) & (g1382)) + ((g73) & (!g985) & (!g1221) & (g1303) & (g1341) & (!g1382)) + ((g73) & (!g985) & (!g1221) & (g1303) & (g1341) & (g1382)) + ((g73) & (!g985) & (g1221) & (!g1303) & (!g1341) & (!g1382)) + ((g73) & (!g985) & (g1221) & (!g1303) & (!g1341) & (g1382)) + ((g73) & (!g985) & (g1221) & (!g1303) & (g1341) & (!g1382)) + ((g73) & (!g985) & (g1221) & (!g1303) & (g1341) & (g1382)) + ((g73) & (!g985) & (g1221) & (g1303) & (!g1341) & (!g1382)) + ((g73) & (!g985) & (g1221) & (g1303) & (!g1341) & (g1382)) + ((g73) & (!g985) & (g1221) & (g1303) & (g1341) & (!g1382)) + ((g73) & (!g985) & (g1221) & (g1303) & (g1341) & (g1382)) + ((g73) & (g985) & (!g1221) & (!g1303) & (!g1341) & (!g1382)) + ((g73) & (g985) & (!g1221) & (!g1303) & (!g1341) & (g1382)) + ((g73) & (g985) & (!g1221) & (!g1303) & (g1341) & (!g1382)) + ((g73) & (g985) & (!g1221) & (!g1303) & (g1341) & (g1382)) + ((g73) & (g985) & (!g1221) & (g1303) & (!g1341) & (!g1382)) + ((g73) & (g985) & (!g1221) & (g1303) & (!g1341) & (g1382)) + ((g73) & (g985) & (!g1221) & (g1303) & (g1341) & (!g1382)) + ((g73) & (g985) & (!g1221) & (g1303) & (g1341) & (g1382)) + ((g73) & (g985) & (g1221) & (!g1303) & (!g1341) & (!g1382)) + ((g73) & (g985) & (g1221) & (!g1303) & (!g1341) & (g1382)) + ((g73) & (g985) & (g1221) & (!g1303) & (g1341) & (!g1382)) + ((g73) & (g985) & (g1221) & (!g1303) & (g1341) & (g1382)) + ((g73) & (g985) & (g1221) & (g1303) & (!g1341) & (!g1382)) + ((g73) & (g985) & (g1221) & (g1303) & (!g1341) & (g1382)) + ((g73) & (g985) & (g1221) & (g1303) & (g1341) & (!g1382)));
	assign g1384 = (((!g203) & (!g678) & (!sk[122]) & (g669) & (g818)) + ((!g203) & (g678) & (!sk[122]) & (!g669) & (!g818)) + ((!g203) & (g678) & (!sk[122]) & (!g669) & (g818)) + ((!g203) & (g678) & (!sk[122]) & (g669) & (!g818)) + ((!g203) & (g678) & (!sk[122]) & (g669) & (g818)) + ((!g203) & (g678) & (sk[122]) & (g669) & (g818)) + ((g203) & (!g678) & (!sk[122]) & (g669) & (!g818)) + ((g203) & (!g678) & (!sk[122]) & (g669) & (g818)) + ((g203) & (g678) & (!sk[122]) & (!g669) & (!g818)) + ((g203) & (g678) & (!sk[122]) & (!g669) & (g818)) + ((g203) & (g678) & (!sk[122]) & (g669) & (!g818)) + ((g203) & (g678) & (!sk[122]) & (g669) & (g818)));
	assign g1385 = (((!sk[123]) & (!g134) & (!g304) & (g270) & (g136)) + ((!sk[123]) & (!g134) & (g304) & (!g270) & (!g136)) + ((!sk[123]) & (!g134) & (g304) & (!g270) & (g136)) + ((!sk[123]) & (!g134) & (g304) & (g270) & (!g136)) + ((!sk[123]) & (!g134) & (g304) & (g270) & (g136)) + ((!sk[123]) & (g134) & (!g304) & (g270) & (!g136)) + ((!sk[123]) & (g134) & (!g304) & (g270) & (g136)) + ((!sk[123]) & (g134) & (g304) & (!g270) & (!g136)) + ((!sk[123]) & (g134) & (g304) & (!g270) & (g136)) + ((!sk[123]) & (g134) & (g304) & (g270) & (!g136)) + ((!sk[123]) & (g134) & (g304) & (g270) & (g136)) + ((sk[123]) & (!g134) & (!g304) & (!g270) & (g136)) + ((sk[123]) & (!g134) & (g304) & (!g270) & (g136)) + ((sk[123]) & (g134) & (!g304) & (!g270) & (g136)) + ((sk[123]) & (g134) & (g304) & (!g270) & (!g136)) + ((sk[123]) & (g134) & (g304) & (!g270) & (g136)) + ((sk[123]) & (g134) & (g304) & (g270) & (!g136)) + ((sk[123]) & (g134) & (g304) & (g270) & (g136)));
	assign g1386 = (((!sk[124]) & (g134) & (!g94) & (!g475)) + ((!sk[124]) & (g134) & (!g94) & (g475)) + ((!sk[124]) & (g134) & (g94) & (!g475)) + ((!sk[124]) & (g134) & (g94) & (g475)) + ((sk[124]) & (g134) & (!g94) & (!g475)) + ((sk[124]) & (g134) & (g94) & (!g475)) + ((sk[124]) & (g134) & (g94) & (g475)));
	assign g1387 = (((!g136) & (!g96) & (!g474) & (!sk[125]) & (!g1385) & (g1386)) + ((!g136) & (!g96) & (!g474) & (!sk[125]) & (g1385) & (g1386)) + ((!g136) & (!g96) & (!g474) & (sk[125]) & (!g1385) & (!g1386)) + ((!g136) & (!g96) & (g474) & (!sk[125]) & (!g1385) & (g1386)) + ((!g136) & (!g96) & (g474) & (!sk[125]) & (g1385) & (g1386)) + ((!g136) & (!g96) & (g474) & (sk[125]) & (!g1385) & (!g1386)) + ((!g136) & (g96) & (!g474) & (!sk[125]) & (!g1385) & (g1386)) + ((!g136) & (g96) & (!g474) & (!sk[125]) & (g1385) & (g1386)) + ((!g136) & (g96) & (!g474) & (sk[125]) & (!g1385) & (!g1386)) + ((!g136) & (g96) & (g474) & (!sk[125]) & (!g1385) & (g1386)) + ((!g136) & (g96) & (g474) & (!sk[125]) & (g1385) & (g1386)) + ((!g136) & (g96) & (g474) & (sk[125]) & (!g1385) & (!g1386)) + ((g136) & (!g96) & (!g474) & (!sk[125]) & (!g1385) & (!g1386)) + ((g136) & (!g96) & (!g474) & (!sk[125]) & (!g1385) & (g1386)) + ((g136) & (!g96) & (!g474) & (!sk[125]) & (g1385) & (!g1386)) + ((g136) & (!g96) & (!g474) & (!sk[125]) & (g1385) & (g1386)) + ((g136) & (!g96) & (g474) & (!sk[125]) & (!g1385) & (!g1386)) + ((g136) & (!g96) & (g474) & (!sk[125]) & (!g1385) & (g1386)) + ((g136) & (!g96) & (g474) & (!sk[125]) & (g1385) & (!g1386)) + ((g136) & (!g96) & (g474) & (!sk[125]) & (g1385) & (g1386)) + ((g136) & (g96) & (!g474) & (!sk[125]) & (!g1385) & (!g1386)) + ((g136) & (g96) & (!g474) & (!sk[125]) & (!g1385) & (g1386)) + ((g136) & (g96) & (!g474) & (!sk[125]) & (g1385) & (!g1386)) + ((g136) & (g96) & (!g474) & (!sk[125]) & (g1385) & (g1386)) + ((g136) & (g96) & (!g474) & (sk[125]) & (!g1385) & (!g1386)) + ((g136) & (g96) & (g474) & (!sk[125]) & (!g1385) & (!g1386)) + ((g136) & (g96) & (g474) & (!sk[125]) & (!g1385) & (g1386)) + ((g136) & (g96) & (g474) & (!sk[125]) & (g1385) & (!g1386)) + ((g136) & (g96) & (g474) & (!sk[125]) & (g1385) & (g1386)));
	assign g1388 = (((!g109) & (!g94) & (!sk[126]) & (g96) & (g678)) + ((!g109) & (g94) & (!sk[126]) & (!g96) & (!g678)) + ((!g109) & (g94) & (!sk[126]) & (!g96) & (g678)) + ((!g109) & (g94) & (!sk[126]) & (g96) & (!g678)) + ((!g109) & (g94) & (!sk[126]) & (g96) & (g678)) + ((g109) & (!g94) & (!sk[126]) & (g96) & (!g678)) + ((g109) & (!g94) & (!sk[126]) & (g96) & (g678)) + ((g109) & (!g94) & (sk[126]) & (!g96) & (!g678)) + ((g109) & (!g94) & (sk[126]) & (!g96) & (g678)) + ((g109) & (!g94) & (sk[126]) & (g96) & (!g678)) + ((g109) & (g94) & (!sk[126]) & (!g96) & (!g678)) + ((g109) & (g94) & (!sk[126]) & (!g96) & (g678)) + ((g109) & (g94) & (!sk[126]) & (g96) & (!g678)) + ((g109) & (g94) & (!sk[126]) & (g96) & (g678)) + ((g109) & (g94) & (sk[126]) & (!g96) & (!g678)) + ((g109) & (g94) & (sk[126]) & (!g96) & (g678)) + ((g109) & (g94) & (sk[126]) & (g96) & (!g678)) + ((g109) & (g94) & (sk[126]) & (g96) & (g678)));
	assign g1389 = (((!sk[127]) & (!i_8_) & (!g108) & (g96) & (g986)) + ((!sk[127]) & (!i_8_) & (g108) & (!g96) & (!g986)) + ((!sk[127]) & (!i_8_) & (g108) & (!g96) & (g986)) + ((!sk[127]) & (!i_8_) & (g108) & (g96) & (!g986)) + ((!sk[127]) & (!i_8_) & (g108) & (g96) & (g986)) + ((!sk[127]) & (i_8_) & (!g108) & (g96) & (!g986)) + ((!sk[127]) & (i_8_) & (!g108) & (g96) & (g986)) + ((!sk[127]) & (i_8_) & (g108) & (!g96) & (!g986)) + ((!sk[127]) & (i_8_) & (g108) & (!g96) & (g986)) + ((!sk[127]) & (i_8_) & (g108) & (g96) & (!g986)) + ((!sk[127]) & (i_8_) & (g108) & (g96) & (g986)) + ((sk[127]) & (!i_8_) & (g108) & (!g96) & (g986)) + ((sk[127]) & (!i_8_) & (g108) & (g96) & (g986)) + ((sk[127]) & (i_8_) & (g108) & (!g96) & (!g986)) + ((sk[127]) & (i_8_) & (g108) & (!g96) & (g986)) + ((sk[127]) & (i_8_) & (g108) & (g96) & (g986)));
	assign g1390 = (((!g109) & (!g203) & (!g183) & (!g268) & (!g1255) & (!g1389)) + ((!g109) & (!g203) & (!g183) & (!g268) & (g1255) & (!g1389)) + ((!g109) & (!g203) & (!g183) & (g268) & (!g1255) & (!g1389)) + ((!g109) & (!g203) & (!g183) & (g268) & (g1255) & (!g1389)) + ((!g109) & (!g203) & (g183) & (!g268) & (!g1255) & (!g1389)) + ((!g109) & (!g203) & (g183) & (!g268) & (g1255) & (!g1389)) + ((!g109) & (!g203) & (g183) & (g268) & (!g1255) & (!g1389)) + ((!g109) & (!g203) & (g183) & (g268) & (g1255) & (!g1389)) + ((!g109) & (g203) & (!g183) & (!g268) & (!g1255) & (!g1389)) + ((!g109) & (g203) & (!g183) & (!g268) & (g1255) & (!g1389)) + ((!g109) & (g203) & (!g183) & (g268) & (!g1255) & (!g1389)) + ((!g109) & (g203) & (!g183) & (g268) & (g1255) & (!g1389)) + ((!g109) & (g203) & (g183) & (!g268) & (!g1255) & (!g1389)) + ((!g109) & (g203) & (g183) & (!g268) & (g1255) & (!g1389)) + ((!g109) & (g203) & (g183) & (g268) & (!g1255) & (!g1389)) + ((!g109) & (g203) & (g183) & (g268) & (g1255) & (!g1389)) + ((g109) & (!g203) & (!g183) & (!g268) & (!g1255) & (!g1389)));
	assign g1391 = (((!i_14_) & (!i_12_) & (i_13_) & (!i_8_) & (g108) & (!g93)) + ((i_14_) & (i_12_) & (i_13_) & (i_8_) & (g108) & (!g93)));
	assign g1392 = (((!g510) & (!sk[2]) & (!g1388) & (!g1390) & (!g1538) & (g1391)) + ((!g510) & (!sk[2]) & (!g1388) & (!g1390) & (g1538) & (g1391)) + ((!g510) & (!sk[2]) & (!g1388) & (g1390) & (!g1538) & (g1391)) + ((!g510) & (!sk[2]) & (!g1388) & (g1390) & (g1538) & (g1391)) + ((!g510) & (!sk[2]) & (g1388) & (!g1390) & (!g1538) & (g1391)) + ((!g510) & (!sk[2]) & (g1388) & (!g1390) & (g1538) & (g1391)) + ((!g510) & (!sk[2]) & (g1388) & (g1390) & (!g1538) & (g1391)) + ((!g510) & (!sk[2]) & (g1388) & (g1390) & (g1538) & (g1391)) + ((!g510) & (sk[2]) & (!g1388) & (g1390) & (g1538) & (!g1391)) + ((g510) & (!sk[2]) & (!g1388) & (!g1390) & (!g1538) & (!g1391)) + ((g510) & (!sk[2]) & (!g1388) & (!g1390) & (!g1538) & (g1391)) + ((g510) & (!sk[2]) & (!g1388) & (!g1390) & (g1538) & (!g1391)) + ((g510) & (!sk[2]) & (!g1388) & (!g1390) & (g1538) & (g1391)) + ((g510) & (!sk[2]) & (!g1388) & (g1390) & (!g1538) & (!g1391)) + ((g510) & (!sk[2]) & (!g1388) & (g1390) & (!g1538) & (g1391)) + ((g510) & (!sk[2]) & (!g1388) & (g1390) & (g1538) & (!g1391)) + ((g510) & (!sk[2]) & (!g1388) & (g1390) & (g1538) & (g1391)) + ((g510) & (!sk[2]) & (g1388) & (!g1390) & (!g1538) & (!g1391)) + ((g510) & (!sk[2]) & (g1388) & (!g1390) & (!g1538) & (g1391)) + ((g510) & (!sk[2]) & (g1388) & (!g1390) & (g1538) & (!g1391)) + ((g510) & (!sk[2]) & (g1388) & (!g1390) & (g1538) & (g1391)) + ((g510) & (!sk[2]) & (g1388) & (g1390) & (!g1538) & (!g1391)) + ((g510) & (!sk[2]) & (g1388) & (g1390) & (!g1538) & (g1391)) + ((g510) & (!sk[2]) & (g1388) & (g1390) & (g1538) & (!g1391)) + ((g510) & (!sk[2]) & (g1388) & (g1390) & (g1538) & (g1391)));
	assign g1393 = (((!sk[3]) & (!g89) & (!g135) & (g268) & (g495)) + ((!sk[3]) & (!g89) & (g135) & (!g268) & (!g495)) + ((!sk[3]) & (!g89) & (g135) & (!g268) & (g495)) + ((!sk[3]) & (!g89) & (g135) & (g268) & (!g495)) + ((!sk[3]) & (!g89) & (g135) & (g268) & (g495)) + ((!sk[3]) & (g89) & (!g135) & (g268) & (!g495)) + ((!sk[3]) & (g89) & (!g135) & (g268) & (g495)) + ((!sk[3]) & (g89) & (g135) & (!g268) & (!g495)) + ((!sk[3]) & (g89) & (g135) & (!g268) & (g495)) + ((!sk[3]) & (g89) & (g135) & (g268) & (!g495)) + ((!sk[3]) & (g89) & (g135) & (g268) & (g495)) + ((sk[3]) & (!g89) & (!g135) & (g268) & (!g495)) + ((sk[3]) & (!g89) & (!g135) & (g268) & (g495)) + ((sk[3]) & (!g89) & (g135) & (g268) & (!g495)) + ((sk[3]) & (!g89) & (g135) & (g268) & (g495)) + ((sk[3]) & (g89) & (!g135) & (g268) & (g495)) + ((sk[3]) & (g89) & (g135) & (g268) & (!g495)) + ((sk[3]) & (g89) & (g135) & (g268) & (g495)));
	assign g1394 = (((g474) & (!sk[4]) & (!g495)) + ((g474) & (!sk[4]) & (g495)) + ((g474) & (sk[4]) & (g495)));
	assign g1395 = (((!sk[5]) & (!i_8_) & (!g270) & (g475) & (g495)) + ((!sk[5]) & (!i_8_) & (g270) & (!g475) & (!g495)) + ((!sk[5]) & (!i_8_) & (g270) & (!g475) & (g495)) + ((!sk[5]) & (!i_8_) & (g270) & (g475) & (!g495)) + ((!sk[5]) & (!i_8_) & (g270) & (g475) & (g495)) + ((!sk[5]) & (i_8_) & (!g270) & (g475) & (!g495)) + ((!sk[5]) & (i_8_) & (!g270) & (g475) & (g495)) + ((!sk[5]) & (i_8_) & (g270) & (!g475) & (!g495)) + ((!sk[5]) & (i_8_) & (g270) & (!g475) & (g495)) + ((!sk[5]) & (i_8_) & (g270) & (g475) & (!g495)) + ((!sk[5]) & (i_8_) & (g270) & (g475) & (g495)) + ((sk[5]) & (!i_8_) & (!g270) & (!g475) & (g495)) + ((sk[5]) & (!i_8_) & (g270) & (!g475) & (g495)) + ((sk[5]) & (i_8_) & (!g270) & (!g475) & (g495)) + ((sk[5]) & (i_8_) & (!g270) & (g475) & (g495)));
	assign g1396 = (((!g118) & (!g270) & (!sk[6]) & (g813) & (g495)) + ((!g118) & (!g270) & (sk[6]) & (g813) & (g495)) + ((!g118) & (g270) & (!sk[6]) & (!g813) & (!g495)) + ((!g118) & (g270) & (!sk[6]) & (!g813) & (g495)) + ((!g118) & (g270) & (!sk[6]) & (g813) & (!g495)) + ((!g118) & (g270) & (!sk[6]) & (g813) & (g495)) + ((!g118) & (g270) & (sk[6]) & (g813) & (g495)) + ((g118) & (!g270) & (!sk[6]) & (g813) & (!g495)) + ((g118) & (!g270) & (!sk[6]) & (g813) & (g495)) + ((g118) & (!g270) & (sk[6]) & (!g813) & (!g495)) + ((g118) & (!g270) & (sk[6]) & (!g813) & (g495)) + ((g118) & (!g270) & (sk[6]) & (g813) & (!g495)) + ((g118) & (!g270) & (sk[6]) & (g813) & (g495)) + ((g118) & (g270) & (!sk[6]) & (!g813) & (!g495)) + ((g118) & (g270) & (!sk[6]) & (!g813) & (g495)) + ((g118) & (g270) & (!sk[6]) & (g813) & (!g495)) + ((g118) & (g270) & (!sk[6]) & (g813) & (g495)) + ((g118) & (g270) & (sk[6]) & (g813) & (g495)));
	assign g1397 = (((!i_14_) & (!i_12_) & (!i_13_) & (g118) & (!g112) & (!g93)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g118) & (g112) & (!g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (!g118) & (g112) & (!g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (g118) & (!g112) & (!g93)) + ((!i_14_) & (i_12_) & (!i_13_) & (g118) & (g112) & (!g93)) + ((!i_14_) & (i_12_) & (i_13_) & (!g118) & (g112) & (!g93)) + ((!i_14_) & (i_12_) & (i_13_) & (g118) & (g112) & (!g93)) + ((i_14_) & (i_12_) & (!i_13_) & (!g118) & (g112) & (!g93)) + ((i_14_) & (i_12_) & (!i_13_) & (g118) & (!g112) & (!g93)) + ((i_14_) & (i_12_) & (!i_13_) & (g118) & (g112) & (!g93)));
	assign g1398 = (((!g659) & (!g682) & (!g1394) & (!g1395) & (!g1396) & (!g1397)));
	assign g1399 = (((!g118) & (!g423) & (!g429) & (!sk[9]) & (!g556) & (g1048)) + ((!g118) & (!g423) & (!g429) & (!sk[9]) & (g556) & (g1048)) + ((!g118) & (!g423) & (g429) & (!sk[9]) & (!g556) & (g1048)) + ((!g118) & (!g423) & (g429) & (!sk[9]) & (g556) & (g1048)) + ((!g118) & (!g423) & (g429) & (sk[9]) & (!g556) & (g1048)) + ((!g118) & (g423) & (!g429) & (!sk[9]) & (!g556) & (g1048)) + ((!g118) & (g423) & (!g429) & (!sk[9]) & (g556) & (g1048)) + ((!g118) & (g423) & (g429) & (!sk[9]) & (!g556) & (g1048)) + ((!g118) & (g423) & (g429) & (!sk[9]) & (g556) & (g1048)) + ((!g118) & (g423) & (g429) & (sk[9]) & (!g556) & (g1048)) + ((!g118) & (g423) & (g429) & (sk[9]) & (g556) & (g1048)) + ((g118) & (!g423) & (!g429) & (!sk[9]) & (!g556) & (!g1048)) + ((g118) & (!g423) & (!g429) & (!sk[9]) & (!g556) & (g1048)) + ((g118) & (!g423) & (!g429) & (!sk[9]) & (g556) & (!g1048)) + ((g118) & (!g423) & (!g429) & (!sk[9]) & (g556) & (g1048)) + ((g118) & (!g423) & (g429) & (!sk[9]) & (!g556) & (!g1048)) + ((g118) & (!g423) & (g429) & (!sk[9]) & (!g556) & (g1048)) + ((g118) & (!g423) & (g429) & (!sk[9]) & (g556) & (!g1048)) + ((g118) & (!g423) & (g429) & (!sk[9]) & (g556) & (g1048)) + ((g118) & (!g423) & (g429) & (sk[9]) & (!g556) & (!g1048)) + ((g118) & (!g423) & (g429) & (sk[9]) & (!g556) & (g1048)) + ((g118) & (g423) & (!g429) & (!sk[9]) & (!g556) & (!g1048)) + ((g118) & (g423) & (!g429) & (!sk[9]) & (!g556) & (g1048)) + ((g118) & (g423) & (!g429) & (!sk[9]) & (g556) & (!g1048)) + ((g118) & (g423) & (!g429) & (!sk[9]) & (g556) & (g1048)) + ((g118) & (g423) & (g429) & (!sk[9]) & (!g556) & (!g1048)) + ((g118) & (g423) & (g429) & (!sk[9]) & (!g556) & (g1048)) + ((g118) & (g423) & (g429) & (!sk[9]) & (g556) & (!g1048)) + ((g118) & (g423) & (g429) & (!sk[9]) & (g556) & (g1048)) + ((g118) & (g423) & (g429) & (sk[9]) & (!g556) & (!g1048)) + ((g118) & (g423) & (g429) & (sk[9]) & (!g556) & (g1048)) + ((g118) & (g423) & (g429) & (sk[9]) & (g556) & (g1048)));
	assign g1400 = (((!g983) & (!sk[10]) & (!g1393) & (g1398) & (g1399)) + ((!g983) & (!sk[10]) & (g1393) & (!g1398) & (!g1399)) + ((!g983) & (!sk[10]) & (g1393) & (!g1398) & (g1399)) + ((!g983) & (!sk[10]) & (g1393) & (g1398) & (!g1399)) + ((!g983) & (!sk[10]) & (g1393) & (g1398) & (g1399)) + ((g983) & (!sk[10]) & (!g1393) & (g1398) & (!g1399)) + ((g983) & (!sk[10]) & (!g1393) & (g1398) & (g1399)) + ((g983) & (!sk[10]) & (g1393) & (!g1398) & (!g1399)) + ((g983) & (!sk[10]) & (g1393) & (!g1398) & (g1399)) + ((g983) & (!sk[10]) & (g1393) & (g1398) & (!g1399)) + ((g983) & (!sk[10]) & (g1393) & (g1398) & (g1399)) + ((g983) & (sk[10]) & (!g1393) & (g1398) & (!g1399)));
	assign g1401 = (((!g145) & (!g268) & (!sk[11]) & (!g555) & (!g474) & (g678)) + ((!g145) & (!g268) & (!sk[11]) & (!g555) & (g474) & (g678)) + ((!g145) & (!g268) & (!sk[11]) & (g555) & (!g474) & (g678)) + ((!g145) & (!g268) & (!sk[11]) & (g555) & (g474) & (g678)) + ((!g145) & (g268) & (!sk[11]) & (!g555) & (!g474) & (g678)) + ((!g145) & (g268) & (!sk[11]) & (!g555) & (g474) & (g678)) + ((!g145) & (g268) & (!sk[11]) & (g555) & (!g474) & (g678)) + ((!g145) & (g268) & (!sk[11]) & (g555) & (g474) & (g678)) + ((g145) & (!g268) & (!sk[11]) & (!g555) & (!g474) & (!g678)) + ((g145) & (!g268) & (!sk[11]) & (!g555) & (!g474) & (g678)) + ((g145) & (!g268) & (!sk[11]) & (!g555) & (g474) & (!g678)) + ((g145) & (!g268) & (!sk[11]) & (!g555) & (g474) & (g678)) + ((g145) & (!g268) & (!sk[11]) & (g555) & (!g474) & (!g678)) + ((g145) & (!g268) & (!sk[11]) & (g555) & (!g474) & (g678)) + ((g145) & (!g268) & (!sk[11]) & (g555) & (g474) & (!g678)) + ((g145) & (!g268) & (!sk[11]) & (g555) & (g474) & (g678)) + ((g145) & (!g268) & (sk[11]) & (!g555) & (!g474) & (!g678)) + ((g145) & (!g268) & (sk[11]) & (!g555) & (g474) & (!g678)) + ((g145) & (!g268) & (sk[11]) & (!g555) & (g474) & (g678)) + ((g145) & (!g268) & (sk[11]) & (g555) & (!g474) & (!g678)) + ((g145) & (!g268) & (sk[11]) & (g555) & (!g474) & (g678)) + ((g145) & (!g268) & (sk[11]) & (g555) & (g474) & (!g678)) + ((g145) & (!g268) & (sk[11]) & (g555) & (g474) & (g678)) + ((g145) & (g268) & (!sk[11]) & (!g555) & (!g474) & (!g678)) + ((g145) & (g268) & (!sk[11]) & (!g555) & (!g474) & (g678)) + ((g145) & (g268) & (!sk[11]) & (!g555) & (g474) & (!g678)) + ((g145) & (g268) & (!sk[11]) & (!g555) & (g474) & (g678)) + ((g145) & (g268) & (!sk[11]) & (g555) & (!g474) & (!g678)) + ((g145) & (g268) & (!sk[11]) & (g555) & (!g474) & (g678)) + ((g145) & (g268) & (!sk[11]) & (g555) & (g474) & (!g678)) + ((g145) & (g268) & (!sk[11]) & (g555) & (g474) & (g678)) + ((g145) & (g268) & (sk[11]) & (!g555) & (!g474) & (!g678)) + ((g145) & (g268) & (sk[11]) & (!g555) & (!g474) & (g678)) + ((g145) & (g268) & (sk[11]) & (!g555) & (g474) & (!g678)) + ((g145) & (g268) & (sk[11]) & (!g555) & (g474) & (g678)) + ((g145) & (g268) & (sk[11]) & (g555) & (!g474) & (!g678)) + ((g145) & (g268) & (sk[11]) & (g555) & (!g474) & (g678)) + ((g145) & (g268) & (sk[11]) & (g555) & (g474) & (!g678)) + ((g145) & (g268) & (sk[11]) & (g555) & (g474) & (g678)));
	assign g1402 = (((!sk[12]) & (!g1002) & (!g1003) & (!g1004) & (!g1005) & (g1401)) + ((!sk[12]) & (!g1002) & (!g1003) & (!g1004) & (g1005) & (g1401)) + ((!sk[12]) & (!g1002) & (!g1003) & (g1004) & (!g1005) & (g1401)) + ((!sk[12]) & (!g1002) & (!g1003) & (g1004) & (g1005) & (g1401)) + ((!sk[12]) & (!g1002) & (g1003) & (!g1004) & (!g1005) & (g1401)) + ((!sk[12]) & (!g1002) & (g1003) & (!g1004) & (g1005) & (g1401)) + ((!sk[12]) & (!g1002) & (g1003) & (g1004) & (!g1005) & (g1401)) + ((!sk[12]) & (!g1002) & (g1003) & (g1004) & (g1005) & (g1401)) + ((!sk[12]) & (g1002) & (!g1003) & (!g1004) & (!g1005) & (!g1401)) + ((!sk[12]) & (g1002) & (!g1003) & (!g1004) & (!g1005) & (g1401)) + ((!sk[12]) & (g1002) & (!g1003) & (!g1004) & (g1005) & (!g1401)) + ((!sk[12]) & (g1002) & (!g1003) & (!g1004) & (g1005) & (g1401)) + ((!sk[12]) & (g1002) & (!g1003) & (g1004) & (!g1005) & (!g1401)) + ((!sk[12]) & (g1002) & (!g1003) & (g1004) & (!g1005) & (g1401)) + ((!sk[12]) & (g1002) & (!g1003) & (g1004) & (g1005) & (!g1401)) + ((!sk[12]) & (g1002) & (!g1003) & (g1004) & (g1005) & (g1401)) + ((!sk[12]) & (g1002) & (g1003) & (!g1004) & (!g1005) & (!g1401)) + ((!sk[12]) & (g1002) & (g1003) & (!g1004) & (!g1005) & (g1401)) + ((!sk[12]) & (g1002) & (g1003) & (!g1004) & (g1005) & (!g1401)) + ((!sk[12]) & (g1002) & (g1003) & (!g1004) & (g1005) & (g1401)) + ((!sk[12]) & (g1002) & (g1003) & (g1004) & (!g1005) & (!g1401)) + ((!sk[12]) & (g1002) & (g1003) & (g1004) & (!g1005) & (g1401)) + ((!sk[12]) & (g1002) & (g1003) & (g1004) & (g1005) & (!g1401)) + ((!sk[12]) & (g1002) & (g1003) & (g1004) & (g1005) & (g1401)) + ((sk[12]) & (!g1002) & (!g1003) & (!g1004) & (!g1005) & (!g1401)));
	assign g1403 = (((!sk[13]) & (g118) & (!g214) & (!g756)) + ((!sk[13]) & (g118) & (!g214) & (g756)) + ((!sk[13]) & (g118) & (g214) & (!g756)) + ((!sk[13]) & (g118) & (g214) & (g756)) + ((sk[13]) & (!g118) & (g214) & (g756)) + ((sk[13]) & (g118) & (!g214) & (g756)) + ((sk[13]) & (g118) & (g214) & (g756)));
	assign g1404 = (((!g7) & (!g95) & (!g461) & (sk[14]) & (!g756)) + ((!g7) & (!g95) & (g461) & (!sk[14]) & (g756)) + ((!g7) & (!g95) & (g461) & (sk[14]) & (!g756)) + ((!g7) & (g95) & (!g461) & (!sk[14]) & (!g756)) + ((!g7) & (g95) & (!g461) & (!sk[14]) & (g756)) + ((!g7) & (g95) & (!g461) & (sk[14]) & (!g756)) + ((!g7) & (g95) & (g461) & (!sk[14]) & (!g756)) + ((!g7) & (g95) & (g461) & (!sk[14]) & (g756)) + ((g7) & (!g95) & (!g461) & (sk[14]) & (!g756)) + ((g7) & (!g95) & (g461) & (!sk[14]) & (!g756)) + ((g7) & (!g95) & (g461) & (!sk[14]) & (g756)) + ((g7) & (!g95) & (g461) & (sk[14]) & (!g756)) + ((g7) & (g95) & (!g461) & (!sk[14]) & (!g756)) + ((g7) & (g95) & (!g461) & (!sk[14]) & (g756)) + ((g7) & (g95) & (g461) & (!sk[14]) & (!g756)) + ((g7) & (g95) & (g461) & (!sk[14]) & (g756)));
	assign g1405 = (((!g99) & (!g330) & (!g251) & (!g986) & (!g1403) & (g1404)) + ((!g99) & (!g330) & (!g251) & (!g986) & (g1403) & (g1404)) + ((!g99) & (!g330) & (!g251) & (g986) & (!g1403) & (g1404)) + ((!g99) & (!g330) & (!g251) & (g986) & (g1403) & (g1404)) + ((!g99) & (!g330) & (g251) & (!g986) & (!g1403) & (g1404)) + ((!g99) & (!g330) & (g251) & (!g986) & (g1403) & (g1404)) + ((!g99) & (g330) & (!g251) & (!g986) & (!g1403) & (!g1404)) + ((!g99) & (g330) & (!g251) & (!g986) & (!g1403) & (g1404)) + ((!g99) & (g330) & (!g251) & (!g986) & (g1403) & (g1404)) + ((!g99) & (g330) & (!g251) & (g986) & (!g1403) & (!g1404)) + ((!g99) & (g330) & (!g251) & (g986) & (!g1403) & (g1404)) + ((!g99) & (g330) & (!g251) & (g986) & (g1403) & (g1404)) + ((!g99) & (g330) & (g251) & (!g986) & (!g1403) & (!g1404)) + ((!g99) & (g330) & (g251) & (!g986) & (!g1403) & (g1404)) + ((!g99) & (g330) & (g251) & (!g986) & (g1403) & (g1404)) + ((g99) & (!g330) & (!g251) & (!g986) & (!g1403) & (g1404)) + ((g99) & (!g330) & (!g251) & (!g986) & (g1403) & (g1404)) + ((g99) & (!g330) & (g251) & (!g986) & (!g1403) & (g1404)) + ((g99) & (!g330) & (g251) & (!g986) & (g1403) & (g1404)) + ((g99) & (g330) & (!g251) & (!g986) & (!g1403) & (!g1404)) + ((g99) & (g330) & (!g251) & (!g986) & (!g1403) & (g1404)) + ((g99) & (g330) & (!g251) & (!g986) & (g1403) & (g1404)) + ((g99) & (g330) & (g251) & (!g986) & (!g1403) & (!g1404)) + ((g99) & (g330) & (g251) & (!g986) & (!g1403) & (g1404)) + ((g99) & (g330) & (g251) & (!g986) & (g1403) & (g1404)));
	assign g1406 = (((!g212) & (!g213) & (!g215) & (!g217) & (!sk[16]) & (g1036)) + ((!g212) & (!g213) & (!g215) & (!g217) & (sk[16]) & (!g1036)) + ((!g212) & (!g213) & (!g215) & (g217) & (!sk[16]) & (g1036)) + ((!g212) & (!g213) & (g215) & (!g217) & (!sk[16]) & (g1036)) + ((!g212) & (!g213) & (g215) & (!g217) & (sk[16]) & (!g1036)) + ((!g212) & (!g213) & (g215) & (g217) & (!sk[16]) & (g1036)) + ((!g212) & (g213) & (!g215) & (!g217) & (!sk[16]) & (g1036)) + ((!g212) & (g213) & (!g215) & (g217) & (!sk[16]) & (g1036)) + ((!g212) & (g213) & (g215) & (!g217) & (!sk[16]) & (g1036)) + ((!g212) & (g213) & (g215) & (g217) & (!sk[16]) & (g1036)) + ((g212) & (!g213) & (!g215) & (!g217) & (!sk[16]) & (!g1036)) + ((g212) & (!g213) & (!g215) & (!g217) & (!sk[16]) & (g1036)) + ((g212) & (!g213) & (!g215) & (!g217) & (sk[16]) & (!g1036)) + ((g212) & (!g213) & (!g215) & (g217) & (!sk[16]) & (!g1036)) + ((g212) & (!g213) & (!g215) & (g217) & (!sk[16]) & (g1036)) + ((g212) & (!g213) & (g215) & (!g217) & (!sk[16]) & (!g1036)) + ((g212) & (!g213) & (g215) & (!g217) & (!sk[16]) & (g1036)) + ((g212) & (!g213) & (g215) & (!g217) & (sk[16]) & (!g1036)) + ((g212) & (!g213) & (g215) & (g217) & (!sk[16]) & (!g1036)) + ((g212) & (!g213) & (g215) & (g217) & (!sk[16]) & (g1036)) + ((g212) & (g213) & (!g215) & (!g217) & (!sk[16]) & (!g1036)) + ((g212) & (g213) & (!g215) & (!g217) & (!sk[16]) & (g1036)) + ((g212) & (g213) & (!g215) & (g217) & (!sk[16]) & (!g1036)) + ((g212) & (g213) & (!g215) & (g217) & (!sk[16]) & (g1036)) + ((g212) & (g213) & (g215) & (!g217) & (!sk[16]) & (!g1036)) + ((g212) & (g213) & (g215) & (!g217) & (!sk[16]) & (g1036)) + ((g212) & (g213) & (g215) & (!g217) & (sk[16]) & (!g1036)) + ((g212) & (g213) & (g215) & (g217) & (!sk[16]) & (!g1036)) + ((g212) & (g213) & (g215) & (g217) & (!sk[16]) & (g1036)));
	assign g1407 = (((!i_8_) & (!g88) & (!g212) & (!g534) & (g555) & (!g1099)) + ((!i_8_) & (!g88) & (!g212) & (!g534) & (g555) & (g1099)) + ((!i_8_) & (!g88) & (!g212) & (g534) & (g555) & (!g1099)) + ((!i_8_) & (!g88) & (!g212) & (g534) & (g555) & (g1099)) + ((!i_8_) & (g88) & (!g212) & (!g534) & (g555) & (!g1099)) + ((!i_8_) & (g88) & (!g212) & (!g534) & (g555) & (g1099)) + ((!i_8_) & (g88) & (!g212) & (g534) & (g555) & (!g1099)) + ((!i_8_) & (g88) & (!g212) & (g534) & (g555) & (g1099)) + ((!i_8_) & (g88) & (g212) & (!g534) & (g555) & (!g1099)) + ((!i_8_) & (g88) & (g212) & (!g534) & (g555) & (g1099)) + ((!i_8_) & (g88) & (g212) & (g534) & (g555) & (!g1099)) + ((!i_8_) & (g88) & (g212) & (g534) & (g555) & (g1099)) + ((i_8_) & (!g88) & (!g212) & (!g534) & (g555) & (!g1099)) + ((i_8_) & (!g88) & (!g212) & (!g534) & (g555) & (g1099)) + ((i_8_) & (!g88) & (!g212) & (g534) & (g555) & (!g1099)) + ((i_8_) & (!g88) & (!g212) & (g534) & (g555) & (g1099)) + ((i_8_) & (g88) & (!g212) & (!g534) & (!g555) & (!g1099)) + ((i_8_) & (g88) & (!g212) & (!g534) & (g555) & (!g1099)) + ((i_8_) & (g88) & (!g212) & (!g534) & (g555) & (g1099)) + ((i_8_) & (g88) & (!g212) & (g534) & (!g555) & (!g1099)) + ((i_8_) & (g88) & (!g212) & (g534) & (!g555) & (g1099)) + ((i_8_) & (g88) & (!g212) & (g534) & (g555) & (!g1099)) + ((i_8_) & (g88) & (!g212) & (g534) & (g555) & (g1099)) + ((i_8_) & (g88) & (g212) & (!g534) & (!g555) & (!g1099)) + ((i_8_) & (g88) & (g212) & (!g534) & (g555) & (!g1099)) + ((i_8_) & (g88) & (g212) & (g534) & (!g555) & (!g1099)) + ((i_8_) & (g88) & (g212) & (g534) & (!g555) & (g1099)) + ((i_8_) & (g88) & (g212) & (g534) & (g555) & (!g1099)) + ((i_8_) & (g88) & (g212) & (g534) & (g555) & (g1099)));
	assign g1408 = (((!g99) & (!g88) & (g554) & (!sk[18]) & (g895)) + ((!g99) & (g88) & (!g554) & (!sk[18]) & (!g895)) + ((!g99) & (g88) & (!g554) & (!sk[18]) & (g895)) + ((!g99) & (g88) & (g554) & (!sk[18]) & (!g895)) + ((!g99) & (g88) & (g554) & (!sk[18]) & (g895)) + ((!g99) & (g88) & (g554) & (sk[18]) & (!g895)) + ((!g99) & (g88) & (g554) & (sk[18]) & (g895)) + ((g99) & (!g88) & (!g554) & (sk[18]) & (g895)) + ((g99) & (!g88) & (g554) & (!sk[18]) & (!g895)) + ((g99) & (!g88) & (g554) & (!sk[18]) & (g895)) + ((g99) & (!g88) & (g554) & (sk[18]) & (g895)) + ((g99) & (g88) & (!g554) & (!sk[18]) & (!g895)) + ((g99) & (g88) & (!g554) & (!sk[18]) & (g895)) + ((g99) & (g88) & (!g554) & (sk[18]) & (g895)) + ((g99) & (g88) & (g554) & (!sk[18]) & (!g895)) + ((g99) & (g88) & (g554) & (!sk[18]) & (g895)) + ((g99) & (g88) & (g554) & (sk[18]) & (!g895)) + ((g99) & (g88) & (g554) & (sk[18]) & (g895)));
	assign g1409 = (((!g99) & (!g101) & (!g756) & (!g991) & (!g1042) & (!g1408)) + ((!g99) & (!g101) & (g756) & (!g991) & (!g1042) & (!g1408)) + ((!g99) & (g101) & (!g756) & (!g991) & (!g1042) & (!g1408)) + ((g99) & (!g101) & (!g756) & (!g991) & (!g1042) & (!g1408)) + ((g99) & (g101) & (!g756) & (!g991) & (!g1042) & (!g1408)));
	assign g1410 = (((!g149) & (!g338) & (!g341) & (g556) & (!g522) & (!g476)) + ((!g149) & (g338) & (!g341) & (!g556) & (!g522) & (!g476)) + ((!g149) & (g338) & (!g341) & (!g556) & (g522) & (!g476)) + ((!g149) & (g338) & (!g341) & (g556) & (!g522) & (!g476)) + ((!g149) & (g338) & (!g341) & (g556) & (g522) & (!g476)) + ((g149) & (!g338) & (!g341) & (g556) & (!g522) & (!g476)) + ((g149) & (g338) & (!g341) & (!g556) & (!g522) & (!g476)) + ((g149) & (g338) & (!g341) & (g556) & (!g522) & (!g476)));
	assign g1411 = (((i_8_) & (g100) & (!g199) & (!g120) & (!g547) & (!g574)) + ((i_8_) & (g100) & (!g199) & (!g120) & (!g547) & (g574)) + ((i_8_) & (g100) & (!g199) & (!g120) & (g547) & (!g574)) + ((i_8_) & (g100) & (!g199) & (!g120) & (g547) & (g574)) + ((i_8_) & (g100) & (!g199) & (g120) & (!g547) & (!g574)) + ((i_8_) & (g100) & (!g199) & (g120) & (!g547) & (g574)) + ((i_8_) & (g100) & (!g199) & (g120) & (g547) & (g574)) + ((i_8_) & (g100) & (g199) & (!g120) & (!g547) & (!g574)) + ((i_8_) & (g100) & (g199) & (!g120) & (!g547) & (g574)) + ((i_8_) & (g100) & (g199) & (!g120) & (g547) & (!g574)) + ((i_8_) & (g100) & (g199) & (!g120) & (g547) & (g574)) + ((i_8_) & (g100) & (g199) & (g120) & (!g547) & (!g574)) + ((i_8_) & (g100) & (g199) & (g120) & (!g547) & (g574)) + ((i_8_) & (g100) & (g199) & (g120) & (g547) & (!g574)) + ((i_8_) & (g100) & (g199) & (g120) & (g547) & (g574)));
	assign g1412 = (((g1405) & (g1406) & (!g1407) & (g1409) & (g1410) & (!g1558)));
	assign g1413 = (((g527) & (g1110) & (g1059) & (g1400) & (g1402) & (g1412)));
	assign o_19_ = (((g73) & (!g1301) & (!g1341) & (!g1568) & (!g1392) & (!g1413)) + ((g73) & (!g1301) & (!g1341) & (!g1568) & (!g1392) & (g1413)) + ((g73) & (!g1301) & (!g1341) & (!g1568) & (g1392) & (!g1413)) + ((g73) & (!g1301) & (!g1341) & (!g1568) & (g1392) & (g1413)) + ((g73) & (!g1301) & (!g1341) & (g1568) & (!g1392) & (!g1413)) + ((g73) & (!g1301) & (!g1341) & (g1568) & (!g1392) & (g1413)) + ((g73) & (!g1301) & (!g1341) & (g1568) & (g1392) & (!g1413)) + ((g73) & (!g1301) & (!g1341) & (g1568) & (g1392) & (g1413)) + ((g73) & (!g1301) & (g1341) & (!g1568) & (!g1392) & (!g1413)) + ((g73) & (!g1301) & (g1341) & (!g1568) & (!g1392) & (g1413)) + ((g73) & (!g1301) & (g1341) & (!g1568) & (g1392) & (!g1413)) + ((g73) & (!g1301) & (g1341) & (!g1568) & (g1392) & (g1413)) + ((g73) & (!g1301) & (g1341) & (g1568) & (!g1392) & (!g1413)) + ((g73) & (!g1301) & (g1341) & (g1568) & (!g1392) & (g1413)) + ((g73) & (!g1301) & (g1341) & (g1568) & (g1392) & (!g1413)) + ((g73) & (!g1301) & (g1341) & (g1568) & (g1392) & (g1413)) + ((g73) & (g1301) & (!g1341) & (!g1568) & (!g1392) & (!g1413)) + ((g73) & (g1301) & (!g1341) & (!g1568) & (!g1392) & (g1413)) + ((g73) & (g1301) & (!g1341) & (!g1568) & (g1392) & (!g1413)) + ((g73) & (g1301) & (!g1341) & (!g1568) & (g1392) & (g1413)) + ((g73) & (g1301) & (!g1341) & (g1568) & (!g1392) & (!g1413)) + ((g73) & (g1301) & (!g1341) & (g1568) & (!g1392) & (g1413)) + ((g73) & (g1301) & (!g1341) & (g1568) & (g1392) & (!g1413)) + ((g73) & (g1301) & (!g1341) & (g1568) & (g1392) & (g1413)) + ((g73) & (g1301) & (g1341) & (!g1568) & (!g1392) & (!g1413)) + ((g73) & (g1301) & (g1341) & (!g1568) & (!g1392) & (g1413)) + ((g73) & (g1301) & (g1341) & (!g1568) & (g1392) & (!g1413)) + ((g73) & (g1301) & (g1341) & (!g1568) & (g1392) & (g1413)) + ((g73) & (g1301) & (g1341) & (g1568) & (!g1392) & (!g1413)) + ((g73) & (g1301) & (g1341) & (g1568) & (!g1392) & (g1413)) + ((g73) & (g1301) & (g1341) & (g1568) & (g1392) & (!g1413)));
	assign g1415 = (((!g1305) & (sk[25]) & (g1314) & (g1317)) + ((g1305) & (!sk[25]) & (!g1314) & (!g1317)) + ((g1305) & (!sk[25]) & (!g1314) & (g1317)) + ((g1305) & (!sk[25]) & (g1314) & (!g1317)) + ((g1305) & (!sk[25]) & (g1314) & (g1317)));
	assign g1416 = (((!i_8_) & (!sk[26]) & (!g222) & (g531) & (g630)) + ((!i_8_) & (!sk[26]) & (g222) & (!g531) & (!g630)) + ((!i_8_) & (!sk[26]) & (g222) & (!g531) & (g630)) + ((!i_8_) & (!sk[26]) & (g222) & (g531) & (!g630)) + ((!i_8_) & (!sk[26]) & (g222) & (g531) & (g630)) + ((!i_8_) & (sk[26]) & (!g222) & (!g531) & (!g630)) + ((i_8_) & (!sk[26]) & (!g222) & (g531) & (!g630)) + ((i_8_) & (!sk[26]) & (!g222) & (g531) & (g630)) + ((i_8_) & (!sk[26]) & (g222) & (!g531) & (!g630)) + ((i_8_) & (!sk[26]) & (g222) & (!g531) & (g630)) + ((i_8_) & (!sk[26]) & (g222) & (g531) & (!g630)) + ((i_8_) & (!sk[26]) & (g222) & (g531) & (g630)));
	assign g1417 = (((!g246) & (!g593) & (g678) & (!sk[27]) & (g1416)) + ((!g246) & (g593) & (!g678) & (!sk[27]) & (!g1416)) + ((!g246) & (g593) & (!g678) & (!sk[27]) & (g1416)) + ((!g246) & (g593) & (g678) & (!sk[27]) & (!g1416)) + ((!g246) & (g593) & (g678) & (!sk[27]) & (g1416)) + ((!g246) & (g593) & (g678) & (sk[27]) & (g1416)) + ((g246) & (!g593) & (g678) & (!sk[27]) & (!g1416)) + ((g246) & (!g593) & (g678) & (!sk[27]) & (g1416)) + ((g246) & (g593) & (!g678) & (!sk[27]) & (!g1416)) + ((g246) & (g593) & (!g678) & (!sk[27]) & (g1416)) + ((g246) & (g593) & (g678) & (!sk[27]) & (!g1416)) + ((g246) & (g593) & (g678) & (!sk[27]) & (g1416)));
	assign g1418 = (((!g339) & (!g613) & (!g465) & (!g506) & (!sk[28]) & (g1417)) + ((!g339) & (!g613) & (!g465) & (g506) & (!sk[28]) & (g1417)) + ((!g339) & (!g613) & (g465) & (!g506) & (!sk[28]) & (g1417)) + ((!g339) & (!g613) & (g465) & (g506) & (!sk[28]) & (g1417)) + ((!g339) & (g613) & (!g465) & (!g506) & (!sk[28]) & (g1417)) + ((!g339) & (g613) & (!g465) & (g506) & (!sk[28]) & (g1417)) + ((!g339) & (g613) & (g465) & (!g506) & (!sk[28]) & (g1417)) + ((!g339) & (g613) & (g465) & (!g506) & (sk[28]) & (g1417)) + ((!g339) & (g613) & (g465) & (g506) & (!sk[28]) & (g1417)) + ((g339) & (!g613) & (!g465) & (!g506) & (!sk[28]) & (!g1417)) + ((g339) & (!g613) & (!g465) & (!g506) & (!sk[28]) & (g1417)) + ((g339) & (!g613) & (!g465) & (g506) & (!sk[28]) & (!g1417)) + ((g339) & (!g613) & (!g465) & (g506) & (!sk[28]) & (g1417)) + ((g339) & (!g613) & (g465) & (!g506) & (!sk[28]) & (!g1417)) + ((g339) & (!g613) & (g465) & (!g506) & (!sk[28]) & (g1417)) + ((g339) & (!g613) & (g465) & (g506) & (!sk[28]) & (!g1417)) + ((g339) & (!g613) & (g465) & (g506) & (!sk[28]) & (g1417)) + ((g339) & (g613) & (!g465) & (!g506) & (!sk[28]) & (!g1417)) + ((g339) & (g613) & (!g465) & (!g506) & (!sk[28]) & (g1417)) + ((g339) & (g613) & (!g465) & (g506) & (!sk[28]) & (!g1417)) + ((g339) & (g613) & (!g465) & (g506) & (!sk[28]) & (g1417)) + ((g339) & (g613) & (g465) & (!g506) & (!sk[28]) & (!g1417)) + ((g339) & (g613) & (g465) & (!g506) & (!sk[28]) & (g1417)) + ((g339) & (g613) & (g465) & (g506) & (!sk[28]) & (!g1417)) + ((g339) & (g613) & (g465) & (g506) & (!sk[28]) & (g1417)));
	assign g1419 = (((!g6) & (!sk[29]) & (!i_15_) & (g7) & (g461)) + ((!g6) & (!sk[29]) & (i_15_) & (!g7) & (!g461)) + ((!g6) & (!sk[29]) & (i_15_) & (!g7) & (g461)) + ((!g6) & (!sk[29]) & (i_15_) & (g7) & (!g461)) + ((!g6) & (!sk[29]) & (i_15_) & (g7) & (g461)) + ((g6) & (!sk[29]) & (!i_15_) & (g7) & (!g461)) + ((g6) & (!sk[29]) & (!i_15_) & (g7) & (g461)) + ((g6) & (!sk[29]) & (i_15_) & (!g7) & (!g461)) + ((g6) & (!sk[29]) & (i_15_) & (!g7) & (g461)) + ((g6) & (!sk[29]) & (i_15_) & (g7) & (!g461)) + ((g6) & (!sk[29]) & (i_15_) & (g7) & (g461)) + ((g6) & (sk[29]) & (!i_15_) & (!g7) & (g461)) + ((g6) & (sk[29]) & (!i_15_) & (g7) & (!g461)) + ((g6) & (sk[29]) & (!i_15_) & (g7) & (g461)));
	assign g1420 = (((!i_8_) & (!g495) & (!g1026) & (!g1111) & (!sk[30]) & (g1419)) + ((!i_8_) & (!g495) & (!g1026) & (g1111) & (!sk[30]) & (g1419)) + ((!i_8_) & (!g495) & (g1026) & (!g1111) & (!sk[30]) & (g1419)) + ((!i_8_) & (!g495) & (g1026) & (g1111) & (!sk[30]) & (g1419)) + ((!i_8_) & (g495) & (!g1026) & (!g1111) & (!sk[30]) & (g1419)) + ((!i_8_) & (g495) & (!g1026) & (!g1111) & (sk[30]) & (!g1419)) + ((!i_8_) & (g495) & (!g1026) & (!g1111) & (sk[30]) & (g1419)) + ((!i_8_) & (g495) & (!g1026) & (g1111) & (!sk[30]) & (g1419)) + ((!i_8_) & (g495) & (!g1026) & (g1111) & (sk[30]) & (!g1419)) + ((!i_8_) & (g495) & (!g1026) & (g1111) & (sk[30]) & (g1419)) + ((!i_8_) & (g495) & (g1026) & (!g1111) & (!sk[30]) & (g1419)) + ((!i_8_) & (g495) & (g1026) & (!g1111) & (sk[30]) & (!g1419)) + ((!i_8_) & (g495) & (g1026) & (!g1111) & (sk[30]) & (g1419)) + ((!i_8_) & (g495) & (g1026) & (g1111) & (!sk[30]) & (g1419)) + ((!i_8_) & (g495) & (g1026) & (g1111) & (sk[30]) & (!g1419)) + ((!i_8_) & (g495) & (g1026) & (g1111) & (sk[30]) & (g1419)) + ((i_8_) & (!g495) & (!g1026) & (!g1111) & (!sk[30]) & (!g1419)) + ((i_8_) & (!g495) & (!g1026) & (!g1111) & (!sk[30]) & (g1419)) + ((i_8_) & (!g495) & (!g1026) & (g1111) & (!sk[30]) & (!g1419)) + ((i_8_) & (!g495) & (!g1026) & (g1111) & (!sk[30]) & (g1419)) + ((i_8_) & (!g495) & (g1026) & (!g1111) & (!sk[30]) & (!g1419)) + ((i_8_) & (!g495) & (g1026) & (!g1111) & (!sk[30]) & (g1419)) + ((i_8_) & (!g495) & (g1026) & (g1111) & (!sk[30]) & (!g1419)) + ((i_8_) & (!g495) & (g1026) & (g1111) & (!sk[30]) & (g1419)) + ((i_8_) & (g495) & (!g1026) & (!g1111) & (!sk[30]) & (!g1419)) + ((i_8_) & (g495) & (!g1026) & (!g1111) & (!sk[30]) & (g1419)) + ((i_8_) & (g495) & (!g1026) & (!g1111) & (sk[30]) & (!g1419)) + ((i_8_) & (g495) & (!g1026) & (!g1111) & (sk[30]) & (g1419)) + ((i_8_) & (g495) & (!g1026) & (g1111) & (!sk[30]) & (!g1419)) + ((i_8_) & (g495) & (!g1026) & (g1111) & (!sk[30]) & (g1419)) + ((i_8_) & (g495) & (!g1026) & (g1111) & (sk[30]) & (g1419)) + ((i_8_) & (g495) & (g1026) & (!g1111) & (!sk[30]) & (!g1419)) + ((i_8_) & (g495) & (g1026) & (!g1111) & (!sk[30]) & (g1419)) + ((i_8_) & (g495) & (g1026) & (!g1111) & (sk[30]) & (!g1419)) + ((i_8_) & (g495) & (g1026) & (!g1111) & (sk[30]) & (g1419)) + ((i_8_) & (g495) & (g1026) & (g1111) & (!sk[30]) & (!g1419)) + ((i_8_) & (g495) & (g1026) & (g1111) & (!sk[30]) & (g1419)) + ((i_8_) & (g495) & (g1026) & (g1111) & (sk[30]) & (!g1419)) + ((i_8_) & (g495) & (g1026) & (g1111) & (sk[30]) & (g1419)));
	assign g1421 = (((!sk[31]) & (!g1112) & (!g1113) & (g1418) & (g1420)) + ((!sk[31]) & (!g1112) & (g1113) & (!g1418) & (!g1420)) + ((!sk[31]) & (!g1112) & (g1113) & (!g1418) & (g1420)) + ((!sk[31]) & (!g1112) & (g1113) & (g1418) & (!g1420)) + ((!sk[31]) & (!g1112) & (g1113) & (g1418) & (g1420)) + ((!sk[31]) & (g1112) & (!g1113) & (g1418) & (!g1420)) + ((!sk[31]) & (g1112) & (!g1113) & (g1418) & (g1420)) + ((!sk[31]) & (g1112) & (g1113) & (!g1418) & (!g1420)) + ((!sk[31]) & (g1112) & (g1113) & (!g1418) & (g1420)) + ((!sk[31]) & (g1112) & (g1113) & (g1418) & (!g1420)) + ((!sk[31]) & (g1112) & (g1113) & (g1418) & (g1420)) + ((sk[31]) & (!g1112) & (!g1113) & (!g1418) & (g1420)) + ((sk[31]) & (!g1112) & (!g1113) & (g1418) & (g1420)) + ((sk[31]) & (!g1112) & (g1113) & (!g1418) & (g1420)) + ((sk[31]) & (!g1112) & (g1113) & (g1418) & (g1420)) + ((sk[31]) & (g1112) & (!g1113) & (!g1418) & (g1420)) + ((sk[31]) & (g1112) & (!g1113) & (g1418) & (g1420)) + ((sk[31]) & (g1112) & (g1113) & (!g1418) & (g1420)));
	assign g1422 = (((!sk[32]) & (g1238) & (!g1270) & (!g1272)) + ((!sk[32]) & (g1238) & (!g1270) & (g1272)) + ((!sk[32]) & (g1238) & (g1270) & (!g1272)) + ((!sk[32]) & (g1238) & (g1270) & (g1272)) + ((sk[32]) & (g1238) & (!g1270) & (g1272)));
	assign g1423 = (((!g237) & (!sk[33]) & (!g661) & (g1224) & (g1200)) + ((!g237) & (!sk[33]) & (g661) & (!g1224) & (!g1200)) + ((!g237) & (!sk[33]) & (g661) & (!g1224) & (g1200)) + ((!g237) & (!sk[33]) & (g661) & (g1224) & (!g1200)) + ((!g237) & (!sk[33]) & (g661) & (g1224) & (g1200)) + ((!g237) & (sk[33]) & (!g661) & (!g1224) & (!g1200)) + ((g237) & (!sk[33]) & (!g661) & (g1224) & (!g1200)) + ((g237) & (!sk[33]) & (!g661) & (g1224) & (g1200)) + ((g237) & (!sk[33]) & (g661) & (!g1224) & (!g1200)) + ((g237) & (!sk[33]) & (g661) & (!g1224) & (g1200)) + ((g237) & (!sk[33]) & (g661) & (g1224) & (!g1200)) + ((g237) & (!sk[33]) & (g661) & (g1224) & (g1200)));
	assign g1424 = (((!g43) & (!sk[34]) & (!g495) & (g1122) & (g1296)) + ((!g43) & (!sk[34]) & (g495) & (!g1122) & (!g1296)) + ((!g43) & (!sk[34]) & (g495) & (!g1122) & (g1296)) + ((!g43) & (!sk[34]) & (g495) & (g1122) & (!g1296)) + ((!g43) & (!sk[34]) & (g495) & (g1122) & (g1296)) + ((!g43) & (sk[34]) & (!g495) & (!g1122) & (!g1296)) + ((!g43) & (sk[34]) & (!g495) & (g1122) & (!g1296)) + ((!g43) & (sk[34]) & (g495) & (g1122) & (!g1296)) + ((g43) & (!sk[34]) & (!g495) & (g1122) & (!g1296)) + ((g43) & (!sk[34]) & (!g495) & (g1122) & (g1296)) + ((g43) & (!sk[34]) & (g495) & (!g1122) & (!g1296)) + ((g43) & (!sk[34]) & (g495) & (!g1122) & (g1296)) + ((g43) & (!sk[34]) & (g495) & (g1122) & (!g1296)) + ((g43) & (!sk[34]) & (g495) & (g1122) & (g1296)) + ((g43) & (sk[34]) & (!g495) & (!g1122) & (!g1296)) + ((g43) & (sk[34]) & (!g495) & (g1122) & (!g1296)));
	assign g1425 = (((!i_14_) & (!i_12_) & (!i_13_) & (g112) & (!g131) & (g158)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g112) & (g131) & (g158)) + ((!i_14_) & (!i_12_) & (i_13_) & (g112) & (!g131) & (g158)) + ((!i_14_) & (!i_12_) & (i_13_) & (g112) & (g131) & (!g158)) + ((!i_14_) & (!i_12_) & (i_13_) & (g112) & (g131) & (g158)) + ((!i_14_) & (i_12_) & (!i_13_) & (g112) & (!g131) & (g158)) + ((!i_14_) & (i_12_) & (!i_13_) & (g112) & (g131) & (!g158)) + ((!i_14_) & (i_12_) & (!i_13_) & (g112) & (g131) & (g158)) + ((!i_14_) & (i_12_) & (i_13_) & (g112) & (!g131) & (g158)) + ((!i_14_) & (i_12_) & (i_13_) & (g112) & (g131) & (!g158)) + ((!i_14_) & (i_12_) & (i_13_) & (g112) & (g131) & (g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (g112) & (!g131) & (g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (g112) & (g131) & (!g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (g112) & (g131) & (g158)) + ((i_14_) & (!i_12_) & (i_13_) & (g112) & (!g131) & (g158)) + ((i_14_) & (!i_12_) & (i_13_) & (g112) & (g131) & (!g158)) + ((i_14_) & (!i_12_) & (i_13_) & (g112) & (g131) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (g112) & (!g131) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (g112) & (g131) & (g158)) + ((i_14_) & (i_12_) & (i_13_) & (g112) & (g131) & (!g158)) + ((i_14_) & (i_12_) & (i_13_) & (g112) & (g131) & (g158)));
	assign g1426 = (((!g8) & (!g10) & (!g112) & (!g1174) & (!sk[36]) & (g1425)) + ((!g8) & (!g10) & (!g112) & (!g1174) & (sk[36]) & (!g1425)) + ((!g8) & (!g10) & (!g112) & (g1174) & (!sk[36]) & (g1425)) + ((!g8) & (!g10) & (g112) & (!g1174) & (!sk[36]) & (g1425)) + ((!g8) & (!g10) & (g112) & (g1174) & (!sk[36]) & (g1425)) + ((!g8) & (g10) & (!g112) & (!g1174) & (!sk[36]) & (g1425)) + ((!g8) & (g10) & (!g112) & (!g1174) & (sk[36]) & (!g1425)) + ((!g8) & (g10) & (!g112) & (g1174) & (!sk[36]) & (g1425)) + ((!g8) & (g10) & (g112) & (!g1174) & (!sk[36]) & (g1425)) + ((!g8) & (g10) & (g112) & (g1174) & (!sk[36]) & (g1425)) + ((g8) & (!g10) & (!g112) & (!g1174) & (!sk[36]) & (!g1425)) + ((g8) & (!g10) & (!g112) & (!g1174) & (!sk[36]) & (g1425)) + ((g8) & (!g10) & (!g112) & (!g1174) & (sk[36]) & (!g1425)) + ((g8) & (!g10) & (!g112) & (g1174) & (!sk[36]) & (!g1425)) + ((g8) & (!g10) & (!g112) & (g1174) & (!sk[36]) & (g1425)) + ((g8) & (!g10) & (g112) & (!g1174) & (!sk[36]) & (!g1425)) + ((g8) & (!g10) & (g112) & (!g1174) & (!sk[36]) & (g1425)) + ((g8) & (!g10) & (g112) & (!g1174) & (sk[36]) & (!g1425)) + ((g8) & (!g10) & (g112) & (g1174) & (!sk[36]) & (!g1425)) + ((g8) & (!g10) & (g112) & (g1174) & (!sk[36]) & (g1425)) + ((g8) & (g10) & (!g112) & (!g1174) & (!sk[36]) & (!g1425)) + ((g8) & (g10) & (!g112) & (!g1174) & (!sk[36]) & (g1425)) + ((g8) & (g10) & (!g112) & (!g1174) & (sk[36]) & (!g1425)) + ((g8) & (g10) & (!g112) & (g1174) & (!sk[36]) & (!g1425)) + ((g8) & (g10) & (!g112) & (g1174) & (!sk[36]) & (g1425)) + ((g8) & (g10) & (g112) & (!g1174) & (!sk[36]) & (!g1425)) + ((g8) & (g10) & (g112) & (!g1174) & (!sk[36]) & (g1425)) + ((g8) & (g10) & (g112) & (g1174) & (!sk[36]) & (!g1425)) + ((g8) & (g10) & (g112) & (g1174) & (!sk[36]) & (g1425)));
	assign g1427 = (((!g381) & (!g1275) & (!g1423) & (!sk[37]) & (!g1424) & (g1426)) + ((!g381) & (!g1275) & (!g1423) & (!sk[37]) & (g1424) & (g1426)) + ((!g381) & (!g1275) & (g1423) & (!sk[37]) & (!g1424) & (g1426)) + ((!g381) & (!g1275) & (g1423) & (!sk[37]) & (g1424) & (g1426)) + ((!g381) & (g1275) & (!g1423) & (!sk[37]) & (!g1424) & (g1426)) + ((!g381) & (g1275) & (!g1423) & (!sk[37]) & (g1424) & (g1426)) + ((!g381) & (g1275) & (g1423) & (!sk[37]) & (!g1424) & (g1426)) + ((!g381) & (g1275) & (g1423) & (!sk[37]) & (g1424) & (g1426)) + ((!g381) & (g1275) & (g1423) & (sk[37]) & (g1424) & (g1426)) + ((g381) & (!g1275) & (!g1423) & (!sk[37]) & (!g1424) & (!g1426)) + ((g381) & (!g1275) & (!g1423) & (!sk[37]) & (!g1424) & (g1426)) + ((g381) & (!g1275) & (!g1423) & (!sk[37]) & (g1424) & (!g1426)) + ((g381) & (!g1275) & (!g1423) & (!sk[37]) & (g1424) & (g1426)) + ((g381) & (!g1275) & (g1423) & (!sk[37]) & (!g1424) & (!g1426)) + ((g381) & (!g1275) & (g1423) & (!sk[37]) & (!g1424) & (g1426)) + ((g381) & (!g1275) & (g1423) & (!sk[37]) & (g1424) & (!g1426)) + ((g381) & (!g1275) & (g1423) & (!sk[37]) & (g1424) & (g1426)) + ((g381) & (g1275) & (!g1423) & (!sk[37]) & (!g1424) & (!g1426)) + ((g381) & (g1275) & (!g1423) & (!sk[37]) & (!g1424) & (g1426)) + ((g381) & (g1275) & (!g1423) & (!sk[37]) & (g1424) & (!g1426)) + ((g381) & (g1275) & (!g1423) & (!sk[37]) & (g1424) & (g1426)) + ((g381) & (g1275) & (g1423) & (!sk[37]) & (!g1424) & (!g1426)) + ((g381) & (g1275) & (g1423) & (!sk[37]) & (!g1424) & (g1426)) + ((g381) & (g1275) & (g1423) & (!sk[37]) & (g1424) & (!g1426)) + ((g381) & (g1275) & (g1423) & (!sk[37]) & (g1424) & (g1426)));
	assign g1428 = (((g1151) & (!g1358) & (!sk[38]) & (!g1398)) + ((g1151) & (!g1358) & (!sk[38]) & (g1398)) + ((g1151) & (g1358) & (!sk[38]) & (!g1398)) + ((g1151) & (g1358) & (!sk[38]) & (g1398)) + ((g1151) & (g1358) & (sk[38]) & (g1398)));
	assign g1429 = (((g1219) & (g1415) & (!g1421) & (g1422) & (g1427) & (g1428)));
	assign g1430 = (((!sk[40]) & (!g560) & (!g561) & (!g549) & (!g540) & (g895)) + ((!sk[40]) & (!g560) & (!g561) & (!g549) & (g540) & (g895)) + ((!sk[40]) & (!g560) & (!g561) & (g549) & (!g540) & (g895)) + ((!sk[40]) & (!g560) & (!g561) & (g549) & (g540) & (g895)) + ((!sk[40]) & (!g560) & (g561) & (!g549) & (!g540) & (g895)) + ((!sk[40]) & (!g560) & (g561) & (!g549) & (g540) & (g895)) + ((!sk[40]) & (!g560) & (g561) & (g549) & (!g540) & (g895)) + ((!sk[40]) & (!g560) & (g561) & (g549) & (g540) & (g895)) + ((!sk[40]) & (g560) & (!g561) & (!g549) & (!g540) & (!g895)) + ((!sk[40]) & (g560) & (!g561) & (!g549) & (!g540) & (g895)) + ((!sk[40]) & (g560) & (!g561) & (!g549) & (g540) & (!g895)) + ((!sk[40]) & (g560) & (!g561) & (!g549) & (g540) & (g895)) + ((!sk[40]) & (g560) & (!g561) & (g549) & (!g540) & (!g895)) + ((!sk[40]) & (g560) & (!g561) & (g549) & (!g540) & (g895)) + ((!sk[40]) & (g560) & (!g561) & (g549) & (g540) & (!g895)) + ((!sk[40]) & (g560) & (!g561) & (g549) & (g540) & (g895)) + ((!sk[40]) & (g560) & (g561) & (!g549) & (!g540) & (!g895)) + ((!sk[40]) & (g560) & (g561) & (!g549) & (!g540) & (g895)) + ((!sk[40]) & (g560) & (g561) & (!g549) & (g540) & (!g895)) + ((!sk[40]) & (g560) & (g561) & (!g549) & (g540) & (g895)) + ((!sk[40]) & (g560) & (g561) & (g549) & (!g540) & (!g895)) + ((!sk[40]) & (g560) & (g561) & (g549) & (!g540) & (g895)) + ((!sk[40]) & (g560) & (g561) & (g549) & (g540) & (!g895)) + ((!sk[40]) & (g560) & (g561) & (g549) & (g540) & (g895)) + ((sk[40]) & (!g560) & (!g561) & (g549) & (!g540) & (!g895)));
	assign g1431 = (((!g134) & (!sk[41]) & (!g824) & (g1300) & (g1430)) + ((!g134) & (!sk[41]) & (g824) & (!g1300) & (!g1430)) + ((!g134) & (!sk[41]) & (g824) & (!g1300) & (g1430)) + ((!g134) & (!sk[41]) & (g824) & (g1300) & (!g1430)) + ((!g134) & (!sk[41]) & (g824) & (g1300) & (g1430)) + ((!g134) & (sk[41]) & (!g824) & (g1300) & (!g1430)) + ((!g134) & (sk[41]) & (!g824) & (g1300) & (g1430)) + ((!g134) & (sk[41]) & (g824) & (g1300) & (!g1430)) + ((!g134) & (sk[41]) & (g824) & (g1300) & (g1430)) + ((g134) & (!sk[41]) & (!g824) & (g1300) & (!g1430)) + ((g134) & (!sk[41]) & (!g824) & (g1300) & (g1430)) + ((g134) & (!sk[41]) & (g824) & (!g1300) & (!g1430)) + ((g134) & (!sk[41]) & (g824) & (!g1300) & (g1430)) + ((g134) & (!sk[41]) & (g824) & (g1300) & (!g1430)) + ((g134) & (!sk[41]) & (g824) & (g1300) & (g1430)) + ((g134) & (sk[41]) & (g824) & (g1300) & (g1430)));
	assign g1432 = (((!g8) & (!g10) & (!g23) & (g136) & (!g132) & (!g462)) + ((!g8) & (!g10) & (!g23) & (g136) & (!g132) & (g462)) + ((!g8) & (!g10) & (!g23) & (g136) & (g132) & (!g462)) + ((!g8) & (!g10) & (!g23) & (g136) & (g132) & (g462)) + ((!g8) & (!g10) & (g23) & (g136) & (!g132) & (!g462)) + ((!g8) & (!g10) & (g23) & (g136) & (!g132) & (g462)) + ((!g8) & (!g10) & (g23) & (g136) & (g132) & (!g462)) + ((!g8) & (!g10) & (g23) & (g136) & (g132) & (g462)) + ((!g8) & (g10) & (!g23) & (g136) & (!g132) & (!g462)) + ((!g8) & (g10) & (!g23) & (g136) & (!g132) & (g462)) + ((!g8) & (g10) & (!g23) & (g136) & (g132) & (!g462)) + ((!g8) & (g10) & (!g23) & (g136) & (g132) & (g462)) + ((!g8) & (g10) & (g23) & (g136) & (!g132) & (!g462)) + ((!g8) & (g10) & (g23) & (g136) & (!g132) & (g462)) + ((!g8) & (g10) & (g23) & (g136) & (g132) & (!g462)) + ((!g8) & (g10) & (g23) & (g136) & (g132) & (g462)) + ((g8) & (!g10) & (!g23) & (g136) & (!g132) & (!g462)) + ((g8) & (!g10) & (!g23) & (g136) & (!g132) & (g462)) + ((g8) & (!g10) & (!g23) & (g136) & (g132) & (!g462)) + ((g8) & (!g10) & (g23) & (g136) & (!g132) & (!g462)) + ((g8) & (!g10) & (g23) & (g136) & (!g132) & (g462)) + ((g8) & (!g10) & (g23) & (g136) & (g132) & (!g462)) + ((g8) & (!g10) & (g23) & (g136) & (g132) & (g462)) + ((g8) & (g10) & (!g23) & (g136) & (!g132) & (!g462)) + ((g8) & (g10) & (!g23) & (g136) & (!g132) & (g462)) + ((g8) & (g10) & (!g23) & (g136) & (g132) & (!g462)) + ((g8) & (g10) & (!g23) & (g136) & (g132) & (g462)) + ((g8) & (g10) & (g23) & (g136) & (!g132) & (!g462)) + ((g8) & (g10) & (g23) & (g136) & (!g132) & (g462)) + ((g8) & (g10) & (g23) & (g136) & (g132) & (!g462)) + ((g8) & (g10) & (g23) & (g136) & (g132) & (g462)));
	assign g1433 = (((!i_14_) & (!i_12_) & (!i_13_) & (g136) & (!g131) & (g158)) + ((!i_14_) & (!i_12_) & (!i_13_) & (g136) & (g131) & (g158)) + ((!i_14_) & (i_12_) & (!i_13_) & (g136) & (!g131) & (g158)) + ((!i_14_) & (i_12_) & (!i_13_) & (g136) & (g131) & (g158)) + ((!i_14_) & (i_12_) & (i_13_) & (g136) & (!g131) & (g158)) + ((!i_14_) & (i_12_) & (i_13_) & (g136) & (g131) & (g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (g136) & (g131) & (!g158)) + ((i_14_) & (!i_12_) & (!i_13_) & (g136) & (g131) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (g136) & (!g131) & (g158)) + ((i_14_) & (i_12_) & (!i_13_) & (g136) & (g131) & (g158)) + ((i_14_) & (i_12_) & (i_13_) & (g136) & (g131) & (!g158)) + ((i_14_) & (i_12_) & (i_13_) & (g136) & (g131) & (g158)));
	assign g1434 = (((!g135) & (!g1112) & (g1263) & (!g1419) & (!g1432) & (!g1433)) + ((!g135) & (!g1112) & (g1263) & (g1419) & (!g1432) & (!g1433)) + ((!g135) & (g1112) & (g1263) & (!g1419) & (!g1432) & (!g1433)) + ((!g135) & (g1112) & (g1263) & (g1419) & (!g1432) & (!g1433)) + ((g135) & (g1112) & (g1263) & (!g1419) & (!g1432) & (!g1433)));
	assign g1435 = (((!g1202) & (!g1229) & (!g1352) & (!sk[45]) & (!g1434) & (g1640)) + ((!g1202) & (!g1229) & (!g1352) & (!sk[45]) & (g1434) & (g1640)) + ((!g1202) & (!g1229) & (g1352) & (!sk[45]) & (!g1434) & (g1640)) + ((!g1202) & (!g1229) & (g1352) & (!sk[45]) & (g1434) & (g1640)) + ((!g1202) & (g1229) & (!g1352) & (!sk[45]) & (!g1434) & (g1640)) + ((!g1202) & (g1229) & (!g1352) & (!sk[45]) & (g1434) & (g1640)) + ((!g1202) & (g1229) & (g1352) & (!sk[45]) & (!g1434) & (g1640)) + ((!g1202) & (g1229) & (g1352) & (!sk[45]) & (g1434) & (g1640)) + ((g1202) & (!g1229) & (!g1352) & (!sk[45]) & (!g1434) & (!g1640)) + ((g1202) & (!g1229) & (!g1352) & (!sk[45]) & (!g1434) & (g1640)) + ((g1202) & (!g1229) & (!g1352) & (!sk[45]) & (g1434) & (!g1640)) + ((g1202) & (!g1229) & (!g1352) & (!sk[45]) & (g1434) & (g1640)) + ((g1202) & (!g1229) & (g1352) & (!sk[45]) & (!g1434) & (!g1640)) + ((g1202) & (!g1229) & (g1352) & (!sk[45]) & (!g1434) & (g1640)) + ((g1202) & (!g1229) & (g1352) & (!sk[45]) & (g1434) & (!g1640)) + ((g1202) & (!g1229) & (g1352) & (!sk[45]) & (g1434) & (g1640)) + ((g1202) & (g1229) & (!g1352) & (!sk[45]) & (!g1434) & (!g1640)) + ((g1202) & (g1229) & (!g1352) & (!sk[45]) & (!g1434) & (g1640)) + ((g1202) & (g1229) & (!g1352) & (!sk[45]) & (g1434) & (!g1640)) + ((g1202) & (g1229) & (!g1352) & (!sk[45]) & (g1434) & (g1640)) + ((g1202) & (g1229) & (g1352) & (!sk[45]) & (!g1434) & (!g1640)) + ((g1202) & (g1229) & (g1352) & (!sk[45]) & (!g1434) & (g1640)) + ((g1202) & (g1229) & (g1352) & (!sk[45]) & (g1434) & (!g1640)) + ((g1202) & (g1229) & (g1352) & (!sk[45]) & (g1434) & (g1640)) + ((g1202) & (g1229) & (g1352) & (sk[45]) & (g1434) & (g1640)));
	assign o_20_ = (((g73) & (!g1329) & (!g1568) & (!g1429) & (!g1431) & (!g1435)) + ((g73) & (!g1329) & (!g1568) & (!g1429) & (!g1431) & (g1435)) + ((g73) & (!g1329) & (!g1568) & (!g1429) & (g1431) & (!g1435)) + ((g73) & (!g1329) & (!g1568) & (!g1429) & (g1431) & (g1435)) + ((g73) & (!g1329) & (!g1568) & (g1429) & (!g1431) & (!g1435)) + ((g73) & (!g1329) & (!g1568) & (g1429) & (!g1431) & (g1435)) + ((g73) & (!g1329) & (!g1568) & (g1429) & (g1431) & (!g1435)) + ((g73) & (!g1329) & (!g1568) & (g1429) & (g1431) & (g1435)) + ((g73) & (!g1329) & (g1568) & (!g1429) & (!g1431) & (!g1435)) + ((g73) & (!g1329) & (g1568) & (!g1429) & (!g1431) & (g1435)) + ((g73) & (!g1329) & (g1568) & (!g1429) & (g1431) & (!g1435)) + ((g73) & (!g1329) & (g1568) & (!g1429) & (g1431) & (g1435)) + ((g73) & (!g1329) & (g1568) & (g1429) & (!g1431) & (!g1435)) + ((g73) & (!g1329) & (g1568) & (g1429) & (!g1431) & (g1435)) + ((g73) & (!g1329) & (g1568) & (g1429) & (g1431) & (!g1435)) + ((g73) & (!g1329) & (g1568) & (g1429) & (g1431) & (g1435)) + ((g73) & (g1329) & (!g1568) & (!g1429) & (!g1431) & (!g1435)) + ((g73) & (g1329) & (!g1568) & (!g1429) & (!g1431) & (g1435)) + ((g73) & (g1329) & (!g1568) & (!g1429) & (g1431) & (!g1435)) + ((g73) & (g1329) & (!g1568) & (!g1429) & (g1431) & (g1435)) + ((g73) & (g1329) & (!g1568) & (g1429) & (!g1431) & (!g1435)) + ((g73) & (g1329) & (!g1568) & (g1429) & (!g1431) & (g1435)) + ((g73) & (g1329) & (!g1568) & (g1429) & (g1431) & (!g1435)) + ((g73) & (g1329) & (!g1568) & (g1429) & (g1431) & (g1435)) + ((g73) & (g1329) & (g1568) & (!g1429) & (!g1431) & (!g1435)) + ((g73) & (g1329) & (g1568) & (!g1429) & (!g1431) & (g1435)) + ((g73) & (g1329) & (g1568) & (!g1429) & (g1431) & (!g1435)) + ((g73) & (g1329) & (g1568) & (!g1429) & (g1431) & (g1435)) + ((g73) & (g1329) & (g1568) & (g1429) & (!g1431) & (!g1435)) + ((g73) & (g1329) & (g1568) & (g1429) & (!g1431) & (g1435)) + ((g73) & (g1329) & (g1568) & (g1429) & (g1431) & (!g1435)));
	assign g1437 = (((!g73) & (sk[47]) & (!g1429)) + ((!g73) & (sk[47]) & (g1429)) + ((g73) & (!sk[47]) & (!g1429)) + ((g73) & (!sk[47]) & (g1429)) + ((g73) & (sk[47]) & (g1429)));
	assign g1438 = (((!i_11_) & (!i_9_) & (!sk[48]) & (i_10_) & (i_8_)) + ((!i_11_) & (!i_9_) & (sk[48]) & (!i_10_) & (i_8_)) + ((!i_11_) & (!i_9_) & (sk[48]) & (i_10_) & (i_8_)) + ((!i_11_) & (i_9_) & (!sk[48]) & (!i_10_) & (!i_8_)) + ((!i_11_) & (i_9_) & (!sk[48]) & (!i_10_) & (i_8_)) + ((!i_11_) & (i_9_) & (!sk[48]) & (i_10_) & (!i_8_)) + ((!i_11_) & (i_9_) & (!sk[48]) & (i_10_) & (i_8_)) + ((!i_11_) & (i_9_) & (sk[48]) & (!i_10_) & (!i_8_)) + ((!i_11_) & (i_9_) & (sk[48]) & (i_10_) & (!i_8_)) + ((i_11_) & (!i_9_) & (!sk[48]) & (i_10_) & (!i_8_)) + ((i_11_) & (!i_9_) & (!sk[48]) & (i_10_) & (i_8_)) + ((i_11_) & (!i_9_) & (sk[48]) & (!i_10_) & (i_8_)) + ((i_11_) & (!i_9_) & (sk[48]) & (i_10_) & (i_8_)) + ((i_11_) & (i_9_) & (!sk[48]) & (!i_10_) & (!i_8_)) + ((i_11_) & (i_9_) & (!sk[48]) & (!i_10_) & (i_8_)) + ((i_11_) & (i_9_) & (!sk[48]) & (i_10_) & (!i_8_)) + ((i_11_) & (i_9_) & (!sk[48]) & (i_10_) & (i_8_)) + ((i_11_) & (i_9_) & (sk[48]) & (i_10_) & (!i_8_)));
	assign g1439 = (((!i_15_) & (!sk[49]) & (!g4) & (!g87) & (!g182) & (g1438)) + ((!i_15_) & (!sk[49]) & (!g4) & (!g87) & (g182) & (g1438)) + ((!i_15_) & (!sk[49]) & (!g4) & (g87) & (!g182) & (g1438)) + ((!i_15_) & (!sk[49]) & (!g4) & (g87) & (g182) & (g1438)) + ((!i_15_) & (!sk[49]) & (g4) & (!g87) & (!g182) & (g1438)) + ((!i_15_) & (!sk[49]) & (g4) & (!g87) & (g182) & (g1438)) + ((!i_15_) & (!sk[49]) & (g4) & (g87) & (!g182) & (g1438)) + ((!i_15_) & (!sk[49]) & (g4) & (g87) & (g182) & (g1438)) + ((i_15_) & (!sk[49]) & (!g4) & (!g87) & (!g182) & (!g1438)) + ((i_15_) & (!sk[49]) & (!g4) & (!g87) & (!g182) & (g1438)) + ((i_15_) & (!sk[49]) & (!g4) & (!g87) & (g182) & (!g1438)) + ((i_15_) & (!sk[49]) & (!g4) & (!g87) & (g182) & (g1438)) + ((i_15_) & (!sk[49]) & (!g4) & (g87) & (!g182) & (!g1438)) + ((i_15_) & (!sk[49]) & (!g4) & (g87) & (!g182) & (g1438)) + ((i_15_) & (!sk[49]) & (!g4) & (g87) & (g182) & (!g1438)) + ((i_15_) & (!sk[49]) & (!g4) & (g87) & (g182) & (g1438)) + ((i_15_) & (!sk[49]) & (g4) & (!g87) & (!g182) & (!g1438)) + ((i_15_) & (!sk[49]) & (g4) & (!g87) & (!g182) & (g1438)) + ((i_15_) & (!sk[49]) & (g4) & (!g87) & (g182) & (!g1438)) + ((i_15_) & (!sk[49]) & (g4) & (!g87) & (g182) & (g1438)) + ((i_15_) & (!sk[49]) & (g4) & (g87) & (!g182) & (!g1438)) + ((i_15_) & (!sk[49]) & (g4) & (g87) & (!g182) & (g1438)) + ((i_15_) & (!sk[49]) & (g4) & (g87) & (g182) & (!g1438)) + ((i_15_) & (!sk[49]) & (g4) & (g87) & (g182) & (g1438)) + ((i_15_) & (sk[49]) & (g4) & (g87) & (g182) & (g1438)));
	assign o_22_ = (((!g227) & (!g349) & (!g1007) & (sk[50]) & (g1439)) + ((!g227) & (!g349) & (g1007) & (!sk[50]) & (g1439)) + ((!g227) & (!g349) & (g1007) & (sk[50]) & (!g1439)) + ((!g227) & (!g349) & (g1007) & (sk[50]) & (g1439)) + ((!g227) & (g349) & (!g1007) & (!sk[50]) & (!g1439)) + ((!g227) & (g349) & (!g1007) & (!sk[50]) & (g1439)) + ((!g227) & (g349) & (!g1007) & (sk[50]) & (g1439)) + ((!g227) & (g349) & (g1007) & (!sk[50]) & (!g1439)) + ((!g227) & (g349) & (g1007) & (!sk[50]) & (g1439)) + ((!g227) & (g349) & (g1007) & (sk[50]) & (!g1439)) + ((!g227) & (g349) & (g1007) & (sk[50]) & (g1439)) + ((g227) & (!g349) & (!g1007) & (sk[50]) & (g1439)) + ((g227) & (!g349) & (g1007) & (!sk[50]) & (!g1439)) + ((g227) & (!g349) & (g1007) & (!sk[50]) & (g1439)) + ((g227) & (!g349) & (g1007) & (sk[50]) & (!g1439)) + ((g227) & (!g349) & (g1007) & (sk[50]) & (g1439)) + ((g227) & (g349) & (!g1007) & (!sk[50]) & (!g1439)) + ((g227) & (g349) & (!g1007) & (!sk[50]) & (g1439)) + ((g227) & (g349) & (!g1007) & (sk[50]) & (!g1439)) + ((g227) & (g349) & (!g1007) & (sk[50]) & (g1439)) + ((g227) & (g349) & (g1007) & (!sk[50]) & (!g1439)) + ((g227) & (g349) & (g1007) & (!sk[50]) & (g1439)) + ((g227) & (g349) & (g1007) & (sk[50]) & (!g1439)) + ((g227) & (g349) & (g1007) & (sk[50]) & (g1439)));
	assign g1441 = (((!i_5_) & (!i_3_) & (!sk[51]) & (i_4_) & (g1)) + ((!i_5_) & (i_3_) & (!sk[51]) & (!i_4_) & (!g1)) + ((!i_5_) & (i_3_) & (!sk[51]) & (!i_4_) & (g1)) + ((!i_5_) & (i_3_) & (!sk[51]) & (i_4_) & (!g1)) + ((!i_5_) & (i_3_) & (!sk[51]) & (i_4_) & (g1)) + ((i_5_) & (!i_3_) & (!sk[51]) & (i_4_) & (!g1)) + ((i_5_) & (!i_3_) & (!sk[51]) & (i_4_) & (g1)) + ((i_5_) & (i_3_) & (!sk[51]) & (!i_4_) & (!g1)) + ((i_5_) & (i_3_) & (!sk[51]) & (!i_4_) & (g1)) + ((i_5_) & (i_3_) & (!sk[51]) & (i_4_) & (!g1)) + ((i_5_) & (i_3_) & (!sk[51]) & (i_4_) & (g1)) + ((i_5_) & (i_3_) & (sk[51]) & (i_4_) & (g1)));
	assign g1442 = (((!sk[52]) & (g30) & (!g1441)) + ((!sk[52]) & (g30) & (g1441)) + ((sk[52]) & (g30) & (g1441)));
	assign g1443 = (((!g1155) & (!g1230) & (!g1231) & (g1234) & (g1307) & (g1309)));
	assign g1444 = (((!g132) & (!sk[54]) & (!g159) & (!g566) & (!g531) & (g522)) + ((!g132) & (!sk[54]) & (!g159) & (!g566) & (g531) & (g522)) + ((!g132) & (!sk[54]) & (!g159) & (g566) & (!g531) & (g522)) + ((!g132) & (!sk[54]) & (!g159) & (g566) & (g531) & (g522)) + ((!g132) & (!sk[54]) & (g159) & (!g566) & (!g531) & (g522)) + ((!g132) & (!sk[54]) & (g159) & (!g566) & (g531) & (g522)) + ((!g132) & (!sk[54]) & (g159) & (g566) & (!g531) & (g522)) + ((!g132) & (!sk[54]) & (g159) & (g566) & (g531) & (g522)) + ((g132) & (!sk[54]) & (!g159) & (!g566) & (!g531) & (!g522)) + ((g132) & (!sk[54]) & (!g159) & (!g566) & (!g531) & (g522)) + ((g132) & (!sk[54]) & (!g159) & (!g566) & (g531) & (!g522)) + ((g132) & (!sk[54]) & (!g159) & (!g566) & (g531) & (g522)) + ((g132) & (!sk[54]) & (!g159) & (g566) & (!g531) & (!g522)) + ((g132) & (!sk[54]) & (!g159) & (g566) & (!g531) & (g522)) + ((g132) & (!sk[54]) & (!g159) & (g566) & (g531) & (!g522)) + ((g132) & (!sk[54]) & (!g159) & (g566) & (g531) & (g522)) + ((g132) & (!sk[54]) & (g159) & (!g566) & (!g531) & (!g522)) + ((g132) & (!sk[54]) & (g159) & (!g566) & (!g531) & (g522)) + ((g132) & (!sk[54]) & (g159) & (!g566) & (g531) & (!g522)) + ((g132) & (!sk[54]) & (g159) & (!g566) & (g531) & (g522)) + ((g132) & (!sk[54]) & (g159) & (g566) & (!g531) & (!g522)) + ((g132) & (!sk[54]) & (g159) & (g566) & (!g531) & (g522)) + ((g132) & (!sk[54]) & (g159) & (g566) & (g531) & (!g522)) + ((g132) & (!sk[54]) & (g159) & (g566) & (g531) & (g522)) + ((g132) & (sk[54]) & (!g159) & (!g566) & (!g531) & (!g522)));
	assign g1445 = (((!i_8_) & (!g66) & (g108) & (!g207) & (!g1085) & (!g1444)) + ((!i_8_) & (!g66) & (g108) & (!g207) & (!g1085) & (g1444)) + ((!i_8_) & (!g66) & (g108) & (!g207) & (g1085) & (!g1444)) + ((!i_8_) & (!g66) & (g108) & (g207) & (!g1085) & (!g1444)) + ((!i_8_) & (!g66) & (g108) & (g207) & (!g1085) & (g1444)) + ((!i_8_) & (!g66) & (g108) & (g207) & (g1085) & (!g1444)) + ((!i_8_) & (g66) & (g108) & (!g207) & (!g1085) & (!g1444)) + ((!i_8_) & (g66) & (g108) & (!g207) & (!g1085) & (g1444)) + ((!i_8_) & (g66) & (g108) & (!g207) & (g1085) & (!g1444)) + ((!i_8_) & (g66) & (g108) & (g207) & (!g1085) & (!g1444)) + ((!i_8_) & (g66) & (g108) & (g207) & (!g1085) & (g1444)) + ((!i_8_) & (g66) & (g108) & (g207) & (g1085) & (!g1444)) + ((i_8_) & (!g66) & (g108) & (g207) & (!g1085) & (!g1444)) + ((i_8_) & (!g66) & (g108) & (g207) & (!g1085) & (g1444)) + ((i_8_) & (!g66) & (g108) & (g207) & (g1085) & (!g1444)) + ((i_8_) & (g66) & (g108) & (!g207) & (!g1085) & (!g1444)) + ((i_8_) & (g66) & (g108) & (!g207) & (!g1085) & (g1444)) + ((i_8_) & (g66) & (g108) & (!g207) & (g1085) & (!g1444)) + ((i_8_) & (g66) & (g108) & (!g207) & (g1085) & (g1444)) + ((i_8_) & (g66) & (g108) & (g207) & (!g1085) & (!g1444)) + ((i_8_) & (g66) & (g108) & (g207) & (!g1085) & (g1444)) + ((i_8_) & (g66) & (g108) & (g207) & (g1085) & (!g1444)) + ((i_8_) & (g66) & (g108) & (g207) & (g1085) & (g1444)));
	assign g1446 = (((!i_14_) & (!i_12_) & (!sk[56]) & (!i_13_) & (!g131) & (g158)) + ((!i_14_) & (!i_12_) & (!sk[56]) & (!i_13_) & (g131) & (g158)) + ((!i_14_) & (!i_12_) & (!sk[56]) & (i_13_) & (!g131) & (g158)) + ((!i_14_) & (!i_12_) & (!sk[56]) & (i_13_) & (g131) & (g158)) + ((!i_14_) & (!i_12_) & (sk[56]) & (!i_13_) & (g131) & (!g158)) + ((!i_14_) & (!i_12_) & (sk[56]) & (!i_13_) & (g131) & (g158)) + ((!i_14_) & (!i_12_) & (sk[56]) & (i_13_) & (!g131) & (g158)) + ((!i_14_) & (!i_12_) & (sk[56]) & (i_13_) & (g131) & (g158)) + ((!i_14_) & (i_12_) & (!sk[56]) & (!i_13_) & (!g131) & (g158)) + ((!i_14_) & (i_12_) & (!sk[56]) & (!i_13_) & (g131) & (g158)) + ((!i_14_) & (i_12_) & (!sk[56]) & (i_13_) & (!g131) & (g158)) + ((!i_14_) & (i_12_) & (!sk[56]) & (i_13_) & (g131) & (g158)) + ((!i_14_) & (i_12_) & (sk[56]) & (i_13_) & (g131) & (!g158)) + ((!i_14_) & (i_12_) & (sk[56]) & (i_13_) & (g131) & (g158)) + ((i_14_) & (!i_12_) & (!sk[56]) & (!i_13_) & (!g131) & (!g158)) + ((i_14_) & (!i_12_) & (!sk[56]) & (!i_13_) & (!g131) & (g158)) + ((i_14_) & (!i_12_) & (!sk[56]) & (!i_13_) & (g131) & (!g158)) + ((i_14_) & (!i_12_) & (!sk[56]) & (!i_13_) & (g131) & (g158)) + ((i_14_) & (!i_12_) & (!sk[56]) & (i_13_) & (!g131) & (!g158)) + ((i_14_) & (!i_12_) & (!sk[56]) & (i_13_) & (!g131) & (g158)) + ((i_14_) & (!i_12_) & (!sk[56]) & (i_13_) & (g131) & (!g158)) + ((i_14_) & (!i_12_) & (!sk[56]) & (i_13_) & (g131) & (g158)) + ((i_14_) & (i_12_) & (!sk[56]) & (!i_13_) & (!g131) & (!g158)) + ((i_14_) & (i_12_) & (!sk[56]) & (!i_13_) & (!g131) & (g158)) + ((i_14_) & (i_12_) & (!sk[56]) & (!i_13_) & (g131) & (!g158)) + ((i_14_) & (i_12_) & (!sk[56]) & (!i_13_) & (g131) & (g158)) + ((i_14_) & (i_12_) & (!sk[56]) & (i_13_) & (!g131) & (!g158)) + ((i_14_) & (i_12_) & (!sk[56]) & (i_13_) & (!g131) & (g158)) + ((i_14_) & (i_12_) & (!sk[56]) & (i_13_) & (g131) & (!g158)) + ((i_14_) & (i_12_) & (!sk[56]) & (i_13_) & (g131) & (g158)) + ((i_14_) & (i_12_) & (sk[56]) & (!i_13_) & (g131) & (!g158)) + ((i_14_) & (i_12_) & (sk[56]) & (!i_13_) & (g131) & (g158)) + ((i_14_) & (i_12_) & (sk[56]) & (i_13_) & (!g131) & (g158)) + ((i_14_) & (i_12_) & (sk[56]) & (i_13_) & (g131) & (g158)));
	assign g1447 = (((!g46) & (!g101) & (!sk[57]) & (!g108) & (!g209) & (g1446)) + ((!g46) & (!g101) & (!sk[57]) & (!g108) & (g209) & (g1446)) + ((!g46) & (!g101) & (!sk[57]) & (g108) & (!g209) & (g1446)) + ((!g46) & (!g101) & (!sk[57]) & (g108) & (g209) & (g1446)) + ((!g46) & (!g101) & (sk[57]) & (!g108) & (!g209) & (!g1446)) + ((!g46) & (!g101) & (sk[57]) & (!g108) & (!g209) & (g1446)) + ((!g46) & (!g101) & (sk[57]) & (!g108) & (g209) & (!g1446)) + ((!g46) & (!g101) & (sk[57]) & (!g108) & (g209) & (g1446)) + ((!g46) & (!g101) & (sk[57]) & (g108) & (!g209) & (!g1446)) + ((!g46) & (!g101) & (sk[57]) & (g108) & (g209) & (!g1446)) + ((!g46) & (g101) & (!sk[57]) & (!g108) & (!g209) & (g1446)) + ((!g46) & (g101) & (!sk[57]) & (!g108) & (g209) & (g1446)) + ((!g46) & (g101) & (!sk[57]) & (g108) & (!g209) & (g1446)) + ((!g46) & (g101) & (!sk[57]) & (g108) & (g209) & (g1446)) + ((!g46) & (g101) & (sk[57]) & (!g108) & (!g209) & (!g1446)) + ((!g46) & (g101) & (sk[57]) & (!g108) & (!g209) & (g1446)) + ((!g46) & (g101) & (sk[57]) & (g108) & (!g209) & (!g1446)) + ((g46) & (!g101) & (!sk[57]) & (!g108) & (!g209) & (!g1446)) + ((g46) & (!g101) & (!sk[57]) & (!g108) & (!g209) & (g1446)) + ((g46) & (!g101) & (!sk[57]) & (!g108) & (g209) & (!g1446)) + ((g46) & (!g101) & (!sk[57]) & (!g108) & (g209) & (g1446)) + ((g46) & (!g101) & (!sk[57]) & (g108) & (!g209) & (!g1446)) + ((g46) & (!g101) & (!sk[57]) & (g108) & (!g209) & (g1446)) + ((g46) & (!g101) & (!sk[57]) & (g108) & (g209) & (!g1446)) + ((g46) & (!g101) & (!sk[57]) & (g108) & (g209) & (g1446)) + ((g46) & (!g101) & (sk[57]) & (!g108) & (!g209) & (!g1446)) + ((g46) & (!g101) & (sk[57]) & (!g108) & (!g209) & (g1446)) + ((g46) & (!g101) & (sk[57]) & (!g108) & (g209) & (!g1446)) + ((g46) & (!g101) & (sk[57]) & (!g108) & (g209) & (g1446)) + ((g46) & (!g101) & (sk[57]) & (g108) & (!g209) & (!g1446)) + ((g46) & (!g101) & (sk[57]) & (g108) & (g209) & (!g1446)) + ((g46) & (g101) & (!sk[57]) & (!g108) & (!g209) & (!g1446)) + ((g46) & (g101) & (!sk[57]) & (!g108) & (!g209) & (g1446)) + ((g46) & (g101) & (!sk[57]) & (!g108) & (g209) & (!g1446)) + ((g46) & (g101) & (!sk[57]) & (!g108) & (g209) & (g1446)) + ((g46) & (g101) & (!sk[57]) & (g108) & (!g209) & (!g1446)) + ((g46) & (g101) & (!sk[57]) & (g108) & (!g209) & (g1446)) + ((g46) & (g101) & (!sk[57]) & (g108) & (g209) & (!g1446)) + ((g46) & (g101) & (!sk[57]) & (g108) & (g209) & (g1446)));
	assign g1448 = (((!g109) & (!g529) & (!g801) & (!g819) & (!sk[58]) & (g1260)) + ((!g109) & (!g529) & (!g801) & (!g819) & (sk[58]) & (!g1260)) + ((!g109) & (!g529) & (!g801) & (!g819) & (sk[58]) & (g1260)) + ((!g109) & (!g529) & (!g801) & (g819) & (!sk[58]) & (g1260)) + ((!g109) & (!g529) & (g801) & (!g819) & (!sk[58]) & (g1260)) + ((!g109) & (!g529) & (g801) & (!g819) & (sk[58]) & (!g1260)) + ((!g109) & (!g529) & (g801) & (!g819) & (sk[58]) & (g1260)) + ((!g109) & (!g529) & (g801) & (g819) & (!sk[58]) & (g1260)) + ((!g109) & (g529) & (!g801) & (!g819) & (!sk[58]) & (g1260)) + ((!g109) & (g529) & (!g801) & (!g819) & (sk[58]) & (!g1260)) + ((!g109) & (g529) & (!g801) & (!g819) & (sk[58]) & (g1260)) + ((!g109) & (g529) & (!g801) & (g819) & (!sk[58]) & (g1260)) + ((!g109) & (g529) & (g801) & (!g819) & (!sk[58]) & (g1260)) + ((!g109) & (g529) & (g801) & (!g819) & (sk[58]) & (!g1260)) + ((!g109) & (g529) & (g801) & (!g819) & (sk[58]) & (g1260)) + ((!g109) & (g529) & (g801) & (g819) & (!sk[58]) & (g1260)) + ((g109) & (!g529) & (!g801) & (!g819) & (!sk[58]) & (!g1260)) + ((g109) & (!g529) & (!g801) & (!g819) & (!sk[58]) & (g1260)) + ((g109) & (!g529) & (!g801) & (g819) & (!sk[58]) & (!g1260)) + ((g109) & (!g529) & (!g801) & (g819) & (!sk[58]) & (g1260)) + ((g109) & (!g529) & (g801) & (!g819) & (!sk[58]) & (!g1260)) + ((g109) & (!g529) & (g801) & (!g819) & (!sk[58]) & (g1260)) + ((g109) & (!g529) & (g801) & (g819) & (!sk[58]) & (!g1260)) + ((g109) & (!g529) & (g801) & (g819) & (!sk[58]) & (g1260)) + ((g109) & (g529) & (!g801) & (!g819) & (!sk[58]) & (!g1260)) + ((g109) & (g529) & (!g801) & (!g819) & (!sk[58]) & (g1260)) + ((g109) & (g529) & (!g801) & (g819) & (!sk[58]) & (!g1260)) + ((g109) & (g529) & (!g801) & (g819) & (!sk[58]) & (g1260)) + ((g109) & (g529) & (g801) & (!g819) & (!sk[58]) & (!g1260)) + ((g109) & (g529) & (g801) & (!g819) & (!sk[58]) & (g1260)) + ((g109) & (g529) & (g801) & (!g819) & (sk[58]) & (g1260)) + ((g109) & (g529) & (g801) & (g819) & (!sk[58]) & (!g1260)) + ((g109) & (g529) & (g801) & (g819) & (!sk[58]) & (g1260)));
	assign g1449 = (((!sk[59]) & (!i_8_) & (!g108) & (g316) & (g132)) + ((!sk[59]) & (!i_8_) & (g108) & (!g316) & (!g132)) + ((!sk[59]) & (!i_8_) & (g108) & (!g316) & (g132)) + ((!sk[59]) & (!i_8_) & (g108) & (g316) & (!g132)) + ((!sk[59]) & (!i_8_) & (g108) & (g316) & (g132)) + ((!sk[59]) & (i_8_) & (!g108) & (g316) & (!g132)) + ((!sk[59]) & (i_8_) & (!g108) & (g316) & (g132)) + ((!sk[59]) & (i_8_) & (g108) & (!g316) & (!g132)) + ((!sk[59]) & (i_8_) & (g108) & (!g316) & (g132)) + ((!sk[59]) & (i_8_) & (g108) & (g316) & (!g132)) + ((!sk[59]) & (i_8_) & (g108) & (g316) & (g132)) + ((sk[59]) & (!i_8_) & (g108) & (g316) & (!g132)) + ((sk[59]) & (!i_8_) & (g108) & (g316) & (g132)) + ((sk[59]) & (i_8_) & (g108) & (!g316) & (!g132)) + ((sk[59]) & (i_8_) & (g108) & (g316) & (!g132)));
	assign g1450 = (((!g8) & (!i_8_) & (!g46) & (!g108) & (!sk[60]) & (g895)) + ((!g8) & (!i_8_) & (!g46) & (!g108) & (sk[60]) & (!g895)) + ((!g8) & (!i_8_) & (!g46) & (!g108) & (sk[60]) & (g895)) + ((!g8) & (!i_8_) & (!g46) & (g108) & (!sk[60]) & (g895)) + ((!g8) & (!i_8_) & (!g46) & (g108) & (sk[60]) & (!g895)) + ((!g8) & (!i_8_) & (!g46) & (g108) & (sk[60]) & (g895)) + ((!g8) & (!i_8_) & (g46) & (!g108) & (!sk[60]) & (g895)) + ((!g8) & (!i_8_) & (g46) & (!g108) & (sk[60]) & (!g895)) + ((!g8) & (!i_8_) & (g46) & (!g108) & (sk[60]) & (g895)) + ((!g8) & (!i_8_) & (g46) & (g108) & (!sk[60]) & (g895)) + ((!g8) & (!i_8_) & (g46) & (g108) & (sk[60]) & (!g895)) + ((!g8) & (!i_8_) & (g46) & (g108) & (sk[60]) & (g895)) + ((!g8) & (i_8_) & (!g46) & (!g108) & (!sk[60]) & (g895)) + ((!g8) & (i_8_) & (!g46) & (!g108) & (sk[60]) & (!g895)) + ((!g8) & (i_8_) & (!g46) & (!g108) & (sk[60]) & (g895)) + ((!g8) & (i_8_) & (!g46) & (g108) & (!sk[60]) & (g895)) + ((!g8) & (i_8_) & (g46) & (!g108) & (!sk[60]) & (g895)) + ((!g8) & (i_8_) & (g46) & (!g108) & (sk[60]) & (!g895)) + ((!g8) & (i_8_) & (g46) & (!g108) & (sk[60]) & (g895)) + ((!g8) & (i_8_) & (g46) & (g108) & (!sk[60]) & (g895)) + ((g8) & (!i_8_) & (!g46) & (!g108) & (!sk[60]) & (!g895)) + ((g8) & (!i_8_) & (!g46) & (!g108) & (!sk[60]) & (g895)) + ((g8) & (!i_8_) & (!g46) & (!g108) & (sk[60]) & (!g895)) + ((g8) & (!i_8_) & (!g46) & (!g108) & (sk[60]) & (g895)) + ((g8) & (!i_8_) & (!g46) & (g108) & (!sk[60]) & (!g895)) + ((g8) & (!i_8_) & (!g46) & (g108) & (!sk[60]) & (g895)) + ((g8) & (!i_8_) & (!g46) & (g108) & (sk[60]) & (!g895)) + ((g8) & (!i_8_) & (!g46) & (g108) & (sk[60]) & (g895)) + ((g8) & (!i_8_) & (g46) & (!g108) & (!sk[60]) & (!g895)) + ((g8) & (!i_8_) & (g46) & (!g108) & (!sk[60]) & (g895)) + ((g8) & (!i_8_) & (g46) & (!g108) & (sk[60]) & (!g895)) + ((g8) & (!i_8_) & (g46) & (!g108) & (sk[60]) & (g895)) + ((g8) & (!i_8_) & (g46) & (g108) & (!sk[60]) & (!g895)) + ((g8) & (!i_8_) & (g46) & (g108) & (!sk[60]) & (g895)) + ((g8) & (!i_8_) & (g46) & (g108) & (sk[60]) & (!g895)) + ((g8) & (!i_8_) & (g46) & (g108) & (sk[60]) & (g895)) + ((g8) & (i_8_) & (!g46) & (!g108) & (!sk[60]) & (!g895)) + ((g8) & (i_8_) & (!g46) & (!g108) & (!sk[60]) & (g895)) + ((g8) & (i_8_) & (!g46) & (!g108) & (sk[60]) & (!g895)) + ((g8) & (i_8_) & (!g46) & (!g108) & (sk[60]) & (g895)) + ((g8) & (i_8_) & (!g46) & (g108) & (!sk[60]) & (!g895)) + ((g8) & (i_8_) & (!g46) & (g108) & (!sk[60]) & (g895)) + ((g8) & (i_8_) & (!g46) & (g108) & (sk[60]) & (!g895)) + ((g8) & (i_8_) & (g46) & (!g108) & (!sk[60]) & (!g895)) + ((g8) & (i_8_) & (g46) & (!g108) & (!sk[60]) & (g895)) + ((g8) & (i_8_) & (g46) & (!g108) & (sk[60]) & (!g895)) + ((g8) & (i_8_) & (g46) & (!g108) & (sk[60]) & (g895)) + ((g8) & (i_8_) & (g46) & (g108) & (!sk[60]) & (!g895)) + ((g8) & (i_8_) & (g46) & (g108) & (!sk[60]) & (g895)));
	assign g1451 = (((!g145) & (!g638) & (!g676) & (!sk[61]) & (!g677) & (g1157)) + ((!g145) & (!g638) & (!g676) & (!sk[61]) & (g677) & (g1157)) + ((!g145) & (!g638) & (g676) & (!sk[61]) & (!g677) & (g1157)) + ((!g145) & (!g638) & (g676) & (!sk[61]) & (g677) & (g1157)) + ((!g145) & (g638) & (!g676) & (!sk[61]) & (!g677) & (g1157)) + ((!g145) & (g638) & (!g676) & (!sk[61]) & (g677) & (g1157)) + ((!g145) & (g638) & (g676) & (!sk[61]) & (!g677) & (g1157)) + ((!g145) & (g638) & (g676) & (!sk[61]) & (g677) & (g1157)) + ((g145) & (!g638) & (!g676) & (!sk[61]) & (!g677) & (!g1157)) + ((g145) & (!g638) & (!g676) & (!sk[61]) & (!g677) & (g1157)) + ((g145) & (!g638) & (!g676) & (!sk[61]) & (g677) & (!g1157)) + ((g145) & (!g638) & (!g676) & (!sk[61]) & (g677) & (g1157)) + ((g145) & (!g638) & (!g676) & (sk[61]) & (!g677) & (!g1157)) + ((g145) & (!g638) & (!g676) & (sk[61]) & (!g677) & (g1157)) + ((g145) & (!g638) & (!g676) & (sk[61]) & (g677) & (!g1157)) + ((g145) & (!g638) & (!g676) & (sk[61]) & (g677) & (g1157)) + ((g145) & (!g638) & (g676) & (!sk[61]) & (!g677) & (!g1157)) + ((g145) & (!g638) & (g676) & (!sk[61]) & (!g677) & (g1157)) + ((g145) & (!g638) & (g676) & (!sk[61]) & (g677) & (!g1157)) + ((g145) & (!g638) & (g676) & (!sk[61]) & (g677) & (g1157)) + ((g145) & (!g638) & (g676) & (sk[61]) & (!g677) & (!g1157)) + ((g145) & (!g638) & (g676) & (sk[61]) & (!g677) & (g1157)) + ((g145) & (!g638) & (g676) & (sk[61]) & (g677) & (!g1157)) + ((g145) & (!g638) & (g676) & (sk[61]) & (g677) & (g1157)) + ((g145) & (g638) & (!g676) & (!sk[61]) & (!g677) & (!g1157)) + ((g145) & (g638) & (!g676) & (!sk[61]) & (!g677) & (g1157)) + ((g145) & (g638) & (!g676) & (!sk[61]) & (g677) & (!g1157)) + ((g145) & (g638) & (!g676) & (!sk[61]) & (g677) & (g1157)) + ((g145) & (g638) & (!g676) & (sk[61]) & (!g677) & (!g1157)) + ((g145) & (g638) & (!g676) & (sk[61]) & (g677) & (!g1157)) + ((g145) & (g638) & (!g676) & (sk[61]) & (g677) & (g1157)) + ((g145) & (g638) & (g676) & (!sk[61]) & (!g677) & (!g1157)) + ((g145) & (g638) & (g676) & (!sk[61]) & (!g677) & (g1157)) + ((g145) & (g638) & (g676) & (!sk[61]) & (g677) & (!g1157)) + ((g145) & (g638) & (g676) & (!sk[61]) & (g677) & (g1157)) + ((g145) & (g638) & (g676) & (sk[61]) & (!g677) & (!g1157)) + ((g145) & (g638) & (g676) & (sk[61]) & (!g677) & (g1157)) + ((g145) & (g638) & (g676) & (sk[61]) & (g677) & (!g1157)) + ((g145) & (g638) & (g676) & (sk[61]) & (g677) & (g1157)));
	assign g1452 = (((!g1445) & (g1447) & (g1448) & (!g1449) & (g1545) & (!g1451)));
	assign g1453 = (((g1028) & (g1206) & (g1347) & (g1392) & (g1443) & (g1452)));
	assign g1454 = (((g613) & (!sk[64]) & (!g555)) + ((g613) & (!sk[64]) & (g555)) + ((g613) & (sk[64]) & (!g555)));
	assign g1455 = (((!i_8_) & (g108) & (!g268) & (!g172) & (!g895) & (!g1454)) + ((!i_8_) & (g108) & (!g268) & (!g172) & (g895) & (!g1454)) + ((!i_8_) & (g108) & (!g268) & (!g172) & (g895) & (g1454)) + ((!i_8_) & (g108) & (!g268) & (g172) & (!g895) & (!g1454)) + ((!i_8_) & (g108) & (!g268) & (g172) & (g895) & (!g1454)) + ((!i_8_) & (g108) & (!g268) & (g172) & (g895) & (g1454)) + ((!i_8_) & (g108) & (g268) & (!g172) & (!g895) & (!g1454)) + ((!i_8_) & (g108) & (g268) & (!g172) & (g895) & (!g1454)) + ((!i_8_) & (g108) & (g268) & (!g172) & (g895) & (g1454)) + ((!i_8_) & (g108) & (g268) & (g172) & (!g895) & (!g1454)) + ((!i_8_) & (g108) & (g268) & (g172) & (g895) & (!g1454)) + ((!i_8_) & (g108) & (g268) & (g172) & (g895) & (g1454)) + ((i_8_) & (g108) & (!g268) & (!g172) & (!g895) & (!g1454)) + ((i_8_) & (g108) & (!g268) & (!g172) & (g895) & (!g1454)) + ((i_8_) & (g108) & (!g268) & (g172) & (!g895) & (!g1454)) + ((i_8_) & (g108) & (!g268) & (g172) & (!g895) & (g1454)) + ((i_8_) & (g108) & (!g268) & (g172) & (g895) & (!g1454)) + ((i_8_) & (g108) & (!g268) & (g172) & (g895) & (g1454)) + ((i_8_) & (g108) & (g268) & (!g172) & (!g895) & (!g1454)) + ((i_8_) & (g108) & (g268) & (!g172) & (!g895) & (g1454)) + ((i_8_) & (g108) & (g268) & (!g172) & (g895) & (!g1454)) + ((i_8_) & (g108) & (g268) & (!g172) & (g895) & (g1454)) + ((i_8_) & (g108) & (g268) & (g172) & (!g895) & (!g1454)) + ((i_8_) & (g108) & (g268) & (g172) & (!g895) & (g1454)) + ((i_8_) & (g108) & (g268) & (g172) & (g895) & (!g1454)) + ((i_8_) & (g108) & (g268) & (g172) & (g895) & (g1454)));
	assign g1456 = (((!i_8_) & (!g100) & (!sk[66]) & (!g270) & (!g554) & (g678)) + ((!i_8_) & (!g100) & (!sk[66]) & (!g270) & (g554) & (g678)) + ((!i_8_) & (!g100) & (!sk[66]) & (g270) & (!g554) & (g678)) + ((!i_8_) & (!g100) & (!sk[66]) & (g270) & (g554) & (g678)) + ((!i_8_) & (g100) & (!sk[66]) & (!g270) & (!g554) & (g678)) + ((!i_8_) & (g100) & (!sk[66]) & (!g270) & (g554) & (g678)) + ((!i_8_) & (g100) & (!sk[66]) & (g270) & (!g554) & (g678)) + ((!i_8_) & (g100) & (!sk[66]) & (g270) & (g554) & (g678)) + ((i_8_) & (!g100) & (!sk[66]) & (!g270) & (!g554) & (!g678)) + ((i_8_) & (!g100) & (!sk[66]) & (!g270) & (!g554) & (g678)) + ((i_8_) & (!g100) & (!sk[66]) & (!g270) & (g554) & (!g678)) + ((i_8_) & (!g100) & (!sk[66]) & (!g270) & (g554) & (g678)) + ((i_8_) & (!g100) & (!sk[66]) & (g270) & (!g554) & (!g678)) + ((i_8_) & (!g100) & (!sk[66]) & (g270) & (!g554) & (g678)) + ((i_8_) & (!g100) & (!sk[66]) & (g270) & (g554) & (!g678)) + ((i_8_) & (!g100) & (!sk[66]) & (g270) & (g554) & (g678)) + ((i_8_) & (g100) & (!sk[66]) & (!g270) & (!g554) & (!g678)) + ((i_8_) & (g100) & (!sk[66]) & (!g270) & (!g554) & (g678)) + ((i_8_) & (g100) & (!sk[66]) & (!g270) & (g554) & (!g678)) + ((i_8_) & (g100) & (!sk[66]) & (!g270) & (g554) & (g678)) + ((i_8_) & (g100) & (!sk[66]) & (g270) & (!g554) & (!g678)) + ((i_8_) & (g100) & (!sk[66]) & (g270) & (!g554) & (g678)) + ((i_8_) & (g100) & (!sk[66]) & (g270) & (g554) & (!g678)) + ((i_8_) & (g100) & (!sk[66]) & (g270) & (g554) & (g678)) + ((i_8_) & (g100) & (sk[66]) & (!g270) & (!g554) & (!g678)) + ((i_8_) & (g100) & (sk[66]) & (!g270) & (!g554) & (g678)) + ((i_8_) & (g100) & (sk[66]) & (!g270) & (g554) & (!g678)) + ((i_8_) & (g100) & (sk[66]) & (!g270) & (g554) & (g678)) + ((i_8_) & (g100) & (sk[66]) & (g270) & (!g554) & (!g678)) + ((i_8_) & (g100) & (sk[66]) & (g270) & (g554) & (!g678)) + ((i_8_) & (g100) & (sk[66]) & (g270) & (g554) & (g678)));
	assign g1457 = (((!g47) & (!sk[67]) & (!g108) & (!g598) & (!g937) & (g1456)) + ((!g47) & (!sk[67]) & (!g108) & (!g598) & (g937) & (g1456)) + ((!g47) & (!sk[67]) & (!g108) & (g598) & (!g937) & (g1456)) + ((!g47) & (!sk[67]) & (!g108) & (g598) & (g937) & (g1456)) + ((!g47) & (!sk[67]) & (g108) & (!g598) & (!g937) & (g1456)) + ((!g47) & (!sk[67]) & (g108) & (!g598) & (g937) & (g1456)) + ((!g47) & (!sk[67]) & (g108) & (g598) & (!g937) & (g1456)) + ((!g47) & (!sk[67]) & (g108) & (g598) & (g937) & (g1456)) + ((!g47) & (sk[67]) & (!g108) & (!g598) & (!g937) & (!g1456)) + ((!g47) & (sk[67]) & (g108) & (!g598) & (!g937) & (!g1456)) + ((g47) & (!sk[67]) & (!g108) & (!g598) & (!g937) & (!g1456)) + ((g47) & (!sk[67]) & (!g108) & (!g598) & (!g937) & (g1456)) + ((g47) & (!sk[67]) & (!g108) & (!g598) & (g937) & (!g1456)) + ((g47) & (!sk[67]) & (!g108) & (!g598) & (g937) & (g1456)) + ((g47) & (!sk[67]) & (!g108) & (g598) & (!g937) & (!g1456)) + ((g47) & (!sk[67]) & (!g108) & (g598) & (!g937) & (g1456)) + ((g47) & (!sk[67]) & (!g108) & (g598) & (g937) & (!g1456)) + ((g47) & (!sk[67]) & (!g108) & (g598) & (g937) & (g1456)) + ((g47) & (!sk[67]) & (g108) & (!g598) & (!g937) & (!g1456)) + ((g47) & (!sk[67]) & (g108) & (!g598) & (!g937) & (g1456)) + ((g47) & (!sk[67]) & (g108) & (!g598) & (g937) & (!g1456)) + ((g47) & (!sk[67]) & (g108) & (!g598) & (g937) & (g1456)) + ((g47) & (!sk[67]) & (g108) & (g598) & (!g937) & (!g1456)) + ((g47) & (!sk[67]) & (g108) & (g598) & (!g937) & (g1456)) + ((g47) & (!sk[67]) & (g108) & (g598) & (g937) & (!g1456)) + ((g47) & (!sk[67]) & (g108) & (g598) & (g937) & (g1456)) + ((g47) & (sk[67]) & (!g108) & (!g598) & (!g937) & (!g1456)));
	assign g1458 = (((!g744) & (g834) & (!g1192) & (!g1359) & (!g1455) & (g1457)));
	assign g1459 = (((!g1003) & (!g1004) & (g1278) & (!g1279) & (g1330) & (g1458)));
	assign g1460 = (((!g101) & (!sk[70]) & (!g531) & (!g996) & (!g997) & (g998)) + ((!g101) & (!sk[70]) & (!g531) & (!g996) & (g997) & (g998)) + ((!g101) & (!sk[70]) & (!g531) & (g996) & (!g997) & (g998)) + ((!g101) & (!sk[70]) & (!g531) & (g996) & (g997) & (g998)) + ((!g101) & (!sk[70]) & (g531) & (!g996) & (!g997) & (g998)) + ((!g101) & (!sk[70]) & (g531) & (!g996) & (g997) & (g998)) + ((!g101) & (!sk[70]) & (g531) & (g996) & (!g997) & (g998)) + ((!g101) & (!sk[70]) & (g531) & (g996) & (g997) & (g998)) + ((!g101) & (sk[70]) & (!g531) & (g996) & (g997) & (!g998)) + ((!g101) & (sk[70]) & (g531) & (g996) & (g997) & (!g998)) + ((g101) & (!sk[70]) & (!g531) & (!g996) & (!g997) & (!g998)) + ((g101) & (!sk[70]) & (!g531) & (!g996) & (!g997) & (g998)) + ((g101) & (!sk[70]) & (!g531) & (!g996) & (g997) & (!g998)) + ((g101) & (!sk[70]) & (!g531) & (!g996) & (g997) & (g998)) + ((g101) & (!sk[70]) & (!g531) & (g996) & (!g997) & (!g998)) + ((g101) & (!sk[70]) & (!g531) & (g996) & (!g997) & (g998)) + ((g101) & (!sk[70]) & (!g531) & (g996) & (g997) & (!g998)) + ((g101) & (!sk[70]) & (!g531) & (g996) & (g997) & (g998)) + ((g101) & (!sk[70]) & (g531) & (!g996) & (!g997) & (!g998)) + ((g101) & (!sk[70]) & (g531) & (!g996) & (!g997) & (g998)) + ((g101) & (!sk[70]) & (g531) & (!g996) & (g997) & (!g998)) + ((g101) & (!sk[70]) & (g531) & (!g996) & (g997) & (g998)) + ((g101) & (!sk[70]) & (g531) & (g996) & (!g997) & (!g998)) + ((g101) & (!sk[70]) & (g531) & (g996) & (!g997) & (g998)) + ((g101) & (!sk[70]) & (g531) & (g996) & (g997) & (!g998)) + ((g101) & (!sk[70]) & (g531) & (g996) & (g997) & (g998)) + ((g101) & (sk[70]) & (!g531) & (g996) & (g997) & (!g998)));
	assign g1461 = (((!i_3_) & (!i_4_) & (g1) & (!i_8_) & (i_6_) & (!i_7_)) + ((!i_3_) & (i_4_) & (g1) & (!i_8_) & (!i_6_) & (!i_7_)) + ((!i_3_) & (i_4_) & (g1) & (!i_8_) & (i_6_) & (!i_7_)));
	assign g1462 = (((!g32) & (!g21) & (!g900) & (sk[72]) & (!g1461)) + ((!g32) & (!g21) & (!g900) & (sk[72]) & (g1461)) + ((!g32) & (!g21) & (g900) & (!sk[72]) & (g1461)) + ((!g32) & (g21) & (!g900) & (!sk[72]) & (!g1461)) + ((!g32) & (g21) & (!g900) & (!sk[72]) & (g1461)) + ((!g32) & (g21) & (!g900) & (sk[72]) & (!g1461)) + ((!g32) & (g21) & (g900) & (!sk[72]) & (!g1461)) + ((!g32) & (g21) & (g900) & (!sk[72]) & (g1461)) + ((g32) & (!g21) & (!g900) & (sk[72]) & (!g1461)) + ((g32) & (!g21) & (!g900) & (sk[72]) & (g1461)) + ((g32) & (!g21) & (g900) & (!sk[72]) & (!g1461)) + ((g32) & (!g21) & (g900) & (!sk[72]) & (g1461)) + ((g32) & (g21) & (!g900) & (!sk[72]) & (!g1461)) + ((g32) & (g21) & (!g900) & (!sk[72]) & (g1461)) + ((g32) & (g21) & (g900) & (!sk[72]) & (!g1461)) + ((g32) & (g21) & (g900) & (!sk[72]) & (g1461)));
	assign g1463 = (((!g101) & (!g534) & (!sk[73]) & (!g983) & (!g984) & (g1462)) + ((!g101) & (!g534) & (!sk[73]) & (!g983) & (g984) & (g1462)) + ((!g101) & (!g534) & (!sk[73]) & (g983) & (!g984) & (g1462)) + ((!g101) & (!g534) & (!sk[73]) & (g983) & (g984) & (g1462)) + ((!g101) & (!g534) & (sk[73]) & (g983) & (g984) & (g1462)) + ((!g101) & (g534) & (!sk[73]) & (!g983) & (!g984) & (g1462)) + ((!g101) & (g534) & (!sk[73]) & (!g983) & (g984) & (g1462)) + ((!g101) & (g534) & (!sk[73]) & (g983) & (!g984) & (g1462)) + ((!g101) & (g534) & (!sk[73]) & (g983) & (g984) & (g1462)) + ((!g101) & (g534) & (sk[73]) & (g983) & (g984) & (g1462)) + ((g101) & (!g534) & (!sk[73]) & (!g983) & (!g984) & (!g1462)) + ((g101) & (!g534) & (!sk[73]) & (!g983) & (!g984) & (g1462)) + ((g101) & (!g534) & (!sk[73]) & (!g983) & (g984) & (!g1462)) + ((g101) & (!g534) & (!sk[73]) & (!g983) & (g984) & (g1462)) + ((g101) & (!g534) & (!sk[73]) & (g983) & (!g984) & (!g1462)) + ((g101) & (!g534) & (!sk[73]) & (g983) & (!g984) & (g1462)) + ((g101) & (!g534) & (!sk[73]) & (g983) & (g984) & (!g1462)) + ((g101) & (!g534) & (!sk[73]) & (g983) & (g984) & (g1462)) + ((g101) & (!g534) & (sk[73]) & (g983) & (g984) & (g1462)) + ((g101) & (g534) & (!sk[73]) & (!g983) & (!g984) & (!g1462)) + ((g101) & (g534) & (!sk[73]) & (!g983) & (!g984) & (g1462)) + ((g101) & (g534) & (!sk[73]) & (!g983) & (g984) & (!g1462)) + ((g101) & (g534) & (!sk[73]) & (!g983) & (g984) & (g1462)) + ((g101) & (g534) & (!sk[73]) & (g983) & (!g984) & (!g1462)) + ((g101) & (g534) & (!sk[73]) & (g983) & (!g984) & (g1462)) + ((g101) & (g534) & (!sk[73]) & (g983) & (g984) & (!g1462)) + ((g101) & (g534) & (!sk[73]) & (g983) & (g984) & (g1462)));
	assign g1464 = (((!g32) & (sk[74]) & (!g1461)) + ((g32) & (!sk[74]) & (!g1461)) + ((g32) & (!sk[74]) & (g1461)));
	assign g1465 = (((!g23) & (!g12) & (g978) & (!sk[75]) & (g1464)) + ((!g23) & (!g12) & (g978) & (sk[75]) & (!g1464)) + ((!g23) & (!g12) & (g978) & (sk[75]) & (g1464)) + ((!g23) & (g12) & (!g978) & (!sk[75]) & (!g1464)) + ((!g23) & (g12) & (!g978) & (!sk[75]) & (g1464)) + ((!g23) & (g12) & (g978) & (!sk[75]) & (!g1464)) + ((!g23) & (g12) & (g978) & (!sk[75]) & (g1464)) + ((!g23) & (g12) & (g978) & (sk[75]) & (g1464)) + ((g23) & (!g12) & (g978) & (!sk[75]) & (!g1464)) + ((g23) & (!g12) & (g978) & (!sk[75]) & (g1464)) + ((g23) & (!g12) & (g978) & (sk[75]) & (g1464)) + ((g23) & (g12) & (!g978) & (!sk[75]) & (!g1464)) + ((g23) & (g12) & (!g978) & (!sk[75]) & (g1464)) + ((g23) & (g12) & (g978) & (!sk[75]) & (!g1464)) + ((g23) & (g12) & (g978) & (!sk[75]) & (g1464)) + ((g23) & (g12) & (g978) & (sk[75]) & (g1464)));
	assign g1466 = (((!sk[76]) & (!g976) & (!g994) & (!g1460) & (!g1463) & (g1465)) + ((!sk[76]) & (!g976) & (!g994) & (!g1460) & (g1463) & (g1465)) + ((!sk[76]) & (!g976) & (!g994) & (g1460) & (!g1463) & (g1465)) + ((!sk[76]) & (!g976) & (!g994) & (g1460) & (g1463) & (g1465)) + ((!sk[76]) & (!g976) & (g994) & (!g1460) & (!g1463) & (g1465)) + ((!sk[76]) & (!g976) & (g994) & (!g1460) & (g1463) & (g1465)) + ((!sk[76]) & (!g976) & (g994) & (g1460) & (!g1463) & (g1465)) + ((!sk[76]) & (!g976) & (g994) & (g1460) & (g1463) & (g1465)) + ((!sk[76]) & (g976) & (!g994) & (!g1460) & (!g1463) & (!g1465)) + ((!sk[76]) & (g976) & (!g994) & (!g1460) & (!g1463) & (g1465)) + ((!sk[76]) & (g976) & (!g994) & (!g1460) & (g1463) & (!g1465)) + ((!sk[76]) & (g976) & (!g994) & (!g1460) & (g1463) & (g1465)) + ((!sk[76]) & (g976) & (!g994) & (g1460) & (!g1463) & (!g1465)) + ((!sk[76]) & (g976) & (!g994) & (g1460) & (!g1463) & (g1465)) + ((!sk[76]) & (g976) & (!g994) & (g1460) & (g1463) & (!g1465)) + ((!sk[76]) & (g976) & (!g994) & (g1460) & (g1463) & (g1465)) + ((!sk[76]) & (g976) & (g994) & (!g1460) & (!g1463) & (!g1465)) + ((!sk[76]) & (g976) & (g994) & (!g1460) & (!g1463) & (g1465)) + ((!sk[76]) & (g976) & (g994) & (!g1460) & (g1463) & (!g1465)) + ((!sk[76]) & (g976) & (g994) & (!g1460) & (g1463) & (g1465)) + ((!sk[76]) & (g976) & (g994) & (g1460) & (!g1463) & (!g1465)) + ((!sk[76]) & (g976) & (g994) & (g1460) & (!g1463) & (g1465)) + ((!sk[76]) & (g976) & (g994) & (g1460) & (g1463) & (!g1465)) + ((!sk[76]) & (g976) & (g994) & (g1460) & (g1463) & (g1465)) + ((sk[76]) & (g976) & (g994) & (g1460) & (g1463) & (g1465)));
	assign g1467 = (((!g73) & (!g1018) & (!g1442) & (!g1453) & (!g1459) & (!g1466)) + ((!g73) & (!g1018) & (!g1442) & (!g1453) & (!g1459) & (g1466)) + ((!g73) & (!g1018) & (!g1442) & (!g1453) & (g1459) & (!g1466)) + ((!g73) & (!g1018) & (!g1442) & (!g1453) & (g1459) & (g1466)) + ((!g73) & (!g1018) & (!g1442) & (g1453) & (!g1459) & (!g1466)) + ((!g73) & (!g1018) & (!g1442) & (g1453) & (!g1459) & (g1466)) + ((!g73) & (!g1018) & (!g1442) & (g1453) & (g1459) & (!g1466)) + ((!g73) & (!g1018) & (!g1442) & (g1453) & (g1459) & (g1466)) + ((!g73) & (!g1018) & (g1442) & (!g1453) & (!g1459) & (!g1466)) + ((!g73) & (!g1018) & (g1442) & (!g1453) & (!g1459) & (g1466)) + ((!g73) & (!g1018) & (g1442) & (!g1453) & (g1459) & (!g1466)) + ((!g73) & (!g1018) & (g1442) & (!g1453) & (g1459) & (g1466)) + ((!g73) & (!g1018) & (g1442) & (g1453) & (!g1459) & (!g1466)) + ((!g73) & (!g1018) & (g1442) & (g1453) & (!g1459) & (g1466)) + ((!g73) & (!g1018) & (g1442) & (g1453) & (g1459) & (!g1466)) + ((!g73) & (!g1018) & (g1442) & (g1453) & (g1459) & (g1466)) + ((!g73) & (g1018) & (!g1442) & (!g1453) & (!g1459) & (!g1466)) + ((!g73) & (g1018) & (!g1442) & (!g1453) & (!g1459) & (g1466)) + ((!g73) & (g1018) & (!g1442) & (!g1453) & (g1459) & (!g1466)) + ((!g73) & (g1018) & (!g1442) & (!g1453) & (g1459) & (g1466)) + ((!g73) & (g1018) & (!g1442) & (g1453) & (!g1459) & (!g1466)) + ((!g73) & (g1018) & (!g1442) & (g1453) & (!g1459) & (g1466)) + ((!g73) & (g1018) & (!g1442) & (g1453) & (g1459) & (!g1466)) + ((!g73) & (g1018) & (!g1442) & (g1453) & (g1459) & (g1466)) + ((!g73) & (g1018) & (g1442) & (!g1453) & (!g1459) & (!g1466)) + ((!g73) & (g1018) & (g1442) & (!g1453) & (!g1459) & (g1466)) + ((!g73) & (g1018) & (g1442) & (!g1453) & (g1459) & (!g1466)) + ((!g73) & (g1018) & (g1442) & (!g1453) & (g1459) & (g1466)) + ((!g73) & (g1018) & (g1442) & (g1453) & (!g1459) & (!g1466)) + ((!g73) & (g1018) & (g1442) & (g1453) & (!g1459) & (g1466)) + ((!g73) & (g1018) & (g1442) & (g1453) & (g1459) & (!g1466)) + ((!g73) & (g1018) & (g1442) & (g1453) & (g1459) & (g1466)) + ((g73) & (g1018) & (!g1442) & (g1453) & (g1459) & (g1466)));
	assign g1468 = (((g31) & (!sk[78]) & (!g64)) + ((g31) & (!sk[78]) & (g64)) + ((g31) & (sk[78]) & (g64)));
	assign g1469 = (((!g7) & (!g25) & (!g3) & (!sk[79]) & (!g131) & (g1468)) + ((!g7) & (!g25) & (!g3) & (!sk[79]) & (g131) & (g1468)) + ((!g7) & (!g25) & (!g3) & (sk[79]) & (!g131) & (!g1468)) + ((!g7) & (!g25) & (!g3) & (sk[79]) & (g131) & (!g1468)) + ((!g7) & (!g25) & (g3) & (!sk[79]) & (!g131) & (g1468)) + ((!g7) & (!g25) & (g3) & (!sk[79]) & (g131) & (g1468)) + ((!g7) & (!g25) & (g3) & (sk[79]) & (!g131) & (!g1468)) + ((!g7) & (!g25) & (g3) & (sk[79]) & (g131) & (!g1468)) + ((!g7) & (g25) & (!g3) & (!sk[79]) & (!g131) & (g1468)) + ((!g7) & (g25) & (!g3) & (!sk[79]) & (g131) & (g1468)) + ((!g7) & (g25) & (!g3) & (sk[79]) & (!g131) & (!g1468)) + ((!g7) & (g25) & (!g3) & (sk[79]) & (!g131) & (g1468)) + ((!g7) & (g25) & (!g3) & (sk[79]) & (g131) & (!g1468)) + ((!g7) & (g25) & (!g3) & (sk[79]) & (g131) & (g1468)) + ((!g7) & (g25) & (g3) & (!sk[79]) & (!g131) & (g1468)) + ((!g7) & (g25) & (g3) & (!sk[79]) & (g131) & (g1468)) + ((!g7) & (g25) & (g3) & (sk[79]) & (!g131) & (!g1468)) + ((!g7) & (g25) & (g3) & (sk[79]) & (!g131) & (g1468)) + ((!g7) & (g25) & (g3) & (sk[79]) & (g131) & (!g1468)) + ((!g7) & (g25) & (g3) & (sk[79]) & (g131) & (g1468)) + ((g7) & (!g25) & (!g3) & (!sk[79]) & (!g131) & (!g1468)) + ((g7) & (!g25) & (!g3) & (!sk[79]) & (!g131) & (g1468)) + ((g7) & (!g25) & (!g3) & (!sk[79]) & (g131) & (!g1468)) + ((g7) & (!g25) & (!g3) & (!sk[79]) & (g131) & (g1468)) + ((g7) & (!g25) & (!g3) & (sk[79]) & (!g131) & (!g1468)) + ((g7) & (!g25) & (!g3) & (sk[79]) & (g131) & (!g1468)) + ((g7) & (!g25) & (g3) & (!sk[79]) & (!g131) & (!g1468)) + ((g7) & (!g25) & (g3) & (!sk[79]) & (!g131) & (g1468)) + ((g7) & (!g25) & (g3) & (!sk[79]) & (g131) & (!g1468)) + ((g7) & (!g25) & (g3) & (!sk[79]) & (g131) & (g1468)) + ((g7) & (!g25) & (g3) & (sk[79]) & (!g131) & (!g1468)) + ((g7) & (g25) & (!g3) & (!sk[79]) & (!g131) & (!g1468)) + ((g7) & (g25) & (!g3) & (!sk[79]) & (!g131) & (g1468)) + ((g7) & (g25) & (!g3) & (!sk[79]) & (g131) & (!g1468)) + ((g7) & (g25) & (!g3) & (!sk[79]) & (g131) & (g1468)) + ((g7) & (g25) & (!g3) & (sk[79]) & (!g131) & (!g1468)) + ((g7) & (g25) & (!g3) & (sk[79]) & (!g131) & (g1468)) + ((g7) & (g25) & (!g3) & (sk[79]) & (g131) & (!g1468)) + ((g7) & (g25) & (!g3) & (sk[79]) & (g131) & (g1468)) + ((g7) & (g25) & (g3) & (!sk[79]) & (!g131) & (!g1468)) + ((g7) & (g25) & (g3) & (!sk[79]) & (!g131) & (g1468)) + ((g7) & (g25) & (g3) & (!sk[79]) & (g131) & (!g1468)) + ((g7) & (g25) & (g3) & (!sk[79]) & (g131) & (g1468)) + ((g7) & (g25) & (g3) & (sk[79]) & (!g131) & (!g1468)) + ((g7) & (g25) & (g3) & (sk[79]) & (!g131) & (g1468)));
	assign g1470 = (((!g12) & (!g101) & (!sk[80]) & (!g971) & (!g974) & (g975)) + ((!g12) & (!g101) & (!sk[80]) & (!g971) & (g974) & (g975)) + ((!g12) & (!g101) & (!sk[80]) & (g971) & (!g974) & (g975)) + ((!g12) & (!g101) & (!sk[80]) & (g971) & (g974) & (g975)) + ((!g12) & (!g101) & (sk[80]) & (g971) & (g974) & (!g975)) + ((!g12) & (g101) & (!sk[80]) & (!g971) & (!g974) & (g975)) + ((!g12) & (g101) & (!sk[80]) & (!g971) & (g974) & (g975)) + ((!g12) & (g101) & (!sk[80]) & (g971) & (!g974) & (g975)) + ((!g12) & (g101) & (!sk[80]) & (g971) & (g974) & (g975)) + ((!g12) & (g101) & (sk[80]) & (g971) & (g974) & (!g975)) + ((g12) & (!g101) & (!sk[80]) & (!g971) & (!g974) & (!g975)) + ((g12) & (!g101) & (!sk[80]) & (!g971) & (!g974) & (g975)) + ((g12) & (!g101) & (!sk[80]) & (!g971) & (g974) & (!g975)) + ((g12) & (!g101) & (!sk[80]) & (!g971) & (g974) & (g975)) + ((g12) & (!g101) & (!sk[80]) & (g971) & (!g974) & (!g975)) + ((g12) & (!g101) & (!sk[80]) & (g971) & (!g974) & (g975)) + ((g12) & (!g101) & (!sk[80]) & (g971) & (g974) & (!g975)) + ((g12) & (!g101) & (!sk[80]) & (g971) & (g974) & (g975)) + ((g12) & (!g101) & (sk[80]) & (g971) & (g974) & (!g975)) + ((g12) & (g101) & (!sk[80]) & (!g971) & (!g974) & (!g975)) + ((g12) & (g101) & (!sk[80]) & (!g971) & (!g974) & (g975)) + ((g12) & (g101) & (!sk[80]) & (!g971) & (g974) & (!g975)) + ((g12) & (g101) & (!sk[80]) & (!g971) & (g974) & (g975)) + ((g12) & (g101) & (!sk[80]) & (g971) & (!g974) & (!g975)) + ((g12) & (g101) & (!sk[80]) & (g971) & (!g974) & (g975)) + ((g12) & (g101) & (!sk[80]) & (g971) & (g974) & (!g975)) + ((g12) & (g101) & (!sk[80]) & (g971) & (g974) & (g975)));
	assign g1471 = (((!sk[81]) & (!g101) & (!g534) & (!g978) & (!g983) & (g984)) + ((!sk[81]) & (!g101) & (!g534) & (!g978) & (g983) & (g984)) + ((!sk[81]) & (!g101) & (!g534) & (g978) & (!g983) & (g984)) + ((!sk[81]) & (!g101) & (!g534) & (g978) & (g983) & (g984)) + ((!sk[81]) & (!g101) & (g534) & (!g978) & (!g983) & (g984)) + ((!sk[81]) & (!g101) & (g534) & (!g978) & (g983) & (g984)) + ((!sk[81]) & (!g101) & (g534) & (g978) & (!g983) & (g984)) + ((!sk[81]) & (!g101) & (g534) & (g978) & (g983) & (g984)) + ((!sk[81]) & (g101) & (!g534) & (!g978) & (!g983) & (!g984)) + ((!sk[81]) & (g101) & (!g534) & (!g978) & (!g983) & (g984)) + ((!sk[81]) & (g101) & (!g534) & (!g978) & (g983) & (!g984)) + ((!sk[81]) & (g101) & (!g534) & (!g978) & (g983) & (g984)) + ((!sk[81]) & (g101) & (!g534) & (g978) & (!g983) & (!g984)) + ((!sk[81]) & (g101) & (!g534) & (g978) & (!g983) & (g984)) + ((!sk[81]) & (g101) & (!g534) & (g978) & (g983) & (!g984)) + ((!sk[81]) & (g101) & (!g534) & (g978) & (g983) & (g984)) + ((!sk[81]) & (g101) & (g534) & (!g978) & (!g983) & (!g984)) + ((!sk[81]) & (g101) & (g534) & (!g978) & (!g983) & (g984)) + ((!sk[81]) & (g101) & (g534) & (!g978) & (g983) & (!g984)) + ((!sk[81]) & (g101) & (g534) & (!g978) & (g983) & (g984)) + ((!sk[81]) & (g101) & (g534) & (g978) & (!g983) & (!g984)) + ((!sk[81]) & (g101) & (g534) & (g978) & (!g983) & (g984)) + ((!sk[81]) & (g101) & (g534) & (g978) & (g983) & (!g984)) + ((!sk[81]) & (g101) & (g534) & (g978) & (g983) & (g984)) + ((sk[81]) & (!g101) & (!g534) & (g978) & (g983) & (g984)) + ((sk[81]) & (!g101) & (g534) & (g978) & (g983) & (g984)) + ((sk[81]) & (g101) & (!g534) & (g978) & (g983) & (g984)));
	assign g1472 = (((!g987) & (g990) & (sk[82]) & (g992)) + ((g987) & (!g990) & (!sk[82]) & (!g992)) + ((g987) & (!g990) & (!sk[82]) & (g992)) + ((g987) & (g990) & (!sk[82]) & (!g992)) + ((g987) & (g990) & (!sk[82]) & (g992)));
	assign g1473 = (((g99) & (!g119) & (!sk[83]) & (!g711)) + ((g99) & (!g119) & (!sk[83]) & (g711)) + ((g99) & (g119) & (!sk[83]) & (!g711)) + ((g99) & (g119) & (!sk[83]) & (g711)) + ((g99) & (g119) & (sk[83]) & (g711)));
	assign g1474 = (((!g101) & (!g299) & (!g745) & (!g898) & (!g1064) & (!g1473)) + ((!g101) & (!g299) & (!g745) & (!g898) & (g1064) & (!g1473)) + ((!g101) & (!g299) & (!g745) & (g898) & (!g1064) & (!g1473)) + ((!g101) & (!g299) & (!g745) & (g898) & (g1064) & (!g1473)) + ((g101) & (!g299) & (!g745) & (!g898) & (g1064) & (!g1473)));
	assign g1475 = (((!g1470) & (!g1471) & (!g1472) & (!g1460) & (!sk[85]) & (g1474)) + ((!g1470) & (!g1471) & (!g1472) & (g1460) & (!sk[85]) & (g1474)) + ((!g1470) & (!g1471) & (g1472) & (!g1460) & (!sk[85]) & (g1474)) + ((!g1470) & (!g1471) & (g1472) & (g1460) & (!sk[85]) & (g1474)) + ((!g1470) & (g1471) & (!g1472) & (!g1460) & (!sk[85]) & (g1474)) + ((!g1470) & (g1471) & (!g1472) & (g1460) & (!sk[85]) & (g1474)) + ((!g1470) & (g1471) & (g1472) & (!g1460) & (!sk[85]) & (g1474)) + ((!g1470) & (g1471) & (g1472) & (g1460) & (!sk[85]) & (g1474)) + ((g1470) & (!g1471) & (!g1472) & (!g1460) & (!sk[85]) & (!g1474)) + ((g1470) & (!g1471) & (!g1472) & (!g1460) & (!sk[85]) & (g1474)) + ((g1470) & (!g1471) & (!g1472) & (g1460) & (!sk[85]) & (!g1474)) + ((g1470) & (!g1471) & (!g1472) & (g1460) & (!sk[85]) & (g1474)) + ((g1470) & (!g1471) & (g1472) & (!g1460) & (!sk[85]) & (!g1474)) + ((g1470) & (!g1471) & (g1472) & (!g1460) & (!sk[85]) & (g1474)) + ((g1470) & (!g1471) & (g1472) & (g1460) & (!sk[85]) & (!g1474)) + ((g1470) & (!g1471) & (g1472) & (g1460) & (!sk[85]) & (g1474)) + ((g1470) & (g1471) & (!g1472) & (!g1460) & (!sk[85]) & (!g1474)) + ((g1470) & (g1471) & (!g1472) & (!g1460) & (!sk[85]) & (g1474)) + ((g1470) & (g1471) & (!g1472) & (g1460) & (!sk[85]) & (!g1474)) + ((g1470) & (g1471) & (!g1472) & (g1460) & (!sk[85]) & (g1474)) + ((g1470) & (g1471) & (g1472) & (!g1460) & (!sk[85]) & (!g1474)) + ((g1470) & (g1471) & (g1472) & (!g1460) & (!sk[85]) & (g1474)) + ((g1470) & (g1471) & (g1472) & (g1460) & (!sk[85]) & (!g1474)) + ((g1470) & (g1471) & (g1472) & (g1460) & (!sk[85]) & (g1474)) + ((g1470) & (g1471) & (g1472) & (g1460) & (sk[85]) & (g1474)));
	assign g1476 = (((!g73) & (!g1018) & (!sk[86]) & (!g1453) & (!g1459) & (g1475)) + ((!g73) & (!g1018) & (!sk[86]) & (!g1453) & (g1459) & (g1475)) + ((!g73) & (!g1018) & (!sk[86]) & (g1453) & (!g1459) & (g1475)) + ((!g73) & (!g1018) & (!sk[86]) & (g1453) & (g1459) & (g1475)) + ((!g73) & (!g1018) & (sk[86]) & (!g1453) & (!g1459) & (!g1475)) + ((!g73) & (!g1018) & (sk[86]) & (!g1453) & (!g1459) & (g1475)) + ((!g73) & (!g1018) & (sk[86]) & (!g1453) & (g1459) & (!g1475)) + ((!g73) & (!g1018) & (sk[86]) & (!g1453) & (g1459) & (g1475)) + ((!g73) & (!g1018) & (sk[86]) & (g1453) & (!g1459) & (!g1475)) + ((!g73) & (!g1018) & (sk[86]) & (g1453) & (!g1459) & (g1475)) + ((!g73) & (!g1018) & (sk[86]) & (g1453) & (g1459) & (!g1475)) + ((!g73) & (!g1018) & (sk[86]) & (g1453) & (g1459) & (g1475)) + ((!g73) & (g1018) & (!sk[86]) & (!g1453) & (!g1459) & (g1475)) + ((!g73) & (g1018) & (!sk[86]) & (!g1453) & (g1459) & (g1475)) + ((!g73) & (g1018) & (!sk[86]) & (g1453) & (!g1459) & (g1475)) + ((!g73) & (g1018) & (!sk[86]) & (g1453) & (g1459) & (g1475)) + ((!g73) & (g1018) & (sk[86]) & (!g1453) & (!g1459) & (!g1475)) + ((!g73) & (g1018) & (sk[86]) & (!g1453) & (!g1459) & (g1475)) + ((!g73) & (g1018) & (sk[86]) & (!g1453) & (g1459) & (!g1475)) + ((!g73) & (g1018) & (sk[86]) & (!g1453) & (g1459) & (g1475)) + ((!g73) & (g1018) & (sk[86]) & (g1453) & (!g1459) & (!g1475)) + ((!g73) & (g1018) & (sk[86]) & (g1453) & (!g1459) & (g1475)) + ((!g73) & (g1018) & (sk[86]) & (g1453) & (g1459) & (!g1475)) + ((!g73) & (g1018) & (sk[86]) & (g1453) & (g1459) & (g1475)) + ((g73) & (!g1018) & (!sk[86]) & (!g1453) & (!g1459) & (!g1475)) + ((g73) & (!g1018) & (!sk[86]) & (!g1453) & (!g1459) & (g1475)) + ((g73) & (!g1018) & (!sk[86]) & (!g1453) & (g1459) & (!g1475)) + ((g73) & (!g1018) & (!sk[86]) & (!g1453) & (g1459) & (g1475)) + ((g73) & (!g1018) & (!sk[86]) & (g1453) & (!g1459) & (!g1475)) + ((g73) & (!g1018) & (!sk[86]) & (g1453) & (!g1459) & (g1475)) + ((g73) & (!g1018) & (!sk[86]) & (g1453) & (g1459) & (!g1475)) + ((g73) & (!g1018) & (!sk[86]) & (g1453) & (g1459) & (g1475)) + ((g73) & (g1018) & (!sk[86]) & (!g1453) & (!g1459) & (!g1475)) + ((g73) & (g1018) & (!sk[86]) & (!g1453) & (!g1459) & (g1475)) + ((g73) & (g1018) & (!sk[86]) & (!g1453) & (g1459) & (!g1475)) + ((g73) & (g1018) & (!sk[86]) & (!g1453) & (g1459) & (g1475)) + ((g73) & (g1018) & (!sk[86]) & (g1453) & (!g1459) & (!g1475)) + ((g73) & (g1018) & (!sk[86]) & (g1453) & (!g1459) & (g1475)) + ((g73) & (g1018) & (!sk[86]) & (g1453) & (g1459) & (!g1475)) + ((g73) & (g1018) & (!sk[86]) & (g1453) & (g1459) & (g1475)) + ((g73) & (g1018) & (sk[86]) & (g1453) & (g1459) & (g1475)));
	assign g1477 = (((!g338) & (!g540) & (!g1286) & (g1607) & (g1353) & (g1410)) + ((g338) & (!g540) & (!g1286) & (g1607) & (g1353) & (g1410)) + ((g338) & (g540) & (!g1286) & (g1607) & (g1353) & (g1410)));
	assign o_27_ = (((!i_1_) & (!i_0_) & (!i_2_) & (!sk[88]) & (!g4) & (g73)) + ((!i_1_) & (!i_0_) & (!i_2_) & (!sk[88]) & (g4) & (g73)) + ((!i_1_) & (!i_0_) & (i_2_) & (!sk[88]) & (!g4) & (g73)) + ((!i_1_) & (!i_0_) & (i_2_) & (!sk[88]) & (g4) & (g73)) + ((!i_1_) & (i_0_) & (!i_2_) & (!sk[88]) & (!g4) & (g73)) + ((!i_1_) & (i_0_) & (!i_2_) & (!sk[88]) & (g4) & (g73)) + ((!i_1_) & (i_0_) & (i_2_) & (!sk[88]) & (!g4) & (g73)) + ((!i_1_) & (i_0_) & (i_2_) & (!sk[88]) & (g4) & (g73)) + ((i_1_) & (!i_0_) & (!i_2_) & (!sk[88]) & (!g4) & (!g73)) + ((i_1_) & (!i_0_) & (!i_2_) & (!sk[88]) & (!g4) & (g73)) + ((i_1_) & (!i_0_) & (!i_2_) & (!sk[88]) & (g4) & (!g73)) + ((i_1_) & (!i_0_) & (!i_2_) & (!sk[88]) & (g4) & (g73)) + ((i_1_) & (!i_0_) & (i_2_) & (!sk[88]) & (!g4) & (!g73)) + ((i_1_) & (!i_0_) & (i_2_) & (!sk[88]) & (!g4) & (g73)) + ((i_1_) & (!i_0_) & (i_2_) & (!sk[88]) & (g4) & (!g73)) + ((i_1_) & (!i_0_) & (i_2_) & (!sk[88]) & (g4) & (g73)) + ((i_1_) & (i_0_) & (!i_2_) & (!sk[88]) & (!g4) & (!g73)) + ((i_1_) & (i_0_) & (!i_2_) & (!sk[88]) & (!g4) & (g73)) + ((i_1_) & (i_0_) & (!i_2_) & (!sk[88]) & (g4) & (!g73)) + ((i_1_) & (i_0_) & (!i_2_) & (!sk[88]) & (g4) & (g73)) + ((i_1_) & (i_0_) & (!i_2_) & (sk[88]) & (g4) & (g73)) + ((i_1_) & (i_0_) & (i_2_) & (!sk[88]) & (!g4) & (!g73)) + ((i_1_) & (i_0_) & (i_2_) & (!sk[88]) & (!g4) & (g73)) + ((i_1_) & (i_0_) & (i_2_) & (!sk[88]) & (g4) & (!g73)) + ((i_1_) & (i_0_) & (i_2_) & (!sk[88]) & (g4) & (g73)));
	assign g1479 = (((!g2) & (!i_8_) & (!i_6_) & (!sk[89]) & (!i_7_) & (g42)) + ((!g2) & (!i_8_) & (!i_6_) & (!sk[89]) & (i_7_) & (g42)) + ((!g2) & (!i_8_) & (i_6_) & (!sk[89]) & (!i_7_) & (g42)) + ((!g2) & (!i_8_) & (i_6_) & (!sk[89]) & (i_7_) & (g42)) + ((!g2) & (!i_8_) & (i_6_) & (sk[89]) & (!i_7_) & (g42)) + ((!g2) & (!i_8_) & (i_6_) & (sk[89]) & (i_7_) & (g42)) + ((!g2) & (i_8_) & (!i_6_) & (!sk[89]) & (!i_7_) & (g42)) + ((!g2) & (i_8_) & (!i_6_) & (!sk[89]) & (i_7_) & (g42)) + ((!g2) & (i_8_) & (i_6_) & (!sk[89]) & (!i_7_) & (g42)) + ((!g2) & (i_8_) & (i_6_) & (!sk[89]) & (i_7_) & (g42)) + ((g2) & (!i_8_) & (!i_6_) & (!sk[89]) & (!i_7_) & (!g42)) + ((g2) & (!i_8_) & (!i_6_) & (!sk[89]) & (!i_7_) & (g42)) + ((g2) & (!i_8_) & (!i_6_) & (!sk[89]) & (i_7_) & (!g42)) + ((g2) & (!i_8_) & (!i_6_) & (!sk[89]) & (i_7_) & (g42)) + ((g2) & (!i_8_) & (i_6_) & (!sk[89]) & (!i_7_) & (!g42)) + ((g2) & (!i_8_) & (i_6_) & (!sk[89]) & (!i_7_) & (g42)) + ((g2) & (!i_8_) & (i_6_) & (!sk[89]) & (i_7_) & (!g42)) + ((g2) & (!i_8_) & (i_6_) & (!sk[89]) & (i_7_) & (g42)) + ((g2) & (!i_8_) & (i_6_) & (sk[89]) & (!i_7_) & (!g42)) + ((g2) & (!i_8_) & (i_6_) & (sk[89]) & (!i_7_) & (g42)) + ((g2) & (!i_8_) & (i_6_) & (sk[89]) & (i_7_) & (g42)) + ((g2) & (i_8_) & (!i_6_) & (!sk[89]) & (!i_7_) & (!g42)) + ((g2) & (i_8_) & (!i_6_) & (!sk[89]) & (!i_7_) & (g42)) + ((g2) & (i_8_) & (!i_6_) & (!sk[89]) & (i_7_) & (!g42)) + ((g2) & (i_8_) & (!i_6_) & (!sk[89]) & (i_7_) & (g42)) + ((g2) & (i_8_) & (i_6_) & (!sk[89]) & (!i_7_) & (!g42)) + ((g2) & (i_8_) & (i_6_) & (!sk[89]) & (!i_7_) & (g42)) + ((g2) & (i_8_) & (i_6_) & (!sk[89]) & (i_7_) & (!g42)) + ((g2) & (i_8_) & (i_6_) & (!sk[89]) & (i_7_) & (g42)));
	assign g1480 = (((!sk[90]) & (!g32) & (!g75) & (g1468) & (g1479)) + ((!sk[90]) & (!g32) & (g75) & (!g1468) & (!g1479)) + ((!sk[90]) & (!g32) & (g75) & (!g1468) & (g1479)) + ((!sk[90]) & (!g32) & (g75) & (g1468) & (!g1479)) + ((!sk[90]) & (!g32) & (g75) & (g1468) & (g1479)) + ((!sk[90]) & (g32) & (!g75) & (g1468) & (!g1479)) + ((!sk[90]) & (g32) & (!g75) & (g1468) & (g1479)) + ((!sk[90]) & (g32) & (g75) & (!g1468) & (!g1479)) + ((!sk[90]) & (g32) & (g75) & (!g1468) & (g1479)) + ((!sk[90]) & (g32) & (g75) & (g1468) & (!g1479)) + ((!sk[90]) & (g32) & (g75) & (g1468) & (g1479)) + ((sk[90]) & (!g32) & (!g75) & (!g1468) & (!g1479)));
	assign g1481 = (((!i_3_) & (!i_4_) & (!i_6_) & (!i_7_) & (!sk[91]) & (g29)) + ((!i_3_) & (!i_4_) & (!i_6_) & (i_7_) & (!sk[91]) & (g29)) + ((!i_3_) & (!i_4_) & (i_6_) & (!i_7_) & (!sk[91]) & (g29)) + ((!i_3_) & (!i_4_) & (i_6_) & (i_7_) & (!sk[91]) & (g29)) + ((!i_3_) & (i_4_) & (!i_6_) & (!i_7_) & (!sk[91]) & (g29)) + ((!i_3_) & (i_4_) & (!i_6_) & (i_7_) & (!sk[91]) & (g29)) + ((!i_3_) & (i_4_) & (i_6_) & (!i_7_) & (!sk[91]) & (g29)) + ((!i_3_) & (i_4_) & (i_6_) & (!i_7_) & (sk[91]) & (g29)) + ((!i_3_) & (i_4_) & (i_6_) & (i_7_) & (!sk[91]) & (g29)) + ((i_3_) & (!i_4_) & (!i_6_) & (!i_7_) & (!sk[91]) & (!g29)) + ((i_3_) & (!i_4_) & (!i_6_) & (!i_7_) & (!sk[91]) & (g29)) + ((i_3_) & (!i_4_) & (!i_6_) & (i_7_) & (!sk[91]) & (!g29)) + ((i_3_) & (!i_4_) & (!i_6_) & (i_7_) & (!sk[91]) & (g29)) + ((i_3_) & (!i_4_) & (i_6_) & (!i_7_) & (!sk[91]) & (!g29)) + ((i_3_) & (!i_4_) & (i_6_) & (!i_7_) & (!sk[91]) & (g29)) + ((i_3_) & (!i_4_) & (i_6_) & (i_7_) & (!sk[91]) & (!g29)) + ((i_3_) & (!i_4_) & (i_6_) & (i_7_) & (!sk[91]) & (g29)) + ((i_3_) & (i_4_) & (!i_6_) & (!i_7_) & (!sk[91]) & (!g29)) + ((i_3_) & (i_4_) & (!i_6_) & (!i_7_) & (!sk[91]) & (g29)) + ((i_3_) & (i_4_) & (!i_6_) & (i_7_) & (!sk[91]) & (!g29)) + ((i_3_) & (i_4_) & (!i_6_) & (i_7_) & (!sk[91]) & (g29)) + ((i_3_) & (i_4_) & (i_6_) & (!i_7_) & (!sk[91]) & (!g29)) + ((i_3_) & (i_4_) & (i_6_) & (!i_7_) & (!sk[91]) & (g29)) + ((i_3_) & (i_4_) & (i_6_) & (i_7_) & (!sk[91]) & (!g29)) + ((i_3_) & (i_4_) & (i_6_) & (i_7_) & (!sk[91]) & (g29)));
	assign g1482 = (((!g32) & (!g20) & (!sk[92]) & (!g75) & (!g1468) & (g1481)) + ((!g32) & (!g20) & (!sk[92]) & (!g75) & (g1468) & (g1481)) + ((!g32) & (!g20) & (!sk[92]) & (g75) & (!g1468) & (g1481)) + ((!g32) & (!g20) & (!sk[92]) & (g75) & (g1468) & (g1481)) + ((!g32) & (!g20) & (sk[92]) & (!g75) & (!g1468) & (!g1481)) + ((!g32) & (g20) & (!sk[92]) & (!g75) & (!g1468) & (g1481)) + ((!g32) & (g20) & (!sk[92]) & (!g75) & (g1468) & (g1481)) + ((!g32) & (g20) & (!sk[92]) & (g75) & (!g1468) & (g1481)) + ((!g32) & (g20) & (!sk[92]) & (g75) & (g1468) & (g1481)) + ((!g32) & (g20) & (sk[92]) & (!g75) & (!g1468) & (!g1481)) + ((!g32) & (g20) & (sk[92]) & (!g75) & (g1468) & (!g1481)) + ((!g32) & (g20) & (sk[92]) & (g75) & (!g1468) & (!g1481)) + ((!g32) & (g20) & (sk[92]) & (g75) & (g1468) & (!g1481)) + ((g32) & (!g20) & (!sk[92]) & (!g75) & (!g1468) & (!g1481)) + ((g32) & (!g20) & (!sk[92]) & (!g75) & (!g1468) & (g1481)) + ((g32) & (!g20) & (!sk[92]) & (!g75) & (g1468) & (!g1481)) + ((g32) & (!g20) & (!sk[92]) & (!g75) & (g1468) & (g1481)) + ((g32) & (!g20) & (!sk[92]) & (g75) & (!g1468) & (!g1481)) + ((g32) & (!g20) & (!sk[92]) & (g75) & (!g1468) & (g1481)) + ((g32) & (!g20) & (!sk[92]) & (g75) & (g1468) & (!g1481)) + ((g32) & (!g20) & (!sk[92]) & (g75) & (g1468) & (g1481)) + ((g32) & (g20) & (!sk[92]) & (!g75) & (!g1468) & (!g1481)) + ((g32) & (g20) & (!sk[92]) & (!g75) & (!g1468) & (g1481)) + ((g32) & (g20) & (!sk[92]) & (!g75) & (g1468) & (!g1481)) + ((g32) & (g20) & (!sk[92]) & (!g75) & (g1468) & (g1481)) + ((g32) & (g20) & (!sk[92]) & (g75) & (!g1468) & (!g1481)) + ((g32) & (g20) & (!sk[92]) & (g75) & (!g1468) & (g1481)) + ((g32) & (g20) & (!sk[92]) & (g75) & (g1468) & (!g1481)) + ((g32) & (g20) & (!sk[92]) & (g75) & (g1468) & (g1481)) + ((g32) & (g20) & (sk[92]) & (!g75) & (!g1468) & (!g1481)) + ((g32) & (g20) & (sk[92]) & (!g75) & (g1468) & (!g1481)) + ((g32) & (g20) & (sk[92]) & (g75) & (!g1468) & (!g1481)) + ((g32) & (g20) & (sk[92]) & (g75) & (g1468) & (!g1481)));
	assign g1483 = (((!i_3_) & (!i_4_) & (!sk[93]) & (g30) & (g29)) + ((!i_3_) & (i_4_) & (!sk[93]) & (!g30) & (!g29)) + ((!i_3_) & (i_4_) & (!sk[93]) & (!g30) & (g29)) + ((!i_3_) & (i_4_) & (!sk[93]) & (g30) & (!g29)) + ((!i_3_) & (i_4_) & (!sk[93]) & (g30) & (g29)) + ((!i_3_) & (i_4_) & (sk[93]) & (g30) & (g29)) + ((i_3_) & (!i_4_) & (!sk[93]) & (g30) & (!g29)) + ((i_3_) & (!i_4_) & (!sk[93]) & (g30) & (g29)) + ((i_3_) & (i_4_) & (!sk[93]) & (!g30) & (!g29)) + ((i_3_) & (i_4_) & (!sk[93]) & (!g30) & (g29)) + ((i_3_) & (i_4_) & (!sk[93]) & (g30) & (!g29)) + ((i_3_) & (i_4_) & (!sk[93]) & (g30) & (g29)));
	assign g1484 = (((!g32) & (!g19) & (!g75) & (!sk[94]) & (!g1468) & (g1483)) + ((!g32) & (!g19) & (!g75) & (!sk[94]) & (g1468) & (g1483)) + ((!g32) & (!g19) & (!g75) & (sk[94]) & (!g1468) & (!g1483)) + ((!g32) & (!g19) & (!g75) & (sk[94]) & (g1468) & (!g1483)) + ((!g32) & (!g19) & (g75) & (!sk[94]) & (!g1468) & (g1483)) + ((!g32) & (!g19) & (g75) & (!sk[94]) & (g1468) & (g1483)) + ((!g32) & (!g19) & (g75) & (sk[94]) & (!g1468) & (!g1483)) + ((!g32) & (!g19) & (g75) & (sk[94]) & (g1468) & (!g1483)) + ((!g32) & (g19) & (!g75) & (!sk[94]) & (!g1468) & (g1483)) + ((!g32) & (g19) & (!g75) & (!sk[94]) & (g1468) & (g1483)) + ((!g32) & (g19) & (!g75) & (sk[94]) & (!g1468) & (!g1483)) + ((!g32) & (g19) & (g75) & (!sk[94]) & (!g1468) & (g1483)) + ((!g32) & (g19) & (g75) & (!sk[94]) & (g1468) & (g1483)) + ((g32) & (!g19) & (!g75) & (!sk[94]) & (!g1468) & (!g1483)) + ((g32) & (!g19) & (!g75) & (!sk[94]) & (!g1468) & (g1483)) + ((g32) & (!g19) & (!g75) & (!sk[94]) & (g1468) & (!g1483)) + ((g32) & (!g19) & (!g75) & (!sk[94]) & (g1468) & (g1483)) + ((g32) & (!g19) & (!g75) & (sk[94]) & (!g1468) & (!g1483)) + ((g32) & (!g19) & (!g75) & (sk[94]) & (g1468) & (!g1483)) + ((g32) & (!g19) & (g75) & (!sk[94]) & (!g1468) & (!g1483)) + ((g32) & (!g19) & (g75) & (!sk[94]) & (!g1468) & (g1483)) + ((g32) & (!g19) & (g75) & (!sk[94]) & (g1468) & (!g1483)) + ((g32) & (!g19) & (g75) & (!sk[94]) & (g1468) & (g1483)) + ((g32) & (!g19) & (g75) & (sk[94]) & (!g1468) & (!g1483)) + ((g32) & (!g19) & (g75) & (sk[94]) & (g1468) & (!g1483)) + ((g32) & (g19) & (!g75) & (!sk[94]) & (!g1468) & (!g1483)) + ((g32) & (g19) & (!g75) & (!sk[94]) & (!g1468) & (g1483)) + ((g32) & (g19) & (!g75) & (!sk[94]) & (g1468) & (!g1483)) + ((g32) & (g19) & (!g75) & (!sk[94]) & (g1468) & (g1483)) + ((g32) & (g19) & (g75) & (!sk[94]) & (!g1468) & (!g1483)) + ((g32) & (g19) & (g75) & (!sk[94]) & (!g1468) & (g1483)) + ((g32) & (g19) & (g75) & (!sk[94]) & (g1468) & (!g1483)) + ((g32) & (g19) & (g75) & (!sk[94]) & (g1468) & (g1483)));
	assign g1485 = (((!sk[95]) & (!g19) & (!g20) & (g1479) & (g1484)) + ((!sk[95]) & (!g19) & (g20) & (!g1479) & (!g1484)) + ((!sk[95]) & (!g19) & (g20) & (!g1479) & (g1484)) + ((!sk[95]) & (!g19) & (g20) & (g1479) & (!g1484)) + ((!sk[95]) & (!g19) & (g20) & (g1479) & (g1484)) + ((!sk[95]) & (g19) & (!g20) & (g1479) & (!g1484)) + ((!sk[95]) & (g19) & (!g20) & (g1479) & (g1484)) + ((!sk[95]) & (g19) & (g20) & (!g1479) & (!g1484)) + ((!sk[95]) & (g19) & (g20) & (!g1479) & (g1484)) + ((!sk[95]) & (g19) & (g20) & (g1479) & (!g1484)) + ((!sk[95]) & (g19) & (g20) & (g1479) & (g1484)) + ((sk[95]) & (!g19) & (!g20) & (!g1479) & (g1484)) + ((sk[95]) & (!g19) & (g20) & (!g1479) & (g1484)) + ((sk[95]) & (!g19) & (g20) & (g1479) & (g1484)) + ((sk[95]) & (g19) & (!g20) & (!g1479) & (g1484)) + ((sk[95]) & (g19) & (g20) & (!g1479) & (g1484)));
	assign g1486 = (((!sk[96]) & (!g16) & (!g1480) & (g1482) & (g1485)) + ((!sk[96]) & (!g16) & (g1480) & (!g1482) & (!g1485)) + ((!sk[96]) & (!g16) & (g1480) & (!g1482) & (g1485)) + ((!sk[96]) & (!g16) & (g1480) & (g1482) & (!g1485)) + ((!sk[96]) & (!g16) & (g1480) & (g1482) & (g1485)) + ((!sk[96]) & (g16) & (!g1480) & (g1482) & (!g1485)) + ((!sk[96]) & (g16) & (!g1480) & (g1482) & (g1485)) + ((!sk[96]) & (g16) & (g1480) & (!g1482) & (!g1485)) + ((!sk[96]) & (g16) & (g1480) & (!g1482) & (g1485)) + ((!sk[96]) & (g16) & (g1480) & (g1482) & (!g1485)) + ((!sk[96]) & (g16) & (g1480) & (g1482) & (g1485)) + ((sk[96]) & (!g16) & (g1480) & (g1482) & (g1485)) + ((sk[96]) & (g16) & (!g1480) & (g1482) & (g1485)) + ((sk[96]) & (g16) & (g1480) & (g1482) & (g1485)));
	assign g1487 = (((!sk[97]) & (i_3_) & (!i_4_) & (!g29)) + ((!sk[97]) & (i_3_) & (!i_4_) & (g29)) + ((!sk[97]) & (i_3_) & (i_4_) & (!g29)) + ((!sk[97]) & (i_3_) & (i_4_) & (g29)) + ((sk[97]) & (!i_3_) & (!i_4_) & (g29)));
	assign g1488 = (((!g5) & (!g61) & (g62) & (!sk[98]) & (g111)) + ((!g5) & (g61) & (!g62) & (!sk[98]) & (!g111)) + ((!g5) & (g61) & (!g62) & (!sk[98]) & (g111)) + ((!g5) & (g61) & (g62) & (!sk[98]) & (!g111)) + ((!g5) & (g61) & (g62) & (!sk[98]) & (g111)) + ((g5) & (!g61) & (g62) & (!sk[98]) & (!g111)) + ((g5) & (!g61) & (g62) & (!sk[98]) & (g111)) + ((g5) & (!g61) & (g62) & (sk[98]) & (g111)) + ((g5) & (g61) & (!g62) & (!sk[98]) & (!g111)) + ((g5) & (g61) & (!g62) & (!sk[98]) & (g111)) + ((g5) & (g61) & (!g62) & (sk[98]) & (g111)) + ((g5) & (g61) & (g62) & (!sk[98]) & (!g111)) + ((g5) & (g61) & (g62) & (!sk[98]) & (g111)) + ((g5) & (g61) & (g62) & (sk[98]) & (g111)));
	assign g1489 = (((!i_7_) & (!sk[99]) & (!g141) & (!g1487) & (!g63) & (g1488)) + ((!i_7_) & (!sk[99]) & (!g141) & (!g1487) & (g63) & (g1488)) + ((!i_7_) & (!sk[99]) & (!g141) & (g1487) & (!g63) & (g1488)) + ((!i_7_) & (!sk[99]) & (!g141) & (g1487) & (g63) & (g1488)) + ((!i_7_) & (!sk[99]) & (g141) & (!g1487) & (!g63) & (g1488)) + ((!i_7_) & (!sk[99]) & (g141) & (!g1487) & (g63) & (g1488)) + ((!i_7_) & (!sk[99]) & (g141) & (g1487) & (!g63) & (g1488)) + ((!i_7_) & (!sk[99]) & (g141) & (g1487) & (g63) & (g1488)) + ((!i_7_) & (sk[99]) & (!g141) & (!g1487) & (!g63) & (!g1488)) + ((!i_7_) & (sk[99]) & (!g141) & (!g1487) & (g63) & (!g1488)) + ((!i_7_) & (sk[99]) & (g141) & (!g1487) & (!g63) & (!g1488)) + ((i_7_) & (!sk[99]) & (!g141) & (!g1487) & (!g63) & (!g1488)) + ((i_7_) & (!sk[99]) & (!g141) & (!g1487) & (!g63) & (g1488)) + ((i_7_) & (!sk[99]) & (!g141) & (!g1487) & (g63) & (!g1488)) + ((i_7_) & (!sk[99]) & (!g141) & (!g1487) & (g63) & (g1488)) + ((i_7_) & (!sk[99]) & (!g141) & (g1487) & (!g63) & (!g1488)) + ((i_7_) & (!sk[99]) & (!g141) & (g1487) & (!g63) & (g1488)) + ((i_7_) & (!sk[99]) & (!g141) & (g1487) & (g63) & (!g1488)) + ((i_7_) & (!sk[99]) & (!g141) & (g1487) & (g63) & (g1488)) + ((i_7_) & (!sk[99]) & (g141) & (!g1487) & (!g63) & (!g1488)) + ((i_7_) & (!sk[99]) & (g141) & (!g1487) & (!g63) & (g1488)) + ((i_7_) & (!sk[99]) & (g141) & (!g1487) & (g63) & (!g1488)) + ((i_7_) & (!sk[99]) & (g141) & (!g1487) & (g63) & (g1488)) + ((i_7_) & (!sk[99]) & (g141) & (g1487) & (!g63) & (!g1488)) + ((i_7_) & (!sk[99]) & (g141) & (g1487) & (!g63) & (g1488)) + ((i_7_) & (!sk[99]) & (g141) & (g1487) & (g63) & (!g1488)) + ((i_7_) & (!sk[99]) & (g141) & (g1487) & (g63) & (g1488)) + ((i_7_) & (sk[99]) & (!g141) & (!g1487) & (!g63) & (!g1488)) + ((i_7_) & (sk[99]) & (!g141) & (!g1487) & (g63) & (!g1488)) + ((i_7_) & (sk[99]) & (!g141) & (g1487) & (!g63) & (!g1488)) + ((i_7_) & (sk[99]) & (!g141) & (g1487) & (g63) & (!g1488)) + ((i_7_) & (sk[99]) & (g141) & (!g1487) & (!g63) & (!g1488)) + ((i_7_) & (sk[99]) & (g141) & (g1487) & (!g63) & (!g1488)));
	assign g1490 = (((!g19) & (!g20) & (!sk[100]) & (!g16) & (!g78) & (g1489)) + ((!g19) & (!g20) & (!sk[100]) & (!g16) & (g78) & (g1489)) + ((!g19) & (!g20) & (!sk[100]) & (g16) & (!g78) & (g1489)) + ((!g19) & (!g20) & (!sk[100]) & (g16) & (g78) & (g1489)) + ((!g19) & (!g20) & (sk[100]) & (!g16) & (!g78) & (g1489)) + ((!g19) & (!g20) & (sk[100]) & (g16) & (!g78) & (g1489)) + ((!g19) & (g20) & (!sk[100]) & (!g16) & (!g78) & (g1489)) + ((!g19) & (g20) & (!sk[100]) & (!g16) & (g78) & (g1489)) + ((!g19) & (g20) & (!sk[100]) & (g16) & (!g78) & (g1489)) + ((!g19) & (g20) & (!sk[100]) & (g16) & (g78) & (g1489)) + ((!g19) & (g20) & (sk[100]) & (!g16) & (!g78) & (g1489)) + ((!g19) & (g20) & (sk[100]) & (g16) & (!g78) & (g1489)) + ((!g19) & (g20) & (sk[100]) & (g16) & (g78) & (g1489)) + ((g19) & (!g20) & (!sk[100]) & (!g16) & (!g78) & (!g1489)) + ((g19) & (!g20) & (!sk[100]) & (!g16) & (!g78) & (g1489)) + ((g19) & (!g20) & (!sk[100]) & (!g16) & (g78) & (!g1489)) + ((g19) & (!g20) & (!sk[100]) & (!g16) & (g78) & (g1489)) + ((g19) & (!g20) & (!sk[100]) & (g16) & (!g78) & (!g1489)) + ((g19) & (!g20) & (!sk[100]) & (g16) & (!g78) & (g1489)) + ((g19) & (!g20) & (!sk[100]) & (g16) & (g78) & (!g1489)) + ((g19) & (!g20) & (!sk[100]) & (g16) & (g78) & (g1489)) + ((g19) & (!g20) & (sk[100]) & (!g16) & (!g78) & (g1489)) + ((g19) & (!g20) & (sk[100]) & (g16) & (!g78) & (g1489)) + ((g19) & (g20) & (!sk[100]) & (!g16) & (!g78) & (!g1489)) + ((g19) & (g20) & (!sk[100]) & (!g16) & (!g78) & (g1489)) + ((g19) & (g20) & (!sk[100]) & (!g16) & (g78) & (!g1489)) + ((g19) & (g20) & (!sk[100]) & (!g16) & (g78) & (g1489)) + ((g19) & (g20) & (!sk[100]) & (g16) & (!g78) & (!g1489)) + ((g19) & (g20) & (!sk[100]) & (g16) & (!g78) & (g1489)) + ((g19) & (g20) & (!sk[100]) & (g16) & (g78) & (!g1489)) + ((g19) & (g20) & (!sk[100]) & (g16) & (g78) & (g1489)) + ((g19) & (g20) & (sk[100]) & (!g16) & (!g78) & (g1489)) + ((g19) & (g20) & (sk[100]) & (g16) & (!g78) & (g1489)));
	assign g1491 = (((!g30) & (!g61) & (!sk[101]) & (!g73) & (!g1486) & (g1490)) + ((!g30) & (!g61) & (!sk[101]) & (!g73) & (g1486) & (g1490)) + ((!g30) & (!g61) & (!sk[101]) & (g73) & (!g1486) & (g1490)) + ((!g30) & (!g61) & (!sk[101]) & (g73) & (g1486) & (g1490)) + ((!g30) & (!g61) & (sk[101]) & (!g73) & (!g1486) & (!g1490)) + ((!g30) & (!g61) & (sk[101]) & (!g73) & (!g1486) & (g1490)) + ((!g30) & (!g61) & (sk[101]) & (!g73) & (g1486) & (!g1490)) + ((!g30) & (!g61) & (sk[101]) & (!g73) & (g1486) & (g1490)) + ((!g30) & (!g61) & (sk[101]) & (g73) & (g1486) & (g1490)) + ((!g30) & (g61) & (!sk[101]) & (!g73) & (!g1486) & (g1490)) + ((!g30) & (g61) & (!sk[101]) & (!g73) & (g1486) & (g1490)) + ((!g30) & (g61) & (!sk[101]) & (g73) & (!g1486) & (g1490)) + ((!g30) & (g61) & (!sk[101]) & (g73) & (g1486) & (g1490)) + ((!g30) & (g61) & (sk[101]) & (!g73) & (!g1486) & (!g1490)) + ((!g30) & (g61) & (sk[101]) & (!g73) & (!g1486) & (g1490)) + ((!g30) & (g61) & (sk[101]) & (!g73) & (g1486) & (!g1490)) + ((!g30) & (g61) & (sk[101]) & (!g73) & (g1486) & (g1490)) + ((g30) & (!g61) & (!sk[101]) & (!g73) & (!g1486) & (!g1490)) + ((g30) & (!g61) & (!sk[101]) & (!g73) & (!g1486) & (g1490)) + ((g30) & (!g61) & (!sk[101]) & (!g73) & (g1486) & (!g1490)) + ((g30) & (!g61) & (!sk[101]) & (!g73) & (g1486) & (g1490)) + ((g30) & (!g61) & (!sk[101]) & (g73) & (!g1486) & (!g1490)) + ((g30) & (!g61) & (!sk[101]) & (g73) & (!g1486) & (g1490)) + ((g30) & (!g61) & (!sk[101]) & (g73) & (g1486) & (!g1490)) + ((g30) & (!g61) & (!sk[101]) & (g73) & (g1486) & (g1490)) + ((g30) & (!g61) & (sk[101]) & (!g73) & (!g1486) & (!g1490)) + ((g30) & (!g61) & (sk[101]) & (!g73) & (!g1486) & (g1490)) + ((g30) & (!g61) & (sk[101]) & (!g73) & (g1486) & (!g1490)) + ((g30) & (!g61) & (sk[101]) & (!g73) & (g1486) & (g1490)) + ((g30) & (!g61) & (sk[101]) & (g73) & (g1486) & (g1490)) + ((g30) & (g61) & (!sk[101]) & (!g73) & (!g1486) & (!g1490)) + ((g30) & (g61) & (!sk[101]) & (!g73) & (!g1486) & (g1490)) + ((g30) & (g61) & (!sk[101]) & (!g73) & (g1486) & (!g1490)) + ((g30) & (g61) & (!sk[101]) & (!g73) & (g1486) & (g1490)) + ((g30) & (g61) & (!sk[101]) & (g73) & (!g1486) & (!g1490)) + ((g30) & (g61) & (!sk[101]) & (g73) & (!g1486) & (g1490)) + ((g30) & (g61) & (!sk[101]) & (g73) & (g1486) & (!g1490)) + ((g30) & (g61) & (!sk[101]) & (g73) & (g1486) & (g1490)) + ((g30) & (g61) & (sk[101]) & (!g73) & (!g1486) & (!g1490)) + ((g30) & (g61) & (sk[101]) & (!g73) & (!g1486) & (g1490)) + ((g30) & (g61) & (sk[101]) & (!g73) & (g1486) & (!g1490)) + ((g30) & (g61) & (sk[101]) & (!g73) & (g1486) & (g1490)) + ((g30) & (g61) & (sk[101]) & (g73) & (g1486) & (g1490)));
	assign g1492 = (((!g14) & (!g4) & (!g29) & (!g39) & (!sk[102]) & (g1480)) + ((!g14) & (!g4) & (!g29) & (g39) & (!sk[102]) & (g1480)) + ((!g14) & (!g4) & (g29) & (!g39) & (!sk[102]) & (g1480)) + ((!g14) & (!g4) & (g29) & (g39) & (!sk[102]) & (g1480)) + ((!g14) & (g4) & (!g29) & (!g39) & (!sk[102]) & (g1480)) + ((!g14) & (g4) & (!g29) & (g39) & (!sk[102]) & (g1480)) + ((!g14) & (g4) & (g29) & (!g39) & (!sk[102]) & (g1480)) + ((!g14) & (g4) & (g29) & (g39) & (!sk[102]) & (g1480)) + ((!g14) & (g4) & (g29) & (g39) & (sk[102]) & (!g1480)) + ((!g14) & (g4) & (g29) & (g39) & (sk[102]) & (g1480)) + ((g14) & (!g4) & (!g29) & (!g39) & (!sk[102]) & (!g1480)) + ((g14) & (!g4) & (!g29) & (!g39) & (!sk[102]) & (g1480)) + ((g14) & (!g4) & (!g29) & (!g39) & (sk[102]) & (!g1480)) + ((g14) & (!g4) & (!g29) & (g39) & (!sk[102]) & (!g1480)) + ((g14) & (!g4) & (!g29) & (g39) & (!sk[102]) & (g1480)) + ((g14) & (!g4) & (!g29) & (g39) & (sk[102]) & (!g1480)) + ((g14) & (!g4) & (g29) & (!g39) & (!sk[102]) & (!g1480)) + ((g14) & (!g4) & (g29) & (!g39) & (!sk[102]) & (g1480)) + ((g14) & (!g4) & (g29) & (!g39) & (sk[102]) & (!g1480)) + ((g14) & (!g4) & (g29) & (g39) & (!sk[102]) & (!g1480)) + ((g14) & (!g4) & (g29) & (g39) & (!sk[102]) & (g1480)) + ((g14) & (!g4) & (g29) & (g39) & (sk[102]) & (!g1480)) + ((g14) & (g4) & (!g29) & (!g39) & (!sk[102]) & (!g1480)) + ((g14) & (g4) & (!g29) & (!g39) & (!sk[102]) & (g1480)) + ((g14) & (g4) & (!g29) & (!g39) & (sk[102]) & (!g1480)) + ((g14) & (g4) & (!g29) & (g39) & (!sk[102]) & (!g1480)) + ((g14) & (g4) & (!g29) & (g39) & (!sk[102]) & (g1480)) + ((g14) & (g4) & (!g29) & (g39) & (sk[102]) & (!g1480)) + ((g14) & (g4) & (g29) & (!g39) & (!sk[102]) & (!g1480)) + ((g14) & (g4) & (g29) & (!g39) & (!sk[102]) & (g1480)) + ((g14) & (g4) & (g29) & (!g39) & (sk[102]) & (!g1480)) + ((g14) & (g4) & (g29) & (g39) & (!sk[102]) & (!g1480)) + ((g14) & (g4) & (g29) & (g39) & (!sk[102]) & (g1480)) + ((g14) & (g4) & (g29) & (g39) & (sk[102]) & (!g1480)) + ((g14) & (g4) & (g29) & (g39) & (sk[102]) & (g1480)));
	assign g1493 = (((!sk[103]) & (!g8) & (!g32) & (!g75) & (!g1468) & (g1479)) + ((!sk[103]) & (!g8) & (!g32) & (!g75) & (g1468) & (g1479)) + ((!sk[103]) & (!g8) & (!g32) & (g75) & (!g1468) & (g1479)) + ((!sk[103]) & (!g8) & (!g32) & (g75) & (g1468) & (g1479)) + ((!sk[103]) & (!g8) & (g32) & (!g75) & (!g1468) & (g1479)) + ((!sk[103]) & (!g8) & (g32) & (!g75) & (g1468) & (g1479)) + ((!sk[103]) & (!g8) & (g32) & (g75) & (!g1468) & (g1479)) + ((!sk[103]) & (!g8) & (g32) & (g75) & (g1468) & (g1479)) + ((!sk[103]) & (g8) & (!g32) & (!g75) & (!g1468) & (!g1479)) + ((!sk[103]) & (g8) & (!g32) & (!g75) & (!g1468) & (g1479)) + ((!sk[103]) & (g8) & (!g32) & (!g75) & (g1468) & (!g1479)) + ((!sk[103]) & (g8) & (!g32) & (!g75) & (g1468) & (g1479)) + ((!sk[103]) & (g8) & (!g32) & (g75) & (!g1468) & (!g1479)) + ((!sk[103]) & (g8) & (!g32) & (g75) & (!g1468) & (g1479)) + ((!sk[103]) & (g8) & (!g32) & (g75) & (g1468) & (!g1479)) + ((!sk[103]) & (g8) & (!g32) & (g75) & (g1468) & (g1479)) + ((!sk[103]) & (g8) & (g32) & (!g75) & (!g1468) & (!g1479)) + ((!sk[103]) & (g8) & (g32) & (!g75) & (!g1468) & (g1479)) + ((!sk[103]) & (g8) & (g32) & (!g75) & (g1468) & (!g1479)) + ((!sk[103]) & (g8) & (g32) & (!g75) & (g1468) & (g1479)) + ((!sk[103]) & (g8) & (g32) & (g75) & (!g1468) & (!g1479)) + ((!sk[103]) & (g8) & (g32) & (g75) & (!g1468) & (g1479)) + ((!sk[103]) & (g8) & (g32) & (g75) & (g1468) & (!g1479)) + ((!sk[103]) & (g8) & (g32) & (g75) & (g1468) & (g1479)) + ((sk[103]) & (!g8) & (!g32) & (!g75) & (!g1468) & (g1479)) + ((sk[103]) & (!g8) & (!g32) & (!g75) & (g1468) & (!g1479)) + ((sk[103]) & (!g8) & (!g32) & (!g75) & (g1468) & (g1479)) + ((sk[103]) & (!g8) & (!g32) & (g75) & (!g1468) & (!g1479)) + ((sk[103]) & (!g8) & (!g32) & (g75) & (!g1468) & (g1479)) + ((sk[103]) & (!g8) & (!g32) & (g75) & (g1468) & (!g1479)) + ((sk[103]) & (!g8) & (!g32) & (g75) & (g1468) & (g1479)) + ((sk[103]) & (!g8) & (g32) & (!g75) & (!g1468) & (!g1479)) + ((sk[103]) & (!g8) & (g32) & (!g75) & (!g1468) & (g1479)) + ((sk[103]) & (!g8) & (g32) & (!g75) & (g1468) & (!g1479)) + ((sk[103]) & (!g8) & (g32) & (!g75) & (g1468) & (g1479)) + ((sk[103]) & (!g8) & (g32) & (g75) & (!g1468) & (!g1479)) + ((sk[103]) & (!g8) & (g32) & (g75) & (!g1468) & (g1479)) + ((sk[103]) & (!g8) & (g32) & (g75) & (g1468) & (!g1479)) + ((sk[103]) & (!g8) & (g32) & (g75) & (g1468) & (g1479)));
	assign g1494 = (((!i_3_) & (!i_4_) & (!sk[104]) & (!g34) & (!g29) & (g1493)) + ((!i_3_) & (!i_4_) & (!sk[104]) & (!g34) & (g29) & (g1493)) + ((!i_3_) & (!i_4_) & (!sk[104]) & (g34) & (!g29) & (g1493)) + ((!i_3_) & (!i_4_) & (!sk[104]) & (g34) & (g29) & (g1493)) + ((!i_3_) & (!i_4_) & (sk[104]) & (!g34) & (!g29) & (!g1493)) + ((!i_3_) & (!i_4_) & (sk[104]) & (!g34) & (g29) & (!g1493)) + ((!i_3_) & (!i_4_) & (sk[104]) & (g34) & (!g29) & (!g1493)) + ((!i_3_) & (!i_4_) & (sk[104]) & (g34) & (g29) & (!g1493)) + ((!i_3_) & (i_4_) & (!sk[104]) & (!g34) & (!g29) & (g1493)) + ((!i_3_) & (i_4_) & (!sk[104]) & (!g34) & (g29) & (g1493)) + ((!i_3_) & (i_4_) & (!sk[104]) & (g34) & (!g29) & (g1493)) + ((!i_3_) & (i_4_) & (!sk[104]) & (g34) & (g29) & (g1493)) + ((!i_3_) & (i_4_) & (sk[104]) & (!g34) & (!g29) & (!g1493)) + ((!i_3_) & (i_4_) & (sk[104]) & (!g34) & (g29) & (!g1493)) + ((!i_3_) & (i_4_) & (sk[104]) & (g34) & (!g29) & (!g1493)) + ((i_3_) & (!i_4_) & (!sk[104]) & (!g34) & (!g29) & (!g1493)) + ((i_3_) & (!i_4_) & (!sk[104]) & (!g34) & (!g29) & (g1493)) + ((i_3_) & (!i_4_) & (!sk[104]) & (!g34) & (g29) & (!g1493)) + ((i_3_) & (!i_4_) & (!sk[104]) & (!g34) & (g29) & (g1493)) + ((i_3_) & (!i_4_) & (!sk[104]) & (g34) & (!g29) & (!g1493)) + ((i_3_) & (!i_4_) & (!sk[104]) & (g34) & (!g29) & (g1493)) + ((i_3_) & (!i_4_) & (!sk[104]) & (g34) & (g29) & (!g1493)) + ((i_3_) & (!i_4_) & (!sk[104]) & (g34) & (g29) & (g1493)) + ((i_3_) & (!i_4_) & (sk[104]) & (!g34) & (!g29) & (!g1493)) + ((i_3_) & (!i_4_) & (sk[104]) & (!g34) & (g29) & (!g1493)) + ((i_3_) & (!i_4_) & (sk[104]) & (g34) & (!g29) & (!g1493)) + ((i_3_) & (!i_4_) & (sk[104]) & (g34) & (g29) & (!g1493)) + ((i_3_) & (i_4_) & (!sk[104]) & (!g34) & (!g29) & (!g1493)) + ((i_3_) & (i_4_) & (!sk[104]) & (!g34) & (!g29) & (g1493)) + ((i_3_) & (i_4_) & (!sk[104]) & (!g34) & (g29) & (!g1493)) + ((i_3_) & (i_4_) & (!sk[104]) & (!g34) & (g29) & (g1493)) + ((i_3_) & (i_4_) & (!sk[104]) & (g34) & (!g29) & (!g1493)) + ((i_3_) & (i_4_) & (!sk[104]) & (g34) & (!g29) & (g1493)) + ((i_3_) & (i_4_) & (!sk[104]) & (g34) & (g29) & (!g1493)) + ((i_3_) & (i_4_) & (!sk[104]) & (g34) & (g29) & (g1493)) + ((i_3_) & (i_4_) & (sk[104]) & (!g34) & (!g29) & (!g1493)) + ((i_3_) & (i_4_) & (sk[104]) & (!g34) & (g29) & (!g1493)) + ((i_3_) & (i_4_) & (sk[104]) & (g34) & (!g29) & (!g1493)) + ((i_3_) & (i_4_) & (sk[104]) & (g34) & (g29) & (!g1493)));
	assign g1495 = (((!g10) & (!g78) & (!g1480) & (!g1492) & (!sk[105]) & (g1494)) + ((!g10) & (!g78) & (!g1480) & (!g1492) & (sk[105]) & (g1494)) + ((!g10) & (!g78) & (!g1480) & (g1492) & (!sk[105]) & (g1494)) + ((!g10) & (!g78) & (g1480) & (!g1492) & (!sk[105]) & (g1494)) + ((!g10) & (!g78) & (g1480) & (!g1492) & (sk[105]) & (g1494)) + ((!g10) & (!g78) & (g1480) & (g1492) & (!sk[105]) & (g1494)) + ((!g10) & (g78) & (!g1480) & (!g1492) & (!sk[105]) & (g1494)) + ((!g10) & (g78) & (!g1480) & (!g1492) & (sk[105]) & (g1494)) + ((!g10) & (g78) & (!g1480) & (g1492) & (!sk[105]) & (g1494)) + ((!g10) & (g78) & (g1480) & (!g1492) & (!sk[105]) & (g1494)) + ((!g10) & (g78) & (g1480) & (!g1492) & (sk[105]) & (g1494)) + ((!g10) & (g78) & (g1480) & (g1492) & (!sk[105]) & (g1494)) + ((g10) & (!g78) & (!g1480) & (!g1492) & (!sk[105]) & (!g1494)) + ((g10) & (!g78) & (!g1480) & (!g1492) & (!sk[105]) & (g1494)) + ((g10) & (!g78) & (!g1480) & (g1492) & (!sk[105]) & (!g1494)) + ((g10) & (!g78) & (!g1480) & (g1492) & (!sk[105]) & (g1494)) + ((g10) & (!g78) & (g1480) & (!g1492) & (!sk[105]) & (!g1494)) + ((g10) & (!g78) & (g1480) & (!g1492) & (!sk[105]) & (g1494)) + ((g10) & (!g78) & (g1480) & (!g1492) & (sk[105]) & (g1494)) + ((g10) & (!g78) & (g1480) & (g1492) & (!sk[105]) & (!g1494)) + ((g10) & (!g78) & (g1480) & (g1492) & (!sk[105]) & (g1494)) + ((g10) & (g78) & (!g1480) & (!g1492) & (!sk[105]) & (!g1494)) + ((g10) & (g78) & (!g1480) & (!g1492) & (!sk[105]) & (g1494)) + ((g10) & (g78) & (!g1480) & (g1492) & (!sk[105]) & (!g1494)) + ((g10) & (g78) & (!g1480) & (g1492) & (!sk[105]) & (g1494)) + ((g10) & (g78) & (g1480) & (!g1492) & (!sk[105]) & (!g1494)) + ((g10) & (g78) & (g1480) & (!g1492) & (!sk[105]) & (g1494)) + ((g10) & (g78) & (g1480) & (g1492) & (!sk[105]) & (!g1494)) + ((g10) & (g78) & (g1480) & (g1492) & (!sk[105]) & (g1494)));
	assign g1496 = (((!i_5_) & (!i_3_) & (!sk[106]) & (i_4_) & (g29)) + ((!i_5_) & (!i_3_) & (sk[106]) & (!i_4_) & (g29)) + ((!i_5_) & (i_3_) & (!sk[106]) & (!i_4_) & (!g29)) + ((!i_5_) & (i_3_) & (!sk[106]) & (!i_4_) & (g29)) + ((!i_5_) & (i_3_) & (!sk[106]) & (i_4_) & (!g29)) + ((!i_5_) & (i_3_) & (!sk[106]) & (i_4_) & (g29)) + ((i_5_) & (!i_3_) & (!sk[106]) & (i_4_) & (!g29)) + ((i_5_) & (!i_3_) & (!sk[106]) & (i_4_) & (g29)) + ((i_5_) & (!i_3_) & (sk[106]) & (!i_4_) & (g29)) + ((i_5_) & (!i_3_) & (sk[106]) & (i_4_) & (g29)) + ((i_5_) & (i_3_) & (!sk[106]) & (!i_4_) & (!g29)) + ((i_5_) & (i_3_) & (!sk[106]) & (!i_4_) & (g29)) + ((i_5_) & (i_3_) & (!sk[106]) & (i_4_) & (!g29)) + ((i_5_) & (i_3_) & (!sk[106]) & (i_4_) & (g29)));
	assign g1497 = (((!g14) & (!g4) & (!sk[107]) & (g78) & (g1496)) + ((!g14) & (g4) & (!sk[107]) & (!g78) & (!g1496)) + ((!g14) & (g4) & (!sk[107]) & (!g78) & (g1496)) + ((!g14) & (g4) & (!sk[107]) & (g78) & (!g1496)) + ((!g14) & (g4) & (!sk[107]) & (g78) & (g1496)) + ((!g14) & (g4) & (sk[107]) & (!g78) & (g1496)) + ((!g14) & (g4) & (sk[107]) & (g78) & (g1496)) + ((g14) & (!g4) & (!sk[107]) & (g78) & (!g1496)) + ((g14) & (!g4) & (!sk[107]) & (g78) & (g1496)) + ((g14) & (!g4) & (sk[107]) & (g78) & (!g1496)) + ((g14) & (!g4) & (sk[107]) & (g78) & (g1496)) + ((g14) & (g4) & (!sk[107]) & (!g78) & (!g1496)) + ((g14) & (g4) & (!sk[107]) & (!g78) & (g1496)) + ((g14) & (g4) & (!sk[107]) & (g78) & (!g1496)) + ((g14) & (g4) & (!sk[107]) & (g78) & (g1496)) + ((g14) & (g4) & (sk[107]) & (!g78) & (g1496)) + ((g14) & (g4) & (sk[107]) & (g78) & (!g1496)) + ((g14) & (g4) & (sk[107]) & (g78) & (g1496)));
	assign g1498 = (((!g8) & (!sk[108]) & (!g34) & (g1487) & (g78)) + ((!g8) & (!sk[108]) & (g34) & (!g1487) & (!g78)) + ((!g8) & (!sk[108]) & (g34) & (!g1487) & (g78)) + ((!g8) & (!sk[108]) & (g34) & (g1487) & (!g78)) + ((!g8) & (!sk[108]) & (g34) & (g1487) & (g78)) + ((!g8) & (sk[108]) & (!g34) & (!g1487) & (g78)) + ((!g8) & (sk[108]) & (!g34) & (g1487) & (g78)) + ((!g8) & (sk[108]) & (g34) & (!g1487) & (g78)) + ((!g8) & (sk[108]) & (g34) & (g1487) & (!g78)) + ((!g8) & (sk[108]) & (g34) & (g1487) & (g78)) + ((g8) & (!sk[108]) & (!g34) & (g1487) & (!g78)) + ((g8) & (!sk[108]) & (!g34) & (g1487) & (g78)) + ((g8) & (!sk[108]) & (g34) & (!g1487) & (!g78)) + ((g8) & (!sk[108]) & (g34) & (!g1487) & (g78)) + ((g8) & (!sk[108]) & (g34) & (g1487) & (!g78)) + ((g8) & (!sk[108]) & (g34) & (g1487) & (g78)) + ((g8) & (sk[108]) & (g34) & (g1487) & (!g78)) + ((g8) & (sk[108]) & (g34) & (g1487) & (g78)));
	assign g1499 = (((!g30) & (!g1441) & (!g1488) & (!g1497) & (!sk[109]) & (g1498)) + ((!g30) & (!g1441) & (!g1488) & (!g1497) & (sk[109]) & (!g1498)) + ((!g30) & (!g1441) & (!g1488) & (g1497) & (!sk[109]) & (g1498)) + ((!g30) & (!g1441) & (g1488) & (!g1497) & (!sk[109]) & (g1498)) + ((!g30) & (!g1441) & (g1488) & (g1497) & (!sk[109]) & (g1498)) + ((!g30) & (g1441) & (!g1488) & (!g1497) & (!sk[109]) & (g1498)) + ((!g30) & (g1441) & (!g1488) & (g1497) & (!sk[109]) & (g1498)) + ((!g30) & (g1441) & (g1488) & (!g1497) & (!sk[109]) & (g1498)) + ((!g30) & (g1441) & (g1488) & (g1497) & (!sk[109]) & (g1498)) + ((g30) & (!g1441) & (!g1488) & (!g1497) & (!sk[109]) & (!g1498)) + ((g30) & (!g1441) & (!g1488) & (!g1497) & (!sk[109]) & (g1498)) + ((g30) & (!g1441) & (!g1488) & (!g1497) & (sk[109]) & (!g1498)) + ((g30) & (!g1441) & (!g1488) & (g1497) & (!sk[109]) & (!g1498)) + ((g30) & (!g1441) & (!g1488) & (g1497) & (!sk[109]) & (g1498)) + ((g30) & (!g1441) & (g1488) & (!g1497) & (!sk[109]) & (!g1498)) + ((g30) & (!g1441) & (g1488) & (!g1497) & (!sk[109]) & (g1498)) + ((g30) & (!g1441) & (g1488) & (g1497) & (!sk[109]) & (!g1498)) + ((g30) & (!g1441) & (g1488) & (g1497) & (!sk[109]) & (g1498)) + ((g30) & (g1441) & (!g1488) & (!g1497) & (!sk[109]) & (!g1498)) + ((g30) & (g1441) & (!g1488) & (!g1497) & (!sk[109]) & (g1498)) + ((g30) & (g1441) & (!g1488) & (!g1497) & (sk[109]) & (!g1498)) + ((g30) & (g1441) & (!g1488) & (g1497) & (!sk[109]) & (!g1498)) + ((g30) & (g1441) & (!g1488) & (g1497) & (!sk[109]) & (g1498)) + ((g30) & (g1441) & (g1488) & (!g1497) & (!sk[109]) & (!g1498)) + ((g30) & (g1441) & (g1488) & (!g1497) & (!sk[109]) & (g1498)) + ((g30) & (g1441) & (g1488) & (g1497) & (!sk[109]) & (!g1498)) + ((g30) & (g1441) & (g1488) & (g1497) & (!sk[109]) & (g1498)));
	assign o_29_ = (((!i_9_) & (!i_10_) & (!g63) & (g73) & (!g1495) & (!g1499)) + ((!i_9_) & (!i_10_) & (!g63) & (g73) & (!g1495) & (g1499)) + ((!i_9_) & (!i_10_) & (!g63) & (g73) & (g1495) & (!g1499)) + ((!i_9_) & (!i_10_) & (g63) & (g73) & (!g1495) & (!g1499)) + ((!i_9_) & (!i_10_) & (g63) & (g73) & (!g1495) & (g1499)) + ((!i_9_) & (!i_10_) & (g63) & (g73) & (g1495) & (!g1499)) + ((!i_9_) & (i_10_) & (!g63) & (g73) & (!g1495) & (!g1499)) + ((!i_9_) & (i_10_) & (!g63) & (g73) & (!g1495) & (g1499)) + ((!i_9_) & (i_10_) & (!g63) & (g73) & (g1495) & (!g1499)) + ((!i_9_) & (i_10_) & (g63) & (g73) & (!g1495) & (!g1499)) + ((!i_9_) & (i_10_) & (g63) & (g73) & (!g1495) & (g1499)) + ((!i_9_) & (i_10_) & (g63) & (g73) & (g1495) & (!g1499)) + ((i_9_) & (!i_10_) & (!g63) & (g73) & (!g1495) & (!g1499)) + ((i_9_) & (!i_10_) & (!g63) & (g73) & (!g1495) & (g1499)) + ((i_9_) & (!i_10_) & (!g63) & (g73) & (g1495) & (!g1499)) + ((i_9_) & (!i_10_) & (g63) & (g73) & (!g1495) & (!g1499)) + ((i_9_) & (!i_10_) & (g63) & (g73) & (!g1495) & (g1499)) + ((i_9_) & (!i_10_) & (g63) & (g73) & (g1495) & (!g1499)) + ((i_9_) & (!i_10_) & (g63) & (g73) & (g1495) & (g1499)) + ((i_9_) & (i_10_) & (!g63) & (g73) & (!g1495) & (!g1499)) + ((i_9_) & (i_10_) & (!g63) & (g73) & (!g1495) & (g1499)) + ((i_9_) & (i_10_) & (!g63) & (g73) & (g1495) & (!g1499)) + ((i_9_) & (i_10_) & (g63) & (g73) & (!g1495) & (!g1499)) + ((i_9_) & (i_10_) & (g63) & (g73) & (!g1495) & (g1499)) + ((i_9_) & (i_10_) & (g63) & (g73) & (g1495) & (!g1499)));
	assign g1501 = (((!g2) & (!i_6_) & (!sk[111]) & (!i_7_) & (!g40) & (g77)) + ((!g2) & (!i_6_) & (!sk[111]) & (!i_7_) & (g40) & (g77)) + ((!g2) & (!i_6_) & (!sk[111]) & (i_7_) & (!g40) & (g77)) + ((!g2) & (!i_6_) & (!sk[111]) & (i_7_) & (g40) & (g77)) + ((!g2) & (i_6_) & (!sk[111]) & (!i_7_) & (!g40) & (g77)) + ((!g2) & (i_6_) & (!sk[111]) & (!i_7_) & (g40) & (g77)) + ((!g2) & (i_6_) & (!sk[111]) & (i_7_) & (!g40) & (g77)) + ((!g2) & (i_6_) & (!sk[111]) & (i_7_) & (g40) & (g77)) + ((!g2) & (i_6_) & (sk[111]) & (i_7_) & (!g40) & (g77)) + ((!g2) & (i_6_) & (sk[111]) & (i_7_) & (g40) & (!g77)) + ((!g2) & (i_6_) & (sk[111]) & (i_7_) & (g40) & (g77)) + ((g2) & (!i_6_) & (!sk[111]) & (!i_7_) & (!g40) & (!g77)) + ((g2) & (!i_6_) & (!sk[111]) & (!i_7_) & (!g40) & (g77)) + ((g2) & (!i_6_) & (!sk[111]) & (!i_7_) & (g40) & (!g77)) + ((g2) & (!i_6_) & (!sk[111]) & (!i_7_) & (g40) & (g77)) + ((g2) & (!i_6_) & (!sk[111]) & (i_7_) & (!g40) & (!g77)) + ((g2) & (!i_6_) & (!sk[111]) & (i_7_) & (!g40) & (g77)) + ((g2) & (!i_6_) & (!sk[111]) & (i_7_) & (g40) & (!g77)) + ((g2) & (!i_6_) & (!sk[111]) & (i_7_) & (g40) & (g77)) + ((g2) & (!i_6_) & (sk[111]) & (i_7_) & (!g40) & (!g77)) + ((g2) & (!i_6_) & (sk[111]) & (i_7_) & (!g40) & (g77)) + ((g2) & (!i_6_) & (sk[111]) & (i_7_) & (g40) & (!g77)) + ((g2) & (!i_6_) & (sk[111]) & (i_7_) & (g40) & (g77)) + ((g2) & (i_6_) & (!sk[111]) & (!i_7_) & (!g40) & (!g77)) + ((g2) & (i_6_) & (!sk[111]) & (!i_7_) & (!g40) & (g77)) + ((g2) & (i_6_) & (!sk[111]) & (!i_7_) & (g40) & (!g77)) + ((g2) & (i_6_) & (!sk[111]) & (!i_7_) & (g40) & (g77)) + ((g2) & (i_6_) & (!sk[111]) & (i_7_) & (!g40) & (!g77)) + ((g2) & (i_6_) & (!sk[111]) & (i_7_) & (!g40) & (g77)) + ((g2) & (i_6_) & (!sk[111]) & (i_7_) & (g40) & (!g77)) + ((g2) & (i_6_) & (!sk[111]) & (i_7_) & (g40) & (g77)) + ((g2) & (i_6_) & (sk[111]) & (i_7_) & (!g40) & (!g77)) + ((g2) & (i_6_) & (sk[111]) & (i_7_) & (!g40) & (g77)) + ((g2) & (i_6_) & (sk[111]) & (i_7_) & (g40) & (!g77)) + ((g2) & (i_6_) & (sk[111]) & (i_7_) & (g40) & (g77)));
	assign g1502 = (((!i_3_) & (!sk[112]) & (!i_4_) & (g29) & (g1501)) + ((!i_3_) & (!sk[112]) & (i_4_) & (!g29) & (!g1501)) + ((!i_3_) & (!sk[112]) & (i_4_) & (!g29) & (g1501)) + ((!i_3_) & (!sk[112]) & (i_4_) & (g29) & (!g1501)) + ((!i_3_) & (!sk[112]) & (i_4_) & (g29) & (g1501)) + ((!i_3_) & (sk[112]) & (!i_4_) & (!g29) & (!g1501)) + ((!i_3_) & (sk[112]) & (i_4_) & (!g29) & (!g1501)) + ((!i_3_) & (sk[112]) & (i_4_) & (g29) & (!g1501)) + ((i_3_) & (!sk[112]) & (!i_4_) & (g29) & (!g1501)) + ((i_3_) & (!sk[112]) & (!i_4_) & (g29) & (g1501)) + ((i_3_) & (!sk[112]) & (i_4_) & (!g29) & (!g1501)) + ((i_3_) & (!sk[112]) & (i_4_) & (!g29) & (g1501)) + ((i_3_) & (!sk[112]) & (i_4_) & (g29) & (!g1501)) + ((i_3_) & (!sk[112]) & (i_4_) & (g29) & (g1501)) + ((i_3_) & (sk[112]) & (!i_4_) & (!g29) & (!g1501)) + ((i_3_) & (sk[112]) & (!i_4_) & (g29) & (!g1501)) + ((i_3_) & (sk[112]) & (i_4_) & (!g29) & (!g1501)) + ((i_3_) & (sk[112]) & (i_4_) & (g29) & (!g1501)));
	assign g1503 = (((!g73) & (!g81) & (!g1486) & (!g1495) & (!sk[113]) & (g1502)) + ((!g73) & (!g81) & (!g1486) & (!g1495) & (sk[113]) & (!g1502)) + ((!g73) & (!g81) & (!g1486) & (!g1495) & (sk[113]) & (g1502)) + ((!g73) & (!g81) & (!g1486) & (g1495) & (!sk[113]) & (g1502)) + ((!g73) & (!g81) & (!g1486) & (g1495) & (sk[113]) & (!g1502)) + ((!g73) & (!g81) & (!g1486) & (g1495) & (sk[113]) & (g1502)) + ((!g73) & (!g81) & (g1486) & (!g1495) & (!sk[113]) & (g1502)) + ((!g73) & (!g81) & (g1486) & (!g1495) & (sk[113]) & (!g1502)) + ((!g73) & (!g81) & (g1486) & (!g1495) & (sk[113]) & (g1502)) + ((!g73) & (!g81) & (g1486) & (g1495) & (!sk[113]) & (g1502)) + ((!g73) & (!g81) & (g1486) & (g1495) & (sk[113]) & (!g1502)) + ((!g73) & (!g81) & (g1486) & (g1495) & (sk[113]) & (g1502)) + ((!g73) & (g81) & (!g1486) & (!g1495) & (!sk[113]) & (g1502)) + ((!g73) & (g81) & (!g1486) & (!g1495) & (sk[113]) & (!g1502)) + ((!g73) & (g81) & (!g1486) & (!g1495) & (sk[113]) & (g1502)) + ((!g73) & (g81) & (!g1486) & (g1495) & (!sk[113]) & (g1502)) + ((!g73) & (g81) & (!g1486) & (g1495) & (sk[113]) & (!g1502)) + ((!g73) & (g81) & (!g1486) & (g1495) & (sk[113]) & (g1502)) + ((!g73) & (g81) & (g1486) & (!g1495) & (!sk[113]) & (g1502)) + ((!g73) & (g81) & (g1486) & (!g1495) & (sk[113]) & (!g1502)) + ((!g73) & (g81) & (g1486) & (!g1495) & (sk[113]) & (g1502)) + ((!g73) & (g81) & (g1486) & (g1495) & (!sk[113]) & (g1502)) + ((!g73) & (g81) & (g1486) & (g1495) & (sk[113]) & (!g1502)) + ((!g73) & (g81) & (g1486) & (g1495) & (sk[113]) & (g1502)) + ((g73) & (!g81) & (!g1486) & (!g1495) & (!sk[113]) & (!g1502)) + ((g73) & (!g81) & (!g1486) & (!g1495) & (!sk[113]) & (g1502)) + ((g73) & (!g81) & (!g1486) & (g1495) & (!sk[113]) & (!g1502)) + ((g73) & (!g81) & (!g1486) & (g1495) & (!sk[113]) & (g1502)) + ((g73) & (!g81) & (g1486) & (!g1495) & (!sk[113]) & (!g1502)) + ((g73) & (!g81) & (g1486) & (!g1495) & (!sk[113]) & (g1502)) + ((g73) & (!g81) & (g1486) & (g1495) & (!sk[113]) & (!g1502)) + ((g73) & (!g81) & (g1486) & (g1495) & (!sk[113]) & (g1502)) + ((g73) & (g81) & (!g1486) & (!g1495) & (!sk[113]) & (!g1502)) + ((g73) & (g81) & (!g1486) & (!g1495) & (!sk[113]) & (g1502)) + ((g73) & (g81) & (!g1486) & (g1495) & (!sk[113]) & (!g1502)) + ((g73) & (g81) & (!g1486) & (g1495) & (!sk[113]) & (g1502)) + ((g73) & (g81) & (g1486) & (!g1495) & (!sk[113]) & (!g1502)) + ((g73) & (g81) & (g1486) & (!g1495) & (!sk[113]) & (g1502)) + ((g73) & (g81) & (g1486) & (g1495) & (!sk[113]) & (!g1502)) + ((g73) & (g81) & (g1486) & (g1495) & (!sk[113]) & (g1502)) + ((g73) & (g81) & (g1486) & (g1495) & (sk[113]) & (g1502)));
	assign g1504 = (((!i_3_) & (!i_4_) & (!sk[114]) & (!g1) & (!g32) & (g27)) + ((!i_3_) & (!i_4_) & (!sk[114]) & (!g1) & (g32) & (g27)) + ((!i_3_) & (!i_4_) & (!sk[114]) & (g1) & (!g32) & (g27)) + ((!i_3_) & (!i_4_) & (!sk[114]) & (g1) & (g32) & (g27)) + ((!i_3_) & (!i_4_) & (sk[114]) & (!g1) & (!g32) & (!g27)) + ((!i_3_) & (!i_4_) & (sk[114]) & (!g1) & (!g32) & (g27)) + ((!i_3_) & (!i_4_) & (sk[114]) & (g1) & (!g32) & (!g27)) + ((!i_3_) & (i_4_) & (!sk[114]) & (!g1) & (!g32) & (g27)) + ((!i_3_) & (i_4_) & (!sk[114]) & (!g1) & (g32) & (g27)) + ((!i_3_) & (i_4_) & (!sk[114]) & (g1) & (!g32) & (g27)) + ((!i_3_) & (i_4_) & (!sk[114]) & (g1) & (g32) & (g27)) + ((!i_3_) & (i_4_) & (sk[114]) & (!g1) & (!g32) & (!g27)) + ((!i_3_) & (i_4_) & (sk[114]) & (!g1) & (!g32) & (g27)) + ((!i_3_) & (i_4_) & (sk[114]) & (g1) & (!g32) & (!g27)) + ((!i_3_) & (i_4_) & (sk[114]) & (g1) & (!g32) & (g27)) + ((i_3_) & (!i_4_) & (!sk[114]) & (!g1) & (!g32) & (!g27)) + ((i_3_) & (!i_4_) & (!sk[114]) & (!g1) & (!g32) & (g27)) + ((i_3_) & (!i_4_) & (!sk[114]) & (!g1) & (g32) & (!g27)) + ((i_3_) & (!i_4_) & (!sk[114]) & (!g1) & (g32) & (g27)) + ((i_3_) & (!i_4_) & (!sk[114]) & (g1) & (!g32) & (!g27)) + ((i_3_) & (!i_4_) & (!sk[114]) & (g1) & (!g32) & (g27)) + ((i_3_) & (!i_4_) & (!sk[114]) & (g1) & (g32) & (!g27)) + ((i_3_) & (!i_4_) & (!sk[114]) & (g1) & (g32) & (g27)) + ((i_3_) & (!i_4_) & (sk[114]) & (!g1) & (!g32) & (!g27)) + ((i_3_) & (!i_4_) & (sk[114]) & (!g1) & (!g32) & (g27)) + ((i_3_) & (!i_4_) & (sk[114]) & (g1) & (!g32) & (!g27)) + ((i_3_) & (!i_4_) & (sk[114]) & (g1) & (!g32) & (g27)) + ((i_3_) & (i_4_) & (!sk[114]) & (!g1) & (!g32) & (!g27)) + ((i_3_) & (i_4_) & (!sk[114]) & (!g1) & (!g32) & (g27)) + ((i_3_) & (i_4_) & (!sk[114]) & (!g1) & (g32) & (!g27)) + ((i_3_) & (i_4_) & (!sk[114]) & (!g1) & (g32) & (g27)) + ((i_3_) & (i_4_) & (!sk[114]) & (g1) & (!g32) & (!g27)) + ((i_3_) & (i_4_) & (!sk[114]) & (g1) & (!g32) & (g27)) + ((i_3_) & (i_4_) & (!sk[114]) & (g1) & (g32) & (!g27)) + ((i_3_) & (i_4_) & (!sk[114]) & (g1) & (g32) & (g27)) + ((i_3_) & (i_4_) & (sk[114]) & (!g1) & (!g32) & (!g27)) + ((i_3_) & (i_4_) & (sk[114]) & (!g1) & (!g32) & (g27)) + ((i_3_) & (i_4_) & (sk[114]) & (g1) & (!g32) & (!g27)) + ((i_3_) & (i_4_) & (sk[114]) & (g1) & (!g32) & (g27)));
	assign o_31_ = (((!i_9_) & (!i_10_) & (!g63) & (!g1488) & (!sk[115]) & (g1504)) + ((!i_9_) & (!i_10_) & (!g63) & (!g1488) & (sk[115]) & (!g1504)) + ((!i_9_) & (!i_10_) & (!g63) & (g1488) & (!sk[115]) & (g1504)) + ((!i_9_) & (!i_10_) & (!g63) & (g1488) & (sk[115]) & (!g1504)) + ((!i_9_) & (!i_10_) & (!g63) & (g1488) & (sk[115]) & (g1504)) + ((!i_9_) & (!i_10_) & (g63) & (!g1488) & (!sk[115]) & (g1504)) + ((!i_9_) & (!i_10_) & (g63) & (!g1488) & (sk[115]) & (!g1504)) + ((!i_9_) & (!i_10_) & (g63) & (g1488) & (!sk[115]) & (g1504)) + ((!i_9_) & (!i_10_) & (g63) & (g1488) & (sk[115]) & (!g1504)) + ((!i_9_) & (!i_10_) & (g63) & (g1488) & (sk[115]) & (g1504)) + ((!i_9_) & (i_10_) & (!g63) & (!g1488) & (!sk[115]) & (g1504)) + ((!i_9_) & (i_10_) & (!g63) & (g1488) & (!sk[115]) & (g1504)) + ((!i_9_) & (i_10_) & (!g63) & (g1488) & (sk[115]) & (!g1504)) + ((!i_9_) & (i_10_) & (!g63) & (g1488) & (sk[115]) & (g1504)) + ((!i_9_) & (i_10_) & (g63) & (!g1488) & (!sk[115]) & (g1504)) + ((!i_9_) & (i_10_) & (g63) & (!g1488) & (sk[115]) & (!g1504)) + ((!i_9_) & (i_10_) & (g63) & (!g1488) & (sk[115]) & (g1504)) + ((!i_9_) & (i_10_) & (g63) & (g1488) & (!sk[115]) & (g1504)) + ((!i_9_) & (i_10_) & (g63) & (g1488) & (sk[115]) & (!g1504)) + ((!i_9_) & (i_10_) & (g63) & (g1488) & (sk[115]) & (g1504)) + ((i_9_) & (!i_10_) & (!g63) & (!g1488) & (!sk[115]) & (!g1504)) + ((i_9_) & (!i_10_) & (!g63) & (!g1488) & (!sk[115]) & (g1504)) + ((i_9_) & (!i_10_) & (!g63) & (g1488) & (!sk[115]) & (!g1504)) + ((i_9_) & (!i_10_) & (!g63) & (g1488) & (!sk[115]) & (g1504)) + ((i_9_) & (!i_10_) & (!g63) & (g1488) & (sk[115]) & (!g1504)) + ((i_9_) & (!i_10_) & (!g63) & (g1488) & (sk[115]) & (g1504)) + ((i_9_) & (!i_10_) & (g63) & (!g1488) & (!sk[115]) & (!g1504)) + ((i_9_) & (!i_10_) & (g63) & (!g1488) & (!sk[115]) & (g1504)) + ((i_9_) & (!i_10_) & (g63) & (!g1488) & (sk[115]) & (!g1504)) + ((i_9_) & (!i_10_) & (g63) & (!g1488) & (sk[115]) & (g1504)) + ((i_9_) & (!i_10_) & (g63) & (g1488) & (!sk[115]) & (!g1504)) + ((i_9_) & (!i_10_) & (g63) & (g1488) & (!sk[115]) & (g1504)) + ((i_9_) & (!i_10_) & (g63) & (g1488) & (sk[115]) & (!g1504)) + ((i_9_) & (!i_10_) & (g63) & (g1488) & (sk[115]) & (g1504)) + ((i_9_) & (i_10_) & (!g63) & (!g1488) & (!sk[115]) & (!g1504)) + ((i_9_) & (i_10_) & (!g63) & (!g1488) & (!sk[115]) & (g1504)) + ((i_9_) & (i_10_) & (!g63) & (g1488) & (!sk[115]) & (!g1504)) + ((i_9_) & (i_10_) & (!g63) & (g1488) & (!sk[115]) & (g1504)) + ((i_9_) & (i_10_) & (!g63) & (g1488) & (sk[115]) & (!g1504)) + ((i_9_) & (i_10_) & (!g63) & (g1488) & (sk[115]) & (g1504)) + ((i_9_) & (i_10_) & (g63) & (!g1488) & (!sk[115]) & (!g1504)) + ((i_9_) & (i_10_) & (g63) & (!g1488) & (!sk[115]) & (g1504)) + ((i_9_) & (i_10_) & (g63) & (g1488) & (!sk[115]) & (!g1504)) + ((i_9_) & (i_10_) & (g63) & (g1488) & (!sk[115]) & (g1504)) + ((i_9_) & (i_10_) & (g63) & (g1488) & (sk[115]) & (!g1504)) + ((i_9_) & (i_10_) & (g63) & (g1488) & (sk[115]) & (g1504)));
	assign g1506 = (((!i_5_) & (!i_3_) & (!i_4_) & (!g1) & (!i_6_) & (!i_7_)) + ((!i_5_) & (!i_3_) & (!i_4_) & (!g1) & (!i_6_) & (i_7_)) + ((!i_5_) & (!i_3_) & (!i_4_) & (!g1) & (i_6_) & (!i_7_)) + ((!i_5_) & (!i_3_) & (!i_4_) & (!g1) & (i_6_) & (i_7_)) + ((!i_5_) & (!i_3_) & (!i_4_) & (g1) & (!i_6_) & (!i_7_)) + ((!i_5_) & (!i_3_) & (!i_4_) & (g1) & (i_6_) & (!i_7_)) + ((!i_5_) & (!i_3_) & (i_4_) & (!g1) & (!i_6_) & (!i_7_)) + ((!i_5_) & (!i_3_) & (i_4_) & (!g1) & (!i_6_) & (i_7_)) + ((!i_5_) & (!i_3_) & (i_4_) & (!g1) & (i_6_) & (!i_7_)) + ((!i_5_) & (!i_3_) & (i_4_) & (!g1) & (i_6_) & (i_7_)) + ((!i_5_) & (!i_3_) & (i_4_) & (g1) & (!i_6_) & (!i_7_)) + ((!i_5_) & (!i_3_) & (i_4_) & (g1) & (i_6_) & (!i_7_)) + ((!i_5_) & (i_3_) & (!i_4_) & (!g1) & (!i_6_) & (!i_7_)) + ((!i_5_) & (i_3_) & (!i_4_) & (!g1) & (!i_6_) & (i_7_)) + ((!i_5_) & (i_3_) & (!i_4_) & (!g1) & (i_6_) & (!i_7_)) + ((!i_5_) & (i_3_) & (!i_4_) & (!g1) & (i_6_) & (i_7_)) + ((!i_5_) & (i_3_) & (!i_4_) & (g1) & (!i_6_) & (!i_7_)) + ((!i_5_) & (i_3_) & (!i_4_) & (g1) & (!i_6_) & (i_7_)) + ((!i_5_) & (i_3_) & (!i_4_) & (g1) & (i_6_) & (!i_7_)) + ((!i_5_) & (i_3_) & (!i_4_) & (g1) & (i_6_) & (i_7_)) + ((!i_5_) & (i_3_) & (i_4_) & (!g1) & (!i_6_) & (!i_7_)) + ((!i_5_) & (i_3_) & (i_4_) & (!g1) & (!i_6_) & (i_7_)) + ((!i_5_) & (i_3_) & (i_4_) & (!g1) & (i_6_) & (!i_7_)) + ((!i_5_) & (i_3_) & (i_4_) & (!g1) & (i_6_) & (i_7_)) + ((!i_5_) & (i_3_) & (i_4_) & (g1) & (!i_6_) & (!i_7_)) + ((!i_5_) & (i_3_) & (i_4_) & (g1) & (!i_6_) & (i_7_)) + ((!i_5_) & (i_3_) & (i_4_) & (g1) & (i_6_) & (!i_7_)) + ((i_5_) & (!i_3_) & (!i_4_) & (!g1) & (!i_6_) & (!i_7_)) + ((i_5_) & (!i_3_) & (!i_4_) & (!g1) & (!i_6_) & (i_7_)) + ((i_5_) & (!i_3_) & (!i_4_) & (!g1) & (i_6_) & (!i_7_)) + ((i_5_) & (!i_3_) & (!i_4_) & (!g1) & (i_6_) & (i_7_)) + ((i_5_) & (!i_3_) & (!i_4_) & (g1) & (!i_6_) & (!i_7_)) + ((i_5_) & (!i_3_) & (!i_4_) & (g1) & (!i_6_) & (i_7_)) + ((i_5_) & (!i_3_) & (!i_4_) & (g1) & (i_6_) & (!i_7_)) + ((i_5_) & (!i_3_) & (!i_4_) & (g1) & (i_6_) & (i_7_)) + ((i_5_) & (!i_3_) & (i_4_) & (!g1) & (!i_6_) & (!i_7_)) + ((i_5_) & (!i_3_) & (i_4_) & (!g1) & (!i_6_) & (i_7_)) + ((i_5_) & (!i_3_) & (i_4_) & (!g1) & (i_6_) & (!i_7_)) + ((i_5_) & (!i_3_) & (i_4_) & (!g1) & (i_6_) & (i_7_)) + ((i_5_) & (!i_3_) & (i_4_) & (g1) & (!i_6_) & (!i_7_)) + ((i_5_) & (!i_3_) & (i_4_) & (g1) & (!i_6_) & (i_7_)) + ((i_5_) & (!i_3_) & (i_4_) & (g1) & (i_6_) & (!i_7_)) + ((i_5_) & (!i_3_) & (i_4_) & (g1) & (i_6_) & (i_7_)) + ((i_5_) & (i_3_) & (!i_4_) & (!g1) & (!i_6_) & (!i_7_)) + ((i_5_) & (i_3_) & (!i_4_) & (!g1) & (!i_6_) & (i_7_)) + ((i_5_) & (i_3_) & (!i_4_) & (!g1) & (i_6_) & (!i_7_)) + ((i_5_) & (i_3_) & (!i_4_) & (!g1) & (i_6_) & (i_7_)) + ((i_5_) & (i_3_) & (!i_4_) & (g1) & (!i_6_) & (!i_7_)) + ((i_5_) & (i_3_) & (!i_4_) & (g1) & (!i_6_) & (i_7_)) + ((i_5_) & (i_3_) & (!i_4_) & (g1) & (i_6_) & (!i_7_)) + ((i_5_) & (i_3_) & (!i_4_) & (g1) & (i_6_) & (i_7_)) + ((i_5_) & (i_3_) & (i_4_) & (!g1) & (!i_6_) & (!i_7_)) + ((i_5_) & (i_3_) & (i_4_) & (!g1) & (!i_6_) & (i_7_)) + ((i_5_) & (i_3_) & (i_4_) & (!g1) & (i_6_) & (!i_7_)) + ((i_5_) & (i_3_) & (i_4_) & (!g1) & (i_6_) & (i_7_)) + ((i_5_) & (i_3_) & (i_4_) & (g1) & (!i_6_) & (i_7_)) + ((i_5_) & (i_3_) & (i_4_) & (g1) & (i_6_) & (!i_7_)));
	assign g1507 = (((!g19) & (!g5) & (!g41) & (!sk[117]) & (!g78) & (g1479)) + ((!g19) & (!g5) & (!g41) & (!sk[117]) & (g78) & (g1479)) + ((!g19) & (!g5) & (g41) & (!sk[117]) & (!g78) & (g1479)) + ((!g19) & (!g5) & (g41) & (!sk[117]) & (g78) & (g1479)) + ((!g19) & (g5) & (!g41) & (!sk[117]) & (!g78) & (g1479)) + ((!g19) & (g5) & (!g41) & (!sk[117]) & (g78) & (g1479)) + ((!g19) & (g5) & (g41) & (!sk[117]) & (!g78) & (g1479)) + ((!g19) & (g5) & (g41) & (!sk[117]) & (g78) & (g1479)) + ((!g19) & (g5) & (g41) & (sk[117]) & (!g78) & (!g1479)) + ((!g19) & (g5) & (g41) & (sk[117]) & (!g78) & (g1479)) + ((!g19) & (g5) & (g41) & (sk[117]) & (g78) & (!g1479)) + ((!g19) & (g5) & (g41) & (sk[117]) & (g78) & (g1479)) + ((g19) & (!g5) & (!g41) & (!sk[117]) & (!g78) & (!g1479)) + ((g19) & (!g5) & (!g41) & (!sk[117]) & (!g78) & (g1479)) + ((g19) & (!g5) & (!g41) & (!sk[117]) & (g78) & (!g1479)) + ((g19) & (!g5) & (!g41) & (!sk[117]) & (g78) & (g1479)) + ((g19) & (!g5) & (!g41) & (sk[117]) & (!g78) & (g1479)) + ((g19) & (!g5) & (!g41) & (sk[117]) & (g78) & (!g1479)) + ((g19) & (!g5) & (!g41) & (sk[117]) & (g78) & (g1479)) + ((g19) & (!g5) & (g41) & (!sk[117]) & (!g78) & (!g1479)) + ((g19) & (!g5) & (g41) & (!sk[117]) & (!g78) & (g1479)) + ((g19) & (!g5) & (g41) & (!sk[117]) & (g78) & (!g1479)) + ((g19) & (!g5) & (g41) & (!sk[117]) & (g78) & (g1479)) + ((g19) & (!g5) & (g41) & (sk[117]) & (!g78) & (g1479)) + ((g19) & (!g5) & (g41) & (sk[117]) & (g78) & (!g1479)) + ((g19) & (!g5) & (g41) & (sk[117]) & (g78) & (g1479)) + ((g19) & (g5) & (!g41) & (!sk[117]) & (!g78) & (!g1479)) + ((g19) & (g5) & (!g41) & (!sk[117]) & (!g78) & (g1479)) + ((g19) & (g5) & (!g41) & (!sk[117]) & (g78) & (!g1479)) + ((g19) & (g5) & (!g41) & (!sk[117]) & (g78) & (g1479)) + ((g19) & (g5) & (g41) & (!sk[117]) & (!g78) & (!g1479)) + ((g19) & (g5) & (g41) & (!sk[117]) & (!g78) & (g1479)) + ((g19) & (g5) & (g41) & (!sk[117]) & (g78) & (!g1479)) + ((g19) & (g5) & (g41) & (!sk[117]) & (g78) & (g1479)) + ((g19) & (g5) & (g41) & (sk[117]) & (!g78) & (!g1479)) + ((g19) & (g5) & (g41) & (sk[117]) & (!g78) & (g1479)) + ((g19) & (g5) & (g41) & (sk[117]) & (g78) & (!g1479)) + ((g19) & (g5) & (g41) & (sk[117]) & (g78) & (g1479)));
	assign g1508 = (((!g30) & (!sk[118]) & (!g23) & (!g1487) & (!g1464) & (g1498)) + ((!g30) & (!sk[118]) & (!g23) & (!g1487) & (g1464) & (g1498)) + ((!g30) & (!sk[118]) & (!g23) & (g1487) & (!g1464) & (g1498)) + ((!g30) & (!sk[118]) & (!g23) & (g1487) & (g1464) & (g1498)) + ((!g30) & (!sk[118]) & (g23) & (!g1487) & (!g1464) & (g1498)) + ((!g30) & (!sk[118]) & (g23) & (!g1487) & (g1464) & (g1498)) + ((!g30) & (!sk[118]) & (g23) & (g1487) & (!g1464) & (g1498)) + ((!g30) & (!sk[118]) & (g23) & (g1487) & (g1464) & (g1498)) + ((!g30) & (sk[118]) & (!g23) & (!g1487) & (!g1464) & (!g1498)) + ((!g30) & (sk[118]) & (!g23) & (!g1487) & (g1464) & (!g1498)) + ((!g30) & (sk[118]) & (!g23) & (g1487) & (!g1464) & (!g1498)) + ((!g30) & (sk[118]) & (!g23) & (g1487) & (g1464) & (!g1498)) + ((!g30) & (sk[118]) & (g23) & (!g1487) & (g1464) & (!g1498)) + ((!g30) & (sk[118]) & (g23) & (g1487) & (g1464) & (!g1498)) + ((g30) & (!sk[118]) & (!g23) & (!g1487) & (!g1464) & (!g1498)) + ((g30) & (!sk[118]) & (!g23) & (!g1487) & (!g1464) & (g1498)) + ((g30) & (!sk[118]) & (!g23) & (!g1487) & (g1464) & (!g1498)) + ((g30) & (!sk[118]) & (!g23) & (!g1487) & (g1464) & (g1498)) + ((g30) & (!sk[118]) & (!g23) & (g1487) & (!g1464) & (!g1498)) + ((g30) & (!sk[118]) & (!g23) & (g1487) & (!g1464) & (g1498)) + ((g30) & (!sk[118]) & (!g23) & (g1487) & (g1464) & (!g1498)) + ((g30) & (!sk[118]) & (!g23) & (g1487) & (g1464) & (g1498)) + ((g30) & (!sk[118]) & (g23) & (!g1487) & (!g1464) & (!g1498)) + ((g30) & (!sk[118]) & (g23) & (!g1487) & (!g1464) & (g1498)) + ((g30) & (!sk[118]) & (g23) & (!g1487) & (g1464) & (!g1498)) + ((g30) & (!sk[118]) & (g23) & (!g1487) & (g1464) & (g1498)) + ((g30) & (!sk[118]) & (g23) & (g1487) & (!g1464) & (!g1498)) + ((g30) & (!sk[118]) & (g23) & (g1487) & (!g1464) & (g1498)) + ((g30) & (!sk[118]) & (g23) & (g1487) & (g1464) & (!g1498)) + ((g30) & (!sk[118]) & (g23) & (g1487) & (g1464) & (g1498)) + ((g30) & (sk[118]) & (!g23) & (!g1487) & (!g1464) & (!g1498)) + ((g30) & (sk[118]) & (!g23) & (!g1487) & (g1464) & (!g1498)) + ((g30) & (sk[118]) & (g23) & (!g1487) & (g1464) & (!g1498)));
	assign g1509 = (((!g73) & (!g1484) & (!sk[119]) & (!g1494) & (!g1507) & (g1508)) + ((!g73) & (!g1484) & (!sk[119]) & (!g1494) & (g1507) & (g1508)) + ((!g73) & (!g1484) & (!sk[119]) & (g1494) & (!g1507) & (g1508)) + ((!g73) & (!g1484) & (!sk[119]) & (g1494) & (g1507) & (g1508)) + ((!g73) & (!g1484) & (sk[119]) & (!g1494) & (!g1507) & (!g1508)) + ((!g73) & (!g1484) & (sk[119]) & (!g1494) & (!g1507) & (g1508)) + ((!g73) & (!g1484) & (sk[119]) & (!g1494) & (g1507) & (!g1508)) + ((!g73) & (!g1484) & (sk[119]) & (!g1494) & (g1507) & (g1508)) + ((!g73) & (!g1484) & (sk[119]) & (g1494) & (!g1507) & (!g1508)) + ((!g73) & (!g1484) & (sk[119]) & (g1494) & (!g1507) & (g1508)) + ((!g73) & (!g1484) & (sk[119]) & (g1494) & (g1507) & (!g1508)) + ((!g73) & (!g1484) & (sk[119]) & (g1494) & (g1507) & (g1508)) + ((!g73) & (g1484) & (!sk[119]) & (!g1494) & (!g1507) & (g1508)) + ((!g73) & (g1484) & (!sk[119]) & (!g1494) & (g1507) & (g1508)) + ((!g73) & (g1484) & (!sk[119]) & (g1494) & (!g1507) & (g1508)) + ((!g73) & (g1484) & (!sk[119]) & (g1494) & (g1507) & (g1508)) + ((!g73) & (g1484) & (sk[119]) & (!g1494) & (!g1507) & (!g1508)) + ((!g73) & (g1484) & (sk[119]) & (!g1494) & (!g1507) & (g1508)) + ((!g73) & (g1484) & (sk[119]) & (!g1494) & (g1507) & (!g1508)) + ((!g73) & (g1484) & (sk[119]) & (!g1494) & (g1507) & (g1508)) + ((!g73) & (g1484) & (sk[119]) & (g1494) & (!g1507) & (!g1508)) + ((!g73) & (g1484) & (sk[119]) & (g1494) & (!g1507) & (g1508)) + ((!g73) & (g1484) & (sk[119]) & (g1494) & (g1507) & (!g1508)) + ((!g73) & (g1484) & (sk[119]) & (g1494) & (g1507) & (g1508)) + ((g73) & (!g1484) & (!sk[119]) & (!g1494) & (!g1507) & (!g1508)) + ((g73) & (!g1484) & (!sk[119]) & (!g1494) & (!g1507) & (g1508)) + ((g73) & (!g1484) & (!sk[119]) & (!g1494) & (g1507) & (!g1508)) + ((g73) & (!g1484) & (!sk[119]) & (!g1494) & (g1507) & (g1508)) + ((g73) & (!g1484) & (!sk[119]) & (g1494) & (!g1507) & (!g1508)) + ((g73) & (!g1484) & (!sk[119]) & (g1494) & (!g1507) & (g1508)) + ((g73) & (!g1484) & (!sk[119]) & (g1494) & (g1507) & (!g1508)) + ((g73) & (!g1484) & (!sk[119]) & (g1494) & (g1507) & (g1508)) + ((g73) & (g1484) & (!sk[119]) & (!g1494) & (!g1507) & (!g1508)) + ((g73) & (g1484) & (!sk[119]) & (!g1494) & (!g1507) & (g1508)) + ((g73) & (g1484) & (!sk[119]) & (!g1494) & (g1507) & (!g1508)) + ((g73) & (g1484) & (!sk[119]) & (!g1494) & (g1507) & (g1508)) + ((g73) & (g1484) & (!sk[119]) & (g1494) & (!g1507) & (!g1508)) + ((g73) & (g1484) & (!sk[119]) & (g1494) & (!g1507) & (g1508)) + ((g73) & (g1484) & (!sk[119]) & (g1494) & (g1507) & (!g1508)) + ((g73) & (g1484) & (!sk[119]) & (g1494) & (g1507) & (g1508)) + ((g73) & (g1484) & (sk[119]) & (g1494) & (!g1507) & (g1508)));
	assign g1510 = (((!g976) & (!g994) & (!sk[120]) & (g1460) & (g1463)) + ((!g976) & (g994) & (!sk[120]) & (!g1460) & (!g1463)) + ((!g976) & (g994) & (!sk[120]) & (!g1460) & (g1463)) + ((!g976) & (g994) & (!sk[120]) & (g1460) & (!g1463)) + ((!g976) & (g994) & (!sk[120]) & (g1460) & (g1463)) + ((g976) & (!g994) & (!sk[120]) & (g1460) & (!g1463)) + ((g976) & (!g994) & (!sk[120]) & (g1460) & (g1463)) + ((g976) & (g994) & (!sk[120]) & (!g1460) & (!g1463)) + ((g976) & (g994) & (!sk[120]) & (!g1460) & (g1463)) + ((g976) & (g994) & (!sk[120]) & (g1460) & (!g1463)) + ((g976) & (g994) & (!sk[120]) & (g1460) & (g1463)) + ((g976) & (g994) & (sk[120]) & (g1460) & (g1463)));
	assign g1511 = (((!g931) & (sk[121]) & (!g1266) & (g1268)) + ((g931) & (!sk[121]) & (!g1266) & (!g1268)) + ((g931) & (!sk[121]) & (!g1266) & (g1268)) + ((g931) & (!sk[121]) & (g1266) & (!g1268)) + ((g931) & (!sk[121]) & (g1266) & (g1268)));
	assign g1512 = (((!g1278) & (!g1279) & (!sk[122]) & (!g1281) & (!g1282) & (g1492)) + ((!g1278) & (!g1279) & (!sk[122]) & (!g1281) & (g1282) & (g1492)) + ((!g1278) & (!g1279) & (!sk[122]) & (g1281) & (!g1282) & (g1492)) + ((!g1278) & (!g1279) & (!sk[122]) & (g1281) & (g1282) & (g1492)) + ((!g1278) & (g1279) & (!sk[122]) & (!g1281) & (!g1282) & (g1492)) + ((!g1278) & (g1279) & (!sk[122]) & (!g1281) & (g1282) & (g1492)) + ((!g1278) & (g1279) & (!sk[122]) & (g1281) & (!g1282) & (g1492)) + ((!g1278) & (g1279) & (!sk[122]) & (g1281) & (g1282) & (g1492)) + ((g1278) & (!g1279) & (!sk[122]) & (!g1281) & (!g1282) & (!g1492)) + ((g1278) & (!g1279) & (!sk[122]) & (!g1281) & (!g1282) & (g1492)) + ((g1278) & (!g1279) & (!sk[122]) & (!g1281) & (g1282) & (!g1492)) + ((g1278) & (!g1279) & (!sk[122]) & (!g1281) & (g1282) & (g1492)) + ((g1278) & (!g1279) & (!sk[122]) & (g1281) & (!g1282) & (!g1492)) + ((g1278) & (!g1279) & (!sk[122]) & (g1281) & (!g1282) & (g1492)) + ((g1278) & (!g1279) & (!sk[122]) & (g1281) & (g1282) & (!g1492)) + ((g1278) & (!g1279) & (!sk[122]) & (g1281) & (g1282) & (g1492)) + ((g1278) & (!g1279) & (sk[122]) & (g1281) & (!g1282) & (!g1492)) + ((g1278) & (g1279) & (!sk[122]) & (!g1281) & (!g1282) & (!g1492)) + ((g1278) & (g1279) & (!sk[122]) & (!g1281) & (!g1282) & (g1492)) + ((g1278) & (g1279) & (!sk[122]) & (!g1281) & (g1282) & (!g1492)) + ((g1278) & (g1279) & (!sk[122]) & (!g1281) & (g1282) & (g1492)) + ((g1278) & (g1279) & (!sk[122]) & (g1281) & (!g1282) & (!g1492)) + ((g1278) & (g1279) & (!sk[122]) & (g1281) & (!g1282) & (g1492)) + ((g1278) & (g1279) & (!sk[122]) & (g1281) & (g1282) & (!g1492)) + ((g1278) & (g1279) & (!sk[122]) & (g1281) & (g1282) & (g1492)));
	assign g1513 = (((!i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (!sk[123]) & (g13)) + ((!i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (!sk[123]) & (g13)) + ((!i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (!sk[123]) & (g13)) + ((!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!sk[123]) & (g13)) + ((!i_11_) & (!i_9_) & (i_10_) & (i_15_) & (sk[123]) & (g13)) + ((!i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (!sk[123]) & (g13)) + ((!i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!sk[123]) & (g13)) + ((!i_11_) & (i_9_) & (i_10_) & (!i_15_) & (!sk[123]) & (g13)) + ((!i_11_) & (i_9_) & (i_10_) & (i_15_) & (!sk[123]) & (g13)) + ((i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (!sk[123]) & (!g13)) + ((i_11_) & (!i_9_) & (!i_10_) & (!i_15_) & (!sk[123]) & (g13)) + ((i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (!sk[123]) & (!g13)) + ((i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (!sk[123]) & (g13)) + ((i_11_) & (!i_9_) & (!i_10_) & (i_15_) & (sk[123]) & (g13)) + ((i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (!sk[123]) & (!g13)) + ((i_11_) & (!i_9_) & (i_10_) & (!i_15_) & (!sk[123]) & (g13)) + ((i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!sk[123]) & (!g13)) + ((i_11_) & (!i_9_) & (i_10_) & (i_15_) & (!sk[123]) & (g13)) + ((i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (!sk[123]) & (!g13)) + ((i_11_) & (i_9_) & (!i_10_) & (!i_15_) & (!sk[123]) & (g13)) + ((i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!sk[123]) & (!g13)) + ((i_11_) & (i_9_) & (!i_10_) & (i_15_) & (!sk[123]) & (g13)) + ((i_11_) & (i_9_) & (i_10_) & (!i_15_) & (!sk[123]) & (!g13)) + ((i_11_) & (i_9_) & (i_10_) & (!i_15_) & (!sk[123]) & (g13)) + ((i_11_) & (i_9_) & (i_10_) & (i_15_) & (!sk[123]) & (!g13)) + ((i_11_) & (i_9_) & (i_10_) & (i_15_) & (!sk[123]) & (g13)));
	assign g1514 = (((!g101) & (!g109) & (!g641) & (!g676) & (!g903) & (!g1513)) + ((!g101) & (!g109) & (!g641) & (!g676) & (!g903) & (g1513)) + ((!g101) & (!g109) & (!g641) & (!g676) & (g903) & (!g1513)) + ((!g101) & (!g109) & (!g641) & (!g676) & (g903) & (g1513)) + ((!g101) & (!g109) & (!g641) & (g676) & (!g903) & (!g1513)) + ((!g101) & (!g109) & (!g641) & (g676) & (!g903) & (g1513)) + ((!g101) & (!g109) & (!g641) & (g676) & (g903) & (!g1513)) + ((!g101) & (!g109) & (!g641) & (g676) & (g903) & (g1513)) + ((!g101) & (!g109) & (g641) & (!g676) & (!g903) & (!g1513)) + ((!g101) & (!g109) & (g641) & (!g676) & (!g903) & (g1513)) + ((!g101) & (!g109) & (g641) & (!g676) & (g903) & (!g1513)) + ((!g101) & (!g109) & (g641) & (!g676) & (g903) & (g1513)) + ((!g101) & (!g109) & (g641) & (g676) & (!g903) & (!g1513)) + ((!g101) & (!g109) & (g641) & (g676) & (!g903) & (g1513)) + ((!g101) & (!g109) & (g641) & (g676) & (g903) & (!g1513)) + ((!g101) & (!g109) & (g641) & (g676) & (g903) & (g1513)) + ((!g101) & (g109) & (!g641) & (!g676) & (!g903) & (!g1513)) + ((!g101) & (g109) & (!g641) & (!g676) & (g903) & (!g1513)) + ((!g101) & (g109) & (!g641) & (g676) & (!g903) & (!g1513)) + ((!g101) & (g109) & (!g641) & (g676) & (g903) & (!g1513)) + ((g101) & (!g109) & (!g641) & (!g676) & (!g903) & (!g1513)) + ((g101) & (!g109) & (!g641) & (!g676) & (!g903) & (g1513)) + ((g101) & (!g109) & (g641) & (!g676) & (!g903) & (!g1513)) + ((g101) & (!g109) & (g641) & (!g676) & (!g903) & (g1513)) + ((g101) & (g109) & (!g641) & (!g676) & (!g903) & (!g1513)));
	assign g1515 = (((!sk[125]) & (!i_14_) & (!i_12_) & (!i_8_) & (!g102) & (g108)) + ((!sk[125]) & (!i_14_) & (!i_12_) & (!i_8_) & (g102) & (g108)) + ((!sk[125]) & (!i_14_) & (!i_12_) & (i_8_) & (!g102) & (g108)) + ((!sk[125]) & (!i_14_) & (!i_12_) & (i_8_) & (g102) & (g108)) + ((!sk[125]) & (!i_14_) & (i_12_) & (!i_8_) & (!g102) & (g108)) + ((!sk[125]) & (!i_14_) & (i_12_) & (!i_8_) & (g102) & (g108)) + ((!sk[125]) & (!i_14_) & (i_12_) & (i_8_) & (!g102) & (g108)) + ((!sk[125]) & (!i_14_) & (i_12_) & (i_8_) & (g102) & (g108)) + ((!sk[125]) & (i_14_) & (!i_12_) & (!i_8_) & (!g102) & (!g108)) + ((!sk[125]) & (i_14_) & (!i_12_) & (!i_8_) & (!g102) & (g108)) + ((!sk[125]) & (i_14_) & (!i_12_) & (!i_8_) & (g102) & (!g108)) + ((!sk[125]) & (i_14_) & (!i_12_) & (!i_8_) & (g102) & (g108)) + ((!sk[125]) & (i_14_) & (!i_12_) & (i_8_) & (!g102) & (!g108)) + ((!sk[125]) & (i_14_) & (!i_12_) & (i_8_) & (!g102) & (g108)) + ((!sk[125]) & (i_14_) & (!i_12_) & (i_8_) & (g102) & (!g108)) + ((!sk[125]) & (i_14_) & (!i_12_) & (i_8_) & (g102) & (g108)) + ((!sk[125]) & (i_14_) & (i_12_) & (!i_8_) & (!g102) & (!g108)) + ((!sk[125]) & (i_14_) & (i_12_) & (!i_8_) & (!g102) & (g108)) + ((!sk[125]) & (i_14_) & (i_12_) & (!i_8_) & (g102) & (!g108)) + ((!sk[125]) & (i_14_) & (i_12_) & (!i_8_) & (g102) & (g108)) + ((!sk[125]) & (i_14_) & (i_12_) & (i_8_) & (!g102) & (!g108)) + ((!sk[125]) & (i_14_) & (i_12_) & (i_8_) & (!g102) & (g108)) + ((!sk[125]) & (i_14_) & (i_12_) & (i_8_) & (g102) & (!g108)) + ((!sk[125]) & (i_14_) & (i_12_) & (i_8_) & (g102) & (g108)) + ((sk[125]) & (i_14_) & (!i_12_) & (i_8_) & (!g102) & (g108)));
	assign g1516 = (((!g20) & (!sk[126]) & (!g78) & (!g1479) & (!g1482) & (g1515)) + ((!g20) & (!sk[126]) & (!g78) & (!g1479) & (g1482) & (g1515)) + ((!g20) & (!sk[126]) & (!g78) & (g1479) & (!g1482) & (g1515)) + ((!g20) & (!sk[126]) & (!g78) & (g1479) & (g1482) & (g1515)) + ((!g20) & (!sk[126]) & (g78) & (!g1479) & (!g1482) & (g1515)) + ((!g20) & (!sk[126]) & (g78) & (!g1479) & (g1482) & (g1515)) + ((!g20) & (!sk[126]) & (g78) & (g1479) & (!g1482) & (g1515)) + ((!g20) & (!sk[126]) & (g78) & (g1479) & (g1482) & (g1515)) + ((!g20) & (sk[126]) & (!g78) & (!g1479) & (g1482) & (!g1515)) + ((g20) & (!sk[126]) & (!g78) & (!g1479) & (!g1482) & (!g1515)) + ((g20) & (!sk[126]) & (!g78) & (!g1479) & (!g1482) & (g1515)) + ((g20) & (!sk[126]) & (!g78) & (!g1479) & (g1482) & (!g1515)) + ((g20) & (!sk[126]) & (!g78) & (!g1479) & (g1482) & (g1515)) + ((g20) & (!sk[126]) & (!g78) & (g1479) & (!g1482) & (!g1515)) + ((g20) & (!sk[126]) & (!g78) & (g1479) & (!g1482) & (g1515)) + ((g20) & (!sk[126]) & (!g78) & (g1479) & (g1482) & (!g1515)) + ((g20) & (!sk[126]) & (!g78) & (g1479) & (g1482) & (g1515)) + ((g20) & (!sk[126]) & (g78) & (!g1479) & (!g1482) & (!g1515)) + ((g20) & (!sk[126]) & (g78) & (!g1479) & (!g1482) & (g1515)) + ((g20) & (!sk[126]) & (g78) & (!g1479) & (g1482) & (!g1515)) + ((g20) & (!sk[126]) & (g78) & (!g1479) & (g1482) & (g1515)) + ((g20) & (!sk[126]) & (g78) & (g1479) & (!g1482) & (!g1515)) + ((g20) & (!sk[126]) & (g78) & (g1479) & (!g1482) & (g1515)) + ((g20) & (!sk[126]) & (g78) & (g1479) & (g1482) & (!g1515)) + ((g20) & (!sk[126]) & (g78) & (g1479) & (g1482) & (g1515)) + ((g20) & (sk[126]) & (!g78) & (!g1479) & (g1482) & (!g1515)) + ((g20) & (sk[126]) & (!g78) & (g1479) & (g1482) & (!g1515)) + ((g20) & (sk[126]) & (g78) & (!g1479) & (g1482) & (!g1515)) + ((g20) & (sk[126]) & (g78) & (g1479) & (g1482) & (!g1515)));
	assign g1517 = (((!i_3_) & (!i_4_) & (!g1) & (!g5) & (!sk[127]) & (g27)) + ((!i_3_) & (!i_4_) & (!g1) & (g5) & (!sk[127]) & (g27)) + ((!i_3_) & (!i_4_) & (g1) & (!g5) & (!sk[127]) & (g27)) + ((!i_3_) & (!i_4_) & (g1) & (g5) & (!sk[127]) & (g27)) + ((!i_3_) & (i_4_) & (!g1) & (!g5) & (!sk[127]) & (g27)) + ((!i_3_) & (i_4_) & (!g1) & (g5) & (!sk[127]) & (g27)) + ((!i_3_) & (i_4_) & (g1) & (!g5) & (!sk[127]) & (g27)) + ((!i_3_) & (i_4_) & (g1) & (g5) & (!sk[127]) & (g27)) + ((!i_3_) & (i_4_) & (g1) & (g5) & (sk[127]) & (g27)) + ((i_3_) & (!i_4_) & (!g1) & (!g5) & (!sk[127]) & (!g27)) + ((i_3_) & (!i_4_) & (!g1) & (!g5) & (!sk[127]) & (g27)) + ((i_3_) & (!i_4_) & (!g1) & (g5) & (!sk[127]) & (!g27)) + ((i_3_) & (!i_4_) & (!g1) & (g5) & (!sk[127]) & (g27)) + ((i_3_) & (!i_4_) & (g1) & (!g5) & (!sk[127]) & (!g27)) + ((i_3_) & (!i_4_) & (g1) & (!g5) & (!sk[127]) & (g27)) + ((i_3_) & (!i_4_) & (g1) & (g5) & (!sk[127]) & (!g27)) + ((i_3_) & (!i_4_) & (g1) & (g5) & (!sk[127]) & (g27)) + ((i_3_) & (i_4_) & (!g1) & (!g5) & (!sk[127]) & (!g27)) + ((i_3_) & (i_4_) & (!g1) & (!g5) & (!sk[127]) & (g27)) + ((i_3_) & (i_4_) & (!g1) & (g5) & (!sk[127]) & (!g27)) + ((i_3_) & (i_4_) & (!g1) & (g5) & (!sk[127]) & (g27)) + ((i_3_) & (i_4_) & (g1) & (!g5) & (!sk[127]) & (!g27)) + ((i_3_) & (i_4_) & (g1) & (!g5) & (!sk[127]) & (g27)) + ((i_3_) & (i_4_) & (g1) & (g5) & (!sk[127]) & (!g27)) + ((i_3_) & (i_4_) & (g1) & (g5) & (!sk[127]) & (g27)));
	assign g1518 = (((!i_6_) & (!i_7_) & (!g1487) & (sk[0]) & (!g1517)) + ((!i_6_) & (!i_7_) & (g1487) & (!sk[0]) & (g1517)) + ((!i_6_) & (!i_7_) & (g1487) & (sk[0]) & (!g1517)) + ((!i_6_) & (i_7_) & (!g1487) & (!sk[0]) & (!g1517)) + ((!i_6_) & (i_7_) & (!g1487) & (!sk[0]) & (g1517)) + ((!i_6_) & (i_7_) & (!g1487) & (sk[0]) & (!g1517)) + ((!i_6_) & (i_7_) & (g1487) & (!sk[0]) & (!g1517)) + ((!i_6_) & (i_7_) & (g1487) & (!sk[0]) & (g1517)) + ((!i_6_) & (i_7_) & (g1487) & (sk[0]) & (!g1517)) + ((i_6_) & (!i_7_) & (!g1487) & (sk[0]) & (!g1517)) + ((i_6_) & (!i_7_) & (g1487) & (!sk[0]) & (!g1517)) + ((i_6_) & (!i_7_) & (g1487) & (!sk[0]) & (g1517)) + ((i_6_) & (i_7_) & (!g1487) & (!sk[0]) & (!g1517)) + ((i_6_) & (i_7_) & (!g1487) & (!sk[0]) & (g1517)) + ((i_6_) & (i_7_) & (!g1487) & (sk[0]) & (!g1517)) + ((i_6_) & (i_7_) & (g1487) & (!sk[0]) & (!g1517)) + ((i_6_) & (i_7_) & (g1487) & (!sk[0]) & (g1517)) + ((i_6_) & (i_7_) & (g1487) & (sk[0]) & (!g1517)));
	assign g1519 = (((i_8_) & (!g10) & (!g100) & (g108) & (!g640) & (!g677)) + ((i_8_) & (!g10) & (!g100) & (g108) & (!g640) & (g677)) + ((i_8_) & (!g10) & (g100) & (!g108) & (!g640) & (g677)) + ((i_8_) & (!g10) & (g100) & (!g108) & (g640) & (g677)) + ((i_8_) & (!g10) & (g100) & (g108) & (!g640) & (!g677)) + ((i_8_) & (!g10) & (g100) & (g108) & (!g640) & (g677)) + ((i_8_) & (!g10) & (g100) & (g108) & (g640) & (g677)) + ((i_8_) & (g10) & (!g100) & (g108) & (!g640) & (!g677)) + ((i_8_) & (g10) & (!g100) & (g108) & (!g640) & (g677)) + ((i_8_) & (g10) & (g100) & (!g108) & (!g640) & (!g677)) + ((i_8_) & (g10) & (g100) & (!g108) & (!g640) & (g677)) + ((i_8_) & (g10) & (g100) & (!g108) & (g640) & (!g677)) + ((i_8_) & (g10) & (g100) & (!g108) & (g640) & (g677)) + ((i_8_) & (g10) & (g100) & (g108) & (!g640) & (!g677)) + ((i_8_) & (g10) & (g100) & (g108) & (!g640) & (g677)) + ((i_8_) & (g10) & (g100) & (g108) & (g640) & (!g677)) + ((i_8_) & (g10) & (g100) & (g108) & (g640) & (g677)));
	assign g1520 = (((!sk[2]) & (!g101) & (!g848) & (!g1497) & (!g1518) & (g1519)) + ((!sk[2]) & (!g101) & (!g848) & (!g1497) & (g1518) & (g1519)) + ((!sk[2]) & (!g101) & (!g848) & (g1497) & (!g1518) & (g1519)) + ((!sk[2]) & (!g101) & (!g848) & (g1497) & (g1518) & (g1519)) + ((!sk[2]) & (!g101) & (g848) & (!g1497) & (!g1518) & (g1519)) + ((!sk[2]) & (!g101) & (g848) & (!g1497) & (g1518) & (g1519)) + ((!sk[2]) & (!g101) & (g848) & (g1497) & (!g1518) & (g1519)) + ((!sk[2]) & (!g101) & (g848) & (g1497) & (g1518) & (g1519)) + ((!sk[2]) & (g101) & (!g848) & (!g1497) & (!g1518) & (!g1519)) + ((!sk[2]) & (g101) & (!g848) & (!g1497) & (!g1518) & (g1519)) + ((!sk[2]) & (g101) & (!g848) & (!g1497) & (g1518) & (!g1519)) + ((!sk[2]) & (g101) & (!g848) & (!g1497) & (g1518) & (g1519)) + ((!sk[2]) & (g101) & (!g848) & (g1497) & (!g1518) & (!g1519)) + ((!sk[2]) & (g101) & (!g848) & (g1497) & (!g1518) & (g1519)) + ((!sk[2]) & (g101) & (!g848) & (g1497) & (g1518) & (!g1519)) + ((!sk[2]) & (g101) & (!g848) & (g1497) & (g1518) & (g1519)) + ((!sk[2]) & (g101) & (g848) & (!g1497) & (!g1518) & (!g1519)) + ((!sk[2]) & (g101) & (g848) & (!g1497) & (!g1518) & (g1519)) + ((!sk[2]) & (g101) & (g848) & (!g1497) & (g1518) & (!g1519)) + ((!sk[2]) & (g101) & (g848) & (!g1497) & (g1518) & (g1519)) + ((!sk[2]) & (g101) & (g848) & (g1497) & (!g1518) & (!g1519)) + ((!sk[2]) & (g101) & (g848) & (g1497) & (!g1518) & (g1519)) + ((!sk[2]) & (g101) & (g848) & (g1497) & (g1518) & (!g1519)) + ((!sk[2]) & (g101) & (g848) & (g1497) & (g1518) & (g1519)) + ((sk[2]) & (!g101) & (!g848) & (!g1497) & (g1518) & (!g1519)) + ((sk[2]) & (!g101) & (g848) & (!g1497) & (g1518) & (!g1519)) + ((sk[2]) & (g101) & (g848) & (!g1497) & (g1518) & (!g1519)));
	assign g1521 = (((!sk[3]) & (!g1589) & (!g1380) & (!g1514) & (!g1516) & (g1520)) + ((!sk[3]) & (!g1589) & (!g1380) & (!g1514) & (g1516) & (g1520)) + ((!sk[3]) & (!g1589) & (!g1380) & (g1514) & (!g1516) & (g1520)) + ((!sk[3]) & (!g1589) & (!g1380) & (g1514) & (g1516) & (g1520)) + ((!sk[3]) & (!g1589) & (g1380) & (!g1514) & (!g1516) & (g1520)) + ((!sk[3]) & (!g1589) & (g1380) & (!g1514) & (g1516) & (g1520)) + ((!sk[3]) & (!g1589) & (g1380) & (g1514) & (!g1516) & (g1520)) + ((!sk[3]) & (!g1589) & (g1380) & (g1514) & (g1516) & (g1520)) + ((!sk[3]) & (g1589) & (!g1380) & (!g1514) & (!g1516) & (!g1520)) + ((!sk[3]) & (g1589) & (!g1380) & (!g1514) & (!g1516) & (g1520)) + ((!sk[3]) & (g1589) & (!g1380) & (!g1514) & (g1516) & (!g1520)) + ((!sk[3]) & (g1589) & (!g1380) & (!g1514) & (g1516) & (g1520)) + ((!sk[3]) & (g1589) & (!g1380) & (g1514) & (!g1516) & (!g1520)) + ((!sk[3]) & (g1589) & (!g1380) & (g1514) & (!g1516) & (g1520)) + ((!sk[3]) & (g1589) & (!g1380) & (g1514) & (g1516) & (!g1520)) + ((!sk[3]) & (g1589) & (!g1380) & (g1514) & (g1516) & (g1520)) + ((!sk[3]) & (g1589) & (g1380) & (!g1514) & (!g1516) & (!g1520)) + ((!sk[3]) & (g1589) & (g1380) & (!g1514) & (!g1516) & (g1520)) + ((!sk[3]) & (g1589) & (g1380) & (!g1514) & (g1516) & (!g1520)) + ((!sk[3]) & (g1589) & (g1380) & (!g1514) & (g1516) & (g1520)) + ((!sk[3]) & (g1589) & (g1380) & (g1514) & (!g1516) & (!g1520)) + ((!sk[3]) & (g1589) & (g1380) & (g1514) & (!g1516) & (g1520)) + ((!sk[3]) & (g1589) & (g1380) & (g1514) & (g1516) & (!g1520)) + ((!sk[3]) & (g1589) & (g1380) & (g1514) & (g1516) & (g1520)) + ((sk[3]) & (g1589) & (!g1380) & (g1514) & (g1516) & (g1520)));
	assign g1522 = (((!g1511) & (!g1321) & (!g1402) & (!sk[4]) & (!g1512) & (g1521)) + ((!g1511) & (!g1321) & (!g1402) & (!sk[4]) & (g1512) & (g1521)) + ((!g1511) & (!g1321) & (g1402) & (!sk[4]) & (!g1512) & (g1521)) + ((!g1511) & (!g1321) & (g1402) & (!sk[4]) & (g1512) & (g1521)) + ((!g1511) & (g1321) & (!g1402) & (!sk[4]) & (!g1512) & (g1521)) + ((!g1511) & (g1321) & (!g1402) & (!sk[4]) & (g1512) & (g1521)) + ((!g1511) & (g1321) & (g1402) & (!sk[4]) & (!g1512) & (g1521)) + ((!g1511) & (g1321) & (g1402) & (!sk[4]) & (g1512) & (g1521)) + ((g1511) & (!g1321) & (!g1402) & (!sk[4]) & (!g1512) & (!g1521)) + ((g1511) & (!g1321) & (!g1402) & (!sk[4]) & (!g1512) & (g1521)) + ((g1511) & (!g1321) & (!g1402) & (!sk[4]) & (g1512) & (!g1521)) + ((g1511) & (!g1321) & (!g1402) & (!sk[4]) & (g1512) & (g1521)) + ((g1511) & (!g1321) & (g1402) & (!sk[4]) & (!g1512) & (!g1521)) + ((g1511) & (!g1321) & (g1402) & (!sk[4]) & (!g1512) & (g1521)) + ((g1511) & (!g1321) & (g1402) & (!sk[4]) & (g1512) & (!g1521)) + ((g1511) & (!g1321) & (g1402) & (!sk[4]) & (g1512) & (g1521)) + ((g1511) & (g1321) & (!g1402) & (!sk[4]) & (!g1512) & (!g1521)) + ((g1511) & (g1321) & (!g1402) & (!sk[4]) & (!g1512) & (g1521)) + ((g1511) & (g1321) & (!g1402) & (!sk[4]) & (g1512) & (!g1521)) + ((g1511) & (g1321) & (!g1402) & (!sk[4]) & (g1512) & (g1521)) + ((g1511) & (g1321) & (g1402) & (!sk[4]) & (!g1512) & (!g1521)) + ((g1511) & (g1321) & (g1402) & (!sk[4]) & (!g1512) & (g1521)) + ((g1511) & (g1321) & (g1402) & (!sk[4]) & (g1512) & (!g1521)) + ((g1511) & (g1321) & (g1402) & (!sk[4]) & (g1512) & (g1521)) + ((g1511) & (g1321) & (g1402) & (sk[4]) & (g1512) & (g1521)));
	assign o_34_ = (((!g73) & (!sk[5]) & (!g1195) & (!g1453) & (!g1510) & (g1522)) + ((!g73) & (!sk[5]) & (!g1195) & (!g1453) & (g1510) & (g1522)) + ((!g73) & (!sk[5]) & (!g1195) & (g1453) & (!g1510) & (g1522)) + ((!g73) & (!sk[5]) & (!g1195) & (g1453) & (g1510) & (g1522)) + ((!g73) & (!sk[5]) & (g1195) & (!g1453) & (!g1510) & (g1522)) + ((!g73) & (!sk[5]) & (g1195) & (!g1453) & (g1510) & (g1522)) + ((!g73) & (!sk[5]) & (g1195) & (g1453) & (!g1510) & (g1522)) + ((!g73) & (!sk[5]) & (g1195) & (g1453) & (g1510) & (g1522)) + ((g73) & (!sk[5]) & (!g1195) & (!g1453) & (!g1510) & (!g1522)) + ((g73) & (!sk[5]) & (!g1195) & (!g1453) & (!g1510) & (g1522)) + ((g73) & (!sk[5]) & (!g1195) & (!g1453) & (g1510) & (!g1522)) + ((g73) & (!sk[5]) & (!g1195) & (!g1453) & (g1510) & (g1522)) + ((g73) & (!sk[5]) & (!g1195) & (g1453) & (!g1510) & (!g1522)) + ((g73) & (!sk[5]) & (!g1195) & (g1453) & (!g1510) & (g1522)) + ((g73) & (!sk[5]) & (!g1195) & (g1453) & (g1510) & (!g1522)) + ((g73) & (!sk[5]) & (!g1195) & (g1453) & (g1510) & (g1522)) + ((g73) & (!sk[5]) & (g1195) & (!g1453) & (!g1510) & (!g1522)) + ((g73) & (!sk[5]) & (g1195) & (!g1453) & (!g1510) & (g1522)) + ((g73) & (!sk[5]) & (g1195) & (!g1453) & (g1510) & (!g1522)) + ((g73) & (!sk[5]) & (g1195) & (!g1453) & (g1510) & (g1522)) + ((g73) & (!sk[5]) & (g1195) & (g1453) & (!g1510) & (!g1522)) + ((g73) & (!sk[5]) & (g1195) & (g1453) & (!g1510) & (g1522)) + ((g73) & (!sk[5]) & (g1195) & (g1453) & (g1510) & (!g1522)) + ((g73) & (!sk[5]) & (g1195) & (g1453) & (g1510) & (g1522)) + ((g73) & (sk[5]) & (!g1195) & (!g1453) & (!g1510) & (!g1522)) + ((g73) & (sk[5]) & (!g1195) & (!g1453) & (!g1510) & (g1522)) + ((g73) & (sk[5]) & (!g1195) & (!g1453) & (g1510) & (!g1522)) + ((g73) & (sk[5]) & (!g1195) & (!g1453) & (g1510) & (g1522)) + ((g73) & (sk[5]) & (!g1195) & (g1453) & (!g1510) & (!g1522)) + ((g73) & (sk[5]) & (!g1195) & (g1453) & (!g1510) & (g1522)) + ((g73) & (sk[5]) & (!g1195) & (g1453) & (g1510) & (!g1522)) + ((g73) & (sk[5]) & (!g1195) & (g1453) & (g1510) & (g1522)) + ((g73) & (sk[5]) & (g1195) & (!g1453) & (!g1510) & (!g1522)) + ((g73) & (sk[5]) & (g1195) & (!g1453) & (!g1510) & (g1522)) + ((g73) & (sk[5]) & (g1195) & (!g1453) & (g1510) & (!g1522)) + ((g73) & (sk[5]) & (g1195) & (!g1453) & (g1510) & (g1522)) + ((g73) & (sk[5]) & (g1195) & (g1453) & (!g1510) & (!g1522)) + ((g73) & (sk[5]) & (g1195) & (g1453) & (!g1510) & (g1522)) + ((g73) & (sk[5]) & (g1195) & (g1453) & (g1510) & (!g1522)));
	assign g1524 = (((!g10) & (!g16) & (!g5) & (!sk[6]) & (!g78) & (g1480)) + ((!g10) & (!g16) & (!g5) & (!sk[6]) & (g78) & (g1480)) + ((!g10) & (!g16) & (!g5) & (sk[6]) & (!g78) & (g1480)) + ((!g10) & (!g16) & (g5) & (!sk[6]) & (!g78) & (g1480)) + ((!g10) & (!g16) & (g5) & (!sk[6]) & (g78) & (g1480)) + ((!g10) & (!g16) & (g5) & (sk[6]) & (!g78) & (g1480)) + ((!g10) & (g16) & (!g5) & (!sk[6]) & (!g78) & (g1480)) + ((!g10) & (g16) & (!g5) & (!sk[6]) & (g78) & (g1480)) + ((!g10) & (g16) & (!g5) & (sk[6]) & (!g78) & (!g1480)) + ((!g10) & (g16) & (!g5) & (sk[6]) & (!g78) & (g1480)) + ((!g10) & (g16) & (!g5) & (sk[6]) & (g78) & (!g1480)) + ((!g10) & (g16) & (!g5) & (sk[6]) & (g78) & (g1480)) + ((!g10) & (g16) & (g5) & (!sk[6]) & (!g78) & (g1480)) + ((!g10) & (g16) & (g5) & (!sk[6]) & (g78) & (g1480)) + ((!g10) & (g16) & (g5) & (sk[6]) & (!g78) & (!g1480)) + ((!g10) & (g16) & (g5) & (sk[6]) & (!g78) & (g1480)) + ((g10) & (!g16) & (!g5) & (!sk[6]) & (!g78) & (!g1480)) + ((g10) & (!g16) & (!g5) & (!sk[6]) & (!g78) & (g1480)) + ((g10) & (!g16) & (!g5) & (!sk[6]) & (g78) & (!g1480)) + ((g10) & (!g16) & (!g5) & (!sk[6]) & (g78) & (g1480)) + ((g10) & (!g16) & (!g5) & (sk[6]) & (!g78) & (g1480)) + ((g10) & (!g16) & (g5) & (!sk[6]) & (!g78) & (!g1480)) + ((g10) & (!g16) & (g5) & (!sk[6]) & (!g78) & (g1480)) + ((g10) & (!g16) & (g5) & (!sk[6]) & (g78) & (!g1480)) + ((g10) & (!g16) & (g5) & (!sk[6]) & (g78) & (g1480)) + ((g10) & (!g16) & (g5) & (sk[6]) & (!g78) & (g1480)) + ((g10) & (g16) & (!g5) & (!sk[6]) & (!g78) & (!g1480)) + ((g10) & (g16) & (!g5) & (!sk[6]) & (!g78) & (g1480)) + ((g10) & (g16) & (!g5) & (!sk[6]) & (g78) & (!g1480)) + ((g10) & (g16) & (!g5) & (!sk[6]) & (g78) & (g1480)) + ((g10) & (g16) & (!g5) & (sk[6]) & (!g78) & (g1480)) + ((g10) & (g16) & (g5) & (!sk[6]) & (!g78) & (!g1480)) + ((g10) & (g16) & (g5) & (!sk[6]) & (!g78) & (g1480)) + ((g10) & (g16) & (g5) & (!sk[6]) & (g78) & (!g1480)) + ((g10) & (g16) & (g5) & (!sk[6]) & (g78) & (g1480)) + ((g10) & (g16) & (g5) & (sk[6]) & (!g78) & (g1480)));
	assign o_35_ = (((!g12) & (!g73) & (!sk[7]) & (g1464) & (g1524)) + ((!g12) & (g73) & (!sk[7]) & (!g1464) & (!g1524)) + ((!g12) & (g73) & (!sk[7]) & (!g1464) & (g1524)) + ((!g12) & (g73) & (!sk[7]) & (g1464) & (!g1524)) + ((!g12) & (g73) & (!sk[7]) & (g1464) & (g1524)) + ((!g12) & (g73) & (sk[7]) & (!g1464) & (!g1524)) + ((!g12) & (g73) & (sk[7]) & (g1464) & (!g1524)) + ((g12) & (!g73) & (!sk[7]) & (g1464) & (!g1524)) + ((g12) & (!g73) & (!sk[7]) & (g1464) & (g1524)) + ((g12) & (g73) & (!sk[7]) & (!g1464) & (!g1524)) + ((g12) & (g73) & (!sk[7]) & (!g1464) & (g1524)) + ((g12) & (g73) & (!sk[7]) & (g1464) & (!g1524)) + ((g12) & (g73) & (!sk[7]) & (g1464) & (g1524)) + ((g12) & (g73) & (sk[7]) & (!g1464) & (!g1524)) + ((g12) & (g73) & (sk[7]) & (!g1464) & (g1524)) + ((g12) & (g73) & (sk[7]) & (g1464) & (!g1524)));
	assign g1526 = (((!i_8_) & (!g30) & (g5) & (!sk[8]) & (g61)) + ((!i_8_) & (g30) & (!g5) & (!sk[8]) & (!g61)) + ((!i_8_) & (g30) & (!g5) & (!sk[8]) & (g61)) + ((!i_8_) & (g30) & (!g5) & (sk[8]) & (g61)) + ((!i_8_) & (g30) & (g5) & (!sk[8]) & (!g61)) + ((!i_8_) & (g30) & (g5) & (!sk[8]) & (g61)) + ((!i_8_) & (g30) & (g5) & (sk[8]) & (g61)) + ((i_8_) & (!g30) & (g5) & (!sk[8]) & (!g61)) + ((i_8_) & (!g30) & (g5) & (!sk[8]) & (g61)) + ((i_8_) & (g30) & (!g5) & (!sk[8]) & (!g61)) + ((i_8_) & (g30) & (!g5) & (!sk[8]) & (g61)) + ((i_8_) & (g30) & (g5) & (!sk[8]) & (!g61)) + ((i_8_) & (g30) & (g5) & (!sk[8]) & (g61)) + ((i_8_) & (g30) & (g5) & (sk[8]) & (g61)));
	assign g1527 = (((!g38) & (!g64) & (!sk[9]) & (!g101) & (!g531) & (g1526)) + ((!g38) & (!g64) & (!sk[9]) & (!g101) & (g531) & (g1526)) + ((!g38) & (!g64) & (!sk[9]) & (g101) & (!g531) & (g1526)) + ((!g38) & (!g64) & (!sk[9]) & (g101) & (g531) & (g1526)) + ((!g38) & (!g64) & (sk[9]) & (!g101) & (!g531) & (!g1526)) + ((!g38) & (!g64) & (sk[9]) & (!g101) & (g531) & (!g1526)) + ((!g38) & (!g64) & (sk[9]) & (g101) & (!g531) & (!g1526)) + ((!g38) & (g64) & (!sk[9]) & (!g101) & (!g531) & (g1526)) + ((!g38) & (g64) & (!sk[9]) & (!g101) & (g531) & (g1526)) + ((!g38) & (g64) & (!sk[9]) & (g101) & (!g531) & (g1526)) + ((!g38) & (g64) & (!sk[9]) & (g101) & (g531) & (g1526)) + ((!g38) & (g64) & (sk[9]) & (!g101) & (!g531) & (!g1526)) + ((!g38) & (g64) & (sk[9]) & (!g101) & (g531) & (!g1526)) + ((!g38) & (g64) & (sk[9]) & (g101) & (!g531) & (!g1526)) + ((g38) & (!g64) & (!sk[9]) & (!g101) & (!g531) & (!g1526)) + ((g38) & (!g64) & (!sk[9]) & (!g101) & (!g531) & (g1526)) + ((g38) & (!g64) & (!sk[9]) & (!g101) & (g531) & (!g1526)) + ((g38) & (!g64) & (!sk[9]) & (!g101) & (g531) & (g1526)) + ((g38) & (!g64) & (!sk[9]) & (g101) & (!g531) & (!g1526)) + ((g38) & (!g64) & (!sk[9]) & (g101) & (!g531) & (g1526)) + ((g38) & (!g64) & (!sk[9]) & (g101) & (g531) & (!g1526)) + ((g38) & (!g64) & (!sk[9]) & (g101) & (g531) & (g1526)) + ((g38) & (!g64) & (sk[9]) & (!g101) & (!g531) & (!g1526)) + ((g38) & (!g64) & (sk[9]) & (!g101) & (g531) & (!g1526)) + ((g38) & (!g64) & (sk[9]) & (g101) & (!g531) & (!g1526)) + ((g38) & (g64) & (!sk[9]) & (!g101) & (!g531) & (!g1526)) + ((g38) & (g64) & (!sk[9]) & (!g101) & (!g531) & (g1526)) + ((g38) & (g64) & (!sk[9]) & (!g101) & (g531) & (!g1526)) + ((g38) & (g64) & (!sk[9]) & (!g101) & (g531) & (g1526)) + ((g38) & (g64) & (!sk[9]) & (g101) & (!g531) & (!g1526)) + ((g38) & (g64) & (!sk[9]) & (g101) & (!g531) & (g1526)) + ((g38) & (g64) & (!sk[9]) & (g101) & (g531) & (!g1526)) + ((g38) & (g64) & (!sk[9]) & (g101) & (g531) & (g1526)));
	assign g1528 = (((!g31) & (!g25) & (!g27) & (!sk[10]) & (!g64) & (g1527)) + ((!g31) & (!g25) & (!g27) & (!sk[10]) & (g64) & (g1527)) + ((!g31) & (!g25) & (!g27) & (sk[10]) & (!g64) & (g1527)) + ((!g31) & (!g25) & (!g27) & (sk[10]) & (g64) & (g1527)) + ((!g31) & (!g25) & (g27) & (!sk[10]) & (!g64) & (g1527)) + ((!g31) & (!g25) & (g27) & (!sk[10]) & (g64) & (g1527)) + ((!g31) & (!g25) & (g27) & (sk[10]) & (!g64) & (g1527)) + ((!g31) & (g25) & (!g27) & (!sk[10]) & (!g64) & (g1527)) + ((!g31) & (g25) & (!g27) & (!sk[10]) & (g64) & (g1527)) + ((!g31) & (g25) & (!g27) & (sk[10]) & (!g64) & (g1527)) + ((!g31) & (g25) & (!g27) & (sk[10]) & (g64) & (g1527)) + ((!g31) & (g25) & (g27) & (!sk[10]) & (!g64) & (g1527)) + ((!g31) & (g25) & (g27) & (!sk[10]) & (g64) & (g1527)) + ((!g31) & (g25) & (g27) & (sk[10]) & (!g64) & (g1527)) + ((!g31) & (g25) & (g27) & (sk[10]) & (g64) & (g1527)) + ((g31) & (!g25) & (!g27) & (!sk[10]) & (!g64) & (!g1527)) + ((g31) & (!g25) & (!g27) & (!sk[10]) & (!g64) & (g1527)) + ((g31) & (!g25) & (!g27) & (!sk[10]) & (g64) & (!g1527)) + ((g31) & (!g25) & (!g27) & (!sk[10]) & (g64) & (g1527)) + ((g31) & (!g25) & (!g27) & (sk[10]) & (!g64) & (g1527)) + ((g31) & (!g25) & (g27) & (!sk[10]) & (!g64) & (!g1527)) + ((g31) & (!g25) & (g27) & (!sk[10]) & (!g64) & (g1527)) + ((g31) & (!g25) & (g27) & (!sk[10]) & (g64) & (!g1527)) + ((g31) & (!g25) & (g27) & (!sk[10]) & (g64) & (g1527)) + ((g31) & (!g25) & (g27) & (sk[10]) & (!g64) & (g1527)) + ((g31) & (g25) & (!g27) & (!sk[10]) & (!g64) & (!g1527)) + ((g31) & (g25) & (!g27) & (!sk[10]) & (!g64) & (g1527)) + ((g31) & (g25) & (!g27) & (!sk[10]) & (g64) & (!g1527)) + ((g31) & (g25) & (!g27) & (!sk[10]) & (g64) & (g1527)) + ((g31) & (g25) & (!g27) & (sk[10]) & (!g64) & (g1527)) + ((g31) & (g25) & (!g27) & (sk[10]) & (g64) & (g1527)) + ((g31) & (g25) & (g27) & (!sk[10]) & (!g64) & (!g1527)) + ((g31) & (g25) & (g27) & (!sk[10]) & (!g64) & (g1527)) + ((g31) & (g25) & (g27) & (!sk[10]) & (g64) & (!g1527)) + ((g31) & (g25) & (g27) & (!sk[10]) & (g64) & (g1527)) + ((g31) & (g25) & (g27) & (sk[10]) & (!g64) & (g1527)) + ((g31) & (g25) & (g27) & (sk[10]) & (g64) & (g1527)));
	assign g1529 = (((g83) & (g976) & (g985) & (g994) & (g999) & (g1528)));
	assign g1530 = (((!g73) & (!g1018) & (!g1442) & (!g1453) & (!g1459) & (!g1529)) + ((!g73) & (!g1018) & (!g1442) & (!g1453) & (!g1459) & (g1529)) + ((!g73) & (!g1018) & (!g1442) & (!g1453) & (g1459) & (!g1529)) + ((!g73) & (!g1018) & (!g1442) & (!g1453) & (g1459) & (g1529)) + ((!g73) & (!g1018) & (!g1442) & (g1453) & (!g1459) & (!g1529)) + ((!g73) & (!g1018) & (!g1442) & (g1453) & (!g1459) & (g1529)) + ((!g73) & (!g1018) & (!g1442) & (g1453) & (g1459) & (!g1529)) + ((!g73) & (!g1018) & (!g1442) & (g1453) & (g1459) & (g1529)) + ((!g73) & (!g1018) & (g1442) & (!g1453) & (!g1459) & (!g1529)) + ((!g73) & (!g1018) & (g1442) & (!g1453) & (!g1459) & (g1529)) + ((!g73) & (!g1018) & (g1442) & (!g1453) & (g1459) & (!g1529)) + ((!g73) & (!g1018) & (g1442) & (!g1453) & (g1459) & (g1529)) + ((!g73) & (!g1018) & (g1442) & (g1453) & (!g1459) & (!g1529)) + ((!g73) & (!g1018) & (g1442) & (g1453) & (!g1459) & (g1529)) + ((!g73) & (!g1018) & (g1442) & (g1453) & (g1459) & (!g1529)) + ((!g73) & (!g1018) & (g1442) & (g1453) & (g1459) & (g1529)) + ((!g73) & (g1018) & (!g1442) & (!g1453) & (!g1459) & (!g1529)) + ((!g73) & (g1018) & (!g1442) & (!g1453) & (!g1459) & (g1529)) + ((!g73) & (g1018) & (!g1442) & (!g1453) & (g1459) & (!g1529)) + ((!g73) & (g1018) & (!g1442) & (!g1453) & (g1459) & (g1529)) + ((!g73) & (g1018) & (!g1442) & (g1453) & (!g1459) & (!g1529)) + ((!g73) & (g1018) & (!g1442) & (g1453) & (!g1459) & (g1529)) + ((!g73) & (g1018) & (!g1442) & (g1453) & (g1459) & (!g1529)) + ((!g73) & (g1018) & (!g1442) & (g1453) & (g1459) & (g1529)) + ((!g73) & (g1018) & (g1442) & (!g1453) & (!g1459) & (!g1529)) + ((!g73) & (g1018) & (g1442) & (!g1453) & (!g1459) & (g1529)) + ((!g73) & (g1018) & (g1442) & (!g1453) & (g1459) & (!g1529)) + ((!g73) & (g1018) & (g1442) & (!g1453) & (g1459) & (g1529)) + ((!g73) & (g1018) & (g1442) & (g1453) & (!g1459) & (!g1529)) + ((!g73) & (g1018) & (g1442) & (g1453) & (!g1459) & (g1529)) + ((!g73) & (g1018) & (g1442) & (g1453) & (g1459) & (!g1529)) + ((!g73) & (g1018) & (g1442) & (g1453) & (g1459) & (g1529)) + ((g73) & (g1018) & (!g1442) & (g1453) & (g1459) & (g1529)));
	assign g1531 = (((!g26) & (sk[13]) & (!g27) & (!g38)) + ((g26) & (!sk[13]) & (!g27) & (!g38)) + ((g26) & (!sk[13]) & (!g27) & (g38)) + ((g26) & (!sk[13]) & (g27) & (!g38)) + ((g26) & (!sk[13]) & (g27) & (g38)) + ((g26) & (sk[13]) & (!g27) & (!g38)) + ((g26) & (sk[13]) & (g27) & (!g38)));
	assign g1532 = (((!i_8_) & (!g30) & (!sk[14]) & (g5) & (g62)) + ((!i_8_) & (g30) & (!sk[14]) & (!g5) & (!g62)) + ((!i_8_) & (g30) & (!sk[14]) & (!g5) & (g62)) + ((!i_8_) & (g30) & (!sk[14]) & (g5) & (!g62)) + ((!i_8_) & (g30) & (!sk[14]) & (g5) & (g62)) + ((!i_8_) & (g30) & (sk[14]) & (!g5) & (g62)) + ((!i_8_) & (g30) & (sk[14]) & (g5) & (g62)) + ((i_8_) & (!g30) & (!sk[14]) & (g5) & (!g62)) + ((i_8_) & (!g30) & (!sk[14]) & (g5) & (g62)) + ((i_8_) & (g30) & (!sk[14]) & (!g5) & (!g62)) + ((i_8_) & (g30) & (!sk[14]) & (!g5) & (g62)) + ((i_8_) & (g30) & (!sk[14]) & (g5) & (!g62)) + ((i_8_) & (g30) & (!sk[14]) & (g5) & (g62)) + ((i_8_) & (g30) & (sk[14]) & (g5) & (g62)));
	assign o_37_ = (((!g37) & (!sk[15]) & (!g65) & (!g73) & (!g1531) & (g1532)) + ((!g37) & (!sk[15]) & (!g65) & (!g73) & (g1531) & (g1532)) + ((!g37) & (!sk[15]) & (!g65) & (g73) & (!g1531) & (g1532)) + ((!g37) & (!sk[15]) & (!g65) & (g73) & (g1531) & (g1532)) + ((!g37) & (!sk[15]) & (g65) & (!g73) & (!g1531) & (g1532)) + ((!g37) & (!sk[15]) & (g65) & (!g73) & (g1531) & (g1532)) + ((!g37) & (!sk[15]) & (g65) & (g73) & (!g1531) & (g1532)) + ((!g37) & (!sk[15]) & (g65) & (g73) & (g1531) & (g1532)) + ((!g37) & (sk[15]) & (!g65) & (g73) & (!g1531) & (!g1532)) + ((!g37) & (sk[15]) & (!g65) & (g73) & (!g1531) & (g1532)) + ((!g37) & (sk[15]) & (!g65) & (g73) & (g1531) & (!g1532)) + ((!g37) & (sk[15]) & (!g65) & (g73) & (g1531) & (g1532)) + ((!g37) & (sk[15]) & (g65) & (g73) & (!g1531) & (!g1532)) + ((!g37) & (sk[15]) & (g65) & (g73) & (!g1531) & (g1532)) + ((!g37) & (sk[15]) & (g65) & (g73) & (g1531) & (!g1532)) + ((!g37) & (sk[15]) & (g65) & (g73) & (g1531) & (g1532)) + ((g37) & (!sk[15]) & (!g65) & (!g73) & (!g1531) & (!g1532)) + ((g37) & (!sk[15]) & (!g65) & (!g73) & (!g1531) & (g1532)) + ((g37) & (!sk[15]) & (!g65) & (!g73) & (g1531) & (!g1532)) + ((g37) & (!sk[15]) & (!g65) & (!g73) & (g1531) & (g1532)) + ((g37) & (!sk[15]) & (!g65) & (g73) & (!g1531) & (!g1532)) + ((g37) & (!sk[15]) & (!g65) & (g73) & (!g1531) & (g1532)) + ((g37) & (!sk[15]) & (!g65) & (g73) & (g1531) & (!g1532)) + ((g37) & (!sk[15]) & (!g65) & (g73) & (g1531) & (g1532)) + ((g37) & (!sk[15]) & (g65) & (!g73) & (!g1531) & (!g1532)) + ((g37) & (!sk[15]) & (g65) & (!g73) & (!g1531) & (g1532)) + ((g37) & (!sk[15]) & (g65) & (!g73) & (g1531) & (!g1532)) + ((g37) & (!sk[15]) & (g65) & (!g73) & (g1531) & (g1532)) + ((g37) & (!sk[15]) & (g65) & (g73) & (!g1531) & (!g1532)) + ((g37) & (!sk[15]) & (g65) & (g73) & (!g1531) & (g1532)) + ((g37) & (!sk[15]) & (g65) & (g73) & (g1531) & (!g1532)) + ((g37) & (!sk[15]) & (g65) & (g73) & (g1531) & (g1532)) + ((g37) & (sk[15]) & (!g65) & (g73) & (!g1531) & (g1532)) + ((g37) & (sk[15]) & (!g65) & (g73) & (g1531) & (g1532)) + ((g37) & (sk[15]) & (g65) & (g73) & (!g1531) & (!g1532)) + ((g37) & (sk[15]) & (g65) & (g73) & (!g1531) & (g1532)) + ((g37) & (sk[15]) & (g65) & (g73) & (g1531) & (g1532)));
	assign o_38_ = (((!i_3_) & (!i_4_) & (!sk[16]) & (g1) & (g34)) + ((!i_3_) & (i_4_) & (!sk[16]) & (!g1) & (!g34)) + ((!i_3_) & (i_4_) & (!sk[16]) & (!g1) & (g34)) + ((!i_3_) & (i_4_) & (!sk[16]) & (g1) & (!g34)) + ((!i_3_) & (i_4_) & (!sk[16]) & (g1) & (g34)) + ((i_3_) & (!i_4_) & (!sk[16]) & (g1) & (!g34)) + ((i_3_) & (!i_4_) & (!sk[16]) & (g1) & (g34)) + ((i_3_) & (i_4_) & (!sk[16]) & (!g1) & (!g34)) + ((i_3_) & (i_4_) & (!sk[16]) & (!g1) & (g34)) + ((i_3_) & (i_4_) & (!sk[16]) & (g1) & (!g34)) + ((i_3_) & (i_4_) & (!sk[16]) & (g1) & (g34)) + ((i_3_) & (i_4_) & (sk[16]) & (g1) & (g34)));
	assign o_39_ = (((!i_3_) & (!i_4_) & (!g1) & (!i_6_) & (!sk[17]) & (i_7_)) + ((!i_3_) & (!i_4_) & (!g1) & (i_6_) & (!sk[17]) & (i_7_)) + ((!i_3_) & (!i_4_) & (g1) & (!i_6_) & (!sk[17]) & (i_7_)) + ((!i_3_) & (!i_4_) & (g1) & (i_6_) & (!sk[17]) & (i_7_)) + ((!i_3_) & (i_4_) & (!g1) & (!i_6_) & (!sk[17]) & (i_7_)) + ((!i_3_) & (i_4_) & (!g1) & (i_6_) & (!sk[17]) & (i_7_)) + ((!i_3_) & (i_4_) & (g1) & (!i_6_) & (!sk[17]) & (i_7_)) + ((!i_3_) & (i_4_) & (g1) & (i_6_) & (!sk[17]) & (i_7_)) + ((i_3_) & (!i_4_) & (!g1) & (!i_6_) & (!sk[17]) & (!i_7_)) + ((i_3_) & (!i_4_) & (!g1) & (!i_6_) & (!sk[17]) & (i_7_)) + ((i_3_) & (!i_4_) & (!g1) & (i_6_) & (!sk[17]) & (!i_7_)) + ((i_3_) & (!i_4_) & (!g1) & (i_6_) & (!sk[17]) & (i_7_)) + ((i_3_) & (!i_4_) & (g1) & (!i_6_) & (!sk[17]) & (!i_7_)) + ((i_3_) & (!i_4_) & (g1) & (!i_6_) & (!sk[17]) & (i_7_)) + ((i_3_) & (!i_4_) & (g1) & (i_6_) & (!sk[17]) & (!i_7_)) + ((i_3_) & (!i_4_) & (g1) & (i_6_) & (!sk[17]) & (i_7_)) + ((i_3_) & (i_4_) & (!g1) & (!i_6_) & (!sk[17]) & (!i_7_)) + ((i_3_) & (i_4_) & (!g1) & (!i_6_) & (!sk[17]) & (i_7_)) + ((i_3_) & (i_4_) & (!g1) & (i_6_) & (!sk[17]) & (!i_7_)) + ((i_3_) & (i_4_) & (!g1) & (i_6_) & (!sk[17]) & (i_7_)) + ((i_3_) & (i_4_) & (g1) & (!i_6_) & (!sk[17]) & (!i_7_)) + ((i_3_) & (i_4_) & (g1) & (!i_6_) & (!sk[17]) & (i_7_)) + ((i_3_) & (i_4_) & (g1) & (i_6_) & (!sk[17]) & (!i_7_)) + ((i_3_) & (i_4_) & (g1) & (i_6_) & (!sk[17]) & (i_7_)) + ((i_3_) & (i_4_) & (g1) & (i_6_) & (sk[17]) & (!i_7_)));
	assign g1536 = (((!g95) & (!i_13_) & (!i_12_) & (!i_14_) & (!g93) & (g108)) + ((g95) & (!i_13_) & (!i_12_) & (!i_14_) & (!g93) & (g108)) + ((g95) & (!i_13_) & (!i_12_) & (i_14_) & (!g93) & (g108)) + ((g95) & (!i_13_) & (!i_12_) & (i_14_) & (g93) & (g108)) + ((g95) & (!i_13_) & (i_12_) & (!i_14_) & (!g93) & (g108)) + ((g95) & (!i_13_) & (i_12_) & (!i_14_) & (g93) & (g108)) + ((g95) & (i_13_) & (i_12_) & (!i_14_) & (!g93) & (g108)) + ((g95) & (i_13_) & (i_12_) & (!i_14_) & (g93) & (g108)));
	assign g1537 = (((!g95) & (!i_13_) & (!i_12_) & (!i_14_) & (!g93) & (g108)) + ((!g95) & (!i_13_) & (i_12_) & (!i_14_) & (!g93) & (g108)) + ((!g95) & (!i_13_) & (i_12_) & (i_14_) & (!g93) & (g108)) + ((!g95) & (i_13_) & (!i_12_) & (!i_14_) & (!g93) & (g108)) + ((!g95) & (i_13_) & (i_12_) & (!i_14_) & (!g93) & (g108)) + ((g95) & (!i_13_) & (!i_12_) & (!i_14_) & (!g93) & (g108)) + ((g95) & (!i_13_) & (!i_12_) & (i_14_) & (!g93) & (g108)) + ((g95) & (!i_13_) & (!i_12_) & (i_14_) & (g93) & (g108)) + ((g95) & (!i_13_) & (i_12_) & (!i_14_) & (!g93) & (g108)) + ((g95) & (!i_13_) & (i_12_) & (!i_14_) & (g93) & (g108)) + ((g95) & (!i_13_) & (i_12_) & (i_14_) & (!g93) & (g108)) + ((g95) & (!i_13_) & (i_12_) & (i_14_) & (g93) & (g108)) + ((g95) & (i_13_) & (!i_12_) & (!i_14_) & (!g93) & (g108)) + ((g95) & (i_13_) & (i_12_) & (!i_14_) & (!g93) & (g108)) + ((g95) & (i_13_) & (i_12_) & (!i_14_) & (g93) & (g108)));
	assign g1538 = (((!sk[20]) & (g1536) & (!g1537) & (!i_8_)) + ((!sk[20]) & (g1536) & (!g1537) & (i_8_)) + ((!sk[20]) & (g1536) & (g1537) & (!i_8_)) + ((!sk[20]) & (g1536) & (g1537) & (i_8_)) + ((sk[20]) & (!g1536) & (!g1537) & (!i_8_)) + ((sk[20]) & (!g1536) & (!g1537) & (i_8_)) + ((sk[20]) & (!g1536) & (g1537) & (!i_8_)) + ((sk[20]) & (g1536) & (!g1537) & (i_8_)));
	assign g1539 = (((!g22) & (!i_13_) & (i_12_) & (!i_14_) & (g11) & (g88)) + ((!g22) & (!i_13_) & (i_12_) & (i_14_) & (g11) & (g88)) + ((!g22) & (i_13_) & (!i_12_) & (!i_14_) & (g11) & (g88)) + ((!g22) & (i_13_) & (i_12_) & (!i_14_) & (g11) & (g88)) + ((g22) & (!i_13_) & (!i_12_) & (!i_14_) & (!g11) & (g88)) + ((g22) & (!i_13_) & (!i_12_) & (!i_14_) & (g11) & (g88)) + ((g22) & (!i_13_) & (i_12_) & (!i_14_) & (!g11) & (g88)) + ((g22) & (!i_13_) & (i_12_) & (!i_14_) & (g11) & (g88)) + ((g22) & (!i_13_) & (i_12_) & (i_14_) & (!g11) & (g88)) + ((g22) & (!i_13_) & (i_12_) & (i_14_) & (g11) & (g88)) + ((g22) & (i_13_) & (!i_12_) & (!i_14_) & (!g11) & (g88)) + ((g22) & (i_13_) & (!i_12_) & (!i_14_) & (g11) & (g88)) + ((g22) & (i_13_) & (i_12_) & (!i_14_) & (!g11) & (g88)) + ((g22) & (i_13_) & (i_12_) & (!i_14_) & (g11) & (g88)) + ((g22) & (i_13_) & (i_12_) & (i_14_) & (!g11) & (g88)) + ((g22) & (i_13_) & (i_12_) & (i_14_) & (g11) & (g88)));
	assign g1540 = (((!g22) & (!i_13_) & (i_12_) & (!i_14_) & (g11) & (g88)) + ((!g22) & (i_13_) & (!i_12_) & (!i_14_) & (g11) & (g88)) + ((g22) & (!i_13_) & (i_12_) & (!i_14_) & (g11) & (g88)) + ((g22) & (!i_13_) & (i_12_) & (i_14_) & (!g11) & (g88)) + ((g22) & (!i_13_) & (i_12_) & (i_14_) & (g11) & (g88)) + ((g22) & (i_13_) & (!i_12_) & (!i_14_) & (g11) & (g88)) + ((g22) & (i_13_) & (i_12_) & (i_14_) & (!g11) & (g88)) + ((g22) & (i_13_) & (i_12_) & (i_14_) & (g11) & (g88)));
	assign g1541 = (((!sk[23]) & (g1539) & (!g1540) & (!i_8_)) + ((!sk[23]) & (g1539) & (!g1540) & (i_8_)) + ((!sk[23]) & (g1539) & (g1540) & (!i_8_)) + ((!sk[23]) & (g1539) & (g1540) & (i_8_)) + ((sk[23]) & (!g1539) & (!g1540) & (!i_8_)) + ((sk[23]) & (!g1539) & (!g1540) & (i_8_)) + ((sk[23]) & (!g1539) & (g1540) & (!i_8_)) + ((sk[23]) & (g1539) & (!g1540) & (i_8_)));
	assign g1542 = (((!sk[24]) & (!g158) & (!g131) & (g1027) & (g99)) + ((!sk[24]) & (!g158) & (g131) & (!g1027) & (!g99)) + ((!sk[24]) & (!g158) & (g131) & (!g1027) & (g99)) + ((!sk[24]) & (!g158) & (g131) & (g1027) & (!g99)) + ((!sk[24]) & (!g158) & (g131) & (g1027) & (g99)) + ((!sk[24]) & (g158) & (!g131) & (g1027) & (!g99)) + ((!sk[24]) & (g158) & (!g131) & (g1027) & (g99)) + ((!sk[24]) & (g158) & (g131) & (!g1027) & (!g99)) + ((!sk[24]) & (g158) & (g131) & (!g1027) & (g99)) + ((!sk[24]) & (g158) & (g131) & (g1027) & (!g99)) + ((!sk[24]) & (g158) & (g131) & (g1027) & (g99)) + ((sk[24]) & (!g158) & (!g131) & (!g1027) & (!g99)) + ((sk[24]) & (!g158) & (!g131) & (!g1027) & (g99)) + ((sk[24]) & (!g158) & (g131) & (!g1027) & (!g99)) + ((sk[24]) & (g158) & (!g131) & (!g1027) & (!g99)) + ((sk[24]) & (g158) & (g131) & (!g1027) & (!g99)));
	assign g1543 = (((!g183) & (!g88) & (!g196) & (!g194) & (!g192) & (!g190)) + ((!g183) & (g88) & (!g196) & (!g194) & (!g192) & (!g190)) + ((g183) & (!g88) & (!g196) & (!g194) & (!g192) & (!g190)));
	assign g1544 = (((!g10) & (!g20) & (!g19) & (!g77) & (!g75) & (!g8)) + ((!g10) & (!g20) & (!g19) & (!g77) & (!g75) & (g8)) + ((!g10) & (!g20) & (g19) & (!g77) & (!g75) & (!g8)) + ((!g10) & (!g20) & (g19) & (!g77) & (!g75) & (g8)) + ((!g10) & (g20) & (!g19) & (!g77) & (!g75) & (!g8)) + ((!g10) & (g20) & (!g19) & (!g77) & (!g75) & (g8)) + ((!g10) & (g20) & (!g19) & (!g77) & (g75) & (g8)) + ((!g10) & (g20) & (g19) & (!g77) & (!g75) & (!g8)) + ((!g10) & (g20) & (g19) & (!g77) & (!g75) & (g8)) + ((g10) & (!g20) & (!g19) & (!g77) & (!g75) & (!g8)) + ((g10) & (!g20) & (!g19) & (!g77) & (!g75) & (g8)) + ((g10) & (!g20) & (g19) & (!g77) & (!g75) & (!g8)) + ((g10) & (!g20) & (g19) & (!g77) & (!g75) & (g8)) + ((g10) & (g20) & (!g19) & (!g77) & (!g75) & (!g8)) + ((g10) & (g20) & (!g19) & (!g77) & (!g75) & (g8)) + ((g10) & (g20) & (g19) & (!g77) & (!g75) & (!g8)) + ((g10) & (g20) & (g19) & (!g77) & (!g75) & (g8)));
	assign g1545 = (((!g1546) & (sk[27]) & (!g1547)) + ((g1546) & (!sk[27]) & (!g1547)) + ((g1546) & (!sk[27]) & (g1547)));
	assign g1546 = (((!sk[28]) & (g544) & (!g1548)) + ((!sk[28]) & (g544) & (g1548)) + ((sk[28]) & (!g544) & (g1548)));
	assign g1547 = (((g544) & (!sk[29]) & (!g1551)) + ((g544) & (!sk[29]) & (g1551)) + ((g544) & (sk[29]) & (g1551)));
	assign g1548 = (((!g1549) & (sk[30]) & (!g1550)) + ((g1549) & (!sk[30]) & (!g1550)) + ((g1549) & (!sk[30]) & (g1550)));
	assign g1549 = (((!sk[31]) & (i_8_) & (!g1554)) + ((!sk[31]) & (i_8_) & (g1554)) + ((sk[31]) & (!i_8_) & (g1554)));
	assign g1550 = (((i_8_) & (!sk[32]) & (!g1555)) + ((i_8_) & (!sk[32]) & (g1555)) + ((i_8_) & (sk[32]) & (g1555)));
	assign g1551 = (((!sk[33]) & (g1552) & (!g1553)) + ((!sk[33]) & (g1552) & (g1553)) + ((sk[33]) & (!g1552) & (!g1553)));
	assign g1552 = (((!i_8_) & (sk[34]) & (g1556)) + ((i_8_) & (!sk[34]) & (!g1556)) + ((i_8_) & (!sk[34]) & (g1556)));
	assign g1553 = (((i_8_) & (!sk[35]) & (!g1557)) + ((i_8_) & (!sk[35]) & (g1557)) + ((i_8_) & (sk[35]) & (g1557)));
	assign g1554 = (((!g108) & (sk[36]) & (g1450) & (!g470)) + ((!g108) & (sk[36]) & (g1450) & (g470)) + ((g108) & (!sk[36]) & (!g1450) & (!g470)) + ((g108) & (!sk[36]) & (!g1450) & (g470)) + ((g108) & (!sk[36]) & (g1450) & (!g470)) + ((g108) & (!sk[36]) & (g1450) & (g470)) + ((g108) & (sk[36]) & (g1450) & (!g470)));
	assign g1555 = (((!sk[37]) & (g108) & (!g1450)) + ((!sk[37]) & (g108) & (g1450)) + ((sk[37]) & (!g108) & (g1450)));
	assign g1556 = (((!g108) & (g1450) & (sk[38]) & (!g470)) + ((!g108) & (g1450) & (sk[38]) & (g470)) + ((g108) & (!g1450) & (!sk[38]) & (!g470)) + ((g108) & (!g1450) & (!sk[38]) & (g470)) + ((g108) & (g1450) & (!sk[38]) & (!g470)) + ((g108) & (g1450) & (!sk[38]) & (g470)) + ((g108) & (g1450) & (sk[38]) & (!g470)));
	assign g1557 = (((!g108) & (!g1450) & (!sk[39]) & (g204) & (g848)) + ((!g108) & (g1450) & (!sk[39]) & (!g204) & (!g848)) + ((!g108) & (g1450) & (!sk[39]) & (!g204) & (g848)) + ((!g108) & (g1450) & (!sk[39]) & (g204) & (!g848)) + ((!g108) & (g1450) & (!sk[39]) & (g204) & (g848)) + ((!g108) & (g1450) & (sk[39]) & (!g204) & (!g848)) + ((!g108) & (g1450) & (sk[39]) & (!g204) & (g848)) + ((!g108) & (g1450) & (sk[39]) & (g204) & (!g848)) + ((!g108) & (g1450) & (sk[39]) & (g204) & (g848)) + ((g108) & (!g1450) & (!sk[39]) & (g204) & (!g848)) + ((g108) & (!g1450) & (!sk[39]) & (g204) & (g848)) + ((g108) & (g1450) & (!sk[39]) & (!g204) & (!g848)) + ((g108) & (g1450) & (!sk[39]) & (!g204) & (g848)) + ((g108) & (g1450) & (!sk[39]) & (g204) & (!g848)) + ((g108) & (g1450) & (!sk[39]) & (g204) & (g848)) + ((g108) & (g1450) & (sk[39]) & (g204) & (g848)));
	assign g1558 = (((!sk[40]) & (g1559) & (!g1560)) + ((!sk[40]) & (g1559) & (g1560)) + ((sk[40]) & (!g1559) & (!g1560)));
	assign g1559 = (((!sk[41]) & (g134) & (!g1561)) + ((!sk[41]) & (g134) & (g1561)) + ((sk[41]) & (!g134) & (g1561)));
	assign g1560 = (((!sk[42]) & (g134) & (!g1564)) + ((!sk[42]) & (g134) & (g1564)) + ((sk[42]) & (g134) & (g1564)));
	assign g1561 = (((!g1562) & (sk[43]) & (!g1563)) + ((g1562) & (!sk[43]) & (!g1563)) + ((g1562) & (!sk[43]) & (g1563)));
	assign g1562 = (((!g678) & (sk[44]) & (g1566)) + ((g678) & (!sk[44]) & (!g1566)) + ((g678) & (!sk[44]) & (g1566)));
	assign g1563 = (((g678) & (!sk[45]) & (!g1411)) + ((g678) & (!sk[45]) & (g1411)) + ((g678) & (sk[45]) & (g1411)));
	assign g1564 = (((!sk[46]) & (g678) & (!g1565)) + ((!sk[46]) & (g678) & (g1565)) + ((sk[46]) & (g678) & (!g1565)));
	assign g1565 = (((!sk[47]) & (g678) & (!g1567)) + ((!sk[47]) & (g678) & (g1567)) + ((sk[47]) & (g678) & (g1567)));
	assign g1566 = (((!sk[48]) & (g118) & (!g1411)) + ((!sk[48]) & (g118) & (g1411)) + ((sk[48]) & (!g118) & (g1411)) + ((sk[48]) & (g118) & (!g1411)) + ((sk[48]) & (g118) & (g1411)));
	assign g1567 = (((!g572) & (!g93) & (!g270) & (sk[49]) & (!g1411)) + ((!g572) & (!g93) & (!g270) & (sk[49]) & (g1411)) + ((!g572) & (!g93) & (g270) & (!sk[49]) & (g1411)) + ((!g572) & (!g93) & (g270) & (sk[49]) & (g1411)) + ((!g572) & (g93) & (!g270) & (!sk[49]) & (!g1411)) + ((!g572) & (g93) & (!g270) & (!sk[49]) & (g1411)) + ((!g572) & (g93) & (!g270) & (sk[49]) & (!g1411)) + ((!g572) & (g93) & (!g270) & (sk[49]) & (g1411)) + ((!g572) & (g93) & (g270) & (!sk[49]) & (!g1411)) + ((!g572) & (g93) & (g270) & (!sk[49]) & (g1411)) + ((!g572) & (g93) & (g270) & (sk[49]) & (g1411)) + ((g572) & (!g93) & (!g270) & (sk[49]) & (!g1411)) + ((g572) & (!g93) & (!g270) & (sk[49]) & (g1411)) + ((g572) & (!g93) & (g270) & (!sk[49]) & (!g1411)) + ((g572) & (!g93) & (g270) & (!sk[49]) & (g1411)) + ((g572) & (!g93) & (g270) & (sk[49]) & (!g1411)) + ((g572) & (!g93) & (g270) & (sk[49]) & (g1411)) + ((g572) & (g93) & (!g270) & (!sk[49]) & (!g1411)) + ((g572) & (g93) & (!g270) & (!sk[49]) & (g1411)) + ((g572) & (g93) & (!g270) & (sk[49]) & (!g1411)) + ((g572) & (g93) & (!g270) & (sk[49]) & (g1411)) + ((g572) & (g93) & (g270) & (!sk[49]) & (!g1411)) + ((g572) & (g93) & (g270) & (!sk[49]) & (g1411)) + ((g572) & (g93) & (g270) & (sk[49]) & (g1411)));
	assign g1568 = (((!sk[50]) & (g1569) & (!g1570)) + ((!sk[50]) & (g1569) & (g1570)) + ((sk[50]) & (!g1569) & (!g1570)));
	assign g1569 = (((!sk[51]) & (g96) & (!g1571)) + ((!sk[51]) & (g96) & (g1571)) + ((sk[51]) & (!g96) & (g1571)));
	assign g1570 = (((g96) & (!sk[52]) & (!g1574)) + ((g96) & (!sk[52]) & (g1574)) + ((g96) & (sk[52]) & (g1574)));
	assign g1571 = (((!g1572) & (sk[53]) & (!g1573)) + ((g1572) & (!sk[53]) & (!g1573)) + ((g1572) & (!sk[53]) & (g1573)));
	assign g1572 = (((!g1384) & (sk[54]) & (g1577)) + ((g1384) & (!sk[54]) & (!g1577)) + ((g1384) & (!sk[54]) & (g1577)));
	assign g1573 = (((!sk[55]) & (g1384) & (!g1578)) + ((!sk[55]) & (g1384) & (g1578)) + ((sk[55]) & (g1384) & (g1578)));
	assign g1574 = (((!g1575) & (sk[56]) & (!g1576)) + ((g1575) & (!sk[56]) & (!g1576)) + ((g1575) & (!sk[56]) & (g1576)));
	assign g1575 = (((!g1384) & (sk[57]) & (g1579)) + ((g1384) & (!sk[57]) & (!g1579)) + ((g1384) & (!sk[57]) & (g1579)));
	assign g1576 = (((!sk[58]) & (g1384) & (!g1387)) + ((!sk[58]) & (g1384) & (g1387)) + ((sk[58]) & (g1384) & (g1387)));
	assign g1577 = (((!sk[59]) & (g135) & (!g1387)) + ((!sk[59]) & (g135) & (g1387)) + ((sk[59]) & (!g135) & (g1387)));
	assign g1578 = (((!g135) & (g1387) & (sk[60]) & (!g134)) + ((!g135) & (g1387) & (sk[60]) & (g134)) + ((g135) & (!g1387) & (!sk[60]) & (!g134)) + ((g135) & (!g1387) & (!sk[60]) & (g134)) + ((g135) & (g1387) & (!sk[60]) & (!g134)) + ((g135) & (g1387) & (!sk[60]) & (g134)) + ((g135) & (g1387) & (sk[60]) & (!g134)));
	assign g1579 = (((!sk[61]) & (!g135) & (!g1387) & (i_8_) & (g669)) + ((!sk[61]) & (!g135) & (g1387) & (!i_8_) & (!g669)) + ((!sk[61]) & (!g135) & (g1387) & (!i_8_) & (g669)) + ((!sk[61]) & (!g135) & (g1387) & (i_8_) & (!g669)) + ((!sk[61]) & (!g135) & (g1387) & (i_8_) & (g669)) + ((!sk[61]) & (g135) & (!g1387) & (i_8_) & (!g669)) + ((!sk[61]) & (g135) & (!g1387) & (i_8_) & (g669)) + ((!sk[61]) & (g135) & (g1387) & (!i_8_) & (!g669)) + ((!sk[61]) & (g135) & (g1387) & (!i_8_) & (g669)) + ((!sk[61]) & (g135) & (g1387) & (i_8_) & (!g669)) + ((!sk[61]) & (g135) & (g1387) & (i_8_) & (g669)) + ((sk[61]) & (!g135) & (g1387) & (!i_8_) & (!g669)) + ((sk[61]) & (!g135) & (g1387) & (!i_8_) & (g669)) + ((sk[61]) & (!g135) & (g1387) & (i_8_) & (!g669)) + ((sk[61]) & (!g135) & (g1387) & (i_8_) & (g669)) + ((sk[61]) & (g135) & (g1387) & (!i_8_) & (g669)));
	assign g1580 = (((!sk[62]) & (g1581) & (!g1582)) + ((!sk[62]) & (g1581) & (g1582)) + ((sk[62]) & (!g1581) & (!g1582)));
	assign g1581 = (((!sk[63]) & (i_14_) & (!g1583)) + ((!sk[63]) & (i_14_) & (g1583)) + ((sk[63]) & (!i_14_) & (g1583)));
	assign g1582 = (((i_14_) & (!sk[64]) & (!g1585)) + ((i_14_) & (!sk[64]) & (g1585)) + ((i_14_) & (sk[64]) & (g1585)));
	assign g1583 = (((i_13_) & (!sk[65]) & (!g1584)) + ((i_13_) & (!sk[65]) & (g1584)) + ((i_13_) & (sk[65]) & (!g1584)));
	assign g1584 = (((!sk[66]) & (i_13_) & (!g1587)) + ((!sk[66]) & (i_13_) & (g1587)) + ((sk[66]) & (i_13_) & (g1587)));
	assign g1585 = (((!i_13_) & (sk[67]) & (!g1586)) + ((i_13_) & (!sk[67]) & (!g1586)) + ((i_13_) & (!sk[67]) & (g1586)));
	assign g1586 = (((!sk[68]) & (i_13_) & (!g1588)) + ((!sk[68]) & (i_13_) & (g1588)) + ((sk[68]) & (!i_13_) & (g1588)));
	assign g1587 = (((!sk[69]) & (g18) & (!i_12_) & (!g135)) + ((!sk[69]) & (g18) & (!i_12_) & (g135)) + ((!sk[69]) & (g18) & (i_12_) & (!g135)) + ((!sk[69]) & (g18) & (i_12_) & (g135)) + ((sk[69]) & (!g18) & (!i_12_) & (!g135)) + ((sk[69]) & (!g18) & (!i_12_) & (g135)) + ((sk[69]) & (!g18) & (i_12_) & (!g135)) + ((sk[69]) & (g18) & (!i_12_) & (!g135)) + ((sk[69]) & (g18) & (!i_12_) & (g135)) + ((sk[69]) & (g18) & (i_12_) & (!g135)) + ((sk[69]) & (g18) & (i_12_) & (g135)));
	assign g1588 = (((!sk[70]) & (!g18) & (!i_12_) & (g212) & (g215)) + ((!sk[70]) & (!g18) & (i_12_) & (!g212) & (!g215)) + ((!sk[70]) & (!g18) & (i_12_) & (!g212) & (g215)) + ((!sk[70]) & (!g18) & (i_12_) & (g212) & (!g215)) + ((!sk[70]) & (!g18) & (i_12_) & (g212) & (g215)) + ((!sk[70]) & (g18) & (!i_12_) & (g212) & (!g215)) + ((!sk[70]) & (g18) & (!i_12_) & (g212) & (g215)) + ((!sk[70]) & (g18) & (i_12_) & (!g212) & (!g215)) + ((!sk[70]) & (g18) & (i_12_) & (!g212) & (g215)) + ((!sk[70]) & (g18) & (i_12_) & (g212) & (!g215)) + ((!sk[70]) & (g18) & (i_12_) & (g212) & (g215)) + ((sk[70]) & (!g18) & (!i_12_) & (g212) & (g215)) + ((sk[70]) & (!g18) & (i_12_) & (!g212) & (!g215)) + ((sk[70]) & (!g18) & (i_12_) & (!g212) & (g215)) + ((sk[70]) & (!g18) & (i_12_) & (g212) & (!g215)) + ((sk[70]) & (!g18) & (i_12_) & (g212) & (g215)) + ((sk[70]) & (g18) & (!i_12_) & (!g212) & (!g215)) + ((sk[70]) & (g18) & (!i_12_) & (!g212) & (g215)) + ((sk[70]) & (g18) & (!i_12_) & (g212) & (!g215)) + ((sk[70]) & (g18) & (!i_12_) & (g212) & (g215)) + ((sk[70]) & (g18) & (i_12_) & (!g212) & (!g215)) + ((sk[70]) & (g18) & (i_12_) & (!g212) & (g215)) + ((sk[70]) & (g18) & (i_12_) & (g212) & (!g215)) + ((sk[70]) & (g18) & (i_12_) & (g212) & (g215)));
	assign g1589 = (((!sk[71]) & (g108) & (!g1590)) + ((!sk[71]) & (g108) & (g1590)) + ((sk[71]) & (g108) & (!g1590)));
	assign g1590 = (((g108) & (!sk[72]) & (!g1591)) + ((g108) & (!sk[72]) & (g1591)) + ((g108) & (sk[72]) & (g1591)));
	assign g1591 = (((!sk[73]) & (g1592) & (!g1593)) + ((!sk[73]) & (g1592) & (g1593)) + ((sk[73]) & (!g1592) & (!g1593)));
	assign g1592 = (((!i_14_) & (sk[74]) & (g1594)) + ((i_14_) & (!sk[74]) & (!g1594)) + ((i_14_) & (!sk[74]) & (g1594)));
	assign g1593 = (((!sk[75]) & (i_14_) & (!g1595)) + ((!sk[75]) & (i_14_) & (g1595)) + ((sk[75]) & (i_14_) & (g1595)));
	assign g1594 = (((!i_13_) & (!i_12_) & (!g102) & (sk[76]) & (g115)) + ((!i_13_) & (!i_12_) & (g102) & (!sk[76]) & (g115)) + ((!i_13_) & (!i_12_) & (g102) & (sk[76]) & (g115)) + ((!i_13_) & (i_12_) & (!g102) & (!sk[76]) & (!g115)) + ((!i_13_) & (i_12_) & (!g102) & (!sk[76]) & (g115)) + ((!i_13_) & (i_12_) & (g102) & (!sk[76]) & (!g115)) + ((!i_13_) & (i_12_) & (g102) & (!sk[76]) & (g115)) + ((!i_13_) & (i_12_) & (g102) & (sk[76]) & (g115)) + ((i_13_) & (!i_12_) & (g102) & (!sk[76]) & (!g115)) + ((i_13_) & (!i_12_) & (g102) & (!sk[76]) & (g115)) + ((i_13_) & (!i_12_) & (g102) & (sk[76]) & (!g115)) + ((i_13_) & (!i_12_) & (g102) & (sk[76]) & (g115)) + ((i_13_) & (i_12_) & (!g102) & (!sk[76]) & (!g115)) + ((i_13_) & (i_12_) & (!g102) & (!sk[76]) & (g115)) + ((i_13_) & (i_12_) & (g102) & (!sk[76]) & (!g115)) + ((i_13_) & (i_12_) & (g102) & (!sk[76]) & (g115)) + ((i_13_) & (i_12_) & (g102) & (sk[76]) & (g115)));
	assign g1595 = (((!i_13_) & (!i_12_) & (!i_8_) & (sk[77]) & (!g115)) + ((!i_13_) & (!i_12_) & (!i_8_) & (sk[77]) & (g115)) + ((!i_13_) & (!i_12_) & (i_8_) & (!sk[77]) & (g115)) + ((!i_13_) & (!i_12_) & (i_8_) & (sk[77]) & (!g115)) + ((!i_13_) & (!i_12_) & (i_8_) & (sk[77]) & (g115)) + ((!i_13_) & (i_12_) & (!i_8_) & (!sk[77]) & (!g115)) + ((!i_13_) & (i_12_) & (!i_8_) & (!sk[77]) & (g115)) + ((!i_13_) & (i_12_) & (!i_8_) & (sk[77]) & (!g115)) + ((!i_13_) & (i_12_) & (!i_8_) & (sk[77]) & (g115)) + ((!i_13_) & (i_12_) & (i_8_) & (!sk[77]) & (!g115)) + ((!i_13_) & (i_12_) & (i_8_) & (!sk[77]) & (g115)) + ((!i_13_) & (i_12_) & (i_8_) & (sk[77]) & (g115)) + ((i_13_) & (!i_12_) & (!i_8_) & (sk[77]) & (!g115)) + ((i_13_) & (!i_12_) & (!i_8_) & (sk[77]) & (g115)) + ((i_13_) & (!i_12_) & (i_8_) & (!sk[77]) & (!g115)) + ((i_13_) & (!i_12_) & (i_8_) & (!sk[77]) & (g115)) + ((i_13_) & (!i_12_) & (i_8_) & (sk[77]) & (!g115)) + ((i_13_) & (!i_12_) & (i_8_) & (sk[77]) & (g115)) + ((i_13_) & (i_12_) & (!i_8_) & (!sk[77]) & (!g115)) + ((i_13_) & (i_12_) & (!i_8_) & (!sk[77]) & (g115)) + ((i_13_) & (i_12_) & (!i_8_) & (sk[77]) & (!g115)) + ((i_13_) & (i_12_) & (!i_8_) & (sk[77]) & (g115)) + ((i_13_) & (i_12_) & (i_8_) & (!sk[77]) & (!g115)) + ((i_13_) & (i_12_) & (i_8_) & (!sk[77]) & (g115)) + ((i_13_) & (i_12_) & (i_8_) & (sk[77]) & (!g115)) + ((i_13_) & (i_12_) & (i_8_) & (sk[77]) & (g115)));
	assign g1596 = (((!sk[78]) & (g1597) & (!g1598)) + ((!sk[78]) & (g1597) & (g1598)) + ((sk[78]) & (!g1597) & (!g1598)));
	assign g1597 = (((!g119) & (sk[79]) & (g1599)) + ((g119) & (!sk[79]) & (!g1599)) + ((g119) & (!sk[79]) & (g1599)));
	assign g1598 = (((!sk[80]) & (g119) & (!g1601)) + ((!sk[80]) & (g119) & (g1601)) + ((sk[80]) & (g119) & (g1601)));
	assign g1599 = (((!sk[81]) & (g134) & (!g1600)) + ((!sk[81]) & (g134) & (g1600)) + ((sk[81]) & (g134) & (!g1600)));
	assign g1600 = (((g134) & (!sk[82]) & (!g1604)) + ((g134) & (!sk[82]) & (g1604)) + ((g134) & (sk[82]) & (g1604)));
	assign g1601 = (((!sk[83]) & (g1602) & (!g1603)) + ((!sk[83]) & (g1602) & (g1603)) + ((sk[83]) & (!g1602) & (!g1603)));
	assign g1602 = (((!sk[84]) & (g134) & (!g1605)) + ((!sk[84]) & (g134) & (g1605)) + ((sk[84]) & (!g134) & (g1605)));
	assign g1603 = (((g134) & (!sk[85]) & (!g1606)) + ((g134) & (!sk[85]) & (g1606)) + ((g134) & (sk[85]) & (g1606)));
	assign g1604 = (((!i_13_) & (!sk[86]) & (!i_12_) & (g122) & (i_14_)) + ((!i_13_) & (!sk[86]) & (i_12_) & (!g122) & (!i_14_)) + ((!i_13_) & (!sk[86]) & (i_12_) & (!g122) & (i_14_)) + ((!i_13_) & (!sk[86]) & (i_12_) & (g122) & (!i_14_)) + ((!i_13_) & (!sk[86]) & (i_12_) & (g122) & (i_14_)) + ((!i_13_) & (sk[86]) & (!i_12_) & (!g122) & (i_14_)) + ((!i_13_) & (sk[86]) & (!i_12_) & (g122) & (!i_14_)) + ((!i_13_) & (sk[86]) & (!i_12_) & (g122) & (i_14_)) + ((!i_13_) & (sk[86]) & (i_12_) & (!g122) & (!i_14_)) + ((!i_13_) & (sk[86]) & (i_12_) & (g122) & (!i_14_)) + ((!i_13_) & (sk[86]) & (i_12_) & (g122) & (i_14_)) + ((i_13_) & (!sk[86]) & (!i_12_) & (g122) & (!i_14_)) + ((i_13_) & (!sk[86]) & (!i_12_) & (g122) & (i_14_)) + ((i_13_) & (!sk[86]) & (i_12_) & (!g122) & (!i_14_)) + ((i_13_) & (!sk[86]) & (i_12_) & (!g122) & (i_14_)) + ((i_13_) & (!sk[86]) & (i_12_) & (g122) & (!i_14_)) + ((i_13_) & (!sk[86]) & (i_12_) & (g122) & (i_14_)) + ((i_13_) & (sk[86]) & (!i_12_) & (g122) & (!i_14_)) + ((i_13_) & (sk[86]) & (!i_12_) & (g122) & (i_14_)) + ((i_13_) & (sk[86]) & (i_12_) & (!g122) & (!i_14_)) + ((i_13_) & (sk[86]) & (i_12_) & (!g122) & (i_14_)) + ((i_13_) & (sk[86]) & (i_12_) & (g122) & (!i_14_)) + ((i_13_) & (sk[86]) & (i_12_) & (g122) & (i_14_)));
	assign g1605 = (((!sk[87]) & (!i_13_) & (!i_12_) & (g136) & (i_14_)) + ((!sk[87]) & (!i_13_) & (i_12_) & (!g136) & (!i_14_)) + ((!sk[87]) & (!i_13_) & (i_12_) & (!g136) & (i_14_)) + ((!sk[87]) & (!i_13_) & (i_12_) & (g136) & (!i_14_)) + ((!sk[87]) & (!i_13_) & (i_12_) & (g136) & (i_14_)) + ((!sk[87]) & (i_13_) & (!i_12_) & (g136) & (!i_14_)) + ((!sk[87]) & (i_13_) & (!i_12_) & (g136) & (i_14_)) + ((!sk[87]) & (i_13_) & (i_12_) & (!g136) & (!i_14_)) + ((!sk[87]) & (i_13_) & (i_12_) & (!g136) & (i_14_)) + ((!sk[87]) & (i_13_) & (i_12_) & (g136) & (!i_14_)) + ((!sk[87]) & (i_13_) & (i_12_) & (g136) & (i_14_)) + ((sk[87]) & (!i_13_) & (!i_12_) & (!g136) & (!i_14_)) + ((sk[87]) & (!i_13_) & (!i_12_) & (!g136) & (i_14_)) + ((sk[87]) & (!i_13_) & (!i_12_) & (g136) & (!i_14_)) + ((sk[87]) & (!i_13_) & (!i_12_) & (g136) & (i_14_)) + ((sk[87]) & (!i_13_) & (i_12_) & (!g136) & (!i_14_)) + ((sk[87]) & (!i_13_) & (i_12_) & (!g136) & (i_14_)) + ((sk[87]) & (!i_13_) & (i_12_) & (g136) & (!i_14_)) + ((sk[87]) & (i_13_) & (!i_12_) & (!g136) & (!i_14_)) + ((sk[87]) & (i_13_) & (!i_12_) & (!g136) & (i_14_)) + ((sk[87]) & (i_13_) & (!i_12_) & (g136) & (!i_14_)) + ((sk[87]) & (i_13_) & (!i_12_) & (g136) & (i_14_)) + ((sk[87]) & (i_13_) & (i_12_) & (!g136) & (!i_14_)) + ((sk[87]) & (i_13_) & (i_12_) & (!g136) & (i_14_)) + ((sk[87]) & (i_13_) & (i_12_) & (g136) & (!i_14_)) + ((sk[87]) & (i_13_) & (i_12_) & (g136) & (i_14_)));
	assign g1606 = (((!sk[88]) & (!i_13_) & (!i_12_) & (g122) & (i_14_)) + ((!sk[88]) & (!i_13_) & (i_12_) & (!g122) & (!i_14_)) + ((!sk[88]) & (!i_13_) & (i_12_) & (!g122) & (i_14_)) + ((!sk[88]) & (!i_13_) & (i_12_) & (g122) & (!i_14_)) + ((!sk[88]) & (!i_13_) & (i_12_) & (g122) & (i_14_)) + ((!sk[88]) & (i_13_) & (!i_12_) & (g122) & (!i_14_)) + ((!sk[88]) & (i_13_) & (!i_12_) & (g122) & (i_14_)) + ((!sk[88]) & (i_13_) & (i_12_) & (!g122) & (!i_14_)) + ((!sk[88]) & (i_13_) & (i_12_) & (!g122) & (i_14_)) + ((!sk[88]) & (i_13_) & (i_12_) & (g122) & (!i_14_)) + ((!sk[88]) & (i_13_) & (i_12_) & (g122) & (i_14_)) + ((sk[88]) & (!i_13_) & (!i_12_) & (!g122) & (i_14_)) + ((sk[88]) & (!i_13_) & (!i_12_) & (g122) & (!i_14_)) + ((sk[88]) & (!i_13_) & (!i_12_) & (g122) & (i_14_)) + ((sk[88]) & (i_13_) & (!i_12_) & (g122) & (i_14_)) + ((sk[88]) & (i_13_) & (i_12_) & (!g122) & (!i_14_)) + ((sk[88]) & (i_13_) & (i_12_) & (!g122) & (i_14_)) + ((sk[88]) & (i_13_) & (i_12_) & (g122) & (!i_14_)) + ((sk[88]) & (i_13_) & (i_12_) & (g122) & (i_14_)));
	assign g1607 = (((!g1608) & (sk[89]) & (!g1609)) + ((g1608) & (!sk[89]) & (!g1609)) + ((g1608) & (!sk[89]) & (g1609)));
	assign g1608 = (((!g149) & (sk[90]) & (g1610)) + ((g149) & (!sk[90]) & (!g1610)) + ((g149) & (!sk[90]) & (g1610)));
	assign g1609 = (((g149) & (!sk[91]) & (!g1613)) + ((g149) & (!sk[91]) & (g1613)) + ((g149) & (sk[91]) & (g1613)));
	assign g1610 = (((!sk[92]) & (g1611) & (!g1612)) + ((!sk[92]) & (g1611) & (g1612)) + ((sk[92]) & (!g1611) & (!g1612)));
	assign g1611 = (((!g201) & (sk[93]) & (g1614)) + ((g201) & (!sk[93]) & (!g1614)) + ((g201) & (!sk[93]) & (g1614)));
	assign g1612 = (((g201) & (!sk[94]) & (!g452)) + ((g201) & (!sk[94]) & (g452)) + ((g201) & (sk[94]) & (g452)));
	assign g1613 = (((!sk[95]) & (g201) & (!g1615)) + ((!sk[95]) & (g201) & (g1615)) + ((sk[95]) & (g201) & (g1615)));
	assign g1614 = (((!sk[96]) & (g452) & (!g338)) + ((!sk[96]) & (g452) & (g338)) + ((sk[96]) & (g452) & (g338)));
	assign g1615 = (((!sk[97]) & (!g1096) & (!g452) & (g206) & (g127)) + ((!sk[97]) & (!g1096) & (g452) & (!g206) & (!g127)) + ((!sk[97]) & (!g1096) & (g452) & (!g206) & (g127)) + ((!sk[97]) & (!g1096) & (g452) & (g206) & (!g127)) + ((!sk[97]) & (!g1096) & (g452) & (g206) & (g127)) + ((!sk[97]) & (g1096) & (!g452) & (g206) & (!g127)) + ((!sk[97]) & (g1096) & (!g452) & (g206) & (g127)) + ((!sk[97]) & (g1096) & (g452) & (!g206) & (!g127)) + ((!sk[97]) & (g1096) & (g452) & (!g206) & (g127)) + ((!sk[97]) & (g1096) & (g452) & (g206) & (!g127)) + ((!sk[97]) & (g1096) & (g452) & (g206) & (g127)) + ((sk[97]) & (g1096) & (g452) & (g206) & (g127)));
	assign g1616 = (((g1116) & (!sk[98]) & (!g1617)) + ((g1116) & (!sk[98]) & (g1617)) + ((g1116) & (sk[98]) & (g1617)));
	assign g1617 = (((!g1618) & (sk[99]) & (!g1619)) + ((g1618) & (!sk[99]) & (!g1619)) + ((g1618) & (!sk[99]) & (g1619)));
	assign g1618 = (((!sk[100]) & (i_8_) & (!g1620)) + ((!sk[100]) & (i_8_) & (g1620)) + ((sk[100]) & (!i_8_) & (g1620)));
	assign g1619 = (((i_8_) & (!sk[101]) & (!g1621)) + ((i_8_) & (!sk[101]) & (g1621)) + ((i_8_) & (sk[101]) & (g1621)));
	assign g1620 = (((!g88) & (sk[102]) & (!g1117) & (g1118)) + ((!g88) & (sk[102]) & (g1117) & (g1118)) + ((g88) & (!sk[102]) & (!g1117) & (!g1118)) + ((g88) & (!sk[102]) & (!g1117) & (g1118)) + ((g88) & (!sk[102]) & (g1117) & (!g1118)) + ((g88) & (!sk[102]) & (g1117) & (g1118)) + ((g88) & (sk[102]) & (!g1117) & (g1118)));
	assign g1621 = (((!sk[103]) & (!g696) & (!g88) & (g185) & (g1118)) + ((!sk[103]) & (!g696) & (g88) & (!g185) & (!g1118)) + ((!sk[103]) & (!g696) & (g88) & (!g185) & (g1118)) + ((!sk[103]) & (!g696) & (g88) & (g185) & (!g1118)) + ((!sk[103]) & (!g696) & (g88) & (g185) & (g1118)) + ((!sk[103]) & (g696) & (!g88) & (g185) & (!g1118)) + ((!sk[103]) & (g696) & (!g88) & (g185) & (g1118)) + ((!sk[103]) & (g696) & (g88) & (!g185) & (!g1118)) + ((!sk[103]) & (g696) & (g88) & (!g185) & (g1118)) + ((!sk[103]) & (g696) & (g88) & (g185) & (!g1118)) + ((!sk[103]) & (g696) & (g88) & (g185) & (g1118)) + ((sk[103]) & (!g696) & (!g88) & (!g185) & (g1118)) + ((sk[103]) & (!g696) & (!g88) & (g185) & (g1118)) + ((sk[103]) & (g696) & (!g88) & (!g185) & (g1118)) + ((sk[103]) & (g696) & (!g88) & (g185) & (g1118)) + ((sk[103]) & (g696) & (g88) & (g185) & (g1118)));
	assign g1622 = (((g1102) & (!sk[104]) & (!g1623)) + ((g1102) & (!sk[104]) & (g1623)) + ((g1102) & (sk[104]) & (g1623)));
	assign g1623 = (((!g1624) & (sk[105]) & (!g1625)) + ((g1624) & (!sk[105]) & (!g1625)) + ((g1624) & (!sk[105]) & (g1625)));
	assign g1624 = (((!i_8_) & (sk[106]) & (g1626)) + ((i_8_) & (!sk[106]) & (!g1626)) + ((i_8_) & (!sk[106]) & (g1626)));
	assign g1625 = (((i_8_) & (!sk[107]) & (!g1627)) + ((i_8_) & (!sk[107]) & (g1627)) + ((i_8_) & (sk[107]) & (g1627)));
	assign g1626 = (((!g8) & (sk[108]) & (!g88)) + ((g8) & (!sk[108]) & (!g88)) + ((g8) & (!sk[108]) & (g88)) + ((g8) & (sk[108]) & (!g88)) + ((g8) & (sk[108]) & (g88)));
	assign g1627 = (((!g92) & (!g221) & (!sk[109]) & (g231) & (g88)) + ((!g92) & (!g221) & (sk[109]) & (!g231) & (!g88)) + ((!g92) & (!g221) & (sk[109]) & (g231) & (!g88)) + ((!g92) & (g221) & (!sk[109]) & (!g231) & (!g88)) + ((!g92) & (g221) & (!sk[109]) & (!g231) & (g88)) + ((!g92) & (g221) & (!sk[109]) & (g231) & (!g88)) + ((!g92) & (g221) & (!sk[109]) & (g231) & (g88)) + ((!g92) & (g221) & (sk[109]) & (!g231) & (!g88)) + ((!g92) & (g221) & (sk[109]) & (g231) & (!g88)) + ((g92) & (!g221) & (!sk[109]) & (g231) & (!g88)) + ((g92) & (!g221) & (!sk[109]) & (g231) & (g88)) + ((g92) & (!g221) & (sk[109]) & (!g231) & (!g88)) + ((g92) & (!g221) & (sk[109]) & (g231) & (!g88)) + ((g92) & (g221) & (!sk[109]) & (!g231) & (!g88)) + ((g92) & (g221) & (!sk[109]) & (!g231) & (g88)) + ((g92) & (g221) & (!sk[109]) & (g231) & (!g88)) + ((g92) & (g221) & (!sk[109]) & (g231) & (g88)) + ((g92) & (g221) & (sk[109]) & (!g231) & (!g88)) + ((g92) & (g221) & (sk[109]) & (g231) & (!g88)) + ((g92) & (g221) & (sk[109]) & (g231) & (g88)));
	assign g1628 = (((!sk[110]) & (g1629) & (!g1630)) + ((!sk[110]) & (g1629) & (g1630)) + ((sk[110]) & (!g1629) & (!g1630)));
	assign g1629 = (((!g90) & (sk[111]) & (g1631)) + ((g90) & (!sk[111]) & (!g1631)) + ((g90) & (!sk[111]) & (g1631)));
	assign g1630 = (((g90) & (!sk[112]) & (!g1634)) + ((g90) & (!sk[112]) & (g1634)) + ((g90) & (sk[112]) & (g1634)));
	assign g1631 = (((!g1632) & (sk[113]) & (!g1633)) + ((g1632) & (!sk[113]) & (!g1633)) + ((g1632) & (!sk[113]) & (g1633)));
	assign g1632 = (((!i_8_) & (sk[114]) & (!g88)) + ((i_8_) & (!sk[114]) & (!g88)) + ((i_8_) & (!sk[114]) & (g88)));
	assign g1633 = (((i_8_) & (!sk[115]) & (!g1637)) + ((i_8_) & (!sk[115]) & (g1637)) + ((i_8_) & (sk[115]) & (g1637)));
	assign g1634 = (((!sk[116]) & (g1635) & (!g1636)) + ((!sk[116]) & (g1635) & (g1636)) + ((sk[116]) & (!g1635) & (!g1636)));
	assign g1635 = (((!i_8_) & (sk[117]) & (g1638)) + ((i_8_) & (!sk[117]) & (!g1638)) + ((i_8_) & (!sk[117]) & (g1638)));
	assign g1636 = (((!sk[118]) & (i_8_) & (!g1639)) + ((!sk[118]) & (i_8_) & (g1639)) + ((sk[118]) & (i_8_) & (g1639)));
	assign g1637 = (((!g467) & (sk[119]) & (!g528) & (!g88)) + ((!g467) & (sk[119]) & (g528) & (!g88)) + ((g467) & (!sk[119]) & (!g528) & (!g88)) + ((g467) & (!sk[119]) & (!g528) & (g88)) + ((g467) & (!sk[119]) & (g528) & (!g88)) + ((g467) & (!sk[119]) & (g528) & (g88)) + ((g467) & (sk[119]) & (!g528) & (!g88)) + ((g467) & (sk[119]) & (g528) & (!g88)) + ((g467) & (sk[119]) & (g528) & (g88)));
	assign g1638 = (((!g468) & (!g467) & (!sk[120]) & (g92) & (g88)) + ((!g468) & (!g467) & (sk[120]) & (!g92) & (!g88)) + ((!g468) & (!g467) & (sk[120]) & (g92) & (!g88)) + ((!g468) & (g467) & (!sk[120]) & (!g92) & (!g88)) + ((!g468) & (g467) & (!sk[120]) & (!g92) & (g88)) + ((!g468) & (g467) & (!sk[120]) & (g92) & (!g88)) + ((!g468) & (g467) & (!sk[120]) & (g92) & (g88)) + ((!g468) & (g467) & (sk[120]) & (!g92) & (!g88)) + ((!g468) & (g467) & (sk[120]) & (g92) & (!g88)) + ((g468) & (!g467) & (!sk[120]) & (g92) & (!g88)) + ((g468) & (!g467) & (!sk[120]) & (g92) & (g88)) + ((g468) & (!g467) & (sk[120]) & (!g92) & (!g88)) + ((g468) & (!g467) & (sk[120]) & (g92) & (!g88)) + ((g468) & (g467) & (!sk[120]) & (!g92) & (!g88)) + ((g468) & (g467) & (!sk[120]) & (!g92) & (g88)) + ((g468) & (g467) & (!sk[120]) & (g92) & (!g88)) + ((g468) & (g467) & (!sk[120]) & (g92) & (g88)) + ((g468) & (g467) & (sk[120]) & (!g92) & (!g88)) + ((g468) & (g467) & (sk[120]) & (g92) & (!g88)) + ((g468) & (g467) & (sk[120]) & (g92) & (g88)));
	assign g1639 = (((!sk[121]) & (g467) & (!g528) & (!g88)) + ((!sk[121]) & (g467) & (!g528) & (g88)) + ((!sk[121]) & (g467) & (g528) & (!g88)) + ((!sk[121]) & (g467) & (g528) & (g88)) + ((sk[121]) & (!g467) & (!g528) & (!g88)) + ((sk[121]) & (!g467) & (g528) & (!g88)) + ((sk[121]) & (g467) & (!g528) & (!g88)) + ((sk[121]) & (g467) & (g528) & (!g88)) + ((sk[121]) & (g467) & (g528) & (g88)));
	assign g1640 = (((!sk[122]) & (g1641) & (!g1642)) + ((!sk[122]) & (g1641) & (g1642)) + ((sk[122]) & (!g1641) & (!g1642)));
	assign g1641 = (((!g1031) & (sk[123]) & (g1643)) + ((g1031) & (!sk[123]) & (!g1643)) + ((g1031) & (!sk[123]) & (g1643)));
	assign g1642 = (((!sk[124]) & (g1031) & (!g1646)) + ((!sk[124]) & (g1031) & (g1646)) + ((sk[124]) & (g1031) & (g1646)));
	assign g1643 = (((!g1644) & (sk[125]) & (!g1645)) + ((g1644) & (!sk[125]) & (!g1645)) + ((g1644) & (!sk[125]) & (g1645)));
	assign g1644 = (((!sk[126]) & (i_8_) & (!g1649)) + ((!sk[126]) & (i_8_) & (g1649)) + ((sk[126]) & (!i_8_) & (g1649)));
	assign g1645 = (((i_8_) & (!sk[127]) & (!g1650)) + ((i_8_) & (!sk[127]) & (g1650)) + ((i_8_) & (sk[127]) & (g1650)));
	assign g1646 = (((!sk[0]) & (g1647) & (!g1648)) + ((!sk[0]) & (g1647) & (g1648)) + ((sk[0]) & (!g1647) & (!g1648)));
	assign g1647 = (((!i_8_) & (sk[1]) & (g1651)) + ((i_8_) & (!sk[1]) & (!g1651)) + ((i_8_) & (!sk[1]) & (g1651)));
	assign g1648 = (((i_8_) & (!sk[2]) & (!g1652)) + ((i_8_) & (!sk[2]) & (g1652)) + ((i_8_) & (sk[2]) & (g1652)));
	assign g1649 = (((!g400) & (!i_7_) & (sk[3]) & (g1038)) + ((!g400) & (i_7_) & (sk[3]) & (g1038)) + ((g400) & (!i_7_) & (!sk[3]) & (!g1038)) + ((g400) & (!i_7_) & (!sk[3]) & (g1038)) + ((g400) & (!i_7_) & (sk[3]) & (g1038)) + ((g400) & (i_7_) & (!sk[3]) & (!g1038)) + ((g400) & (i_7_) & (!sk[3]) & (g1038)));
	assign g1650 = (((!g400) & (!sk[4]) & (!i_7_) & (g1032) & (g1038)) + ((!g400) & (!sk[4]) & (i_7_) & (!g1032) & (!g1038)) + ((!g400) & (!sk[4]) & (i_7_) & (!g1032) & (g1038)) + ((!g400) & (!sk[4]) & (i_7_) & (g1032) & (!g1038)) + ((!g400) & (!sk[4]) & (i_7_) & (g1032) & (g1038)) + ((!g400) & (sk[4]) & (!i_7_) & (!g1032) & (g1038)) + ((!g400) & (sk[4]) & (!i_7_) & (g1032) & (g1038)) + ((!g400) & (sk[4]) & (i_7_) & (!g1032) & (g1038)) + ((!g400) & (sk[4]) & (i_7_) & (g1032) & (g1038)) + ((g400) & (!sk[4]) & (!i_7_) & (g1032) & (!g1038)) + ((g400) & (!sk[4]) & (!i_7_) & (g1032) & (g1038)) + ((g400) & (!sk[4]) & (i_7_) & (!g1032) & (!g1038)) + ((g400) & (!sk[4]) & (i_7_) & (!g1032) & (g1038)) + ((g400) & (!sk[4]) & (i_7_) & (g1032) & (!g1038)) + ((g400) & (!sk[4]) & (i_7_) & (g1032) & (g1038)) + ((g400) & (sk[4]) & (!i_7_) & (!g1032) & (g1038)) + ((g400) & (sk[4]) & (!i_7_) & (g1032) & (g1038)) + ((g400) & (sk[4]) & (i_7_) & (g1032) & (g1038)));
	assign g1651 = (((!sk[5]) & (!g400) & (!i_7_) & (g20) & (g1038)) + ((!sk[5]) & (!g400) & (i_7_) & (!g20) & (!g1038)) + ((!sk[5]) & (!g400) & (i_7_) & (!g20) & (g1038)) + ((!sk[5]) & (!g400) & (i_7_) & (g20) & (!g1038)) + ((!sk[5]) & (!g400) & (i_7_) & (g20) & (g1038)) + ((!sk[5]) & (g400) & (!i_7_) & (g20) & (!g1038)) + ((!sk[5]) & (g400) & (!i_7_) & (g20) & (g1038)) + ((!sk[5]) & (g400) & (i_7_) & (!g20) & (!g1038)) + ((!sk[5]) & (g400) & (i_7_) & (!g20) & (g1038)) + ((!sk[5]) & (g400) & (i_7_) & (g20) & (!g1038)) + ((!sk[5]) & (g400) & (i_7_) & (g20) & (g1038)) + ((sk[5]) & (!g400) & (!i_7_) & (!g20) & (g1038)) + ((sk[5]) & (!g400) & (!i_7_) & (g20) & (g1038)) + ((sk[5]) & (!g400) & (i_7_) & (!g20) & (g1038)) + ((sk[5]) & (!g400) & (i_7_) & (g20) & (g1038)) + ((sk[5]) & (g400) & (!i_7_) & (!g20) & (g1038)) + ((sk[5]) & (g400) & (!i_7_) & (g20) & (g1038)) + ((sk[5]) & (g400) & (i_7_) & (g20) & (g1038)));
	assign g1652 = (((!g400) & (!sk[6]) & (!i_7_) & (g1032) & (g1038)) + ((!g400) & (!sk[6]) & (i_7_) & (!g1032) & (!g1038)) + ((!g400) & (!sk[6]) & (i_7_) & (!g1032) & (g1038)) + ((!g400) & (!sk[6]) & (i_7_) & (g1032) & (!g1038)) + ((!g400) & (!sk[6]) & (i_7_) & (g1032) & (g1038)) + ((!g400) & (sk[6]) & (!i_7_) & (!g1032) & (g1038)) + ((!g400) & (sk[6]) & (!i_7_) & (g1032) & (g1038)) + ((!g400) & (sk[6]) & (i_7_) & (!g1032) & (g1038)) + ((!g400) & (sk[6]) & (i_7_) & (g1032) & (g1038)) + ((g400) & (!sk[6]) & (!i_7_) & (g1032) & (!g1038)) + ((g400) & (!sk[6]) & (!i_7_) & (g1032) & (g1038)) + ((g400) & (!sk[6]) & (i_7_) & (!g1032) & (!g1038)) + ((g400) & (!sk[6]) & (i_7_) & (!g1032) & (g1038)) + ((g400) & (!sk[6]) & (i_7_) & (g1032) & (!g1038)) + ((g400) & (!sk[6]) & (i_7_) & (g1032) & (g1038)) + ((g400) & (sk[6]) & (!i_7_) & (!g1032) & (g1038)) + ((g400) & (sk[6]) & (!i_7_) & (g1032) & (g1038)) + ((g400) & (sk[6]) & (i_7_) & (g1032) & (g1038)));
	assign g1653 = (((!g1654) & (sk[7]) & (!g1655)) + ((g1654) & (!sk[7]) & (!g1655)) + ((g1654) & (!sk[7]) & (g1655)));
	assign g1654 = (((!g118) & (sk[8]) & (g1656)) + ((g118) & (!sk[8]) & (!g1656)) + ((g118) & (!sk[8]) & (g1656)));
	assign g1655 = (((g118) & (!sk[9]) & (!g1659)) + ((g118) & (!sk[9]) & (g1659)) + ((g118) & (sk[9]) & (g1659)));
	assign g1656 = (((!g1657) & (sk[10]) & (!g1658)) + ((g1657) & (!sk[10]) & (!g1658)) + ((g1657) & (!sk[10]) & (g1658)));
	assign g1657 = (((!sk[11]) & (i_13_) & (!g1662)) + ((!sk[11]) & (i_13_) & (g1662)) + ((sk[11]) & (!i_13_) & (g1662)));
	assign g1658 = (((i_13_) & (!sk[12]) & (!g1663)) + ((i_13_) & (!sk[12]) & (g1663)) + ((i_13_) & (sk[12]) & (g1663)));
	assign g1659 = (((!g1660) & (sk[13]) & (!g1661)) + ((g1660) & (!sk[13]) & (!g1661)) + ((g1660) & (!sk[13]) & (g1661)));
	assign g1660 = (((!i_13_) & (sk[14]) & (g1664)) + ((i_13_) & (!sk[14]) & (!g1664)) + ((i_13_) & (!sk[14]) & (g1664)));
	assign g1661 = (((i_13_) & (!sk[15]) & (!g1665)) + ((i_13_) & (!sk[15]) & (g1665)) + ((i_13_) & (sk[15]) & (g1665)));
	assign g1662 = (((!i_12_) & (!i_14_) & (!sk[16]) & (g134) & (g102)) + ((!i_12_) & (!i_14_) & (sk[16]) & (!g134) & (!g102)) + ((!i_12_) & (!i_14_) & (sk[16]) & (!g134) & (g102)) + ((!i_12_) & (!i_14_) & (sk[16]) & (g134) & (!g102)) + ((!i_12_) & (!i_14_) & (sk[16]) & (g134) & (g102)) + ((!i_12_) & (i_14_) & (!sk[16]) & (!g134) & (!g102)) + ((!i_12_) & (i_14_) & (!sk[16]) & (!g134) & (g102)) + ((!i_12_) & (i_14_) & (!sk[16]) & (g134) & (!g102)) + ((!i_12_) & (i_14_) & (!sk[16]) & (g134) & (g102)) + ((!i_12_) & (i_14_) & (sk[16]) & (!g134) & (!g102)) + ((!i_12_) & (i_14_) & (sk[16]) & (!g134) & (g102)) + ((!i_12_) & (i_14_) & (sk[16]) & (g134) & (g102)) + ((i_12_) & (!i_14_) & (!sk[16]) & (g134) & (!g102)) + ((i_12_) & (!i_14_) & (!sk[16]) & (g134) & (g102)) + ((i_12_) & (!i_14_) & (sk[16]) & (!g134) & (!g102)) + ((i_12_) & (!i_14_) & (sk[16]) & (!g134) & (g102)) + ((i_12_) & (!i_14_) & (sk[16]) & (g134) & (!g102)) + ((i_12_) & (!i_14_) & (sk[16]) & (g134) & (g102)) + ((i_12_) & (i_14_) & (!sk[16]) & (!g134) & (!g102)) + ((i_12_) & (i_14_) & (!sk[16]) & (!g134) & (g102)) + ((i_12_) & (i_14_) & (!sk[16]) & (g134) & (!g102)) + ((i_12_) & (i_14_) & (!sk[16]) & (g134) & (g102)) + ((i_12_) & (i_14_) & (sk[16]) & (!g134) & (!g102)) + ((i_12_) & (i_14_) & (sk[16]) & (!g134) & (g102)) + ((i_12_) & (i_14_) & (sk[16]) & (g134) & (!g102)) + ((i_12_) & (i_14_) & (sk[16]) & (g134) & (g102)));
	assign g1663 = (((!i_12_) & (!i_14_) & (!g186) & (sk[17]) & (!g102)) + ((!i_12_) & (!i_14_) & (!g186) & (sk[17]) & (g102)) + ((!i_12_) & (!i_14_) & (g186) & (!sk[17]) & (g102)) + ((!i_12_) & (!i_14_) & (g186) & (sk[17]) & (g102)) + ((!i_12_) & (i_14_) & (!g186) & (!sk[17]) & (!g102)) + ((!i_12_) & (i_14_) & (!g186) & (!sk[17]) & (g102)) + ((!i_12_) & (i_14_) & (!g186) & (sk[17]) & (!g102)) + ((!i_12_) & (i_14_) & (!g186) & (sk[17]) & (g102)) + ((!i_12_) & (i_14_) & (g186) & (!sk[17]) & (!g102)) + ((!i_12_) & (i_14_) & (g186) & (!sk[17]) & (g102)) + ((!i_12_) & (i_14_) & (g186) & (sk[17]) & (!g102)) + ((!i_12_) & (i_14_) & (g186) & (sk[17]) & (g102)) + ((i_12_) & (!i_14_) & (!g186) & (sk[17]) & (!g102)) + ((i_12_) & (!i_14_) & (!g186) & (sk[17]) & (g102)) + ((i_12_) & (!i_14_) & (g186) & (!sk[17]) & (!g102)) + ((i_12_) & (!i_14_) & (g186) & (!sk[17]) & (g102)) + ((i_12_) & (!i_14_) & (g186) & (sk[17]) & (!g102)) + ((i_12_) & (!i_14_) & (g186) & (sk[17]) & (g102)) + ((i_12_) & (i_14_) & (!g186) & (!sk[17]) & (!g102)) + ((i_12_) & (i_14_) & (!g186) & (!sk[17]) & (g102)) + ((i_12_) & (i_14_) & (!g186) & (sk[17]) & (!g102)) + ((i_12_) & (i_14_) & (!g186) & (sk[17]) & (g102)) + ((i_12_) & (i_14_) & (g186) & (!sk[17]) & (!g102)) + ((i_12_) & (i_14_) & (g186) & (!sk[17]) & (g102)) + ((i_12_) & (i_14_) & (g186) & (sk[17]) & (!g102)) + ((i_12_) & (i_14_) & (g186) & (sk[17]) & (g102)));
	assign g1664 = (((!i_12_) & (!i_14_) & (sk[18]) & (!g102)) + ((!i_12_) & (!i_14_) & (sk[18]) & (g102)) + ((!i_12_) & (i_14_) & (sk[18]) & (g102)) + ((i_12_) & (!i_14_) & (!sk[18]) & (!g102)) + ((i_12_) & (!i_14_) & (!sk[18]) & (g102)) + ((i_12_) & (!i_14_) & (sk[18]) & (!g102)) + ((i_12_) & (!i_14_) & (sk[18]) & (g102)) + ((i_12_) & (i_14_) & (!sk[18]) & (!g102)) + ((i_12_) & (i_14_) & (!sk[18]) & (g102)) + ((i_12_) & (i_14_) & (sk[18]) & (!g102)) + ((i_12_) & (i_14_) & (sk[18]) & (g102)));
	assign g1665 = (((!i_12_) & (sk[19]) & (!i_14_) & (g102)) + ((!i_12_) & (sk[19]) & (i_14_) & (!g102)) + ((!i_12_) & (sk[19]) & (i_14_) & (g102)) + ((i_12_) & (!sk[19]) & (!i_14_) & (!g102)) + ((i_12_) & (!sk[19]) & (!i_14_) & (g102)) + ((i_12_) & (!sk[19]) & (i_14_) & (!g102)) + ((i_12_) & (!sk[19]) & (i_14_) & (g102)) + ((i_12_) & (sk[19]) & (!i_14_) & (!g102)) + ((i_12_) & (sk[19]) & (!i_14_) & (g102)) + ((i_12_) & (sk[19]) & (i_14_) & (!g102)) + ((i_12_) & (sk[19]) & (i_14_) & (g102)));
	assign g1666 = (((i_14_) & (!sk[20]) & (!g1667)) + ((i_14_) & (!sk[20]) & (g1667)) + ((i_14_) & (sk[20]) & (!g1667)));
	assign g1667 = (((!sk[21]) & (i_14_) & (!g1668)) + ((!sk[21]) & (i_14_) & (g1668)) + ((sk[21]) & (i_14_) & (g1668)));
	assign g1668 = (((!g1669) & (sk[22]) & (!g1670)) + ((g1669) & (!sk[22]) & (!g1670)) + ((g1669) & (!sk[22]) & (g1670)));
	assign g1669 = (((!i_13_) & (sk[23]) & (g1671)) + ((i_13_) & (!sk[23]) & (!g1671)) + ((i_13_) & (!sk[23]) & (g1671)));
	assign g1670 = (((!sk[24]) & (i_13_) & (!g1672)) + ((!sk[24]) & (i_13_) & (g1672)) + ((sk[24]) & (i_13_) & (g1672)));
	assign g1671 = (((!g495) & (!sk[25]) & (!i_12_) & (g186) & (g15)) + ((!g495) & (!sk[25]) & (i_12_) & (!g186) & (!g15)) + ((!g495) & (!sk[25]) & (i_12_) & (!g186) & (g15)) + ((!g495) & (!sk[25]) & (i_12_) & (g186) & (!g15)) + ((!g495) & (!sk[25]) & (i_12_) & (g186) & (g15)) + ((!g495) & (sk[25]) & (!i_12_) & (!g186) & (!g15)) + ((!g495) & (sk[25]) & (!i_12_) & (!g186) & (g15)) + ((!g495) & (sk[25]) & (!i_12_) & (g186) & (!g15)) + ((!g495) & (sk[25]) & (!i_12_) & (g186) & (g15)) + ((!g495) & (sk[25]) & (i_12_) & (!g186) & (!g15)) + ((!g495) & (sk[25]) & (i_12_) & (!g186) & (g15)) + ((!g495) & (sk[25]) & (i_12_) & (g186) & (g15)) + ((g495) & (!sk[25]) & (!i_12_) & (g186) & (!g15)) + ((g495) & (!sk[25]) & (!i_12_) & (g186) & (g15)) + ((g495) & (!sk[25]) & (i_12_) & (!g186) & (!g15)) + ((g495) & (!sk[25]) & (i_12_) & (!g186) & (g15)) + ((g495) & (!sk[25]) & (i_12_) & (g186) & (!g15)) + ((g495) & (!sk[25]) & (i_12_) & (g186) & (g15)) + ((g495) & (sk[25]) & (!i_12_) & (!g186) & (!g15)) + ((g495) & (sk[25]) & (!i_12_) & (!g186) & (g15)) + ((g495) & (sk[25]) & (!i_12_) & (g186) & (!g15)) + ((g495) & (sk[25]) & (!i_12_) & (g186) & (g15)) + ((g495) & (sk[25]) & (i_12_) & (!g186) & (g15)) + ((g495) & (sk[25]) & (i_12_) & (g186) & (g15)));
	assign g1672 = (((!sk[26]) & (i_12_) & (!g135) & (!g15)) + ((!sk[26]) & (i_12_) & (!g135) & (g15)) + ((!sk[26]) & (i_12_) & (g135) & (!g15)) + ((!sk[26]) & (i_12_) & (g135) & (g15)) + ((sk[26]) & (!i_12_) & (!g135) & (!g15)) + ((sk[26]) & (!i_12_) & (!g135) & (g15)) + ((sk[26]) & (!i_12_) & (g135) & (!g15)) + ((sk[26]) & (!i_12_) & (g135) & (g15)) + ((sk[26]) & (i_12_) & (!g135) & (!g15)) + ((sk[26]) & (i_12_) & (!g135) & (g15)) + ((sk[26]) & (i_12_) & (g135) & (g15)));
	assign g1673 = (((!g1674) & (sk[27]) & (!g1675)) + ((g1674) & (!sk[27]) & (!g1675)) + ((g1674) & (!sk[27]) & (g1675)));
	assign g1674 = (((!sk[28]) & (g807) & (!g1676)) + ((!sk[28]) & (g807) & (g1676)) + ((sk[28]) & (!g807) & (g1676)));
	assign g1675 = (((g807) & (!sk[29]) & (!g1679)) + ((g807) & (!sk[29]) & (g1679)) + ((g807) & (sk[29]) & (g1679)));
	assign g1676 = (((!g1677) & (sk[30]) & (!g1678)) + ((g1677) & (!sk[30]) & (!g1678)) + ((g1677) & (!sk[30]) & (g1678)));
	assign g1677 = (((!sk[31]) & (i_8_) & (!g1682)) + ((!sk[31]) & (i_8_) & (g1682)) + ((sk[31]) & (!i_8_) & (g1682)));
	assign g1678 = (((i_8_) & (!sk[32]) & (!g1683)) + ((i_8_) & (!sk[32]) & (g1683)) + ((i_8_) & (sk[32]) & (g1683)));
	assign g1679 = (((!g1680) & (sk[33]) & (!g1681)) + ((g1680) & (!sk[33]) & (!g1681)) + ((g1680) & (!sk[33]) & (g1681)));
	assign g1680 = (((!sk[34]) & (i_8_) & (!g1684)) + ((!sk[34]) & (i_8_) & (g1684)) + ((sk[34]) & (!i_8_) & (g1684)));
	assign g1681 = (((i_8_) & (!sk[35]) & (!g1685)) + ((i_8_) & (!sk[35]) & (g1685)) + ((i_8_) & (sk[35]) & (g1685)));
	assign g1682 = (((!g30) & (sk[36]) & (!g87)) + ((!g30) & (sk[36]) & (g87)) + ((g30) & (!sk[36]) & (!g87)) + ((g30) & (!sk[36]) & (g87)) + ((g30) & (sk[36]) & (!g87)));
	assign g1683 = (((!g30) & (sk[37]) & (!g16) & (!g87)) + ((!g30) & (sk[37]) & (!g16) & (g87)) + ((!g30) & (sk[37]) & (g16) & (!g87)) + ((!g30) & (sk[37]) & (g16) & (g87)) + ((g30) & (!sk[37]) & (!g16) & (!g87)) + ((g30) & (!sk[37]) & (!g16) & (g87)) + ((g30) & (!sk[37]) & (g16) & (!g87)) + ((g30) & (!sk[37]) & (g16) & (g87)) + ((g30) & (sk[37]) & (!g16) & (!g87)) + ((g30) & (sk[37]) & (g16) & (!g87)) + ((g30) & (sk[37]) & (g16) & (g87)));
	assign g1684 = (((!g30) & (!g464) & (!sk[38]) & (g226) & (g87)) + ((!g30) & (!g464) & (sk[38]) & (!g226) & (!g87)) + ((!g30) & (!g464) & (sk[38]) & (!g226) & (g87)) + ((!g30) & (!g464) & (sk[38]) & (g226) & (!g87)) + ((!g30) & (!g464) & (sk[38]) & (g226) & (g87)) + ((!g30) & (g464) & (!sk[38]) & (!g226) & (!g87)) + ((!g30) & (g464) & (!sk[38]) & (!g226) & (g87)) + ((!g30) & (g464) & (!sk[38]) & (g226) & (!g87)) + ((!g30) & (g464) & (!sk[38]) & (g226) & (g87)) + ((!g30) & (g464) & (sk[38]) & (!g226) & (!g87)) + ((!g30) & (g464) & (sk[38]) & (!g226) & (g87)) + ((!g30) & (g464) & (sk[38]) & (g226) & (!g87)) + ((!g30) & (g464) & (sk[38]) & (g226) & (g87)) + ((g30) & (!g464) & (!sk[38]) & (g226) & (!g87)) + ((g30) & (!g464) & (!sk[38]) & (g226) & (g87)) + ((g30) & (!g464) & (sk[38]) & (!g226) & (!g87)) + ((g30) & (!g464) & (sk[38]) & (g226) & (!g87)) + ((g30) & (g464) & (!sk[38]) & (!g226) & (!g87)) + ((g30) & (g464) & (!sk[38]) & (!g226) & (g87)) + ((g30) & (g464) & (!sk[38]) & (g226) & (!g87)) + ((g30) & (g464) & (!sk[38]) & (g226) & (g87)) + ((g30) & (g464) & (sk[38]) & (!g226) & (!g87)) + ((g30) & (g464) & (sk[38]) & (g226) & (!g87)) + ((g30) & (g464) & (sk[38]) & (g226) & (g87)));
	assign g1685 = (((!g30) & (sk[39]) & (!g16) & (!g87)) + ((!g30) & (sk[39]) & (!g16) & (g87)) + ((!g30) & (sk[39]) & (g16) & (!g87)) + ((!g30) & (sk[39]) & (g16) & (g87)) + ((g30) & (!sk[39]) & (!g16) & (!g87)) + ((g30) & (!sk[39]) & (!g16) & (g87)) + ((g30) & (!sk[39]) & (g16) & (!g87)) + ((g30) & (!sk[39]) & (g16) & (g87)) + ((g30) & (sk[39]) & (!g16) & (!g87)) + ((g30) & (sk[39]) & (g16) & (!g87)) + ((g30) & (sk[39]) & (g16) & (g87)));
	assign g1686 = (((!sk[40]) & (g1687) & (!g1688)) + ((!sk[40]) & (g1687) & (g1688)) + ((sk[40]) & (!g1687) & (!g1688)));
	assign g1687 = (((!sk[41]) & (i_6_) & (!g1689)) + ((!sk[41]) & (i_6_) & (g1689)) + ((sk[41]) & (!i_6_) & (g1689)));
	assign g1688 = (((i_6_) & (!sk[42]) & (!g1691)) + ((i_6_) & (!sk[42]) & (g1691)) + ((i_6_) & (sk[42]) & (g1691)));
	assign g1689 = (((!i_7_) & (sk[43]) & (!g1690)) + ((i_7_) & (!sk[43]) & (!g1690)) + ((i_7_) & (!sk[43]) & (g1690)));
	assign g1690 = (((!sk[44]) & (i_7_) & (!g1693)) + ((!sk[44]) & (i_7_) & (g1693)) + ((sk[44]) & (!i_7_) & (g1693)));
	assign g1691 = (((i_7_) & (!sk[45]) & (!g1692)) + ((i_7_) & (!sk[45]) & (g1692)) + ((i_7_) & (sk[45]) & (!g1692)));
	assign g1692 = (((i_7_) & (!sk[46]) & (!g1694)) + ((i_7_) & (!sk[46]) & (g1694)) + ((i_7_) & (sk[46]) & (g1694)));
	assign g1693 = (((!sk[47]) & (g87) & (!g615) & (!g528)) + ((!sk[47]) & (g87) & (!g615) & (g528)) + ((!sk[47]) & (g87) & (g615) & (!g528)) + ((!sk[47]) & (g87) & (g615) & (g528)) + ((sk[47]) & (!g87) & (!g615) & (!g528)) + ((sk[47]) & (!g87) & (!g615) & (g528)) + ((sk[47]) & (!g87) & (g615) & (!g528)) + ((sk[47]) & (!g87) & (g615) & (g528)) + ((sk[47]) & (g87) & (g615) & (g528)));
	assign g1694 = (((!g98) & (sk[48]) & (!g616)) + ((!g98) & (sk[48]) & (g616)) + ((g98) & (!sk[48]) & (!g616)) + ((g98) & (!sk[48]) & (g616)) + ((g98) & (sk[48]) & (g616)));
	assign g1695 = (((!g1696) & (sk[49]) & (!g1697)) + ((g1696) & (!sk[49]) & (!g1697)) + ((g1696) & (!sk[49]) & (g1697)));
	assign g1696 = (((!sk[50]) & (g100) & (!g1698)) + ((!sk[50]) & (g100) & (g1698)) + ((sk[50]) & (!g100) & (g1698)));
	assign g1697 = (((g100) & (!sk[51]) & (!g1701)) + ((g100) & (!sk[51]) & (g1701)) + ((g100) & (sk[51]) & (g1701)));
	assign g1698 = (((!g1699) & (sk[52]) & (!g1700)) + ((g1699) & (!sk[52]) & (!g1700)) + ((g1699) & (!sk[52]) & (g1700)));
	assign g1699 = (((!i_8_) & (sk[53]) & (g1704)) + ((i_8_) & (!sk[53]) & (!g1704)) + ((i_8_) & (!sk[53]) & (g1704)));
	assign g1700 = (((!sk[54]) & (i_8_) & (!g1705)) + ((!sk[54]) & (i_8_) & (g1705)) + ((sk[54]) & (i_8_) & (g1705)));
	assign g1701 = (((!sk[55]) & (g1702) & (!g1703)) + ((!sk[55]) & (g1702) & (g1703)) + ((sk[55]) & (!g1702) & (!g1703)));
	assign g1702 = (((!sk[56]) & (i_8_) & (!g1706)) + ((!sk[56]) & (i_8_) & (g1706)) + ((sk[56]) & (!i_8_) & (g1706)));
	assign g1703 = (((!sk[57]) & (i_8_) & (!g1707)) + ((!sk[57]) & (i_8_) & (g1707)) + ((sk[57]) & (i_8_) & (g1707)));
	assign g1704 = (((!g592) & (sk[58]) & (!g590) & (g251)) + ((g592) & (!sk[58]) & (!g590) & (!g251)) + ((g592) & (!sk[58]) & (!g590) & (g251)) + ((g592) & (!sk[58]) & (g590) & (!g251)) + ((g592) & (!sk[58]) & (g590) & (g251)) + ((g592) & (sk[58]) & (!g590) & (g251)) + ((g592) & (sk[58]) & (g590) & (g251)));
	assign g1705 = (((!g592) & (!g590) & (sk[59]) & (g251)) + ((g592) & (!g590) & (!sk[59]) & (!g251)) + ((g592) & (!g590) & (!sk[59]) & (g251)) + ((g592) & (!g590) & (sk[59]) & (g251)) + ((g592) & (g590) & (!sk[59]) & (!g251)) + ((g592) & (g590) & (!sk[59]) & (g251)) + ((g592) & (g590) & (sk[59]) & (g251)));
	assign g1706 = (((!sk[60]) & (!g592) & (!g590) & (g547) & (g251)) + ((!sk[60]) & (!g592) & (g590) & (!g547) & (!g251)) + ((!sk[60]) & (!g592) & (g590) & (!g547) & (g251)) + ((!sk[60]) & (!g592) & (g590) & (g547) & (!g251)) + ((!sk[60]) & (!g592) & (g590) & (g547) & (g251)) + ((!sk[60]) & (g592) & (!g590) & (g547) & (!g251)) + ((!sk[60]) & (g592) & (!g590) & (g547) & (g251)) + ((!sk[60]) & (g592) & (g590) & (!g547) & (!g251)) + ((!sk[60]) & (g592) & (g590) & (!g547) & (g251)) + ((!sk[60]) & (g592) & (g590) & (g547) & (!g251)) + ((!sk[60]) & (g592) & (g590) & (g547) & (g251)) + ((sk[60]) & (!g592) & (!g590) & (!g547) & (!g251)) + ((sk[60]) & (!g592) & (!g590) & (!g547) & (g251)) + ((sk[60]) & (!g592) & (!g590) & (g547) & (!g251)) + ((sk[60]) & (!g592) & (!g590) & (g547) & (g251)) + ((sk[60]) & (!g592) & (g590) & (!g547) & (!g251)) + ((sk[60]) & (!g592) & (g590) & (!g547) & (g251)) + ((sk[60]) & (g592) & (!g590) & (!g547) & (!g251)) + ((sk[60]) & (g592) & (!g590) & (!g547) & (g251)) + ((sk[60]) & (g592) & (!g590) & (g547) & (!g251)) + ((sk[60]) & (g592) & (!g590) & (g547) & (g251)) + ((sk[60]) & (g592) & (g590) & (!g547) & (!g251)) + ((sk[60]) & (g592) & (g590) & (!g547) & (g251)) + ((sk[60]) & (g592) & (g590) & (g547) & (g251)));
	assign g1707 = (((!g592) & (!sk[61]) & (!g590) & (g462) & (g251)) + ((!g592) & (!sk[61]) & (g590) & (!g462) & (!g251)) + ((!g592) & (!sk[61]) & (g590) & (!g462) & (g251)) + ((!g592) & (!sk[61]) & (g590) & (g462) & (!g251)) + ((!g592) & (!sk[61]) & (g590) & (g462) & (g251)) + ((!g592) & (sk[61]) & (!g590) & (!g462) & (!g251)) + ((!g592) & (sk[61]) & (!g590) & (!g462) & (g251)) + ((!g592) & (sk[61]) & (!g590) & (g462) & (!g251)) + ((!g592) & (sk[61]) & (!g590) & (g462) & (g251)) + ((!g592) & (sk[61]) & (g590) & (!g462) & (!g251)) + ((!g592) & (sk[61]) & (g590) & (!g462) & (g251)) + ((g592) & (!sk[61]) & (!g590) & (g462) & (!g251)) + ((g592) & (!sk[61]) & (!g590) & (g462) & (g251)) + ((g592) & (!sk[61]) & (g590) & (!g462) & (!g251)) + ((g592) & (!sk[61]) & (g590) & (!g462) & (g251)) + ((g592) & (!sk[61]) & (g590) & (g462) & (!g251)) + ((g592) & (!sk[61]) & (g590) & (g462) & (g251)) + ((g592) & (sk[61]) & (!g590) & (!g462) & (!g251)) + ((g592) & (sk[61]) & (!g590) & (!g462) & (g251)) + ((g592) & (sk[61]) & (!g590) & (g462) & (!g251)) + ((g592) & (sk[61]) & (!g590) & (g462) & (g251)) + ((g592) & (sk[61]) & (g590) & (!g462) & (!g251)) + ((g592) & (sk[61]) & (g590) & (!g462) & (g251)) + ((g592) & (sk[61]) & (g590) & (g462) & (g251)));
	assign g1708 = (((!g1709) & (sk[62]) & (!g1710)) + ((g1709) & (!sk[62]) & (!g1710)) + ((g1709) & (!sk[62]) & (g1710)));
	assign g1709 = (((!g134) & (sk[63]) & (g1711)) + ((g134) & (!sk[63]) & (!g1711)) + ((g134) & (!sk[63]) & (g1711)));
	assign g1710 = (((g134) & (!sk[64]) & (!g1714)) + ((g134) & (!sk[64]) & (g1714)) + ((g134) & (sk[64]) & (g1714)));
	assign g1711 = (((!sk[65]) & (g1712) & (!g1713)) + ((!sk[65]) & (g1712) & (g1713)) + ((sk[65]) & (!g1712) & (!g1713)));
	assign g1712 = (((!g100) & (sk[66]) & (g1717)) + ((g100) & (!sk[66]) & (!g1717)) + ((g100) & (!sk[66]) & (g1717)));
	assign g1713 = (((g100) & (!sk[67]) & (!g1718)) + ((g100) & (!sk[67]) & (g1718)) + ((g100) & (sk[67]) & (g1718)));
	assign g1714 = (((!sk[68]) & (g1715) & (!g1716)) + ((!sk[68]) & (g1715) & (g1716)) + ((sk[68]) & (!g1715) & (!g1716)));
	assign g1715 = (((!g100) & (sk[69]) & (g1719)) + ((g100) & (!sk[69]) & (!g1719)) + ((g100) & (!sk[69]) & (g1719)));
	assign g1716 = (((g100) & (!sk[70]) & (!g1720)) + ((g100) & (!sk[70]) & (g1720)) + ((g100) & (sk[70]) & (g1720)));
	assign g1717 = (((!sk[71]) & (g164) & (!g13) & (!g251)) + ((!sk[71]) & (g164) & (!g13) & (g251)) + ((!sk[71]) & (g164) & (g13) & (!g251)) + ((!sk[71]) & (g164) & (g13) & (g251)) + ((sk[71]) & (!g164) & (!g13) & (!g251)) + ((sk[71]) & (!g164) & (!g13) & (g251)) + ((sk[71]) & (!g164) & (g13) & (!g251)) + ((sk[71]) & (!g164) & (g13) & (g251)) + ((sk[71]) & (g164) & (!g13) & (!g251)) + ((sk[71]) & (g164) & (!g13) & (g251)) + ((sk[71]) & (g164) & (g13) & (!g251)));
	assign g1718 = (((!sk[72]) & (!g164) & (!g13) & (g18) & (g251)) + ((!sk[72]) & (!g164) & (g13) & (!g18) & (!g251)) + ((!sk[72]) & (!g164) & (g13) & (!g18) & (g251)) + ((!sk[72]) & (!g164) & (g13) & (g18) & (!g251)) + ((!sk[72]) & (!g164) & (g13) & (g18) & (g251)) + ((!sk[72]) & (g164) & (!g13) & (g18) & (!g251)) + ((!sk[72]) & (g164) & (!g13) & (g18) & (g251)) + ((!sk[72]) & (g164) & (g13) & (!g18) & (!g251)) + ((!sk[72]) & (g164) & (g13) & (!g18) & (g251)) + ((!sk[72]) & (g164) & (g13) & (g18) & (!g251)) + ((!sk[72]) & (g164) & (g13) & (g18) & (g251)) + ((sk[72]) & (!g164) & (!g13) & (!g18) & (!g251)) + ((sk[72]) & (!g164) & (!g13) & (!g18) & (g251)) + ((sk[72]) & (!g164) & (!g13) & (g18) & (!g251)) + ((sk[72]) & (!g164) & (!g13) & (g18) & (g251)) + ((sk[72]) & (!g164) & (g13) & (!g18) & (!g251)) + ((sk[72]) & (!g164) & (g13) & (!g18) & (g251)) + ((sk[72]) & (!g164) & (g13) & (g18) & (!g251)) + ((sk[72]) & (!g164) & (g13) & (g18) & (g251)) + ((sk[72]) & (g164) & (!g13) & (!g18) & (!g251)) + ((sk[72]) & (g164) & (!g13) & (!g18) & (g251)) + ((sk[72]) & (g164) & (!g13) & (g18) & (!g251)) + ((sk[72]) & (g164) & (!g13) & (g18) & (g251)) + ((sk[72]) & (g164) & (g13) & (g18) & (!g251)));
	assign g1719 = (((!g164) & (!sk[73]) & (!g13) & (g115) & (g251)) + ((!g164) & (!sk[73]) & (g13) & (!g115) & (!g251)) + ((!g164) & (!sk[73]) & (g13) & (!g115) & (g251)) + ((!g164) & (!sk[73]) & (g13) & (g115) & (!g251)) + ((!g164) & (!sk[73]) & (g13) & (g115) & (g251)) + ((!g164) & (sk[73]) & (!g13) & (!g115) & (!g251)) + ((!g164) & (sk[73]) & (!g13) & (!g115) & (g251)) + ((!g164) & (sk[73]) & (!g13) & (g115) & (!g251)) + ((!g164) & (sk[73]) & (!g13) & (g115) & (g251)) + ((!g164) & (sk[73]) & (g13) & (!g115) & (!g251)) + ((!g164) & (sk[73]) & (g13) & (!g115) & (g251)) + ((!g164) & (sk[73]) & (g13) & (g115) & (!g251)) + ((!g164) & (sk[73]) & (g13) & (g115) & (g251)) + ((g164) & (!sk[73]) & (!g13) & (g115) & (!g251)) + ((g164) & (!sk[73]) & (!g13) & (g115) & (g251)) + ((g164) & (!sk[73]) & (g13) & (!g115) & (!g251)) + ((g164) & (!sk[73]) & (g13) & (!g115) & (g251)) + ((g164) & (!sk[73]) & (g13) & (g115) & (!g251)) + ((g164) & (!sk[73]) & (g13) & (g115) & (g251)) + ((g164) & (sk[73]) & (!g13) & (!g115) & (!g251)) + ((g164) & (sk[73]) & (!g13) & (!g115) & (g251)) + ((g164) & (sk[73]) & (!g13) & (g115) & (!g251)) + ((g164) & (sk[73]) & (!g13) & (g115) & (g251)) + ((g164) & (sk[73]) & (g13) & (g115) & (!g251)));
	assign g1720 = (((!sk[74]) & (g164) & (!g13)) + ((!sk[74]) & (g164) & (g13)) + ((sk[74]) & (!g164) & (!g13)) + ((sk[74]) & (!g164) & (g13)) + ((sk[74]) & (g164) & (!g13)));
	assign g1721 = (((!g171) & (sk[75]) & (!g1722)) + ((g171) & (!sk[75]) & (!g1722)) + ((g171) & (!sk[75]) & (g1722)));
	assign g1722 = (((!sk[76]) & (g171) & (!g1723)) + ((!sk[76]) & (g171) & (g1723)) + ((sk[76]) & (!g171) & (g1723)));
	assign g1723 = (((!g1724) & (sk[77]) & (!g1725)) + ((g1724) & (!sk[77]) & (!g1725)) + ((g1724) & (!sk[77]) & (g1725)));
	assign g1724 = (((!sk[78]) & (i_10_) & (!g1726)) + ((!sk[78]) & (i_10_) & (g1726)) + ((sk[78]) & (!i_10_) & (g1726)));
	assign g1725 = (((!sk[79]) & (i_10_) & (!g1727)) + ((!sk[79]) & (i_10_) & (g1727)) + ((sk[79]) & (i_10_) & (g1727)));
	assign g1726 = (((!i_9_) & (!i_11_) & (!sk[80]) & (g251) & (i_15_)) + ((!i_9_) & (!i_11_) & (sk[80]) & (!g251) & (!i_15_)) + ((!i_9_) & (!i_11_) & (sk[80]) & (!g251) & (i_15_)) + ((!i_9_) & (!i_11_) & (sk[80]) & (g251) & (!i_15_)) + ((!i_9_) & (!i_11_) & (sk[80]) & (g251) & (i_15_)) + ((!i_9_) & (i_11_) & (!sk[80]) & (!g251) & (!i_15_)) + ((!i_9_) & (i_11_) & (!sk[80]) & (!g251) & (i_15_)) + ((!i_9_) & (i_11_) & (!sk[80]) & (g251) & (!i_15_)) + ((!i_9_) & (i_11_) & (!sk[80]) & (g251) & (i_15_)) + ((!i_9_) & (i_11_) & (sk[80]) & (!g251) & (!i_15_)) + ((!i_9_) & (i_11_) & (sk[80]) & (!g251) & (i_15_)) + ((!i_9_) & (i_11_) & (sk[80]) & (g251) & (!i_15_)) + ((!i_9_) & (i_11_) & (sk[80]) & (g251) & (i_15_)) + ((i_9_) & (!i_11_) & (!sk[80]) & (g251) & (!i_15_)) + ((i_9_) & (!i_11_) & (!sk[80]) & (g251) & (i_15_)) + ((i_9_) & (!i_11_) & (sk[80]) & (!g251) & (!i_15_)) + ((i_9_) & (!i_11_) & (sk[80]) & (!g251) & (i_15_)) + ((i_9_) & (!i_11_) & (sk[80]) & (g251) & (!i_15_)) + ((i_9_) & (i_11_) & (!sk[80]) & (!g251) & (!i_15_)) + ((i_9_) & (i_11_) & (!sk[80]) & (!g251) & (i_15_)) + ((i_9_) & (i_11_) & (!sk[80]) & (g251) & (!i_15_)) + ((i_9_) & (i_11_) & (!sk[80]) & (g251) & (i_15_)) + ((i_9_) & (i_11_) & (sk[80]) & (!g251) & (!i_15_)) + ((i_9_) & (i_11_) & (sk[80]) & (!g251) & (i_15_)) + ((i_9_) & (i_11_) & (sk[80]) & (g251) & (!i_15_)) + ((i_9_) & (i_11_) & (sk[80]) & (g251) & (i_15_)));
	assign g1727 = (((!sk[81]) & (!i_9_) & (!i_11_) & (g285) & (i_15_)) + ((!sk[81]) & (!i_9_) & (i_11_) & (!g285) & (!i_15_)) + ((!sk[81]) & (!i_9_) & (i_11_) & (!g285) & (i_15_)) + ((!sk[81]) & (!i_9_) & (i_11_) & (g285) & (!i_15_)) + ((!sk[81]) & (!i_9_) & (i_11_) & (g285) & (i_15_)) + ((!sk[81]) & (i_9_) & (!i_11_) & (g285) & (!i_15_)) + ((!sk[81]) & (i_9_) & (!i_11_) & (g285) & (i_15_)) + ((!sk[81]) & (i_9_) & (i_11_) & (!g285) & (!i_15_)) + ((!sk[81]) & (i_9_) & (i_11_) & (!g285) & (i_15_)) + ((!sk[81]) & (i_9_) & (i_11_) & (g285) & (!i_15_)) + ((!sk[81]) & (i_9_) & (i_11_) & (g285) & (i_15_)) + ((sk[81]) & (!i_9_) & (!i_11_) & (!g285) & (!i_15_)) + ((sk[81]) & (!i_9_) & (!i_11_) & (!g285) & (i_15_)) + ((sk[81]) & (!i_9_) & (!i_11_) & (g285) & (!i_15_)) + ((sk[81]) & (!i_9_) & (!i_11_) & (g285) & (i_15_)) + ((sk[81]) & (!i_9_) & (i_11_) & (!g285) & (!i_15_)) + ((sk[81]) & (!i_9_) & (i_11_) & (!g285) & (i_15_)) + ((sk[81]) & (!i_9_) & (i_11_) & (g285) & (!i_15_)) + ((sk[81]) & (!i_9_) & (i_11_) & (g285) & (i_15_)) + ((sk[81]) & (i_9_) & (!i_11_) & (!g285) & (!i_15_)) + ((sk[81]) & (i_9_) & (!i_11_) & (g285) & (!i_15_)) + ((sk[81]) & (i_9_) & (!i_11_) & (g285) & (i_15_)) + ((sk[81]) & (i_9_) & (i_11_) & (!g285) & (!i_15_)) + ((sk[81]) & (i_9_) & (i_11_) & (!g285) & (i_15_)) + ((sk[81]) & (i_9_) & (i_11_) & (g285) & (!i_15_)) + ((sk[81]) & (i_9_) & (i_11_) & (g285) & (i_15_)));
	assign g1728 = (((!sk[82]) & (g1729) & (!g1730)) + ((!sk[82]) & (g1729) & (g1730)) + ((sk[82]) & (!g1729) & (!g1730)));
	assign g1729 = (((!sk[83]) & (g465) & (!g1731)) + ((!sk[83]) & (g465) & (g1731)) + ((sk[83]) & (!g465) & (g1731)));
	assign g1730 = (((g465) & (!sk[84]) & (!g1732)) + ((g465) & (!sk[84]) & (g1732)) + ((g465) & (sk[84]) & (g1732)));
	assign g1731 = (((!sk[85]) & (g89) & (!g99)) + ((!sk[85]) & (g89) & (g99)) + ((sk[85]) & (g89) & (!g99)));
	assign g1732 = (((!sk[86]) & (g1733) & (!g1734)) + ((!sk[86]) & (g1733) & (g1734)) + ((sk[86]) & (!g1733) & (!g1734)));
	assign g1733 = (((!g89) & (sk[87]) & (g1735)) + ((g89) & (!sk[87]) & (!g1735)) + ((g89) & (!sk[87]) & (g1735)));
	assign g1734 = (((g89) & (!sk[88]) & (!g1736)) + ((g89) & (!sk[88]) & (g1736)) + ((g89) & (sk[88]) & (g1736)));
	assign g1735 = (((!sk[89]) & (!g468) & (!g467) & (g475) & (g462)) + ((!sk[89]) & (!g468) & (g467) & (!g475) & (!g462)) + ((!sk[89]) & (!g468) & (g467) & (!g475) & (g462)) + ((!sk[89]) & (!g468) & (g467) & (g475) & (!g462)) + ((!sk[89]) & (!g468) & (g467) & (g475) & (g462)) + ((!sk[89]) & (g468) & (!g467) & (g475) & (!g462)) + ((!sk[89]) & (g468) & (!g467) & (g475) & (g462)) + ((!sk[89]) & (g468) & (g467) & (!g475) & (!g462)) + ((!sk[89]) & (g468) & (g467) & (!g475) & (g462)) + ((!sk[89]) & (g468) & (g467) & (g475) & (!g462)) + ((!sk[89]) & (g468) & (g467) & (g475) & (g462)) + ((sk[89]) & (g468) & (g467) & (g475) & (g462)));
	assign g1736 = (((!sk[90]) & (g99) & (!g462)) + ((!sk[90]) & (g99) & (g462)) + ((sk[90]) & (!g99) & (!g462)) + ((sk[90]) & (!g99) & (g462)) + ((sk[90]) & (g99) & (g462)));
	assign g1737 = (((!sk[91]) & (g1738) & (!g1739)) + ((!sk[91]) & (g1738) & (g1739)) + ((sk[91]) & (!g1738) & (!g1739)));
	assign g1738 = (((!sk[92]) & (g477) & (!g1740)) + ((!sk[92]) & (g477) & (g1740)) + ((sk[92]) & (!g477) & (g1740)));
	assign g1739 = (((g477) & (!sk[93]) & (!g1741)) + ((g477) & (!sk[93]) & (g1741)) + ((g477) & (sk[93]) & (g1741)));
	assign g1740 = (((!sk[94]) & (g118) & (!g1744)) + ((!sk[94]) & (g118) & (g1744)) + ((sk[94]) & (!g118) & (g1744)));
	assign g1741 = (((!g1742) & (sk[95]) & (!g1743)) + ((g1742) & (!sk[95]) & (!g1743)) + ((g1742) & (!sk[95]) & (g1743)));
	assign g1742 = (((!g118) & (sk[96]) & (g1745)) + ((g118) & (!sk[96]) & (!g1745)) + ((g118) & (!sk[96]) & (g1745)));
	assign g1743 = (((!sk[97]) & (g118) & (!g1746)) + ((!sk[97]) & (g118) & (g1746)) + ((sk[97]) & (g118) & (g1746)));
	assign g1744 = (((!g491) & (!g494) & (g134) & (!sk[98]) & (g492)) + ((!g491) & (g494) & (!g134) & (!sk[98]) & (!g492)) + ((!g491) & (g494) & (!g134) & (!sk[98]) & (g492)) + ((!g491) & (g494) & (g134) & (!sk[98]) & (!g492)) + ((!g491) & (g494) & (g134) & (!sk[98]) & (g492)) + ((g491) & (!g494) & (g134) & (!sk[98]) & (!g492)) + ((g491) & (!g494) & (g134) & (!sk[98]) & (g492)) + ((g491) & (g494) & (!g134) & (!sk[98]) & (!g492)) + ((g491) & (g494) & (!g134) & (!sk[98]) & (g492)) + ((g491) & (g494) & (!g134) & (sk[98]) & (g492)) + ((g491) & (g494) & (g134) & (!sk[98]) & (!g492)) + ((g491) & (g494) & (g134) & (!sk[98]) & (g492)));
	assign g1745 = (((g491) & (!g494) & (!sk[99]) & (!g492)) + ((g491) & (!g494) & (!sk[99]) & (g492)) + ((g491) & (g494) & (!sk[99]) & (!g492)) + ((g491) & (g494) & (!sk[99]) & (g492)) + ((g491) & (g494) & (sk[99]) & (g492)));
	assign g1746 = (((!sk[100]) & (!g491) & (!g494) & (g481) & (g492)) + ((!sk[100]) & (!g491) & (g494) & (!g481) & (!g492)) + ((!sk[100]) & (!g491) & (g494) & (!g481) & (g492)) + ((!sk[100]) & (!g491) & (g494) & (g481) & (!g492)) + ((!sk[100]) & (!g491) & (g494) & (g481) & (g492)) + ((!sk[100]) & (g491) & (!g494) & (g481) & (!g492)) + ((!sk[100]) & (g491) & (!g494) & (g481) & (g492)) + ((!sk[100]) & (g491) & (g494) & (!g481) & (!g492)) + ((!sk[100]) & (g491) & (g494) & (!g481) & (g492)) + ((!sk[100]) & (g491) & (g494) & (g481) & (!g492)) + ((!sk[100]) & (g491) & (g494) & (g481) & (g492)) + ((sk[100]) & (g491) & (g494) & (g481) & (g492)));
	assign g1747 = (((g145) & (!sk[101]) & (!g1748)) + ((g145) & (!sk[101]) & (g1748)) + ((g145) & (sk[101]) & (!g1748)));
	assign g1748 = (((g145) & (!sk[102]) & (!g1749)) + ((g145) & (!sk[102]) & (g1749)) + ((g145) & (sk[102]) & (g1749)));
	assign g1749 = (((!g1750) & (sk[103]) & (!g1751)) + ((g1750) & (!sk[103]) & (!g1751)) + ((g1750) & (!sk[103]) & (g1751)));
	assign g1750 = (((!i_15_) & (sk[104]) & (g1752)) + ((i_15_) & (!sk[104]) & (!g1752)) + ((i_15_) & (!sk[104]) & (g1752)));
	assign g1751 = (((!sk[105]) & (i_15_) & (!g1753)) + ((!sk[105]) & (i_15_) & (g1753)) + ((sk[105]) & (i_15_) & (g1753)));
	assign g1752 = (((!i_10_) & (!sk[106]) & (!i_9_) & (g48) & (i_11_)) + ((!i_10_) & (!sk[106]) & (i_9_) & (!g48) & (!i_11_)) + ((!i_10_) & (!sk[106]) & (i_9_) & (!g48) & (i_11_)) + ((!i_10_) & (!sk[106]) & (i_9_) & (g48) & (!i_11_)) + ((!i_10_) & (!sk[106]) & (i_9_) & (g48) & (i_11_)) + ((!i_10_) & (sk[106]) & (!i_9_) & (!g48) & (!i_11_)) + ((!i_10_) & (sk[106]) & (!i_9_) & (g48) & (!i_11_)) + ((!i_10_) & (sk[106]) & (!i_9_) & (g48) & (i_11_)) + ((!i_10_) & (sk[106]) & (i_9_) & (!g48) & (!i_11_)) + ((!i_10_) & (sk[106]) & (i_9_) & (g48) & (!i_11_)) + ((!i_10_) & (sk[106]) & (i_9_) & (g48) & (i_11_)) + ((i_10_) & (!sk[106]) & (!i_9_) & (g48) & (!i_11_)) + ((i_10_) & (!sk[106]) & (!i_9_) & (g48) & (i_11_)) + ((i_10_) & (!sk[106]) & (i_9_) & (!g48) & (!i_11_)) + ((i_10_) & (!sk[106]) & (i_9_) & (!g48) & (i_11_)) + ((i_10_) & (!sk[106]) & (i_9_) & (g48) & (!i_11_)) + ((i_10_) & (!sk[106]) & (i_9_) & (g48) & (i_11_)) + ((i_10_) & (sk[106]) & (!i_9_) & (!g48) & (i_11_)) + ((i_10_) & (sk[106]) & (!i_9_) & (g48) & (!i_11_)) + ((i_10_) & (sk[106]) & (!i_9_) & (g48) & (i_11_)) + ((i_10_) & (sk[106]) & (i_9_) & (!g48) & (!i_11_)) + ((i_10_) & (sk[106]) & (i_9_) & (!g48) & (i_11_)) + ((i_10_) & (sk[106]) & (i_9_) & (g48) & (!i_11_)) + ((i_10_) & (sk[106]) & (i_9_) & (g48) & (i_11_)));
	assign g1753 = (((!i_10_) & (!i_9_) & (!sk[107]) & (g91) & (i_11_)) + ((!i_10_) & (!i_9_) & (sk[107]) & (!g91) & (!i_11_)) + ((!i_10_) & (!i_9_) & (sk[107]) & (!g91) & (i_11_)) + ((!i_10_) & (!i_9_) & (sk[107]) & (g91) & (!i_11_)) + ((!i_10_) & (!i_9_) & (sk[107]) & (g91) & (i_11_)) + ((!i_10_) & (i_9_) & (!sk[107]) & (!g91) & (!i_11_)) + ((!i_10_) & (i_9_) & (!sk[107]) & (!g91) & (i_11_)) + ((!i_10_) & (i_9_) & (!sk[107]) & (g91) & (!i_11_)) + ((!i_10_) & (i_9_) & (!sk[107]) & (g91) & (i_11_)) + ((!i_10_) & (i_9_) & (sk[107]) & (g91) & (!i_11_)) + ((!i_10_) & (i_9_) & (sk[107]) & (g91) & (i_11_)) + ((i_10_) & (!i_9_) & (!sk[107]) & (g91) & (!i_11_)) + ((i_10_) & (!i_9_) & (!sk[107]) & (g91) & (i_11_)) + ((i_10_) & (!i_9_) & (sk[107]) & (!g91) & (i_11_)) + ((i_10_) & (!i_9_) & (sk[107]) & (g91) & (!i_11_)) + ((i_10_) & (!i_9_) & (sk[107]) & (g91) & (i_11_)) + ((i_10_) & (i_9_) & (!sk[107]) & (!g91) & (!i_11_)) + ((i_10_) & (i_9_) & (!sk[107]) & (!g91) & (i_11_)) + ((i_10_) & (i_9_) & (!sk[107]) & (g91) & (!i_11_)) + ((i_10_) & (i_9_) & (!sk[107]) & (g91) & (i_11_)) + ((i_10_) & (i_9_) & (sk[107]) & (!g91) & (!i_11_)) + ((i_10_) & (i_9_) & (sk[107]) & (!g91) & (i_11_)) + ((i_10_) & (i_9_) & (sk[107]) & (g91) & (!i_11_)) + ((i_10_) & (i_9_) & (sk[107]) & (g91) & (i_11_)));
	assign g1754 = (((!sk[108]) & (g91) & (!g1755)) + ((!sk[108]) & (g91) & (g1755)) + ((sk[108]) & (!g91) & (!g1755)));
	assign g1755 = (((!g91) & (sk[109]) & (g1756)) + ((g91) & (!sk[109]) & (!g1756)) + ((g91) & (!sk[109]) & (g1756)));
	assign g1756 = (((!g1757) & (sk[110]) & (!g1758)) + ((g1757) & (!sk[110]) & (!g1758)) + ((g1757) & (!sk[110]) & (g1758)));
	assign g1757 = (((!sk[111]) & (i_10_) & (!g1759)) + ((!sk[111]) & (i_10_) & (g1759)) + ((sk[111]) & (!i_10_) & (g1759)));
	assign g1758 = (((i_10_) & (!sk[112]) & (!g1760)) + ((i_10_) & (!sk[112]) & (g1760)) + ((i_10_) & (sk[112]) & (g1760)));
	assign g1759 = (((!sk[113]) & (!i_15_) & (!i_11_) & (g145) & (i_9_)) + ((!sk[113]) & (!i_15_) & (i_11_) & (!g145) & (!i_9_)) + ((!sk[113]) & (!i_15_) & (i_11_) & (!g145) & (i_9_)) + ((!sk[113]) & (!i_15_) & (i_11_) & (g145) & (!i_9_)) + ((!sk[113]) & (!i_15_) & (i_11_) & (g145) & (i_9_)) + ((!sk[113]) & (i_15_) & (!i_11_) & (g145) & (!i_9_)) + ((!sk[113]) & (i_15_) & (!i_11_) & (g145) & (i_9_)) + ((!sk[113]) & (i_15_) & (i_11_) & (!g145) & (!i_9_)) + ((!sk[113]) & (i_15_) & (i_11_) & (!g145) & (i_9_)) + ((!sk[113]) & (i_15_) & (i_11_) & (g145) & (!i_9_)) + ((!sk[113]) & (i_15_) & (i_11_) & (g145) & (i_9_)) + ((sk[113]) & (!i_15_) & (!i_11_) & (!g145) & (i_9_)) + ((sk[113]) & (!i_15_) & (i_11_) & (!g145) & (!i_9_)) + ((sk[113]) & (!i_15_) & (i_11_) & (!g145) & (i_9_)) + ((sk[113]) & (!i_15_) & (i_11_) & (g145) & (!i_9_)) + ((sk[113]) & (i_15_) & (!i_11_) & (!g145) & (!i_9_)) + ((sk[113]) & (i_15_) & (!i_11_) & (!g145) & (i_9_)) + ((sk[113]) & (i_15_) & (!i_11_) & (g145) & (!i_9_)) + ((sk[113]) & (i_15_) & (!i_11_) & (g145) & (i_9_)) + ((sk[113]) & (i_15_) & (i_11_) & (!g145) & (!i_9_)) + ((sk[113]) & (i_15_) & (i_11_) & (!g145) & (i_9_)) + ((sk[113]) & (i_15_) & (i_11_) & (g145) & (!i_9_)) + ((sk[113]) & (i_15_) & (i_11_) & (g145) & (i_9_)));
	assign g1760 = (((!i_15_) & (!sk[114]) & (!i_11_) & (g151) & (i_9_)) + ((!i_15_) & (!sk[114]) & (i_11_) & (!g151) & (!i_9_)) + ((!i_15_) & (!sk[114]) & (i_11_) & (!g151) & (i_9_)) + ((!i_15_) & (!sk[114]) & (i_11_) & (g151) & (!i_9_)) + ((!i_15_) & (!sk[114]) & (i_11_) & (g151) & (i_9_)) + ((!i_15_) & (sk[114]) & (!i_11_) & (!g151) & (!i_9_)) + ((!i_15_) & (sk[114]) & (!i_11_) & (!g151) & (i_9_)) + ((!i_15_) & (sk[114]) & (!i_11_) & (g151) & (!i_9_)) + ((!i_15_) & (sk[114]) & (!i_11_) & (g151) & (i_9_)) + ((!i_15_) & (sk[114]) & (i_11_) & (!g151) & (!i_9_)) + ((!i_15_) & (sk[114]) & (i_11_) & (!g151) & (i_9_)) + ((!i_15_) & (sk[114]) & (i_11_) & (g151) & (!i_9_)) + ((i_15_) & (!sk[114]) & (!i_11_) & (g151) & (!i_9_)) + ((i_15_) & (!sk[114]) & (!i_11_) & (g151) & (i_9_)) + ((i_15_) & (!sk[114]) & (i_11_) & (!g151) & (!i_9_)) + ((i_15_) & (!sk[114]) & (i_11_) & (!g151) & (i_9_)) + ((i_15_) & (!sk[114]) & (i_11_) & (g151) & (!i_9_)) + ((i_15_) & (!sk[114]) & (i_11_) & (g151) & (i_9_)) + ((i_15_) & (sk[114]) & (!i_11_) & (!g151) & (!i_9_)) + ((i_15_) & (sk[114]) & (!i_11_) & (!g151) & (i_9_)) + ((i_15_) & (sk[114]) & (!i_11_) & (g151) & (!i_9_)) + ((i_15_) & (sk[114]) & (!i_11_) & (g151) & (i_9_)) + ((i_15_) & (sk[114]) & (i_11_) & (!g151) & (!i_9_)) + ((i_15_) & (sk[114]) & (i_11_) & (!g151) & (i_9_)) + ((i_15_) & (sk[114]) & (i_11_) & (g151) & (!i_9_)) + ((i_15_) & (sk[114]) & (i_11_) & (g151) & (i_9_)));
	assign g1761 = (((g13) & (!sk[115]) & (!g1762)) + ((g13) & (!sk[115]) & (g1762)) + ((g13) & (sk[115]) & (!g1762)));
	assign g1762 = (((!sk[116]) & (g13) & (!g1763)) + ((!sk[116]) & (g13) & (g1763)) + ((sk[116]) & (g13) & (g1763)));
	assign g1763 = (((!sk[117]) & (g1764) & (!g1765)) + ((!sk[117]) & (g1764) & (g1765)) + ((sk[117]) & (!g1764) & (!g1765)));
	assign g1764 = (((!i_9_) & (sk[118]) & (g1766)) + ((i_9_) & (!sk[118]) & (!g1766)) + ((i_9_) & (!sk[118]) & (g1766)));
	assign g1765 = (((i_9_) & (!sk[119]) & (!g1767)) + ((i_9_) & (!sk[119]) & (g1767)) + ((i_9_) & (sk[119]) & (g1767)));
	assign g1766 = (((!sk[120]) & (!i_15_) & (!i_10_) & (g112) & (i_11_)) + ((!sk[120]) & (!i_15_) & (i_10_) & (!g112) & (!i_11_)) + ((!sk[120]) & (!i_15_) & (i_10_) & (!g112) & (i_11_)) + ((!sk[120]) & (!i_15_) & (i_10_) & (g112) & (!i_11_)) + ((!sk[120]) & (!i_15_) & (i_10_) & (g112) & (i_11_)) + ((!sk[120]) & (i_15_) & (!i_10_) & (g112) & (!i_11_)) + ((!sk[120]) & (i_15_) & (!i_10_) & (g112) & (i_11_)) + ((!sk[120]) & (i_15_) & (i_10_) & (!g112) & (!i_11_)) + ((!sk[120]) & (i_15_) & (i_10_) & (!g112) & (i_11_)) + ((!sk[120]) & (i_15_) & (i_10_) & (g112) & (!i_11_)) + ((!sk[120]) & (i_15_) & (i_10_) & (g112) & (i_11_)) + ((sk[120]) & (!i_15_) & (!i_10_) & (!g112) & (!i_11_)) + ((sk[120]) & (!i_15_) & (!i_10_) & (!g112) & (i_11_)) + ((sk[120]) & (!i_15_) & (!i_10_) & (g112) & (!i_11_)) + ((sk[120]) & (!i_15_) & (!i_10_) & (g112) & (i_11_)) + ((sk[120]) & (!i_15_) & (i_10_) & (!g112) & (!i_11_)) + ((sk[120]) & (!i_15_) & (i_10_) & (!g112) & (i_11_)) + ((sk[120]) & (!i_15_) & (i_10_) & (g112) & (!i_11_)) + ((sk[120]) & (i_15_) & (!i_10_) & (!g112) & (!i_11_)) + ((sk[120]) & (i_15_) & (!i_10_) & (!g112) & (i_11_)) + ((sk[120]) & (i_15_) & (!i_10_) & (g112) & (!i_11_)) + ((sk[120]) & (i_15_) & (!i_10_) & (g112) & (i_11_)) + ((sk[120]) & (i_15_) & (i_10_) & (!g112) & (!i_11_)) + ((sk[120]) & (i_15_) & (i_10_) & (!g112) & (i_11_)) + ((sk[120]) & (i_15_) & (i_10_) & (g112) & (!i_11_)) + ((sk[120]) & (i_15_) & (i_10_) & (g112) & (i_11_)));
	assign g1767 = (((!i_15_) & (!i_10_) & (!sk[121]) & (g151) & (i_11_)) + ((!i_15_) & (!i_10_) & (sk[121]) & (!g151) & (!i_11_)) + ((!i_15_) & (!i_10_) & (sk[121]) & (!g151) & (i_11_)) + ((!i_15_) & (!i_10_) & (sk[121]) & (g151) & (!i_11_)) + ((!i_15_) & (!i_10_) & (sk[121]) & (g151) & (i_11_)) + ((!i_15_) & (i_10_) & (!sk[121]) & (!g151) & (!i_11_)) + ((!i_15_) & (i_10_) & (!sk[121]) & (!g151) & (i_11_)) + ((!i_15_) & (i_10_) & (!sk[121]) & (g151) & (!i_11_)) + ((!i_15_) & (i_10_) & (!sk[121]) & (g151) & (i_11_)) + ((!i_15_) & (i_10_) & (sk[121]) & (!g151) & (!i_11_)) + ((!i_15_) & (i_10_) & (sk[121]) & (!g151) & (i_11_)) + ((!i_15_) & (i_10_) & (sk[121]) & (g151) & (i_11_)) + ((i_15_) & (!i_10_) & (!sk[121]) & (g151) & (!i_11_)) + ((i_15_) & (!i_10_) & (!sk[121]) & (g151) & (i_11_)) + ((i_15_) & (!i_10_) & (sk[121]) & (!g151) & (!i_11_)) + ((i_15_) & (!i_10_) & (sk[121]) & (!g151) & (i_11_)) + ((i_15_) & (!i_10_) & (sk[121]) & (g151) & (!i_11_)) + ((i_15_) & (!i_10_) & (sk[121]) & (g151) & (i_11_)) + ((i_15_) & (i_10_) & (!sk[121]) & (!g151) & (!i_11_)) + ((i_15_) & (i_10_) & (!sk[121]) & (!g151) & (i_11_)) + ((i_15_) & (i_10_) & (!sk[121]) & (g151) & (!i_11_)) + ((i_15_) & (i_10_) & (!sk[121]) & (g151) & (i_11_)) + ((i_15_) & (i_10_) & (sk[121]) & (!g151) & (!i_11_)) + ((i_15_) & (i_10_) & (sk[121]) & (!g151) & (i_11_)) + ((i_15_) & (i_10_) & (sk[121]) & (g151) & (!i_11_)) + ((i_15_) & (i_10_) & (sk[121]) & (g151) & (i_11_)));
	assign g1768 = (((!sk[122]) & (g91) & (!g1769)) + ((!sk[122]) & (g91) & (g1769)) + ((sk[122]) & (!g91) & (!g1769)));
	assign g1769 = (((!sk[123]) & (g91) & (!g1770)) + ((!sk[123]) & (g91) & (g1770)) + ((sk[123]) & (!g91) & (g1770)));
	assign g1770 = (((!g1771) & (sk[124]) & (!g1772)) + ((g1771) & (!sk[124]) & (!g1772)) + ((g1771) & (!sk[124]) & (g1772)));
	assign g1771 = (((!sk[125]) & (i_10_) & (!g1773)) + ((!sk[125]) & (i_10_) & (g1773)) + ((sk[125]) & (!i_10_) & (g1773)));
	assign g1772 = (((!sk[126]) & (i_10_) & (!g1774)) + ((!sk[126]) & (i_10_) & (g1774)) + ((sk[126]) & (i_10_) & (g1774)));
	assign g1773 = (((!i_15_) & (!sk[127]) & (!i_9_) & (g109) & (i_11_)) + ((!i_15_) & (!sk[127]) & (i_9_) & (!g109) & (!i_11_)) + ((!i_15_) & (!sk[127]) & (i_9_) & (!g109) & (i_11_)) + ((!i_15_) & (!sk[127]) & (i_9_) & (g109) & (!i_11_)) + ((!i_15_) & (!sk[127]) & (i_9_) & (g109) & (i_11_)) + ((!i_15_) & (sk[127]) & (!i_9_) & (!g109) & (!i_11_)) + ((!i_15_) & (sk[127]) & (!i_9_) & (!g109) & (i_11_)) + ((!i_15_) & (sk[127]) & (!i_9_) & (g109) & (i_11_)) + ((!i_15_) & (sk[127]) & (i_9_) & (!g109) & (!i_11_)) + ((!i_15_) & (sk[127]) & (i_9_) & (!g109) & (i_11_)) + ((!i_15_) & (sk[127]) & (i_9_) & (g109) & (!i_11_)) + ((!i_15_) & (sk[127]) & (i_9_) & (g109) & (i_11_)) + ((i_15_) & (!sk[127]) & (!i_9_) & (g109) & (!i_11_)) + ((i_15_) & (!sk[127]) & (!i_9_) & (g109) & (i_11_)) + ((i_15_) & (!sk[127]) & (i_9_) & (!g109) & (!i_11_)) + ((i_15_) & (!sk[127]) & (i_9_) & (!g109) & (i_11_)) + ((i_15_) & (!sk[127]) & (i_9_) & (g109) & (!i_11_)) + ((i_15_) & (!sk[127]) & (i_9_) & (g109) & (i_11_)) + ((i_15_) & (sk[127]) & (!i_9_) & (!g109) & (!i_11_)) + ((i_15_) & (sk[127]) & (!i_9_) & (!g109) & (i_11_)) + ((i_15_) & (sk[127]) & (!i_9_) & (g109) & (!i_11_)) + ((i_15_) & (sk[127]) & (!i_9_) & (g109) & (i_11_)) + ((i_15_) & (sk[127]) & (i_9_) & (!g109) & (!i_11_)) + ((i_15_) & (sk[127]) & (i_9_) & (!g109) & (i_11_)) + ((i_15_) & (sk[127]) & (i_9_) & (g109) & (!i_11_)) + ((i_15_) & (sk[127]) & (i_9_) & (g109) & (i_11_)));
	assign g1774 = (((!i_15_) & (!i_9_) & (!g136) & (sk[0]) & (!i_11_)) + ((!i_15_) & (!i_9_) & (!g136) & (sk[0]) & (i_11_)) + ((!i_15_) & (!i_9_) & (g136) & (!sk[0]) & (i_11_)) + ((!i_15_) & (!i_9_) & (g136) & (sk[0]) & (!i_11_)) + ((!i_15_) & (!i_9_) & (g136) & (sk[0]) & (i_11_)) + ((!i_15_) & (i_9_) & (!g136) & (!sk[0]) & (!i_11_)) + ((!i_15_) & (i_9_) & (!g136) & (!sk[0]) & (i_11_)) + ((!i_15_) & (i_9_) & (!g136) & (sk[0]) & (!i_11_)) + ((!i_15_) & (i_9_) & (!g136) & (sk[0]) & (i_11_)) + ((!i_15_) & (i_9_) & (g136) & (!sk[0]) & (!i_11_)) + ((!i_15_) & (i_9_) & (g136) & (!sk[0]) & (i_11_)) + ((!i_15_) & (i_9_) & (g136) & (sk[0]) & (!i_11_)) + ((i_15_) & (!i_9_) & (!g136) & (sk[0]) & (!i_11_)) + ((i_15_) & (!i_9_) & (!g136) & (sk[0]) & (i_11_)) + ((i_15_) & (!i_9_) & (g136) & (!sk[0]) & (!i_11_)) + ((i_15_) & (!i_9_) & (g136) & (!sk[0]) & (i_11_)) + ((i_15_) & (!i_9_) & (g136) & (sk[0]) & (!i_11_)) + ((i_15_) & (!i_9_) & (g136) & (sk[0]) & (i_11_)) + ((i_15_) & (i_9_) & (!g136) & (!sk[0]) & (!i_11_)) + ((i_15_) & (i_9_) & (!g136) & (!sk[0]) & (i_11_)) + ((i_15_) & (i_9_) & (!g136) & (sk[0]) & (!i_11_)) + ((i_15_) & (i_9_) & (!g136) & (sk[0]) & (i_11_)) + ((i_15_) & (i_9_) & (g136) & (!sk[0]) & (!i_11_)) + ((i_15_) & (i_9_) & (g136) & (!sk[0]) & (i_11_)) + ((i_15_) & (i_9_) & (g136) & (sk[0]) & (!i_11_)) + ((i_15_) & (i_9_) & (g136) & (sk[0]) & (i_11_)));
	assign g1775 = (((!sk[1]) & (g91) & (!g1776)) + ((!sk[1]) & (g91) & (g1776)) + ((sk[1]) & (!g91) & (!g1776)));
	assign g1776 = (((!g91) & (sk[2]) & (g1777)) + ((g91) & (!sk[2]) & (!g1777)) + ((g91) & (!sk[2]) & (g1777)));
	assign g1777 = (((!g1778) & (sk[3]) & (!g1779)) + ((g1778) & (!sk[3]) & (!g1779)) + ((g1778) & (!sk[3]) & (g1779)));
	assign g1778 = (((!i_9_) & (sk[4]) & (g1780)) + ((i_9_) & (!sk[4]) & (!g1780)) + ((i_9_) & (!sk[4]) & (g1780)));
	assign g1779 = (((i_9_) & (!sk[5]) & (!g1781)) + ((i_9_) & (!sk[5]) & (g1781)) + ((i_9_) & (sk[5]) & (g1781)));
	assign g1780 = (((!sk[6]) & (!i_15_) & (!i_10_) & (g136) & (i_11_)) + ((!sk[6]) & (!i_15_) & (i_10_) & (!g136) & (!i_11_)) + ((!sk[6]) & (!i_15_) & (i_10_) & (!g136) & (i_11_)) + ((!sk[6]) & (!i_15_) & (i_10_) & (g136) & (!i_11_)) + ((!sk[6]) & (!i_15_) & (i_10_) & (g136) & (i_11_)) + ((!sk[6]) & (i_15_) & (!i_10_) & (g136) & (!i_11_)) + ((!sk[6]) & (i_15_) & (!i_10_) & (g136) & (i_11_)) + ((!sk[6]) & (i_15_) & (i_10_) & (!g136) & (!i_11_)) + ((!sk[6]) & (i_15_) & (i_10_) & (!g136) & (i_11_)) + ((!sk[6]) & (i_15_) & (i_10_) & (g136) & (!i_11_)) + ((!sk[6]) & (i_15_) & (i_10_) & (g136) & (i_11_)) + ((sk[6]) & (!i_15_) & (!i_10_) & (!g136) & (!i_11_)) + ((sk[6]) & (!i_15_) & (!i_10_) & (!g136) & (i_11_)) + ((sk[6]) & (!i_15_) & (!i_10_) & (g136) & (!i_11_)) + ((sk[6]) & (!i_15_) & (!i_10_) & (g136) & (i_11_)) + ((sk[6]) & (!i_15_) & (i_10_) & (!g136) & (!i_11_)) + ((sk[6]) & (!i_15_) & (i_10_) & (!g136) & (i_11_)) + ((sk[6]) & (!i_15_) & (i_10_) & (g136) & (!i_11_)) + ((sk[6]) & (!i_15_) & (i_10_) & (g136) & (i_11_)) + ((sk[6]) & (i_15_) & (!i_10_) & (!g136) & (!i_11_)) + ((sk[6]) & (i_15_) & (!i_10_) & (!g136) & (i_11_)) + ((sk[6]) & (i_15_) & (!i_10_) & (g136) & (!i_11_)) + ((sk[6]) & (i_15_) & (i_10_) & (!g136) & (!i_11_)) + ((sk[6]) & (i_15_) & (i_10_) & (!g136) & (i_11_)) + ((sk[6]) & (i_15_) & (i_10_) & (g136) & (!i_11_)) + ((sk[6]) & (i_15_) & (i_10_) & (g136) & (i_11_)));
	assign g1781 = (((!i_15_) & (!i_10_) & (!sk[7]) & (g151) & (i_11_)) + ((!i_15_) & (!i_10_) & (sk[7]) & (!g151) & (!i_11_)) + ((!i_15_) & (!i_10_) & (sk[7]) & (!g151) & (i_11_)) + ((!i_15_) & (!i_10_) & (sk[7]) & (g151) & (!i_11_)) + ((!i_15_) & (!i_10_) & (sk[7]) & (g151) & (i_11_)) + ((!i_15_) & (i_10_) & (!sk[7]) & (!g151) & (!i_11_)) + ((!i_15_) & (i_10_) & (!sk[7]) & (!g151) & (i_11_)) + ((!i_15_) & (i_10_) & (!sk[7]) & (g151) & (!i_11_)) + ((!i_15_) & (i_10_) & (!sk[7]) & (g151) & (i_11_)) + ((!i_15_) & (i_10_) & (sk[7]) & (!g151) & (!i_11_)) + ((!i_15_) & (i_10_) & (sk[7]) & (!g151) & (i_11_)) + ((!i_15_) & (i_10_) & (sk[7]) & (g151) & (!i_11_)) + ((!i_15_) & (i_10_) & (sk[7]) & (g151) & (i_11_)) + ((i_15_) & (!i_10_) & (!sk[7]) & (g151) & (!i_11_)) + ((i_15_) & (!i_10_) & (!sk[7]) & (g151) & (i_11_)) + ((i_15_) & (!i_10_) & (sk[7]) & (!g151) & (!i_11_)) + ((i_15_) & (!i_10_) & (sk[7]) & (!g151) & (i_11_)) + ((i_15_) & (!i_10_) & (sk[7]) & (g151) & (!i_11_)) + ((i_15_) & (i_10_) & (!sk[7]) & (!g151) & (!i_11_)) + ((i_15_) & (i_10_) & (!sk[7]) & (!g151) & (i_11_)) + ((i_15_) & (i_10_) & (!sk[7]) & (g151) & (!i_11_)) + ((i_15_) & (i_10_) & (!sk[7]) & (g151) & (i_11_)) + ((i_15_) & (i_10_) & (sk[7]) & (!g151) & (!i_11_)) + ((i_15_) & (i_10_) & (sk[7]) & (!g151) & (i_11_)) + ((i_15_) & (i_10_) & (sk[7]) & (g151) & (!i_11_)) + ((i_15_) & (i_10_) & (sk[7]) & (g151) & (i_11_)));
	assign g1782 = (((!sk[8]) & (g1783) & (!g1784)) + ((!sk[8]) & (g1783) & (g1784)) + ((sk[8]) & (!g1783) & (!g1784)));
	assign g1783 = (((!sk[9]) & (g132) & (!g1785)) + ((!sk[9]) & (g132) & (g1785)) + ((sk[9]) & (!g132) & (g1785)));
	assign g1784 = (((!sk[10]) & (g132) & (!g1786)) + ((!sk[10]) & (g132) & (g1786)) + ((sk[10]) & (g132) & (g1786)));
	assign g1785 = (((!g109) & (sk[11]) & (g1789)) + ((g109) & (!sk[11]) & (!g1789)) + ((g109) & (!sk[11]) & (g1789)));
	assign g1786 = (((!g1787) & (sk[12]) & (!g1788)) + ((g1787) & (!sk[12]) & (!g1788)) + ((g1787) & (!sk[12]) & (g1788)));
	assign g1787 = (((!g109) & (sk[13]) & (g1790)) + ((g109) & (!sk[13]) & (!g1790)) + ((g109) & (!sk[13]) & (g1790)));
	assign g1788 = (((!sk[14]) & (g109) & (!g1791)) + ((!sk[14]) & (g109) & (g1791)) + ((sk[14]) & (g109) & (g1791)));
	assign g1789 = (((!g96) & (!g133) & (g99) & (!sk[15]) & (g120)) + ((!g96) & (g133) & (!g99) & (!sk[15]) & (!g120)) + ((!g96) & (g133) & (!g99) & (!sk[15]) & (g120)) + ((!g96) & (g133) & (!g99) & (sk[15]) & (!g120)) + ((!g96) & (g133) & (!g99) & (sk[15]) & (g120)) + ((!g96) & (g133) & (g99) & (!sk[15]) & (!g120)) + ((!g96) & (g133) & (g99) & (!sk[15]) & (g120)) + ((g96) & (!g133) & (g99) & (!sk[15]) & (!g120)) + ((g96) & (!g133) & (g99) & (!sk[15]) & (g120)) + ((g96) & (g133) & (!g99) & (!sk[15]) & (!g120)) + ((g96) & (g133) & (!g99) & (!sk[15]) & (g120)) + ((g96) & (g133) & (!g99) & (sk[15]) & (!g120)) + ((g96) & (g133) & (!g99) & (sk[15]) & (g120)) + ((g96) & (g133) & (g99) & (!sk[15]) & (!g120)) + ((g96) & (g133) & (g99) & (!sk[15]) & (g120)) + ((g96) & (g133) & (g99) & (sk[15]) & (g120)));
	assign g1790 = (((!sk[16]) & (!g96) & (!g133) & (g99) & (g120)) + ((!sk[16]) & (!g96) & (g133) & (!g99) & (!g120)) + ((!sk[16]) & (!g96) & (g133) & (!g99) & (g120)) + ((!sk[16]) & (!g96) & (g133) & (g99) & (!g120)) + ((!sk[16]) & (!g96) & (g133) & (g99) & (g120)) + ((!sk[16]) & (g96) & (!g133) & (g99) & (!g120)) + ((!sk[16]) & (g96) & (!g133) & (g99) & (g120)) + ((!sk[16]) & (g96) & (g133) & (!g99) & (!g120)) + ((!sk[16]) & (g96) & (g133) & (!g99) & (g120)) + ((!sk[16]) & (g96) & (g133) & (g99) & (!g120)) + ((!sk[16]) & (g96) & (g133) & (g99) & (g120)) + ((sk[16]) & (!g96) & (g133) & (!g99) & (!g120)) + ((sk[16]) & (!g96) & (g133) & (!g99) & (g120)) + ((sk[16]) & (g96) & (g133) & (!g99) & (!g120)) + ((sk[16]) & (g96) & (g133) & (!g99) & (g120)) + ((sk[16]) & (g96) & (g133) & (g99) & (g120)));
	assign g1791 = (((!sk[17]) & (!g96) & (!g133) & (g103) & (g120)) + ((!sk[17]) & (!g96) & (g133) & (!g103) & (!g120)) + ((!sk[17]) & (!g96) & (g133) & (!g103) & (g120)) + ((!sk[17]) & (!g96) & (g133) & (g103) & (!g120)) + ((!sk[17]) & (!g96) & (g133) & (g103) & (g120)) + ((!sk[17]) & (g96) & (!g133) & (g103) & (!g120)) + ((!sk[17]) & (g96) & (!g133) & (g103) & (g120)) + ((!sk[17]) & (g96) & (g133) & (!g103) & (!g120)) + ((!sk[17]) & (g96) & (g133) & (!g103) & (g120)) + ((!sk[17]) & (g96) & (g133) & (g103) & (!g120)) + ((!sk[17]) & (g96) & (g133) & (g103) & (g120)) + ((sk[17]) & (g96) & (g133) & (g103) & (g120)));

endmodule