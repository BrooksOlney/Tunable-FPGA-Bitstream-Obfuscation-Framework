module des (
	Preset_0_, Poutreg_63_, Poutreg_62_, Poutreg_61_, Poutreg_60_, Poutreg_59_, Poutreg_58_, Poutreg_57_, 
	Poutreg_56_, Poutreg_55_, Poutreg_54_, Poutreg_53_, Poutreg_52_, Poutreg_51_, Poutreg_50_, Poutreg_49_, Poutreg_48_, Poutreg_47_, 
	Poutreg_46_, Poutreg_45_, Poutreg_44_, Poutreg_43_, Poutreg_42_, Poutreg_41_, Poutreg_40_, Poutreg_39_, Poutreg_38_, Poutreg_37_, 
	Poutreg_36_, Poutreg_35_, Poutreg_34_, Poutreg_33_, Poutreg_32_, Poutreg_31_, Poutreg_30_, Poutreg_29_, Poutreg_28_, Poutreg_27_, 
	Poutreg_26_, Poutreg_25_, Poutreg_24_, Poutreg_23_, Poutreg_22_, Poutreg_21_, Poutreg_20_, Poutreg_19_, Poutreg_18_, Poutreg_17_, 
	Poutreg_16_, Poutreg_15_, Poutreg_14_, Poutreg_13_, Poutreg_12_, Poutreg_11_, Poutreg_10_, Poutreg_9_, Poutreg_8_, Poutreg_7_, 
	Poutreg_6_, Poutreg_5_, Poutreg_4_, Poutreg_3_, Poutreg_2_, Poutreg_1_, Poutreg_0_, Pload_key_0_, Pinreg_55_, Pinreg_54_, 
	Pinreg_53_, Pinreg_52_, Pinreg_51_, Pinreg_50_, Pinreg_49_, Pinreg_48_, Pinreg_47_, Pinreg_46_, Pinreg_45_, Pinreg_44_, 
	Pinreg_43_, Pinreg_42_, Pinreg_41_, Pinreg_40_, Pinreg_39_, Pinreg_38_, Pinreg_37_, Pinreg_36_, Pinreg_35_, Pinreg_34_, 
	Pinreg_33_, Pinreg_32_, Pinreg_31_, Pinreg_30_, Pinreg_29_, Pinreg_28_, Pinreg_27_, Pinreg_26_, Pinreg_25_, Pinreg_24_, 
	Pinreg_23_, Pinreg_22_, Pinreg_21_, Pinreg_20_, Pinreg_19_, Pinreg_18_, Pinreg_17_, Pinreg_16_, Pinreg_15_, Pinreg_14_, 
	Pinreg_13_, Pinreg_12_, Pinreg_11_, Pinreg_10_, Pinreg_9_, Pinreg_8_, Pinreg_7_, Pinreg_6_, Pinreg_5_, Pinreg_4_, 
	Pinreg_3_, Pinreg_2_, Pinreg_1_, Pinreg_0_, Pencrypt_mode_0_, Pencrypt_0_, Pdata_in_7_, Pdata_in_6_, Pdata_in_5_, Pdata_in_4_, 
	Pdata_in_3_, Pdata_in_2_, Pdata_in_1_, Pdata_in_0_, Pdata_63_, Pdata_62_, Pdata_61_, Pdata_60_, Pdata_59_, Pdata_58_, 
	Pdata_57_, Pdata_56_, Pdata_55_, Pdata_54_, Pdata_53_, Pdata_52_, Pdata_51_, Pdata_50_, Pdata_49_, Pdata_48_, 
	Pdata_47_, Pdata_46_, Pdata_45_, Pdata_44_, Pdata_43_, Pdata_42_, Pdata_41_, Pdata_40_, Pdata_39_, Pdata_38_, 
	Pdata_37_, Pdata_36_, Pdata_35_, Pdata_34_, Pdata_33_, Pdata_32_, Pdata_31_, Pdata_30_, Pdata_29_, Pdata_28_, 
	Pdata_27_, Pdata_26_, Pdata_25_, Pdata_24_, Pdata_23_, Pdata_22_, Pdata_21_, Pdata_20_, Pdata_19_, Pdata_18_, 
	Pdata_17_, Pdata_16_, Pdata_15_, Pdata_14_, Pdata_13_, Pdata_12_, Pdata_11_, Pdata_10_, Pdata_9_, Pdata_8_, 
	Pdata_7_, Pdata_6_, Pdata_5_, Pdata_4_, Pdata_3_, Pdata_2_, Pdata_1_, Pdata_0_, Pcount_3_, Pcount_2_, 
	Pcount_1_, Pcount_0_, PD_27_, PD_26_, PD_25_, PD_24_, PD_23_, PD_22_, PD_21_, PD_20_, 
	PD_19_, PD_18_, PD_17_, PD_16_, PD_15_, PD_14_, PD_13_, PD_12_, PD_11_, PD_10_, 
	PD_9_, PD_8_, PD_7_, PD_6_, PD_5_, PD_4_, PD_3_, PD_2_, PD_1_, PD_0_, 
	PC_27_, PC_26_, PC_25_, PC_24_, PC_23_, PC_22_, PC_21_, PC_20_, PC_19_, PC_18_, 
	PC_17_, PC_16_, PC_15_, PC_14_, PC_13_, PC_12_, PC_11_, PC_10_, PC_9_, PC_8_, 
	PC_7_, PC_6_, PC_5_, PC_4_, PC_3_, PC_2_, PC_1_, PC_0_, Poutreg_new_63_, Poutreg_new_62_, 
	Poutreg_new_61_, Poutreg_new_60_, Poutreg_new_59_, Poutreg_new_58_, Poutreg_new_57_, Poutreg_new_56_, Poutreg_new_55_, Poutreg_new_54_, Poutreg_new_53_, Poutreg_new_52_, 
	Poutreg_new_51_, Poutreg_new_50_, Poutreg_new_49_, Poutreg_new_48_, Poutreg_new_47_, Poutreg_new_46_, Poutreg_new_45_, Poutreg_new_44_, Poutreg_new_43_, Poutreg_new_42_, 
	Poutreg_new_41_, Poutreg_new_40_, Poutreg_new_39_, Poutreg_new_38_, Poutreg_new_37_, Poutreg_new_36_, Poutreg_new_35_, Poutreg_new_34_, Poutreg_new_33_, Poutreg_new_32_, 
	Poutreg_new_31_, Poutreg_new_30_, Poutreg_new_29_, Poutreg_new_28_, Poutreg_new_27_, Poutreg_new_26_, Poutreg_new_25_, Poutreg_new_24_, Poutreg_new_23_, Poutreg_new_22_, 
	Poutreg_new_21_, Poutreg_new_20_, Poutreg_new_19_, Poutreg_new_18_, Poutreg_new_17_, Poutreg_new_16_, Poutreg_new_15_, Poutreg_new_14_, Poutreg_new_13_, Poutreg_new_12_, 
	Poutreg_new_11_, Poutreg_new_10_, Poutreg_new_9_, Poutreg_new_8_, Poutreg_new_7_, Poutreg_new_6_, Poutreg_new_5_, Poutreg_new_4_, Poutreg_new_3_, Poutreg_new_2_, 
	Poutreg_new_1_, Poutreg_new_0_, Pinreg_new_55_, Pinreg_new_54_, Pinreg_new_53_, Pinreg_new_52_, Pinreg_new_51_, Pinreg_new_50_, Pinreg_new_49_, Pinreg_new_48_, 
	Pinreg_new_47_, Pinreg_new_46_, Pinreg_new_45_, Pinreg_new_44_, Pinreg_new_43_, Pinreg_new_42_, Pinreg_new_41_, Pinreg_new_40_, Pinreg_new_39_, Pinreg_new_38_, 
	Pinreg_new_37_, Pinreg_new_36_, Pinreg_new_35_, Pinreg_new_34_, Pinreg_new_33_, Pinreg_new_32_, Pinreg_new_31_, Pinreg_new_30_, Pinreg_new_29_, Pinreg_new_28_, 
	Pinreg_new_27_, Pinreg_new_26_, Pinreg_new_25_, Pinreg_new_24_, Pinreg_new_23_, Pinreg_new_22_, Pinreg_new_21_, Pinreg_new_20_, Pinreg_new_19_, Pinreg_new_18_, 
	Pinreg_new_17_, Pinreg_new_16_, Pinreg_new_15_, Pinreg_new_14_, Pinreg_new_13_, Pinreg_new_12_, Pinreg_new_11_, Pinreg_new_10_, Pinreg_new_9_, Pinreg_new_8_, 
	Pinreg_new_7_, Pinreg_new_6_, Pinreg_new_5_, Pinreg_new_4_, Pinreg_new_3_, Pinreg_new_2_, Pinreg_new_1_, Pinreg_new_0_, Pencrypt_mode_new_0_, Pdata_new_63_, 
	Pdata_new_62_, Pdata_new_61_, Pdata_new_60_, Pdata_new_59_, Pdata_new_58_, Pdata_new_57_, Pdata_new_56_, Pdata_new_55_, Pdata_new_54_, Pdata_new_53_, 
	Pdata_new_52_, Pdata_new_51_, Pdata_new_50_, Pdata_new_49_, Pdata_new_48_, Pdata_new_47_, Pdata_new_46_, Pdata_new_45_, Pdata_new_44_, Pdata_new_43_, 
	Pdata_new_42_, Pdata_new_41_, Pdata_new_40_, Pdata_new_39_, Pdata_new_38_, Pdata_new_37_, Pdata_new_36_, Pdata_new_35_, Pdata_new_34_, Pdata_new_33_, 
	Pdata_new_32_, Pdata_new_31_, Pdata_new_30_, Pdata_new_29_, Pdata_new_28_, Pdata_new_27_, Pdata_new_26_, Pdata_new_25_, Pdata_new_24_, Pdata_new_23_, 
	Pdata_new_22_, Pdata_new_21_, Pdata_new_20_, Pdata_new_19_, Pdata_new_18_, Pdata_new_17_, Pdata_new_16_, Pdata_new_15_, Pdata_new_14_, Pdata_new_13_, 
	Pdata_new_12_, Pdata_new_11_, Pdata_new_10_, Pdata_new_9_, Pdata_new_8_, Pdata_new_7_, Pdata_new_6_, Pdata_new_5_, Pdata_new_4_, Pdata_new_3_, 
	Pdata_new_2_, Pdata_new_1_, Pdata_new_0_, Pcount_new_3_, Pcount_new_2_, Pcount_new_1_, Pcount_new_0_, PD_new_27_, PD_new_26_, PD_new_25_, 
	PD_new_24_, PD_new_23_, PD_new_22_, PD_new_21_, PD_new_20_, PD_new_19_, PD_new_18_, PD_new_17_, PD_new_16_, PD_new_15_, 
	PD_new_14_, PD_new_13_, PD_new_12_, PD_new_11_, PD_new_10_, PD_new_9_, PD_new_8_, PD_new_7_, PD_new_6_, PD_new_5_, 
	PD_new_4_, PD_new_3_, PD_new_2_, PD_new_1_, PD_new_0_, PC_new_27_, PC_new_26_, PC_new_25_, PC_new_24_, PC_new_23_, 
	PC_new_22_, PC_new_21_, PC_new_20_, PC_new_19_, PC_new_18_, PC_new_17_, PC_new_16_, PC_new_15_, PC_new_14_, PC_new_13_, 
	PC_new_12_, PC_new_11_, PC_new_10_, PC_new_9_, PC_new_8_, PC_new_7_, PC_new_6_, PC_new_5_, PC_new_4_, PC_new_3_, 
	PC_new_2_, PC_new_1_, PC_new_0_);

input Preset_0_, Poutreg_63_, Poutreg_62_, Poutreg_61_, Poutreg_60_, Poutreg_59_, Poutreg_58_, Poutreg_57_, Poutreg_56_, Poutreg_55_, Poutreg_54_, Poutreg_53_, Poutreg_52_, Poutreg_51_, Poutreg_50_, Poutreg_49_, Poutreg_48_, Poutreg_47_, Poutreg_46_, Poutreg_45_, Poutreg_44_, Poutreg_43_, Poutreg_42_, Poutreg_41_, Poutreg_40_, Poutreg_39_, Poutreg_38_, Poutreg_37_, Poutreg_36_, Poutreg_35_, Poutreg_34_, Poutreg_33_, Poutreg_32_, Poutreg_31_, Poutreg_30_, Poutreg_29_, Poutreg_28_, Poutreg_27_, Poutreg_26_, Poutreg_25_, Poutreg_24_, Poutreg_23_, Poutreg_22_, Poutreg_21_, Poutreg_20_, Poutreg_19_, Poutreg_18_, Poutreg_17_, Poutreg_16_, Poutreg_15_, Poutreg_14_, Poutreg_13_, Poutreg_12_, Poutreg_11_, Poutreg_10_, Poutreg_9_, Poutreg_8_, Poutreg_7_, Poutreg_6_, Poutreg_5_, Poutreg_4_, Poutreg_3_, Poutreg_2_, Poutreg_1_, Poutreg_0_, Pload_key_0_, Pinreg_55_, Pinreg_54_, Pinreg_53_, Pinreg_52_, Pinreg_51_, Pinreg_50_, Pinreg_49_, Pinreg_48_, Pinreg_47_, Pinreg_46_, Pinreg_45_, Pinreg_44_, Pinreg_43_, Pinreg_42_, Pinreg_41_, Pinreg_40_, Pinreg_39_, Pinreg_38_, Pinreg_37_, Pinreg_36_, Pinreg_35_, Pinreg_34_, Pinreg_33_, Pinreg_32_, Pinreg_31_, Pinreg_30_, Pinreg_29_, Pinreg_28_, Pinreg_27_, Pinreg_26_, Pinreg_25_, Pinreg_24_, Pinreg_23_, Pinreg_22_, Pinreg_21_, Pinreg_20_, Pinreg_19_, Pinreg_18_, Pinreg_17_, Pinreg_16_, Pinreg_15_, Pinreg_14_, Pinreg_13_, Pinreg_12_, Pinreg_11_, Pinreg_10_, Pinreg_9_, Pinreg_8_, Pinreg_7_, Pinreg_6_, Pinreg_5_, Pinreg_4_, Pinreg_3_, Pinreg_2_, Pinreg_1_, Pinreg_0_, Pencrypt_mode_0_, Pencrypt_0_, Pdata_in_7_, Pdata_in_6_, Pdata_in_5_, Pdata_in_4_, Pdata_in_3_, Pdata_in_2_, Pdata_in_1_, Pdata_in_0_, Pdata_63_, Pdata_62_, Pdata_61_, Pdata_60_, Pdata_59_, Pdata_58_, Pdata_57_, Pdata_56_, Pdata_55_, Pdata_54_, Pdata_53_, Pdata_52_, Pdata_51_, Pdata_50_, Pdata_49_, Pdata_48_, Pdata_47_, Pdata_46_, Pdata_45_, Pdata_44_, Pdata_43_, Pdata_42_, Pdata_41_, Pdata_40_, Pdata_39_, Pdata_38_, Pdata_37_, Pdata_36_, Pdata_35_, Pdata_34_, Pdata_33_, Pdata_32_, Pdata_31_, Pdata_30_, Pdata_29_, Pdata_28_, Pdata_27_, Pdata_26_, Pdata_25_, Pdata_24_, Pdata_23_, Pdata_22_, Pdata_21_, Pdata_20_, Pdata_19_, Pdata_18_, Pdata_17_, Pdata_16_, Pdata_15_, Pdata_14_, Pdata_13_, Pdata_12_, Pdata_11_, Pdata_10_, Pdata_9_, Pdata_8_, Pdata_7_, Pdata_6_, Pdata_5_, Pdata_4_, Pdata_3_, Pdata_2_, Pdata_1_, Pdata_0_, Pcount_3_, Pcount_2_, Pcount_1_, Pcount_0_, PD_27_, PD_26_, PD_25_, PD_24_, PD_23_, PD_22_, PD_21_, PD_20_, PD_19_, PD_18_, PD_17_, PD_16_, PD_15_, PD_14_, PD_13_, PD_12_, PD_11_, PD_10_, PD_9_, PD_8_, PD_7_, PD_6_, PD_5_, PD_4_, PD_3_, PD_2_, PD_1_, PD_0_, PC_27_, PC_26_, PC_25_, PC_24_, PC_23_, PC_22_, PC_21_, PC_20_, PC_19_, PC_18_, PC_17_, PC_16_, PC_15_, PC_14_, PC_13_, PC_12_, PC_11_, PC_10_, PC_9_, PC_8_, PC_7_, PC_6_, PC_5_, PC_4_, PC_3_, PC_2_, PC_1_, PC_0_;

output Poutreg_new_63_, Poutreg_new_62_, Poutreg_new_61_, Poutreg_new_60_, Poutreg_new_59_, Poutreg_new_58_, Poutreg_new_57_, Poutreg_new_56_, Poutreg_new_55_, Poutreg_new_54_, Poutreg_new_53_, Poutreg_new_52_, Poutreg_new_51_, Poutreg_new_50_, Poutreg_new_49_, Poutreg_new_48_, Poutreg_new_47_, Poutreg_new_46_, Poutreg_new_45_, Poutreg_new_44_, Poutreg_new_43_, Poutreg_new_42_, Poutreg_new_41_, Poutreg_new_40_, Poutreg_new_39_, Poutreg_new_38_, Poutreg_new_37_, Poutreg_new_36_, Poutreg_new_35_, Poutreg_new_34_, Poutreg_new_33_, Poutreg_new_32_, Poutreg_new_31_, Poutreg_new_30_, Poutreg_new_29_, Poutreg_new_28_, Poutreg_new_27_, Poutreg_new_26_, Poutreg_new_25_, Poutreg_new_24_, Poutreg_new_23_, Poutreg_new_22_, Poutreg_new_21_, Poutreg_new_20_, Poutreg_new_19_, Poutreg_new_18_, Poutreg_new_17_, Poutreg_new_16_, Poutreg_new_15_, Poutreg_new_14_, Poutreg_new_13_, Poutreg_new_12_, Poutreg_new_11_, Poutreg_new_10_, Poutreg_new_9_, Poutreg_new_8_, Poutreg_new_7_, Poutreg_new_6_, Poutreg_new_5_, Poutreg_new_4_, Poutreg_new_3_, Poutreg_new_2_, Poutreg_new_1_, Poutreg_new_0_, Pinreg_new_55_, Pinreg_new_54_, Pinreg_new_53_, Pinreg_new_52_, Pinreg_new_51_, Pinreg_new_50_, Pinreg_new_49_, Pinreg_new_48_, Pinreg_new_47_, Pinreg_new_46_, Pinreg_new_45_, Pinreg_new_44_, Pinreg_new_43_, Pinreg_new_42_, Pinreg_new_41_, Pinreg_new_40_, Pinreg_new_39_, Pinreg_new_38_, Pinreg_new_37_, Pinreg_new_36_, Pinreg_new_35_, Pinreg_new_34_, Pinreg_new_33_, Pinreg_new_32_, Pinreg_new_31_, Pinreg_new_30_, Pinreg_new_29_, Pinreg_new_28_, Pinreg_new_27_, Pinreg_new_26_, Pinreg_new_25_, Pinreg_new_24_, Pinreg_new_23_, Pinreg_new_22_, Pinreg_new_21_, Pinreg_new_20_, Pinreg_new_19_, Pinreg_new_18_, Pinreg_new_17_, Pinreg_new_16_, Pinreg_new_15_, Pinreg_new_14_, Pinreg_new_13_, Pinreg_new_12_, Pinreg_new_11_, Pinreg_new_10_, Pinreg_new_9_, Pinreg_new_8_, Pinreg_new_7_, Pinreg_new_6_, Pinreg_new_5_, Pinreg_new_4_, Pinreg_new_3_, Pinreg_new_2_, Pinreg_new_1_, Pinreg_new_0_, Pencrypt_mode_new_0_, Pdata_new_63_, Pdata_new_62_, Pdata_new_61_, Pdata_new_60_, Pdata_new_59_, Pdata_new_58_, Pdata_new_57_, Pdata_new_56_, Pdata_new_55_, Pdata_new_54_, Pdata_new_53_, Pdata_new_52_, Pdata_new_51_, Pdata_new_50_, Pdata_new_49_, Pdata_new_48_, Pdata_new_47_, Pdata_new_46_, Pdata_new_45_, Pdata_new_44_, Pdata_new_43_, Pdata_new_42_, Pdata_new_41_, Pdata_new_40_, Pdata_new_39_, Pdata_new_38_, Pdata_new_37_, Pdata_new_36_, Pdata_new_35_, Pdata_new_34_, Pdata_new_33_, Pdata_new_32_, Pdata_new_31_, Pdata_new_30_, Pdata_new_29_, Pdata_new_28_, Pdata_new_27_, Pdata_new_26_, Pdata_new_25_, Pdata_new_24_, Pdata_new_23_, Pdata_new_22_, Pdata_new_21_, Pdata_new_20_, Pdata_new_19_, Pdata_new_18_, Pdata_new_17_, Pdata_new_16_, Pdata_new_15_, Pdata_new_14_, Pdata_new_13_, Pdata_new_12_, Pdata_new_11_, Pdata_new_10_, Pdata_new_9_, Pdata_new_8_, Pdata_new_7_, Pdata_new_6_, Pdata_new_5_, Pdata_new_4_, Pdata_new_3_, Pdata_new_2_, Pdata_new_1_, Pdata_new_0_, Pcount_new_3_, Pcount_new_2_, Pcount_new_1_, Pcount_new_0_, PD_new_27_, PD_new_26_, PD_new_25_, PD_new_24_, PD_new_23_, PD_new_22_, PD_new_21_, PD_new_20_, PD_new_19_, PD_new_18_, PD_new_17_, PD_new_16_, PD_new_15_, PD_new_14_, PD_new_13_, PD_new_12_, PD_new_11_, PD_new_10_, PD_new_9_, PD_new_8_, PD_new_7_, PD_new_6_, PD_new_5_, PD_new_4_, PD_new_3_, PD_new_2_, PD_new_1_, PD_new_0_, PC_new_27_, PC_new_26_, PC_new_25_, PC_new_24_, PC_new_23_, PC_new_22_, PC_new_21_, PC_new_20_, PC_new_19_, PC_new_18_, PC_new_17_, PC_new_16_, PC_new_15_, PC_new_14_, PC_new_13_, PC_new_12_, PC_new_11_, PC_new_10_, PC_new_9_, PC_new_8_, PC_new_7_, PC_new_6_, PC_new_5_, PC_new_4_, PC_new_3_, PC_new_2_, PC_new_1_, PC_new_0_;

wire n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n126, n191, n196, n201, n199, n204, n202, n209, n208, n207, n205, n214, n212, n210, n217, n218, n216, n215, n220, n222, n219, n224, n223, n228, n227, n226, n225, n230, n231, n229, n234, n243, n240, n239, n244, n252, n249, n254, n253, n259, n260, n257, n263, n262, n261, n266, n264, n269, n268, n272, n270, n275, n274, n273, n276, n279, n278, n281, n280, n283, n285, n282, n287, n292, n291, n294, n295, n293, n299, n297, n296, n300, n304, n305, n303, n301, n307, n308, n306, n309, n314, n315, n317, n313, n321, n319, n318, n323, n325, n326, n322, n329, n328, n327, n331, n334, n335, n333, n339, n337, n336, n341, n342, n343, n340, n345, n344, n346, n351, n352, n350, n357, n355, n353, n359, n358, n360, n365, n367, n371, n369, n368, n373, n372, n375, n377, n374, n382, n380, n378, n386, n387, n384, n385, n383, n389, n392, n388, n395, n396, n393, n398, n399, n397, n401, n400, n405, n406, n403, n404, n402, n409, n410, n408, n407, n412, n414, n416, n417, n415, n421, n420, n418, n423, n424, n425, n426, n422, n428, n430, n432, n431, n436, n434, n433, n438, n437, n441, n442, n439, n447, n444, n445, n443, n449, n450, n448, n452, n453, n451, n455, n457, n459, n460, n461, n458, n464, n463, n462, n467, n468, n466, n470, n471, n472, n473, n469, n475, n476, n477, n474, n480, n481, n479, n483, n482, n484, n487, n491, n489, n495, n493, n497, n498, n499, n500, n501, n502, n503, n496, n505, n507, n511, n510, n508, n515, n513, n512, n519, n520, n517, n516, n523, n522, n521, n527, n528, n525, n526, n524, n532, n531, n529, n534, n535, n536, n533, n538, n540, n544, n542, n543, n541, n549, n546, n545, n551, n553, n556, n557, n554, n559, n558, n561, n560, n564, n566, n570, n569, n567, n572, n571, n574, n573, n576, n577, n578, n575, n580, n582, n585, n583, n588, n587, n591, n590, n594, n593, n596, n598, n602, n600, n599, n607, n604, n605, n603, n612, n609, n608, n615, n613, n620, n621, n618, n622, n626, n627, n625, n631, n632, n629, n628, n634, n635, n636, n637, n633, n639, n641, n642, n648, n647, n646, n650, n652, n655, n656, n654, n653, n659, n660, n658, n657, n662, n663, n661, n665, n667, n671, n672, n670, n668, n675, n673, n678, n679, n676, n681, n682, n683, n684, n685, n680, n687, n689, n691, n692, n690, n694, n695, n696, n693, n698, n700, n702, n703, n704, n701, n706, n708, n710, n711, n709, n716, n717, n714, n722, n721, n719, n720, n718, n727, n724, n725, n723, n729, n730, n728, n732, n731, n735, n738, n740, n737, n744, n745, n742, n743, n741, n748, n746, n751, n749, n754, n752, n756, n755, n759, n757, n760, n762, n764, n766, n765, n769, n773, n772, n771, n777, n775, n776, n774, n780, n781, n779, n783, n785, n786, n789, n788, n790, n795, n794, n797, n799, n802, n803, n801, n800, n806, n804, n808, n809, n811, n810, n814, n813, n817, n816, n819, n821, n824, n822, n827, n829, n826, n831, n833, n835, n834, n837, n838, n839, n841, n836, n843, n845, n847, n846, n849, n848, n851, n852, n850, n855, n857, n858, n859, n862, n863, n860, n866, n864, n869, n871, n874, n875, n873, n872, n877, n878, n876, n879, n880, n884, n886, n888, n887, n889, n891, n893, n896, n895, n894, n898, n897, n901, n902, n903, n904, n905, n900, n907, n909, n912, n911, n910, n914, n915, n913, n917, n920, n922, n925, n924, n923, n926, n928, n929, n932, n933, n934, n931, n936, n937, n938, n935, n940, n941, n942, n939, n944, n945, n946, n943, n948, n949, n950, n947, n952, n953, n954, n951, n956, n957, n958, n955, n960, n961, n962, n959, n964, n965, n966, n963, n968, n969, n970, n967, n972, n973, n974, n971, n976, n977, n978, n975, n980, n981, n982, n979, n984, n985, n986, n983, n988, n989, n990, n987, n992, n993, n994, n991, n996, n997, n998, n995, n1000, n1001, n1002, n999, n1004, n1005, n1006, n1003, n1008, n1009, n1010, n1007, n1012, n1013, n1014, n1011, n1016, n1017, n1018, n1015, n1020, n1021, n1022, n1019, n1024, n1025, n1026, n1023, n1028, n1029, n1030, n1027, n1032, n1033, n1034, n1031, n1036, n1037, n1038, n1035, n1040, n1041, n1042, n1039, n1044, n1045, n1046, n1043, n1048, n1049, n1050, n1047, n1052, n1053, n1054, n1051, n1056, n1057, n1058, n1055, n1060, n1061, n1062, n1059, n1064, n1065, n1066, n1063, n1068, n1069, n1070, n1067, n1072, n1073, n1074, n1071, n1076, n1077, n1078, n1075, n1080, n1081, n1082, n1079, n1084, n1085, n1086, n1083, n1088, n1089, n1090, n1087, n1092, n1093, n1094, n1091, n1096, n1097, n1098, n1095, n1100, n1101, n1102, n1099, n1104, n1105, n1106, n1103, n1108, n1109, n1110, n1107, n1112, n1113, n1114, n1111, n1116, n1117, n1118, n1115, n1120, n1121, n1122, n1119, n1124, n1125, n1126, n1123, n1128, n1129, n1130, n1127, n1132, n1133, n1134, n1131, n1136, n1137, n1138, n1135, n1140, n1141, n1142, n1139, n1144, n1145, n1146, n1143, n1148, n1149, n1150, n1147, n1152, n1153, n1154, n1151, n1155, n1156, n1158, n1159, n1160, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1172, n1173, n1177, n1184, n1185, n1186, n1187, n1188, n1189, n1198, n1199, n1200, n1201, n1202, n1204, n1205, n1203, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1232, n1234, n1246, n1248, n1249, n1250, n1251, n1252, n1254, n1257, n1258, n1265, n1270, n1272, n1273, n1274, n1275, n1281, n1289, n1292, n1293, n1295, n1297, n1298, n1300, n1301, n1303, n1318, n1319, n1321, n1323, n1324, n1325, n1326, n1329, n1340, n1341, n1345, n1347, n1348, n1350, n1351, n1352, n1353, n1354, n1356, n1357, n1358, n1359, n1369, n1371, n1372, n1373, n1375, n1376, n1378, n1380, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1457, n1458, n1459, n1464, n1465, n1466, n1468, n1470, n1469, n1471, n1472, n1473, n1475, n1474, n1476, n1477, n1478, n1479, n1480, n1482, n1483, n1486, n1484, n1487, n1488, n1489, n1490, n1493, n1492, n1494, n1495, n1497, n1496, n1499, n1500, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1514, n1515, n1516, n1517, n1520, n1518, n1521, n1522, n1524, n1525, n1528, n1529, n1530, n1532, n1533, n1534, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1602, n1604, n1605, n1607, n1609, n1610, n1611, n1614, n1615, n1616, n1617, n1619, n1620, n1622, n1621, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1633, n1632, n1635, n1636, n1638, n1639, n1640, n1641, n1642, n1643, n1645, n1647, n1648, n1649, n1651, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1663, n1664, n1665, n1666, n1668, n1669, n1672, n1675, n1678, n1680, n1683, n1684, n1688, n1690, n1692, n1695, n1698, n1702, n1703, n1706, n1709, n1711, n1714, n1717, n1718, n1719;

assign Poutreg_new_63_ = ( (~ n2) ) ;
 assign Poutreg_new_62_ = ( (~ n105) ) ;
 assign Poutreg_new_61_ = ( (~ n3) ) ;
 assign Poutreg_new_60_ = ( (~ n101) ) ;
 assign Poutreg_new_59_ = ( (~ n4) ) ;
 assign Poutreg_new_58_ = ( (~ n97) ) ;
 assign Poutreg_new_57_ = ( (~ n5) ) ;
 assign Poutreg_new_56_ = ( (~ n91) ) ;
 assign Poutreg_new_55_ = ( (~ n6) ) ;
 assign Poutreg_new_54_ = ( (~ n124) ) ;
 assign Poutreg_new_53_ = ( (~ n7) ) ;
 assign Poutreg_new_52_ = ( (~ n94) ) ;
 assign Poutreg_new_51_ = ( (~ n8) ) ;
 assign Poutreg_new_50_ = ( (~ n123) ) ;
 assign Poutreg_new_49_ = ( (~ n9) ) ;
 assign Poutreg_new_48_ = ( (~ n122) ) ;
 assign Poutreg_new_47_ = ( (~ n10) ) ;
 assign Poutreg_new_46_ = ( (~ n121) ) ;
 assign Poutreg_new_45_ = ( (~ n11) ) ;
 assign Poutreg_new_44_ = ( (~ n120) ) ;
 assign Poutreg_new_43_ = ( (~ n12) ) ;
 assign Poutreg_new_42_ = ( (~ n119) ) ;
 assign Poutreg_new_41_ = ( (~ n13) ) ;
 assign Poutreg_new_40_ = ( (~ n118) ) ;
 assign Poutreg_new_39_ = ( (~ n14) ) ;
 assign Poutreg_new_38_ = ( (~ n117) ) ;
 assign Poutreg_new_37_ = ( (~ n15) ) ;
 assign Poutreg_new_36_ = ( (~ n116) ) ;
 assign Poutreg_new_35_ = ( (~ n16) ) ;
 assign Poutreg_new_34_ = ( (~ n115) ) ;
 assign Poutreg_new_33_ = ( (~ n17) ) ;
 assign Poutreg_new_32_ = ( (~ n114) ) ;
 assign Poutreg_new_31_ = ( (~ n18) ) ;
 assign Poutreg_new_30_ = ( (~ n113) ) ;
 assign Poutreg_new_29_ = ( (~ n19) ) ;
 assign Poutreg_new_28_ = ( (~ n112) ) ;
 assign Poutreg_new_27_ = ( (~ n20) ) ;
 assign Poutreg_new_26_ = ( (~ n111) ) ;
 assign Poutreg_new_25_ = ( (~ n21) ) ;
 assign Poutreg_new_24_ = ( (~ n110) ) ;
 assign Poutreg_new_23_ = ( (~ n22) ) ;
 assign Poutreg_new_22_ = ( (~ n109) ) ;
 assign Poutreg_new_21_ = ( (~ n23) ) ;
 assign Poutreg_new_20_ = ( (~ n108) ) ;
 assign Poutreg_new_19_ = ( (~ n24) ) ;
 assign Poutreg_new_18_ = ( (~ n107) ) ;
 assign Poutreg_new_17_ = ( (~ n25) ) ;
 assign Poutreg_new_16_ = ( (~ n106) ) ;
 assign Poutreg_new_15_ = ( (~ n26) ) ;
 assign Poutreg_new_14_ = ( (~ n104) ) ;
 assign Poutreg_new_13_ = ( (~ n27) ) ;
 assign Poutreg_new_12_ = ( (~ n103) ) ;
 assign Poutreg_new_11_ = ( (~ n28) ) ;
 assign Poutreg_new_10_ = ( (~ n102) ) ;
 assign Poutreg_new_9_ = ( (~ n29) ) ;
 assign Poutreg_new_8_ = ( (~ n100) ) ;
 assign Poutreg_new_7_ = ( (~ n30) ) ;
 assign Poutreg_new_6_ = ( (~ n99) ) ;
 assign Poutreg_new_5_ = ( (~ n31) ) ;
 assign Poutreg_new_4_ = ( (~ n98) ) ;
 assign Poutreg_new_3_ = ( (~ n32) ) ;
 assign Poutreg_new_2_ = ( (~ n96) ) ;
 assign Poutreg_new_1_ = ( (~ n33) ) ;
 assign Poutreg_new_0_ = ( (~ n95) ) ;
 assign Pinreg_new_55_ = ( (~ n35) ) ;
 assign Pinreg_new_54_ = ( (~ n36) ) ;
 assign Pinreg_new_53_ = ( (~ n37) ) ;
 assign Pinreg_new_52_ = ( (~ n38) ) ;
 assign Pinreg_new_51_ = ( (~ n39) ) ;
 assign Pinreg_new_50_ = ( (~ n40) ) ;
 assign Pinreg_new_49_ = ( (~ n41) ) ;
 assign Pinreg_new_48_ = ( (~ n42) ) ;
 assign Pinreg_new_47_ = ( (~ n43) ) ;
 assign Pinreg_new_46_ = ( (~ n44) ) ;
 assign Pinreg_new_45_ = ( (~ n45) ) ;
 assign Pinreg_new_44_ = ( (~ n46) ) ;
 assign Pinreg_new_43_ = ( (~ n47) ) ;
 assign Pinreg_new_42_ = ( (~ n48) ) ;
 assign Pinreg_new_41_ = ( (~ n49) ) ;
 assign Pinreg_new_40_ = ( (~ n50) ) ;
 assign Pinreg_new_39_ = ( (~ n51) ) ;
 assign Pinreg_new_38_ = ( (~ n52) ) ;
 assign Pinreg_new_37_ = ( (~ n53) ) ;
 assign Pinreg_new_36_ = ( (~ n54) ) ;
 assign Pinreg_new_35_ = ( (~ n55) ) ;
 assign Pinreg_new_34_ = ( (~ n56) ) ;
 assign Pinreg_new_33_ = ( (~ n57) ) ;
 assign Pinreg_new_32_ = ( (~ n58) ) ;
 assign Pinreg_new_31_ = ( (~ n59) ) ;
 assign Pinreg_new_30_ = ( (~ n60) ) ;
 assign Pinreg_new_29_ = ( (~ n61) ) ;
 assign Pinreg_new_28_ = ( (~ n62) ) ;
 assign Pinreg_new_27_ = ( (~ n63) ) ;
 assign Pinreg_new_26_ = ( (~ n64) ) ;
 assign Pinreg_new_25_ = ( (~ n65) ) ;
 assign Pinreg_new_24_ = ( (~ n66) ) ;
 assign Pinreg_new_23_ = ( (~ n67) ) ;
 assign Pinreg_new_22_ = ( (~ n68) ) ;
 assign Pinreg_new_21_ = ( (~ n69) ) ;
 assign Pinreg_new_20_ = ( (~ n70) ) ;
 assign Pinreg_new_19_ = ( (~ n71) ) ;
 assign Pinreg_new_18_ = ( (~ n72) ) ;
 assign Pinreg_new_17_ = ( (~ n73) ) ;
 assign Pinreg_new_16_ = ( (~ n74) ) ;
 assign Pinreg_new_15_ = ( (~ n75) ) ;
 assign Pinreg_new_14_ = ( (~ n76) ) ;
 assign Pinreg_new_13_ = ( (~ n77) ) ;
 assign Pinreg_new_12_ = ( (~ n78) ) ;
 assign Pinreg_new_11_ = ( (~ n79) ) ;
 assign Pinreg_new_10_ = ( (~ n80) ) ;
 assign Pinreg_new_9_ = ( (~ n81) ) ;
 assign Pinreg_new_8_ = ( (~ n82) ) ;
 assign Pinreg_new_7_ = ( (~ n83) ) ;
 assign Pinreg_new_6_ = ( (~ n84) ) ;
 assign Pinreg_new_5_ = ( (~ n85) ) ;
 assign Pinreg_new_4_ = ( (~ n86) ) ;
 assign Pinreg_new_3_ = ( (~ n87) ) ;
 assign Pinreg_new_2_ = ( (~ n88) ) ;
 assign Pinreg_new_1_ = ( (~ n89) ) ;
 assign Pinreg_new_0_ = ( (~ n90) ) ;
 assign Pencrypt_mode_new_0_ = ( (~ n1454) ) ;
 assign Pdata_new_63_ = ( (~ n1387) ) ;
 assign Pdata_new_62_ = ( (~ n1388) ) ;
 assign Pdata_new_61_ = ( (~ n1389) ) ;
 assign Pdata_new_60_ = ( (~ n1390) ) ;
 assign Pdata_new_59_ = ( (~ n1391) ) ;
 assign Pdata_new_58_ = ( (~ n1392) ) ;
 assign Pdata_new_57_ = ( (~ n1393) ) ;
 assign Pdata_new_56_ = ( (~ n1394) ) ;
 assign Pdata_new_55_ = ( (~ n1395) ) ;
 assign Pdata_new_54_ = ( (~ n1396) ) ;
 assign Pdata_new_53_ = ( (~ n1397) ) ;
 assign Pdata_new_52_ = ( (~ n1398) ) ;
 assign Pdata_new_51_ = ( (~ n1399) ) ;
 assign Pdata_new_50_ = ( (~ n1400) ) ;
 assign Pdata_new_49_ = ( (~ n1401) ) ;
 assign Pdata_new_48_ = ( (~ n1402) ) ;
 assign Pdata_new_47_ = ( (~ n1403) ) ;
 assign Pdata_new_46_ = ( (~ n1404) ) ;
 assign Pdata_new_45_ = ( (~ n1405) ) ;
 assign Pdata_new_44_ = ( (~ n1406) ) ;
 assign Pdata_new_43_ = ( (~ n1407) ) ;
 assign Pdata_new_42_ = ( (~ n1408) ) ;
 assign Pdata_new_41_ = ( (~ n1409) ) ;
 assign Pdata_new_40_ = ( (~ n1410) ) ;
 assign Pdata_new_39_ = ( (~ n1411) ) ;
 assign Pdata_new_38_ = ( (~ n1412) ) ;
 assign Pdata_new_37_ = ( (~ n1413) ) ;
 assign Pdata_new_36_ = ( (~ n1414) ) ;
 assign Pdata_new_35_ = ( (~ n1415) ) ;
 assign Pdata_new_34_ = ( (~ n1416) ) ;
 assign Pdata_new_33_ = ( (~ n1417) ) ;
 assign Pdata_new_32_ = ( (~ n1418) ) ;
 assign Pdata_new_31_ = ( (~ n1419) ) ;
 assign Pdata_new_30_ = ( (~ n1420) ) ;
 assign Pdata_new_29_ = ( (~ n1421) ) ;
 assign Pdata_new_28_ = ( (~ n1422) ) ;
 assign Pdata_new_27_ = ( (~ n1423) ) ;
 assign Pdata_new_26_ = ( (~ n1424) ) ;
 assign Pdata_new_25_ = ( (~ n1425) ) ;
 assign Pdata_new_24_ = ( (~ n1426) ) ;
 assign Pdata_new_23_ = ( (~ n1427) ) ;
 assign Pdata_new_22_ = ( (~ n1428) ) ;
 assign Pdata_new_21_ = ( (~ n1429) ) ;
 assign Pdata_new_20_ = ( (~ n1430) ) ;
 assign Pdata_new_19_ = ( (~ n1431) ) ;
 assign Pdata_new_18_ = ( (~ n1432) ) ;
 assign Pdata_new_17_ = ( (~ n1433) ) ;
 assign Pdata_new_16_ = ( (~ n1434) ) ;
 assign Pdata_new_15_ = ( (~ n1435) ) ;
 assign Pdata_new_14_ = ( (~ n1436) ) ;
 assign Pdata_new_13_ = ( (~ n1437) ) ;
 assign Pdata_new_12_ = ( (~ n1438) ) ;
 assign Pdata_new_11_ = ( (~ n1439) ) ;
 assign Pdata_new_10_ = ( (~ n1440) ) ;
 assign Pdata_new_9_ = ( (~ n1441) ) ;
 assign Pdata_new_8_ = ( (~ n1442) ) ;
 assign Pdata_new_7_ = ( (~ n1443) ) ;
 assign Pdata_new_6_ = ( (~ n1444) ) ;
 assign Pdata_new_5_ = ( (~ n1445) ) ;
 assign Pdata_new_4_ = ( (~ n1446) ) ;
 assign Pdata_new_3_ = ( (~ n1447) ) ;
 assign Pdata_new_2_ = ( (~ n1448) ) ;
 assign Pdata_new_1_ = ( (~ n1449) ) ;
 assign Pdata_new_0_ = ( (~ n1450) ) ;
 assign Pcount_new_3_ = ( (~ n34) ) ;
 assign Pcount_new_2_ = ( (~ n1451) ) ;
 assign Pcount_new_1_ = ( (~ n1452) ) ;
 assign Pcount_new_0_ = ( (~ n925) ) ;
 assign PD_new_27_ = ( (~ n1043) ) ;
 assign PD_new_26_ = ( (~ n1047) ) ;
 assign PD_new_25_ = ( (~ n1051) ) ;
 assign PD_new_24_ = ( (~ n1055) ) ;
 assign PD_new_23_ = ( (~ n1059) ) ;
 assign PD_new_22_ = ( (~ n1063) ) ;
 assign PD_new_21_ = ( (~ n1067) ) ;
 assign PD_new_20_ = ( (~ n1071) ) ;
 assign PD_new_19_ = ( (~ n1075) ) ;
 assign PD_new_18_ = ( (~ n1079) ) ;
 assign PD_new_17_ = ( (~ n1083) ) ;
 assign PD_new_16_ = ( (~ n1087) ) ;
 assign PD_new_15_ = ( (~ n1091) ) ;
 assign PD_new_14_ = ( (~ n1095) ) ;
 assign PD_new_13_ = ( (~ n1099) ) ;
 assign PD_new_12_ = ( (~ n1103) ) ;
 assign PD_new_11_ = ( (~ n1107) ) ;
 assign PD_new_10_ = ( (~ n1111) ) ;
 assign PD_new_9_ = ( (~ n1115) ) ;
 assign PD_new_8_ = ( (~ n1119) ) ;
 assign PD_new_7_ = ( (~ n1123) ) ;
 assign PD_new_6_ = ( (~ n1127) ) ;
 assign PD_new_5_ = ( (~ n1131) ) ;
 assign PD_new_4_ = ( (~ n1135) ) ;
 assign PD_new_3_ = ( (~ n1139) ) ;
 assign PD_new_2_ = ( (~ n1143) ) ;
 assign PD_new_1_ = ( (~ n1147) ) ;
 assign PD_new_0_ = ( (~ n1151) ) ;
 assign PC_new_27_ = ( (~ n931) ) ;
 assign PC_new_26_ = ( (~ n935) ) ;
 assign PC_new_25_ = ( (~ n939) ) ;
 assign PC_new_24_ = ( (~ n943) ) ;
 assign PC_new_23_ = ( (~ n947) ) ;
 assign PC_new_22_ = ( (~ n951) ) ;
 assign PC_new_21_ = ( (~ n955) ) ;
 assign PC_new_20_ = ( (~ n959) ) ;
 assign PC_new_19_ = ( (~ n963) ) ;
 assign PC_new_18_ = ( (~ n967) ) ;
 assign PC_new_17_ = ( (~ n971) ) ;
 assign PC_new_16_ = ( (~ n975) ) ;
 assign PC_new_15_ = ( (~ n979) ) ;
 assign PC_new_14_ = ( (~ n983) ) ;
 assign PC_new_13_ = ( (~ n987) ) ;
 assign PC_new_12_ = ( (~ n991) ) ;
 assign PC_new_11_ = ( (~ n995) ) ;
 assign PC_new_10_ = ( (~ n999) ) ;
 assign PC_new_9_ = ( (~ n1003) ) ;
 assign PC_new_8_ = ( (~ n1007) ) ;
 assign PC_new_7_ = ( (~ n1011) ) ;
 assign PC_new_6_ = ( (~ n1015) ) ;
 assign PC_new_5_ = ( (~ n1019) ) ;
 assign PC_new_4_ = ( (~ n1023) ) ;
 assign PC_new_3_ = ( (~ n1027) ) ;
 assign PC_new_2_ = ( (~ n1031) ) ;
 assign PC_new_1_ = ( (~ n1035) ) ;
 assign PC_new_0_ = ( (~ n1039) ) ;
 assign n1 = ( (~ Pcount_3_) ) | ( n1177 ) ;
 assign n2 = ( (~ Poutreg_63_)  &  n1 ) | ( Pcount_0_  &  n1 ) | ( (~ Poutreg_63_)  &  n234 ) | ( Pcount_0_  &  n234 ) ;
 assign n3 = ( (~ Poutreg_61_)  &  n1 ) | ( Pcount_0_  &  n1 ) | ( (~ Poutreg_61_)  &  n287 ) | ( Pcount_0_  &  n287 ) ;
 assign n4 = ( (~ Poutreg_59_)  &  n1 ) | ( Pcount_0_  &  n1 ) | ( (~ Poutreg_59_)  &  n309 ) | ( Pcount_0_  &  n309 ) ;
 assign n5 = ( (~ Poutreg_57_)  &  n1 ) | ( Pcount_0_  &  n1 ) | ( (~ Poutreg_57_)  &  n346 ) | ( Pcount_0_  &  n346 ) ;
 assign n6 = ( (~ Poutreg_55_)  &  n365 ) | ( Pcount_0_  &  n365 ) ;
 assign n7 = ( (~ Poutreg_53_)  &  n412 ) | ( Pcount_0_  &  n412 ) ;
 assign n8 = ( (~ Poutreg_51_)  &  n428 ) | ( Pcount_0_  &  n428 ) ;
 assign n9 = ( (~ Poutreg_49_)  &  n455 ) | ( Pcount_0_  &  n455 ) ;
 assign n10 = ( (~ Poutreg_47_)  &  n505 ) | ( Pcount_0_  &  n505 ) ;
 assign n11 = ( (~ Poutreg_45_)  &  n538 ) | ( Pcount_0_  &  n538 ) ;
 assign n12 = ( (~ Poutreg_43_)  &  n551 ) | ( Pcount_0_  &  n551 ) ;
 assign n13 = ( (~ Poutreg_41_)  &  n564 ) | ( Pcount_0_  &  n564 ) ;
 assign n14 = ( (~ Poutreg_39_)  &  n580 ) | ( Pcount_0_  &  n580 ) ;
 assign n15 = ( (~ Poutreg_37_)  &  n596 ) | ( Pcount_0_  &  n596 ) ;
 assign n16 = ( (~ Poutreg_35_)  &  n639 ) | ( Pcount_0_  &  n639 ) ;
 assign n17 = ( (~ Poutreg_33_)  &  n650 ) | ( Pcount_0_  &  n650 ) ;
 assign n18 = ( (~ Poutreg_31_)  &  n665 ) | ( Pcount_0_  &  n665 ) ;
 assign n19 = ( (~ Poutreg_29_)  &  n687 ) | ( Pcount_0_  &  n687 ) ;
 assign n20 = ( (~ Poutreg_27_)  &  n698 ) | ( Pcount_0_  &  n698 ) ;
 assign n21 = ( (~ Poutreg_25_)  &  n706 ) | ( Pcount_0_  &  n706 ) ;
 assign n22 = ( (~ Poutreg_23_)  &  n762 ) | ( Pcount_0_  &  n762 ) ;
 assign n23 = ( (~ Poutreg_21_)  &  n783 ) | ( Pcount_0_  &  n783 ) ;
 assign n24 = ( (~ Poutreg_19_)  &  n797 ) | ( Pcount_0_  &  n797 ) ;
 assign n25 = ( (~ Poutreg_17_)  &  n819 ) | ( Pcount_0_  &  n819 ) ;
 assign n26 = ( (~ Poutreg_15_)  &  n831 ) | ( Pcount_0_  &  n831 ) ;
 assign n27 = ( (~ Poutreg_13_)  &  n843 ) | ( Pcount_0_  &  n843 ) ;
 assign n28 = ( (~ Poutreg_11_)  &  n855 ) | ( Pcount_0_  &  n855 ) ;
 assign n29 = ( (~ Poutreg_9_)  &  n869 ) | ( Pcount_0_  &  n869 ) ;
 assign n30 = ( (~ Poutreg_7_)  &  n884 ) | ( Pcount_0_  &  n884 ) ;
 assign n31 = ( (~ Poutreg_5_)  &  n891 ) | ( Pcount_0_  &  n891 ) ;
 assign n32 = ( (~ Poutreg_3_)  &  n907 ) | ( Pcount_0_  &  n907 ) ;
 assign n33 = ( (~ Poutreg_1_)  &  n920 ) | ( Pcount_0_  &  n920 ) ;
 assign n34 = ( (~ Pcount_3_)  &  n924 ) | ( n924  &  n926 ) | ( (~ Pcount_3_)  &  n928 ) | ( n926  &  n928 ) ;
 assign n35 = ( (~ Pinreg_55_)  &  (~ Pinreg_47_) ) | ( (~ Pinreg_47_)  &  Pcount_0_ ) | ( (~ Pinreg_55_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n36 = ( (~ Pinreg_54_)  &  (~ Pinreg_46_) ) | ( (~ Pinreg_46_)  &  Pcount_0_ ) | ( (~ Pinreg_54_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n37 = ( (~ Pinreg_53_)  &  (~ Pinreg_45_) ) | ( (~ Pinreg_45_)  &  Pcount_0_ ) | ( (~ Pinreg_53_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n38 = ( (~ Pinreg_52_)  &  (~ Pinreg_44_) ) | ( (~ Pinreg_44_)  &  Pcount_0_ ) | ( (~ Pinreg_52_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n39 = ( (~ Pinreg_51_)  &  (~ Pinreg_43_) ) | ( (~ Pinreg_43_)  &  Pcount_0_ ) | ( (~ Pinreg_51_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n40 = ( (~ Pinreg_50_)  &  (~ Pinreg_42_) ) | ( (~ Pinreg_42_)  &  Pcount_0_ ) | ( (~ Pinreg_50_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n41 = ( (~ Pinreg_49_)  &  (~ Pinreg_41_) ) | ( (~ Pinreg_41_)  &  Pcount_0_ ) | ( (~ Pinreg_49_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n42 = ( (~ Pinreg_48_)  &  (~ Pinreg_40_) ) | ( (~ Pinreg_40_)  &  Pcount_0_ ) | ( (~ Pinreg_48_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n43 = ( (~ Pinreg_47_)  &  (~ Pinreg_39_) ) | ( (~ Pinreg_39_)  &  Pcount_0_ ) | ( (~ Pinreg_47_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n44 = ( (~ Pinreg_46_)  &  (~ Pinreg_38_) ) | ( (~ Pinreg_38_)  &  Pcount_0_ ) | ( (~ Pinreg_46_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n45 = ( (~ Pinreg_45_)  &  (~ Pinreg_37_) ) | ( (~ Pinreg_37_)  &  Pcount_0_ ) | ( (~ Pinreg_45_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n46 = ( (~ Pinreg_44_)  &  (~ Pinreg_36_) ) | ( (~ Pinreg_36_)  &  Pcount_0_ ) | ( (~ Pinreg_44_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n47 = ( (~ Pinreg_43_)  &  (~ Pinreg_35_) ) | ( (~ Pinreg_35_)  &  Pcount_0_ ) | ( (~ Pinreg_43_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n48 = ( (~ Pinreg_42_)  &  (~ Pinreg_34_) ) | ( (~ Pinreg_34_)  &  Pcount_0_ ) | ( (~ Pinreg_42_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n49 = ( (~ Pinreg_41_)  &  (~ Pinreg_33_) ) | ( (~ Pinreg_33_)  &  Pcount_0_ ) | ( (~ Pinreg_41_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n50 = ( (~ Pinreg_40_)  &  (~ Pinreg_32_) ) | ( (~ Pinreg_32_)  &  Pcount_0_ ) | ( (~ Pinreg_40_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n51 = ( (~ Pinreg_39_)  &  (~ Pinreg_31_) ) | ( (~ Pinreg_31_)  &  Pcount_0_ ) | ( (~ Pinreg_39_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n52 = ( (~ Pinreg_38_)  &  (~ Pinreg_30_) ) | ( (~ Pinreg_30_)  &  Pcount_0_ ) | ( (~ Pinreg_38_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n53 = ( (~ Pinreg_37_)  &  (~ Pinreg_29_) ) | ( (~ Pinreg_29_)  &  Pcount_0_ ) | ( (~ Pinreg_37_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n54 = ( (~ Pinreg_36_)  &  (~ Pinreg_28_) ) | ( (~ Pinreg_28_)  &  Pcount_0_ ) | ( (~ Pinreg_36_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n55 = ( (~ Pinreg_35_)  &  (~ Pinreg_27_) ) | ( (~ Pinreg_27_)  &  Pcount_0_ ) | ( (~ Pinreg_35_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n56 = ( (~ Pinreg_34_)  &  (~ Pinreg_26_) ) | ( (~ Pinreg_26_)  &  Pcount_0_ ) | ( (~ Pinreg_34_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n57 = ( (~ Pinreg_33_)  &  (~ Pinreg_25_) ) | ( (~ Pinreg_25_)  &  Pcount_0_ ) | ( (~ Pinreg_33_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n58 = ( (~ Pinreg_32_)  &  (~ Pinreg_24_) ) | ( (~ Pinreg_24_)  &  Pcount_0_ ) | ( (~ Pinreg_32_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n59 = ( (~ Pinreg_31_)  &  (~ Pinreg_23_) ) | ( (~ Pinreg_23_)  &  Pcount_0_ ) | ( (~ Pinreg_31_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n60 = ( (~ Pinreg_30_)  &  (~ Pinreg_22_) ) | ( (~ Pinreg_22_)  &  Pcount_0_ ) | ( (~ Pinreg_30_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n61 = ( (~ Pinreg_29_)  &  (~ Pinreg_21_) ) | ( (~ Pinreg_21_)  &  Pcount_0_ ) | ( (~ Pinreg_29_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n62 = ( (~ Pinreg_28_)  &  (~ Pinreg_20_) ) | ( (~ Pinreg_20_)  &  Pcount_0_ ) | ( (~ Pinreg_28_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n63 = ( (~ Pinreg_27_)  &  (~ Pinreg_19_) ) | ( (~ Pinreg_19_)  &  Pcount_0_ ) | ( (~ Pinreg_27_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n64 = ( (~ Pinreg_26_)  &  (~ Pinreg_18_) ) | ( (~ Pinreg_18_)  &  Pcount_0_ ) | ( (~ Pinreg_26_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n65 = ( (~ Pinreg_25_)  &  (~ Pinreg_17_) ) | ( (~ Pinreg_17_)  &  Pcount_0_ ) | ( (~ Pinreg_25_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n66 = ( (~ Pinreg_24_)  &  (~ Pinreg_16_) ) | ( (~ Pinreg_16_)  &  Pcount_0_ ) | ( (~ Pinreg_24_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n67 = ( (~ Pinreg_23_)  &  (~ Pinreg_15_) ) | ( (~ Pinreg_15_)  &  Pcount_0_ ) | ( (~ Pinreg_23_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n68 = ( (~ Pinreg_22_)  &  (~ Pinreg_14_) ) | ( (~ Pinreg_14_)  &  Pcount_0_ ) | ( (~ Pinreg_22_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n69 = ( (~ Pinreg_21_)  &  (~ Pinreg_13_) ) | ( (~ Pinreg_13_)  &  Pcount_0_ ) | ( (~ Pinreg_21_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n70 = ( (~ Pinreg_20_)  &  (~ Pinreg_12_) ) | ( (~ Pinreg_12_)  &  Pcount_0_ ) | ( (~ Pinreg_20_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n71 = ( (~ Pinreg_19_)  &  (~ Pinreg_11_) ) | ( (~ Pinreg_11_)  &  Pcount_0_ ) | ( (~ Pinreg_19_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n72 = ( (~ Pinreg_18_)  &  (~ Pinreg_10_) ) | ( (~ Pinreg_10_)  &  Pcount_0_ ) | ( (~ Pinreg_18_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n73 = ( (~ Pinreg_17_)  &  (~ Pinreg_9_) ) | ( (~ Pinreg_9_)  &  Pcount_0_ ) | ( (~ Pinreg_17_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n74 = ( (~ Pinreg_16_)  &  (~ Pinreg_8_) ) | ( (~ Pinreg_8_)  &  Pcount_0_ ) | ( (~ Pinreg_16_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n75 = ( (~ Pinreg_15_)  &  (~ Pinreg_7_) ) | ( (~ Pinreg_7_)  &  Pcount_0_ ) | ( (~ Pinreg_15_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n76 = ( (~ Pinreg_14_)  &  (~ Pinreg_6_) ) | ( (~ Pinreg_6_)  &  Pcount_0_ ) | ( (~ Pinreg_14_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n77 = ( (~ Pinreg_13_)  &  (~ Pinreg_5_) ) | ( (~ Pinreg_5_)  &  Pcount_0_ ) | ( (~ Pinreg_13_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n78 = ( (~ Pinreg_12_)  &  (~ Pinreg_4_) ) | ( (~ Pinreg_4_)  &  Pcount_0_ ) | ( (~ Pinreg_12_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n79 = ( (~ Pinreg_11_)  &  (~ Pinreg_3_) ) | ( (~ Pinreg_3_)  &  Pcount_0_ ) | ( (~ Pinreg_11_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n80 = ( (~ Pinreg_10_)  &  (~ Pinreg_2_) ) | ( (~ Pinreg_2_)  &  Pcount_0_ ) | ( (~ Pinreg_10_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n81 = ( (~ Pinreg_9_)  &  (~ Pinreg_1_) ) | ( (~ Pinreg_1_)  &  Pcount_0_ ) | ( (~ Pinreg_9_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n82 = ( (~ Pinreg_8_)  &  (~ Pinreg_0_) ) | ( (~ Pinreg_0_)  &  Pcount_0_ ) | ( (~ Pinreg_8_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n83 = ( (~ Pinreg_7_)  &  (~ Pdata_in_7_) ) | ( (~ Pdata_in_7_)  &  Pcount_0_ ) | ( (~ Pinreg_7_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n84 = ( (~ Pinreg_6_)  &  (~ Pdata_in_6_) ) | ( (~ Pdata_in_6_)  &  Pcount_0_ ) | ( (~ Pinreg_6_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n85 = ( (~ Pinreg_5_)  &  (~ Pdata_in_5_) ) | ( (~ Pdata_in_5_)  &  Pcount_0_ ) | ( (~ Pinreg_5_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n86 = ( (~ Pinreg_4_)  &  (~ Pdata_in_4_) ) | ( (~ Pdata_in_4_)  &  Pcount_0_ ) | ( (~ Pinreg_4_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n87 = ( (~ Pinreg_3_)  &  (~ Pdata_in_3_) ) | ( (~ Pdata_in_3_)  &  Pcount_0_ ) | ( (~ Pinreg_3_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n88 = ( (~ Pinreg_2_)  &  (~ Pdata_in_2_) ) | ( (~ Pdata_in_2_)  &  Pcount_0_ ) | ( (~ Pinreg_2_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n89 = ( (~ Pinreg_1_)  &  (~ Pdata_in_1_) ) | ( (~ Pdata_in_1_)  &  Pcount_0_ ) | ( (~ Pinreg_1_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n90 = ( (~ Pinreg_0_)  &  (~ Pdata_in_0_) ) | ( (~ Pdata_in_0_)  &  Pcount_0_ ) | ( (~ Pinreg_0_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n91 = ( (~ Poutreg_56_)  &  (~ Pdata_32_) ) | ( (~ Pdata_32_)  &  Pcount_0_ ) | ( (~ Poutreg_56_)  &  n1 ) | ( Pcount_0_  &  n1 ) ;
 assign n92 = ( Pload_key_0_  &  (~ n1) ) ;
 assign n94 = ( (~ Pdata_49_)  &  n414 ) | ( n1  &  n414 ) ;
 assign n95 = ( (~ Pdata_39_)  &  n922 ) | ( n1  &  n922 ) ;
 assign n96 = ( (~ Pdata_47_)  &  n909 ) | ( n1  &  n909 ) ;
 assign n97 = ( (~ Poutreg_58_)  &  (~ Pdata_40_) ) | ( (~ Pdata_40_)  &  Pcount_0_ ) | ( (~ Poutreg_58_)  &  n1 ) | ( Pcount_0_  &  n1 ) ;
 assign n98 = ( (~ Pdata_55_)  &  n893 ) | ( n1  &  n893 ) ;
 assign n99 = ( (~ Pdata_63_)  &  n886 ) | ( n1  &  n886 ) ;
 assign n100 = ( (~ Pdata_38_)  &  n871 ) | ( n1  &  n871 ) ;
 assign n101 = ( (~ Poutreg_60_)  &  (~ Pdata_48_) ) | ( (~ Pdata_48_)  &  Pcount_0_ ) | ( (~ Poutreg_60_)  &  n1 ) | ( Pcount_0_  &  n1 ) ;
 assign n102 = ( (~ Pdata_46_)  &  n857 ) | ( n1  &  n857 ) ;
 assign n103 = ( (~ Pdata_54_)  &  n845 ) | ( n1  &  n845 ) ;
 assign n104 = ( (~ Pdata_62_)  &  n833 ) | ( n1  &  n833 ) ;
 assign n105 = ( (~ Poutreg_62_)  &  (~ Pdata_56_) ) | ( (~ Pdata_56_)  &  Pcount_0_ ) | ( (~ Poutreg_62_)  &  n1 ) | ( Pcount_0_  &  n1 ) ;
 assign n106 = ( (~ Pdata_37_)  &  n821 ) | ( n1  &  n821 ) ;
 assign n107 = ( (~ Pdata_45_)  &  n799 ) | ( n1  &  n799 ) ;
 assign n108 = ( (~ Pdata_53_)  &  n785 ) | ( n1  &  n785 ) ;
 assign n109 = ( (~ Pdata_61_)  &  n764 ) | ( n1  &  n764 ) ;
 assign n110 = ( (~ Pdata_36_)  &  n708 ) | ( n1  &  n708 ) ;
 assign n111 = ( (~ Pdata_44_)  &  n700 ) | ( n1  &  n700 ) ;
 assign n112 = ( (~ Pdata_52_)  &  n689 ) | ( n1  &  n689 ) ;
 assign n113 = ( (~ Pdata_60_)  &  n667 ) | ( n1  &  n667 ) ;
 assign n114 = ( (~ Pdata_35_)  &  n652 ) | ( n1  &  n652 ) ;
 assign n115 = ( (~ Pdata_43_)  &  n641 ) | ( n1  &  n641 ) ;
 assign n116 = ( (~ Pdata_51_)  &  n598 ) | ( n1  &  n598 ) ;
 assign n117 = ( (~ Pdata_59_)  &  n582 ) | ( n1  &  n582 ) ;
 assign n118 = ( (~ Pdata_34_)  &  n566 ) | ( n1  &  n566 ) ;
 assign n119 = ( (~ Pdata_42_)  &  n553 ) | ( n1  &  n553 ) ;
 assign n120 = ( (~ Pdata_50_)  &  n540 ) | ( n1  &  n540 ) ;
 assign n121 = ( (~ Pdata_58_)  &  n507 ) | ( n1  &  n507 ) ;
 assign n122 = ( (~ Pdata_33_)  &  n457 ) | ( n1  &  n457 ) ;
 assign n123 = ( (~ Pdata_41_)  &  n430 ) | ( n1  &  n430 ) ;
 assign n124 = ( (~ Pdata_57_)  &  n367 ) | ( n1  &  n367 ) ;
 assign n126 = ( (~ Pcount_0_) ) | ( (~ n1) ) ;
 assign n191 = ( (~ n228)  &  (~ n227) ) | ( (~ n227)  &  (~ n230) ) | ( (~ n228)  &  (~ n559) ) | ( (~ n230)  &  (~ n559) ) ;
 assign n196 = ( (~ n207)  &  (~ n559) ) | ( (~ n228)  &  (~ n559) ) | ( (~ n207)  &  (~ n1184) ) | ( (~ n228)  &  (~ n1184) ) ;
 assign n201 = ( (~ Pdata_49_)  &  PD_2_ ) | ( Pdata_49_  &  (~ PD_2_) ) ;
 assign n199 = ( n191  &  n196 ) | ( n196  &  n201 ) | ( n191  &  (~ n912) ) | ( n201  &  (~ n912) ) ;
 assign n204 = ( (~ n1186)  &  n1457 ) | ( (~ n208)  &  n216  &  n1457 ) ;
 assign n202 = ( n199  &  n204  &  (~ n912) ) | ( n199  &  n204  &  (~ n1187) ) ;
 assign n209 = ( n915  &  (~ n1155) ) ;
 assign n208 = ( n912  &  n1185 ) ;
 assign n207 = ( (~ n220)  &  n1156 ) ;
 assign n205 = ( n209  &  n208 ) | ( n209  &  n207  &  (~ n224) ) ;
 assign n214 = ( n224 ) | ( (~ n1184) ) | ( (~ n1186) ) ;
 assign n212 = ( n1155 ) | ( n1188 ) ;
 assign n210 = ( (~ n205)  &  n214  &  n212 ) | ( (~ n205)  &  n214  &  (~ n911) ) ;
 assign n217 = ( n201 ) | ( n914 ) | ( (~ n1187) ) ;
 assign n218 = ( (~ n207)  &  n795 ) | ( (~ n207)  &  (~ n1185) ) | ( n795  &  n1189 ) | ( (~ n1185)  &  n1189 ) ;
 assign n216 = ( (~ n201) ) | ( (~ n230) ) ;
 assign n215 = ( n217  &  n218  &  n216 ) | ( n217  &  n218  &  (~ n559) ) ;
 assign n220 = ( (~ Pdata_50_)  &  PD_8_ ) | ( Pdata_50_  &  (~ PD_8_) ) ;
 assign n222 = ( (~ n914)  &  n1156 ) | ( n914  &  (~ n1156) ) ;
 assign n219 = ( n220 ) | ( n222 ) | ( (~ n1186) ) ;
 assign n224 = ( (~ n201) ) | ( n914 ) ;
 assign n223 = ( n224 ) | ( (~ n1186) ) ;
 assign n228 = ( n915  &  n1155 ) ;
 assign n227 = ( (~ n914)  &  n1185 ) ;
 assign n226 = ( n1185 ) | ( n1184 ) ;
 assign n225 = ( n228  &  n227 ) | ( n228  &  n201  &  n226 ) ;
 assign n230 = ( n911  &  (~ n914) ) ;
 assign n231 = ( n559 ) | ( n209 ) ;
 assign n229 = ( (~ n201)  &  (~ n219) ) | ( (~ n201)  &  n230  &  n231 ) ;
 assign n234 = ( (~ Pdata_24_)  &  n1669 ) | ( Pdata_24_  &  (~ n1669) ) ;
 assign n243 = ( n266  &  (~ n275) ) ;
 assign n240 = ( (~ n262)  &  (~ n269)  &  (~ n835) ) ;
 assign n239 = ( n243  &  n240  &  (~ n1602) ) | ( n243  &  (~ n254)  &  (~ n1602) ) ;
 assign n244 = ( (~ n239)  &  (~ n262) ) | ( (~ n239)  &  (~ n272) ) | ( (~ n239)  &  (~ n1372) ) ;
 assign n252 = ( (~ n294)  &  (~ n835) ) | ( n297  &  (~ n835) ) | ( (~ n294)  &  (~ n1371) ) | ( n297  &  (~ n1371) ) ;
 assign n249 = ( n244  &  n252  &  (~ n281) ) | ( n244  &  n252  &  (~ n1199) ) ;
 assign n254 = ( (~ Pdata_36_)  &  PC_4_ ) | ( Pdata_36_  &  (~ PC_4_) ) ;
 assign n253 = ( n254  &  (~ n281) ) | ( n254  &  (~ n835) ) | ( (~ n281)  &  (~ n1200) ) | ( (~ n835)  &  (~ n1200) ) ;
 assign n259 = ( (~ n266) ) | ( (~ n292) ) | ( n1198 ) ;
 assign n260 = ( (~ n294) ) | ( (~ n1199) ) ;
 assign n257 = ( n253  &  n259  &  n260 ) | ( n259  &  n260  &  (~ n295) ) ;
 assign n263 = ( n254 ) | ( (~ n262) ) ;
 assign n262 = ( (~ Pdata_35_)  &  PC_0_ ) | ( Pdata_35_  &  (~ PC_0_) ) ;
 assign n261 = ( (~ n254)  &  n263 ) | ( n263  &  n262 ) ;
 assign n266 = ( (~ Pdata_63_)  &  PC_13_ ) | ( Pdata_63_  &  (~ PC_13_) ) ;
 assign n264 = ( (~ n243)  &  n266 ) | ( (~ n243)  &  (~ n275) ) ;
 assign n269 = ( (~ Pdata_32_)  &  PC_16_ ) | ( Pdata_32_  &  (~ PC_16_) ) ;
 assign n268 = ( (~ n254)  &  n269 ) ;
 assign n272 = ( (~ n269)  &  (~ n275) ) ;
 assign n270 = ( (~ n254)  &  (~ n262)  &  n272 ) | ( (~ n254)  &  (~ n266)  &  n272 ) ;
 assign n275 = ( (~ Pdata_34_)  &  PC_23_ ) | ( Pdata_34_  &  (~ PC_23_) ) ;
 assign n274 = ( (~ n262)  &  n269 ) ;
 assign n273 = ( (~ n266)  &  n268  &  n275 ) | ( (~ n266)  &  n275  &  n274 ) ;
 assign n276 = ( n261  &  (~ n275) ) | ( (~ n272)  &  (~ n275) ) | ( n261  &  (~ n274) ) | ( (~ n272)  &  (~ n274) ) ;
 assign n279 = ( n835  &  n294 ) ;
 assign n278 = ( (~ n262)  &  n272  &  n279 ) ;
 assign n281 = ( (~ n254)  &  (~ n266) ) ;
 assign n280 = ( n240  &  (~ n275)  &  n281 ) ;
 assign n283 = ( (~ n266) ) | ( n276 ) | ( (~ n835) ) ;
 assign n285 = ( (~ n281)  &  (~ n292) ) | ( (~ n281)  &  (~ n1201) ) | ( (~ n292)  &  n1202 ) | ( (~ n1201)  &  n1202 ) ;
 assign n282 = ( n249  &  n257  &  n283  &  n285  &  (~ n1203)  &  (~ n1599) ) ;
 assign n287 = ( (~ n282)  &  Pdata_16_ ) | ( n282  &  (~ Pdata_16_) ) ;
 assign n292 = ( n262  &  n254 ) ;
 assign n291 = ( n243  &  n269  &  n292 ) ;
 assign n294 = ( n254  &  (~ n266) ) ;
 assign n295 = ( n269  &  n262  &  n275 ) ;
 assign n293 = ( n291  &  (~ n835) ) | ( n294  &  n295  &  (~ n835) ) ;
 assign n299 = ( n263 ) | ( (~ n266) ) | ( n1198 ) ;
 assign n297 = ( n262 ) | ( n1198 ) ;
 assign n296 = ( (~ n281)  &  (~ n293)  &  n299 ) | ( (~ n293)  &  n299  &  n297 ) ;
 assign n300 = ( n254  &  n261 ) | ( n254  &  n269 ) | ( n261  &  (~ n274) ) | ( n269  &  (~ n274) ) ;
 assign n304 = ( (~ n243) ) | ( (~ n254) ) | ( n269 ) ;
 assign n305 = ( (~ n281) ) | ( n1198 ) ;
 assign n303 = ( n254  &  (~ n275) ) | ( n254  &  (~ n279) ) | ( n275  &  (~ n279) ) ;
 assign n301 = ( (~ n269)  &  n304  &  n305 ) | ( n304  &  n305  &  n303 ) ;
 assign n307 = ( (~ n275)  &  n1464 ) | ( n300  &  n1464 ) | ( (~ n1200)  &  n1464 ) ;
 assign n308 = ( n249  &  (~ n254)  &  n838 ) | ( n249  &  n838  &  n1202 ) ;
 assign n306 = ( (~ n262)  &  n307  &  n308 ) | ( n301  &  n307  &  n308 ) ;
 assign n309 = ( (~ n306)  &  Pdata_8_ ) | ( n306  &  (~ Pdata_8_) ) ;
 assign n314 = ( n357 ) | ( n1158 ) ;
 assign n315 = ( (~ n323) ) | ( n420 ) ;
 assign n317 = ( n325 ) | ( (~ n357) ) ;
 assign n313 = ( n314  &  n317 ) | ( n315  &  n317 ) | ( n314  &  (~ n591) ) | ( n315  &  (~ n591) ) ;
 assign n321 = ( n313  &  n359 ) | ( n326  &  n359 ) | ( n313  &  n1215 ) | ( n326  &  n1215 ) ;
 assign n319 = ( n314 ) | ( n355 ) ;
 assign n318 = ( n321  &  n319 ) | ( n321  &  (~ n588) ) ;
 assign n323 = ( (~ Pdata_43_)  &  PC_15_ ) | ( Pdata_43_  &  (~ PC_15_) ) ;
 assign n325 = ( n323 ) | ( (~ n585) ) ;
 assign n326 = ( (~ Pdata_48_)  &  PC_1_ ) | ( Pdata_48_  &  (~ PC_1_) ) ;
 assign n322 = ( n323  &  n325 ) | ( n323  &  n326 ) | ( n325  &  (~ n328) ) | ( n326  &  (~ n328) ) ;
 assign n329 = ( n323  &  (~ n326)  &  n585 ) ;
 assign n328 = ( n326  &  (~ n585) ) ;
 assign n327 = ( n329  &  (~ n1216) ) | ( n323  &  n328  &  (~ n1216) ) ;
 assign n331 = ( n319  &  n318  &  (~ n327) ) | ( n318  &  n322  &  (~ n327) ) ;
 assign n334 = ( (~ n329)  &  (~ n328) ) | ( (~ n328)  &  n1215 ) | ( (~ n329)  &  n1219 ) | ( n1215  &  n1219 ) ;
 assign n335 = ( n326  &  n1466 ) | ( (~ n1158)  &  n1466 ) | ( n1218  &  n1466 ) ;
 assign n333 = ( n334  &  n335 ) ;
 assign n339 = ( n314  &  n1465 ) | ( (~ n355)  &  n1465 ) | ( n359  &  n1465 ) ;
 assign n337 = ( n585 ) | ( n326 ) ;
 assign n336 = ( n339  &  n337 ) | ( n339  &  (~ n1376) ) ;
 assign n341 = ( (~ n323)  &  n1158 ) | ( n323  &  (~ n1158) ) ;
 assign n342 = ( n420 ) | ( n326 ) ;
 assign n343 = ( n355 ) | ( (~ n1158) ) ;
 assign n340 = ( n341  &  n343 ) | ( n342  &  n343 ) | ( n341  &  (~ n588) ) | ( n342  &  (~ n588) ) ;
 assign n345 = ( (~ n323) ) | ( n337 ) ;
 assign n344 = ( n345  &  n315  &  n325 ) | ( n345  &  n315  &  n326 ) ;
 assign n346 = ( (~ Pdata_0_)  &  n1672 ) | ( Pdata_0_  &  (~ n1672) ) ;
 assign n351 = ( (~ n326)  &  n337 ) | ( (~ n326)  &  n1219 ) | ( n337  &  n1221 ) | ( n1219  &  n1221 ) ;
 assign n352 = ( (~ n329)  &  n1471 ) | ( (~ n355)  &  n1471 ) | ( n1217  &  n1471 ) ;
 assign n350 = ( n351  &  n352 ) ;
 assign n357 = ( (~ Pdata_46_)  &  PC_19_ ) | ( Pdata_46_  &  (~ PC_19_) ) ;
 assign n355 = ( (~ Pdata_44_)  &  PC_6_ ) | ( Pdata_44_  &  (~ PC_6_) ) ;
 assign n353 = ( (~ n340)  &  n357 ) | ( n357  &  n355  &  (~ n359) ) ;
 assign n359 = ( n325 ) | ( (~ n326) ) ;
 assign n358 = ( n319 ) | ( n359 ) ;
 assign n360 = ( n323  &  (~ n1469) ) | ( n323  &  (~ n585)  &  (~ n1215) ) ;
 assign n365 = ( (~ Poutreg_63_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_63_)  &  n1472 ) | ( n126  &  n1472 ) ;
 assign n367 = ( (~ Poutreg_62_)  &  (~ Poutreg_54_) ) | ( (~ Poutreg_62_)  &  Pcount_0_ ) | ( (~ Poutreg_54_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n371 = ( (~ n382)  &  n403 ) | ( (~ n380)  &  n403 ) | ( (~ n382)  &  n692 ) | ( (~ n380)  &  n692 ) ;
 assign n369 = ( (~ n403) ) | ( n572 ) ;
 assign n368 = ( n371  &  n369 ) | ( n371  &  (~ n432) ) ;
 assign n373 = ( (~ n375) ) | ( (~ n570) ) ;
 assign n372 = ( n369 ) | ( n373 ) | ( (~ n432) ) ;
 assign n375 = ( (~ Pdata_36_)  &  PC_27_ ) | ( Pdata_36_  &  (~ PC_27_) ) ;
 assign n377 = ( n389 ) | ( (~ n570) ) ;
 assign n374 = ( n375 ) | ( n377 ) | ( (~ n380) ) ;
 assign n382 = ( (~ n450)  &  (~ n1159) ) ;
 assign n380 = ( n403  &  n572 ) ;
 assign n378 = ( n382  &  (~ n408) ) | ( n382  &  n380  &  (~ n1232) ) ;
 assign n386 = ( n372  &  n374  &  (~ n378) ) ;
 assign n387 = ( (~ n444)  &  n1474 ) | ( (~ n570)  &  n1474 ) | ( n1234  &  n1474 ) ;
 assign n384 = ( n1232 ) | ( n403 ) ;
 assign n385 = ( n389 ) | ( (~ n572) ) ;
 assign n383 = ( n386  &  n387  &  n384 ) | ( n386  &  n387  &  n385 ) ;
 assign n389 = ( (~ n450) ) | ( n1159 ) ;
 assign n392 = ( n375 ) | ( (~ n570) ) ;
 assign n388 = ( n389  &  n392 ) | ( n392  &  (~ n447) ) | ( n389  &  (~ n444) ) | ( (~ n447)  &  (~ n444) ) ;
 assign n395 = ( (~ n375) ) | ( n404 ) | ( n452 ) ;
 assign n396 = ( n384 ) | ( n692 ) ;
 assign n393 = ( n388  &  n395  &  n396 ) | ( n395  &  n396  &  (~ n445) ) ;
 assign n398 = ( n389  &  n434 ) | ( n389  &  (~ n447) ) | ( n434  &  n449 ) | ( (~ n447)  &  n449 ) ;
 assign n399 = ( (~ n375)  &  n1473 ) | ( n401  &  n1473 ) | ( n452  &  n1473 ) ;
 assign n397 = ( n398  &  n399 ) ;
 assign n401 = ( (~ n382) ) | ( (~ n572) ) ;
 assign n400 = ( n397  &  n393  &  n384 ) | ( n397  &  n393  &  n401 ) ;
 assign n405 = ( n369 ) | ( (~ n570) ) | ( n1159 ) ;
 assign n406 = ( (~ n382)  &  (~ n380) ) | ( (~ n380)  &  (~ n445) ) | ( (~ n382)  &  (~ n450) ) | ( (~ n445)  &  (~ n450) ) ;
 assign n403 = ( (~ Pdata_37_)  &  PC_14_ ) | ( Pdata_37_  &  (~ PC_14_) ) ;
 assign n404 = ( (~ n444) ) | ( (~ n572) ) ;
 assign n402 = ( n405  &  n406  &  n403 ) | ( n405  &  n406  &  n404 ) ;
 assign n409 = ( n1476  &  n368 ) | ( n1476  &  n392 ) ;
 assign n410 = ( (~ n375)  &  n383  &  n400 ) | ( n383  &  n400  &  n402 ) ;
 assign n408 = ( n572 ) | ( n384 ) ;
 assign n407 = ( n409  &  n410  &  n389 ) | ( n409  &  n410  &  n408 ) ;
 assign n412 = ( (~ Poutreg_61_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_61_)  &  n1477 ) | ( n126  &  n1477 ) ;
 assign n414 = ( (~ Poutreg_60_)  &  (~ Poutreg_52_) ) | ( (~ Poutreg_60_)  &  Pcount_0_ ) | ( (~ Poutreg_52_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n416 = ( n341 ) | ( n357 ) | ( (~ n355) ) | ( (~ n585) ) ;
 assign n417 = ( n315  &  n325 ) | ( n1217  &  n325 ) | ( n315  &  n343 ) | ( n1217  &  n343 ) ;
 assign n415 = ( n416  &  n417  &  n317 ) | ( n416  &  n417  &  n355 ) ;
 assign n421 = ( n325 ) | ( n357 ) | ( (~ n591) ) ;
 assign n420 = ( (~ n355) ) | ( n585 ) ;
 assign n418 = ( n341  &  n421 ) | ( (~ n357)  &  n421 ) | ( n421  &  n420 ) ;
 assign n423 = ( (~ n326)  &  n415 ) | ( n326  &  n418 ) | ( n415  &  n418 ) ;
 assign n424 = ( n336  &  n333 ) ;
 assign n425 = ( n317  &  n319 ) | ( n317  &  (~ n323) ) | ( n319  &  n343 ) | ( (~ n323)  &  n343 ) ;
 assign n426 = ( (~ n588)  &  n594 ) | ( n594  &  n1217 ) ;
 assign n422 = ( n423  &  n350  &  n424  &  n318  &  n425  &  n426 ) ;
 assign n428 = ( (~ Poutreg_59_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_59_)  &  n1478 ) | ( n126  &  n1478 ) ;
 assign n430 = ( (~ Poutreg_58_)  &  (~ Poutreg_50_) ) | ( (~ Poutreg_58_)  &  Pcount_0_ ) | ( (~ Poutreg_50_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n432 = ( n450  &  n1159 ) ;
 assign n431 = ( (~ n408)  &  n432 ) | ( n380  &  n432  &  (~ n1232) ) ;
 assign n436 = ( n375 ) | ( n377 ) | ( (~ n445) ) ;
 assign n434 = ( (~ n403) ) | ( n404 ) ;
 assign n433 = ( n373  &  (~ n431)  &  n436 ) | ( (~ n431)  &  n436  &  n434 ) ;
 assign n438 = ( n389  &  (~ n444) ) ;
 assign n437 = ( n373 ) | ( n438 ) | ( n369 ) ;
 assign n441 = ( (~ n382)  &  n570  &  n692 ) ;
 assign n442 = ( n385  &  (~ n570) ) ;
 assign n439 = ( n375 ) | ( (~ n403) ) | ( n441 ) | ( n442 ) ;
 assign n447 = ( n375  &  (~ n570) ) ;
 assign n444 = ( (~ n450)  &  n1159 ) ;
 assign n445 = ( (~ n403)  &  (~ n572) ) ;
 assign n443 = ( (~ n368)  &  n447 ) | ( n447  &  n444  &  n445 ) ;
 assign n449 = ( n570 ) | ( n1234 ) ;
 assign n450 = ( (~ Pdata_39_)  &  PC_20_ ) | ( Pdata_39_  &  (~ PC_20_) ) ;
 assign n448 = ( n449 ) | ( n450 ) ;
 assign n452 = ( n403 ) | ( (~ n570) ) ;
 assign n453 = ( n404  &  (~ n1160) ) ;
 assign n451 = ( n452 ) | ( n453 ) ;
 assign n455 = ( (~ Poutreg_57_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_57_)  &  n1479 ) | ( n126  &  n1479 ) ;
 assign n457 = ( (~ Poutreg_56_)  &  (~ Poutreg_48_) ) | ( (~ Poutreg_56_)  &  Pcount_0_ ) | ( (~ Poutreg_48_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n459 = ( (~ Pdata_63_)  &  PD_0_ ) | ( Pdata_63_  &  (~ PD_0_) ) ;
 assign n460 = ( (~ Pdata_61_)  &  PD_21_ ) | ( Pdata_61_  &  (~ PD_21_) ) ;
 assign n461 = ( (~ n491) ) | ( (~ n1246) ) ;
 assign n458 = ( n459 ) | ( n460 ) | ( n461 ) ;
 assign n464 = ( n475 ) | ( n1248 ) | ( n477 ) ;
 assign n463 = ( n459 ) | ( (~ n460) ) | ( n477 ) ;
 assign n462 = ( n461  &  n464  &  (~ n1607) ) | ( n464  &  n463  &  (~ n1607) ) ;
 assign n467 = ( n477  &  n1609 ) | ( n483  &  n1609 ) | ( (~ n852)  &  n1609 ) ;
 assign n468 = ( n472  &  (~ n849) ) | ( n472  &  n1251 ) | ( (~ n849)  &  n1480 ) | ( n1251  &  n1480 ) ;
 assign n466 = ( n467  &  n462  &  n468 ) ;
 assign n470 = ( (~ n460) ) | ( n491 ) | ( n675 ) ;
 assign n471 = ( n459 ) | ( (~ n477) ) ;
 assign n472 = ( n460 ) | ( n483 ) ;
 assign n473 = ( n477 ) | ( (~ n675) ) ;
 assign n469 = ( n470  &  n472 ) | ( n471  &  n472 ) | ( n470  &  n473 ) | ( n471  &  n473 ) ;
 assign n475 = ( (~ Pdata_59_)  &  PD_17_ ) | ( Pdata_59_  &  (~ PD_17_) ) ;
 assign n476 = ( (~ n477) ) | ( (~ n675) ) ;
 assign n477 = ( (~ Pdata_32_)  &  PD_3_ ) | ( Pdata_32_  &  (~ PD_3_) ) ;
 assign n474 = ( n475  &  n477 ) | ( n476  &  n477 ) | ( n475  &  (~ n851) ) | ( n476  &  (~ n851) ) ;
 assign n480 = ( (~ n459) ) | ( n473 ) | ( (~ n475) ) | ( (~ n849) ) ;
 assign n481 = ( n1249 ) | ( n670 ) ;
 assign n479 = ( n480  &  n481  &  n474 ) | ( n480  &  n481  &  n472 ) ;
 assign n483 = ( n459 ) | ( n491 ) ;
 assign n482 = ( n475 ) | ( n483 ) | ( n476 ) ;
 assign n484 = ( (~ n475) ) | ( n476 ) | ( (~ n1250) ) ;
 assign n487 = ( n472 ) | ( n477 ) | ( (~ n1246) ) ;
 assign n491 = ( (~ Pdata_60_)  &  PD_13_ ) | ( Pdata_60_  &  (~ PD_13_) ) ;
 assign n489 = ( n460  &  (~ n482) ) | ( n460  &  n491  &  (~ n1251) ) ;
 assign n495 = ( n459 ) | ( n475 ) | ( (~ n849) ) ;
 assign n493 = ( (~ n459)  &  n495 ) | ( n461  &  n495 ) ;
 assign n497 = ( n459 ) | ( (~ n491) ) | ( (~ n852) ) ;
 assign n498 = ( n463 ) | ( (~ n851) ) ;
 assign n499 = ( (~ n459) ) | ( n460 ) | ( n461 ) ;
 assign n500 = ( (~ n477)  &  n1482 ) | ( n493  &  n1482  &  (~ n1633) ) ;
 assign n501 = ( (~ n460)  &  n1251 ) | ( n460  &  n1258 ) | ( n1251  &  n1258 ) ;
 assign n502 = ( n463  &  n469 ) | ( n463  &  (~ n475) ) | ( n469  &  (~ n491) ) | ( (~ n475)  &  (~ n491) ) ;
 assign n503 = ( n1254  &  n479 ) ;
 assign n496 = ( n497  &  n498  &  n499  &  n500  &  n501  &  n466  &  n502  &  n503 ) ;
 assign n505 = ( (~ Poutreg_55_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_55_)  &  n1483 ) | ( n126  &  n1483 ) ;
 assign n507 = ( (~ Poutreg_54_)  &  (~ Poutreg_46_) ) | ( (~ Poutreg_54_)  &  Pcount_0_ ) | ( (~ Poutreg_46_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n511 = ( (~ n510) ) | ( n531 ) ;
 assign n510 = ( (~ Pdata_55_)  &  PD_4_ ) | ( Pdata_55_  &  (~ PD_4_) ) ;
 assign n508 = ( n511  &  n510 ) | ( n511  &  (~ n531) ) ;
 assign n515 = ( (~ n1163)  &  (~ n1164) ) ;
 assign n513 = ( (~ n510)  &  n1270 ) ;
 assign n512 = ( n515  &  n513 ) | ( n515  &  (~ n1484) ) ;
 assign n519 = ( (~ n513)  &  (~ n1611) ) | ( (~ n549)  &  (~ n1611) ) | ( (~ n647)  &  (~ n1611) ) ;
 assign n520 = ( n1487  &  n1488  &  n543 ) | ( n1487  &  n1488  &  n526 ) ;
 assign n517 = ( n647 ) | ( n654 ) ;
 assign n516 = ( n519  &  n520  &  n517 ) | ( n519  &  n520  &  (~ n1272) ) ;
 assign n523 = ( n543  &  n1486 ) | ( (~ n513)  &  n1486  &  n1484 ) ;
 assign n522 = ( n510 ) | ( n532 ) ;
 assign n521 = ( n523  &  n522 ) | ( n523  &  n517 ) ;
 assign n527 = ( (~ n647) ) | ( n654 ) | ( (~ n1272) ) ;
 assign n528 = ( n543  &  n517 ) | ( n1273  &  n517 ) | ( n543  &  n1274 ) | ( n1273  &  n1274 ) ;
 assign n525 = ( n647 ) | ( n658 ) ;
 assign n526 = ( n546 ) | ( n511 ) ;
 assign n524 = ( n527  &  n528  &  n525 ) | ( n527  &  n528  &  n526 ) ;
 assign n532 = ( (~ n531) ) | ( n546 ) ;
 assign n531 = ( (~ Pdata_51_)  &  PD_1_ ) | ( Pdata_51_  &  (~ PD_1_) ) ;
 assign n529 = ( n532  &  n531 ) | ( n532  &  (~ n546) ) ;
 assign n534 = ( n524  &  n521 ) ;
 assign n535 = ( (~ n647)  &  n1610 ) | ( n1489  &  n1490  &  n1610 ) ;
 assign n536 = ( n1492  &  n658 ) | ( n1492  &  n1274 ) ;
 assign n533 = ( n516  &  n534  &  n535  &  n536 ) ;
 assign n538 = ( (~ Poutreg_53_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_53_)  &  n1494 ) | ( n126  &  n1494 ) ;
 assign n540 = ( (~ Poutreg_52_)  &  (~ Poutreg_44_) ) | ( (~ Poutreg_52_)  &  Pcount_0_ ) | ( (~ Poutreg_44_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n544 = ( n1495  &  n517 ) | ( n1495  &  n1484  &  n1273 ) ;
 assign n542 = ( n546 ) | ( (~ n1265) ) ;
 assign n543 = ( (~ n647) ) | ( n658 ) ;
 assign n541 = ( n544  &  n542 ) | ( n544  &  n543 ) ;
 assign n549 = ( (~ n1163)  &  n1164 ) ;
 assign n546 = ( (~ Pdata_54_)  &  PD_16_ ) | ( Pdata_54_  &  (~ PD_16_) ) ;
 assign n545 = ( n549  &  (~ n1273) ) | ( (~ n508)  &  n549  &  n546 ) ;
 assign n551 = ( (~ Poutreg_51_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_51_)  &  n1500 ) | ( n126  &  n1500 ) ;
 assign n553 = ( (~ Poutreg_50_)  &  (~ Poutreg_42_) ) | ( (~ Poutreg_50_)  &  Pcount_0_ ) | ( (~ Poutreg_42_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n556 = ( n224 ) | ( (~ n559) ) | ( (~ n1184) ) ;
 assign n557 = ( (~ n207)  &  (~ n1185) ) | ( n212  &  (~ n1185) ) | ( (~ n207)  &  n1189 ) | ( n212  &  n1189 ) ;
 assign n554 = ( (~ n209)  &  n556  &  n557 ) | ( n216  &  n556  &  n557 ) ;
 assign n559 = ( (~ n915)  &  n1155 ) ;
 assign n558 = ( n559  &  n224  &  n207 ) ;
 assign n561 = ( n1184  &  n228 ) ;
 assign n560 = ( n561  &  (~ n914) ) ;
 assign n564 = ( (~ Poutreg_49_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_49_)  &  (~ n1717) ) | ( n126  &  (~ n1717) ) ;
 assign n566 = ( (~ Poutreg_48_)  &  (~ Poutreg_40_) ) | ( (~ Poutreg_48_)  &  Pcount_0_ ) | ( (~ Poutreg_40_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n570 = ( (~ Pdata_35_)  &  PC_2_ ) | ( Pdata_35_  &  (~ PC_2_) ) ;
 assign n569 = ( (~ n403) ) | ( (~ n432) ) ;
 assign n567 = ( n377  &  n570 ) | ( n377  &  (~ n382)  &  n569 ) ;
 assign n572 = ( (~ Pdata_40_)  &  PC_9_ ) | ( Pdata_40_  &  (~ PC_9_) ) ;
 assign n571 = ( n572  &  n369 ) | ( n452  &  n369 ) | ( n572  &  n570 ) | ( n452  &  n570 ) ;
 assign n574 = ( n450  &  n567 ) | ( n450  &  (~ n572) ) | ( n567  &  n571 ) | ( (~ n572)  &  n571 ) ;
 assign n573 = ( (~ n432)  &  n574 ) | ( n452  &  n574 ) ;
 assign n576 = ( n384 ) | ( n404 ) ;
 assign n577 = ( (~ n375)  &  n570 ) | ( n570  &  n573 ) | ( (~ n375)  &  n1281 ) | ( n573  &  n1281 ) ;
 assign n578 = ( n1502  &  n377 ) | ( n1502  &  n1234 ) ;
 assign n575 = ( n433  &  n383  &  n393  &  n576  &  n577  &  n578 ) ;
 assign n580 = ( (~ Poutreg_47_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_47_)  &  n1503 ) | ( n126  &  n1503 ) ;
 assign n582 = ( (~ Poutreg_46_)  &  (~ Poutreg_38_) ) | ( (~ Poutreg_46_)  &  Pcount_0_ ) | ( (~ Poutreg_38_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n585 = ( (~ Pdata_47_)  &  PC_12_ ) | ( Pdata_47_  &  (~ PC_12_) ) ;
 assign n583 = ( (~ n315)  &  n357 ) | ( n357  &  (~ n355)  &  n585 ) ;
 assign n588 = ( n323  &  n326  &  n585 ) ;
 assign n587 = ( (~ n317)  &  n355 ) | ( (~ n357)  &  n355  &  n588 ) ;
 assign n591 = ( n355  &  n1158 ) ;
 assign n590 = ( (~ n319)  &  n329 ) | ( n329  &  n357  &  n591 ) ;
 assign n594 = ( (~ n328) ) | ( n1215 ) ;
 assign n593 = ( n594 ) | ( n323 ) ;
 assign n596 = ( (~ Poutreg_45_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_45_)  &  n1504 ) | ( n126  &  n1504 ) ;
 assign n598 = ( (~ Poutreg_44_)  &  (~ Poutreg_36_) ) | ( (~ Poutreg_44_)  &  Pcount_0_ ) | ( (~ Poutreg_36_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n602 = ( n609  &  (~ n766) ) | ( (~ n766)  &  (~ n862) ) | ( n609  &  (~ n1380) ) | ( (~ n862)  &  (~ n1380) ) ;
 assign n600 = ( n873 ) | ( (~ n1167) ) ;
 assign n599 = ( n602  &  n600 ) | ( n602  &  (~ n781) ) ;
 assign n607 = ( (~ n629)  &  n1166 ) ;
 assign n604 = ( (~ n775)  &  (~ n1167) ) ;
 assign n605 = ( (~ n766)  &  (~ n776) ) ;
 assign n603 = ( (~ n600)  &  n607 ) | ( n607  &  n604  &  n605 ) ;
 assign n612 = ( (~ n772) ) | ( (~ n781) ) | ( n1292 ) ;
 assign n609 = ( n1292 ) | ( (~ n1293) ) ;
 assign n608 = ( (~ n603)  &  n612  &  n609 ) | ( (~ n603)  &  n612  &  (~ n773) ) ;
 assign n615 = ( n766 ) | ( (~ n776) ) ;
 assign n613 = ( (~ n607)  &  n615 ) | ( (~ n605)  &  n615 ) | ( (~ n607)  &  (~ n862) ) | ( (~ n605)  &  (~ n862) ) ;
 assign n620 = ( (~ n766) ) | ( n1166 ) | ( (~ n1295) ) ;
 assign n621 = ( n609 ) | ( (~ n781) ) ;
 assign n618 = ( n613  &  n620  &  n621 ) | ( n620  &  n621  &  (~ n777) ) ;
 assign n622 = ( (~ n773)  &  (~ n772) ) | ( (~ n773)  &  (~ n862) ) | ( (~ n772)  &  (~ n1293) ) | ( (~ n862)  &  (~ n1293) ) ;
 assign n626 = ( (~ n607) ) | ( (~ n780) ) | ( (~ n1293) ) ;
 assign n627 = ( (~ n604) ) | ( n1297 ) ;
 assign n625 = ( n622  &  n626  &  n627 ) | ( n626  &  n627  &  (~ n777) ) ;
 assign n631 = ( (~ n780) ) | ( (~ n862) ) ;
 assign n632 = ( (~ n777) ) | ( (~ n776) ) | ( n1300 ) ;
 assign n629 = ( (~ Pdata_57_)  &  PD_10_ ) | ( Pdata_57_  &  (~ PD_10_) ) ;
 assign n628 = ( n631  &  n632  &  n629 ) | ( n631  &  n632  &  (~ n866) ) ;
 assign n634 = ( n1624  &  n1300 ) | ( n1624  &  n1301 ) ;
 assign n635 = ( n608  &  n599 ) ;
 assign n636 = ( n628  &  (~ n775) ) | ( (~ n766)  &  (~ n775) ) | ( n628  &  n1297 ) | ( (~ n766)  &  n1297 ) ;
 assign n637 = ( (~ n773)  &  n878 ) | ( (~ n773)  &  (~ n1166) ) | ( n878  &  n1298 ) | ( (~ n1166)  &  n1298 ) ;
 assign n633 = ( n634  &  n635  &  n618  &  n625  &  n636  &  n637 ) ;
 assign n639 = ( (~ Poutreg_43_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_43_)  &  n1505 ) | ( n126  &  n1505 ) ;
 assign n641 = ( (~ Poutreg_42_)  &  (~ Poutreg_34_) ) | ( (~ Poutreg_42_)  &  Pcount_0_ ) | ( (~ Poutreg_34_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n642 = ( n508  &  (~ n1265) ) | ( (~ n1165)  &  (~ n1265) ) | ( n508  &  (~ n1303) ) | ( (~ n1165)  &  (~ n1303) ) ;
 assign n648 = ( (~ n510) ) | ( (~ n531) ) ;
 assign n647 = ( (~ Pdata_53_)  &  PD_22_ ) | ( Pdata_53_  &  (~ PD_22_) ) ;
 assign n646 = ( n510  &  n648  &  (~ n1265) ) | ( n648  &  n647  &  (~ n1265) ) ;
 assign n650 = ( (~ Poutreg_41_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_41_)  &  n1507 ) | ( n126  &  n1507 ) ;
 assign n652 = ( (~ Poutreg_40_)  &  (~ Poutreg_32_) ) | ( (~ Poutreg_40_)  &  Pcount_0_ ) | ( (~ Poutreg_32_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n655 = ( n1164 ) | ( n1274 ) ;
 assign n656 = ( n658  &  n1508  &  n1509 ) | ( (~ n1272)  &  n1508  &  n1509 ) ;
 assign n654 = ( (~ n1163) ) | ( (~ n1164) ) ;
 assign n653 = ( n655  &  n656  &  n522 ) | ( n655  &  n656  &  n654 ) ;
 assign n659 = ( n510 ) | ( n529 ) | ( (~ n549) ) ;
 assign n660 = ( n1163  &  (~ n1265) ) | ( (~ n1265)  &  (~ n1272) ) | ( n1163  &  n1275 ) | ( (~ n1272)  &  n1275 ) ;
 assign n658 = ( (~ n1163) ) | ( n1164 ) ;
 assign n657 = ( n659  &  n660  &  n508 ) | ( n659  &  n660  &  n658 ) ;
 assign n662 = ( n647  &  n653 ) | ( (~ n647)  &  n657 ) | ( n653  &  n657 ) ;
 assign n663 = ( n524  &  n542 ) | ( n524  &  n517 ) ;
 assign n661 = ( n662  &  n541  &  n663  &  n516 ) ;
 assign n665 = ( (~ Poutreg_39_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_39_)  &  n1510 ) | ( n126  &  n1510 ) ;
 assign n667 = ( (~ Poutreg_38_)  &  (~ Poutreg_30_) ) | ( (~ Poutreg_38_)  &  Pcount_0_ ) | ( (~ Poutreg_30_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n671 = ( n463 ) | ( n475 ) | ( n491 ) | ( (~ n675) ) ;
 assign n672 = ( n477  &  n1628 ) | ( (~ n1246)  &  n1628 ) | ( (~ n1250)  &  n1628 ) ;
 assign n670 = ( (~ n477) ) | ( (~ n852) ) ;
 assign n668 = ( n671  &  n672  &  n670 ) | ( n671  &  n672  &  (~ n1252) ) ;
 assign n675 = ( (~ Pdata_62_)  &  PD_7_ ) | ( Pdata_62_  &  (~ PD_7_) ) ;
 assign n673 = ( n473  &  (~ n477) ) | ( n473  &  n675 ) ;
 assign n678 = ( n472 ) | ( (~ n851) ) ;
 assign n679 = ( n459 ) | ( (~ n491) ) | ( (~ n675) ) | ( n1168 ) ;
 assign n676 = ( (~ n460)  &  n678  &  n679 ) | ( n461  &  n678  &  n679 ) ;
 assign n681 = ( n673 ) | ( n1249 ) | ( n1168 ) ;
 assign n682 = ( n675 ) | ( (~ n1168) ) | ( (~ n1252) ) ;
 assign n683 = ( (~ n477)  &  n497 ) | ( n477  &  n676 ) | ( n497  &  n676 ) ;
 assign n684 = ( n459 ) | ( n1257 ) ;
 assign n685 = ( n473  &  (~ n491) ) | ( (~ n491)  &  n495 ) | ( n473  &  n498 ) | ( n495  &  n498 ) ;
 assign n680 = ( n681  &  n682  &  n683  &  n668  &  n503  &  n462  &  n684  &  n685 ) ;
 assign n687 = ( (~ Poutreg_37_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_37_)  &  n1511 ) | ( n126  &  n1511 ) ;
 assign n689 = ( (~ Poutreg_36_)  &  (~ Poutreg_28_) ) | ( (~ Poutreg_36_)  &  Pcount_0_ ) | ( (~ Poutreg_28_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n691 = ( n438 ) | ( (~ n570) ) | ( n572 ) ;
 assign n692 = ( (~ n432) ) | ( (~ n572) ) ;
 assign n690 = ( (~ n382)  &  n691  &  n692 ) | ( n570  &  n691  &  n692 ) ;
 assign n694 = ( (~ n403)  &  n1631 ) | ( n453  &  n1631 ) | ( n570  &  n1631 ) ;
 assign n695 = ( (~ n375) ) | ( n403 ) | ( n690 ) ;
 assign n696 = ( n408  &  (~ n1232) ) | ( (~ n444)  &  (~ n1232) ) | ( n408  &  n1281 ) | ( (~ n444)  &  n1281 ) ;
 assign n693 = ( n433  &  n383  &  n694  &  n397  &  n695  &  n696 ) ;
 assign n698 = ( (~ Poutreg_35_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_35_)  &  n1512 ) | ( n126  &  n1512 ) ;
 assign n700 = ( (~ Poutreg_34_)  &  (~ Poutreg_26_) ) | ( (~ Poutreg_34_)  &  Pcount_0_ ) | ( (~ Poutreg_26_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n702 = ( (~ n477)  &  n1514  &  (~ n1632) ) | ( n499  &  n1514  &  (~ n1632) ) ;
 assign n703 = ( n460  &  n675 ) | ( n1258  &  n675 ) | ( n460  &  n495 ) | ( n1258  &  n495 ) ;
 assign n704 = ( n679  &  n1257  &  n483 ) | ( n679  &  n1257  &  n670 ) ;
 assign n701 = ( n466  &  n479  &  n668  &  n702  &  n703  &  n704 ) ;
 assign n706 = ( (~ Poutreg_33_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_33_)  &  n1515 ) | ( n126  &  n1515 ) ;
 assign n708 = ( (~ Poutreg_32_)  &  (~ Poutreg_24_) ) | ( (~ Poutreg_32_)  &  Pcount_0_ ) | ( (~ Poutreg_24_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n710 = ( n742 ) | ( n895 ) ;
 assign n711 = ( (~ n751) ) | ( (~ n756) ) ;
 assign n709 = ( n710  &  (~ n719) ) | ( n711  &  (~ n719) ) | ( n710  &  (~ n720) ) | ( n711  &  (~ n720) ) ;
 assign n716 = ( n711 ) | ( (~ n742) ) | ( n1318 ) ;
 assign n717 = ( n729 ) | ( n898 ) | ( n742 ) ;
 assign n714 = ( n709  &  n716  &  n717 ) | ( n716  &  n717  &  (~ n801) ) ;
 assign n722 = ( n1169  &  n738 ) ;
 assign n721 = ( n719  &  (~ n742)  &  n895 ) ;
 assign n719 = ( (~ n751)  &  n756 ) ;
 assign n720 = ( n742  &  (~ n895) ) ;
 assign n718 = ( n722  &  n721 ) | ( n722  &  n719  &  n720 ) ;
 assign n727 = ( n711 ) | ( (~ n720) ) | ( n732 ) ;
 assign n724 = ( (~ n814) ) | ( (~ n895) ) ;
 assign n725 = ( n751 ) | ( n732 ) ;
 assign n723 = ( (~ n718)  &  n727  &  n724 ) | ( (~ n718)  &  n727  &  n725 ) ;
 assign n729 = ( (~ n738) ) | ( n1169 ) ;
 assign n730 = ( (~ n742) ) | ( (~ n895) ) ;
 assign n728 = ( (~ n719) ) | ( n729 ) | ( n730 ) ;
 assign n732 = ( n738 ) | ( (~ n1169) ) ;
 assign n731 = ( n732 ) | ( (~ n814) ) | ( (~ n888) ) ;
 assign n735 = ( n710 ) | ( n711 ) | ( (~ n722) ) ;
 assign n738 = ( (~ Pdata_44_)  &  PC_7_ ) | ( Pdata_44_  &  (~ PC_7_) ) ;
 assign n740 = ( (~ n802) ) | ( (~ n895) ) | ( n1169 ) ;
 assign n737 = ( n738 ) | ( n740 ) | ( (~ n751) ) ;
 assign n744 = ( n732 ) | ( (~ n742) ) | ( n898 ) ;
 assign n745 = ( n1635  &  n729 ) | ( n1635  &  n724 ) | ( n1635  &  n751 ) ;
 assign n742 = ( (~ Pdata_39_)  &  PC_22_ ) | ( Pdata_39_  &  (~ PC_22_) ) ;
 assign n743 = ( n725 ) | ( (~ n756) ) | ( (~ n895) ) ;
 assign n741 = ( n744  &  n745  &  n742 ) | ( n744  &  n745  &  n743 ) ;
 assign n748 = ( n711  &  (~ n719) ) | ( (~ n719)  &  n742 ) | ( n711  &  (~ n742) ) ;
 assign n746 = ( n748  &  (~ n751) ) | ( n748  &  (~ n802) ) ;
 assign n751 = ( (~ Pdata_41_)  &  PC_11_ ) | ( Pdata_41_  &  (~ PC_11_) ) ;
 assign n749 = ( n751  &  (~ n888) ) | ( (~ n888)  &  (~ n895) ) ;
 assign n754 = ( (~ n801) ) | ( n898 ) ;
 assign n752 = ( (~ n722)  &  n754 ) | ( n749  &  n754 ) | ( n754  &  (~ n756) ) ;
 assign n756 = ( (~ Pdata_40_)  &  PC_18_ ) | ( Pdata_40_  &  (~ PC_18_) ) ;
 assign n755 = ( (~ n719)  &  (~ n751) ) | ( n742  &  (~ n751) ) | ( (~ n719)  &  n756 ) | ( n742  &  n756 ) ;
 assign n759 = ( (~ n746)  &  n814 ) | ( (~ n746)  &  n1169 ) | ( n814  &  (~ n1169) ) ;
 assign n757 = ( (~ n738)  &  n759  &  (~ n895) ) ;
 assign n760 = ( n740 ) | ( n751 ) ;
 assign n762 = ( (~ Poutreg_31_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_31_)  &  n1517 ) | ( n126  &  n1517 ) ;
 assign n764 = ( (~ Poutreg_30_)  &  (~ Poutreg_22_) ) | ( (~ Poutreg_30_)  &  Pcount_0_ ) | ( (~ Poutreg_22_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n766 = ( (~ Pdata_59_)  &  PD_5_ ) | ( Pdata_59_  &  (~ PD_5_) ) ;
 assign n765 = ( n766 ) | ( (~ n1166) ) | ( (~ n1295) ) ;
 assign n769 = ( (~ n607) ) | ( (~ n604) ) | ( (~ n1293) ) ;
 assign n773 = ( (~ n629)  &  (~ n1166) ) ;
 assign n772 = ( n766  &  (~ n776) ) ;
 assign n771 = ( (~ n600)  &  n773 ) | ( n604  &  n773  &  n772 ) ;
 assign n777 = ( n775  &  (~ n1167) ) ;
 assign n775 = ( (~ Pdata_56_)  &  PD_20_ ) | ( Pdata_56_  &  (~ PD_20_) ) ;
 assign n776 = ( (~ Pdata_55_)  &  PD_15_ ) | ( Pdata_55_  &  (~ PD_15_) ) ;
 assign n774 = ( (~ n629)  &  n777 ) | ( (~ n629)  &  n775  &  n776 ) ;
 assign n780 = ( n775  &  n1167 ) ;
 assign n781 = ( n629  &  (~ n1166) ) ;
 assign n779 = ( n780  &  n781 ) ;
 assign n783 = ( (~ Poutreg_29_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_29_)  &  n1521 ) | ( n126  &  n1521 ) ;
 assign n785 = ( (~ Poutreg_28_)  &  (~ Poutreg_20_) ) | ( (~ Poutreg_28_)  &  Pcount_0_ ) | ( (~ Poutreg_20_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n786 = ( (~ n207)  &  (~ n789) ) | ( (~ n789)  &  (~ n914) ) ;
 assign n789 = ( n220  &  n222 ) ;
 assign n788 = ( n789  &  n209 ) ;
 assign n790 = ( (~ n915)  &  (~ n1383) ) | ( n230  &  (~ n915)  &  (~ n1155) ) ;
 assign n795 = ( (~ n1155) ) | ( n1188 ) ;
 assign n794 = ( n795 ) | ( (~ n1184) ) ;
 assign n797 = ( (~ Poutreg_27_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_27_)  &  n1524 ) | ( n126  &  n1524 ) ;
 assign n799 = ( (~ Poutreg_26_)  &  (~ Poutreg_18_) ) | ( (~ Poutreg_26_)  &  Pcount_0_ ) | ( (~ Poutreg_18_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n802 = ( n742  &  (~ n756) ) ;
 assign n803 = ( (~ n751)  &  (~ n895) ) ;
 assign n801 = ( (~ n738)  &  (~ n1169) ) ;
 assign n800 = ( n802  &  n803  &  n801 ) | ( n802  &  n803  &  n722 ) ;
 assign n806 = ( n751 ) | ( (~ n814) ) | ( n1318 ) ;
 assign n804 = ( (~ n721)  &  (~ n800)  &  n806 ) | ( (~ n801)  &  (~ n800)  &  n806 ) ;
 assign n808 = ( n711 ) | ( (~ n720) ) | ( (~ n801) ) ;
 assign n809 = ( n732 ) | ( n749 ) | ( (~ n802) ) ;
 assign n811 = ( n730  &  n710 ) ;
 assign n810 = ( (~ n719) ) | ( n811 ) | ( (~ n1340) ) ;
 assign n814 = ( (~ n742)  &  (~ n756) ) ;
 assign n813 = ( (~ n725)  &  n814  &  (~ n895) ) ;
 assign n817 = ( (~ n742)  &  (~ n898)  &  n1169 ) ;
 assign n816 = ( n817  &  n738 ) ;
 assign n819 = ( (~ Poutreg_25_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_25_)  &  (~ n1718) ) | ( n126  &  (~ n1718) ) ;
 assign n821 = ( (~ Poutreg_24_)  &  (~ Poutreg_16_) ) | ( (~ Poutreg_24_)  &  Pcount_0_ ) | ( (~ Poutreg_16_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n824 = ( (~ n266) ) | ( n1172 ) ;
 assign n822 = ( n254  &  (~ n279)  &  n824 ) | ( (~ n264)  &  (~ n279)  &  n824 ) ;
 assign n827 = ( (~ n254) ) | ( n297 ) ;
 assign n829 = ( (~ n274)  &  (~ n835) ) | ( n822  &  (~ n835) ) | ( (~ n274)  &  (~ n1201) ) | ( n822  &  (~ n1201) ) ;
 assign n826 = ( n249  &  n257  &  n296  &  n827  &  n829  &  (~ n1702) ) ;
 assign n831 = ( (~ Poutreg_23_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_23_)  &  n1528 ) | ( n126  &  n1528 ) ;
 assign n833 = ( (~ Poutreg_22_)  &  (~ Poutreg_14_) ) | ( (~ Poutreg_22_)  &  Pcount_0_ ) | ( (~ Poutreg_14_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n835 = ( (~ Pdata_33_)  &  PC_10_ ) | ( Pdata_33_  &  (~ PC_10_) ) ;
 assign n834 = ( n274  &  n266 ) | ( n274  &  n835 ) ;
 assign n837 = ( (~ n254)  &  n297 ) | ( n254  &  (~ n1384) ) | ( n297  &  (~ n1384) ) ;
 assign n838 = ( n296  &  (~ n1203) ) ;
 assign n839 = ( n275 ) | ( (~ n835) ) | ( n1647 ) | ( n1648 ) ;
 assign n841 = ( n244  &  (~ n266) ) | ( n244  &  n1202 ) ;
 assign n836 = ( n257  &  n837  &  n838  &  n839  &  n841  &  (~ n1649) ) ;
 assign n843 = ( (~ Poutreg_21_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_21_)  &  n1529 ) | ( n126  &  n1529 ) ;
 assign n845 = ( (~ Poutreg_20_)  &  (~ Poutreg_12_) ) | ( (~ Poutreg_20_)  &  Pcount_0_ ) | ( (~ Poutreg_12_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n847 = ( (~ n459) ) | ( n475 ) | ( (~ n675) ) ;
 assign n846 = ( n459  &  n847 ) | ( (~ n475)  &  n847 ) ;
 assign n849 = ( (~ n460)  &  n491 ) ;
 assign n848 = ( (~ n459)  &  n675  &  n849 ) ;
 assign n851 = ( (~ n475)  &  (~ n675) ) ;
 assign n852 = ( n460  &  n675  &  n475 ) ;
 assign n850 = ( n851  &  (~ n1249) ) | ( n852  &  (~ n1249) ) ;
 assign n855 = ( (~ Poutreg_19_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_19_)  &  n1533 ) | ( n126  &  n1533 ) ;
 assign n857 = ( (~ Poutreg_18_)  &  (~ Poutreg_10_) ) | ( (~ Poutreg_18_)  &  Pcount_0_ ) | ( (~ Poutreg_10_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n858 = ( n772  &  n781  &  n780 ) ;
 assign n859 = ( n607  &  (~ n605)  &  n777 ) ;
 assign n862 = ( n1166  &  n629 ) ;
 assign n863 = ( n605  &  n1167 ) | ( n605  &  n1325 ) | ( (~ n1167)  &  n1325 ) ;
 assign n860 = ( (~ n775)  &  n862  &  n863 ) ;
 assign n866 = ( n777  &  (~ n776)  &  (~ n1166) ) ;
 assign n864 = ( (~ n766)  &  n866 ) | ( (~ n766)  &  (~ n878) ) ;
 assign n869 = ( (~ Poutreg_17_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_17_)  &  (~ n1719) ) | ( n126  &  (~ n1719) ) ;
 assign n871 = ( (~ Poutreg_16_)  &  (~ Poutreg_8_) ) | ( (~ Poutreg_16_)  &  Pcount_0_ ) | ( (~ Poutreg_8_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n874 = ( (~ n775) ) | ( (~ n1300) ) | ( n1325 ) ;
 assign n875 = ( n1297 ) | ( n775 ) ;
 assign n873 = ( n775 ) | ( n615 ) ;
 assign n872 = ( (~ n862)  &  n874  &  n875 ) | ( n874  &  n875  &  n873 ) ;
 assign n877 = ( n629  &  n1654 ) | ( (~ n776)  &  n1654 ) | ( n1292  &  n1654 ) ;
 assign n878 = ( (~ n775) ) | ( n1289 ) ;
 assign n876 = ( (~ n866)  &  (~ n1166) ) | ( (~ n866)  &  n877  &  n878 ) ;
 assign n879 = ( n615 ) | ( n629 ) | ( (~ n777) ) ;
 assign n880 = ( n781  &  (~ n1298) ) | ( n781  &  (~ n1301) ) ;
 assign n884 = ( (~ Poutreg_15_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_15_)  &  n1538 ) | ( n126  &  n1538 ) ;
 assign n886 = ( (~ Poutreg_14_)  &  (~ Poutreg_6_) ) | ( (~ Poutreg_14_)  &  Pcount_0_ ) | ( (~ Poutreg_6_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n888 = ( n751  &  (~ n895) ) ;
 assign n887 = ( (~ n756)  &  n888 ) ;
 assign n889 = ( n725 ) | ( n811 ) ;
 assign n891 = ( (~ Poutreg_13_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_13_)  &  n1539 ) | ( n126  &  n1539 ) ;
 assign n893 = ( (~ Poutreg_12_)  &  (~ Poutreg_4_) ) | ( (~ Poutreg_12_)  &  Pcount_0_ ) | ( (~ Poutreg_4_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n896 = ( n801 ) | ( (~ n895) ) ;
 assign n895 = ( (~ Pdata_43_)  &  PC_25_ ) | ( Pdata_43_  &  (~ PC_25_) ) ;
 assign n894 = ( (~ n725)  &  (~ n756)  &  n896 ) | ( (~ n756)  &  n896  &  n895 ) ;
 assign n898 = ( n711 ) | ( (~ n895) ) ;
 assign n897 = ( (~ n738)  &  n743  &  (~ n894) ) | ( n743  &  (~ n894)  &  n898 ) ;
 assign n901 = ( n741  &  n804  &  n808  &  n1319 ) ;
 assign n902 = ( (~ n742)  &  n754 ) | ( n742  &  n897 ) | ( n754  &  n897 ) ;
 assign n903 = ( n724 ) | ( (~ n751) ) | ( n1340 ) ;
 assign n904 = ( n710 ) | ( (~ n719) ) | ( (~ n1169) ) ;
 assign n905 = ( n895  &  n746 ) | ( n1341  &  n746 ) | ( n895  &  n1318 ) | ( n1341  &  n1318 ) ;
 assign n900 = ( n901  &  n723  &  n902  &  n903  &  n904  &  n905 ) ;
 assign n907 = ( (~ Poutreg_11_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_11_)  &  n1540 ) | ( n126  &  n1540 ) ;
 assign n909 = ( (~ Poutreg_10_)  &  (~ Poutreg_2_) ) | ( (~ Poutreg_10_)  &  Pcount_0_ ) | ( (~ Poutreg_2_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n912 = ( (~ n201)  &  n914 ) ;
 assign n911 = ( n220  &  (~ n1156) ) ;
 assign n910 = ( n231  &  n912  &  n911 ) | ( n231  &  n912  &  n207 ) ;
 assign n914 = ( (~ Pdata_47_)  &  PD_12_ ) | ( Pdata_47_  &  (~ PD_12_) ) ;
 assign n915 = ( (~ Pdata_52_)  &  PD_26_ ) | ( Pdata_52_  &  (~ PD_26_) ) ;
 assign n913 = ( n914 ) | ( n915 ) | ( (~ n1660) ) ;
 assign n917 = ( n212 ) | ( (~ n226) ) ;
 assign n920 = ( (~ Poutreg_9_)  &  n1 ) | ( n1  &  n126 ) | ( (~ Poutreg_9_)  &  n1541 ) | ( n126  &  n1541 ) ;
 assign n922 = ( (~ Poutreg_8_)  &  (~ Poutreg_0_) ) | ( (~ Poutreg_8_)  &  Pcount_0_ ) | ( (~ Poutreg_0_)  &  n126 ) | ( Pcount_0_  &  n126 ) ;
 assign n925 = ( Pcount_0_ ) | ( n924 ) ;
 assign n924 = ( n92 ) | ( Preset_0_ ) ;
 assign n923 = ( n925  &  Pcount_1_ ) | ( n925  &  n924 ) ;
 assign n926 = ( n923  &  Pcount_2_ ) | ( n923  &  n924 ) ;
 assign n928 = ( Pcount_3_ ) | ( n1177 ) ;
 assign n929 = ( Pcount_0_  &  n1  &  n928 ) | ( n1  &  n928  &  (~ n1453) ) ;
 assign n932 = ( (~ PC_26_)  &  (~ PC_0_) ) | ( (~ PC_0_)  &  n1352 ) | ( (~ PC_26_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n933 = ( (~ PC_25_)  &  (~ PC_1_) ) | ( (~ PC_1_)  &  n1348 ) | ( (~ PC_25_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n934 = ( (~ PC_27_)  &  n1542 ) | ( n1359  &  n1542 ) ;
 assign n931 = ( n932  &  n933  &  n934 ) ;
 assign n936 = ( (~ PC_27_)  &  (~ PC_25_) ) | ( (~ PC_27_)  &  n1352 ) | ( (~ PC_25_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n937 = ( (~ PC_24_)  &  (~ PC_0_) ) | ( (~ PC_0_)  &  n1348 ) | ( (~ PC_24_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n938 = ( (~ PC_26_)  &  n1543 ) | ( n1359  &  n1543 ) ;
 assign n935 = ( n936  &  n937  &  n938 ) ;
 assign n940 = ( (~ PC_26_)  &  (~ PC_24_) ) | ( (~ PC_26_)  &  n1352 ) | ( (~ PC_24_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n941 = ( (~ PC_27_)  &  (~ PC_23_) ) | ( (~ PC_27_)  &  n1348 ) | ( (~ PC_23_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n942 = ( (~ PC_25_)  &  n1544 ) | ( n1359  &  n1544 ) ;
 assign n939 = ( n940  &  n941  &  n942 ) ;
 assign n944 = ( (~ PC_25_)  &  (~ PC_23_) ) | ( (~ PC_25_)  &  n1352 ) | ( (~ PC_23_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n945 = ( (~ PC_26_)  &  (~ PC_22_) ) | ( (~ PC_26_)  &  n1348 ) | ( (~ PC_22_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n946 = ( (~ PC_24_)  &  n1545 ) | ( n1359  &  n1545 ) ;
 assign n943 = ( n944  &  n945  &  n946 ) ;
 assign n948 = ( (~ PC_24_)  &  (~ PC_22_) ) | ( (~ PC_24_)  &  n1352 ) | ( (~ PC_22_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n949 = ( (~ PC_25_)  &  (~ PC_21_) ) | ( (~ PC_25_)  &  n1348 ) | ( (~ PC_21_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n950 = ( (~ PC_23_)  &  n1546 ) | ( n1359  &  n1546 ) ;
 assign n947 = ( n948  &  n949  &  n950 ) ;
 assign n952 = ( (~ PC_23_)  &  (~ PC_21_) ) | ( (~ PC_23_)  &  n1352 ) | ( (~ PC_21_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n953 = ( (~ PC_24_)  &  (~ PC_20_) ) | ( (~ PC_24_)  &  n1348 ) | ( (~ PC_20_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n954 = ( (~ PC_22_)  &  n1547 ) | ( n1359  &  n1547 ) ;
 assign n951 = ( n952  &  n953  &  n954 ) ;
 assign n956 = ( (~ PC_22_)  &  (~ PC_20_) ) | ( (~ PC_22_)  &  n1352 ) | ( (~ PC_20_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n957 = ( (~ PC_23_)  &  (~ PC_19_) ) | ( (~ PC_23_)  &  n1348 ) | ( (~ PC_19_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n958 = ( (~ PC_21_)  &  n1548 ) | ( n1359  &  n1548 ) ;
 assign n955 = ( n956  &  n957  &  n958 ) ;
 assign n960 = ( (~ PC_21_)  &  (~ PC_19_) ) | ( (~ PC_21_)  &  n1352 ) | ( (~ PC_19_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n961 = ( (~ PC_22_)  &  (~ PC_18_) ) | ( (~ PC_22_)  &  n1348 ) | ( (~ PC_18_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n962 = ( (~ PC_20_)  &  n1549 ) | ( n1359  &  n1549 ) ;
 assign n959 = ( n960  &  n961  &  n962 ) ;
 assign n964 = ( (~ PC_20_)  &  (~ PC_18_) ) | ( (~ PC_20_)  &  n1352 ) | ( (~ PC_18_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n965 = ( (~ PC_21_)  &  (~ PC_17_) ) | ( (~ PC_21_)  &  n1348 ) | ( (~ PC_17_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n966 = ( (~ PC_19_)  &  n1550 ) | ( n1359  &  n1550 ) ;
 assign n963 = ( n964  &  n965  &  n966 ) ;
 assign n968 = ( (~ PC_19_)  &  (~ PC_17_) ) | ( (~ PC_19_)  &  n1352 ) | ( (~ PC_17_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n969 = ( (~ PC_20_)  &  (~ PC_16_) ) | ( (~ PC_20_)  &  n1348 ) | ( (~ PC_16_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n970 = ( (~ PC_18_)  &  n1551 ) | ( n1359  &  n1551 ) ;
 assign n967 = ( n968  &  n969  &  n970 ) ;
 assign n972 = ( (~ PC_18_)  &  (~ PC_16_) ) | ( (~ PC_18_)  &  n1352 ) | ( (~ PC_16_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n973 = ( (~ PC_19_)  &  (~ PC_15_) ) | ( (~ PC_19_)  &  n1348 ) | ( (~ PC_15_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n974 = ( (~ PC_17_)  &  n1552 ) | ( n1359  &  n1552 ) ;
 assign n971 = ( n972  &  n973  &  n974 ) ;
 assign n976 = ( (~ PC_17_)  &  (~ PC_15_) ) | ( (~ PC_17_)  &  n1352 ) | ( (~ PC_15_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n977 = ( (~ PC_18_)  &  (~ PC_14_) ) | ( (~ PC_18_)  &  n1348 ) | ( (~ PC_14_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n978 = ( (~ PC_16_)  &  n1553 ) | ( n1359  &  n1553 ) ;
 assign n975 = ( n976  &  n977  &  n978 ) ;
 assign n980 = ( (~ PC_16_)  &  (~ PC_14_) ) | ( (~ PC_16_)  &  n1352 ) | ( (~ PC_14_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n981 = ( (~ PC_17_)  &  (~ PC_13_) ) | ( (~ PC_17_)  &  n1348 ) | ( (~ PC_13_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n982 = ( (~ PC_15_)  &  n1554 ) | ( n1359  &  n1554 ) ;
 assign n979 = ( n980  &  n981  &  n982 ) ;
 assign n984 = ( (~ PC_15_)  &  (~ PC_13_) ) | ( (~ PC_15_)  &  n1352 ) | ( (~ PC_13_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n985 = ( (~ PC_16_)  &  (~ PC_12_) ) | ( (~ PC_16_)  &  n1348 ) | ( (~ PC_12_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n986 = ( (~ PC_14_)  &  n1555 ) | ( n1359  &  n1555 ) ;
 assign n983 = ( n984  &  n985  &  n986 ) ;
 assign n988 = ( (~ PC_14_)  &  (~ PC_12_) ) | ( (~ PC_14_)  &  n1352 ) | ( (~ PC_12_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n989 = ( (~ PC_15_)  &  (~ PC_11_) ) | ( (~ PC_15_)  &  n1348 ) | ( (~ PC_11_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n990 = ( (~ PC_13_)  &  n1556 ) | ( n1359  &  n1556 ) ;
 assign n987 = ( n988  &  n989  &  n990 ) ;
 assign n992 = ( (~ PC_13_)  &  (~ PC_11_) ) | ( (~ PC_13_)  &  n1352 ) | ( (~ PC_11_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n993 = ( (~ PC_14_)  &  (~ PC_10_) ) | ( (~ PC_14_)  &  n1348 ) | ( (~ PC_10_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n994 = ( (~ PC_12_)  &  n1557 ) | ( n1359  &  n1557 ) ;
 assign n991 = ( n992  &  n993  &  n994 ) ;
 assign n996 = ( (~ PC_12_)  &  (~ PC_10_) ) | ( (~ PC_12_)  &  n1352 ) | ( (~ PC_10_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n997 = ( (~ PC_13_)  &  (~ PC_9_) ) | ( (~ PC_13_)  &  n1348 ) | ( (~ PC_9_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n998 = ( (~ PC_11_)  &  n1558 ) | ( n1359  &  n1558 ) ;
 assign n995 = ( n996  &  n997  &  n998 ) ;
 assign n1000 = ( (~ PC_11_)  &  (~ PC_9_) ) | ( (~ PC_11_)  &  n1352 ) | ( (~ PC_9_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1001 = ( (~ PC_12_)  &  (~ PC_8_) ) | ( (~ PC_12_)  &  n1348 ) | ( (~ PC_8_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1002 = ( (~ PC_10_)  &  n1559 ) | ( n1359  &  n1559 ) ;
 assign n999 = ( n1000  &  n1001  &  n1002 ) ;
 assign n1004 = ( (~ PC_10_)  &  (~ PC_8_) ) | ( (~ PC_10_)  &  n1352 ) | ( (~ PC_8_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1005 = ( (~ PC_11_)  &  (~ PC_7_) ) | ( (~ PC_11_)  &  n1348 ) | ( (~ PC_7_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1006 = ( (~ PC_9_)  &  n1560 ) | ( n1359  &  n1560 ) ;
 assign n1003 = ( n1004  &  n1005  &  n1006 ) ;
 assign n1008 = ( (~ PC_9_)  &  (~ PC_7_) ) | ( (~ PC_9_)  &  n1352 ) | ( (~ PC_7_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1009 = ( (~ PC_10_)  &  (~ PC_6_) ) | ( (~ PC_10_)  &  n1348 ) | ( (~ PC_6_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1010 = ( (~ PC_8_)  &  n1561 ) | ( n1359  &  n1561 ) ;
 assign n1007 = ( n1008  &  n1009  &  n1010 ) ;
 assign n1012 = ( (~ PC_8_)  &  (~ PC_6_) ) | ( (~ PC_8_)  &  n1352 ) | ( (~ PC_6_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1013 = ( (~ PC_9_)  &  (~ PC_5_) ) | ( (~ PC_9_)  &  n1348 ) | ( (~ PC_5_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1014 = ( (~ PC_7_)  &  n1562 ) | ( n1359  &  n1562 ) ;
 assign n1011 = ( n1012  &  n1013  &  n1014 ) ;
 assign n1016 = ( (~ PC_7_)  &  (~ PC_5_) ) | ( (~ PC_7_)  &  n1352 ) | ( (~ PC_5_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1017 = ( (~ PC_8_)  &  (~ PC_4_) ) | ( (~ PC_8_)  &  n1348 ) | ( (~ PC_4_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1018 = ( (~ PC_6_)  &  n1563 ) | ( n1359  &  n1563 ) ;
 assign n1015 = ( n1016  &  n1017  &  n1018 ) ;
 assign n1020 = ( (~ PC_6_)  &  (~ PC_4_) ) | ( (~ PC_6_)  &  n1352 ) | ( (~ PC_4_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1021 = ( (~ PC_7_)  &  (~ PC_3_) ) | ( (~ PC_7_)  &  n1348 ) | ( (~ PC_3_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1022 = ( (~ PC_5_)  &  n1564 ) | ( n1359  &  n1564 ) ;
 assign n1019 = ( n1020  &  n1021  &  n1022 ) ;
 assign n1024 = ( (~ PC_5_)  &  (~ PC_3_) ) | ( (~ PC_5_)  &  n1352 ) | ( (~ PC_3_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1025 = ( (~ PC_6_)  &  (~ PC_2_) ) | ( (~ PC_6_)  &  n1348 ) | ( (~ PC_2_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1026 = ( (~ PC_4_)  &  n1565 ) | ( n1359  &  n1565 ) ;
 assign n1023 = ( n1024  &  n1025  &  n1026 ) ;
 assign n1028 = ( (~ PC_4_)  &  (~ PC_2_) ) | ( (~ PC_4_)  &  n1352 ) | ( (~ PC_2_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1029 = ( (~ PC_5_)  &  (~ PC_1_) ) | ( (~ PC_5_)  &  n1348 ) | ( (~ PC_1_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1030 = ( (~ PC_3_)  &  n1566 ) | ( n1359  &  n1566 ) ;
 assign n1027 = ( n1028  &  n1029  &  n1030 ) ;
 assign n1032 = ( (~ PC_3_)  &  (~ PC_1_) ) | ( (~ PC_3_)  &  n1352 ) | ( (~ PC_1_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1033 = ( (~ PC_4_)  &  (~ PC_0_) ) | ( (~ PC_4_)  &  n1348 ) | ( (~ PC_0_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1034 = ( (~ PC_2_)  &  n1567 ) | ( n1359  &  n1567 ) ;
 assign n1031 = ( n1032  &  n1033  &  n1034 ) ;
 assign n1036 = ( (~ PC_2_)  &  (~ PC_0_) ) | ( (~ PC_2_)  &  n1352 ) | ( (~ PC_0_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1037 = ( (~ PC_27_)  &  (~ PC_3_) ) | ( (~ PC_3_)  &  n1348 ) | ( (~ PC_27_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1038 = ( (~ PC_1_)  &  n1568 ) | ( n1359  &  n1568 ) ;
 assign n1035 = ( n1036  &  n1037  &  n1038 ) ;
 assign n1040 = ( (~ PC_27_)  &  (~ PC_1_) ) | ( (~ PC_1_)  &  n1352 ) | ( (~ PC_27_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1041 = ( (~ PC_26_)  &  (~ PC_2_) ) | ( (~ PC_2_)  &  n1348 ) | ( (~ PC_26_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1042 = ( (~ PC_0_)  &  n1569 ) | ( n1359  &  n1569 ) ;
 assign n1039 = ( n1040  &  n1041  &  n1042 ) ;
 assign n1044 = ( (~ PD_26_)  &  (~ PD_0_) ) | ( (~ PD_0_)  &  n1352 ) | ( (~ PD_26_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1045 = ( (~ PD_25_)  &  (~ PD_1_) ) | ( (~ PD_1_)  &  n1348 ) | ( (~ PD_25_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1046 = ( (~ PD_27_)  &  n1570 ) | ( n1359  &  n1570 ) ;
 assign n1043 = ( n1044  &  n1045  &  n1046 ) ;
 assign n1048 = ( (~ PD_27_)  &  (~ PD_25_) ) | ( (~ PD_27_)  &  n1352 ) | ( (~ PD_25_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1049 = ( (~ PD_24_)  &  (~ PD_0_) ) | ( (~ PD_0_)  &  n1348 ) | ( (~ PD_24_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1050 = ( (~ PD_26_)  &  n1571 ) | ( n1359  &  n1571 ) ;
 assign n1047 = ( n1048  &  n1049  &  n1050 ) ;
 assign n1052 = ( (~ PD_26_)  &  (~ PD_24_) ) | ( (~ PD_26_)  &  n1352 ) | ( (~ PD_24_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1053 = ( (~ PD_27_)  &  (~ PD_23_) ) | ( (~ PD_27_)  &  n1348 ) | ( (~ PD_23_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1054 = ( (~ PD_25_)  &  n1572 ) | ( n1359  &  n1572 ) ;
 assign n1051 = ( n1052  &  n1053  &  n1054 ) ;
 assign n1056 = ( (~ PD_25_)  &  (~ PD_23_) ) | ( (~ PD_25_)  &  n1352 ) | ( (~ PD_23_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1057 = ( (~ PD_26_)  &  (~ PD_22_) ) | ( (~ PD_26_)  &  n1348 ) | ( (~ PD_22_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1058 = ( (~ PD_24_)  &  n1573 ) | ( n1359  &  n1573 ) ;
 assign n1055 = ( n1056  &  n1057  &  n1058 ) ;
 assign n1060 = ( (~ PD_24_)  &  (~ PD_22_) ) | ( (~ PD_24_)  &  n1352 ) | ( (~ PD_22_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1061 = ( (~ PD_25_)  &  (~ PD_21_) ) | ( (~ PD_25_)  &  n1348 ) | ( (~ PD_21_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1062 = ( (~ PD_23_)  &  n1574 ) | ( n1359  &  n1574 ) ;
 assign n1059 = ( n1060  &  n1061  &  n1062 ) ;
 assign n1064 = ( (~ PD_23_)  &  (~ PD_21_) ) | ( (~ PD_23_)  &  n1352 ) | ( (~ PD_21_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1065 = ( (~ PD_24_)  &  (~ PD_20_) ) | ( (~ PD_24_)  &  n1348 ) | ( (~ PD_20_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1066 = ( (~ PD_22_)  &  n1575 ) | ( n1359  &  n1575 ) ;
 assign n1063 = ( n1064  &  n1065  &  n1066 ) ;
 assign n1068 = ( (~ PD_22_)  &  (~ PD_20_) ) | ( (~ PD_22_)  &  n1352 ) | ( (~ PD_20_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1069 = ( (~ PD_23_)  &  (~ PD_19_) ) | ( (~ PD_23_)  &  n1348 ) | ( (~ PD_19_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1070 = ( (~ PD_21_)  &  n1576 ) | ( n1359  &  n1576 ) ;
 assign n1067 = ( n1068  &  n1069  &  n1070 ) ;
 assign n1072 = ( (~ PD_21_)  &  (~ PD_19_) ) | ( (~ PD_21_)  &  n1352 ) | ( (~ PD_19_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1073 = ( (~ PD_22_)  &  (~ PD_18_) ) | ( (~ PD_22_)  &  n1348 ) | ( (~ PD_18_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1074 = ( (~ PD_20_)  &  n1577 ) | ( n1359  &  n1577 ) ;
 assign n1071 = ( n1072  &  n1073  &  n1074 ) ;
 assign n1076 = ( (~ PD_20_)  &  (~ PD_18_) ) | ( (~ PD_20_)  &  n1352 ) | ( (~ PD_18_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1077 = ( (~ PD_21_)  &  (~ PD_17_) ) | ( (~ PD_21_)  &  n1348 ) | ( (~ PD_17_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1078 = ( (~ PD_19_)  &  n1578 ) | ( n1359  &  n1578 ) ;
 assign n1075 = ( n1076  &  n1077  &  n1078 ) ;
 assign n1080 = ( (~ PD_19_)  &  (~ PD_17_) ) | ( (~ PD_19_)  &  n1352 ) | ( (~ PD_17_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1081 = ( (~ PD_20_)  &  (~ PD_16_) ) | ( (~ PD_20_)  &  n1348 ) | ( (~ PD_16_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1082 = ( (~ PD_18_)  &  n1579 ) | ( n1359  &  n1579 ) ;
 assign n1079 = ( n1080  &  n1081  &  n1082 ) ;
 assign n1084 = ( (~ PD_18_)  &  (~ PD_16_) ) | ( (~ PD_18_)  &  n1352 ) | ( (~ PD_16_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1085 = ( (~ PD_19_)  &  (~ PD_15_) ) | ( (~ PD_19_)  &  n1348 ) | ( (~ PD_15_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1086 = ( (~ PD_17_)  &  n1580 ) | ( n1359  &  n1580 ) ;
 assign n1083 = ( n1084  &  n1085  &  n1086 ) ;
 assign n1088 = ( (~ PD_17_)  &  (~ PD_15_) ) | ( (~ PD_17_)  &  n1352 ) | ( (~ PD_15_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1089 = ( (~ PD_18_)  &  (~ PD_14_) ) | ( (~ PD_18_)  &  n1348 ) | ( (~ PD_14_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1090 = ( (~ PD_16_)  &  n1581 ) | ( n1359  &  n1581 ) ;
 assign n1087 = ( n1088  &  n1089  &  n1090 ) ;
 assign n1092 = ( (~ PD_16_)  &  (~ PD_14_) ) | ( (~ PD_16_)  &  n1352 ) | ( (~ PD_14_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1093 = ( (~ PD_17_)  &  (~ PD_13_) ) | ( (~ PD_17_)  &  n1348 ) | ( (~ PD_13_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1094 = ( (~ PD_15_)  &  n1582 ) | ( n1359  &  n1582 ) ;
 assign n1091 = ( n1092  &  n1093  &  n1094 ) ;
 assign n1096 = ( (~ PD_15_)  &  (~ PD_13_) ) | ( (~ PD_15_)  &  n1352 ) | ( (~ PD_13_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1097 = ( (~ PD_16_)  &  (~ PD_12_) ) | ( (~ PD_16_)  &  n1348 ) | ( (~ PD_12_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1098 = ( (~ PD_14_)  &  n1583 ) | ( n1359  &  n1583 ) ;
 assign n1095 = ( n1096  &  n1097  &  n1098 ) ;
 assign n1100 = ( (~ PD_14_)  &  (~ PD_12_) ) | ( (~ PD_14_)  &  n1352 ) | ( (~ PD_12_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1101 = ( (~ PD_15_)  &  (~ PD_11_) ) | ( (~ PD_15_)  &  n1348 ) | ( (~ PD_11_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1102 = ( (~ PD_13_)  &  n1584 ) | ( n1359  &  n1584 ) ;
 assign n1099 = ( n1100  &  n1101  &  n1102 ) ;
 assign n1104 = ( (~ PD_13_)  &  (~ PD_11_) ) | ( (~ PD_13_)  &  n1352 ) | ( (~ PD_11_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1105 = ( (~ PD_14_)  &  (~ PD_10_) ) | ( (~ PD_14_)  &  n1348 ) | ( (~ PD_10_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1106 = ( (~ PD_12_)  &  n1585 ) | ( n1359  &  n1585 ) ;
 assign n1103 = ( n1104  &  n1105  &  n1106 ) ;
 assign n1108 = ( (~ PD_12_)  &  (~ PD_10_) ) | ( (~ PD_12_)  &  n1352 ) | ( (~ PD_10_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1109 = ( (~ PD_13_)  &  (~ PD_9_) ) | ( (~ PD_13_)  &  n1348 ) | ( (~ PD_9_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1110 = ( (~ PD_11_)  &  n1586 ) | ( n1359  &  n1586 ) ;
 assign n1107 = ( n1108  &  n1109  &  n1110 ) ;
 assign n1112 = ( (~ PD_11_)  &  (~ PD_9_) ) | ( (~ PD_11_)  &  n1352 ) | ( (~ PD_9_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1113 = ( (~ PD_12_)  &  (~ PD_8_) ) | ( (~ PD_12_)  &  n1348 ) | ( (~ PD_8_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1114 = ( (~ PD_10_)  &  n1587 ) | ( n1359  &  n1587 ) ;
 assign n1111 = ( n1112  &  n1113  &  n1114 ) ;
 assign n1116 = ( (~ PD_10_)  &  (~ PD_8_) ) | ( (~ PD_10_)  &  n1352 ) | ( (~ PD_8_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1117 = ( (~ PD_11_)  &  (~ PD_7_) ) | ( (~ PD_11_)  &  n1348 ) | ( (~ PD_7_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1118 = ( (~ PD_9_)  &  n1588 ) | ( n1359  &  n1588 ) ;
 assign n1115 = ( n1116  &  n1117  &  n1118 ) ;
 assign n1120 = ( (~ PD_9_)  &  (~ PD_7_) ) | ( (~ PD_9_)  &  n1352 ) | ( (~ PD_7_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1121 = ( (~ PD_10_)  &  (~ PD_6_) ) | ( (~ PD_10_)  &  n1348 ) | ( (~ PD_6_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1122 = ( (~ PD_8_)  &  n1589 ) | ( n1359  &  n1589 ) ;
 assign n1119 = ( n1120  &  n1121  &  n1122 ) ;
 assign n1124 = ( (~ PD_8_)  &  (~ PD_6_) ) | ( (~ PD_8_)  &  n1352 ) | ( (~ PD_6_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1125 = ( (~ PD_9_)  &  (~ PD_5_) ) | ( (~ PD_9_)  &  n1348 ) | ( (~ PD_5_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1126 = ( (~ PD_7_)  &  n1590 ) | ( n1359  &  n1590 ) ;
 assign n1123 = ( n1124  &  n1125  &  n1126 ) ;
 assign n1128 = ( (~ PD_7_)  &  (~ PD_5_) ) | ( (~ PD_7_)  &  n1352 ) | ( (~ PD_5_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1129 = ( (~ PD_8_)  &  (~ PD_4_) ) | ( (~ PD_8_)  &  n1348 ) | ( (~ PD_4_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1130 = ( (~ PD_6_)  &  n1591 ) | ( n1359  &  n1591 ) ;
 assign n1127 = ( n1128  &  n1129  &  n1130 ) ;
 assign n1132 = ( (~ PD_6_)  &  (~ PD_4_) ) | ( (~ PD_6_)  &  n1352 ) | ( (~ PD_4_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1133 = ( (~ PD_7_)  &  (~ PD_3_) ) | ( (~ PD_7_)  &  n1348 ) | ( (~ PD_3_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1134 = ( (~ PD_5_)  &  n1592 ) | ( n1359  &  n1592 ) ;
 assign n1131 = ( n1132  &  n1133  &  n1134 ) ;
 assign n1136 = ( (~ PD_5_)  &  (~ PD_3_) ) | ( (~ PD_5_)  &  n1352 ) | ( (~ PD_3_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1137 = ( (~ PD_6_)  &  (~ PD_2_) ) | ( (~ PD_6_)  &  n1348 ) | ( (~ PD_2_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1138 = ( (~ PD_4_)  &  n1593 ) | ( n1359  &  n1593 ) ;
 assign n1135 = ( n1136  &  n1137  &  n1138 ) ;
 assign n1140 = ( (~ PD_4_)  &  (~ PD_2_) ) | ( (~ PD_4_)  &  n1352 ) | ( (~ PD_2_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1141 = ( (~ PD_5_)  &  (~ PD_1_) ) | ( (~ PD_5_)  &  n1348 ) | ( (~ PD_1_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1142 = ( (~ PD_3_)  &  n1594 ) | ( n1359  &  n1594 ) ;
 assign n1139 = ( n1140  &  n1141  &  n1142 ) ;
 assign n1144 = ( (~ PD_3_)  &  (~ PD_1_) ) | ( (~ PD_3_)  &  n1352 ) | ( (~ PD_1_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1145 = ( (~ PD_4_)  &  (~ PD_0_) ) | ( (~ PD_4_)  &  n1348 ) | ( (~ PD_0_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1146 = ( (~ PD_2_)  &  n1595 ) | ( n1359  &  n1595 ) ;
 assign n1143 = ( n1144  &  n1145  &  n1146 ) ;
 assign n1148 = ( (~ PD_2_)  &  (~ PD_0_) ) | ( (~ PD_2_)  &  n1352 ) | ( (~ PD_0_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1149 = ( (~ PD_27_)  &  (~ PD_3_) ) | ( (~ PD_3_)  &  n1348 ) | ( (~ PD_27_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1150 = ( (~ PD_1_)  &  n1596 ) | ( n1359  &  n1596 ) ;
 assign n1147 = ( n1148  &  n1149  &  n1150 ) ;
 assign n1152 = ( (~ PD_27_)  &  (~ PD_1_) ) | ( (~ PD_1_)  &  n1352 ) | ( (~ PD_27_)  &  n1353 ) | ( n1352  &  n1353 ) ;
 assign n1153 = ( (~ PD_26_)  &  (~ PD_2_) ) | ( (~ PD_2_)  &  n1348 ) | ( (~ PD_26_)  &  n1351 ) | ( n1348  &  n1351 ) ;
 assign n1154 = ( (~ PD_0_)  &  n1597 ) | ( n1359  &  n1597 ) ;
 assign n1151 = ( n1152  &  n1153  &  n1154 ) ;
 assign n1155 = ( (~ Pdata_48_)  &  PD_23_ ) | ( Pdata_48_  &  (~ PD_23_) ) ;
 assign n1156 = ( (~ Pdata_51_)  &  PD_18_ ) | ( Pdata_51_  &  (~ PD_18_) ) ;
 assign n1158 = ( (~ Pdata_45_)  &  PC_26_ ) | ( Pdata_45_  &  (~ PC_26_) ) ;
 assign n1159 = ( (~ Pdata_38_)  &  PC_5_ ) | ( Pdata_38_  &  (~ PC_5_) ) ;
 assign n1160 = ( n375  &  (~ n385) ) | ( n375  &  n432  &  (~ n572) ) ;
 assign n1163 = ( (~ Pdata_52_)  &  PD_11_ ) | ( Pdata_52_  &  (~ PD_11_) ) ;
 assign n1164 = ( (~ Pdata_56_)  &  PD_19_ ) | ( Pdata_56_  &  (~ PD_19_) ) ;
 assign n1165 = ( (~ n1164)  &  n546 ) | ( n1164  &  (~ n546) ) ;
 assign n1166 = ( (~ Pdata_60_)  &  PD_24_ ) | ( Pdata_60_  &  (~ PD_24_) ) ;
 assign n1167 = ( (~ Pdata_58_)  &  PD_27_ ) | ( Pdata_58_  &  (~ PD_27_) ) ;
 assign n1168 = ( n460  &  n475 ) | ( (~ n460)  &  (~ n475) ) ;
 assign n1169 = ( (~ Pdata_42_)  &  PC_3_ ) | ( Pdata_42_  &  (~ PC_3_) ) ;
 assign n1170 = ( (~ n220)  &  (~ n1184) ) | ( (~ n1155)  &  (~ n1184) ) ;
 assign n1172 = ( n254  &  n835 ) | ( (~ n254)  &  (~ n835) ) ;
 assign n1173 = ( Pencrypt_mode_0_  &  Pencrypt_0_ ) | ( (~ Pencrypt_mode_0_)  &  (~ Pencrypt_0_) ) ;
 assign n1177 = ( (~ Pcount_2_) ) | ( (~ Pcount_1_) ) | ( (~ Pcount_0_) ) ;
 assign n1184 = ( (~ n220)  &  (~ n1156) ) ;
 assign n1185 = ( n220  &  n1156 ) ;
 assign n1186 = ( (~ n915)  &  (~ n1155) ) ;
 assign n1187 = ( n1184  &  n209 ) ;
 assign n1188 = ( (~ n201) ) | ( (~ n914) ) | ( n915 ) ;
 assign n1189 = ( (~ n201) ) | ( (~ n209) ) | ( (~ n914) ) ;
 assign n1198 = ( n269 ) | ( (~ n275) ) | ( (~ n835) ) ;
 assign n1199 = ( n275  &  n240 ) ;
 assign n1200 = ( n266  &  (~ n835) ) ;
 assign n1201 = ( (~ n266)  &  n269  &  (~ n275) ) ;
 assign n1202 = ( n275 ) | ( (~ n274) ) | ( (~ n835) ) ;
 assign n1204 = ( (~ n254)  &  n266  &  n1199 ) ;
 assign n1205 = ( n1200  &  n295  &  n254 ) ;
 assign n1203 = ( n278 ) | ( n280 ) | ( n1204 ) | ( n1205 ) ;
 assign n1215 = ( n357 ) | ( n343 ) ;
 assign n1216 = ( n343 ) | ( (~ n357) ) ;
 assign n1217 = ( (~ n357) ) | ( n1158 ) ;
 assign n1218 = ( n420 ) | ( n357 ) | ( n323 ) ;
 assign n1219 = ( n323 ) | ( n355 ) | ( n1217 ) ;
 assign n1220 = ( n323 ) | ( n326 ) | ( n1216 ) ;
 assign n1221 = ( n323 ) | ( (~ n357) ) | ( n420 ) | ( (~ n1158) ) ;
 assign n1232 = ( n375 ) | ( n570 ) ;
 assign n1234 = ( n369 ) | ( n375 ) ;
 assign n1246 = ( n475  &  (~ n675) ) ;
 assign n1248 = ( (~ n459) ) | ( n470 ) ;
 assign n1249 = ( (~ n459) ) | ( n491 ) ;
 assign n1250 = ( (~ n460)  &  (~ n1249) ) ;
 assign n1251 = ( n477 ) | ( n847 ) ;
 assign n1252 = ( n459  &  n491 ) ;
 assign n1254 = ( n484  &  n487  &  (~ n489) ) ;
 assign n1257 = ( n470 ) | ( (~ n475) ) | ( n477 ) ;
 assign n1258 = ( (~ n477) ) | ( n491 ) | ( n847 ) ;
 assign n1265 = ( (~ n510)  &  (~ n531) ) ;
 assign n1270 = ( n531  &  n546 ) ;
 assign n1272 = ( n510  &  n1270 ) ;
 assign n1273 = ( (~ n510) ) | ( n532 ) ;
 assign n1274 = ( (~ n546) ) | ( (~ n1265) ) ;
 assign n1275 = ( (~ n515) ) | ( n546 ) ;
 assign n1281 = ( n369 ) | ( (~ n382) ) ;
 assign n1289 = ( n629 ) | ( n776 ) | ( (~ n1167) ) ;
 assign n1292 = ( n775 ) | ( (~ n1167) ) ;
 assign n1293 = ( n776  &  n766 ) ;
 assign n1295 = ( (~ n775)  &  (~ n1289) ) ;
 assign n1297 = ( (~ n605) ) | ( (~ n781) ) ;
 assign n1298 = ( n615 ) | ( (~ n780) ) ;
 assign n1300 = ( (~ n607)  &  (~ n781) ) ;
 assign n1301 = ( n873 ) | ( n1167 ) ;
 assign n1303 = ( n1164  &  n546 ) ;
 assign n1318 = ( n895 ) | ( n729 ) ;
 assign n1319 = ( n735  &  n737  &  n728  &  n731 ) ;
 assign n1321 = ( n1319  &  n723  &  n714 ) ;
 assign n1323 = ( n781  &  (~ n1167)  &  n1293 ) ;
 assign n1324 = ( n629 ) | ( n1301 ) ;
 assign n1325 = ( (~ n605)  &  (~ n1293) ) ;
 assign n1326 = ( n625  &  n765  &  n769  &  (~ n771) ) ;
 assign n1329 = ( n215  &  n554 ) ;
 assign n1340 = ( n801 ) | ( n722 ) ;
 assign n1341 = ( (~ n751) ) | ( (~ n814) ) | ( (~ n1340) ) ;
 assign n1345 = ( n924 ) | ( (~ n1358) ) ;
 assign n1347 = ( Pencrypt_mode_0_ ) | ( n1345 ) ;
 assign n1348 = ( (~ n929) ) | ( n1347 ) ;
 assign n1350 = ( (~ Pencrypt_mode_0_) ) | ( n1345 ) ;
 assign n1351 = ( (~ n929) ) | ( n1350 ) ;
 assign n1352 = ( n929 ) | ( n1347 ) ;
 assign n1353 = ( n929 ) | ( n1350 ) ;
 assign n1354 = ( Preset_0_ ) | ( (~ n92) ) ;
 assign n1356 = ( Pencrypt_0_ ) | ( n1354 ) ;
 assign n1357 = ( (~ Pencrypt_0_) ) | ( n1354 ) ;
 assign n1358 = ( n1173 ) | ( n1 ) ;
 assign n1359 = ( n924 ) | ( n1358 ) ;
 assign n1369 = ( (~ n243)  &  n1598 ) | ( n261  &  n1598 ) | ( (~ n269)  &  n1598 ) ;
 assign n1371 = ( (~ n254)  &  (~ n1600) ) | ( n266  &  n295  &  (~ n1600) ) ;
 assign n1372 = ( n281  &  n294 ) | ( n281  &  n835 ) | ( n294  &  (~ n835) ) ;
 assign n1373 = ( n323  &  n328 ) | ( n323  &  (~ n326)  &  n355 ) ;
 assign n1375 = ( n344  &  n357 ) | ( n344  &  (~ n1373) ) | ( (~ n357)  &  (~ n1373) ) ;
 assign n1376 = ( (~ n319)  &  (~ n323) ) | ( (~ n319)  &  (~ n1216) ) | ( n323  &  (~ n1216) ) ;
 assign n1378 = ( n220  &  (~ n1617) ) | ( (~ n228)  &  (~ n1617) ) | ( n914  &  (~ n1617) ) ;
 assign n1380 = ( (~ n878)  &  (~ n1166) ) | ( (~ n878)  &  n1295 ) | ( n1166  &  n1295 ) ;
 assign n1382 = ( n642  &  n1625 ) | ( (~ n647)  &  n1625 ) ;
 assign n1383 = ( (~ n207)  &  (~ n914) ) | ( (~ n207)  &  n1170 ) | ( n914  &  n1170 ) ;
 assign n1384 = ( n275  &  n834 ) | ( n275  &  n1200  &  n262 ) ;
 assign n1385 = ( n228  &  n230 ) | ( (~ n220)  &  n222  &  n228 ) ;
 assign n1386 = ( n228  &  n1185 ) | ( (~ n914)  &  n915  &  n1185 ) ;
 assign n1387 = ( (~ Pdata_in_6_)  &  (~ n1) ) | ( (~ Pdata_in_6_)  &  n1538 ) | ( n1  &  n1538 ) ;
 assign n1388 = ( (~ Pinreg_6_)  &  (~ n1) ) | ( (~ Pinreg_6_)  &  n1528 ) | ( n1  &  n1528 ) ;
 assign n1389 = ( (~ Pinreg_14_)  &  (~ n1) ) | ( (~ Pinreg_14_)  &  n1517 ) | ( n1  &  n1517 ) ;
 assign n1390 = ( (~ Pinreg_22_)  &  (~ n1) ) | ( (~ Pinreg_22_)  &  n1510 ) | ( n1  &  n1510 ) ;
 assign n1391 = ( (~ Pinreg_30_)  &  (~ n1) ) | ( (~ Pinreg_30_)  &  n1503 ) | ( n1  &  n1503 ) ;
 assign n1392 = ( (~ Pinreg_38_)  &  (~ n1) ) | ( (~ Pinreg_38_)  &  n1483 ) | ( n1  &  n1483 ) ;
 assign n1393 = ( (~ Pinreg_46_)  &  (~ n1) ) | ( (~ Pinreg_46_)  &  n1472 ) | ( n1  &  n1472 ) ;
 assign n1394 = ( (~ Pinreg_54_)  &  (~ n1) ) | ( (~ Pinreg_54_)  &  n234 ) | ( n1  &  n234 ) ;
 assign n1395 = ( (~ Pdata_in_4_)  &  (~ n1) ) | ( (~ Pdata_in_4_)  &  n1539 ) | ( n1  &  n1539 ) ;
 assign n1396 = ( (~ Pinreg_4_)  &  (~ n1) ) | ( (~ Pinreg_4_)  &  n1529 ) | ( n1  &  n1529 ) ;
 assign n1397 = ( (~ Pinreg_12_)  &  (~ n1) ) | ( (~ Pinreg_12_)  &  n1521 ) | ( n1  &  n1521 ) ;
 assign n1398 = ( (~ Pinreg_20_)  &  (~ n1) ) | ( (~ Pinreg_20_)  &  n1511 ) | ( n1  &  n1511 ) ;
 assign n1399 = ( (~ Pinreg_28_)  &  (~ n1) ) | ( (~ Pinreg_28_)  &  n1504 ) | ( n1  &  n1504 ) ;
 assign n1400 = ( (~ Pinreg_36_)  &  (~ n1) ) | ( (~ Pinreg_36_)  &  n1494 ) | ( n1  &  n1494 ) ;
 assign n1401 = ( (~ Pinreg_44_)  &  (~ n1) ) | ( (~ Pinreg_44_)  &  n1477 ) | ( n1  &  n1477 ) ;
 assign n1402 = ( (~ Pinreg_52_)  &  (~ n1) ) | ( (~ Pinreg_52_)  &  n287 ) | ( n1  &  n287 ) ;
 assign n1403 = ( (~ Pdata_in_2_)  &  (~ n1) ) | ( (~ Pdata_in_2_)  &  n1540 ) | ( n1  &  n1540 ) ;
 assign n1404 = ( (~ Pinreg_2_)  &  (~ n1) ) | ( (~ Pinreg_2_)  &  n1533 ) | ( n1  &  n1533 ) ;
 assign n1405 = ( (~ Pinreg_10_)  &  (~ n1) ) | ( (~ Pinreg_10_)  &  n1524 ) | ( n1  &  n1524 ) ;
 assign n1406 = ( (~ Pinreg_18_)  &  (~ n1) ) | ( (~ Pinreg_18_)  &  n1512 ) | ( n1  &  n1512 ) ;
 assign n1407 = ( (~ Pinreg_26_)  &  (~ n1) ) | ( (~ Pinreg_26_)  &  n1505 ) | ( n1  &  n1505 ) ;
 assign n1408 = ( (~ Pinreg_34_)  &  (~ n1) ) | ( (~ Pinreg_34_)  &  n1500 ) | ( n1  &  n1500 ) ;
 assign n1409 = ( (~ Pinreg_42_)  &  (~ n1) ) | ( (~ Pinreg_42_)  &  n1478 ) | ( n1  &  n1478 ) ;
 assign n1410 = ( (~ Pinreg_50_)  &  (~ n1) ) | ( (~ Pinreg_50_)  &  n309 ) | ( n1  &  n309 ) ;
 assign n1411 = ( (~ Pdata_in_0_)  &  (~ n1) ) | ( (~ Pdata_in_0_)  &  n1541 ) | ( n1  &  n1541 ) ;
 assign n1412 = ( (~ Pinreg_0_)  &  (~ n1) ) | ( (~ Pinreg_0_)  &  (~ n1719) ) | ( n1  &  (~ n1719) ) ;
 assign n1413 = ( (~ Pinreg_8_)  &  (~ n1) ) | ( (~ Pinreg_8_)  &  (~ n1718) ) | ( n1  &  (~ n1718) ) ;
 assign n1414 = ( (~ Pinreg_16_)  &  (~ n1) ) | ( (~ Pinreg_16_)  &  n1515 ) | ( n1  &  n1515 ) ;
 assign n1415 = ( (~ Pinreg_24_)  &  (~ n1) ) | ( (~ Pinreg_24_)  &  n1507 ) | ( n1  &  n1507 ) ;
 assign n1416 = ( (~ Pinreg_32_)  &  (~ n1) ) | ( (~ Pinreg_32_)  &  (~ n1717) ) | ( n1  &  (~ n1717) ) ;
 assign n1417 = ( (~ Pinreg_40_)  &  (~ n1) ) | ( (~ Pinreg_40_)  &  n1479 ) | ( n1  &  n1479 ) ;
 assign n1418 = ( (~ Pinreg_48_)  &  (~ n1) ) | ( (~ Pinreg_48_)  &  n346 ) | ( n1  &  n346 ) ;
 assign n1419 = ( (~ Pdata_in_7_)  &  (~ Pdata_63_) ) | ( (~ Pdata_63_)  &  n1 ) | ( (~ Pdata_in_7_)  &  (~ n1) ) ;
 assign n1420 = ( (~ Pinreg_7_)  &  (~ Pdata_62_) ) | ( (~ Pdata_62_)  &  n1 ) | ( (~ Pinreg_7_)  &  (~ n1) ) ;
 assign n1421 = ( (~ Pinreg_15_)  &  (~ Pdata_61_) ) | ( (~ Pdata_61_)  &  n1 ) | ( (~ Pinreg_15_)  &  (~ n1) ) ;
 assign n1422 = ( (~ Pinreg_23_)  &  (~ Pdata_60_) ) | ( (~ Pdata_60_)  &  n1 ) | ( (~ Pinreg_23_)  &  (~ n1) ) ;
 assign n1423 = ( (~ Pinreg_31_)  &  (~ Pdata_59_) ) | ( (~ Pdata_59_)  &  n1 ) | ( (~ Pinreg_31_)  &  (~ n1) ) ;
 assign n1424 = ( (~ Pinreg_39_)  &  (~ Pdata_58_) ) | ( (~ Pdata_58_)  &  n1 ) | ( (~ Pinreg_39_)  &  (~ n1) ) ;
 assign n1425 = ( (~ Pinreg_47_)  &  (~ Pdata_57_) ) | ( (~ Pdata_57_)  &  n1 ) | ( (~ Pinreg_47_)  &  (~ n1) ) ;
 assign n1426 = ( (~ Pinreg_55_)  &  (~ Pdata_56_) ) | ( (~ Pdata_56_)  &  n1 ) | ( (~ Pinreg_55_)  &  (~ n1) ) ;
 assign n1427 = ( (~ Pdata_in_5_)  &  (~ Pdata_55_) ) | ( (~ Pdata_55_)  &  n1 ) | ( (~ Pdata_in_5_)  &  (~ n1) ) ;
 assign n1428 = ( (~ Pinreg_5_)  &  (~ Pdata_54_) ) | ( (~ Pdata_54_)  &  n1 ) | ( (~ Pinreg_5_)  &  (~ n1) ) ;
 assign n1429 = ( (~ Pinreg_13_)  &  (~ Pdata_53_) ) | ( (~ Pdata_53_)  &  n1 ) | ( (~ Pinreg_13_)  &  (~ n1) ) ;
 assign n1430 = ( (~ Pinreg_21_)  &  (~ Pdata_52_) ) | ( (~ Pdata_52_)  &  n1 ) | ( (~ Pinreg_21_)  &  (~ n1) ) ;
 assign n1431 = ( (~ Pinreg_29_)  &  (~ Pdata_51_) ) | ( (~ Pdata_51_)  &  n1 ) | ( (~ Pinreg_29_)  &  (~ n1) ) ;
 assign n1432 = ( (~ Pinreg_37_)  &  (~ Pdata_50_) ) | ( (~ Pdata_50_)  &  n1 ) | ( (~ Pinreg_37_)  &  (~ n1) ) ;
 assign n1433 = ( (~ Pinreg_45_)  &  (~ Pdata_49_) ) | ( (~ Pdata_49_)  &  n1 ) | ( (~ Pinreg_45_)  &  (~ n1) ) ;
 assign n1434 = ( (~ Pinreg_53_)  &  (~ Pdata_48_) ) | ( (~ Pdata_48_)  &  n1 ) | ( (~ Pinreg_53_)  &  (~ n1) ) ;
 assign n1435 = ( (~ Pdata_in_3_)  &  (~ Pdata_47_) ) | ( (~ Pdata_47_)  &  n1 ) | ( (~ Pdata_in_3_)  &  (~ n1) ) ;
 assign n1436 = ( (~ Pinreg_3_)  &  (~ Pdata_46_) ) | ( (~ Pdata_46_)  &  n1 ) | ( (~ Pinreg_3_)  &  (~ n1) ) ;
 assign n1437 = ( (~ Pinreg_11_)  &  (~ Pdata_45_) ) | ( (~ Pdata_45_)  &  n1 ) | ( (~ Pinreg_11_)  &  (~ n1) ) ;
 assign n1438 = ( (~ Pinreg_19_)  &  (~ Pdata_44_) ) | ( (~ Pdata_44_)  &  n1 ) | ( (~ Pinreg_19_)  &  (~ n1) ) ;
 assign n1439 = ( (~ Pinreg_27_)  &  (~ Pdata_43_) ) | ( (~ Pdata_43_)  &  n1 ) | ( (~ Pinreg_27_)  &  (~ n1) ) ;
 assign n1440 = ( (~ Pinreg_35_)  &  (~ Pdata_42_) ) | ( (~ Pdata_42_)  &  n1 ) | ( (~ Pinreg_35_)  &  (~ n1) ) ;
 assign n1441 = ( (~ Pinreg_43_)  &  (~ Pdata_41_) ) | ( (~ Pdata_41_)  &  n1 ) | ( (~ Pinreg_43_)  &  (~ n1) ) ;
 assign n1442 = ( (~ Pinreg_51_)  &  (~ Pdata_40_) ) | ( (~ Pdata_40_)  &  n1 ) | ( (~ Pinreg_51_)  &  (~ n1) ) ;
 assign n1443 = ( (~ Pdata_in_1_)  &  (~ Pdata_39_) ) | ( (~ Pdata_39_)  &  n1 ) | ( (~ Pdata_in_1_)  &  (~ n1) ) ;
 assign n1444 = ( (~ Pinreg_1_)  &  (~ Pdata_38_) ) | ( (~ Pdata_38_)  &  n1 ) | ( (~ Pinreg_1_)  &  (~ n1) ) ;
 assign n1445 = ( (~ Pinreg_9_)  &  (~ Pdata_37_) ) | ( (~ Pdata_37_)  &  n1 ) | ( (~ Pinreg_9_)  &  (~ n1) ) ;
 assign n1446 = ( (~ Pinreg_17_)  &  (~ Pdata_36_) ) | ( (~ Pdata_36_)  &  n1 ) | ( (~ Pinreg_17_)  &  (~ n1) ) ;
 assign n1447 = ( (~ Pinreg_25_)  &  (~ Pdata_35_) ) | ( (~ Pdata_35_)  &  n1 ) | ( (~ Pinreg_25_)  &  (~ n1) ) ;
 assign n1448 = ( (~ Pinreg_33_)  &  (~ Pdata_34_) ) | ( (~ Pdata_34_)  &  n1 ) | ( (~ Pinreg_33_)  &  (~ n1) ) ;
 assign n1449 = ( (~ Pinreg_41_)  &  (~ Pdata_33_) ) | ( (~ Pdata_33_)  &  n1 ) | ( (~ Pinreg_41_)  &  (~ n1) ) ;
 assign n1450 = ( (~ Pinreg_49_)  &  (~ Pdata_32_) ) | ( (~ Pdata_32_)  &  n1 ) | ( (~ Pinreg_49_)  &  (~ n1) ) ;
 assign n1451 = ( (~ Pcount_2_)  &  n1664 ) | ( n923  &  n1664 ) ;
 assign n1452 = ( (~ Pcount_1_)  &  n1665 ) | ( n925  &  n1665 ) ;
 assign n1453 = ( (~ Pcount_1_)  &  (~ n1666) ) | ( Pcount_3_  &  Pcount_2_  &  (~ n1666) ) ;
 assign n1454 = ( (~ Pencrypt_mode_0_)  &  (~ Pencrypt_0_) ) | ( (~ Pencrypt_mode_0_)  &  n1 ) | ( (~ Pencrypt_0_)  &  (~ n1) ) ;
 assign n1457 = ( n201 ) | ( (~ n209) ) | ( (~ n207) ) | ( n914 ) ;
 assign n1458 = ( n220  &  (~ n911) ) | ( n795  &  (~ n911) ) | ( n220  &  n1189 ) | ( n795  &  n1189 ) ;
 assign n1459 = ( (~ n561)  &  (~ n1184) ) | ( (~ n914)  &  (~ n1184) ) | ( (~ n561)  &  n1188 ) | ( (~ n914)  &  n1188 ) ;
 assign n1464 = ( n261 ) | ( n266 ) | ( (~ n269) ) | ( n835 ) ;
 assign n1465 = ( n357 ) | ( (~ n588) ) | ( (~ n591) ) ;
 assign n1466 = ( (~ n355) ) | ( (~ n588) ) | ( n1217 ) ;
 assign n1468 = ( n585  &  n340 ) | ( n1220  &  n340 ) | ( n585  &  n357 ) | ( n1220  &  n357 ) ;
 assign n1470 = ( n1158 ) | ( n355 ) | ( n337 ) ;
 assign n1469 = ( (~ n326)  &  n1470 ) | ( n357  &  n1470 ) | ( n420  &  n1470 ) ;
 assign n1471 = ( (~ n357) ) | ( (~ n588) ) | ( (~ n591) ) ;
 assign n1472 = ( (~ Pdata_25_)  &  n1675 ) | ( Pdata_25_  &  (~ n1675) ) ;
 assign n1473 = ( n392 ) | ( (~ n432) ) | ( (~ n445) ) ;
 assign n1475 = ( (~ n432) ) | ( (~ n447) ) | ( (~ n445) ) ;
 assign n1474 = ( n1475  &  n401 ) | ( n1475  &  n375 ) | ( n1475  &  n452 ) ;
 assign n1476 = ( n369 ) | ( (~ n444) ) | ( n570 ) ;
 assign n1477 = ( (~ n407)  &  Pdata_17_ ) | ( n407  &  (~ Pdata_17_) ) ;
 assign n1478 = ( (~ n422)  &  Pdata_9_ ) | ( n422  &  (~ Pdata_9_) ) ;
 assign n1479 = ( (~ Pdata_1_)  &  n1678 ) | ( Pdata_1_  &  (~ n1678) ) ;
 assign n1480 = ( (~ n475) ) | ( n476 ) ;
 assign n1482 = ( (~ n459) ) | ( n1257 ) ;
 assign n1483 = ( (~ n496)  &  Pdata_26_ ) | ( n496  &  (~ Pdata_26_) ) ;
 assign n1486 = ( n526 ) | ( (~ n647) ) | ( n654 ) ;
 assign n1484 = ( n511 ) | ( (~ n546) ) ;
 assign n1487 = ( n525 ) | ( n522 ) ;
 assign n1488 = ( n542 ) | ( (~ n549) ) | ( (~ n647) ) ;
 assign n1489 = ( n522  &  (~ n1163) ) | ( n658  &  (~ n1163) ) | ( n522  &  n1274 ) | ( n658  &  n1274 ) ;
 assign n1490 = ( n529  &  (~ n1265) ) | ( (~ n549)  &  (~ n1265) ) | ( n529  &  n1275 ) | ( (~ n549)  &  n1275 ) ;
 assign n1493 = ( n648 ) | ( n1163 ) | ( (~ n1165) ) ;
 assign n1492 = ( n517  &  n1493 ) | ( (~ n513)  &  n526  &  n1493 ) ;
 assign n1494 = ( (~ n533)  &  Pdata_18_ ) | ( n533  &  (~ Pdata_18_) ) ;
 assign n1495 = ( n648 ) | ( n647 ) | ( n1275 ) ;
 assign n1497 = ( n529 ) | ( n510 ) | ( n654 ) ;
 assign n1496 = ( n1497  &  n508 ) | ( n1497  &  n1275 ) ;
 assign n1499 = ( n655  &  n658 ) | ( n658  &  n1163 ) | ( n655  &  (~ n1272) ) | ( n1163  &  (~ n1272) ) ;
 assign n1500 = ( (~ Pdata_10_)  &  n1680 ) | ( Pdata_10_  &  (~ n1680) ) ;
 assign n1502 = ( n392  &  (~ n432) ) | ( (~ n432)  &  n434 ) | ( n392  &  n449 ) | ( n434  &  n449 ) ;
 assign n1503 = ( (~ n575)  &  Pdata_27_ ) | ( n575  &  (~ Pdata_27_) ) ;
 assign n1504 = ( (~ Pdata_19_)  &  n1684 ) | ( Pdata_19_  &  (~ n1684) ) ;
 assign n1505 = ( (~ n633)  &  Pdata_11_ ) | ( n633  &  (~ Pdata_11_) ) ;
 assign n1506 = ( n525  &  n646 ) | ( n646  &  (~ n1272) ) | ( n525  &  n1275 ) | ( (~ n1272)  &  n1275 ) ;
 assign n1507 = ( (~ Pdata_3_)  &  n1688 ) | ( Pdata_3_  &  (~ n1688) ) ;
 assign n1508 = ( (~ n510) ) | ( (~ n549) ) | ( n1270 ) ;
 assign n1509 = ( n510 ) | ( (~ n515) ) | ( (~ n546) ) ;
 assign n1510 = ( (~ n661)  &  Pdata_28_ ) | ( n661  &  (~ Pdata_28_) ) ;
 assign n1511 = ( (~ n680)  &  Pdata_20_ ) | ( n680  &  (~ Pdata_20_) ) ;
 assign n1512 = ( (~ n693)  &  Pdata_12_ ) | ( n693  &  (~ Pdata_12_) ) ;
 assign n1514 = ( n469  &  (~ n475) ) | ( n469  &  n1248 ) | ( n475  &  n1248 ) ;
 assign n1515 = ( (~ n701)  &  Pdata_4_ ) | ( n701  &  (~ Pdata_4_) ) ;
 assign n1516 = ( (~ n742)  &  n755 ) | ( n752  &  n755 ) | ( (~ n742)  &  n1318 ) | ( n752  &  n1318 ) ;
 assign n1517 = ( (~ Pdata_29_)  &  n1690 ) | ( Pdata_29_  &  (~ n1690) ) ;
 assign n1520 = ( (~ n772) ) | ( (~ n777) ) | ( n1300 ) ;
 assign n1518 = ( n775  &  n1520 ) | ( (~ n1323)  &  n1520 ) ;
 assign n1521 = ( (~ Pdata_21_)  &  n1692 ) | ( Pdata_21_  &  (~ n1692) ) ;
 assign n1522 = ( (~ n228)  &  n914 ) | ( n786  &  n914 ) | ( (~ n228)  &  (~ n1187) ) | ( n786  &  (~ n1187) ) ;
 assign n1524 = ( (~ Pdata_13_)  &  n1695 ) | ( Pdata_13_  &  (~ n1695) ) ;
 assign n1525 = ( n729  &  n738 ) | ( n730  &  n738 ) | ( n729  &  n724 ) | ( n730  &  n724 ) ;
 assign n1528 = ( (~ n826)  &  Pdata_30_ ) | ( n826  &  (~ Pdata_30_) ) ;
 assign n1529 = ( (~ n836)  &  Pdata_22_ ) | ( n836  &  (~ Pdata_22_) ) ;
 assign n1530 = ( (~ n460)  &  n1248 ) | ( (~ n491)  &  n1248 ) | ( n846  &  n1248 ) ;
 assign n1532 = ( n470  &  n495 ) | ( n475  &  n495 ) | ( n470  &  (~ n675) ) | ( n475  &  (~ n675) ) ;
 assign n1533 = ( (~ Pdata_14_)  &  n1703 ) | ( Pdata_14_  &  (~ n1703) ) ;
 assign n1534 = ( (~ n629)  &  n1166 ) | ( n1166  &  n1298 ) | ( (~ n629)  &  n1324 ) | ( n1298  &  n1324 ) ;
 assign n1537 = ( (~ n766)  &  n872 ) | ( n872  &  n876 ) | ( (~ n766)  &  (~ n1167) ) | ( n876  &  (~ n1167) ) ;
 assign n1538 = ( (~ Pdata_31_)  &  n1709 ) | ( Pdata_31_  &  (~ n1709) ) ;
 assign n1539 = ( (~ Pdata_23_)  &  n1711 ) | ( Pdata_23_  &  (~ n1711) ) ;
 assign n1540 = ( (~ n900)  &  Pdata_15_ ) | ( n900  &  (~ Pdata_15_) ) ;
 assign n1541 = ( (~ Pdata_7_)  &  n1714 ) | ( Pdata_7_  &  (~ n1714) ) ;
 assign n1542 = ( (~ Pinreg_48_)  &  (~ Pinreg_27_) ) | ( (~ Pinreg_48_)  &  n1356 ) | ( (~ Pinreg_27_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1543 = ( (~ Pinreg_35_)  &  (~ Pinreg_27_) ) | ( (~ Pinreg_27_)  &  n1356 ) | ( (~ Pinreg_35_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1544 = ( (~ Pinreg_43_)  &  (~ Pinreg_35_) ) | ( (~ Pinreg_35_)  &  n1356 ) | ( (~ Pinreg_43_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1545 = ( (~ Pinreg_51_)  &  (~ Pinreg_43_) ) | ( (~ Pinreg_43_)  &  n1356 ) | ( (~ Pinreg_51_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1546 = ( (~ Pinreg_51_)  &  (~ Pdata_in_2_) ) | ( (~ Pinreg_51_)  &  n1356 ) | ( (~ Pdata_in_2_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1547 = ( (~ Pinreg_2_)  &  (~ Pdata_in_2_) ) | ( (~ Pdata_in_2_)  &  n1356 ) | ( (~ Pinreg_2_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1548 = ( (~ Pinreg_10_)  &  (~ Pinreg_2_) ) | ( (~ Pinreg_2_)  &  n1356 ) | ( (~ Pinreg_10_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1549 = ( (~ Pinreg_18_)  &  (~ Pinreg_10_) ) | ( (~ Pinreg_10_)  &  n1356 ) | ( (~ Pinreg_18_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1550 = ( (~ Pinreg_26_)  &  (~ Pinreg_18_) ) | ( (~ Pinreg_18_)  &  n1356 ) | ( (~ Pinreg_26_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1551 = ( (~ Pinreg_34_)  &  (~ Pinreg_26_) ) | ( (~ Pinreg_26_)  &  n1356 ) | ( (~ Pinreg_34_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1552 = ( (~ Pinreg_42_)  &  (~ Pinreg_34_) ) | ( (~ Pinreg_34_)  &  n1356 ) | ( (~ Pinreg_42_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1553 = ( (~ Pinreg_50_)  &  (~ Pinreg_42_) ) | ( (~ Pinreg_42_)  &  n1356 ) | ( (~ Pinreg_50_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1554 = ( (~ Pinreg_50_)  &  (~ Pdata_in_1_) ) | ( (~ Pinreg_50_)  &  n1356 ) | ( (~ Pdata_in_1_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1555 = ( (~ Pinreg_1_)  &  (~ Pdata_in_1_) ) | ( (~ Pdata_in_1_)  &  n1356 ) | ( (~ Pinreg_1_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1556 = ( (~ Pinreg_9_)  &  (~ Pinreg_1_) ) | ( (~ Pinreg_1_)  &  n1356 ) | ( (~ Pinreg_9_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1557 = ( (~ Pinreg_17_)  &  (~ Pinreg_9_) ) | ( (~ Pinreg_9_)  &  n1356 ) | ( (~ Pinreg_17_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1558 = ( (~ Pinreg_25_)  &  (~ Pinreg_17_) ) | ( (~ Pinreg_17_)  &  n1356 ) | ( (~ Pinreg_25_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1559 = ( (~ Pinreg_33_)  &  (~ Pinreg_25_) ) | ( (~ Pinreg_25_)  &  n1356 ) | ( (~ Pinreg_33_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1560 = ( (~ Pinreg_41_)  &  (~ Pinreg_33_) ) | ( (~ Pinreg_33_)  &  n1356 ) | ( (~ Pinreg_41_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1561 = ( (~ Pinreg_49_)  &  (~ Pinreg_41_) ) | ( (~ Pinreg_41_)  &  n1356 ) | ( (~ Pinreg_49_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1562 = ( (~ Pinreg_49_)  &  (~ Pdata_in_0_) ) | ( (~ Pinreg_49_)  &  n1356 ) | ( (~ Pdata_in_0_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1563 = ( (~ Pinreg_0_)  &  (~ Pdata_in_0_) ) | ( (~ Pdata_in_0_)  &  n1356 ) | ( (~ Pinreg_0_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1564 = ( (~ Pinreg_8_)  &  (~ Pinreg_0_) ) | ( (~ Pinreg_0_)  &  n1356 ) | ( (~ Pinreg_8_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1565 = ( (~ Pinreg_16_)  &  (~ Pinreg_8_) ) | ( (~ Pinreg_8_)  &  n1356 ) | ( (~ Pinreg_16_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1566 = ( (~ Pinreg_24_)  &  (~ Pinreg_16_) ) | ( (~ Pinreg_16_)  &  n1356 ) | ( (~ Pinreg_24_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1567 = ( (~ Pinreg_32_)  &  (~ Pinreg_24_) ) | ( (~ Pinreg_24_)  &  n1356 ) | ( (~ Pinreg_32_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1568 = ( (~ Pinreg_40_)  &  (~ Pinreg_32_) ) | ( (~ Pinreg_32_)  &  n1356 ) | ( (~ Pinreg_40_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1569 = ( (~ Pinreg_48_)  &  (~ Pinreg_40_) ) | ( (~ Pinreg_40_)  &  n1356 ) | ( (~ Pinreg_48_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1570 = ( (~ Pinreg_54_)  &  (~ Pdata_in_3_) ) | ( (~ Pinreg_54_)  &  n1356 ) | ( (~ Pdata_in_3_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1571 = ( (~ Pinreg_3_)  &  (~ Pdata_in_3_) ) | ( (~ Pdata_in_3_)  &  n1356 ) | ( (~ Pinreg_3_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1572 = ( (~ Pinreg_11_)  &  (~ Pinreg_3_) ) | ( (~ Pinreg_3_)  &  n1356 ) | ( (~ Pinreg_11_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1573 = ( (~ Pinreg_19_)  &  (~ Pinreg_11_) ) | ( (~ Pinreg_11_)  &  n1356 ) | ( (~ Pinreg_19_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1574 = ( (~ Pinreg_19_)  &  (~ Pdata_in_4_) ) | ( (~ Pinreg_19_)  &  n1356 ) | ( (~ Pdata_in_4_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1575 = ( (~ Pinreg_4_)  &  (~ Pdata_in_4_) ) | ( (~ Pdata_in_4_)  &  n1356 ) | ( (~ Pinreg_4_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1576 = ( (~ Pinreg_12_)  &  (~ Pinreg_4_) ) | ( (~ Pinreg_4_)  &  n1356 ) | ( (~ Pinreg_12_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1577 = ( (~ Pinreg_20_)  &  (~ Pinreg_12_) ) | ( (~ Pinreg_12_)  &  n1356 ) | ( (~ Pinreg_20_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1578 = ( (~ Pinreg_28_)  &  (~ Pinreg_20_) ) | ( (~ Pinreg_20_)  &  n1356 ) | ( (~ Pinreg_28_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1579 = ( (~ Pinreg_36_)  &  (~ Pinreg_28_) ) | ( (~ Pinreg_28_)  &  n1356 ) | ( (~ Pinreg_36_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1580 = ( (~ Pinreg_44_)  &  (~ Pinreg_36_) ) | ( (~ Pinreg_36_)  &  n1356 ) | ( (~ Pinreg_44_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1581 = ( (~ Pinreg_52_)  &  (~ Pinreg_44_) ) | ( (~ Pinreg_44_)  &  n1356 ) | ( (~ Pinreg_52_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1582 = ( (~ Pinreg_52_)  &  (~ Pdata_in_5_) ) | ( (~ Pinreg_52_)  &  n1356 ) | ( (~ Pdata_in_5_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1583 = ( (~ Pinreg_5_)  &  (~ Pdata_in_5_) ) | ( (~ Pdata_in_5_)  &  n1356 ) | ( (~ Pinreg_5_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1584 = ( (~ Pinreg_13_)  &  (~ Pinreg_5_) ) | ( (~ Pinreg_5_)  &  n1356 ) | ( (~ Pinreg_13_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1585 = ( (~ Pinreg_21_)  &  (~ Pinreg_13_) ) | ( (~ Pinreg_13_)  &  n1356 ) | ( (~ Pinreg_21_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1586 = ( (~ Pinreg_29_)  &  (~ Pinreg_21_) ) | ( (~ Pinreg_21_)  &  n1356 ) | ( (~ Pinreg_29_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1587 = ( (~ Pinreg_37_)  &  (~ Pinreg_29_) ) | ( (~ Pinreg_29_)  &  n1356 ) | ( (~ Pinreg_37_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1588 = ( (~ Pinreg_45_)  &  (~ Pinreg_37_) ) | ( (~ Pinreg_37_)  &  n1356 ) | ( (~ Pinreg_45_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1589 = ( (~ Pinreg_53_)  &  (~ Pinreg_45_) ) | ( (~ Pinreg_45_)  &  n1356 ) | ( (~ Pinreg_53_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1590 = ( (~ Pinreg_53_)  &  (~ Pdata_in_6_) ) | ( (~ Pinreg_53_)  &  n1356 ) | ( (~ Pdata_in_6_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1591 = ( (~ Pinreg_6_)  &  (~ Pdata_in_6_) ) | ( (~ Pdata_in_6_)  &  n1356 ) | ( (~ Pinreg_6_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1592 = ( (~ Pinreg_14_)  &  (~ Pinreg_6_) ) | ( (~ Pinreg_6_)  &  n1356 ) | ( (~ Pinreg_14_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1593 = ( (~ Pinreg_22_)  &  (~ Pinreg_14_) ) | ( (~ Pinreg_14_)  &  n1356 ) | ( (~ Pinreg_22_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1594 = ( (~ Pinreg_30_)  &  (~ Pinreg_22_) ) | ( (~ Pinreg_22_)  &  n1356 ) | ( (~ Pinreg_30_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1595 = ( (~ Pinreg_38_)  &  (~ Pinreg_30_) ) | ( (~ Pinreg_30_)  &  n1356 ) | ( (~ Pinreg_38_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1596 = ( (~ Pinreg_46_)  &  (~ Pinreg_38_) ) | ( (~ Pinreg_38_)  &  n1356 ) | ( (~ Pinreg_46_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1597 = ( (~ Pinreg_54_)  &  (~ Pinreg_46_) ) | ( (~ Pinreg_46_)  &  n1356 ) | ( (~ Pinreg_54_)  &  n1357 ) | ( n1356  &  n1357 ) ;
 assign n1598 = ( n264 ) | ( n269 ) | ( (~ n292) ) ;
 assign n1599 = ( n270  &  (~ n835) ) | ( n273  &  (~ n835) ) | ( (~ n835)  &  (~ n1369) ) ;
 assign n1600 = ( (~ n243)  &  (~ n254) ) | ( (~ n254)  &  n262 ) | ( (~ n254)  &  n269 ) ;
 assign n1602 = ( (~ n254)  &  (~ n274) ) | ( (~ n254)  &  n835 ) ;
 assign n1604 = ( (~ n1158)  &  (~ n1375) ) | ( (~ n317)  &  (~ n355)  &  (~ n1158) ) ;
 assign n1605 = ( (~ n317)  &  n326  &  n1158 ) | ( n326  &  n1158  &  (~ n1218) ) ;
 assign n1607 = ( (~ n458)  &  n477 ) | ( n477  &  n851  &  n1250 ) ;
 assign n1609 = ( (~ n460) ) | ( (~ n477) ) | ( (~ n851) ) | ( (~ n1252) ) ;
 assign n1610 = ( n508 ) | ( n1275 ) | ( n647 ) ;
 assign n1611 = ( n512  &  (~ n647) ) | ( (~ n526)  &  n549  &  (~ n647) ) ;
 assign n1614 = ( n647  &  (~ n1496) ) | ( n647  &  (~ n1163)  &  n1272 ) ;
 assign n1615 = ( n545  &  (~ n647) ) | ( (~ n647)  &  n1165  &  n1265 ) ;
 assign n1616 = ( n230  &  n789 ) | ( n230  &  n1155 ) | ( n789  &  (~ n1155) ) ;
 assign n1617 = ( n914  &  n1187 ) | ( n914  &  n228  &  n220 ) ;
 assign n1619 = ( n201  &  (~ n1378) ) | ( n201  &  n227  &  n231 ) ;
 assign n1620 = ( (~ n201)  &  (~ n915)  &  n1616 ) ;
 assign n1622 = ( n583 ) | ( (~ n1218) ) ;
 assign n1621 = ( n587  &  (~ n1158) ) | ( n326  &  (~ n1158)  &  n1622 ) ;
 assign n1623 = ( n344 ) | ( n357 ) | ( (~ n1158) ) ;
 assign n1624 = ( (~ n604) ) | ( (~ n1300) ) | ( n1325 ) ;
 assign n1625 = ( n647 ) | ( (~ n1265) ) | ( n1303 ) ;
 assign n1626 = ( (~ n1163)  &  (~ n1382) ) | ( (~ n1163)  &  n1164  &  n1272 ) ;
 assign n1627 = ( n508 ) | ( (~ n647) ) | ( (~ n1163) ) | ( (~ n1303) ) ;
 assign n1628 = ( (~ n477) ) | ( n847 ) | ( (~ n849) ) ;
 assign n1629 = ( n375  &  (~ n432) ) ;
 assign n1630 = ( (~ n375)  &  n403 ) | ( (~ n375)  &  n438 ) ;
 assign n1631 = ( (~ n570) ) | ( (~ n572) ) | ( n1629 ) | ( n1630 ) ;
 assign n1633 = ( n851  &  n849 ) ;
 assign n1632 = ( (~ n477)  &  n1633 ) | ( (~ n477)  &  n852  &  n1252 ) ;
 assign n1635 = ( (~ n722) ) | ( (~ n751) ) | ( (~ n802) ) | ( (~ n895) ) ;
 assign n1636 = ( n779  &  (~ n1325) ) | ( n777  &  n862  &  (~ n1325) ) ;
 assign n1638 = ( (~ n862) ) | ( (~ n1167) ) | ( (~ n1325) ) ;
 assign n1639 = ( (~ n766)  &  n774  &  (~ n1166) ) | ( (~ n766)  &  (~ n1166)  &  n1295 ) ;
 assign n1640 = ( (~ n1166) ) | ( n1324 ) ;
 assign n1641 = ( n201  &  (~ n1522) ) | ( n201  &  n227  &  n1186 ) ;
 assign n1642 = ( (~ n201)  &  n561 ) | ( (~ n201)  &  n788 ) | ( (~ n201)  &  n790 ) ;
 assign n1643 = ( n751  &  (~ n1525) ) | ( n751  &  n814  &  (~ n1318) ) ;
 assign n1645 = ( (~ n751)  &  (~ n1668) ) | ( (~ n751)  &  n802  &  (~ n1318) ) ;
 assign n1647 = ( n266  &  n263 ) ;
 assign n1648 = ( (~ n261)  &  (~ n266) ) | ( (~ n266)  &  n269 ) ;
 assign n1649 = ( (~ n835)  &  n1201 ) | ( n274  &  n281  &  (~ n835) ) ;
 assign n1651 = ( n477  &  (~ n1530) ) | ( (~ n472)  &  n477  &  n1246 ) ;
 assign n1653 = ( (~ n477)  &  (~ n493) ) | ( (~ n477)  &  n848 ) | ( (~ n477)  &  n850 ) ;
 assign n1654 = ( (~ n629) ) | ( n775 ) | ( n776 ) ;
 assign n1655 = ( n729 ) | ( n742 ) | ( n749 ) | ( (~ n756) ) ;
 assign n1656 = ( n742  &  n887  &  n1340 ) | ( n742  &  (~ n898)  &  n1340 ) ;
 assign n1657 = ( (~ n738) ) | ( n740 ) ;
 assign n1658 = ( (~ n738)  &  n817 ) | ( (~ n738)  &  n803  &  n814 ) ;
 assign n1659 = ( (~ n201)  &  n1184 ) | ( n201  &  n1185 ) | ( n1184  &  n1185 ) ;
 assign n1660 = ( n207  &  (~ n1155) ) | ( n207  &  n1659 ) | ( n1155  &  n1659 ) ;
 assign n1663 = ( n201  &  (~ n1385) ) | ( (~ n201)  &  (~ n1386) ) | ( (~ n1385)  &  (~ n1386) ) ;
 assign n1664 = ( Pcount_2_ ) | ( (~ Pcount_1_) ) | ( (~ Pcount_0_) ) | ( n924 ) ;
 assign n1665 = ( Pcount_1_ ) | ( (~ Pcount_0_) ) | ( n924 ) ;
 assign n1666 = ( Pcount_3_  &  (~ Pcount_1_) ) | ( Pcount_2_  &  (~ Pcount_1_) ) ;
 assign n1668 = ( (~ n722) ) | ( n724 ) ;
 assign n1669 = ( n202  &  n210  &  n215  &  n223  &  (~ n225)  &  (~ n229)  &  n1458  &  n1459 ) ;
 assign n1672 = ( n331  &  n424  &  n1468  &  (~ n1604)  &  (~ n1605) ) ;
 assign n1675 = ( n331  &  n333  &  n350  &  (~ n353)  &  n358  &  (~ n360)  &  n421  &  n1220 ) ;
 assign n1678 = ( n386  &  n400  &  n433  &  n437  &  n439  &  (~ n443)  &  n448  &  n451 ) ;
 assign n1680 = ( n516  &  n521  &  n541  &  n1499  &  (~ n1614)  &  (~ n1615) ) ;
 assign n1683 = ( (~ n202) ) | ( n208 ) | ( (~ n210) ) | ( (~ n554) ) | ( n558 ) | ( n560 ) | ( n1619 ) | ( n1620 ) ;
 assign n1684 = ( n331  &  n336  &  n350  &  (~ n590)  &  n593  &  n1221  &  (~ n1621)  &  n1623 ) ;
 assign n1688 = ( n519  &  n534  &  n541  &  n1506  &  (~ n1626)  &  n1627 ) ;
 assign n1690 = ( n741  &  (~ n757)  &  n760  &  n1321  &  n1341  &  n1516 ) ;
 assign n1692 = ( n599  &  n618  &  n1326  &  n1518  &  (~ n1636)  &  n1638  &  (~ n1639)  &  n1640 ) ;
 assign n1695 = ( n199  &  n210  &  n794  &  n1329  &  (~ n1641)  &  (~ n1642) ) ;
 assign n1698 = ( (~ n714) ) | ( (~ n809) ) | ( (~ n810) ) | ( n813 ) | ( n816 ) | ( (~ n901) ) | ( n1643 ) | ( n1645 ) ;
 assign n1702 = ( n262  &  (~ n264)  &  (~ n269)  &  n1172 ) ;
 assign n1703 = ( n466  &  n668  &  n1254  &  n1532  &  (~ n1651)  &  (~ n1653) ) ;
 assign n1706 = ( (~ n635) ) | ( n858 ) | ( n859 ) | ( n860 ) | ( n864 ) | ( n1323 ) | ( (~ n1326) ) | ( (~ n1534) ) ;
 assign n1709 = ( n608  &  n618  &  n879  &  (~ n880)  &  n1326  &  n1537 ) ;
 assign n1711 = ( n804  &  n889  &  n1321  &  n1655  &  (~ n1656)  &  n1657  &  (~ n1658)  &  n1668 ) ;
 assign n1714 = ( n202  &  (~ n910)  &  n913  &  n917  &  n1329  &  n1663 ) ;
 assign n1717 = ( (~ Pdata_2_)  &  n1683 ) | ( Pdata_2_  &  (~ n1683) ) ;
 assign n1718 = ( (~ Pdata_5_)  &  n1698 ) | ( Pdata_5_  &  (~ n1698) ) ;
 assign n1719 = ( (~ Pdata_6_)  &  n1706 ) | ( Pdata_6_  &  (~ n1706) ) ;


endmodule

