module s38584 (
	Pg6753, Pg6752, Pg6751, Pg6750, Pg6749, Pg6748, Pg6747, Pg6746, 
	Pg6745, Pg6744, Pg135, Pg134, Pg127, Pg126, Pg125, Pg124, Pg120, Pg116, 
	Pg115, Pg114, Pg113, Pg100, Pg99, Pg92, Pg91, Pg90, Pg84, Pg73, 
	Pg72, Pg64, Pg57, Pg56, Pg54, Pg53, Pg44, Pg36, Pg35, Pg5, 
	PCLK, Pg34972, Pg34956, Pg34927, Pg34925, Pg34923, Pg34921, Pg34919, Pg34917, Pg34915, 
	Pg34913, Pg34839, Pg34788, Pg34597, Pg34437, Pg34436, Pg34435, Pg34425, Pg34383, Pg34240, 
	Pg34239, Pg34238, Pg34237, Pg34236, Pg34235, Pg34234, Pg34233, Pg34232, Pg34221, Pg34201, 
	Pg33959, Pg33950, Pg33949, Pg33948, Pg33947, Pg33946, Pg33945, Pg33935, Pg33894, Pg33874, 
	Pg33659, Pg33636, Pg33533, Pg33435, Pg33079, Pg32975, Pg32454, Pg32429, Pg32185, Pg31863, 
	Pg31862, Pg31861, Pg31860, Pg31793, Pg31665, Pg31656, Pg31521, Pg30332, Pg30331, Pg30330, 
	Pg30329, Pg30327, Pg29221, Pg29220, Pg29219, Pg29218, Pg29217, Pg29216, Pg29215, Pg29214, 
	Pg29213, Pg29212, Pg29211, Pg29210, Pg28753, Pg28042, Pg28041, Pg28030, Pg27831, Pg26877, 
	Pg26876, Pg26875, Pg26801, Pg25590, Pg25589, Pg25588, Pg25587, Pg25586, Pg25585, Pg25584, 
	Pg25583, Pg25582, Pg25259, Pg25219, Pg25167, Pg25114, Pg24185, Pg24184, Pg24183, Pg24182, 
	Pg24181, Pg24180, Pg24179, Pg24178, Pg24177, Pg24176, Pg24175, Pg24174, Pg24173, Pg24172, 
	Pg24171, Pg24170, Pg24169, Pg24168, Pg24167, Pg24166, Pg24165, Pg24164, Pg24163, Pg24162, 
	Pg24161, Pg24151, Pg23759, Pg23683, Pg23652, Pg23612, Pg23190, Pg23002, Pg21727, Pg21698, 
	Pg21292, Pg21270, Pg21245, Pg21176, Pg20901, Pg20899, Pg20763, Pg20654, Pg20652, Pg20557, 
	Pg20049, Pg19357, Pg19334, Pg18881, Pg18101, Pg18100, Pg18099, Pg18098, Pg18097, Pg18096, 
	Pg18095, Pg18094, Pg18092, Pg17871, Pg17845, Pg17819, Pg17813, Pg17787, Pg17778, Pg17764, 
	Pg17760, Pg17743, Pg17739, Pg17722, Pg17715, Pg17711, Pg17688, Pg17685, Pg17678, Pg17674, 
	Pg17649, Pg17646, Pg17639, Pg17607, Pg17604, Pg17580, Pg17577, Pg17519, Pg17423, Pg17404, 
	Pg17400, Pg17320, Pg17316, Pg17291, Pg16955, Pg16924, Pg16874, Pg16775, Pg16748, Pg16744, 
	Pg16722, Pg16718, Pg16693, Pg16686, Pg16659, Pg16656, Pg16627, Pg16624, Pg16603, Pg14828, 
	Pg14779, Pg14749, Pg14738, Pg14705, Pg14694, Pg14673, Pg14662, Pg14635, Pg14597, Pg14518, 
	Pg14451, Pg14421, Pg14217, Pg14201, Pg14189, Pg14167, Pg14147, Pg14125, Pg14096, Pg13966, 
	Pg13926, Pg13906, Pg13895, Pg13881, Pg13865, Pg13272, Pg13259, Pg13099, Pg13085, Pg13068, 
	Pg13049, Pg13039, Pg12923, Pg12919, Pg12833, Pg12832, Pg12470, Pg12422, Pg12368, Pg12350, 
	Pg12300, Pg12238, Pg12184, Pg11770, Pg11678, Pg11447, Pg11418, Pg11388, Pg11349, Pg10527, 
	Pg10500, Pg10306, Pg10122, Pg9817, Pg9743, Pg9741, Pg9682, Pg9680, Pg9617, Pg9615, 
	Pg9555, Pg9553, Pg9497, Pg9251, Pg9048, Pg9019, Pg8920, Pg8919, Pg8918, Pg8917, 
	Pg8916, Pg8915, Pg8870, Pg8839, Pg8789, Pg8788, Pg8787, Pg8786, Pg8785, Pg8784, 
	Pg8783, Pg8719, Pg8475, Pg8416, Pg8403, Pg8398, Pg8358, Pg8353, Pg8344, Pg8342, 
	Pg8291, Pg8283, Pg8279, Pg8277, Pg8235, Pg8215, Pg8178, Pg8132, Pg7946, Pg7916, 
	Pg7540, Pg7260, Pg7257, Pg7245, Pg7243);

input Pg6753, Pg6752, Pg6751, Pg6750, Pg6749, Pg6748, Pg6747, Pg6746, Pg6745, Pg6744, Pg135, Pg134, Pg127, Pg126, Pg125, Pg124, Pg120, Pg116, Pg115, Pg114, Pg113, Pg100, Pg99, Pg92, Pg91, Pg90, Pg84, Pg73, Pg72, Pg64, Pg57, Pg56, Pg54, Pg53, Pg44, Pg36, Pg35, Pg5, PCLK;

output Pg34972, Pg34956, Pg34927, Pg34925, Pg34923, Pg34921, Pg34919, Pg34917, Pg34915, Pg34913, Pg34839, Pg34788, Pg34597, Pg34437, Pg34436, Pg34435, Pg34425, Pg34383, Pg34240, Pg34239, Pg34238, Pg34237, Pg34236, Pg34235, Pg34234, Pg34233, Pg34232, Pg34221, Pg34201, Pg33959, Pg33950, Pg33949, Pg33948, Pg33947, Pg33946, Pg33945, Pg33935, Pg33894, Pg33874, Pg33659, Pg33636, Pg33533, Pg33435, Pg33079, Pg32975, Pg32454, Pg32429, Pg32185, Pg31863, Pg31862, Pg31861, Pg31860, Pg31793, Pg31665, Pg31656, Pg31521, Pg30332, Pg30331, Pg30330, Pg30329, Pg30327, Pg29221, Pg29220, Pg29219, Pg29218, Pg29217, Pg29216, Pg29215, Pg29214, Pg29213, Pg29212, Pg29211, Pg29210, Pg28753, Pg28042, Pg28041, Pg28030, Pg27831, Pg26877, Pg26876, Pg26875, Pg26801, Pg25590, Pg25589, Pg25588, Pg25587, Pg25586, Pg25585, Pg25584, Pg25583, Pg25582, Pg25259, Pg25219, Pg25167, Pg25114, Pg24185, Pg24184, Pg24183, Pg24182, Pg24181, Pg24180, Pg24179, Pg24178, Pg24177, Pg24176, Pg24175, Pg24174, Pg24173, Pg24172, Pg24171, Pg24170, Pg24169, Pg24168, Pg24167, Pg24166, Pg24165, Pg24164, Pg24163, Pg24162, Pg24161, Pg24151, Pg23759, Pg23683, Pg23652, Pg23612, Pg23190, Pg23002, Pg21727, Pg21698, Pg21292, Pg21270, Pg21245, Pg21176, Pg20901, Pg20899, Pg20763, Pg20654, Pg20652, Pg20557, Pg20049, Pg19357, Pg19334, Pg18881, Pg18101, Pg18100, Pg18099, Pg18098, Pg18097, Pg18096, Pg18095, Pg18094, Pg18092, Pg17871, Pg17845, Pg17819, Pg17813, Pg17787, Pg17778, Pg17764, Pg17760, Pg17743, Pg17739, Pg17722, Pg17715, Pg17711, Pg17688, Pg17685, Pg17678, Pg17674, Pg17649, Pg17646, Pg17639, Pg17607, Pg17604, Pg17580, Pg17577, Pg17519, Pg17423, Pg17404, Pg17400, Pg17320, Pg17316, Pg17291, Pg16955, Pg16924, Pg16874, Pg16775, Pg16748, Pg16744, Pg16722, Pg16718, Pg16693, Pg16686, Pg16659, Pg16656, Pg16627, Pg16624, Pg16603, Pg14828, Pg14779, Pg14749, Pg14738, Pg14705, Pg14694, Pg14673, Pg14662, Pg14635, Pg14597, Pg14518, Pg14451, Pg14421, Pg14217, Pg14201, Pg14189, Pg14167, Pg14147, Pg14125, Pg14096, Pg13966, Pg13926, Pg13906, Pg13895, Pg13881, Pg13865, Pg13272, Pg13259, Pg13099, Pg13085, Pg13068, Pg13049, Pg13039, Pg12923, Pg12919, Pg12833, Pg12832, Pg12470, Pg12422, Pg12368, Pg12350, Pg12300, Pg12238, Pg12184, Pg11770, Pg11678, Pg11447, Pg11418, Pg11388, Pg11349, Pg10527, Pg10500, Pg10306, Pg10122, Pg9817, Pg9743, Pg9741, Pg9682, Pg9680, Pg9617, Pg9615, Pg9555, Pg9553, Pg9497, Pg9251, Pg9048, Pg9019, Pg8920, Pg8919, Pg8918, Pg8917, Pg8916, Pg8915, Pg8870, Pg8839, Pg8789, Pg8788, Pg8787, Pg8786, Pg8785, Pg8784, Pg8783, Pg8719, Pg8475, Pg8416, Pg8403, Pg8398, Pg8358, Pg8353, Pg8344, Pg8342, Pg8291, Pg8283, Pg8279, Pg8277, Pg8235, Pg8215, Pg8178, Pg8132, Pg7946, Pg7916, Pg7540, Pg7260, Pg7257, Pg7245, Pg7243;

wire wire4366, wire4376, wire4378, wire4379, wire4394, wire4406, n160, n172, n173, n171, n175, n176, n174, n178, n179, n177, n180, n181, n182, n184, n185, n186, n188, Ng33046, n189, Ng34441, n190, Ng33982, n191, Ng34007, n192, Ng30405, n193, Ng30416, n194, Ng30466, n195, Ng34617, n196, Ng33974, n197, Ng30505, n198, Ng33554, n199, Ng30432, n200, Ng33064, n201, Ng34881, n202, Ng24232, n206, n204, Ng34733, n207, Ng33026, n208, Ng31867, n212, Ng24344, n213, Ng33966, n214, Ng33550, Ng30393, n217, Ng29248, n218, Ng24274, n219, Ng33973, n220, Ng30360, n221, Ng34460, n222, Ng30494, n223, Ng30384, n227, Ng24340, n228, Ng29223, n229, Ng34252, n230, Ng30489, n231, Ng29301, n232, Ng33022, n233, Ng30496, n234, Ng33043, n235, Ng29263, n236, Ng30533, n237, Ng34015, n238, Ng34031, n239, Ng34452, n240, Ng34646, n241, Ng34001, n242, Ng25633, n243, Ng24259, n244, Ng33049, n245, Ng34609, n246, Ng31869, n247, Ng30490, n248, Ng30427, n249, Ng21894, n250, Ng33965, n251, Ng34645, n252, Ng34267, n253, Ng34644, n254, Ng30534, n255, Ng33535, n256, Ng30498, n257, Ng25613, n258, Ng34438, n259, Ng30439, n260, Ng30541, n261, Ng30519, n262, Ng25621, n263, Ng34036, n264, Ng30476, n265, Ng30429, n266, Ng32997, n267, Ng33063, n268, Ng30424, n269, Ng32977, n270, Ng34026, n271, Ng30420, n272, Ng33560, n273, Ng29226, n274, Ng25619, n275, Ng34455, n276, Ng33625, n277, Ng34790, Ng30414, n280, Ng30390, n282, n281, Ng25594, Ng34034, n283, Ng33541, n284, Ng28093, n285, Ng30404, n286, Ng29303, n287, Ng26917, n288, Ng33624, n289, Ng34911, n290, Ng34627, n291, Ng33013, n292, Ng32981, n293, Ng30483, n294, Ng32994, n295, Ng28070, n296, Ng30453, n297, Ng33539, n298, Ng30526, n299, Ng26951, Ng34035, n300, Ng34636, n301, Ng32978, n302, Ng30348, n306, Ng24336, n307, Ng29298, n308, Ng30499, n309, Ng33976, n310, Ng30335, n311, Ng34637, n312, Ng30528, n313, Ng30521, n314, Ng24239, Ng34259, n317, Ng30474, n318, Ng34643, n319, Ng30510, n320, Ng34729, n321, Ng34625, n322, Ng33029, n323, Ng33615, n324, Ng24281, n325, Ng33997, n326, Ng33584, n327, Ng24280, n328, Ng26920, n329, Ng29296, n330, n331, Ng30338, n332, Ng21895, n333, Ng34041, n334, Ng30495, n335, Ng29279, n338, Ng25655, n339, Ng30403, n340, Ng33042, n341, Ng30419, n342, Ng28090, n343, Ng34642, n344, Ng30370, n345, Ng34448, n346, Ng26946, n347, Ng34610, n348, Ng24209, n349, Ng30504, n350, Ng25669, Ng30480, n353, Ng33027, n354, Ng33972, n355, Ng28099, n356, Ng26947, n359, n357, n358, Ng24210, n360, Ng30455, n361, Ng28084, n362, Ng33993, n363, Ng30444, n364, Ng25625, n366, Ng33593, n367, Ng30502, n368, Ng33036, Ng25595, n371, Ng33024, n372, Ng33552, n373, Ng34014, n374, Ng29273, n375, Ng34638, n376, Ng30341, n377, Ng26899, n378, Ng30336, n380, n379, Ng25622, n381, Ng34447, n382, Ng33613, n383, Ng25749, Ng25704, n384, Ng33053, n385, Ng30555, n386, Ng33971, n387, Ng26915, n388, Ng30538, n389, Ng30369, n390, Ng34446, n391, Ng29230, n392, Ng33975, n393, Ng30497, n394, Ng30418, n395, Ng25721, n396, Ng34622, n397, Ng30438, n398, Ng30540, n399, Ng32986, n400, Ng33960, n401, Ng34442, n402, Ng30421, n403, Ng33573, n404, Ng24205, n405, Ng32979, n406, Ng25763, n407, Ng30481, n408, Ng30517, n409, Ng30539, n410, Ng34880, n411, Ng30436, n412, Ng32990, n413, Ng24245, n414, Ng30553, n415, Ng26907, n416, Ng24278, n417, Ng26955, n418, Ng29276, n419, Ng29277, n422, Ng31894, n423, Ng33037, n424, Ng34451, n425, Ng34250, n426, Ng29295, n427, Ng26905, n428, Ng32983, n429, Ng30402, n430, Ng33999, n431, Ng24262, n432, Ng30558, n433, Ng26901, n434, Ng33039, n435, Ng33059, n436, Ng31899, n437, Ng33007, n438, Ng30462, n439, Ng30487, n440, Ng33058, n441, Ng24261, n442, Ng30531, n443, Ng30506, n444, Ng25747, n445, Ng33601, n446, Ng26922, n447, Ng29250, Ng30459, n450, Ng33534, Ng30543, n453, Ng29275, n454, Ng34030, n455, Ng30451, n456, Ng30552, n457, Ng30337, n461, Ng24254, n462, Ng30378, n463, Ng33019, n464, Ng33623, n465, Ng29235, n466, Ng31902, n467, Ng33978, n468, Ng29278, Ng34253, n472, Ng29272, n473, Ng33610, n474, Ng33589, n475, Ng34605, n476, Ng30350, n477, Ng25611, n478, Ng33619, n479, Ng34022, n480, Ng34033, n481, Ng34726, n482, Ng31870, n483, Ng33985, n484, Ng29283, n485, Ng34003, n486, Ng34463, n487, Ng33006, n488, Ng29292, n489, Ng30557, n490, Ng33989, n491, Ng33033, n492, Ng34005, n493, Ng26932, n494, Ng30516, n495, Ng33575, n496, Ng33032, n497, Ng30486, n498, Ng30440, n499, Ng26949, n500, Ng30530, n501, Ng30542, n502, Ng25624, n503, Ng30383, n504, Ng33597, n505, Ng26957, n506, Ng28102, n507, Ng30524, n508, Ng26903, n509, Ng30475, n510, Ng34647, n511, Ng30377, n512, Ng33553, n513, Ng31903, n514, Ng33984, n515, Ng33602, n516, Ng28045, n517, Ng34603, n518, Ng33035, n519, Ng24208, n520, Ng24213, n521, Ng33614, n522, Ng33060, n523, Ng30362, n524, Ng33023, n525, Ng26898, n526, Ng25618, n527, Ng30518, n528, Ng26884, n529, Ng26933, n530, Ng28066, n531, Ng33612, n532, Ng26906, n533, Ng29269, n534, Ng34255, n535, Ng30450, n536, Ng30456, n537, Ng32991, n541, Ng24348, n542, Ng34249, n543, Ng29268, n544, Ng29224, n545, Ng33017, n546, Ng30339, n547, Ng33967, n548, Ng33559, n549, Ng29255, n550, Ng30368, n551, Ng30375, n552, Ng28089, n553, Ng33055, n554, Ng30392, n555, Ng30343, n556, Ng30523, n559, n557, Ng24233, n560, Ng33018, n561, Ng32976, n562, Ng30349, n563, Ng33067, Ng26900, n564, Ng33034, n565, Ng30551, n566, Ng25667, n567, Ng30452, n568, Ng25612, n571, n569, Ng34719, n572, Ng33607, n573, Ng26923, n574, Ng24211, n575, Ng33050, n576, Ng30463, n577, Ng34464, n578, Ng24243, n579, Ng24335, n580, Ng34611, n581, Ng34262, n582, Ng30546, n583, Ng30347, n584, Ng30556, n585, Ng33562, n586, Ng25610, n587, Ng33015, n588, Ng31896, n589, Ng34004, n590, Ng30428, n591, Ng30485, n592, Ng30422, n593, Ng30423, n594, Ng30529, Ng34028, n595, Ng30460, n596, Ng30401, n597, Ng33990, n598, Ng29309, n599, Ng30411, n600, Ng33546, n601, Ng28085, n602, Ng26904, n603, Ng25605, n604, Ng33062, n605, Ng26893, n606, Ng34626, n607, Ng33583, n608, Ng30472, n609, Ng34454, n610, Ng34850, n611, Ng24214, n612, Ng30406, n613, Ng33569, n614, Ng34628, n615, Ng34458, n616, Ng34634, n617, Ng29293, n618, Ng33009, n619, Ng24355, n620, Ng25691, n621, Ng29264, n622, Ng28072, n623, Ng31900, n624, Ng26956, n625, Ng29304, n626, Ng29261, n627, Ng28063, Ng34027, n628, Ng33961, n629, Ng32995, n630, Ng34624, n631, Ng30415, Ng33536, n633, Ng28055, n634, Ng24238, n637, Ng33600, n638, Ng28105, n639, Ng29307, n640, Ng30345, n641, Ng34453, n644, n642, n643, Ng32980, n645, Ng29238, n646, Ng34639, Ng25695, n648, Ng33057, n649, Ng29253, n650, Ng34021, n651, Ng26895, n652, Ng30413, n653, Ng30549, n654, Ng24347, Ng30501, n657, Ng33969, n658, Ng30433, n659, Ng29270, n660, Ng33038, n661, Ng26926, n662, Ng28083, n663, Ng30478, n664, Ng34724, n665, Ng26883, n666, n667, Ng32985, n668, Ng25761, n669, Ng26886, n670, Ng32982, n672, Ng33561, Ng26880, n673, Ng26931, n674, Ng34641, n675, Ng34629, n676, Ng33598, n677, Ng33576, n678, Ng26902, n679, Ng29244, n680, Ng30468, n681, Ng26924, n682, Ng33031, n683, Ng29245, n684, Ng29266, n685, Ng30559, n686, Ng28087, Ng30435, n689, n690, Ng25609, n691, Ng28057, n692, Ng34439, Ng34260, n697, Ng32989, n698, Ng34006, n699, Ng28043, n700, Ng33021, n701, Ng29251, n702, Ng34456, n703, Ng33991, n704, Ng26930, n705, Ng34599, n706, Ng33557, n707, Ng30511, n708, Ng33045, n709, Ng30379, n713, Ng24267, n714, Ng34020, n717, n715, Ng24249, n718, Ng30382, n719, Ng29285, n720, Ng33622, n721, Ng33582, n722, Ng28086, n723, Ng29262, n724, Ng24270, n725, Ng33581, n726, Ng34849, n727, Ng28060, n728, Ng33618, n729, Ng34038, n730, Ng34032, n731, Ng30509, n732, Ng34640, n733, Ng28069, n734, Ng31868, n735, Ng26938, n736, Ng30363, n737, Ng30334, n738, Ng33970, n739, Ng30391, n740, Ng33540, n741, Ng30445, n742, Ng25617, n743, Ng24215, n744, Ng33964, n745, Ng25719, n746, Ng29228, n747, Ng30514, n748, Ng33627, n749, Ng34615, n750, Ng25696, n751, Ng30493, n752, Ng33594, n753, Ng34009, n754, Ng30365, n755, Ng34018, n756, Ng34040, n757, Ng34029, n758, Ng30488, n759, Ng34600, n760, Ng25614, n761, Ng28058, n762, Ng29225, n763, Ng30532, n764, Ng33054, n765, Ng32984, n766, Ng34039, n767, Ng33065, n768, Ng30443, n769, Ng29291, n770, Ng30508, n771, Ng30464, n772, Ng33988, Ng30522, n775, Ng30374, n776, Ng34008, n777, Ng34444, n778, Ng34731, n779, Ng33606, n780, Ng24334, Ng34265, n785, Ng30482, n786, Ng34604, n787, Ng33591, n788, Ng30525, n789, Ng26929, n790, Ng30448, n791, Ng30513, n792, Ng30469, n793, Ng33608, n794, Ng33626, n795, Ng34725, n796, Ng30342, n797, Ng29267, n798, Ng30548, n799, Ng33052, n800, Ng34012, n801, Ng34017, n802, Ng26912, n803, Ng30364, n804, Ng34254, n805, Ng34251, n806, Ng30560, n807, Ng33983, n808, Ng33980, n809, Ng34631, n810, Ng29243, n811, Ng25623, n812, Ng26950, n813, Ng30431, n814, Ng30467, n815, Ng30353, n816, Ng34467, n817, Ng30442, n818, Ng29305, Ng25616, n820, Ng29252, n821, Ng33003, Ng34613, n823, Ng33570, n827, Ng24275, n828, Ng29302, n829, Ng30484, n830, Ng25634, n832, Ng33567, n833, Ng33585, n834, Ng30527, n835, Ng30447, n836, Ng25630, n837, Ng29290, n838, Ng29227, n839, Ng31872, n840, Ng29287, n841, Ng31897, n842, Ng30562, n843, Ng34011, n844, Ng33996, n845, Ng33014, n846, Ng34465, n847, Ng33995, n848, Ng30372, n849, Ng30545, n850, Ng30389, n851, Ng33590, n852, Ng34616, n853, Ng26927, n855, n854, Ng25631, n856, Ng30477, n857, Ng34632, n858, Ng28046, n859, Ng26896, n860, Ng25602, n861, Ng26916, n862, Ng33578, n863, Ng30354, n864, Ng30425, n865, Ng24200, n866, Ng33544, n867, Ng24246, n868, Ng30507, n869, Ng30333, n870, Ng32998, n871, Ng32987, n872, Ng29286, n873, Ng34606, n874, Ng33070, n875, Ng29240, n876, Ng32999, n877, Ng33605, n878, Ng24255, n879, Ng26945, n880, Ng33558, n881, Ng25699, n882, Ng29289, n883, Ng30388, n884, Ng29254, n885, Ng28074, n886, Ng34450, n887, Ng30512, n888, Ng33551, n889, Ng33538, n890, Ng33005, n891, Ng24248, n893, Ng33002, n894, Ng30471, n895, Ng34000, n896, Ng34016, n897, Ng33048, n898, Ng26934, n899, Ng34468, n900, Ng33542, n901, Ng34445, n902, Ng34013, n903, Ng26919, n904, Ng30554, n905, Ng29281, n906, Ng30537, n907, Ng34732, n908, Ng28049, n909, Ng33545, n910, Ng30441, n911, Ng29247, n912, Ng26914, n913, Ng33998, n914, Ng25626, n915, Ng33977, n916, Ng29297, n917, Ng30387, n918, Ng33577, n919, Ng33592, n920, Ng26913, n921, Ng28044, n922, Ng26948, n923, n924, Ng30344, n925, Ng33069, n926, Ng34621, n927, Ng28059, n928, Ng34633, n932, Ng24352, n933, Ng30446, n934, Ng30357, n935, Ng26908, n936, Ng30399, n937, Ng29242, n938, Ng30547, n939, Ng34010, n940, Ng33986, n941, Ng30544, n942, Ng30561, n943, Ng30430, n944, Ng33565, n945, Ng33968, n946, Ng33566, n947, Ng30465, n948, Ng28073, n949, Ng24351, n950, Ng31904, n951, Ng34635, n952, Ng29274, n953, Ng30396, n954, Ng25735, n955, Ng34037, n956, Ng34791, n957, Ng30520, n958, Ng30358, n959, Ng29299, n960, Ng28096, n961, Ng28088, n962, Ng30397, n963, Ng30409, n964, Ng29284, n965, Ng30470, n966, Ng30367, n967, Ng30359, n968, Ng25698, n969, Ng30398, n970, Ng26952, n971, Ng26928, n972, Ng26954, n973, Ng31871, n974, Ng33994, n975, Ng33586, n976, Ng31866, n977, Ng30373, n978, Ng28056, n979, Ng30355, n980, Ng30426, n983, n981, Ng34805, n984, Ng34002, n985, Ng28053, n986, Ng29229, n987, Ng33620, n988, Ng33599, n989, Ng30515, n990, Ng33979, n991, Ng30417, n992, Ng25683, n993, Ng33574, n994, Ng30410, n995, Ng30454, n996, Ng34607, n997, Ng31895, n998, Ng33068, n999, Ng29233, n1000, Ng33549, n1001, Ng29308, n1002, Ng30408, n1003, Ng29241, n1004, Ng34620, n1005, Ng25707, n1006, Ng24339, n1007, Ng34443, n1008, Ng34619, n1009, Ng30503, n1010, Ng30550, n1011, Ng33001, n1012, Ng30492, n1013, n1014, n1015, Ng26944, n1016, Ng29260, n1017, Ng33047, n1018, Ng25733, n1019, Ng30536, n1020, Ng29246, n1021, Ng33611, n1022, Ng34728, n1023, Ng29222, n1024, Ng30449, n1025, Ng34608, n1026, Ng25635, n1027, Ng30461, n1028, Ng31901, n1029, Ng29249, n1030, Ng33041, n1031, Ng33011, n1032, Ng34618, n1033, Ng33010, n1034, Ng31864, n1035, Ng34630, n1036, Ng31898, n1037, Ng25653, n1038, Ng25632, n1039, Ng29280, n1040, Ng33609, n1041, Ng30563, n1042, Ng30437, n1043, Ng30412, n1044, Ng30491, n1045, Ng30434, n1046, Ng34612, n1047, Ng25681, n1048, Ng25687, n1049, Ng30479, n1050, Ng29256, n1051, Ng30535, n1052, Ng30385, n1053, Ng25705, n1054, Ng29257, n1055, Ng34461, n1056, Ng34258, n1057, Ng32993, n1058, Ng33992, n1059, Ng30394, n1061, Ng34449, n1062, Ng34019, n1063, Ng30395, n1064, Ng25598, n1065, Ng33987, n1066, Ng30380, n1067, Ng30400, n1068, Ng34623, n1069, Ng24343, n1070, Ng30473, n1071, Ng33028, n1072, Ng29258, n1073, Ng30407, n1074, Ng26958, n1075, Ng34457, n1076, Ng33568, n1077, Ng26964, n1078, Ng30352, n1079, Ng33543, n1083, Ng24271, n1084, Ng33981, n1085, Ng30500, n1086, n1090, n1088, n1087, n1092, Ng34992, n1094, n1093, n1096, n1099, n1100, n1097, n1101, n1104, Ng34991, n1107, n1108, n1110, n1111, n1109, n1112, n1114, n1113, n1118, n1116, Ng34994, Ng34990, n1119, Ng34993, n1120, n1121, Ng34996, n1124, n1122, n1126, Ng34879, n1129, n1131, n1132, Ng34997, n1133, n1134, n1136, n1135, n1139, n1138, n1140, n1141, Ng34995, n1142, n1145, n1146, Ng34847, n1150, n1151, n1153, n1155, n1158, n1156, n1160, n1162, n1166, n1165, Ng34878, n1168, n1169, n1170, Ng21726, n1173, n1172, n1176, n1175, Ng34848, n1178, n1180, n1179, n1182, n1184, Ng35002, n1187, n1189, Ng34789, n1191, n1192, n1195, n1194, n1197, n1196, n1199, n1201, Ng25692, n1203, n1205, n1209, n1211, n1215, n1216, n1212, n1219, n1217, n1218, n1221, n1222, n1220, n1224, n1223, n1226, n1228, n1229, n1230, n1231, n1227, n1233, n1234, n1235, n1236, n1232, n1240, n1238, n1239, n1237, Ng34787, Ng34786, n1242, n1243, n1245, n1248, n1250, n1253, n1255, n1256, n1254, n1258, n1257, n1261, n1260, n1264, n1263, n1266, n1265, n1268, n1267, n1270, n1269, n1272, n1271, n1274, n1273, n1278, n1279, n1277, n1275, n1282, n1283, n1281, n1280, n1284, n1285, n1286, n1287, n1291, n1292, n1289, n1288, n1296, n1297, n1294, n1293, n1298, n1299, n1300, n1303, n1304, n1301, n1305, n1306, n1307, n1308, n1312, n1313, n1310, n1309, n1314, n1315, n1316, n1317, n1320, n1321, n1318, n1325, n1326, n1323, n1322, n1327, n1328, n1329, n1333, n1334, n1331, n1330, n1335, n1336, n1337, n1338, n1341, n1342, n1339, n1345, n1346, n1343, n1347, n1348, n1349, n1353, n1354, n1351, n1350, n1355, n1356, n1357, n1358, n1362, n1359, n1363, n1366, n1368, n1369, n1372, n1371, n1376, n1374, n1375, n1373, n1377, n1378, n1380, n1381, n1379, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1392, n1393, n1396, n1397, n1395, n1399, n1400, n1398, n1402, n1403, n1404, n1405, n1401, n1409, n1406, n1407, n1408, n1410, n1411, n1413, n1414, n1412, n1416, n1417, n1415, n1418, n1419, n1421, n1422, n1425, n1426, n1428, n1429, n1432, n1433, n1435, n1437, n1438, n1436, n1440, n1441, n1439, n1452, n1454, n1456, n1458, n1462, n1464, n1466, n1468, n1472, n1474, n1476, n1478, n1480, n1485, n1487, n1489, n1491, n1493, n1495, n1497, n1499, n1501, n1502, n1505, n1507, n1508, n1510, n1512, n1514, n1516, n1518, n1520, n1522, n1523, n1521, n1525, n1526, n1524, n1531, n1530, n1532, n1533, n1537, n1541, n1540, n1542, n1543, n1547, n1549, n1548, n1551, n1552, n1555, n1557, n1556, n1558, n1560, n1559, n1562, n1563, n1564, n1570, n1569, n1574, n1572, n1576, n1577, n1578, n1579, n1582, n1583, n1584, n1587, n1588, n1589, n1593, n1591, n1592, n1594, n1596, n1595, n1597, n1599, n1598, n1600, n1602, n1601, n1603, n1605, n1604, n1606, n1607, n1608, n1609, n1610, n1611, n1613, n1614, n1612, n1617, n1621, n1620, n1622, n1627, n1628, n1626, n1631, n1629, n1635, n1633, n1634, n1632, n1638, n1636, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1651, n1653, n1656, n1657, n1655, n1658, n1663, n1660, n1664, n1666, n1669, n1670, n1668, n1671, n1675, n1679, n1677, n1681, n1683, n1684, n1682, n1687, n1685, n1689, n1690, n1691, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1706, n1709, n1713, n1710, n1711, n1715, n1716, n1717, n1718, n1719, n1720, n1722, n1725, n1729, n1726, n1727, n1731, n1732, n1733, n1734, n1736, n1737, n1735, n1739, n1742, n1743, n1747, n1745, n1750, n1751, n1749, n1753, n1754, n1756, n1757, n1755, n1759, n1760, n1758, n1762, n1763, n1761, n1765, n1767, n1768, n1773, n1771, n1776, n1775, n1779, n1780, n1782, n1783, n1781, n1785, n1786, n1784, n1788, n1789, n1787, n1791, n1793, n1794, n1798, n1796, n1801, n1800, n1804, n1805, n1807, n1808, n1806, n1810, n1811, n1809, n1813, n1814, n1812, n1816, n1818, n1819, n1823, n1821, n1826, n1827, n1825, n1829, n1830, n1832, n1833, n1831, n1835, n1836, n1834, n1838, n1839, n1837, n1841, n1844, n1845, n1849, n1847, n1852, n1853, n1851, n1855, n1856, n1858, n1859, n1857, n1861, n1862, n1860, n1864, n1865, n1863, n1867, n1869, n1870, n1875, n1873, n1878, n1879, n1877, n1881, n1882, n1884, n1885, n1883, n1887, n1888, n1886, n1890, n1891, n1889, n1893, n1895, n1896, n1900, n1898, n1903, n1902, n1906, n1907, n1909, n1910, n1908, n1912, n1913, n1911, n1915, n1916, n1914, n1918, n1920, n1921, n1925, n1923, n1928, n1929, n1927, n1931, n1932, n1930, n1934, n1935, n1933, n1937, n1938, n1936, n1940, n1941, n1939, n1943, n1944, n1942, n1947, n1945, n1949, n1950, n1952, n1953, n1957, n1956, n1954, n1961, n1962, n1960, n1966, n1965, n1963, n1970, n1971, n1969, n1975, n1974, n1972, n1979, n1980, n1978, n1982, n1983, n1987, n1986, n1984, n1991, n1992, n1990, n1994, n1995, n1993, n1999, n1998, n1996, n2003, n2004, n2002, n2008, n2007, n2005, n2012, n2013, n2011, n2017, n2016, n2014, n2021, n2022, n2024, n2023, n2027, n2025, n2030, n2033, n2034, n2036, n2038, n2037, n2042, n2043, n2044, n2046, n2047, n2051, n2054, n2055, n2057, n2059, n2058, n2063, n2064, n2065, n2067, n2068, n2072, n2075, n2076, n2078, n2080, n2079, n2084, n2085, n2086, n2088, n2089, n2093, n2096, n2097, n2099, n2101, n2100, n2105, n2106, n2107, n2109, n2110, n2114, n2117, n2118, n2120, n2122, n2121, n2126, n2127, n2128, n2130, n2131, n2135, n2138, n2139, n2141, n2143, n2142, n2147, n2148, n2149, n2151, n2152, n2156, n2159, n2160, n2162, n2164, n2163, n2168, n2169, n2170, n2172, n2173, n2177, n2180, n2181, n2183, n2185, n2186, n2187, n2188, n2191, n2194, n2192, n2195, n2196, n2197, n2203, n2204, n2207, n2205, n2208, n2209, n2210, n2216, n2217, n2219, n2220, n2218, n2223, n2221, n2225, n2226, n2228, n2229, n2232, n2230, n2233, n2235, n2237, n2238, n2242, n2241, n2240, n2245, n2244, n2243, n2246, n2248, n2250, n2251, n2255, n2254, n2253, n2258, n2256, n2259, n2261, n2263, n2264, n2268, n2267, n2266, n2271, n2270, n2269, n2272, n2274, n2276, n2277, n2281, n2280, n2279, n2284, n2283, n2282, n2285, n2287, n2289, n2290, n2294, n2293, n2292, n2296, n2297, n2302, n2301, n2304, n2309, n2310, n2308, n2312, n2317, n2316, n2320, n2319, n2318, n2321, n2323, n2325, n2326, n2330, n2329, n2328, n2333, n2332, n2331, n2334, n2336, n2338, n2339, n2343, n2342, n2341, n2346, n2345, n2344, n2347, n2349, n2351, n2352, n2356, n2355, n2354, n2358, n2357, n2361, n2359, n2363, n2364, n2366, n2367, n2369, n2368, n2370, n2371, n2374, n2372, n2376, n2377, n2379, n2380, n2382, n2381, n2384, n2385, n2388, n2386, n2390, n2391, n2393, n2394, n2396, n2395, n2397, n2398, n2401, n2399, n2403, n2404, n2406, n2407, n2409, n2408, n2410, n2411, n2414, n2412, n2416, n2417, n2419, n2420, n2422, n2421, n2424, n2425, n2428, n2426, n2430, n2431, n2433, n2434, n2436, n2435, n2437, n2438, n2441, n2439, n2443, n2444, n2446, n2447, n2449, n2448, n2450, n2451, n2454, n2452, n2456, n2457, n2459, n2460, n2462, n2461, n2463, n2464, n2466, n2467, n2469, n2470, n2468, n2472, n2473, n2475, n2476, n2474, n2478, n2479, n2477, n2482, n2480, n2484, n2485, n2487, n2488, n2489, n2490, n2491, n2492, n2498, n2501, n2505, n2503, n2507, n2508, n2511, n2509, n2514, n2517, n2519, n2522, n2521, n2520, n2527, n2526, n2532, n2533, n2535, n2536, n2538, n2539, n2541, n2542, n2544, n2545, n2547, n2548, n2546, n2550, n2551, n2549, n2553, n2554, n2555, n2563, n2562, n2560, n2561, n2559, n2567, n2564, n2565, n2569, n2572, n2573, n2571, n2574, n2577, n2578, n2576, n2580, n2579, n2583, n2584, n2582, n2586, n2587, n2585, n2589, n2590, n2588, n2592, n2593, n2591, n2595, n2594, n2598, n2599, n2597, n2601, n2602, n2600, n2604, n2605, n2603, n2607, n2608, n2606, n2610, n2611, n2609, n2613, n2614, n2612, n2616, n2617, n2615, n2619, n2620, n2618, n2622, n2623, n2621, n2625, n2626, n2624, n2628, n2630, n2631, n2629, n2632, n2633, n2635, n2636, n2634, n2638, n2639, n2637, n2641, n2642, n2640, n2644, n2645, n2643, n2647, n2648, n2646, n2650, n2651, n2649, n2653, n2652, n2656, n2655, n2659, n2660, n2658, n2662, n2661, n2665, n2666, n2664, n2668, n2669, n2667, n2671, n2672, n2670, n2674, n2675, n2673, n2677, n2678, n2676, n2680, n2681, n2679, n2683, n2684, n2682, n2686, n2688, n2689, n2687, n2690, n2693, n2694, n2692, n2696, n2695, n2699, n2700, n2698, n2702, n2703, n2701, n2705, n2706, n2704, n2708, n2709, n2707, n2711, n2710, n2714, n2715, n2713, n2717, n2718, n2716, n2720, n2721, n2719, n2723, n2724, n2722, n2726, n2727, n2725, n2729, n2730, n2728, n2732, n2733, n2731, n2735, n2736, n2734, n2738, n2739, n2737, n2741, n2742, n2740, n2744, n2746, n2747, n2745, n2748, n2751, n2752, n2750, n2754, n2755, n2753, n2757, n2758, n2756, n2760, n2761, n2759, n2763, n2764, n2762, n2766, n2767, n2765, n2769, n2768, n2772, n2773, n2771, n2775, n2776, n2774, n2778, n2779, n2777, n2781, n2782, n2780, n2784, n2785, n2783, n2787, n2788, n2786, n2790, n2791, n2789, n2793, n2794, n2792, n2796, n2797, n2795, n2799, n2800, n2798, n2802, n2804, n2805, n2803, n2806, n2807, n2809, n2810, n2808, n2812, n2813, n2811, n2815, n2816, n2814, n2818, n2817, n2821, n2822, n2820, n2824, n2823, n2827, n2826, n2830, n2831, n2829, n2833, n2834, n2832, n2836, n2837, n2835, n2839, n2840, n2838, n2842, n2843, n2841, n2845, n2846, n2844, n2848, n2849, n2847, n2851, n2852, n2850, n2854, n2855, n2853, n2857, n2858, n2856, n2860, n2859, n2862, n2863, n2864, n2865, n2861, n2867, n2868, n2870, n2872, n2873, n2871, n2874, n2875, n2877, n2878, n2876, n2880, n2881, n2879, n2883, n2884, n2882, n2886, n2885, n2889, n2890, n2888, n2892, n2891, n2895, n2894, n2898, n2899, n2897, n2901, n2902, n2900, n2904, n2905, n2903, n2907, n2908, n2906, n2910, n2911, n2909, n2913, n2914, n2912, n2916, n2917, n2915, n2919, n2920, n2918, n2922, n2923, n2921, n2925, n2926, n2924, n2928, n2930, n2931, n2929, n2932, n2933, n2935, n2936, n2934, n2938, n2939, n2937, n2941, n2942, n2940, n2944, n2943, n2947, n2948, n2946, n2950, n2951, n2949, n2953, n2952, n2956, n2957, n2955, n2959, n2960, n2958, n2962, n2961, n2965, n2966, n2964, n2968, n2969, n2967, n2971, n2972, n2970, n2974, n2975, n2973, n2977, n2978, n2976, n2980, n2981, n2979, n2983, n2984, n2982, n2986, n2988, n2989, n2987, n2990, n2991, n2993, n2994, n2992, n2996, n2997, n2995, n2999, n3000, n2998, n3002, n3003, n3001, n3005, n3006, n3004, n3008, n3009, n3007, n3011, n3010, n3014, n3013, n3017, n3018, n3016, n3020, n3019, n3023, n3024, n3022, n3026, n3027, n3025, n3029, n3030, n3028, n3032, n3033, n3031, n3035, n3036, n3034, n3038, n3039, n3037, n3041, n3042, n3040, n3043, n3044, n3045, n3046, n3050, n3048, n3053, n3056, n3059, n3062, n3060, n3065, n3068, n3071, n3074, n3072, n3077, n3080, n3083, n3086, n3084, n3089, n3092, n3095, n3098, n3096, n3101, n3104, n3107, n3110, n3108, n3113, n3116, n3119, n3122, n3120, n3125, n3128, n3131, n3134, n3132, n3137, n3140, n3141, n3148, n3152, n3151, n3154, n3155, n3157, n3158, n3156, n3160, n3159, n3163, n3168, n3167, n3170, n3171, n3173, n3174, n3172, n3176, n3177, n3175, n3179, n3180, n3178, n3181, n3182, n3185, n3184, n3187, n3189, n3188, n3192, n3194, n3198, n3202, n3209, n3210, n3208, n3207, n3211, n3214, n3218, n3219, n3220, n3217, n3225, n3223, n3221, n3229, n3227, n3226, n3233, n3234, n3232, n3230, n3236, n3235, n3239, n3238, n3241, n3243, n3242, n3247, n3249, n3253, n3257, n3264, n3265, n3263, n3262, n3266, n3269, n3273, n3274, n3275, n3272, n3278, n3277, n3276, n3282, n3281, n3279, n3286, n3287, n3285, n3283, n3289, n3288, n3292, n3291, n3294, n3296, n3295, n3300, n3302, n3306, n3310, n3317, n3318, n3316, n3315, n3319, n3322, n3326, n3327, n3328, n3325, n3333, n3331, n3329, n3337, n3335, n3334, n3341, n3342, n3340, n3338, n3344, n3343, n3347, n3346, n3349, n3351, n3350, n3355, n3357, n3361, n3365, n3372, n3373, n3371, n3370, n3374, n3377, n3381, n3382, n3383, n3380, n3388, n3386, n3384, n3392, n3391, n3389, n3396, n3397, n3395, n3393, n3400, n3402, n3401, n3404, n3406, n3405, n3410, n3412, n3417, n3421, n3426, n3427, n3425, n3428, n3431, n3435, n3436, n3437, n3434, n3442, n3440, n3438, n3446, n3444, n3443, n3450, n3451, n3447, n3453, n3452, n3455, n3457, n3458, n3456, n3459, n3464, n3466, n3467, n3465, n3468, n3473, n3474, n3477, n3476, n3479, n3481, n3480, n3485, n3487, n3491, n3495, n3502, n3503, n3501, n3500, n3504, n3507, n3511, n3512, n3513, n3510, n3518, n3516, n3514, n3522, n3520, n3519, n3526, n3527, n3525, n3523, n3529, n3528, n3532, n3531, n3534, n3536, n3535, n3539, n3541, n3546, n3550, n3555, n3556, n3554, n3557, n3560, n3564, n3565, n3566, n3563, n3570, n3567, n3574, n3572, n3571, n3578, n3579, n3577, n3575, n3581, n3580, n3584, n3583, n3585, n3587, n3586, n3591, n3593, n3597, n3602, n3608, n3609, n3607, n3606, n3610, n3613, n3617, n3618, n3619, n3616, n3621, n3620, n3625, n3624, n3622, n3629, n3630, n3628, n3626, n3633, n3635, n3634, n3636, n3640, n3639, n3642, n3647, n3648, n3646, n3651, n3652, n3653, n3657, n3656, n3659, n3664, n3665, n3663, n3668, n3669, n3672, n3670, n3673, n3676, n3681, n3682, n3680, n3685, n3686, n3689, n3687, n3690, n3693, n3698, n3699, n3697, n3702, n3703, n3706, n3704, n3707, n3710, n3715, n3716, n3714, n3719, n3720, n3723, n3721, n3724, n3727, n3732, n3733, n3731, n3736, n3737, n3738, n3742, n3741, n3744, n3749, n3750, n3748, n3753, n3754, n3755, n3759, n3758, n3761, n3766, n3767, n3765, n3770, n3771, n3774, n3772, n3776, n3777, n3780, n3778, n3782, n3783, n3786, n3784, n3788, n3789, n3790, n3791, n3794, n3793, n3797, n3798, n3800, n3801, n3802, n3803, n3806, n3807, n3805, n3809, n3810, n3813, n3812, n3815, n3816, n3817, n3818, n3819, n3821, n3822, n3820, n3824, n3823, n3826, n3827, n3825, n3829, n3828, n3830, n3832, n3834, n3835, n3833, n3836, n3838, n3839, n3837, n3841, n3840, n3843, n3844, n3842, n3846, n3845, n3847, n3849, n3851, n3852, n3850, n3854, n3853, n3858, n3861, n3862, n3855, n3860, n3863, n3864, n3865, n3866, n3868, n3867, n3869, n3870, n3871, n3873, n3872, n3876, n3875, n3878, n3879, n3877, n3882, n3881, n3884, n3885, n3883, n3887, n3888, n3890, n3891, n3893, n3894, n3900, n3901, n3899, n3903, n3902, n3904, n3907, n3906, n3911, n3914, n3915, n3916, n3918, n3923, n3920, n3926, n3925, n3929, n3933, n3934, n3935, n3937, n3936, n3940, n3943, n3942, n3948, n3949, n3950, n3952, n3953, n3955, n3954, n3957, n3959, n3961, n3963, n3965, n3967, n3969, n3971, n3973, n3974, n3976, n3977, n3979, n3980, n3983, n3984, n3985, n3986, n3990, n3993, n3994, n3996, n3997, n3999, n4000, n4003, n4004, n4005, n4010, n4014, n4017, n4018, n4019, n4021, n4023, n4025, n4027, n4029, n4031, n4033, n4035, n4036, n4037, n4039, n4044, n4047, n4048, n4046, n4049, n4052, n4055, n4059, n4060, n4058, n4063, n4061, n4064, n4067, n4070, n4071, n4073, n4076, n4077, n4079, n4082, n4083, n4085, n4088, n4089, n4091, n4094, n4095, n4092, n4097, n4096, n4100, n4101, n4102, n4106, n4103, n4110, n4107, n4112, n4113, n4115, n4114, n4117, n4120, n4121, n4123, n4126, n4127, n4129, n4132, n4133, n4135, n4136, n4134, n4138, n4139, n4140, n4141, n4144, n4142, n4149, n4152, n4154, n4155, n4156, n4157, n4160, n4158, n4165, n4168, n4170, n4169, n4176, n4177, n4178, n4182, n4183, n4180, n4186, n4184, n4192, n4190, n4196, n4198, n4200, n4202, n4203, n4201, n4204, n4205, n4208, n4210, n4209, n4211, n4212, n4218, n4217, n4220, n4221, n4222, n4223, n4226, n4225, n4227, n4228, n4231, n4233, n4234, n4235, n4236, n4239, n4238, n4241, n4242, n4245, n4246, n4248, n4247, n4251, n4253, n4256, n4259, n4261, n4263, n4265, n4266, n4267, n4268, n4271, n4270, n4272, n4275, n4274, n4276, n4277, n4279, n4280, n4281, n4283, n4285, n4286, n4288, n4287, n4290, n4289, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, Ng25599, n4300, n4301, n4303, n4302, n4304, n4307, n4305, n4309, n4308, n4311, n4310, n4313, n4312, n4315, n4314, n4317, n4316, n4319, n4318, n4321, n4320, n4322, n4323, n4325, n4324, n4327, n4326, n4329, n4328, n4331, n4330, n4333, n4332, n4335, n4334, n4337, n4336, n4339, n4338, n4341, n4340, n4343, n4342, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4356, n4355, n4358, n4357, n4359, n4360, n4361, n4363, n4365, n4364, n4366, n4368, n4367, n4371, n4374, n4376, n4379, n4380, n4382, n4381, n4385, n4384, n4387, n4388, n4389, n4392, n4393, n4394, n4397, n4398, n4401, n4402, n4403, n4404, n4406, n4407, n4411, Ng29209, n4412, n4414, n4416, n4417, n4419, n4418, n4421, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4441, n4442, n4443, n4444, n4449, n4464, n4465, n4486, n4487, n4488, n4490, n4492, n4503, n4508, n4509, n4510, n4511, n4512, n4515, n4516, n4518, n4521, n4527, n4531, n4532, n4530, n4533, n4535, n4536, n4538, n4540, n4542, n4544, n4546, n4548, n4550, n4551, n4553, n4556, n4559, n4561, n4564, n4567, n4569, n4568, n4570, n4577, n4581, n4582, n4584, n4585, n4587, n4588, n4590, n4593, n4595, n4596, n4597, n4630, n4632, n4633, n4635, n4637, n4638, n4640, n4641, n4642, n4652, n4653, n4654, n4659, n4657, n4660, n4661, n4663, n4664, n4666, n4667, n4669, n4670, n4672, n4673, n4674, n4676, n4677, n4689, n4690, n4691, n4692, n4695, n4696, n4697, n4699, n4700, n4702, n4703, n4704, n4706, n4707, n4709, n4710, n4712, n4713, n4714, n4716, n4717, n4719, n4720, n4722, n4723, n4724, n4726, n4727, n4729, n4730, n4731, n4733, n4734, n4736, n4737, n4738, n4740, n4741, n4742, n4744, n4745, n4747, n4748, n4750, n4751, n4752, n4754, n4755, n4757, n4758, n4760, n4761, n4763, n4764, n4765, n4767, n4768, n4770, n4771, n4773, n4774, n4776, n4777, n4778, n4779, n4781, n4783, n4784, n4786, n4787, n4790, n4791, n4792, n4793, n4794, n4796, n4806, n4807, n4805, n4808, n4810, n4813, n4819, n4820, n4818, n4821, n4823, n4826, n4830, n4832, Ng25756, n4833, n4835, n4836, Ng25728, n4837, n4838, n4839, n4840, n4842, n4844, n4845, n4846, n4848, n4849, n4851, n4852, n4853, n4854, n4850, n4855, n4856, n4857, n4859, n4860, n4862, n4864, n4866, n4868, n4870, n4873, n4875, n4878, n4881, n4883, n4884, n4886, n4887, n4888, n4889, n4893, n4894, n4895, n4896, n4900, n4901, n4902, n4903, n4907, n4908, n4909, n4910, n4914, n4915, n4916, n4919, n4922, n4923, n4924, n4927, n4928, n4929, n4930, n4933, n4934, n4935, n4936, n4940, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4977, n4983, n4984, n4990, n4991, n4998, n4999, n5005, n5006, n5011, n5012, n5013, n5023, n5024, n5030, n5031, n5034, n5038, n5039, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5051, n5052, n5054, n5056, n5057, n5058, n5068, n5070, n5071, n5075, n5074, n5076, n5077, n5079, n5081, n5083, n5084, n5085, n5086, n5088, n5089, n5090, n5091, n5092, n5093, n5095, n5094, n5096, n5109, n5122, n5130, n5132, n5133, n5135, n5136, n5137, n5139, n5140, n5142, n5143, n5145, n5147, n5149, n5150, n5151, n5152, n5154, n5160, n5162, n5163, n5165, n5167, n5168, n5170, n5172, n5175, n5174, n5176, n5177, n5178, n5180, n5179, n5181, n5182, n5183, Ng26965, Ng26910, Ng25697, n5184, n5185, n5186, Ng24260, Ng24257, Ng24244, Ng24241, n5189, n5187, n5192, n5190, n5193, Ng34980, n5194, Ng34882, n5195, Ng34808, n5196, Ng34807, n5197, Ng34806, n5198, Ng34804, n5199, Ng34803, n5200, Ng34802, n5201, Ng34801, n5202, n5203, Ng34800, n5204, n5205, Ng34799, n5206, n5207, Ng34798, n5208, n5209, Ng34797, n5210, Ng34796, n5211, n5213, Ng34795, n5214, n5215, Ng34794, n5216, Ng34793, n5217, Ng34792, n5218, n5219, Ng34735, n5220, n5221, Ng34734, n5222, n5223, Ng34730, n5224, n5225, Ng34727, n5226, n5227, Ng34723, n5228, n5229, Ng34722, n5230, n5231, Ng34721, n5232, n5233, Ng34720, n5234, Ng34614, Ng34602, Ng34601, n5237, Ng34598, n5238, Ng34466, n5239, Ng34462, n5240, Ng34459, n5241, Ng34440, n5242, Ng34269, n5243, Ng34268, n5244, Ng34266, n5245, Ng34264, n5246, Ng34263, n5247, Ng34261, n5248, n5249, Ng34257, n5250, Ng34256, n5252, n5253, Ng34024, n5255, n5256, Ng34023, n5259, n5257, n5262, n5260, n5265, n5263, n5268, n5266, n5271, n5269, n5274, n5272, n5277, n5275, n5280, n5278, n5282, n5281, n5283, Ng33963, n5286, n5287, n5285, n5284, n5288, Ng33962, n5290, n5291, Ng33621, n5292, Ng33617, n5293, Ng33616, n5295, n5296, Ng33604, n5297, Ng33603, n5299, n5300, Ng33596, n5301, Ng33595, n5303, n5304, Ng33588, n5305, Ng33587, n5307, n5308, Ng33580, n5309, Ng33579, n5311, n5312, Ng33572, n5313, Ng33571, n5315, n5316, Ng33564, n5317, Ng33563, n5319, n5320, Ng33556, n5321, Ng33555, n5323, n5324, Ng33548, n5325, Ng33547, n5326, Ng33537, n5327, n5328, n5329, Ng31865, n5330, Ng30457, n5331, Ng30386, n5332, Ng30381, n5333, Ng30376, n5334, Ng30371, n5335, Ng30366, n5336, Ng30361, n5337, Ng30356, n5338, Ng30351, n5339, n5340, Ng30346, n5341, n5342, Ng30340, n5343, Ng29306, n5344, Ng29300, n5345, Ng29294, n5346, Ng29288, n5347, Ng29282, n5348, n5350, n5352, Ng29271, n5353, Ng29265, n5354, Ng29259, n5355, Ng29239, n5357, n5356, n5358, Ng29237, n5359, Ng29236, n5360, Ng29234, n5362, n5361, n5363, Ng29232, n5364, Ng29231, n5365, Ng28092, n5366, Ng28091, n5367, Ng28082, n5368, Ng28081, n5369, Ng28071, n5370, Ng28054, n5371, Ng28052, n5372, Ng28051, n5373, Ng28050, n5374, Ng28048, n5375, Ng28047, n5376, Ng26971, n5377, Ng26970, n5378, Ng26969, n5379, Ng26968, n5380, Ng26967, n5381, Ng26966, n5382, Ng26963, n5383, Ng26962, n5384, Ng26961, n5385, Ng26940, n5386, Ng26939, n5387, Ng26937, n5388, Ng26925, n5389, Ng26921, n5390, Ng26918, n5391, Ng26909, n5392, n5393, Ng26897, n5394, n5396, Ng26894, n5397, n5398, Ng26892, n5399, Ng26891, n5400, Ng26890, n5402, Ng26889, n5403, Ng26888, n5404, Ng26887, n5405, Ng26882, n5406, Ng26881, n5407, Ng25764, n5409, n5410, Ng25762, n5411, n5413, Ng25758, n5414, Ng25757, n5415, Ng25750, n5417, n5418, Ng25748, n5419, n5421, Ng25744, n5422, Ng25743, n5423, Ng25736, n5425, n5426, Ng25734, n5427, n5429, Ng25730, n5430, Ng25729, n5431, Ng25722, n5433, n5434, Ng25720, n5435, n5437, Ng25716, n5438, Ng25715, n5439, Ng25708, n5441, n5442, Ng25706, n5443, n5445, Ng25703, n5446, n5448, Ng25702, n5449, Ng25701, n5450, n5451, Ng25686, n5452, Ng25684, n5454, n5455, Ng25682, n5456, n5458, Ng25678, n5459, Ng25677, n5460, Ng25670, n5462, n5463, Ng25668, n5464, n5466, Ng25664, n5467, Ng25663, n5468, Ng25656, n5470, n5471, Ng25654, n5472, n5474, Ng25650, n5475, Ng25649, n5476, Ng25638, n5477, n5479, Ng25637, n5480, Ng25636, n5481, Ng25629, n5482, n5483, Ng25628, n5484, Ng25627, n5485, n5486, Ng25615, n5487, Ng25604, n5488, Ng25601, n5489, Ng25600, n5490, Ng25597, n5491, Ng25596, n5492, Ng25593, n5493, Ng25592, n5494, Ng25591, n5495, Ng24354, n5496, Ng24353, n5497, Ng24350, n5498, Ng24349, n5499, Ng24346, n5500, Ng24345, n5501, Ng24342, n5502, Ng24341, n5503, Ng24338, n5504, Ng24337, n5505, Ng24282, n5506, Ng24279, n5507, Ng24277, n5508, Ng24276, n5509, Ng24273, n5510, Ng24272, n5511, Ng24269, n5512, Ng24268, n5513, Ng24258, n5514, Ng24256, n5515, Ng24253, n5516, Ng24252, n5517, Ng24251, n5518, Ng24250, n5519, Ng24242, n5520, Ng24240, n5521, Ng24237, n5522, Ng24236, n5523, Ng24235, n5524, Ng24234, n5525, Ng24216, n5526, Ng24207, n5527, Ng24206, n5528, Ng24204, n5529, Ng24203, n5530, Ng24202, n5531, Ng24201, n5532, Ng21901, n5533, Ng21900, n5534, Ng21899, n5535, Ng21898, n5536, Ng21897, n5537, Ng21896, n5538, Ng21892, n5539, Ng21891, n5540, n5541, n5543, n5545, n5544, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5554, n5553, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5576, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5593, n5595, n5597, n5599, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5622, n5623, n5621, n5626, n5627, n5625, n5630, n5631, n5634, n5635, n5636, n5637, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5648, n5649, n5652, n5651, n5655, n5654, n5658, n5657, n5660, n5664, n5663, n5666, n5670, n5669, n5677, n5676, n5682, n5681, n5685, n5684, n5687, n5688, n5698, n5699, n5700, n5701, n5704, n5705, n5706, n5710, n5712, n5715, n5717, n5719, n5721, n5723, n5724, n5725, n5726, n5727, n5730, n5731, n5732, n5733, n5734, n5735, n5737, n5738, n5740, n5741, n5743, n5744, n5746, n5747, n5749, n5750, n5752, n5754, n5755, n5756, n5757, n5758, n5760, n5777, n5775, n5781, n5785, n5793, n5794, n5795, n5799, n5809, n5812, n5815, n5816, n5817, n5818, n5819, n5821, n5825, n5828, n5829, n5830, n5831, n5832, n5833, n5835, n5836, n5837, n5838, n5840, n5842, n5843, n5845, n5847, n5848, n5850, n5852, n5853, n5855, n5857, n5858, n5860, n5862, n5863, n5865, n5867, n5868, n5870, n5872, n5873, n5875, n5877, n5878, n5879, n5880, n5883, n5885, n5886, n5888, n5891, n5893, n5894, n5896, n5900, n5902, n5903, n5905, n5908, n5910, n5911, n5913, n5916, n5918, n5919, n5921, n5922, n5923, n5924, n5925, n5928, n5930, n5931, n5933, n5936, n5938, n5939, n5941, n5944, n5946, n5947, n5949, n5951, n5952, n5953, n5957, n5958, n5961, n5962, n5965, n5966, n5970, n5971, n5974, n5975, n5978, n5980, n5982, n5984, n5983, n5985, n5986, n5988, n5987, n5989, n5992, n5993, n5994, n5995, n5999, n6001, n6002, n6003, n6004, n6005, n6007, n6010, n6011, n6013, n6022, n6023, n6029, n6032, n6033, n6036, n6035, n6037, n6040, n6041, n6044, n6043, n6047, n6048, n6050, n6052, n6057, n6055, n6059, n6060, n6062, n6063, n6065, n6066, n6068, n6069, n6071, n6072, n6074, n6075, n6078, n6077, n6076, n6079, n6082, n6083, n6085, n6086, n6088, n6089, n6093, n6092, n6094, n6095, n6098, n6097, n6099, n6100, n6102, n6107, n6106, n6105, n6109, Ng25676, Ng25694, Ng25648, Ng34025, Ng25714, Ng25700, Ng24212, Ng25662, Ng24247, Ng24231, Ng26953, Ng21893, Ng25742, Ng28079, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6123, n6124, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6174, n6186, n6188, n6200, n6201, n6203, n6207, n6214, n6218, n6234, n6244, n6251, n6256, n6261, n6263, n6268, n6287, n6288, n6290, n6299, n6301, n6306, n6318, n6325, n6341, n6343, n6344, n6364, n6366, n6367, n6383, n6386, n6389, n6405, n6406, n6408, n6431, n6435, n6444, Ng32996, Ng32992, Ng32988, Ng24263, Ng33040, Ng33016, Ng33012, Ng33008, Ng33004, Ng33000, Ng25685, Ng25639, Ng33044, Ng30458;

reg Ng5057, Ng2771, Ng1882, Ng2299, Ng4040, Ng2547, Ng559, Ng3243, Ng452, Ng3542, Ng5232, Ng5813, Ng2907, Ng1744, Ng5909, Ng1802, Ng3554, Ng6219, Ng807, Ng6031, Ng847, Ng976, Ng4172, Ng4372, Ng3512, Ng749, Ng3490, Pg12350, Ng4235, Ng1600, Ng1714, Pg14451, Ng3155, Ng2236, Ng4555, Ng3698, Ng1736, Ng1968, Ng4621, Ng5607, Ng2657, Pg12300, Ng490, Ng311, Ng772, Ng5587, Ng6177, Ng6377, Ng3167, Ng5615, Ng4567, Ng3457, Ng6287, Pg7946, Ng2563, Ng4776, Ng4593, Ng6199, Ng2295, Ng1384, Ng1339, Ng5180, Ng2844, Ng1024, Ng5591, Ng3598, Ng4264, Ng767, Ng5853, Pg13865, Ng2089, Ng4933, Ng4521, Ng5507, Pg16656, Ng6291, Ng294, Ng5559, Pg9617, Pg9741, Ng3813, Ng562, Ng608, Ng1205, Ng3909, Ng6259, Ng5905, Ng921, Ng2955, Ng203, Ng1099, Ng4878, Ng5204, Pg17604, Ng3606, Ng1926, Ng6215, Ng3586, Ng291, Ng4674, Ng3570, Pg9048, Pg17607, Ng1862, Ng676, Ng843, Ng4332, Ng4153, Pg17711, Ng6336, Ng622, Ng3506, Ng4558, Pg17685, Ng3111, wire4430, Ng26936, Ng939, Ng278, Ng4492, Ng4864, Ng1036, wire4427, Ng1178, Ng3239, Ng718, Ng6195, Ng1135, Ng6395, wire4415, Ng554, Ng496, Ng3853, Ng5134, Pg17404, Pg8344, Ng2485, Ng925, Ng48, Ng5555, Pg14096, Ng1798, Ng4076, Ng2941, Ng3905, Ng763, Ng6255, Ng4375, Ng4871, Ng4722, Ng590, Pg13099, Ng1632, Pg12238, Ng3100, Ng1495, Ng1437, Ng6154, Ng1579, Ng5567, Ng1752, Ng1917, Ng744, Ng4737, wire4661, Ng6267, Pg16659, Ng1442, Ng5965, Ng4477, Pg10500, Ng4643, Ng5264, Pg14779, Ng2610, Ng5160, Ng5933, Ng1454, Ng753, Ng1296, Ng3151, Ng2980, Ng6727, Ng3530, Ng4104, Ng1532, Pg9251, Ng2177, Ng52, Ng4754, Ng1189, Ng2287, Ng4273, Ng1389, Ng1706, Ng5835, Ng1171, Ng4269, Ng2399, Ng4983, Ng5611, Pg16627, Ng4572, Ng3143, Ng2898, Ng3343, Ng3235, Ng4543, Ng3566, Ng4534, Ng4961, Ng4927, Ng2259, Ng2819, Pg7257, Ng5802, Ng2852, Ng417, Ng681, Ng437, Ng351, Ng5901, Ng2886, Ng3494, Ng5511, Ng3518, Ng1604, Ng5092, Ng4831, Ng4382, Ng6386, Ng479, Ng3965, Ng4749, Ng2008, Ng736, Ng3933, Ng222, Ng3050, Ng1052, Pg17580, Ng2122, Ng2465, Ng5889, Ng4495, Pg8719, Ng4653, Ng3179, Ng1728, Ng2433, Ng3835, Ng6187, Ng4917, Ng1070, Ng822, Pg17715, Ng914, Ng5339, Ng4164, Ng969, Ng2807, Ng4054, Ng6191, Ng5077, Ng5523, Ng3680, Ng6637, Ng174, Ng1682, Ng355, Ng1087, Ng1105, Ng2342, Ng6307, Ng3802, Ng6159, Ng2255, Ng2815, Ng911, Ng43, Pg16775, Ng1748, Ng5551, Ng3558, Ng5499, Ng2960, Ng3901, Ng4888, Ng6251, Pg17649, Ng1373, Pg8215, Ng157, Ng2783, Ng4281, Ng3574, Ng2112, Ng1283, Ng433, Ng4297, Pg14738, Pg13272, Ng758, Ng4639, Ng6537, Ng5543, Pg8475, Ng5961, Ng6243, Ng632, Pg12919, Ng3889, Ng3476, Ng1664, Ng1246, Ng6629, Ng246, Ng4049, Pg7260, Ng2932, Ng4575, Ng4098, Ng4498, Ng528, Ng16, Ng3139, wire4432, Ng4584, Ng142, Pg17639, Ng5831, Ng239, Ng1216, Ng2848, Ng5022, Pg16955, Ng1030, Pg13881, Ng3231, Pg9817, Ng1430, Ng4452, Ng2241, Ng1564, Pg9680, Ng6148, Ng6649, Ng110, Pg14147, Ng225, Ng4486, Ng4504, Ng5873, Ng5037, Ng2319, Ng5495, Pg11770, Ng5208, Ng5579, Ng5869, Ng1589, Ng5752, Ng6279, Ng5917, Ng2975, Ng6167, Pg13966, Ng2599, Ng1448, Pg14125, Ng2370, Ng5164, Ng1333, Ng153, Ng6549, Ng4087, Ng4801, Ng2984, Ng3961, Ng962, Ng101, Pg8918, Ng6625, Ng51, Ng1018, Pg17320, Ng4045, Ng1467, Ng2461, Ng2756, Ng5990, Ng1256, Ng5029, Ng6519, Ng1816, Ng4369, Ng4578, Ng4459, Ng3831, Ng2514, Ng3288, Ng2403, Ng2145, Ng1700, Ng513, Ng2841, Ng5297, Ng2763, Ng4793, Ng952, Ng1263, Ng1950, Ng5138, Ng2307, Ng5109, Pg8398, Ng4664, Ng2223, Ng5808, Ng6645, Ng2016, Ng3873, Pg13926, Ng2315, Ng2811, Ng5957, Ng2047, Ng3869, Pg17760, Ng5575, Ng46, Ng3752, Ng3917, Pg8783, Ng1585, Ng4388, Ng6275, Ng6311, Pg8916, Ng1041, Ng2595, Ng2537, wire4426, Ng4430, Ng4564, Ng4826, Ng6239, Ng232, Ng5268, Ng6545, Ng2417, Ng1772, Ng5052, Pg9615, Ng1890, Ng2629, Ng572, Ng2130, Ng4108, Ng4308, Ng475, Ng990, Ng45, Pg12184, Ng3990, Ng5881, Ng1992, Ng3171, Ng812, Ng832, Ng5897, Ng4571, Pg13895, Ng4455, Ng2902, Ng333, Ng168, Ng2823, Ng3684, Ng3639, Pg14597, Ng3338, Ng5406, Ng269, Ng401, Ng6040, Ng441, Pg9553, Ng3808, Ng10384, Ng3957, Ng4093, Ng1760, Pg12422, Ng160, Ng2279, Ng3498, Ng586, Pg14201, Ng2619, Ng1183, Ng1608, Pg8785, Pg17577, Ng1779, Ng2652, Ng2193, Ng2393, Ng661, Ng4950, Ng5535, Ng2834, Ng1361, Ng6235, Ng1146, Ng2625, Ng150, Ng1696, Ng6555, Pg14189, Ng3881, Ng6621, Ng3470, Ng3897, Ng518, Ng538, Ng2606, Ng1472, Ng542, Ng5188, Ng5689, Pg13259, Ng405, Ng5216, Ng6494, Ng4669, Ng996, Ng4531, Ng2860, Ng4743, Ng6593, Pg8291, Ng4411, Ng1413, Ng26960, Pg13039, Ng6641, Ng1936, Ng55, Ng504, Ng2587, Ng4480, Ng2311, Ng3602, Ng5571, Ng3578, Pg9555, Ng5827, Ng3582, Ng6271, Ng4688, Ng2380, Ng5196, Ng3227, Ng2020, Pg14518, Pg17316, Ng6541, Ng3203, Ng1668, Ng4760, Ng262, Ng1840, Ng5467, Ng460, Ng6209, wire4436, Pg14662, Ng655, Ng3502, Ng2204, Ng5256, Ng4608, Ng794, Pg13906, Ng4423, Ng3689, Ng5685, Ng703, Ng862, Ng3247, Ng2040, Ng4146, Ng4633, Pg7916, Ng4732, Pg9497, Ng5817, Ng2351, Ng2648, Ng6736, Ng4944, Ng4072, Pg7540, Ng4443, Ng3466, Ng4116, Ng5041, Ng4434, Ng3827, Ng6500, Pg17813, Ng3133, Ng3333, Ng979, Ng4681, Ng298, Ng2667, Pg8789, Ng1894, Ng2988, Ng3538, Ng301, Ng341, Ng827, Pg17291, Ng2555, Ng5011, Ng199, Ng6523, Ng1526, Ng4601, Ng854, Ng1484, Ng4922, Ng5080, Ng5863, Ng4581, Ng2518, Ng2567, Ng568, Ng3263, Ng6613, Ng6044, Ng6444, Ng2965, Ng5857, Ng1616, Ng890, Pg17646, Ng3562, Pg10122, Ng1404, Ng3817, Ng93, Ng4501, Ng287, Ng2724, Ng4704, Ng22, Ng2878, Ng5220, Ng617, Pg12368, Ng316, Ng1277, Ng6513, Ng336, Ng2882, Ng933, Ng1906, Ng305, Ng8, Ng2799, Pg14167, Pg17787, Ng4912, Ng4157, Ng2541, Ng2153, Ng550, Ng255, Ng1945, Ng5240, Ng1478, Ng3863, Ng1959, Ng3480, Ng6653, Pg17764, Ng2864, Ng4894, Pg17678, Ng3857, Pg16693, Ng499, Ng1002, Ng776, Ng1236, Ng4646, Ng2476, Ng1657, Ng2375, Ng63, Pg17739, Ng358, Ng896, Ng283, Ng3161, Ng2384, Pg14828, Ng4616, Ng4561, Ng2024, Ng3451, Ng2795, Ng613, Ng4527, Ng1844, Ng5937, Ng4546, Ng2523, Pg11349, Ng2643, Ng1489, Pg8358, Ng2551, Ng5156, wire4421, Pg8279, Pg8839, Ng1955, Ng6049, Ng2273, Pg14749, Ng4771, Ng6098, Ng3147, Ng3347, Ng2269, Ng191, Ng2712, Ng626, Ng2729, Ng5357, Ng4991, Pg17819, Ng4709, Ng2927, Ng4340, Ng5929, Ng4907, Pg16874, Ng4035, Ng2946, Ng918, Ng4082, Pg9743, Ng2036, Ng577, Ng1620, Ng2831, Ng667, Ng930, Ng3937, Ng817, Ng1249, Ng837, Pg16924, Ng599, Ng5475, Ng739, Ng5949, Ng6682, Ng904, Ng2873, Ng1854, Ng5084, Ng5603, Pg8870, Ng2495, Ng2437, Ng2102, Ng2208, Ng2579, Ng4064, Ng4899, Ng2719, Ng4785, Ng5583, Ng781, Ng6173, Pg17743, Ng2917, Ng686, Ng1252, Ng671, Ng2265, Ng6283, Pg14705, Pg17519, Pg8784, Ng5527, Ng4489, Ng1974, Ng1270, Ng4966, Ng6227, Ng3929, Ng5503, Ng4242, Ng5925, Ng1124, Ng4955, Ng5224, Ng2012, Ng6203, Ng5120, Pg17674, Ng2389, Ng4438, Ng2429, Ng2787, Ng1287, Ng2675, wire4507, Ng4836, Ng1199, Pg19357, Ng5547, Ng2138, Pg16744, Ng2338, Pg8919, Ng6247, Ng2791, Ng3949, Ng1291, Ng5945, Ng5244, Ng2759, Ng6741, Ng785, Ng1259, Ng3484, Ng209, Ng6609, Ng5517, Ng2449, Ng2575, Ng65, Ng2715, Ng936, Ng2098, Ng4462, Ng604, Ng6589, Ng1886, Pg17845, Pg17871, Ng429, Ng1870, Ng4249, Ng1825, Ng1008, Ng4392, Ng3546, Ng5236, Ng1768, Ng4854, Ng3925, Ng6509, Ng732, Ng2504, Ng1322, Ng4520, Pg8917, Ng2185, Ng37, Ng4031, Ng2070, wire4658, Ng4176, Pg11418, Ng4405, Ng872, Ng6181, Ng6381, Ng4765, Ng5563, Ng1395, Ng1913, Ng2331, Ng6263, Ng50, Ng3945, Ng347, Ng4473, Ng1266, Ng5489, Ng714, Ng2748, Ng5471, Ng4540, Ng6723, Ng6605, Ng2445, Ng2173, Pg9019, Ng2491, Ng4849, Ng2169, Ng2283, Ng6585, wire4428, Ng2407, Ng2868, Ng2767, Ng1783, Pg16718, Ng1312, Ng5212, Ng4245, Ng645, Ng4291, wire4435, Ng182, Ng1129, Ng2227, Pg8788, Ng2246, Ng1830, Ng3590, Ng392, Ng1592, Ng6505, Ng1221, Ng5921, wire4431, Ng146, Ng218, Ng1932, Ng1624, Ng5062, Ng5462, Ng2689, Ng6573, Ng1677, Ng2028, Ng2671, Pg10527, Pg7243, Ng1848, wire4434, Ng5485, Ng2741, Pg11678, Ng2638, Ng4122, Ng4322, Ng5941, Ng2108, Pg13068, Ng25, Ng1644, Ng595, Ng2217, Ng1319, Ng2066, Ng1152, Ng5252, Ng2165, Ng2571, Ng5176, Pg14673, Ng1211, Ng2827, Pg14217, Ng4859, Ng424, Ng1274, Pg17423, Ng85, Ng2803, Ng1821, Ng2509, Ng5073, Ng1280, wire4651, Pg13085, Ng6633, Ng5124, Pg17400, Ng6303, Ng5069, Ng2994, Ng650, Ng1636, Ng3921, Ng2093, Ng6732, Ng1306, Ng1061, Ng3462, Ng2181, Ng956, Ng1756, Ng5849, Ng4112, Ng2685, Ng2197, Ng2421, Ng1046, Ng482, Ng4401, Ng1514, Ng329, Ng6565, Ng2950, Ng1345, Ng6533, Pg14421, Ng4727, Pg12470, Ng1536, Ng3941, Ng370, Ng5694, Ng1858, Ng446, Ng3219, Ng1811, Ng6601, Ng2441, Ng1874, Ng4349, Ng6581, Ng6597, Ng3610, Ng2890, Ng1978, Ng1612, Ng112, Ng2856, Ng1982, Pg17722, Ng5228, Ng4119, Ng6390, Ng1542, Ng4258, Ng4818, Ng5033, Ng4717, Ng1554, Ng3849, Pg17778, Ng3199, Ng5845, Ng4975, Ng790, Ng5913, Ng1902, Ng6163, Ng4125, Ng4821, Ng4939, Pg19334, Ng3207, Ng4483, Ng3259, Ng5142, Ng5248, Ng2126, Ng3694, Ng5481, Ng1964, Ng5097, Ng3215, Pg16748, Ng111, Ng4427, Ng2779, Pg8786, Pg7245, Ng1720, Ng1367, Ng5112, Ng4145, Ng2161, Ng376, Ng2361, Pg11447, Ng582, Ng2051, Ng1193, Ng2327, Ng907, Ng947, Ng1834, Ng3594, Ng2999, Ng2303, Pg17688, Ng699, Ng723, Ng5703, Ng546, Ng2472, Ng5953, Pg8277, Ng1740, Ng3550, Ng3845, Ng2116, Pg14635, Ng3195, Ng3913, Pg10306, Ng1687, Ng2681, Ng2533, Ng324, Ng2697, Ng4417, Ng6561, Ng1141, Pg12923, Ng2413, Ng1710, Ng6527, Ng3255, Ng1691, Ng2936, Ng5644, Ng5152, Ng5352, Pg8915, Ng2775, Ng2922, Ng1111, Ng5893, Pg16603, Ng6617, Ng2060, Ng4512, Ng5599, Ng3401, Ng4366, Pg16722, wire4433, Ng3129, Ng3329, Ng5170, Ng26959, Ng5821, Ng6299, Pg8416, Ng2079, Ng4698, Ng3703, Ng1559, Ng943, Ng411, Pg9682, Ng3953, Ng2704, Ng6035, Ng1300, Ng4057, Ng5200, Ng4843, Ng5046, Ng2250, Ng26885, Ng4549, Ng2453, Ng5841, Pg14694, Ng2912, Ng2357, Pg8920, Ng164, Ng4253, Ng5016, Ng3119, Ng1351, Ng1648, Ng6972, Ng5115, Ng3352, Ng6657, Ng4552, Ng3893, Ng3211, Pg13049, Pg16624, Ng5595, Ng3614, Ng2894, Ng3125, Pg16686, Ng3821, Ng4141, Ng6974, Ng5272, Ng2735, Ng728, Ng6295, Ng2661, Ng1988, Ng5128, Ng1548, Ng3106, Ng4659, Ng4358, Ng1792, Ng2084, Ng3187, Ng4311, Ng2583, Ng3003, Ng1094, Ng3841, Ng4284, Ng3191, Ng4239, Ng4180, Ng691, Ng534, Ng385, Ng2004, Ng2527, Ng5456, Ng4420, Ng5148, Ng4507, Ng5348, Ng3223, Ng2970, Ng5698, Ng5260, Ng1521, Ng3522, Ng3115, Ng3251, Pg12832, Ng4628, Ng1996, Pg8342, Ng4515, Pg8787, Ng4300, Ng1724, Ng1379, Pg11388, Ng1878, Ng5619, Ng71, wire4437;

always  @(posedge PCLK)
	Ng5057<=Ng33046;

 always  @(posedge PCLK)
	Ng2771<=Ng34441;

 always  @(posedge PCLK)
	Ng1882<=Ng33982;

 always  @(posedge PCLK)
	Ng2299<=Ng34007;

 always  @(posedge PCLK)
	Ng4040<=Ng24276;

 always  @(posedge PCLK)
	Ng2547<=Ng30381;

 always  @(posedge PCLK)
	Ng559<=Pg9048;

 always  @(posedge PCLK)
	Ng3243<=Ng30405;

 always  @(posedge PCLK)
	Ng452<=Ng25604;

 always  @(posedge PCLK)
	Ng3542<=Ng30416;

 always  @(posedge PCLK)
	Ng5232<=Ng30466;

 always  @(posedge PCLK)
	Ng5813<=Ng25736;

 always  @(posedge PCLK)
	Ng2907<=Ng34617;

 always  @(posedge PCLK)
	Ng1744<=Ng33974;

 always  @(posedge PCLK)
	Ng5909<=Ng30505;

 always  @(posedge PCLK)
	Ng1802<=Ng33554;

 always  @(posedge PCLK)
	Ng3554<=Ng30432;

 always  @(posedge PCLK)
	Ng6219<=Ng33064;

 always  @(posedge PCLK)
	Ng807<=Ng34881;

 always  @(posedge PCLK)
	Ng6031<=Pg17715;

 always  @(posedge PCLK)
	Ng847<=Ng24216;

 always  @(posedge PCLK)
	Ng976<=Ng24232;

 always  @(posedge PCLK)
	Ng4172<=Ng34733;

 always  @(posedge PCLK)
	Ng4372<=Ng34882;

 always  @(posedge PCLK)
	Ng3512<=Ng33026;

 always  @(posedge PCLK)
	Ng749<=Ng31867;

 always  @(posedge PCLK)
	Ng3490<=Ng25668;

 always  @(posedge PCLK)
	Pg12350<=Ng24344;

 always  @(posedge PCLK)
	Ng4235<=Pg8920;

 always  @(posedge PCLK)
	Ng1600<=Ng33966;

 always  @(posedge PCLK)
	Ng1714<=Ng33550;

 always  @(posedge PCLK)
	Pg14451<=Pg16656;

 always  @(posedge PCLK)
	Ng3155<=Ng30393;

 always  @(posedge PCLK)
	Ng2236<=Ng29248;

 always  @(posedge PCLK)
	Ng4555<=Ng4571;

 always  @(posedge PCLK)
	Ng3698<=Ng24274;

 always  @(posedge PCLK)
	Ng1736<=Ng33973;

 always  @(posedge PCLK)
	Ng1968<=Ng30360;

 always  @(posedge PCLK)
	Ng4621<=Ng34460;

 always  @(posedge PCLK)
	Ng5607<=Ng30494;

 always  @(posedge PCLK)
	Ng2657<=Ng30384;

 always  @(posedge PCLK)
	Pg12300<=Ng24340;

 always  @(posedge PCLK)
	Ng490<=Ng29223;

 always  @(posedge PCLK)
	Ng311<=Ng26881;

 always  @(posedge PCLK)
	Ng772<=Ng34252;

 always  @(posedge PCLK)
	Ng5587<=Ng30489;

 always  @(posedge PCLK)
	Ng6177<=Ng29301;

 always  @(posedge PCLK)
	Ng6377<=Pg17743;

 always  @(posedge PCLK)
	Ng3167<=Ng33022;

 always  @(posedge PCLK)
	Ng5615<=Ng30496;

 always  @(posedge PCLK)
	Ng4567<=Ng33043;

 always  @(posedge PCLK)
	Ng3457<=Ng29263;

 always  @(posedge PCLK)
	Ng6287<=Ng30533;

 always  @(posedge PCLK)
	Pg7946<=Ng24256;

 always  @(posedge PCLK)
	Ng2563<=Ng34015;

 always  @(posedge PCLK)
	Ng4776<=Ng34031;

 always  @(posedge PCLK)
	Ng4593<=Ng34452;

 always  @(posedge PCLK)
	Ng6199<=Ng34646;

 always  @(posedge PCLK)
	Ng2295<=Ng34001;

 always  @(posedge PCLK)
	Ng1384<=Ng25633;

 always  @(posedge PCLK)
	Ng1339<=Ng24259;

 always  @(posedge PCLK)
	Ng5180<=Ng33049;

 always  @(posedge PCLK)
	Ng2844<=Ng34609;

 always  @(posedge PCLK)
	Ng1024<=Ng31869;

 always  @(posedge PCLK)
	Ng5591<=Ng30490;

 always  @(posedge PCLK)
	Ng3598<=Ng30427;

 always  @(posedge PCLK)
	Ng4264<=Ng21894;

 always  @(posedge PCLK)
	Ng767<=Ng33965;

 always  @(posedge PCLK)
	Ng5853<=Ng34645;

 always  @(posedge PCLK)
	Pg13865<=Pg16874;

 always  @(posedge PCLK)
	Ng2089<=Ng33571;

 always  @(posedge PCLK)
	Ng4933<=Ng34267;

 always  @(posedge PCLK)
	Ng4521<=Ng26971;

 always  @(posedge PCLK)
	Ng5507<=Ng34644;

 always  @(posedge PCLK)
	Pg16656<=Pg16627;

 always  @(posedge PCLK)
	Ng6291<=Ng30534;

 always  @(posedge PCLK)
	Ng294<=Ng33535;

 always  @(posedge PCLK)
	Ng5559<=Ng30498;

 always  @(posedge PCLK)
	Pg9617<=Ng25728;

 always  @(posedge PCLK)
	Pg9741<=Ng25743;

 always  @(posedge PCLK)
	Ng3813<=Ng25684;

 always  @(posedge PCLK)
	Ng562<=Ng25613;

 always  @(posedge PCLK)
	Ng608<=Ng34438;

 always  @(posedge PCLK)
	Ng1205<=Ng24244;

 always  @(posedge PCLK)
	Ng3909<=Ng30439;

 always  @(posedge PCLK)
	Ng6259<=Ng30541;

 always  @(posedge PCLK)
	Ng5905<=Ng30519;

 always  @(posedge PCLK)
	Ng921<=Ng25621;

 always  @(posedge PCLK)
	Ng2955<=Ng34807;

 always  @(posedge PCLK)
	Ng203<=Ng25599;

 always  @(posedge PCLK)
	Ng1099<=Ng24235;

 always  @(posedge PCLK)
	Ng4878<=Ng34036;

 always  @(posedge PCLK)
	Ng5204<=Ng30476;

 always  @(posedge PCLK)
	Pg17604<=Pg17580;

 always  @(posedge PCLK)
	Ng3606<=Ng30429;

 always  @(posedge PCLK)
	Ng1926<=Ng32997;

 always  @(posedge PCLK)
	Ng6215<=Ng33063;

 always  @(posedge PCLK)
	Ng3586<=Ng30424;

 always  @(posedge PCLK)
	Ng291<=Ng32977;

 always  @(posedge PCLK)
	Ng4674<=Ng34026;

 always  @(posedge PCLK)
	Ng3570<=Ng30420;

 always  @(posedge PCLK)
	Pg9048<=Pg12368;

 always  @(posedge PCLK)
	Pg17607<=Pg17739;

 always  @(posedge PCLK)
	Ng1862<=Ng33560;

 always  @(posedge PCLK)
	Ng676<=Ng29226;

 always  @(posedge PCLK)
	Ng843<=Ng25619;

 always  @(posedge PCLK)
	Ng4332<=Ng34455;

 always  @(posedge PCLK)
	Ng4153<=Ng30457;

 always  @(posedge PCLK)
	Pg17711<=Pg14694;

 always  @(posedge PCLK)
	Ng6336<=Ng33625;

 always  @(posedge PCLK)
	Ng622<=Ng34790;

 always  @(posedge PCLK)
	Ng3506<=Ng30414;

 always  @(posedge PCLK)
	Ng4558<=Ng26966;

 always  @(posedge PCLK)
	Pg17685<=Pg17649;

 always  @(posedge PCLK)
	Ng3111<=Ng25656;

 always  @(posedge PCLK)
	wire4430<=Ng30390;

 always  @(posedge PCLK)
	Ng26936<=Ng28079;

 always  @(posedge PCLK)
	Ng939<=Ng34727;

 always  @(posedge PCLK)
	Ng278<=Ng25594;

 always  @(posedge PCLK)
	Ng4492<=Ng26963;

 always  @(posedge PCLK)
	Ng4864<=Ng34034;

 always  @(posedge PCLK)
	Ng1036<=Ng33541;

 always  @(posedge PCLK)
	wire4427<=Ng28093;

 always  @(posedge PCLK)
	Ng1178<=Ng24236;

 always  @(posedge PCLK)
	Ng3239<=Ng30404;

 always  @(posedge PCLK)
	Ng718<=Ng28051;

 always  @(posedge PCLK)
	Ng6195<=Ng29303;

 always  @(posedge PCLK)
	Ng1135<=Ng26917;

 always  @(posedge PCLK)
	Ng6395<=Ng33624;

 always  @(posedge PCLK)
	wire4415<=Ng24337;

 always  @(posedge PCLK)
	Ng554<=Ng34911;

 always  @(posedge PCLK)
	Ng496<=Ng33963;

 always  @(posedge PCLK)
	Ng3853<=Ng34627;

 always  @(posedge PCLK)
	Ng5134<=Ng29282;

 always  @(posedge PCLK)
	Pg17404<=Pg17320;

 always  @(posedge PCLK)
	Pg8344<=Ng25676;

 always  @(posedge PCLK)
	Ng2485<=Ng33013;

 always  @(posedge PCLK)
	Ng925<=Ng32981;

 always  @(posedge PCLK)
	Ng48<=Ng34993;

 always  @(posedge PCLK)
	Ng5555<=Ng30483;

 always  @(posedge PCLK)
	Pg14096<=Pg14217;

 always  @(posedge PCLK)
	Ng1798<=Ng32994;

 always  @(posedge PCLK)
	Ng4076<=Ng28070;

 always  @(posedge PCLK)
	Ng2941<=Ng34806;

 always  @(posedge PCLK)
	Ng3905<=Ng30453;

 always  @(posedge PCLK)
	Ng763<=Ng33539;

 always  @(posedge PCLK)
	Ng6255<=Ng30526;

 always  @(posedge PCLK)
	Ng4375<=Ng26951;

 always  @(posedge PCLK)
	Ng4871<=Ng34035;

 always  @(posedge PCLK)
	Ng4722<=Ng34636;

 always  @(posedge PCLK)
	Ng590<=Ng32978;

 always  @(posedge PCLK)
	Pg13099<=Pg17722;

 always  @(posedge PCLK)
	Ng1632<=Ng30348;

 always  @(posedge PCLK)
	Pg12238<=Ng24336;

 always  @(posedge PCLK)
	Ng3100<=Pg8215;

 always  @(posedge PCLK)
	Ng1495<=Ng24250;

 always  @(posedge PCLK)
	Ng1437<=Ng29236;

 always  @(posedge PCLK)
	Ng6154<=Ng29298;

 always  @(posedge PCLK)
	Ng1579<=Pg10527;

 always  @(posedge PCLK)
	Ng5567<=Ng30499;

 always  @(posedge PCLK)
	Ng1752<=Ng33976;

 always  @(posedge PCLK)
	Ng1917<=Ng32996;

 always  @(posedge PCLK)
	Ng744<=Ng30335;

 always  @(posedge PCLK)
	Ng4737<=Ng34637;

 always  @(posedge PCLK)
	wire4661<=Ng25694;

 always  @(posedge PCLK)
	Ng6267<=Ng30528;

 always  @(posedge PCLK)
	Pg16659<=Pg16775;

 always  @(posedge PCLK)
	Ng1442<=Ng24251;

 always  @(posedge PCLK)
	Ng5965<=Ng30521;

 always  @(posedge PCLK)
	Ng4477<=Ng26960;

 always  @(posedge PCLK)
	Pg10500<=Ng24239;

 always  @(posedge PCLK)
	Ng4643<=Ng34259;

 always  @(posedge PCLK)
	Ng5264<=Ng30474;

 always  @(posedge PCLK)
	Pg14779<=Pg12422;

 always  @(posedge PCLK)
	Ng2610<=Ng33016;

 always  @(posedge PCLK)
	Ng5160<=Ng34643;

 always  @(posedge PCLK)
	Ng5933<=Ng30510;

 always  @(posedge PCLK)
	Ng1454<=Ng29239;

 always  @(posedge PCLK)
	Ng753<=Ng26897;

 always  @(posedge PCLK)
	Ng1296<=Ng34729;

 always  @(posedge PCLK)
	Ng3151<=Ng34625;

 always  @(posedge PCLK)
	Ng2980<=Ng34800;

 always  @(posedge PCLK)
	Ng6727<=Ng24353;

 always  @(posedge PCLK)
	Ng3530<=Ng33029;

 always  @(posedge PCLK)
	Ng4104<=Ng33615;

 always  @(posedge PCLK)
	Ng1532<=Ng24253;

 always  @(posedge PCLK)
	Pg9251<=Ng24281;

 always  @(posedge PCLK)
	Ng2177<=Ng33997;

 always  @(posedge PCLK)
	Ng52<=Ng34997;

 always  @(posedge PCLK)
	Ng4754<=Ng34263;

 always  @(posedge PCLK)
	Ng1189<=Ng24237;

 always  @(posedge PCLK)
	Ng2287<=Ng33584;

 always  @(posedge PCLK)
	Ng4273<=Ng24280;

 always  @(posedge PCLK)
	Ng1389<=Ng26920;

 always  @(posedge PCLK)
	Ng1706<=Ng33548;

 always  @(posedge PCLK)
	Ng5835<=Ng29296;

 always  @(posedge PCLK)
	Ng1171<=Ng30338;

 always  @(posedge PCLK)
	Ng4269<=Ng21895;

 always  @(posedge PCLK)
	Ng2399<=Ng33588;

 always  @(posedge PCLK)
	Ng4983<=Ng34041;

 always  @(posedge PCLK)
	Ng5611<=Ng30495;

 always  @(posedge PCLK)
	Pg16627<=Pg16744;

 always  @(posedge PCLK)
	Ng4572<=Ng29279;

 always  @(posedge PCLK)
	Ng3143<=Ng25655;

 always  @(posedge PCLK)
	Ng2898<=Ng34795;

 always  @(posedge PCLK)
	Ng3343<=Ng24269;

 always  @(posedge PCLK)
	Ng3235<=Ng30403;

 always  @(posedge PCLK)
	Ng4543<=Ng33042;

 always  @(posedge PCLK)
	Ng3566<=Ng30419;

 always  @(posedge PCLK)
	Ng4534<=Ng34023;

 always  @(posedge PCLK)
	Ng4961<=Ng28090;

 always  @(posedge PCLK)
	Ng4927<=Ng34642;

 always  @(posedge PCLK)
	Ng2259<=Ng30370;

 always  @(posedge PCLK)
	Ng2819<=Ng34448;

 always  @(posedge PCLK)
	Pg7257<=Ng26946;

 always  @(posedge PCLK)
	Ng5802<=Pg9617;

 always  @(posedge PCLK)
	Ng2852<=Ng34610;

 always  @(posedge PCLK)
	Ng417<=Ng24209;

 always  @(posedge PCLK)
	Ng681<=Ng28047;

 always  @(posedge PCLK)
	Ng437<=Ng24206;

 always  @(posedge PCLK)
	Ng351<=Ng26891;

 always  @(posedge PCLK)
	Ng5901<=Ng30504;

 always  @(posedge PCLK)
	Ng2886<=Ng34798;

 always  @(posedge PCLK)
	Ng3494<=Ng25669;

 always  @(posedge PCLK)
	Ng5511<=Ng30480;

 always  @(posedge PCLK)
	Ng3518<=Ng33027;

 always  @(posedge PCLK)
	Ng1604<=Ng33972;

 always  @(posedge PCLK)
	Ng5092<=Ng25697;

 always  @(posedge PCLK)
	Ng4831<=Ng28099;

 always  @(posedge PCLK)
	Ng4382<=Ng26947;

 always  @(posedge PCLK)
	Ng6386<=Ng24350;

 always  @(posedge PCLK)
	Ng479<=Ng24210;

 always  @(posedge PCLK)
	Ng3965<=Ng30455;

 always  @(posedge PCLK)
	Ng4749<=Ng28084;

 always  @(posedge PCLK)
	Ng2008<=Ng33993;

 always  @(posedge PCLK)
	Ng736<=Pg11678;

 always  @(posedge PCLK)
	Ng3933<=Ng30444;

 always  @(posedge PCLK)
	Ng222<=Ng33537;

 always  @(posedge PCLK)
	Ng3050<=Ng25650;

 always  @(posedge PCLK)
	Ng1052<=Ng25625;

 always  @(posedge PCLK)
	Pg17580<=Pg17711;

 always  @(posedge PCLK)
	Ng2122<=Ng30366;

 always  @(posedge PCLK)
	Ng2465<=Ng33593;

 always  @(posedge PCLK)
	Ng5889<=Ng30502;

 always  @(posedge PCLK)
	Ng4495<=Ng33036;

 always  @(posedge PCLK)
	Pg8719<=Ng25595;

 always  @(posedge PCLK)
	Ng4653<=Ng34462;

 always  @(posedge PCLK)
	Ng3179<=Ng33024;

 always  @(posedge PCLK)
	Ng1728<=Ng33552;

 always  @(posedge PCLK)
	Ng2433<=Ng34014;

 always  @(posedge PCLK)
	Ng3835<=Ng29273;

 always  @(posedge PCLK)
	Ng6187<=Ng25748;

 always  @(posedge PCLK)
	Ng4917<=Ng34638;

 always  @(posedge PCLK)
	Ng1070<=Ng30341;

 always  @(posedge PCLK)
	Ng822<=Ng26899;

 always  @(posedge PCLK)
	Pg17715<=Pg14673;

 always  @(posedge PCLK)
	Ng914<=Ng30336;

 always  @(posedge PCLK)
	Ng5339<=Pg17639;

 always  @(posedge PCLK)
	Ng4164<=Ng26940;

 always  @(posedge PCLK)
	Ng969<=Ng25622;

 always  @(posedge PCLK)
	Ng2807<=Ng34447;

 always  @(posedge PCLK)
	Ng4054<=Ng33613;

 always  @(posedge PCLK)
	Ng6191<=Ng25749;

 always  @(posedge PCLK)
	Ng5077<=Ng25704;

 always  @(posedge PCLK)
	Ng5523<=Ng33053;

 always  @(posedge PCLK)
	Ng3680<=Pg16722;

 always  @(posedge PCLK)
	Ng6637<=Ng30555;

 always  @(posedge PCLK)
	Ng174<=Ng25601;

 always  @(posedge PCLK)
	Ng1682<=Ng33971;

 always  @(posedge PCLK)
	Ng355<=Ng26892;

 always  @(posedge PCLK)
	Ng1087<=Pg17400;

 always  @(posedge PCLK)
	Ng1105<=Ng26915;

 always  @(posedge PCLK)
	Ng2342<=Ng33008;

 always  @(posedge PCLK)
	Ng6307<=Ng30538;

 always  @(posedge PCLK)
	Ng3802<=Pg8344;

 always  @(posedge PCLK)
	Ng6159<=Ng25750;

 always  @(posedge PCLK)
	Ng2255<=Ng30369;

 always  @(posedge PCLK)
	Ng2815<=Ng34446;

 always  @(posedge PCLK)
	Ng911<=Ng29230;

 always  @(posedge PCLK)
	Ng43<=Ng34789;

 always  @(posedge PCLK)
	Pg16775<=Pg13966;

 always  @(posedge PCLK)
	Ng1748<=Ng33975;

 always  @(posedge PCLK)
	Ng5551<=Ng30497;

 always  @(posedge PCLK)
	Ng3558<=Ng30418;

 always  @(posedge PCLK)
	Ng5499<=Ng25721;

 always  @(posedge PCLK)
	Ng2960<=Ng34622;

 always  @(posedge PCLK)
	Ng3901<=Ng30438;

 always  @(posedge PCLK)
	Ng4888<=Ng34266;

 always  @(posedge PCLK)
	Ng6251<=Ng30540;

 always  @(posedge PCLK)
	Pg17649<=Pg17760;

 always  @(posedge PCLK)
	Ng1373<=Ng32986;

 always  @(posedge PCLK)
	Pg8215<=Ng25648;

 always  @(posedge PCLK)
	Ng157<=Ng33960;

 always  @(posedge PCLK)
	Ng2783<=Ng34442;

 always  @(posedge PCLK)
	Ng4281<=Pg8839;

 always  @(posedge PCLK)
	Ng3574<=Ng30421;

 always  @(posedge PCLK)
	Ng2112<=Ng33573;

 always  @(posedge PCLK)
	Ng1283<=Ng34730;

 always  @(posedge PCLK)
	Ng433<=Ng24205;

 always  @(posedge PCLK)
	Ng4297<=Pg10122;

 always  @(posedge PCLK)
	Pg14738<=Pg12350;

 always  @(posedge PCLK)
	Pg13272<=Pg19357;

 always  @(posedge PCLK)
	Ng758<=Ng32979;

 always  @(posedge PCLK)
	Ng4639<=Ng34025;

 always  @(posedge PCLK)
	Ng6537<=Ng25763;

 always  @(posedge PCLK)
	Ng5543<=Ng30481;

 always  @(posedge PCLK)
	Pg8475<=Pg7946;

 always  @(posedge PCLK)
	Ng5961<=Ng30517;

 always  @(posedge PCLK)
	Ng6243<=Ng30539;

 always  @(posedge PCLK)
	Ng632<=Ng34880;

 always  @(posedge PCLK)
	Pg12919<=Ng24242;

 always  @(posedge PCLK)
	Ng3889<=Ng30436;

 always  @(posedge PCLK)
	Ng3476<=Ng29265;

 always  @(posedge PCLK)
	Ng1664<=Ng32990;

 always  @(posedge PCLK)
	Ng1246<=Ng24245;

 always  @(posedge PCLK)
	Ng6629<=Ng30553;

 always  @(posedge PCLK)
	Ng246<=Ng26907;

 always  @(posedge PCLK)
	Ng4049<=Ng24278;

 always  @(posedge PCLK)
	Pg7260<=Ng26955;

 always  @(posedge PCLK)
	Ng2932<=Ng24282;

 always  @(posedge PCLK)
	Ng4575<=Ng29276;

 always  @(posedge PCLK)
	Ng4098<=Ng31894;

 always  @(posedge PCLK)
	Ng4498<=Ng33037;

 always  @(posedge PCLK)
	Ng528<=Ng26894;

 always  @(posedge PCLK)
	Ng16<=Ng34994;

 always  @(posedge PCLK)
	Ng3139<=Ng25654;

 always  @(posedge PCLK)
	wire4432<=Ng33962;

 always  @(posedge PCLK)
	Ng4584<=Ng34451;

 always  @(posedge PCLK)
	Ng142<=Ng34250;

 always  @(posedge PCLK)
	Pg17639<=Pg14597;

 always  @(posedge PCLK)
	Ng5831<=Ng29295;

 always  @(posedge PCLK)
	Ng239<=Ng26905;

 always  @(posedge PCLK)
	Ng1216<=Ng25629;

 always  @(posedge PCLK)
	Ng2848<=Ng34792;

 always  @(posedge PCLK)
	Ng5022<=Ng25703;

 always  @(posedge PCLK)
	Pg16955<=Pg14518;

 always  @(posedge PCLK)
	Ng1030<=Ng32983;

 always  @(posedge PCLK)
	Pg13881<=Pg16924;

 always  @(posedge PCLK)
	Ng3231<=Ng30402;

 always  @(posedge PCLK)
	Pg9817<=Ng25757;

 always  @(posedge PCLK)
	Ng1430<=Pg17423;

 always  @(posedge PCLK)
	Ng4452<=Pg7245;

 always  @(posedge PCLK)
	Ng2241<=Ng33999;

 always  @(posedge PCLK)
	Ng1564<=Ng24262;

 always  @(posedge PCLK)
	Pg9680<=Ng25729;

 always  @(posedge PCLK)
	Ng6148<=Pg9682;

 always  @(posedge PCLK)
	Ng6649<=Ng30558;

 always  @(posedge PCLK)
	Ng110<=Ng34848;

 always  @(posedge PCLK)
	Pg14147<=Pg14125;

 always  @(posedge PCLK)
	Ng225<=Ng26901;

 always  @(posedge PCLK)
	Ng4486<=Ng26961;

 always  @(posedge PCLK)
	Ng4504<=Ng33039;

 always  @(posedge PCLK)
	Ng5873<=Ng33059;

 always  @(posedge PCLK)
	Ng5037<=Ng31899;

 always  @(posedge PCLK)
	Ng2319<=Ng33007;

 always  @(posedge PCLK)
	Ng5495<=Ng25720;

 always  @(posedge PCLK)
	Pg11770<=Ng21891;

 always  @(posedge PCLK)
	Ng5208<=Ng30462;

 always  @(posedge PCLK)
	Ng5579<=Ng30487;

 always  @(posedge PCLK)
	Ng5869<=Ng33058;

 always  @(posedge PCLK)
	Ng1589<=Ng24261;

 always  @(posedge PCLK)
	Ng5752<=Ng25730;

 always  @(posedge PCLK)
	Ng6279<=Ng30531;

 always  @(posedge PCLK)
	Ng5917<=Ng30506;

 always  @(posedge PCLK)
	Ng2975<=Ng34804;

 always  @(posedge PCLK)
	Ng6167<=Ng25747;

 always  @(posedge PCLK)
	Pg13966<=Pg11418;

 always  @(posedge PCLK)
	Ng2599<=Ng33601;

 always  @(posedge PCLK)
	Ng1448<=Ng26922;

 always  @(posedge PCLK)
	Pg14125<=Pg14096;

 always  @(posedge PCLK)
	Ng2370<=Ng29250;

 always  @(posedge PCLK)
	Ng5164<=Ng30459;

 always  @(posedge PCLK)
	Ng1333<=Pg8475;

 always  @(posedge PCLK)
	Ng153<=Ng33534;

 always  @(posedge PCLK)
	Ng6549<=Ng30543;

 always  @(posedge PCLK)
	Ng4087<=Ng29275;

 always  @(posedge PCLK)
	Ng4801<=Ng34030;

 always  @(posedge PCLK)
	Ng2984<=Ng34980;

 always  @(posedge PCLK)
	Ng3961<=Ng30451;

 always  @(posedge PCLK)
	Ng962<=Ng25627;

 always  @(posedge PCLK)
	Ng101<=Ng34787;

 always  @(posedge PCLK)
	Pg8918<=Pg8870;

 always  @(posedge PCLK)
	Ng6625<=Ng30552;

 always  @(posedge PCLK)
	Ng51<=Ng34996;

 always  @(posedge PCLK)
	Ng1018<=Ng30337;

 always  @(posedge PCLK)
	Pg17320<=Ng24254;

 always  @(posedge PCLK)
	Ng4045<=Ng24277;

 always  @(posedge PCLK)
	Ng1467<=Ng29237;

 always  @(posedge PCLK)
	Ng2461<=Ng30378;

 always  @(posedge PCLK)
	Ng2756<=Ng33019;

 always  @(posedge PCLK)
	Ng5990<=Ng33623;

 always  @(posedge PCLK)
	Ng1256<=Ng29235;

 always  @(posedge PCLK)
	Ng5029<=Ng31902;

 always  @(posedge PCLK)
	Ng6519<=Ng29306;

 always  @(posedge PCLK)
	Ng1816<=Ng33978;

 always  @(posedge PCLK)
	Ng4369<=Ng26970;

 always  @(posedge PCLK)
	Ng4578<=Ng29278;

 always  @(posedge PCLK)
	Ng4459<=Ng34253;

 always  @(posedge PCLK)
	Ng3831<=Ng29272;

 always  @(posedge PCLK)
	Ng2514<=Ng33595;

 always  @(posedge PCLK)
	Ng3288<=Ng33610;

 always  @(posedge PCLK)
	Ng2403<=Ng33589;

 always  @(posedge PCLK)
	Ng2145<=Ng34605;

 always  @(posedge PCLK)
	Ng1700<=Ng30350;

 always  @(posedge PCLK)
	Ng513<=Ng25611;

 always  @(posedge PCLK)
	Ng2841<=Ng26936;

 always  @(posedge PCLK)
	Ng5297<=Ng33619;

 always  @(posedge PCLK)
	Ng2763<=Ng34022;

 always  @(posedge PCLK)
	Ng4793<=Ng34033;

 always  @(posedge PCLK)
	Ng952<=Ng34726;

 always  @(posedge PCLK)
	Ng1263<=Ng31870;

 always  @(posedge PCLK)
	Ng1950<=Ng33985;

 always  @(posedge PCLK)
	Ng5138<=Ng29283;

 always  @(posedge PCLK)
	Ng2307<=Ng34003;

 always  @(posedge PCLK)
	Ng5109<=Pg9497;

 always  @(posedge PCLK)
	Pg8398<=Ng25677;

 always  @(posedge PCLK)
	Ng4664<=Ng34463;

 always  @(posedge PCLK)
	Ng2223<=Ng33006;

 always  @(posedge PCLK)
	Ng5808<=Ng29292;

 always  @(posedge PCLK)
	Ng6645<=Ng30557;

 always  @(posedge PCLK)
	Ng2016<=Ng33989;

 always  @(posedge PCLK)
	Ng3873<=Ng33033;

 always  @(posedge PCLK)
	Pg13926<=Pg11388;

 always  @(posedge PCLK)
	Ng2315<=Ng34005;

 always  @(posedge PCLK)
	Ng2811<=Ng26932;

 always  @(posedge PCLK)
	Ng5957<=Ng30516;

 always  @(posedge PCLK)
	Ng2047<=Ng33575;

 always  @(posedge PCLK)
	Ng3869<=Ng33032;

 always  @(posedge PCLK)
	Pg17760<=Pg14779;

 always  @(posedge PCLK)
	Ng5575<=Ng30486;

 always  @(posedge PCLK)
	Ng46<=Ng34991;

 always  @(posedge PCLK)
	Ng3752<=Ng25678;

 always  @(posedge PCLK)
	Ng3917<=Ng30440;

 always  @(posedge PCLK)
	Pg8783<=Pg11447;

 always  @(posedge PCLK)
	Ng1585<=Pg12923;

 always  @(posedge PCLK)
	Ng4388<=Ng26949;

 always  @(posedge PCLK)
	Ng6275<=Ng30530;

 always  @(posedge PCLK)
	Ng6311<=Ng30542;

 always  @(posedge PCLK)
	Pg8916<=Pg8915;

 always  @(posedge PCLK)
	Ng1041<=Ng25624;

 always  @(posedge PCLK)
	Ng2595<=Ng30383;

 always  @(posedge PCLK)
	Ng2537<=Ng33597;

 always  @(posedge PCLK)
	wire4426<=Ng34598;

 always  @(posedge PCLK)
	Ng4430<=Ng26957;

 always  @(posedge PCLK)
	Ng4564<=Ng26967;

 always  @(posedge PCLK)
	Ng4826<=Ng28102;

 always  @(posedge PCLK)
	Ng6239<=Ng30524;

 always  @(posedge PCLK)
	Ng232<=Ng26903;

 always  @(posedge PCLK)
	Ng5268<=Ng30475;

 always  @(posedge PCLK)
	Ng6545<=Ng34647;

 always  @(posedge PCLK)
	Ng2417<=Ng30377;

 always  @(posedge PCLK)
	Ng1772<=Ng33553;

 always  @(posedge PCLK)
	Ng5052<=Ng31903;

 always  @(posedge PCLK)
	Pg9615<=Ng25715;

 always  @(posedge PCLK)
	Ng1890<=Ng33984;

 always  @(posedge PCLK)
	Ng2629<=Ng33602;

 always  @(posedge PCLK)
	Ng572<=Ng28045;

 always  @(posedge PCLK)
	Ng2130<=Ng34603;

 always  @(posedge PCLK)
	Ng4108<=Ng33035;

 always  @(posedge PCLK)
	Ng4308<=Pg9251;

 always  @(posedge PCLK)
	Ng475<=Ng24208;

 always  @(posedge PCLK)
	Ng990<=Pg8416;

 always  @(posedge PCLK)
	Ng45<=Ng34990;

 always  @(posedge PCLK)
	Pg12184<=Ng24213;

 always  @(posedge PCLK)
	Ng3990<=Ng33614;

 always  @(posedge PCLK)
	Ng5881<=Ng33060;

 always  @(posedge PCLK)
	Ng1992<=Ng30362;

 always  @(posedge PCLK)
	Ng3171<=Ng33023;

 always  @(posedge PCLK)
	Ng812<=Ng26898;

 always  @(posedge PCLK)
	Ng832<=Ng25618;

 always  @(posedge PCLK)
	Ng5897<=Ng30518;

 always  @(posedge PCLK)
	Ng4571<=Ng6974;

 always  @(posedge PCLK)
	Pg13895<=Pg11349;

 always  @(posedge PCLK)
	Ng4455<=Ng26959;

 always  @(posedge PCLK)
	Ng2902<=Ng34801;

 always  @(posedge PCLK)
	Ng333<=Ng26884;

 always  @(posedge PCLK)
	Ng168<=Ng25600;

 always  @(posedge PCLK)
	Ng2823<=Ng26933;

 always  @(posedge PCLK)
	Ng3684<=Ng28066;

 always  @(posedge PCLK)
	Ng3639<=Ng33612;

 always  @(posedge PCLK)
	Pg14597<=Pg17787;

 always  @(posedge PCLK)
	Ng3338<=Ng24268;

 always  @(posedge PCLK)
	Ng5406<=Ng25716;

 always  @(posedge PCLK)
	Ng269<=Ng26906;

 always  @(posedge PCLK)
	Ng401<=Ng24203;

 always  @(posedge PCLK)
	Ng6040<=Ng24346;

 always  @(posedge PCLK)
	Ng441<=Ng24207;

 always  @(posedge PCLK)
	Pg9553<=Ng25701;

 always  @(posedge PCLK)
	Ng3808<=Ng29269;

 always  @(posedge PCLK)
	Ng10384<=Ng34255;

 always  @(posedge PCLK)
	Ng3957<=Ng30450;

 always  @(posedge PCLK)
	Ng4093<=Ng30456;

 always  @(posedge PCLK)
	Ng1760<=Ng32991;

 always  @(posedge PCLK)
	Pg12422<=Ng24348;

 always  @(posedge PCLK)
	Ng160<=Ng34249;

 always  @(posedge PCLK)
	Ng2279<=Ng30371;

 always  @(posedge PCLK)
	Ng3498<=Ng29268;

 always  @(posedge PCLK)
	Ng586<=Ng29224;

 always  @(posedge PCLK)
	Pg14201<=Pg14189;

 always  @(posedge PCLK)
	Ng2619<=Ng33017;

 always  @(posedge PCLK)
	Ng1183<=Ng30339;

 always  @(posedge PCLK)
	Ng1608<=Ng33967;

 always  @(posedge PCLK)
	Pg8785<=Pg8784;

 always  @(posedge PCLK)
	Pg17577<=Pg17519;

 always  @(posedge PCLK)
	Ng1779<=Ng33559;

 always  @(posedge PCLK)
	Ng2652<=Ng29255;

 always  @(posedge PCLK)
	Ng2193<=Ng30368;

 always  @(posedge PCLK)
	Ng2393<=Ng30375;

 always  @(posedge PCLK)
	Ng661<=Ng28052;

 always  @(posedge PCLK)
	Ng4950<=Ng28089;

 always  @(posedge PCLK)
	Ng5535<=Ng33055;

 always  @(posedge PCLK)
	Ng2834<=Ng30392;

 always  @(posedge PCLK)
	Ng1361<=Ng30343;

 always  @(posedge PCLK)
	Ng6235<=Ng30523;

 always  @(posedge PCLK)
	Ng1146<=Ng24233;

 always  @(posedge PCLK)
	Ng2625<=Ng33018;

 always  @(posedge PCLK)
	Ng150<=Ng32976;

 always  @(posedge PCLK)
	Ng1696<=Ng30349;

 always  @(posedge PCLK)
	Ng6555<=Ng33067;

 always  @(posedge PCLK)
	Pg14189<=Ng26900;

 always  @(posedge PCLK)
	Ng3881<=Ng33034;

 always  @(posedge PCLK)
	Ng6621<=Ng30551;

 always  @(posedge PCLK)
	Ng3470<=Ng25667;

 always  @(posedge PCLK)
	Ng3897<=Ng30452;

 always  @(posedge PCLK)
	Ng518<=Ng25612;

 always  @(posedge PCLK)
	Ng538<=Ng34719;

 always  @(posedge PCLK)
	Ng2606<=Ng33607;

 always  @(posedge PCLK)
	Ng1472<=Ng26923;

 always  @(posedge PCLK)
	Ng542<=Ng24211;

 always  @(posedge PCLK)
	Ng5188<=Ng33050;

 always  @(posedge PCLK)
	Ng5689<=Ng24341;

 always  @(posedge PCLK)
	Pg13259<=Pg19334;

 always  @(posedge PCLK)
	Ng405<=Ng24201;

 always  @(posedge PCLK)
	Ng5216<=Ng30463;

 always  @(posedge PCLK)
	Ng6494<=Pg9743;

 always  @(posedge PCLK)
	Ng4669<=Ng34464;

 always  @(posedge PCLK)
	Ng996<=Ng24243;

 always  @(posedge PCLK)
	Ng4531<=Ng24335;

 always  @(posedge PCLK)
	Ng2860<=Ng34611;

 always  @(posedge PCLK)
	Ng4743<=Ng34262;

 always  @(posedge PCLK)
	Ng6593<=Ng30546;

 always  @(posedge PCLK)
	Pg8291<=Ng25591;

 always  @(posedge PCLK)
	Ng4411<=Pg7257;

 always  @(posedge PCLK)
	Ng1413<=Ng30347;

 always  @(posedge PCLK)
	Ng26960<=Ng10384;

 always  @(posedge PCLK)
	Pg13039<=Pg17577;

 always  @(posedge PCLK)
	Ng6641<=Ng30556;

 always  @(posedge PCLK)
	Ng1936<=Ng33562;

 always  @(posedge PCLK)
	Ng55<=Ng35002;

 always  @(posedge PCLK)
	Ng504<=Ng25610;

 always  @(posedge PCLK)
	Ng2587<=Ng33015;

 always  @(posedge PCLK)
	Ng4480<=Ng31896;

 always  @(posedge PCLK)
	Ng2311<=Ng34004;

 always  @(posedge PCLK)
	Ng3602<=Ng30428;

 always  @(posedge PCLK)
	Ng5571<=Ng30485;

 always  @(posedge PCLK)
	Ng3578<=Ng30422;

 always  @(posedge PCLK)
	Pg9555<=Ng25714;

 always  @(posedge PCLK)
	Ng5827<=Ng29294;

 always  @(posedge PCLK)
	Ng3582<=Ng30423;

 always  @(posedge PCLK)
	Ng6271<=Ng30529;

 always  @(posedge PCLK)
	Ng4688<=Ng34028;

 always  @(posedge PCLK)
	Ng2380<=Ng33587;

 always  @(posedge PCLK)
	Ng5196<=Ng30460;

 always  @(posedge PCLK)
	Ng3227<=Ng30401;

 always  @(posedge PCLK)
	Ng2020<=Ng33990;

 always  @(posedge PCLK)
	Pg14518<=Pg16693;

 always  @(posedge PCLK)
	Pg17316<=Pg17291;

 always  @(posedge PCLK)
	Ng6541<=Ng29309;

 always  @(posedge PCLK)
	Ng3203<=Ng30411;

 always  @(posedge PCLK)
	Ng1668<=Ng33546;

 always  @(posedge PCLK)
	Ng4760<=Ng28085;

 always  @(posedge PCLK)
	Ng262<=Ng26904;

 always  @(posedge PCLK)
	Ng1840<=Ng33556;

 always  @(posedge PCLK)
	Ng5467<=Ng25722;

 always  @(posedge PCLK)
	Ng460<=Ng25605;

 always  @(posedge PCLK)
	Ng6209<=Ng33062;

 always  @(posedge PCLK)
	wire4436<=Ng26893;

 always  @(posedge PCLK)
	Pg14662<=Pg12238;

 always  @(posedge PCLK)
	Ng655<=Ng28050;

 always  @(posedge PCLK)
	Ng3502<=Ng34626;

 always  @(posedge PCLK)
	Ng2204<=Ng33583;

 always  @(posedge PCLK)
	Ng5256<=Ng30472;

 always  @(posedge PCLK)
	Ng4608<=Ng34454;

 always  @(posedge PCLK)
	Ng794<=Ng34850;

 always  @(posedge PCLK)
	Pg13906<=Pg16955;

 always  @(posedge PCLK)
	Ng4423<=Pg10306;

 always  @(posedge PCLK)
	Ng3689<=Ng24272;

 always  @(posedge PCLK)
	Ng5685<=Pg17678;

 always  @(posedge PCLK)
	Ng703<=Ng24214;

 always  @(posedge PCLK)
	Ng862<=Ng26909;

 always  @(posedge PCLK)
	Ng3247<=Ng30406;

 always  @(posedge PCLK)
	Ng2040<=Ng33569;

 always  @(posedge PCLK)
	Ng4146<=Ng34628;

 always  @(posedge PCLK)
	Ng4633<=Ng34458;

 always  @(posedge PCLK)
	Pg7916<=Ng24240;

 always  @(posedge PCLK)
	Ng4732<=Ng34634;

 always  @(posedge PCLK)
	Pg9497<=Ng25700;

 always  @(posedge PCLK)
	Ng5817<=Ng29293;

 always  @(posedge PCLK)
	Ng2351<=Ng33009;

 always  @(posedge PCLK)
	Ng2648<=Ng33603;

 always  @(posedge PCLK)
	Ng6736<=Ng24355;

 always  @(posedge PCLK)
	Ng4944<=Ng34268;

 always  @(posedge PCLK)
	Ng4072<=Ng25691;

 always  @(posedge PCLK)
	Pg7540<=Ng26890;

 always  @(posedge PCLK)
	Ng4443<=Pg7260;

 always  @(posedge PCLK)
	Ng3466<=Ng29264;

 always  @(posedge PCLK)
	Ng4116<=Ng28072;

 always  @(posedge PCLK)
	Ng5041<=Ng31900;

 always  @(posedge PCLK)
	Ng4434<=Ng26956;

 always  @(posedge PCLK)
	Ng3827<=Ng29271;

 always  @(posedge PCLK)
	Ng6500<=Ng29304;

 always  @(posedge PCLK)
	Pg17813<=Pg13049;

 always  @(posedge PCLK)
	Ng3133<=Ng29261;

 always  @(posedge PCLK)
	Ng3333<=Ng28063;

 always  @(posedge PCLK)
	Ng979<=Pg13259;

 always  @(posedge PCLK)
	Ng4681<=Ng34027;

 always  @(posedge PCLK)
	Ng298<=Ng33961;

 always  @(posedge PCLK)
	Ng2667<=Ng33604;

 always  @(posedge PCLK)
	Pg8789<=Pg8788;

 always  @(posedge PCLK)
	Ng1894<=Ng32995;

 always  @(posedge PCLK)
	Ng2988<=Ng34624;

 always  @(posedge PCLK)
	Ng3538<=Ng30415;

 always  @(posedge PCLK)
	Ng301<=Ng33536;

 always  @(posedge PCLK)
	Ng341<=Ng26888;

 always  @(posedge PCLK)
	Ng827<=Ng28055;

 always  @(posedge PCLK)
	Pg17291<=Ng24238;

 always  @(posedge PCLK)
	Ng2555<=Ng33600;

 always  @(posedge PCLK)
	Ng5011<=Ng28105;

 always  @(posedge PCLK)
	Ng199<=Ng34721;

 always  @(posedge PCLK)
	Ng6523<=Ng29307;

 always  @(posedge PCLK)
	Ng1526<=Ng30345;

 always  @(posedge PCLK)
	Ng4601<=Ng34453;

 always  @(posedge PCLK)
	Ng854<=Ng32980;

 always  @(posedge PCLK)
	Ng1484<=Ng29238;

 always  @(posedge PCLK)
	Ng4922<=Ng34639;

 always  @(posedge PCLK)
	Ng5080<=Ng25695;

 always  @(posedge PCLK)
	Ng5863<=Ng33057;

 always  @(posedge PCLK)
	Ng4581<=Ng26969;

 always  @(posedge PCLK)
	Ng2518<=Ng29253;

 always  @(posedge PCLK)
	Ng2567<=Ng34021;

 always  @(posedge PCLK)
	Ng568<=Ng26895;

 always  @(posedge PCLK)
	Ng3263<=Ng30413;

 always  @(posedge PCLK)
	Ng6613<=Ng30549;

 always  @(posedge PCLK)
	Ng6044<=Ng24347;

 always  @(posedge PCLK)
	Ng6444<=Ng25758;

 always  @(posedge PCLK)
	Ng2965<=Ng34808;

 always  @(posedge PCLK)
	Ng5857<=Ng30501;

 always  @(posedge PCLK)
	Ng1616<=Ng33969;

 always  @(posedge PCLK)
	Ng890<=Ng34440;

 always  @(posedge PCLK)
	Pg17646<=Pg17607;

 always  @(posedge PCLK)
	Ng3562<=Ng30433;

 always  @(posedge PCLK)
	Pg10122<=Ng21900;

 always  @(posedge PCLK)
	Ng1404<=Ng26921;

 always  @(posedge PCLK)
	Ng3817<=Ng29270;

 always  @(posedge PCLK)
	Ng93<=Ng34878;

 always  @(posedge PCLK)
	Ng4501<=Ng33038;

 always  @(posedge PCLK)
	Ng287<=Ng31865;

 always  @(posedge PCLK)
	Ng2724<=Ng26926;

 always  @(posedge PCLK)
	Ng4704<=Ng28083;

 always  @(posedge PCLK)
	Ng22<=Ng29209;

 always  @(posedge PCLK)
	Ng2878<=Ng34797;

 always  @(posedge PCLK)
	Ng5220<=Ng30478;

 always  @(posedge PCLK)
	Ng617<=Ng34724;

 always  @(posedge PCLK)
	Pg12368<=Ng24212;

 always  @(posedge PCLK)
	Ng316<=Ng26883;

 always  @(posedge PCLK)
	Ng1277<=Ng32985;

 always  @(posedge PCLK)
	Ng6513<=Ng25761;

 always  @(posedge PCLK)
	Ng336<=Ng26886;

 always  @(posedge PCLK)
	Ng2882<=Ng34796;

 always  @(posedge PCLK)
	Ng933<=Ng32982;

 always  @(posedge PCLK)
	Ng1906<=Ng33561;

 always  @(posedge PCLK)
	Ng305<=Ng26880;

 always  @(posedge PCLK)
	Ng8<=Ng34992;

 always  @(posedge PCLK)
	Ng2799<=Ng26931;

 always  @(posedge PCLK)
	Pg14167<=Pg14147;

 always  @(posedge PCLK)
	Pg17787<=Pg13039;

 always  @(posedge PCLK)
	Ng4912<=Ng34641;

 always  @(posedge PCLK)
	Ng4157<=Ng34629;

 always  @(posedge PCLK)
	Ng2541<=Ng33598;

 always  @(posedge PCLK)
	Ng2153<=Ng33576;

 always  @(posedge PCLK)
	Ng550<=Ng34720;

 always  @(posedge PCLK)
	Ng255<=Ng26902;

 always  @(posedge PCLK)
	Ng1945<=Ng29244;

 always  @(posedge PCLK)
	Ng5240<=Ng30468;

 always  @(posedge PCLK)
	Ng1478<=Ng26924;

 always  @(posedge PCLK)
	Ng3863<=Ng33031;

 always  @(posedge PCLK)
	Ng1959<=Ng29245;

 always  @(posedge PCLK)
	Ng3480<=Ng29266;

 always  @(posedge PCLK)
	Ng6653<=Ng30559;

 always  @(posedge PCLK)
	Pg17764<=Pg14749;

 always  @(posedge PCLK)
	Ng2864<=Ng34794;

 always  @(posedge PCLK)
	Ng4894<=Ng28087;

 always  @(posedge PCLK)
	Pg17678<=Pg14635;

 always  @(posedge PCLK)
	Ng3857<=Ng30435;

 always  @(posedge PCLK)
	Pg16693<=Pg16659;

 always  @(posedge PCLK)
	Ng499<=Ng25609;

 always  @(posedge PCLK)
	Ng1002<=Ng28057;

 always  @(posedge PCLK)
	Ng776<=Ng34439;

 always  @(posedge PCLK)
	Ng1236<=Pg10500;

 always  @(posedge PCLK)
	Ng4646<=Ng34260;

 always  @(posedge PCLK)
	Ng2476<=Ng33012;

 always  @(posedge PCLK)
	Ng1657<=Ng32989;

 always  @(posedge PCLK)
	Ng2375<=Ng34006;

 always  @(posedge PCLK)
	Ng63<=Ng34847;

 always  @(posedge PCLK)
	Pg17739<=Pg14738;

 always  @(posedge PCLK)
	Ng358<=Pg8719;

 always  @(posedge PCLK)
	Ng896<=Ng26910;

 always  @(posedge PCLK)
	Ng283<=Ng28043;

 always  @(posedge PCLK)
	Ng3161<=Ng33021;

 always  @(posedge PCLK)
	Ng2384<=Ng29251;

 always  @(posedge PCLK)
	Pg14828<=Pg12470;

 always  @(posedge PCLK)
	Ng4616<=Ng34456;

 always  @(posedge PCLK)
	Ng4561<=Ng26968;

 always  @(posedge PCLK)
	Ng2024<=Ng33991;

 always  @(posedge PCLK)
	Ng3451<=Pg8279;

 always  @(posedge PCLK)
	Ng2795<=Ng26930;

 always  @(posedge PCLK)
	Ng613<=Ng34599;

 always  @(posedge PCLK)
	Ng4527<=Ng28082;

 always  @(posedge PCLK)
	Ng1844<=Ng33557;

 always  @(posedge PCLK)
	Ng5937<=Ng30511;

 always  @(posedge PCLK)
	Ng4546<=Ng33045;

 always  @(posedge PCLK)
	Ng2523<=Ng30379;

 always  @(posedge PCLK)
	Pg11349<=Ng24267;

 always  @(posedge PCLK)
	Ng2643<=Ng34020;

 always  @(posedge PCLK)
	Ng1489<=Ng24249;

 always  @(posedge PCLK)
	Pg8358<=Ng25592;

 always  @(posedge PCLK)
	Ng2551<=Ng30382;

 always  @(posedge PCLK)
	Ng5156<=Ng29285;

 always  @(posedge PCLK)
	wire4421<=Pg12919;

 always  @(posedge PCLK)
	Pg8279<=Ng25662;

 always  @(posedge PCLK)
	Pg8839<=Ng21896;

 always  @(posedge PCLK)
	Ng1955<=Ng33563;

 always  @(posedge PCLK)
	Ng6049<=Ng33622;

 always  @(posedge PCLK)
	Ng2273<=Ng33582;

 always  @(posedge PCLK)
	Pg14749<=Pg17871;

 always  @(posedge PCLK)
	Ng4771<=Ng28086;

 always  @(posedge PCLK)
	Ng6098<=Ng25744;

 always  @(posedge PCLK)
	Ng3147<=Ng29262;

 always  @(posedge PCLK)
	Ng3347<=Ng24270;

 always  @(posedge PCLK)
	Ng2269<=Ng33581;

 always  @(posedge PCLK)
	Ng191<=Pg8358;

 always  @(posedge PCLK)
	Ng2712<=Ng26937;

 always  @(posedge PCLK)
	Ng626<=Ng34849;

 always  @(posedge PCLK)
	Ng2729<=Ng28060;

 always  @(posedge PCLK)
	Ng5357<=Ng33618;

 always  @(posedge PCLK)
	Ng4991<=Ng34038;

 always  @(posedge PCLK)
	Pg17819<=Pg13068;

 always  @(posedge PCLK)
	Ng4709<=Ng34032;

 always  @(posedge PCLK)
	Ng2927<=Ng34803;

 always  @(posedge PCLK)
	Ng4340<=Ng34459;

 always  @(posedge PCLK)
	Ng5929<=Ng30509;

 always  @(posedge PCLK)
	Ng4907<=Ng34640;

 always  @(posedge PCLK)
	Pg16874<=Pg14421;

 always  @(posedge PCLK)
	Ng4035<=Ng28069;

 always  @(posedge PCLK)
	Ng2946<=Ng21899;

 always  @(posedge PCLK)
	Ng918<=Ng31868;

 always  @(posedge PCLK)
	Ng4082<=Ng26938;

 always  @(posedge PCLK)
	Pg9743<=Ng25756;

 always  @(posedge PCLK)
	Ng2036<=Ng30363;

 always  @(posedge PCLK)
	Ng577<=Ng30334;

 always  @(posedge PCLK)
	Ng1620<=Ng33970;

 always  @(posedge PCLK)
	Ng2831<=Ng30391;

 always  @(posedge PCLK)
	Ng667<=Ng25615;

 always  @(posedge PCLK)
	Ng930<=Ng33540;

 always  @(posedge PCLK)
	Ng3937<=Ng30445;

 always  @(posedge PCLK)
	Ng817<=Ng25617;

 always  @(posedge PCLK)
	Ng1249<=Ng24247;

 always  @(posedge PCLK)
	Ng837<=Ng24215;

 always  @(posedge PCLK)
	Pg16924<=Pg14451;

 always  @(posedge PCLK)
	Ng599<=Ng33964;

 always  @(posedge PCLK)
	Ng5475<=Ng25719;

 always  @(posedge PCLK)
	Ng739<=Ng29228;

 always  @(posedge PCLK)
	Ng5949<=Ng30514;

 always  @(posedge PCLK)
	Ng6682<=Ng33627;

 always  @(posedge PCLK)
	Ng904<=Ng24231;

 always  @(posedge PCLK)
	Ng2873<=Ng34615;

 always  @(posedge PCLK)
	Ng1854<=Ng30356;

 always  @(posedge PCLK)
	Ng5084<=Ng25696;

 always  @(posedge PCLK)
	Ng5603<=Ng30493;

 always  @(posedge PCLK)
	Pg8870<=Pg8917;

 always  @(posedge PCLK)
	Ng2495<=Ng33594;

 always  @(posedge PCLK)
	Ng2437<=Ng34009;

 always  @(posedge PCLK)
	Ng2102<=Ng30365;

 always  @(posedge PCLK)
	Ng2208<=Ng33004;

 always  @(posedge PCLK)
	Ng2579<=Ng34018;

 always  @(posedge PCLK)
	Ng4064<=Ng25685;

 always  @(posedge PCLK)
	Ng4899<=Ng34040;

 always  @(posedge PCLK)
	Ng2719<=Ng25639;

 always  @(posedge PCLK)
	Ng4785<=Ng34029;

 always  @(posedge PCLK)
	Ng5583<=Ng30488;

 always  @(posedge PCLK)
	Ng781<=Ng34600;

 always  @(posedge PCLK)
	Ng6173<=Ng29300;

 always  @(posedge PCLK)
	Pg17743<=Pg14705;

 always  @(posedge PCLK)
	Ng2917<=Ng34802;

 always  @(posedge PCLK)
	Ng686<=Ng25614;

 always  @(posedge PCLK)
	Ng1252<=Ng28058;

 always  @(posedge PCLK)
	Ng671<=Ng29225;

 always  @(posedge PCLK)
	Ng2265<=Ng33580;

 always  @(posedge PCLK)
	Ng6283<=Ng30532;

 always  @(posedge PCLK)
	Pg14705<=Pg17845;

 always  @(posedge PCLK)
	Pg17519<=Pg17674;

 always  @(posedge PCLK)
	Pg8784<=Pg8783;

 always  @(posedge PCLK)
	Ng5527<=Ng33054;

 always  @(posedge PCLK)
	Ng4489<=Ng26962;

 always  @(posedge PCLK)
	Ng1974<=Ng33564;

 always  @(posedge PCLK)
	Ng1270<=Ng32984;

 always  @(posedge PCLK)
	Ng4966<=Ng34039;

 always  @(posedge PCLK)
	Ng6227<=Ng33065;

 always  @(posedge PCLK)
	Ng3929<=Ng30443;

 always  @(posedge PCLK)
	Ng5503<=Ng29291;

 always  @(posedge PCLK)
	Ng4242<=Ng24279;

 always  @(posedge PCLK)
	Ng5925<=Ng30508;

 always  @(posedge PCLK)
	Ng1124<=Ng29232;

 always  @(posedge PCLK)
	Ng4955<=Ng34269;

 always  @(posedge PCLK)
	Ng5224<=Ng30464;

 always  @(posedge PCLK)
	Ng2012<=Ng33988;

 always  @(posedge PCLK)
	Ng6203<=Ng30522;

 always  @(posedge PCLK)
	Ng5120<=Ng25708;

 always  @(posedge PCLK)
	Pg17674<=Pg14662;

 always  @(posedge PCLK)
	Ng2389<=Ng30374;

 always  @(posedge PCLK)
	Ng4438<=Ng26953;

 always  @(posedge PCLK)
	Ng2429<=Ng34008;

 always  @(posedge PCLK)
	Ng2787<=Ng34444;

 always  @(posedge PCLK)
	Ng1287<=Ng34731;

 always  @(posedge PCLK)
	Ng2675<=Ng33606;

 always  @(posedge PCLK)
	wire4507<=Ng24334;

 always  @(posedge PCLK)
	Ng4836<=Ng34265;

 always  @(posedge PCLK)
	Ng1199<=Ng30340;

 always  @(posedge PCLK)
	Pg19357<=Ng24257;

 always  @(posedge PCLK)
	Ng5547<=Ng30482;

 always  @(posedge PCLK)
	Ng2138<=Ng34604;

 always  @(posedge PCLK)
	Pg16744<=Pg13926;

 always  @(posedge PCLK)
	Ng2338<=Ng33591;

 always  @(posedge PCLK)
	Pg8919<=Pg8918;

 always  @(posedge PCLK)
	Ng6247<=Ng30525;

 always  @(posedge PCLK)
	Ng2791<=Ng26929;

 always  @(posedge PCLK)
	Ng3949<=Ng30448;

 always  @(posedge PCLK)
	Ng1291<=Ng34602;

 always  @(posedge PCLK)
	Ng5945<=Ng30513;

 always  @(posedge PCLK)
	Ng5244<=Ng30469;

 always  @(posedge PCLK)
	Ng2759<=Ng33608;

 always  @(posedge PCLK)
	Ng6741<=Ng33626;

 always  @(posedge PCLK)
	Ng785<=Ng34725;

 always  @(posedge PCLK)
	Ng1259<=Ng30342;

 always  @(posedge PCLK)
	Ng3484<=Ng29267;

 always  @(posedge PCLK)
	Ng209<=Ng25593;

 always  @(posedge PCLK)
	Ng6609<=Ng30548;

 always  @(posedge PCLK)
	Ng5517<=Ng33052;

 always  @(posedge PCLK)
	Ng2449<=Ng34012;

 always  @(posedge PCLK)
	Ng2575<=Ng34017;

 always  @(posedge PCLK)
	Ng65<=wire4507;

 always  @(posedge PCLK)
	Ng2715<=Ng24263;

 always  @(posedge PCLK)
	Ng936<=Ng26912;

 always  @(posedge PCLK)
	Ng2098<=Ng30364;

 always  @(posedge PCLK)
	Ng4462<=Ng34254;

 always  @(posedge PCLK)
	Ng604<=Ng34251;

 always  @(posedge PCLK)
	Ng6589<=Ng30560;

 always  @(posedge PCLK)
	Ng1886<=Ng33983;

 always  @(posedge PCLK)
	Pg17845<=Pg13085;

 always  @(posedge PCLK)
	Pg17871<=Pg13099;

 always  @(posedge PCLK)
	Ng429<=Ng24204;

 always  @(posedge PCLK)
	Ng1870<=Ng33980;

 always  @(posedge PCLK)
	Ng4249<=Ng34631;

 always  @(posedge PCLK)
	Ng1825<=Ng29243;

 always  @(posedge PCLK)
	Ng1008<=Ng25623;

 always  @(posedge PCLK)
	Ng4392<=Ng26950;

 always  @(posedge PCLK)
	Ng3546<=Ng30431;

 always  @(posedge PCLK)
	Ng5236<=Ng30467;

 always  @(posedge PCLK)
	Ng1768<=Ng30353;

 always  @(posedge PCLK)
	Ng4854<=Ng34467;

 always  @(posedge PCLK)
	Ng3925<=Ng30442;

 always  @(posedge PCLK)
	Ng6509<=Ng29305;

 always  @(posedge PCLK)
	Ng732<=Ng25616;

 always  @(posedge PCLK)
	Ng2504<=Ng29252;

 always  @(posedge PCLK)
	Ng1322<=Pg13272;

 always  @(posedge PCLK)
	Ng4520<=Ng6972;

 always  @(posedge PCLK)
	Pg8917<=Pg8916;

 always  @(posedge PCLK)
	Ng2185<=Ng33003;

 always  @(posedge PCLK)
	Ng37<=Ng34613;

 always  @(posedge PCLK)
	Ng4031<=Pg16748;

 always  @(posedge PCLK)
	Ng2070<=Ng33570;

 always  @(posedge PCLK)
	wire4658<=wire4661;

 always  @(posedge PCLK)
	Ng4176<=Ng34734;

 always  @(posedge PCLK)
	Pg11418<=Ng24275;

 always  @(posedge PCLK)
	Ng4405<=Pg7243;

 always  @(posedge PCLK)
	Ng872<=Pg14167;

 always  @(posedge PCLK)
	Ng6181<=Ng29302;

 always  @(posedge PCLK)
	Ng6381<=Ng24349;

 always  @(posedge PCLK)
	Ng4765<=Ng34264;

 always  @(posedge PCLK)
	Ng5563<=Ng30484;

 always  @(posedge PCLK)
	Ng1395<=Ng25634;

 always  @(posedge PCLK)
	Ng1913<=Ng33567;

 always  @(posedge PCLK)
	Ng2331<=Ng33585;

 always  @(posedge PCLK)
	Ng6263<=Ng30527;

 always  @(posedge PCLK)
	Ng50<=Ng34995;

 always  @(posedge PCLK)
	Ng3945<=Ng30447;

 always  @(posedge PCLK)
	Ng347<=Pg7540;

 always  @(posedge PCLK)
	Ng4473<=Ng34256;

 always  @(posedge PCLK)
	Ng1266<=Ng25630;

 always  @(posedge PCLK)
	Ng5489<=Ng29290;

 always  @(posedge PCLK)
	Ng714<=Ng29227;

 always  @(posedge PCLK)
	Ng2748<=Ng31872;

 always  @(posedge PCLK)
	Ng5471<=Ng29287;

 always  @(posedge PCLK)
	Ng4540<=Ng31897;

 always  @(posedge PCLK)
	Ng6723<=Pg17764;

 always  @(posedge PCLK)
	Ng6605<=Ng30562;

 always  @(posedge PCLK)
	Ng2445<=Ng34011;

 always  @(posedge PCLK)
	Ng2173<=Ng33996;

 always  @(posedge PCLK)
	Pg9019<=Ng21898;

 always  @(posedge PCLK)
	Ng2491<=Ng33014;

 always  @(posedge PCLK)
	Ng4849<=Ng34465;

 always  @(posedge PCLK)
	Ng2169<=Ng33995;

 always  @(posedge PCLK)
	Ng2283<=Ng30372;

 always  @(posedge PCLK)
	Ng6585<=Ng30545;

 always  @(posedge PCLK)
	wire4428<=Ng30389;

 always  @(posedge PCLK)
	Ng2407<=Ng33590;

 always  @(posedge PCLK)
	Ng2868<=Ng34616;

 always  @(posedge PCLK)
	Ng2767<=Ng26927;

 always  @(posedge PCLK)
	Ng1783<=Ng32992;

 always  @(posedge PCLK)
	Pg16718<=Pg13895;

 always  @(posedge PCLK)
	Ng1312<=Ng25631;

 always  @(posedge PCLK)
	Ng5212<=Ng30477;

 always  @(posedge PCLK)
	Ng4245<=Ng34632;

 always  @(posedge PCLK)
	Ng645<=Ng28046;

 always  @(posedge PCLK)
	Ng4291<=Pg9019;

 always  @(posedge PCLK)
	wire4435<=Ng26896;

 always  @(posedge PCLK)
	Ng182<=Ng25602;

 always  @(posedge PCLK)
	Ng1129<=Ng26916;

 always  @(posedge PCLK)
	Ng2227<=Ng33578;

 always  @(posedge PCLK)
	Pg8788<=Pg8787;

 always  @(posedge PCLK)
	Ng2246<=Ng33579;

 always  @(posedge PCLK)
	Ng1830<=Ng30354;

 always  @(posedge PCLK)
	Ng3590<=Ng30425;

 always  @(posedge PCLK)
	Ng392<=Ng24200;

 always  @(posedge PCLK)
	Ng1592<=Ng33544;

 always  @(posedge PCLK)
	Ng6505<=Ng25764;

 always  @(posedge PCLK)
	Ng1221<=Ng24246;

 always  @(posedge PCLK)
	Ng5921<=Ng30507;

 always  @(posedge PCLK)
	wire4431<=Ng26889;

 always  @(posedge PCLK)
	Ng146<=Ng30333;

 always  @(posedge PCLK)
	Ng218<=Pg8291;

 always  @(posedge PCLK)
	Ng1932<=Ng32998;

 always  @(posedge PCLK)
	Ng1624<=Ng32987;

 always  @(posedge PCLK)
	Ng5062<=Ng25702;

 always  @(posedge PCLK)
	Ng5462<=Ng29286;

 always  @(posedge PCLK)
	Ng2689<=Ng34606;

 always  @(posedge PCLK)
	Ng6573<=Ng33070;

 always  @(posedge PCLK)
	Ng1677<=Ng29240;

 always  @(posedge PCLK)
	Ng2028<=Ng32999;

 always  @(posedge PCLK)
	Ng2671<=Ng33605;

 always  @(posedge PCLK)
	Pg10527<=Ng24255;

 always  @(posedge PCLK)
	Pg7243<=Ng26945;

 always  @(posedge PCLK)
	Ng1848<=Ng33558;

 always  @(posedge PCLK)
	wire4434<=Ng25699;

 always  @(posedge PCLK)
	Ng5485<=Ng29289;

 always  @(posedge PCLK)
	Ng2741<=Ng30388;

 always  @(posedge PCLK)
	Pg11678<=Pg12184;

 always  @(posedge PCLK)
	Ng2638<=Ng29254;

 always  @(posedge PCLK)
	Ng4122<=Ng28074;

 always  @(posedge PCLK)
	Ng4322<=Ng34450;

 always  @(posedge PCLK)
	Ng5941<=Ng30512;

 always  @(posedge PCLK)
	Ng2108<=Ng33572;

 always  @(posedge PCLK)
	Pg13068<=Pg17646;

 always  @(posedge PCLK)
	Ng25<=Ng25;

 always  @(posedge PCLK)
	Ng1644<=Ng33551;

 always  @(posedge PCLK)
	Ng595<=Ng33538;

 always  @(posedge PCLK)
	Ng2217<=Ng33005;

 always  @(posedge PCLK)
	Ng1319<=Ng24248;

 always  @(posedge PCLK)
	Ng2066<=Ng33002;

 always  @(posedge PCLK)
	Ng1152<=Ng24234;

 always  @(posedge PCLK)
	Ng5252<=Ng30471;

 always  @(posedge PCLK)
	Ng2165<=Ng34000;

 always  @(posedge PCLK)
	Ng2571<=Ng34016;

 always  @(posedge PCLK)
	Ng5176<=Ng33048;

 always  @(posedge PCLK)
	Pg14673<=Pg17819;

 always  @(posedge PCLK)
	Ng1211<=Ng25628;

 always  @(posedge PCLK)
	Ng2827<=Ng26934;

 always  @(posedge PCLK)
	Pg14217<=Pg14201;

 always  @(posedge PCLK)
	Ng4859<=Ng34468;

 always  @(posedge PCLK)
	Ng424<=Ng24202;

 always  @(posedge PCLK)
	Ng1274<=Ng33542;

 always  @(posedge PCLK)
	Pg17423<=Pg17404;

 always  @(posedge PCLK)
	Ng85<=Pg33435;

 always  @(posedge PCLK)
	Ng2803<=Ng34445;

 always  @(posedge PCLK)
	Ng1821<=Ng33555;

 always  @(posedge PCLK)
	Ng2509<=Ng34013;

 always  @(posedge PCLK)
	Ng5073<=Ng28091;

 always  @(posedge PCLK)
	Ng1280<=Ng26919;

 always  @(posedge PCLK)
	wire4651<=wire4658;

 always  @(posedge PCLK)
	Pg13085<=Pg17685;

 always  @(posedge PCLK)
	Ng6633<=Ng30554;

 always  @(posedge PCLK)
	Ng5124<=Ng29281;

 always  @(posedge PCLK)
	Pg17400<=Pg17316;

 always  @(posedge PCLK)
	Ng6303<=Ng30537;

 always  @(posedge PCLK)
	Ng5069<=Ng28092;

 always  @(posedge PCLK)
	Ng2994<=Ng34732;

 always  @(posedge PCLK)
	Ng650<=Ng28049;

 always  @(posedge PCLK)
	Ng1636<=Ng33545;

 always  @(posedge PCLK)
	Ng3921<=Ng30441;

 always  @(posedge PCLK)
	Ng2093<=Ng29247;

 always  @(posedge PCLK)
	Ng6732<=Ng24354;

 always  @(posedge PCLK)
	Ng1306<=Ng25636;

 always  @(posedge PCLK)
	Ng1061<=Ng26914;

 always  @(posedge PCLK)
	Ng3462<=Ng25670;

 always  @(posedge PCLK)
	Ng2181<=Ng33998;

 always  @(posedge PCLK)
	Ng956<=Ng25626;

 always  @(posedge PCLK)
	Ng1756<=Ng33977;

 always  @(posedge PCLK)
	Ng5849<=Ng29297;

 always  @(posedge PCLK)
	Ng4112<=Ng28071;

 always  @(posedge PCLK)
	Ng2685<=Ng30387;

 always  @(posedge PCLK)
	Ng2197<=Ng33577;

 always  @(posedge PCLK)
	Ng2421<=Ng33592;

 always  @(posedge PCLK)
	Ng1046<=Ng26913;

 always  @(posedge PCLK)
	Ng482<=Ng28044;

 always  @(posedge PCLK)
	Ng4401<=Ng26948;

 always  @(posedge PCLK)
	Ng1514<=Ng30344;

 always  @(posedge PCLK)
	Ng329<=Ng26885;

 always  @(posedge PCLK)
	Ng6565<=Ng33069;

 always  @(posedge PCLK)
	Ng2950<=Ng34621;

 always  @(posedge PCLK)
	Ng1345<=Ng28059;

 always  @(posedge PCLK)
	Ng6533<=Ng25762;

 always  @(posedge PCLK)
	Pg14421<=Pg16624;

 always  @(posedge PCLK)
	Ng4727<=Ng34633;

 always  @(posedge PCLK)
	Pg12470<=Ng24352;

 always  @(posedge PCLK)
	Ng1536<=Ng26925;

 always  @(posedge PCLK)
	Ng3941<=Ng30446;

 always  @(posedge PCLK)
	Ng370<=Ng25597;

 always  @(posedge PCLK)
	Ng5694<=Ng24342;

 always  @(posedge PCLK)
	Ng1858<=Ng30357;

 always  @(posedge PCLK)
	Ng446<=Ng26908;

 always  @(posedge PCLK)
	Ng3219<=Ng30399;

 always  @(posedge PCLK)
	Ng1811<=Ng29242;

 always  @(posedge PCLK)
	Ng6601<=Ng30547;

 always  @(posedge PCLK)
	Ng2441<=Ng34010;

 always  @(posedge PCLK)
	Ng1874<=Ng33986;

 always  @(posedge PCLK)
	Ng4349<=Ng34257;

 always  @(posedge PCLK)
	Ng6581<=Ng30544;

 always  @(posedge PCLK)
	Ng6597<=Ng30561;

 always  @(posedge PCLK)
	Ng3610<=Ng30430;

 always  @(posedge PCLK)
	Ng2890<=Ng34799;

 always  @(posedge PCLK)
	Ng1978<=Ng33565;

 always  @(posedge PCLK)
	Ng1612<=Ng33968;

 always  @(posedge PCLK)
	Ng112<=Ng34879;

 always  @(posedge PCLK)
	Ng2856<=Ng34793;

 always  @(posedge PCLK)
	Ng1982<=Ng33566;

 always  @(posedge PCLK)
	Pg17722<=Pg17688;

 always  @(posedge PCLK)
	Ng5228<=Ng30465;

 always  @(posedge PCLK)
	Ng4119<=Ng28073;

 always  @(posedge PCLK)
	Ng6390<=Ng24351;

 always  @(posedge PCLK)
	Ng1542<=Ng30346;

 always  @(posedge PCLK)
	Ng4258<=Ng21893;

 always  @(posedge PCLK)
	Ng4818<=wire4651;

 always  @(posedge PCLK)
	Ng5033<=Ng31904;

 always  @(posedge PCLK)
	Ng4717<=Ng34635;

 always  @(posedge PCLK)
	Ng1554<=Ng25637;

 always  @(posedge PCLK)
	Ng3849<=Ng29274;

 always  @(posedge PCLK)
	Pg17778<=Pg14828;

 always  @(posedge PCLK)
	Ng3199<=Ng30396;

 always  @(posedge PCLK)
	Ng5845<=Ng25735;

 always  @(posedge PCLK)
	Ng4975<=Ng34037;

 always  @(posedge PCLK)
	Ng790<=Ng34791;

 always  @(posedge PCLK)
	Ng5913<=Ng30520;

 always  @(posedge PCLK)
	Ng1902<=Ng30358;

 always  @(posedge PCLK)
	Ng6163<=Ng29299;

 always  @(posedge PCLK)
	Ng4125<=Ng28081;

 always  @(posedge PCLK)
	Ng4821<=Ng28096;

 always  @(posedge PCLK)
	Ng4939<=Ng28088;

 always  @(posedge PCLK)
	Pg19334<=Ng24241;

 always  @(posedge PCLK)
	Ng3207<=Ng30397;

 always  @(posedge PCLK)
	Ng4483<=Ng4520;

 always  @(posedge PCLK)
	Ng3259<=Ng30409;

 always  @(posedge PCLK)
	Ng5142<=Ng29284;

 always  @(posedge PCLK)
	Ng5248<=Ng30470;

 always  @(posedge PCLK)
	Ng2126<=Ng30367;

 always  @(posedge PCLK)
	Ng3694<=Ng24273;

 always  @(posedge PCLK)
	Ng5481<=Ng29288;

 always  @(posedge PCLK)
	Ng1964<=Ng30359;

 always  @(posedge PCLK)
	Ng5097<=Ng25698;

 always  @(posedge PCLK)
	Ng3215<=Ng30398;

 always  @(posedge PCLK)
	Pg16748<=Pg13906;

 always  @(posedge PCLK)
	Ng111<=Pg33079;

 always  @(posedge PCLK)
	Ng4427<=Ng26952;

 always  @(posedge PCLK)
	Ng2779<=Ng26928;

 always  @(posedge PCLK)
	Pg8786<=Pg8785;

 always  @(posedge PCLK)
	Pg7245<=Ng26954;

 always  @(posedge PCLK)
	Ng1720<=Ng30351;

 always  @(posedge PCLK)
	Ng1367<=Ng31871;

 always  @(posedge PCLK)
	Ng5112<=Pg9553;

 always  @(posedge PCLK)
	Ng4145<=Ng26939;

 always  @(posedge PCLK)
	Ng2161<=Ng33994;

 always  @(posedge PCLK)
	Ng376<=Ng25596;

 always  @(posedge PCLK)
	Ng2361<=Ng33586;

 always  @(posedge PCLK)
	Pg11447<=Ng21901;

 always  @(posedge PCLK)
	Ng582<=Ng31866;

 always  @(posedge PCLK)
	Ng2051<=Ng33000;

 always  @(posedge PCLK)
	Ng1193<=Ng26918;

 always  @(posedge PCLK)
	Ng2327<=Ng30373;

 always  @(posedge PCLK)
	Ng907<=Ng28056;

 always  @(posedge PCLK)
	Ng947<=Ng34601;

 always  @(posedge PCLK)
	Ng1834<=Ng30355;

 always  @(posedge PCLK)
	Ng3594<=Ng30426;

 always  @(posedge PCLK)
	Ng2999<=Ng34805;

 always  @(posedge PCLK)
	Ng2303<=Ng34002;

 always  @(posedge PCLK)
	Pg17688<=Pg17778;

 always  @(posedge PCLK)
	Ng699<=Ng28053;

 always  @(posedge PCLK)
	Ng723<=Ng29229;

 always  @(posedge PCLK)
	Ng5703<=Ng33620;

 always  @(posedge PCLK)
	Ng546<=Ng34722;

 always  @(posedge PCLK)
	Ng2472<=Ng33599;

 always  @(posedge PCLK)
	Ng5953<=Ng30515;

 always  @(posedge PCLK)
	Pg8277<=Ng25649;

 always  @(posedge PCLK)
	Ng1740<=Ng33979;

 always  @(posedge PCLK)
	Ng3550<=Ng30417;

 always  @(posedge PCLK)
	Ng3845<=Ng25683;

 always  @(posedge PCLK)
	Ng2116<=Ng33574;

 always  @(posedge PCLK)
	Pg14635<=Pg17813;

 always  @(posedge PCLK)
	Ng3195<=Ng30410;

 always  @(posedge PCLK)
	Ng3913<=Ng30454;

 always  @(posedge PCLK)
	Pg10306<=Ng34024;

 always  @(posedge PCLK)
	Ng1687<=Ng33547;

 always  @(posedge PCLK)
	Ng2681<=Ng30386;

 always  @(posedge PCLK)
	Ng2533<=Ng33596;

 always  @(posedge PCLK)
	Ng324<=Ng26887;

 always  @(posedge PCLK)
	Ng2697<=Ng34607;

 always  @(posedge PCLK)
	Ng4417<=Ng31895;

 always  @(posedge PCLK)
	Ng6561<=Ng33068;

 always  @(posedge PCLK)
	Ng1141<=Ng29233;

 always  @(posedge PCLK)
	Pg12923<=Ng24258;

 always  @(posedge PCLK)
	Ng2413<=Ng30376;

 always  @(posedge PCLK)
	Ng1710<=Ng33549;

 always  @(posedge PCLK)
	Ng6527<=Ng29308;

 always  @(posedge PCLK)
	Ng3255<=Ng30408;

 always  @(posedge PCLK)
	Ng1691<=Ng29241;

 always  @(posedge PCLK)
	Ng2936<=Ng34620;

 always  @(posedge PCLK)
	Ng5644<=Ng33621;

 always  @(posedge PCLK)
	Ng5152<=Ng25707;

 always  @(posedge PCLK)
	Ng5352<=Ng24339;

 always  @(posedge PCLK)
	Pg8915<=Pg11770;

 always  @(posedge PCLK)
	Ng2775<=Ng34443;

 always  @(posedge PCLK)
	Ng2922<=Ng34619;

 always  @(posedge PCLK)
	Ng1111<=Ng29234;

 always  @(posedge PCLK)
	Ng5893<=Ng30503;

 always  @(posedge PCLK)
	Pg16603<=Pg16718;

 always  @(posedge PCLK)
	Ng6617<=Ng30550;

 always  @(posedge PCLK)
	Ng2060<=Ng33001;

 always  @(posedge PCLK)
	Ng4512<=Ng33040;

 always  @(posedge PCLK)
	Ng5599<=Ng30492;

 always  @(posedge PCLK)
	Ng3401<=Ng25664;

 always  @(posedge PCLK)
	Ng4366<=Ng26944;

 always  @(posedge PCLK)
	Pg16722<=Pg13881;

 always  @(posedge PCLK)
	wire4433<=Ng34614;

 always  @(posedge PCLK)
	Ng3129<=Ng29260;

 always  @(posedge PCLK)
	Ng3329<=Pg16686;

 always  @(posedge PCLK)
	Ng5170<=Ng33047;

 always  @(posedge PCLK)
	Ng26959<=Ng25692;

 always  @(posedge PCLK)
	Ng5821<=Ng25733;

 always  @(posedge PCLK)
	Ng6299<=Ng30536;

 always  @(posedge PCLK)
	Pg8416<=Pg7916;

 always  @(posedge PCLK)
	Ng2079<=Ng29246;

 always  @(posedge PCLK)
	Ng4698<=Ng34261;

 always  @(posedge PCLK)
	Ng3703<=Ng33611;

 always  @(posedge PCLK)
	Ng1559<=Ng25638;

 always  @(posedge PCLK)
	Ng943<=Ng34728;

 always  @(posedge PCLK)
	Ng411<=Ng29222;

 always  @(posedge PCLK)
	Pg9682<=Ng25742;

 always  @(posedge PCLK)
	Ng3953<=Ng30449;

 always  @(posedge PCLK)
	Ng2704<=Ng34608;

 always  @(posedge PCLK)
	Ng6035<=Ng24345;

 always  @(posedge PCLK)
	Ng1300<=Ng25635;

 always  @(posedge PCLK)
	Ng4057<=Ng25686;

 always  @(posedge PCLK)
	Ng5200<=Ng30461;

 always  @(posedge PCLK)
	Ng4843<=Ng34466;

 always  @(posedge PCLK)
	Ng5046<=Ng31901;

 always  @(posedge PCLK)
	Ng2250<=Ng29249;

 always  @(posedge PCLK)
	Ng26885<=Ng26882;

 always  @(posedge PCLK)
	Ng4549<=Ng33041;

 always  @(posedge PCLK)
	Ng2453<=Ng33011;

 always  @(posedge PCLK)
	Ng5841<=Ng25734;

 always  @(posedge PCLK)
	Pg14694<=Pg12300;

 always  @(posedge PCLK)
	Ng2912<=Ng34618;

 always  @(posedge PCLK)
	Ng2357<=Ng33010;

 always  @(posedge PCLK)
	Pg8920<=Pg8919;

 always  @(posedge PCLK)
	Ng164<=Ng31864;

 always  @(posedge PCLK)
	Ng4253<=Ng34630;

 always  @(posedge PCLK)
	Ng5016<=Ng31898;

 always  @(posedge PCLK)
	Ng3119<=Ng25653;

 always  @(posedge PCLK)
	Ng1351<=Ng25632;

 always  @(posedge PCLK)
	Ng1648<=Ng32988;

 always  @(posedge PCLK)
	Ng6972<=Ng33616;

 always  @(posedge PCLK)
	Ng5115<=Ng29280;

 always  @(posedge PCLK)
	Ng3352<=Ng33609;

 always  @(posedge PCLK)
	Ng6657<=Ng30563;

 always  @(posedge PCLK)
	Ng4552<=Ng33044;

 always  @(posedge PCLK)
	Ng3893<=Ng30437;

 always  @(posedge PCLK)
	Ng3211<=Ng30412;

 always  @(posedge PCLK)
	Pg13049<=Pg17604;

 always  @(posedge PCLK)
	Pg16624<=Pg16603;

 always  @(posedge PCLK)
	Ng5595<=Ng30491;

 always  @(posedge PCLK)
	Ng3614<=Ng30434;

 always  @(posedge PCLK)
	Ng2894<=Ng34612;

 always  @(posedge PCLK)
	Ng3125<=Ng29259;

 always  @(posedge PCLK)
	Pg16686<=Pg13865;

 always  @(posedge PCLK)
	Ng3821<=Ng25681;

 always  @(posedge PCLK)
	Ng4141<=Ng25687;

 always  @(posedge PCLK)
	Ng6974<=Ng33617;

 always  @(posedge PCLK)
	Ng5272<=Ng30479;

 always  @(posedge PCLK)
	Ng2735<=Ng29256;

 always  @(posedge PCLK)
	Ng728<=Ng28054;

 always  @(posedge PCLK)
	Ng6295<=Ng30535;

 always  @(posedge PCLK)
	Ng2661<=Ng30385;

 always  @(posedge PCLK)
	Ng1988<=Ng30361;

 always  @(posedge PCLK)
	Ng5128<=Ng25705;

 always  @(posedge PCLK)
	Ng1548<=Ng24260;

 always  @(posedge PCLK)
	Ng3106<=Ng29257;

 always  @(posedge PCLK)
	Ng4659<=Ng34461;

 always  @(posedge PCLK)
	Ng4358<=Ng34258;

 always  @(posedge PCLK)
	Ng1792<=Ng32993;

 always  @(posedge PCLK)
	Ng2084<=Ng33992;

 always  @(posedge PCLK)
	Ng3187<=Ng30394;

 always  @(posedge PCLK)
	Ng4311<=Ng34449;

 always  @(posedge PCLK)
	Ng2583<=Ng34019;

 always  @(posedge PCLK)
	Ng3003<=Ng21726;

 always  @(posedge PCLK)
	Ng1094<=Ng29231;

 always  @(posedge PCLK)
	Ng3841<=Ng25682;

 always  @(posedge PCLK)
	Ng4284<=Ng21897;

 always  @(posedge PCLK)
	Ng3191<=Ng30395;

 always  @(posedge PCLK)
	Ng4239<=Ng21892;

 always  @(posedge PCLK)
	Ng4180<=Pg8789;

 always  @(posedge PCLK)
	Ng691<=Ng28048;

 always  @(posedge PCLK)
	Ng534<=Ng34723;

 always  @(posedge PCLK)
	Ng385<=Ng25598;

 always  @(posedge PCLK)
	Ng2004<=Ng33987;

 always  @(posedge PCLK)
	Ng2527<=Ng30380;

 always  @(posedge PCLK)
	Ng5456<=Pg9555;

 always  @(posedge PCLK)
	Ng4420<=Ng26965;

 always  @(posedge PCLK)
	Ng5148<=Ng25706;

 always  @(posedge PCLK)
	Ng4507<=Ng30458;

 always  @(posedge PCLK)
	Ng5348<=Ng24338;

 always  @(posedge PCLK)
	Ng3223<=Ng30400;

 always  @(posedge PCLK)
	Ng2970<=Ng34623;

 always  @(posedge PCLK)
	Ng5698<=Ng24343;

 always  @(posedge PCLK)
	Ng5260<=Ng30473;

 always  @(posedge PCLK)
	Ng1521<=Ng24252;

 always  @(posedge PCLK)
	Ng3522<=Ng33028;

 always  @(posedge PCLK)
	Ng3115<=Ng29258;

 always  @(posedge PCLK)
	Ng3251<=Ng30407;

 always  @(posedge PCLK)
	Pg12832<=Ng26958;

 always  @(posedge PCLK)
	Ng4628<=Ng34457;

 always  @(posedge PCLK)
	Ng1996<=Ng33568;

 always  @(posedge PCLK)
	Pg8342<=Ng25663;

 always  @(posedge PCLK)
	Ng4515<=Ng26964;

 always  @(posedge PCLK)
	Pg8787<=Pg8786;

 always  @(posedge PCLK)
	Ng4300<=Ng34735;

 always  @(posedge PCLK)
	Ng1724<=Ng30352;

 always  @(posedge PCLK)
	Ng1379<=Ng33543;

 always  @(posedge PCLK)
	Pg11388<=Ng24271;

 always  @(posedge PCLK)
	Ng1878<=Ng33981;

 always  @(posedge PCLK)
	Ng5619<=Ng30500;

 always  @(posedge PCLK)
	Ng71<=Ng34786;

 always  @(posedge PCLK)
	wire4437<=Ng29277;

 assign Pg34972 = ( (~ n4486) ) | ( (~ Ng22) ) ;
 assign wire4366 = ( Ng4369  &  Ng4366 ) | ( Ng4369  &  n1368 ) ;
 assign Pg34927 = ( (~ n1121) ) | ( (~ Ng22) ) ;
 assign Pg34925 = ( (~ n1141) ) | ( (~ Ng22) ) ;
 assign Pg34923 = ( (~ n204) ) | ( (~ Ng22) ) ;
 assign Pg34921 = ( (~ n1119) ) | ( (~ Ng22) ) ;
 assign Pg34919 = ( (~ n1092) ) | ( (~ Ng22) ) ;
 assign Pg34917 = ( (~ n981) ) | ( (~ Ng22) ) ;
 assign Pg34915 = ( (~ n1132) ) | ( (~ Ng22) ) ;
 assign Pg34913 = ( (~ n569) ) | ( (~ Ng22) ) ;
 assign wire4376 = ( Ng890  &  Ng528 ) | ( Ng890  &  n1170 ) | ( Ng890  &  (~ Ng479) ) ;
 assign Pg34597 =((~ Pg6753) & Pg6753);
 assign wire4378 = ( (~ Pg113) ) | ( (~ Ng2868) ) ;
 assign wire4379 = ( (~ Pg113) ) | ( (~ Ng2873) ) ;
 assign Pg34435 = ( (~ n6112) ) ;
 assign Pg34425 = ( (~ n1189) ) | ( (~ n1636) ) ;
 assign Pg34383 = ( n1129 ) | ( (~ n1169) ) | ( (~ n1638) ) ;
 assign Pg34240 =((~ Pg6753) & Pg6753);
 assign Pg34239 =((~ Pg6753) & Pg6753);
 assign Pg34238 =((~ Pg6753) & Pg6753);
 assign Pg34237 =((~ Pg6753) & Pg6753);
 assign Pg34236 =((~ Pg6753) & Pg6753);
 assign Pg34235 =((~ Pg6753) & Pg6753);
 assign Pg34234 =((~ Pg6753) & Pg6753);
 assign Pg34233 =((~ Pg6753) & Pg6753);
 assign Pg34232 =((~ Pg6753) & Pg6753);
 assign Pg34221 = ( (~ n1168) ) | ( (~ n1636) ) ;
 assign Pg34201 = ( n1178 ) | ( (~ n1401) ) | ( (~ n1638) ) ;
 assign wire4394 = ( Ng4646  &  n1100 ) | ( Ng4646  &  n1145 ) ;
 assign Pg33950 =((~ Pg6753) & Pg6753);
 assign Pg33949 =((~ Pg6753) & Pg6753);
 assign Pg33948 =((~ Pg6753) & Pg6753);
 assign Pg33947 =((~ Pg6753) & Pg6753);
 assign Pg33946 =((~ Pg6753) & Pg6753);
 assign Pg33945 =((~ Pg6753) & Pg6753);
 assign Pg33935 = ( (~ n1175) ) ;
 assign Pg33874 = ( wire4507 ) | ( n1160 ) | ( (~ Ng4507) ) ;
 assign Pg33659 = ( n1191 ) | ( (~ n1638) ) | ( (~ n6113) ) ;
 assign Pg33636 = ( (~ n1194) ) ;
 assign wire4406 = ( Pg17291  &  (~ Ng1171) ) | ( Pg17291  &  n1142 ) ;
 assign Pg33435 = ( (~ Ng2729)  &  n5700 ) | ( Ng2729  &  n5701 ) | ( n5700  &  n5701 ) ;
 assign Pg33079 = ( (~ Ng2729)  &  n5698 ) | ( Ng2729  &  n5699 ) | ( n5698  &  n5699 ) ;
 assign Pg32975 = ( (~ n3401) ) ;
 assign Pg32454 =((~ Pg6753) & Pg6753);
 assign Pg32429 =((~ Pg6753) & Pg6753);
 assign Pg32185 = ( n2489  &  n2490  &  n2491  &  n2492 ) ;
 assign Pg31863 = ( (~ n4553) ) ;
 assign Pg31862 = ( (~ n4321) ) ;
 assign Pg31860 = ( (~ n4527) ) ;
 assign Pg31793 = ( (~ n186) ) ;
 assign Pg31521 = ( (~ n6112) ) ;
 assign Pg30331 = ( (~ Ng2831) ) ;
 assign Pg30330 = ( (~ Ng2834) ) ;
 assign Pg30329 = ( (~ wire4426) ) ;
 assign Pg30327 = ( (~ Ng37) ) ;
 assign Pg28042 = ( n184 ) | ( n185 ) ;
 assign Pg28041 = ( n182 ) | ( (~ n5079) ) ;
 assign Pg28030 = ( n180 ) | ( n181 ) ;
 assign Pg26877 = ( (~ n177) ) ;
 assign Pg26876 = ( (~ n174) ) ;
 assign Pg26875 = ( (~ n171) ) ;
 assign Pg26801 = ( (~ n3401) ) ;
 assign Pg25590 =((~ Pg6753) & Pg6753);
 assign Pg25589 =((~ Pg6753) & Pg6753);
 assign Pg25588 =((~ Pg6753) & Pg6753);
 assign Pg25587 =((~ Pg6753) & Pg6753);
 assign Pg25586 =((~ Pg6753) & Pg6753);
 assign Pg25585 =((~ Pg6753) & Pg6753);
 assign Pg25584 =((~ Pg6753) & Pg6753);
 assign Pg25583 =((~ Pg6753) & Pg6753);
 assign Pg25582 =((~ Pg6753) & Pg6753);
 assign Pg25259 = ( (~ n4321) ) ;
 assign Pg25167 = ( (~ n4553) ) ;
 assign Pg25114 = ( (~ n4527) ) ;
 assign Pg24151 =((~ Pg6753) & Pg6753);
 assign Pg23759 = ( (~ Ng2831) ) ;
 assign Pg23652 = ( (~ Ng2834) ) ;
 assign Pg23612 = ( (~ wire4426) ) ;
 assign Pg23190 = ( (~ Ng25)  &  (~ Ng22) ) ;
 assign Pg23002 = ( (~ Ng37) ) ;
 assign Pg21727 = ( (~ Pg35)  &  Ng3003 ) ;
 assign Pg12833 = ( (~ Pg5) ) ;
 assign n160 = ( (~ Pg35) ) | ( n4887 ) ;
 assign n172 = ( Ng1830 ) | ( Ng2098 ) | ( Ng1696 ) | ( Ng1964 ) ;
 assign n173 = ( n1410  &  Pg35 ) ;
 assign n171 = ( n172  &  n173 ) ;
 assign n175 = ( Ng1710 ) | ( Ng1858 ) | ( Ng1844 ) | ( Ng2126 ) | ( Ng1992 ) | ( Ng1978 ) | ( Ng1724 ) | ( Ng2112 ) ;
 assign n176 = ( n1243  &  Pg35 ) ;
 assign n174 = ( n175  &  n176 ) ;
 assign n178 = ( Ng1913 ) | ( Ng2047 ) | ( Ng1932 ) | ( Ng1798 ) | ( Ng1644 ) | ( Ng2066 ) | ( Ng1664 ) | ( Ng1779 ) ;
 assign n179 = ( n1242  &  Pg35 ) ;
 assign n177 = ( n178  &  n179 ) ;
 assign n180 = ( (~ n1134)  &  n3911  &  (~ n4366) ) | ( n3911  &  (~ n4366)  &  (~ n4567) ) ;
 assign n181 = ( (~ n1131)  &  (~ n1134)  &  n3914 ) | ( (~ n1133)  &  (~ n1134)  &  n3914 ) ;
 assign n182 = ( (~ Pg35) ) | ( n1411 ) ;
 assign n184 = ( (~ Pg35) ) | ( Ng962 ) ;
 assign n185 = ( (~ Pg35) ) | ( Ng1306 ) ;
 assign n186 = ( n2567  &  n2564 ) | ( n2567  &  n2565 ) | ( n2567  &  (~ n5591) ) ;
 assign n188 = ( Pg35  &  n2296  &  n2297 ) | ( n2296  &  n2297  &  (~ Ng5052) ) ;
 assign Ng33046 = ( (~ n188) ) ;
 assign n189 = ( n1611  &  n1604 ) | ( n1611  &  n1610 ) | ( n1611  &  n1601 ) ;
 assign Ng34441 = ( (~ n189) ) ;
 assign n190 = ( (~ n1267)  &  n1884  &  n1885 ) | ( n1884  &  n1885  &  n1883 ) ;
 assign Ng33982 = ( (~ n190) ) ;
 assign n191 = ( Pg35  &  n1793 ) | ( n1793  &  (~ Ng2380) ) ;
 assign Ng34007 = ( (~ n191) ) ;
 assign n192 = ( n3008  &  n3009  &  n160 ) | ( n3008  &  n3009  &  n3007 ) ;
 assign Ng30405 = ( (~ n192) ) ;
 assign n193 = ( n2980  &  n2981  &  n160 ) | ( n2980  &  n2981  &  n2979 ) ;
 assign Ng30416 = ( (~ n193) ) ;
 assign n194 = ( n2839  &  n2840  &  n160 ) | ( n2839  &  n2840  &  n2838 ) ;
 assign Ng30466 = ( (~ n194) ) ;
 assign n195 = ( Pg35  &  n1499 ) | ( n1499  &  (~ Ng2984) ) ;
 assign Ng34617 = ( (~ n195) ) ;
 assign n196 = ( (~ n1257)  &  n1912  &  n1913 ) | ( n1912  &  n1913  &  n1911 ) ;
 assign Ng33974 = ( (~ n196) ) ;
 assign n197 = ( n160  &  n2732  &  n2733 ) | ( n2732  &  n2733  &  n2731 ) ;
 assign Ng30505 = ( (~ n197) ) ;
 assign n198 = ( n1898  &  n2163 ) | ( n1898  &  (~ Ng1772) ) | ( n2163  &  (~ Ng1802) ) | ( (~ Ng1772)  &  (~ Ng1802) ) ;
 assign Ng33554 = ( (~ n198) ) ;
 assign n199 = ( n2932  &  n2933  &  n160 ) | ( n2932  &  n2933  &  n2333 ) ;
 assign Ng30432 = ( (~ n199) ) ;
 assign n200 = ( (~ Ng6215)  &  (~ Ng6219) ) | ( (~ Ng6219)  &  n2248 ) | ( (~ Ng6215)  &  n2250 ) | ( n2248  &  n2250 ) ;
 assign Ng33064 = ( (~ n200) ) ;
 assign n201 = ( n1377  &  n1378  &  Ng807 ) | ( n1377  &  n1378  &  n1371 ) ;
 assign Ng34881 = ( (~ n201) ) ;
 assign n202 = ( (~ Ng1061)  &  n4245 ) | ( Ng1061  &  (~ n4245) ) ;
 assign Ng24232 = ( n202 ) | ( (~ n5636) ) ;
 assign n206 = ( Ng4172 ) | ( Ng4153 ) ;
 assign n204 = ( n1284  &  n1285  &  n1286  &  n1287 ) ;
 assign Ng34733 = ( n206  &  Pg35 ) ;
 assign n207 = ( Pg35  &  n2334 ) | ( Pg35  &  n2341 ) | ( n2334  &  (~ Ng3506) ) | ( n2341  &  (~ Ng3506) ) ;
 assign Ng33026 = ( (~ n207) ) ;
 assign n208 = ( n2547  &  n2548  &  Ng749 ) | ( n2547  &  n2548  &  n2546 ) ;
 assign Ng31867 = ( (~ n208) ) ;
 assign n212 = ( (~ Pg17739)  &  (~ Pg14738) ) | ( (~ Pg17739)  &  Pg12350 ) | ( Pg14738  &  Pg12350 ) ;
 assign Ng24344 = ( Pg35  &  (~ Pg17646)  &  (~ Pg17607)  &  (~ Pg13068)  &  n212 ) ;
 assign n213 = ( (~ n1271)  &  n1940  &  n1941 ) | ( n1940  &  n1941  &  n1939 ) ;
 assign Ng33966 = ( (~ n213) ) ;
 assign n214 = ( n2180  &  n2181  &  (~ n4770) ) | ( n2180  &  n2181  &  (~ Ng1714) ) ;
 assign Ng33550 = ( (~ n214) ) ;
 assign Ng30393 = ( (~ n2351)  &  (~ Ng3155) ) ;
 assign n217 = ( n3702  &  n3703  &  (~ Ng2165) ) | ( n3702  &  n3703  &  (~ n4956) ) ;
 assign Ng29248 = ( (~ n217) ) ;
 assign n218 = ( (~ Ng3689) ) | ( n5150 ) ;
 assign Ng24274 = ( (~ Pg35)  &  Ng3694 ) | ( Ng3694  &  n218 ) ;
 assign n219 = ( (~ n1257)  &  n1915  &  n1916 ) | ( n1915  &  n1916  &  n1914 ) ;
 assign Ng33973 = ( (~ n219) ) ;
 assign n220 = ( Pg35  &  n3113 ) | ( (~ Ng1964)  &  n3113 ) ;
 assign Ng30360 = ( (~ n220) ) ;
 assign n221 = ( (~ Ng4621)  &  n1548 ) | ( n1548  &  n1551 ) | ( (~ Ng4621)  &  (~ Ng4639) ) | ( n1551  &  (~ Ng4639) ) ;
 assign Ng34460 = ( (~ n221) ) ;
 assign n222 = ( n160  &  n2760  &  n2761 ) | ( n2760  &  n2761  &  n2759 ) ;
 assign Ng30494 = ( (~ n222) ) ;
 assign n223 = ( Pg35  &  n3056  &  (~ n5842) ) | ( n3056  &  (~ Ng2652)  &  (~ n5842) ) ;
 assign Ng30384 = ( (~ n223) ) ;
 assign n227 = ( (~ Pg17711)  &  (~ Pg14694) ) | ( (~ Pg17711)  &  Pg12300 ) | ( Pg14694  &  Pg12300 ) ;
 assign Ng24340 = ( Pg35  &  (~ Pg17604)  &  (~ Pg17580)  &  (~ Pg13049)  &  n227 ) ;
 assign n228 = ( n3809  &  n3810  &  Ng490 ) | ( n3809  &  n3810  &  (~ n5058) ) ;
 assign Ng29223 = ( (~ n228) ) ;
 assign n229 = ( n1683  &  n1684  &  Ng772 ) | ( n1683  &  n1684  &  n1682 ) ;
 assign Ng34252 = ( (~ n229) ) ;
 assign n230 = ( n160  &  n2775  &  n2776 ) | ( n2775  &  n2776  &  n2774 ) ;
 assign Ng30489 = ( (~ n230) ) ;
 assign n231 = ( (~ Ng6177)  &  n3243  &  (~ n5891) ) | ( n3243  &  n3242  &  (~ n5891) ) ;
 assign Ng29301 = ( (~ n231) ) ;
 assign n232 = ( Pg35  &  n2351 ) | ( Pg35  &  n2352 ) | ( n2351  &  (~ Ng3161) ) | ( n2352  &  (~ Ng3161) ) ;
 assign Ng33022 = ( (~ n232) ) ;
 assign n233 = ( n160  &  n2754  &  n2755 ) | ( n2754  &  n2755  &  n2753 ) ;
 assign Ng30496 = ( (~ n233) ) ;
 assign n234 = ( (~ n1245)  &  n2304  &  (~ n2521) ) | ( (~ n1245)  &  n2304  &  (~ Ng4543) ) ;
 assign Ng33043 = ( (~ n234) ) ;
 assign n235 = ( n3581  &  Ng3457  &  (~ n5941) ) | ( n3581  &  n3580  &  (~ n5941) ) ;
 assign Ng29263 = ( (~ n235) ) ;
 assign n236 = ( n160  &  n2653  &  (~ n6287) ) | ( n2653  &  n2652  &  (~ n6287) ) ;
 assign Ng30533 = ( (~ n236) ) ;
 assign n237 = ( (~ n1260)  &  n1762  &  n1763 ) | ( n1762  &  n1763  &  n1761 ) ;
 assign Ng34015 = ( (~ n237) ) ;
 assign n238 = ( n1729  &  n1726 ) | ( n1729  &  n1727 ) | ( n1729  &  (~ Ng4801) ) ;
 assign Ng34031 = ( (~ n238) ) ;
 assign n239 = ( Pg35  &  n1582  &  n1583 ) | ( n1582  &  n1583  &  (~ Ng4584) ) ;
 assign Ng34452 = ( (~ n239) ) ;
 assign n240 = ( (~ Pg35) ) | ( (~ Ng6199) ) ;
 assign Ng34646 = ( (~ n240) ) ;
 assign n241 = ( (~ n1273)  &  n1813  &  n1814 ) | ( n1813  &  n1814  &  n1812 ) ;
 assign Ng34001 = ( (~ n241) ) ;
 assign n242 = ( Pg35  &  n4140  &  n4141 ) | ( (~ Ng1379)  &  n4140  &  n4141 ) ;
 assign Ng25633 = ( (~ n242) ) ;
 assign n243 = ( Pg35  &  n4222 ) | ( n4222  &  (~ Ng1579) ) ;
 assign Ng24259 = ( (~ n243) ) ;
 assign n244 = ( (~ Ng5176)  &  (~ Ng5180) ) | ( (~ Ng5180)  &  n2287 ) | ( (~ Ng5176)  &  n2289 ) | ( n2287  &  n2289 ) ;
 assign Ng33049 = ( (~ n244) ) ;
 assign n245 = ( Pg35  &  n1512 ) | ( n1512  &  (~ Ng2890) ) ;
 assign Ng34609 = ( (~ n245) ) ;
 assign n246 = ( Pg35  &  n2541  &  n2542 ) | ( (~ Ng1018)  &  n2541  &  n2542 ) ;
 assign Ng31869 = ( (~ n246) ) ;
 assign n247 = ( n160  &  n2772  &  n2773 ) | ( n2772  &  n2773  &  n2771 ) ;
 assign Ng30490 = ( (~ n247) ) ;
 assign n248 = ( n2947  &  n2948  &  n160 ) | ( n2947  &  n2948  &  n2946 ) ;
 assign Ng30427 = ( (~ n248) ) ;
 assign n249 = ( n4210  &  n4268 ) | ( (~ Ng4264)  &  n4268 ) | ( n4210  &  (~ Ng4258) ) | ( (~ Ng4264)  &  (~ Ng4258) ) ;
 assign Ng21894 = ( (~ n249) ) ;
 assign n250 = ( n1943  &  n1944  &  Ng767 ) | ( n1943  &  n1944  &  n1942 ) ;
 assign Ng33965 = ( (~ n250) ) ;
 assign n251 = ( (~ Pg35) ) | ( (~ Ng5853) ) ;
 assign Ng34645 = ( (~ n251) ) ;
 assign n252 = ( n1656  &  n1657  &  n1655 ) | ( n1656  &  n1657  &  n1653 ) ;
 assign Ng34267 = ( (~ n252) ) ;
 assign n253 = ( (~ Pg35) ) | ( (~ Ng5507) ) ;
 assign Ng34644 = ( (~ n253) ) ;
 assign n254 = ( n160  &  n2650  &  n2651 ) | ( n2650  &  n2651  &  n2649 ) ;
 assign Ng30534 = ( (~ n254) ) ;
 assign n255 = ( Pg35  &  n2225  &  n2226 ) | ( n2225  &  n2226  &  (~ Ng291) ) ;
 assign Ng33535 = ( (~ n255) ) ;
 assign n256 = ( n160  &  n2748  &  (~ n6318) ) | ( n2271  &  n2748  &  (~ n6318) ) ;
 assign Ng30498 = ( (~ n256) ) ;
 assign n257 = ( Pg35  &  (~ n4184) ) | ( (~ n4184)  &  (~ Ng559) ) ;
 assign Ng25613 = ( (~ n257) ) ;
 assign n258 = ( n1631  &  Ng608  &  (~ n6203) ) | ( n1631  &  n1629  &  (~ n6203) ) ;
 assign Ng34438 = ( (~ n258) ) ;
 assign n259 = ( n2916  &  n2917  &  n160 ) | ( n2916  &  n2917  &  n2915 ) ;
 assign Ng30439 = ( (~ n259) ) ;
 assign n260 = ( n160  &  n2630  &  n2631 ) | ( n2630  &  n2631  &  n2629 ) ;
 assign Ng30541 = ( (~ n260) ) ;
 assign n261 = ( n160  &  n2690  &  (~ n6299) ) | ( n2258  &  n2690  &  (~ n6299) ) ;
 assign Ng30519 = ( (~ n261) ) ;
 assign n262 = ( (~ Ng921)  &  n4165 ) | ( n4165  &  n4168 ) | ( (~ Ng921)  &  (~ Ng904) ) | ( n4168  &  (~ Ng904) ) ;
 assign Ng25621 = ( (~ n262) ) ;
 assign n263 = ( (~ Pg35) ) | ( (~ n4673) ) ;
 assign Ng34036 = ( Ng4871  &  n263 ) ;
 assign n264 = ( n160  &  n2809  &  n2810 ) | ( n2809  &  n2810  &  n2808 ) ;
 assign Ng30476 = ( (~ n264) ) ;
 assign n265 = ( n2941  &  n2942  &  n160 ) | ( n2941  &  n2942  &  n2940 ) ;
 assign Ng30429 = ( (~ n265) ) ;
 assign n266 = ( n2428  &  n2433  &  n2434 ) | ( n2433  &  n2434  &  (~ Ng1926) ) ;
 assign Ng32997 = ( (~ n266) ) ;
 assign n267 = ( Pg35  &  n2250 ) | ( Pg35  &  n2251 ) | ( n2250  &  (~ Ng6209) ) | ( n2251  &  (~ Ng6209) ) ;
 assign Ng33063 = ( (~ n267) ) ;
 assign n268 = ( n2956  &  n2957  &  n160 ) | ( n2956  &  n2957  &  n2955 ) ;
 assign Ng30424 = ( (~ n268) ) ;
 assign n269 = ( Pg35  &  n2484  &  n2485 ) | ( n2484  &  n2485  &  (~ Ng287) ) ;
 assign Ng32977 = ( (~ n269) ) ;
 assign n270 = ( (~ Pg35) ) | ( (~ n4676) ) ;
 assign Ng34026 = ( Ng4646  &  n270 ) ;
 assign n271 = ( n2968  &  n2969  &  n160 ) | ( n2968  &  n2969  &  n2967 ) ;
 assign Ng30420 = ( (~ n271) ) ;
 assign n272 = ( n1873  &  n2151 ) | ( n2151  &  (~ Ng1862) ) ;
 assign Ng33560 = ( (~ n272) ) ;
 assign n273 = ( Pg35  &  n3800  &  n3801 ) | ( n3800  &  n3801  &  (~ Ng671) ) ;
 assign Ng29226 = ( (~ n273) ) ;
 assign n274 = ( (~ Ng843)  &  n4248 ) | ( Ng843  &  (~ n4248) ) ;
 assign Ng25619 = ( (~ Pg35)  &  Ng837 ) | ( Ng837  &  n274 ) ;
 assign n275 = ( n1574  &  n1572 ) | ( n1574  &  (~ Ng4322) ) | ( n1574  &  (~ n4642) ) ;
 assign Ng34455 = ( (~ n275) ) ;
 assign n276 = ( Pg35  &  n1963 ) | ( n1963  &  (~ Ng6395) ) | ( Pg35  &  (~ n6116) ) | ( (~ Ng6395)  &  (~ n6116) ) ;
 assign Ng33625 = ( (~ n276) ) ;
 assign n277 = ( n1416  &  n1417  &  Ng622 ) | ( n1416  &  n1417  &  n1415 ) ;
 assign Ng34790 = ( (~ n277) ) ;
 assign Ng30414 = ( (~ n2338)  &  (~ Ng3506) ) ;
 assign n280 = ( Pg35  &  n3043 ) | ( (~ Ng2834)  &  n3043 ) ;
 assign Ng30390 = ( (~ n280) ) ;
 assign n282 = ( (~ Ng246) ) | ( (~ Ng239) ) | ( (~ Ng232) ) | ( (~ Ng225) ) | ( Ng269 ) | ( Ng262 ) | ( Ng255 ) ;
 assign n281 = ( (~ Ng246)  &  (~ Ng239)  &  (~ Ng232)  &  (~ Ng225)  &  Ng269  &  Ng262  &  Ng255 ) ;
 assign Ng25594 = ( n282  &  Pg35  &  Ng278 ) | ( n282  &  Pg35  &  n281 ) ;
 assign Ng34034 = ( Ng4836  &  n263 ) ;
 assign n283 = ( (~ Ng1036)  &  n2210 ) | ( (~ Ng1036)  &  (~ Ng1030) ) | ( n2210  &  (~ n5590) ) | ( (~ Ng1030)  &  (~ n5590) ) ;
 assign Ng33541 = ( (~ n283) ) ;
 assign n284 = ( Pg35  &  n3452  &  n3819 ) | ( n3452  &  n3819  &  (~ Ng5272) ) ;
 assign Ng28093 = ( (~ n284) ) ;
 assign n285 = ( n160  &  n3011  &  (~ n6405) ) | ( n3011  &  n3010  &  (~ n6405) ) ;
 assign Ng30404 = ( (~ n285) ) ;
 assign n286 = ( n3239  &  n160 ) | ( n3239  &  Ng6195  &  n3238 ) ;
 assign Ng29303 = ( (~ n286) ) ;
 assign n287 = ( Ng1135  &  n3996  &  n3997 ) | ( n3996  &  n3997  &  (~ n5090) ) ;
 assign Ng26917 = ( (~ n287) ) ;
 assign n288 = ( n1970  &  n1971  &  n1969 ) | ( n1970  &  n1971  &  (~ Ng6395) ) ;
 assign Ng33624 = ( (~ n288) ) ;
 assign n289 = ( n1372  &  n1371 ) | ( n1372  &  (~ Ng807) ) ;
 assign Ng34911 = ( (~ n289) ) ;
 assign n290 = ( (~ Pg35) ) | ( (~ Ng3853) ) ;
 assign Ng34627 = ( (~ n290) ) ;
 assign n291 = ( n2374  &  n2379  &  n2380 ) | ( n2379  &  n2380  &  (~ Ng2485) ) ;
 assign Ng33013 = ( (~ n291) ) ;
 assign n292 = ( n2475  &  n2476  &  Ng925 ) | ( n2475  &  n2476  &  n2474 ) ;
 assign Ng32981 = ( (~ n292) ) ;
 assign n293 = ( n160  &  n2793  &  n2794 ) | ( n2793  &  n2794  &  n2792 ) ;
 assign Ng30483 = ( (~ n293) ) ;
 assign n294 = ( (~ Ng1798)  &  n2443  &  n2444 ) | ( n2439  &  n2443  &  n2444 ) ;
 assign Ng32994 = ( (~ n294) ) ;
 assign n295 = ( n1994  &  n3868  &  Ng4076 ) | ( n1994  &  n3868  &  n3867 ) ;
 assign Ng28070 = ( (~ n295) ) ;
 assign n296 = ( n2874  &  n2875  &  n160 ) | ( n2874  &  n2875  &  n2320 ) ;
 assign Ng30453 = ( (~ n296) ) ;
 assign n297 = ( n2219  &  n2220  &  Ng763 ) | ( n2219  &  n2220  &  n2218 ) ;
 assign Ng33539 = ( (~ n297) ) ;
 assign n298 = ( n160  &  n2674  &  n2675 ) | ( n2674  &  n2675  &  n2673 ) ;
 assign Ng30526 = ( (~ n298) ) ;
 assign n299 = ( Pg35  &  n3940 ) | ( (~ Ng4427)  &  n3940 ) ;
 assign Ng26951 = ( (~ n299) ) ;
 assign Ng34035 = ( Ng4864  &  n263 ) ;
 assign n300 = ( Pg35  &  n1464 ) | ( n1464  &  (~ Ng4717) ) ;
 assign Ng34636 = ( (~ n300) ) ;
 assign n301 = ( n2482  &  Ng590  &  (~ n6256) ) | ( n2482  &  n2480  &  (~ n6256) ) ;
 assign Ng32978 = ( (~ n301) ) ;
 assign n302 = ( Pg35  &  (~ n3141)  &  (~ n5878) ) | ( (~ n3141)  &  (~ Ng1612)  &  (~ n5878) ) ;
 assign Ng30348 = ( (~ n302) ) ;
 assign n306 = ( (~ Pg17674)  &  (~ Pg14662) ) | ( (~ Pg17674)  &  Pg12238 ) | ( Pg14662  &  Pg12238 ) ;
 assign Ng24336 = ( Pg35  &  (~ Pg17577)  &  (~ Pg17519)  &  (~ Pg13039)  &  n306 ) ;
 assign n307 = ( n3289  &  Ng6154  &  (~ n5896) ) | ( n3289  &  n3288  &  (~ n5896) ) ;
 assign Ng29298 = ( (~ n307) ) ;
 assign n308 = ( n160  &  n2746  &  n2747 ) | ( n2746  &  n2747  &  n2745 ) ;
 assign Ng30499 = ( (~ n308) ) ;
 assign n309 = ( (~ n1257)  &  n1906  &  n1907 ) | ( n1906  &  n1907  &  (~ n4764) ) ;
 assign Ng33976 = ( (~ n309) ) ;
 assign n310 = ( n3176  &  n3177  &  Ng744 ) | ( n3176  &  n3177  &  n3175 ) ;
 assign Ng30335 = ( (~ n310) ) ;
 assign n311 = ( Pg35  &  n1462 ) | ( n1462  &  (~ Ng4722) ) ;
 assign Ng34637 = ( (~ n311) ) ;
 assign n312 = ( n160  &  n2668  &  n2669 ) | ( n2668  &  n2669  &  n2667 ) ;
 assign Ng30528 = ( (~ n312) ) ;
 assign n313 = ( Pg35  &  n2686 ) | ( n2686  &  (~ Ng5961) ) ;
 assign Ng30521 = ( (~ n313) ) ;
 assign n314 = ( (~ Pg17400)  &  n4241  &  n4242 ) | ( n4235  &  n4241  &  n4242 ) ;
 assign Ng24239 = ( (~ n314) ) ;
 assign Ng34259 = ( (~ Pg35)  &  Ng4633 ) | ( Ng4633  &  (~ Ng4639)  &  (~ n1560) ) ;
 assign n317 = ( n160  &  n2815  &  n2816 ) | ( n2815  &  n2816  &  n2814 ) ;
 assign Ng30474 = ( (~ n317) ) ;
 assign n318 = ( (~ Pg35) ) | ( (~ Ng5160) ) ;
 assign Ng34643 = ( (~ n318) ) ;
 assign n319 = ( n160  &  n2717  &  n2718 ) | ( n2717  &  n2718  &  n2716 ) ;
 assign Ng30510 = ( (~ n319) ) ;
 assign n320 = ( n1426  &  n1428 ) ;
 assign Ng34729 = ( (~ n320) ) ;
 assign n321 = ( (~ Pg35) ) | ( (~ Ng3151) ) ;
 assign Ng34625 = ( (~ n321) ) ;
 assign n322 = ( Pg35  &  n2331 ) | ( (~ Ng3522)  &  n2331 ) | ( Pg35  &  n2334 ) | ( (~ Ng3522)  &  n2334 ) ;
 assign Ng33029 = ( (~ n322) ) ;
 assign n323 = ( n1994  &  n1995  &  Ng4104 ) | ( n1994  &  n1995  &  n1993 ) ;
 assign Ng33615 = ( (~ n323) ) ;
 assign n324 = ( (~ n6074)  &  Pg9251 ) | ( n6074  &  (~ Pg9251) ) ;
 assign Ng24281 = ( n324  &  Pg35 ) ;
 assign n325 = ( (~ n1269)  &  n1829  &  n1830 ) | ( n1829  &  n1830  &  (~ n4734) ) ;
 assign Ng33997 = ( (~ n325) ) ;
 assign n326 = ( n1796  &  n2088 ) | ( n2088  &  (~ Ng2287) ) ;
 assign Ng33584 = ( (~ n326) ) ;
 assign n327 = ( (~ Ng4269)  &  n4211 ) | ( (~ Ng4269)  &  (~ Ng4273) ) | ( n4211  &  n4212 ) | ( (~ Ng4273)  &  n4212 ) ;
 assign Ng24280 = ( (~ n327) ) ;
 assign n328 = ( Pg35  &  n3990  &  (~ n6186) ) | ( (~ Ng1384)  &  n3990  &  (~ n6186) ) ;
 assign Ng26920 = ( (~ n328) ) ;
 assign n329 = ( Pg35  &  n3294 ) | ( (~ Ng5831)  &  n3294 ) ;
 assign Ng29296 = ( (~ n329) ) ;
 assign n330 = ( n1211  &  (~ Ng1193) ) | ( (~ Ng1171)  &  n1211  &  Ng1183 ) ;
 assign n331 = ( (~ Pg7916)  &  Ng1171 ) | ( Pg7916  &  (~ Ng1171) ) ;
 assign Ng30338 = ( Pg35  &  n330 ) | ( Pg35  &  n331 ) ;
 assign n332 = ( (~ Ng4264)  &  n4209 ) | ( (~ Ng4264)  &  (~ Ng4269) ) | ( n4209  &  n4267 ) | ( (~ Ng4269)  &  n4267 ) ;
 assign Ng21895 = ( (~ n332) ) ;
 assign n333 = ( Pg35  &  n1703 ) | ( Pg35  &  n1704 ) | ( n1703  &  (~ Ng4818) ) | ( n1704  &  (~ Ng4818) ) ;
 assign Ng34041 = ( (~ n333) ) ;
 assign n334 = ( n160  &  n2757  &  n2758 ) | ( n2757  &  n2758  &  n2756 ) ;
 assign Ng30495 = ( (~ n334) ) ;
 assign n335 = ( Ng4864 ) | ( Ng4878 ) | ( Ng4836 ) | ( Ng4871 ) ;
 assign Ng29279 = ( Pg35  &  n335  &  (~ n5923) ) | ( Pg35  &  (~ n5348)  &  (~ n5923) ) ;
 assign n338 = ( Pg35  &  n4129 ) | ( n4129  &  (~ Ng3139) ) ;
 assign Ng25655 = ( (~ n338) ) ;
 assign n339 = ( n160  &  n3014  &  (~ n6406) ) | ( n3014  &  n3013  &  (~ n6406) ) ;
 assign Ng30403 = ( (~ n339) ) ;
 assign n340 = ( (~ n1245)  &  (~ n1253)  &  (~ n2521) ) | ( (~ n1245)  &  (~ n1253)  &  (~ Ng4540) ) ;
 assign Ng33042 = ( (~ n340) ) ;
 assign n341 = ( n2971  &  n2972  &  n160 ) | ( n2971  &  n2972  &  n2970 ) ;
 assign Ng30419 = ( (~ n341) ) ;
 assign n342 = ( (~ Pg35)  &  n3824 ) | ( n3820  &  n3824 ) | ( n3824  &  n3823 ) ;
 assign Ng28090 = ( (~ n342) ) ;
 assign n343 = ( Pg35  &  n1452 ) | ( n1452  &  (~ Ng4912) ) ;
 assign Ng34642 = ( (~ n343) ) ;
 assign n344 = ( Pg35  &  n3089 ) | ( (~ Ng2255)  &  n3089 ) ;
 assign Ng30370 = ( (~ n344) ) ;
 assign n345 = ( n1593  &  n1591 ) | ( n1593  &  n1589 ) | ( n1593  &  n1592 ) ;
 assign Ng34448 = ( (~ n345) ) ;
 assign n346 = ( n3952  &  (~ Ng4375) ) | ( Pg35  &  n3952  &  (~ Ng4382) ) ;
 assign Ng26946 = ( (~ n346) ) ;
 assign n347 = ( Pg35  &  n1510 ) | ( n1510  &  (~ Ng2844) ) ;
 assign Ng34610 = ( (~ n347) ) ;
 assign n348 = ( n3812  &  n4259 ) | ( n4259  &  (~ Ng417) ) | ( n3812  &  (~ Ng446) ) | ( (~ Ng417)  &  (~ Ng446) ) ;
 assign Ng24209 = ( (~ n348) ) ;
 assign n349 = ( n160  &  n2735  &  n2736 ) | ( n2735  &  n2736  &  n2734 ) ;
 assign Ng30504 = ( (~ n349) ) ;
 assign n350 = ( Pg35  &  n4123 ) | ( n4123  &  (~ Ng3490) ) ;
 assign Ng25669 = ( (~ n350) ) ;
 assign Ng30480 = ( (~ n2276)  &  (~ Ng5511) ) ;
 assign n353 = ( Pg35  &  n2338 ) | ( Pg35  &  n2339 ) | ( n2338  &  (~ Ng3512) ) | ( n2339  &  (~ Ng3512) ) ;
 assign Ng33027 = ( (~ n353) ) ;
 assign n354 = ( Pg35  &  n1920 ) | ( n1920  &  (~ Ng1687) ) ;
 assign Ng33972 = ( (~ n354) ) ;
 assign n355 = ( Pg35  &  n3343  &  n3817 ) | ( n3343  &  n3817  &  (~ Ng5965) ) ;
 assign Ng28099 = ( (~ n355) ) ;
 assign n356 = ( n3948  &  n3949  &  n3950 ) ;
 assign Ng26947 = ( (~ n356) ) ;
 assign n359 = ( Ng518  &  Ng203  &  (~ Ng513) ) ;
 assign n357 = ( Ng182  &  Ng168 ) | ( Ng182  &  Ng174 ) ;
 assign n358 = ( Ng168  &  Ng174 ) ;
 assign Ng24210 = ( Pg35  &  n359  &  n357 ) | ( Pg35  &  n359  &  n358 ) ;
 assign n360 = ( Pg35  &  n2870 ) | ( n2870  &  (~ Ng3961) ) ;
 assign Ng30455 = ( (~ n360) ) ;
 assign n361 = ( n3847  &  n3849 ) | ( n3847  &  (~ Ng4749) ) | ( n3849  &  (~ n5625) ) | ( (~ Ng4749)  &  (~ n5625) ) ;
 assign Ng28084 = ( (~ n361) ) ;
 assign n362 = ( Pg35  &  n1844 ) | ( n1844  &  (~ Ng2089) ) ;
 assign Ng33993 = ( (~ n362) ) ;
 assign n363 = ( n2901  &  n2902  &  n160 ) | ( n2901  &  n2902  &  n2900 ) ;
 assign Ng30444 = ( (~ n363) ) ;
 assign n364 = ( (~ Ng1052)  &  n4004 ) | ( Ng1052  &  (~ n4004) ) ;
 assign Ng25625 = ( Pg35  &  n364  &  (~ Ng979) ) ;
 assign n366 = ( n1771  &  n2063  &  n2064 ) | ( n2063  &  n2064  &  (~ Ng2465) ) ;
 assign Ng33593 = ( (~ n366) ) ;
 assign n367 = ( n160  &  n2741  &  n2742 ) | ( n2741  &  n2742  &  n2740 ) ;
 assign Ng30502 = ( (~ n367) ) ;
 assign n368 = ( (~ n1245)  &  n2310  &  (~ n2521) ) | ( (~ n1245)  &  n2310  &  (~ Ng4480) ) ;
 assign Ng33036 = ( (~ n368) ) ;
 assign Ng25595 = ( Pg35  &  (~ Pg8719)  &  (~ Ng358) ) ;
 assign n371 = ( Pg35  &  n2344 ) | ( (~ Ng3171)  &  n2344 ) | ( Pg35  &  n2347 ) | ( (~ Ng3171)  &  n2347 ) ;
 assign Ng33024 = ( (~ n371) ) ;
 assign n372 = ( n1898  &  n2172 ) | ( n2172  &  (~ Ng1728) ) ;
 assign Ng33552 = ( (~ n372) ) ;
 assign n373 = ( Pg35  &  n1767 ) | ( n1767  &  (~ Ng2514) ) ;
 assign Ng34014 = ( (~ n373) ) ;
 assign n374 = ( Pg35  &  n3479 ) | ( (~ Ng3831)  &  n3479 ) ;
 assign Ng29273 = ( (~ n374) ) ;
 assign n375 = ( (~ Pg35) ) | ( (~ Ng4917) ) ;
 assign Ng34638 = ( (~ n375) ) ;
 assign n376 = ( Pg35  &  n330 ) | ( n330  &  (~ Ng1199) ) | ( Pg35  &  (~ n5341) ) | ( (~ Ng1199)  &  (~ n5341) ) ;
 assign Ng30341 = ( (~ n376) ) ;
 assign n377 = ( Pg35  &  n4036 ) | ( Pg35  &  n4037 ) | ( n4036  &  (~ Ng832) ) | ( n4037  &  (~ Ng832) ) ;
 assign Ng26899 = ( (~ n377) ) ;
 assign n378 = ( n3173  &  n3174  &  Ng914 ) | ( n3173  &  n3174  &  n3172 ) ;
 assign Ng30336 = ( (~ n378) ) ;
 assign n380 = ( Ng1008  &  n2207  &  (~ n6043) ) | ( n2207  &  n3160  &  (~ n6043) ) ;
 assign n379 = ( (~ n2207) ) | ( n4323 ) ;
 assign Ng25622 = ( Pg35  &  n380 ) | ( Pg35  &  Ng969  &  n379 ) ;
 assign n381 = ( n1596  &  n1591 ) | ( n1596  &  n1594 ) | ( n1596  &  n1595 ) ;
 assign Ng34447 = ( (~ n381) ) ;
 assign n382 = ( n2003  &  n2004  &  n2002 ) | ( n2003  &  n2004  &  (~ Ng4054) ) ;
 assign Ng33613 = ( (~ n382) ) ;
 assign n383 = ( Pg35  &  n4073 ) | ( n4073  &  (~ Ng6187) ) ;
 assign Ng25749 = ( (~ n383) ) ;
 assign Ng25704 = ( (~ Pg35)  &  Ng5073 ) | ( Ng5073  &  Ng5069 ) ;
 assign n384 = ( Pg35  &  n2276 ) | ( Pg35  &  n2277 ) | ( n2276  &  (~ Ng5517) ) | ( n2277  &  (~ Ng5517) ) ;
 assign Ng33053 = ( (~ n384) ) ;
 assign n385 = ( n160  &  n2592  &  n2593 ) | ( n2592  &  n2593  &  n2591 ) ;
 assign Ng30555 = ( (~ n385) ) ;
 assign n386 = ( n1925  &  n1923 ) | ( n1925  &  (~ Ng1682) ) ;
 assign Ng33971 = ( (~ n386) ) ;
 assign n387 = ( Ng1105  &  n4003  &  (~ n6435) ) | ( n4003  &  (~ n5092)  &  (~ n6435) ) ;
 assign Ng26915 = ( (~ n387) ) ;
 assign n388 = ( n160  &  n2638  &  n2639 ) | ( n2638  &  n2639  &  n2637 ) ;
 assign Ng30538 = ( (~ n388) ) ;
 assign n389 = ( Pg35  &  n3092  &  (~ n5857) ) | ( n3092  &  (~ Ng2250)  &  (~ n5857) ) ;
 assign Ng30369 = ( (~ n389) ) ;
 assign n390 = ( n1599  &  n1591 ) | ( n1599  &  n1597 ) | ( n1599  &  n1598 ) ;
 assign Ng34446 = ( (~ n390) ) ;
 assign n391 = ( n3782  &  n3783  &  Ng911 ) | ( n3782  &  n3783  &  (~ n4823) ) ;
 assign Ng29230 = ( (~ n391) ) ;
 assign n392 = ( (~ n1257)  &  n1909  &  n1910 ) | ( n1909  &  n1910  &  n1908 ) ;
 assign Ng33975 = ( (~ n392) ) ;
 assign n393 = ( n160  &  n2751  &  n2752 ) | ( n2751  &  n2752  &  n2750 ) ;
 assign Ng30497 = ( (~ n393) ) ;
 assign n394 = ( n2974  &  n2975  &  n160 ) | ( n2974  &  n2975  &  n2973 ) ;
 assign Ng30418 = ( (~ n394) ) ;
 assign n395 = ( Pg35  &  n4085 ) | ( n4085  &  (~ Ng5495) ) ;
 assign Ng25721 = ( (~ n395) ) ;
 assign n396 = ( Pg35  &  n1489 ) | ( n1489  &  (~ Ng2950) ) ;
 assign Ng34622 = ( (~ n396) ) ;
 assign n397 = ( n2919  &  n2920  &  n160 ) | ( n2919  &  n2920  &  n2918 ) ;
 assign Ng30438 = ( (~ n397) ) ;
 assign n398 = ( n160  &  n2632  &  n2633 ) | ( n2245  &  n2632  &  n2633 ) ;
 assign Ng30540 = ( (~ n398) ) ;
 assign n399 = ( Pg35  &  n2466  &  n2467 ) | ( (~ Ng1367)  &  n2466  &  n2467 ) ;
 assign Ng32986 = ( (~ n399) ) ;
 assign n400 = ( Pg35  &  n1952  &  n1953 ) | ( n1952  &  n1953  &  (~ Ng153) ) ;
 assign Ng33960 = ( (~ n400) ) ;
 assign n401 = ( n1609  &  n1604 ) | ( n1609  &  n1608 ) | ( n1609  &  n1598 ) ;
 assign Ng34442 = ( (~ n401) ) ;
 assign n402 = ( n2965  &  n2966  &  n160 ) | ( n2965  &  n2966  &  n2964 ) ;
 assign Ng30421 = ( (~ n402) ) ;
 assign n403 = ( Pg35  &  n2120 ) | ( n2120  &  (~ Ng2108) ) ;
 assign Ng33573 = ( (~ n403) ) ;
 assign n404 = ( Pg35  &  n4263 ) | ( n4263  &  (~ Ng437) ) ;
 assign Ng24205 = ( (~ n404) ) ;
 assign n405 = ( n2478  &  n2479  &  Ng758 ) | ( n2478  &  n2479  &  n2477 ) ;
 assign Ng32979 = ( (~ n405) ) ;
 assign n406 = ( Pg35  &  n4067 ) | ( n4067  &  (~ Ng6533) ) ;
 assign Ng25763 = ( (~ n406) ) ;
 assign n407 = ( n160  &  n2799  &  n2800 ) | ( n2799  &  n2800  &  n2798 ) ;
 assign Ng30481 = ( (~ n407) ) ;
 assign n408 = ( n160  &  n2696  &  (~ n6301) ) | ( n2696  &  n2695  &  (~ n6301) ) ;
 assign Ng30517 = ( (~ n408) ) ;
 assign n409 = ( n160  &  n2635  &  n2636 ) | ( n2635  &  n2636  &  n2634 ) ;
 assign Ng30539 = ( (~ n409) ) ;
 assign n410 = ( n1380  &  n1381  &  Ng632 ) | ( n1380  &  n1381  &  n1379 ) ;
 assign Ng34880 = ( (~ n410) ) ;
 assign n411 = ( n2925  &  n2926  &  n160 ) | ( n2925  &  n2926  &  n2924 ) ;
 assign Ng30436 = ( (~ n411) ) ;
 assign n412 = ( (~ Ng1664)  &  n2456  &  n2457 ) | ( n2452  &  n2456  &  n2457 ) ;
 assign Ng32990 = ( (~ n412) ) ;
 assign n413 = ( Pg35  &  n4235 ) | ( (~ wire4421)  &  n4235 ) ;
 assign Ng24245 = ( (~ n413) ) ;
 assign n414 = ( n160  &  n2598  &  n2599 ) | ( n2598  &  n2599  &  n2597 ) ;
 assign Ng30553 = ( (~ n414) ) ;
 assign n415 = ( Pg35  &  n4023 ) | ( n4023  &  (~ Ng269) ) ;
 assign Ng26907 = ( (~ n415) ) ;
 assign n416 = ( (~ Ng4040) ) | ( n5149 ) ;
 assign Ng24278 = ( (~ Pg35)  &  Ng4045 ) | ( Ng4045  &  n416 ) ;
 assign n417 = ( n3933  &  (~ Ng4438) ) | ( Pg35  &  n3933  &  (~ Ng4382) ) ;
 assign Ng26955 = ( (~ n417) ) ;
 assign n418 = ( Pg35  &  (~ Ng29277) ) | ( (~ wire4437)  &  (~ Ng29277) ) ;
 assign Ng29276 = ( (~ n418) ) ;
 assign n419 = ( Ng4681 ) | ( Ng4688 ) | ( Ng4674 ) | ( Ng4646 ) ;
 assign Ng29277 = ( Pg35  &  n419  &  (~ n5925) ) | ( Pg35  &  (~ n5350)  &  (~ n5925) ) ;
 assign n422 = ( (~ Pg35)  &  n1994  &  n2527 ) | ( n1994  &  n2527  &  n2526 ) ;
 assign Ng31894 = ( (~ n422) ) ;
 assign n423 = ( (~ n1245)  &  n2312  &  (~ n2521) ) | ( (~ n1245)  &  n2312  &  (~ Ng4495) ) ;
 assign Ng33037 = ( (~ n423) ) ;
 assign n424 = ( Pg35  &  n1579 ) | ( Pg35  &  n1584 ) | ( n1579  &  (~ Ng4332) ) | ( n1584  &  (~ Ng4332) ) ;
 assign Ng34451 = ( (~ n424) ) ;
 assign n425 = ( Pg35  &  n1689  &  n1690 ) | ( n1689  &  n1690  &  (~ Ng298) ) ;
 assign Ng34250 = ( (~ n425) ) ;
 assign n426 = ( (~ Ng5831)  &  n3296  &  (~ n5900) ) | ( n3296  &  n3295  &  (~ n5900) ) ;
 assign Ng29295 = ( (~ n426) ) ;
 assign n427 = ( Pg35  &  n4027 ) | ( n4027  &  (~ Ng262) ) ;
 assign Ng26905 = ( (~ n427) ) ;
 assign n428 = ( Pg35  &  n2472  &  n2473 ) | ( (~ Ng1024)  &  n2472  &  n2473 ) ;
 assign Ng32983 = ( (~ n428) ) ;
 assign n429 = ( n3017  &  n3018  &  n160 ) | ( n3017  &  n3018  &  n3016 ) ;
 assign Ng30402 = ( (~ n429) ) ;
 assign n430 = ( n1823  &  n1821 ) | ( n1823  &  (~ Ng2241) ) ;
 assign Ng33999 = ( (~ n430) ) ;
 assign n431 = ( n4220  &  n4221  &  Ng1564 ) | ( n4220  &  n4221  &  (~ n5130) ) ;
 assign Ng24262 = ( (~ n431) ) ;
 assign n432 = ( n160  &  n2583  &  n2584 ) | ( n2583  &  n2584  &  n2582 ) ;
 assign Ng30558 = ( (~ n432) ) ;
 assign n433 = ( Pg35  &  n4035 ) | ( n4035  &  (~ Ng872) ) ;
 assign Ng26901 = ( (~ n433) ) ;
 assign n434 = ( (~ n1248)  &  n2312  &  (~ n2521) ) | ( (~ n1248)  &  n2312  &  (~ Ng4501) ) ;
 assign Ng33039 = ( (~ n434) ) ;
 assign n435 = ( (~ Ng5869)  &  (~ Ng5873) ) | ( (~ Ng5873)  &  n2261 ) | ( (~ Ng5869)  &  n2263 ) | ( n2261  &  n2263 ) ;
 assign Ng33059 = ( (~ n435) ) ;
 assign n436 = ( n2509  &  n2517 ) | ( n2517  &  (~ Ng5037) ) | ( n2517  &  (~ n5328) ) ;
 assign Ng31899 = ( (~ n436) ) ;
 assign n437 = ( n2397  &  n2393  &  n2398 ) ;
 assign Ng33007 = ( (~ n437) ) ;
 assign n438 = ( n2851  &  n2852  &  n160 ) | ( n2851  &  n2852  &  n2850 ) ;
 assign Ng30462 = ( (~ n438) ) ;
 assign n439 = ( n160  &  n2781  &  n2782 ) | ( n2781  &  n2782  &  n2780 ) ;
 assign Ng30487 = ( (~ n439) ) ;
 assign n440 = ( Pg35  &  n2263 ) | ( Pg35  &  n2264 ) | ( n2263  &  (~ Ng5863) ) | ( n2264  &  (~ Ng5863) ) ;
 assign Ng33058 = ( (~ n440) ) ;
 assign n441 = ( Pg35  &  n4222 ) | ( (~ Ng1585)  &  n4222 ) ;
 assign Ng24261 = ( (~ n441) ) ;
 assign n442 = ( n160  &  n2659  &  n2660 ) | ( n2659  &  n2660  &  n2658 ) ;
 assign Ng30531 = ( (~ n442) ) ;
 assign n443 = ( n160  &  n2729  &  n2730 ) | ( n2729  &  n2730  &  n2728 ) ;
 assign Ng30506 = ( (~ n443) ) ;
 assign n444 = ( n4076  &  n4077  &  (~ n4894) ) | ( n4076  &  n4077  &  (~ Ng6167) ) ;
 assign Ng25747 = ( (~ n444) ) ;
 assign n445 = ( n1745  &  n2042  &  n2043 ) | ( n2042  &  n2043  &  (~ Ng2599) ) ;
 assign Ng33601 = ( (~ n445) ) ;
 assign n446 = ( Ng1448  &  n3983  &  (~ n6431) ) | ( n3983  &  (~ n5086)  &  (~ n6431) ) ;
 assign Ng26922 = ( (~ n446) ) ;
 assign n447 = ( n3685  &  n3686  &  (~ Ng2299) ) | ( n3685  &  n3686  &  (~ n4953) ) ;
 assign Ng29250 = ( (~ n447) ) ;
 assign Ng30459 = ( (~ n2289)  &  (~ Ng5164) ) ;
 assign n450 = ( Pg35  &  n2228  &  n2229 ) | ( n2228  &  n2229  &  (~ Ng150) ) ;
 assign Ng33534 = ( (~ n450) ) ;
 assign Ng30543 = ( (~ n2237)  &  (~ Ng6549) ) ;
 assign n453 = ( Pg35  &  n3473 ) | ( Pg35  &  n3474 ) | ( n3473  &  (~ Ng4076) ) | ( n3474  &  (~ Ng4076) ) ;
 assign Ng29275 = ( (~ n453) ) ;
 assign n454 = ( Pg35  &  n1731  &  n1732 ) | ( n1731  &  n1732  &  (~ Ng4793) ) ;
 assign Ng34030 = ( (~ n454) ) ;
 assign n455 = ( n2880  &  n2881  &  n160 ) | ( n2880  &  n2881  &  n2879 ) ;
 assign Ng30451 = ( (~ n455) ) ;
 assign n456 = ( n160  &  n2601  &  n2602 ) | ( n2601  &  n2602  &  n2600 ) ;
 assign Ng30552 = ( (~ n456) ) ;
 assign n457 = ( Pg35  &  n3170  &  n3171 ) | ( (~ Ng1002)  &  n3170  &  n3171 ) ;
 assign Ng30337 = ( (~ n457) ) ;
 assign n461 = ( Pg35  &  (~ n5152) ) | ( Pg35  &  (~ n854)  &  (~ n1218) ) ;
 assign Ng24254 = ( (~ Pg17423)  &  (~ Pg17404)  &  (~ Pg17320)  &  n461 ) ;
 assign n462 = ( Pg35  &  n3071  &  (~ n5848) ) | ( n3071  &  (~ Ng2441)  &  (~ n5848) ) ;
 assign Ng30378 = ( (~ n462) ) ;
 assign n463 = ( (~ Pg35)  &  n1736  &  n2358 ) | ( n1736  &  n2358  &  n2357 ) ;
 assign Ng33019 = ( (~ n463) ) ;
 assign n464 = ( Pg35  &  n1972 ) | ( n1972  &  (~ Ng6049) ) | ( Pg35  &  (~ n6118) ) | ( (~ Ng6049)  &  (~ n6118) ) ;
 assign Ng33623 = ( (~ n464) ) ;
 assign n465 = ( n3776  &  n3777  &  Ng1256 ) | ( n3776  &  n3777  &  (~ n4810) ) ;
 assign Ng29235 = ( (~ n465) ) ;
 assign n466 = ( n2503  &  n2507  &  n2508 ) | ( n2507  &  n2508  &  (~ Ng5016) ) ;
 assign Ng31902 = ( (~ n466) ) ;
 assign n467 = ( n1900  &  n1898 ) | ( n1900  &  (~ Ng1816) ) ;
 assign Ng33978 = ( (~ n467) ) ;
 assign n468 = ( Pg35  &  (~ Ng29279) ) | ( (~ Ng29279)  &  (~ Ng4572) ) ;
 assign Ng29278 = ( (~ n468) ) ;
 assign Ng34253 = ( Pg35  &  (~ Ng4462) ) | ( Pg35  &  (~ n1679) ) | ( Pg35  &  (~ Ng10384) ) ;
 assign n472 = ( (~ Ng3831)  &  n3481  &  (~ n5928) ) | ( n3481  &  n3480  &  (~ n5928) ) ;
 assign Ng29272 = ( (~ n472) ) ;
 assign n473 = ( Pg35  &  n2014 ) | ( n2014  &  (~ Ng3352) ) | ( Pg35  &  (~ n6120) ) | ( (~ Ng3352)  &  (~ n6120) ) ;
 assign Ng33610 = ( (~ n473) ) ;
 assign n474 = ( Pg35  &  n2078 ) | ( n2078  &  (~ Ng2399) ) ;
 assign Ng33589 = ( (~ n474) ) ;
 assign n475 = ( Pg35  &  n1518 ) | ( n1518  &  (~ Ng2138) ) ;
 assign Ng34605 = ( (~ n475) ) ;
 assign n476 = ( Pg35  &  n3137 ) | ( (~ Ng1696)  &  n3137 ) ;
 assign Ng30350 = ( (~ n476) ) ;
 assign n477 = ( n4180  &  n4190 ) | ( n4180  &  (~ Ng504) ) | ( n4190  &  (~ Ng513) ) | ( (~ Ng504)  &  (~ Ng513) ) ;
 assign Ng25611 = ( (~ n477) ) ;
 assign n478 = ( Pg35  &  n1984 ) | ( n1984  &  (~ Ng5357) ) | ( Pg35  &  (~ n6117) ) | ( (~ Ng5357)  &  (~ n6117) ) ;
 assign Ng33619 = ( (~ n478) ) ;
 assign n479 = ( n1736  &  n1737  &  Ng2763 ) | ( n1736  &  n1737  &  n1735 ) ;
 assign Ng34022 = ( (~ n479) ) ;
 assign n480 = ( Pg35  &  n1719 ) | ( Pg35  &  n1720 ) | ( n1719  &  (~ Ng4818) ) | ( n1720  &  (~ Ng4818) ) ;
 assign Ng34033 = ( (~ n480) ) ;
 assign n481 = ( n1433  &  n1435 ) ;
 assign Ng34726 = ( (~ n481) ) ;
 assign n482 = ( n2538  &  n2539  &  Ng1263 ) | ( n2538  &  n2539  &  (~ n4813) ) ;
 assign Ng31870 = ( (~ n482) ) ;
 assign n483 = ( n1875  &  n1873 ) | ( n1875  &  (~ Ng1950) ) ;
 assign Ng33985 = ( (~ n483) ) ;
 assign n484 = ( (~ Ng5138)  &  n3406  &  (~ n5916) ) | ( n3406  &  n3405  &  (~ n5916) ) ;
 assign Ng29283 = ( (~ n484) ) ;
 assign n485 = ( (~ n1273)  &  n1807  &  n1808 ) | ( n1807  &  n1808  &  n1806 ) ;
 assign Ng34003 = ( (~ n485) ) ;
 assign n486 = ( Pg35  &  n1542 ) | ( Pg35  &  n1543 ) | ( n1542  &  (~ Ng4659) ) | ( n1543  &  (~ Ng4659) ) ;
 assign Ng34463 = ( (~ n486) ) ;
 assign n487 = ( (~ Ng2223)  &  n2403  &  n2404 ) | ( n2399  &  n2403  &  n2404 ) ;
 assign Ng33006 = ( (~ n487) ) ;
 assign n488 = ( n3344  &  Ng5808  &  (~ n5905) ) | ( n3344  &  n3343  &  (~ n5905) ) ;
 assign Ng29292 = ( (~ n488) ) ;
 assign n489 = ( n160  &  n2586  &  n2587 ) | ( n2586  &  n2587  &  n2585 ) ;
 assign Ng30557 = ( (~ n489) ) ;
 assign n490 = ( (~ n1265)  &  n1858  &  n1859 ) | ( n1858  &  n1859  &  n1857 ) ;
 assign Ng33989 = ( (~ n490) ) ;
 assign n491 = ( (~ Ng3869)  &  (~ Ng3873) ) | ( (~ Ng3873)  &  n2323 ) | ( (~ Ng3869)  &  n2325 ) | ( n2323  &  n2325 ) ;
 assign Ng33033 = ( (~ n491) ) ;
 assign n492 = ( (~ n1273)  &  n1801  &  (~ n6218) ) | ( n1801  &  n1800  &  (~ n6218) ) ;
 assign Ng34005 = ( (~ n492) ) ;
 assign n493 = ( Pg35  &  n3961 ) | ( (~ Ng2799)  &  n3961 ) ;
 assign Ng26932 = ( (~ n493) ) ;
 assign n494 = ( n160  &  n2699  &  n2700 ) | ( n2699  &  n2700  &  n2698 ) ;
 assign Ng30516 = ( (~ n494) ) ;
 assign n495 = ( (~ Ng2047)  &  n2114  &  (~ n6132) ) | ( n2110  &  n2114  &  (~ n6132) ) ;
 assign Ng33575 = ( (~ n495) ) ;
 assign n496 = ( Pg35  &  n2325 ) | ( Pg35  &  n2326 ) | ( n2325  &  (~ Ng3863) ) | ( n2326  &  (~ Ng3863) ) ;
 assign Ng33032 = ( (~ n496) ) ;
 assign n497 = ( n160  &  n2784  &  n2785 ) | ( n2784  &  n2785  &  n2783 ) ;
 assign Ng30486 = ( (~ n497) ) ;
 assign n498 = ( n2913  &  n2914  &  n160 ) | ( n2913  &  n2914  &  n2912 ) ;
 assign Ng30440 = ( (~ n498) ) ;
 assign n499 = ( (~ Pg35)  &  n3942 ) | ( n3942  &  (~ Ng4411) ) | ( (~ Pg35)  &  (~ Ng4401) ) | ( (~ Ng4411)  &  (~ Ng4401) ) ;
 assign Ng26949 = ( (~ n499) ) ;
 assign n500 = ( n160  &  n2662  &  (~ n6290) ) | ( n2662  &  n2661  &  (~ n6290) ) ;
 assign Ng30530 = ( (~ n500) ) ;
 assign n501 = ( Pg35  &  n2628 ) | ( n2628  &  (~ Ng6307) ) ;
 assign Ng30542 = ( (~ n501) ) ;
 assign n502 = ( Pg35  &  n4156  &  n4157 ) | ( (~ Ng1036)  &  n4156  &  n4157 ) ;
 assign Ng25624 = ( (~ n502) ) ;
 assign n503 = ( Pg35  &  n3059  &  (~ n5843) ) | ( n3059  &  (~ Ng2575)  &  (~ n5843) ) ;
 assign Ng30383 = ( (~ n503) ) ;
 assign n504 = ( Pg35  &  n2057 ) | ( n2057  &  (~ Ng2533) ) ;
 assign Ng33597 = ( (~ n504) ) ;
 assign n505 = ( (~ Pg35)  &  n3925 ) | ( n3925  &  (~ Ng4443) ) | ( (~ Pg35)  &  (~ Ng4434) ) | ( (~ Ng4443)  &  (~ Ng4434) ) ;
 assign Ng26957 = ( (~ n505) ) ;
 assign n506 = ( Pg35  &  n3288  &  n3816 ) | ( n3288  &  n3816  &  (~ Ng6311) ) ;
 assign Ng28102 = ( (~ n506) ) ;
 assign n507 = ( n160  &  n2680  &  n2681 ) | ( n2680  &  n2681  &  n2679 ) ;
 assign Ng30524 = ( (~ n507) ) ;
 assign n508 = ( Pg35  &  n4031 ) | ( n4031  &  (~ Ng255) ) ;
 assign Ng26903 = ( (~ n508) ) ;
 assign n509 = ( n160  &  n2812  &  n2813 ) | ( n2812  &  n2813  &  n2811 ) ;
 assign Ng30475 = ( (~ n509) ) ;
 assign n510 = ( (~ Pg35) ) | ( (~ Ng6545) ) ;
 assign Ng34647 = ( (~ n510) ) ;
 assign n511 = ( (~ Ng2417)  &  n3074  &  (~ n5850) ) | ( n3074  &  n3072  &  (~ n5850) ) ;
 assign Ng30377 = ( (~ n511) ) ;
 assign n512 = ( n1898  &  n2168  &  n2169 ) | ( n2168  &  n2169  &  (~ Ng1772) ) ;
 assign Ng33553 = ( (~ n512) ) ;
 assign n513 = ( Pg35  &  n2501  &  (~ n5812) ) | ( n2501  &  (~ Ng5046)  &  (~ n5812) ) ;
 assign Ng31903 = ( (~ n513) ) ;
 assign n514 = ( (~ n1267)  &  n1878  &  n1879 ) | ( n1878  &  n1879  &  n1877 ) ;
 assign Ng33984 = ( (~ n514) ) ;
 assign n515 = ( n1745  &  n2037 ) | ( n1745  &  (~ Ng2599) ) | ( n2037  &  (~ Ng2629) ) | ( (~ Ng2599)  &  (~ Ng2629) ) ;
 assign Ng33602 = ( (~ n515) ) ;
 assign n516 = ( n3900  &  n3901  &  Ng572 ) | ( n3900  &  n3901  &  n3899 ) ;
 assign Ng28045 = ( (~ n516) ) ;
 assign n517 = ( (~ Pg35) ) | ( (~ Ng2130) ) ;
 assign Ng34603 = ( (~ n517) ) ;
 assign n518 = ( n1994  &  n2317  &  Ng4108 ) | ( n1994  &  n2317  &  n2316 ) ;
 assign Ng33035 = ( (~ n518) ) ;
 assign n519 = ( Pg35  &  n4261 ) | ( n4261  &  (~ Ng424) ) ;
 assign Ng24208 = ( (~ n519) ) ;
 assign n520 = ( Pg35  &  (~ Ng24212) ) | ( (~ Ng753)  &  (~ Ng24212) ) ;
 assign Ng24213 = ( (~ n520) ) ;
 assign n521 = ( Pg35  &  n1996 ) | ( n1996  &  (~ Ng4054) ) | ( Pg35  &  (~ n6114) ) | ( (~ Ng4054)  &  (~ n6114) ) ;
 assign Ng33614 = ( (~ n521) ) ;
 assign n522 = ( Pg35  &  n2256 ) | ( (~ Ng5873)  &  n2256 ) | ( Pg35  &  n2259 ) | ( (~ Ng5873)  &  n2259 ) ;
 assign Ng33060 = ( (~ n522) ) ;
 assign n523 = ( (~ Ng1992)  &  n3110  &  (~ n5865) ) | ( n3110  &  n3108  &  (~ n5865) ) ;
 assign Ng30362 = ( (~ n523) ) ;
 assign n524 = ( (~ Ng3167)  &  (~ Ng3171) ) | ( (~ Ng3171)  &  n2349 ) | ( (~ Ng3167)  &  n2351 ) | ( n2349  &  n2351 ) ;
 assign Ng33023 = ( (~ n524) ) ;
 assign n525 = ( Pg35  &  (~ Ng837) ) | ( (~ Ng837)  &  (~ Ng843) ) | ( Pg35  &  (~ n5392) ) | ( (~ Ng843)  &  (~ n5392) ) ;
 assign Ng26898 = ( (~ n525) ) ;
 assign n526 = ( (~ n3784)  &  n4169 ) | ( (~ n3784)  &  (~ Ng817) ) | ( n4169  &  (~ n5631) ) | ( (~ Ng817)  &  (~ n5631) ) ;
 assign Ng25618 = ( (~ n526) ) ;
 assign n527 = ( n160  &  n2693  &  n2694 ) | ( n2693  &  n2694  &  n2692 ) ;
 assign Ng30518 = ( (~ n527) ) ;
 assign n528 = ( n4058  &  n4063 ) | ( n4063  &  n4061  &  (~ Ng26885) ) ;
 assign Ng26884 = ( (~ n528) ) ;
 assign n529 = ( Pg35  &  n3959 ) | ( (~ Ng2811)  &  n3959 ) ;
 assign Ng26933 = ( (~ n529) ) ;
 assign n530 = ( Pg35  &  n3580  &  n3870 ) | ( n3580  &  n3870  &  (~ Ng3614) ) ;
 assign Ng28066 = ( (~ n530) ) ;
 assign n531 = ( Pg35  &  n2005 ) | ( n2005  &  (~ Ng3703) ) | ( Pg35  &  (~ n6119) ) | ( (~ Ng3703)  &  (~ n6119) ) ;
 assign Ng33612 = ( (~ n531) ) ;
 assign n532 = ( Pg35  &  n4025 ) | ( n4025  &  (~ Ng239) ) ;
 assign Ng26906 = ( (~ n532) ) ;
 assign n533 = ( n3529  &  Ng3808  &  (~ n5933) ) | ( n3529  &  n3528  &  (~ n5933) ) ;
 assign Ng29269 = ( (~ n533) ) ;
 assign n534 = ( Ng10384  &  Ng4473 ) ;
 assign Ng34255 = ( (~ Pg35) ) | ( n534 ) | ( Ng4462 ) | ( (~ n1679) ) ;
 assign n535 = ( n2883  &  n2884  &  n160 ) | ( n2883  &  n2884  &  n2882 ) ;
 assign Ng30450 = ( (~ n535) ) ;
 assign n536 = ( Pg35  &  n2867  &  n2868 ) | ( (~ Ng4087)  &  n2867  &  n2868 ) ;
 assign Ng30456 = ( (~ n536) ) ;
 assign n537 = ( n2450  &  n2446  &  n2451 ) ;
 assign Ng32991 = ( (~ n537) ) ;
 assign n541 = ( (~ Pg17760)  &  (~ Pg14779) ) | ( (~ Pg17760)  &  Pg12422 ) | ( Pg14779  &  Pg12422 ) ;
 assign Ng24348 = ( Pg35  &  (~ Pg17685)  &  (~ Pg17649)  &  (~ Pg13085)  &  n541 ) ;
 assign n542 = ( Pg35  &  n1693  &  n1694 ) | ( n1693  &  n1694  &  (~ Ng157) ) ;
 assign Ng34249 = ( (~ n542) ) ;
 assign n543 = ( n3532  &  n160 ) | ( n3532  &  Ng3498  &  n3531 ) ;
 assign Ng29268 = ( (~ n543) ) ;
 assign n544 = ( n3806  &  n3807  &  Ng586 ) | ( n3806  &  n3807  &  n3805 ) ;
 assign Ng29224 = ( (~ n544) ) ;
 assign n545 = ( n2361  &  n2366  &  n2367 ) | ( n2366  &  n2367  &  (~ Ng2619) ) ;
 assign Ng33017 = ( (~ n545) ) ;
 assign n546 = ( n3168  &  Ng1183 ) | ( n3168  &  n3167 ) ;
 assign Ng30339 = ( (~ n546) ) ;
 assign n547 = ( (~ n1271)  &  n1937  &  n1938 ) | ( n1937  &  n1938  &  n1936 ) ;
 assign Ng33967 = ( (~ n547) ) ;
 assign n548 = ( (~ Ng1779)  &  n2156  &  (~ n6134) ) | ( n2152  &  n2156  &  (~ n6134) ) ;
 assign Ng33559 = ( (~ n548) ) ;
 assign n549 = ( (~ Pg35)  &  (~ n3639) ) | ( n3636  &  (~ n3639) ) | ( (~ n3639)  &  (~ Ng2652) ) ;
 assign Ng29255 = ( (~ n549) ) ;
 assign n550 = ( Pg35  &  n3095  &  (~ n5858) ) | ( n3095  &  (~ Ng2173)  &  (~ n5858) ) ;
 assign Ng30368 = ( (~ n550) ) ;
 assign n551 = ( Pg35  &  n3077 ) | ( (~ Ng2389)  &  n3077 ) ;
 assign Ng30375 = ( (~ n551) ) ;
 assign n552 = ( (~ Pg35)  &  n3829 ) | ( n3825  &  n3829 ) | ( n3829  &  n3828 ) ;
 assign Ng28089 = ( (~ n552) ) ;
 assign n553 = ( Pg35  &  n2269 ) | ( (~ Ng5527)  &  n2269 ) | ( Pg35  &  n2272 ) | ( (~ Ng5527)  &  n2272 ) ;
 assign Ng33055 = ( (~ n553) ) ;
 assign n554 = ( Pg35  &  n3043 ) | ( n3043  &  (~ Ng2803) ) ;
 assign Ng30392 = ( (~ n554) ) ;
 assign n555 = ( Pg35  &  n3154  &  n3155 ) | ( (~ Ng1345)  &  n3154  &  n3155 ) ;
 assign Ng30343 = ( (~ n555) ) ;
 assign n556 = ( n160  &  n2683  &  n2684 ) | ( n2683  &  n2684  &  n2682 ) ;
 assign Ng30523 = ( (~ n556) ) ;
 assign n559 = ( (~ n557)  &  Ng1146 ) | ( Ng1146  &  (~ Ng1152) ) ;
 assign n557 = ( Pg13259  &  (~ Ng1171)  &  (~ Ng1183) ) ;
 assign Ng24233 = ( Pg35  &  n559 ) | ( Pg35  &  n557  &  (~ Ng1099) ) ;
 assign n560 = ( (~ Ng2625)  &  n2363  &  n2364 ) | ( n2359  &  n2363  &  n2364 ) ;
 assign Ng33018 = ( (~ n560) ) ;
 assign n561 = ( Pg35  &  n2487  &  n2488 ) | ( n2487  &  n2488  &  (~ Ng164) ) ;
 assign Ng32976 = ( (~ n561) ) ;
 assign n562 = ( Pg35  &  n3140  &  (~ n5877) ) | ( n3140  &  (~ Ng1691)  &  (~ n5877) ) ;
 assign Ng30349 = ( (~ n562) ) ;
 assign n563 = ( Pg35  &  n2233 ) | ( Pg35  &  n2240 ) | ( n2233  &  (~ Ng6549) ) | ( n2240  &  (~ Ng6549) ) ;
 assign Ng33067 = ( (~ n563) ) ;
 assign Ng26900 = ( wire4431  &  Pg35 ) ;
 assign n564 = ( Pg35  &  n2318 ) | ( (~ Ng3873)  &  n2318 ) | ( Pg35  &  n2321 ) | ( (~ Ng3873)  &  n2321 ) ;
 assign Ng33034 = ( (~ n564) ) ;
 assign n565 = ( n160  &  n2604  &  n2605 ) | ( n2604  &  n2605  &  n2603 ) ;
 assign Ng30551 = ( (~ n565) ) ;
 assign n566 = ( n4126  &  n4127  &  (~ n4928) ) | ( n4126  &  n4127  &  (~ Ng3470) ) ;
 assign Ng25667 = ( (~ n566) ) ;
 assign n567 = ( n2877  &  n2878  &  n160 ) | ( n2877  &  n2878  &  n2876 ) ;
 assign Ng30452 = ( (~ n567) ) ;
 assign n568 = ( n4180  &  n4190 ) | ( n4190  &  (~ Ng518) ) | ( n4180  &  (~ Ng513) ) | ( (~ Ng518)  &  (~ Ng513) ) ;
 assign Ng25612 = ( (~ n568) ) ;
 assign n571 = ( Ng538 ) | ( Ng209 ) ;
 assign n569 = ( n1335  &  n1336  &  n1337  &  n1338 ) ;
 assign Ng34719 = ( n571  &  Pg35 ) ;
 assign n572 = ( (~ Ng2606)  &  n2030  &  (~ n6128) ) | ( n2025  &  n2030  &  (~ n6128) ) ;
 assign Ng33607 = ( (~ n572) ) ;
 assign n573 = ( Ng1472  &  n3979  &  n3980 ) | ( n3979  &  n3980  &  (~ n5085) ) ;
 assign Ng26923 = ( (~ n573) ) ;
 assign n574 = ( Pg35  &  n3791 ) | ( Pg35  &  n4256 ) | ( n3791  &  (~ Ng546) ) | ( n4256  &  (~ Ng546) ) ;
 assign Ng24211 = ( (~ n574) ) ;
 assign n575 = ( Pg35  &  n2282 ) | ( (~ Ng5180)  &  n2282 ) | ( Pg35  &  n2285 ) | ( (~ Ng5180)  &  n2285 ) ;
 assign Ng33050 = ( (~ n575) ) ;
 assign n576 = ( n2848  &  n2849  &  n160 ) | ( n2848  &  n2849  &  n2847 ) ;
 assign Ng30463 = ( (~ n576) ) ;
 assign n577 = ( n1541  &  n1540 ) | ( n1541  &  (~ Ng4664) ) | ( n1541  &  (~ n4633) ) ;
 assign Ng34464 = ( (~ n577) ) ;
 assign n578 = ( Pg35  &  n4235 ) | ( n4235  &  (~ Ng1236) ) ;
 assign Ng24243 = ( (~ n578) ) ;
 assign n579 = ( Pg35  &  n4204 ) | ( (~ wire4507)  &  n4204 ) | ( Pg35  &  n4205 ) | ( (~ wire4507)  &  n4205 ) ;
 assign Ng24335 = ( (~ n579) ) ;
 assign n580 = ( Pg35  &  n1508 ) | ( n1508  &  (~ Ng2852) ) ;
 assign Ng34611 = ( (~ n580) ) ;
 assign n581 = ( n1669  &  n1670  &  n1668 ) | ( n1669  &  n1670  &  n1666 ) ;
 assign Ng34262 = ( (~ n581) ) ;
 assign n582 = ( n160  &  n2619  &  n2620 ) | ( n2619  &  n2620  &  n2618 ) ;
 assign Ng30546 = ( (~ n582) ) ;
 assign n583 = ( Pg35  &  n923 ) | ( n923  &  (~ Ng1542) ) | ( Pg35  &  (~ n5339) ) | ( (~ Ng1542)  &  (~ n5339) ) ;
 assign Ng30347 = ( (~ n583) ) ;
 assign n584 = ( n160  &  n2589  &  n2590 ) | ( n2589  &  n2590  &  n2588 ) ;
 assign Ng30556 = ( (~ n584) ) ;
 assign n585 = ( n1873  &  n2142 ) | ( n1873  &  (~ Ng1906) ) | ( n2142  &  (~ Ng1936) ) | ( (~ Ng1906)  &  (~ Ng1936) ) ;
 assign Ng33562 = ( (~ n585) ) ;
 assign n586 = ( n4196  &  n4192 ) | ( n4196  &  n3809 ) ;
 assign Ng25610 = ( (~ n586) ) ;
 assign n587 = ( n2370  &  n2366  &  n2371 ) ;
 assign Ng33015 = ( (~ n587) ) ;
 assign n588 = ( Pg35  &  n2312  &  n2520 ) | ( n2312  &  n2520  &  (~ Ng4477) ) ;
 assign Ng31896 = ( (~ n588) ) ;
 assign n589 = ( (~ n1273)  &  n1804  &  n1805 ) | ( n1804  &  n1805  &  (~ n4723) ) ;
 assign Ng34004 = ( (~ n589) ) ;
 assign n590 = ( n160  &  n2944  &  (~ n6383) ) | ( n2944  &  n2943  &  (~ n6383) ) ;
 assign Ng30428 = ( (~ n590) ) ;
 assign n591 = ( n160  &  n2787  &  n2788 ) | ( n2787  &  n2788  &  n2786 ) ;
 assign Ng30485 = ( (~ n591) ) ;
 assign n592 = ( n160  &  n2962  &  (~ n6389) ) | ( n2962  &  n2961  &  (~ n6389) ) ;
 assign Ng30422 = ( (~ n592) ) ;
 assign n593 = ( n2959  &  n2960  &  n160 ) | ( n2959  &  n2960  &  n2958 ) ;
 assign Ng30423 = ( (~ n593) ) ;
 assign n594 = ( n160  &  n2665  &  n2666 ) | ( n2665  &  n2666  &  n2664 ) ;
 assign Ng30529 = ( (~ n594) ) ;
 assign Ng34028 = ( Ng4681  &  n270 ) ;
 assign n595 = ( n2857  &  n2858  &  n160 ) | ( n2857  &  n2858  &  n2856 ) ;
 assign Ng30460 = ( (~ n595) ) ;
 assign n596 = ( n160  &  n3020  &  (~ n6408) ) | ( n3020  &  n3019  &  (~ n6408) ) ;
 assign Ng30401 = ( (~ n596) ) ;
 assign n597 = ( (~ n1265)  &  n1855  &  n1856 ) | ( n1855  &  n1856  &  (~ n4745) ) ;
 assign Ng33990 = ( (~ n597) ) ;
 assign n598 = ( n3185  &  n160 ) | ( n3185  &  Ng6541  &  n3184 ) ;
 assign Ng29309 = ( (~ n598) ) ;
 assign n599 = ( n2990  &  n2991  &  n160 ) | ( n2990  &  n2991  &  n2346 ) ;
 assign Ng30411 = ( (~ n599) ) ;
 assign n600 = ( Pg35  &  n2185 ) | ( n2185  &  (~ Ng1636) ) ;
 assign Ng33546 = ( (~ n600) ) ;
 assign n601 = ( (~ Pg35)  &  n3846 ) | ( n3842  &  n3846 ) | ( n3846  &  n3845 ) ;
 assign Ng28085 = ( (~ n601) ) ;
 assign n602 = ( Pg35  &  n4029 ) | ( n4029  &  (~ Ng232) ) ;
 assign Ng26904 = ( (~ n602) ) ;
 assign n603 = ( Pg35  &  n4198 ) | ( (~ Ng168)  &  n4198 ) ;
 assign Ng25605 = ( (~ n603) ) ;
 assign n604 = ( Pg35  &  n2246 ) | ( Pg35  &  n2253 ) | ( n2246  &  (~ Ng6203) ) | ( n2253  &  (~ Ng6203) ) ;
 assign Ng33062 = ( (~ n604) ) ;
 assign n605 = ( Pg35  &  n4049 ) | ( Pg35  &  n4052 ) | ( n4049  &  (~ Ng355) ) | ( n4052  &  (~ Ng355) ) ;
 assign Ng26893 = ( (~ n605) ) ;
 assign n606 = ( (~ Pg35) ) | ( (~ Ng3502) ) ;
 assign Ng34626 = ( (~ n606) ) ;
 assign n607 = ( (~ Ng2204)  &  n2093  &  (~ n6131) ) | ( n2089  &  n2093  &  (~ n6131) ) ;
 assign Ng33583 = ( (~ n607) ) ;
 assign n608 = ( n160  &  n2821  &  n2822 ) | ( n2821  &  n2822  &  n2820 ) ;
 assign Ng30472 = ( (~ n608) ) ;
 assign n609 = ( Pg35  &  n1576  &  n1577 ) | ( n1576  &  n1577  &  (~ Ng4601) ) ;
 assign Ng34454 = ( (~ n609) ) ;
 assign n610 = ( n1396  &  n1397  &  Ng794 ) | ( n1396  &  n1397  &  n1395 ) ;
 assign Ng34850 = ( (~ n610) ) ;
 assign n611 = ( (~ Ng703)  &  n4253 ) | ( n4251  &  n4253 ) ;
 assign Ng24214 = ( (~ n611) ) ;
 assign n612 = ( n3005  &  n3006  &  n160 ) | ( n3005  &  n3006  &  n3004 ) ;
 assign Ng30406 = ( (~ n612) ) ;
 assign n613 = ( n1847  &  n2126  &  n2127 ) | ( n2126  &  n2127  &  (~ Ng2040) ) ;
 assign Ng33569 = ( (~ n613) ) ;
 assign n614 = ( Pg35  &  n1480 ) | ( n1480  &  (~ Ng4176) ) ;
 assign Ng34628 = ( (~ n614) ) ;
 assign n615 = ( (~ Ng4633)  &  (~ Ng4628) ) | ( (~ Ng4628)  &  n1558 ) | ( (~ Ng4633)  &  n1559 ) | ( n1558  &  n1559 ) ;
 assign Ng34458 = ( (~ n615) ) ;
 assign n616 = ( Pg35  &  n1468 ) | ( n1468  &  (~ Ng4727) ) ;
 assign Ng34634 = ( (~ n616) ) ;
 assign n617 = ( (~ n2562)  &  n3300  &  (~ n5902) ) | ( n3300  &  (~ n4998)  &  (~ n5902) ) ;
 assign Ng29293 = ( (~ n617) ) ;
 assign n618 = ( n2388  &  n2393  &  n2394 ) | ( n2393  &  n2394  &  (~ Ng2351) ) ;
 assign Ng33009 = ( (~ n618) ) ;
 assign n619 = ( (~ Ng6727) ) | ( (~ n5140) ) ;
 assign Ng24355 = ( (~ Pg35)  &  Ng6732 ) | ( Ng6732  &  n619 ) ;
 assign n620 = ( Pg35  &  n1994 ) | ( Pg35  &  n4107 ) | ( n1994  &  (~ Ng4125) ) | ( n4107  &  (~ Ng4125) ) ;
 assign Ng25691 = ( (~ n620) ) ;
 assign n621 = ( n3539  &  (~ n4345)  &  (~ n5938) ) | ( n3539  &  (~ n5030)  &  (~ n5938) ) ;
 assign Ng29264 = ( (~ n621) ) ;
 assign n622 = ( n3860  &  n3865  &  n3866 ) | ( n3865  &  n3866  &  (~ n5071) ) ;
 assign Ng28072 = ( (~ n622) ) ;
 assign n623 = ( n2509  &  n2514 ) | ( n2514  &  (~ Ng5041) ) | ( n2514  &  (~ n4883) ) ;
 assign Ng31900 = ( (~ n623) ) ;
 assign n624 = ( n3926  &  (~ Ng4452) ) | ( n3929  &  (~ Ng4452) ) | ( (~ Ng4452)  &  (~ Ng4430) ) ;
 assign Ng26956 = ( (~ n624) ) ;
 assign n625 = ( n3236  &  Ng6500  &  (~ n5888) ) | ( n3236  &  n3235  &  (~ n5888) ) ;
 assign Ng29304 = ( (~ n625) ) ;
 assign n626 = ( Pg35  &  n3585 ) | ( n3585  &  (~ Ng3129) ) ;
 assign Ng29261 = ( (~ n626) ) ;
 assign n627 = ( Pg35  &  n3871 ) | ( n3871  &  (~ Ng3263) ) ;
 assign Ng28063 = ( (~ n627) ) ;
 assign Ng34027 = ( Ng4674  &  n270 ) ;
 assign n628 = ( Pg35  &  n1949  &  n1950 ) | ( n1949  &  n1950  &  (~ Ng294) ) ;
 assign Ng33961 = ( (~ n628) ) ;
 assign n629 = ( n2437  &  n2433  &  n2438 ) ;
 assign Ng32995 = ( (~ n629) ) ;
 assign n630 = ( Pg35  &  n1485 ) | ( n1485  &  (~ Ng2994) ) ;
 assign Ng34624 = ( (~ n630) ) ;
 assign n631 = ( n2983  &  n2984  &  n160 ) | ( n2983  &  n2984  &  n2982 ) ;
 assign Ng30415 = ( (~ n631) ) ;
 assign Ng33536 = ( (~ Pg35)  &  Ng160 ) | ( Ng160  &  (~ n5754) ) ;
 assign n633 = ( Pg35  &  n3887  &  n3888 ) | ( n3887  &  n3888  &  (~ Ng822) ) ;
 assign Ng28055 = ( (~ n633) ) ;
 assign n634 = ( (~ Ng969)  &  (~ n379)  &  (~ Ng1008) ) ;
 assign Ng24238 = ( Pg35  &  n634  &  (~ n5635) ) | ( Pg35  &  (~ n5154)  &  (~ n5635) ) ;
 assign n637 = ( n1745  &  n2046 ) | ( n2046  &  (~ Ng2555) ) ;
 assign Ng33600 = ( (~ n637) ) ;
 assign n638 = ( Pg35  &  n3235  &  n3815 ) | ( n3235  &  n3815  &  (~ Ng6657) ) ;
 assign Ng28105 = ( (~ n638) ) ;
 assign n639 = ( (~ Ng6523)  &  n3189  &  (~ n5883) ) | ( n3189  &  n3188  &  (~ n5883) ) ;
 assign Ng29307 = ( (~ n639) ) ;
 assign n640 = ( n3152  &  Ng1526 ) | ( n3152  &  n3151 ) ;
 assign Ng30345 = ( (~ n640) ) ;
 assign n641 = ( Pg35  &  n1578 ) | ( Pg35  &  n1579 ) | ( n1578  &  (~ Ng4593) ) | ( n1579  &  (~ Ng4593) ) ;
 assign Ng34453 = ( (~ n641) ) ;
 assign n644 = ( (~ n642) ) | ( Ng854 ) ;
 assign n642 = ( (~ Pg8719) ) | ( Ng385 ) | ( (~ Ng376) ) | ( (~ Ng370) ) ;
 assign n643 = ( n1612 ) | ( (~ n5984) ) ;
 assign Ng32980 = ( n644  &  Pg35  &  n642 ) | ( n644  &  Pg35  &  n643 ) ;
 assign n645 = ( n3774  &  n3772 ) | ( n3774  &  (~ Ng1484) ) ;
 assign Ng29238 = ( (~ n645) ) ;
 assign n646 = ( Pg35  &  n1458 ) | ( n1458  &  (~ Ng4917) ) ;
 assign Ng34639 = ( (~ n646) ) ;
 assign Ng25695 = ( (~ Pg35)  &  Ng5077 ) | ( Ng5077  &  (~ n5450) ) ;
 assign n648 = ( Pg35  &  n2259 ) | ( Pg35  &  n2266 ) | ( n2259  &  (~ Ng5857) ) | ( n2266  &  (~ Ng5857) ) ;
 assign Ng33057 = ( (~ n648) ) ;
 assign n649 = ( (~ Pg35)  &  (~ n3656) ) | ( n3653  &  (~ n3656) ) | ( (~ n3656)  &  (~ Ng2518) ) ;
 assign Ng29253 = ( (~ n649) ) ;
 assign n650 = ( Pg35  &  n1742 ) | ( n1742  &  (~ Ng2648) ) ;
 assign Ng34021 = ( (~ n650) ) ;
 assign n651 = ( n4047  &  n4048  &  Ng568 ) | ( n4047  &  n4048  &  n4046 ) ;
 assign Ng26895 = ( (~ n651) ) ;
 assign n652 = ( Pg35  &  n2986 ) | ( n2986  &  (~ Ng3259) ) ;
 assign Ng30413 = ( (~ n652) ) ;
 assign n653 = ( n160  &  n2610  &  n2611 ) | ( n2610  &  n2611  &  n2609 ) ;
 assign Ng30549 = ( (~ n653) ) ;
 assign n654 = ( (~ Ng6035) ) | ( (~ n5143) ) ;
 assign Ng24347 = ( (~ Pg35)  &  Ng6040 ) | ( Ng6040  &  n654 ) ;
 assign Ng30501 = ( (~ n2263)  &  (~ Ng5857) ) ;
 assign n657 = ( (~ n1271)  &  n1931  &  n1932 ) | ( n1931  &  n1932  &  n1930 ) ;
 assign Ng33969 = ( (~ n657) ) ;
 assign n658 = ( n2930  &  n2931  &  n160 ) | ( n2930  &  n2931  &  n2929 ) ;
 assign Ng30433 = ( (~ n658) ) ;
 assign n659 = ( (~ n2564)  &  n3485  &  (~ n5930) ) | ( n3485  &  (~ n5023)  &  (~ n5930) ) ;
 assign Ng29270 = ( (~ n659) ) ;
 assign n660 = ( (~ n1248)  &  n2310  &  (~ n2521) ) | ( (~ n1248)  &  n2310  &  (~ Ng4498) ) ;
 assign Ng33038 = ( (~ n660) ) ;
 assign n661 = ( Pg35  &  n3973  &  n3974 ) | ( n3973  &  n3974  &  (~ Ng2719) ) ;
 assign Ng26926 = ( (~ n661) ) ;
 assign n662 = ( (~ Pg35)  &  n3854 ) | ( n3850  &  n3854 ) | ( n3854  &  n3853 ) ;
 assign Ng28083 = ( (~ n662) ) ;
 assign n663 = ( n160  &  n2804  &  n2805 ) | ( n2804  &  n2805  &  n2803 ) ;
 assign Ng30478 = ( (~ n663) ) ;
 assign n664 = ( n1440  &  n1441  &  Ng617 ) | ( n1440  &  n1441  &  n1439 ) ;
 assign Ng34724 = ( (~ n664) ) ;
 assign n665 = ( Pg35  &  n4058 ) | ( n4058  &  (~ Ng324) ) ;
 assign Ng26883 = ( (~ n665) ) ;
 assign n666 = ( Ng1270  &  (~ n2468) ) ;
 assign n667 = ( (~ n1218) ) | ( (~ Ng1536) ) ;
 assign Ng32985 = ( (~ Pg35)  &  Ng1274 ) | ( Ng1274  &  n666  &  n667 ) ;
 assign n668 = ( n4070  &  n4071  &  (~ n4886) ) | ( n4070  &  n4071  &  (~ Ng6513) ) ;
 assign Ng25761 = ( (~ n668) ) ;
 assign n669 = ( n4059  &  n4060  &  n4058 ) | ( n4059  &  n4060  &  (~ Ng305) ) ;
 assign Ng26886 = ( (~ n669) ) ;
 assign n670 = ( Ng925  &  (~ n2474) ) ;
 assign Ng32982 = ( (~ Pg35)  &  Ng930 ) | ( Ng930  &  n670  &  (~ n1411) ) ;
 assign n672 = ( n1873  &  n2147  &  n2148 ) | ( n2147  &  n2148  &  (~ Ng1906) ) ;
 assign Ng33561 = ( (~ n672) ) ;
 assign Ng26880 = ( Pg6745  &  Pg35 ) ;
 assign n673 = ( Pg35  &  n3963 ) | ( (~ wire4428)  &  n3963 ) ;
 assign Ng26931 = ( (~ n673) ) ;
 assign n674 = ( Pg35  &  n1454 ) | ( n1454  &  (~ Ng4907) ) ;
 assign Ng34641 = ( (~ n674) ) ;
 assign n675 = ( Pg35  &  n1478 ) | ( n1478  &  (~ Ng4146) ) ;
 assign Ng34629 = ( (~ n675) ) ;
 assign n676 = ( n2054  &  n2055  &  (~ n4709) ) | ( n2054  &  n2055  &  (~ Ng2541) ) ;
 assign Ng33598 = ( (~ n676) ) ;
 assign n677 = ( n1821  &  n2109 ) | ( n2109  &  (~ Ng2153) ) ;
 assign Ng33576 = ( (~ n677) ) ;
 assign n678 = ( Pg35  &  n4033 ) | ( n4033  &  (~ Ng225) ) ;
 assign Ng26902 = ( (~ n678) ) ;
 assign n679 = ( n3736  &  n3737  &  (~ Ng1874) ) | ( n3736  &  n3737  &  (~ n4963) ) ;
 assign Ng29244 = ( (~ n679) ) ;
 assign n680 = ( n2833  &  n2834  &  n160 ) | ( n2833  &  n2834  &  n2832 ) ;
 assign Ng30468 = ( (~ n680) ) ;
 assign n681 = ( Ng1478  &  n3976  &  n3977 ) | ( n3976  &  n3977  &  (~ n5084) ) ;
 assign Ng26924 = ( (~ n681) ) ;
 assign n682 = ( Pg35  &  n2321 ) | ( Pg35  &  n2328 ) | ( n2321  &  (~ Ng3857) ) | ( n2328  &  (~ Ng3857) ) ;
 assign Ng33031 = ( (~ n682) ) ;
 assign n683 = ( (~ Pg35)  &  (~ n3724) ) | ( n3721  &  (~ n3724) ) | ( (~ n3724)  &  (~ Ng1959) ) ;
 assign Ng29245 = ( (~ n683) ) ;
 assign n684 = ( (~ Ng3480)  &  n3536  &  (~ n5936) ) | ( n3536  &  n3535  &  (~ n5936) ) ;
 assign Ng29266 = ( (~ n684) ) ;
 assign n685 = ( n160  &  n2580  &  (~ n6263) ) | ( n2580  &  n2579  &  (~ n6263) ) ;
 assign Ng30559 = ( (~ n685) ) ;
 assign n686 = ( (~ Pg35)  &  n3836 ) | ( n1407  &  n3836 ) | ( n3833  &  n3836 ) ;
 assign Ng28087 = ( (~ n686) ) ;
 assign Ng30435 = ( (~ n2325)  &  (~ Ng3857) ) ;
 assign n689 = ( n4192  &  Ng499 ) | ( Ng499  &  (~ Ng513) ) ;
 assign n690 = ( (~ n4192)  &  (~ Ng518) ) | ( (~ n4192)  &  (~ n5056) ) ;
 assign Ng25609 = ( Pg35  &  n689 ) | ( Pg35  &  n690 ) ;
 assign n691 = ( (~ n2207)  &  n3882 ) | ( Ng1002  &  n3882 ) | ( n3882  &  n3881 ) ;
 assign Ng28057 = ( (~ n691) ) ;
 assign n692 = ( n1627  &  n1628  &  Ng776 ) | ( n1627  &  n1628  &  n1626 ) ;
 assign Ng34439 = ( (~ n692) ) ;
 assign Ng34260 = ( (~ Ng4646)  &  (~ Ng4681)  &  (~ Ng4674)  &  (~ n1543) ) ;
 assign n697 = ( n2454  &  n2459  &  n2460 ) | ( n2459  &  n2460  &  (~ Ng1657) ) ;
 assign Ng32989 = ( (~ n697) ) ;
 assign n698 = ( n1798  &  n1796 ) | ( n1798  &  (~ Ng2375) ) ;
 assign Ng34006 = ( (~ n698) ) ;
 assign n699 = ( Pg35  &  Ng283 ) | ( (~ Ng278)  &  Ng283 ) | ( Pg35  &  n3904 ) | ( (~ Ng278)  &  n3904 ) ;
 assign Ng28043 = ( (~ n699) ) ;
 assign n700 = ( Pg35  &  n2347 ) | ( Pg35  &  n2354 ) | ( n2347  &  (~ Ng3155) ) | ( n2354  &  (~ Ng3155) ) ;
 assign Ng33021 = ( (~ n700) ) ;
 assign n701 = ( (~ Pg35)  &  (~ n3673) ) | ( n3670  &  (~ n3673) ) | ( (~ n3673)  &  (~ Ng2384) ) ;
 assign Ng29251 = ( (~ n701) ) ;
 assign n702 = ( (~ n1564)  &  n1570 ) | ( n1570  &  n1569 ) | ( n1570  &  (~ Ng4608) ) ;
 assign Ng34456 = ( (~ n702) ) ;
 assign n703 = ( (~ n1265)  &  n1852  &  n1853 ) | ( n1852  &  n1853  &  n1851 ) ;
 assign Ng33991 = ( (~ n703) ) ;
 assign n704 = ( Pg35  &  n3965 ) | ( (~ Ng2791)  &  n3965 ) ;
 assign Ng26930 = ( (~ n704) ) ;
 assign n705 = ( n1525  &  n1526  &  Ng613 ) | ( n1525  &  n1526  &  n1524 ) ;
 assign Ng34599 = ( (~ n705) ) ;
 assign n706 = ( Pg35  &  n2162 ) | ( n2162  &  (~ Ng1840) ) ;
 assign Ng33557 = ( (~ n706) ) ;
 assign n707 = ( n160  &  n2714  &  n2715 ) | ( n2714  &  n2715  &  n2713 ) ;
 assign Ng30511 = ( (~ n707) ) ;
 assign n708 = ( (~ n1248)  &  (~ n1253)  &  (~ n2521) ) | ( (~ n1248)  &  (~ n1253)  &  (~ Ng4567) ) ;
 assign Ng33045 = ( (~ n708) ) ;
 assign n709 = ( Pg35  &  n3068  &  (~ n5847) ) | ( n3068  &  (~ Ng2518)  &  (~ n5847) ) ;
 assign Ng30379 = ( (~ n709) ) ;
 assign n713 = ( (~ Pg16718)  &  (~ Pg13895) ) | ( (~ Pg16718)  &  Pg11349 ) | ( Pg13895  &  Pg11349 ) ;
 assign Ng24267 = ( Pg35  &  (~ Pg16624)  &  (~ Pg16603)  &  (~ Pg14421)  &  n713 ) ;
 assign n714 = ( n1747  &  n1745 ) | ( n1747  &  (~ Ng2643) ) ;
 assign Ng34020 = ( (~ n714) ) ;
 assign n717 = ( (~ n715)  &  Ng1489 ) | ( Ng1489  &  (~ Ng1495) ) ;
 assign n715 = ( Pg13272  &  (~ Ng1526)  &  (~ Ng1514) ) ;
 assign Ng24249 = ( Pg35  &  n717 ) | ( Pg35  &  n715  &  (~ Ng1442) ) ;
 assign n718 = ( (~ Ng2551)  &  n3062  &  (~ n5845) ) | ( n3062  &  n3060  &  (~ n5845) ) ;
 assign Ng30382 = ( (~ n718) ) ;
 assign n719 = ( n3402  &  n160 ) | ( n3402  &  Ng5156  &  n3401 ) ;
 assign Ng29285 = ( (~ n719) ) ;
 assign n720 = ( n1979  &  n1980  &  n1978 ) | ( n1979  &  n1980  &  (~ Ng6049) ) ;
 assign Ng33622 = ( (~ n720) ) ;
 assign n721 = ( n2096  &  n2097  &  (~ n4729) ) | ( n2096  &  n2097  &  (~ Ng2273) ) ;
 assign Ng33582 = ( (~ n721) ) ;
 assign n722 = ( (~ Pg35)  &  n3841 ) | ( n3837  &  n3841 ) | ( n3841  &  n3840 ) ;
 assign Ng28086 = ( (~ n722) ) ;
 assign n723 = ( n3584  &  n160 ) | ( n3584  &  Ng3147  &  n3583 ) ;
 assign Ng29262 = ( (~ n723) ) ;
 assign n724 = ( (~ Ng3338) ) | ( n5151 ) ;
 assign Ng24270 = ( (~ Pg35)  &  Ng3343 ) | ( Ng3343  &  n724 ) ;
 assign n725 = ( Pg35  &  n2099 ) | ( n2099  &  (~ Ng2265) ) ;
 assign Ng33581 = ( (~ n725) ) ;
 assign n726 = ( n1399  &  n1400  &  Ng626 ) | ( n1399  &  n1400  &  n1398 ) ;
 assign Ng34849 = ( (~ n726) ) ;
 assign n727 = ( (~ Pg35)  &  n1736  &  n3873 ) | ( n1736  &  n3873  &  n3872 ) ;
 assign Ng28060 = ( (~ n727) ) ;
 assign n728 = ( n1991  &  n1992  &  n1990 ) | ( n1991  &  n1992  &  (~ Ng5357) ) ;
 assign Ng33618 = ( (~ n728) ) ;
 assign n729 = ( Pg35  &  n1715  &  n1716 ) | ( n1715  &  n1716  &  (~ Ng4983) ) ;
 assign Ng34038 = ( (~ n729) ) ;
 assign n730 = ( Pg35  &  n1725 ) | ( n1725  &  (~ Ng4785) ) ;
 assign Ng34032 = ( (~ n730) ) ;
 assign n731 = ( n160  &  n2720  &  n2721 ) | ( n2720  &  n2721  &  n2719 ) ;
 assign Ng30509 = ( (~ n731) ) ;
 assign n732 = ( Pg35  &  n1456 ) | ( n1456  &  (~ Ng4922) ) ;
 assign Ng34640 = ( (~ n732) ) ;
 assign n733 = ( Pg35  &  n3528  &  n3869 ) | ( n3528  &  n3869  &  (~ Ng3965) ) ;
 assign Ng28069 = ( (~ n733) ) ;
 assign n734 = ( n2544  &  n2545  &  Ng918 ) | ( n2544  &  n2545  &  (~ n4826) ) ;
 assign Ng31868 = ( (~ n734) ) ;
 assign n735 = ( (~ Pg35)  &  n1994  &  n3955 ) | ( n1994  &  n3955  &  n3954 ) ;
 assign Ng26938 = ( (~ n735) ) ;
 assign n736 = ( Pg35  &  n3107  &  (~ n5863) ) | ( n3107  &  (~ Ng2016)  &  (~ n5863) ) ;
 assign Ng30363 = ( (~ n736) ) ;
 assign n737 = ( n3179  &  n3180  &  Ng577 ) | ( n3179  &  n3180  &  n3178 ) ;
 assign Ng30334 = ( (~ n737) ) ;
 assign n738 = ( (~ n1271)  &  n1928  &  n1929 ) | ( n1928  &  n1929  &  n1927 ) ;
 assign Ng33970 = ( (~ n738) ) ;
 assign n739 = ( Pg35  &  n3044 ) | ( n3044  &  (~ Ng2771) ) ;
 assign Ng30391 = ( (~ n739) ) ;
 assign n740 = ( Ng930  &  n2216  &  n2217 ) | ( (~ n670)  &  n2216  &  n2217 ) ;
 assign Ng33540 = ( (~ n740) ) ;
 assign n741 = ( n2898  &  n2899  &  n160 ) | ( n2898  &  n2899  &  n2897 ) ;
 assign Ng30445 = ( (~ n741) ) ;
 assign n742 = ( Pg35  &  (~ n3784) ) | ( (~ n3784)  &  (~ Ng812) ) | ( Pg35  &  (~ n5485) ) | ( (~ Ng812)  &  (~ n5485) ) ;
 assign Ng25617 = ( (~ n742) ) ;
 assign n743 = ( (~ Ng837)  &  (~ n4247) ) | ( n3812  &  (~ n4246)  &  (~ n4247) ) ;
 assign Ng24215 = ( (~ n743) ) ;
 assign n744 = ( n1947  &  Ng599  &  (~ n6244) ) | ( n1947  &  n1945  &  (~ n6244) ) ;
 assign Ng33964 = ( (~ n744) ) ;
 assign n745 = ( n4088  &  n4089  &  (~ n4908) ) | ( n4088  &  n4089  &  (~ Ng5475) ) ;
 assign Ng25719 = ( (~ n745) ) ;
 assign n746 = ( Pg35  &  n3790 ) | ( Pg35  &  n3791 ) | ( n3790  &  (~ Ng736) ) | ( n3791  &  (~ Ng736) ) ;
 assign Ng29228 = ( (~ n746) ) ;
 assign n747 = ( n160  &  n2705  &  n2706 ) | ( n2705  &  n2706  &  n2704 ) ;
 assign Ng30514 = ( (~ n747) ) ;
 assign n748 = ( Pg35  &  n1954 ) | ( n1954  &  (~ Ng6741) ) | ( Pg35  &  (~ n6115) ) | ( (~ Ng6741)  &  (~ n6115) ) ;
 assign Ng33627 = ( (~ n748) ) ;
 assign n749 = ( Pg35  &  n1502 ) | ( n1502  &  (~ Ng2868) ) ;
 assign Ng34615 = ( (~ n749) ) ;
 assign n750 = ( n4106  &  n4103  &  (~ n6022) ) | ( n4106  &  (~ Ng5080)  &  (~ n6022) ) ;
 assign Ng25696 = ( (~ n750) ) ;
 assign n751 = ( n160  &  n2763  &  n2764 ) | ( n2763  &  n2764  &  n2762 ) ;
 assign Ng30493 = ( (~ n751) ) ;
 assign n752 = ( n1771  &  n2058 ) | ( n1771  &  (~ Ng2465) ) | ( n2058  &  (~ Ng2495) ) | ( (~ Ng2465)  &  (~ Ng2495) ) ;
 assign Ng33594 = ( (~ n752) ) ;
 assign n753 = ( (~ n1263)  &  n1785  &  n1786 ) | ( n1785  &  n1786  &  n1784 ) ;
 assign Ng34009 = ( (~ n753) ) ;
 assign n754 = ( Pg35  &  n3101 ) | ( (~ Ng2098)  &  n3101 ) ;
 assign Ng30365 = ( (~ n754) ) ;
 assign n755 = ( (~ n1260)  &  n1753  &  n1754 ) | ( n1753  &  n1754  &  (~ n4703) ) ;
 assign Ng34018 = ( (~ n755) ) ;
 assign n756 = ( Pg35  &  n1709 ) | ( n1709  &  (~ Ng4975) ) ;
 assign Ng34040 = ( (~ n756) ) ;
 assign n757 = ( n1720  &  n1733  &  n1734 ) | ( n1733  &  n1734  &  (~ Ng4785) ) ;
 assign Ng34029 = ( (~ n757) ) ;
 assign n758 = ( n160  &  n2778  &  n2779 ) | ( n2778  &  n2779  &  n2777 ) ;
 assign Ng30488 = ( (~ n758) ) ;
 assign n759 = ( n1522  &  n1523  &  Ng781 ) | ( n1522  &  n1523  &  n1521 ) ;
 assign Ng34600 = ( (~ n759) ) ;
 assign n760 = ( n4182  &  n4183  &  n4180 ) | ( n4182  &  n4183  &  (~ Ng686) ) ;
 assign Ng25614 = ( (~ n760) ) ;
 assign n761 = ( n3878  &  n3879  &  Ng1252 ) | ( n3878  &  n3879  &  n3877 ) ;
 assign Ng28058 = ( (~ n761) ) ;
 assign n762 = ( Pg35  &  n3802 ) | ( Pg35  &  n3803 ) | ( n3802  &  (~ Ng667) ) | ( n3803  &  (~ Ng667) ) ;
 assign Ng29225 = ( (~ n762) ) ;
 assign n763 = ( n160  &  n2656  &  (~ n6288) ) | ( n2656  &  n2655  &  (~ n6288) ) ;
 assign Ng30532 = ( (~ n763) ) ;
 assign n764 = ( (~ Ng5523)  &  (~ Ng5527) ) | ( (~ Ng5527)  &  n2274 ) | ( (~ Ng5523)  &  n2276 ) | ( n2274  &  n2276 ) ;
 assign Ng33054 = ( (~ n764) ) ;
 assign n765 = ( n2469  &  n2470  &  Ng1270 ) | ( n2469  &  n2470  &  n2468 ) ;
 assign Ng32984 = ( (~ n765) ) ;
 assign n766 = ( n1713  &  n1710 ) | ( n1713  &  n1711 ) | ( n1713  &  (~ Ng4991) ) ;
 assign Ng34039 = ( (~ n766) ) ;
 assign n767 = ( Pg35  &  n2243 ) | ( (~ Ng6219)  &  n2243 ) | ( Pg35  &  n2246 ) | ( (~ Ng6219)  &  n2246 ) ;
 assign Ng33065 = ( (~ n767) ) ;
 assign n768 = ( n2904  &  n2905  &  n160 ) | ( n2904  &  n2905  &  n2903 ) ;
 assign Ng30443 = ( (~ n768) ) ;
 assign n769 = ( n3347  &  n160 ) | ( n3347  &  Ng5503  &  n3346 ) ;
 assign Ng29291 = ( (~ n769) ) ;
 assign n770 = ( n160  &  n2723  &  n2724 ) | ( n2723  &  n2724  &  n2722 ) ;
 assign Ng30508 = ( (~ n770) ) ;
 assign n771 = ( n2845  &  n2846  &  n160 ) | ( n2845  &  n2846  &  n2844 ) ;
 assign Ng30464 = ( (~ n771) ) ;
 assign n772 = ( (~ n1265)  &  n1861  &  n1862 ) | ( n1861  &  n1862  &  n1860 ) ;
 assign Ng33988 = ( (~ n772) ) ;
 assign Ng30522 = ( (~ n2250)  &  (~ Ng6203) ) ;
 assign n775 = ( Pg35  &  n3080  &  (~ n5852) ) | ( n3080  &  (~ Ng2384)  &  (~ n5852) ) ;
 assign Ng30374 = ( (~ n775) ) ;
 assign n776 = ( (~ n1263)  &  n1788  &  n1789 ) | ( n1788  &  n1789  &  n1787 ) ;
 assign Ng34008 = ( (~ n776) ) ;
 assign n777 = ( n1605  &  n1604 ) | ( n1605  &  n1603 ) | ( n1605  &  n1592 ) ;
 assign Ng34444 = ( (~ n777) ) ;
 assign n778 = ( n1422  &  n1425 ) ;
 assign Ng34731 = ( (~ n778) ) ;
 assign n779 = ( n2033  &  n2034  &  (~ n4699) ) | ( n2033  &  n2034  &  (~ Ng2675) ) ;
 assign Ng33606 = ( (~ n779) ) ;
 assign n780 = ( Pg35  &  n4208 ) | ( n4208  &  (~ Ng4358) ) ;
 assign Ng24334 = ( (~ n780) ) ;
 assign Ng34265 = ( (~ Ng4871)  &  (~ Ng4836)  &  (~ Ng4864)  &  (~ n1533) ) ;
 assign n785 = ( n160  &  n2796  &  n2797 ) | ( n2796  &  n2797  &  n2795 ) ;
 assign Ng30482 = ( (~ n785) ) ;
 assign n786 = ( Pg35  &  n1520 ) | ( n1520  &  (~ Ng2130) ) ;
 assign Ng34604 = ( (~ n786) ) ;
 assign n787 = ( (~ Ng2338)  &  n2072  &  (~ n6130) ) | ( n2068  &  n2072  &  (~ n6130) ) ;
 assign Ng33591 = ( (~ n787) ) ;
 assign n788 = ( n160  &  n2677  &  n2678 ) | ( n2677  &  n2678  &  n2676 ) ;
 assign Ng30525 = ( (~ n788) ) ;
 assign n789 = ( Pg35  &  n3967 ) | ( (~ Ng2779)  &  n3967 ) ;
 assign Ng26929 = ( (~ n789) ) ;
 assign n790 = ( n2889  &  n2890  &  n160 ) | ( n2889  &  n2890  &  n2888 ) ;
 assign Ng30448 = ( (~ n790) ) ;
 assign n791 = ( n160  &  n2708  &  n2709 ) | ( n2708  &  n2709  &  n2707 ) ;
 assign Ng30513 = ( (~ n791) ) ;
 assign n792 = ( n2830  &  n2831  &  n160 ) | ( n2830  &  n2831  &  n2829 ) ;
 assign Ng30469 = ( (~ n792) ) ;
 assign n793 = ( n1736  &  n2024  &  Ng2759 ) | ( n1736  &  n2024  &  n2023 ) ;
 assign Ng33608 = ( (~ n793) ) ;
 assign n794 = ( n1961  &  n1962  &  n1960 ) | ( n1961  &  n1962  &  (~ Ng6741) ) ;
 assign Ng33626 = ( (~ n794) ) ;
 assign n795 = ( n1437  &  n1438  &  Ng785 ) | ( n1437  &  n1438  &  n1436 ) ;
 assign Ng34725 = ( (~ n795) ) ;
 assign n796 = ( n3157  &  n3158  &  Ng1259 ) | ( n3157  &  n3158  &  n3156 ) ;
 assign Ng30342 = ( (~ n796) ) ;
 assign n797 = ( Pg35  &  n3534 ) | ( (~ Ng3480)  &  n3534 ) ;
 assign Ng29267 = ( (~ n797) ) ;
 assign n798 = ( n160  &  n2613  &  n2614 ) | ( n2613  &  n2614  &  n2612 ) ;
 assign Ng30548 = ( (~ n798) ) ;
 assign n799 = ( Pg35  &  n2272 ) | ( Pg35  &  n2279 ) | ( n2272  &  (~ Ng5511) ) | ( n2279  &  (~ Ng5511) ) ;
 assign Ng33052 = ( (~ n799) ) ;
 assign n800 = ( (~ n1263)  &  n1776  &  (~ n6214) ) | ( n1776  &  n1775  &  (~ n6214) ) ;
 assign Ng34012 = ( (~ n800) ) ;
 assign n801 = ( (~ n1260)  &  n1756  &  n1757 ) | ( n1756  &  n1757  &  n1755 ) ;
 assign Ng34017 = ( (~ n801) ) ;
 assign n802 = ( Pg35  &  n4017  &  n4018 ) | ( n4017  &  n4018  &  (~ Ng921) ) ;
 assign Ng26912 = ( (~ n802) ) ;
 assign n803 = ( Pg35  &  n3104  &  (~ n5862) ) | ( n3104  &  (~ Ng2093)  &  (~ n5862) ) ;
 assign Ng30364 = ( (~ n803) ) ;
 assign n804 = ( (~ Pg35)  &  (~ Ng4473) ) | ( n1679  &  (~ Ng4473) ) | ( (~ Pg35)  &  n1681 ) | ( n1679  &  n1681 ) ;
 assign Ng34254 = ( (~ n804) ) ;
 assign n805 = ( n1687  &  Ng604  &  (~ n6207) ) | ( n1687  &  n1685  &  (~ n6207) ) ;
 assign Ng34251 = ( (~ n805) ) ;
 assign n806 = ( n160  &  n2577  &  n2578 ) | ( n2577  &  n2578  &  n2576 ) ;
 assign Ng30560 = ( (~ n806) ) ;
 assign n807 = ( (~ n1267)  &  n1881  &  n1882 ) | ( n1881  &  n1882  &  (~ n4755) ) ;
 assign Ng33983 = ( (~ n807) ) ;
 assign n808 = ( (~ n1267)  &  n1890  &  n1891 ) | ( n1890  &  n1891  &  n1889 ) ;
 assign Ng33980 = ( (~ n808) ) ;
 assign n809 = ( Pg35  &  n1474 ) | ( n1474  &  (~ Ng4253) ) ;
 assign Ng34631 = ( (~ n809) ) ;
 assign n810 = ( (~ Pg35)  &  (~ n3741) ) | ( n3738  &  (~ n3741) ) | ( (~ n3741)  &  (~ Ng1825) ) ;
 assign Ng29243 = ( (~ n810) ) ;
 assign n811 = ( (~ Ng969)  &  (~ n4158) ) | ( Pg35  &  n379  &  (~ n4158) ) ;
 assign Ng25623 = ( (~ n811) ) ;
 assign n812 = ( Pg35  &  n3920 ) | ( n3920  &  (~ Ng4417) ) ;
 assign Ng26950 = ( (~ n812) ) ;
 assign n813 = ( n2935  &  n2936  &  n160 ) | ( n2935  &  n2936  &  n2934 ) ;
 assign Ng30431 = ( (~ n813) ) ;
 assign n814 = ( n2836  &  n2837  &  n160 ) | ( n2836  &  n2837  &  n2835 ) ;
 assign Ng30467 = ( (~ n814) ) ;
 assign n815 = ( Pg35  &  n3131  &  (~ n5873) ) | ( n3131  &  (~ Ng1748)  &  (~ n5873) ) ;
 assign Ng30353 = ( (~ n815) ) ;
 assign n816 = ( Pg35  &  n1532 ) | ( Pg35  &  n1533 ) | ( n1532  &  (~ Ng4849) ) | ( n1533  &  (~ Ng4849) ) ;
 assign Ng34467 = ( (~ n816) ) ;
 assign n817 = ( n2907  &  n2908  &  n160 ) | ( n2907  &  n2908  &  n2906 ) ;
 assign Ng30442 = ( (~ n817) ) ;
 assign n818 = ( n3192  &  (~ n4569)  &  (~ n5885) ) | ( n3192  &  (~ n4983)  &  (~ n5885) ) ;
 assign Ng29305 = ( (~ n818) ) ;
 assign Ng25616 = ( Pg35  &  (~ n5186) ) ;
 assign n820 = ( n3668  &  n3669  &  (~ Ng2433) ) | ( n3668  &  n3669  &  (~ n4950) ) ;
 assign Ng29252 = ( (~ n820) ) ;
 assign n821 = ( n2410  &  n2406  &  n2411 ) ;
 assign Ng33003 = ( (~ n821) ) ;
 assign Ng34613 = ( (~ n1505) ) ;
 assign n823 = ( n1847  &  n2121 ) | ( n1847  &  (~ Ng2040) ) | ( n2121  &  (~ Ng2070) ) | ( (~ Ng2040)  &  (~ Ng2070) ) ;
 assign Ng33570 = ( (~ n823) ) ;
 assign n827 = ( (~ Pg16775)  &  (~ Pg13966) ) | ( (~ Pg16775)  &  Pg11418 ) | ( Pg13966  &  Pg11418 ) ;
 assign Ng24275 = ( Pg35  &  (~ Pg16693)  &  (~ Pg16659)  &  (~ Pg14518)  &  n827 ) ;
 assign n828 = ( Pg35  &  n3241 ) | ( (~ Ng6177)  &  n3241 ) ;
 assign Ng29302 = ( (~ n828) ) ;
 assign n829 = ( n160  &  n2790  &  n2791 ) | ( n2790  &  n2791  &  n2789 ) ;
 assign Ng30484 = ( (~ n829) ) ;
 assign n830 = ( (~ Ng1395)  &  n3984 ) | ( Ng1395  &  (~ n3984) ) ;
 assign Ng25634 = ( Pg35  &  n830  &  (~ Ng1322) ) ;
 assign n832 = ( (~ Ng1913)  &  n2135  &  (~ n6133) ) | ( n2131  &  n2135  &  (~ n6133) ) ;
 assign Ng33567 = ( (~ n832) ) ;
 assign n833 = ( n1796  &  n2084  &  n2085 ) | ( n2084  &  n2085  &  (~ Ng2331) ) ;
 assign Ng33585 = ( (~ n833) ) ;
 assign n834 = ( n160  &  n2671  &  n2672 ) | ( n2671  &  n2672  &  n2670 ) ;
 assign Ng30527 = ( (~ n834) ) ;
 assign n835 = ( n160  &  n2892  &  (~ n6366) ) | ( n2892  &  n2891  &  (~ n6366) ) ;
 assign Ng30447 = ( (~ n835) ) ;
 assign n836 = ( (~ Ng1266)  &  n4149 ) | ( n4149  &  n4152 ) | ( (~ Ng1266)  &  (~ Ng1249) ) | ( n4152  &  (~ Ng1249) ) ;
 assign Ng25630 = ( (~ n836) ) ;
 assign n837 = ( Pg35  &  n3349 ) | ( (~ Ng5485)  &  n3349 ) ;
 assign Ng29290 = ( (~ n837) ) ;
 assign n838 = ( Pg35  &  n3797  &  n3798 ) | ( n3797  &  n3798  &  (~ Ng676) ) ;
 assign Ng29227 = ( (~ n838) ) ;
 assign n839 = ( Pg35  &  n2532  &  n2533 ) | ( n2532  &  n2533  &  (~ Ng2741) ) ;
 assign Ng31872 = ( (~ n839) ) ;
 assign n840 = ( n3355  &  (~ n4341)  &  (~ n5910) ) | ( n3355  &  (~ n5005)  &  (~ n5910) ) ;
 assign Ng29287 = ( (~ n840) ) ;
 assign n841 = ( Pg35  &  n2304  &  n2520 ) | ( n2304  &  n2520  &  (~ Ng4423) ) ;
 assign Ng31897 = ( (~ n841) ) ;
 assign n842 = ( n160  &  n2572  &  n2573 ) | ( n2572  &  n2573  &  n2571 ) ;
 assign Ng30562 = ( (~ n842) ) ;
 assign n843 = ( (~ n1263)  &  n1779  &  n1780 ) | ( n1779  &  n1780  &  (~ n4713) ) ;
 assign Ng34011 = ( (~ n843) ) ;
 assign n844 = ( (~ n1269)  &  n1832  &  n1833 ) | ( n1832  &  n1833  &  n1831 ) ;
 assign Ng33996 = ( (~ n844) ) ;
 assign n845 = ( (~ Ng2491)  &  n2376  &  n2377 ) | ( n2372  &  n2376  &  n2377 ) ;
 assign Ng33014 = ( (~ n845) ) ;
 assign n846 = ( Pg35  &  n1537  &  (~ n6200) ) | ( n1537  &  (~ Ng4843)  &  (~ n6200) ) ;
 assign Ng34465 = ( (~ n846) ) ;
 assign n847 = ( (~ n1269)  &  n1835  &  n1836 ) | ( n1835  &  n1836  &  n1834 ) ;
 assign Ng33995 = ( (~ n847) ) ;
 assign n848 = ( (~ Ng2283)  &  n3086  &  (~ n5855) ) | ( n3086  &  n3084  &  (~ n5855) ) ;
 assign Ng30372 = ( (~ n848) ) ;
 assign n849 = ( n160  &  n2622  &  n2623 ) | ( n2622  &  n2623  &  n2621 ) ;
 assign Ng30545 = ( (~ n849) ) ;
 assign n850 = ( Pg35  &  n3044 ) | ( (~ Ng2831)  &  n3044 ) ;
 assign Ng30389 = ( (~ n850) ) ;
 assign n851 = ( n2075  &  n2076  &  (~ n4719) ) | ( n2075  &  n2076  &  (~ Ng2407) ) ;
 assign Ng33590 = ( (~ n851) ) ;
 assign n852 = ( Pg35  &  n1501 ) | ( n1501  &  (~ Ng2988) ) ;
 assign Ng34616 = ( (~ n852) ) ;
 assign n853 = ( Pg35  &  n3971 ) | ( (~ Ng2763)  &  n3971 ) ;
 assign Ng26927 = ( (~ n853) ) ;
 assign n855 = ( n1217  &  n2194  &  (~ n6035) ) | ( n2194  &  Ng1351  &  (~ n6035) ) ;
 assign n854 = ( (~ n2194) ) | ( n4322 ) ;
 assign Ng25631 = ( Pg35  &  n855 ) | ( Pg35  &  Ng1312  &  n854 ) ;
 assign n856 = ( n160  &  n2806  &  n2807 ) | ( n2284  &  n2806  &  n2807 ) ;
 assign Ng30477 = ( (~ n856) ) ;
 assign n857 = ( Pg35  &  n1472 ) | ( n1472  &  (~ Ng4249) ) ;
 assign Ng34632 = ( (~ n857) ) ;
 assign n858 = ( n3891  &  (~ Ng645) ) | ( (~ Ng446)  &  (~ Ng645) ) | ( n3891  &  (~ n5074) ) | ( (~ Ng446)  &  (~ n5074) ) ;
 assign Ng28046 = ( (~ n858) ) ;
 assign n859 = ( Pg35  &  n4044  &  (~ n4380) ) | ( n4044  &  (~ Ng728)  &  (~ n4380) ) ;
 assign Ng26896 = ( (~ n859) ) ;
 assign n860 = ( Pg35  &  n4200 ) | ( n4200  &  (~ Ng405) ) ;
 assign Ng25602 = ( (~ n860) ) ;
 assign n861 = ( Ng1129  &  n3999  &  n4000 ) | ( n3999  &  n4000  &  (~ n5091) ) ;
 assign Ng26916 = ( (~ n861) ) ;
 assign n862 = ( n1821  &  n2100 ) | ( n1821  &  (~ Ng2197) ) | ( n2100  &  (~ Ng2227) ) | ( (~ Ng2197)  &  (~ Ng2227) ) ;
 assign Ng33578 = ( (~ n862) ) ;
 assign n863 = ( Pg35  &  n3128  &  (~ n5872) ) | ( n3128  &  (~ Ng1825)  &  (~ n5872) ) ;
 assign Ng30354 = ( (~ n863) ) ;
 assign n864 = ( n160  &  n2953  &  (~ n6386) ) | ( n2953  &  n2952  &  (~ n6386) ) ;
 assign Ng30425 = ( (~ n864) ) ;
 assign n865 = ( Pg35  &  n4265  &  n4266 ) | ( n4265  &  n4266  &  (~ Ng401) ) ;
 assign Ng24200 = ( (~ n865) ) ;
 assign n866 = ( n1923  &  n2191 ) | ( n2191  &  (~ Ng1592) ) ;
 assign Ng33544 = ( (~ n866) ) ;
 assign n867 = ( n4233  &  n4234  &  Ng1221 ) | ( n4233  &  n4234  &  (~ n5133) ) ;
 assign Ng24246 = ( (~ n867) ) ;
 assign n868 = ( n160  &  n2726  &  n2727 ) | ( n2726  &  n2727  &  n2725 ) ;
 assign Ng30507 = ( (~ n868) ) ;
 assign n869 = ( Pg35  &  n3181 ) | ( Pg35  &  n3182 ) | ( n3181  &  (~ Ng142) ) | ( n3182  &  (~ Ng142) ) ;
 assign Ng30333 = ( (~ n869) ) ;
 assign n870 = ( (~ Ng1932)  &  n2430  &  n2431 ) | ( n2426  &  n2430  &  n2431 ) ;
 assign Ng32998 = ( (~ n870) ) ;
 assign n871 = ( n2463  &  n2459  &  n2464 ) ;
 assign Ng32987 = ( (~ n871) ) ;
 assign n872 = ( Pg35  &  n3400  &  (~ n5913) ) | ( n3400  &  (~ Ng5467)  &  (~ n5913) ) ;
 assign Ng29286 = ( (~ n872) ) ;
 assign n873 = ( (~ Pg35) ) | ( (~ Ng2689) ) ;
 assign Ng34606 = ( (~ n873) ) ;
 assign n874 = ( Pg35  &  n2230 ) | ( (~ Ng6565)  &  n2230 ) | ( Pg35  &  n2233 ) | ( (~ Ng6565)  &  n2233 ) ;
 assign Ng33070 = ( (~ n874) ) ;
 assign n875 = ( n3770  &  n3771  &  (~ Ng1604) ) | ( n3770  &  n3771  &  (~ n4969) ) ;
 assign Ng29240 = ( (~ n875) ) ;
 assign n876 = ( Pg35  &  n2424  &  n2425 ) | ( n2424  &  n2425  &  (~ Ng2036) ) ;
 assign Ng32999 = ( (~ n876) ) ;
 assign n877 = ( Pg35  &  n2036 ) | ( n2036  &  (~ Ng2667) ) ;
 assign Ng33605 = ( (~ n877) ) ;
 assign n878 = ( (~ Pg17423)  &  n4227  &  n4228 ) | ( n4222  &  n4227  &  n4228 ) ;
 assign Ng24255 = ( (~ n878) ) ;
 assign n879 = ( Pg35  &  n3949  &  n3953 ) | ( n3949  &  n3953  &  (~ Ng4411) ) ;
 assign Ng26945 = ( (~ n879) ) ;
 assign n880 = ( n2159  &  n2160  &  (~ n4760) ) | ( n2159  &  n2160  &  (~ Ng1848) ) ;
 assign Ng33558 = ( (~ n880) ) ;
 assign n881 = ( wire4434  &  n4097  &  (~ n6444) ) | ( n4097  &  n4096  &  (~ n6444) ) ;
 assign Ng25699 = ( (~ n881) ) ;
 assign n882 = ( (~ Ng5485)  &  n3351  &  (~ n5908) ) | ( n3351  &  n3350  &  (~ n5908) ) ;
 assign Ng29289 = ( (~ n882) ) ;
 assign n883 = ( Pg35  &  n3045 ) | ( Pg35  &  n3046 ) | ( n3045  &  (~ Ng2735) ) | ( n3046  &  (~ Ng2735) ) ;
 assign Ng30388 = ( (~ n883) ) ;
 assign n884 = ( n3651  &  n3652  &  (~ Ng2567) ) | ( n3651  &  n3652  &  (~ n4946) ) ;
 assign Ng29254 = ( (~ n884) ) ;
 assign n885 = ( n3861  &  n3862  &  n3855 ) | ( n3861  &  n3862  &  n3860 ) ;
 assign Ng28074 = ( (~ n885) ) ;
 assign n886 = ( Pg35  &  n1587  &  n1588 ) | ( n1587  &  n1588  &  (~ Ng4311) ) ;
 assign Ng34450 = ( (~ n886) ) ;
 assign n887 = ( n160  &  n2711  &  (~ n6306) ) | ( n2711  &  n2710  &  (~ n6306) ) ;
 assign Ng30512 = ( (~ n887) ) ;
 assign n888 = ( (~ Ng1644)  &  n2177  &  (~ n6135) ) | ( n2173  &  n2177  &  (~ n6135) ) ;
 assign Ng33551 = ( (~ n888) ) ;
 assign n889 = ( n2223  &  Ng595  &  (~ n6251) ) | ( n2223  &  n2221  &  (~ n6251) ) ;
 assign Ng33538 = ( (~ n889) ) ;
 assign n890 = ( n2401  &  n2406  &  n2407 ) | ( n2406  &  n2407  &  (~ Ng2217) ) ;
 assign Ng33005 = ( (~ n890) ) ;
 assign n891 = ( (~ Ng1404)  &  n4231 ) | ( Ng1404  &  (~ n4231) ) ;
 assign Ng24248 = ( n891 ) | ( (~ n5634) ) ;
 assign n893 = ( (~ Ng2066)  &  n2416  &  n2417 ) | ( n2412  &  n2416  &  n2417 ) ;
 assign Ng33002 = ( (~ n893) ) ;
 assign n894 = ( n160  &  n2824  &  (~ n6343) ) | ( n2824  &  n2823  &  (~ n6343) ) ;
 assign Ng30471 = ( (~ n894) ) ;
 assign n895 = ( Pg35  &  n1818 ) | ( n1818  &  (~ Ng2246) ) ;
 assign Ng34000 = ( (~ n895) ) ;
 assign n896 = ( (~ n1260)  &  n1759  &  n1760 ) | ( n1759  &  n1760  &  n1758 ) ;
 assign Ng34016 = ( (~ n896) ) ;
 assign n897 = ( Pg35  &  n2289 ) | ( Pg35  &  n2290 ) | ( n2289  &  (~ Ng5170) ) | ( n2290  &  (~ Ng5170) ) ;
 assign Ng33048 = ( (~ n897) ) ;
 assign n898 = ( Pg35  &  n3957 ) | ( (~ Ng2823)  &  n3957 ) ;
 assign Ng26934 = ( (~ n898) ) ;
 assign n899 = ( n1531  &  n1530 ) | ( n1531  &  (~ Ng4854) ) | ( n1531  &  (~ n4630) ) ;
 assign Ng34468 = ( (~ n899) ) ;
 assign n900 = ( Ng1274  &  n2203  &  n2204 ) | ( (~ n666)  &  n2203  &  n2204 ) ;
 assign Ng33542 = ( (~ n900) ) ;
 assign n901 = ( n1602  &  n1591 ) | ( n1602  &  n1600 ) | ( n1602  &  n1601 ) ;
 assign Ng34445 = ( (~ n901) ) ;
 assign n902 = ( n1773  &  n1771 ) | ( n1773  &  (~ Ng2509) ) ;
 assign Ng34013 = ( (~ n902) ) ;
 assign n903 = ( Pg35  &  n3993  &  n3994 ) | ( n3993  &  n3994  &  (~ Ng1266) ) ;
 assign Ng26919 = ( (~ n903) ) ;
 assign n904 = ( n160  &  n2595  &  (~ n6268) ) | ( n2595  &  n2594  &  (~ n6268) ) ;
 assign Ng30554 = ( (~ n904) ) ;
 assign n905 = ( (~ n2560)  &  n3410  &  (~ n5918) ) | ( n3410  &  (~ n5012)  &  (~ n5918) ) ;
 assign Ng29281 = ( (~ n905) ) ;
 assign n906 = ( n160  &  n2641  &  n2642 ) | ( n2641  &  n2642  &  n2640 ) ;
 assign Ng30537 = ( (~ n906) ) ;
 assign n907 = ( Pg35  &  n1421 ) | ( n1421  &  (~ Ng2999) ) ;
 assign Ng34732 = ( (~ n907) ) ;
 assign n908 = ( Pg35  &  n3893 ) | ( n3893  &  (~ Ng699) ) ;
 assign Ng28049 = ( (~ n908) ) ;
 assign n909 = ( n1923  &  n2186  &  n2187 ) | ( n2186  &  n2187  &  (~ Ng1636) ) ;
 assign Ng33545 = ( (~ n909) ) ;
 assign n910 = ( n2910  &  n2911  &  n160 ) | ( n2910  &  n2911  &  n2909 ) ;
 assign Ng30441 = ( (~ n910) ) ;
 assign n911 = ( (~ Pg35)  &  (~ n3707) ) | ( n3704  &  (~ n3707) ) | ( (~ n3707)  &  (~ Ng2093) ) ;
 assign Ng29247 = ( (~ n911) ) ;
 assign n912 = ( Pg35  &  n4005 ) | ( n4005  &  (~ Ng1052) ) | ( Pg35  &  (~ n5630) ) | ( (~ Ng1052)  &  (~ n5630) ) ;
 assign Ng26914 = ( (~ n912) ) ;
 assign n913 = ( (~ n1269)  &  n1826  &  n1827 ) | ( n1826  &  n1827  &  n1825 ) ;
 assign Ng33998 = ( (~ n913) ) ;
 assign n914 = ( Ng956  &  n4154  &  n4155 ) | ( n4154  &  n4155  &  (~ n5135) ) ;
 assign Ng25626 = ( (~ n914) ) ;
 assign n915 = ( (~ n1257)  &  n1903  &  (~ n6234) ) | ( n1903  &  n1902  &  (~ n6234) ) ;
 assign Ng33977 = ( (~ n915) ) ;
 assign n916 = ( n3292  &  n160 ) | ( n3292  &  Ng5849  &  n3291 ) ;
 assign Ng29297 = ( (~ n916) ) ;
 assign n917 = ( (~ Ng2685)  &  n3050  &  (~ n5840) ) | ( n3050  &  n3048  &  (~ n5840) ) ;
 assign Ng30387 = ( (~ n917) ) ;
 assign n918 = ( n1821  &  n2105  &  n2106 ) | ( n2105  &  n2106  &  (~ Ng2197) ) ;
 assign Ng33577 = ( (~ n918) ) ;
 assign n919 = ( n1771  &  n2067 ) | ( n2067  &  (~ Ng2421) ) ;
 assign Ng33592 = ( (~ n919) ) ;
 assign n920 = ( Pg35  &  n4014  &  (~ n6188) ) | ( (~ Ng1041)  &  n4014  &  (~ n6188) ) ;
 assign Ng26913 = ( (~ n920) ) ;
 assign n921 = ( (~ Pg35)  &  n3809  &  n3903 ) | ( n3809  &  n3903  &  n3902 ) ;
 assign Ng28044 = ( (~ n921) ) ;
 assign n922 = ( n3929  &  (~ Ng4405) ) | ( (~ Ng4388)  &  (~ Ng4405) ) | ( n3943  &  (~ Ng4405) ) ;
 assign Ng26948 = ( (~ n922) ) ;
 assign n923 = ( n1209  &  (~ Ng1536) ) | ( Ng1526  &  n1209  &  (~ Ng1514) ) ;
 assign n924 = ( (~ Pg7946)  &  Ng1514 ) | ( Pg7946  &  (~ Ng1514) ) ;
 assign Ng30344 = ( Pg35  &  n923 ) | ( Pg35  &  n924 ) ;
 assign n925 = ( (~ Ng6561)  &  (~ Ng6565) ) | ( (~ Ng6565)  &  n2235 ) | ( (~ Ng6561)  &  n2237 ) | ( n2235  &  n2237 ) ;
 assign Ng33069 = ( (~ n925) ) ;
 assign n926 = ( Pg35  &  n1491 ) | ( n1491  &  (~ Ng2936) ) ;
 assign Ng34621 = ( (~ n926) ) ;
 assign n927 = ( (~ n2194)  &  n3876 ) | ( Ng1345  &  n3876 ) | ( n3876  &  n3875 ) ;
 assign Ng28059 = ( (~ n927) ) ;
 assign n928 = ( (~ Pg35) ) | ( (~ Ng4727) ) ;
 assign Ng34633 = ( (~ n928) ) ;
 assign n932 = ( (~ Pg17778)  &  (~ Pg14828) ) | ( (~ Pg17778)  &  Pg12470 ) | ( Pg14828  &  Pg12470 ) ;
 assign Ng24352 = ( Pg35  &  (~ Pg17722)  &  (~ Pg17688)  &  (~ Pg13099)  &  n932 ) ;
 assign n933 = ( n160  &  n2895  &  (~ n6367) ) | ( n2895  &  n2894  &  (~ n6367) ) ;
 assign Ng30446 = ( (~ n933) ) ;
 assign n934 = ( (~ Ng1858)  &  n3122  &  (~ n5870) ) | ( n3122  &  n3120  &  (~ n5870) ) ;
 assign Ng30357 = ( (~ n934) ) ;
 assign n935 = ( Pg35  &  n4021 ) | ( n4021  &  (~ Ng246) ) ;
 assign Ng26908 = ( (~ n935) ) ;
 assign n936 = ( n3026  &  n3027  &  n160 ) | ( n3026  &  n3027  &  n3025 ) ;
 assign Ng30399 = ( (~ n936) ) ;
 assign n937 = ( n3753  &  n3754  &  (~ Ng1740) ) | ( n3753  &  n3754  &  (~ n4966) ) ;
 assign Ng29242 = ( (~ n937) ) ;
 assign n938 = ( n160  &  n2616  &  n2617 ) | ( n2616  &  n2617  &  n2615 ) ;
 assign Ng30547 = ( (~ n938) ) ;
 assign n939 = ( (~ n1263)  &  n1782  &  n1783 ) | ( n1782  &  n1783  &  n1781 ) ;
 assign Ng34010 = ( (~ n939) ) ;
 assign n940 = ( Pg35  &  n1869 ) | ( n1869  &  (~ Ng1955) ) ;
 assign Ng33986 = ( (~ n940) ) ;
 assign n941 = ( n160  &  n2625  &  n2626 ) | ( n2625  &  n2626  &  n2624 ) ;
 assign Ng30544 = ( (~ n941) ) ;
 assign n942 = ( n160  &  n2574  &  (~ n6261) ) | ( n2232  &  n2574  &  (~ n6261) ) ;
 assign Ng30561 = ( (~ n942) ) ;
 assign n943 = ( n2938  &  n2939  &  n160 ) | ( n2938  &  n2939  &  n2937 ) ;
 assign Ng30430 = ( (~ n943) ) ;
 assign n944 = ( Pg35  &  n2141 ) | ( n2141  &  (~ Ng1974) ) ;
 assign Ng33565 = ( (~ n944) ) ;
 assign n945 = ( (~ n1271)  &  n1934  &  n1935 ) | ( n1934  &  n1935  &  n1933 ) ;
 assign Ng33968 = ( (~ n945) ) ;
 assign n946 = ( n2138  &  n2139  &  (~ n4750) ) | ( n2138  &  n2139  &  (~ Ng1982) ) ;
 assign Ng33566 = ( (~ n946) ) ;
 assign n947 = ( n2842  &  n2843  &  n160 ) | ( n2842  &  n2843  &  n2841 ) ;
 assign Ng30465 = ( (~ n947) ) ;
 assign n948 = ( n3860  &  n3863  &  n3864 ) | ( n3863  &  n3864  &  (~ n5070) ) ;
 assign Ng28073 = ( (~ n948) ) ;
 assign n949 = ( (~ Ng6381) ) | ( n5142 ) ;
 assign Ng24351 = ( (~ Pg35)  &  Ng6386 ) | ( Ng6386  &  n949 ) ;
 assign n950 = ( Pg35  &  n2498  &  (~ n5809) ) | ( n2498  &  (~ Ng5029)  &  (~ n5809) ) ;
 assign Ng31904 = ( (~ n950) ) ;
 assign n951 = ( Pg35  &  n1466 ) | ( n1466  &  (~ Ng4732) ) ;
 assign Ng34635 = ( (~ n951) ) ;
 assign n952 = ( n3477  &  n160 ) | ( n3477  &  Ng3849  &  n3476 ) ;
 assign Ng29274 = ( (~ n952) ) ;
 assign n953 = ( n3035  &  n3036  &  n160 ) | ( n3035  &  n3036  &  n3034 ) ;
 assign Ng30396 = ( (~ n953) ) ;
 assign n954 = ( Pg35  &  n4079 ) | ( n4079  &  (~ Ng5841) ) ;
 assign Ng25735 = ( (~ n954) ) ;
 assign n955 = ( n1704  &  n1717  &  n1718 ) | ( n1717  &  n1718  &  (~ Ng4975) ) ;
 assign Ng34037 = ( (~ n955) ) ;
 assign n956 = ( n1413  &  n1414  &  Ng790 ) | ( n1413  &  n1414  &  n1412 ) ;
 assign Ng34791 = ( (~ n956) ) ;
 assign n957 = ( n160  &  n2688  &  n2689 ) | ( n2688  &  n2689  &  n2687 ) ;
 assign Ng30520 = ( (~ n957) ) ;
 assign n958 = ( Pg35  &  n3119  &  (~ n5868) ) | ( n3119  &  (~ Ng1882)  &  (~ n5868) ) ;
 assign Ng30358 = ( (~ n958) ) ;
 assign n959 = ( (~ n2561)  &  n3247  &  (~ n5893) ) | ( n3247  &  (~ n4990)  &  (~ n5893) ) ;
 assign Ng29299 = ( (~ n959) ) ;
 assign n960 = ( Pg35  &  n3818 ) | ( n3818  &  (~ Ng5619) ) ;
 assign Ng28096 = ( (~ n960) ) ;
 assign n961 = ( n3830  &  n3832 ) | ( n3830  &  (~ Ng4939) ) | ( n3832  &  (~ n5621) ) | ( (~ Ng4939)  &  (~ n5621) ) ;
 assign Ng28088 = ( (~ n961) ) ;
 assign n962 = ( n3032  &  n3033  &  n160 ) | ( n3032  &  n3033  &  n3031 ) ;
 assign Ng30397 = ( (~ n962) ) ;
 assign n963 = ( n2996  &  n2997  &  n160 ) | ( n2996  &  n2997  &  n2995 ) ;
 assign Ng30409 = ( (~ n963) ) ;
 assign n964 = ( Pg35  &  n3404 ) | ( (~ Ng5138)  &  n3404 ) ;
 assign Ng29284 = ( (~ n964) ) ;
 assign n965 = ( n160  &  n2827  &  (~ n6344) ) | ( n2827  &  n2826  &  (~ n6344) ) ;
 assign Ng30470 = ( (~ n965) ) ;
 assign n966 = ( (~ Ng2126)  &  n3098  &  (~ n5860) ) | ( n3098  &  n3096  &  (~ n5860) ) ;
 assign Ng30367 = ( (~ n966) ) ;
 assign n967 = ( Pg35  &  n3116  &  (~ n5867) ) | ( n3116  &  (~ Ng1959)  &  (~ n5867) ) ;
 assign Ng30359 = ( (~ n967) ) ;
 assign n968 = ( n4100  &  n4101  &  Ng5097 ) | ( n4100  &  n4101  &  (~ n5122) ) ;
 assign Ng25698 = ( (~ n968) ) ;
 assign n969 = ( n3029  &  n3030  &  n160 ) | ( n3029  &  n3030  &  n3028 ) ;
 assign Ng30398 = ( (~ n969) ) ;
 assign n970 = ( (~ n3936)  &  (~ Ng4430) ) | ( Pg35  &  Ng4388  &  (~ n3936) ) ;
 assign Ng26952 = ( (~ n970) ) ;
 assign n971 = ( Pg35  &  n3969 ) | ( (~ Ng2767)  &  n3969 ) ;
 assign Ng26928 = ( (~ n971) ) ;
 assign n972 = ( n3934  &  n3935  &  n3926 ) | ( n3934  &  n3935  &  n3929 ) ;
 assign Ng26954 = ( (~ n972) ) ;
 assign n973 = ( Pg35  &  n2535  &  n2536 ) | ( (~ Ng1361)  &  n2535  &  n2536 ) ;
 assign Ng31871 = ( (~ n973) ) ;
 assign n974 = ( (~ n1269)  &  n1838  &  n1839 ) | ( n1838  &  n1839  &  n1837 ) ;
 assign Ng33994 = ( (~ n974) ) ;
 assign n975 = ( n1796  &  n2079 ) | ( n1796  &  (~ Ng2331) ) | ( n2079  &  (~ Ng2361) ) | ( (~ Ng2331)  &  (~ Ng2361) ) ;
 assign Ng33586 = ( (~ n975) ) ;
 assign n976 = ( n2550  &  n2551  &  Ng582 ) | ( n2550  &  n2551  &  n2549 ) ;
 assign Ng31866 = ( (~ n976) ) ;
 assign n977 = ( Pg35  &  n3083  &  (~ n5853) ) | ( n3083  &  (~ Ng2307)  &  (~ n5853) ) ;
 assign Ng30373 = ( (~ n977) ) ;
 assign n978 = ( n3884  &  n3885  &  Ng907 ) | ( n3884  &  n3885  &  n3883 ) ;
 assign Ng28056 = ( (~ n978) ) ;
 assign n979 = ( Pg35  &  n3125 ) | ( (~ Ng1830)  &  n3125 ) ;
 assign Ng30355 = ( (~ n979) ) ;
 assign n980 = ( n2950  &  n2951  &  n160 ) | ( n2950  &  n2951  &  n2949 ) ;
 assign Ng30426 = ( (~ n980) ) ;
 assign n983 = ( Ng2932 ) | ( Ng2999 ) ;
 assign n981 = ( n1355  &  n1356  &  n1357  &  n1358 ) ;
 assign Ng34805 = ( n983  &  Pg35 ) ;
 assign n984 = ( (~ n1273)  &  n1810  &  n1811 ) | ( n1810  &  n1811  &  n1809 ) ;
 assign Ng34002 = ( (~ n984) ) ;
 assign n985 = ( Pg35  &  n3890  &  n3891 ) | ( n3890  &  n3891  &  (~ Ng681) ) ;
 assign Ng28053 = ( (~ n985) ) ;
 assign n986 = ( Pg35  &  n3788  &  n3789 ) | ( n3788  &  n3789  &  (~ Ng827) ) ;
 assign Ng29229 = ( (~ n986) ) ;
 assign n987 = ( Pg35  &  n1982  &  n1983 ) | ( n1982  &  n1983  &  (~ Ng5698) ) ;
 assign Ng33620 = ( (~ n987) ) ;
 assign n988 = ( (~ Ng2472)  &  n2051  &  (~ n6129) ) | ( n2047  &  n2051  &  (~ n6129) ) ;
 assign Ng33599 = ( (~ n988) ) ;
 assign n989 = ( n160  &  n2702  &  n2703 ) | ( n2702  &  n2703  &  n2701 ) ;
 assign Ng30515 = ( (~ n989) ) ;
 assign n990 = ( Pg35  &  n1895 ) | ( n1895  &  (~ Ng1821) ) ;
 assign Ng33979 = ( (~ n990) ) ;
 assign n991 = ( n2977  &  n2978  &  n160 ) | ( n2977  &  n2978  &  n2976 ) ;
 assign Ng30417 = ( (~ n991) ) ;
 assign n992 = ( Pg35  &  n4117 ) | ( n4117  &  (~ Ng3841) ) ;
 assign Ng25683 = ( (~ n992) ) ;
 assign n993 = ( n2117  &  n2118  &  (~ n4740) ) | ( n2117  &  n2118  &  (~ Ng2116) ) ;
 assign Ng33574 = ( (~ n993) ) ;
 assign n994 = ( n2993  &  n2994  &  n160 ) | ( n2993  &  n2994  &  n2992 ) ;
 assign Ng30410 = ( (~ n994) ) ;
 assign n995 = ( n2872  &  n2873  &  n160 ) | ( n2872  &  n2873  &  n2871 ) ;
 assign Ng30454 = ( (~ n995) ) ;
 assign n996 = ( Pg35  &  n1516 ) | ( n1516  &  (~ Ng2689) ) ;
 assign Ng34607 = ( (~ n996) ) ;
 assign n997 = ( Pg35  &  (~ n4794) ) | ( (~ n4794)  &  (~ Ng4382) ) ;
 assign Ng31895 = ( (~ n997) ) ;
 assign n998 = ( Pg35  &  n2237 ) | ( Pg35  &  n2238 ) | ( n2237  &  (~ Ng6555) ) | ( n2238  &  (~ Ng6555) ) ;
 assign Ng33068 = ( (~ n998) ) ;
 assign n999 = ( n3780  &  n3778 ) | ( n3780  &  (~ Ng1141) ) ;
 assign Ng29233 = ( (~ n999) ) ;
 assign n1000 = ( Pg35  &  n2183 ) | ( n2183  &  (~ Ng1706) ) ;
 assign Ng33549 = ( (~ n1000) ) ;
 assign n1001 = ( Pg35  &  n3187 ) | ( (~ Ng6523)  &  n3187 ) ;
 assign Ng29308 = ( (~ n1001) ) ;
 assign n1002 = ( n2999  &  n3000  &  n160 ) | ( n2999  &  n3000  &  n2998 ) ;
 assign Ng30408 = ( (~ n1002) ) ;
 assign n1003 = ( (~ Pg35)  &  (~ n3758) ) | ( n3755  &  (~ n3758) ) | ( (~ n3758)  &  (~ Ng1691) ) ;
 assign Ng29241 = ( (~ n1003) ) ;
 assign n1004 = ( Pg35  &  n1493 ) | ( n1493  &  (~ Ng2922) ) ;
 assign Ng34620 = ( (~ n1004) ) ;
 assign n1005 = ( Pg35  &  n4091 ) | ( n4091  &  (~ Ng5148) ) ;
 assign Ng25707 = ( (~ n1005) ) ;
 assign n1006 = ( (~ wire4415) ) | ( n5147 ) ;
 assign Ng24339 = ( (~ Pg35)  &  Ng5348 ) | ( Ng5348  &  n1006 ) ;
 assign n1007 = ( n1607  &  n1604 ) | ( n1607  &  n1606 ) | ( n1607  &  n1595 ) ;
 assign Ng34443 = ( (~ n1007) ) ;
 assign n1008 = ( Pg35  &  n1495 ) | ( n1495  &  (~ Ng2912) ) ;
 assign Ng34619 = ( (~ n1008) ) ;
 assign n1009 = ( n160  &  n2738  &  n2739 ) | ( n2738  &  n2739  &  n2737 ) ;
 assign Ng30503 = ( (~ n1009) ) ;
 assign n1010 = ( n160  &  n2607  &  n2608 ) | ( n2607  &  n2608  &  n2606 ) ;
 assign Ng30550 = ( (~ n1010) ) ;
 assign n1011 = ( n2414  &  n2419  &  n2420 ) | ( n2419  &  n2420  &  (~ Ng2060) ) ;
 assign Ng33001 = ( (~ n1011) ) ;
 assign n1012 = ( n160  &  n2766  &  n2767 ) | ( n2766  &  n2767  &  n2765 ) ;
 assign Ng30492 = ( (~ n1012) ) ;
 assign n1013 = ( Pg135 ) | ( n1373 ) ;
 assign n1014 = ( (~ Ng4349) ) | ( (~ Ng4358) ) ;
 assign n1015 = ( (~ Ng4633) ) | ( n4637 ) ;
 assign Ng26944 = ( Pg35  &  n1013 ) | ( Pg35  &  n1014 ) | ( Pg35  &  n1015 ) ;
 assign n1016 = ( n3587  &  n3586  &  (~ n5944) ) | ( n3587  &  (~ Ng3129)  &  (~ n5944) ) ;
 assign Ng29260 = ( (~ n1016) ) ;
 assign n1017 = ( Pg35  &  n2285 ) | ( Pg35  &  n2292 ) | ( n2285  &  (~ Ng5164) ) | ( n2292  &  (~ Ng5164) ) ;
 assign Ng33047 = ( (~ n1017) ) ;
 assign n1018 = ( n4082  &  n4083  &  (~ n4901) ) | ( n4082  &  n4083  &  (~ Ng5821) ) ;
 assign Ng25733 = ( (~ n1018) ) ;
 assign n1019 = ( n160  &  n2644  &  n2645 ) | ( n2644  &  n2645  &  n2643 ) ;
 assign Ng30536 = ( (~ n1019) ) ;
 assign n1020 = ( n3719  &  n3720  &  (~ Ng2008) ) | ( n3719  &  n3720  &  (~ n4960) ) ;
 assign Ng29246 = ( (~ n1020) ) ;
 assign n1021 = ( n2012  &  n2013  &  n2011 ) | ( n2012  &  n2013  &  (~ Ng3703) ) ;
 assign Ng33611 = ( (~ n1021) ) ;
 assign n1022 = ( n1429  &  n1432 ) ;
 assign Ng34728 = ( (~ n1022) ) ;
 assign n1023 = ( n3813  &  n3812  &  (~ n5983) ) | ( n3813  &  (~ Ng411)  &  (~ n5983) ) ;
 assign Ng29222 = ( (~ n1023) ) ;
 assign n1024 = ( n160  &  n2886  &  (~ n6364) ) | ( n2886  &  n2885  &  (~ n6364) ) ;
 assign Ng30449 = ( (~ n1024) ) ;
 assign n1025 = ( Pg35  &  n1514 ) | ( n1514  &  (~ Ng2697) ) ;
 assign Ng34608 = ( (~ n1025) ) ;
 assign n1026 = ( Ng1300  &  n4138  &  n4139 ) | ( n4138  &  n4139  &  (~ n5132) ) ;
 assign Ng25635 = ( (~ n1026) ) ;
 assign n1027 = ( n2854  &  n2855  &  n160 ) | ( n2854  &  n2855  &  n2853 ) ;
 assign Ng30461 = ( (~ n1027) ) ;
 assign n1028 = ( n2511  &  n2509 ) | ( n2511  &  (~ Ng5046) ) | ( n2511  &  (~ n5327) ) ;
 assign Ng31901 = ( (~ n1028) ) ;
 assign n1029 = ( (~ Pg35)  &  (~ n3690) ) | ( n3687  &  (~ n3690) ) | ( (~ n3690)  &  (~ Ng2250) ) ;
 assign Ng29249 = ( (~ n1029) ) ;
 assign n1030 = ( (~ n1248)  &  n2304  &  (~ n2521) ) | ( (~ n1248)  &  n2304  &  (~ Ng4546) ) ;
 assign Ng33041 = ( (~ n1030) ) ;
 assign n1031 = ( Pg35  &  n2384  &  n2385 ) | ( n2384  &  n2385  &  (~ Ng2461) ) ;
 assign Ng33011 = ( (~ n1031) ) ;
 assign n1032 = ( Pg35  &  n1497 ) | ( n1497  &  (~ Ng2907) ) ;
 assign Ng34618 = ( (~ n1032) ) ;
 assign n1033 = ( (~ Ng2357)  &  n2390  &  n2391 ) | ( n2386  &  n2390  &  n2391 ) ;
 assign Ng33010 = ( (~ n1033) ) ;
 assign n1034 = ( Pg35  &  n2553  &  n2554 ) | ( n2553  &  n2554  &  (~ Ng146) ) ;
 assign Ng31864 = ( (~ n1034) ) ;
 assign n1035 = ( Pg35  &  n1476 ) | ( n1476  &  (~ Ng4300) ) ;
 assign Ng34630 = ( (~ n1035) ) ;
 assign n1036 = ( n2509  &  n2519 ) | ( n2519  &  Ng5016 ) | ( n2519  &  (~ n4884) ) ;
 assign Ng31898 = ( (~ n1036) ) ;
 assign n1037 = ( n4132  &  n4133  &  (~ n4934) ) | ( n4132  &  n4133  &  (~ Ng3119) ) ;
 assign Ng25653 = ( (~ n1037) ) ;
 assign n1038 = ( (~ Ng1312)  &  (~ n4142) ) | ( Pg35  &  n854  &  (~ n4142) ) ;
 assign Ng25632 = ( (~ n1038) ) ;
 assign n1039 = ( n3453  &  Ng5115  &  (~ n5921) ) | ( n3453  &  n3452  &  (~ n5921) ) ;
 assign Ng29280 = ( (~ n1039) ) ;
 assign n1040 = ( Pg35  &  n2021  &  n2022 ) | ( n2021  &  n2022  &  (~ Ng3347) ) ;
 assign Ng33609 = ( (~ n1040) ) ;
 assign n1041 = ( Pg35  &  n2569 ) | ( n2569  &  (~ Ng6653) ) ;
 assign Ng30563 = ( (~ n1041) ) ;
 assign n1042 = ( n2922  &  n2923  &  n160 ) | ( n2922  &  n2923  &  n2921 ) ;
 assign Ng30437 = ( (~ n1042) ) ;
 assign n1043 = ( n2988  &  n2989  &  n160 ) | ( n2988  &  n2989  &  n2987 ) ;
 assign Ng30412 = ( (~ n1043) ) ;
 assign n1044 = ( n160  &  n2769  &  (~ n6325) ) | ( n2769  &  n2768  &  (~ n6325) ) ;
 assign Ng30491 = ( (~ n1044) ) ;
 assign n1045 = ( Pg35  &  n2928 ) | ( n2928  &  (~ Ng3610) ) ;
 assign Ng30434 = ( (~ n1045) ) ;
 assign n1046 = ( Pg35  &  n1507 ) | ( n1507  &  (~ Ng2860) ) ;
 assign Ng34612 = ( (~ n1046) ) ;
 assign n1047 = ( n4120  &  n4121  &  (~ n4922) ) | ( n4120  &  n4121  &  (~ Ng3821) ) ;
 assign Ng25681 = ( (~ n1047) ) ;
 assign n1048 = ( Pg35  &  n4112  &  n4113 ) | ( (~ Ng4057)  &  n4112  &  n4113 ) ;
 assign Ng25687 = ( (~ n1048) ) ;
 assign n1049 = ( Pg35  &  n2802 ) | ( n2802  &  (~ Ng5268) ) ;
 assign Ng30479 = ( (~ n1049) ) ;
 assign n1050 = ( n1736  &  n3635  &  Ng2735 ) | ( n1736  &  n3635  &  n3634 ) ;
 assign Ng29256 = ( (~ n1050) ) ;
 assign n1051 = ( n160  &  n2647  &  n2648 ) | ( n2647  &  n2648  &  n2646 ) ;
 assign Ng30535 = ( (~ n1051) ) ;
 assign n1052 = ( Pg35  &  n3053 ) | ( (~ Ng2657)  &  n3053 ) ;
 assign Ng30385 = ( (~ n1052) ) ;
 assign n1053 = ( n4094  &  n4095  &  n4092 ) | ( n4094  &  n4095  &  (~ Ng5128) ) ;
 assign Ng25705 = ( (~ n1053) ) ;
 assign n1054 = ( Pg35  &  n3633  &  (~ n5949) ) | ( n3633  &  (~ Ng3111)  &  (~ n5949) ) ;
 assign Ng29257 = ( (~ n1054) ) ;
 assign n1055 = ( Pg35  &  n1547  &  (~ n6201) ) | ( n1547  &  (~ Ng4653)  &  (~ n6201) ) ;
 assign Ng34461 = ( (~ n1055) ) ;
 assign n1056 = ( Pg35  &  n1220 ) | ( n1220  &  (~ Ng4349) ) | ( Pg35  &  (~ n5248) ) | ( (~ Ng4349)  &  (~ n5248) ) ;
 assign Ng34258 = ( (~ n1056) ) ;
 assign n1057 = ( n2441  &  n2446  &  n2447 ) | ( n2446  &  n2447  &  (~ Ng1792) ) ;
 assign Ng32993 = ( (~ n1057) ) ;
 assign n1058 = ( n1849  &  n1847 ) | ( n1849  &  (~ Ng2084) ) ;
 assign Ng33992 = ( (~ n1058) ) ;
 assign n1059 = ( n3041  &  n3042  &  n160 ) | ( n3041  &  n3042  &  n3040 ) ;
 assign Ng30394 = ( (~ n1059) ) ;
 assign n1061 = ( (~ n4638)  &  Ng4311 ) | ( n4638  &  (~ Ng4311) ) ;
 assign Ng34449 = ( n1061  &  (~ n4641) ) ;
 assign n1062 = ( (~ n1260)  &  n1750  &  n1751 ) | ( n1750  &  n1751  &  n1749 ) ;
 assign Ng34019 = ( (~ n1062) ) ;
 assign n1063 = ( n3038  &  n3039  &  n160 ) | ( n3038  &  n3039  &  n3037 ) ;
 assign Ng30395 = ( (~ n1063) ) ;
 assign n1064 = ( n4202  &  n4203  &  Ng385 ) | ( n4202  &  n4203  &  n4201 ) ;
 assign Ng25598 = ( (~ n1064) ) ;
 assign n1065 = ( (~ n1265)  &  n1864  &  n1865 ) | ( n1864  &  n1865  &  n1863 ) ;
 assign Ng33987 = ( (~ n1065) ) ;
 assign n1066 = ( Pg35  &  n3065 ) | ( (~ Ng2523)  &  n3065 ) ;
 assign Ng30380 = ( (~ n1066) ) ;
 assign n1067 = ( n3023  &  n3024  &  n160 ) | ( n3023  &  n3024  &  n3022 ) ;
 assign Ng30400 = ( (~ n1067) ) ;
 assign n1068 = ( Pg35  &  n1487 ) | ( n1487  &  (~ Ng2960) ) ;
 assign Ng34623 = ( (~ n1068) ) ;
 assign n1069 = ( (~ Ng5689) ) | ( (~ n5145) ) ;
 assign Ng24343 = ( (~ Pg35)  &  Ng5694 ) | ( Ng5694  &  n1069 ) ;
 assign n1070 = ( n160  &  n2818  &  (~ n6341) ) | ( n2818  &  n2817  &  (~ n6341) ) ;
 assign Ng30473 = ( (~ n1070) ) ;
 assign n1071 = ( (~ Ng3518)  &  (~ Ng3522) ) | ( (~ Ng3522)  &  n2336 ) | ( (~ Ng3518)  &  n2338 ) | ( n2336  &  n2338 ) ;
 assign Ng33028 = ( (~ n1071) ) ;
 assign n1072 = ( (~ n2565)  &  n3591  &  (~ n5946) ) | ( n3591  &  (~ n5038)  &  (~ n5946) ) ;
 assign Ng29258 = ( (~ n1072) ) ;
 assign n1073 = ( n3002  &  n3003  &  n160 ) | ( n3002  &  n3003  &  n3001 ) ;
 assign Ng30407 = ( (~ n1073) ) ;
 assign n1074 = ( Pg35  &  n3920 ) | ( n3920  &  (~ Ng4455) ) ;
 assign Ng26958 = ( (~ n1074) ) ;
 assign n1075 = ( n1556  &  n1562  &  n1563 ) | ( (~ Ng4628)  &  n1562  &  n1563 ) ;
 assign Ng34457 = ( (~ n1075) ) ;
 assign n1076 = ( n1847  &  n2130 ) | ( n2130  &  (~ Ng1996) ) ;
 assign Ng33568 = ( (~ n1076) ) ;
 assign n1077 = ( Pg35  &  n3918  &  (~ n4367) ) | ( n3918  &  (~ Ng4527)  &  (~ n4367) ) ;
 assign Ng26964 = ( (~ n1077) ) ;
 assign n1078 = ( (~ Ng1724)  &  n3134  &  (~ n5875) ) | ( n3134  &  n3132  &  (~ n5875) ) ;
 assign Ng30352 = ( (~ n1078) ) ;
 assign n1079 = ( (~ Ng1379)  &  n2197 ) | ( (~ Ng1379)  &  (~ Ng1373) ) | ( n2197  &  (~ n5589) ) | ( (~ Ng1373)  &  (~ n5589) ) ;
 assign Ng33543 = ( (~ n1079) ) ;
 assign n1083 = ( (~ Pg16744)  &  (~ Pg13926) ) | ( (~ Pg16744)  &  Pg11388 ) | ( Pg13926  &  Pg11388 ) ;
 assign Ng24271 = ( Pg35  &  (~ Pg16656)  &  (~ Pg16627)  &  (~ Pg14451)  &  n1083 ) ;
 assign n1084 = ( (~ n1267)  &  n1887  &  n1888 ) | ( n1887  &  n1888  &  n1886 ) ;
 assign Ng33981 = ( (~ n1084) ) ;
 assign n1085 = ( Pg35  &  n2744 ) | ( n2744  &  (~ Ng5615) ) ;
 assign Ng30500 = ( (~ n1085) ) ;
 assign n1086 = ( Pg35  &  Ng5845 ) | ( Pg35  &  Ng5831 ) ;
 assign n1090 = ( Ng2724 ) | ( Ng2729 ) ;
 assign n1088 = ( n4551  &  Ng2735 ) ;
 assign n1087 = ( n1090  &  (~ n4868) ) | ( n1088  &  (~ Ng2771)  &  (~ n4868) ) ;
 assign n1092 = ( n1327  &  n1328  &  n1329 ) ;
 assign Ng34992 = ( (~ n1092) ) ;
 assign n1094 = ( n4695 ) | ( (~ Ng1514) ) ;
 assign n1093 = ( Pg17423  &  n1094 ) | ( Pg17423  &  (~ Ng1526) ) ;
 assign n1096 = ( Pg17320  &  Ng1526 ) | ( Pg17320  &  n1094 ) ;
 assign n1099 = ( Ng4709 ) | ( (~ Ng4785) ) ;
 assign n1100 = ( n4556 ) | ( n4776 ) ;
 assign n1097 = ( Ng4674  &  n1099 ) | ( Ng4674  &  n1100 ) | ( Ng4674  &  (~ Ng4743) ) ;
 assign n1101 = ( (~ Ng3129)  &  (~ Ng3143) ) ;
 assign n1104 = ( n1090  &  (~ n4868) ) | ( n1088  &  (~ Ng2803)  &  (~ n4868) ) ;
 assign Ng34991 = ( (~ n981) ) ;
 assign n1107 = ( Ng4420 ) | ( Ng4427 ) ;
 assign n1108 = ( Pg35  &  Ng6537 ) | ( Pg35  &  Ng6523 ) ;
 assign n1110 = ( n4561 ) | ( n4777 ) ;
 assign n1111 = ( Ng4899 ) | ( Ng4975 ) | ( (~ Ng4888) ) ;
 assign n1109 = ( Ng4836  &  n1110 ) | ( Ng4836  &  n1111 ) ;
 assign n1112 = ( Pg35  &  Ng6191 ) | ( Pg35  &  Ng6177 ) ;
 assign n1114 = ( (~ Ng1183) ) | ( n4736 ) ;
 assign n1113 = ( Pg17400  &  n1114 ) | ( Pg17400  &  (~ Ng1171) ) ;
 assign n1118 = ( (~ Ng4899) ) | ( Ng4975 ) ;
 assign n1116 = ( Ng4871  &  n1110 ) | ( Ng4871  &  n1118 ) | ( Ng4871  &  (~ Ng4944) ) ;
 assign Ng34994 = ( (~ n204) ) ;
 assign Ng34990 = ( (~ n569) ) ;
 assign n1119 = ( n1347  &  n1348  &  n1349 ) ;
 assign Ng34993 = ( (~ n1119) ) ;
 assign n1120 = ( Pg17316  &  Ng1171 ) | ( Pg17316  &  n1114 ) ;
 assign n1121 = ( n1298  &  n1299  &  n1300 ) ;
 assign Ng34996 = ( (~ n1121) ) ;
 assign n1124 = ( n1223 ) | ( (~ Ng4180) ) ;
 assign n1122 = ( n1124  &  (~ n1258) ) | ( Ng1105  &  (~ n1258)  &  (~ Ng947) ) ;
 assign n1126 = ( n1090  &  (~ n4862) ) | ( n1088  &  (~ Ng2783)  &  (~ n4862) ) ;
 assign Ng34879 = ( (~ n1169) ) ;
 assign n1129 = ( n1639  &  n1640  &  n1641  &  n1642  &  n1643  &  n1644  &  n1645  &  n1646 ) ;
 assign n1131 = ( Pg35  &  Ng3480 ) | ( Pg35  &  Ng3494 ) ;
 assign n1132 = ( n1305  &  n1306  &  n1307  &  n1308 ) ;
 assign Ng34997 = ( (~ n1132) ) ;
 assign n1133 = ( Pg35  &  Ng5152 ) | ( Pg35  &  Ng5138 ) ;
 assign n1134 = ( Pg35  &  Ng3845 ) | ( Pg35  &  Ng3831 ) ;
 assign n1136 = ( Ng4899 ) | ( (~ Ng4975) ) ;
 assign n1135 = ( Ng4864  &  n1110 ) | ( Ng4864  &  n1136 ) | ( Ng4864  &  (~ Ng4933) ) ;
 assign n1139 = ( Ng1514 ) | ( n4695 ) ;
 assign n1138 = ( Pg17404  &  (~ Ng1526) ) | ( Pg17404  &  n1139 ) ;
 assign n1140 = ( Ng1430  &  Ng1526 ) | ( Ng1430  &  n1139 ) ;
 assign n1141 = ( n1314  &  n1315  &  n1316  &  n1317 ) ;
 assign Ng34995 = ( (~ n1141) ) ;
 assign n1142 = ( Ng1183 ) | ( n4736 ) ;
 assign n1145 = ( Ng4709 ) | ( Ng4785 ) | ( (~ Ng4698) ) ;
 assign n1146 = ( n1090  &  (~ n4689) ) | ( n1088  &  (~ Ng2787)  &  (~ n4689) ) ;
 assign Ng34847 = ( (~ n1168) ) ;
 assign n1150 = ( Pg35  &  Ng5499 ) | ( Pg35  &  Ng5485 ) ;
 assign n1151 = ( n1090  &  (~ n4862) ) | ( n1088  &  (~ Ng2815)  &  (~ n4862) ) ;
 assign n1153 = ( n1090  &  (~ n4689) ) | ( n1088  &  (~ Ng2819)  &  (~ n4689) ) ;
 assign n1155 = ( Ng1087  &  Ng1171 ) | ( Ng1087  &  n1142 ) ;
 assign n1158 = ( n1226 ) | ( (~ Ng4180) ) ;
 assign n1156 = ( n1158  &  (~ n1261) ) | ( Ng1300  &  (~ n1261)  &  (~ Ng1291) ) ;
 assign n1160 = ( (~ Pg134)  &  (~ Pg99) ) | ( (~ Pg134)  &  (~ Ng37) ) ;
 assign n1162 = ( n1090  &  (~ n4135) ) | ( n1088  &  (~ n4135)  &  (~ Ng2807) ) ;
 assign n1166 = ( (~ Ng4899) ) | ( (~ Ng4975) ) ;
 assign n1165 = ( n1110  &  Ng4878 ) | ( Ng4878  &  n1166 ) | ( Ng4878  &  (~ Ng4955) ) ;
 assign Ng34878 = ( (~ n1189) ) ;
 assign n1168 = ( n1409  &  n1406 ) | ( n1409  &  n1407 ) | ( n1409  &  n1408 ) ;
 assign n1169 = ( n1382  &  n1383  &  n1384  &  n1385  &  n1386  &  n1387 ) ;
 assign n1170 = ( n4509 ) | ( n4510 ) ;
 assign Ng21726 = ( (~ Pg35)  &  Ng2975 ) ;
 assign n1173 = ( (~ Ng528)  &  Ng490  &  Ng482 ) ;
 assign n1172 = ( Ng528  &  (~ n5057) ) | ( n1173  &  (~ n5057) ) ;
 assign n1176 = ( n1111  &  n1136  &  n1419 ) | ( n1111  &  n1419  &  (~ Ng4933) ) ;
 assign n1175 = ( wire4651  &  wire4658  &  (~ n1160)  &  n1176 ) ;
 assign Ng34848 = ( (~ n1401) ) ;
 assign n1178 = ( n1695  &  n1696  &  n1697  &  n1698  &  n1699  &  n1700  &  n1701  &  n1702 ) ;
 assign n1180 = ( (~ Ng4709) ) | ( Ng4785 ) ;
 assign n1179 = ( Ng4681  &  n1100 ) | ( Ng4681  &  n1180 ) | ( Ng4681  &  (~ Ng4754) ) ;
 assign n1182 = ( n1090  &  (~ n4135) ) | ( n1088  &  (~ n4135)  &  (~ Ng2775) ) ;
 assign n1184 = ( n1158  &  (~ n1264) ) | ( Ng1472  &  (~ n1264)  &  (~ Ng1291) ) ;
 assign Ng35002 = ( (~ n4486) ) ;
 assign n1187 = ( n1124  &  (~ n1266) ) | ( Ng956  &  (~ n1266)  &  (~ Ng947) ) ;
 assign n1189 = ( n1368  &  (~ n1388) ) | ( (~ n1388)  &  n1392  &  n1393 ) ;
 assign Ng34789 = ( (~ n6113) ) ;
 assign n1191 = ( n4596 ) | ( n4597 ) ;
 assign n1192 = ( n1124  &  (~ n1268) ) | ( Ng1129  &  (~ n1268)  &  (~ Ng947) ) ;
 assign n1195 = ( n1145  &  n1180  &  n1418 ) | ( n1145  &  n1418  &  (~ Ng4754) ) ;
 assign n1194 = ( wire4651  &  wire4658  &  (~ n1160)  &  n1195 ) ;
 assign n1197 = ( (~ Ng4709) ) | ( (~ Ng4785) ) ;
 assign n1196 = ( n1100  &  Ng4688 ) | ( Ng4688  &  n1197 ) | ( Ng4688  &  (~ Ng4765) ) ;
 assign n1199 = ( n1158  &  (~ n1270) ) | ( Ng1478  &  (~ n1270)  &  (~ Ng1291) ) ;
 assign n1201 = ( n1124  &  (~ n1272) ) | ( Ng1135  &  (~ n1272)  &  (~ Ng947) ) ;
 assign Ng25692 = ( (~ Pg35)  &  Ng4392 ) ;
 assign n1203 = ( n1158  &  (~ n1274) ) | ( Ng1448  &  (~ n1274)  &  (~ Ng1291) ) ;
 assign n1205 = ( wire4436  &  (~ Pg12368) ) | ( wire4436  &  Pg9048 ) ;
 assign n1209 = ( n1219  &  Pg7946  &  n1217 ) | ( n1219  &  Pg7946  &  n1218 ) ;
 assign n1211 = ( n3159  &  Pg7916  &  n4977 ) ;
 assign n1215 = ( (~ Ng528)  &  (~ Ng490)  &  (~ Ng499)  &  (~ n4492)  &  (~ Ng482)  &  (~ Ng518) ) ;
 assign n1216 = ( (~ Ng718)  &  n5640 ) | ( (~ Ng655)  &  n5640 ) | ( (~ Ng753)  &  n5640 ) ;
 assign n1212 = ( n1215  &  n1216  &  (~ Ng807) ) | ( n1215  &  n1216  &  (~ Ng554) ) ;
 assign n1219 = ( Ng1339  &  Ng1521  &  (~ Ng1532) ) ;
 assign n1217 = ( Ng1367  &  Ng1345  &  Ng1379  &  n4322 ) ;
 assign n1218 = ( Ng1351 ) | ( Ng1312 ) ;
 assign n1221 = ( (~ Pg113)  &  (~ n1160) ) ;
 assign n1222 = ( Pg72 ) | ( Pg73 ) ;
 assign n1220 = ( Ng65  &  n1221 ) | ( Ng65  &  n1222 ) ;
 assign n1224 = ( (~ Ng691) ) | ( Ng209 ) ;
 assign n1223 = ( (~ Pg134)  &  n1224 ) | ( (~ Pg134)  &  (~ n1411) ) ;
 assign n1226 = ( (~ Pg134)  &  n667 ) | ( (~ Pg134)  &  n1224 ) ;
 assign n1228 = ( n204  &  n1141 ) | ( (~ n204)  &  (~ n1141) ) ;
 assign n1229 = ( n1121  &  n1132 ) | ( (~ n1121)  &  (~ n1132) ) ;
 assign n1230 = ( (~ n204)  &  n1141 ) | ( n204  &  (~ n1141) ) ;
 assign n1231 = ( (~ n1121)  &  n1132 ) | ( n1121  &  (~ n1132) ) ;
 assign n1227 = ( n1228  &  n1230 ) | ( n1229  &  n1230 ) | ( n1228  &  n1231 ) | ( n1229  &  n1231 ) ;
 assign n1233 = ( n569  &  n981 ) | ( (~ n569)  &  (~ n981) ) ;
 assign n1234 = ( n1092  &  n1119 ) | ( (~ n1092)  &  (~ n1119) ) ;
 assign n1235 = ( (~ n569)  &  n981 ) | ( n569  &  (~ n981) ) ;
 assign n1236 = ( (~ n1092)  &  n1119 ) | ( n1092  &  (~ n1119) ) ;
 assign n1232 = ( n1233  &  n1235 ) | ( n1234  &  n1235 ) | ( n1233  &  n1236 ) | ( n1234  &  n1236 ) ;
 assign n1240 = ( n4176  &  n4177 ) ;
 assign n1238 = ( Ng225 ) | ( n4387 ) ;
 assign n1239 = ( (~ n4387) ) | ( (~ Ng225) ) ;
 assign n1237 = ( n1240  &  (~ n6174) ) | ( n1238  &  n1239  &  (~ n6174) ) ;
 assign Ng34787 = ( (~ n1195) ) ;
 assign Ng34786 = ( (~ n1176) ) ;
 assign n1242 = ( Ng2357 ) | ( Ng2491 ) | ( Ng2223 ) | ( Ng2472 ) | ( Ng2338 ) | ( Ng2606 ) | ( Ng2204 ) | ( Ng2625 ) ;
 assign n1243 = ( Ng2283 ) | ( Ng2685 ) | ( Ng2417 ) | ( Ng2537 ) | ( Ng2403 ) | ( Ng2269 ) | ( Ng2671 ) | ( Ng2551 ) ;
 assign n1245 = ( (~ Pg73)  &  (~ n2521) ) | ( Pg72  &  (~ n2521) ) ;
 assign n1248 = ( Pg73  &  (~ n2521) ) | ( (~ Pg72)  &  (~ n2521) ) ;
 assign n1250 = ( (~ Pg35)  &  (~ n1277) ) | ( (~ Pg35)  &  (~ n4418) ) ;
 assign n1253 = ( Ng4578  &  (~ n2521) ) ;
 assign n1255 = ( (~ Ng2756) ) | ( (~ Ng2748) ) | ( (~ Ng2735) ) | ( (~ Ng2741) ) ;
 assign n1256 = ( n4536  &  Pg35 ) ;
 assign n1254 = ( n1255  &  n1256  &  Ng2756 ) | ( n1255  &  n1256  &  Ng2748 ) ;
 assign n1258 = ( (~ Ng1105)  &  (~ n1223)  &  n1893 ) | ( (~ n1223)  &  Ng947  &  n1893 ) ;
 assign n1257 = ( Pg35  &  n1122 ) | ( Pg35  &  (~ wire4421)  &  n1258 ) ;
 assign n1261 = ( (~ Ng1300)  &  (~ n1226)  &  n1739 ) | ( (~ n1226)  &  n1739  &  Ng1291 ) ;
 assign n1260 = ( Pg35  &  n1156 ) | ( Pg35  &  n1261  &  (~ Ng1585) ) ;
 assign n1264 = ( (~ Ng1472)  &  (~ n1226)  &  n1765 ) | ( (~ n1226)  &  Ng1291  &  n1765 ) ;
 assign n1263 = ( Pg35  &  n1184 ) | ( Pg35  &  Ng1585  &  n1264 ) ;
 assign n1266 = ( (~ Ng956)  &  (~ n1223)  &  n1841 ) | ( (~ n1223)  &  n1841  &  Ng947 ) ;
 assign n1265 = ( Pg35  &  n1187 ) | ( Pg35  &  (~ wire4421)  &  n1266 ) ;
 assign n1268 = ( (~ Ng1129)  &  (~ n1223)  &  n1867 ) | ( (~ n1223)  &  Ng947  &  n1867 ) ;
 assign n1267 = ( Pg35  &  n1192 ) | ( Pg35  &  wire4421  &  n1268 ) ;
 assign n1270 = ( (~ Ng1478)  &  (~ n1226)  &  n1816 ) | ( (~ n1226)  &  Ng1291  &  n1816 ) ;
 assign n1269 = ( Pg35  &  n1199 ) | ( Pg35  &  n1270  &  Ng1585 ) ;
 assign n1272 = ( (~ Ng1135)  &  (~ n1223)  &  n1918 ) | ( (~ n1223)  &  Ng947  &  n1918 ) ;
 assign n1271 = ( Pg35  &  n1201 ) | ( Pg35  &  n1272  &  wire4421 ) ;
 assign n1274 = ( (~ Ng1448)  &  (~ n1226)  &  n1791 ) | ( (~ n1226)  &  Ng1291  &  n1791 ) ;
 assign n1273 = ( Pg35  &  n1203 ) | ( Pg35  &  (~ Ng1585)  &  n1274 ) ;
 assign n1278 = ( n1289  &  (~ Ng586) ) | ( (~ Ng758)  &  (~ Ng586) ) | ( n1289  &  n4419 ) | ( (~ Ng758)  &  n4419 ) ;
 assign n1279 = ( (~ n1250)  &  n1331  &  n5541 ) | ( (~ n1250)  &  (~ Ng613)  &  n5541 ) ;
 assign n1277 = ( n4403 ) | ( n4407 ) ;
 assign n1275 = ( n1278  &  n1279  &  n1277 ) | ( n1278  &  n1279  &  (~ Ng794) ) ;
 assign n1282 = ( n1294  &  n1323 ) | ( n1323  &  (~ Ng2950) ) | ( n1294  &  (~ Ng2955) ) | ( (~ Ng2950)  &  (~ Ng2955) ) ;
 assign n1283 = ( n1303  &  (~ Ng2868)  &  n5540 ) | ( n1303  &  n4406  &  n5540 ) ;
 assign n1281 = ( (~ Ng51) ) | ( n4404 ) | ( n4411 ) ;
 assign n1280 = ( (~ Ng37)  &  n1282  &  n1283 ) | ( n1282  &  n1283  &  n1281 ) ;
 assign n1284 = ( Ng4927  &  Ng4737 ) | ( n4433  &  Ng4737 ) | ( Ng4927  &  n4434 ) | ( n4433  &  n4434 ) ;
 assign n1285 = ( (~ Ng947)  &  (~ Ng4300) ) | ( n4428  &  (~ Ng4300) ) | ( (~ Ng947)  &  n4431 ) | ( n4428  &  n4431 ) ;
 assign n1286 = ( n1275  &  (~ Ng1291) ) | ( (~ Ng1291)  &  n4394 ) | ( n1275  &  n4426 ) | ( n4394  &  n4426 ) ;
 assign n1287 = ( (~ Ng4172)  &  n5543 ) | ( n4416  &  n5543 ) ;
 assign n1291 = ( n1277  &  (~ Ng568) ) | ( (~ Ng785)  &  (~ Ng568) ) | ( n1277  &  n4419 ) | ( (~ Ng785)  &  n4419 ) ;
 assign n1292 = ( (~ wire4426)  &  (~ n1250)  &  n5550 ) | ( (~ n1250)  &  n4421  &  n5550 ) ;
 assign n1289 = ( (~ Ng51) ) | ( n4407 ) | ( n4411 ) ;
 assign n1288 = ( n1291  &  n1292  &  n1289 ) | ( n1291  &  n1292  &  (~ Ng744) ) ;
 assign n1296 = ( (~ Pg127)  &  (~ Pg92) ) | ( (~ Pg127)  &  n1281 ) | ( (~ Pg92)  &  n4406 ) | ( n1281  &  n4406 ) ;
 assign n1297 = ( (~ Ng2975)  &  n5549 ) | ( n1323  &  n5549 ) ;
 assign n1294 = ( (~ n4398) ) | ( (~ Ng51) ) | ( n4407 ) ;
 assign n1293 = ( n1296  &  n1297  &  n1294 ) | ( n1296  &  n1297  &  (~ Ng2970) ) ;
 assign n1298 = ( n4416  &  n4431 ) | ( n4431  &  (~ Ng4146) ) | ( n4416  &  (~ Ng4249) ) | ( (~ Ng4146)  &  (~ Ng4249) ) ;
 assign n1299 = ( n1288  &  n4444 ) | ( n4394  &  n4444 ) | ( n1288  &  (~ Ng2697) ) | ( n4394  &  (~ Ng2697) ) ;
 assign n1300 = ( n4428  &  n5551  &  n5552 ) | ( (~ Ng939)  &  n5551  &  n5552 ) ;
 assign n1303 = ( n4397 ) | ( (~ n4398) ) | ( (~ Ng51) ) ;
 assign n1304 = ( n4406  &  n4449 ) | ( n4449  &  (~ Ng2890) ) | ( n4406  &  (~ Ng2984) ) | ( (~ Ng2890)  &  (~ Ng2984) ) ;
 assign n1301 = ( (~ Pg100)  &  n1303  &  n1304 ) | ( n1281  &  n1303  &  n1304 ) ;
 assign n1305 = ( n4426  &  n4428 ) | ( n4428  &  (~ Ng1287) ) | ( n4426  &  (~ Ng943) ) | ( (~ Ng1287)  &  (~ Ng943) ) ;
 assign n1306 = ( n4431  &  n4442 ) | ( n4442  &  (~ Ng4245) ) | ( n4431  &  (~ Ng2145) ) | ( (~ Ng4245)  &  (~ Ng2145) ) ;
 assign n1307 = ( n4416  &  n4444 ) | ( n4444  &  (~ Ng4157) ) | ( n4416  &  (~ Ng2704) ) | ( (~ Ng4157)  &  (~ Ng2704) ) ;
 assign n1308 = ( n5557  &  n4394 ) | ( n5557  &  n5556  &  n5553 ) ;
 assign n1312 = ( n1294  &  n1323 ) | ( n1294  &  (~ Ng2965) ) | ( n1323  &  (~ Ng2960) ) | ( (~ Ng2965)  &  (~ Ng2960) ) ;
 assign n1313 = ( (~ wire4433)  &  n4406 ) | ( n1281  &  n4406 ) | ( (~ wire4433)  &  (~ Ng2873) ) | ( n1281  &  (~ Ng2873) ) ;
 assign n1310 = ( (~ Ng48) ) | ( n4402 ) | ( n4407 ) ;
 assign n1309 = ( n1312  &  n1313  &  n1310 ) | ( n1312  &  n1313  &  (~ Ng2878) ) ;
 assign n1314 = ( n4428  &  (~ Ng2689) ) | ( n4428  &  n4444 ) | ( (~ Ng2689)  &  Ng952 ) | ( n4444  &  Ng952 ) ;
 assign n1315 = ( n4416  &  (~ Ng2130) ) | ( (~ Ng4176)  &  (~ Ng2130) ) | ( n4416  &  n4442 ) | ( (~ Ng4176)  &  n4442 ) ;
 assign n1316 = ( n4426  &  n4431 ) | ( n4426  &  (~ Ng4253) ) | ( n4431  &  Ng1296 ) | ( (~ Ng4253)  &  Ng1296 ) ;
 assign n1317 = ( n5548  &  n4394 ) | ( n5548  &  n5547  &  n5544 ) ;
 assign n1320 = ( (~ Ng582)  &  n4421 ) | ( n4419  &  n4421 ) | ( (~ Ng582)  &  (~ Ng546) ) | ( n4419  &  (~ Ng546) ) ;
 assign n1321 = ( (~ n1250)  &  n1331  &  n5564 ) | ( (~ n1250)  &  (~ Ng622)  &  n5564 ) ;
 assign n1318 = ( n1289  &  n1320  &  n1321 ) | ( n1320  &  n1321  &  (~ Ng767) ) ;
 assign n1325 = ( n1310  &  n1351 ) | ( n1351  &  (~ Ng2864) ) | ( n1310  &  (~ Ng2860) ) | ( (~ Ng2864)  &  (~ Ng2860) ) ;
 assign n1326 = ( n1294  &  n4406 ) | ( n4406  &  (~ Ng2922) ) | ( n1294  &  Ng2994 ) | ( (~ Ng2922)  &  Ng2994 ) ;
 assign n1323 = ( (~ n4398) ) | ( Ng51 ) | ( n4407 ) ;
 assign n1322 = ( n1325  &  n1326  &  n1323 ) | ( n1325  &  n1326  &  (~ Ng2927) ) ;
 assign n1327 = ( n4433  &  n4444 ) | ( n4444  &  (~ Ng4907) ) | ( n4433  &  (~ Ng3151) ) | ( (~ Ng4907)  &  (~ Ng3151) ) ;
 assign n1328 = ( n1318  &  n4434 ) | ( n4394  &  n4434 ) | ( n1318  &  (~ Ng4717) ) | ( n4394  &  (~ Ng4717) ) ;
 assign n1329 = ( n5565  &  n5566  &  n1322 ) | ( n5565  &  n5566  &  n4394 ) ;
 assign n1333 = ( Pg35  &  (~ Ng595) ) | ( Pg35  &  n4419 ) | ( (~ Ng595)  &  n4418 ) | ( n4419  &  n4418 ) ;
 assign n1334 = ( n1289  &  n4421 ) | ( (~ Ng776)  &  n4421 ) | ( n1289  &  (~ Ng538) ) | ( (~ Ng776)  &  (~ Ng538) ) ;
 assign n1331 = ( n4397 ) | ( n4417 ) ;
 assign n1330 = ( n1333  &  n1334  &  n1331 ) | ( n1333  &  n1334  &  (~ Ng632) ) ;
 assign n1335 = ( n4434  &  n4442 ) | ( n4434  &  (~ Ng6199) ) | ( n4442  &  (~ Ng4727) ) | ( (~ Ng6199)  &  (~ Ng4727) ) ;
 assign n1336 = ( n4433  &  n4444 ) | ( n4433  &  (~ Ng3853) ) | ( n4444  &  (~ Ng4917) ) | ( (~ Ng3853)  &  (~ Ng4917) ) ;
 assign n1337 = ( n1330  &  n4412 ) | ( n4394  &  n4412 ) | ( n1330  &  (~ Ng45) ) | ( n4394  &  (~ Ng45) ) ;
 assign n1338 = ( n5560  &  n4394 ) | ( n5560  &  n5559  &  n5558 ) ;
 assign n1341 = ( n1277  &  (~ Ng577) ) | ( (~ Ng807)  &  (~ Ng577) ) | ( n1277  &  n4419 ) | ( (~ Ng807)  &  n4419 ) ;
 assign n1342 = ( (~ n1250)  &  n4421  &  n5568 ) | ( (~ n1250)  &  (~ Ng542)  &  n5568 ) ;
 assign n1339 = ( n1289  &  n1341  &  n1342 ) | ( n1341  &  n1342  &  (~ Ng763) ) ;
 assign n1345 = ( n1294  &  n1351 ) | ( n1294  &  (~ Ng2894) ) | ( n1351  &  (~ Ng2936) ) | ( (~ Ng2894)  &  (~ Ng2936) ) ;
 assign n1346 = ( n1303  &  n4406  &  n5567 ) | ( n1303  &  (~ Ng2988)  &  n5567 ) ;
 assign n1343 = ( n1323  &  n1345  &  n1346 ) | ( n1345  &  n1346  &  (~ Ng2941) ) ;
 assign n1347 = ( n1339  &  n4434 ) | ( n4394  &  n4434 ) | ( n1339  &  (~ Ng4722) ) | ( n4394  &  (~ Ng4722) ) ;
 assign n1348 = ( n4442  &  n4444 ) | ( n4444  &  (~ Ng5160) ) | ( n4442  &  (~ Ng6545) ) | ( (~ Ng5160)  &  (~ Ng6545) ) ;
 assign n1349 = ( n5569  &  n5570  &  n1343 ) | ( n5569  &  n5570  &  n4394 ) ;
 assign n1353 = ( n1310  &  n1323 ) | ( n1310  &  (~ Ng2917) ) | ( n1323  &  (~ Ng2856) ) | ( (~ Ng2917)  &  (~ Ng2856) ) ;
 assign n1354 = ( n1294  &  n4406 ) | ( n1294  &  (~ Ng2999) ) | ( n4406  &  (~ Ng2912) ) | ( (~ Ng2999)  &  (~ Ng2912) ) ;
 assign n1351 = ( (~ Ng48) ) | ( n4407 ) | ( n4414 ) ;
 assign n1350 = ( n1353  &  n1354  &  n1351 ) | ( n1353  &  n1354  &  (~ Ng2852) ) ;
 assign n1355 = ( n4433  &  n4444 ) | ( n4444  &  (~ Ng4922) ) | ( n4433  &  (~ Ng3502) ) | ( (~ Ng4922)  &  (~ Ng3502) ) ;
 assign n1356 = ( n4434  &  n4442 ) | ( n4442  &  (~ Ng4732) ) | ( n4434  &  (~ Ng5853) ) | ( (~ Ng4732)  &  (~ Ng5853) ) ;
 assign n1357 = ( n1350  &  n4412 ) | ( n4394  &  n4412 ) | ( n1350  &  (~ Ng46) ) | ( n4394  &  (~ Ng46) ) ;
 assign n1358 = ( n5563  &  n4394 ) | ( n5563  &  n5562  &  n5561 ) ;
 assign n1362 = ( (~ n1232)  &  n1227 ) | ( n1232  &  (~ n1227) ) ;
 assign n1359 = ( n1362  &  (~ Ng55) ) | ( (~ Pg56)  &  Pg54  &  n1362 ) ;
 assign n1363 = ( Pg56  &  (~ n1362)  &  Ng55 ) | ( (~ Pg54)  &  (~ n1362)  &  Ng55 ) ;
 assign n1366 = ( (~ Pg56)  &  (~ Pg54)  &  (~ Pg53)  &  (~ n4486) ) ;
 assign n1368 = ( Ng4311 ) | ( n4487 ) | ( n4488 ) ;
 assign n1369 = ( (~ Pg12184)  &  n1212 ) | ( Pg11678  &  n1212 ) ;
 assign n1372 = ( Pg35  &  n3791 ) | ( (~ Ng807)  &  n3791 ) | ( Pg35  &  (~ Ng554) ) | ( (~ Ng807)  &  (~ Ng554) ) ;
 assign n1371 = ( (~ Ng794) ) | ( n1395 ) ;
 assign n1376 = ( Ng4584  &  n5644 ) | ( (~ Ng4608)  &  n5644 ) | ( Ng4593  &  n5644 ) ;
 assign n1374 = ( (~ Ng4584)  &  Ng4608 ) | ( Ng4584  &  (~ Ng4608) ) ;
 assign n1375 = ( (~ Ng4601)  &  Ng4593 ) | ( Ng4601  &  (~ Ng4593) ) ;
 assign n1373 = ( n1376  &  Ng4616 ) | ( n1376  &  n1374 ) | ( n1376  &  n1375 ) ;
 assign n1377 = ( (~ n1371) ) | ( (~ Ng807) ) | ( n3791 ) ;
 assign n1378 = ( Pg35 ) | ( (~ Ng794) ) ;
 assign n1380 = ( (~ Ng632) ) | ( (~ n1379) ) | ( n4508 ) ;
 assign n1381 = ( Pg35 ) | ( (~ Ng626) ) ;
 assign n1379 = ( (~ Ng626) ) | ( n1398 ) ;
 assign n1382 = ( n4309 ) | ( n1642 ) ;
 assign n1383 = ( n1640 ) | ( Ng2040 ) | ( (~ Ng2070) ) ;
 assign n1384 = ( n1645 ) | ( Ng1906 ) | ( (~ Ng1936) ) ;
 assign n1385 = ( n1644 ) | ( Ng2197 ) | ( (~ Ng2227) ) ;
 assign n1386 = ( n4319  &  n4321 ) | ( n1639  &  n4321 ) | ( n4319  &  n1641 ) | ( n1639  &  n1641 ) ;
 assign n1387 = ( n4311  &  n4307 ) | ( n1643  &  n4307 ) | ( n4311  &  n1646 ) | ( n1643  &  n1646 ) ;
 assign n1388 = ( (~ n1406)  &  (~ n5571) ) | ( (~ n1406)  &  (~ n5572) ) ;
 assign n1392 = ( n1014  &  n4521 ) | ( n3263  &  n4521 ) | ( n1014  &  n4527 ) | ( n3263  &  n4527 ) ;
 assign n1393 = ( n4515  &  n4518 ) | ( n3371  &  n4518 ) | ( n4515  &  n3316 ) | ( n3371  &  n3316 ) ;
 assign n1396 = ( (~ Ng794) ) | ( (~ n1395) ) | ( n3791 ) ;
 assign n1397 = ( Pg35 ) | ( (~ Ng790) ) ;
 assign n1395 = ( (~ Ng790) ) | ( n1412 ) ;
 assign n1399 = ( (~ Ng626) ) | ( (~ n1398) ) | ( n4508 ) ;
 assign n1400 = ( Pg35 ) | ( (~ Ng622) ) ;
 assign n1398 = ( (~ Ng622) ) | ( n1415 ) ;
 assign n1402 = ( n4550  &  n4553 ) | ( n1698  &  n4553 ) | ( n4550  &  n1702 ) | ( n1698  &  n1702 ) ;
 assign n1403 = ( n4546  &  n4548 ) | ( n1695  &  n4548 ) | ( n4546  &  n1697 ) | ( n1695  &  n1697 ) ;
 assign n1404 = ( n4542  &  n4544 ) | ( n1701  &  n4544 ) | ( n4542  &  n1700 ) | ( n1701  &  n1700 ) ;
 assign n1405 = ( n4535  &  n4538 ) | ( n1699  &  n4538 ) | ( n4535  &  n1696 ) | ( n1699  &  n1696 ) ;
 assign n1401 = ( n1402  &  n1403  &  n1404  &  n1405 ) ;
 assign n1409 = ( n1368 ) | ( n3853 ) | ( n4304 ) ;
 assign n1406 = ( (~ Ng4311) ) | ( n4487 ) | ( n4488 ) ;
 assign n1407 = ( n1166 ) | ( n4564 ) ;
 assign n1408 = ( (~ Ng4878) ) | ( n4561 ) ;
 assign n1410 = ( Ng2389 ) | ( Ng2657 ) | ( Ng2523 ) | ( Ng2255 ) ;
 assign n1411 = ( Ng1193  &  Ng969 ) | ( Ng1193  &  Ng1008 ) ;
 assign n1413 = ( (~ Ng790) ) | ( (~ n1412) ) | ( n3791 ) ;
 assign n1414 = ( Pg35 ) | ( (~ Ng785) ) ;
 assign n1412 = ( (~ Ng785) ) | ( n1436 ) ;
 assign n1416 = ( (~ Ng622) ) | ( (~ n1415) ) | ( n4508 ) ;
 assign n1417 = ( Pg35 ) | ( (~ Ng617) ) ;
 assign n1415 = ( (~ Ng617) ) | ( n1439 ) ;
 assign n1418 = ( n1099  &  n1197 ) | ( n1197  &  (~ Ng4743) ) | ( n1099  &  (~ Ng4765) ) | ( (~ Ng4743)  &  (~ Ng4765) ) ;
 assign n1419 = ( n1118  &  n1166 ) | ( n1166  &  (~ Ng4944) ) | ( n1118  &  (~ Ng4955) ) | ( (~ Ng4944)  &  (~ Ng4955) ) ;
 assign n1421 = ( (~ Pg35) ) | ( (~ Ng2994) ) ;
 assign n1422 = ( (~ Pg35)  &  (~ n5079) ) | ( (~ Ng1287)  &  (~ n5079) ) ;
 assign n1425 = ( Pg35 ) | ( (~ Ng1283) ) ;
 assign n1426 = ( (~ Pg35)  &  n185 ) | ( n185  &  (~ Ng1296) ) ;
 assign n1428 = ( Pg35 ) | ( (~ Ng1291) ) ;
 assign n1429 = ( (~ Pg35)  &  n182 ) | ( n182  &  (~ Ng943) ) ;
 assign n1432 = ( Pg35 ) | ( (~ Ng939) ) ;
 assign n1433 = ( (~ Pg35)  &  n184 ) | ( n184  &  (~ Ng952) ) ;
 assign n1435 = ( Pg35 ) | ( (~ Ng947) ) ;
 assign n1437 = ( (~ Ng785) ) | ( (~ n1436) ) | ( n3791 ) ;
 assign n1438 = ( Pg35 ) | ( (~ Ng781) ) ;
 assign n1436 = ( (~ Ng781) ) | ( n1521 ) ;
 assign n1440 = ( (~ Ng617) ) | ( (~ n1439) ) | ( n4508 ) ;
 assign n1441 = ( Pg35 ) | ( (~ Ng613) ) ;
 assign n1439 = ( (~ Ng613) ) | ( n1524 ) ;
 assign n1452 = ( (~ Pg35) ) | ( (~ Ng4927) ) ;
 assign n1454 = ( (~ Pg35) ) | ( (~ Ng4912) ) ;
 assign n1456 = ( (~ Pg35) ) | ( (~ Ng4907) ) ;
 assign n1458 = ( (~ Pg35) ) | ( (~ Ng4922) ) ;
 assign n1462 = ( (~ Pg35) ) | ( (~ Ng4737) ) ;
 assign n1464 = ( (~ Pg35) ) | ( (~ Ng4722) ) ;
 assign n1466 = ( (~ Pg35) ) | ( (~ Ng4717) ) ;
 assign n1468 = ( (~ Pg35) ) | ( (~ Ng4732) ) ;
 assign n1472 = ( (~ Pg35) ) | ( (~ Ng4245) ) ;
 assign n1474 = ( (~ Pg35) ) | ( (~ Ng4249) ) ;
 assign n1476 = ( (~ Pg35) ) | ( (~ Ng4253) ) ;
 assign n1478 = ( (~ Pg35) ) | ( (~ Ng4157) ) ;
 assign n1480 = ( (~ Pg35) ) | ( (~ Ng4146) ) ;
 assign n1485 = ( (~ Pg35) ) | ( (~ Ng2988) ) ;
 assign n1487 = ( (~ Pg35) ) | ( (~ Ng2970) ) ;
 assign n1489 = ( (~ Pg35) ) | ( (~ Ng2960) ) ;
 assign n1491 = ( (~ Pg35) ) | ( (~ Ng2950) ) ;
 assign n1493 = ( (~ Pg35) ) | ( (~ Ng2936) ) ;
 assign n1495 = ( (~ Pg35) ) | ( (~ Ng2922) ) ;
 assign n1497 = ( (~ Pg35) ) | ( (~ Ng2912) ) ;
 assign n1499 = ( (~ Pg35) ) | ( (~ Ng2907) ) ;
 assign n1501 = ( (~ Pg35) ) | ( (~ Ng2868) ) ;
 assign n1502 = ( (~ Pg35) ) | ( (~ Ng2873) ) ;
 assign n1505 = ( (~ Pg35)  &  n5704 ) | ( (~ Ng37)  &  n5704 ) ;
 assign n1507 = ( (~ Pg35) ) | ( (~ Ng2894) ) ;
 assign n1508 = ( (~ Pg35) ) | ( (~ Ng2860) ) ;
 assign n1510 = ( (~ Pg35) ) | ( (~ Ng2852) ) ;
 assign n1512 = ( (~ Pg35) ) | ( (~ Ng2844) ) ;
 assign n1514 = ( (~ Pg35) ) | ( (~ Ng2704) ) ;
 assign n1516 = ( (~ Pg35) ) | ( (~ Ng2697) ) ;
 assign n1518 = ( (~ Pg35) ) | ( (~ Ng2145) ) ;
 assign n1520 = ( (~ Pg35) ) | ( (~ Ng2138) ) ;
 assign n1522 = ( (~ Ng781) ) | ( (~ n1521) ) | ( n3791 ) ;
 assign n1523 = ( Pg35 ) | ( (~ Ng776) ) ;
 assign n1521 = ( (~ Ng776) ) | ( n1626 ) ;
 assign n1525 = ( (~ Ng613) ) | ( (~ n1524) ) | ( n4508 ) ;
 assign n1526 = ( Pg35 ) | ( (~ Ng608) ) ;
 assign n1524 = ( (~ Ng608) ) | ( n1629 ) ;
 assign n1531 = ( Pg35  &  n1533 ) | ( n1533  &  (~ Ng4854) ) | ( Pg35  &  (~ Ng4859) ) | ( (~ Ng4854)  &  (~ Ng4859) ) ;
 assign n1530 = ( (~ Ng4849) ) | ( n4632 ) ;
 assign n1532 = ( (~ n1530)  &  Ng4854 ) | ( n1530  &  (~ Ng4854) ) ;
 assign n1533 = ( (~ Pg35) ) | ( (~ n4630) ) ;
 assign n1537 = ( Ng4849 ) | ( (~ n4630) ) | ( n4632 ) ;
 assign n1541 = ( Pg35  &  n1543 ) | ( n1543  &  (~ Ng4664) ) | ( Pg35  &  (~ Ng4669) ) | ( (~ Ng4664)  &  (~ Ng4669) ) ;
 assign n1540 = ( (~ Ng4659) ) | ( n4635 ) ;
 assign n1542 = ( (~ n1540)  &  Ng4664 ) | ( n1540  &  (~ Ng4664) ) ;
 assign n1543 = ( (~ Pg35) ) | ( (~ n4633) ) ;
 assign n1547 = ( Ng4659 ) | ( (~ n4633) ) | ( n4635 ) ;
 assign n1549 = ( n1220 ) | ( Ng4643 ) ;
 assign n1548 = ( Pg35  &  Ng4621 ) | ( Pg35  &  n1549 ) ;
 assign n1551 = ( Ng4639 ) | ( n1557 ) ;
 assign n1552 = ( (~ n1220)  &  (~ Ng4621) ) | ( (~ n1220)  &  Ng4639 ) | ( (~ n1220)  &  (~ Ng4628) ) ;
 assign n1555 = ( (~ n1220)  &  Ng4340 ) ;
 assign n1557 = ( (~ Pg35) ) | ( n1549 ) ;
 assign n1556 = ( n1551  &  Ng4621 ) | ( n1551  &  n1557 ) ;
 assign n1558 = ( n1556  &  Ng4628 ) | ( n1556  &  n1557 ) ;
 assign n1560 = ( (~ Ng4621) ) | ( n1549 ) ;
 assign n1559 = ( Pg35  &  Ng4633 ) | ( Pg35  &  (~ Ng4639) ) | ( Pg35  &  n1560 ) ;
 assign n1562 = ( (~ Ng4639) ) | ( Ng4628 ) | ( n1560 ) ;
 assign n1563 = ( Pg35 ) | ( (~ Ng4621) ) ;
 assign n1564 = ( (~ n1220)  &  (~ Ng4616) ) | ( (~ n1220)  &  (~ n4640) ) ;
 assign n1570 = ( Pg35  &  (~ Ng4616) ) | ( Pg35  &  n1579 ) | ( (~ Ng4616)  &  (~ Ng4608) ) | ( n1579  &  (~ Ng4608) ) ;
 assign n1569 = ( (~ Ng4601) ) | ( n4300 ) ;
 assign n1574 = ( Pg35  &  (~ Ng4332) ) | ( (~ Ng4332)  &  (~ Ng4322) ) | ( Pg35  &  n4641 ) | ( (~ Ng4322)  &  n4641 ) ;
 assign n1572 = ( n1220 ) | ( n4301 ) ;
 assign n1576 = ( (~ n1569) ) | ( n1579 ) | ( (~ Ng4608) ) ;
 assign n1577 = ( (~ n1564) ) | ( n1569 ) | ( Ng4608 ) ;
 assign n1578 = ( (~ Ng4601)  &  n4300 ) | ( Ng4601  &  (~ n4300) ) ;
 assign n1579 = ( (~ Pg35) ) | ( (~ n1564) ) ;
 assign n1582 = ( n1579 ) | ( (~ Ng4593) ) | ( n4640 ) ;
 assign n1583 = ( (~ n1564) ) | ( Ng4593 ) | ( (~ n4640) ) ;
 assign n1584 = ( n4301  &  Ng4584 ) | ( (~ n4301)  &  (~ Ng4584) ) ;
 assign n1587 = ( (~ Ng4322) ) | ( n4641 ) | ( n4642 ) ;
 assign n1588 = ( n1572 ) | ( Ng4322 ) | ( (~ n4642) ) ;
 assign n1589 = ( (~ Pg35)  &  (~ n4794) ) | ( Ng2827  &  (~ n4794) ) ;
 assign n1593 = ( (~ Pg35)  &  n5717 ) | ( (~ n1592)  &  n5717 ) | ( (~ Ng2819)  &  n5717 ) ;
 assign n1591 = ( n1221  &  Ng111 ) ;
 assign n1592 = ( n1255 ) | ( (~ Ng2724) ) | ( (~ Ng2729) ) ;
 assign n1594 = ( (~ Pg35)  &  (~ n4794) ) | ( Ng2811  &  (~ n4794) ) ;
 assign n1596 = ( (~ Pg35)  &  n5719 ) | ( (~ n1595)  &  n5719 ) | ( (~ Ng2807)  &  n5719 ) ;
 assign n1595 = ( n1255 ) | ( (~ Ng2724) ) | ( Ng2729 ) ;
 assign n1597 = ( (~ Pg35)  &  (~ n4794) ) | ( Ng2823  &  (~ n4794) ) ;
 assign n1599 = ( (~ Pg35)  &  n5721 ) | ( (~ n1598)  &  n5721 ) | ( (~ Ng2815)  &  n5721 ) ;
 assign n1598 = ( n1255 ) | ( Ng2724 ) | ( (~ Ng2729) ) ;
 assign n1600 = ( (~ Pg35)  &  (~ n4794) ) | ( Ng2799  &  (~ n4794) ) ;
 assign n1602 = ( (~ Pg35)  &  n5723 ) | ( (~ n1601)  &  n5723 ) | ( (~ Ng2803)  &  n5723 ) ;
 assign n1601 = ( n1255 ) | ( n1090 ) ;
 assign n1603 = ( (~ Pg35)  &  (~ n4794) ) | ( Ng2795  &  (~ n4794) ) ;
 assign n1605 = ( (~ Pg35)  &  n5724 ) | ( (~ n1592)  &  n5724 ) | ( (~ Ng2787)  &  n5724 ) ;
 assign n1604 = ( n1221  &  Ng85 ) ;
 assign n1606 = ( (~ Pg35)  &  (~ n4794) ) | ( Ng2779  &  (~ n4794) ) ;
 assign n1607 = ( (~ Pg35)  &  n5725 ) | ( (~ n1595)  &  n5725 ) | ( (~ Ng2775)  &  n5725 ) ;
 assign n1608 = ( (~ Pg35)  &  (~ n4794) ) | ( Ng2791  &  (~ n4794) ) ;
 assign n1609 = ( (~ Pg35)  &  n5726 ) | ( (~ n1598)  &  n5726 ) | ( (~ Ng2783)  &  n5726 ) ;
 assign n1610 = ( (~ Pg35)  &  (~ n4794) ) | ( Ng2767  &  (~ n4794) ) ;
 assign n1611 = ( (~ Pg35)  &  n5727 ) | ( (~ n1601)  &  n5727 ) | ( (~ Ng2771)  &  n5727 ) ;
 assign n1613 = ( Ng182  &  n5730 ) | ( (~ Ng182)  &  (~ n5730) ) ;
 assign n1614 = ( (~ Ng392)  &  (~ Ng411) ) | ( Ng392  &  (~ Ng441) ) | ( (~ Ng411)  &  (~ Ng441) ) ;
 assign n1612 = ( n1613  &  n1614  &  (~ Ng691)  &  (~ Ng417) ) ;
 assign n1617 = ( (~ n642)  &  n643  &  (~ Ng703) ) ;
 assign n1621 = ( Ng376  &  Ng385  &  Pg8719 ) ;
 assign n1620 = ( Ng896  &  n1621 ) | ( Ng896  &  n1617 ) ;
 assign n1622 = ( (~ Ng890)  &  n1620 ) | ( (~ Ng896)  &  n1620 ) | ( (~ Ng890)  &  (~ Ng862) ) | ( (~ Ng896)  &  (~ Ng862) ) ;
 assign n1627 = ( (~ Ng776) ) | ( (~ n1626) ) | ( n3791 ) ;
 assign n1628 = ( Pg35 ) | ( (~ Ng772) ) ;
 assign n1626 = ( (~ Ng772) ) | ( n1682 ) ;
 assign n1631 = ( Pg35 ) | ( (~ Ng604) ) ;
 assign n1629 = ( (~ Ng604) ) | ( n1685 ) ;
 assign n1635 = ( (~ Ng4141)  &  (~ Ng4082) ) ;
 assign n1633 = ( Ng4093 ) | ( Ng4098 ) ;
 assign n1634 = ( (~ Ng4076) ) | ( (~ Ng4112) ) ;
 assign n1632 = ( n1635  &  Ng4087 ) | ( n1635  &  n1633 ) | ( n1635  &  n1634 ) ;
 assign n1638 = ( Pg113  &  (~ n1160) ) ;
 assign n1636 = ( (~ n1368)  &  n1638 ) | ( (~ n1406)  &  n1638 ) ;
 assign n1639 = ( Ng528 ) | ( n4511 ) | ( (~ Ng504) ) ;
 assign n1640 = ( Ng504 ) | ( Ng528 ) | ( n4512 ) ;
 assign n1641 = ( Ng504 ) | ( Ng528 ) | ( n4511 ) ;
 assign n1642 = ( (~ Ng528) ) | ( (~ Ng504) ) | ( n4512 ) ;
 assign n1643 = ( (~ Ng528) ) | ( n4511 ) | ( (~ Ng504) ) ;
 assign n1644 = ( (~ Ng528) ) | ( n4511 ) | ( Ng504 ) ;
 assign n1645 = ( Ng528 ) | ( (~ Ng504) ) | ( n4512 ) ;
 assign n1646 = ( (~ Ng528) ) | ( Ng504 ) | ( n4512 ) ;
 assign n1647 = ( (~ Ng4961)  &  (~ n4653) ) | ( (~ n4652)  &  (~ n4653) ) ;
 assign n1651 = ( (~ n4652)  &  (~ n4653) ) | ( (~ Ng4950)  &  (~ n4653) ) ;
 assign n1653 = ( (~ Pg35)  &  (~ n4652) ) | ( (~ Pg35)  &  (~ Ng4939) ) | ( (~ n4652)  &  (~ n4653) ) | ( (~ Ng4939)  &  (~ n4653) ) ;
 assign n1656 = ( Pg35 ) | ( (~ Ng4939) ) ;
 assign n1657 = ( (~ Pg35) ) | ( (~ n1655) ) | ( (~ Ng4933) ) ;
 assign n1655 = ( n3830  &  n4652 ) ;
 assign n1658 = ( (~ n4652)  &  (~ n4653) ) | ( (~ n4653)  &  (~ Ng4894) ) ;
 assign n1663 = ( n4654 ) | ( (~ Ng101) ) ;
 assign n1660 = ( n1663  &  (~ Ng4771) ) | ( n1663  &  (~ n4654) ) ;
 assign n1664 = ( n1663  &  (~ n4654) ) | ( n1663  &  (~ Ng4760) ) ;
 assign n1666 = ( (~ Pg35)  &  (~ n4654) ) | ( n1663  &  (~ n4654) ) | ( (~ Pg35)  &  (~ Ng4749) ) | ( n1663  &  (~ Ng4749) ) ;
 assign n1669 = ( Pg35 ) | ( (~ Ng4749) ) ;
 assign n1670 = ( (~ Pg35) ) | ( (~ n1668) ) | ( (~ Ng4743) ) ;
 assign n1668 = ( n3847  &  n4654 ) ;
 assign n1671 = ( n1663  &  (~ n4654) ) | ( n1663  &  (~ Ng4704) ) ;
 assign n1675 = ( n1160  &  (~ n1222) ) | ( (~ n1222)  &  Ng4507 ) ;
 assign n1679 = ( n1675 ) | ( Ng4477 ) | ( (~ Ng26960) ) ;
 assign n1677 = ( Ng4462  &  n1679  &  (~ Ng4459) ) | ( n1679  &  (~ Ng4473)  &  (~ Ng4459) ) ;
 assign n1681 = ( Pg35  &  Ng4462  &  (~ Ng10384)  &  Ng4643 ) ;
 assign n1683 = ( (~ Ng772) ) | ( (~ n1682) ) | ( n3791 ) ;
 assign n1684 = ( Pg35 ) | ( (~ Ng767) ) ;
 assign n1682 = ( (~ Ng767) ) | ( n1942 ) ;
 assign n1687 = ( Pg35 ) | ( (~ Ng599) ) ;
 assign n1685 = ( (~ Ng599) ) | ( n1945 ) ;
 assign n1689 = ( Ng142 ) | ( n4664 ) ;
 assign n1690 = ( n3904 ) | ( (~ n4664) ) | ( (~ Ng142) ) ;
 assign n1691 = ( n359  &  Ng182 ) | ( n359  &  Ng174 ) | ( n359  &  Ng168 ) ;
 assign n1693 = ( Ng160 ) | ( n5754 ) ;
 assign n1694 = ( (~ Ng160) ) | ( n3182 ) | ( (~ n5754) ) ;
 assign n1695 = ( (~ Ng2756) ) | ( Ng2741 ) | ( n4540 ) ;
 assign n1696 = ( n4530 ) | ( n4536 ) ;
 assign n1697 = ( (~ Ng2741) ) | ( n4533 ) ;
 assign n1698 = ( (~ Ng2756) ) | ( (~ Ng2741) ) | ( n4540 ) ;
 assign n1699 = ( Ng2741 ) | ( n4533 ) ;
 assign n1700 = ( Ng2741 ) | ( Ng2756 ) | ( n4540 ) ;
 assign n1701 = ( Ng2756 ) | ( (~ Ng2741) ) | ( n4540 ) ;
 assign n1702 = ( n4530 ) | ( (~ n4551) ) ;
 assign n1703 = ( (~ n1408)  &  Ng4983 ) | ( n1408  &  (~ Ng4983) ) ;
 assign n1704 = ( (~ Pg35) ) | ( n1711 ) ;
 assign n1706 = ( (~ Pg35)  &  n1136 ) | ( n1118  &  n1136 ) | ( (~ Pg35)  &  (~ n4674) ) | ( n1118  &  (~ n4674) ) ;
 assign n1709 = ( n1704  &  n1706 ) | ( n1706  &  (~ Ng4899) ) | ( n1704  &  n4673 ) | ( (~ Ng4899)  &  n4673 ) ;
 assign n1713 = ( Pg35  &  n1704 ) | ( Pg35  &  (~ Ng4966) ) | ( n1704  &  (~ Ng4991) ) | ( (~ Ng4966)  &  (~ Ng4991) ) ;
 assign n1710 = ( n1408 ) | ( (~ Ng4983) ) ;
 assign n1711 = ( n4673 ) | ( n4674 ) ;
 assign n1715 = ( Ng4991 ) | ( n1711 ) | ( n1710 ) ;
 assign n1716 = ( n1704 ) | ( (~ n1710) ) | ( (~ Ng4991) ) ;
 assign n1717 = ( Ng4975 ) | ( n4673 ) | ( (~ n4674) ) ;
 assign n1718 = ( Pg35 ) | ( (~ Ng4966) ) ;
 assign n1719 = ( (~ n4304)  &  Ng4793 ) | ( n4304  &  (~ Ng4793) ) ;
 assign n1720 = ( (~ Pg35) ) | ( n1727 ) ;
 assign n1722 = ( (~ Pg35)  &  n1099 ) | ( n1099  &  n1180 ) | ( (~ Pg35)  &  (~ n4677) ) | ( n1180  &  (~ n4677) ) ;
 assign n1725 = ( n1720  &  n1722 ) | ( n1722  &  (~ Ng4709) ) | ( n1720  &  n4676 ) | ( (~ Ng4709)  &  n4676 ) ;
 assign n1729 = ( Pg35  &  n1720 ) | ( Pg35  &  (~ Ng4776) ) | ( n1720  &  (~ Ng4801) ) | ( (~ Ng4776)  &  (~ Ng4801) ) ;
 assign n1726 = ( n4304 ) | ( (~ Ng4793) ) ;
 assign n1727 = ( n4676 ) | ( n4677 ) ;
 assign n1731 = ( Ng4801 ) | ( n1727 ) | ( n1726 ) ;
 assign n1732 = ( n1720 ) | ( (~ n1726) ) | ( (~ Ng4801) ) ;
 assign n1733 = ( Ng4785 ) | ( n4676 ) | ( (~ n4677) ) ;
 assign n1734 = ( Pg35 ) | ( (~ Ng4776) ) ;
 assign n1736 = ( (~ Pg35) ) | ( Ng2841 ) ;
 assign n1737 = ( (~ Pg35)  &  n5760 ) | ( (~ Ng2763)  &  n5760 ) | ( (~ n1735)  &  n5760 ) ;
 assign n1735 = ( (~ Ng2759) ) | ( n2023 ) ;
 assign n1739 = ( (~ Ng2689) ) | ( (~ Ng2697) ) | ( (~ Ng2704) ) ;
 assign n1742 = ( (~ n1260)  &  (~ n4699) ) | ( n4697  &  (~ n4699) ) | ( (~ n1260)  &  (~ Ng2567) ) | ( n4697  &  (~ Ng2567) ) ;
 assign n1743 = ( (~ n1156)  &  (~ n1261) ) | ( (~ n1156)  &  Ng1589 ) ;
 assign n1747 = ( (~ Pg35)  &  (~ Ng2629) ) | ( Pg35  &  (~ n5257) ) | ( (~ Ng2629)  &  (~ n5257) ) ;
 assign n1745 = ( (~ Pg35) ) | ( n4700 ) ;
 assign n1750 = ( Pg35 ) | ( (~ Ng2571) ) ;
 assign n1751 = ( (~ Pg35) ) | ( (~ n1749) ) | ( (~ Ng2583) ) ;
 assign n1749 = ( n4307 ) | ( (~ n4700) ) ;
 assign n1753 = ( Pg35 ) | ( (~ Ng2583) ) ;
 assign n1754 = ( (~ Pg35) ) | ( (~ Ng2579) ) | ( n4703 ) ;
 assign n1756 = ( Pg35 ) | ( (~ Ng2579) ) ;
 assign n1757 = ( (~ Pg35) ) | ( (~ n1755) ) | ( (~ Ng2575) ) ;
 assign n1755 = ( (~ Ng2629) ) | ( n4704 ) ;
 assign n1759 = ( Pg35 ) | ( (~ Ng2563) ) ;
 assign n1760 = ( (~ Pg35) ) | ( (~ n1758) ) | ( (~ Ng2571) ) ;
 assign n1758 = ( (~ Ng2599) ) | ( Ng2629 ) | ( (~ n4700) ) ;
 assign n1762 = ( Pg35 ) | ( (~ Ng2567) ) ;
 assign n1763 = ( (~ Pg35) ) | ( (~ n1761) ) | ( (~ Ng2563) ) ;
 assign n1761 = ( Ng2599 ) | ( n4704 ) ;
 assign n1765 = ( (~ Ng2689) ) | ( (~ Ng2697) ) | ( Ng2704 ) ;
 assign n1767 = ( (~ n1263)  &  (~ n4709) ) | ( n4707  &  (~ n4709) ) | ( (~ n1263)  &  (~ Ng2433) ) | ( n4707  &  (~ Ng2433) ) ;
 assign n1768 = ( (~ n1184)  &  (~ n1264) ) | ( (~ n1184)  &  (~ Ng1589) ) ;
 assign n1773 = ( (~ Pg35)  &  (~ Ng2495) ) | ( Pg35  &  (~ n5260) ) | ( (~ Ng2495)  &  (~ n5260) ) ;
 assign n1771 = ( (~ Pg35) ) | ( n4710 ) ;
 assign n1776 = ( Pg35 ) | ( (~ Ng2437) ) ;
 assign n1775 = ( n4309 ) | ( (~ n4710) ) ;
 assign n1779 = ( Pg35 ) | ( (~ Ng2449) ) ;
 assign n1780 = ( (~ Pg35) ) | ( (~ Ng2445) ) | ( n4713 ) ;
 assign n1782 = ( Pg35 ) | ( (~ Ng2445) ) ;
 assign n1783 = ( (~ Pg35) ) | ( (~ n1781) ) | ( (~ Ng2441) ) ;
 assign n1781 = ( (~ Ng2495) ) | ( n4714 ) ;
 assign n1785 = ( Pg35 ) | ( (~ Ng2429) ) ;
 assign n1786 = ( (~ Pg35) ) | ( (~ n1784) ) | ( (~ Ng2437) ) ;
 assign n1784 = ( (~ Ng2465) ) | ( Ng2495 ) | ( (~ n4710) ) ;
 assign n1788 = ( Pg35 ) | ( (~ Ng2433) ) ;
 assign n1789 = ( (~ Pg35) ) | ( (~ n1787) ) | ( (~ Ng2429) ) ;
 assign n1787 = ( Ng2465 ) | ( n4714 ) ;
 assign n1791 = ( (~ Ng2689) ) | ( Ng2697 ) | ( (~ Ng2704) ) ;
 assign n1793 = ( (~ n1273)  &  (~ n4719) ) | ( n4717  &  (~ n4719) ) | ( (~ n1273)  &  (~ Ng2299) ) | ( n4717  &  (~ Ng2299) ) ;
 assign n1794 = ( (~ n1203)  &  (~ n1274) ) | ( (~ n1203)  &  Ng1589 ) ;
 assign n1798 = ( (~ Pg35)  &  (~ Ng2361) ) | ( Pg35  &  (~ n5263) ) | ( (~ Ng2361)  &  (~ n5263) ) ;
 assign n1796 = ( (~ Pg35) ) | ( n4720 ) ;
 assign n1801 = ( Pg35 ) | ( (~ Ng2303) ) ;
 assign n1800 = ( n4311 ) | ( (~ n4720) ) ;
 assign n1804 = ( Pg35 ) | ( (~ Ng2315) ) ;
 assign n1805 = ( (~ Pg35) ) | ( (~ Ng2311) ) | ( n4723 ) ;
 assign n1807 = ( Pg35 ) | ( (~ Ng2311) ) ;
 assign n1808 = ( (~ Pg35) ) | ( (~ n1806) ) | ( (~ Ng2307) ) ;
 assign n1806 = ( (~ Ng2361) ) | ( n4724 ) ;
 assign n1810 = ( Pg35 ) | ( (~ Ng2295) ) ;
 assign n1811 = ( (~ Pg35) ) | ( (~ n1809) ) | ( (~ Ng2303) ) ;
 assign n1809 = ( (~ Ng2331) ) | ( Ng2361 ) | ( (~ n4720) ) ;
 assign n1813 = ( Pg35 ) | ( (~ Ng2299) ) ;
 assign n1814 = ( (~ Pg35) ) | ( (~ n1812) ) | ( (~ Ng2295) ) ;
 assign n1812 = ( Ng2331 ) | ( n4724 ) ;
 assign n1816 = ( (~ Ng2689) ) | ( Ng2697 ) | ( Ng2704 ) ;
 assign n1818 = ( (~ n1269)  &  (~ n4729) ) | ( n4727  &  (~ n4729) ) | ( (~ n1269)  &  (~ Ng2165) ) | ( n4727  &  (~ Ng2165) ) ;
 assign n1819 = ( (~ n1199)  &  (~ n1270) ) | ( (~ n1199)  &  (~ Ng1589) ) ;
 assign n1823 = ( (~ Pg35)  &  (~ Ng2227) ) | ( Pg35  &  (~ n5266) ) | ( (~ Ng2227)  &  (~ n5266) ) ;
 assign n1821 = ( (~ Pg35) ) | ( n4730 ) ;
 assign n1826 = ( Pg35 ) | ( (~ Ng2169) ) ;
 assign n1827 = ( (~ Pg35) ) | ( (~ n1825) ) | ( (~ Ng2181) ) ;
 assign n1825 = ( Ng2197 ) | ( n4731 ) ;
 assign n1829 = ( Pg35 ) | ( (~ Ng2181) ) ;
 assign n1830 = ( (~ Pg35) ) | ( (~ Ng2177) ) | ( n4734 ) ;
 assign n1832 = ( Pg35 ) | ( (~ Ng2177) ) ;
 assign n1833 = ( (~ Pg35) ) | ( (~ n1831) ) | ( (~ Ng2173) ) ;
 assign n1831 = ( n4731 ) | ( (~ Ng2153) ) ;
 assign n1835 = ( Pg35 ) | ( (~ Ng2161) ) ;
 assign n1836 = ( (~ Pg35) ) | ( (~ n1834) ) | ( (~ Ng2169) ) ;
 assign n1834 = ( (~ Ng2197) ) | ( Ng2227 ) | ( (~ n4730) ) ;
 assign n1838 = ( Pg35 ) | ( (~ Ng2165) ) ;
 assign n1839 = ( (~ Pg35) ) | ( (~ n1837) ) | ( (~ Ng2161) ) ;
 assign n1837 = ( Ng2197 ) | ( (~ n4730) ) | ( (~ Ng2153) ) ;
 assign n1841 = ( (~ Ng2130) ) | ( (~ Ng2138) ) | ( (~ Ng2145) ) ;
 assign n1844 = ( (~ n1265)  &  (~ n4740) ) | ( n4738  &  (~ n4740) ) | ( (~ n1265)  &  (~ Ng2008) ) | ( n4738  &  (~ Ng2008) ) ;
 assign n1845 = ( (~ n1187)  &  (~ n1266) ) | ( (~ n1187)  &  Ng1246 ) ;
 assign n1849 = ( (~ Pg35)  &  (~ Ng2070) ) | ( Pg35  &  (~ n5269) ) | ( (~ Ng2070)  &  (~ n5269) ) ;
 assign n1847 = ( (~ Pg35) ) | ( n4741 ) ;
 assign n1852 = ( Pg35 ) | ( (~ Ng2012) ) ;
 assign n1853 = ( (~ Pg35) ) | ( (~ n1851) ) | ( (~ Ng2024) ) ;
 assign n1851 = ( Ng2040 ) | ( n4742 ) ;
 assign n1855 = ( Pg35 ) | ( (~ Ng2024) ) ;
 assign n1856 = ( (~ Pg35) ) | ( (~ Ng2020) ) | ( n4745 ) ;
 assign n1858 = ( Pg35 ) | ( (~ Ng2020) ) ;
 assign n1859 = ( (~ Pg35) ) | ( (~ n1857) ) | ( (~ Ng2016) ) ;
 assign n1857 = ( n4742 ) | ( (~ Ng1996) ) ;
 assign n1861 = ( Pg35 ) | ( (~ Ng2004) ) ;
 assign n1862 = ( (~ Pg35) ) | ( (~ n1860) ) | ( (~ Ng2012) ) ;
 assign n1860 = ( (~ Ng2040) ) | ( Ng2070 ) | ( (~ n4741) ) ;
 assign n1864 = ( Pg35 ) | ( (~ Ng2008) ) ;
 assign n1865 = ( (~ Pg35) ) | ( (~ n1863) ) | ( (~ Ng2004) ) ;
 assign n1863 = ( Ng2040 ) | ( (~ n4741) ) | ( (~ Ng1996) ) ;
 assign n1867 = ( (~ Ng2130) ) | ( (~ Ng2138) ) | ( Ng2145 ) ;
 assign n1869 = ( (~ n1267)  &  (~ n4750) ) | ( n4748  &  (~ n4750) ) | ( (~ n1267)  &  (~ Ng1874) ) | ( n4748  &  (~ Ng1874) ) ;
 assign n1870 = ( (~ n1192)  &  (~ n1268) ) | ( (~ n1192)  &  (~ Ng1246) ) ;
 assign n1875 = ( (~ Pg35)  &  (~ Ng1936) ) | ( Pg35  &  (~ n5272) ) | ( (~ Ng1936)  &  (~ n5272) ) ;
 assign n1873 = ( (~ Pg35) ) | ( n4751 ) ;
 assign n1878 = ( Pg35 ) | ( (~ Ng1878) ) ;
 assign n1879 = ( (~ Pg35) ) | ( (~ n1877) ) | ( (~ Ng1890) ) ;
 assign n1877 = ( Ng1906 ) | ( n4752 ) ;
 assign n1881 = ( Pg35 ) | ( (~ Ng1890) ) ;
 assign n1882 = ( (~ Pg35) ) | ( (~ Ng1886) ) | ( n4755 ) ;
 assign n1884 = ( Pg35 ) | ( (~ Ng1886) ) ;
 assign n1885 = ( (~ Pg35) ) | ( (~ n1883) ) | ( (~ Ng1882) ) ;
 assign n1883 = ( n4752 ) | ( (~ Ng1862) ) ;
 assign n1887 = ( Pg35 ) | ( (~ Ng1870) ) ;
 assign n1888 = ( (~ Pg35) ) | ( (~ n1886) ) | ( (~ Ng1878) ) ;
 assign n1886 = ( (~ Ng1906) ) | ( Ng1936 ) | ( (~ n4751) ) ;
 assign n1890 = ( Pg35 ) | ( (~ Ng1874) ) ;
 assign n1891 = ( (~ Pg35) ) | ( (~ n1889) ) | ( (~ Ng1870) ) ;
 assign n1889 = ( Ng1906 ) | ( (~ n4751) ) | ( (~ Ng1862) ) ;
 assign n1893 = ( (~ Ng2130) ) | ( Ng2138 ) | ( (~ Ng2145) ) ;
 assign n1895 = ( (~ n1257)  &  (~ n4760) ) | ( n4758  &  (~ n4760) ) | ( (~ n1257)  &  (~ Ng1740) ) | ( n4758  &  (~ Ng1740) ) ;
 assign n1896 = ( (~ n1122)  &  (~ n1258) ) | ( (~ n1122)  &  Ng1246 ) ;
 assign n1900 = ( (~ Pg35)  &  (~ Ng1802) ) | ( Pg35  &  (~ n5275) ) | ( (~ Ng1802)  &  (~ n5275) ) ;
 assign n1898 = ( (~ Pg35) ) | ( n4761 ) ;
 assign n1903 = ( Pg35 ) | ( (~ Ng1744) ) ;
 assign n1902 = ( n4319 ) | ( (~ n4761) ) ;
 assign n1906 = ( Pg35 ) | ( (~ Ng1756) ) ;
 assign n1907 = ( (~ Pg35) ) | ( (~ Ng1752) ) | ( n4764 ) ;
 assign n1909 = ( Pg35 ) | ( (~ Ng1752) ) ;
 assign n1910 = ( (~ Pg35) ) | ( (~ n1908) ) | ( (~ Ng1748) ) ;
 assign n1908 = ( (~ Ng1802) ) | ( n4765 ) ;
 assign n1912 = ( Pg35 ) | ( (~ Ng1736) ) ;
 assign n1913 = ( (~ Pg35) ) | ( (~ n1911) ) | ( (~ Ng1744) ) ;
 assign n1911 = ( (~ Ng1772) ) | ( Ng1802 ) | ( (~ n4761) ) ;
 assign n1915 = ( Pg35 ) | ( (~ Ng1740) ) ;
 assign n1916 = ( (~ Pg35) ) | ( (~ n1914) ) | ( (~ Ng1736) ) ;
 assign n1914 = ( Ng1772 ) | ( n4765 ) ;
 assign n1918 = ( (~ Ng2130) ) | ( Ng2138 ) | ( Ng2145 ) ;
 assign n1920 = ( (~ n1271)  &  (~ n4770) ) | ( n4768  &  (~ n4770) ) | ( (~ n1271)  &  (~ Ng1604) ) | ( n4768  &  (~ Ng1604) ) ;
 assign n1921 = ( (~ n1201)  &  (~ n1272) ) | ( (~ n1201)  &  (~ Ng1246) ) ;
 assign n1925 = ( (~ Pg35)  &  (~ Ng1668) ) | ( Pg35  &  (~ n5278) ) | ( (~ Ng1668)  &  (~ n5278) ) ;
 assign n1923 = ( (~ Pg35) ) | ( n4771 ) ;
 assign n1928 = ( Pg35 ) | ( (~ Ng1608) ) ;
 assign n1929 = ( (~ Pg35) ) | ( (~ n1927) ) | ( (~ Ng1620) ) ;
 assign n1927 = ( n4321 ) | ( (~ n4771) ) ;
 assign n1931 = ( Pg35 ) | ( (~ Ng1620) ) ;
 assign n1932 = ( (~ Pg35) ) | ( (~ n1930) ) | ( (~ Ng1616) ) ;
 assign n1930 = ( Ng1592 ) | ( n4773 ) ;
 assign n1934 = ( Pg35 ) | ( (~ Ng1616) ) ;
 assign n1935 = ( (~ Pg35) ) | ( (~ n1933) ) | ( (~ Ng1612) ) ;
 assign n1933 = ( (~ Ng1668) ) | ( n4774 ) ;
 assign n1937 = ( Pg35 ) | ( (~ Ng1600) ) ;
 assign n1938 = ( (~ Pg35) ) | ( (~ n1936) ) | ( (~ Ng1608) ) ;
 assign n1936 = ( Ng1668 ) | ( n4773 ) ;
 assign n1940 = ( Pg35 ) | ( (~ Ng1604) ) ;
 assign n1941 = ( (~ Pg35) ) | ( (~ n1939) ) | ( (~ Ng1600) ) ;
 assign n1939 = ( Ng1636 ) | ( n4774 ) ;
 assign n1943 = ( (~ Ng767) ) | ( (~ n1942) ) | ( n3791 ) ;
 assign n1944 = ( Pg35 ) | ( (~ Ng763) ) ;
 assign n1942 = ( (~ Ng763) ) | ( n2218 ) ;
 assign n1947 = ( Pg35 ) | ( (~ Ng595) ) ;
 assign n1945 = ( (~ Ng595) ) | ( n2221 ) ;
 assign n1949 = ( Ng298 ) | ( n4663 ) ;
 assign n1950 = ( n3904 ) | ( (~ Ng298) ) | ( (~ n4663) ) ;
 assign n1952 = ( Ng157 ) | ( n4672 ) ;
 assign n1953 = ( n3182 ) | ( (~ Ng157) ) | ( (~ n4672) ) ;
 assign n1957 = ( (~ Pg35)  &  n1960 ) | ( n1960  &  n3227 ) | ( (~ Pg35)  &  (~ Ng6682) ) | ( n3227  &  (~ Ng6682) ) ;
 assign n1956 = ( (~ Ng6741) ) | ( Ng6682 ) ;
 assign n1954 = ( (~ n1109)  &  n1957 ) | ( n1957  &  n1956 ) ;
 assign n1961 = ( Pg35 ) | ( (~ Ng6736) ) ;
 assign n1962 = ( (~ Pg35) ) | ( (~ n1109) ) | ( Ng6741 ) | ( (~ n6115) ) ;
 assign n1960 = ( (~ Pg35) ) | ( n1109 ) ;
 assign n1966 = ( (~ Pg35)  &  n1969 ) | ( n1969  &  n3277 ) | ( (~ Pg35)  &  (~ Ng6336) ) | ( n3277  &  (~ Ng6336) ) ;
 assign n1965 = ( (~ Ng6395) ) | ( Ng6336 ) ;
 assign n1963 = ( (~ n1196)  &  n1966 ) | ( n1966  &  n1965 ) ;
 assign n1970 = ( Pg35 ) | ( (~ Ng6390) ) ;
 assign n1971 = ( (~ Pg35) ) | ( (~ n1196) ) | ( Ng6395 ) | ( (~ n6116) ) ;
 assign n1969 = ( (~ Pg35) ) | ( n1196 ) ;
 assign n1975 = ( (~ Pg35)  &  n1978 ) | ( n1978  &  n3335 ) | ( (~ Pg35)  &  (~ Ng5990) ) | ( n3335  &  (~ Ng5990) ) ;
 assign n1974 = ( (~ Ng6049) ) | ( Ng5990 ) ;
 assign n1972 = ( (~ n1179)  &  n1975 ) | ( n1975  &  n1974 ) ;
 assign n1979 = ( Pg35 ) | ( (~ Ng6044) ) ;
 assign n1980 = ( (~ Pg35) ) | ( (~ n1179) ) | ( Ng6049 ) | ( (~ n6118) ) ;
 assign n1978 = ( (~ Pg35) ) | ( n1179 ) ;
 assign n1982 = ( n3849 ) | ( (~ Ng5703) ) ;
 assign n1983 = ( Ng5703 ) | ( n4784 ) | ( (~ n5777) ) ;
 assign n1987 = ( (~ Pg35)  &  n1990 ) | ( n1990  &  n3444 ) | ( (~ Pg35)  &  (~ Ng5297) ) | ( n3444  &  (~ Ng5297) ) ;
 assign n1986 = ( (~ Ng5357) ) | ( Ng5297 ) ;
 assign n1984 = ( (~ wire4394)  &  n1987 ) | ( n1987  &  n1986 ) ;
 assign n1991 = ( Pg35 ) | ( (~ Ng5352) ) ;
 assign n1992 = ( (~ Pg35) ) | ( (~ wire4394) ) | ( Ng5357 ) | ( (~ n6117) ) ;
 assign n1990 = ( (~ Pg35) ) | ( wire4394 ) ;
 assign n1994 = ( (~ Pg35) ) | ( Ng2841 ) ;
 assign n1995 = ( (~ Pg35)  &  n5781 ) | ( (~ Ng4104)  &  n5781 ) | ( (~ n1993)  &  n5781 ) ;
 assign n1993 = ( (~ Ng4108) ) | ( n2316 ) ;
 assign n1999 = ( (~ Pg35)  &  n2002 ) | ( n2002  &  n3520 ) | ( (~ Pg35)  &  (~ Ng3990) ) | ( n3520  &  (~ Ng3990) ) ;
 assign n1998 = ( (~ Ng4054) ) | ( Ng3990 ) ;
 assign n1996 = ( (~ n1165)  &  n1999 ) | ( n1999  &  n1998 ) ;
 assign n2003 = ( Pg35 ) | ( (~ Ng4049) ) ;
 assign n2004 = ( (~ Pg35) ) | ( (~ n1165) ) | ( Ng4054 ) | ( (~ n6114) ) ;
 assign n2002 = ( (~ Pg35) ) | ( n1165 ) ;
 assign n2008 = ( (~ Pg35)  &  n2011 ) | ( (~ Pg35)  &  (~ Ng3639) ) | ( n2011  &  n4792 ) | ( (~ Ng3639)  &  n4792 ) ;
 assign n2007 = ( (~ Ng3703) ) | ( Ng3639 ) ;
 assign n2005 = ( (~ n1116)  &  n2008 ) | ( n2008  &  n2007 ) ;
 assign n2012 = ( Pg35 ) | ( (~ Ng3698) ) ;
 assign n2013 = ( (~ Pg35) ) | ( (~ n1116) ) | ( Ng3703 ) | ( (~ n6119) ) ;
 assign n2011 = ( (~ Pg35) ) | ( n1116 ) ;
 assign n2017 = ( (~ Pg35)  &  n3832 ) | ( n3607  &  n3832 ) | ( (~ Pg35)  &  (~ Ng3288) ) | ( n3607  &  (~ Ng3288) ) ;
 assign n2016 = ( (~ Ng3352) ) | ( Ng3288 ) ;
 assign n2014 = ( (~ n1135)  &  n2017 ) | ( n2017  &  n2016 ) ;
 assign n2021 = ( n3832 ) | ( (~ Ng3352) ) ;
 assign n2022 = ( Ng3352 ) | ( n4793 ) | ( (~ n6120) ) ;
 assign n2024 = ( (~ Pg35)  &  n5785 ) | ( (~ Ng2759)  &  n5785 ) | ( (~ n2023)  &  n5785 ) ;
 assign n2023 = ( (~ Ng2756) ) | ( n4692 ) ;
 assign n2027 = ( (~ Pg35) ) | ( n1221 ) ;
 assign n2025 = ( (~ Pg35)  &  n2027 ) | ( n1140  &  (~ n1646)  &  n2027 ) ;
 assign n2030 = ( Pg35 ) | ( (~ Ng2555) ) ;
 assign n2033 = ( Pg35 ) | ( (~ Ng2671) ) ;
 assign n2034 = ( (~ Pg35) ) | ( n4697 ) | ( Ng2675 ) ;
 assign n2036 = ( (~ Ng2671)  &  n4697 ) | ( n4697  &  (~ n4699) ) | ( (~ Ng2671)  &  (~ n5295) ) | ( (~ n4699)  &  (~ n5295) ) ;
 assign n2038 = ( (~ n1646)  &  n4796 ) ;
 assign n2037 = ( Pg35  &  n2038 ) | ( Pg35  &  (~ n4700) ) ;
 assign n2042 = ( (~ Pg35) ) | ( n2038 ) | ( n4704 ) ;
 assign n2043 = ( Pg35 ) | ( (~ Ng2606) ) ;
 assign n2044 = ( Ng2599  &  (~ Ng2555) ) | ( (~ n4700)  &  (~ Ng2555) ) ;
 assign n2046 = ( (~ Pg35) ) | ( n2038 ) | ( n2044 ) | ( Ng2629 ) ;
 assign n2047 = ( (~ Pg35)  &  n2027 ) | ( n1093  &  (~ n1642)  &  n2027 ) ;
 assign n2051 = ( Pg35 ) | ( (~ Ng2421) ) ;
 assign n2054 = ( Pg35 ) | ( (~ Ng2537) ) ;
 assign n2055 = ( (~ Pg35) ) | ( n4707 ) | ( Ng2541 ) ;
 assign n2057 = ( (~ Ng2537)  &  n4707 ) | ( n4707  &  (~ n4709) ) | ( (~ Ng2537)  &  (~ n5299) ) | ( (~ n4709)  &  (~ n5299) ) ;
 assign n2059 = ( (~ n1642)  &  n4796 ) ;
 assign n2058 = ( Pg35  &  n2059 ) | ( Pg35  &  (~ n4710) ) ;
 assign n2063 = ( (~ Pg35) ) | ( n2059 ) | ( n4714 ) ;
 assign n2064 = ( Pg35 ) | ( (~ Ng2472) ) ;
 assign n2065 = ( Ng2465  &  (~ Ng2421) ) | ( (~ n4710)  &  (~ Ng2421) ) ;
 assign n2067 = ( (~ Pg35) ) | ( n2059 ) | ( n2065 ) | ( Ng2495 ) ;
 assign n2068 = ( (~ Pg35)  &  n2027 ) | ( n1138  &  (~ n1643)  &  n2027 ) ;
 assign n2072 = ( Pg35 ) | ( (~ Ng2287) ) ;
 assign n2075 = ( Pg35 ) | ( (~ Ng2403) ) ;
 assign n2076 = ( (~ Pg35) ) | ( n4717 ) | ( Ng2407 ) ;
 assign n2078 = ( (~ Ng2403)  &  n4717 ) | ( n4717  &  (~ n4719) ) | ( (~ Ng2403)  &  (~ n5303) ) | ( (~ n4719)  &  (~ n5303) ) ;
 assign n2080 = ( (~ n1643)  &  n4796 ) ;
 assign n2079 = ( Pg35  &  n2080 ) | ( Pg35  &  (~ n4720) ) ;
 assign n2084 = ( (~ Pg35) ) | ( n2080 ) | ( n4724 ) ;
 assign n2085 = ( Pg35 ) | ( (~ Ng2338) ) ;
 assign n2086 = ( Ng2331  &  (~ Ng2287) ) | ( (~ n4720)  &  (~ Ng2287) ) ;
 assign n2088 = ( (~ Pg35) ) | ( n2080 ) | ( n2086 ) | ( Ng2361 ) ;
 assign n2089 = ( (~ Pg35)  &  n2027 ) | ( n1096  &  (~ n1644)  &  n2027 ) ;
 assign n2093 = ( Pg35 ) | ( (~ Ng2153) ) ;
 assign n2096 = ( Pg35 ) | ( (~ Ng2269) ) ;
 assign n2097 = ( (~ Pg35) ) | ( n4727 ) | ( Ng2273 ) ;
 assign n2099 = ( (~ Ng2269)  &  n4727 ) | ( n4727  &  (~ n4729) ) | ( (~ Ng2269)  &  (~ n5307) ) | ( (~ n4729)  &  (~ n5307) ) ;
 assign n2101 = ( (~ n1644)  &  n4796 ) ;
 assign n2100 = ( Pg35  &  n2101 ) | ( Pg35  &  (~ n4730) ) ;
 assign n2105 = ( (~ Pg35) ) | ( n2101 ) | ( (~ n4730) ) | ( (~ Ng2153) ) ;
 assign n2106 = ( Pg35 ) | ( (~ Ng2204) ) ;
 assign n2107 = ( Ng2197  &  (~ Ng2153) ) | ( (~ n4730)  &  (~ Ng2153) ) ;
 assign n2109 = ( (~ Pg35) ) | ( n2101 ) | ( n2107 ) | ( Ng2227 ) ;
 assign n2110 = ( (~ Pg35)  &  n2027 ) | ( n1155  &  (~ n1640)  &  n2027 ) ;
 assign n2114 = ( Pg35 ) | ( (~ Ng1996) ) ;
 assign n2117 = ( Pg35 ) | ( (~ Ng2112) ) ;
 assign n2118 = ( (~ Pg35) ) | ( n4738 ) | ( Ng2116 ) ;
 assign n2120 = ( (~ Ng2112)  &  n4738 ) | ( n4738  &  (~ n4740) ) | ( (~ Ng2112)  &  (~ n5311) ) | ( (~ n4740)  &  (~ n5311) ) ;
 assign n2122 = ( (~ n1640)  &  n4796 ) ;
 assign n2121 = ( Pg35  &  n2122 ) | ( Pg35  &  (~ n4741) ) ;
 assign n2126 = ( (~ Pg35) ) | ( n2122 ) | ( (~ n4741) ) | ( (~ Ng1996) ) ;
 assign n2127 = ( Pg35 ) | ( (~ Ng2047) ) ;
 assign n2128 = ( Ng2040  &  (~ Ng1996) ) | ( (~ n4741)  &  (~ Ng1996) ) ;
 assign n2130 = ( (~ Pg35) ) | ( n2122 ) | ( n2128 ) | ( Ng2070 ) ;
 assign n2131 = ( (~ Pg35)  &  n2027 ) | ( n1113  &  (~ n1645)  &  n2027 ) ;
 assign n2135 = ( Pg35 ) | ( (~ Ng1862) ) ;
 assign n2138 = ( Pg35 ) | ( (~ Ng1978) ) ;
 assign n2139 = ( (~ Pg35) ) | ( n4748 ) | ( Ng1982 ) ;
 assign n2141 = ( (~ Ng1978)  &  n4748 ) | ( n4748  &  (~ n4750) ) | ( (~ Ng1978)  &  (~ n5315) ) | ( (~ n4750)  &  (~ n5315) ) ;
 assign n2143 = ( (~ n1645)  &  n4796 ) ;
 assign n2142 = ( Pg35  &  n2143 ) | ( Pg35  &  (~ n4751) ) ;
 assign n2147 = ( (~ Pg35) ) | ( n2143 ) | ( (~ n4751) ) | ( (~ Ng1862) ) ;
 assign n2148 = ( Pg35 ) | ( (~ Ng1913) ) ;
 assign n2149 = ( Ng1906  &  (~ Ng1862) ) | ( (~ n4751)  &  (~ Ng1862) ) ;
 assign n2151 = ( (~ Pg35) ) | ( n2143 ) | ( n2149 ) | ( Ng1936 ) ;
 assign n2152 = ( (~ Pg35)  &  n2027 ) | ( n1120  &  (~ n1639)  &  n2027 ) ;
 assign n2156 = ( Pg35 ) | ( (~ Ng1728) ) ;
 assign n2159 = ( Pg35 ) | ( (~ Ng1844) ) ;
 assign n2160 = ( (~ Pg35) ) | ( n4758 ) | ( Ng1848 ) ;
 assign n2162 = ( (~ Ng1844)  &  n4758 ) | ( n4758  &  (~ n4760) ) | ( (~ Ng1844)  &  (~ n5319) ) | ( (~ n4760)  &  (~ n5319) ) ;
 assign n2164 = ( (~ n1639)  &  n4796 ) ;
 assign n2163 = ( Pg35  &  n2164 ) | ( Pg35  &  (~ n4761) ) ;
 assign n2168 = ( (~ Pg35) ) | ( n2164 ) | ( n4765 ) ;
 assign n2169 = ( Pg35 ) | ( (~ Ng1779) ) ;
 assign n2170 = ( Ng1772  &  (~ Ng1728) ) | ( (~ n4761)  &  (~ Ng1728) ) ;
 assign n2172 = ( (~ Pg35) ) | ( n2164 ) | ( n2170 ) | ( Ng1802 ) ;
 assign n2173 = ( (~ Pg35)  &  n2027 ) | ( wire4406  &  (~ n1641)  &  n2027 ) ;
 assign n2177 = ( Pg35 ) | ( (~ Ng1592) ) ;
 assign n2180 = ( Pg35 ) | ( (~ Ng1710) ) ;
 assign n2181 = ( (~ Pg35) ) | ( n4768 ) | ( Ng1714 ) ;
 assign n2183 = ( (~ Ng1710)  &  n4768 ) | ( n4768  &  (~ n4770) ) | ( (~ Ng1710)  &  (~ n5323) ) | ( (~ n4770)  &  (~ n5323) ) ;
 assign n2185 = ( n1923  &  n4773 ) | ( (~ Ng1668)  &  n4773 ) | ( n1923  &  n5588 ) | ( (~ Ng1668)  &  n5588 ) ;
 assign n2186 = ( (~ Pg35) ) | ( n4774 ) | ( n5588 ) ;
 assign n2187 = ( Pg35 ) | ( (~ Ng1644) ) ;
 assign n2188 = ( Ng1636  &  (~ Ng1592) ) | ( (~ Ng1592)  &  (~ n4771) ) ;
 assign n2191 = ( (~ Pg35) ) | ( n2188 ) | ( Ng1668 ) | ( n5588 ) ;
 assign n2194 = ( Ng1333 ) | ( Ng1322 ) ;
 assign n2192 = ( n2194  &  Ng1345 ) | ( n2194  &  (~ n4805) ) ;
 assign n2195 = ( n2192  &  Ng1361 ) | ( n2192  &  (~ n4805) ) ;
 assign n2196 = ( n2195  &  Ng1367 ) | ( n2195  &  (~ n4805) ) ;
 assign n2197 = ( Pg35  &  (~ n2196) ) | ( Pg35  &  Ng1379 ) | ( Pg35  &  (~ n4805) ) ;
 assign n2203 = ( (~ Ng1274) ) | ( n666 ) | ( n4222 ) ;
 assign n2204 = ( Pg35 ) | ( (~ Ng1270) ) ;
 assign n2207 = ( Ng990 ) | ( Ng979 ) ;
 assign n2205 = ( n2207  &  Ng1002 ) | ( n2207  &  (~ n4818) ) ;
 assign n2208 = ( n2205  &  Ng1018 ) | ( n2205  &  (~ n4818) ) ;
 assign n2209 = ( n2208  &  Ng1024 ) | ( n2208  &  (~ n4818) ) ;
 assign n2210 = ( Pg35  &  (~ n2209) ) | ( Pg35  &  Ng1036 ) | ( Pg35  &  (~ n4818) ) ;
 assign n2216 = ( (~ Ng930) ) | ( n670 ) | ( n4235 ) ;
 assign n2217 = ( Pg35 ) | ( (~ Ng925) ) ;
 assign n2219 = ( (~ Ng763) ) | ( (~ n2218) ) | ( n3791 ) ;
 assign n2220 = ( Pg35 ) | ( (~ Ng758) ) ;
 assign n2218 = ( (~ Ng758) ) | ( n2477 ) ;
 assign n2223 = ( Pg35 ) | ( (~ Ng590) ) ;
 assign n2221 = ( (~ Ng590) ) | ( n2480 ) ;
 assign n2225 = ( Ng294 ) | ( n4661 ) ;
 assign n2226 = ( n3904 ) | ( (~ Ng294) ) | ( (~ n4661) ) ;
 assign n2228 = ( Ng153 ) | ( n4670 ) ;
 assign n2229 = ( n3182 ) | ( (~ Ng153) ) | ( (~ n4670) ) ;
 assign n2232 = ( (~ Ng6561) ) | ( n4833 ) ;
 assign n2230 = ( n2232  &  (~ Ng25756) ) | ( n2232  &  Ng6561  &  Ng6565 ) ;
 assign n2233 = ( n4110  &  n4832 ) ;
 assign n2235 = ( Pg35  &  Ng6565 ) | ( Pg35  &  n2233 ) ;
 assign n2237 = ( (~ Pg35) ) | ( Ng6561 ) | ( n2233 ) ;
 assign n2238 = ( (~ Ng6555) ) | ( (~ Ng6549) ) ;
 assign n2242 = ( Ng6555 ) | ( (~ Ng6549) ) ;
 assign n2241 = ( (~ Ng6555) ) | ( Ng6549 ) ;
 assign n2240 = ( (~ Pg35)  &  n2242 ) | ( n2242  &  n2241 ) ;
 assign n2245 = ( (~ Ng6215) ) | ( n4836 ) ;
 assign n2244 = ( (~ Pg35) ) | ( (~ Ng6227) ) ;
 assign n2243 = ( n2245  &  n2244 ) | ( n2245  &  Ng6215  &  Ng6219 ) ;
 assign n2246 = ( n4582  &  n4835 ) ;
 assign n2248 = ( Pg35  &  Ng6219 ) | ( Pg35  &  n2246 ) ;
 assign n2250 = ( (~ Pg35) ) | ( Ng6215 ) | ( n2246 ) ;
 assign n2251 = ( (~ Ng6203) ) | ( (~ Ng6209) ) ;
 assign n2255 = ( (~ Ng6203) ) | ( Ng6209 ) ;
 assign n2254 = ( Ng6203 ) | ( (~ Ng6209) ) ;
 assign n2253 = ( (~ Pg35)  &  n2255 ) | ( n2255  &  n2254 ) ;
 assign n2258 = ( (~ Ng5869) ) | ( n4837 ) ;
 assign n2256 = ( n2258  &  (~ Ng25728) ) | ( n2258  &  Ng5869  &  Ng5873 ) ;
 assign n2259 = ( n4582  &  n4832 ) ;
 assign n2261 = ( Pg35  &  Ng5873 ) | ( Pg35  &  n2259 ) ;
 assign n2263 = ( (~ Pg35) ) | ( Ng5869 ) | ( n2259 ) ;
 assign n2264 = ( (~ Ng5863) ) | ( (~ Ng5857) ) ;
 assign n2268 = ( Ng5863 ) | ( (~ Ng5857) ) ;
 assign n2267 = ( (~ Ng5863) ) | ( Ng5857 ) ;
 assign n2266 = ( (~ Pg35)  &  n2268 ) | ( n2268  &  n2267 ) ;
 assign n2271 = ( (~ Ng5523) ) | ( n4838 ) ;
 assign n2270 = ( (~ Pg35) ) | ( (~ Ng5535) ) ;
 assign n2269 = ( n2271  &  n2270 ) | ( n2271  &  Ng5523  &  Ng5527 ) ;
 assign n2272 = ( (~ n1633)  &  n4835 ) ;
 assign n2274 = ( Pg35  &  Ng5527 ) | ( Pg35  &  n2272 ) ;
 assign n2276 = ( (~ Pg35) ) | ( Ng5523 ) | ( n2272 ) ;
 assign n2277 = ( (~ Ng5517) ) | ( (~ Ng5511) ) ;
 assign n2281 = ( Ng5517 ) | ( (~ Ng5511) ) ;
 assign n2280 = ( (~ Ng5517) ) | ( Ng5511 ) ;
 assign n2279 = ( (~ Pg35)  &  n2281 ) | ( n2281  &  n2280 ) ;
 assign n2284 = ( (~ Ng5176) ) | ( n4839 ) ;
 assign n2283 = ( (~ Pg35) ) | ( (~ Ng5188) ) ;
 assign n2282 = ( n2284  &  n2283 ) | ( n2284  &  Ng5176  &  Ng5180 ) ;
 assign n2285 = ( (~ n1633)  &  n4832 ) ;
 assign n2287 = ( Pg35  &  Ng5180 ) | ( Pg35  &  n2285 ) ;
 assign n2289 = ( (~ Pg35) ) | ( Ng5176 ) | ( n2285 ) ;
 assign n2290 = ( (~ Ng5170) ) | ( (~ Ng5164) ) ;
 assign n2294 = ( Ng5170 ) | ( (~ Ng5164) ) ;
 assign n2293 = ( (~ Ng5170) ) | ( Ng5164 ) ;
 assign n2292 = ( (~ Pg35)  &  n2294 ) | ( n2294  &  n2293 ) ;
 assign n2296 = ( (~ Pg35) ) | ( Ng5057 ) | ( n5795 ) ;
 assign n2297 = ( n2509 ) | ( (~ Ng5057) ) | ( (~ n5795) ) ;
 assign n2302 = ( (~ n1222)  &  (~ n2521) ) | ( (~ n1222)  &  (~ Ng4549) ) | ( n2521  &  (~ Ng4549) ) ;
 assign n2301 = ( (~ n1253)  &  n2302 ) ;
 assign n2304 = ( n2521 ) | ( (~ Ng4575) ) ;
 assign n2309 = ( (~ n1222)  &  (~ n2521) ) | ( (~ n1222)  &  (~ Ng4504) ) | ( n2521  &  (~ Ng4504) ) ;
 assign n2310 = ( n2521 ) | ( (~ Ng4572) ) ;
 assign n2308 = ( n2309  &  n2310 ) ;
 assign n2312 = ( (~ wire4437) ) | ( n2521 ) ;
 assign n2317 = ( (~ Pg35)  &  n5799 ) | ( (~ Ng4108)  &  n5799 ) | ( (~ n2316)  &  n5799 ) ;
 assign n2316 = ( (~ Ng4098) ) | ( n4791 ) ;
 assign n2320 = ( (~ Ng3869) ) | ( n4855 ) ;
 assign n2319 = ( (~ Pg35) ) | ( (~ Ng3881) ) ;
 assign n2318 = ( n2320  &  n2319 ) | ( n2320  &  Ng3869  &  Ng3873 ) ;
 assign n2321 = ( n4585  &  n4835 ) ;
 assign n2323 = ( Pg35  &  Ng3873 ) | ( Pg35  &  n2321 ) ;
 assign n2325 = ( (~ Pg35) ) | ( Ng3869 ) | ( n2321 ) ;
 assign n2326 = ( (~ Ng3857) ) | ( (~ Ng3863) ) ;
 assign n2330 = ( (~ Ng3857) ) | ( Ng3863 ) ;
 assign n2329 = ( Ng3857 ) | ( (~ Ng3863) ) ;
 assign n2328 = ( (~ Pg35)  &  n2330 ) | ( n2330  &  n2329 ) ;
 assign n2333 = ( (~ Ng3518) ) | ( n4856 ) ;
 assign n2332 = ( (~ Pg35) ) | ( (~ Ng3530) ) ;
 assign n2331 = ( n2333  &  n2332 ) | ( n2333  &  Ng3518  &  Ng3522 ) ;
 assign n2334 = ( n4585  &  n4832 ) ;
 assign n2336 = ( Pg35  &  Ng3522 ) | ( Pg35  &  n2334 ) ;
 assign n2338 = ( (~ Pg35) ) | ( Ng3518 ) | ( n2334 ) ;
 assign n2339 = ( (~ Ng3512) ) | ( (~ Ng3506) ) ;
 assign n2343 = ( Ng3512 ) | ( (~ Ng3506) ) ;
 assign n2342 = ( (~ Ng3512) ) | ( Ng3506 ) ;
 assign n2341 = ( (~ Pg35)  &  n2343 ) | ( n2343  &  n2342 ) ;
 assign n2346 = ( (~ Ng3167) ) | ( n4857 ) ;
 assign n2345 = ( (~ Pg35) ) | ( (~ Ng3179) ) ;
 assign n2344 = ( n2346  &  n2345 ) | ( n2346  &  Ng3167  &  Ng3171 ) ;
 assign n2347 = ( n4110  &  n4835 ) ;
 assign n2349 = ( Pg35  &  Ng3171 ) | ( Pg35  &  n2347 ) ;
 assign n2351 = ( (~ Pg35) ) | ( Ng3167 ) | ( n2347 ) ;
 assign n2352 = ( (~ Ng3161) ) | ( (~ Ng3155) ) ;
 assign n2356 = ( Ng3161 ) | ( (~ Ng3155) ) ;
 assign n2355 = ( (~ Ng3161) ) | ( Ng3155 ) ;
 assign n2354 = ( (~ Pg35)  &  n2356 ) | ( n2356  &  n2355 ) ;
 assign n2358 = ( Pg35 ) | ( (~ Ng2748) ) ;
 assign n2357 = ( (~ n4692)  &  Ng2756 ) | ( n4692  &  (~ Ng2756) ) ;
 assign n2361 = ( (~ Pg35) ) | ( n1153 ) ;
 assign n2359 = ( (~ Pg35)  &  n2027  &  n2361 ) | ( (~ n1698)  &  n2027  &  n2361 ) ;
 assign n2363 = ( (~ n1153) ) | ( n1698 ) | ( n4324 ) | ( (~ n4794) ) ;
 assign n2364 = ( Pg35 ) | ( (~ Ng2610) ) ;
 assign n2366 = ( n1698 ) | ( (~ n4859) ) | ( n4860 ) ;
 assign n2367 = ( Pg35  &  (~ Ng2610) ) | ( (~ Ng2625)  &  (~ Ng2610) ) | ( Pg35  &  n4860 ) | ( (~ Ng2625)  &  n4860 ) ;
 assign n2369 = ( (~ n2361)  &  (~ Ng2610) ) | ( n2361  &  (~ Ng2587) ) | ( (~ Ng2610)  &  (~ Ng2587) ) ;
 assign n2368 = ( n2369  &  n2366 ) ;
 assign n2370 = ( Ng2619 ) | ( n4860 ) | ( (~ n4947) ) ;
 assign n2371 = ( Pg35  &  n2361 ) | ( Pg35  &  (~ Ng2587) ) | ( n2361  &  (~ Ng2595) ) | ( (~ Ng2587)  &  (~ Ng2595) ) ;
 assign n2374 = ( (~ Pg35) ) | ( n1151 ) ;
 assign n2372 = ( (~ Pg35)  &  n2027  &  n2374 ) | ( (~ n1695)  &  n2027  &  n2374 ) ;
 assign n2376 = ( (~ n1151) ) | ( n1695 ) | ( n4326 ) | ( (~ n4794) ) ;
 assign n2377 = ( Pg35 ) | ( (~ Ng2476) ) ;
 assign n2379 = ( n1695 ) | ( (~ n4859) ) | ( n4864 ) ;
 assign n2380 = ( Pg35  &  (~ Ng2476) ) | ( (~ Ng2491)  &  (~ Ng2476) ) | ( Pg35  &  n4864 ) | ( (~ Ng2491)  &  n4864 ) ;
 assign n2382 = ( (~ n2374)  &  (~ Ng2476) ) | ( n2374  &  (~ Ng2453) ) | ( (~ Ng2476)  &  (~ Ng2453) ) ;
 assign n2381 = ( n2382  &  n2379 ) ;
 assign n2384 = ( (~ Pg35) ) | ( (~ Ng2453) ) | ( n4948 ) ;
 assign n2385 = ( n2379  &  Ng2485 ) | ( n2379  &  Ng2476 ) | ( n2379  &  n4864 ) ;
 assign n2388 = ( (~ Pg35) ) | ( n1162 ) ;
 assign n2386 = ( (~ Pg35)  &  n2027  &  n2388 ) | ( (~ n1697)  &  n2027  &  n2388 ) ;
 assign n2390 = ( (~ n1162) ) | ( n1697 ) | ( n4328 ) | ( (~ n4794) ) ;
 assign n2391 = ( Pg35 ) | ( (~ Ng2342) ) ;
 assign n2393 = ( n1697 ) | ( (~ n4859) ) | ( n4866 ) ;
 assign n2394 = ( Pg35  &  (~ Ng2342) ) | ( (~ Ng2357)  &  (~ Ng2342) ) | ( Pg35  &  n4866 ) | ( (~ Ng2357)  &  n4866 ) ;
 assign n2396 = ( (~ n2388)  &  (~ Ng2342) ) | ( n2388  &  (~ Ng2319) ) | ( (~ Ng2342)  &  (~ Ng2319) ) ;
 assign n2395 = ( n2396  &  n2393 ) ;
 assign n2397 = ( Ng2351 ) | ( n4866 ) | ( (~ n4954) ) ;
 assign n2398 = ( Pg35  &  n2388 ) | ( Pg35  &  (~ Ng2319) ) | ( n2388  &  (~ Ng2327) ) | ( (~ Ng2319)  &  (~ Ng2327) ) ;
 assign n2401 = ( (~ Pg35) ) | ( n1104 ) ;
 assign n2399 = ( (~ Pg35)  &  n2027  &  n2401 ) | ( (~ n1699)  &  n2027  &  n2401 ) ;
 assign n2403 = ( (~ n1104) ) | ( n1699 ) | ( n4330 ) | ( (~ n4794) ) ;
 assign n2404 = ( Pg35 ) | ( (~ Ng2208) ) ;
 assign n2406 = ( n1699 ) | ( (~ n4859) ) | ( n4870 ) ;
 assign n2407 = ( Pg35  &  (~ Ng2208) ) | ( (~ Ng2223)  &  (~ Ng2208) ) | ( Pg35  &  n4870 ) | ( (~ Ng2223)  &  n4870 ) ;
 assign n2409 = ( (~ n2401)  &  (~ Ng2208) ) | ( n2401  &  (~ Ng2185) ) | ( (~ Ng2208)  &  (~ Ng2185) ) ;
 assign n2408 = ( n2409  &  n2406 ) ;
 assign n2410 = ( Ng2217 ) | ( n4870 ) | ( (~ n4957) ) ;
 assign n2411 = ( Pg35  &  n2401 ) | ( Pg35  &  (~ Ng2185) ) | ( n2401  &  (~ Ng2193) ) | ( (~ Ng2185)  &  (~ Ng2193) ) ;
 assign n2414 = ( (~ Pg35) ) | ( n1146 ) ;
 assign n2412 = ( (~ Pg35)  &  n2027  &  n2414 ) | ( (~ n1701)  &  n2027  &  n2414 ) ;
 assign n2416 = ( (~ n1146) ) | ( n1701 ) | ( n4332 ) | ( (~ n4794) ) ;
 assign n2417 = ( Pg35 ) | ( (~ Ng2051) ) ;
 assign n2419 = ( n1701 ) | ( (~ n4859) ) | ( n4873 ) ;
 assign n2420 = ( Pg35  &  (~ Ng2051) ) | ( (~ Ng2066)  &  (~ Ng2051) ) | ( Pg35  &  n4873 ) | ( (~ Ng2066)  &  n4873 ) ;
 assign n2422 = ( (~ n2414)  &  (~ Ng2051) ) | ( n2414  &  (~ Ng2028) ) | ( (~ Ng2051)  &  (~ Ng2028) ) ;
 assign n2421 = ( n2422  &  n2419 ) ;
 assign n2424 = ( (~ Pg35) ) | ( (~ Ng2028) ) | ( n4958 ) ;
 assign n2425 = ( n2419  &  Ng2051 ) | ( n2419  &  Ng2060 ) | ( n2419  &  n4873 ) ;
 assign n2428 = ( (~ Pg35) ) | ( n1126 ) ;
 assign n2426 = ( (~ Pg35)  &  n2027  &  n2428 ) | ( (~ n1700)  &  n2027  &  n2428 ) ;
 assign n2430 = ( (~ n1126) ) | ( n1700 ) | ( n4334 ) | ( (~ n4794) ) ;
 assign n2431 = ( Pg35 ) | ( (~ Ng1917) ) ;
 assign n2433 = ( n1700 ) | ( (~ n4859) ) | ( n4875 ) ;
 assign n2434 = ( Pg35  &  (~ Ng1917) ) | ( (~ Ng1932)  &  (~ Ng1917) ) | ( Pg35  &  n4875 ) | ( (~ Ng1932)  &  n4875 ) ;
 assign n2436 = ( (~ n2428)  &  (~ Ng1917) ) | ( n2428  &  (~ Ng1894) ) | ( (~ Ng1917)  &  (~ Ng1894) ) ;
 assign n2435 = ( n2436  &  n2433 ) ;
 assign n2437 = ( Ng1926 ) | ( n4875 ) | ( (~ n4964) ) ;
 assign n2438 = ( Pg35  &  n2428 ) | ( Pg35  &  (~ Ng1894) ) | ( n2428  &  (~ Ng1902) ) | ( (~ Ng1894)  &  (~ Ng1902) ) ;
 assign n2441 = ( (~ Pg35) ) | ( n1182 ) ;
 assign n2439 = ( (~ Pg35)  &  n2027  &  n2441 ) | ( (~ n1696)  &  n2027  &  n2441 ) ;
 assign n2443 = ( (~ n1182) ) | ( n1696 ) | ( n4336 ) | ( (~ n4794) ) ;
 assign n2444 = ( Pg35 ) | ( (~ Ng1783) ) ;
 assign n2446 = ( n1696 ) | ( (~ n4859) ) | ( n4878 ) ;
 assign n2447 = ( Pg35  &  (~ Ng1783) ) | ( (~ Ng1798)  &  (~ Ng1783) ) | ( Pg35  &  n4878 ) | ( (~ Ng1798)  &  n4878 ) ;
 assign n2449 = ( (~ n2441)  &  (~ Ng1783) ) | ( n2441  &  (~ Ng1760) ) | ( (~ Ng1783)  &  (~ Ng1760) ) ;
 assign n2448 = ( n2449  &  n2446 ) ;
 assign n2450 = ( Ng1792 ) | ( n4878 ) | ( (~ n4967) ) ;
 assign n2451 = ( Pg35  &  n2441 ) | ( Pg35  &  (~ Ng1760) ) | ( n2441  &  (~ Ng1768) ) | ( (~ Ng1760)  &  (~ Ng1768) ) ;
 assign n2454 = ( (~ Pg35) ) | ( n1087 ) ;
 assign n2452 = ( (~ Pg35)  &  n2027  &  n2454 ) | ( (~ n1702)  &  n2027  &  n2454 ) ;
 assign n2456 = ( (~ n1087) ) | ( n1702 ) | ( n4338 ) | ( (~ n4794) ) ;
 assign n2457 = ( Pg35 ) | ( (~ Ng1648) ) ;
 assign n2459 = ( n1702 ) | ( (~ n4859) ) | ( n4881 ) ;
 assign n2460 = ( Pg35  &  (~ Ng1648) ) | ( (~ Ng1664)  &  (~ Ng1648) ) | ( Pg35  &  n4881 ) | ( (~ Ng1664)  &  n4881 ) ;
 assign n2462 = ( (~ n2454)  &  (~ Ng1648) ) | ( n2454  &  (~ Ng1624) ) | ( (~ Ng1648)  &  (~ Ng1624) ) ;
 assign n2461 = ( n2462  &  n2459 ) ;
 assign n2463 = ( Ng1657 ) | ( n4881 ) | ( (~ n4970) ) ;
 assign n2464 = ( Pg35  &  n2454 ) | ( Pg35  &  (~ Ng1624) ) | ( n2454  &  (~ Ng1632) ) | ( (~ Ng1624)  &  (~ Ng1632) ) ;
 assign n2466 = ( (~ Pg35) ) | ( n2196 ) | ( (~ Ng1373) ) ;
 assign n2467 = ( (~ n2196) ) | ( n3875 ) | ( Ng1373 ) ;
 assign n2469 = ( (~ Ng1270) ) | ( (~ n2468) ) | ( n4222 ) ;
 assign n2470 = ( Pg35 ) | ( (~ Ng1263) ) ;
 assign n2468 = ( (~ Ng1263) ) | ( (~ n4813) ) ;
 assign n2472 = ( (~ Pg35) ) | ( n2209 ) | ( (~ Ng1030) ) ;
 assign n2473 = ( (~ n2209) ) | ( n3881 ) | ( Ng1030 ) ;
 assign n2475 = ( (~ Ng925) ) | ( (~ n2474) ) | ( n4235 ) ;
 assign n2476 = ( Pg35 ) | ( (~ Ng918) ) ;
 assign n2474 = ( (~ Ng918) ) | ( (~ n4826) ) ;
 assign n2478 = ( (~ Ng758) ) | ( (~ n2477) ) | ( n3791 ) ;
 assign n2479 = ( Pg35 ) | ( (~ Ng749) ) ;
 assign n2477 = ( (~ Ng749) ) | ( n2546 ) ;
 assign n2482 = ( Pg35 ) | ( (~ Ng582) ) ;
 assign n2480 = ( (~ Ng582) ) | ( n2549 ) ;
 assign n2484 = ( (~ n4660) ) | ( Ng291 ) ;
 assign n2485 = ( n3904 ) | ( n4660 ) | ( (~ Ng291) ) ;
 assign n2487 = ( (~ n4669) ) | ( Ng150 ) ;
 assign n2488 = ( n3182 ) | ( n4669 ) | ( (~ Ng150) ) ;
 assign n2489 = ( (~ Ng2950)  &  (~ Ng2927) ) | ( (~ Ng2955)  &  (~ Ng2927) ) | ( (~ Ng2950)  &  (~ Ng2922) ) | ( (~ Ng2955)  &  (~ Ng2922) ) ;
 assign n2490 = ( (~ Ng2936) ) | ( (~ Ng2941) ) ;
 assign n2491 = ( (~ Ng2975)  &  (~ Ng2902) ) | ( (~ Ng2970)  &  (~ Ng2902) ) | ( (~ Ng2975)  &  (~ Ng2907) ) | ( (~ Ng2970)  &  (~ Ng2907) ) ;
 assign n2492 = ( (~ Ng2965)  &  (~ Ng2917) ) | ( (~ Ng2960)  &  (~ Ng2917) ) | ( (~ Ng2965)  &  (~ Ng2912) ) | ( (~ Ng2960)  &  (~ Ng2912) ) ;
 assign n2498 = ( n2509 ) | ( (~ n4840) ) | ( (~ Ng5033) ) | ( (~ n4844) ) ;
 assign n2501 = ( n2509 ) | ( (~ Ng5052) ) | ( (~ n4846) ) | ( (~ n5794) ) ;
 assign n2505 = ( (~ Ng5029) ) | ( Ng5062 ) | ( n4850 ) ;
 assign n2503 = ( Pg35  &  n2505  &  Ng5029 ) | ( Pg35  &  n2505  &  (~ Ng5062) ) ;
 assign n2507 = ( (~ Ng5029) ) | ( n2509 ) | ( Ng5016 ) | ( Ng5022 ) ;
 assign n2508 = ( (~ Pg35) ) | ( n4844 ) ;
 assign n2511 = ( (~ Pg35)  &  n5815 ) | ( Ng5046  &  n5815 ) | ( n5327  &  n5815 ) ;
 assign n2509 = ( (~ Pg35) ) | ( n4850 ) ;
 assign n2514 = ( (~ Pg35)  &  n5816 ) | ( Ng5041  &  n5816 ) | ( n4883  &  n5816 ) ;
 assign n2517 = ( (~ Pg35)  &  n5817 ) | ( Ng5037  &  n5817 ) | ( n5328  &  n5817 ) ;
 assign n2519 = ( (~ Pg35)  &  n5818 ) | ( (~ Ng5016)  &  n5818 ) | ( n4884  &  n5818 ) ;
 assign n2522 = ( (~ Pg35) ) | ( Ng4581 ) | ( (~ Ng4372) ) ;
 assign n2521 = ( (~ Pg35) ) | ( (~ Ng4581) ) ;
 assign n2520 = ( n2522  &  n2521 ) | ( n2522  &  Pg72  &  Pg73 ) ;
 assign n2527 = ( Pg35 ) | ( (~ Ng4093) ) ;
 assign n2526 = ( (~ n4791)  &  Ng4098 ) | ( n4791  &  (~ Ng4098) ) ;
 assign n2532 = ( (~ Ng2748) ) | ( n3046 ) | ( (~ n4691) ) ;
 assign n2533 = ( Ng2748 ) | ( n4691 ) | ( (~ Ng2841) ) ;
 assign n2535 = ( (~ Pg35) ) | ( n2195 ) | ( (~ Ng1367) ) ;
 assign n2536 = ( (~ n2195) ) | ( Ng1367 ) | ( n3875 ) ;
 assign n2538 = ( (~ Ng1263) ) | ( n4222 ) | ( n4813 ) ;
 assign n2539 = ( Pg35 ) | ( (~ Ng1259) ) ;
 assign n2541 = ( (~ Pg35) ) | ( n2208 ) | ( (~ Ng1024) ) ;
 assign n2542 = ( (~ n2208) ) | ( Ng1024 ) | ( n3881 ) ;
 assign n2544 = ( (~ Ng918) ) | ( n4235 ) | ( n4826 ) ;
 assign n2545 = ( Pg35 ) | ( (~ Ng914) ) ;
 assign n2547 = ( (~ Ng749) ) | ( (~ n2546) ) | ( n3791 ) ;
 assign n2548 = ( Pg35 ) | ( (~ Ng744) ) ;
 assign n2546 = ( (~ Ng744) ) | ( n3175 ) ;
 assign n2550 = ( (~ Ng582) ) | ( (~ n2549) ) | ( n4508 ) ;
 assign n2551 = ( Pg35 ) | ( (~ Ng577) ) ;
 assign n2549 = ( (~ Ng577) ) | ( n3178 ) ;
 assign n2553 = ( Ng164 ) | ( (~ n4667) ) ;
 assign n2554 = ( n3182 ) | ( (~ Ng164) ) | ( n4667 ) ;
 assign n2555 = ( (~ n1107)  &  (~ n4569) ) | ( (~ n4345)  &  (~ n4569) ) ;
 assign n2563 = ( n2560 ) | ( n2561 ) ;
 assign n2562 = ( Pg35  &  Ng5817 ) ;
 assign n2560 = ( Pg35  &  Ng5124 ) ;
 assign n2561 = ( Pg35  &  Ng6163 ) ;
 assign n2559 = ( n2563  &  n2562 ) | ( n2563  &  n2560  &  n2561 ) ;
 assign n2567 = ( n4340 ) | ( n4342 ) | ( n4344 ) | ( n4569 ) | ( n4345 ) | ( n1107 ) ;
 assign n2564 = ( Pg35  &  Ng3817 ) ;
 assign n2565 = ( Pg35  &  Ng3115 ) ;
 assign n2569 = ( n160  &  (~ n4886) ) | ( n3184  &  (~ n4886) ) | ( n160  &  (~ Ng6657) ) | ( n3184  &  (~ Ng6657) ) ;
 assign n2572 = ( Pg35 ) | ( (~ Ng6649) ) ;
 assign n2573 = ( (~ Pg35) ) | ( (~ n2571) ) | ( (~ Ng6605) ) ;
 assign n2571 = ( (~ Ng6561) ) | ( n4888 ) ;
 assign n2574 = ( Pg35 ) | ( (~ Ng6645) ) ;
 assign n2577 = ( Pg35 ) | ( (~ Ng6641) ) ;
 assign n2578 = ( (~ Pg35) ) | ( (~ n2576) ) | ( (~ Ng6589) ) ;
 assign n2576 = ( (~ Ng6561) ) | ( n4889 ) ;
 assign n2580 = ( Pg35 ) | ( (~ Ng6637) ) ;
 assign n2579 = ( n4588 ) | ( n2238 ) ;
 assign n2583 = ( Pg35 ) | ( (~ Ng6633) ) ;
 assign n2584 = ( (~ Pg35) ) | ( (~ n2582) ) | ( (~ Ng6649) ) ;
 assign n2582 = ( n2238 ) | ( n4888 ) ;
 assign n2586 = ( Pg35 ) | ( (~ Ng6629) ) ;
 assign n2587 = ( (~ Pg35) ) | ( (~ n2585) ) | ( (~ Ng6645) ) ;
 assign n2585 = ( n4833 ) | ( n2238 ) ;
 assign n2589 = ( Pg35 ) | ( (~ Ng6625) ) ;
 assign n2590 = ( (~ Pg35) ) | ( (~ n2588) ) | ( (~ Ng6641) ) ;
 assign n2588 = ( n2238 ) | ( n4889 ) ;
 assign n2592 = ( Pg35 ) | ( (~ Ng6621) ) ;
 assign n2593 = ( (~ Pg35) ) | ( (~ n2591) ) | ( (~ Ng6637) ) ;
 assign n2591 = ( n4588 ) | ( n2241 ) ;
 assign n2595 = ( Pg35 ) | ( (~ Ng6617) ) ;
 assign n2594 = ( n2241 ) | ( n4888 ) ;
 assign n2598 = ( Pg35 ) | ( (~ Ng6613) ) ;
 assign n2599 = ( (~ Pg35) ) | ( (~ n2597) ) | ( (~ Ng6629) ) ;
 assign n2597 = ( n4833 ) | ( n2241 ) ;
 assign n2601 = ( Pg35 ) | ( (~ Ng6609) ) ;
 assign n2602 = ( (~ Pg35) ) | ( (~ n2600) ) | ( (~ Ng6625) ) ;
 assign n2600 = ( n2241 ) | ( n4889 ) ;
 assign n2604 = ( Pg35 ) | ( (~ Ng6601) ) ;
 assign n2605 = ( (~ Pg35) ) | ( (~ n2603) ) | ( (~ Ng6621) ) ;
 assign n2603 = ( n4588 ) | ( n2242 ) ;
 assign n2607 = ( Pg35 ) | ( (~ Ng6593) ) ;
 assign n2608 = ( (~ Pg35) ) | ( (~ n2606) ) | ( (~ Ng6617) ) ;
 assign n2606 = ( n4888 ) | ( n2242 ) ;
 assign n2610 = ( Pg35 ) | ( (~ Ng6585) ) ;
 assign n2611 = ( (~ Pg35) ) | ( (~ n2609) ) | ( (~ Ng6613) ) ;
 assign n2609 = ( n4833 ) | ( n2242 ) ;
 assign n2613 = ( Pg35 ) | ( (~ Ng6581) ) ;
 assign n2614 = ( (~ Pg35) ) | ( (~ n2612) ) | ( (~ Ng6609) ) ;
 assign n2612 = ( n4889 ) | ( n2242 ) ;
 assign n2616 = ( Pg35 ) | ( (~ Ng6605) ) ;
 assign n2617 = ( (~ Pg35) ) | ( (~ n2615) ) | ( (~ Ng6601) ) ;
 assign n2615 = ( n4588 ) | ( n4893 ) ;
 assign n2619 = ( Pg35 ) | ( (~ Ng6597) ) ;
 assign n2620 = ( (~ Pg35) ) | ( (~ n2618) ) | ( (~ Ng6593) ) ;
 assign n2618 = ( n4888 ) | ( n4893 ) ;
 assign n2622 = ( Pg35 ) | ( (~ Ng6589) ) ;
 assign n2623 = ( (~ Pg35) ) | ( (~ n2621) ) | ( (~ Ng6585) ) ;
 assign n2621 = ( n4833 ) | ( n4893 ) ;
 assign n2625 = ( Pg35 ) | ( (~ Ng6573) ) ;
 assign n2626 = ( (~ Pg35) ) | ( (~ n2624) ) | ( (~ Ng6581) ) ;
 assign n2624 = ( n4889 ) | ( n4893 ) ;
 assign n2628 = ( n160  &  (~ n4894) ) | ( n3238  &  (~ n4894) ) | ( n160  &  (~ Ng6311) ) | ( n3238  &  (~ Ng6311) ) ;
 assign n2630 = ( Pg35 ) | ( (~ Ng6303) ) ;
 assign n2631 = ( (~ Pg35) ) | ( (~ n2629) ) | ( (~ Ng6259) ) ;
 assign n2629 = ( (~ Ng6215) ) | ( n4895 ) ;
 assign n2632 = ( Pg35 ) | ( (~ Ng6299) ) ;
 assign n2633 = ( (~ Pg35) ) | ( (~ n2245) ) | ( (~ Ng6251) ) ;
 assign n2635 = ( Pg35 ) | ( (~ Ng6295) ) ;
 assign n2636 = ( (~ Pg35) ) | ( (~ n2634) ) | ( (~ Ng6243) ) ;
 assign n2634 = ( (~ Ng6215) ) | ( n4896 ) ;
 assign n2638 = ( Pg35 ) | ( (~ Ng6291) ) ;
 assign n2639 = ( (~ Pg35) ) | ( (~ n2637) ) | ( (~ Ng6307) ) ;
 assign n2637 = ( n4581 ) | ( n2251 ) ;
 assign n2641 = ( Pg35 ) | ( (~ Ng6287) ) ;
 assign n2642 = ( (~ Pg35) ) | ( (~ n2640) ) | ( (~ Ng6303) ) ;
 assign n2640 = ( n2251 ) | ( n4895 ) ;
 assign n2644 = ( Pg35 ) | ( (~ Ng6283) ) ;
 assign n2645 = ( (~ Pg35) ) | ( (~ n2643) ) | ( (~ Ng6299) ) ;
 assign n2643 = ( n4836 ) | ( n2251 ) ;
 assign n2647 = ( Pg35 ) | ( (~ Ng6279) ) ;
 assign n2648 = ( (~ Pg35) ) | ( (~ n2646) ) | ( (~ Ng6295) ) ;
 assign n2646 = ( n2251 ) | ( n4896 ) ;
 assign n2650 = ( Pg35 ) | ( (~ Ng6275) ) ;
 assign n2651 = ( (~ Pg35) ) | ( (~ n2649) ) | ( (~ Ng6291) ) ;
 assign n2649 = ( n4581 ) | ( n2254 ) ;
 assign n2653 = ( Pg35 ) | ( (~ Ng6271) ) ;
 assign n2652 = ( n2254 ) | ( n4895 ) ;
 assign n2656 = ( Pg35 ) | ( (~ Ng6267) ) ;
 assign n2655 = ( n4836 ) | ( n2254 ) ;
 assign n2659 = ( Pg35 ) | ( (~ Ng6263) ) ;
 assign n2660 = ( (~ Pg35) ) | ( (~ n2658) ) | ( (~ Ng6279) ) ;
 assign n2658 = ( n2254 ) | ( n4896 ) ;
 assign n2662 = ( Pg35 ) | ( (~ Ng6255) ) ;
 assign n2661 = ( n4581 ) | ( n2255 ) ;
 assign n2665 = ( Pg35 ) | ( (~ Ng6247) ) ;
 assign n2666 = ( (~ Pg35) ) | ( (~ n2664) ) | ( (~ Ng6271) ) ;
 assign n2664 = ( n4895 ) | ( n2255 ) ;
 assign n2668 = ( Pg35 ) | ( (~ Ng6239) ) ;
 assign n2669 = ( (~ Pg35) ) | ( (~ n2667) ) | ( (~ Ng6267) ) ;
 assign n2667 = ( n4836 ) | ( n2255 ) ;
 assign n2671 = ( Pg35 ) | ( (~ Ng6235) ) ;
 assign n2672 = ( (~ Pg35) ) | ( (~ n2670) ) | ( (~ Ng6263) ) ;
 assign n2670 = ( n4896 ) | ( n2255 ) ;
 assign n2674 = ( Pg35 ) | ( (~ Ng6259) ) ;
 assign n2675 = ( (~ Pg35) ) | ( (~ n2673) ) | ( (~ Ng6255) ) ;
 assign n2673 = ( n4581 ) | ( n4900 ) ;
 assign n2677 = ( Pg35 ) | ( (~ Ng6251) ) ;
 assign n2678 = ( (~ Pg35) ) | ( (~ n2676) ) | ( (~ Ng6247) ) ;
 assign n2676 = ( n4895 ) | ( n4900 ) ;
 assign n2680 = ( Pg35 ) | ( (~ Ng6243) ) ;
 assign n2681 = ( (~ Pg35) ) | ( (~ n2679) ) | ( (~ Ng6239) ) ;
 assign n2679 = ( n4836 ) | ( n4900 ) ;
 assign n2683 = ( Pg35 ) | ( (~ Ng6227) ) ;
 assign n2684 = ( (~ Pg35) ) | ( (~ n2682) ) | ( (~ Ng6235) ) ;
 assign n2682 = ( n4896 ) | ( n4900 ) ;
 assign n2686 = ( n160  &  (~ n4901) ) | ( n3291  &  (~ n4901) ) | ( n160  &  (~ Ng5965) ) | ( n3291  &  (~ Ng5965) ) ;
 assign n2688 = ( Pg35 ) | ( (~ Ng5957) ) ;
 assign n2689 = ( (~ Pg35) ) | ( (~ n2687) ) | ( (~ Ng5913) ) ;
 assign n2687 = ( (~ Ng5869) ) | ( n4902 ) ;
 assign n2690 = ( Pg35 ) | ( (~ Ng5953) ) ;
 assign n2693 = ( Pg35 ) | ( (~ Ng5949) ) ;
 assign n2694 = ( (~ Pg35) ) | ( (~ n2692) ) | ( (~ Ng5897) ) ;
 assign n2692 = ( (~ Ng5869) ) | ( n4903 ) ;
 assign n2696 = ( Pg35 ) | ( (~ Ng5945) ) ;
 assign n2695 = ( n4590 ) | ( n2264 ) ;
 assign n2699 = ( Pg35 ) | ( (~ Ng5941) ) ;
 assign n2700 = ( (~ Pg35) ) | ( (~ n2698) ) | ( (~ Ng5957) ) ;
 assign n2698 = ( n2264 ) | ( n4902 ) ;
 assign n2702 = ( Pg35 ) | ( (~ Ng5937) ) ;
 assign n2703 = ( (~ Pg35) ) | ( (~ n2701) ) | ( (~ Ng5953) ) ;
 assign n2701 = ( n4837 ) | ( n2264 ) ;
 assign n2705 = ( Pg35 ) | ( (~ Ng5933) ) ;
 assign n2706 = ( (~ Pg35) ) | ( (~ n2704) ) | ( (~ Ng5949) ) ;
 assign n2704 = ( n2264 ) | ( n4903 ) ;
 assign n2708 = ( Pg35 ) | ( (~ Ng5929) ) ;
 assign n2709 = ( (~ Pg35) ) | ( (~ n2707) ) | ( (~ Ng5945) ) ;
 assign n2707 = ( n4590 ) | ( n2267 ) ;
 assign n2711 = ( Pg35 ) | ( (~ Ng5925) ) ;
 assign n2710 = ( n2267 ) | ( n4902 ) ;
 assign n2714 = ( Pg35 ) | ( (~ Ng5921) ) ;
 assign n2715 = ( (~ Pg35) ) | ( (~ n2713) ) | ( (~ Ng5937) ) ;
 assign n2713 = ( n4837 ) | ( n2267 ) ;
 assign n2717 = ( Pg35 ) | ( (~ Ng5917) ) ;
 assign n2718 = ( (~ Pg35) ) | ( (~ n2716) ) | ( (~ Ng5933) ) ;
 assign n2716 = ( n2267 ) | ( n4903 ) ;
 assign n2720 = ( Pg35 ) | ( (~ Ng5909) ) ;
 assign n2721 = ( (~ Pg35) ) | ( (~ n2719) ) | ( (~ Ng5929) ) ;
 assign n2719 = ( n4590 ) | ( n2268 ) ;
 assign n2723 = ( Pg35 ) | ( (~ Ng5901) ) ;
 assign n2724 = ( (~ Pg35) ) | ( (~ n2722) ) | ( (~ Ng5925) ) ;
 assign n2722 = ( n4902 ) | ( n2268 ) ;
 assign n2726 = ( Pg35 ) | ( (~ Ng5893) ) ;
 assign n2727 = ( (~ Pg35) ) | ( (~ n2725) ) | ( (~ Ng5921) ) ;
 assign n2725 = ( n4837 ) | ( n2268 ) ;
 assign n2729 = ( Pg35 ) | ( (~ Ng5889) ) ;
 assign n2730 = ( (~ Pg35) ) | ( (~ n2728) ) | ( (~ Ng5917) ) ;
 assign n2728 = ( n4903 ) | ( n2268 ) ;
 assign n2732 = ( Pg35 ) | ( (~ Ng5913) ) ;
 assign n2733 = ( (~ Pg35) ) | ( (~ n2731) ) | ( (~ Ng5909) ) ;
 assign n2731 = ( n4590 ) | ( n4907 ) ;
 assign n2735 = ( Pg35 ) | ( (~ Ng5905) ) ;
 assign n2736 = ( (~ Pg35) ) | ( (~ n2734) ) | ( (~ Ng5901) ) ;
 assign n2734 = ( n4902 ) | ( n4907 ) ;
 assign n2738 = ( Pg35 ) | ( (~ Ng5897) ) ;
 assign n2739 = ( (~ Pg35) ) | ( (~ n2737) ) | ( (~ Ng5893) ) ;
 assign n2737 = ( n4837 ) | ( n4907 ) ;
 assign n2741 = ( Pg35 ) | ( (~ Ng5881) ) ;
 assign n2742 = ( (~ Pg35) ) | ( (~ n2740) ) | ( (~ Ng5889) ) ;
 assign n2740 = ( n4903 ) | ( n4907 ) ;
 assign n2744 = ( n160  &  (~ n4908) ) | ( n3346  &  (~ n4908) ) | ( n160  &  (~ Ng5619) ) | ( n3346  &  (~ Ng5619) ) ;
 assign n2746 = ( Pg35 ) | ( (~ Ng5611) ) ;
 assign n2747 = ( (~ Pg35) ) | ( (~ n2745) ) | ( (~ Ng5567) ) ;
 assign n2745 = ( (~ Ng5523) ) | ( n4909 ) ;
 assign n2748 = ( Pg35 ) | ( (~ Ng5607) ) ;
 assign n2751 = ( Pg35 ) | ( (~ Ng5603) ) ;
 assign n2752 = ( (~ Pg35) ) | ( (~ n2750) ) | ( (~ Ng5551) ) ;
 assign n2750 = ( (~ Ng5523) ) | ( n4910 ) ;
 assign n2754 = ( Pg35 ) | ( (~ Ng5599) ) ;
 assign n2755 = ( (~ Pg35) ) | ( (~ n2753) ) | ( (~ Ng5615) ) ;
 assign n2753 = ( n4587 ) | ( n2277 ) ;
 assign n2757 = ( Pg35 ) | ( (~ Ng5595) ) ;
 assign n2758 = ( (~ Pg35) ) | ( (~ n2756) ) | ( (~ Ng5611) ) ;
 assign n2756 = ( n2277 ) | ( n4909 ) ;
 assign n2760 = ( Pg35 ) | ( (~ Ng5591) ) ;
 assign n2761 = ( (~ Pg35) ) | ( (~ n2759) ) | ( (~ Ng5607) ) ;
 assign n2759 = ( n4838 ) | ( n2277 ) ;
 assign n2763 = ( Pg35 ) | ( (~ Ng5587) ) ;
 assign n2764 = ( (~ Pg35) ) | ( (~ n2762) ) | ( (~ Ng5603) ) ;
 assign n2762 = ( n2277 ) | ( n4910 ) ;
 assign n2766 = ( Pg35 ) | ( (~ Ng5583) ) ;
 assign n2767 = ( (~ Pg35) ) | ( (~ n2765) ) | ( (~ Ng5599) ) ;
 assign n2765 = ( n4587 ) | ( n2280 ) ;
 assign n2769 = ( Pg35 ) | ( (~ Ng5579) ) ;
 assign n2768 = ( n2280 ) | ( n4909 ) ;
 assign n2772 = ( Pg35 ) | ( (~ Ng5575) ) ;
 assign n2773 = ( (~ Pg35) ) | ( (~ n2771) ) | ( (~ Ng5591) ) ;
 assign n2771 = ( n4838 ) | ( n2280 ) ;
 assign n2775 = ( Pg35 ) | ( (~ Ng5571) ) ;
 assign n2776 = ( (~ Pg35) ) | ( (~ n2774) ) | ( (~ Ng5587) ) ;
 assign n2774 = ( n2280 ) | ( n4910 ) ;
 assign n2778 = ( Pg35 ) | ( (~ Ng5563) ) ;
 assign n2779 = ( (~ Pg35) ) | ( (~ n2777) ) | ( (~ Ng5583) ) ;
 assign n2777 = ( n4587 ) | ( n2281 ) ;
 assign n2781 = ( Pg35 ) | ( (~ Ng5555) ) ;
 assign n2782 = ( (~ Pg35) ) | ( (~ n2780) ) | ( (~ Ng5579) ) ;
 assign n2780 = ( n4909 ) | ( n2281 ) ;
 assign n2784 = ( Pg35 ) | ( (~ Ng5547) ) ;
 assign n2785 = ( (~ Pg35) ) | ( (~ n2783) ) | ( (~ Ng5575) ) ;
 assign n2783 = ( n4838 ) | ( n2281 ) ;
 assign n2787 = ( Pg35 ) | ( (~ Ng5543) ) ;
 assign n2788 = ( (~ Pg35) ) | ( (~ n2786) ) | ( (~ Ng5571) ) ;
 assign n2786 = ( n4910 ) | ( n2281 ) ;
 assign n2790 = ( Pg35 ) | ( (~ Ng5567) ) ;
 assign n2791 = ( (~ Pg35) ) | ( (~ n2789) ) | ( (~ Ng5563) ) ;
 assign n2789 = ( n4587 ) | ( n4914 ) ;
 assign n2793 = ( Pg35 ) | ( (~ Ng5559) ) ;
 assign n2794 = ( (~ Pg35) ) | ( (~ n2792) ) | ( (~ Ng5555) ) ;
 assign n2792 = ( n4909 ) | ( n4914 ) ;
 assign n2796 = ( Pg35 ) | ( (~ Ng5551) ) ;
 assign n2797 = ( (~ Pg35) ) | ( (~ n2795) ) | ( (~ Ng5547) ) ;
 assign n2795 = ( n4838 ) | ( n4914 ) ;
 assign n2799 = ( Pg35 ) | ( (~ Ng5535) ) ;
 assign n2800 = ( (~ Pg35) ) | ( (~ n2798) ) | ( (~ Ng5543) ) ;
 assign n2798 = ( n4910 ) | ( n4914 ) ;
 assign n2802 = ( n160  &  n4092 ) | ( n3401  &  n4092 ) | ( n160  &  (~ Ng5272) ) | ( n3401  &  (~ Ng5272) ) ;
 assign n2804 = ( Pg35 ) | ( (~ Ng5264) ) ;
 assign n2805 = ( (~ Pg35) ) | ( (~ n2803) ) | ( (~ Ng5220) ) ;
 assign n2803 = ( (~ Ng5176) ) | ( n4915 ) ;
 assign n2806 = ( Pg35 ) | ( (~ Ng5260) ) ;
 assign n2807 = ( (~ Pg35) ) | ( (~ n2284) ) | ( (~ Ng5212) ) ;
 assign n2809 = ( Pg35 ) | ( (~ Ng5256) ) ;
 assign n2810 = ( (~ Pg35) ) | ( (~ n2808) ) | ( (~ Ng5204) ) ;
 assign n2808 = ( (~ Ng5176) ) | ( n4916 ) ;
 assign n2812 = ( Pg35 ) | ( (~ Ng5252) ) ;
 assign n2813 = ( (~ Pg35) ) | ( (~ n2811) ) | ( (~ Ng5268) ) ;
 assign n2811 = ( n4595 ) | ( n2290 ) ;
 assign n2815 = ( Pg35 ) | ( (~ Ng5248) ) ;
 assign n2816 = ( (~ Pg35) ) | ( (~ n2814) ) | ( (~ Ng5264) ) ;
 assign n2814 = ( n2290 ) | ( n4915 ) ;
 assign n2818 = ( Pg35 ) | ( (~ Ng5244) ) ;
 assign n2817 = ( n4839 ) | ( n2290 ) ;
 assign n2821 = ( Pg35 ) | ( (~ Ng5240) ) ;
 assign n2822 = ( (~ Pg35) ) | ( (~ n2820) ) | ( (~ Ng5256) ) ;
 assign n2820 = ( n2290 ) | ( n4916 ) ;
 assign n2824 = ( Pg35 ) | ( (~ Ng5236) ) ;
 assign n2823 = ( n4595 ) | ( n2293 ) ;
 assign n2827 = ( Pg35 ) | ( (~ Ng5232) ) ;
 assign n2826 = ( n2293 ) | ( n4915 ) ;
 assign n2830 = ( Pg35 ) | ( (~ Ng5228) ) ;
 assign n2831 = ( (~ Pg35) ) | ( (~ n2829) ) | ( (~ Ng5244) ) ;
 assign n2829 = ( n4839 ) | ( n2293 ) ;
 assign n2833 = ( Pg35 ) | ( (~ Ng5224) ) ;
 assign n2834 = ( (~ Pg35) ) | ( (~ n2832) ) | ( (~ Ng5240) ) ;
 assign n2832 = ( n2293 ) | ( n4916 ) ;
 assign n2836 = ( Pg35 ) | ( (~ Ng5216) ) ;
 assign n2837 = ( (~ Pg35) ) | ( (~ n2835) ) | ( (~ Ng5236) ) ;
 assign n2835 = ( n4595 ) | ( n2294 ) ;
 assign n2839 = ( Pg35 ) | ( (~ Ng5208) ) ;
 assign n2840 = ( (~ Pg35) ) | ( (~ n2838) ) | ( (~ Ng5232) ) ;
 assign n2838 = ( n4915 ) | ( n2294 ) ;
 assign n2842 = ( Pg35 ) | ( (~ Ng5200) ) ;
 assign n2843 = ( (~ Pg35) ) | ( (~ n2841) ) | ( (~ Ng5228) ) ;
 assign n2841 = ( n4839 ) | ( n2294 ) ;
 assign n2845 = ( Pg35 ) | ( (~ Ng5196) ) ;
 assign n2846 = ( (~ Pg35) ) | ( (~ n2844) ) | ( (~ Ng5224) ) ;
 assign n2844 = ( n4916 ) | ( n2294 ) ;
 assign n2848 = ( Pg35 ) | ( (~ Ng5220) ) ;
 assign n2849 = ( (~ Pg35) ) | ( (~ n2847) ) | ( (~ Ng5216) ) ;
 assign n2847 = ( n4595 ) | ( n4919 ) ;
 assign n2851 = ( Pg35 ) | ( (~ Ng5212) ) ;
 assign n2852 = ( (~ Pg35) ) | ( (~ n2850) ) | ( (~ Ng5208) ) ;
 assign n2850 = ( n4915 ) | ( n4919 ) ;
 assign n2854 = ( Pg35 ) | ( (~ Ng5204) ) ;
 assign n2855 = ( (~ Pg35) ) | ( (~ n2853) ) | ( (~ Ng5200) ) ;
 assign n2853 = ( n4839 ) | ( n4919 ) ;
 assign n2857 = ( Pg35 ) | ( (~ Ng5188) ) ;
 assign n2858 = ( (~ Pg35) ) | ( (~ n2856) ) | ( (~ Ng5196) ) ;
 assign n2856 = ( n4916 ) | ( n4919 ) ;
 assign n2860 = ( (~ Pg113)  &  (~ Ng4507) ) | ( (~ Ng4507)  &  n5821 ) | ( (~ Pg113)  &  (~ n5821) ) ;
 assign n2859 = ( n2860  &  Pg35 ) ;
 assign n2862 = ( (~ Pg115) ) | ( Ng4157 ) | ( n5828 ) ;
 assign n2863 = ( Pg115 ) | ( Ng4157 ) | ( (~ n5828) ) ;
 assign n2864 = ( (~ Pg126) ) | ( Ng4146 ) | ( n5825 ) ;
 assign n2865 = ( Pg126 ) | ( Ng4146 ) | ( (~ n5825) ) ;
 assign n2861 = ( n2862  &  n2863  &  n2864  &  n2865 ) ;
 assign n2867 = ( n3474 ) | ( (~ Ng4093) ) | ( (~ n4790) ) ;
 assign n2868 = ( Ng4093 ) | ( n4790 ) | ( (~ Ng2841) ) ;
 assign n2870 = ( n160  &  (~ n4922) ) | ( n3476  &  (~ n4922) ) | ( n160  &  (~ Ng3965) ) | ( n3476  &  (~ Ng3965) ) ;
 assign n2872 = ( Pg35 ) | ( (~ Ng3957) ) ;
 assign n2873 = ( (~ Pg35) ) | ( (~ n2871) ) | ( (~ Ng3913) ) ;
 assign n2871 = ( (~ Ng3869) ) | ( n4923 ) ;
 assign n2874 = ( Pg35 ) | ( (~ Ng3953) ) ;
 assign n2875 = ( (~ Pg35) ) | ( (~ n2320) ) | ( (~ Ng3905) ) ;
 assign n2877 = ( Pg35 ) | ( (~ Ng3949) ) ;
 assign n2878 = ( (~ Pg35) ) | ( (~ n2876) ) | ( (~ Ng3897) ) ;
 assign n2876 = ( (~ Ng3869) ) | ( n4924 ) ;
 assign n2880 = ( Pg35 ) | ( (~ Ng3945) ) ;
 assign n2881 = ( (~ Pg35) ) | ( (~ n2879) ) | ( (~ Ng3961) ) ;
 assign n2879 = ( n4584 ) | ( n2326 ) ;
 assign n2883 = ( Pg35 ) | ( (~ Ng3941) ) ;
 assign n2884 = ( (~ Pg35) ) | ( (~ n2882) ) | ( (~ Ng3957) ) ;
 assign n2882 = ( n2326 ) | ( n4923 ) ;
 assign n2886 = ( Pg35 ) | ( (~ Ng3937) ) ;
 assign n2885 = ( n4855 ) | ( n2326 ) ;
 assign n2889 = ( Pg35 ) | ( (~ Ng3933) ) ;
 assign n2890 = ( (~ Pg35) ) | ( (~ n2888) ) | ( (~ Ng3949) ) ;
 assign n2888 = ( n2326 ) | ( n4924 ) ;
 assign n2892 = ( Pg35 ) | ( (~ Ng3929) ) ;
 assign n2891 = ( n4584 ) | ( n2329 ) ;
 assign n2895 = ( Pg35 ) | ( (~ Ng3925) ) ;
 assign n2894 = ( n2329 ) | ( n4923 ) ;
 assign n2898 = ( Pg35 ) | ( (~ Ng3921) ) ;
 assign n2899 = ( (~ Pg35) ) | ( (~ n2897) ) | ( (~ Ng3937) ) ;
 assign n2897 = ( n4855 ) | ( n2329 ) ;
 assign n2901 = ( Pg35 ) | ( (~ Ng3917) ) ;
 assign n2902 = ( (~ Pg35) ) | ( (~ n2900) ) | ( (~ Ng3933) ) ;
 assign n2900 = ( n2329 ) | ( n4924 ) ;
 assign n2904 = ( Pg35 ) | ( (~ Ng3909) ) ;
 assign n2905 = ( (~ Pg35) ) | ( (~ n2903) ) | ( (~ Ng3929) ) ;
 assign n2903 = ( n4584 ) | ( n2330 ) ;
 assign n2907 = ( Pg35 ) | ( (~ Ng3901) ) ;
 assign n2908 = ( (~ Pg35) ) | ( (~ n2906) ) | ( (~ Ng3925) ) ;
 assign n2906 = ( n4923 ) | ( n2330 ) ;
 assign n2910 = ( Pg35 ) | ( (~ Ng3893) ) ;
 assign n2911 = ( (~ Pg35) ) | ( (~ n2909) ) | ( (~ Ng3921) ) ;
 assign n2909 = ( n4855 ) | ( n2330 ) ;
 assign n2913 = ( Pg35 ) | ( (~ Ng3889) ) ;
 assign n2914 = ( (~ Pg35) ) | ( (~ n2912) ) | ( (~ Ng3917) ) ;
 assign n2912 = ( n4924 ) | ( n2330 ) ;
 assign n2916 = ( Pg35 ) | ( (~ Ng3913) ) ;
 assign n2917 = ( (~ Pg35) ) | ( (~ n2915) ) | ( (~ Ng3909) ) ;
 assign n2915 = ( n4584 ) | ( n4927 ) ;
 assign n2919 = ( Pg35 ) | ( (~ Ng3905) ) ;
 assign n2920 = ( (~ Pg35) ) | ( (~ n2918) ) | ( (~ Ng3901) ) ;
 assign n2918 = ( n4923 ) | ( n4927 ) ;
 assign n2922 = ( Pg35 ) | ( (~ Ng3897) ) ;
 assign n2923 = ( (~ Pg35) ) | ( (~ n2921) ) | ( (~ Ng3893) ) ;
 assign n2921 = ( n4855 ) | ( n4927 ) ;
 assign n2925 = ( Pg35 ) | ( (~ Ng3881) ) ;
 assign n2926 = ( (~ Pg35) ) | ( (~ n2924) ) | ( (~ Ng3889) ) ;
 assign n2924 = ( n4924 ) | ( n4927 ) ;
 assign n2928 = ( n160  &  (~ n4928) ) | ( n3531  &  (~ n4928) ) | ( n160  &  (~ Ng3614) ) | ( n3531  &  (~ Ng3614) ) ;
 assign n2930 = ( Pg35 ) | ( (~ Ng3606) ) ;
 assign n2931 = ( (~ Pg35) ) | ( (~ n2929) ) | ( (~ Ng3562) ) ;
 assign n2929 = ( (~ Ng3518) ) | ( n4929 ) ;
 assign n2932 = ( Pg35 ) | ( (~ Ng3602) ) ;
 assign n2933 = ( (~ Pg35) ) | ( (~ n2333) ) | ( (~ Ng3554) ) ;
 assign n2935 = ( Pg35 ) | ( (~ Ng3598) ) ;
 assign n2936 = ( (~ Pg35) ) | ( (~ n2934) ) | ( (~ Ng3546) ) ;
 assign n2934 = ( (~ Ng3518) ) | ( n4930 ) ;
 assign n2938 = ( Pg35 ) | ( (~ Ng3594) ) ;
 assign n2939 = ( (~ Pg35) ) | ( (~ n2937) ) | ( (~ Ng3610) ) ;
 assign n2937 = ( n4593 ) | ( n2339 ) ;
 assign n2941 = ( Pg35 ) | ( (~ Ng3590) ) ;
 assign n2942 = ( (~ Pg35) ) | ( (~ n2940) ) | ( (~ Ng3606) ) ;
 assign n2940 = ( n2339 ) | ( n4929 ) ;
 assign n2944 = ( Pg35 ) | ( (~ Ng3586) ) ;
 assign n2943 = ( n4856 ) | ( n2339 ) ;
 assign n2947 = ( Pg35 ) | ( (~ Ng3582) ) ;
 assign n2948 = ( (~ Pg35) ) | ( (~ n2946) ) | ( (~ Ng3598) ) ;
 assign n2946 = ( n2339 ) | ( n4930 ) ;
 assign n2950 = ( Pg35 ) | ( (~ Ng3578) ) ;
 assign n2951 = ( (~ Pg35) ) | ( (~ n2949) ) | ( (~ Ng3594) ) ;
 assign n2949 = ( n4593 ) | ( n2342 ) ;
 assign n2953 = ( Pg35 ) | ( (~ Ng3574) ) ;
 assign n2952 = ( n2342 ) | ( n4929 ) ;
 assign n2956 = ( Pg35 ) | ( (~ Ng3570) ) ;
 assign n2957 = ( (~ Pg35) ) | ( (~ n2955) ) | ( (~ Ng3586) ) ;
 assign n2955 = ( n4856 ) | ( n2342 ) ;
 assign n2959 = ( Pg35 ) | ( (~ Ng3566) ) ;
 assign n2960 = ( (~ Pg35) ) | ( (~ n2958) ) | ( (~ Ng3582) ) ;
 assign n2958 = ( n2342 ) | ( n4930 ) ;
 assign n2962 = ( Pg35 ) | ( (~ Ng3558) ) ;
 assign n2961 = ( n4593 ) | ( n2343 ) ;
 assign n2965 = ( Pg35 ) | ( (~ Ng3550) ) ;
 assign n2966 = ( (~ Pg35) ) | ( (~ n2964) ) | ( (~ Ng3574) ) ;
 assign n2964 = ( n4929 ) | ( n2343 ) ;
 assign n2968 = ( Pg35 ) | ( (~ Ng3542) ) ;
 assign n2969 = ( (~ Pg35) ) | ( (~ n2967) ) | ( (~ Ng3570) ) ;
 assign n2967 = ( n4856 ) | ( n2343 ) ;
 assign n2971 = ( Pg35 ) | ( (~ Ng3538) ) ;
 assign n2972 = ( (~ Pg35) ) | ( (~ n2970) ) | ( (~ Ng3566) ) ;
 assign n2970 = ( n4930 ) | ( n2343 ) ;
 assign n2974 = ( Pg35 ) | ( (~ Ng3562) ) ;
 assign n2975 = ( (~ Pg35) ) | ( (~ n2973) ) | ( (~ Ng3558) ) ;
 assign n2973 = ( n4593 ) | ( n4933 ) ;
 assign n2977 = ( Pg35 ) | ( (~ Ng3554) ) ;
 assign n2978 = ( (~ Pg35) ) | ( (~ n2976) ) | ( (~ Ng3550) ) ;
 assign n2976 = ( n4929 ) | ( n4933 ) ;
 assign n2980 = ( Pg35 ) | ( (~ Ng3546) ) ;
 assign n2981 = ( (~ Pg35) ) | ( (~ n2979) ) | ( (~ Ng3542) ) ;
 assign n2979 = ( n4856 ) | ( n4933 ) ;
 assign n2983 = ( Pg35 ) | ( (~ Ng3530) ) ;
 assign n2984 = ( (~ Pg35) ) | ( (~ n2982) ) | ( (~ Ng3538) ) ;
 assign n2982 = ( n4930 ) | ( n4933 ) ;
 assign n2986 = ( n160  &  (~ n4934) ) | ( n3583  &  (~ n4934) ) | ( n160  &  (~ Ng3263) ) | ( n3583  &  (~ Ng3263) ) ;
 assign n2988 = ( Pg35 ) | ( (~ Ng3255) ) ;
 assign n2989 = ( (~ Pg35) ) | ( (~ n2987) ) | ( (~ Ng3211) ) ;
 assign n2987 = ( (~ Ng3167) ) | ( n4935 ) ;
 assign n2990 = ( Pg35 ) | ( (~ Ng3251) ) ;
 assign n2991 = ( (~ Pg35) ) | ( (~ n2346) ) | ( (~ Ng3203) ) ;
 assign n2993 = ( Pg35 ) | ( (~ Ng3247) ) ;
 assign n2994 = ( (~ Pg35) ) | ( (~ n2992) ) | ( (~ Ng3195) ) ;
 assign n2992 = ( (~ Ng3167) ) | ( n4936 ) ;
 assign n2996 = ( Pg35 ) | ( (~ Ng3243) ) ;
 assign n2997 = ( (~ Pg35) ) | ( (~ n2995) ) | ( (~ Ng3259) ) ;
 assign n2995 = ( n4577 ) | ( n2352 ) ;
 assign n2999 = ( Pg35 ) | ( (~ Ng3239) ) ;
 assign n3000 = ( (~ Pg35) ) | ( (~ n2998) ) | ( (~ Ng3255) ) ;
 assign n2998 = ( n2352 ) | ( n4935 ) ;
 assign n3002 = ( Pg35 ) | ( (~ Ng3235) ) ;
 assign n3003 = ( (~ Pg35) ) | ( (~ n3001) ) | ( (~ Ng3251) ) ;
 assign n3001 = ( n4857 ) | ( n2352 ) ;
 assign n3005 = ( Pg35 ) | ( (~ Ng3231) ) ;
 assign n3006 = ( (~ Pg35) ) | ( (~ n3004) ) | ( (~ Ng3247) ) ;
 assign n3004 = ( n2352 ) | ( n4936 ) ;
 assign n3008 = ( Pg35 ) | ( (~ Ng3227) ) ;
 assign n3009 = ( (~ Pg35) ) | ( (~ n3007) ) | ( (~ Ng3243) ) ;
 assign n3007 = ( n4577 ) | ( n2355 ) ;
 assign n3011 = ( Pg35 ) | ( (~ Ng3223) ) ;
 assign n3010 = ( n2355 ) | ( n4935 ) ;
 assign n3014 = ( Pg35 ) | ( (~ Ng3219) ) ;
 assign n3013 = ( n4857 ) | ( n2355 ) ;
 assign n3017 = ( Pg35 ) | ( (~ Ng3215) ) ;
 assign n3018 = ( (~ Pg35) ) | ( (~ n3016) ) | ( (~ Ng3231) ) ;
 assign n3016 = ( n2355 ) | ( n4936 ) ;
 assign n3020 = ( Pg35 ) | ( (~ Ng3207) ) ;
 assign n3019 = ( n4577 ) | ( n2356 ) ;
 assign n3023 = ( Pg35 ) | ( (~ Ng3199) ) ;
 assign n3024 = ( (~ Pg35) ) | ( (~ n3022) ) | ( (~ Ng3223) ) ;
 assign n3022 = ( n4935 ) | ( n2356 ) ;
 assign n3026 = ( Pg35 ) | ( (~ Ng3191) ) ;
 assign n3027 = ( (~ Pg35) ) | ( (~ n3025) ) | ( (~ Ng3219) ) ;
 assign n3025 = ( n4857 ) | ( n2356 ) ;
 assign n3029 = ( Pg35 ) | ( (~ Ng3187) ) ;
 assign n3030 = ( (~ Pg35) ) | ( (~ n3028) ) | ( (~ Ng3215) ) ;
 assign n3028 = ( n4936 ) | ( n2356 ) ;
 assign n3032 = ( Pg35 ) | ( (~ Ng3211) ) ;
 assign n3033 = ( (~ Pg35) ) | ( (~ n3031) ) | ( (~ Ng3207) ) ;
 assign n3031 = ( n4577 ) | ( n4940 ) ;
 assign n3035 = ( Pg35 ) | ( (~ Ng3203) ) ;
 assign n3036 = ( (~ Pg35) ) | ( (~ n3034) ) | ( (~ Ng3199) ) ;
 assign n3034 = ( n4935 ) | ( n4940 ) ;
 assign n3038 = ( Pg35 ) | ( (~ Ng3195) ) ;
 assign n3039 = ( (~ Pg35) ) | ( (~ n3037) ) | ( (~ Ng3191) ) ;
 assign n3037 = ( n4857 ) | ( n4940 ) ;
 assign n3041 = ( Pg35 ) | ( (~ Ng3179) ) ;
 assign n3042 = ( (~ Pg35) ) | ( (~ n3040) ) | ( (~ Ng3187) ) ;
 assign n3040 = ( n4936 ) | ( n4940 ) ;
 assign n3043 = ( (~ Pg35) ) | ( n5832 ) | ( n5833 ) ;
 assign n3044 = ( (~ Pg35) ) | ( n5837 ) | ( n5838 ) ;
 assign n3045 = ( (~ n4346)  &  Ng2741 ) | ( n4346  &  (~ Ng2741) ) ;
 assign n3046 = ( (~ Pg35) ) | ( (~ Ng2841) ) ;
 assign n3050 = ( Ng2675 ) | ( (~ n4946) ) | ( Ng2681 ) ;
 assign n3048 = ( (~ Pg35) ) | ( n4945 ) ;
 assign n3053 = ( n3048  &  (~ n4946) ) | ( n3048  &  Ng2661 ) | ( (~ n4946)  &  (~ Ng2661) ) ;
 assign n3056 = ( n4347 ) | ( n4860 ) | ( n4947 ) ;
 assign n3059 = ( n4702 ) | ( n4550 ) | ( n4860 ) ;
 assign n3062 = ( Ng2541 ) | ( (~ n4950) ) | ( Ng2547 ) ;
 assign n3060 = ( (~ Pg35) ) | ( n4949 ) ;
 assign n3065 = ( n3060  &  Ng2527 ) | ( n3060  &  (~ n4950) ) | ( (~ Ng2527)  &  (~ n4950) ) ;
 assign n3068 = ( n4348 ) | ( n4864 ) | ( n4951 ) ;
 assign n3071 = ( n4712 ) | ( n4546 ) | ( n4864 ) ;
 assign n3074 = ( Ng2407 ) | ( (~ n4953) ) | ( Ng2413 ) ;
 assign n3072 = ( (~ Pg35) ) | ( n4952 ) ;
 assign n3077 = ( n3072  &  (~ n4953) ) | ( n3072  &  Ng2393 ) | ( (~ n4953)  &  (~ Ng2393) ) ;
 assign n3080 = ( n4349 ) | ( n4866 ) | ( n4954 ) ;
 assign n3083 = ( n4722 ) | ( n4548 ) | ( n4866 ) ;
 assign n3086 = ( Ng2273 ) | ( (~ n4956) ) | ( Ng2279 ) ;
 assign n3084 = ( (~ Pg35) ) | ( n4955 ) ;
 assign n3089 = ( n3084  &  (~ n4956) ) | ( n3084  &  Ng2259 ) | ( (~ n4956)  &  (~ Ng2259) ) ;
 assign n3092 = ( n4350 ) | ( n4870 ) | ( n4957 ) ;
 assign n3095 = ( n4733 ) | ( n4535 ) | ( n4870 ) ;
 assign n3098 = ( Ng2116 ) | ( (~ n4960) ) | ( Ng2122 ) ;
 assign n3096 = ( (~ Pg35) ) | ( n4959 ) ;
 assign n3101 = ( n3096  &  Ng2102 ) | ( n3096  &  (~ n4960) ) | ( (~ Ng2102)  &  (~ n4960) ) ;
 assign n3104 = ( n4351 ) | ( n4873 ) | ( n4961 ) ;
 assign n3107 = ( n4744 ) | ( n4542 ) | ( n4873 ) ;
 assign n3110 = ( Ng1982 ) | ( (~ n4963) ) | ( Ng1988 ) ;
 assign n3108 = ( (~ Pg35) ) | ( n4962 ) ;
 assign n3113 = ( n3108  &  Ng1968 ) | ( n3108  &  (~ n4963) ) | ( (~ Ng1968)  &  (~ n4963) ) ;
 assign n3116 = ( n4352 ) | ( n4875 ) | ( n4964 ) ;
 assign n3119 = ( n4754 ) | ( n4544 ) | ( n4875 ) ;
 assign n3122 = ( Ng1848 ) | ( (~ n4966) ) | ( Ng1854 ) ;
 assign n3120 = ( (~ Pg35) ) | ( n4965 ) ;
 assign n3125 = ( n3120  &  (~ n4966) ) | ( n3120  &  Ng1834 ) | ( (~ n4966)  &  (~ Ng1834) ) ;
 assign n3128 = ( n4353 ) | ( n4878 ) | ( n4967 ) ;
 assign n3131 = ( n4763 ) | ( n4538 ) | ( n4878 ) ;
 assign n3134 = ( Ng1714 ) | ( (~ n4969) ) | ( Ng1720 ) ;
 assign n3132 = ( (~ Pg35) ) | ( n4968 ) ;
 assign n3137 = ( n3132  &  (~ n4969) ) | ( n3132  &  Ng1700 ) | ( (~ n4969)  &  (~ Ng1700) ) ;
 assign n3140 = ( n4354 ) | ( n4881 ) | ( n4970 ) ;
 assign n3141 = ( (~ Ng1636)  &  (~ n4553)  &  (~ n4881) ) | ( Ng1592  &  (~ n4553)  &  (~ n4881) ) ;
 assign n3148 = ( (~ n923)  &  (~ Ng1526) ) | ( (~ n923)  &  (~ n3151) ) ;
 assign n3152 = ( Pg35  &  n3148 ) | ( (~ Pg35)  &  (~ Ng1514) ) | ( n3148  &  (~ Ng1514) ) ;
 assign n3151 = ( (~ Pg7946) ) | ( (~ Ng1514) ) ;
 assign n3154 = ( (~ Pg35) ) | ( n2192 ) | ( (~ Ng1361) ) ;
 assign n3155 = ( (~ n2192) ) | ( Ng1361 ) | ( n3875 ) ;
 assign n3157 = ( (~ Ng1259) ) | ( (~ n3156) ) | ( n4222 ) ;
 assign n3158 = ( Pg35 ) | ( (~ Ng1256) ) ;
 assign n3156 = ( (~ Ng1256) ) | ( (~ n4810) ) ;
 assign n3160 = ( Ng1024  &  Ng1002  &  Ng1036  &  n4323 ) ;
 assign n3159 = ( Ng1008 ) | ( Ng969 ) | ( n3160 ) ;
 assign n3163 = ( (~ n330)  &  (~ Ng1183) ) | ( (~ n330)  &  (~ n3167) ) ;
 assign n3168 = ( (~ Pg35)  &  (~ Ng1171) ) | ( Pg35  &  n3163 ) | ( (~ Ng1171)  &  n3163 ) ;
 assign n3167 = ( (~ Pg7916) ) | ( (~ Ng1171) ) ;
 assign n3170 = ( (~ Pg35) ) | ( n2205 ) | ( (~ Ng1018) ) ;
 assign n3171 = ( (~ n2205) ) | ( Ng1018 ) | ( n3881 ) ;
 assign n3173 = ( (~ Ng914) ) | ( (~ n3172) ) | ( n4235 ) ;
 assign n3174 = ( Pg35 ) | ( (~ Ng911) ) ;
 assign n3172 = ( (~ Ng911) ) | ( (~ n4823) ) ;
 assign n3176 = ( (~ Ng744) ) | ( (~ n3175) ) | ( n3791 ) ;
 assign n3177 = ( Pg35 ) | ( (~ Ng739) ) ;
 assign n3175 = ( (~ n1369) ) | ( (~ Ng739) ) | ( n4490 ) ;
 assign n3179 = ( (~ Ng577) ) | ( (~ n3178) ) | ( n4508 ) ;
 assign n3180 = ( Pg35 ) | ( (~ Ng586) ) ;
 assign n3178 = ( (~ Ng586) ) | ( n3805 ) ;
 assign n3181 = ( n359  &  Ng146 ) | ( (~ n359)  &  (~ Ng146) ) ;
 assign n3182 = ( (~ Pg35) ) | ( n4666 ) ;
 assign n3185 = ( (~ Ng6541) ) | ( (~ n4886) ) | ( (~ n4887) ) ;
 assign n3184 = ( (~ Ng6561) ) | ( n4588 ) ;
 assign n3187 = ( n3188  &  n4984 ) | ( n3188  &  Ng6527 ) | ( n4984  &  (~ Ng6527) ) ;
 assign n3189 = ( Ng6513 ) | ( n4984 ) | ( Ng6519 ) ;
 assign n3188 = ( (~ Pg35) ) | ( (~ n4983) ) ;
 assign n3192 = ( Ng6500 ) | ( n4984 ) | ( (~ Ng6505) ) ;
 assign n3194 = ( (~ Pg13099)  &  (~ Ng6605) ) | ( (~ Ng6605)  &  (~ Ng6593) ) | ( (~ Pg13099)  &  (~ Ng6723) ) | ( (~ Ng6593)  &  (~ Ng6723) ) ;
 assign n3198 = ( (~ Pg17764)  &  (~ Pg17722) ) | ( (~ Pg17722)  &  (~ Ng6649) ) | ( (~ Pg17764)  &  (~ Ng6597) ) | ( (~ Ng6649)  &  (~ Ng6597) ) ;
 assign n3202 = ( (~ Pg17871)  &  (~ Pg12470) ) | ( (~ Pg12470)  &  (~ Ng6617) ) | ( (~ Pg17871)  &  (~ Ng6601) ) | ( (~ Ng6617)  &  (~ Ng6601) ) ;
 assign n3209 = ( (~ Pg14749) ) | ( n3223 ) | ( (~ Ng6633) ) ;
 assign n3210 = ( n3198  &  n3194 ) | ( n1956  &  n3194 ) | ( n3198  &  n3227 ) | ( n1956  &  n3227 ) ;
 assign n3208 = ( (~ Ng6741) ) | ( (~ Ng6682) ) ;
 assign n3207 = ( n3209  &  n3210  &  n3202 ) | ( n3209  &  n3210  &  n3208 ) ;
 assign n3211 = ( (~ Pg13099)  &  (~ Ng6589) ) | ( (~ Ng6589)  &  (~ Ng6581) ) | ( (~ Pg13099)  &  (~ Ng6723) ) | ( (~ Ng6581)  &  (~ Ng6723) ) ;
 assign n3214 = ( (~ Pg17871)  &  (~ Pg12470) ) | ( (~ Pg12470)  &  (~ Ng6609) ) | ( (~ Pg17871)  &  (~ Ng6585) ) | ( (~ Ng6609)  &  (~ Ng6585) ) ;
 assign n3218 = ( (~ Pg17764) ) | ( n3208 ) | ( (~ Ng6641) ) ;
 assign n3219 = ( (~ Pg14749) ) | ( n3227 ) | ( (~ Ng6625) ) ;
 assign n3220 = ( n3214  &  n3211 ) | ( n1956  &  n3211 ) | ( n3214  &  n3223 ) | ( n1956  &  n3223 ) ;
 assign n3217 = ( n3218  &  n3219  &  n3220 ) ;
 assign n3225 = ( (~ Pg17778)  &  n5602 ) | ( n1956  &  n5602 ) | ( (~ Ng6637)  &  n5602 ) ;
 assign n3223 = ( Ng6682 ) | ( Ng6741 ) ;
 assign n3221 = ( (~ Pg14828)  &  n3225 ) | ( n3225  &  n3223 ) | ( n3225  &  (~ Ng6621) ) ;
 assign n3229 = ( (~ Pg17778)  &  n5601 ) | ( n3208  &  n5601 ) | ( (~ Ng6629)  &  n5601 ) ;
 assign n3227 = ( Ng6741 ) | ( (~ Ng6682) ) ;
 assign n3226 = ( (~ Pg14828)  &  n3229 ) | ( n3229  &  n3227 ) | ( n3229  &  (~ Ng6613) ) ;
 assign n3233 = ( n3207  &  n3217 ) | ( n3217  &  Ng6727 ) | ( n3207  &  (~ Ng6727) ) ;
 assign n3234 = ( n3221  &  n3226 ) | ( n3226  &  n5886 ) | ( n3221  &  (~ n5886) ) ;
 assign n3232 = ( (~ Pg17722) ) | ( n3208 ) | ( (~ Ng6727) ) ;
 assign n3230 = ( n3233  &  n3234  &  n3232 ) | ( n3233  &  n3234  &  (~ Ng6657) ) ;
 assign n3236 = ( Pg35 ) | ( (~ Ng6505) ) ;
 assign n3235 = ( (~ Pg35) ) | ( (~ n1109) ) | ( n3230 ) ;
 assign n3239 = ( (~ Ng6195) ) | ( (~ n4887) ) | ( (~ n4894) ) ;
 assign n3238 = ( (~ Ng6215) ) | ( n4581 ) ;
 assign n3241 = ( n3242  &  n4991 ) | ( n3242  &  Ng6181 ) | ( n4991  &  (~ Ng6181) ) ;
 assign n3243 = ( Ng6167 ) | ( n4991 ) | ( Ng6173 ) ;
 assign n3242 = ( (~ Pg35) ) | ( (~ n4990) ) ;
 assign n3247 = ( Ng6154 ) | ( n4991 ) | ( (~ Ng6159) ) ;
 assign n3249 = ( (~ Pg17743)  &  (~ Pg17685) ) | ( (~ Pg17685)  &  (~ Ng6303) ) | ( (~ Pg17743)  &  (~ Ng6251) ) | ( (~ Ng6303)  &  (~ Ng6251) ) ;
 assign n3253 = ( (~ Pg13085)  &  (~ Ng6259) ) | ( (~ Ng6259)  &  (~ Ng6247) ) | ( (~ Pg13085)  &  (~ Ng6377) ) | ( (~ Ng6247)  &  (~ Ng6377) ) ;
 assign n3257 = ( (~ Pg17845)  &  (~ Pg12422) ) | ( (~ Pg12422)  &  (~ Ng6271) ) | ( (~ Pg17845)  &  (~ Ng6255) ) | ( (~ Ng6271)  &  (~ Ng6255) ) ;
 assign n3264 = ( (~ Pg14705) ) | ( n3281 ) | ( (~ Ng6287) ) ;
 assign n3265 = ( n3253  &  n3249 ) | ( n3277  &  n3249 ) | ( n3253  &  n1965 ) | ( n3277  &  n1965 ) ;
 assign n3263 = ( (~ Ng6395) ) | ( (~ Ng6336) ) ;
 assign n3262 = ( n3264  &  n3265  &  n3257 ) | ( n3264  &  n3265  &  n3263 ) ;
 assign n3266 = ( (~ Pg13085)  &  (~ Ng6243) ) | ( (~ Ng6243)  &  (~ Ng6235) ) | ( (~ Pg13085)  &  (~ Ng6377) ) | ( (~ Ng6235)  &  (~ Ng6377) ) ;
 assign n3269 = ( (~ Pg17845)  &  (~ Pg12422) ) | ( (~ Pg12422)  &  (~ Ng6263) ) | ( (~ Pg17845)  &  (~ Ng6239) ) | ( (~ Ng6263)  &  (~ Ng6239) ) ;
 assign n3273 = ( (~ Pg17743) ) | ( n3263 ) | ( (~ Ng6295) ) ;
 assign n3274 = ( (~ Pg14705) ) | ( n3277 ) | ( (~ Ng6279) ) ;
 assign n3275 = ( n3269  &  n3266 ) | ( n1965  &  n3266 ) | ( n3269  &  n3281 ) | ( n1965  &  n3281 ) ;
 assign n3272 = ( n3273  &  n3274  &  n3275 ) ;
 assign n3278 = ( (~ Pg17760)  &  n5604 ) | ( n1965  &  n5604 ) | ( (~ Ng6291)  &  n5604 ) ;
 assign n3277 = ( Ng6395 ) | ( (~ Ng6336) ) ;
 assign n3276 = ( (~ Pg17649)  &  n3278 ) | ( n3278  &  n3277 ) | ( n3278  &  (~ Ng6307) ) ;
 assign n3282 = ( (~ Pg14779)  &  n5603 ) | ( n3277  &  n5603 ) | ( (~ Ng6267)  &  n5603 ) ;
 assign n3281 = ( Ng6336 ) | ( Ng6395 ) ;
 assign n3279 = ( (~ Pg17649)  &  n3282 ) | ( n3282  &  n3281 ) | ( n3282  &  (~ Ng6299) ) ;
 assign n3286 = ( n3262  &  n3272 ) | ( n3272  &  Ng6381 ) | ( n3262  &  (~ Ng6381) ) ;
 assign n3287 = ( n3276  &  n3279 ) | ( n3279  &  n5894 ) | ( n3276  &  (~ n5894) ) ;
 assign n3285 = ( (~ Pg17685) ) | ( n3263 ) | ( (~ Ng6381) ) ;
 assign n3283 = ( n3286  &  n3287  &  n3285 ) | ( n3286  &  n3287  &  (~ Ng6311) ) ;
 assign n3289 = ( Pg35 ) | ( (~ Ng6159) ) ;
 assign n3288 = ( (~ Pg35) ) | ( (~ n1196) ) | ( n3283 ) ;
 assign n3292 = ( (~ Ng5849) ) | ( (~ n4887) ) | ( (~ n4901) ) ;
 assign n3291 = ( (~ Ng5869) ) | ( n4590 ) ;
 assign n3294 = ( n3295  &  n4999 ) | ( n3295  &  Ng5835 ) | ( n4999  &  (~ Ng5835) ) ;
 assign n3296 = ( Ng5821 ) | ( n4999 ) | ( Ng5827 ) ;
 assign n3295 = ( (~ Pg35) ) | ( (~ n4998) ) ;
 assign n3300 = ( Ng5808 ) | ( n4999 ) | ( (~ Ng5813) ) ;
 assign n3302 = ( (~ Pg13068)  &  (~ Ng5913) ) | ( (~ Ng5913)  &  (~ Ng5901) ) | ( (~ Pg13068)  &  (~ Ng6031) ) | ( (~ Ng5901)  &  (~ Ng6031) ) ;
 assign n3306 = ( (~ Pg17715)  &  (~ Pg17646) ) | ( (~ Pg17646)  &  (~ Ng5957) ) | ( (~ Pg17715)  &  (~ Ng5905) ) | ( (~ Ng5957)  &  (~ Ng5905) ) ;
 assign n3310 = ( (~ Pg17819)  &  (~ Pg12350) ) | ( (~ Pg12350)  &  (~ Ng5925) ) | ( (~ Pg17819)  &  (~ Ng5909) ) | ( (~ Ng5925)  &  (~ Ng5909) ) ;
 assign n3317 = ( (~ Pg14673) ) | ( n3331 ) | ( (~ Ng5941) ) ;
 assign n3318 = ( n3306  &  n3302 ) | ( n1974  &  n3302 ) | ( n3306  &  n3335 ) | ( n1974  &  n3335 ) ;
 assign n3316 = ( (~ Ng6049) ) | ( (~ Ng5990) ) ;
 assign n3315 = ( n3317  &  n3318  &  n3310 ) | ( n3317  &  n3318  &  n3316 ) ;
 assign n3319 = ( (~ Pg13068)  &  (~ Ng5897) ) | ( (~ Ng5897)  &  (~ Ng5889) ) | ( (~ Pg13068)  &  (~ Ng6031) ) | ( (~ Ng5889)  &  (~ Ng6031) ) ;
 assign n3322 = ( (~ Pg17819)  &  (~ Pg12350) ) | ( (~ Pg12350)  &  (~ Ng5917) ) | ( (~ Pg17819)  &  (~ Ng5893) ) | ( (~ Ng5917)  &  (~ Ng5893) ) ;
 assign n3326 = ( (~ Pg14673) ) | ( n3335 ) | ( (~ Ng5933) ) ;
 assign n3327 = ( (~ Pg17715) ) | ( n3316 ) | ( (~ Ng5949) ) ;
 assign n3328 = ( n3322  &  n3319 ) | ( n1974  &  n3319 ) | ( n3322  &  n3331 ) | ( n1974  &  n3331 ) ;
 assign n3325 = ( n3326  &  n3327  &  n3328 ) ;
 assign n3333 = ( (~ Pg17739)  &  n5606 ) | ( n1974  &  n5606 ) | ( (~ Ng5945)  &  n5606 ) ;
 assign n3331 = ( Ng5990 ) | ( Ng6049 ) ;
 assign n3329 = ( (~ Pg14738)  &  n3333 ) | ( n3333  &  n3331 ) | ( n3333  &  (~ Ng5929) ) ;
 assign n3337 = ( (~ Pg17739)  &  n5605 ) | ( n3316  &  n5605 ) | ( (~ Ng5937)  &  n5605 ) ;
 assign n3335 = ( Ng6049 ) | ( (~ Ng5990) ) ;
 assign n3334 = ( (~ Pg14738)  &  n3337 ) | ( n3337  &  n3335 ) | ( n3337  &  (~ Ng5921) ) ;
 assign n3341 = ( n3315  &  n3325 ) | ( n3325  &  Ng6035 ) | ( n3315  &  (~ Ng6035) ) ;
 assign n3342 = ( n3329  &  n3334 ) | ( n3334  &  n5903 ) | ( n3329  &  (~ n5903) ) ;
 assign n3340 = ( (~ Pg17646) ) | ( n3316 ) | ( (~ Ng6035) ) ;
 assign n3338 = ( n3341  &  n3342  &  n3340 ) | ( n3341  &  n3342  &  (~ Ng5965) ) ;
 assign n3344 = ( Pg35 ) | ( (~ Ng5813) ) ;
 assign n3343 = ( (~ Pg35) ) | ( (~ n1179) ) | ( n3338 ) ;
 assign n3347 = ( (~ Ng5503) ) | ( (~ n4887) ) | ( (~ n4908) ) ;
 assign n3346 = ( (~ Ng5523) ) | ( n4587 ) ;
 assign n3349 = ( n3350  &  n5006 ) | ( n3350  &  Ng5489 ) | ( n5006  &  (~ Ng5489) ) ;
 assign n3351 = ( Ng5475 ) | ( n5006 ) | ( Ng5481 ) ;
 assign n3350 = ( (~ Pg35) ) | ( (~ n5005) ) ;
 assign n3355 = ( n5006 ) | ( (~ Ng5467) ) | ( Ng5462 ) ;
 assign n3357 = ( (~ Pg17678)  &  (~ Pg17604) ) | ( (~ Pg17604)  &  (~ Ng5611) ) | ( (~ Pg17678)  &  (~ Ng5559) ) | ( (~ Ng5611)  &  (~ Ng5559) ) ;
 assign n3361 = ( (~ Pg13049)  &  (~ Ng5567) ) | ( (~ Ng5567)  &  (~ Ng5555) ) | ( (~ Pg13049)  &  (~ Ng5685) ) | ( (~ Ng5555)  &  (~ Ng5685) ) ;
 assign n3365 = ( (~ Pg17813)  &  (~ Pg12300) ) | ( (~ Pg12300)  &  (~ Ng5579) ) | ( (~ Pg17813)  &  (~ Ng5563) ) | ( (~ Ng5579)  &  (~ Ng5563) ) ;
 assign n3372 = ( (~ Pg14635) ) | ( n3386 ) | ( (~ Ng5595) ) ;
 assign n3373 = ( n3361  &  n3357 ) | ( n3391  &  n3357 ) | ( n3361  &  n4783 ) | ( n3391  &  n4783 ) ;
 assign n3371 = ( (~ Ng5703) ) | ( (~ Ng5644) ) ;
 assign n3370 = ( n3372  &  n3373  &  n3365 ) | ( n3372  &  n3373  &  n3371 ) ;
 assign n3374 = ( (~ Pg17813)  &  (~ Pg12300) ) | ( (~ Pg12300)  &  (~ Ng5571) ) | ( (~ Pg17813)  &  (~ Ng5547) ) | ( (~ Ng5571)  &  (~ Ng5547) ) ;
 assign n3377 = ( (~ Pg13049)  &  (~ Ng5551) ) | ( (~ Ng5551)  &  (~ Ng5543) ) | ( (~ Pg13049)  &  (~ Ng5685) ) | ( (~ Ng5543)  &  (~ Ng5685) ) ;
 assign n3381 = ( (~ Pg17678) ) | ( n3371 ) | ( (~ Ng5603) ) ;
 assign n3382 = ( (~ Pg14635) ) | ( n3391 ) | ( (~ Ng5587) ) ;
 assign n3383 = ( n3377  &  n3374 ) | ( n3386  &  n3374 ) | ( n3377  &  n4783 ) | ( n3386  &  n4783 ) ;
 assign n3380 = ( n3381  &  n3382  &  n3383 ) ;
 assign n3388 = ( (~ Pg17711)  &  n5608 ) | ( n4783  &  n5608 ) | ( (~ Ng5599)  &  n5608 ) ;
 assign n3386 = ( Ng5644 ) | ( Ng5703 ) ;
 assign n3384 = ( (~ Pg14694)  &  n3388 ) | ( n3388  &  n3386 ) | ( n3388  &  (~ Ng5583) ) ;
 assign n3392 = ( (~ Pg17711)  &  n5607 ) | ( n3371  &  n5607 ) | ( (~ Ng5591)  &  n5607 ) ;
 assign n3391 = ( Ng5703 ) | ( (~ Ng5644) ) ;
 assign n3389 = ( (~ Pg14694)  &  n3392 ) | ( n3392  &  n3391 ) | ( n3392  &  (~ Ng5575) ) ;
 assign n3396 = ( n3370  &  n3380 ) | ( n3380  &  Ng5689 ) | ( n3370  &  (~ Ng5689) ) ;
 assign n3397 = ( n3384  &  n3389 ) | ( n3389  &  n5911 ) | ( n3384  &  (~ n5911) ) ;
 assign n3395 = ( (~ Pg17604) ) | ( n3371 ) | ( (~ Ng5689) ) ;
 assign n3393 = ( n3396  &  n3397  &  n3395 ) | ( n3396  &  n3397  &  (~ Ng5619) ) ;
 assign n3400 = ( Ng5462 ) | ( n3393 ) | ( n4784 ) ;
 assign n3402 = ( (~ Ng5156) ) | ( n4092 ) | ( (~ n4887) ) ;
 assign n3401 = ( (~ Ng5176) ) | ( n4595 ) ;
 assign n3404 = ( n3405  &  n5013 ) | ( n3405  &  Ng5142 ) | ( n5013  &  (~ Ng5142) ) ;
 assign n3406 = ( Ng5128 ) | ( n5013 ) | ( Ng5134 ) ;
 assign n3405 = ( (~ Pg35) ) | ( (~ n5012) ) ;
 assign n3410 = ( Ng5115 ) | ( n5013 ) | ( (~ Ng5120) ) ;
 assign n3412 = ( (~ Pg17787)  &  (~ Pg12238) ) | ( (~ Pg12238)  &  (~ Ng5232) ) | ( (~ Pg17787)  &  (~ Ng5216) ) | ( (~ Ng5232)  &  (~ Ng5216) ) ;
 assign n3417 = ( (~ Pg13039)  &  (~ Ng5220) ) | ( (~ Ng5220)  &  (~ Ng5208) ) | ( (~ Pg13039)  &  (~ Ng5339) ) | ( (~ Ng5208)  &  (~ Ng5339) ) ;
 assign n3421 = ( (~ Pg17639)  &  (~ Pg17577) ) | ( (~ Pg17577)  &  (~ Ng5264) ) | ( (~ Pg17639)  &  (~ Ng5212) ) | ( (~ Ng5264)  &  (~ Ng5212) ) ;
 assign n3426 = ( (~ Pg14597) ) | ( n3440 ) | ( (~ Ng5248) ) ;
 assign n3427 = ( n3417  &  n3412 ) | ( n3444  &  n3412 ) | ( n3417  &  n4527 ) | ( n3444  &  n4527 ) ;
 assign n3425 = ( n3426  &  n3427  &  n3421 ) | ( n3426  &  n3427  &  n1986 ) ;
 assign n3428 = ( (~ Pg17787)  &  (~ Pg12238) ) | ( (~ Pg12238)  &  (~ Ng5224) ) | ( (~ Pg17787)  &  (~ Ng5200) ) | ( (~ Ng5224)  &  (~ Ng5200) ) ;
 assign n3431 = ( (~ Pg13039)  &  (~ Ng5204) ) | ( (~ Ng5204)  &  (~ Ng5196) ) | ( (~ Pg13039)  &  (~ Ng5339) ) | ( (~ Ng5196)  &  (~ Ng5339) ) ;
 assign n3435 = ( (~ Pg14597) ) | ( n3444 ) | ( (~ Ng5240) ) ;
 assign n3436 = ( (~ Pg17639) ) | ( n4527 ) | ( (~ Ng5256) ) ;
 assign n3437 = ( n3431  &  n3428 ) | ( n3440  &  n3428 ) | ( n3431  &  n1986 ) | ( n3440  &  n1986 ) ;
 assign n3434 = ( n3435  &  n3436  &  n3437 ) ;
 assign n3442 = ( (~ Pg17519)  &  n5610 ) | ( n3444  &  n5610 ) | ( (~ Ng5268)  &  n5610 ) ;
 assign n3440 = ( Ng5297 ) | ( Ng5357 ) ;
 assign n3438 = ( (~ Pg14662)  &  n3442 ) | ( n3442  &  n3440 ) | ( n3442  &  (~ Ng5236) ) ;
 assign n3446 = ( (~ Pg17674)  &  n5609 ) | ( n4527  &  n5609 ) | ( (~ Ng5244)  &  n5609 ) ;
 assign n3444 = ( Ng5357 ) | ( (~ Ng5297) ) ;
 assign n3443 = ( (~ Pg14662)  &  n3446 ) | ( n3446  &  n3444 ) | ( n3446  &  (~ Ng5228) ) ;
 assign n3450 = ( (~ wire4415)  &  n3425 ) | ( wire4415  &  n3434 ) | ( n3425  &  n3434 ) ;
 assign n3451 = ( n3438  &  n3443 ) | ( n3443  &  n5919 ) | ( n3438  &  (~ n5919) ) ;
 assign n3447 = ( n3450  &  n3451  &  (~ Ng5272) ) | ( n3450  &  n3451  &  (~ n5011) ) ;
 assign n3453 = ( Pg35 ) | ( (~ Ng5120) ) ;
 assign n3452 = ( (~ Pg35) ) | ( (~ wire4394) ) | ( n3447 ) ;
 assign n3455 = ( n1136  &  n1118  &  Ng4927 ) | ( n1136  &  n1118  &  n1166 ) ;
 assign n3457 = ( (~ Ng4912) ) | ( Ng4899 ) | ( Ng4975 ) ;
 assign n3458 = ( n1118  &  n1166 ) | ( n1118  &  (~ Ng4917) ) | ( n1166  &  (~ Ng4922) ) | ( (~ Ng4917)  &  (~ Ng4922) ) ;
 assign n3456 = ( n1136  &  n3457  &  n3458 ) | ( n3457  &  n3458  &  (~ Ng4907) ) ;
 assign n3459 = ( (~ n1176)  &  (~ Ng4966)  &  (~ n5922) ) | ( (~ Ng4983)  &  (~ Ng4966)  &  (~ n5922) ) ;
 assign n3464 = ( n1180  &  n1099  &  Ng4737 ) | ( n1180  &  n1099  &  n1197 ) ;
 assign n3466 = ( (~ Ng4722) ) | ( Ng4709 ) | ( Ng4785 ) ;
 assign n3467 = ( n1099  &  n1197 ) | ( n1099  &  (~ Ng4727) ) | ( n1197  &  (~ Ng4717) ) | ( (~ Ng4727)  &  (~ Ng4717) ) ;
 assign n3465 = ( n1180  &  n3466  &  n3467 ) | ( n3466  &  n3467  &  (~ Ng4732) ) ;
 assign n3468 = ( (~ n1195)  &  (~ Ng4776)  &  (~ n5924) ) | ( (~ Ng4793)  &  (~ Ng4776)  &  (~ n5924) ) ;
 assign n3473 = ( (~ n4361)  &  Ng4087 ) | ( n4361  &  (~ Ng4087) ) ;
 assign n3474 = ( (~ Pg35) ) | ( (~ Ng2841) ) ;
 assign n3477 = ( (~ Ng3849) ) | ( (~ n4887) ) | ( (~ n4922) ) ;
 assign n3476 = ( (~ Ng3869) ) | ( n4584 ) ;
 assign n3479 = ( n3480  &  n5024 ) | ( n3480  &  Ng3835 ) | ( n5024  &  (~ Ng3835) ) ;
 assign n3481 = ( Ng3821 ) | ( n5024 ) | ( Ng3827 ) ;
 assign n3480 = ( (~ Pg35) ) | ( (~ n5023) ) ;
 assign n3485 = ( Ng3808 ) | ( n5024 ) | ( (~ Ng3813) ) ;
 assign n3487 = ( (~ Pg14518)  &  (~ Ng3913) ) | ( (~ Ng3913)  &  (~ Ng3901) ) | ( (~ Pg14518)  &  (~ Ng4031) ) | ( (~ Ng3901)  &  (~ Ng4031) ) ;
 assign n3491 = ( (~ Pg16748)  &  (~ Pg16693) ) | ( (~ Pg16693)  &  (~ Ng3957) ) | ( (~ Pg16748)  &  (~ Ng3905) ) | ( (~ Ng3957)  &  (~ Ng3905) ) ;
 assign n3495 = ( (~ Pg16955)  &  (~ Pg11418) ) | ( (~ Pg11418)  &  (~ Ng3925) ) | ( (~ Pg16955)  &  (~ Ng3909) ) | ( (~ Ng3925)  &  (~ Ng3909) ) ;
 assign n3502 = ( (~ Pg13906) ) | ( n3516 ) | ( (~ Ng3941) ) ;
 assign n3503 = ( n3491  &  n3487 ) | ( n1998  &  n3487 ) | ( n3491  &  n3520 ) | ( n1998  &  n3520 ) ;
 assign n3501 = ( (~ Ng4054) ) | ( (~ Ng3990) ) ;
 assign n3500 = ( n3502  &  n3503  &  n3495 ) | ( n3502  &  n3503  &  n3501 ) ;
 assign n3504 = ( (~ Pg16955)  &  (~ Pg11418) ) | ( (~ Pg11418)  &  (~ Ng3917) ) | ( (~ Pg16955)  &  (~ Ng3893) ) | ( (~ Ng3917)  &  (~ Ng3893) ) ;
 assign n3507 = ( (~ Pg14518)  &  (~ Ng3897) ) | ( (~ Ng3897)  &  (~ Ng3889) ) | ( (~ Pg14518)  &  (~ Ng4031) ) | ( (~ Ng3889)  &  (~ Ng4031) ) ;
 assign n3511 = ( (~ Pg16748) ) | ( n3501 ) | ( (~ Ng3949) ) ;
 assign n3512 = ( (~ Pg13906) ) | ( n3520 ) | ( (~ Ng3933) ) ;
 assign n3513 = ( n3507  &  n3504 ) | ( n3516  &  n3504 ) | ( n3507  &  n1998 ) | ( n3516  &  n1998 ) ;
 assign n3510 = ( n3511  &  n3512  &  n3513 ) ;
 assign n3518 = ( (~ Pg16659)  &  n5616 ) | ( n3520  &  n5616 ) | ( (~ Ng3961)  &  n5616 ) ;
 assign n3516 = ( Ng3990 ) | ( Ng4054 ) ;
 assign n3514 = ( (~ Pg13966)  &  n3518 ) | ( n3518  &  n3516 ) | ( n3518  &  (~ Ng3929) ) ;
 assign n3522 = ( (~ Pg16775)  &  n5615 ) | ( n3501  &  n5615 ) | ( (~ Ng3937)  &  n5615 ) ;
 assign n3520 = ( Ng4054 ) | ( (~ Ng3990) ) ;
 assign n3519 = ( (~ Pg13966)  &  n3522 ) | ( n3522  &  n3520 ) | ( n3522  &  (~ Ng3921) ) ;
 assign n3526 = ( n3500  &  n3510 ) | ( n3510  &  Ng4040 ) | ( n3500  &  (~ Ng4040) ) ;
 assign n3527 = ( n3514  &  n3519 ) | ( n3519  &  n5931 ) | ( n3514  &  (~ n5931) ) ;
 assign n3525 = ( (~ Pg16693) ) | ( n3501 ) | ( (~ Ng4040) ) ;
 assign n3523 = ( n3526  &  n3527  &  n3525 ) | ( n3526  &  n3527  &  (~ Ng3965) ) ;
 assign n3529 = ( Pg35 ) | ( (~ Ng3813) ) ;
 assign n3528 = ( (~ Pg35) ) | ( (~ n1165) ) | ( n3523 ) ;
 assign n3532 = ( (~ Ng3498) ) | ( (~ n4887) ) | ( (~ n4928) ) ;
 assign n3531 = ( (~ Ng3518) ) | ( n4593 ) ;
 assign n3534 = ( n3535  &  n5031 ) | ( n3535  &  Ng3484 ) | ( n5031  &  (~ Ng3484) ) ;
 assign n3536 = ( Ng3470 ) | ( n5031 ) | ( Ng3476 ) ;
 assign n3535 = ( (~ Pg35) ) | ( (~ n5030) ) ;
 assign n3539 = ( Ng3457 ) | ( n5031 ) | ( (~ Ng3462) ) ;
 assign n3541 = ( (~ Pg16924)  &  (~ Pg11388) ) | ( (~ Pg11388)  &  (~ Ng3574) ) | ( (~ Pg16924)  &  (~ Ng3558) ) | ( (~ Ng3574)  &  (~ Ng3558) ) ;
 assign n3546 = ( (~ Pg14451)  &  (~ Ng3562) ) | ( (~ Ng3562)  &  (~ Ng3550) ) | ( (~ Pg14451)  &  (~ Ng3680) ) | ( (~ Ng3550)  &  (~ Ng3680) ) ;
 assign n3550 = ( (~ Pg16722)  &  (~ Pg16656) ) | ( (~ Pg16656)  &  (~ Ng3606) ) | ( (~ Pg16722)  &  (~ Ng3554) ) | ( (~ Ng3606)  &  (~ Ng3554) ) ;
 assign n3555 = ( (~ Pg13881) ) | ( n5034 ) | ( (~ Ng3590) ) ;
 assign n3556 = ( n3546  &  n3541 ) | ( n4792  &  n3541 ) | ( n3546  &  n3572 ) | ( n4792  &  n3572 ) ;
 assign n3554 = ( n3555  &  n3556  &  n3550 ) | ( n3555  &  n3556  &  n2007 ) ;
 assign n3557 = ( (~ Pg14451)  &  (~ Ng3546) ) | ( (~ Ng3546)  &  (~ Ng3538) ) | ( (~ Pg14451)  &  (~ Ng3680) ) | ( (~ Ng3538)  &  (~ Ng3680) ) ;
 assign n3560 = ( (~ Pg16924)  &  (~ Pg11388) ) | ( (~ Pg11388)  &  (~ Ng3566) ) | ( (~ Pg16924)  &  (~ Ng3542) ) | ( (~ Ng3566)  &  (~ Ng3542) ) ;
 assign n3564 = ( (~ Pg13881) ) | ( n4792 ) | ( (~ Ng3582) ) ;
 assign n3565 = ( (~ Pg16722) ) | ( n3572 ) | ( (~ Ng3598) ) ;
 assign n3566 = ( n3560  &  n3557 ) | ( n2007  &  n3557 ) | ( n3560  &  n5034 ) | ( n2007  &  n5034 ) ;
 assign n3563 = ( n3564  &  n3565  &  n3566 ) ;
 assign n3570 = ( (~ Pg16627)  &  n5618 ) | ( n4792  &  n5618 ) | ( (~ Ng3610)  &  n5618 ) ;
 assign n3567 = ( (~ Pg16744)  &  n3570 ) | ( n2007  &  n3570 ) | ( n3570  &  (~ Ng3594) ) ;
 assign n3574 = ( (~ Pg13926)  &  n5617 ) | ( n4792  &  n5617 ) | ( (~ Ng3570)  &  n5617 ) ;
 assign n3572 = ( (~ Ng3703) ) | ( (~ Ng3639) ) ;
 assign n3571 = ( (~ Pg16744)  &  n3574 ) | ( n3574  &  n3572 ) | ( n3574  &  (~ Ng3586) ) ;
 assign n3578 = ( n3554  &  n3563 ) | ( n3563  &  Ng3689 ) | ( n3554  &  (~ Ng3689) ) ;
 assign n3579 = ( n3567  &  n3571 ) | ( n3571  &  n5939 ) | ( n3567  &  (~ n5939) ) ;
 assign n3577 = ( (~ Pg16656) ) | ( n3572 ) | ( (~ Ng3689) ) ;
 assign n3575 = ( n3578  &  n3579  &  n3577 ) | ( n3578  &  n3579  &  (~ Ng3614) ) ;
 assign n3581 = ( Pg35 ) | ( (~ Ng3462) ) ;
 assign n3580 = ( (~ Pg35) ) | ( (~ n1116) ) | ( n3575 ) ;
 assign n3584 = ( (~ Ng3147) ) | ( (~ n4887) ) | ( (~ n4934) ) ;
 assign n3583 = ( (~ Ng3167) ) | ( n4577 ) ;
 assign n3585 = ( n3586  &  n5039 ) | ( n3586  &  Ng3133 ) | ( n5039  &  (~ Ng3133) ) ;
 assign n3587 = ( Ng3119 ) | ( n5039 ) | ( Ng3125 ) ;
 assign n3586 = ( (~ Pg35) ) | ( (~ n5038) ) ;
 assign n3591 = ( n5039 ) | ( (~ Ng3111) ) | ( Ng3106 ) ;
 assign n3593 = ( (~ Pg16686)  &  (~ Pg16624) ) | ( (~ Pg16624)  &  (~ Ng3255) ) | ( (~ Pg16686)  &  (~ Ng3203) ) | ( (~ Ng3255)  &  (~ Ng3203) ) ;
 assign n3597 = ( (~ Pg16874)  &  (~ Pg11349) ) | ( (~ Pg11349)  &  (~ Ng3223) ) | ( (~ Pg16874)  &  (~ Ng3207) ) | ( (~ Ng3223)  &  (~ Ng3207) ) ;
 assign n3602 = ( (~ Pg14421)  &  (~ Ng3211) ) | ( (~ Ng3211)  &  (~ Ng3199) ) | ( (~ Pg14421)  &  (~ Ng3329) ) | ( (~ Ng3199)  &  (~ Ng3329) ) ;
 assign n3608 = ( (~ Pg13865) ) | ( n3624 ) | ( (~ Ng3239) ) ;
 assign n3609 = ( n3597  &  n3593 ) | ( n4516  &  n3593 ) | ( n3597  &  n2016 ) | ( n4516  &  n2016 ) ;
 assign n3607 = ( Ng3352 ) | ( (~ Ng3288) ) ;
 assign n3606 = ( n3608  &  n3609  &  n3602 ) | ( n3608  &  n3609  &  n3607 ) ;
 assign n3610 = ( (~ Pg16874)  &  (~ Pg11349) ) | ( (~ Pg11349)  &  (~ Ng3215) ) | ( (~ Pg16874)  &  (~ Ng3191) ) | ( (~ Ng3215)  &  (~ Ng3191) ) ;
 assign n3613 = ( (~ Pg14421)  &  (~ Ng3195) ) | ( (~ Ng3195)  &  (~ Ng3187) ) | ( (~ Pg14421)  &  (~ Ng3329) ) | ( (~ Ng3187)  &  (~ Ng3329) ) ;
 assign n3617 = ( (~ Pg16686) ) | ( n4516 ) | ( (~ Ng3247) ) ;
 assign n3618 = ( (~ Pg13865) ) | ( n3607 ) | ( (~ Ng3231) ) ;
 assign n3619 = ( n3613  &  n3610 ) | ( n3624  &  n3610 ) | ( n3613  &  n2016 ) | ( n3624  &  n2016 ) ;
 assign n3616 = ( n3617  &  n3618  &  n3619 ) ;
 assign n3621 = ( (~ Pg16718)  &  n5620 ) | ( n2016  &  n5620 ) | ( (~ Ng3243)  &  n5620 ) ;
 assign n3620 = ( (~ Pg16603)  &  n3621 ) | ( n3607  &  n3621 ) | ( n3621  &  (~ Ng3259) ) ;
 assign n3625 = ( (~ Pg13895)  &  n5619 ) | ( n3607  &  n5619 ) | ( (~ Ng3219)  &  n5619 ) ;
 assign n3624 = ( Ng3288 ) | ( Ng3352 ) ;
 assign n3622 = ( (~ Pg16603)  &  n3625 ) | ( n3625  &  n3624 ) | ( n3625  &  (~ Ng3251) ) ;
 assign n3629 = ( n3606  &  n3616 ) | ( n3616  &  Ng3338 ) | ( n3606  &  (~ Ng3338) ) ;
 assign n3630 = ( n3620  &  n3622 ) | ( n3622  &  n5947 ) | ( n3620  &  (~ n5947) ) ;
 assign n3628 = ( (~ Pg16624) ) | ( n4516 ) | ( (~ Ng3338) ) ;
 assign n3626 = ( n3629  &  n3630  &  n3628 ) | ( n3629  &  n3630  &  (~ Ng3263) ) ;
 assign n3633 = ( Ng3106 ) | ( n3626 ) | ( n4793 ) ;
 assign n3635 = ( (~ Pg35)  &  n5951 ) | ( (~ Ng2735)  &  n5951 ) | ( (~ n3634)  &  n5951 ) ;
 assign n3634 = ( (~ Ng2729) ) | ( n4690 ) ;
 assign n3636 = ( n1153  &  (~ n3640) ) | ( n1153  &  (~ n4947) ) ;
 assign n3640 = ( (~ Ng2638) ) | ( (~ Ng2652) ) | ( (~ n4947) ) ;
 assign n3639 = ( (~ Pg35)  &  Ng2638 ) | ( n1153  &  Ng2638  &  n3640 ) ;
 assign n3642 = ( (~ Ng2619)  &  (~ Ng2579) ) | ( (~ Ng2571)  &  (~ Ng2579) ) | ( (~ Ng2619)  &  (~ Ng2587) ) | ( (~ Ng2571)  &  (~ Ng2587) ) ;
 assign n3647 = ( Ng2619 ) | ( (~ Ng2575) ) | ( Ng2587 ) ;
 assign n3648 = ( n4550  &  (~ Ng2563) ) | ( (~ Ng2583)  &  (~ Ng2563) ) | ( n4550  &  n4947 ) | ( (~ Ng2583)  &  n4947 ) ;
 assign n3646 = ( n3647  &  n3648  &  Ng2610 ) | ( n3647  &  n3648  &  n3642 ) ;
 assign n3651 = ( n2361 ) | ( (~ Ng2638) ) ;
 assign n3652 = ( Pg35  &  n3646 ) | ( n3646  &  (~ Ng2619) ) | ( Pg35  &  n4860 ) | ( (~ Ng2619)  &  n4860 ) ;
 assign n3653 = ( n1151  &  (~ n3657) ) | ( n1151  &  (~ n4951) ) ;
 assign n3657 = ( (~ Ng2504) ) | ( (~ Ng2518) ) | ( (~ n4951) ) ;
 assign n3656 = ( (~ Pg35)  &  Ng2504 ) | ( n1151  &  Ng2504  &  n3657 ) ;
 assign n3659 = ( (~ Ng2485)  &  (~ Ng2445) ) | ( (~ Ng2437)  &  (~ Ng2445) ) | ( (~ Ng2485)  &  (~ Ng2453) ) | ( (~ Ng2437)  &  (~ Ng2453) ) ;
 assign n3664 = ( Ng2485 ) | ( (~ Ng2441) ) | ( Ng2453 ) ;
 assign n3665 = ( n4546  &  (~ Ng2429) ) | ( (~ Ng2449)  &  (~ Ng2429) ) | ( n4546  &  n4951 ) | ( (~ Ng2449)  &  n4951 ) ;
 assign n3663 = ( n3664  &  n3665  &  Ng2476 ) | ( n3664  &  n3665  &  n3659 ) ;
 assign n3668 = ( n2374 ) | ( (~ Ng2504) ) ;
 assign n3669 = ( Pg35  &  n3663 ) | ( n3663  &  (~ Ng2485) ) | ( Pg35  &  n4864 ) | ( (~ Ng2485)  &  n4864 ) ;
 assign n3672 = ( n4954  &  Ng2384  &  Ng2370 ) ;
 assign n3670 = ( n1162  &  n3672 ) | ( n1162  &  (~ n4954) ) ;
 assign n3673 = ( (~ Pg35)  &  Ng2370 ) | ( n1162  &  (~ n3672)  &  Ng2370 ) ;
 assign n3676 = ( (~ Ng2351)  &  (~ Ng2311) ) | ( (~ Ng2303)  &  (~ Ng2311) ) | ( (~ Ng2351)  &  (~ Ng2319) ) | ( (~ Ng2303)  &  (~ Ng2319) ) ;
 assign n3681 = ( Ng2351 ) | ( (~ Ng2307) ) | ( Ng2319 ) ;
 assign n3682 = ( n4548  &  (~ Ng2295) ) | ( (~ Ng2315)  &  (~ Ng2295) ) | ( n4548  &  n4954 ) | ( (~ Ng2315)  &  n4954 ) ;
 assign n3680 = ( n3681  &  n3682  &  Ng2342 ) | ( n3681  &  n3682  &  n3676 ) ;
 assign n3685 = ( n2388 ) | ( (~ Ng2370) ) ;
 assign n3686 = ( Pg35  &  n3680 ) | ( n3680  &  (~ Ng2351) ) | ( Pg35  &  n4866 ) | ( (~ Ng2351)  &  n4866 ) ;
 assign n3689 = ( n4957  &  Ng2250  &  Ng2236 ) ;
 assign n3687 = ( n1104  &  n3689 ) | ( n1104  &  (~ n4957) ) ;
 assign n3690 = ( (~ Pg35)  &  Ng2236 ) | ( n1104  &  (~ n3689)  &  Ng2236 ) ;
 assign n3693 = ( (~ Ng2217)  &  (~ Ng2177) ) | ( (~ Ng2169)  &  (~ Ng2177) ) | ( (~ Ng2217)  &  (~ Ng2185) ) | ( (~ Ng2169)  &  (~ Ng2185) ) ;
 assign n3698 = ( Ng2217 ) | ( (~ Ng2173) ) | ( Ng2185 ) ;
 assign n3699 = ( n4535  &  (~ Ng2161) ) | ( (~ Ng2181)  &  (~ Ng2161) ) | ( n4535  &  n4957 ) | ( (~ Ng2181)  &  n4957 ) ;
 assign n3697 = ( n3698  &  n3699  &  Ng2208 ) | ( n3698  &  n3699  &  n3693 ) ;
 assign n3702 = ( n2401 ) | ( (~ Ng2236) ) ;
 assign n3703 = ( Pg35  &  n3697 ) | ( n3697  &  (~ Ng2217) ) | ( Pg35  &  n4870 ) | ( (~ Ng2217)  &  n4870 ) ;
 assign n3706 = ( n4961  &  Ng2093  &  Ng2079 ) ;
 assign n3704 = ( n1146  &  n3706 ) | ( n1146  &  (~ n4961) ) ;
 assign n3707 = ( (~ Pg35)  &  Ng2079 ) | ( n1146  &  (~ n3706)  &  Ng2079 ) ;
 assign n3710 = ( (~ Ng2060)  &  (~ Ng2020) ) | ( (~ Ng2012)  &  (~ Ng2020) ) | ( (~ Ng2060)  &  (~ Ng2028) ) | ( (~ Ng2012)  &  (~ Ng2028) ) ;
 assign n3715 = ( Ng2060 ) | ( (~ Ng2016) ) | ( Ng2028 ) ;
 assign n3716 = ( n4542  &  (~ Ng2004) ) | ( (~ Ng2024)  &  (~ Ng2004) ) | ( n4542  &  n4961 ) | ( (~ Ng2024)  &  n4961 ) ;
 assign n3714 = ( n3715  &  n3716  &  Ng2051 ) | ( n3715  &  n3716  &  n3710 ) ;
 assign n3719 = ( n2414 ) | ( (~ Ng2079) ) ;
 assign n3720 = ( Pg35  &  n3714 ) | ( n3714  &  (~ Ng2060) ) | ( Pg35  &  n4873 ) | ( (~ Ng2060)  &  n4873 ) ;
 assign n3723 = ( n4964  &  Ng1959  &  Ng1945 ) ;
 assign n3721 = ( n1126  &  n3723 ) | ( n1126  &  (~ n4964) ) ;
 assign n3724 = ( (~ Pg35)  &  Ng1945 ) | ( n1126  &  (~ n3723)  &  Ng1945 ) ;
 assign n3727 = ( (~ Ng1926)  &  (~ Ng1886) ) | ( (~ Ng1878)  &  (~ Ng1886) ) | ( (~ Ng1926)  &  (~ Ng1894) ) | ( (~ Ng1878)  &  (~ Ng1894) ) ;
 assign n3732 = ( Ng1926 ) | ( (~ Ng1882) ) | ( Ng1894 ) ;
 assign n3733 = ( n4544  &  (~ Ng1870) ) | ( (~ Ng1890)  &  (~ Ng1870) ) | ( n4544  &  n4964 ) | ( (~ Ng1890)  &  n4964 ) ;
 assign n3731 = ( n3732  &  n3733  &  Ng1917 ) | ( n3732  &  n3733  &  n3727 ) ;
 assign n3736 = ( n2428 ) | ( (~ Ng1945) ) ;
 assign n3737 = ( Pg35  &  n3731 ) | ( n3731  &  (~ Ng1926) ) | ( Pg35  &  n4875 ) | ( (~ Ng1926)  &  n4875 ) ;
 assign n3738 = ( n1182  &  (~ n3742) ) | ( n1182  &  (~ n4967) ) ;
 assign n3742 = ( (~ Ng1811) ) | ( (~ Ng1825) ) | ( (~ n4967) ) ;
 assign n3741 = ( (~ Pg35)  &  Ng1811 ) | ( n1182  &  Ng1811  &  n3742 ) ;
 assign n3744 = ( (~ Ng1792)  &  (~ Ng1752) ) | ( (~ Ng1744)  &  (~ Ng1752) ) | ( (~ Ng1792)  &  (~ Ng1760) ) | ( (~ Ng1744)  &  (~ Ng1760) ) ;
 assign n3749 = ( Ng1792 ) | ( (~ Ng1748) ) | ( Ng1760 ) ;
 assign n3750 = ( n4538  &  (~ Ng1736) ) | ( (~ Ng1756)  &  (~ Ng1736) ) | ( n4538  &  n4967 ) | ( (~ Ng1756)  &  n4967 ) ;
 assign n3748 = ( n3749  &  n3750  &  Ng1783 ) | ( n3749  &  n3750  &  n3744 ) ;
 assign n3753 = ( n2441 ) | ( (~ Ng1811) ) ;
 assign n3754 = ( Pg35  &  n3748 ) | ( n3748  &  (~ Ng1792) ) | ( Pg35  &  n4878 ) | ( (~ Ng1792)  &  n4878 ) ;
 assign n3755 = ( n1087  &  (~ n3759) ) | ( n1087  &  (~ n4970) ) ;
 assign n3759 = ( (~ Ng1677) ) | ( (~ Ng1691) ) | ( (~ n4970) ) ;
 assign n3758 = ( (~ Pg35)  &  Ng1677 ) | ( n1087  &  Ng1677  &  n3759 ) ;
 assign n3761 = ( (~ Ng1657)  &  (~ Ng1616) ) | ( (~ Ng1608)  &  (~ Ng1616) ) | ( (~ Ng1657)  &  (~ Ng1624) ) | ( (~ Ng1608)  &  (~ Ng1624) ) ;
 assign n3766 = ( Ng1657 ) | ( (~ Ng1612) ) | ( Ng1624 ) ;
 assign n3767 = ( n4553  &  (~ Ng1600) ) | ( (~ Ng1620)  &  (~ Ng1600) ) | ( n4553  &  n4970 ) | ( (~ Ng1620)  &  n4970 ) ;
 assign n3765 = ( n3766  &  n3767  &  Ng1648 ) | ( n3766  &  n3767  &  n3761 ) ;
 assign n3770 = ( n2454 ) | ( (~ Ng1677) ) ;
 assign n3771 = ( Pg35  &  n3765 ) | ( n3765  &  (~ Ng1657) ) | ( Pg35  &  n4881 ) | ( (~ Ng1657)  &  n4881 ) ;
 assign n3774 = ( (~ Pg35)  &  (~ Ng1472) ) | ( Pg35  &  (~ n5356) ) | ( (~ Ng1472)  &  (~ n5356) ) ;
 assign n3772 = ( (~ Pg35) ) | ( n715 ) ;
 assign n3776 = ( (~ Ng1256) ) | ( n4222 ) | ( n4810 ) ;
 assign n3777 = ( Pg35 ) | ( (~ Ng1252) ) ;
 assign n3780 = ( (~ Pg35)  &  (~ Ng1129) ) | ( Pg35  &  (~ n5361) ) | ( (~ Ng1129)  &  (~ n5361) ) ;
 assign n3778 = ( (~ Pg35) ) | ( n557 ) ;
 assign n3782 = ( (~ Ng911) ) | ( n4235 ) | ( n4823 ) ;
 assign n3783 = ( Pg35 ) | ( (~ Ng907) ) ;
 assign n3786 = ( (~ Ng847) ) | ( (~ Ng812) ) ;
 assign n3784 = ( Ng837  &  n3786 ) | ( n3786  &  (~ Ng847) ) ;
 assign n3788 = ( (~ n3784) ) | ( (~ n5978) ) | ( Ng723 ) ;
 assign n3789 = ( n4037 ) | ( n5978 ) | ( (~ Ng723) ) ;
 assign n3790 = ( n1369  &  Ng739 ) | ( (~ n1369)  &  (~ Ng739) ) ;
 assign n3791 = ( (~ Pg35) ) | ( n4490 ) ;
 assign n3794 = ( (~ Ng699) ) | ( (~ Ng681) ) | ( n5051 ) | ( n5052 ) | ( Ng650 ) | ( Ng645 ) ;
 assign n3793 = ( Ng703  &  n3794 ) | ( Ng703  &  (~ n4363) ) ;
 assign n3797 = ( (~ n3793) ) | ( Ng714 ) | ( n5980 ) ;
 assign n3798 = ( n3803 ) | ( (~ Ng714) ) | ( (~ n5980) ) ;
 assign n3800 = ( (~ n3793) ) | ( Ng676 ) | ( (~ n5054) ) ;
 assign n3801 = ( n3803 ) | ( (~ Ng676) ) | ( n5054 ) ;
 assign n3802 = ( n4363  &  Ng671 ) | ( (~ n4363)  &  (~ Ng671) ) ;
 assign n3803 = ( (~ Pg35) ) | ( (~ n3793) ) ;
 assign n3806 = ( (~ Ng586) ) | ( (~ n3805) ) | ( n4508 ) ;
 assign n3807 = ( Pg35 ) | ( (~ Ng572) ) ;
 assign n3805 = ( (~ Ng572) ) | ( n3899 ) ;
 assign n3809 = ( (~ Pg35) ) | ( n5056 ) ;
 assign n3810 = ( (~ Pg35)  &  n5982 ) | ( (~ Ng490)  &  n5982 ) | ( n5058  &  n5982 ) ;
 assign n3813 = ( n5984 ) | ( n4259 ) | ( Ng417 ) ;
 assign n3812 = ( (~ Pg35) ) | ( (~ n4170) ) ;
 assign n3815 = ( n1960 ) | ( (~ Ng5011) ) ;
 assign n3816 = ( n1969 ) | ( (~ Ng4826) ) ;
 assign n3817 = ( n1978 ) | ( (~ Ng4831) ) ;
 assign n3818 = ( n3393  &  n3849 ) | ( n3849  &  n4784 ) | ( n3393  &  (~ Ng4821) ) | ( n4784  &  (~ Ng4821) ) ;
 assign n3819 = ( (~ wire4427) ) | ( n1990 ) ;
 assign n3821 = ( n1998  &  n3501 ) | ( n3501  &  Ng4049 ) | ( n1998  &  (~ Ng4049) ) ;
 assign n3822 = ( (~ Ng4045)  &  n3516 ) | ( Ng4045  &  n3520 ) | ( n3516  &  n3520 ) ;
 assign n3820 = ( (~ n1165)  &  (~ Ng4961) ) | ( n3821  &  n3822  &  (~ Ng4961) ) ;
 assign n3824 = ( n2002 ) | ( (~ Ng4961) ) ;
 assign n3823 = ( n4564 ) | ( n1118 ) ;
 assign n3826 = ( Ng3694  &  n4792 ) | ( (~ Ng3694)  &  n5034 ) | ( n4792  &  n5034 ) ;
 assign n3827 = ( n2007  &  n3572 ) | ( n3572  &  Ng3698 ) | ( n2007  &  (~ Ng3698) ) ;
 assign n3825 = ( (~ n1116)  &  (~ Ng4950) ) | ( n3826  &  n3827  &  (~ Ng4950) ) ;
 assign n3829 = ( n2011 ) | ( (~ Ng4950) ) ;
 assign n3828 = ( n4564 ) | ( n1136 ) ;
 assign n3830 = ( Ng4975 ) | ( Ng4899 ) | ( n4564 ) ;
 assign n3832 = ( (~ Pg35) ) | ( n1135 ) ;
 assign n3834 = ( (~ Ng6732)  &  n3223 ) | ( Ng6732  &  n3227 ) | ( n3223  &  n3227 ) ;
 assign n3835 = ( n1956  &  n3208 ) | ( n3208  &  Ng6736 ) | ( n1956  &  (~ Ng6736) ) ;
 assign n3833 = ( (~ n1109)  &  (~ Ng4894) ) | ( n3834  &  n3835  &  (~ Ng4894) ) ;
 assign n3836 = ( n1960 ) | ( (~ Ng4894) ) ;
 assign n3838 = ( Ng6386  &  n3277 ) | ( (~ Ng6386)  &  n3281 ) | ( n3277  &  n3281 ) ;
 assign n3839 = ( n1965  &  n3263 ) | ( n3263  &  Ng6390 ) | ( n1965  &  (~ Ng6390) ) ;
 assign n3837 = ( (~ n1196)  &  (~ Ng4771) ) | ( n3838  &  n3839  &  (~ Ng4771) ) ;
 assign n3841 = ( n1969 ) | ( (~ Ng4771) ) ;
 assign n3840 = ( n4559 ) | ( n1180 ) ;
 assign n3843 = ( (~ Ng6040)  &  n3331 ) | ( Ng6040  &  n3335 ) | ( n3331  &  n3335 ) ;
 assign n3844 = ( n1974  &  n3316 ) | ( n3316  &  Ng6044 ) | ( n1974  &  (~ Ng6044) ) ;
 assign n3842 = ( (~ n1179)  &  (~ Ng4760) ) | ( n3843  &  n3844  &  (~ Ng4760) ) ;
 assign n3846 = ( n1978 ) | ( (~ Ng4760) ) ;
 assign n3845 = ( n4559 ) | ( n1099 ) ;
 assign n3847 = ( Ng4785 ) | ( Ng4709 ) | ( n4559 ) ;
 assign n3849 = ( (~ Pg35) ) | ( n1097 ) ;
 assign n3851 = ( n1986  &  n4527 ) | ( n4527  &  Ng5352 ) | ( n1986  &  (~ Ng5352) ) ;
 assign n3852 = ( (~ Ng5348)  &  n3440 ) | ( Ng5348  &  n3444 ) | ( n3440  &  n3444 ) ;
 assign n3850 = ( (~ wire4394)  &  (~ Ng4704) ) | ( n3851  &  n3852  &  (~ Ng4704) ) ;
 assign n3854 = ( n1990 ) | ( (~ Ng4704) ) ;
 assign n3853 = ( n1197 ) | ( n4559 ) ;
 assign n3858 = ( Pg35  &  Ng4057 ) | ( Pg35  &  Ng4064 ) | ( Pg35  &  (~ n5068) ) ;
 assign n3861 = ( Pg35 ) | ( (~ Ng4119) ) ;
 assign n3862 = ( (~ Pg35) ) | ( (~ n3855) ) | ( (~ Ng4122) ) ;
 assign n3855 = ( n4786 ) | ( (~ n5068) ) ;
 assign n3860 = ( (~ Pg35) ) | ( (~ Ng4145) ) ;
 assign n3863 = ( Pg35 ) | ( (~ Ng4116) ) ;
 assign n3864 = ( (~ Pg35) ) | ( n5070 ) | ( (~ Ng4119) ) ;
 assign n3865 = ( Pg35 ) | ( (~ Ng4112) ) ;
 assign n3866 = ( (~ Pg35) ) | ( n5071 ) | ( (~ Ng4116) ) ;
 assign n3868 = ( (~ Pg35)  &  n5992 ) | ( (~ Ng4076)  &  n5992 ) | ( (~ n3867)  &  n5992 ) ;
 assign n3867 = ( (~ n4787) ) | ( (~ Ng4082) ) ;
 assign n3869 = ( n2002 ) | ( (~ Ng4035) ) ;
 assign n3870 = ( n2011 ) | ( (~ Ng3684) ) ;
 assign n3871 = ( n3626  &  n3832 ) | ( n3832  &  n4793 ) | ( n3626  &  (~ Ng3333) ) | ( n4793  &  (~ Ng3333) ) ;
 assign n3873 = ( Pg35 ) | ( (~ Ng2724) ) ;
 assign n3872 = ( (~ n4690)  &  Ng2729 ) | ( n4690  &  (~ Ng2729) ) ;
 assign n3876 = ( (~ Pg35)  &  n5993 ) | ( n2194  &  n5993 ) | ( (~ Ng1345)  &  n5993 ) ;
 assign n3875 = ( (~ Pg35) ) | ( (~ n4805) ) ;
 assign n3878 = ( (~ Ng1252) ) | ( (~ n3877) ) | ( n4222 ) ;
 assign n3879 = ( Pg35 ) | ( (~ Ng1280) ) ;
 assign n3877 = ( n4808 ) | ( (~ Ng1280) ) ;
 assign n3882 = ( (~ Pg35)  &  n5994 ) | ( n2207  &  n5994 ) | ( (~ Ng1002)  &  n5994 ) ;
 assign n3881 = ( (~ Pg35) ) | ( (~ n4818) ) ;
 assign n3884 = ( (~ Ng907) ) | ( (~ n3883) ) | ( n4235 ) ;
 assign n3885 = ( Pg35 ) | ( (~ Ng936) ) ;
 assign n3883 = ( n4821 ) | ( (~ Ng936) ) ;
 assign n3887 = ( (~ n3784) ) | ( Ng827 ) | ( n5049 ) ;
 assign n3888 = ( n4037 ) | ( (~ Ng827) ) | ( (~ n5049) ) ;
 assign n3890 = ( n3812 ) | ( (~ Ng699) ) ;
 assign n3891 = ( (~ Pg35) ) | ( n5075 ) ;
 assign n3893 = ( n3891  &  (~ Ng650) ) | ( (~ Ng681)  &  (~ Ng650) ) | ( n3891  &  (~ n5074) ) | ( (~ Ng681)  &  (~ n5074) ) ;
 assign n3894 = ( (~ Ng703)  &  (~ n4192) ) | ( Ng714  &  (~ n4192) ) ;
 assign n3900 = ( (~ Ng572) ) | ( (~ n3899) ) | ( n4508 ) ;
 assign n3901 = ( Pg35 ) | ( (~ Ng568) ) ;
 assign n3899 = ( (~ Ng568) ) | ( n4046 ) ;
 assign n3903 = ( Pg35 ) | ( (~ Ng528) ) ;
 assign n3902 = ( n1172  &  Ng482 ) | ( (~ n1172)  &  (~ Ng482) ) ;
 assign n3904 = ( (~ Pg35) ) | ( (~ n4657) ) ;
 assign n3907 = ( n1108 ) | ( n1112 ) ;
 assign n3906 = ( n3907  &  n1150 ) | ( n3907  &  n1108  &  n1112 ) ;
 assign n3911 = ( n1101  &  (~ n1131)  &  (~ n1133) ) ;
 assign n3914 = ( n1101  &  (~ n4567) ) | ( (~ n1131)  &  (~ n1133)  &  (~ n4567) ) ;
 assign n3915 = ( Ng4531  &  Ng4581 ) ;
 assign n3916 = ( Pg10306  &  Pg35 ) ;
 assign n3918 = ( (~ Pg35) ) | ( (~ Ng4515) ) | ( (~ Ng4521) ) ;
 assign n3923 = ( Ng4392 ) | ( Ng4417 ) | ( n3943 ) ;
 assign n3920 = ( (~ Pg35)  &  (~ Ng4392) ) | ( (~ Ng4392)  &  n3923 ) | ( (~ Pg35)  &  (~ n5081) ) | ( n3923  &  (~ n5081) ) ;
 assign n3926 = ( Ng4438 ) | ( Ng4443 ) | ( Ng4452 ) | ( Pg7245 ) | ( Pg7260 ) ;
 assign n3925 = ( Pg35  &  (~ Ng4392) ) | ( Pg35  &  n3926 ) ;
 assign n3929 = ( (~ Pg35) ) | ( Ng4392 ) ;
 assign n3933 = ( (~ Pg35) ) | ( (~ Ng4392) ) | ( n3926 ) ;
 assign n3934 = ( Pg35 ) | ( (~ Ng4443) ) ;
 assign n3935 = ( (~ Pg35) ) | ( Ng4382 ) | ( (~ Ng4438) ) ;
 assign n3937 = ( (~ Ng4401)  &  Ng4434 ) | ( Ng4401  &  (~ Ng4434) ) ;
 assign n3936 = ( Pg35  &  n3937 ) | ( Pg35  &  Ng4388  &  (~ Ng4430) ) ;
 assign n3940 = ( (~ Pg35) ) | ( (~ Ng4423) ) ;
 assign n3943 = ( Ng4405 ) | ( Ng4375 ) | ( Ng4411 ) | ( Pg7257 ) | ( Pg7243 ) ;
 assign n3942 = ( Pg35  &  (~ Ng4392) ) | ( Pg35  &  n3943 ) ;
 assign n3948 = ( (~ Ng4382) ) | ( (~ n5081) ) | ( Ng4375 ) ;
 assign n3949 = ( Ng4382 ) | ( (~ n5081) ) | ( (~ Ng4375) ) ;
 assign n3950 = ( Pg35  &  n3923 ) | ( (~ Pg35)  &  (~ Ng4388) ) | ( n3923  &  (~ Ng4388) ) ;
 assign n3952 = ( (~ Pg35) ) | ( (~ Ng4392) ) | ( n3943 ) ;
 assign n3953 = ( n3943 ) | ( n3929 ) ;
 assign n3955 = ( Pg35 ) | ( (~ Ng4141) ) ;
 assign n3954 = ( n4787  &  Ng4082 ) | ( (~ n4787)  &  (~ Ng4082) ) ;
 assign n3957 = ( (~ n1256)  &  (~ n1254) ) | ( (~ n1254)  &  (~ Ng2827) ) | ( (~ n1256)  &  Ng2595 ) | ( (~ Ng2827)  &  Ng2595 ) ;
 assign n3959 = ( (~ n1256)  &  (~ n1254) ) | ( (~ n1254)  &  (~ Ng2823) ) | ( (~ n1256)  &  Ng2461 ) | ( (~ Ng2823)  &  Ng2461 ) ;
 assign n3961 = ( (~ n1256)  &  (~ n1254) ) | ( (~ n1254)  &  (~ Ng2811) ) | ( (~ n1256)  &  Ng2327 ) | ( (~ Ng2811)  &  Ng2327 ) ;
 assign n3963 = ( (~ n1256)  &  (~ n1254) ) | ( (~ n1254)  &  (~ Ng2799) ) | ( (~ n1256)  &  Ng2193 ) | ( (~ Ng2799)  &  Ng2193 ) ;
 assign n3965 = ( (~ n1256)  &  (~ n1254) ) | ( (~ n1254)  &  (~ Ng2795) ) | ( (~ n1256)  &  Ng2036 ) | ( (~ Ng2795)  &  Ng2036 ) ;
 assign n3967 = ( (~ n1256)  &  (~ n1254) ) | ( (~ n1254)  &  (~ Ng2791) ) | ( (~ n1256)  &  Ng1902 ) | ( (~ Ng2791)  &  Ng1902 ) ;
 assign n3969 = ( (~ n1256)  &  (~ n1254) ) | ( (~ n1254)  &  (~ Ng2779) ) | ( (~ n1256)  &  Ng1768 ) | ( (~ Ng2779)  &  Ng1768 ) ;
 assign n3971 = ( (~ n1256)  &  (~ n1254) ) | ( (~ n1254)  &  (~ Ng2767) ) | ( (~ n1256)  &  Ng1632 ) | ( (~ Ng2767)  &  Ng1632 ) ;
 assign n3973 = ( n3046 ) | ( (~ Ng2724) ) | ( (~ n4689) ) ;
 assign n3974 = ( Ng2724 ) | ( n4689 ) | ( (~ Ng2841) ) ;
 assign n3976 = ( Pg35 ) | ( (~ Ng1437) ) ;
 assign n3977 = ( (~ Pg35) ) | ( (~ Ng1478) ) | ( n5084 ) ;
 assign n3979 = ( Pg35 ) | ( (~ Ng1467) ) ;
 assign n3980 = ( (~ Pg35) ) | ( (~ Ng1472) ) | ( n5085 ) ;
 assign n3983 = ( (~ Pg35) ) | ( (~ Ng1448) ) | ( n5086 ) ;
 assign n3984 = ( Pg12923  &  Pg7946 ) | ( Pg12923  &  Pg19357 ) | ( Pg12923  &  Ng1333 ) ;
 assign n3985 = ( Ng1395  &  n3984 ) ;
 assign n3986 = ( (~ n854)  &  Ng1384 ) | ( (~ n854)  &  (~ Ng1351) ) ;
 assign n3990 = ( (~ Pg35) ) | ( n3986 ) | ( (~ Ng1389) ) ;
 assign n3993 = ( Ng1280 ) | ( n4808 ) ;
 assign n3994 = ( n4222 ) | ( (~ n4808) ) | ( (~ Ng1280) ) ;
 assign n3996 = ( Pg35 ) | ( (~ Ng1094) ) ;
 assign n3997 = ( (~ Pg35) ) | ( (~ Ng1135) ) | ( n5090 ) ;
 assign n3999 = ( Pg35 ) | ( (~ Ng1124) ) ;
 assign n4000 = ( (~ Pg35) ) | ( (~ Ng1129) ) | ( n5091 ) ;
 assign n4003 = ( (~ Pg35) ) | ( (~ Ng1105) ) | ( n5092 ) ;
 assign n4004 = ( Pg12919  &  Pg7916 ) | ( Pg12919  &  Pg19334 ) | ( Pg12919  &  Ng990 ) ;
 assign n4005 = ( (~ Pg35)  &  (~ n4004) ) | ( (~ n4004)  &  (~ Ng1061) ) | ( (~ Pg35)  &  (~ Ng1052) ) | ( (~ Ng1061)  &  (~ Ng1052) ) ;
 assign n4010 = ( (~ n379)  &  (~ Ng1008) ) | ( (~ n379)  &  Ng1041 ) ;
 assign n4014 = ( (~ Pg35) ) | ( n4010 ) | ( (~ Ng1046) ) ;
 assign n4017 = ( Ng936 ) | ( n4821 ) ;
 assign n4018 = ( n4235 ) | ( (~ n4821) ) | ( (~ Ng936) ) ;
 assign n4019 = ( Pg35  &  (~ Ng890) ) ;
 assign n4021 = ( (~ Ng446)  &  n5096 ) | ( n5094  &  n5096 ) | ( (~ Ng446)  &  (~ Ng872) ) | ( n5094  &  (~ Ng872) ) ;
 assign n4023 = ( (~ Pg14167)  &  (~ Ng246) ) | ( (~ Pg14167)  &  n5094 ) | ( (~ Ng246)  &  n5096 ) | ( n5094  &  n5096 ) ;
 assign n4025 = ( (~ Pg14147)  &  (~ Ng269) ) | ( (~ Pg14147)  &  n5094 ) | ( (~ Ng269)  &  n5096 ) | ( n5094  &  n5096 ) ;
 assign n4027 = ( (~ Pg14125)  &  (~ Ng239) ) | ( (~ Pg14125)  &  n5094 ) | ( (~ Ng239)  &  n5096 ) | ( n5094  &  n5096 ) ;
 assign n4029 = ( (~ Pg14096)  &  (~ Ng262) ) | ( (~ Pg14096)  &  n5094 ) | ( (~ Ng262)  &  n5096 ) | ( n5094  &  n5096 ) ;
 assign n4031 = ( (~ Pg14217)  &  (~ Ng232) ) | ( (~ Pg14217)  &  n5094 ) | ( (~ Ng232)  &  n5096 ) | ( n5094  &  n5096 ) ;
 assign n4033 = ( (~ Pg14201)  &  (~ Ng255) ) | ( (~ Pg14201)  &  n5094 ) | ( (~ Ng255)  &  n5096 ) | ( n5094  &  n5096 ) ;
 assign n4035 = ( (~ Pg14189)  &  (~ Ng225) ) | ( (~ Pg14189)  &  n5094 ) | ( (~ Ng225)  &  n5096 ) | ( n5094  &  n5096 ) ;
 assign n4036 = ( (~ n4379)  &  Ng822 ) | ( n4379  &  (~ Ng822) ) ;
 assign n4037 = ( (~ Pg35) ) | ( (~ n3784) ) ;
 assign n4039 = ( Pg35  &  (~ Ng847) ) | ( Pg35  &  (~ Ng843) ) ;
 assign n4044 = ( (~ Pg35) ) | ( (~ wire4435) ) | ( n4363 ) ;
 assign n4047 = ( (~ Ng568) ) | ( (~ n4046) ) | ( n4508 ) ;
 assign n4048 = ( Pg35 ) | ( (~ Ng562) ) ;
 assign n4046 = ( (~ n1205) ) | ( (~ Ng562) ) | ( n4503 ) ;
 assign n4049 = ( (~ Pg35)  &  (~ Ng355) ) | ( Ng351  &  (~ Ng355)  &  (~ Ng333) ) ;
 assign n4052 = ( (~ wire4436)  &  (~ Ng351) ) ;
 assign n4055 = ( Ng311  &  (~ Ng305) ) | ( (~ Ng324)  &  (~ Ng305) ) ;
 assign n4059 = ( (~ Pg35) ) | ( (~ Ng336) ) | ( (~ n5109) ) ;
 assign n4060 = ( Pg35 ) | ( (~ Ng311) ) ;
 assign n4058 = ( (~ Pg35) ) | ( n5109 ) ;
 assign n4063 = ( Pg35  &  Ng329 ) | ( Pg35  &  n6013 ) | ( (~ Ng329)  &  n6013 ) ;
 assign n4061 = ( (~ Ng311)  &  (~ Ng305) ) | ( (~ Ng305)  &  Ng336 ) | ( (~ Ng311)  &  (~ Ng336) ) ;
 assign n4064 = ( (~ Ng311)  &  (~ Ng305) ) ;
 assign n4067 = ( (~ Ng6537)  &  n3184 ) | ( n3184  &  (~ n4886) ) | ( (~ Ng6537)  &  (~ n5409) ) | ( (~ n4886)  &  (~ n5409) ) ;
 assign n4070 = ( Pg35 ) | ( (~ Ng6509) ) ;
 assign n4071 = ( (~ Pg35) ) | ( n3184 ) | ( Ng6513 ) ;
 assign n4073 = ( (~ Ng6191)  &  n3238 ) | ( n3238  &  (~ n4894) ) | ( (~ Ng6191)  &  (~ n5417) ) | ( (~ n4894)  &  (~ n5417) ) ;
 assign n4076 = ( Pg35 ) | ( (~ Ng6163) ) ;
 assign n4077 = ( (~ Pg35) ) | ( n3238 ) | ( Ng6167 ) ;
 assign n4079 = ( (~ Ng5845)  &  n3291 ) | ( n3291  &  (~ n4901) ) | ( (~ Ng5845)  &  (~ n5425) ) | ( (~ n4901)  &  (~ n5425) ) ;
 assign n4082 = ( Pg35 ) | ( (~ Ng5817) ) ;
 assign n4083 = ( (~ Pg35) ) | ( n3291 ) | ( Ng5821 ) ;
 assign n4085 = ( (~ Ng5499)  &  n3346 ) | ( n3346  &  (~ n4908) ) | ( (~ Ng5499)  &  (~ n5433) ) | ( (~ n4908)  &  (~ n5433) ) ;
 assign n4088 = ( Pg35 ) | ( (~ Ng5471) ) ;
 assign n4089 = ( (~ Pg35) ) | ( n3346 ) | ( Ng5475 ) ;
 assign n4091 = ( (~ Ng5152)  &  n3401 ) | ( n3401  &  n4092 ) | ( (~ Ng5152)  &  (~ n5441) ) | ( n4092  &  (~ n5441) ) ;
 assign n4094 = ( Pg35 ) | ( (~ Ng5124) ) ;
 assign n4095 = ( (~ Pg35) ) | ( n3401 ) | ( Ng5128 ) ;
 assign n4092 = ( (~ Pg35) ) | ( (~ n3401) ) ;
 assign n4097 = ( Pg35 ) | ( (~ Ng5097) ) ;
 assign n4096 = ( (~ Ng5097) ) | ( (~ n5122) ) ;
 assign n4100 = ( Pg35 ) | ( (~ Ng5092) ) ;
 assign n4101 = ( (~ Pg35) ) | ( (~ Ng5097) ) | ( n5122 ) ;
 assign n4102 = ( Ng5092  &  Pg35 ) ;
 assign n4106 = ( (~ Pg35) ) | ( Ng5073 ) | ( (~ Ng5077) ) ;
 assign n4103 = ( Pg35  &  (~ Ng5084) ) ;
 assign n4110 = ( Ng4098  &  (~ Ng4093) ) ;
 assign n4107 = ( n1635  &  Ng4087  &  (~ Ng4057)  &  (~ Ng4064)  &  Ng4076  &  n4110 ) ;
 assign n4112 = ( n4786 ) | ( Ng4141 ) | ( (~ Ng2841) ) ;
 assign n4113 = ( n3474 ) | ( (~ n4786) ) | ( (~ Ng4141) ) ;
 assign n4115 = ( Pg35  &  Ng4064 ) | ( (~ Pg35)  &  (~ Ng4072) ) | ( Ng4064  &  (~ Ng4072) ) ;
 assign n4114 = ( n4115  &  n1994 ) ;
 assign n4117 = ( (~ Ng3845)  &  n3476 ) | ( n3476  &  (~ n4922) ) | ( (~ Ng3845)  &  (~ n5454) ) | ( (~ n4922)  &  (~ n5454) ) ;
 assign n4120 = ( Pg35 ) | ( (~ Ng3817) ) ;
 assign n4121 = ( (~ Pg35) ) | ( n3476 ) | ( Ng3821 ) ;
 assign n4123 = ( (~ Ng3494)  &  n3531 ) | ( n3531  &  (~ n4928) ) | ( (~ Ng3494)  &  (~ n5462) ) | ( (~ n4928)  &  (~ n5462) ) ;
 assign n4126 = ( Pg35 ) | ( (~ Ng3466) ) ;
 assign n4127 = ( (~ Pg35) ) | ( n3531 ) | ( Ng3470 ) ;
 assign n4129 = ( n3583  &  (~ n4934) ) | ( n3583  &  (~ Ng3143) ) | ( (~ n4934)  &  (~ n5470) ) | ( (~ Ng3143)  &  (~ n5470) ) ;
 assign n4132 = ( Pg35 ) | ( (~ Ng3115) ) ;
 assign n4133 = ( (~ Pg35) ) | ( n3583 ) | ( Ng3119 ) ;
 assign n4135 = ( (~ Ng2715) ) | ( Ng2719 ) ;
 assign n4136 = ( (~ Pg35)  &  (~ Ng2715) ) | ( Pg35  &  n4862 ) | ( (~ Ng2715)  &  n4862 ) ;
 assign n4134 = ( n4135  &  n1736  &  n4136 ) ;
 assign n4138 = ( Pg35 ) | ( (~ Ng1484) ) ;
 assign n4139 = ( (~ Pg35) ) | ( (~ Ng1300) ) | ( n5132 ) ;
 assign n4140 = ( (~ Pg35) ) | ( (~ n854) ) | ( (~ Ng1384) ) ;
 assign n4141 = ( Ng1384 ) | ( n854 ) | ( n5088 ) ;
 assign n4144 = ( (~ Ng1361) ) | ( (~ Ng1373) ) ;
 assign n4142 = ( (~ n2194)  &  (~ n5088) ) | ( n4144  &  (~ n5088)  &  (~ n6036) ) ;
 assign n4149 = ( Pg35  &  (~ Pg12923) ) | ( Pg35  &  Ng1266 ) ;
 assign n4152 = ( Ng1249 ) | ( n4222 ) ;
 assign n4154 = ( Pg35 ) | ( (~ Ng1141) ) ;
 assign n4155 = ( (~ Pg35) ) | ( (~ Ng956) ) | ( n5135 ) ;
 assign n4156 = ( (~ Pg35) ) | ( (~ n379) ) | ( (~ Ng1041) ) ;
 assign n4157 = ( Ng1041 ) | ( n379 ) | ( n5093 ) ;
 assign n4160 = ( (~ Ng1018) ) | ( (~ Ng1030) ) ;
 assign n4158 = ( (~ n2207)  &  (~ n5093) ) | ( n4160  &  (~ n5093)  &  (~ n6044) ) ;
 assign n4165 = ( Pg35  &  (~ Pg12919) ) | ( Pg35  &  Ng921 ) ;
 assign n4168 = ( Ng904 ) | ( n4235 ) ;
 assign n4170 = ( (~ Ng385) ) | ( n4201 ) | ( (~ Ng370) ) ;
 assign n4169 = ( Pg35  &  (~ n3784) ) | ( Pg35  &  Ng832 ) | ( Pg35  &  n4170 ) ;
 assign n4176 = ( n5184 ) | ( n5185 ) ;
 assign n4177 = ( n4388 ) | ( n4389 ) ;
 assign n4178 = ( n1215 ) | ( (~ Ng732) ) ;
 assign n4182 = ( (~ Pg35) ) | ( n4192 ) | ( (~ n4365) ) ;
 assign n4183 = ( Pg35 ) | ( (~ Ng691) ) ;
 assign n4180 = ( (~ Pg35) ) | ( (~ n4192) ) ;
 assign n4186 = ( (~ n1205)  &  Ng562 ) | ( n1205  &  (~ Ng562) ) ;
 assign n4184 = ( (~ Ng632)  &  n4186  &  (~ n4508) ) | ( (~ Ng626)  &  n4186  &  (~ n4508) ) ;
 assign n4192 = ( (~ Ng385) ) | ( Ng376 ) | ( (~ Ng358) ) ;
 assign n4190 = ( Pg35  &  n4192 ) | ( Pg35  &  (~ n5056) ) ;
 assign n4196 = ( n4180  &  (~ Ng499) ) | ( (~ n4180)  &  (~ Ng504) ) | ( (~ Ng499)  &  (~ Ng504) ) ;
 assign n4198 = ( (~ Ng246)  &  (~ n5137) ) | ( n5136  &  (~ n5137) ) | ( (~ Ng246)  &  (~ Ng460) ) | ( n5136  &  (~ Ng460) ) ;
 assign n4200 = ( (~ Ng182)  &  (~ Ng446) ) | ( (~ Ng182)  &  n5136 ) | ( (~ Ng446)  &  (~ n5137) ) | ( n5136  &  (~ n5137) ) ;
 assign n4202 = ( Pg35 ) | ( (~ Ng376) ) ;
 assign n4203 = ( (~ Pg35) ) | ( (~ Ng385) ) | ( (~ n4201) ) ;
 assign n4201 = ( (~ Ng376) ) | ( (~ Ng358) ) ;
 assign n4204 = ( (~ Pg35) ) | ( Ng4332 ) | ( Ng4322 ) | ( Ng4311 ) | ( n4521 ) ;
 assign n4205 = ( Ng4340 ) | ( (~ Ng4643) ) ;
 assign n4208 = ( (~ Ng4633) ) | ( Ng4616 ) | ( n4204 ) | ( Ng4601 ) | ( Ng4584 ) | ( Ng4608 ) | ( Ng4593 ) | ( n4637 ) ;
 assign n4210 = ( (~ Pg35) ) | ( Ng4258 ) ;
 assign n4209 = ( (~ Pg35)  &  n4210 ) | ( n4210  &  Ng4264 ) ;
 assign n4211 = ( (~ Pg35)  &  n4209 ) | ( n4209  &  Ng4269 ) ;
 assign n4212 = ( Pg35  &  (~ Ng4264) ) | ( Pg35  &  Ng4273 ) | ( Pg35  &  (~ Ng4258) ) ;
 assign n4218 = ( Pg35  &  Ng2715 ) | ( (~ Pg35)  &  (~ Ng2712) ) | ( Ng2715  &  (~ Ng2712) ) ;
 assign n4217 = ( n4218  &  n1736 ) ;
 assign n4220 = ( Pg35 ) | ( (~ Ng1548) ) ;
 assign n4221 = ( (~ Pg35) ) | ( (~ Ng1564) ) | ( n5130 ) ;
 assign n4222 = ( (~ Pg35) ) | ( (~ Pg12923) ) ;
 assign n4223 = ( Ng1548  &  Pg35 ) ;
 assign n4226 = ( (~ n854)  &  (~ n1218)  &  n4392 ) ;
 assign n4225 = ( n4226  &  Pg35 ) ;
 assign n4227 = ( Pg35 ) | ( (~ Ng1589) ) ;
 assign n4228 = ( (~ Pg35) ) | ( Pg17423 ) | ( (~ Pg10527) ) ;
 assign n4231 = ( Pg35  &  (~ Pg12923) ) ;
 assign n4233 = ( Pg35 ) | ( (~ Ng1205) ) ;
 assign n4234 = ( (~ Pg35) ) | ( (~ Ng1221) ) | ( n5133 ) ;
 assign n4235 = ( (~ Pg35) ) | ( (~ Pg12919) ) ;
 assign n4236 = ( Ng1205  &  Pg35 ) ;
 assign n4239 = ( n4393  &  n634 ) ;
 assign n4238 = ( n4239  &  Pg35 ) ;
 assign n4241 = ( Pg35 ) | ( (~ Ng1246) ) ;
 assign n4242 = ( (~ Pg35) ) | ( Pg17400 ) | ( (~ Pg10500) ) ;
 assign n4245 = ( Pg35  &  (~ Pg12919) ) ;
 assign n4246 = ( Pg35  &  n3786  &  (~ Ng832) ) | ( Pg35  &  n3786  &  (~ Ng827) ) ;
 assign n4248 = ( (~ n4170)  &  Ng847 ) ;
 assign n4247 = ( (~ Pg35)  &  Ng703 ) | ( (~ Ng837)  &  Ng703  &  n4248 ) ;
 assign n4251 = ( (~ Pg35)  &  n3812 ) | ( Ng837  &  (~ n3786)  &  n3812 ) ;
 assign n4253 = ( Pg35  &  Ng847 ) | ( Pg35  &  n6102 ) | ( (~ Ng847)  &  n6102 ) ;
 assign n4256 = ( Ng691  &  (~ Ng542) ) ;
 assign n4259 = ( (~ Pg35) ) | ( n4170 ) ;
 assign n4261 = ( n3812  &  n4259 ) | ( n3812  &  (~ Ng246) ) | ( n4259  &  (~ Ng475) ) | ( (~ Ng246)  &  (~ Ng475) ) ;
 assign n4263 = ( n3812  &  n4259 ) | ( n3812  &  (~ Ng269) ) | ( n4259  &  (~ Ng433) ) | ( (~ Ng269)  &  (~ Ng433) ) ;
 assign n4265 = ( n3812 ) | ( (~ Ng392) ) ;
 assign n4266 = ( Ng703 ) | ( n4259 ) | ( (~ Ng854) ) ;
 assign n4267 = ( Pg35  &  Ng4269 ) | ( Pg35  &  (~ Ng4258) ) ;
 assign n4268 = ( Ng4264  &  Pg35 ) ;
 assign n4271 = ( (~ Ng4349) ) | ( n4303 ) ;
 assign n4270 = ( Pg35  &  n4271 ) ;
 assign n4272 = ( (~ n4368)  &  (~ Ng2988) ) ;
 assign n4275 = ( (~ Ng4564) ) | ( (~ Ng4555) ) | ( (~ Ng4561) ) | ( (~ Ng4558) ) ;
 assign n4274 = ( n4275  &  (~ Ng2988) ) ;
 assign n4276 = ( Pg35  &  (~ Ng2667) ) ;
 assign n4277 = ( Pg35  &  (~ Ng2527) ) ;
 assign n4279 = ( Pg35  &  (~ Ng2399) ) ;
 assign n4280 = ( Pg35  &  (~ Ng2265) ) ;
 assign n4281 = ( Pg35  &  (~ Ng2102) ) ;
 assign n4283 = ( Pg35  &  (~ Ng1968) ) ;
 assign n4285 = ( Pg35  &  (~ Ng1840) ) ;
 assign n4286 = ( Pg35  &  (~ Ng1706) ) ;
 assign n4288 = ( n4356 ) | ( (~ Ng1542) ) ;
 assign n4287 = ( Pg35  &  n4288 ) ;
 assign n4290 = ( n4358 ) | ( (~ Ng1199) ) ;
 assign n4289 = ( Pg35  &  n4290 ) ;
 assign n4291 = ( Pg35  &  (~ Ng6533) ) ;
 assign n4292 = ( Pg35  &  (~ Ng6187) ) ;
 assign n4293 = ( Pg35  &  (~ Ng5841) ) ;
 assign n4294 = ( Pg35  &  (~ Ng5495) ) ;
 assign n4295 = ( Pg35  &  (~ Ng5148) ) ;
 assign n4296 = ( Pg35  &  (~ Ng3841) ) ;
 assign n4297 = ( Pg35  &  (~ Ng3490) ) ;
 assign n4298 = ( Pg35  &  (~ Ng3139) ) ;
 assign n4299 = ( Pg35  &  (~ n1621) ) | ( (~ n1621)  &  (~ Ng385) ) ;
 assign Ng25599 = ( (~ n4299) ) ;
 assign n4300 = ( (~ Ng4593) ) | ( (~ n4640) ) ;
 assign n4301 = ( Ng4332  &  Ng4322  &  n4638 ) ;
 assign n4303 = ( (~ Ng4628) ) | ( n4637 ) ;
 assign n4302 = ( (~ Ng4349)  &  n4303 ) | ( Ng4349  &  (~ n4303) ) ;
 assign n4304 = ( (~ Ng4688) ) | ( n4556 ) ;
 assign n4307 = ( Ng2599 ) | ( (~ Ng2629) ) ;
 assign n4305 = ( n4307  &  Ng112 ) | ( (~ n4307)  &  (~ Ng112) ) ;
 assign n4309 = ( Ng2465 ) | ( (~ Ng2495) ) ;
 assign n4308 = ( n4309  &  Ng112 ) | ( (~ n4309)  &  (~ Ng112) ) ;
 assign n4311 = ( Ng2331 ) | ( (~ Ng2361) ) ;
 assign n4310 = ( n4311  &  Ng112 ) | ( (~ n4311)  &  (~ Ng112) ) ;
 assign n4313 = ( Ng2197 ) | ( (~ Ng2227) ) ;
 assign n4312 = ( n4313  &  Ng112 ) | ( (~ n4313)  &  (~ Ng112) ) ;
 assign n4315 = ( Ng2040 ) | ( (~ Ng2070) ) ;
 assign n4314 = ( n4315  &  Ng112 ) | ( (~ n4315)  &  (~ Ng112) ) ;
 assign n4317 = ( Ng1906 ) | ( (~ Ng1936) ) ;
 assign n4316 = ( n4317  &  Ng112 ) | ( (~ n4317)  &  (~ Ng112) ) ;
 assign n4319 = ( Ng1772 ) | ( (~ Ng1802) ) ;
 assign n4318 = ( n4319  &  Ng112 ) | ( (~ n4319)  &  (~ Ng112) ) ;
 assign n4321 = ( Ng1636 ) | ( (~ Ng1668) ) ;
 assign n4320 = ( n4321  &  Ng112 ) | ( (~ n4321)  &  (~ Ng112) ) ;
 assign n4322 = ( Ng1339  &  Ng1322 ) | ( (~ Ng1339)  &  (~ Ng1322) ) ;
 assign n4323 = ( Ng996  &  Ng979 ) | ( (~ Ng996)  &  (~ Ng979) ) ;
 assign n4325 = ( Ng2610 ) | ( (~ Ng2619) ) ;
 assign n4324 = ( (~ Ng110)  &  n4325 ) | ( Ng110  &  (~ n4325) ) ;
 assign n4327 = ( Ng2476 ) | ( (~ Ng2485) ) ;
 assign n4326 = ( (~ Ng110)  &  n4327 ) | ( Ng110  &  (~ n4327) ) ;
 assign n4329 = ( Ng2342 ) | ( (~ Ng2351) ) ;
 assign n4328 = ( (~ Ng110)  &  n4329 ) | ( Ng110  &  (~ n4329) ) ;
 assign n4331 = ( Ng2208 ) | ( (~ Ng2217) ) ;
 assign n4330 = ( (~ Ng110)  &  n4331 ) | ( Ng110  &  (~ n4331) ) ;
 assign n4333 = ( Ng2051 ) | ( (~ Ng2060) ) ;
 assign n4332 = ( (~ Ng110)  &  n4333 ) | ( Ng110  &  (~ n4333) ) ;
 assign n4335 = ( Ng1917 ) | ( (~ Ng1926) ) ;
 assign n4334 = ( (~ Ng110)  &  n4335 ) | ( Ng110  &  (~ n4335) ) ;
 assign n4337 = ( Ng1783 ) | ( (~ Ng1792) ) ;
 assign n4336 = ( (~ Ng110)  &  n4337 ) | ( Ng110  &  (~ n4337) ) ;
 assign n4339 = ( Ng1648 ) | ( (~ Ng1657) ) ;
 assign n4338 = ( (~ Ng110)  &  n4339 ) | ( Ng110  &  (~ n4339) ) ;
 assign n4341 = ( Pg35  &  Ng5471 ) ;
 assign n4340 = ( n2562  &  n4341 ) | ( n2563  &  n4341 ) | ( n2562  &  n2559 ) | ( n2563  &  n2559 ) ;
 assign n4343 = ( n4341 ) | ( n2562 ) | ( n2563 ) ;
 assign n4342 = ( n2565  &  n4343 ) ;
 assign n4344 = ( n2564  &  n2565 ) | ( n2564  &  n4343 ) ;
 assign n4345 = ( Pg35  &  Ng3466 ) ;
 assign n4346 = ( (~ Ng2735) ) | ( n3634 ) ;
 assign n4347 = ( Ng2652  &  Ng2648 ) | ( (~ Ng2652)  &  (~ Ng2648) ) ;
 assign n4348 = ( Ng2514  &  Ng2518 ) | ( (~ Ng2514)  &  (~ Ng2518) ) ;
 assign n4349 = ( Ng2384  &  Ng2380 ) | ( (~ Ng2384)  &  (~ Ng2380) ) ;
 assign n4350 = ( Ng2250  &  Ng2246 ) | ( (~ Ng2250)  &  (~ Ng2246) ) ;
 assign n4351 = ( Ng2089  &  Ng2093 ) | ( (~ Ng2089)  &  (~ Ng2093) ) ;
 assign n4352 = ( Ng1955  &  Ng1959 ) | ( (~ Ng1955)  &  (~ Ng1959) ) ;
 assign n4353 = ( Ng1821  &  Ng1825 ) | ( (~ Ng1821)  &  (~ Ng1825) ) ;
 assign n4354 = ( Ng1687  &  Ng1691 ) | ( (~ Ng1687)  &  (~ Ng1691) ) ;
 assign n4356 = ( (~ Pg7946) ) | ( (~ Ng1526) ) | ( n1219 ) | ( Ng1514 ) ;
 assign n4355 = ( (~ n4356)  &  Ng1542 ) | ( n4356  &  (~ Ng1542) ) ;
 assign n4358 = ( (~ Pg7916) ) | ( Ng1171 ) | ( (~ Ng1183) ) | ( n4977 ) ;
 assign n4357 = ( (~ n4358)  &  Ng1199 ) | ( n4358  &  (~ Ng1199) ) ;
 assign n4359 = ( n1176  &  n3456 ) | ( (~ n1176)  &  (~ n3456) ) ;
 assign n4360 = ( n1195  &  n3465 ) | ( (~ n1195)  &  (~ n3465) ) ;
 assign n4361 = ( (~ Ng4076) ) | ( n3867 ) ;
 assign n4363 = ( n1173  &  (~ n4170)  &  Ng499  &  (~ Ng504) ) ;
 assign n4365 = ( (~ Ng703) ) | ( n3794 ) | ( Ng691 ) ;
 assign n4364 = ( n3894  &  n4192 ) | ( n4192  &  (~ Ng691) ) | ( n3894  &  n4365 ) | ( (~ Ng691)  &  n4365 ) ;
 assign n4366 = ( n1150  &  n1086 ) | ( n3907  &  n1086 ) | ( n1150  &  n3906 ) | ( n3907  &  n3906 ) ;
 assign n4368 = ( Ng4483  &  Ng4486  &  Ng4492  &  Ng4489 ) ;
 assign n4367 = ( n4368  &  (~ Ng4521)  &  (~ n5999) ) | ( Ng4527  &  (~ Ng4521)  &  (~ n5999) ) ;
 assign n4371 = ( (~ n1209)  &  (~ Ng1536) ) | ( (~ n1209)  &  (~ n4288)  &  Ng1413 ) ;
 assign n4374 = ( n3985  &  Ng1404 ) | ( (~ n3985)  &  (~ Ng1404) ) ;
 assign n4376 = ( (~ n1211)  &  (~ Ng1193) ) | ( (~ n1211)  &  (~ n4290)  &  Ng1070 ) ;
 assign n4379 = ( (~ Ng832) ) | ( n4170 ) | ( (~ Ng817) ) ;
 assign n4380 = ( n4363  &  Ng728 ) | ( n4363  &  Ng661  &  Pg35 ) ;
 assign n4382 = ( n5130  &  Ng1564 ) ;
 assign n4381 = ( n4382  &  Ng1559 ) | ( (~ n4382)  &  (~ Ng1559) ) ;
 assign n4385 = ( n5133  &  Ng1221 ) ;
 assign n4384 = ( n4385  &  Ng1216 ) | ( (~ n4385)  &  (~ Ng1216) ) ;
 assign n4387 = ( (~ Ng232)  &  Ng255 ) | ( Ng232  &  (~ Ng255) ) ;
 assign n4388 = ( Ng246  &  Ng269 ) | ( (~ Ng246)  &  (~ Ng269) ) ;
 assign n4389 = ( Ng239  &  Ng262 ) | ( (~ Ng239)  &  (~ Ng262) ) ;
 assign n4392 = ( (~ Ng1322)  &  Ng1579 ) | ( Ng1322  &  (~ Ng1579) ) ;
 assign n4393 = ( (~ Ng1236)  &  Ng979 ) | ( Ng1236  &  (~ Ng979) ) ;
 assign n4394 = ( Pg57 ) | ( Pg56 ) | ( (~ Pg54) ) | ( Pg53 ) | ( Ng55 ) ;
 assign n4397 = ( (~ Ng50) ) | ( Ng16 ) ;
 assign n4398 = ( Ng48  &  Ng45  &  Ng8  &  Ng46  &  (~ Ng52) ) ;
 assign n4401 = ( Ng46 ) | ( Ng8 ) | ( Ng45 ) ;
 assign n4402 = ( (~ Ng51) ) | ( n4401 ) | ( Ng52 ) ;
 assign n4403 = ( Ng48 ) | ( n4402 ) ;
 assign n4404 = ( Ng50 ) | ( (~ Ng16) ) ;
 assign n4406 = ( n4403 ) | ( n4404 ) ;
 assign n4407 = ( Ng16 ) | ( Ng50 ) ;
 assign n4411 = ( Ng48 ) | ( n4401 ) | ( (~ Ng52) ) ;
 assign Ng29209 = ( (~ n4394) ) ;
 assign n4412 = ( Pg53 ) | ( (~ n4394) ) ;
 assign n4414 = ( Ng51 ) | ( Ng52 ) | ( n4401 ) ;
 assign n4416 = ( n4394 ) | ( n1351 ) ;
 assign n4417 = ( Ng48 ) | ( n4414 ) ;
 assign n4419 = ( Ng51 ) | ( n4397 ) | ( n4411 ) ;
 assign n4418 = ( n4419  &  n1331  &  n1289 ) ;
 assign n4421 = ( n4407 ) | ( n4417 ) ;
 assign n4425 = ( n4404 ) | ( n4417 ) ;
 assign n4426 = ( n4394 ) | ( n4425 ) ;
 assign n4427 = ( n4397 ) | ( n4403 ) ;
 assign n4428 = ( n4394 ) | ( n4427 ) ;
 assign n4429 = ( (~ Ng48) ) | ( n4397 ) ;
 assign n4430 = ( n4402 ) | ( n4429 ) ;
 assign n4431 = ( n4394 ) | ( n4430 ) ;
 assign n4432 = ( n4394 ) | ( Ng48 ) | ( (~ Ng50) ) | ( (~ Ng16) ) ;
 assign n4433 = ( n4402 ) | ( n4432 ) ;
 assign n4434 = ( n4414 ) | ( n4432 ) ;
 assign n4441 = ( n4414 ) | ( n4429 ) ;
 assign n4442 = ( n4394 ) | ( n4441 ) ;
 assign n4443 = ( Ng51 ) | ( n4401 ) | ( (~ Ng52) ) | ( n4429 ) ;
 assign n4444 = ( n4394 ) | ( n4443 ) ;
 assign n4449 = ( (~ n4398) ) | ( Ng51 ) | ( n4404 ) ;
 assign n4464 = ( Ng1291 ) | ( n4426 ) ;
 assign n4465 = ( Ng947 ) | ( n4428 ) ;
 assign n4486 = ( n1359 ) | ( n1363 ) ;
 assign n4487 = ( (~ Ng4322)  &  Pg72 ) | ( Ng4322  &  (~ Pg72) ) ;
 assign n4488 = ( (~ Ng4332)  &  Pg73 ) | ( Ng4332  &  (~ Pg73) ) ;
 assign n4490 = ( Pg11678  &  (~ Ng736) ) ;
 assign n4492 = ( (~ Ng385) ) | ( n4201 ) | ( Ng370 ) ;
 assign n4503 = ( Pg9048  &  (~ Ng559) ) ;
 assign n4508 = ( (~ Pg35) ) | ( n4503 ) ;
 assign n4509 = ( (~ Ng490)  &  Pg73 ) | ( Ng490  &  (~ Pg73) ) ;
 assign n4510 = ( (~ Ng482)  &  Pg72 ) | ( Ng482  &  (~ Pg72) ) ;
 assign n4511 = ( Ng518 ) | ( n1170 ) ;
 assign n4512 = ( n1170 ) | ( (~ Ng518) ) ;
 assign n4515 = ( (~ Ng4349) ) | ( Ng4358 ) ;
 assign n4516 = ( (~ Ng3352) ) | ( (~ Ng3288) ) ;
 assign n4518 = ( Ng4349 ) | ( (~ Ng4358) ) ;
 assign n4521 = ( Ng4358 ) | ( Ng4349 ) ;
 assign n4527 = ( (~ Ng5357) ) | ( (~ Ng5297) ) ;
 assign n4531 = ( (~ Ng2759)  &  Pg72 ) | ( Ng2759  &  (~ Pg72) ) ;
 assign n4532 = ( (~ Ng2763)  &  Pg73 ) | ( Ng2763  &  (~ Pg73) ) ;
 assign n4530 = ( n4531 ) | ( n4532 ) ;
 assign n4533 = ( (~ Ng2756) ) | ( Ng2748 ) | ( n4530 ) ;
 assign n4535 = ( (~ Ng2208) ) | ( Ng2217 ) ;
 assign n4536 = ( Ng2756 ) | ( Ng2748 ) | ( (~ Ng2741) ) ;
 assign n4538 = ( (~ Ng1783) ) | ( Ng1792 ) ;
 assign n4540 = ( (~ Ng2748) ) | ( n4530 ) ;
 assign n4542 = ( (~ Ng2051) ) | ( Ng2060 ) ;
 assign n4544 = ( (~ Ng1917) ) | ( Ng1926 ) ;
 assign n4546 = ( (~ Ng2476) ) | ( Ng2485 ) ;
 assign n4548 = ( (~ Ng2342) ) | ( Ng2351 ) ;
 assign n4550 = ( (~ Ng2610) ) | ( Ng2619 ) ;
 assign n4551 = ( (~ Ng2756)  &  (~ Ng2748)  &  (~ Ng2741) ) ;
 assign n4553 = ( (~ Ng1648) ) | ( Ng1657 ) ;
 assign n4556 = ( (~ Ng4669) ) | ( (~ Ng4659) ) | ( (~ Ng4653) ) ;
 assign n4559 = ( (~ Ng4793) ) | ( (~ Ng4776) ) | ( Ng4801 ) ;
 assign n4561 = ( (~ Ng4859) ) | ( (~ Ng4843) ) | ( (~ Ng4849) ) ;
 assign n4564 = ( (~ Ng4983) ) | ( (~ Ng4966) ) | ( Ng4991 ) ;
 assign n4567 = ( n1086 ) | ( n1150 ) | ( n3907 ) ;
 assign n4569 = ( Pg35  &  Ng6509 ) ;
 assign n4568 = ( n1107 ) | ( n2565 ) | ( n4343 ) | ( n2564 ) | ( n4569 ) | ( n4345 ) ;
 assign n4570 = ( n1101  &  (~ n1131)  &  (~ n1133)  &  (~ n1134)  &  (~ n4567) ) ;
 assign n4577 = ( (~ Ng3171) ) | ( (~ Ng3179) ) ;
 assign n4581 = ( (~ Ng6219) ) | ( (~ Ng6227) ) ;
 assign n4582 = ( (~ Ng4098)  &  Ng4093 ) ;
 assign n4584 = ( (~ Ng3873) ) | ( (~ Ng3881) ) ;
 assign n4585 = ( Ng4098  &  Ng4093 ) ;
 assign n4587 = ( (~ Ng5527) ) | ( (~ Ng5535) ) ;
 assign n4588 = ( (~ Ng6565) ) | ( (~ Ng6573) ) ;
 assign n4590 = ( (~ Ng5873) ) | ( (~ Ng5881) ) ;
 assign n4593 = ( (~ Ng3522) ) | ( (~ Ng3530) ) ;
 assign n4595 = ( (~ Ng5180) ) | ( (~ Ng5188) ) ;
 assign n4596 = ( (~ Ng4108)  &  Pg72 ) | ( Ng4108  &  (~ Pg72) ) ;
 assign n4597 = ( (~ Ng4104)  &  Pg73 ) | ( Ng4104  &  (~ Pg73) ) ;
 assign n4630 = ( n1408  &  (~ n4673) ) ;
 assign n4632 = ( (~ Ng4878) ) | ( (~ Ng4843) ) ;
 assign n4633 = ( n4304  &  (~ n4676) ) ;
 assign n4635 = ( (~ Ng4688) ) | ( (~ Ng4653) ) ;
 assign n4637 = ( (~ Ng4621) ) | ( Ng4639 ) | ( (~ Ng4340) ) ;
 assign n4638 = ( (~ n4271)  &  Ng4358 ) ;
 assign n4640 = ( Ng4584  &  n4301 ) ;
 assign n4641 = ( (~ Pg35) ) | ( n1572 ) ;
 assign n4642 = ( Ng4311  &  n4638 ) ;
 assign n4652 = ( Ng4818 ) | ( wire4661 ) | ( n1160 ) ;
 assign n4653 = ( (~ n4652)  &  Ng71 ) ;
 assign n4654 = ( Ng4818 ) | ( wire4661 ) | ( n1160 ) ;
 assign n4659 = ( (~ n282)  &  Ng278 ) | ( (~ n282)  &  n281 ) | ( (~ Ng278)  &  n281 ) ;
 assign n4657 = ( (~ n1212)  &  Ng691  &  n4659 ) ;
 assign n4660 = ( Ng287  &  Ng283  &  n4657 ) ;
 assign n4661 = ( (~ n4660) ) | ( (~ Ng291) ) ;
 assign n4663 = ( (~ Ng294) ) | ( n4661 ) ;
 assign n4664 = ( (~ Ng298) ) | ( n4663 ) ;
 assign n4666 = ( n1212 ) | ( n1691 ) | ( (~ Ng691) ) ;
 assign n4667 = ( n359  &  Ng146  &  (~ n4666) ) ;
 assign n4669 = ( Ng164  &  n4667 ) ;
 assign n4670 = ( (~ n4669) ) | ( (~ Ng150) ) ;
 assign n4672 = ( (~ Ng153) ) | ( n4670 ) ;
 assign n4673 = ( n1221  &  (~ n1406)  &  Ng63 ) ;
 assign n4674 = ( (~ n1710)  &  Ng4966 ) ;
 assign n4676 = ( n1221  &  (~ n1368)  &  Ng63 ) ;
 assign n4677 = ( (~ n1726)  &  Ng4776 ) ;
 assign n4689 = ( (~ Ng2715) ) | ( (~ Ng2719) ) ;
 assign n4690 = ( (~ Ng2724) ) | ( n4689 ) ;
 assign n4691 = ( n4346 ) | ( (~ Ng2741) ) ;
 assign n4692 = ( (~ Ng2748) ) | ( n4691 ) ;
 assign n4695 = ( Ng1564 ) | ( Ng1548 ) | ( (~ Ng1322) ) | ( Ng1559 ) | ( Ng1554 ) | ( (~ Ng1404) ) ;
 assign n4696 = ( (~ Ng2629)  &  (~ Ng2555) ) ;
 assign n4697 = ( (~ n4696) ) | ( (~ n4700) ) ;
 assign n4699 = ( n4697  &  Pg35 ) ;
 assign n4700 = ( n1140 ) | ( (~ n1261) ) ;
 assign n4702 = ( Ng2599  &  (~ Ng2555) ) ;
 assign n4703 = ( n4700  &  n4702 ) ;
 assign n4704 = ( (~ n4700) ) | ( (~ Ng2555) ) ;
 assign n4706 = ( (~ Ng2495)  &  (~ Ng2421) ) ;
 assign n4707 = ( (~ n4706) ) | ( (~ n4710) ) ;
 assign n4709 = ( n4707  &  Pg35 ) ;
 assign n4710 = ( n1093 ) | ( (~ n1264) ) ;
 assign n4712 = ( Ng2465  &  (~ Ng2421) ) ;
 assign n4713 = ( n4710  &  n4712 ) ;
 assign n4714 = ( (~ n4710) ) | ( (~ Ng2421) ) ;
 assign n4716 = ( (~ Ng2361)  &  (~ Ng2287) ) ;
 assign n4717 = ( (~ n4716) ) | ( (~ n4720) ) ;
 assign n4719 = ( n4717  &  Pg35 ) ;
 assign n4720 = ( n1138 ) | ( (~ n1274) ) ;
 assign n4722 = ( Ng2331  &  (~ Ng2287) ) ;
 assign n4723 = ( n4720  &  n4722 ) ;
 assign n4724 = ( (~ n4720) ) | ( (~ Ng2287) ) ;
 assign n4726 = ( (~ Ng2227)  &  (~ Ng2153) ) ;
 assign n4727 = ( (~ n4726) ) | ( (~ n4730) ) ;
 assign n4729 = ( n4727  &  Pg35 ) ;
 assign n4730 = ( n1096 ) | ( (~ n1270) ) ;
 assign n4731 = ( (~ Ng2227) ) | ( (~ n4730) ) ;
 assign n4733 = ( Ng2197  &  (~ Ng2153) ) ;
 assign n4734 = ( n4730  &  n4733 ) ;
 assign n4736 = ( Ng1221 ) | ( Ng1205 ) | ( (~ Ng979) ) | ( (~ Ng1061) ) | ( Ng1216 ) | ( Ng1211 ) ;
 assign n4737 = ( (~ Ng2070)  &  (~ Ng1996) ) ;
 assign n4738 = ( (~ n4737) ) | ( (~ n4741) ) ;
 assign n4740 = ( n4738  &  Pg35 ) ;
 assign n4741 = ( n1155 ) | ( (~ n1266) ) ;
 assign n4742 = ( (~ Ng2070) ) | ( (~ n4741) ) ;
 assign n4744 = ( Ng2040  &  (~ Ng1996) ) ;
 assign n4745 = ( n4741  &  n4744 ) ;
 assign n4747 = ( (~ Ng1936)  &  (~ Ng1862) ) ;
 assign n4748 = ( (~ n4747) ) | ( (~ n4751) ) ;
 assign n4750 = ( n4748  &  Pg35 ) ;
 assign n4751 = ( n1113 ) | ( (~ n1268) ) ;
 assign n4752 = ( (~ Ng1936) ) | ( (~ n4751) ) ;
 assign n4754 = ( Ng1906  &  (~ Ng1862) ) ;
 assign n4755 = ( n4751  &  n4754 ) ;
 assign n4757 = ( (~ Ng1802)  &  (~ Ng1728) ) ;
 assign n4758 = ( (~ n4757) ) | ( (~ n4761) ) ;
 assign n4760 = ( n4758  &  Pg35 ) ;
 assign n4761 = ( n1120 ) | ( (~ n1258) ) ;
 assign n4763 = ( Ng1772  &  (~ Ng1728) ) ;
 assign n4764 = ( n4761  &  n4763 ) ;
 assign n4765 = ( (~ n4761) ) | ( (~ Ng1728) ) ;
 assign n4767 = ( (~ Ng1592)  &  (~ Ng1668) ) ;
 assign n4768 = ( (~ n4767) ) | ( (~ n4771) ) ;
 assign n4770 = ( n4768  &  Pg35 ) ;
 assign n4771 = ( wire4406 ) | ( (~ n1272) ) ;
 assign n4773 = ( (~ Ng1636) ) | ( (~ n4771) ) ;
 assign n4774 = ( (~ Ng1592) ) | ( (~ n4771) ) ;
 assign n4776 = ( Ng4793 ) | ( (~ Ng4776) ) | ( Ng4801 ) ;
 assign n4777 = ( Ng4983 ) | ( (~ Ng4966) ) | ( Ng4991 ) ;
 assign n4778 = ( n1221  &  Ng93 ) ;
 assign n4779 = ( n1406 ) | ( (~ n4778) ) ;
 assign n4781 = ( n1368 ) | ( (~ n4778) ) ;
 assign n4783 = ( (~ Ng5703) ) | ( Ng5644 ) ;
 assign n4784 = ( (~ Pg35) ) | ( (~ n1097) ) ;
 assign n4786 = ( (~ Ng4057) ) | ( (~ Ng4064) ) ;
 assign n4787 = ( (~ n4786)  &  Ng4141 ) ;
 assign n4790 = ( (~ Ng4087) ) | ( n4361 ) ;
 assign n4791 = ( (~ Ng4093) ) | ( n4790 ) ;
 assign n4792 = ( Ng3703 ) | ( (~ Ng3639) ) ;
 assign n4793 = ( (~ Pg35) ) | ( (~ n1135) ) ;
 assign n4794 = ( Pg35  &  n1221 ) ;
 assign n4796 = ( n1221  &  Ng112 ) ;
 assign n4806 = ( n4322 ) | ( Ng1351 ) ;
 assign n4807 = ( n4144 ) | ( (~ Ng1351) ) | ( (~ n4322) ) ;
 assign n4805 = ( (~ Ng1312)  &  n4806  &  n4807  &  (~ n6036) ) ;
 assign n4808 = ( (~ Pg12923) ) | ( (~ Ng1266) ) | ( (~ Ng1249) ) ;
 assign n4810 = ( Ng1252  &  (~ n3877) ) ;
 assign n4813 = ( Ng1259  &  (~ n3156) ) ;
 assign n4819 = ( n4323 ) | ( Ng1008 ) ;
 assign n4820 = ( (~ Ng1008) ) | ( n4160 ) | ( (~ n4323) ) ;
 assign n4818 = ( (~ Ng969)  &  n4819  &  n4820  &  (~ n6044) ) ;
 assign n4821 = ( (~ Pg12919) ) | ( (~ Ng921) ) | ( (~ Ng904) ) ;
 assign n4823 = ( Ng907  &  (~ n3883) ) ;
 assign n4826 = ( Ng914  &  (~ n3172) ) ;
 assign n4830 = ( (~ n1191)  &  n1221  &  Ng43 ) ;
 assign n4832 = ( (~ Ng4087)  &  n4830 ) ;
 assign Ng25756 = ( Pg35  &  Ng6573 ) ;
 assign n4833 = ( (~ Ng6565) ) | ( Ng6573 ) ;
 assign n4835 = ( Ng4087  &  n4830 ) ;
 assign n4836 = ( (~ Ng6219) ) | ( Ng6227 ) ;
 assign Ng25728 = ( Pg35  &  Ng5881 ) ;
 assign n4837 = ( (~ Ng5873) ) | ( Ng5881 ) ;
 assign n4838 = ( (~ Ng5527) ) | ( Ng5535 ) ;
 assign n4839 = ( (~ Ng5180) ) | ( Ng5188 ) ;
 assign n4840 = ( (~ Ng5029) ) | ( (~ Ng5016) ) | ( (~ Ng5062) ) ;
 assign n4842 = ( n4840 ) | ( (~ Ng5037) ) | ( (~ Ng5033) ) ;
 assign n4844 = ( Ng5029 ) | ( Ng5016 ) | ( (~ Ng5022) ) ;
 assign n4845 = ( Ng5033 ) | ( Ng5037 ) | ( n4844 ) ;
 assign n4846 = ( Ng5046 ) | ( Ng5041 ) | ( n4845 ) ;
 assign n4848 = ( (~ Ng5046)  &  Ng5022  &  Ng5057 ) ;
 assign n4849 = ( Ng5062  &  Ng5046  &  (~ Ng5057) ) ;
 assign n4851 = ( Pg84  &  (~ Ng5041)  &  n4848 ) ;
 assign n4852 = ( (~ Pg84)  &  Ng5052  &  n4849 ) ;
 assign n4853 = ( (~ Pg84)  &  (~ Ng5052)  &  n4848 ) ;
 assign n4854 = ( Pg84  &  Ng5041  &  n4849 ) ;
 assign n4850 = ( n4851 ) | ( n4852 ) | ( n4853 ) | ( n4854 ) ;
 assign n4855 = ( (~ Ng3873) ) | ( Ng3881 ) ;
 assign n4856 = ( (~ Ng3522) ) | ( Ng3530 ) ;
 assign n4857 = ( (~ Ng3171) ) | ( Ng3179 ) ;
 assign n4859 = ( n1221  &  Ng110 ) ;
 assign n4860 = ( (~ Pg35) ) | ( (~ n1153) ) ;
 assign n4862 = ( Ng2715 ) | ( (~ Ng2719) ) ;
 assign n4864 = ( (~ Pg35) ) | ( (~ n1151) ) ;
 assign n4866 = ( (~ Pg35) ) | ( (~ n1162) ) ;
 assign n4868 = ( Ng2719 ) | ( Ng2715 ) ;
 assign n4870 = ( (~ Pg35) ) | ( (~ n1104) ) ;
 assign n4873 = ( (~ Pg35) ) | ( (~ n1146) ) ;
 assign n4875 = ( (~ Pg35) ) | ( (~ n1126) ) ;
 assign n4878 = ( (~ Pg35) ) | ( (~ n1182) ) ;
 assign n4881 = ( (~ Pg35) ) | ( (~ n1087) ) ;
 assign n4883 = ( n4845  &  n4842 ) ;
 assign n4884 = ( Ng5062 ) | ( Ng5022 ) ;
 assign n4886 = ( n3184  &  Pg35 ) ;
 assign n4887 = ( Ng4180  &  (~ Ng4284) ) ;
 assign n4888 = ( Ng6565 ) | ( (~ Ng6573) ) ;
 assign n4889 = ( Ng6565 ) | ( Ng6573 ) ;
 assign n4893 = ( Ng6549 ) | ( Ng6561 ) | ( Ng6555 ) ;
 assign n4894 = ( n3238  &  Pg35 ) ;
 assign n4895 = ( Ng6219 ) | ( (~ Ng6227) ) ;
 assign n4896 = ( Ng6219 ) | ( Ng6227 ) ;
 assign n4900 = ( Ng6215 ) | ( Ng6209 ) | ( Ng6203 ) ;
 assign n4901 = ( n3291  &  Pg35 ) ;
 assign n4902 = ( Ng5873 ) | ( (~ Ng5881) ) ;
 assign n4903 = ( Ng5873 ) | ( Ng5881 ) ;
 assign n4907 = ( Ng5857 ) | ( Ng5869 ) | ( Ng5863 ) ;
 assign n4908 = ( n3346  &  Pg35 ) ;
 assign n4909 = ( Ng5527 ) | ( (~ Ng5535) ) ;
 assign n4910 = ( Ng5527 ) | ( Ng5535 ) ;
 assign n4914 = ( Ng5511 ) | ( Ng5523 ) | ( Ng5517 ) ;
 assign n4915 = ( Ng5180 ) | ( (~ Ng5188) ) ;
 assign n4916 = ( Ng5180 ) | ( Ng5188 ) ;
 assign n4919 = ( Ng5164 ) | ( Ng5176 ) | ( Ng5170 ) ;
 assign n4922 = ( n3476  &  Pg35 ) ;
 assign n4923 = ( Ng3873 ) | ( (~ Ng3881) ) ;
 assign n4924 = ( Ng3873 ) | ( Ng3881 ) ;
 assign n4927 = ( Ng3869 ) | ( Ng3863 ) | ( Ng3857 ) ;
 assign n4928 = ( n3531  &  Pg35 ) ;
 assign n4929 = ( Ng3522 ) | ( (~ Ng3530) ) ;
 assign n4930 = ( Ng3522 ) | ( Ng3530 ) ;
 assign n4933 = ( Ng3506 ) | ( Ng3518 ) | ( Ng3512 ) ;
 assign n4934 = ( n3583  &  Pg35 ) ;
 assign n4935 = ( Ng3171 ) | ( (~ Ng3179) ) ;
 assign n4936 = ( Ng3171 ) | ( Ng3179 ) ;
 assign n4940 = ( Ng3155 ) | ( Ng3167 ) | ( Ng3161 ) ;
 assign n4945 = ( Ng2619  &  n1153  &  Ng2587 ) ;
 assign n4946 = ( Pg35  &  n4945 ) ;
 assign n4947 = ( (~ Ng2610) ) | ( Ng2587 ) ;
 assign n4948 = ( Ng2485  &  n1151 ) ;
 assign n4949 = ( Ng2453  &  n4948 ) ;
 assign n4950 = ( Pg35  &  n4949 ) ;
 assign n4951 = ( (~ Ng2476) ) | ( Ng2453 ) ;
 assign n4952 = ( Ng2351  &  n1162  &  Ng2319 ) ;
 assign n4953 = ( Pg35  &  n4952 ) ;
 assign n4954 = ( (~ Ng2342) ) | ( Ng2319 ) ;
 assign n4955 = ( Ng2217  &  n1104  &  Ng2185 ) ;
 assign n4956 = ( Pg35  &  n4955 ) ;
 assign n4957 = ( (~ Ng2208) ) | ( Ng2185 ) ;
 assign n4958 = ( Ng2060  &  n1146 ) ;
 assign n4959 = ( Ng2028  &  n4958 ) ;
 assign n4960 = ( Pg35  &  n4959 ) ;
 assign n4961 = ( (~ Ng2051) ) | ( Ng2028 ) ;
 assign n4962 = ( Ng1926  &  n1126  &  Ng1894 ) ;
 assign n4963 = ( Pg35  &  n4962 ) ;
 assign n4964 = ( (~ Ng1917) ) | ( Ng1894 ) ;
 assign n4965 = ( Ng1792  &  n1182  &  Ng1760 ) ;
 assign n4966 = ( Pg35  &  n4965 ) ;
 assign n4967 = ( (~ Ng1783) ) | ( Ng1760 ) ;
 assign n4968 = ( Ng1657  &  n1087  &  Ng1624 ) ;
 assign n4969 = ( Pg35  &  n4968 ) ;
 assign n4970 = ( (~ Ng1648) ) | ( Ng1624 ) ;
 assign n4977 = ( Ng996  &  Ng1178  &  (~ Ng1189) ) ;
 assign n4983 = ( (~ n1109) ) | ( n3232 ) ;
 assign n4984 = ( (~ Pg35) ) | ( n4983 ) ;
 assign n4990 = ( (~ n1196) ) | ( n3285 ) ;
 assign n4991 = ( (~ Pg35) ) | ( n4990 ) ;
 assign n4998 = ( (~ n1179) ) | ( n3340 ) ;
 assign n4999 = ( (~ Pg35) ) | ( n4998 ) ;
 assign n5005 = ( (~ n1097) ) | ( n3395 ) ;
 assign n5006 = ( (~ Pg35) ) | ( n5005 ) ;
 assign n5011 = ( wire4415  &  Pg17577  &  (~ n4527) ) ;
 assign n5012 = ( (~ wire4394) ) | ( (~ n5011) ) ;
 assign n5013 = ( (~ Pg35) ) | ( n5012 ) ;
 assign n5023 = ( (~ n1165) ) | ( n3525 ) ;
 assign n5024 = ( (~ Pg35) ) | ( n5023 ) ;
 assign n5030 = ( (~ n1116) ) | ( n3577 ) ;
 assign n5031 = ( (~ Pg35) ) | ( n5030 ) ;
 assign n5034 = ( Ng3639 ) | ( Ng3703 ) ;
 assign n5038 = ( (~ n1135) ) | ( n3628 ) ;
 assign n5039 = ( (~ Pg35) ) | ( n5038 ) ;
 assign n5043 = ( Pg13272  &  Ng1526  &  (~ Ng1514) ) ;
 assign n5044 = ( Ng1514  &  Ng1526  &  Pg13272 ) ;
 assign n5045 = ( Pg13272  &  (~ Ng1526)  &  Ng1514 ) ;
 assign n5046 = ( Pg13259  &  (~ Ng1171)  &  Ng1183 ) ;
 assign n5047 = ( Ng1183  &  Ng1171  &  Pg13259 ) ;
 assign n5048 = ( Pg13259  &  Ng1171  &  (~ Ng1183) ) ;
 assign n5049 = ( n4379 ) | ( (~ Ng822) ) ;
 assign n5051 = ( (~ Ng661)  &  Ng728 ) | ( Ng661  &  (~ Ng728) ) ;
 assign n5052 = ( (~ Ng655)  &  Ng718 ) | ( Ng655  &  (~ Ng718) ) ;
 assign n5054 = ( n4363  &  Ng671 ) ;
 assign n5056 = ( (~ Ng667) ) | ( Ng686 ) ;
 assign n5057 = ( n4192 ) | ( (~ Ng518) ) | ( Ng513 ) ;
 assign n5058 = ( Ng482  &  n1172 ) ;
 assign n5068 = ( n1635  &  (~ Ng4087)  &  (~ n1633)  &  (~ Ng4076) ) ;
 assign n5070 = ( Ng4057  &  (~ Ng4064)  &  n5068 ) ;
 assign n5071 = ( (~ Ng4057)  &  Ng4064  &  n5068 ) ;
 assign n5075 = ( n5076 ) | ( n5077 ) | ( n4492 ) ;
 assign n5074 = ( n5075  &  Pg35 ) ;
 assign n5076 = ( (~ Ng691)  &  Ng411 ) | ( (~ Ng691)  &  Ng424 ) | ( (~ Ng691)  &  (~ Ng417) ) ;
 assign n5077 = ( Ng691  &  Ng499 ) | ( Ng691  &  Ng518 ) ;
 assign n5079 = ( n667  &  Pg35 ) ;
 assign n5081 = ( n3943  &  Pg35 ) ;
 assign n5083 = ( Ng1442  &  (~ Ng1495) ) ;
 assign n5084 = ( Ng1437  &  n5045  &  n5083 ) ;
 assign n5085 = ( Ng1467  &  n5044  &  n5083 ) ;
 assign n5086 = ( Ng1454  &  n5043  &  n5083 ) ;
 assign n5088 = ( (~ Pg35) ) | ( (~ Ng1351) ) ;
 assign n5089 = ( Ng1099  &  (~ Ng1152) ) ;
 assign n5090 = ( Ng1094  &  n5048  &  n5089 ) ;
 assign n5091 = ( Ng1124  &  n5047  &  n5089 ) ;
 assign n5092 = ( Ng1111  &  n5046  &  n5089 ) ;
 assign n5093 = ( (~ Pg35) ) | ( (~ Ng1008) ) ;
 assign n5095 = ( Ng890  &  (~ Ng896)  &  (~ Ng862) ) ;
 assign n5094 = ( (~ Pg35) ) | ( n5095 ) ;
 assign n5096 = ( (~ Pg35) ) | ( (~ n5095) ) ;
 assign n5109 = ( (~ Ng311)  &  (~ Ng324) ) | ( (~ Ng311)  &  (~ Ng305) ) | ( Ng324  &  (~ Ng305) ) ;
 assign n5122 = ( Ng5084  &  Ng5092 ) ;
 assign n5130 = ( Ng1430  &  Ng1548 ) ;
 assign n5132 = ( Ng1484  &  n715  &  n5083 ) ;
 assign n5133 = ( Ng1087  &  Ng1205 ) ;
 assign n5135 = ( Ng1141  &  n557  &  n5089 ) ;
 assign n5136 = ( (~ Pg35) ) | ( n4492 ) ;
 assign n5137 = ( n4492  &  Pg35 ) ;
 assign n5139 = ( Pg8291  &  Ng218 ) ;
 assign n5140 = ( Pg17778  &  Pg14828  &  Pg12470  &  Pg17688 ) ;
 assign n5142 = ( (~ Pg17760) ) | ( (~ Pg17649) ) | ( (~ Pg14779) ) | ( (~ Pg12422) ) ;
 assign n5143 = ( Pg17739  &  Pg14738  &  Pg12350  &  Pg17607 ) ;
 assign n5145 = ( Pg17711  &  Pg14694  &  Pg12300  &  Pg17580 ) ;
 assign n5147 = ( (~ Pg17674) ) | ( (~ Pg17519) ) | ( (~ Pg14662) ) | ( (~ Pg12238) ) ;
 assign n5149 = ( (~ Pg16775) ) | ( (~ Pg16659) ) | ( (~ Pg13966) ) | ( (~ Pg11418) ) ;
 assign n5150 = ( (~ Pg16744) ) | ( (~ Pg16627) ) | ( (~ Pg13926) ) | ( (~ Pg11388) ) ;
 assign n5151 = ( (~ Pg16718) ) | ( (~ Pg16603) ) | ( (~ Pg13895) ) | ( (~ Pg11349) ) ;
 assign n5152 = ( n4382  &  Ng1554 ) ;
 assign n5154 = ( n4385  &  Ng1211 ) ;
 assign n5160 = ( n3232  &  n3230 ) | ( (~ n3232)  &  (~ n3230) ) ;
 assign n5162 = ( (~ n3285)  &  n3283 ) | ( n3285  &  (~ n3283) ) ;
 assign n5163 = ( n3340  &  n3338 ) | ( (~ n3340)  &  (~ n3338) ) ;
 assign n5165 = ( n3395  &  n3393 ) | ( (~ n3395)  &  (~ n3393) ) ;
 assign n5167 = ( (~ n5011)  &  n3447 ) | ( n5011  &  (~ n3447) ) ;
 assign n5168 = ( n3525  &  n3523 ) | ( (~ n3525)  &  (~ n3523) ) ;
 assign n5170 = ( n3577  &  n3575 ) | ( (~ n3577)  &  (~ n3575) ) ;
 assign n5172 = ( n3628  &  n3626 ) | ( (~ n3628)  &  (~ n3626) ) ;
 assign n5175 = ( Ng1319 ) | ( n667 ) ;
 assign n5174 = ( Ng1448  &  n5175 ) | ( (~ Ng1448)  &  (~ n5175) ) ;
 assign n5176 = ( Ng1300  &  n5175 ) | ( (~ Ng1300)  &  (~ n5175) ) ;
 assign n5177 = ( Ng1472  &  n5175 ) | ( (~ Ng1472)  &  (~ n5175) ) ;
 assign n5178 = ( Ng1478  &  n5175 ) | ( (~ Ng1478)  &  (~ n5175) ) ;
 assign n5180 = ( (~ n1411) ) | ( Ng976 ) ;
 assign n5179 = ( Ng1105  &  n5180 ) | ( (~ Ng1105)  &  (~ n5180) ) ;
 assign n5181 = ( Ng956  &  n5180 ) | ( (~ Ng956)  &  (~ n5180) ) ;
 assign n5182 = ( Ng1129  &  n5180 ) | ( (~ Ng1129)  &  (~ n5180) ) ;
 assign n5183 = ( Ng1135  &  n5180 ) | ( (~ Ng1135)  &  (~ n5180) ) ;
 assign Ng26965 = ( (~ Ng4534)  &  n3916 ) | ( Ng4534  &  (~ n3916) ) ;
 assign Ng26910 = ( (~ Ng862)  &  n4019 ) | ( Ng862  &  (~ n4019) ) ;
 assign Ng25697 = ( (~ Ng5084)  &  n4102 ) | ( Ng5084  &  (~ n4102) ) ;
 assign n5184 = ( (~ Ng246)  &  Ng269 ) | ( Ng246  &  (~ Ng269) ) ;
 assign n5185 = ( (~ Ng239)  &  Ng262 ) | ( Ng239  &  (~ Ng262) ) ;
 assign n5186 = ( (~ n1237)  &  n4178 ) | ( n1237  &  (~ n4178) ) ;
 assign Ng24260 = ( (~ Ng1430)  &  n4223 ) | ( Ng1430  &  (~ n4223) ) ;
 assign Ng24257 = ( (~ Ng1333)  &  n4225 ) | ( Ng1333  &  (~ n4225) ) ;
 assign Ng24244 = ( (~ Ng1087)  &  n4236 ) | ( Ng1087  &  (~ n4236) ) ;
 assign Ng24241 = ( (~ Ng990)  &  n4238 ) | ( Ng990  &  (~ n4238) ) ;
 assign n5189 = ( Pg9019  &  Ng4291 ) | ( (~ Pg9019)  &  (~ Ng4291) ) ;
 assign n5187 = ( Pg9019  &  n5189 ) | ( (~ Pg9019)  &  (~ n5189) ) ;
 assign n5192 = ( Pg8839  &  Ng4281 ) | ( (~ Pg8839)  &  (~ Ng4281) ) ;
 assign n5190 = ( Pg8839  &  n5192 ) | ( (~ Pg8839)  &  (~ n5192) ) ;
 assign n5193 = ( Pg35  &  (~ n5637) ) | ( (~ Ng2980)  &  (~ n5637) ) ;
 assign Ng34980 = ( (~ n5193) ) ;
 assign n5194 = ( (~ Pg35)  &  (~ Ng4366) ) | ( Pg35  &  n5649 ) | ( (~ Ng4366)  &  n5649 ) ;
 assign Ng34882 = ( (~ n5194) ) ;
 assign n5195 = ( Pg35  &  (~ n5651) ) | ( (~ Ng2955)  &  (~ n5651) ) ;
 assign Ng34808 = ( (~ n5195) ) ;
 assign n5196 = ( Pg35  &  (~ n5654) ) | ( (~ Ng2941)  &  (~ n5654) ) ;
 assign Ng34807 = ( (~ n5196) ) ;
 assign n5197 = ( Pg35  &  (~ n5657) ) | ( (~ Ng2927)  &  (~ n5657) ) ;
 assign Ng34806 = ( (~ n5197) ) ;
 assign n5198 = ( Pg35  &  (~ n5660) ) | ( (~ Ng2965)  &  (~ n5660) ) ;
 assign Ng34804 = ( (~ n5198) ) ;
 assign n5199 = ( Pg35  &  (~ n5663) ) | ( (~ Ng2917)  &  (~ n5663) ) ;
 assign Ng34803 = ( (~ n5199) ) ;
 assign n5200 = ( Pg35  &  (~ n5666) ) | ( (~ Ng2902)  &  (~ n5666) ) ;
 assign Ng34802 = ( (~ n5200) ) ;
 assign n5201 = ( Pg35  &  (~ n5669) ) | ( (~ Ng2970)  &  (~ n5669) ) ;
 assign Ng34801 = ( (~ n5201) ) ;
 assign n5202 = ( Ng55 ) | ( Ng2980 ) ;
 assign n5203 = ( (~ Pg35)  &  (~ Ng2886) ) | ( Pg35  &  (~ n5202) ) | ( (~ Ng2886)  &  (~ n5202) ) ;
 assign Ng34800 = ( (~ n5203) ) ;
 assign n5204 = ( (~ Pg44) ) | ( Ng2890 ) ;
 assign n5205 = ( (~ Pg35)  &  (~ Ng2873) ) | ( Pg35  &  (~ n5204) ) | ( (~ Ng2873)  &  (~ n5204) ) ;
 assign Ng34799 = ( (~ n5205) ) ;
 assign n5206 = ( Ng2946 ) | ( Ng2886 ) ;
 assign n5207 = ( (~ Pg35)  &  (~ Ng2878) ) | ( Pg35  &  (~ n5206) ) | ( (~ Ng2878)  &  (~ n5206) ) ;
 assign Ng34798 = ( (~ n5207) ) ;
 assign n5208 = ( (~ Pg91) ) | ( Ng2878 ) ;
 assign n5209 = ( (~ Pg35)  &  (~ Ng2882) ) | ( Pg35  &  (~ n5208) ) | ( (~ Ng2882)  &  (~ n5208) ) ;
 assign Ng34797 = ( (~ n5209) ) ;
 assign n5210 = ( Pg35  &  (~ n5676) ) | ( (~ Ng2898)  &  (~ n5676) ) ;
 assign Ng34796 = ( (~ n5210) ) ;
 assign n5211 = ( Ng2898 ) | ( (~ n4570) ) ;
 assign n5213 = ( (~ Pg35)  &  (~ Ng2864) ) | ( Pg35  &  (~ n5211) ) | ( (~ Ng2864)  &  (~ n5211) ) ;
 assign Ng34795 = ( (~ n5213) ) ;
 assign n5214 = ( Ng2864 ) | ( n4568 ) ;
 assign n5215 = ( (~ Pg35)  &  (~ Ng2856) ) | ( Pg35  &  (~ n5214) ) | ( (~ Ng2856)  &  (~ n5214) ) ;
 assign Ng34794 = ( (~ n5215) ) ;
 assign n5216 = ( Pg35  &  (~ n5681) ) | ( (~ Ng2848)  &  (~ n5681) ) ;
 assign Ng34793 = ( (~ n5216) ) ;
 assign n5217 = ( Pg35  &  (~ n5684) ) | ( (~ wire4433)  &  (~ n5684) ) ;
 assign Ng34792 = ( (~ n5217) ) ;
 assign n5218 = ( Ng4242 ) | ( Ng4300 ) ;
 assign n5219 = ( Pg35  &  (~ n5218) ) | ( (~ Pg35)  &  (~ Ng4297) ) | ( (~ n5218)  &  (~ Ng4297) ) ;
 assign Ng34735 = ( (~ n5219) ) ;
 assign n5220 = ( Ng4176 ) | ( Ng4072 ) ;
 assign n5221 = ( (~ Pg35)  &  (~ Ng4172) ) | ( Pg35  &  (~ n5220) ) | ( (~ Ng4172)  &  (~ n5220) ) ;
 assign Ng34734 = ( (~ n5221) ) ;
 assign n5222 = ( Ng1283 ) | ( Ng1277 ) ;
 assign n5223 = ( (~ Pg35)  &  (~ Ng1296) ) | ( Pg35  &  (~ n5222) ) | ( (~ Ng1296)  &  (~ n5222) ) ;
 assign Ng34730 = ( (~ n5223) ) ;
 assign n5224 = ( Ng933 ) | ( Ng939 ) ;
 assign n5225 = ( (~ Pg35)  &  (~ Ng952) ) | ( Pg35  &  (~ n5224) ) | ( (~ Ng952)  &  (~ n5224) ) ;
 assign Ng34727 = ( (~ n5225) ) ;
 assign n5226 = ( Ng534 ) | ( Ng301 ) ;
 assign n5227 = ( (~ Pg35)  &  (~ Ng542) ) | ( Pg35  &  (~ n5226) ) | ( (~ Ng542)  &  (~ n5226) ) ;
 assign Ng34723 = ( (~ n5227) ) ;
 assign n5228 = ( (~ Ng691) ) | ( Ng546 ) ;
 assign n5229 = ( (~ Pg35)  &  (~ Ng538) ) | ( Pg35  &  (~ n5228) ) | ( (~ Ng538)  &  (~ n5228) ) ;
 assign Ng34722 = ( (~ n5229) ) ;
 assign n5230 = ( Ng199 ) | ( Ng222 ) ;
 assign n5231 = ( (~ Pg35)  &  (~ wire4426) ) | ( Pg35  &  (~ n5230) ) | ( (~ wire4426)  &  (~ n5230) ) ;
 assign Ng34721 = ( (~ n5231) ) ;
 assign n5232 = ( (~ wire4435) ) | ( Ng550 ) ;
 assign n5233 = ( (~ Pg35)  &  (~ Ng534) ) | ( Pg35  &  (~ n5232) ) | ( (~ Ng534)  &  (~ n5232) ) ;
 assign Ng34720 = ( (~ n5233) ) ;
 assign n5234 = ( Pg35  &  (~ wire4433) ) | ( (~ Pg35)  &  (~ Ng37) ) | ( (~ wire4433)  &  (~ Ng37) ) ;
 assign Ng34614 = ( (~ n5234) ) ;
 assign Ng34602 = ( (~ n5705) ) ;
 assign Ng34601 = ( (~ n5706) ) ;
 assign n5237 = ( Pg35  &  (~ wire4426) ) | ( (~ Pg35)  &  (~ Ng550) ) | ( (~ wire4426)  &  (~ Ng550) ) ;
 assign Ng34598 = ( (~ n5237) ) ;
 assign n5238 = ( Ng4878  &  (~ n5710) ) | ( n1533  &  (~ n5710) ) | ( (~ Ng4843)  &  (~ n5710) ) ;
 assign Ng34466 = ( (~ n5238) ) ;
 assign n5239 = ( Ng4688  &  (~ n5712) ) | ( n1543  &  (~ n5712) ) | ( (~ Ng4653)  &  (~ n5712) ) ;
 assign Ng34462 = ( (~ n5239) ) ;
 assign n5240 = ( (~ Pg35)  &  (~ Ng4643) ) | ( Pg35  &  n5715 ) | ( (~ Ng4643)  &  n5715 ) ;
 assign Ng34459 = ( (~ n5240) ) ;
 assign n5241 = ( Pg35  &  n1622 ) | ( (~ Pg35)  &  (~ Ng446) ) | ( n1622  &  (~ Ng446) ) ;
 assign Ng34440 = ( (~ n5241) ) ;
 assign n5242 = ( (~ Pg35)  &  (~ Ng4961) ) | ( Pg35  &  n5735 ) | ( (~ Ng4961)  &  n5735 ) ;
 assign Ng34269 = ( (~ n5242) ) ;
 assign n5243 = ( (~ Pg35)  &  (~ Ng4950) ) | ( Pg35  &  n5738 ) | ( (~ Ng4950)  &  n5738 ) ;
 assign Ng34268 = ( (~ n5243) ) ;
 assign n5244 = ( (~ Pg35)  &  (~ Ng4894) ) | ( Pg35  &  n5741 ) | ( (~ Ng4894)  &  n5741 ) ;
 assign Ng34266 = ( (~ n5244) ) ;
 assign n5245 = ( (~ Pg35)  &  (~ Ng4771) ) | ( Pg35  &  n5744 ) | ( (~ Ng4771)  &  n5744 ) ;
 assign Ng34264 = ( (~ n5245) ) ;
 assign n5246 = ( (~ Pg35)  &  (~ Ng4760) ) | ( Pg35  &  n5747 ) | ( (~ Ng4760)  &  n5747 ) ;
 assign Ng34263 = ( (~ n5246) ) ;
 assign n5247 = ( (~ Pg35)  &  (~ Ng4704) ) | ( Pg35  &  n5750 ) | ( (~ Ng4704)  &  n5750 ) ;
 assign Ng34261 = ( (~ n5247) ) ;
 assign n5248 = ( (~ n4271)  &  n4270 ) | ( n4270  &  Ng4358 ) | ( (~ n4271)  &  (~ Ng4358) ) ;
 assign n5249 = ( (~ Pg35)  &  n5752 ) | ( n1220  &  n5752 ) | ( n4302  &  n5752 ) ;
 assign Ng34257 = ( (~ n5249) ) ;
 assign n5250 = ( (~ Pg35)  &  (~ Ng4369) ) | ( Pg35  &  n1677 ) | ( (~ Ng4369)  &  n1677 ) ;
 assign Ng34256 = ( (~ n5250) ) ;
 assign n5252 = ( wire4437  &  n5755 ) | ( n1222  &  n5755 ) | ( (~ Ng4581)  &  n5755 ) ;
 assign n5253 = ( (~ Pg35)  &  (~ Ng4492) ) | ( Pg35  &  n5756 ) | ( (~ Ng4492)  &  n5756 ) ;
 assign Ng34024 = ( (~ n5253) ) ;
 assign n5255 = ( n1222  &  n5757 ) | ( (~ Ng4581)  &  n5757 ) | ( n5757  &  Ng4575 ) ;
 assign n5256 = ( (~ Pg35)  &  (~ Ng4564) ) | ( Pg35  &  n5758 ) | ( (~ Ng4564)  &  n5758 ) ;
 assign Ng34023 = ( (~ n5256) ) ;
 assign n5259 = ( n1743  &  n4700 ) | ( n4696  &  n4700 ) | ( n4700  &  (~ Ng2643) ) ;
 assign n5257 = ( n5259  &  (~ n5580) ) | ( n1261  &  (~ Ng1589)  &  n5259 ) ;
 assign n5262 = ( n1768  &  n4710 ) | ( n4706  &  n4710 ) | ( n4710  &  (~ Ng2509) ) ;
 assign n5260 = ( n5262  &  (~ n5581) ) | ( n1264  &  Ng1589  &  n5262 ) ;
 assign n5265 = ( n1794  &  n4720 ) | ( n4716  &  n4720 ) | ( n4720  &  (~ Ng2375) ) ;
 assign n5263 = ( n5265  &  (~ n5582) ) | ( n1274  &  (~ Ng1589)  &  n5265 ) ;
 assign n5268 = ( n1819  &  n4730 ) | ( n4726  &  n4730 ) | ( n4730  &  (~ Ng2241) ) ;
 assign n5266 = ( n5268  &  (~ n5583) ) | ( n1270  &  Ng1589  &  n5268 ) ;
 assign n5271 = ( n1845  &  n4741 ) | ( n4737  &  n4741 ) | ( n4741  &  (~ Ng2084) ) ;
 assign n5269 = ( n5271  &  (~ n5584) ) | ( n1266  &  (~ Ng1246)  &  n5271 ) ;
 assign n5274 = ( n1870  &  n4751 ) | ( n4747  &  n4751 ) | ( n4751  &  (~ Ng1950) ) ;
 assign n5272 = ( n5274  &  (~ n5585) ) | ( n1268  &  Ng1246  &  n5274 ) ;
 assign n5277 = ( n1896  &  n4761 ) | ( n4757  &  n4761 ) | ( n4761  &  (~ Ng1816) ) ;
 assign n5275 = ( n5277  &  (~ n5586) ) | ( n1258  &  (~ Ng1246)  &  n5277 ) ;
 assign n5280 = ( n1921  &  n4771 ) | ( n4767  &  n4771 ) | ( n4771  &  (~ Ng1682) ) ;
 assign n5278 = ( n5280  &  (~ n5587) ) | ( n1272  &  Ng1246  &  n5280 ) ;
 assign n5282 = ( (~ Pg72)  &  n1222 ) | ( (~ Pg72)  &  Ng269 ) | ( n1222  &  Ng262 ) | ( Ng269  &  Ng262 ) ;
 assign n5281 = ( (~ Pg73)  &  n5282 ) | ( (~ Pg72)  &  Ng255  &  n5282 ) ;
 assign n5283 = ( (~ Pg35)  &  (~ wire4432) ) | ( Pg35  &  (~ n5281) ) | ( (~ wire4432)  &  (~ n5281) ) ;
 assign Ng33963 = ( (~ n5283) ) ;
 assign n5286 = ( Pg73 ) | ( (~ Pg72) ) | ( Ng239 ) ;
 assign n5287 = ( Ng246 ) | ( n1222 ) ;
 assign n5285 = ( (~ Pg72)  &  Ng232 ) | ( Pg72  &  Ng225 ) | ( Ng232  &  Ng225 ) ;
 assign n5284 = ( (~ Pg73)  &  n5286  &  n5287 ) | ( n5286  &  n5287  &  n5285 ) ;
 assign n5288 = ( (~ Pg35)  &  (~ Ng479) ) | ( Pg35  &  (~ n5284) ) | ( (~ Ng479)  &  (~ n5284) ) ;
 assign Ng33962 = ( (~ n5288) ) ;
 assign n5290 = ( (~ n1097)  &  (~ Ng5644) ) | ( n1097  &  n4783 ) | ( (~ Ng5644)  &  n4783 ) ;
 assign n5291 = ( Pg35  &  (~ n5775) ) | ( (~ Ng5703)  &  (~ n5775) ) ;
 assign Ng33621 = ( (~ n5291) ) ;
 assign n5292 = ( (~ Pg35)  &  (~ Ng4552) ) | ( Pg35  &  (~ n5255) ) | ( (~ Ng4552)  &  (~ n5255) ) ;
 assign Ng33617 = ( (~ n5292) ) ;
 assign n5293 = ( (~ Pg35)  &  (~ Ng4515) ) | ( Pg35  &  (~ n5252) ) | ( (~ Ng4515)  &  (~ n5252) ) ;
 assign Ng33616 = ( (~ n5293) ) ;
 assign n5295 = ( n4276  &  Ng2667 ) | ( Ng2667  &  Ng2661 ) | ( n4276  &  (~ Ng2661) ) ;
 assign n5296 = ( n4699  &  (~ Ng2667) ) | ( (~ n4699)  &  (~ Ng2661) ) | ( (~ Ng2667)  &  (~ Ng2661) ) ;
 assign Ng33604 = ( (~ n5296) ) ;
 assign n5297 = ( n4699  &  (~ Ng2648) ) | ( (~ n4699)  &  (~ Ng2643) ) | ( (~ Ng2648)  &  (~ Ng2643) ) ;
 assign Ng33603 = ( (~ n5297) ) ;
 assign n5299 = ( n4277  &  (~ Ng2533) ) | ( n4277  &  Ng2527 ) | ( Ng2533  &  Ng2527 ) ;
 assign n5300 = ( n4709  &  (~ Ng2533) ) | ( (~ n4709)  &  (~ Ng2527) ) | ( (~ Ng2533)  &  (~ Ng2527) ) ;
 assign Ng33596 = ( (~ n5300) ) ;
 assign n5301 = ( (~ Ng2514)  &  n4709 ) | ( (~ Ng2514)  &  (~ Ng2509) ) | ( (~ n4709)  &  (~ Ng2509) ) ;
 assign Ng33595 = ( (~ n5301) ) ;
 assign n5303 = ( n4279  &  Ng2399 ) | ( Ng2399  &  Ng2393 ) | ( n4279  &  (~ Ng2393) ) ;
 assign n5304 = ( n4719  &  (~ Ng2399) ) | ( (~ n4719)  &  (~ Ng2393) ) | ( (~ Ng2399)  &  (~ Ng2393) ) ;
 assign Ng33588 = ( (~ n5304) ) ;
 assign n5305 = ( n4719  &  (~ Ng2380) ) | ( (~ n4719)  &  (~ Ng2375) ) | ( (~ Ng2380)  &  (~ Ng2375) ) ;
 assign Ng33587 = ( (~ n5305) ) ;
 assign n5307 = ( n4280  &  Ng2265 ) | ( Ng2265  &  Ng2259 ) | ( n4280  &  (~ Ng2259) ) ;
 assign n5308 = ( n4729  &  (~ Ng2265) ) | ( (~ n4729)  &  (~ Ng2259) ) | ( (~ Ng2265)  &  (~ Ng2259) ) ;
 assign Ng33580 = ( (~ n5308) ) ;
 assign n5309 = ( n4729  &  (~ Ng2246) ) | ( (~ n4729)  &  (~ Ng2241) ) | ( (~ Ng2246)  &  (~ Ng2241) ) ;
 assign Ng33579 = ( (~ n5309) ) ;
 assign n5311 = ( n4281  &  (~ Ng2108) ) | ( n4281  &  Ng2102 ) | ( Ng2108  &  Ng2102 ) ;
 assign n5312 = ( n4740  &  (~ Ng2108) ) | ( (~ n4740)  &  (~ Ng2102) ) | ( (~ Ng2108)  &  (~ Ng2102) ) ;
 assign Ng33572 = ( (~ n5312) ) ;
 assign n5313 = ( (~ Ng2089)  &  n4740 ) | ( (~ Ng2089)  &  (~ Ng2084) ) | ( (~ n4740)  &  (~ Ng2084) ) ;
 assign Ng33571 = ( (~ n5313) ) ;
 assign n5315 = ( n4283  &  (~ Ng1974) ) | ( n4283  &  Ng1968 ) | ( Ng1974  &  Ng1968 ) ;
 assign n5316 = ( n4750  &  (~ Ng1974) ) | ( (~ n4750)  &  (~ Ng1968) ) | ( (~ Ng1974)  &  (~ Ng1968) ) ;
 assign Ng33564 = ( (~ n5316) ) ;
 assign n5317 = ( (~ Ng1955)  &  n4750 ) | ( (~ Ng1955)  &  (~ Ng1950) ) | ( (~ n4750)  &  (~ Ng1950) ) ;
 assign Ng33563 = ( (~ n5317) ) ;
 assign n5319 = ( n4285  &  Ng1840 ) | ( Ng1840  &  Ng1834 ) | ( n4285  &  (~ Ng1834) ) ;
 assign n5320 = ( n4760  &  (~ Ng1840) ) | ( (~ n4760)  &  (~ Ng1834) ) | ( (~ Ng1840)  &  (~ Ng1834) ) ;
 assign Ng33556 = ( (~ n5320) ) ;
 assign n5321 = ( (~ Ng1821)  &  n4760 ) | ( (~ Ng1821)  &  (~ Ng1816) ) | ( (~ n4760)  &  (~ Ng1816) ) ;
 assign Ng33555 = ( (~ n5321) ) ;
 assign n5323 = ( n4286  &  Ng1706 ) | ( Ng1706  &  Ng1700 ) | ( n4286  &  (~ Ng1700) ) ;
 assign n5324 = ( n4770  &  (~ Ng1706) ) | ( (~ n4770)  &  (~ Ng1700) ) | ( (~ Ng1706)  &  (~ Ng1700) ) ;
 assign Ng33548 = ( (~ n5324) ) ;
 assign n5325 = ( (~ Ng1687)  &  n4770 ) | ( (~ Ng1687)  &  (~ Ng1682) ) | ( (~ n4770)  &  (~ Ng1682) ) ;
 assign Ng33547 = ( (~ n5325) ) ;
 assign n5326 = ( (~ Pg35)  &  n5793 ) | ( n4664  &  n5793 ) | ( (~ Ng142)  &  n5793 ) ;
 assign Ng33537 = ( (~ n5326) ) ;
 assign n5327 = ( n4842  &  Ng5041 ) | ( n4842  &  n4845 ) | ( (~ Ng5041)  &  n4845 ) ;
 assign n5328 = ( n4840  &  Ng5033 ) | ( n4840  &  n4844 ) | ( (~ Ng5033)  &  n4844 ) ;
 assign n5329 = ( Ng283  &  (~ n5819) ) | ( n3904  &  (~ n5819) ) | ( (~ Ng287)  &  (~ n5819) ) ;
 assign Ng31865 = ( (~ n5329) ) ;
 assign n5330 = ( Pg35  &  n2861 ) | ( (~ Pg35)  &  (~ Ng4122) ) | ( n2861  &  (~ Ng4122) ) ;
 assign Ng30457 = ( (~ n5330) ) ;
 assign n5331 = ( n3048  &  (~ Ng2675) ) | ( (~ n3048)  &  (~ Ng2681) ) | ( (~ Ng2675)  &  (~ Ng2681) ) ;
 assign Ng30386 = ( (~ n5331) ) ;
 assign n5332 = ( n3060  &  (~ Ng2541) ) | ( (~ n3060)  &  (~ Ng2547) ) | ( (~ Ng2541)  &  (~ Ng2547) ) ;
 assign Ng30381 = ( (~ n5332) ) ;
 assign n5333 = ( n3072  &  (~ Ng2407) ) | ( (~ n3072)  &  (~ Ng2413) ) | ( (~ Ng2407)  &  (~ Ng2413) ) ;
 assign Ng30376 = ( (~ n5333) ) ;
 assign n5334 = ( n3084  &  (~ Ng2273) ) | ( (~ n3084)  &  (~ Ng2279) ) | ( (~ Ng2273)  &  (~ Ng2279) ) ;
 assign Ng30371 = ( (~ n5334) ) ;
 assign n5335 = ( n3096  &  (~ Ng2116) ) | ( (~ n3096)  &  (~ Ng2122) ) | ( (~ Ng2116)  &  (~ Ng2122) ) ;
 assign Ng30366 = ( (~ n5335) ) ;
 assign n5336 = ( n3108  &  (~ Ng1982) ) | ( (~ n3108)  &  (~ Ng1988) ) | ( (~ Ng1982)  &  (~ Ng1988) ) ;
 assign Ng30361 = ( (~ n5336) ) ;
 assign n5337 = ( n3120  &  (~ Ng1848) ) | ( (~ n3120)  &  (~ Ng1854) ) | ( (~ Ng1848)  &  (~ Ng1854) ) ;
 assign Ng30356 = ( (~ n5337) ) ;
 assign n5338 = ( n3132  &  (~ Ng1714) ) | ( (~ n3132)  &  (~ Ng1720) ) | ( (~ Ng1714)  &  (~ Ng1720) ) ;
 assign Ng30351 = ( (~ n5338) ) ;
 assign n5339 = ( (~ n4288)  &  n4287 ) | ( n4287  &  Ng1413 ) | ( (~ n4288)  &  (~ Ng1413) ) ;
 assign n5340 = ( (~ Pg35)  &  n5879 ) | ( n923  &  n5879 ) | ( n4355  &  n5879 ) ;
 assign Ng30346 = ( (~ n5340) ) ;
 assign n5341 = ( (~ n4290)  &  n4289 ) | ( n4289  &  Ng1070 ) | ( (~ n4290)  &  (~ Ng1070) ) ;
 assign n5342 = ( (~ Pg35)  &  n5880 ) | ( n330  &  n5880 ) | ( n4357  &  n5880 ) ;
 assign Ng30340 = ( (~ n5342) ) ;
 assign n5343 = ( n3188  &  (~ Ng6513) ) | ( (~ n3188)  &  (~ Ng6519) ) | ( (~ Ng6513)  &  (~ Ng6519) ) ;
 assign Ng29306 = ( (~ n5343) ) ;
 assign n5344 = ( n3242  &  (~ Ng6167) ) | ( (~ n3242)  &  (~ Ng6173) ) | ( (~ Ng6167)  &  (~ Ng6173) ) ;
 assign Ng29300 = ( (~ n5344) ) ;
 assign n5345 = ( n3295  &  (~ Ng5821) ) | ( (~ n3295)  &  (~ Ng5827) ) | ( (~ Ng5821)  &  (~ Ng5827) ) ;
 assign Ng29294 = ( (~ n5345) ) ;
 assign n5346 = ( n3350  &  (~ Ng5475) ) | ( (~ n3350)  &  (~ Ng5481) ) | ( (~ Ng5475)  &  (~ Ng5481) ) ;
 assign Ng29288 = ( (~ n5346) ) ;
 assign n5347 = ( n3405  &  (~ Ng5128) ) | ( (~ n3405)  &  (~ Ng5134) ) | ( (~ Ng5128)  &  (~ Ng5134) ) ;
 assign Ng29282 = ( (~ n5347) ) ;
 assign n5348 = ( (~ n3459)  &  n4359  &  n4564 ) | ( (~ n3459)  &  n4564  &  n4777 ) ;
 assign n5350 = ( (~ n3468)  &  n4360  &  n4559 ) | ( (~ n3468)  &  n4559  &  n4776 ) ;
 assign n5352 = ( n3480  &  (~ Ng3821) ) | ( (~ n3480)  &  (~ Ng3827) ) | ( (~ Ng3821)  &  (~ Ng3827) ) ;
 assign Ng29271 = ( (~ n5352) ) ;
 assign n5353 = ( n3535  &  (~ Ng3470) ) | ( (~ n3535)  &  (~ Ng3476) ) | ( (~ Ng3470)  &  (~ Ng3476) ) ;
 assign Ng29265 = ( (~ n5353) ) ;
 assign n5354 = ( n3586  &  (~ Ng3119) ) | ( (~ n3586)  &  (~ Ng3125) ) | ( (~ Ng3119)  &  (~ Ng3125) ) ;
 assign Ng29259 = ( (~ n5354) ) ;
 assign n5355 = ( Pg35  &  (~ n5953) ) | ( (~ Ng1478)  &  (~ n5953) ) ;
 assign Ng29239 = ( (~ n5355) ) ;
 assign n5357 = ( (~ Ng1489)  &  (~ Ng1442) ) ;
 assign n5356 = ( n5176  &  n715  &  Ng1484 ) | ( n5176  &  n715  &  n5357 ) ;
 assign n5358 = ( Pg35  &  (~ n5958) ) | ( (~ Ng1448)  &  (~ n5958) ) ;
 assign Ng29237 = ( (~ n5358) ) ;
 assign n5359 = ( Pg35  &  (~ n5962) ) | ( (~ Ng1442)  &  (~ n5962) ) ;
 assign Ng29236 = ( (~ n5359) ) ;
 assign n5360 = ( Pg35  &  (~ n5966) ) | ( (~ Ng1135)  &  (~ n5966) ) ;
 assign Ng29234 = ( (~ n5360) ) ;
 assign n5362 = ( (~ Ng1146)  &  (~ Ng1099) ) ;
 assign n5361 = ( n5181  &  n557  &  Ng1141 ) | ( n5181  &  n557  &  n5362 ) ;
 assign n5363 = ( Pg35  &  (~ n5971) ) | ( (~ Ng1105)  &  (~ n5971) ) ;
 assign Ng29232 = ( (~ n5363) ) ;
 assign n5364 = ( Pg35  &  (~ n5975) ) | ( (~ Ng1099)  &  (~ n5975) ) ;
 assign Ng29231 = ( (~ n5364) ) ;
 assign n5365 = ( (~ Pg35)  &  n5985 ) | ( n4851  &  n5985 ) | ( n4853  &  n5985 ) ;
 assign Ng28092 = ( (~ n5365) ) ;
 assign n5366 = ( (~ Pg35)  &  n5986 ) | ( n4852  &  n5986 ) | ( n4854  &  n5986 ) ;
 assign Ng28091 = ( (~ n5366) ) ;
 assign n5367 = ( (~ Ng4521)  &  n5988 ) | ( Pg35  &  n5988  &  n5987 ) ;
 assign Ng28082 = ( (~ n5367) ) ;
 assign n5368 = ( Pg35  &  n5989 ) | ( (~ Ng2841)  &  n5989 ) ;
 assign Ng28081 = ( (~ n5368) ) ;
 assign n5369 = ( n3858  &  (~ Ng4112) ) | ( (~ n3858)  &  (~ Ng4145) ) | ( (~ Ng4112)  &  (~ Ng4145) ) ;
 assign Ng28071 = ( (~ n5369) ) ;
 assign n5370 = ( (~ Ng728)  &  (~ Ng661) ) | ( (~ Ng728)  &  n5074 ) | ( (~ Ng661)  &  (~ n5074) ) ;
 assign Ng28054 = ( (~ n5370) ) ;
 assign n5371 = ( (~ Ng661)  &  (~ Ng718) ) | ( (~ Ng661)  &  n5074 ) | ( (~ Ng718)  &  (~ n5074) ) ;
 assign Ng28052 = ( (~ n5371) ) ;
 assign n5372 = ( (~ Ng718)  &  (~ Ng655) ) | ( (~ Ng718)  &  n5074 ) | ( (~ Ng655)  &  (~ n5074) ) ;
 assign Ng28051 = ( (~ n5372) ) ;
 assign n5373 = ( (~ Ng655)  &  (~ Ng650) ) | ( (~ Ng655)  &  n5074 ) | ( (~ Ng650)  &  (~ n5074) ) ;
 assign Ng28050 = ( (~ n5373) ) ;
 assign n5374 = ( (~ Pg35)  &  (~ wire4435) ) | ( Pg35  &  n4364 ) | ( (~ wire4435)  &  n4364 ) ;
 assign Ng28048 = ( (~ n5374) ) ;
 assign n5375 = ( (~ Ng681)  &  (~ Ng645) ) | ( (~ Ng681)  &  n5074 ) | ( (~ Ng645)  &  (~ n5074) ) ;
 assign Ng28047 = ( (~ n5375) ) ;
 assign n5376 = ( Pg35  &  n3915 ) | ( (~ Pg35)  &  (~ Ng4512) ) | ( n3915  &  (~ Ng4512) ) ;
 assign Ng26971 = ( (~ n5376) ) ;
 assign n5377 = ( Pg35  &  (~ Ng4473) ) | ( (~ Pg35)  &  (~ Ng4459) ) | ( (~ Ng4473)  &  (~ Ng4459) ) ;
 assign Ng26970 = ( (~ n5377) ) ;
 assign n5378 = ( (~ Pg35)  &  (~ Ng4462) ) | ( Pg35  &  n5995 ) | ( (~ Ng4462)  &  n5995 ) ;
 assign Ng26969 = ( (~ n5378) ) ;
 assign n5379 = ( (~ Pg6749)  &  Pg35 ) | ( (~ Pg6749)  &  (~ Ng4558) ) | ( (~ Pg35)  &  (~ Ng4558) ) ;
 assign Ng26968 = ( (~ n5379) ) ;
 assign n5380 = ( (~ Pg6750)  &  Pg35 ) | ( (~ Pg6750)  &  (~ Ng4561) ) | ( (~ Pg35)  &  (~ Ng4561) ) ;
 assign Ng26967 = ( (~ n5380) ) ;
 assign n5381 = ( (~ Pg6748)  &  Pg35 ) | ( (~ Pg6748)  &  (~ Ng4555) ) | ( (~ Pg35)  &  (~ Ng4555) ) ;
 assign Ng26966 = ( (~ n5381) ) ;
 assign n5382 = ( (~ Pg6750)  &  Pg35 ) | ( (~ Pg6750)  &  (~ Ng4489) ) | ( (~ Pg35)  &  (~ Ng4489) ) ;
 assign Ng26963 = ( (~ n5382) ) ;
 assign n5383 = ( (~ Pg6749)  &  Pg35 ) | ( (~ Pg6749)  &  (~ Ng4486) ) | ( (~ Pg35)  &  (~ Ng4486) ) ;
 assign Ng26962 = ( (~ n5383) ) ;
 assign n5384 = ( (~ Pg6748)  &  Pg35 ) | ( (~ Pg6748)  &  (~ Ng4483) ) | ( (~ Pg35)  &  (~ Ng4483) ) ;
 assign Ng26961 = ( (~ n5384) ) ;
 assign n5385 = ( Pg35  &  n5828 ) | ( (~ Pg35)  &  (~ Ng4153) ) | ( n5828  &  (~ Ng4153) ) ;
 assign Ng26940 = ( (~ n5385) ) ;
 assign n5386 = ( (~ Pg35)  &  (~ Ng4104) ) | ( Pg35  &  n5825 ) | ( (~ Ng4104)  &  n5825 ) ;
 assign Ng26939 = ( (~ n5386) ) ;
 assign n5387 = ( Pg35  &  n6001 ) | ( (~ Ng2841)  &  n6001 ) ;
 assign Ng26937 = ( (~ n5387) ) ;
 assign n5388 = ( Pg35  &  n4371 ) | ( (~ Pg35)  &  (~ Ng1532) ) | ( n4371  &  (~ Ng1532) ) ;
 assign Ng26925 = ( (~ n5388) ) ;
 assign n5389 = ( (~ Pg35)  &  n6002 ) | ( n4374  &  n6002 ) | ( Ng1322  &  n6002 ) ;
 assign Ng26921 = ( (~ n5389) ) ;
 assign n5390 = ( Pg35  &  n4376 ) | ( (~ Pg35)  &  (~ Ng1189) ) | ( n4376  &  (~ Ng1189) ) ;
 assign Ng26918 = ( (~ n5390) ) ;
 assign n5391 = ( (~ Pg35)  &  (~ Ng890) ) | ( Pg35  &  n6003 ) | ( (~ Ng890)  &  n6003 ) ;
 assign Ng26909 = ( (~ n5391) ) ;
 assign n5392 = ( n6004  &  Ng812 ) | ( n6004  &  n4248  &  Ng843 ) ;
 assign n5393 = ( (~ Ng753)  &  (~ Ng732) ) | ( (~ Ng732)  &  n6005 ) | ( (~ Ng753)  &  (~ n6005) ) ;
 assign Ng26897 = ( (~ n5393) ) ;
 assign n5394 = ( (~ Ng528)  &  n5056  &  (~ n6007) ) | ( n5056  &  n5057  &  (~ n6007) ) ;
 assign n5396 = ( (~ Pg35)  &  (~ Ng518) ) | ( Pg35  &  (~ n5394) ) | ( (~ Ng518)  &  (~ n5394) ) ;
 assign Ng26894 = ( (~ n5396) ) ;
 assign n5397 = ( Pg35  &  Ng333 ) | ( Pg35  &  Ng355 ) ;
 assign n5398 = ( Pg35  &  Ng351 ) | ( Pg35  &  (~ n5397) ) | ( (~ Ng351)  &  (~ n5397) ) ;
 assign Ng26892 = ( (~ n5398) ) ;
 assign n5399 = ( Pg35  &  n6010 ) | ( (~ Ng347)  &  n6010 ) ;
 assign Ng26891 = ( (~ n5399) ) ;
 assign n5400 = ( Pg35  &  Ng347 ) | ( (~ Pg35)  &  (~ Ng333) ) | ( Ng347  &  (~ Ng333) ) ;
 assign Ng26890 = ( (~ n5400) ) ;
 assign n5402 = ( Pg35  &  n6011 ) | ( (~ wire4436)  &  n6011 ) ;
 assign Ng26889 = ( (~ n5402) ) ;
 assign n5403 = ( (~ Pg35)  &  (~ wire4431) ) | ( Pg35  &  (~ Ng316) ) | ( (~ wire4431)  &  (~ Ng316) ) ;
 assign Ng26888 = ( (~ n5403) ) ;
 assign n5404 = ( Pg35  &  n4055 ) | ( (~ Pg35)  &  (~ Ng336) ) | ( n4055  &  (~ Ng336) ) ;
 assign Ng26887 = ( (~ n5404) ) ;
 assign n5405 = ( Pg35  &  n4064 ) | ( (~ Pg35)  &  (~ Ng316) ) | ( n4064  &  (~ Ng316) ) ;
 assign Ng26882 = ( (~ n5405) ) ;
 assign n5406 = ( (~ Pg6744)  &  Pg35 ) | ( (~ Pg6744)  &  (~ Ng305) ) | ( (~ Pg35)  &  (~ Ng305) ) ;
 assign Ng26881 = ( (~ n5406) ) ;
 assign n5407 = ( (~ Ng6541)  &  (~ n4886) ) | ( (~ Ng6541)  &  (~ Ng6505) ) | ( n4886  &  (~ Ng6505) ) ;
 assign Ng25764 = ( (~ n5407) ) ;
 assign n5409 = ( n4291  &  Ng6533 ) | ( Ng6533  &  Ng6527 ) | ( n4291  &  (~ Ng6527) ) ;
 assign n5410 = ( n4886  &  (~ Ng6533) ) | ( (~ n4886)  &  (~ Ng6527) ) | ( (~ Ng6533)  &  (~ Ng6527) ) ;
 assign Ng25762 = ( (~ n5410) ) ;
 assign n5411 = ( (~ Pg9817)  &  Ng6444 ) | ( (~ Pg9817)  &  Pg9743  &  (~ Ng6494) ) ;
 assign n5413 = ( Pg35  &  (~ n5411) ) | ( (~ Pg35)  &  (~ Ng6494) ) | ( (~ n5411)  &  (~ Ng6494) ) ;
 assign Ng25758 = ( (~ n5413) ) ;
 assign n5414 = ( (~ Pg35)  &  (~ Ng6444) ) | ( Pg35  &  (~ Ng6727) ) | ( (~ Ng6444)  &  (~ Ng6727) ) ;
 assign Ng25757 = ( (~ n5414) ) ;
 assign n5415 = ( (~ Ng6195)  &  (~ n4894) ) | ( (~ Ng6195)  &  (~ Ng6159) ) | ( n4894  &  (~ Ng6159) ) ;
 assign Ng25750 = ( (~ n5415) ) ;
 assign n5417 = ( n4292  &  Ng6187 ) | ( Ng6187  &  Ng6181 ) | ( n4292  &  (~ Ng6181) ) ;
 assign n5418 = ( n4894  &  (~ Ng6187) ) | ( (~ n4894)  &  (~ Ng6181) ) | ( (~ Ng6187)  &  (~ Ng6181) ) ;
 assign Ng25748 = ( (~ n5418) ) ;
 assign n5419 = ( (~ Pg9741)  &  Ng6098 ) | ( (~ Pg9741)  &  Pg9682  &  (~ Ng6148) ) ;
 assign n5421 = ( Pg35  &  (~ n5419) ) | ( (~ Pg35)  &  (~ Ng6148) ) | ( (~ n5419)  &  (~ Ng6148) ) ;
 assign Ng25744 = ( (~ n5421) ) ;
 assign n5422 = ( (~ Pg35)  &  (~ Ng6098) ) | ( Pg35  &  (~ Ng6381) ) | ( (~ Ng6098)  &  (~ Ng6381) ) ;
 assign Ng25743 = ( (~ n5422) ) ;
 assign n5423 = ( (~ Ng5849)  &  (~ n4901) ) | ( (~ Ng5849)  &  (~ Ng5813) ) | ( n4901  &  (~ Ng5813) ) ;
 assign Ng25736 = ( (~ n5423) ) ;
 assign n5425 = ( n4293  &  Ng5841 ) | ( Ng5841  &  Ng5835 ) | ( n4293  &  (~ Ng5835) ) ;
 assign n5426 = ( n4901  &  (~ Ng5841) ) | ( (~ n4901)  &  (~ Ng5835) ) | ( (~ Ng5841)  &  (~ Ng5835) ) ;
 assign Ng25734 = ( (~ n5426) ) ;
 assign n5427 = ( (~ Pg9680)  &  Ng5752 ) | ( (~ Pg9680)  &  Pg9617  &  (~ Ng5802) ) ;
 assign n5429 = ( Pg35  &  (~ n5427) ) | ( (~ Pg35)  &  (~ Ng5802) ) | ( (~ n5427)  &  (~ Ng5802) ) ;
 assign Ng25730 = ( (~ n5429) ) ;
 assign n5430 = ( (~ Pg35)  &  (~ Ng5752) ) | ( Pg35  &  (~ Ng6035) ) | ( (~ Ng5752)  &  (~ Ng6035) ) ;
 assign Ng25729 = ( (~ n5430) ) ;
 assign n5431 = ( (~ Ng5503)  &  (~ n4908) ) | ( (~ Ng5503)  &  (~ Ng5467) ) | ( n4908  &  (~ Ng5467) ) ;
 assign Ng25722 = ( (~ n5431) ) ;
 assign n5433 = ( n4294  &  Ng5495 ) | ( Ng5495  &  Ng5489 ) | ( n4294  &  (~ Ng5489) ) ;
 assign n5434 = ( n4908  &  (~ Ng5495) ) | ( (~ n4908)  &  (~ Ng5489) ) | ( (~ Ng5495)  &  (~ Ng5489) ) ;
 assign Ng25720 = ( (~ n5434) ) ;
 assign n5435 = ( (~ Pg9615)  &  Ng5406 ) | ( (~ Pg9615)  &  Pg9555  &  (~ Ng5456) ) ;
 assign n5437 = ( Pg35  &  (~ n5435) ) | ( (~ Pg35)  &  (~ Ng5456) ) | ( (~ n5435)  &  (~ Ng5456) ) ;
 assign Ng25716 = ( (~ n5437) ) ;
 assign n5438 = ( (~ Pg35)  &  (~ Ng5406) ) | ( Pg35  &  (~ Ng5689) ) | ( (~ Ng5406)  &  (~ Ng5689) ) ;
 assign Ng25715 = ( (~ n5438) ) ;
 assign n5439 = ( (~ Ng5156)  &  n4092 ) | ( (~ Ng5156)  &  (~ Ng5120) ) | ( (~ n4092)  &  (~ Ng5120) ) ;
 assign Ng25708 = ( (~ n5439) ) ;
 assign n5441 = ( n4295  &  Ng5148 ) | ( Ng5148  &  Ng5142 ) | ( n4295  &  (~ Ng5142) ) ;
 assign n5442 = ( (~ n4092)  &  (~ Ng5148) ) | ( n4092  &  (~ Ng5142) ) | ( (~ Ng5148)  &  (~ Ng5142) ) ;
 assign Ng25706 = ( (~ n5442) ) ;
 assign n5443 = ( (~ Pg9497)  &  Ng5022 ) | ( Pg9553  &  (~ Pg9497)  &  (~ Ng5112) ) ;
 assign n5445 = ( Pg35  &  (~ n5443) ) | ( (~ Pg35)  &  (~ Ng5112) ) | ( (~ n5443)  &  (~ Ng5112) ) ;
 assign Ng25703 = ( (~ n5445) ) ;
 assign n5446 = ( (~ Pg9553)  &  Ng5062 ) | ( (~ Pg9553)  &  Pg9497  &  (~ Ng5109) ) ;
 assign n5448 = ( Pg35  &  (~ n5446) ) | ( (~ Pg35)  &  (~ Ng5109) ) | ( (~ n5446)  &  (~ Ng5109) ) ;
 assign Ng25702 = ( (~ n5448) ) ;
 assign n5449 = ( Pg35  &  (~ wire4415) ) | ( (~ Pg35)  &  (~ Ng5062) ) | ( (~ wire4415)  &  (~ Ng5062) ) ;
 assign Ng25701 = ( (~ n5449) ) ;
 assign n5450 = ( Ng5073  &  Ng5069 ) | ( Ng5069  &  Ng5084 ) | ( Ng5073  &  (~ Ng5084) ) ;
 assign n5451 = ( n3474  &  (~ n6023) ) | ( (~ Ng4057)  &  (~ n6023) ) | ( Ng4064  &  (~ n6023) ) ;
 assign Ng25686 = ( (~ n5451) ) ;
 assign n5452 = ( (~ Ng3849)  &  (~ n4922) ) | ( (~ Ng3849)  &  (~ Ng3813) ) | ( n4922  &  (~ Ng3813) ) ;
 assign Ng25684 = ( (~ n5452) ) ;
 assign n5454 = ( n4296  &  Ng3841 ) | ( Ng3841  &  Ng3835 ) | ( n4296  &  (~ Ng3835) ) ;
 assign n5455 = ( n4922  &  (~ Ng3841) ) | ( (~ n4922)  &  (~ Ng3835) ) | ( (~ Ng3841)  &  (~ Ng3835) ) ;
 assign Ng25682 = ( (~ n5455) ) ;
 assign n5456 = ( (~ Pg8398)  &  Ng3752 ) | ( (~ Pg8398)  &  Pg8344  &  (~ Ng3802) ) ;
 assign n5458 = ( Pg35  &  (~ n5456) ) | ( (~ Pg35)  &  (~ Ng3802) ) | ( (~ n5456)  &  (~ Ng3802) ) ;
 assign Ng25678 = ( (~ n5458) ) ;
 assign n5459 = ( (~ Pg35)  &  (~ Ng3752) ) | ( Pg35  &  (~ Ng4040) ) | ( (~ Ng3752)  &  (~ Ng4040) ) ;
 assign Ng25677 = ( (~ n5459) ) ;
 assign n5460 = ( (~ Ng3498)  &  (~ n4928) ) | ( (~ Ng3498)  &  (~ Ng3462) ) | ( n4928  &  (~ Ng3462) ) ;
 assign Ng25670 = ( (~ n5460) ) ;
 assign n5462 = ( n4297  &  Ng3490 ) | ( Ng3490  &  Ng3484 ) | ( n4297  &  (~ Ng3484) ) ;
 assign n5463 = ( n4928  &  (~ Ng3490) ) | ( (~ n4928)  &  (~ Ng3484) ) | ( (~ Ng3490)  &  (~ Ng3484) ) ;
 assign Ng25668 = ( (~ n5463) ) ;
 assign n5464 = ( (~ Pg8342)  &  Ng3401 ) | ( (~ Pg8342)  &  Pg8279  &  (~ Ng3451) ) ;
 assign n5466 = ( Pg35  &  (~ n5464) ) | ( (~ Pg35)  &  (~ Ng3451) ) | ( (~ n5464)  &  (~ Ng3451) ) ;
 assign Ng25664 = ( (~ n5466) ) ;
 assign n5467 = ( (~ Pg35)  &  (~ Ng3401) ) | ( Pg35  &  (~ Ng3689) ) | ( (~ Ng3401)  &  (~ Ng3689) ) ;
 assign Ng25663 = ( (~ n5467) ) ;
 assign n5468 = ( (~ Ng3147)  &  (~ n4934) ) | ( (~ Ng3147)  &  (~ Ng3111) ) | ( n4934  &  (~ Ng3111) ) ;
 assign Ng25656 = ( (~ n5468) ) ;
 assign n5470 = ( n4298  &  Ng3139 ) | ( Ng3139  &  Ng3133 ) | ( n4298  &  (~ Ng3133) ) ;
 assign n5471 = ( n4934  &  (~ Ng3139) ) | ( (~ n4934)  &  (~ Ng3133) ) | ( (~ Ng3139)  &  (~ Ng3133) ) ;
 assign Ng25654 = ( (~ n5471) ) ;
 assign n5472 = ( (~ Pg8277)  &  Ng3050 ) | ( (~ Pg8277)  &  Pg8215  &  (~ Ng3100) ) ;
 assign n5474 = ( Pg35  &  (~ n5472) ) | ( (~ Pg35)  &  (~ Ng3100) ) | ( (~ n5472)  &  (~ Ng3100) ) ;
 assign Ng25650 = ( (~ n5474) ) ;
 assign n5475 = ( (~ Pg35)  &  (~ Ng3050) ) | ( Pg35  &  (~ Ng3338) ) | ( (~ Ng3050)  &  (~ Ng3338) ) ;
 assign Ng25649 = ( (~ n5475) ) ;
 assign n5476 = ( (~ Pg35)  &  n6029 ) | ( n4381  &  n6029 ) | ( n5152  &  n6029 ) ;
 assign Ng25638 = ( (~ n5476) ) ;
 assign n5477 = ( Ng1554  &  (~ n5152) ) | ( n4382  &  Ng1559  &  (~ n5152) ) ;
 assign n5479 = ( (~ Pg35)  &  (~ Ng1559) ) | ( Pg35  &  (~ n5477) ) | ( (~ Ng1559)  &  (~ n5477) ) ;
 assign Ng25637 = ( (~ n5479) ) ;
 assign n5480 = ( (~ Pg35)  &  (~ Ng1521) ) | ( Pg35  &  n6033 ) | ( (~ Ng1521)  &  n6033 ) ;
 assign Ng25636 = ( (~ n5480) ) ;
 assign n5481 = ( (~ Pg35)  &  n6037 ) | ( n4384  &  n6037 ) | ( n5154  &  n6037 ) ;
 assign Ng25629 = ( (~ n5481) ) ;
 assign n5482 = ( Ng1211  &  (~ n5154) ) | ( n4385  &  Ng1216  &  (~ n5154) ) ;
 assign n5483 = ( (~ Pg35)  &  (~ Ng1216) ) | ( Pg35  &  (~ n5482) ) | ( (~ Ng1216)  &  (~ n5482) ) ;
 assign Ng25628 = ( (~ n5483) ) ;
 assign n5484 = ( (~ Pg35)  &  (~ Ng1178) ) | ( Pg35  &  n6041 ) | ( (~ Ng1178)  &  n6041 ) ;
 assign Ng25627 = ( (~ n5484) ) ;
 assign n5485 = ( (~ n3812)  &  (~ n4259) ) | ( (~ n3812)  &  Ng817 ) | ( (~ n4259)  &  (~ Ng817) ) ;
 assign n5486 = ( (~ n4180)  &  (~ Ng667) ) | ( n4180  &  (~ Ng686) ) | ( (~ Ng667)  &  (~ Ng686) ) ;
 assign Ng25615 = ( (~ n5486) ) ;
 assign n5487 = ( (~ n5137)  &  (~ Ng460) ) | ( n5137  &  (~ Ng452) ) | ( (~ Ng460)  &  (~ Ng452) ) ;
 assign Ng25604 = ( (~ n5487) ) ;
 assign n5488 = ( (~ Ng182)  &  (~ Ng174) ) | ( (~ Ng174)  &  n5137 ) | ( (~ Ng182)  &  (~ n5137) ) ;
 assign Ng25601 = ( (~ n5488) ) ;
 assign n5489 = ( (~ Ng174)  &  (~ Ng168) ) | ( (~ Ng168)  &  n5137 ) | ( (~ Ng174)  &  (~ n5137) ) ;
 assign Ng25600 = ( (~ n5489) ) ;
 assign n5490 = ( (~ Pg35)  &  (~ Ng358) ) | ( Pg35  &  n6047 ) | ( (~ Ng358)  &  n6047 ) ;
 assign Ng25597 = ( (~ n5490) ) ;
 assign n5491 = ( (~ Pg35)  &  (~ Ng370) ) | ( Pg35  &  n6048 ) | ( (~ Ng370)  &  n6048 ) ;
 assign Ng25596 = ( (~ n5491) ) ;
 assign n5492 = ( Pg35  &  n6052 ) | ( (~ Pg35)  &  (~ Ng191) ) | ( n6052  &  (~ Ng191) ) ;
 assign Ng25593 = ( (~ n5492) ) ;
 assign n5493 = ( (~ Pg35)  &  (~ Ng222) ) | ( Pg35  &  n6055 ) | ( (~ Ng222)  &  n6055 ) ;
 assign Ng25592 = ( (~ n5493) ) ;
 assign n5494 = ( (~ Pg35)  &  (~ Ng209) ) | ( Pg35  &  Ng218 ) | ( (~ Ng209)  &  Ng218 ) ;
 assign Ng25591 = ( (~ n5494) ) ;
 assign n5495 = ( (~ Pg35)  &  n6059 ) | ( (~ n619)  &  n6059 ) | ( Ng6736  &  n6059 ) ;
 assign Ng24354 = ( (~ n5495) ) ;
 assign n5496 = ( (~ Pg35)  &  (~ Ng6723) ) | ( Pg35  &  n6060 ) | ( (~ Ng6723)  &  n6060 ) ;
 assign Ng24353 = ( (~ n5496) ) ;
 assign n5497 = ( (~ Pg35)  &  n6062 ) | ( (~ n949)  &  n6062 ) | ( Ng6390  &  n6062 ) ;
 assign Ng24350 = ( (~ n5497) ) ;
 assign n5498 = ( (~ Pg35)  &  (~ Ng6377) ) | ( Pg35  &  n6063 ) | ( (~ Ng6377)  &  n6063 ) ;
 assign Ng24349 = ( (~ n5498) ) ;
 assign n5499 = ( (~ Pg35)  &  n6065 ) | ( (~ n654)  &  n6065 ) | ( Ng6044  &  n6065 ) ;
 assign Ng24346 = ( (~ n5499) ) ;
 assign n5500 = ( (~ Pg35)  &  (~ Ng6031) ) | ( Pg35  &  n6066 ) | ( (~ Ng6031)  &  n6066 ) ;
 assign Ng24345 = ( (~ n5500) ) ;
 assign n5501 = ( (~ Pg35)  &  n6068 ) | ( (~ n1069)  &  n6068 ) | ( Ng5698  &  n6068 ) ;
 assign Ng24342 = ( (~ n5501) ) ;
 assign n5502 = ( (~ Pg35)  &  (~ Ng5685) ) | ( Pg35  &  n6069 ) | ( (~ Ng5685)  &  n6069 ) ;
 assign Ng24341 = ( (~ n5502) ) ;
 assign n5503 = ( (~ Pg35)  &  n6071 ) | ( (~ n1006)  &  n6071 ) | ( Ng5352  &  n6071 ) ;
 assign Ng24338 = ( (~ n5503) ) ;
 assign n5504 = ( (~ Pg35)  &  (~ Ng5339) ) | ( Pg35  &  n6072 ) | ( (~ Ng5339)  &  n6072 ) ;
 assign Ng24337 = ( (~ n5504) ) ;
 assign n5505 = ( (~ Pg35)  &  (~ Ng4308) ) | ( Pg35  &  n6074 ) | ( (~ Ng4308)  &  n6074 ) ;
 assign Ng24282 = ( (~ n5505) ) ;
 assign n5506 = ( (~ Pg35)  &  (~ Ng4235) ) | ( Pg35  &  (~ n6079) ) | ( (~ Ng4235)  &  (~ n6079) ) ;
 assign Ng24279 = ( (~ n5506) ) ;
 assign n5507 = ( (~ Pg35)  &  n6082 ) | ( (~ n416)  &  n6082 ) | ( Ng4049  &  n6082 ) ;
 assign Ng24277 = ( (~ n5507) ) ;
 assign n5508 = ( (~ Pg35)  &  (~ Ng4031) ) | ( Pg35  &  n6083 ) | ( (~ Ng4031)  &  n6083 ) ;
 assign Ng24276 = ( (~ n5508) ) ;
 assign n5509 = ( (~ Pg35)  &  n6085 ) | ( (~ n218)  &  n6085 ) | ( Ng3698  &  n6085 ) ;
 assign Ng24273 = ( (~ n5509) ) ;
 assign n5510 = ( (~ Pg35)  &  (~ Ng3680) ) | ( Pg35  &  n6086 ) | ( (~ Ng3680)  &  n6086 ) ;
 assign Ng24272 = ( (~ n5510) ) ;
 assign n5511 = ( (~ Pg35)  &  n6088 ) | ( (~ n724)  &  n6088 ) | ( Ng3347  &  n6088 ) ;
 assign Ng24269 = ( (~ n5511) ) ;
 assign n5512 = ( (~ Pg35)  &  (~ Ng3329) ) | ( Pg35  &  n6089 ) | ( (~ Ng3329)  &  n6089 ) ;
 assign Ng24268 = ( (~ n5512) ) ;
 assign n5513 = ( (~ Pg35)  &  (~ Ng1554) ) | ( Pg35  &  (~ Ng496) ) | ( (~ Ng1554)  &  (~ Ng496) ) ;
 assign Ng24258 = ( (~ n5513) ) ;
 assign n5514 = ( (~ Pg35)  &  (~ Ng1339) ) | ( Pg35  &  n6092 ) | ( (~ Ng1339)  &  n6092 ) ;
 assign Ng24256 = ( (~ n5514) ) ;
 assign n5515 = ( (~ Pg35)  &  (~ Ng1306) ) | ( Pg35  &  n6094 ) | ( (~ Ng1306)  &  n6094 ) ;
 assign Ng24253 = ( (~ n5515) ) ;
 assign n5516 = ( (~ Pg35)  &  (~ Ng1526) ) | ( Pg35  &  n6095 ) | ( (~ Ng1526)  &  n6095 ) ;
 assign Ng24252 = ( (~ n5516) ) ;
 assign n5517 = ( (~ n3772)  &  (~ Ng1442) ) | ( n3772  &  (~ Ng1495) ) | ( (~ Ng1442)  &  (~ Ng1495) ) ;
 assign Ng24251 = ( (~ n5517) ) ;
 assign n5518 = ( n3772  &  (~ Ng1489) ) | ( (~ n3772)  &  (~ Ng1495) ) | ( (~ Ng1489)  &  (~ Ng1495) ) ;
 assign Ng24250 = ( (~ n5518) ) ;
 assign n5519 = ( Pg35  &  (~ wire4432) ) | ( (~ Pg35)  &  (~ Ng1211) ) | ( (~ wire4432)  &  (~ Ng1211) ) ;
 assign Ng24242 = ( (~ n5519) ) ;
 assign n5520 = ( (~ Pg35)  &  (~ Ng996) ) | ( Pg35  &  n6097 ) | ( (~ Ng996)  &  n6097 ) ;
 assign Ng24240 = ( (~ n5520) ) ;
 assign n5521 = ( (~ Pg35)  &  (~ Ng962) ) | ( Pg35  &  n6099 ) | ( (~ Ng962)  &  n6099 ) ;
 assign Ng24237 = ( (~ n5521) ) ;
 assign n5522 = ( (~ Pg35)  &  (~ Ng1183) ) | ( Pg35  &  n6100 ) | ( (~ Ng1183)  &  n6100 ) ;
 assign Ng24236 = ( (~ n5522) ) ;
 assign n5523 = ( (~ n3778)  &  (~ Ng1099) ) | ( n3778  &  (~ Ng1152) ) | ( (~ Ng1099)  &  (~ Ng1152) ) ;
 assign Ng24235 = ( (~ n5523) ) ;
 assign n5524 = ( n3778  &  (~ Ng1146) ) | ( (~ n3778)  &  (~ Ng1152) ) | ( (~ Ng1146)  &  (~ Ng1152) ) ;
 assign Ng24234 = ( (~ n5524) ) ;
 assign n5525 = ( (~ n3812)  &  (~ Ng847) ) | ( n3812  &  (~ Ng854) ) | ( (~ Ng847)  &  (~ Ng854) ) ;
 assign Ng24216 = ( (~ n5525) ) ;
 assign n5526 = ( n3812  &  (~ Ng475) ) | ( (~ n3812)  &  (~ Ng441) ) | ( (~ Ng475)  &  (~ Ng441) ) ;
 assign Ng24207 = ( (~ n5526) ) ;
 assign n5527 = ( (~ n3812)  &  (~ Ng437) ) | ( n3812  &  (~ Ng441) ) | ( (~ Ng437)  &  (~ Ng441) ) ;
 assign Ng24206 = ( (~ n5527) ) ;
 assign n5528 = ( n3812  &  (~ Ng433) ) | ( (~ n3812)  &  (~ Ng429) ) | ( (~ Ng433)  &  (~ Ng429) ) ;
 assign Ng24204 = ( (~ n5528) ) ;
 assign n5529 = ( (~ n3812)  &  (~ Ng401) ) | ( n3812  &  (~ Ng429) ) | ( (~ Ng401)  &  (~ Ng429) ) ;
 assign Ng24203 = ( (~ n5529) ) ;
 assign n5530 = ( n3812  &  (~ Ng411) ) | ( (~ n3812)  &  (~ Ng424) ) | ( (~ Ng411)  &  (~ Ng424) ) ;
 assign Ng24202 = ( (~ n5530) ) ;
 assign n5531 = ( n3812  &  (~ Ng392) ) | ( (~ n3812)  &  (~ Ng405) ) | ( (~ Ng392)  &  (~ Ng405) ) ;
 assign Ng24201 = ( (~ n5531) ) ;
 assign n5532 = ( (~ Pg35)  &  (~ Ng2946) ) | ( Pg35  &  n6105 ) | ( (~ Ng2946)  &  n6105 ) ;
 assign Ng21901 = ( (~ n5532) ) ;
 assign n5533 = ( (~ Pg35)  &  (~ Ng4239) ) | ( Pg35  &  n6109 ) | ( (~ Ng4239)  &  n6109 ) ;
 assign Ng21900 = ( (~ n5533) ) ;
 assign n5534 = ( Pg35  &  n5189 ) | ( (~ Pg35)  &  (~ Ng4291) ) | ( n5189  &  (~ Ng4291) ) ;
 assign Ng21899 = ( (~ n5534) ) ;
 assign n5535 = ( Pg35  &  n5187 ) | ( (~ Pg35)  &  (~ Ng4284) ) | ( n5187  &  (~ Ng4284) ) ;
 assign Ng21898 = ( (~ n5535) ) ;
 assign n5536 = ( Pg35  &  n5192 ) | ( (~ Pg35)  &  (~ Ng4281) ) | ( n5192  &  (~ Ng4281) ) ;
 assign Ng21897 = ( (~ n5536) ) ;
 assign n5537 = ( (~ Pg35)  &  (~ Ng4245) ) | ( Pg35  &  n5190 ) | ( (~ Ng4245)  &  n5190 ) ;
 assign Ng21896 = ( (~ n5537) ) ;
 assign n5538 = ( (~ Pg35)  &  (~ Ng4273) ) | ( Pg35  &  Ng4239 ) | ( (~ Ng4273)  &  Ng4239 ) ;
 assign Ng21892 = ( (~ n5538) ) ;
 assign n5539 = ( (~ Pg35)  &  (~ Ng4180) ) | ( Pg35  &  n6075 ) | ( (~ Ng4180)  &  n6075 ) ;
 assign Ng21891 = ( (~ n5539) ) ;
 assign n5540 = ( n1310 ) | ( (~ Ng2882) ) ;
 assign n5541 = ( (~ Ng534) ) | ( n4421 ) ;
 assign n5543 = ( n1280  &  n4412 ) | ( n4394  &  n4412 ) | ( n1280  &  (~ Ng16) ) | ( n4394  &  (~ Ng16) ) ;
 assign n5545 = ( n1277 ) | ( (~ Ng790) ) ;
 assign n5544 = ( (~ n1250)  &  n1289  &  n5545 ) | ( (~ n1250)  &  (~ Ng749)  &  n5545 ) ;
 assign n5546 = ( n1331  &  n4421 ) | ( (~ Ng608)  &  n4421 ) | ( n1331  &  Ng550 ) | ( (~ Ng608)  &  Ng550 ) ;
 assign n5547 = ( (~ Ng572)  &  n5546 ) | ( n4419  &  n5546 ) ;
 assign n5548 = ( n1309  &  n4412 ) | ( n4394  &  n4412 ) | ( n1309  &  (~ Ng50) ) | ( n4394  &  (~ Ng50) ) ;
 assign n5549 = ( n1310  &  (~ Ng2980) ) | ( (~ Ng2886)  &  (~ Ng2980) ) | ( n1310  &  n4449 ) | ( (~ Ng2886)  &  n4449 ) ;
 assign n5550 = ( n1331 ) | ( (~ Ng604) ) ;
 assign n5551 = ( n1293  &  n4412 ) | ( n4394  &  n4412 ) | ( n1293  &  (~ Ng51) ) | ( n4394  &  (~ Ng51) ) ;
 assign n5552 = ( n4426  &  n4442 ) | ( n4442  &  (~ Ng1283) ) | ( n4426  &  (~ Ng2138) ) | ( (~ Ng1283)  &  (~ Ng2138) ) ;
 assign n5554 = ( n1331 ) | ( (~ Ng599) ) ;
 assign n5553 = ( (~ n1250)  &  n4419  &  n5554 ) | ( (~ n1250)  &  (~ Ng562)  &  n5554 ) ;
 assign n5555 = ( n1277  &  n1289 ) | ( n1289  &  (~ Ng781) ) | ( n1277  &  (~ Ng739) ) | ( (~ Ng781)  &  (~ Ng739) ) ;
 assign n5556 = ( n4421  &  n5555 ) | ( (~ Ng199)  &  n5555 ) ;
 assign n5557 = ( n1301  &  n4412 ) | ( n4394  &  n4412 ) | ( n1301  &  (~ Ng52) ) | ( n4394  &  (~ Ng52) ) ;
 assign n5558 = ( n1310  &  n1323 ) | ( n1310  &  (~ Ng2902) ) | ( n1323  &  (~ Ng2848) ) | ( (~ Ng2902)  &  (~ Ng2848) ) ;
 assign n5559 = ( n1294  &  n1351 ) | ( n1294  &  (~ Ng2844) ) | ( n1351  &  (~ Ng2907) ) | ( (~ Ng2844)  &  (~ Ng2907) ) ;
 assign n5560 = ( (~ Ng1300)  &  (~ Ng956) ) | ( (~ Ng956)  &  n4464 ) | ( (~ Ng1300)  &  n4465 ) | ( n4464  &  n4465 ) ;
 assign n5561 = ( Pg35  &  n1289 ) | ( Pg35  &  (~ Ng772) ) | ( n1289  &  n4418 ) | ( (~ Ng772)  &  n4418 ) ;
 assign n5562 = ( n1331  &  (~ Ng590) ) | ( (~ Ng626)  &  (~ Ng590) ) | ( n1331  &  n4419 ) | ( (~ Ng626)  &  n4419 ) ;
 assign n5563 = ( (~ Ng1472)  &  (~ Ng1129) ) | ( (~ Ng1129)  &  n4464 ) | ( (~ Ng1472)  &  n4465 ) | ( n4464  &  n4465 ) ;
 assign n5564 = ( n1277 ) | ( (~ Ng554) ) ;
 assign n5565 = ( (~ Ng1105)  &  (~ Ng1448) ) | ( (~ Ng1105)  &  n4464 ) | ( (~ Ng1448)  &  n4465 ) | ( n4464  &  n4465 ) ;
 assign n5566 = ( n4412  &  n4442 ) | ( n4442  &  (~ Ng8) ) | ( n4412  &  (~ Ng5507) ) | ( (~ Ng8)  &  (~ Ng5507) ) ;
 assign n5567 = ( n1310 ) | ( (~ Ng2898) ) ;
 assign n5568 = ( n1331 ) | ( (~ Ng617) ) ;
 assign n5569 = ( (~ Ng1478)  &  (~ Ng1135) ) | ( (~ Ng1135)  &  n4464 ) | ( (~ Ng1478)  &  n4465 ) | ( n4464  &  n4465 ) ;
 assign n5570 = ( n4412  &  n4433 ) | ( n4433  &  (~ Ng48) ) | ( n4412  &  (~ Ng4912) ) | ( (~ Ng48)  &  (~ Ng4912) ) ;
 assign n5571 = ( n4515  &  n4518 ) | ( n4516  &  n4518 ) | ( n4515  &  n3572 ) | ( n4516  &  n3572 ) ;
 assign n5572 = ( n1014  &  n4521 ) | ( n3501  &  n4521 ) | ( n1014  &  n3208 ) | ( n3501  &  n3208 ) ;
 assign n5573 = ( n3184  &  n3291 ) | ( n3291  &  (~ n4110) ) | ( n3184  &  (~ n4582) ) | ( (~ n4110)  &  (~ n4582) ) ;
 assign n5576 = ( n1633  &  n3531 ) | ( n3401  &  n3531 ) | ( n1633  &  (~ n4585) ) | ( n3401  &  (~ n4585) ) ;
 assign n5578 = ( n3238  &  n3583 ) | ( n3238  &  (~ n4110) ) | ( n3583  &  (~ n4582) ) | ( (~ n4110)  &  (~ n4582) ) ;
 assign n5579 = ( n1633  &  n3476 ) | ( n3346  &  n3476 ) | ( n1633  &  (~ n4585) ) | ( n3346  &  (~ n4585) ) ;
 assign n5580 = ( (~ n1156)  &  n4696 ) | ( (~ n1156)  &  (~ Ng2643) ) ;
 assign n5581 = ( (~ n1184)  &  n4706 ) | ( (~ n1184)  &  (~ Ng2509) ) ;
 assign n5582 = ( (~ n1203)  &  n4716 ) | ( (~ n1203)  &  (~ Ng2375) ) ;
 assign n5583 = ( (~ n1199)  &  n4726 ) | ( (~ n1199)  &  (~ Ng2241) ) ;
 assign n5584 = ( (~ n1187)  &  n4737 ) | ( (~ n1187)  &  (~ Ng2084) ) ;
 assign n5585 = ( (~ n1192)  &  n4747 ) | ( (~ n1192)  &  (~ Ng1950) ) ;
 assign n5586 = ( (~ n1122)  &  n4757 ) | ( (~ n1122)  &  (~ Ng1816) ) ;
 assign n5587 = ( (~ n1201)  &  n4767 ) | ( (~ n1201)  &  (~ Ng1682) ) ;
 assign n5588 = ( (~ n1641)  &  n4796 ) ;
 assign n5589 = ( Pg35  &  (~ n2196) ) | ( Pg35  &  (~ Ng1373)  &  n4805 ) ;
 assign n5590 = ( Pg35  &  (~ n2209) ) | ( Pg35  &  (~ Ng1030)  &  n4818 ) ;
 assign n5591 = ( n2555  &  (~ n4343) ) | ( (~ n1107)  &  (~ n4343)  &  (~ n4345) ) ;
 assign n5593 = ( Ng2236  &  Ng2370 ) | ( n4868  &  Ng2370 ) | ( Ng2236  &  n4135 ) | ( n4868  &  n4135 ) ;
 assign n5595 = ( n4135  &  (~ Ng2803) ) | ( (~ Ng2807)  &  (~ Ng2803) ) | ( n4135  &  n4868 ) | ( (~ Ng2807)  &  n4868 ) ;
 assign n5597 = ( Ng1945  &  Ng2079 ) | ( n4862  &  Ng2079 ) | ( Ng1945  &  n4689 ) | ( n4862  &  n4689 ) ;
 assign n5599 = ( n4135  &  (~ Ng2771) ) | ( (~ Ng2775)  &  (~ Ng2771) ) | ( n4135  &  n4868 ) | ( (~ Ng2775)  &  n4868 ) ;
 assign n5601 = ( (~ Pg17688) ) | ( n3223 ) | ( (~ Ng6645) ) ;
 assign n5602 = ( (~ Pg17688) ) | ( n3227 ) | ( (~ Ng6653) ) ;
 assign n5603 = ( (~ Pg17760) ) | ( n3263 ) | ( (~ Ng6283) ) ;
 assign n5604 = ( (~ Pg14779) ) | ( n3281 ) | ( (~ Ng6275) ) ;
 assign n5605 = ( (~ Pg17607) ) | ( n3331 ) | ( (~ Ng5953) ) ;
 assign n5606 = ( (~ Pg17607) ) | ( n3335 ) | ( (~ Ng5961) ) ;
 assign n5607 = ( (~ Pg17580) ) | ( n3386 ) | ( (~ Ng5607) ) ;
 assign n5608 = ( (~ Pg17580) ) | ( n3391 ) | ( (~ Ng5615) ) ;
 assign n5609 = ( (~ Pg17519) ) | ( n3440 ) | ( (~ Ng5260) ) ;
 assign n5610 = ( (~ Pg17674) ) | ( n1986 ) | ( (~ Ng5252) ) ;
 assign n5611 = ( (~ Ng4836)  &  (~ Ng4864) ) | ( (~ Ng4864)  &  (~ Ng5011) ) | ( (~ Ng4836)  &  Ng3333 ) | ( (~ Ng5011)  &  Ng3333 ) ;
 assign n5612 = ( (~ Ng4871)  &  (~ Ng4878) ) | ( (~ Ng4878)  &  (~ Ng3684) ) | ( (~ Ng4871)  &  Ng4035 ) | ( (~ Ng3684)  &  Ng4035 ) ;
 assign n5613 = ( (~ wire4427)  &  (~ Ng4674) ) | ( (~ Ng4646)  &  (~ Ng4674) ) | ( (~ wire4427)  &  Ng4821 ) | ( (~ Ng4646)  &  Ng4821 ) ;
 assign n5614 = ( (~ Ng4681)  &  (~ Ng4688) ) | ( (~ Ng4688)  &  (~ Ng4831) ) | ( (~ Ng4681)  &  Ng4826 ) | ( (~ Ng4831)  &  Ng4826 ) ;
 assign n5615 = ( (~ Pg16659) ) | ( n3516 ) | ( (~ Ng3953) ) ;
 assign n5616 = ( (~ Pg16775) ) | ( n1998 ) | ( (~ Ng3945) ) ;
 assign n5617 = ( (~ Pg16627) ) | ( n5034 ) | ( (~ Ng3602) ) ;
 assign n5618 = ( (~ Pg13926) ) | ( n5034 ) | ( (~ Ng3578) ) ;
 assign n5619 = ( (~ Pg16718) ) | ( n4516 ) | ( (~ Ng3235) ) ;
 assign n5620 = ( (~ Pg13895) ) | ( n3624 ) | ( (~ Ng3227) ) ;
 assign n5622 = ( n2016  &  n4516 ) | ( n2016  &  Ng3347 ) | ( n4516  &  (~ Ng3347) ) ;
 assign n5623 = ( (~ Ng3343)  &  n3607 ) | ( Ng3343  &  n3624 ) | ( n3607  &  n3624 ) ;
 assign n5621 = ( Ng4939  &  (~ n4793) ) | ( (~ n4793)  &  n5622  &  n5623 ) ;
 assign n5626 = ( Ng5694  &  n3386 ) | ( (~ Ng5694)  &  n3391 ) | ( n3386  &  n3391 ) ;
 assign n5627 = ( n3371  &  n4783 ) | ( n4783  &  Ng5698 ) | ( n3371  &  (~ Ng5698) ) ;
 assign n5625 = ( Ng4749  &  (~ n4784) ) | ( (~ n4784)  &  n5626  &  n5627 ) ;
 assign n5630 = ( (~ n4004)  &  (~ Ng979) ) | ( (~ Ng979)  &  (~ Ng1061) ) | ( (~ Ng979)  &  (~ Ng1052) ) ;
 assign n5631 = ( (~ n3812)  &  Ng832 ) | ( Pg35  &  Ng832  &  (~ Ng817) ) ;
 assign n5634 = ( (~ Pg35)  &  (~ Ng1395) ) | ( Pg19357  &  (~ Ng1395) ) | ( (~ Pg35)  &  n4222 ) | ( Pg19357  &  n4222 ) ;
 assign n5635 = ( Pg17400 ) | ( Pg17291 ) | ( Pg17316 ) ;
 assign n5636 = ( (~ Pg35)  &  n4235 ) | ( Pg19334  &  n4235 ) | ( (~ Pg35)  &  (~ Ng1052) ) | ( Pg19334  &  (~ Ng1052) ) ;
 assign n5637 = ( Pg35  &  n1366 ) | ( Pg35  &  Ng2984 ) ;
 assign n5640 = ( Ng655 ) | ( Ng718 ) | ( Ng753 ) ;
 assign n5641 = ( n1222  &  (~ Ng4332) ) | ( Pg90  &  (~ Ng4332)  &  (~ Ng2994) ) ;
 assign n5642 = ( (~ Ng4322)  &  n5641 ) | ( Ng4332  &  (~ Ng4322)  &  Ng4311 ) ;
 assign n5643 = ( n1222  &  (~ Ng4332)  &  Ng4322 ) | ( (~ Ng4332)  &  Ng4322  &  (~ Ng4515) ) ;
 assign n5644 = ( Ng4601 ) | ( (~ Ng4584) ) | ( Ng4608 ) | ( (~ Ng4593) ) ;
 assign n5645 = ( Ng4340  &  (~ Ng4349) ) | ( (~ Ng4349)  &  n5642 ) | ( (~ Ng4349)  &  n5643 ) ;
 assign n5646 = ( n1013  &  (~ n5645) ) | ( Ng4340  &  (~ n5645) ) | ( (~ Ng4349)  &  (~ n5645) ) ;
 assign n5648 = ( n1013  &  (~ Ng4340) ) | ( n1013  &  (~ Ng4349) ) | ( Ng4340  &  (~ Ng4349) ) ;
 assign n5649 = ( (~ Ng4358)  &  n5646 ) | ( Ng4358  &  n5648 ) | ( n5646  &  n5648 ) ;
 assign n5652 = ( (~ Pg91) ) | ( n178 ) | ( n179 ) | ( Ng2965 ) ;
 assign n5651 = ( n5652  &  Pg35 ) ;
 assign n5655 = ( n172 ) | ( n173 ) | ( n175 ) | ( n176 ) | ( Ng2955 ) | ( n4568 ) | ( (~ n4570) ) | ( Ng2946 ) ;
 assign n5654 = ( n5655  &  Pg35 ) ;
 assign n5658 = ( Ng4072 ) | ( Ng4153 ) | ( Ng2941 ) ;
 assign n5657 = ( n5658  &  Pg35 ) ;
 assign n5660 = ( Pg35  &  (~ n6123) ) ;
 assign n5664 = ( (~ Pg44) ) | ( Ng2927 ) | ( Ng2932 ) ;
 assign n5663 = ( n5664  &  Pg35 ) ;
 assign n5666 = ( Pg35  &  (~ n6124) ) ;
 assign n5670 = ( Ng301 ) | ( Ng2902 ) | ( n1224 ) ;
 assign n5669 = ( n5670  &  Pg35 ) ;
 assign n5677 = ( n179 ) | ( n178 ) | ( Ng2882 ) ;
 assign n5676 = ( n5677  &  Pg35 ) ;
 assign n5682 = ( n175 ) | ( n176 ) | ( Ng2856 ) ;
 assign n5681 = ( n5682  &  Pg35 ) ;
 assign n5685 = ( n173 ) | ( n172 ) | ( Ng2848 ) ;
 assign n5684 = ( n5685  &  Pg35 ) ;
 assign n5687 = ( (~ Ng4087)  &  n5573  &  n5576 ) ;
 assign n5688 = ( n5579  &  n5578  &  Ng4087 ) ;
 assign n5698 = ( Ng2724  &  (~ Ng2807) ) | ( (~ Ng2724)  &  (~ Ng2803) ) | ( (~ Ng2807)  &  (~ Ng2803) ) ;
 assign n5699 = ( Ng2724  &  (~ Ng2819) ) | ( (~ Ng2724)  &  (~ Ng2815) ) | ( (~ Ng2819)  &  (~ Ng2815) ) ;
 assign n5700 = ( Ng2724  &  (~ Ng2775) ) | ( (~ Ng2724)  &  (~ Ng2771) ) | ( (~ Ng2775)  &  (~ Ng2771) ) ;
 assign n5701 = ( Ng2724  &  (~ Ng2787) ) | ( (~ Ng2724)  &  (~ Ng2783) ) | ( (~ Ng2787)  &  (~ Ng2783) ) ;
 assign n5704 = ( Pg35 ) | ( (~ Ng2894) ) ;
 assign n5705 = ( (~ Pg35) ) | ( (~ Ng1291) ) ;
 assign n5706 = ( (~ Pg35) ) | ( (~ Ng947) ) ;
 assign n5710 = ( (~ Pg35)  &  Ng4878 ) | ( Ng4878  &  (~ Ng4843)  &  n4630 ) ;
 assign n5712 = ( (~ Pg35)  &  Ng4688 ) | ( Ng4688  &  (~ Ng4653)  &  n4633 ) ;
 assign n5715 = ( n1552  &  (~ Ng4340) ) | ( (~ n1552)  &  n1555 ) | ( (~ Ng4340)  &  n1555 ) ;
 assign n5717 = ( Pg35 ) | ( (~ Ng2827) ) ;
 assign n5719 = ( Pg35 ) | ( (~ Ng2815) ) ;
 assign n5721 = ( Pg35 ) | ( (~ Ng2819) ) ;
 assign n5723 = ( Pg35 ) | ( (~ Ng2807) ) ;
 assign n5724 = ( Pg35 ) | ( (~ Ng2795) ) ;
 assign n5725 = ( Pg35 ) | ( (~ Ng2783) ) ;
 assign n5726 = ( Pg35 ) | ( (~ Ng2787) ) ;
 assign n5727 = ( Pg35 ) | ( (~ Ng2775) ) ;
 assign n5730 = ( (~ Ng174)  &  (~ Ng392) ) | ( (~ Ng174)  &  (~ Ng452) ) | ( Ng392  &  (~ Ng452) ) ;
 assign n5731 = ( Ng405  &  (~ Ng437) ) | ( (~ Ng405)  &  (~ Ng424) ) | ( (~ Ng437)  &  (~ Ng424) ) ;
 assign n5732 = ( (~ Ng401)  &  Ng405 ) | ( (~ Ng401)  &  (~ Ng437) ) | ( (~ Ng405)  &  (~ Ng437) ) ;
 assign n5733 = ( (~ Ng392)  &  n5731 ) | ( Ng392  &  n5732 ) | ( n5731  &  n5732 ) ;
 assign n5734 = ( n3823  &  n4652 ) ;
 assign n5735 = ( n1647  &  (~ Ng4955) ) | ( (~ Ng4955)  &  n5734 ) | ( n1647  &  (~ n5734) ) ;
 assign n5737 = ( n3828  &  n4652 ) ;
 assign n5738 = ( n1651  &  (~ Ng4944) ) | ( (~ Ng4944)  &  n5737 ) | ( n1651  &  (~ n5737) ) ;
 assign n5740 = ( n1407  &  n4652 ) ;
 assign n5741 = ( n1658  &  (~ Ng4888) ) | ( (~ Ng4888)  &  n5740 ) | ( n1658  &  (~ n5740) ) ;
 assign n5743 = ( n3840  &  n4654 ) ;
 assign n5744 = ( n1660  &  (~ Ng4765) ) | ( (~ Ng4765)  &  n5743 ) | ( n1660  &  (~ n5743) ) ;
 assign n5746 = ( n3845  &  n4654 ) ;
 assign n5747 = ( n1664  &  (~ Ng4754) ) | ( (~ Ng4754)  &  n5746 ) | ( n1664  &  (~ n5746) ) ;
 assign n5749 = ( n3853  &  n4654 ) ;
 assign n5750 = ( n1671  &  (~ Ng4698) ) | ( (~ Ng4698)  &  n5749 ) | ( n1671  &  (~ n5749) ) ;
 assign n5752 = ( Pg35 ) | ( (~ Ng4340) ) ;
 assign n5754 = ( (~ Ng157) ) | ( n4672 ) ;
 assign n5755 = ( Ng4512 ) | ( Ng4581 ) ;
 assign n5756 = ( (~ n1222)  &  n4272 ) | ( n1222  &  (~ n5252) ) | ( n4272  &  (~ n5252) ) ;
 assign n5757 = ( Ng4552 ) | ( Ng4581 ) ;
 assign n5758 = ( (~ n1222)  &  n4274 ) | ( n1222  &  (~ n5255) ) | ( n4274  &  (~ n5255) ) ;
 assign n5760 = ( Pg35 ) | ( (~ Ng2759) ) ;
 assign n5777 = ( (~ n1097) ) | ( n4515 ) | ( n4781 ) ;
 assign n5775 = ( Pg35  &  (~ n3391)  &  n5777 ) | ( Pg35  &  (~ n5290)  &  n5777 ) ;
 assign n5781 = ( Pg35 ) | ( (~ Ng4108) ) ;
 assign n5785 = ( Pg35 ) | ( (~ Ng2756) ) ;
 assign n5793 = ( Pg35 ) | ( (~ Ng301) ) ;
 assign n5794 = ( n4842 ) | ( (~ Ng5041) ) | ( (~ Ng5046) ) ;
 assign n5795 = ( (~ Ng5052)  &  n4846 ) | ( Ng5052  &  n5794 ) | ( n4846  &  n5794 ) ;
 assign n5799 = ( Pg35 ) | ( (~ Ng4098) ) ;
 assign n5809 = ( (~ n4840)  &  (~ Ng5033) ) | ( Pg35  &  (~ Ng5033)  &  (~ n4844) ) ;
 assign n5812 = ( (~ Ng5052)  &  (~ n5794) ) | ( Pg35  &  (~ Ng5052)  &  (~ n4846) ) ;
 assign n5815 = ( Pg35 ) | ( (~ Ng5041) ) ;
 assign n5816 = ( Pg35 ) | ( (~ Ng5037) ) ;
 assign n5817 = ( Pg35 ) | ( (~ Ng5033) ) ;
 assign n5818 = ( Pg35 ) | ( (~ Ng5022) ) ;
 assign n5819 = ( (~ Pg35)  &  Ng283 ) | ( Ng283  &  (~ Ng287)  &  n4657 ) ;
 assign n5821 = ( (~ Ng4473) ) | ( Ng4459 ) ;
 assign n5825 = ( (~ Pg124)  &  (~ Pg120) ) | ( (~ Pg124)  &  Ng4146 ) | ( (~ Pg120)  &  (~ Ng4146) ) ;
 assign n5828 = ( (~ Pg116)  &  (~ Pg114) ) | ( (~ Pg116)  &  Ng4157 ) | ( (~ Pg114)  &  (~ Ng4157) ) ;
 assign n5829 = ( (~ Ng2638)  &  (~ Ng2504) ) | ( (~ Ng2638)  &  Ng2715 ) | ( (~ Ng2504)  &  (~ Ng2715) ) ;
 assign n5830 = ( Ng2819  &  Ng2815 ) | ( Ng2819  &  Ng2715 ) | ( Ng2815  &  (~ Ng2715) ) ;
 assign n5831 = ( n1090 ) | ( Ng2735 ) | ( (~ n4551) ) ;
 assign n5832 = ( (~ n5593)  &  n5831 ) | ( Ng2719  &  n5829  &  n5831 ) ;
 assign n5833 = ( (~ n5595)  &  (~ n5831) ) | ( Ng2719  &  n5830  &  (~ n5831) ) ;
 assign n5835 = ( (~ Ng1811)  &  (~ Ng1677) ) | ( (~ Ng1811)  &  Ng2715 ) | ( (~ Ng1677)  &  (~ Ng2715) ) ;
 assign n5836 = ( Ng2787  &  Ng2783 ) | ( Ng2787  &  Ng2715 ) | ( Ng2783  &  (~ Ng2715) ) ;
 assign n5837 = ( (~ n5597)  &  n5831 ) | ( (~ Ng2719)  &  n5831  &  n5835 ) ;
 assign n5838 = ( (~ n5599)  &  (~ n5831) ) | ( Ng2719  &  (~ n5831)  &  n5836 ) ;
 assign n5840 = ( (~ Pg35)  &  Ng2681 ) | ( Ng2675  &  n4945  &  Ng2681 ) ;
 assign n5842 = ( Pg35  &  (~ n1153)  &  Ng2657 ) | ( Pg35  &  Ng2657  &  n4947 ) ;
 assign n5843 = ( Pg35  &  (~ n1153)  &  Ng2595 ) | ( Pg35  &  n4550  &  Ng2595 ) ;
 assign n5845 = ( (~ Pg35)  &  Ng2547 ) | ( Ng2541  &  n4949  &  Ng2547 ) ;
 assign n5847 = ( Pg35  &  (~ n1151)  &  Ng2523 ) | ( Pg35  &  Ng2523  &  n4951 ) ;
 assign n5848 = ( Pg35  &  (~ n1151)  &  Ng2461 ) | ( Pg35  &  n4546  &  Ng2461 ) ;
 assign n5850 = ( (~ Pg35)  &  Ng2413 ) | ( Ng2407  &  n4952  &  Ng2413 ) ;
 assign n5852 = ( Pg35  &  (~ n1162)  &  Ng2389 ) | ( Pg35  &  Ng2389  &  n4954 ) ;
 assign n5853 = ( Pg35  &  (~ n1162)  &  Ng2327 ) | ( Pg35  &  n4548  &  Ng2327 ) ;
 assign n5855 = ( (~ Pg35)  &  Ng2279 ) | ( Ng2273  &  n4955  &  Ng2279 ) ;
 assign n5857 = ( Pg35  &  (~ n1104)  &  Ng2255 ) | ( Pg35  &  Ng2255  &  n4957 ) ;
 assign n5858 = ( Pg35  &  (~ n1104)  &  Ng2193 ) | ( Pg35  &  n4535  &  Ng2193 ) ;
 assign n5860 = ( (~ Pg35)  &  Ng2122 ) | ( Ng2116  &  n4959  &  Ng2122 ) ;
 assign n5862 = ( Pg35  &  (~ n1146)  &  Ng2098 ) | ( Pg35  &  Ng2098  &  n4961 ) ;
 assign n5863 = ( Pg35  &  (~ n1146)  &  Ng2036 ) | ( Pg35  &  n4542  &  Ng2036 ) ;
 assign n5865 = ( (~ Pg35)  &  Ng1988 ) | ( Ng1982  &  n4962  &  Ng1988 ) ;
 assign n5867 = ( Pg35  &  (~ n1126)  &  Ng1964 ) | ( Pg35  &  Ng1964  &  n4964 ) ;
 assign n5868 = ( Pg35  &  (~ n1126)  &  Ng1902 ) | ( Pg35  &  n4544  &  Ng1902 ) ;
 assign n5870 = ( (~ Pg35)  &  Ng1854 ) | ( Ng1848  &  n4965  &  Ng1854 ) ;
 assign n5872 = ( Pg35  &  (~ n1182)  &  Ng1830 ) | ( Pg35  &  Ng1830  &  n4967 ) ;
 assign n5873 = ( Pg35  &  (~ n1182)  &  Ng1768 ) | ( Pg35  &  n4538  &  Ng1768 ) ;
 assign n5875 = ( (~ Pg35)  &  Ng1720 ) | ( Ng1714  &  n4968  &  Ng1720 ) ;
 assign n5877 = ( Pg35  &  (~ n1087)  &  Ng1696 ) | ( Pg35  &  Ng1696  &  n4970 ) ;
 assign n5878 = ( Pg35  &  (~ n1087)  &  Ng1632 ) | ( Pg35  &  n4553  &  Ng1632 ) ;
 assign n5879 = ( Pg35 ) | ( (~ Ng1536) ) ;
 assign n5880 = ( Pg35 ) | ( (~ Ng1193) ) ;
 assign n5883 = ( (~ Pg35)  &  Ng6519 ) | ( (~ n4983)  &  Ng6513  &  Ng6519 ) ;
 assign n5885 = ( (~ Pg35)  &  Ng6500 ) | ( Ng6500  &  (~ n4983)  &  (~ Ng6505) ) ;
 assign n5886 = ( Pg12470  &  Ng6727 ) | ( (~ Pg12470)  &  (~ Ng6727) ) ;
 assign n5888 = ( Pg35  &  (~ n1109)  &  Ng6500 ) | ( Pg35  &  Ng6500  &  n5160 ) ;
 assign n5891 = ( (~ Pg35)  &  Ng6173 ) | ( (~ n4990)  &  Ng6167  &  Ng6173 ) ;
 assign n5893 = ( (~ Pg35)  &  Ng6154 ) | ( Ng6154  &  (~ n4990)  &  (~ Ng6159) ) ;
 assign n5894 = ( Pg12422  &  Ng6381 ) | ( (~ Pg12422)  &  (~ Ng6381) ) ;
 assign n5896 = ( Pg35  &  (~ n1196)  &  Ng6154 ) | ( Pg35  &  Ng6154  &  (~ n5162) ) ;
 assign n5900 = ( (~ Pg35)  &  Ng5827 ) | ( (~ n4998)  &  Ng5821  &  Ng5827 ) ;
 assign n5902 = ( (~ Pg35)  &  Ng5808 ) | ( Ng5808  &  (~ n4998)  &  (~ Ng5813) ) ;
 assign n5903 = ( Pg12350  &  Ng6035 ) | ( (~ Pg12350)  &  (~ Ng6035) ) ;
 assign n5905 = ( Pg35  &  (~ n1179)  &  Ng5808 ) | ( Pg35  &  Ng5808  &  n5163 ) ;
 assign n5908 = ( (~ Pg35)  &  Ng5481 ) | ( (~ n5005)  &  Ng5475  &  Ng5481 ) ;
 assign n5910 = ( (~ Pg35)  &  Ng5462 ) | ( (~ n5005)  &  (~ Ng5467)  &  Ng5462 ) ;
 assign n5911 = ( Pg12300  &  Ng5689 ) | ( (~ Pg12300)  &  (~ Ng5689) ) ;
 assign n5913 = ( Pg35  &  (~ n1097)  &  Ng5462 ) | ( Pg35  &  n5165  &  Ng5462 ) ;
 assign n5916 = ( (~ Pg35)  &  Ng5134 ) | ( (~ n5012)  &  Ng5128  &  Ng5134 ) ;
 assign n5918 = ( (~ Pg35)  &  Ng5115 ) | ( Ng5115  &  (~ n5012)  &  (~ Ng5120) ) ;
 assign n5919 = ( wire4415  &  Pg12238 ) | ( (~ wire4415)  &  (~ Pg12238) ) ;
 assign n5921 = ( Pg35  &  (~ wire4394)  &  Ng5115 ) | ( Pg35  &  Ng5115  &  n5167 ) ;
 assign n5922 = ( n3455  &  (~ Ng4983) ) | ( (~ Ng4983)  &  Ng4991 ) ;
 assign n5923 = ( n5612  &  n5611  &  n335 ) ;
 assign n5924 = ( n3464  &  (~ Ng4793) ) | ( (~ Ng4793)  &  Ng4801 ) ;
 assign n5925 = ( n5614  &  n5613  &  n419 ) ;
 assign n5928 = ( (~ Pg35)  &  Ng3827 ) | ( (~ n5023)  &  Ng3821  &  Ng3827 ) ;
 assign n5930 = ( (~ Pg35)  &  Ng3808 ) | ( Ng3808  &  (~ n5023)  &  (~ Ng3813) ) ;
 assign n5931 = ( Pg11418  &  Ng4040 ) | ( (~ Pg11418)  &  (~ Ng4040) ) ;
 assign n5933 = ( Pg35  &  (~ n1165)  &  Ng3808 ) | ( Pg35  &  Ng3808  &  n5168 ) ;
 assign n5936 = ( (~ Pg35)  &  Ng3476 ) | ( (~ n5030)  &  Ng3470  &  Ng3476 ) ;
 assign n5938 = ( (~ Pg35)  &  Ng3457 ) | ( Ng3457  &  (~ n5030)  &  (~ Ng3462) ) ;
 assign n5939 = ( Pg11388  &  Ng3689 ) | ( (~ Pg11388)  &  (~ Ng3689) ) ;
 assign n5941 = ( Pg35  &  (~ n1116)  &  Ng3457 ) | ( Pg35  &  Ng3457  &  n5170 ) ;
 assign n5944 = ( (~ Pg35)  &  Ng3125 ) | ( (~ n5038)  &  Ng3119  &  Ng3125 ) ;
 assign n5946 = ( (~ Pg35)  &  Ng3106 ) | ( (~ n5038)  &  (~ Ng3111)  &  Ng3106 ) ;
 assign n5947 = ( Pg11349  &  Ng3338 ) | ( (~ Pg11349)  &  (~ Ng3338) ) ;
 assign n5949 = ( Pg35  &  (~ n1135)  &  Ng3106 ) | ( Pg35  &  n5172  &  Ng3106 ) ;
 assign n5951 = ( Pg35 ) | ( (~ Ng2729) ) ;
 assign n5952 = ( n5174  &  n5043  &  Ng1454 ) | ( n5174  &  n5043  &  n5357 ) ;
 assign n5953 = ( Pg35  &  n5952 ) | ( Pg35  &  (~ n5043)  &  Ng1454 ) ;
 assign n5957 = ( n5177  &  n5044  &  Ng1467 ) | ( n5177  &  n5044  &  n5357 ) ;
 assign n5958 = ( Pg35  &  n5957 ) | ( Pg35  &  (~ n5044)  &  Ng1467 ) ;
 assign n5961 = ( n5178  &  n5045  &  Ng1437 ) | ( n5178  &  n5045  &  n5357 ) ;
 assign n5962 = ( Pg35  &  n5961 ) | ( Pg35  &  (~ n5045)  &  Ng1437 ) ;
 assign n5965 = ( n5179  &  n5046  &  Ng1111 ) | ( n5179  &  n5046  &  n5362 ) ;
 assign n5966 = ( Pg35  &  n5965 ) | ( Pg35  &  (~ n5046)  &  Ng1111 ) ;
 assign n5970 = ( n5182  &  n5047  &  Ng1124 ) | ( n5182  &  n5047  &  n5362 ) ;
 assign n5971 = ( Pg35  &  n5970 ) | ( Pg35  &  (~ n5047)  &  Ng1124 ) ;
 assign n5974 = ( n5183  &  n5048  &  Ng1094 ) | ( n5183  &  n5048  &  n5362 ) ;
 assign n5975 = ( Pg35  &  n5974 ) | ( Pg35  &  (~ n5048)  &  Ng1094 ) ;
 assign n5978 = ( Ng827  &  (~ n5049) ) ;
 assign n5980 = ( (~ Ng676) ) | ( (~ n5054) ) ;
 assign n5982 = ( Pg35 ) | ( (~ Ng482) ) ;
 assign n5984 = ( Ng417  &  n5733 ) | ( (~ Ng417)  &  (~ n5733) ) ;
 assign n5983 = ( (~ Pg35)  &  Ng417 ) | ( (~ n4170)  &  Ng417  &  n5984 ) ;
 assign n5985 = ( Pg35 ) | ( (~ Ng5057) ) ;
 assign n5986 = ( Pg35 ) | ( (~ Ng5069) ) ;
 assign n5988 = ( (~ Pg35) ) | ( n1013 ) | ( Ng4521 ) ;
 assign n5987 = ( n4368  &  Ng4527 ) | ( (~ n4368)  &  (~ Ng4527) ) ;
 assign n5989 = ( (~ Pg35) ) | ( Ng4125 ) | ( (~ Ng26936) ) ;
 assign n5992 = ( Pg35 ) | ( (~ Ng4082) ) ;
 assign n5993 = ( Pg35 ) | ( (~ Ng1351) ) ;
 assign n5994 = ( Pg35 ) | ( (~ Ng1008) ) ;
 assign n5995 = ( Ng10384 ) | ( Ng4473 ) ;
 assign n5999 = ( (~ Pg35)  &  n4368 ) | ( n4368  &  Ng4527 ) ;
 assign n6001 = ( (~ Pg35) ) | ( Ng2712 ) | ( (~ Ng26936) ) ;
 assign n6002 = ( Pg35 ) | ( (~ Ng1395) ) ;
 assign n6003 = ( Ng890  &  Ng896 ) | ( Ng890  &  (~ Ng862) ) | ( (~ Ng896)  &  (~ Ng862) ) ;
 assign n6004 = ( (~ n3812) ) | ( n4039 ) | ( (~ Ng812) ) ;
 assign n6005 = ( (~ Pg35) ) | ( n1215 ) ;
 assign n6007 = ( (~ Ng528)  &  n1173 ) | ( (~ Ng528)  &  n5057 ) ;
 assign n6010 = ( (~ Pg35) ) | ( (~ Pg7540) ) | ( Ng347 ) ;
 assign n6011 = ( (~ Pg35) ) | ( (~ Ng329) ) | ( (~ n5109) ) | ( Ng341 ) ;
 assign n6013 = ( (~ Pg35) ) | ( Ng311 ) | ( Ng305 ) | ( Ng26885 ) ;
 assign n6022 = ( Ng5069  &  n4103  &  (~ Ng5080) ) | ( (~ Ng5077)  &  n4103  &  (~ Ng5080) ) ;
 assign n6023 = ( (~ Pg35)  &  Ng4064 ) | ( (~ Ng4057)  &  Ng4064  &  Ng2841 ) ;
 assign n6029 = ( Pg35 ) | ( (~ Ng1564) ) ;
 assign n6032 = ( (~ Ng1526) ) | ( n3151 ) ;
 assign n6033 = ( (~ Ng1339)  &  (~ Ng1306) ) | ( (~ Ng1306)  &  n6032 ) | ( (~ Ng1339)  &  (~ n6032) ) ;
 assign n6036 = ( (~ n4322)  &  Ng1389 ) ;
 assign n6035 = ( Ng1351  &  n6036 ) | ( Ng1351  &  n4144 ) ;
 assign n6037 = ( Pg35 ) | ( (~ Ng1221) ) ;
 assign n6040 = ( (~ Ng1183) ) | ( n3167 ) ;
 assign n6041 = ( (~ Ng996)  &  (~ Ng962) ) | ( (~ Ng962)  &  n6040 ) | ( (~ Ng996)  &  (~ n6040) ) ;
 assign n6044 = ( (~ n4323)  &  Ng1046 ) ;
 assign n6043 = ( Ng1008  &  n6044 ) | ( Ng1008  &  n4160 ) ;
 assign n6047 = ( n1621  &  Ng370 ) | ( (~ n1621)  &  (~ Ng370) ) ;
 assign n6048 = ( Ng376  &  Ng358 ) | ( (~ Ng376)  &  (~ Ng358) ) ;
 assign n6050 = ( Pg8358  &  Ng191 ) | ( (~ Pg8358)  &  (~ Ng191) ) ;
 assign n6052 = ( (~ Ng209)  &  (~ n5139) ) | ( (~ Ng209)  &  n6050 ) | ( n5139  &  n6050 ) ;
 assign n6057 = ( n5139  &  n6050 ) ;
 assign n6055 = ( Pg8358  &  n6057 ) | ( (~ Pg8358)  &  (~ n6057) ) ;
 assign n6059 = ( Pg35 ) | ( (~ Ng6727) ) ;
 assign n6060 = ( Ng6727  &  n5140 ) | ( (~ Ng6727)  &  (~ n5140) ) ;
 assign n6062 = ( Pg35 ) | ( (~ Ng6381) ) ;
 assign n6063 = ( (~ n5142)  &  Ng6381 ) | ( n5142  &  (~ Ng6381) ) ;
 assign n6065 = ( Pg35 ) | ( (~ Ng6035) ) ;
 assign n6066 = ( Ng6035  &  n5143 ) | ( (~ Ng6035)  &  (~ n5143) ) ;
 assign n6068 = ( Pg35 ) | ( (~ Ng5689) ) ;
 assign n6069 = ( Ng5689  &  n5145 ) | ( (~ Ng5689)  &  (~ n5145) ) ;
 assign n6071 = ( Pg35 ) | ( (~ wire4415) ) ;
 assign n6072 = ( (~ n5147)  &  wire4415 ) | ( n5147  &  (~ wire4415) ) ;
 assign n6074 = ( Pg9251  &  Ng4308 ) | ( (~ Pg9251)  &  (~ Ng4308) ) ;
 assign n6075 = ( (~ Ng4253)  &  Ng4145 ) | ( Ng4253  &  Ng4164 ) | ( Ng4145  &  Ng4164 ) ;
 assign n6078 = ( (~ Pg8870) ) | ( Ng4235 ) ;
 assign n6077 = ( Pg8918 ) | ( Pg8917 ) | ( Pg8920 ) | ( Pg8919 ) | ( Pg8916 ) | ( Pg8915 ) | ( Pg11770 ) ;
 assign n6076 = ( Pg8870  &  n6078 ) | ( (~ Ng4235)  &  n6078  &  n6077 ) ;
 assign n6079 = ( (~ n6076)  &  n6075 ) | ( n6076  &  (~ n6075) ) ;
 assign n6082 = ( Pg35 ) | ( (~ Ng4040) ) ;
 assign n6083 = ( (~ n5149)  &  Ng4040 ) | ( n5149  &  (~ Ng4040) ) ;
 assign n6085 = ( Pg35 ) | ( (~ Ng3689) ) ;
 assign n6086 = ( (~ n5150)  &  Ng3689 ) | ( n5150  &  (~ Ng3689) ) ;
 assign n6088 = ( Pg35 ) | ( (~ Ng3338) ) ;
 assign n6089 = ( (~ n5151)  &  Ng3338 ) | ( n5151  &  (~ Ng3338) ) ;
 assign n6093 = ( Pg7946 ) | ( Pg19357 ) | ( Pg13272 ) | ( Ng1333 ) | ( Pg8475 ) ;
 assign n6092 = ( (~ n4226)  &  n6093 ) | ( n4226  &  (~ n6093) ) ;
 assign n6094 = ( Pg7946  &  (~ Ng1521) ) | ( (~ Pg7946)  &  (~ Ng1532) ) | ( (~ Ng1521)  &  (~ Ng1532) ) ;
 assign n6095 = ( Pg7946  &  (~ Ng1339) ) | ( (~ Pg7946)  &  (~ Ng1521) ) | ( (~ Ng1339)  &  (~ Ng1521) ) ;
 assign n6098 = ( Pg7916 ) | ( Pg19334 ) | ( Pg13259 ) | ( Ng990 ) | ( Pg8416 ) ;
 assign n6097 = ( (~ n4239)  &  n6098 ) | ( n4239  &  (~ n6098) ) ;
 assign n6099 = ( Pg7916  &  (~ Ng1178) ) | ( (~ Pg7916)  &  (~ Ng1189) ) | ( (~ Ng1178)  &  (~ Ng1189) ) ;
 assign n6100 = ( Pg7916  &  (~ Ng996) ) | ( (~ Pg7916)  &  (~ Ng1178) ) | ( (~ Ng996)  &  (~ Ng1178) ) ;
 assign n6102 = ( n4259 ) | ( (~ Ng822) ) | ( (~ Ng817) ) | ( (~ Ng723) ) ;
 assign n6107 = ( (~ Pg8786) ) | ( Ng4180 ) ;
 assign n6106 = ( Pg8785 ) | ( Pg8787 ) | ( Pg8783 ) | ( Pg8784 ) | ( Pg8788 ) | ( Pg8789 ) | ( Pg11447 ) ;
 assign n6105 = ( Pg8786  &  n6107 ) | ( (~ Ng4180)  &  n6107  &  n6106 ) ;
 assign n6109 = ( Ng4297 ) | ( Pg10122 ) ;
 assign Ng25676 = ( (~ n2319) ) ;
 assign Ng25694 = ( Pg35  &  Pg113 ) ;
 assign Ng25648 = ( (~ n2345) ) ;
 assign Ng34025 = ( (~ n1551) ) ;
 assign Ng25714 = ( (~ n2270) ) ;
 assign Ng25700 = ( (~ n2283) ) ;
 assign Ng24212 = ( Pg35  &  Pg64 ) ;
 assign Ng25662 = ( (~ n2332) ) ;
 assign Ng24247 = ( (~ n4152) ) ;
 assign Ng24231 = ( (~ n4168) ) ;
 assign Ng26953 = ( (~ n3940) ) ;
 assign Ng21893 = ( (~ n4210) ) ;
 assign Ng25742 = ( (~ n2244) ) ;
 assign Ng28079 = ( Pg35  &  Pg125 ) ;
 assign n6112 = ( Ng4125 ) | ( n1632 ) | ( Ng4057 ) | ( Ng4064 ) ;
 assign n6113 = ( n5687 ) | ( n5688 ) | ( n1191 ) ;
 assign n6114 = ( n1014 ) | ( (~ n1165) ) | ( n4779 ) ;
 assign n6115 = ( (~ n1109) ) | ( n4521 ) | ( n4779 ) ;
 assign n6116 = ( n1014 ) | ( (~ n1196) ) | ( n4781 ) ;
 assign n6117 = ( (~ wire4394) ) | ( n4521 ) | ( n4781 ) ;
 assign n6118 = ( (~ n1179) ) | ( n4518 ) | ( n4781 ) ;
 assign n6119 = ( (~ n1116) ) | ( n4518 ) | ( n4779 ) ;
 assign n6120 = ( (~ n1135) ) | ( n4515 ) | ( n4779 ) ;
 assign n6123 = ( n184  &  n185  &  (~ Ng2975) ) ;
 assign n6124 = ( n182  &  (~ Ng2917)  &  (~ n5079) ) ;
 assign n6128 = ( n1140  &  (~ n1646)  &  n4305  &  n4794 ) ;
 assign n6129 = ( n1093  &  (~ n1642)  &  n4308  &  n4794 ) ;
 assign n6130 = ( n1138  &  (~ n1643)  &  n4310  &  n4794 ) ;
 assign n6131 = ( n1096  &  (~ n1644)  &  n4312  &  n4794 ) ;
 assign n6132 = ( n1155  &  (~ n1640)  &  n4314  &  n4794 ) ;
 assign n6133 = ( n1113  &  (~ n1645)  &  n4316  &  n4794 ) ;
 assign n6134 = ( n1120  &  (~ n1639)  &  n4318  &  n4794 ) ;
 assign n6135 = ( wire4406  &  (~ n1641)  &  n4320  &  n4794 ) ;
 assign n6174 = ( n1238  &  n4176  &  n1239  &  n4177 ) ;
 assign n6186 = ( n3986  &  (~ n5088)  &  (~ Ng1389) ) ;
 assign n6188 = ( n4010  &  (~ n5093)  &  (~ Ng1046) ) ;
 assign n6200 = ( (~ n1533)  &  Ng4849  &  n4632 ) ;
 assign n6201 = ( (~ n1543)  &  Ng4659  &  n4635 ) ;
 assign n6203 = ( Ng608  &  n1629  &  (~ n4508) ) ;
 assign n6207 = ( Ng604  &  n1685  &  (~ n4508) ) ;
 assign n6214 = ( n1775  &  Ng2449  &  Pg35 ) ;
 assign n6218 = ( n1800  &  Ng2315  &  Pg35 ) ;
 assign n6234 = ( n1902  &  Ng1756  &  Pg35 ) ;
 assign n6244 = ( Ng599  &  n1945  &  (~ n4508) ) ;
 assign n6251 = ( Ng595  &  n2221  &  (~ n4508) ) ;
 assign n6256 = ( Ng590  &  n2480  &  (~ n4508) ) ;
 assign n6261 = ( n2232  &  Ng6597  &  Pg35 ) ;
 assign n6263 = ( n2579  &  Ng6653  &  Pg35 ) ;
 assign n6268 = ( n2594  &  Ng6633  &  Pg35 ) ;
 assign n6287 = ( n2652  &  Ng6287  &  Pg35 ) ;
 assign n6288 = ( n2655  &  Ng6283  &  Pg35 ) ;
 assign n6290 = ( n2661  &  Ng6275  &  Pg35 ) ;
 assign n6299 = ( n2258  &  Ng5905  &  Pg35 ) ;
 assign n6301 = ( n2695  &  Ng5961  &  Pg35 ) ;
 assign n6306 = ( n2710  &  Ng5941  &  Pg35 ) ;
 assign n6318 = ( n2271  &  Ng5559  &  Pg35 ) ;
 assign n6325 = ( n2768  &  Ng5595  &  Pg35 ) ;
 assign n6341 = ( n2817  &  Ng5260  &  Pg35 ) ;
 assign n6343 = ( n2823  &  Ng5252  &  Pg35 ) ;
 assign n6344 = ( n2826  &  Ng5248  &  Pg35 ) ;
 assign n6364 = ( n2885  &  Ng3953  &  Pg35 ) ;
 assign n6366 = ( n2891  &  Ng3945  &  Pg35 ) ;
 assign n6367 = ( n2894  &  Ng3941  &  Pg35 ) ;
 assign n6383 = ( n2943  &  Ng3602  &  Pg35 ) ;
 assign n6386 = ( n2952  &  Ng3590  &  Pg35 ) ;
 assign n6389 = ( n2961  &  Ng3578  &  Pg35 ) ;
 assign n6405 = ( n3010  &  Ng3239  &  Pg35 ) ;
 assign n6406 = ( n3013  &  Ng3235  &  Pg35 ) ;
 assign n6408 = ( n3019  &  Ng3227  &  Pg35 ) ;
 assign n6431 = ( (~ Pg35)  &  Ng1454 ) ;
 assign n6435 = ( (~ Pg35)  &  Ng1111 ) ;
 assign n6444 = ( n4096  &  wire4434  &  Pg35 ) ;
 assign Ng32996 = ( (~ n2435) ) ;
 assign Ng32992 = ( (~ n2448) ) ;
 assign Ng32988 = ( (~ n2461) ) ;
 assign Ng24263 = ( (~ n4217) ) ;
 assign Ng33040 = ( (~ n2308) ) ;
 assign Ng33016 = ( (~ n2368) ) ;
 assign Ng33012 = ( (~ n2381) ) ;
 assign Ng33008 = ( (~ n2395) ) ;
 assign Ng33004 = ( (~ n2408) ) ;
 assign Ng33000 = ( (~ n2421) ) ;
 assign Ng25685 = ( (~ n4114) ) ;
 assign Ng25639 = ( (~ n4134) ) ;
 assign Ng33044 = ( (~ n2301) ) ;
 assign Ng30458 = ( (~ n2859) ) ;
 assign Pg34956 = ( wire4366 ) ;
 assign Pg34839 = ( wire4366 ) ;
 assign Pg34788 = ( wire4376 ) ;
 assign Pg34437 = ( wire4378 ) ;
 assign Pg34436 = ( wire4379 ) ;
 assign Pg33959 = ( wire4394 ) ;
 assign Pg33894 = ( wire4376 ) ;
 assign Pg33533 = ( wire4406 ) ;
 assign Pg31861 = ( wire4415 ) ;
 assign Pg31665 = ( wire4378 ) ;
 assign Pg31656 = ( wire4379 ) ;
 assign Pg30332 = ( wire4421 ) ;
 assign Pg29221 = ( wire4426 ) ;
 assign Pg29220 = ( wire4427 ) ;
 assign Pg29219 = ( wire4428 ) ;
 assign Pg29218 = ( wire4507 ) ;
 assign Pg29217 = ( wire4430 ) ;
 assign Pg29216 = ( wire4431 ) ;
 assign Pg29215 = ( wire4432 ) ;
 assign Pg29214 = ( wire4433 ) ;
 assign Pg29213 = ( wire4434 ) ;
 assign Pg29212 = ( wire4435 ) ;
 assign Pg29211 = ( wire4436 ) ;
 assign Pg29210 = ( wire4437 ) ;
 assign Pg28753 = ( wire4394 ) ;
 assign Pg27831 = ( wire4406 ) ;
 assign Pg25219 = ( wire4415 ) ;
 assign Pg24185 = ( Pg44 ) ;
 assign Pg24184 = ( Pg135 ) ;
 assign Pg24183 = ( Pg134 ) ;
 assign Pg24182 = ( Pg127 ) ;
 assign Pg24181 = ( Pg126 ) ;
 assign Pg24180 = ( Pg125 ) ;
 assign Pg24179 = ( Pg124 ) ;
 assign Pg24178 = ( Pg120 ) ;
 assign Pg24177 = ( Pg116 ) ;
 assign Pg24176 = ( Pg115 ) ;
 assign Pg24175 = ( Pg114 ) ;
 assign Pg24174 = ( Pg113 ) ;
 assign Pg24173 = ( Pg100 ) ;
 assign Pg24172 = ( Pg99 ) ;
 assign Pg24171 = ( Pg92 ) ;
 assign Pg24170 = ( Pg91 ) ;
 assign Pg24169 = ( Pg90 ) ;
 assign Pg24168 = ( Pg84 ) ;
 assign Pg24167 = ( Pg73 ) ;
 assign Pg24166 = ( Pg72 ) ;
 assign Pg24165 = ( Pg64 ) ;
 assign Pg24164 = ( Pg57 ) ;
 assign Pg24163 = ( Pg56 ) ;
 assign Pg24162 = ( Pg54 ) ;
 assign Pg24161 = ( Pg53 ) ;
 assign Pg23683 = ( wire4421 ) ;
 assign Pg21698 = ( Pg36 ) ;
 assign Pg21292 = ( wire4426 ) ;
 assign Pg21270 = ( wire4430 ) ;
 assign Pg21245 = ( wire4427 ) ;
 assign Pg21176 = ( wire4431 ) ;
 assign Pg20901 = ( wire4432 ) ;
 assign Pg20899 = ( wire4435 ) ;
 assign Pg20763 = ( wire4436 ) ;
 assign Pg20654 = ( wire4428 ) ;
 assign Pg20652 = ( wire4433 ) ;
 assign Pg20557 = ( wire4434 ) ;
 assign Pg20049 = ( wire4437 ) ;
 assign Pg18881 = ( wire4507 ) ;
 assign Pg18101 = ( Pg6746 ) ;
 assign Pg18100 = ( Pg6751 ) ;
 assign Pg18099 = ( Pg6745 ) ;
 assign Pg18098 = ( Pg6744 ) ;
 assign Pg18097 = ( Pg6747 ) ;
 assign Pg18096 = ( Pg6750 ) ;
 assign Pg18095 = ( Pg6749 ) ;
 assign Pg18094 = ( Pg6748 ) ;
 assign Pg18092 = ( Pg6753 ) ;
 assign Pg8403 = ( wire4651 ) ;
 assign Pg8353 = ( wire4651 ) ;
 assign Pg8283 = ( wire4658 ) ;
 assign Pg8235 = ( wire4658 ) ;
 assign Pg8178 = ( wire4661 ) ;
 assign Pg8132 = ( wire4661 ) ;


endmodule

