module ex5p_qmap_map (sk, i_4_, i_5_, i_6_, i_7_, i_3_, i_1_, i_0_, i_2_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_, o_41_, o_42_, o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_, o_51_, o_52_, o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_, o_61_, o_62_);

	input i_4_;
	input i_5_;
	input i_6_;
	input i_7_;
	input i_3_;
	input i_1_;
	input i_0_;
	input i_2_;
	output o_0_;
	output o_1_;
	output o_2_;
	output o_3_;
	output o_4_;
	output o_5_;
	output o_6_;
	output o_7_;
	output o_8_;
	output o_9_;
	output o_10_;
	output o_11_;
	output o_12_;
	output o_13_;
	output o_14_;
	output o_15_;
	output o_16_;
	output o_17_;
	output o_18_;
	output o_19_;
	output o_20_;
	output o_21_;
	output o_22_;
	output o_23_;
	output o_24_;
	output o_25_;
	output o_26_;
	output o_27_;
	output o_28_;
	output o_29_;
	output o_30_;
	output o_31_;
	output o_32_;
	output o_33_;
	output o_34_;
	output o_35_;
	output o_36_;
	output o_37_;
	output o_38_;
	output o_39_;
	output o_40_;
	output o_41_;
	output o_42_;
	output o_43_;
	output o_44_;
	output o_45_;
	output o_46_;
	output o_47_;
	output o_48_;
	output o_49_;
	output o_50_;
	output o_51_;
	output o_52_;
	output o_53_;
	output o_54_;
	output o_55_;
	output o_56_;
	output o_57_;
	output o_58_;
	output o_59_;
	output o_60_;
	output o_61_;
	output o_62_;



	wire g1, g3, g5, g7, g10, g14, g18, g20, g22, g24, g26, g28, g30, g32, g33, g34, g35, g37, g40, g41, g42;
	wire g45, g46, g47, g48, g49, g51, g52, g53, g365, g92, g94, g121, g122, g124, g152, g165, g175, g188, g194, g207, g214;
	wire g215, g223, g224, g235, g236, g237, g239, g247, g257, g262, g270, g276, g281, g288, g291, g298, g300, g303, g307, g2, g4;
	wire g6, g8, g9, g12, g13, g15, g16, g17, g19, g21, g23, g25, g27, g29, g31, g36, g38, g39, g44, g50, g54;
	wire g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73, g74, g75;
	wire g76, g77, g78, g79, g80, g81, g82, g83, g354, g84, g85, g86, g87, g88, g89, g90, g91, g93, g95, g96, g97;
	wire g98, g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118;
	wire g119, g120, g123, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g310, g136, g137, g138, g139, g140, g141;
	wire g142, g143, g144, g145, g146, g147, g148, g149, g150, g343, g333, g151, g153, g154, g155, g156, g157, g158, g159, g160, g161;
	wire g162, g163, g164, g166, g167, g168, g169, g170, g171, g172, g173, g174, g176, g177, g178, g179, g180, g181, g182, g183, g184;
	wire g185, g186, g187, g189, g190, g191, g192, g193, g322, g195, g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206;
	wire g311, g208, g209, g210, g211, g212, g213, g216, g217, g218, g219, g220, g221, g222, g225, g226, g227, g228, g229, g230, g231;
	wire g232, g233, g234, g238, g240, g241, g242, g243, g244, g245, g246, g309, g248, g249, g250, g251, g252, g253, g254, g255, g256;
	wire g258, g259, g260, g261, g263, g264, g265, g266, g267, g268, g269, g271, g272, g273, g274, g275, g277, g278, g279, g280, g282;
	wire g283, g284, g285, g286, g287, g289, g290, g292, g293, g294, g295, g296, g297, g299, g308, g301, g302, g304, g305, g306, g312;
	wire g313, g314, g317, g315, g316, g319, g320, g318, g321, g323, g324, g325, g328, g326, g327, g330, g331, g329, g332, g334, g335;
	wire g336, g339, g337, g338, g340, g341, g342, g344, g345, g346, g349, g347, g348, g352, g350, g351, g353, g355, g356, g357, g360;
	wire g358, g359, g362, g363, g361, g364, g366, g367, g368, g369, g370;

	lut_sub lut_5 ({g1}, o_0_);
	defparam lut_5.LUT_SIZE = 1;
	defparam lut_5.mask = 2'b01;

	lut_sub lut_9 ({g3}, o_1_);
	defparam lut_9.LUT_SIZE = 1;
	defparam lut_9.mask = 2'b10;

	lut_sub lut_13 ({g5}, o_2_);
	defparam lut_13.LUT_SIZE = 1;
	defparam lut_13.mask = 2'b10;

	lut_sub lut_17 ({g7}, o_3_);
	defparam lut_17.LUT_SIZE = 1;
	defparam lut_17.mask = 2'b10;

	lut_sub lut_21 ({g10}, o_4_);
	defparam lut_21.LUT_SIZE = 1;
	defparam lut_21.mask = 2'b10;

	lut_sub lut_25 ({g14}, o_6_);
	defparam lut_25.LUT_SIZE = 1;
	defparam lut_25.mask = 2'b10;

	lut_sub lut_29 ({g18}, o_7_);
	defparam lut_29.LUT_SIZE = 1;
	defparam lut_29.mask = 2'b10;

	lut_sub lut_33 ({g20}, o_8_);
	defparam lut_33.LUT_SIZE = 1;
	defparam lut_33.mask = 2'b10;

	lut_sub lut_37 ({g22}, o_9_);
	defparam lut_37.LUT_SIZE = 1;
	defparam lut_37.mask = 2'b10;

	lut_sub lut_41 ({g24}, o_10_);
	defparam lut_41.LUT_SIZE = 1;
	defparam lut_41.mask = 2'b01;

	lut_sub lut_45 ({g26}, o_11_);
	defparam lut_45.LUT_SIZE = 1;
	defparam lut_45.mask = 2'b10;

	lut_sub lut_49 ({g28}, o_12_);
	defparam lut_49.LUT_SIZE = 1;
	defparam lut_49.mask = 2'b10;

	lut_sub lut_53 ({g30}, o_13_);
	defparam lut_53.LUT_SIZE = 1;
	defparam lut_53.mask = 2'b10;

	lut_sub lut_57 ({g32}, o_14_);
	defparam lut_57.LUT_SIZE = 1;
	defparam lut_57.mask = 2'b10;

	lut_sub lut_61 ({g33}, o_15_);
	defparam lut_61.LUT_SIZE = 1;
	defparam lut_61.mask = 2'b10;

	lut_sub lut_65 ({g34}, o_16_);
	defparam lut_65.LUT_SIZE = 1;
	defparam lut_65.mask = 2'b10;

	lut_sub lut_69 ({g35}, o_17_);
	defparam lut_69.LUT_SIZE = 1;
	defparam lut_69.mask = 2'b01;

	lut_sub lut_73 ({g37}, o_18_);
	defparam lut_73.LUT_SIZE = 1;
	defparam lut_73.mask = 2'b10;

	lut_sub lut_77 ({g40}, o_19_);
	defparam lut_77.LUT_SIZE = 1;
	defparam lut_77.mask = 2'b10;

	lut_sub lut_81 ({g41}, o_20_);
	defparam lut_81.LUT_SIZE = 1;
	defparam lut_81.mask = 2'b10;

	lut_sub lut_85 ({g42}, o_21_);
	defparam lut_85.LUT_SIZE = 1;
	defparam lut_85.mask = 2'b10;

	lut_sub lut_89 ({g45}, o_23_);
	defparam lut_89.LUT_SIZE = 1;
	defparam lut_89.mask = 2'b10;

	lut_sub lut_93 ({g46}, o_24_);
	defparam lut_93.LUT_SIZE = 1;
	defparam lut_93.mask = 2'b10;

	lut_sub lut_97 ({g47}, o_25_);
	defparam lut_97.LUT_SIZE = 1;
	defparam lut_97.mask = 2'b10;

	lut_sub lut_101 ({g48}, o_26_);
	defparam lut_101.LUT_SIZE = 1;
	defparam lut_101.mask = 2'b01;

	lut_sub lut_105 ({g49}, o_27_);
	defparam lut_105.LUT_SIZE = 1;
	defparam lut_105.mask = 2'b10;

	lut_sub lut_109 ({g51}, o_28_);
	defparam lut_109.LUT_SIZE = 1;
	defparam lut_109.mask = 2'b10;

	lut_sub lut_113 ({g52}, o_29_);
	defparam lut_113.LUT_SIZE = 1;
	defparam lut_113.mask = 2'b10;

	lut_sub lut_117 ({g53}, o_30_);
	defparam lut_117.LUT_SIZE = 1;
	defparam lut_117.mask = 2'b10;

	lut_sub lut_121 ({g365}, o_31_);
	defparam lut_121.LUT_SIZE = 1;
	defparam lut_121.mask = 2'b10;

	lut_sub lut_125 ({g92}, o_32_);
	defparam lut_125.LUT_SIZE = 1;
	defparam lut_125.mask = 2'b10;

	lut_sub lut_129 ({g94}, o_33_);
	defparam lut_129.LUT_SIZE = 1;
	defparam lut_129.mask = 2'b10;

	lut_sub lut_133 ({g121}, o_34_);
	defparam lut_133.LUT_SIZE = 1;
	defparam lut_133.mask = 2'b10;

	lut_sub lut_137 ({g122}, o_35_);
	defparam lut_137.LUT_SIZE = 1;
	defparam lut_137.mask = 2'b10;

	lut_sub lut_141 ({g124}, o_36_);
	defparam lut_141.LUT_SIZE = 1;
	defparam lut_141.mask = 2'b10;

	lut_sub lut_145 ({g152}, o_37_);
	defparam lut_145.LUT_SIZE = 1;
	defparam lut_145.mask = 2'b10;

	lut_sub lut_149 ({g165}, o_38_);
	defparam lut_149.LUT_SIZE = 1;
	defparam lut_149.mask = 2'b10;

	lut_sub lut_153 ({g175}, o_39_);
	defparam lut_153.LUT_SIZE = 1;
	defparam lut_153.mask = 2'b10;

	lut_sub lut_157 ({g188}, o_40_);
	defparam lut_157.LUT_SIZE = 1;
	defparam lut_157.mask = 2'b10;

	lut_sub lut_161 ({g194}, o_41_);
	defparam lut_161.LUT_SIZE = 1;
	defparam lut_161.mask = 2'b10;

	lut_sub lut_165 ({g207}, o_42_);
	defparam lut_165.LUT_SIZE = 1;
	defparam lut_165.mask = 2'b10;

	lut_sub lut_169 ({g214}, o_43_);
	defparam lut_169.LUT_SIZE = 1;
	defparam lut_169.mask = 2'b10;

	lut_sub lut_173 ({g215}, o_44_);
	defparam lut_173.LUT_SIZE = 1;
	defparam lut_173.mask = 2'b10;

	lut_sub lut_177 ({g223}, o_45_);
	defparam lut_177.LUT_SIZE = 1;
	defparam lut_177.mask = 2'b10;

	lut_sub lut_181 ({g224}, o_46_);
	defparam lut_181.LUT_SIZE = 1;
	defparam lut_181.mask = 2'b10;

	lut_sub lut_185 ({g235}, o_47_);
	defparam lut_185.LUT_SIZE = 1;
	defparam lut_185.mask = 2'b10;

	lut_sub lut_189 ({g236}, o_48_);
	defparam lut_189.LUT_SIZE = 1;
	defparam lut_189.mask = 2'b10;

	lut_sub lut_193 ({g237}, o_49_);
	defparam lut_193.LUT_SIZE = 1;
	defparam lut_193.mask = 2'b10;

	lut_sub lut_197 ({g239}, o_50_);
	defparam lut_197.LUT_SIZE = 1;
	defparam lut_197.mask = 2'b10;

	lut_sub lut_201 ({g247}, o_51_);
	defparam lut_201.LUT_SIZE = 1;
	defparam lut_201.mask = 2'b10;

	lut_sub lut_205 ({g257}, o_52_);
	defparam lut_205.LUT_SIZE = 1;
	defparam lut_205.mask = 2'b10;

	lut_sub lut_209 ({g262}, o_53_);
	defparam lut_209.LUT_SIZE = 1;
	defparam lut_209.mask = 2'b10;

	lut_sub lut_213 ({g270}, o_54_);
	defparam lut_213.LUT_SIZE = 1;
	defparam lut_213.mask = 2'b10;

	lut_sub lut_217 ({g276}, o_55_);
	defparam lut_217.LUT_SIZE = 1;
	defparam lut_217.mask = 2'b10;

	lut_sub lut_221 ({g281}, o_56_);
	defparam lut_221.LUT_SIZE = 1;
	defparam lut_221.mask = 2'b10;

	lut_sub lut_225 ({g288}, o_57_);
	defparam lut_225.LUT_SIZE = 1;
	defparam lut_225.mask = 2'b10;

	lut_sub lut_229 ({g291}, o_58_);
	defparam lut_229.LUT_SIZE = 1;
	defparam lut_229.mask = 2'b10;

	lut_sub lut_233 ({g298}, o_59_);
	defparam lut_233.LUT_SIZE = 1;
	defparam lut_233.mask = 2'b10;

	lut_sub lut_237 ({g300}, o_60_);
	defparam lut_237.LUT_SIZE = 1;
	defparam lut_237.mask = 2'b10;

	lut_sub lut_241 ({g303}, o_61_);
	defparam lut_241.LUT_SIZE = 1;
	defparam lut_241.mask = 2'b10;

	lut_sub lut_245 ({g307}, o_62_);
	defparam lut_245.LUT_SIZE = 1;
	defparam lut_245.mask = 2'b10;

	lut_sub lut_249 ({i_4_, i_5_, i_6_}, g1);
	defparam lut_249.LUT_SIZE = 3;
	defparam lut_249.mask = 8'h80;

	lut_sub lut_253 ({i_6_, i_7_}, g2);
	defparam lut_253.LUT_SIZE = 2;
	defparam lut_253.mask = 4'b1000;

	lut_sub lut_258 ({i_5_, g2}, g3);
	defparam lut_258.LUT_SIZE = 2;
	defparam lut_258.mask = 4'b1011;

	lut_sub lut_264 ({i_4_, i_5_, i_3_}, g4);
	defparam lut_264.LUT_SIZE = 3;
	defparam lut_264.mask = 8'h20;

	lut_sub lut_270 ({g2, g4}, g5);
	defparam lut_270.LUT_SIZE = 2;
	defparam lut_270.mask = 4'b1110;

	lut_sub lut_276 ({i_4_, i_5_, i_3_}, g6);
	defparam lut_276.LUT_SIZE = 3;
	defparam lut_276.mask = 8'h10;

	lut_sub lut_282 ({g2, g6}, g7);
	defparam lut_282.LUT_SIZE = 2;
	defparam lut_282.mask = 4'b1110;

	lut_sub lut_288 ({i_4_, i_5_, i_3_}, g8);
	defparam lut_288.LUT_SIZE = 3;
	defparam lut_288.mask = 8'h40;

	lut_sub lut_292 ({i_6_, i_7_}, g9);
	defparam lut_292.LUT_SIZE = 2;
	defparam lut_292.mask = 4'b0010;

	lut_sub lut_298 ({g8, g9}, g10);
	defparam lut_298.LUT_SIZE = 2;
	defparam lut_298.mask = 4'b1110;

	lut_sub lut_305 ({i_4_, i_5_, g9}, o_5_);
	defparam lut_305.LUT_SIZE = 3;
	defparam lut_305.mask = 8'h10;

	lut_sub lut_310 ({i_6_, g8}, g12);
	defparam lut_310.LUT_SIZE = 2;
	defparam lut_310.mask = 4'b0100;

	lut_sub lut_314 ({i_1_, i_0_, i_2_}, g13);
	defparam lut_314.LUT_SIZE = 3;
	defparam lut_314.mask = 8'h40;

	lut_sub lut_320 ({g12, g13}, g14);
	defparam lut_320.LUT_SIZE = 2;
	defparam lut_320.mask = 4'b1110;

	lut_sub lut_326 ({i_6_, i_7_}, g15);
	defparam lut_326.LUT_SIZE = 2;
	defparam lut_326.mask = 4'b0001;

	lut_sub lut_332 ({g4, g15}, g16);
	defparam lut_332.LUT_SIZE = 2;
	defparam lut_332.mask = 4'b0001;

	lut_sub lut_336 ({i_1_, i_0_, i_2_}, g17);
	defparam lut_336.LUT_SIZE = 3;
	defparam lut_336.mask = 8'h08;

	lut_sub lut_342 ({g16, g17}, g18);
	defparam lut_342.LUT_SIZE = 2;
	defparam lut_342.mask = 4'b1110;

	lut_sub lut_348 ({i_1_, i_0_, i_2_}, g19);
	defparam lut_348.LUT_SIZE = 3;
	defparam lut_348.mask = 8'h01;

	lut_sub lut_354 ({g16, g19}, g20);
	defparam lut_354.LUT_SIZE = 2;
	defparam lut_354.mask = 4'b1110;

	lut_sub lut_360 ({i_4_, i_5_, i_3_}, g21);
	defparam lut_360.LUT_SIZE = 3;
	defparam lut_360.mask = 8'h80;

	lut_sub lut_367 ({g13, g15, g21}, g22);
	defparam lut_367.LUT_SIZE = 3;
	defparam lut_367.mask = 8'hfe;

	lut_sub lut_377 ({i_1_, i_0_, i_2_}, g23);
	defparam lut_377.LUT_SIZE = 3;
	defparam lut_377.mask = 8'hfb;

	lut_sub lut_389 ({i_4_, i_5_, g15, g23}, g24);
	defparam lut_389.LUT_SIZE = 4;
	defparam lut_389.mask = 16'h0200;

	lut_sub lut_393 ({i_1_, i_0_, i_2_}, g25);
	defparam lut_393.LUT_SIZE = 3;
	defparam lut_393.mask = 8'hfd;

	lut_sub lut_405 ({g16, g25}, g26);
	defparam lut_405.LUT_SIZE = 2;
	defparam lut_405.mask = 4'b1101;

	lut_sub lut_411 ({i_1_, i_0_, i_2_}, g27);
	defparam lut_411.LUT_SIZE = 3;
	defparam lut_411.mask = 8'hef;

	lut_sub lut_423 ({g16, g27}, g28);
	defparam lut_423.LUT_SIZE = 2;
	defparam lut_423.mask = 4'b1101;

	lut_sub lut_431 ({g6, g15}, g29);
	defparam lut_431.LUT_SIZE = 2;
	defparam lut_431.mask = 4'b0001;

	lut_sub lut_437 ({g17, g29}, g30);
	defparam lut_437.LUT_SIZE = 2;
	defparam lut_437.mask = 4'b1110;

	lut_sub lut_443 ({i_1_, i_0_, i_2_}, g31);
	defparam lut_443.LUT_SIZE = 3;
	defparam lut_443.mask = 8'hdf;

	lut_sub lut_455 ({g29, g31}, g32);
	defparam lut_455.LUT_SIZE = 2;
	defparam lut_455.mask = 4'b1101;

	lut_sub lut_463 ({g23, g29}, g33);
	defparam lut_463.LUT_SIZE = 2;
	defparam lut_463.mask = 4'b1011;

	lut_sub lut_471 ({g25, g29}, g34);
	defparam lut_471.LUT_SIZE = 2;
	defparam lut_471.mask = 4'b1011;

	lut_sub lut_478 ({i_4_, i_5_, g31}, g35);
	defparam lut_478.LUT_SIZE = 3;
	defparam lut_478.mask = 8'h08;

	lut_sub lut_482 ({i_4_, i_3_}, g36);
	defparam lut_482.LUT_SIZE = 2;
	defparam lut_482.mask = 4'b0001;

	lut_sub lut_488 ({i_5_, g13, g36}, g37);
	defparam lut_488.LUT_SIZE = 3;
	defparam lut_488.mask = 8'hef;

	lut_sub lut_498 ({i_4_, i_3_}, g38);
	defparam lut_498.LUT_SIZE = 2;
	defparam lut_498.mask = 4'b0010;

	lut_sub lut_502 ({i_1_, i_0_, i_2_}, g39);
	defparam lut_502.LUT_SIZE = 3;
	defparam lut_502.mask = 8'h80;

	lut_sub lut_508 ({g38, g39}, g40);
	defparam lut_508.LUT_SIZE = 2;
	defparam lut_508.mask = 4'b1110;

	lut_sub lut_516 ({i_6_, g21, g31}, g41);
	defparam lut_516.LUT_SIZE = 3;
	defparam lut_516.mask = 8'hdf;

	lut_sub lut_528 ({g12, g31}, g42);
	defparam lut_528.LUT_SIZE = 2;
	defparam lut_528.mask = 4'b1101;

	lut_sub lut_536 ({i_4_, i_5_, g15, g31}, o_22_);
	defparam lut_536.LUT_SIZE = 4;
	defparam lut_536.mask = 16'h2000;

	lut_sub lut_540 ({i_4_, i_5_, i_3_}, g44);
	defparam lut_540.LUT_SIZE = 3;
	defparam lut_540.mask = 8'h01;

	lut_sub lut_547 ({g6, g39, g44}, g45);
	defparam lut_547.LUT_SIZE = 3;
	defparam lut_547.mask = 8'hec;

	lut_sub lut_558 ({g9, g21, g39}, g46);
	defparam lut_558.LUT_SIZE = 3;
	defparam lut_558.mask = 8'hfe;

	lut_sub lut_571 ({g9, g17, g21}, g47);
	defparam lut_571.LUT_SIZE = 3;
	defparam lut_571.mask = 8'hfe;

	lut_sub lut_583 ({i_0_, i_2_, g15, g21}, g48);
	defparam lut_583.LUT_SIZE = 4;
	defparam lut_583.mask = 16'h0001;

	lut_sub lut_590 ({g9, g21, g23}, g49);
	defparam lut_590.LUT_SIZE = 3;
	defparam lut_590.mask = 8'hfd;

	lut_sub lut_602 ({g8, g15}, g50);
	defparam lut_602.LUT_SIZE = 2;
	defparam lut_602.mask = 4'b0001;

	lut_sub lut_608 ({g27, g50}, g51);
	defparam lut_608.LUT_SIZE = 2;
	defparam lut_608.mask = 4'b1011;

	lut_sub lut_616 ({i_6_, i_7_, g21, g39}, g52);
	defparam lut_616.LUT_SIZE = 4;
	defparam lut_616.mask = 16'hfeff;

	lut_sub lut_637 ({g15, g19, g21}, g53);
	defparam lut_637.LUT_SIZE = 3;
	defparam lut_637.mask = 8'hfe;

	lut_sub lut_650 ({i_6_, i_7_, g6, g21, g27}, g54);
	defparam lut_650.LUT_SIZE = 5;
	defparam lut_650.mask = 32'h2f2f2f00;

	lut_sub lut_671 ({i_6_, g6, g36, g39}, g55);
	defparam lut_671.LUT_SIZE = 4;
	defparam lut_671.mask = 16'h1115;

	lut_sub lut_680 ({i_4_, i_5_, i_6_, i_7_, i_3_, g13}, g56);
	defparam lut_680.LUT_SIZE = 6;
	defparam lut_680.mask = 64'h1145444444444444;

	lut_sub lut_703 ({i_6_, g13, g21, g56}, g57);
	defparam lut_703.LUT_SIZE = 4;
	defparam lut_703.mask = 16'ha8aa;

	lut_sub lut_715 ({g55, g57}, g58);
	defparam lut_715.LUT_SIZE = 2;
	defparam lut_715.mask = 4'b0100;

	lut_sub lut_722 ({g27, g29, g36}, g59);
	defparam lut_722.LUT_SIZE = 3;
	defparam lut_722.mask = 8'h70;

	lut_sub lut_730 ({i_5_, g12, g38}, g60);
	defparam lut_730.LUT_SIZE = 3;
	defparam lut_730.mask = 8'hc8;

	lut_sub lut_739 ({i_6_, i_7_, g4, g21, g25}, g61);
	defparam lut_739.LUT_SIZE = 5;
	defparam lut_739.mask = 32'h000f2f22;

	lut_sub lut_755 ({g5, g61}, g62);
	defparam lut_755.LUT_SIZE = 2;
	defparam lut_755.mask = 4'b0010;

	lut_sub lut_760 ({i_4_, i_5_, i_6_, i_7_, i_3_, g19}, g63);
	defparam lut_760.LUT_SIZE = 6;
	defparam lut_760.mask = 64'h5571000044444444;

	lut_sub lut_785 ({g27, g50, g53, g60, g62, g63}, g64);
	defparam lut_785.LUT_SIZE = 6;
	defparam lut_785.mask = 64'h0002000000220022;

	lut_sub lut_795 ({i_6_, i_7_, g6, g27}, g65);
	defparam lut_795.LUT_SIZE = 4;
	defparam lut_795.mask = 16'h0220;

	lut_sub lut_801 ({i_4_, i_5_, i_6_, i_7_, i_3_, g25}, g66);
	defparam lut_801.LUT_SIZE = 6;
	defparam lut_801.mask = 64'haa02222aaaaa8888;

	lut_sub lut_831 ({g15, g21, g25, g27, g44}, g67);
	defparam lut_831.LUT_SIZE = 5;
	defparam lut_831.mask = 32'h505050dc;

	lut_sub lut_846 ({i_4_, i_5_, i_6_, i_7_, i_3_, g19}, g68);
	defparam lut_846.LUT_SIZE = 6;
	defparam lut_846.mask = 64'h0000111511111111;

	lut_sub lut_866 ({i_5_, g16, g27, g38, g68}, g69);
	defparam lut_866.LUT_SIZE = 5;
	defparam lut_866.mask = 32'h8a0aaa0a;

	lut_sub lut_886 ({g59, g64, g65, g66, g67, g69}, g70);
	defparam lut_886.LUT_SIZE = 6;
	defparam lut_886.mask = 64'h0000400000000000;

	lut_sub lut_893 ({i_6_, i_7_, g4, g21, g31}, g71);
	defparam lut_893.LUT_SIZE = 5;
	defparam lut_893.mask = 32'h000a2a22;

	lut_sub lut_906 ({g5, g31, g71}, g72);
	defparam lut_906.LUT_SIZE = 3;
	defparam lut_906.mask = 8'h2a;

	lut_sub lut_915 ({g15, g21, g23}, g73);
	defparam lut_915.LUT_SIZE = 3;
	defparam lut_915.mask = 8'h02;

	lut_sub lut_922 ({i_6_, g21, g23, g30}, g74);
	defparam lut_922.LUT_SIZE = 4;
	defparam lut_922.mask = 16'h5155;

	lut_sub lut_935 ({g17, g36, g49}, g75);
	defparam lut_935.LUT_SIZE = 3;
	defparam lut_935.mask = 8'h54;

	lut_sub lut_945 ({i_6_, i_7_, g6, g21, g23, g31}, g76);
	defparam lut_945.LUT_SIZE = 6;
	defparam lut_945.mask = 64'h0a0a0ace00000000;

	lut_sub lut_960 ({i_4_, i_5_, i_3_, g15}, g77);
	defparam lut_960.LUT_SIZE = 4;
	defparam lut_960.mask = 16'h04c0;

	lut_sub lut_968 ({g31, g77}, g78);
	defparam lut_968.LUT_SIZE = 2;
	defparam lut_968.mask = 4'b0100;

	lut_sub lut_974 ({g2, g8}, g79);
	defparam lut_974.LUT_SIZE = 2;
	defparam lut_974.mask = 4'b1110;

	lut_sub lut_981 ({i_7_, g8}, g80);
	defparam lut_981.LUT_SIZE = 2;
	defparam lut_981.mask = 4'b0001;

	lut_sub lut_989 ({g17, g38, g79, g80}, g81);
	defparam lut_989.LUT_SIZE = 4;
	defparam lut_989.mask = 16'h00df;

	lut_sub lut_1003 ({g12, g16, g23, g38}, g82);
	defparam lut_1003.LUT_SIZE = 4;
	defparam lut_1003.mask = 16'h4ccc;

	lut_sub lut_1016 ({g78, g81, g82}, g83);
	defparam lut_1016.LUT_SIZE = 3;
	defparam lut_1016.mask = 8'h80;

	lut_sub lut_1026 ({g72, g73, g74, g75, g354, g83}, g84);
	defparam lut_1026.LUT_SIZE = 6;
	defparam lut_1026.mask = 64'h0000000000010000;

	lut_sub lut_1032 ({i_6_, i_7_, g4, g39}, g85);
	defparam lut_1032.LUT_SIZE = 4;
	defparam lut_1032.mask = 16'h0111;

	lut_sub lut_1041 ({g5, g39, g85}, g86);
	defparam lut_1041.LUT_SIZE = 3;
	defparam lut_1041.mask = 8'h8a;

	lut_sub lut_1051 ({g12, g38, g39, g86}, g87);
	defparam lut_1051.LUT_SIZE = 4;
	defparam lut_1051.mask = 16'h5444;

	lut_sub lut_1062 ({i_6_, i_7_, g6, g8, g39}, g88);
	defparam lut_1062.LUT_SIZE = 5;
	defparam lut_1062.mask = 32'h05050011;

	lut_sub lut_1074 ({i_6_, i_7_, g17, g21, g39}, g89);
	defparam lut_1074.LUT_SIZE = 5;
	defparam lut_1074.mask = 32'h13130313;

	lut_sub lut_1093 ({g13, g29, g31, g50, g89}, g90);
	defparam lut_1093.LUT_SIZE = 5;
	defparam lut_1093.mask = 32'h8a8a8a00;

	lut_sub lut_1110 ({g18, g35, g87, g88, g90}, g91);
	defparam lut_1110.LUT_SIZE = 5;
	defparam lut_1110.mask = 32'h00000400;

	lut_sub lut_1120 ({g32, g54, g58, g70, g84, g91}, g92);
	defparam lut_1120.LUT_SIZE = 6;
	defparam lut_1120.mask = 64'h0000000000010000;

	lut_sub lut_1124 ({i_5_, i_3_, i_1_}, g93);
	defparam lut_1124.LUT_SIZE = 3;
	defparam lut_1124.mask = 8'h1a;

	lut_sub lut_1132 ({i_4_, i_0_, i_2_, g15, g93}, g94);
	defparam lut_1132.LUT_SIZE = 5;
	defparam lut_1132.mask = 32'h00020000;

	lut_sub lut_1138 ({g17, g21}, g95);
	defparam lut_1138.LUT_SIZE = 2;
	defparam lut_1138.mask = 4'b0001;

	lut_sub lut_1146 ({g13, g29, g36, g95}, g96);
	defparam lut_1146.LUT_SIZE = 4;
	defparam lut_1146.mask = 16'haa80;

	lut_sub lut_1156 ({g18, g96}, g97);
	defparam lut_1156.LUT_SIZE = 2;
	defparam lut_1156.mask = 4'b0001;

	lut_sub lut_1165 ({g12, g16, g25, g31, g44}, g98);
	defparam lut_1165.LUT_SIZE = 5;
	defparam lut_1165.mask = 32'hbb0b0b0b;

	lut_sub lut_1186 ({i_6_, i_7_, g13, g21, g39}, g99);
	defparam lut_1186.LUT_SIZE = 5;
	defparam lut_1186.mask = 32'h13131100;

	lut_sub lut_1200 ({g55, g98, g99}, g100);
	defparam lut_1200.LUT_SIZE = 3;
	defparam lut_1200.mask = 8'h20;

	lut_sub lut_1206 ({i_6_, g21, g25}, g101);
	defparam lut_1206.LUT_SIZE = 3;
	defparam lut_1206.mask = 8'h20;

	lut_sub lut_1212 ({i_1_, i_0_, i_2_, g50, g101}, g102);
	defparam lut_1212.LUT_SIZE = 5;
	defparam lut_1212.mask = 32'h8aaaa88a;

	lut_sub lut_1233 ({g16, g19, g29, g36, g102}, g103);
	defparam lut_1233.LUT_SIZE = 5;
	defparam lut_1233.mask = 32'h55405500;

	lut_sub lut_1246 ({i_4_, i_5_, i_6_, i_7_, i_3_, g39}, g104);
	defparam lut_1246.LUT_SIZE = 6;
	defparam lut_1246.mask = 64'h1104044444444444;

	lut_sub lut_1265 ({i_4_, i_5_, i_3_, g15, g27}, g105);
	defparam lut_1265.LUT_SIZE = 5;
	defparam lut_1265.mask = 32'h2020a000;

	lut_sub lut_1274 ({i_4_, i_5_, g2, i_3_, g25}, g106);
	defparam lut_1274.LUT_SIZE = 5;
	defparam lut_1274.mask = 32'h0020aaee;

	lut_sub lut_1293 ({g27, g29, g36, g105, g106}, g107);
	defparam lut_1293.LUT_SIZE = 5;
	defparam lut_1293.mask = 32'h80008888;

	lut_sub lut_1306 ({g64, g100, g103, g104, g107}, g108);
	defparam lut_1306.LUT_SIZE = 5;
	defparam lut_1306.mask = 32'h00000004;

	lut_sub lut_1314 ({i_6_, g17, g21, g23, g44}, g109);
	defparam lut_1314.LUT_SIZE = 5;
	defparam lut_1314.mask = 32'h0c5d0055;

	lut_sub lut_1331 ({i_5_, g17, g36, g109}, g110);
	defparam lut_1331.LUT_SIZE = 4;
	defparam lut_1331.mask = 16'ha8aa;

	lut_sub lut_1343 ({i_6_, i_7_, g6, g17}, g111);
	defparam lut_1343.LUT_SIZE = 4;
	defparam lut_1343.mask = 16'h0111;

	lut_sub lut_1350 ({i_4_, i_5_, i_6_, i_7_, i_3_, g23}, g112);
	defparam lut_1350.LUT_SIZE = 6;
	defparam lut_1350.mask = 64'h2288000888880000;

	lut_sub lut_1363 ({i_4_, i_5_, i_6_, i_7_, i_3_, g31}, g113);
	defparam lut_1363.LUT_SIZE = 6;
	defparam lut_1363.mask = 64'h0200033800000000;

	lut_sub lut_1376 ({g110, g111, g112, g113}, g114);
	defparam lut_1376.LUT_SIZE = 4;
	defparam lut_1376.mask = 16'h0080;

	lut_sub lut_1382 ({g15, g21}, g115);
	defparam lut_1382.LUT_SIZE = 2;
	defparam lut_1382.mask = 4'b0100;

	lut_sub lut_1390 ({i_4_, g23, g29, g31, g115}, g116);
	defparam lut_1390.LUT_SIZE = 5;
	defparam lut_1390.mask = 32'hb0bb00bb;

	lut_sub lut_1410 ({g27, g115}, g117);
	defparam lut_1410.LUT_SIZE = 2;
	defparam lut_1410.mask = 4'b0100;

	lut_sub lut_1418 ({g12, g13, g38, g50}, g118);
	defparam lut_1418.LUT_SIZE = 4;
	defparam lut_1418.mask = 16'h070f;

	lut_sub lut_1433 ({g13, g16, g29, g31, g79}, g119);
	defparam lut_1433.LUT_SIZE = 5;
	defparam lut_1433.mask = 32'h73737300;

	lut_sub lut_1456 ({g22, g117, g118, g81, g119}, g120);
	defparam lut_1456.LUT_SIZE = 5;
	defparam lut_1456.mask = 32'h00004000;

	lut_sub lut_1465 ({g97, g108, g114, g116, g120}, g121);
	defparam lut_1465.LUT_SIZE = 5;
	defparam lut_1465.mask = 32'h00000001;

	lut_sub lut_1469 ({i_4_, i_5_, i_3_, i_1_, i_0_, i_2_}, g122);
	defparam lut_1469.LUT_SIZE = 6;
	defparam lut_1469.mask = 64'h000000008000a060;

	lut_sub lut_1478 ({i_4_, i_3_, g9, i_0_, i_2_}, g123);
	defparam lut_1478.LUT_SIZE = 5;
	defparam lut_1478.mask = 32'h04002222;

	lut_sub lut_1487 ({i_5_, i_1_, g123}, g124);
	defparam lut_1487.LUT_SIZE = 3;
	defparam lut_1487.mask = 8'h40;

	lut_sub lut_1495 ({i_6_, g5, g21, g23, g38}, g125);
	defparam lut_1495.LUT_SIZE = 5;
	defparam lut_1495.mask = 32'hcc44cc4c;

	lut_sub lut_1514 ({i_6_, i_7_, g4, g23, g109}, g126);
	defparam lut_1514.LUT_SIZE = 5;
	defparam lut_1514.mask = 32'haaa2a2aa;

	lut_sub lut_1535 ({g16, g23, g125, g126}, g127);
	defparam lut_1535.LUT_SIZE = 4;
	defparam lut_1535.mask = 16'h4404;

	lut_sub lut_1544 ({g23, g79, g127}, g128);
	defparam lut_1544.LUT_SIZE = 3;
	defparam lut_1544.mask = 8'h15;

	lut_sub lut_1552 ({i_6_, i_7_, g19, g21}, g129);
	defparam lut_1552.LUT_SIZE = 4;
	defparam lut_1552.mask = 16'h1110;

	lut_sub lut_1560 ({g53, g129}, g130);
	defparam lut_1560.LUT_SIZE = 2;
	defparam lut_1560.mask = 4'b0010;

	lut_sub lut_1568 ({g27, g31, g50, g59}, g131);
	defparam lut_1568.LUT_SIZE = 4;
	defparam lut_1568.mask = 16'h888a;

	lut_sub lut_1582 ({g19, g38, g72, g130, g354, g131}, g132);
	defparam lut_1582.LUT_SIZE = 6;
	defparam lut_1582.mask = 64'h0001000100010000;

	lut_sub lut_1590 ({i_6_, i_7_, g6, g13}, g133);
	defparam lut_1590.LUT_SIZE = 4;
	defparam lut_1590.mask = 16'h1110;

	lut_sub lut_1599 ({i_6_, g4, g17, g38}, g134);
	defparam lut_1599.LUT_SIZE = 4;
	defparam lut_1599.mask = 16'h1113;

	lut_sub lut_1609 ({i_6_, g8, g17}, g135);
	defparam lut_1609.LUT_SIZE = 3;
	defparam lut_1609.mask = 8'h10;

	lut_sub lut_1615 ({g133, g310}, g136);
	defparam lut_1615.LUT_SIZE = 2;
	defparam lut_1615.mask = 4'b1000;

	lut_sub lut_1622 ({g13, g29, g36}, g137);
	defparam lut_1622.LUT_SIZE = 3;
	defparam lut_1622.mask = 8'h07;

	lut_sub lut_1631 ({i_6_, i_7_, g4, g21, g27}, g138);
	defparam lut_1631.LUT_SIZE = 5;
	defparam lut_1631.mask = 32'h0a002222;

	lut_sub lut_1644 ({i_5_, g31, g36, g137, g138}, g139);
	defparam lut_1644.LUT_SIZE = 5;
	defparam lut_1644.mask = 32'h80888888;

	lut_sub lut_1657 ({i_6_, i_7_, g6, g8, g27}, g140);
	defparam lut_1657.LUT_SIZE = 5;
	defparam lut_1657.mask = 32'h2a220000;

	lut_sub lut_1669 ({i_1_, i_0_, g50, g136, g139, g140}, g141);
	defparam lut_1669.LUT_SIZE = 6;
	defparam lut_1669.mask = 64'h0200020202020202;

	lut_sub lut_1683 ({g2, g6, g25, g50}, g142);
	defparam lut_1683.LUT_SIZE = 4;
	defparam lut_1683.mask = 16'h4c44;

	lut_sub lut_1696 ({g7, g23, g78, g65, g142}, g143);
	defparam lut_1696.LUT_SIZE = 5;
	defparam lut_1696.mask = 32'h00808080;

	lut_sub lut_1706 ({g2, g4, g27, g38}, g144);
	defparam lut_1706.LUT_SIZE = 4;
	defparam lut_1706.mask = 16'h4c44;

	lut_sub lut_1718 ({i_5_, g12, g31, g38, g144}, g145);
	defparam lut_1718.LUT_SIZE = 5;
	defparam lut_1718.mask = 32'haa0a8a0a;

	lut_sub lut_1733 ({i_6_, i_7_, g8, i_1_, i_0_, i_2_}, g146);
	defparam lut_1733.LUT_SIZE = 6;
	defparam lut_1733.mask = 64'h004300c700000000;

	lut_sub lut_1745 ({i_4_, i_5_, i_6_, i_7_, i_3_, g17}, g147);
	defparam lut_1745.LUT_SIZE = 6;
	defparam lut_1745.mask = 64'h0001111111110000;

	lut_sub lut_1760 ({i_6_, g21, g27, g147}, g148);
	defparam lut_1760.LUT_SIZE = 4;
	defparam lut_1760.mask = 16'ha2aa;

	lut_sub lut_1770 ({i_4_, i_5_, i_3_, i_1_, i_0_, i_2_}, g149);
	defparam lut_1770.LUT_SIZE = 6;
	defparam lut_1770.mask = 64'h7fff7ffffffdbffd;

	lut_sub lut_1833 ({i_4_, i_5_, i_6_, i_7_, i_3_, g19}, g150);
	defparam lut_1833.LUT_SIZE = 6;
	defparam lut_1833.mask = 64'hfffeaaaaeeeeeeee;

	lut_sub lut_1888 ({g343, g145, g146, g148, g333}, g151);
	defparam lut_1888.LUT_SIZE = 5;
	defparam lut_1888.mask = 32'h00000010;

	lut_sub lut_1897 ({g128, g132, g141, g143, g151}, g152);
	defparam lut_1897.LUT_SIZE = 5;
	defparam lut_1897.mask = 32'h00000001;

	lut_sub lut_1905 ({g5, g16, g31, g71}, g153);
	defparam lut_1905.LUT_SIZE = 4;
	defparam lut_1905.mask = 16'h22a2;

	lut_sub lut_1918 ({g7, g17, g36, g50, g111}, g154);
	defparam lut_1918.LUT_SIZE = 5;
	defparam lut_1918.mask = 32'haa00aa80;

	lut_sub lut_1931 ({i_4_, i_5_, i_6_, i_3_, g23}, g155);
	defparam lut_1931.LUT_SIZE = 5;
	defparam lut_1931.mask = 32'h000222aa;

	lut_sub lut_1945 ({g31, g41, g50, g155}, g156);
	defparam lut_1945.LUT_SIZE = 4;
	defparam lut_1945.mask = 16'h080a;

	lut_sub lut_1952 ({i_4_, i_5_, i_6_, i_7_, i_3_, g23}, g157);
	defparam lut_1952.LUT_SIZE = 6;
	defparam lut_1952.mask = 64'h228aa20888880000;

	lut_sub lut_1974 ({g126, g310, g153, g154, g156, g157}, g158);
	defparam lut_1974.LUT_SIZE = 6;
	defparam lut_1974.mask = 64'h0000000000020000;

	lut_sub lut_1982 ({g15, g21, g39, g86}, g159);
	defparam lut_1982.LUT_SIZE = 4;
	defparam lut_1982.mask = 16'h5554;

	lut_sub lut_1994 ({i_4_, i_3_, g13, g15}, g160);
	defparam lut_1994.LUT_SIZE = 4;
	defparam lut_1994.mask = 16'h0100;

	lut_sub lut_2002 ({g38, g39, g79, g80}, g161);
	defparam lut_2002.LUT_SIZE = 4;
	defparam lut_2002.mask = 16'h0d0f;

	lut_sub lut_2015 ({i_4_, i_5_, i_3_, g13, g15, g39}, g162);
	defparam lut_2015.LUT_SIZE = 6;
	defparam lut_2015.mask = 64'h0f00031100550055;

	lut_sub lut_2039 ({g12, g13, g38, g161, g162}, g163);
	defparam lut_2039.LUT_SIZE = 5;
	defparam lut_2039.mask = 32'h88808800;

	lut_sub lut_2052 ({i_6_, g21, g39, g159, g160, g163}, g164);
	defparam lut_2052.LUT_SIZE = 6;
	defparam lut_2052.mask = 64'h0404040004040404;

	lut_sub lut_2067 ({g32, g54, g70, g158, g164}, g165);
	defparam lut_2067.LUT_SIZE = 5;
	defparam lut_2067.mask = 32'h00000100;

	lut_sub lut_2075 ({g17, g74, g75, g60}, g166);
	defparam lut_2075.LUT_SIZE = 4;
	defparam lut_2075.mask = 16'h0301;

	lut_sub lut_2084 ({i_6_, i_7_, g6, g21, g31}, g167);
	defparam lut_2084.LUT_SIZE = 5;
	defparam lut_2084.mask = 32'h000f2f00;

	lut_sub lut_2100 ({i_6_, g6, g23, g36, g117}, g168);
	defparam lut_2100.LUT_SIZE = 5;
	defparam lut_2100.mask = 32'h8a8a8a0a;

	lut_sub lut_2119 ({g13, g29, g82, g167, g168}, g169);
	defparam lut_2119.LUT_SIZE = 5;
	defparam lut_2119.mask = 32'h40404000;

	lut_sub lut_2128 ({g13, g36, g95}, g170);
	defparam lut_2128.LUT_SIZE = 3;
	defparam lut_2128.mask = 8'ha8;

	lut_sub lut_2137 ({g17, g77, g170}, g171);
	defparam lut_2137.LUT_SIZE = 3;
	defparam lut_2137.mask = 8'h54;

	lut_sub lut_2146 ({g17, g50, g73}, g172);
	defparam lut_2146.LUT_SIZE = 3;
	defparam lut_2146.mask = 8'ha8;

	lut_sub lut_2153 ({i_4_, i_5_, i_6_, i_7_, g31}, g173);
	defparam lut_2153.LUT_SIZE = 5;
	defparam lut_2153.mask = 32'ha002aa00;

	lut_sub lut_2167 ({g56, g171, g172, g173}, g174);
	defparam lut_2167.LUT_SIZE = 4;
	defparam lut_2167.mask = 16'h0200;

	lut_sub lut_2175 ({g166, g108, g169, g174}, g175);
	defparam lut_2175.LUT_SIZE = 4;
	defparam lut_2175.mask = 16'h0001;

	lut_sub lut_2183 ({i_5_, g29, g31, g36, g54}, g176);
	defparam lut_2183.LUT_SIZE = 5;
	defparam lut_2183.mask = 32'h8a0aaa0a;

	lut_sub lut_2200 ({g39, g50, g343}, g177);
	defparam lut_2200.LUT_SIZE = 3;
	defparam lut_2200.mask = 8'h54;

	lut_sub lut_2207 ({i_4_, i_5_, i_6_, i_7_, i_3_, g19}, g178);
	defparam lut_2207.LUT_SIZE = 6;
	defparam lut_2207.mask = 64'h1131155155555555;

	lut_sub lut_2241 ({g20, g62, g177, g178}, g179);
	defparam lut_2241.LUT_SIZE = 4;
	defparam lut_2241.mask = 16'h0002;

	lut_sub lut_2250 ({g12, g13, g38, g39, g50}, g180);
	defparam lut_2250.LUT_SIZE = 5;
	defparam lut_2250.mask = 32'hffa0cc00;

	lut_sub lut_2268 ({i_4_, i_5_, i_6_, i_7_, i_3_, g27}, g181);
	defparam lut_2268.LUT_SIZE = 6;
	defparam lut_2268.mask = 64'h2232222222222222;

	lut_sub lut_2290 ({g144, g181}, g182);
	defparam lut_2290.LUT_SIZE = 2;
	defparam lut_2290.mask = 4'b1000;

	lut_sub lut_2297 ({i_6_, i_7_, g6, g8, g17}, g183);
	defparam lut_2297.LUT_SIZE = 5;
	defparam lut_2297.mask = 32'h05050515;

	lut_sub lut_2313 ({g16, g17, g39, g77}, g184);
	defparam lut_2313.LUT_SIZE = 4;
	defparam lut_2313.mask = 16'h0537;

	lut_sub lut_2323 ({i_4_, i_5_, i_3_, i_1_, i_0_, i_2_}, g185);
	defparam lut_2323.LUT_SIZE = 6;
	defparam lut_2323.mask = 64'h06060606260e0606;

	lut_sub lut_2349 ({g17, g60, g183, g184, g185}, g186);
	defparam lut_2349.LUT_SIZE = 5;
	defparam lut_2349.mask = 32'h80800080;

	lut_sub lut_2360 ({g129, g153, g180, g182, g186}, g187);
	defparam lut_2360.LUT_SIZE = 5;
	defparam lut_2360.mask = 32'h00010000;

	lut_sub lut_2369 ({g128, g176, g90, g179, g187}, g188);
	defparam lut_2369.LUT_SIZE = 5;
	defparam lut_2369.mask = 32'h00000001;

	lut_sub lut_2376 ({i_6_, g8, g31, g38}, g189);
	defparam lut_2376.LUT_SIZE = 4;
	defparam lut_2376.mask = 16'h4c44;

	lut_sub lut_2388 ({g57, g189, g88, g158}, g190);
	defparam lut_2388.LUT_SIZE = 4;
	defparam lut_2388.mask = 16'h0040;

	lut_sub lut_2396 ({g21, g39, g87, g178}, g191);
	defparam lut_2396.LUT_SIZE = 4;
	defparam lut_2396.mask = 16'h2220;

	lut_sub lut_2407 ({g5, g19, g25, g44, g130}, g192);
	defparam lut_2407.LUT_SIZE = 5;
	defparam lut_2407.mask = 32'h45004545;

	lut_sub lut_2424 ({g20, g55, g133, g182, g192}, g193);
	defparam lut_2424.LUT_SIZE = 5;
	defparam lut_2424.mask = 32'h00001000;

	lut_sub lut_2433 ({g139, g190, g191, g322, g193}, g194);
	defparam lut_2433.LUT_SIZE = 5;
	defparam lut_2433.mask = 32'h00000001;

	lut_sub lut_2439 ({i_4_, i_5_, i_3_, g13, g39}, g195);
	defparam lut_2439.LUT_SIZE = 5;
	defparam lut_2439.mask = 32'h30000505;

	lut_sub lut_2453 ({g16, g29, g31, g39, g195}, g196);
	defparam lut_2453.LUT_SIZE = 5;
	defparam lut_2453.mask = 32'haa880a08;

	lut_sub lut_2467 ({i_6_, i_7_, g4, g31}, g197);
	defparam lut_2467.LUT_SIZE = 4;
	defparam lut_2467.mask = 16'h0220;

	lut_sub lut_2477 ({g13, g77, g197, g63, g180}, g198);
	defparam lut_2477.LUT_SIZE = 5;
	defparam lut_2477.mask = 32'h40404000;

	lut_sub lut_2488 ({g61, g172, g103, g196, g198}, g199);
	defparam lut_2488.LUT_SIZE = 5;
	defparam lut_2488.mask = 32'h00010000;

	lut_sub lut_2496 ({g12, g23, g27, g60}, g200);
	defparam lut_2496.LUT_SIZE = 4;
	defparam lut_2496.mask = 16'h88f8;

	lut_sub lut_2511 ({g16, g25, g38, g189, g200}, g201);
	defparam lut_2511.LUT_SIZE = 5;
	defparam lut_2511.mask = 32'h80880088;

	lut_sub lut_2523 ({i_6_, i_7_, g6, g21, g27, g137}, g202);
	defparam lut_2523.LUT_SIZE = 6;
	defparam lut_2523.mask = 64'haaaaaa00a2a2aaaa;

	lut_sub lut_2555 ({g21, g38, g39}, g203);
	defparam lut_2555.LUT_SIZE = 3;
	defparam lut_2555.mask = 8'h15;

	lut_sub lut_2566 ({i_5_, g16, g23, g27, g38, g203}, g204);
	defparam lut_2566.LUT_SIZE = 6;
	defparam lut_2566.mask = 64'h888a000aaaaa000a;

	lut_sub lut_2592 ({g12, g25, g27, g29, g36, g204}, g205);
	defparam lut_2592.LUT_SIZE = 6;
	defparam lut_2592.mask = 64'h4040405500004055;

	lut_sub lut_2612 ({g48, g95, g184, g116, g205}, g206);
	defparam lut_2612.LUT_SIZE = 5;
	defparam lut_2612.mask = 32'h10000000;

	lut_sub lut_2622 ({g166, g199, g311, g201, g202, g206}, g207);
	defparam lut_2622.LUT_SIZE = 6;
	defparam lut_2622.mask = 64'h0000000000000001;

	lut_sub lut_2629 ({g12, g25, g38}, g208);
	defparam lut_2629.LUT_SIZE = 3;
	defparam lut_2629.mask = 8'h4c;

	lut_sub lut_2638 ({g110, g135, g208}, g209);
	defparam lut_2638.LUT_SIZE = 3;
	defparam lut_2638.mask = 8'h08;

	lut_sub lut_2645 ({g49, g144, g111}, g210);
	defparam lut_2645.LUT_SIZE = 3;
	defparam lut_2645.mask = 8'h08;

	lut_sub lut_2653 ({g12, g27, g29, g36}, g211);
	defparam lut_2653.LUT_SIZE = 4;
	defparam lut_2653.mask = 16'h70f0;

	lut_sub lut_2665 ({i_4_, i_5_, i_6_, i_3_, g25, g32}, g212);
	defparam lut_2665.LUT_SIZE = 6;
	defparam lut_2665.mask = 64'h5555555151515151;

	lut_sub lut_2701 ({g26, g85, g134, g211, g89, g212}, g213);
	defparam lut_2701.LUT_SIZE = 6;
	defparam lut_2701.mask = 64'h0000000040000000;

	lut_sub lut_2710 ({g169, g199, g209, g210, g213}, g214);
	defparam lut_2710.LUT_SIZE = 5;
	defparam lut_2710.mask = 32'h00000001;

	lut_sub lut_2715 ({i_4_, i_3_, i_1_, i_0_, i_2_, g1}, g215);
	defparam lut_2715.LUT_SIZE = 6;
	defparam lut_2715.mask = 64'h04000000c4000000;

	lut_sub lut_2725 ({i_4_, i_3_, g12, g13, g15}, g216);
	defparam lut_2725.LUT_SIZE = 5;
	defparam lut_2725.mask = 32'h03130303;

	lut_sub lut_2740 ({g13, g38, g216}, g217);
	defparam lut_2740.LUT_SIZE = 3;
	defparam lut_2740.mask = 8'ha8;

	lut_sub lut_2750 ({g171, g87, g162, g217}, g218);
	defparam lut_2750.LUT_SIZE = 4;
	defparam lut_2750.mask = 16'h0004;

	lut_sub lut_2757 ({g31, g44, g176}, g219);
	defparam lut_2757.LUT_SIZE = 3;
	defparam lut_2757.mask = 8'h45;

	lut_sub lut_2767 ({g23, g31, g41, g50}, g220);
	defparam lut_2767.LUT_SIZE = 4;
	defparam lut_2767.mask = 16'h2223;

	lut_sub lut_2779 ({g39, g115, g189, g220}, g221);
	defparam lut_2779.LUT_SIZE = 4;
	defparam lut_2779.mask = 16'h4440;

	lut_sub lut_2789 ({i_6_, g21, g23, g153, g24}, g222);
	defparam lut_2789.LUT_SIZE = 5;
	defparam lut_2789.mask = 32'h22222202;

	lut_sub lut_2805 ({g17, g218, g219, g70, g221, g222}, g223);
	defparam lut_2805.LUT_SIZE = 6;
	defparam lut_2805.mask = 64'h0000000100000000;

	lut_sub lut_2811 ({i_4_, i_5_, i_3_, g9, g17}, g224);
	defparam lut_2811.LUT_SIZE = 5;
	defparam lut_2811.mask = 32'h40005050;

	lut_sub lut_2821 ({g51, g53}, g225);
	defparam lut_2821.LUT_SIZE = 2;
	defparam lut_2821.mask = 4'b0001;

	lut_sub lut_2827 ({g62, g101}, g226);
	defparam lut_2827.LUT_SIZE = 2;
	defparam lut_2827.mask = 4'b0010;

	lut_sub lut_2836 ({g20, g23, g25, g36, g50}, g227);
	defparam lut_2836.LUT_SIZE = 5;
	defparam lut_2836.mask = 32'h00008acf;

	lut_sub lut_2852 ({g7, g19, g27, g36}, g228);
	defparam lut_2852.LUT_SIZE = 4;
	defparam lut_2852.mask = 16'hcd05;

	lut_sub lut_2868 ({g26, g63, g211, g208, g76, g228}, g229);
	defparam lut_2868.LUT_SIZE = 6;
	defparam lut_2868.mask = 64'h0000000080000000;

	lut_sub lut_2878 ({g71, g225, g226, g143, g227, g229}, g230);
	defparam lut_2878.LUT_SIZE = 6;
	defparam lut_2878.mask = 64'h0000000100000000;

	lut_sub lut_2885 ({i_6_, i_7_, g6, g8, g31}, g231);
	defparam lut_2885.LUT_SIZE = 5;
	defparam lut_2885.mask = 32'h0f0f0022;

	lut_sub lut_2902 ({g12, g38, g39, g115}, g232);
	defparam lut_2902.LUT_SIZE = 4;
	defparam lut_2902.mask = 16'h1333;

	lut_sub lut_2917 ({g138, g145, g311, g231, g232}, g233);
	defparam lut_2917.LUT_SIZE = 5;
	defparam lut_2917.mask = 32'h00080000;

	lut_sub lut_2927 ({g49, g86, g73, g137, g24, g154}, g234);
	defparam lut_2927.LUT_SIZE = 6;
	defparam lut_2927.mask = 64'h0000000000004000;

	lut_sub lut_2936 ({g58, g136, g230, g233, g234}, g235);
	defparam lut_2936.LUT_SIZE = 5;
	defparam lut_2936.mask = 32'h00000001;

	lut_sub lut_2945 ({i_3_, g39, g137, g219, g70, g190}, g236);
	defparam lut_2945.LUT_SIZE = 6;
	defparam lut_2945.mask = 64'h0100000001000100;

	lut_sub lut_2954 ({g13, g38, g1}, g237);
	defparam lut_2954.LUT_SIZE = 3;
	defparam lut_2954.mask = 8'h07;

	lut_sub lut_2960 ({i_3_, i_1_, i_0_}, g238);
	defparam lut_2960.LUT_SIZE = 3;
	defparam lut_2960.mask = 8'h54;

	lut_sub lut_2968 ({i_4_, i_5_, i_2_, g15, g238}, g239);
	defparam lut_2968.LUT_SIZE = 5;
	defparam lut_2968.mask = 32'h20000000;

	lut_sub lut_2976 ({g138, g145, g311, g231}, g240);
	defparam lut_2976.LUT_SIZE = 4;
	defparam lut_2976.mask = 16'h0200;

	lut_sub lut_2983 ({i_6_, g19, g21, g62}, g241);
	defparam lut_2983.LUT_SIZE = 4;
	defparam lut_2983.mask = 16'h5554;

	lut_sub lut_2998 ({g12, g25, g29, g36, g50}, g242);
	defparam lut_2998.LUT_SIZE = 5;
	defparam lut_2998.mask = 32'h7f00ff00;

	lut_sub lut_3019 ({g181, g241, g242}, g243);
	defparam lut_3019.LUT_SIZE = 3;
	defparam lut_3019.mask = 8'h20;

	lut_sub lut_3026 ({g16, g21, g38}, g244);
	defparam lut_3026.LUT_SIZE = 3;
	defparam lut_3026.mask = 8'h80;

	lut_sub lut_3032 ({i_4_, i_5_, i_3_, g15, g19}, g245);
	defparam lut_3032.LUT_SIZE = 5;
	defparam lut_3032.mask = 32'h01100000;

	lut_sub lut_3042 ({g19, g29, g39, g244, g245}, g246);
	defparam lut_3042.LUT_SIZE = 5;
	defparam lut_3042.mask = 32'ha2a0a200;

	lut_sub lut_3058 ({g97, g84, g240, g243, g309}, g247);
	defparam lut_3058.LUT_SIZE = 5;
	defparam lut_3058.mask = 32'h00000001;

	lut_sub lut_3064 ({i_4_, i_3_, g13, g15}, g248);
	defparam lut_3064.LUT_SIZE = 4;
	defparam lut_3064.mask = 16'h1000;

	lut_sub lut_3069 ({i_4_, i_5_, i_6_, i_7_, i_3_, g19}, g249);
	defparam lut_3069.LUT_SIZE = 6;
	defparam lut_3069.mask = 64'h1131000111111111;

	lut_sub lut_3087 ({i_4_, i_5_, i_6_, i_7_, i_3_, g31}, g250);
	defparam lut_3087.LUT_SIZE = 6;
	defparam lut_3087.mask = 64'h2000b002aaaa8888;

	lut_sub lut_3111 ({g9, g13, g19, g21}, g251);
	defparam lut_3111.LUT_SIZE = 4;
	defparam lut_3111.mask = 16'h0015;

	lut_sub lut_3121 ({g249, g156, g250, g251}, g252);
	defparam lut_3121.LUT_SIZE = 4;
	defparam lut_3121.mask = 16'h0800;

	lut_sub lut_3130 ({g71, g225, g114, g227, g252}, g253);
	defparam lut_3130.LUT_SIZE = 5;
	defparam lut_3130.mask = 32'h00010000;

	lut_sub lut_3139 ({g7, g17, g50, g62, g142}, g254);
	defparam lut_3139.LUT_SIZE = 5;
	defparam lut_3139.mask = 32'h22002220;

	lut_sub lut_3152 ({g2, g4, g27, g29, g36}, g255);
	defparam lut_3152.LUT_SIZE = 5;
	defparam lut_3152.mask = 32'h70f07070;

	lut_sub lut_3172 ({g29, g39, g244, g255}, g256);
	defparam lut_3172.LUT_SIZE = 4;
	defparam lut_3172.mask = 16'ha2a0;

	lut_sub lut_3186 ({g248, g98, g141, g253, g254, g256}, g257);
	defparam lut_3186.LUT_SIZE = 6;
	defparam lut_3186.mask = 64'h0000000100000000;

	lut_sub lut_3196 ({g13, g21, g39, g50, g170, g163}, g258);
	defparam lut_3196.LUT_SIZE = 6;
	defparam lut_3196.mask = 64'h1111110010101000;

	lut_sub lut_3213 ({g10, g17, g38, g183, g142}, g259);
	defparam lut_3213.LUT_SIZE = 5;
	defparam lut_3213.mask = 32'h00008880;

	lut_sub lut_3222 ({i_6_, g16, g21, g23}, g260);
	defparam lut_3222.LUT_SIZE = 4;
	defparam lut_3222.mask = 16'h0a2a;

	lut_sub lut_3235 ({g219, g226, g245, g259, g260}, g261);
	defparam lut_3235.LUT_SIZE = 5;
	defparam lut_3235.mask = 32'h00000020;

	lut_sub lut_3244 ({g105, g132, g201, g258, g261}, g262);
	defparam lut_3244.LUT_SIZE = 5;
	defparam lut_3244.mask = 32'h00010000;

	lut_sub lut_3251 ({i_6_, i_7_, g6, g27, g31}, g263);
	defparam lut_3251.LUT_SIZE = 5;
	defparam lut_3251.mask = 32'h10101011;

	lut_sub lut_3263 ({i_6_, i_7_, g8, g21, g27, g263}, g264);
	defparam lut_3263.LUT_SIZE = 6;
	defparam lut_3263.mask = 64'h5111511151515555;

	lut_sub lut_3293 ({g25, g36, g264}, g265);
	defparam lut_3293.LUT_SIZE = 3;
	defparam lut_3293.mask = 8'h45;

	lut_sub lut_3302 ({g18, g47, g118}, g266);
	defparam lut_3302.LUT_SIZE = 3;
	defparam lut_3302.mask = 8'h02;

	lut_sub lut_3311 ({g23, g50, g101, g130, g266}, g267);
	defparam lut_3311.LUT_SIZE = 5;
	defparam lut_3311.mask = 32'h10001010;

	lut_sub lut_3320 ({i_4_, i_5_, i_3_, g13, g15, g17}, g268);
	defparam lut_3320.LUT_SIZE = 6;
	defparam lut_3320.mask = 64'h11000003000f000f;

	lut_sub lut_3340 ({g125, g88, g195, g209, g268}, g269);
	defparam lut_3340.LUT_SIZE = 5;
	defparam lut_3340.mask = 32'h20000000;

	lut_sub lut_3349 ({g265, g191, g254, g267, g269}, g270);
	defparam lut_3349.LUT_SIZE = 5;
	defparam lut_3349.mask = 32'h00000001;

	lut_sub lut_3357 ({g15, g21, g39, g268}, g271);
	defparam lut_3357.LUT_SIZE = 4;
	defparam lut_3357.mask = 16'haaa8;

	lut_sub lut_3371 ({g219, g221, g266, g271}, g272);
	defparam lut_3371.LUT_SIZE = 4;
	defparam lut_3371.mask = 16'h0001;

	lut_sub lut_3381 ({g16, g38, g39, g60, g105, g101}, g273);
	defparam lut_3381.LUT_SIZE = 6;
	defparam lut_3381.mask = 64'h8808880088008800;

	lut_sub lut_3396 ({i_4_, i_3_, g16, g19, g25}, g274);
	defparam lut_3396.LUT_SIZE = 5;
	defparam lut_3396.mask = 32'h0a0aaa3b;

	lut_sub lut_3417 ({g142, g183, g222, g273, g274}, g275);
	defparam lut_3417.LUT_SIZE = 5;
	defparam lut_3417.mask = 32'h02000000;

	lut_sub lut_3426 ({g59, g64, g177, g272, g275}, g276);
	defparam lut_3426.LUT_SIZE = 5;
	defparam lut_3426.mask = 32'h00010000;

	lut_sub lut_3432 ({i_6_, g17, g21}, g277);
	defparam lut_3432.LUT_SIZE = 3;
	defparam lut_3432.mask = 8'h10;

	lut_sub lut_3437 ({i_4_, i_3_, i_1_, i_0_, i_2_, g79}, g278);
	defparam lut_3437.LUT_SIZE = 6;
	defparam lut_3437.mask = 64'h80008000c0c08030;

	lut_sub lut_3454 ({g12, g23, g39, g80, g278}, g279);
	defparam lut_3454.LUT_SIZE = 5;
	defparam lut_3454.mask = 32'ha8a800a8;

	lut_sub lut_3471 ({g85, g71, g277, g125, g279}, g280);
	defparam lut_3471.LUT_SIZE = 5;
	defparam lut_3471.mask = 32'h40000000;

	lut_sub lut_3480 ({g74, g70, g196, g272, g280}, g281);
	defparam lut_3480.LUT_SIZE = 5;
	defparam lut_3480.mask = 32'h00000001;

	lut_sub lut_3487 ({g73, g74, g75}, g282);
	defparam lut_3487.LUT_SIZE = 3;
	defparam lut_3487.mask = 8'h10;

	lut_sub lut_3495 ({g2, g6, g25, g38}, g283);
	defparam lut_3495.LUT_SIZE = 4;
	defparam lut_3495.mask = 16'h4c44;

	lut_sub lut_3505 ({i_4_, i_3_, g13, g23}, g284);
	defparam lut_3505.LUT_SIZE = 4;
	defparam lut_3505.mask = 16'h00ab;

	lut_sub lut_3516 ({g26, g283, g284}, g285);
	defparam lut_3516.LUT_SIZE = 3;
	defparam lut_3516.mask = 8'h08;

	lut_sub lut_3524 ({i_6_, i_7_, g6, g8, g17, g23}, g286);
	defparam lut_3524.LUT_SIZE = 6;
	defparam lut_3524.mask = 64'h0bab0bab00000303;

	lut_sub lut_3552 ({g39, g60, g244, g285, g286}, g287);
	defparam lut_3552.LUT_SIZE = 5;
	defparam lut_3552.mask = 32'h22220002;

	lut_sub lut_3565 ({g282, g264, g179, g267, g287}, g288);
	defparam lut_3565.LUT_SIZE = 5;
	defparam lut_3565.mask = 32'h00000001;

	lut_sub lut_3573 ({g17, g60, g127, g147}, g289);
	defparam lut_3573.LUT_SIZE = 4;
	defparam lut_3573.mask = 16'h2202;

	lut_sub lut_3582 ({g21, g33, g39}, g290);
	defparam lut_3582.LUT_SIZE = 3;
	defparam lut_3582.mask = 8'h32;

	lut_sub lut_3593 ({g218, g230, g240, g289, g290}, g291);
	defparam lut_3593.LUT_SIZE = 5;
	defparam lut_3593.mask = 32'h00000001;

	lut_sub lut_3600 ({i_6_, i_7_, g8, g17, g21}, g292);
	defparam lut_3600.LUT_SIZE = 5;
	defparam lut_3600.mask = 32'h11131100;

	lut_sub lut_3613 ({i_5_, g17, g38, g79}, g293);
	defparam lut_3613.LUT_SIZE = 4;
	defparam lut_3613.mask = 16'h0a0b;

	lut_sub lut_3624 ({i_4_, i_5_, i_3_, g15, g17, g27}, g294);
	defparam lut_3624.LUT_SIZE = 6;
	defparam lut_3624.mask = 64'h0000030a0000aa00;

	lut_sub lut_3638 ({i_4_, i_5_, i_3_, g13, g15, g17}, g295);
	defparam lut_3638.LUT_SIZE = 6;
	defparam lut_3638.mask = 64'h000003005f0f5f0f;

	lut_sub lut_3667 ({g293, g216, g294, g295}, g296);
	defparam lut_3667.LUT_SIZE = 4;
	defparam lut_3667.mask = 16'h8000;

	lut_sub lut_3676 ({g117, g62, g283, g292, g296}, g297);
	defparam lut_3676.LUT_SIZE = 5;
	defparam lut_3676.mask = 32'h00400000;

	lut_sub lut_3684 ({g100, g253, g273, g297}, g298);
	defparam lut_3684.LUT_SIZE = 4;
	defparam lut_3684.mask = 16'h0001;

	lut_sub lut_3691 ({g20, g26, g249}, g299);
	defparam lut_3691.LUT_SIZE = 3;
	defparam lut_3691.mask = 8'h02;

	lut_sub lut_3700 ({g84, g240, g243, g258, g308}, g300);
	defparam lut_3700.LUT_SIZE = 5;
	defparam lut_3700.mask = 32'h00000001;

	lut_sub lut_3707 ({g10, g51, g118}, g301);
	defparam lut_3707.LUT_SIZE = 3;
	defparam lut_3707.mask = 8'h02;

	lut_sub lut_3716 ({g159, g66, g192, g294, g301}, g302);
	defparam lut_3716.LUT_SIZE = 5;
	defparam lut_3716.mask = 32'h00000400;

	lut_sub lut_3725 ({g96, g84, g179, g233, g302}, g303);
	defparam lut_3725.LUT_SIZE = 5;
	defparam lut_3725.mask = 32'h00000001;

	lut_sub lut_3732 ({g171, g162, g217}, g304);
	defparam lut_3732.LUT_SIZE = 3;
	defparam lut_3732.mask = 8'h04;

	lut_sub lut_3738 ({i_3_, g12, i_1_, i_0_, i_2_, g142}, g305);
	defparam lut_3738.LUT_SIZE = 6;
	defparam lut_3738.mask = 64'h2a8a2a82aa8aaa82;

	lut_sub lut_3770 ({g39, g79, g80, g241, g305}, g306);
	defparam lut_3770.LUT_SIZE = 5;
	defparam lut_3770.mask = 32'h11110010;

	lut_sub lut_3783 ({g304, g265, g289, g299, g306}, g307);
	defparam lut_3783.LUT_SIZE = 5;
	defparam lut_3783.mask = 32'h00000001;

	lut_sub lut_3792 ({g25, g21, g19, i_6_, g299, g18}, g308);
	defparam lut_3792.LUT_SIZE = 6;
	defparam lut_3792.mask = 64'h1111010111111101;

	lut_sub lut_3810 ({i_2_, i_3_, g246, g50, i_0_, i_1_}, g309);
	defparam lut_3810.LUT_SIZE = 6;
	defparam lut_3810.mask = 64'h00f700f7007700f7;

	lut_sub lut_3841 ({i_3_, i_5_, i_4_, i_6_, g17}, g310);
	defparam lut_3841.LUT_SIZE = 5;
	defparam lut_3841.mask = 32'h55554000;

	lut_sub lut_3855 ({g312, g313}, g311);
	defparam lut_3855.LUT_SIZE = 2;
	defparam lut_3855.mask = 4'b1000;

	lut_sub lut_3860 ({i_6_, g314}, g312);
	defparam lut_3860.LUT_SIZE = 2;
	defparam lut_3860.mask = 4'b0100;

	lut_sub lut_3865 ({i_6_, g317}, g313);
	defparam lut_3865.LUT_SIZE = 2;
	defparam lut_3865.mask = 4'b0001;

	lut_sub lut_3871 ({g315, g316}, g314);
	defparam lut_3871.LUT_SIZE = 2;
	defparam lut_3871.mask = 4'b1000;

	lut_sub lut_3876 ({i_3_, g319}, g315);
	defparam lut_3876.LUT_SIZE = 2;
	defparam lut_3876.mask = 4'b0100;

	lut_sub lut_3881 ({i_3_, g320}, g316);
	defparam lut_3881.LUT_SIZE = 2;
	defparam lut_3881.mask = 4'b0001;

	lut_sub lut_3886 ({i_3_, g318}, g317);
	defparam lut_3886.LUT_SIZE = 2;
	defparam lut_3886.mask = 4'b0010;

	lut_sub lut_3891 ({i_3_, g321}, g318);
	defparam lut_3891.LUT_SIZE = 2;
	defparam lut_3891.mask = 4'b0001;

	lut_sub lut_3896 ({i_5_, g27, i_4_}, g319);
	defparam lut_3896.LUT_SIZE = 3;
	defparam lut_3896.mask = 8'h7f;

	lut_sub lut_3907 ({g31, i_4_}, g320);
	defparam lut_3907.LUT_SIZE = 2;
	defparam lut_3907.mask = 4'b1011;

	lut_sub lut_3914 ({i_7_, i_5_, g31, i_4_}, g321);
	defparam lut_3914.LUT_SIZE = 4;
	defparam lut_3914.mask = 16'hb1b3;

	lut_sub lut_3928 ({g323, g324}, g322);
	defparam lut_3928.LUT_SIZE = 2;
	defparam lut_3928.mask = 4'b1000;

	lut_sub lut_3933 ({i_6_, g325}, g323);
	defparam lut_3933.LUT_SIZE = 2;
	defparam lut_3933.mask = 4'b0100;

	lut_sub lut_3938 ({i_6_, g328}, g324);
	defparam lut_3938.LUT_SIZE = 2;
	defparam lut_3938.mask = 4'b0001;

	lut_sub lut_3944 ({g326, g327}, g325);
	defparam lut_3944.LUT_SIZE = 2;
	defparam lut_3944.mask = 4'b1000;

	lut_sub lut_3949 ({i_3_, g330}, g326);
	defparam lut_3949.LUT_SIZE = 2;
	defparam lut_3949.mask = 4'b0100;

	lut_sub lut_3954 ({i_3_, g331}, g327);
	defparam lut_3954.LUT_SIZE = 2;
	defparam lut_3954.mask = 4'b0001;

	lut_sub lut_3959 ({i_3_, g329}, g328);
	defparam lut_3959.LUT_SIZE = 2;
	defparam lut_3959.mask = 4'b0010;

	lut_sub lut_3964 ({i_3_, g332}, g329);
	defparam lut_3964.LUT_SIZE = 2;
	defparam lut_3964.mask = 4'b0001;

	lut_sub lut_3969 ({i_5_, i_4_, g27}, g330);
	defparam lut_3969.LUT_SIZE = 3;
	defparam lut_3969.mask = 8'h7f;

	lut_sub lut_3980 ({i_5_, i_4_, g25}, g331);
	defparam lut_3980.LUT_SIZE = 3;
	defparam lut_3980.mask = 8'h57;

	lut_sub lut_3989 ({i_5_, i_4_, i_7_, g25}, g332);
	defparam lut_3989.LUT_SIZE = 4;
	defparam lut_3989.mask = 16'hd55f;

	lut_sub lut_4005 ({g334, g335}, g333);
	defparam lut_4005.LUT_SIZE = 2;
	defparam lut_4005.mask = 4'b1000;

	lut_sub lut_4011 ({g39, g336}, g334);
	defparam lut_4011.LUT_SIZE = 2;
	defparam lut_4011.mask = 4'b0100;

	lut_sub lut_4017 ({g39, g339}, g335);
	defparam lut_4017.LUT_SIZE = 2;
	defparam lut_4017.mask = 4'b0001;

	lut_sub lut_4023 ({g337, g338}, g336);
	defparam lut_4023.LUT_SIZE = 2;
	defparam lut_4023.mask = 4'b1000;

	lut_sub lut_4029 ({g7, g340}, g337);
	defparam lut_4029.LUT_SIZE = 2;
	defparam lut_4029.mask = 4'b0100;

	lut_sub lut_4035 ({g7, g341}, g338);
	defparam lut_4035.LUT_SIZE = 2;
	defparam lut_4035.mask = 4'b0001;

	lut_sub lut_4041 ({g7, g342}, g339);
	defparam lut_4041.LUT_SIZE = 2;
	defparam lut_4041.mask = 4'b0001;

	lut_sub lut_4048 ({g149, g150, g25}, g340);
	defparam lut_4048.LUT_SIZE = 3;
	defparam lut_4048.mask = 8'h01;

	lut_sub lut_4054 ({g149, g150}, g341);
	defparam lut_4054.LUT_SIZE = 2;
	defparam lut_4054.mask = 4'b0001;

	lut_sub lut_4062 ({g149, g150, g38, g79}, g342);
	defparam lut_4062.LUT_SIZE = 4;
	defparam lut_4062.mask = 16'h0004;

	lut_sub lut_4068 ({g344, g345}, g343);
	defparam lut_4068.LUT_SIZE = 2;
	defparam lut_4068.mask = 4'b1000;

	lut_sub lut_4073 ({i_4_, g346}, g344);
	defparam lut_4073.LUT_SIZE = 2;
	defparam lut_4073.mask = 4'b0100;

	lut_sub lut_4078 ({i_4_, g349}, g345);
	defparam lut_4078.LUT_SIZE = 2;
	defparam lut_4078.mask = 4'b0001;

	lut_sub lut_4084 ({g347, g348}, g346);
	defparam lut_4084.LUT_SIZE = 2;
	defparam lut_4084.mask = 4'b1000;

	lut_sub lut_4089 ({i_3_, g13}, g347);
	defparam lut_4089.LUT_SIZE = 2;
	defparam lut_4089.mask = 4'b1000;

	lut_sub lut_4094 ({i_3_, g352}, g348);
	defparam lut_4094.LUT_SIZE = 2;
	defparam lut_4094.mask = 4'b0001;

	lut_sub lut_4100 ({g350, g351}, g349);
	defparam lut_4100.LUT_SIZE = 2;
	defparam lut_4100.mask = 4'b1000;

	lut_sub lut_4105 ({i_3_, g353}, g350);
	defparam lut_4105.LUT_SIZE = 2;
	defparam lut_4105.mask = 4'b0100;

	lut_sub lut_4110 ({i_3_, g39}, g351);
	defparam lut_4110.LUT_SIZE = 2;
	defparam lut_4110.mask = 4'b0010;

	lut_sub lut_4115 ({g39, i_7_, i_6_, i_5_}, g352);
	defparam lut_4115.LUT_SIZE = 4;
	defparam lut_4115.mask = 16'hffea;

	lut_sub lut_4132 ({g13, i_5_}, g353);
	defparam lut_4132.LUT_SIZE = 2;
	defparam lut_4132.mask = 4'b1101;

	lut_sub lut_4140 ({g355, g356}, g354);
	defparam lut_4140.LUT_SIZE = 2;
	defparam lut_4140.mask = 4'b1000;

	lut_sub lut_4146 ({g23, g357}, g355);
	defparam lut_4146.LUT_SIZE = 2;
	defparam lut_4146.mask = 4'b0100;

	lut_sub lut_4152 ({g23, g360}, g356);
	defparam lut_4152.LUT_SIZE = 2;
	defparam lut_4152.mask = 4'b0001;

	lut_sub lut_4158 ({g358, g359}, g357);
	defparam lut_4158.LUT_SIZE = 2;
	defparam lut_4158.mask = 4'b1000;

	lut_sub lut_4163 ({i_3_, g362}, g358);
	defparam lut_4163.LUT_SIZE = 2;
	defparam lut_4163.mask = 4'b0100;

	lut_sub lut_4168 ({i_3_, g363}, g359);
	defparam lut_4168.LUT_SIZE = 2;
	defparam lut_4168.mask = 4'b0001;

	lut_sub lut_4173 ({i_3_, g361}, g360);
	defparam lut_4173.LUT_SIZE = 2;
	defparam lut_4173.mask = 4'b1000;

	lut_sub lut_4178 ({i_3_, g364}, g361);
	defparam lut_4178.LUT_SIZE = 2;
	defparam lut_4178.mask = 4'b0100;

	lut_sub lut_4183 ({i_5_, i_6_, g31, i_4_}, g362);
	defparam lut_4183.LUT_SIZE = 4;
	defparam lut_4183.mask = 16'h7fff;

	lut_sub lut_4201 ({i_5_, i_6_, i_7_, i_4_}, g363);
	defparam lut_4201.LUT_SIZE = 4;
	defparam lut_4201.mask = 16'ha880;

	lut_sub lut_4209 ({i_5_, i_6_, g31, i_4_}, g364);
	defparam lut_4209.LUT_SIZE = 4;
	defparam lut_4209.mask = 16'h7fff;

	lut_sub lut_4228 ({i_1_, g366}, g365);
	defparam lut_4228.LUT_SIZE = 2;
	defparam lut_4228.mask = 4'b0100;

	lut_sub lut_4234 ({g367, g368}, g366);
	defparam lut_4234.LUT_SIZE = 2;
	defparam lut_4234.mask = 4'b1000;

	lut_sub lut_4239 ({i_5_, g369}, g367);
	defparam lut_4239.LUT_SIZE = 2;
	defparam lut_4239.mask = 4'b0100;

	lut_sub lut_4244 ({i_5_, g370}, g368);
	defparam lut_4244.LUT_SIZE = 2;
	defparam lut_4244.mask = 4'b0001;

	lut_sub lut_4248 ({i_4_, i_2_, i_6_, i_0_}, g369);
	defparam lut_4248.LUT_SIZE = 4;
	defparam lut_4248.mask = 16'h4000;

	lut_sub lut_4252 ({i_4_, i_2_, i_3_, i_0_}, g370);
	defparam lut_4252.LUT_SIZE = 4;
	defparam lut_4252.mask = 16'h00d2;


endmodule