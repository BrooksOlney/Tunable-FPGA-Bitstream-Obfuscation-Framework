module apex2 (
	i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, 
	i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, 
	i_18_, i_19_, i_20_, i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, 
	i_28_, i_29_, i_30_, i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, 
	i_38_, o_0_, o_1_, o_2_);

input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, i_18_, i_19_, i_20_, i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_, i_30_, i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_;

output o_0_, o_1_, o_2_;

wire n1, n2, n3, n5, n8, n10, n11, n9, n15, n13, n19, n17, n24, n23, n22, n26, n30, n31, n29, n33, n32, n35, n38, n39, n40, n36, n44, n41, n48, n45, n52, n50, n49, n56, n53, n60, n59, n57, n64, n63, n61, n67, n66, n65, n69, n70, n68, n72, n73, n74, n71, n75, n78, n81, n82, n84, n80, n87, n88, n86, n85, n90, n91, n89, n93, n94, n92, n96, n97, n98, n95, n100, n101, n99, n104, n102, n107, n105, n112, n110, n111, n109, n113, n121, n117, n125, n126, n124, n122, n129, n130, n131, n127, n133, n134, n135, n132, n139, n138, n136, n140, n144, n145, n143, n147, n148, n146, n150, n151, n149, n152, n155, n159, n160, n157, n162, n163, n161, n167, n165, n166, n164, n170, n168, n171, n175, n176, n174, n173, n180, n179, n177, n183, n184, n182, n181, n185, n188, n189, n190, n186, n193, n192, n191, n197, n195, n196, n194, n199, n200, n198, n203, n204, n201, n206, n205, n211, n207, n213, n215, n216, n212, n219, n217, n222, n221, n224, n225, n227, n229, n226, n232, n230, n236, n234, n233, n239, n238, n237, n241, n240, n243, n242, n246, n245, n244, n248, n249, n247, n250, n253, n252, n256, n255, n258, n261, n260, n263, n266, n265, n264, n268, n267, n269, n272, n273, n274, n282, n279, n278, n283, n284, n288, n287, n290, n289, n293, n299, n296, n300, n304, n301, n308, n307, n306, n305, n313, n311, n309, n315, n314, n317, n319, n322, n320, n324, n323, n326, n325, n328, n331, n335, n336, n334, n332, n337, n341, n340, n339, n342, n345, n346, n347, n344, n349, n350, n348, n352, n356, n355, n358, n362, n363, n364, n361, n367, n365, n368, n371, n372, n373, n374, n370, n376, n375, n377, n378, n382, n385, n394, n390, n395, n397, n402, n399, n404, n403, n407, n406, n408, n413, n414, n412, n415, n418, n421, n425, n429, n428, n436, n437, n438, n439, n440, n441, n433, n443, n444, n446, n442, n449, n448, n447, n451, n450, n455, n453, n454, n452, n459, n457, n458, n456, n462, n461, n460, n467, n463, n471, n469, n470, n468, n474, n473, n479, n477, n482, n481, n480, n485, n483, n487, n488, n489, n490, n486, n494, n495, n491, n497, n498, n496, n501, n500, n503, n505, n502, n506, n512, n513, n511, n516, n515, n514, n519, n518, n517, n520, n522, n521, n524, n523, n526, n527, n528, n525, n531, n529, n534, n533, n539, n535, n543, n540, n545, n544, n547, n548, n546, n550, n549, n554, n552, n556, n557, n558, n559, n555, n562, n561, n560, n563, n569, n567, n573, n572, n570, n576, n575, n574, n578, n579, n577, n580, n583, n584, n582, n586, n587, n585, n590, n588, n591, n595, n594, n596, n601, n607, n608, n609, n605, n611, n612, n610, n614, n615, n613, n617, n616, n619, n620, n618, n623, n622, n621, n626, n624, n628, n629, n627, n631, n630, n632, n633, n634, n639, n640, n638, n641, n644, n643, n642, n646, n645, n648, n649, n647, n651, n650, n653, n654, n652, n657, n655, n660, n661, n659, n658, n664, n662, n665, n670, n668, n669, n667, n672, n673, n671, n676, n674, n677, n680, n681, n682, n679, n684, n685, n683, n689, n688, n686, n692, n691, n695, n696, n694, n698, n699, n697, n700, n703, n704, n702, n705, n710, n709, n712, n714, n713, n718, n716, n717, n715, n720, n721, n719, n723, n724, n722, n725, n727, n728, n726, n729, n731, n734, n735, n733, n739, n737, n741, n740, n743, n744, n747, n746, n745, n749, n748, n750, n754, n755, n756, n757, n758, n759, n760, n761, n753, n763, n762, n764, n765, n767, n766, n769, n768, n771, n773, n777, n778, n776, n782, n781, n779, n784, n785, n783, n789, n787, n790, n792, n791, n794, n793, n795, n797, n798, n796, n801, n800, n799, n802, n806, n809, n810, n813, n812, n811, n814, n818, n821, n826, n824, n823, n829, n828, n827, n830, n832, n833, n831, n834, n837, n841, n840, n843, n845, n847, n849, n848, n851, n850, n853, n854, n852, n855, n856, n857, n859, n861, n866, n864, n868, n867, n870, n872, n871, n875, n874, n873, n880, n876, n882, n881, n884, n883, n886, n885, n888, n889, n887, n891, n890, n892, n893, n895, n894, n897, n896, n898, n899, n901, n904, n907, n906, n909, n908, n911, n910, n912, n916, n914, n915, n913, n917, n919, n918, n920, n922, n921, n926, n924, n927, n931, n929, n939, n942, n944, n947, n951, n950, n953, n954, n957, n960, n961, n962, n963, n964, n965, n966, n968, n969, n970, n972, n973, n974, n975, n977, n978, n979, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1033, n1035, n1036, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1050, n1049, n1051, n1053, n1055, n1057, n1056, n1058, n1060, n1062, n1063, n1065, n1066, n1068, n1067, n1070, n1069, n1072, n1071, n1073, n1074, n1076, n1079, n1082, n1081, n1083, n1084, n1085, n1087, n1088, n1089, n1092, n1091, n1094, n1093, n1097, n1100, n1099, n1101, n1102, n1107, n1106, n1108, n1109, n1112, n1114, n1113, n1115, n1116, n1117, n1120, n1118, n1122, n1121, n1124, n1123, n1128, n1127, n1126, n1130, n1129, n1131, n1132, n1134, n1133, n1135, n1136, n1140, n1139, n1141, n1143, n1147, n1146, n1149, n1152, n1153, n1155, n1157, n1159, n1160, n1163, n1164, n1169, n1171, n1170, n1173, n1172, n1174, n1175, n1179, n1180, n1181, n1183, n1182, n1186, n1187, n1189, n1188, n1191, n1190, n1192, n1193, n1195, n1194, n1197, n1196, n1198, n1200, n1199, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1209, n1208, n1210, n1214, n1213, n1215, n1216, n1222, n1220, n1223, n1225, n1226, n1224, n1228, n1227, n1230, n1229, n1231, n1232, n1237, n1236, n1238, n1239, n1242, n1241, n1244, n1243, n1245, n1247, n1246, n1248, n1249, n1250, n1251, n1253, n1256, n1257, n1258, n1259, n1260, n1261, n1263, n1264, n1268, n1272, n1273, n1276, n1279, n1280, n1281;

assign o_0_ = ( n1 ) | ( n2 ) | ( n3 ) | ( n5 ) | ( n8 ) | ( (~ n1248) ) | ( (~ n1249) ) | ( (~ n1250) ) ;
 assign o_1_ = ( (~ n753) ) ;
 assign o_2_ = ( (~ n433) ) ;
 assign n1 = ( n245  &  (~ n479)  &  n880  &  (~ n1025) ) ;
 assign n2 = ( i_35_  &  n670  &  n669  &  (~ n874) ) ;
 assign n3 = ( (~ i_13_)  &  (~ n885)  &  (~ n1035) ) | ( (~ i_14_)  &  (~ n885)  &  (~ n1035) ) ;
 assign n5 = ( (~ n662)  &  (~ n1215) ) | ( (~ n216)  &  (~ n608)  &  (~ n662) ) ;
 assign n8 = ( (~ n217) ) | ( n939 ) | ( n942 ) | ( n944 ) | ( n947 ) | ( n950 ) | ( n1033 ) | ( (~ n1253) ) ;
 assign n10 = ( (~ i_27_)  &  (~ n163) ) ;
 assign n11 = ( (~ i_30_)  &  n350 ) ;
 assign n9 = ( i_36_  &  (~ n1213) ) | ( i_36_  &  n10  &  n11 ) ;
 assign n15 = ( (~ i_12_)  &  (~ i_13_) ) ;
 assign n13 = ( (~ i_7_)  &  n15 ) | ( (~ i_7_)  &  (~ n1030) ) ;
 assign n19 = ( (~ i_11_)  &  (~ i_19_) ) ;
 assign n17 = ( (~ i_24_)  &  (~ n60) ) | ( (~ i_24_)  &  n19  &  (~ n59) ) ;
 assign n24 = ( (~ i_13_)  &  i_18_  &  i_19_ ) ;
 assign n23 = ( (~ i_13_)  &  i_18_ ) ;
 assign n22 = ( (~ i_22_)  &  n24 ) | ( i_11_  &  (~ i_22_)  &  n23 ) ;
 assign n26 = ( (~ i_24_)  &  (~ n67) ) | ( (~ i_24_)  &  n19  &  (~ n66) ) ;
 assign n30 = ( i_17_  &  i_12_ ) ;
 assign n31 = ( i_14_  &  i_13_ ) ;
 assign n29 = ( i_22_  &  n30 ) | ( i_22_  &  n31 ) ;
 assign n33 = ( (~ i_10_)  &  (~ i_24_) ) ;
 assign n32 = ( n33  &  (~ n70) ) | ( i_13_  &  (~ i_24_)  &  (~ n70) ) ;
 assign n35 = ( (~ i_24_)  &  n30 ) | ( (~ i_24_)  &  n31 ) ;
 assign n38 = ( i_1_ ) | ( n966 ) | ( n769 ) ;
 assign n39 = ( (~ i_18_) ) | ( (~ n256) ) ;
 assign n40 = ( i_6_ ) | ( n97 ) ;
 assign n36 = ( n38  &  n39 ) | ( n38  &  n40 ) | ( n39  &  (~ n256) ) | ( n40  &  (~ n256) ) ;
 assign n44 = ( i_11_  &  (~ i_13_) ) ;
 assign n41 = ( n44  &  (~ n1000) ) | ( i_18_  &  n44  &  (~ n147) ) ;
 assign n48 = ( i_9_  &  n44 ) ;
 assign n45 = ( (~ n38)  &  n48 ) | ( i_18_  &  (~ n40)  &  n48 ) ;
 assign n52 = ( (~ n324) ) | ( (~ n394) ) | ( (~ n800) ) ;
 assign n50 = ( (~ n394) ) | ( n968 ) ;
 assign n49 = ( n52  &  n50 ) | ( n52  &  (~ n121) ) ;
 assign n56 = ( n90 ) | ( n135 ) | ( (~ n324) ) ;
 assign n53 = ( n56  &  (~ n121) ) | ( n56  &  (~ n290) ) | ( n56  &  (~ n402) ) ;
 assign n60 = ( i_9_ ) | ( i_18_ ) | ( n990 ) ;
 assign n59 = ( n371 ) | ( n84 ) ;
 assign n57 = ( (~ n19)  &  n60 ) | ( n60  &  n59 ) ;
 assign n64 = ( i_6_ ) | ( n964 ) | ( n97 ) ;
 assign n63 = ( n374 ) | ( n965 ) ;
 assign n61 = ( (~ i_9_)  &  n64 ) | ( n64  &  n63 ) ;
 assign n67 = ( i_18_ ) | ( n985 ) ;
 assign n66 = ( n371 ) | ( n81 ) ;
 assign n65 = ( (~ n19)  &  n67 ) | ( n67  &  n66 ) ;
 assign n69 = ( i_10_  &  (~ i_13_) ) ;
 assign n70 = ( i_9_ ) | ( n986 ) ;
 assign n68 = ( n69  &  i_32_ ) | ( n70  &  i_32_ ) | ( n69  &  n65 ) | ( n70  &  n65 ) ;
 assign n72 = ( (~ i_9_) ) | ( n965 ) | ( n977 ) ;
 assign n73 = ( (~ i_11_) ) | ( i_12_ ) ;
 assign n74 = ( (~ i_11_) ) | ( n964 ) ;
 assign n71 = ( n72  &  n38 ) | ( n73  &  n38 ) | ( n72  &  n74 ) | ( n73  &  n74 ) ;
 assign n75 = ( (~ n44)  &  (~ n48) ) | ( (~ n48)  &  n64 ) | ( (~ n44)  &  n63 ) | ( n64  &  n63 ) ;
 assign n78 = ( i_13_  &  (~ i_18_) ) | ( (~ i_18_)  &  n71 ) | ( i_13_  &  n75 ) | ( n71  &  n75 ) ;
 assign n81 = ( i_7_ ) | ( n989 ) ;
 assign n82 = ( i_32_ ) | ( (~ i_38_) ) ;
 assign n84 = ( i_8_ ) | ( n989 ) ;
 assign n80 = ( n81  &  n84 ) | ( n82  &  n84 ) | ( n81  &  (~ n299) ) | ( n82  &  (~ n299) ) ;
 assign n87 = ( n81 ) | ( n91 ) | ( (~ n322) ) ;
 assign n88 = ( n84 ) | ( n100 ) | ( (~ n402) ) ;
 assign n86 = ( i_25_ ) | ( n963 ) ;
 assign n85 = ( n87  &  n88  &  n80 ) | ( n87  &  n88  &  n86 ) ;
 assign n90 = ( i_32_ ) | ( (~ n394) ) ;
 assign n91 = ( i_32_ ) | ( n963 ) ;
 assign n89 = ( n86  &  n91 ) | ( n90  &  n91 ) | ( n86  &  (~ n402) ) | ( n90  &  (~ n402) ) ;
 assign n93 = ( n983 ) | ( n528 ) ;
 assign n94 = ( n371 ) | ( n991 ) ;
 assign n92 = ( i_18_  &  i_19_ ) | ( n93  &  i_19_ ) | ( i_18_  &  n94 ) | ( n93  &  n94 ) ;
 assign n96 = ( n374 ) | ( n595 ) ;
 assign n97 = ( i_12_ ) | ( n371 ) ;
 assign n98 = ( i_6_ ) | ( (~ n229) ) ;
 assign n95 = ( i_8_  &  n97 ) | ( n96  &  n97 ) | ( i_8_  &  n98 ) | ( n96  &  n98 ) ;
 assign n100 = ( i_31_ ) | ( n963 ) ;
 assign n101 = ( i_35_ ) | ( n970 ) ;
 assign n99 = ( n100 ) | ( n92 ) | ( n101 ) ;
 assign n104 = ( i_32_ ) | ( n92 ) | ( (~ n299) ) ;
 assign n102 = ( i_2_  &  n104 ) | ( n104  &  (~ n290) ) | ( n104  &  (~ n394) ) ;
 assign n107 = ( (~ n86) ) | ( (~ n1258) ) ;
 assign n105 = ( i_38_  &  (~ n99) ) | ( i_38_  &  (~ n95)  &  n107 ) ;
 assign n112 = ( (~ n800)  &  n1117 ) | ( n1001  &  n1117 ) ;
 assign n110 = ( (~ i_38_)  &  n57 ) | ( n57  &  n68 ) | ( (~ i_38_)  &  (~ n299) ) | ( n68  &  (~ n299) ) ;
 assign n111 = ( i_10_  &  n1116 ) | ( n61  &  n1116 ) | ( (~ n394)  &  n1116 ) ;
 assign n109 = ( n112  &  i_28_ ) | ( n112  &  n110  &  n111 ) ;
 assign n113 = ( (~ i_24_)  &  (~ n1118) ) | ( (~ i_24_)  &  (~ n1121) ) | ( (~ i_24_)  &  (~ n1123) ) ;
 assign n121 = ( (~ i_28_)  &  (~ n163) ) ;
 assign n117 = ( n121  &  (~ n1126) ) | ( n121  &  (~ n1129) ) | ( n121  &  (~ n1132) ) ;
 assign n125 = ( i_30_ ) | ( n162 ) | ( (~ n313) ) ;
 assign n126 = ( n86  &  n195 ) | ( n86  &  (~ n306) ) | ( n195  &  n994 ) | ( (~ n306)  &  n994 ) ;
 assign n124 = ( (~ i_38_) ) | ( n988 ) ;
 assign n122 = ( (~ n11)  &  n125  &  n126 ) | ( n125  &  n126  &  n124 ) ;
 assign n129 = ( i_28_ ) | ( n179 ) ;
 assign n130 = ( i_22_ ) | ( (~ n288) ) ;
 assign n131 = ( n138 ) | ( (~ n394) ) ;
 assign n127 = ( n129  &  n130 ) | ( n129  &  n131 ) | ( n130  &  (~ n306) ) | ( n131  &  (~ n306) ) ;
 assign n133 = ( n130 ) | ( n138 ) ;
 assign n134 = ( n179 ) | ( (~ n402) ) ;
 assign n135 = ( i_31_ ) | ( i_30_ ) | ( i_28_ ) ;
 assign n132 = ( n133  &  n134 ) | ( n133  &  n135 ) | ( n134  &  (~ n299) ) | ( n135  &  (~ n299) ) ;
 assign n139 = ( i_30_ ) | ( (~ i_38_) ) | ( n86 ) ;
 assign n138 = ( i_30_ ) | ( n963 ) ;
 assign n136 = ( n139  &  n138 ) | ( n139  &  (~ n322) ) ;
 assign n140 = ( (~ n33)  &  n63 ) | ( n64  &  n63 ) | ( (~ n33)  &  (~ n311) ) | ( n64  &  (~ n311) ) ;
 assign n144 = ( (~ i_18_) ) | ( (~ n288) ) ;
 assign n145 = ( i_13_ ) | ( (~ n288) ) ;
 assign n143 = ( n75  &  n71 ) | ( n144  &  n71 ) | ( n75  &  n145 ) | ( n144  &  n145 ) ;
 assign n147 = ( n962 ) | ( n374 ) ;
 assign n148 = ( i_6_ ) | ( (~ i_9_) ) | ( i_10_ ) ;
 assign n146 = ( i_10_  &  n97 ) | ( n147  &  n97 ) | ( i_10_  &  n148 ) | ( n147  &  n148 ) ;
 assign n150 = ( i_8_ ) | ( i_30_ ) | ( (~ n299) ) ;
 assign n151 = ( n104  &  n69 ) | ( n104  &  n80 ) | ( n104  &  n371 ) ;
 assign n149 = ( n150  &  n151  &  n146 ) | ( n150  &  n151  &  n90 ) ;
 assign n152 = ( i_32_  &  (~ n32) ) | ( (~ n26)  &  (~ n32) ) ;
 assign n155 = ( i_30_  &  n152 ) | ( n152  &  (~ n414) ) ;
 assign n159 = ( (~ n17)  &  n155 ) | ( (~ n17)  &  (~ n322) ) | ( n155  &  n326 ) | ( (~ n322)  &  n326 ) ;
 assign n160 = ( n50  &  n1115 ) | ( (~ n311)  &  n1115 ) ;
 assign n157 = ( n149  &  n159  &  n160 ) | ( n159  &  n160  &  (~ n288) ) ;
 assign n162 = ( (~ i_34_) ) | ( (~ n394) ) ;
 assign n163 = ( i_24_ ) | ( i_26_ ) ;
 assign n161 = ( n162  &  n163 ) | ( n163  &  (~ n288) ) | ( n162  &  (~ n402) ) | ( (~ n288)  &  (~ n402) ) ;
 assign n167 = ( n81 ) | ( n163 ) | ( (~ n322) ) | ( (~ n367) ) ;
 assign n165 = ( n161 ) | ( n170 ) ;
 assign n166 = ( i_31_ ) | ( i_33_ ) | ( n162 ) | ( (~ n308) ) ;
 assign n164 = ( n167  &  n84 ) | ( n167  &  n165  &  n166 ) ;
 assign n170 = ( i_31_ ) | ( (~ n350) ) ;
 assign n168 = ( n100  &  n170 ) | ( n130  &  n170 ) | ( n100  &  (~ n324) ) | ( n130  &  (~ n324) ) ;
 assign n171 = ( (~ n121)  &  n162 ) | ( (~ n121)  &  (~ n304) ) | ( n162  &  (~ n402) ) | ( (~ n304)  &  (~ n402) ) ;
 assign n175 = ( n162 ) | ( (~ n308) ) | ( n972 ) ;
 assign n176 = ( n168  &  i_31_ ) | ( n90  &  i_31_ ) | ( n168  &  n206 ) | ( n90  &  n206 ) ;
 assign n174 = ( i_29_ ) | ( n685 ) ;
 assign n173 = ( n175  &  n176  &  n171 ) | ( n175  &  n176  &  n174 ) ;
 assign n180 = ( i_32_ ) | ( (~ i_38_) ) | ( n130 ) | ( n138 ) ;
 assign n179 = ( i_22_ ) | ( n163 ) ;
 assign n177 = ( n180  &  n179 ) | ( n180  &  (~ n322) ) | ( n180  &  (~ n800) ) ;
 assign n183 = ( n177 ) | ( n987 ) ;
 assign n184 = ( i_3_ ) | ( i_8_ ) | ( (~ i_10_) ) | ( n132 ) ;
 assign n182 = ( i_3_ ) | ( n964 ) ;
 assign n181 = ( n183  &  n184  &  n127 ) | ( n183  &  n184  &  n182 ) ;
 assign n185 = ( i_28_  &  i_29_ ) | ( i_28_  &  (~ n121) ) | ( i_29_  &  n179 ) | ( (~ n121)  &  n179 ) ;
 assign n188 = ( i_2_ ) | ( n964 ) ;
 assign n189 = ( (~ i_12_) ) | ( i_22_ ) | ( i_24_ ) ;
 assign n190 = ( i_10_ ) | ( n964 ) ;
 assign n186 = ( n188  &  n189 ) | ( n188  &  n190 ) | ( n189  &  (~ n429) ) | ( n190  &  (~ n429) ) ;
 assign n193 = ( i_26_ ) | ( (~ i_38_) ) | ( (~ n11) ) | ( n101 ) ;
 assign n192 = ( i_29_ ) | ( (~ n234) ) ;
 assign n191 = ( n193  &  i_28_ ) | ( n193  &  n192 ) | ( n193  &  n124 ) ;
 assign n197 = ( (~ i_38_) ) | ( (~ n11) ) | ( (~ n832) ) ;
 assign n195 = ( i_26_ ) | ( (~ n350) ) ;
 assign n196 = ( i_30_ ) | ( n90 ) ;
 assign n194 = ( n197  &  n195 ) | ( n197  &  n196 ) ;
 assign n199 = ( (~ i_19_) ) | ( i_24_ ) ;
 assign n200 = ( (~ i_19_) ) | ( (~ n288) ) ;
 assign n198 = ( n191  &  n194 ) | ( n199  &  n194 ) | ( n191  &  n200 ) | ( n199  &  n200 ) ;
 assign n203 = ( n91  &  (~ n304) ) | ( n130  &  (~ n304) ) | ( n91  &  n648 ) | ( n130  &  n648 ) ;
 assign n204 = ( (~ n121)  &  (~ n308) ) | ( n241  &  (~ n308) ) | ( (~ n121)  &  n376 ) | ( n241  &  n376 ) ;
 assign n201 = ( n203  &  n204  &  (~ n324) ) | ( n203  &  n204  &  (~ n367) ) ;
 assign n206 = ( i_32_ ) | ( i_28_ ) | ( n134 ) ;
 assign n205 = ( n201  &  n206 ) | ( n206  &  (~ n394) ) ;
 assign n211 = ( (~ i_31_) ) | ( (~ n253) ) ;
 assign n207 = ( n211  &  (~ n253) ) | ( (~ i_30_)  &  (~ i_32_)  &  n211 ) ;
 assign n213 = ( i_23_ ) | ( (~ n957) ) ;
 assign n215 = ( i_27_ ) | ( n960 ) ;
 assign n216 = ( (~ i_14_) ) | ( n734 ) ;
 assign n212 = ( n213  &  n215 ) | ( n213  &  n216 ) | ( n215  &  (~ n363) ) | ( n216  &  (~ n363) ) ;
 assign n219 = ( (~ i_20_) ) | ( (~ n681) ) | ( n874 ) | ( n954 ) ;
 assign n217 = ( n212  &  n219 ) | ( n219  &  (~ n253) ) | ( n219  &  (~ n673) ) ;
 assign n222 = ( i_22_ ) | ( (~ n256) ) ;
 assign n221 = ( i_3_  &  (~ n22) ) | ( (~ n22)  &  n222 ) ;
 assign n224 = ( i_7_  &  i_8_ ) | ( n177  &  i_8_ ) | ( i_7_  &  n132 ) | ( n177  &  n132 ) ;
 assign n225 = ( n224  &  n53 ) | ( n39  &  n53 ) | ( n224  &  n221 ) | ( n39  &  n221 ) ;
 assign n227 = ( (~ i_22_)  &  (~ n199) ) ;
 assign n229 = ( (~ i_7_)  &  (~ i_8_) ) ;
 assign n226 = ( (~ n136)  &  n227  &  n229 ) ;
 assign n232 = ( i_12_  &  n23 ) ;
 assign n230 = ( n226  &  n232 ) | ( i_11_  &  (~ n224)  &  n232 ) ;
 assign n236 = ( (~ i_34_) ) | ( n995 ) ;
 assign n234 = ( (~ i_30_)  &  (~ i_32_) ) ;
 assign n233 = ( i_28_  &  n236 ) | ( (~ i_34_)  &  n236 ) | ( n236  &  n234 ) ;
 assign n239 = ( (~ i_22_)  &  n234 ) | ( n234  &  n233 ) | ( (~ i_22_)  &  (~ n356) ) | ( n233  &  (~ n356) ) ;
 assign n238 = ( i_29_ ) | ( n724 ) ;
 assign n237 = ( n239  &  i_28_ ) | ( n239  &  n238 ) ;
 assign n241 = ( i_29_ ) | ( n970 ) ;
 assign n240 = ( i_25_  &  i_28_ ) | ( i_25_  &  n241 ) | ( i_28_  &  (~ n367) ) | ( n241  &  (~ n367) ) ;
 assign n243 = ( i_31_ ) | ( n974 ) ;
 assign n242 = ( n92  &  i_8_ ) | ( n174  &  i_8_ ) | ( n92  &  n243 ) | ( n174  &  n243 ) ;
 assign n246 = ( i_33_  &  n253 ) ;
 assign n245 = ( i_33_  &  i_34_ ) ;
 assign n244 = ( i_14_  &  n246 ) | ( i_14_  &  (~ i_24_)  &  n245 ) ;
 assign n248 = ( n1012  &  n96 ) ;
 assign n249 = ( i_2_ ) | ( (~ n229) ) ;
 assign n247 = ( i_32_  &  i_30_ ) | ( n248  &  i_30_ ) | ( i_32_  &  n249 ) | ( n248  &  n249 ) ;
 assign n250 = ( i_22_  &  n244 ) | ( i_22_  &  (~ n207)  &  n213 ) ;
 assign n253 = ( (~ i_34_)  &  i_35_ ) ;
 assign n252 = ( (~ n290)  &  (~ n1097) ) | ( n29  &  n253  &  (~ n290) ) ;
 assign n256 = ( (~ i_13_)  &  i_19_ ) ;
 assign n255 = ( n44  &  (~ n182) ) | ( (~ n182)  &  n256 ) ;
 assign n258 = ( (~ i_24_)  &  n255 ) | ( (~ i_24_)  &  n23  &  (~ n74) ) ;
 assign n261 = ( i_13_ ) | ( n964 ) ;
 assign n260 = ( (~ i_18_)  &  (~ n258) ) | ( n199  &  (~ n258) ) | ( (~ n258)  &  n261 ) ;
 assign n263 = ( (~ i_18_)  &  n39 ) | ( n39  &  (~ n44) ) ;
 assign n266 = ( n74  &  n188 ) | ( n188  &  (~ n232) ) | ( n74  &  n263 ) | ( (~ n232)  &  n263 ) ;
 assign n265 = ( (~ i_12_) ) | ( n964 ) ;
 assign n264 = ( n266  &  n39 ) | ( n266  &  n265 ) ;
 assign n268 = ( i_12_  &  n44 ) ;
 assign n267 = ( i_18_  &  (~ i_22_)  &  n268 ) ;
 assign n269 = ( (~ i_8_)  &  i_12_  &  (~ i_13_)  &  n227  &  (~ n987) ) ;
 assign n272 = ( n90  &  n134 ) | ( n133  &  n134 ) | ( n90  &  (~ n800) ) | ( n133  &  (~ n800) ) ;
 assign n273 = ( i_7_  &  n49 ) | ( n177  &  n49 ) | ( i_7_  &  n221 ) | ( n177  &  n221 ) ;
 assign n274 = ( (~ i_2_)  &  (~ i_10_)  &  (~ n272) ) | ( (~ i_10_)  &  i_12_  &  (~ n272) ) ;
 assign n282 = ( (~ i_3_)  &  i_11_ ) ;
 assign n279 = ( i_12_  &  (~ i_13_)  &  (~ i_22_) ) ;
 assign n278 = ( n282  &  (~ n1088) ) | ( (~ n49)  &  n282  &  n279 ) ;
 assign n283 = ( i_8_  &  (~ n19) ) | ( (~ n19)  &  n67 ) | ( i_8_  &  n70 ) | ( n67  &  n70 ) ;
 assign n284 = ( (~ i_24_)  &  (~ n66)  &  (~ n69)  &  (~ n240) ) ;
 assign n288 = ( (~ i_24_)  &  (~ i_25_) ) ;
 assign n287 = ( (~ i_7_)  &  (~ i_32_)  &  n11  &  n288 ) ;
 assign n290 = ( (~ i_31_)  &  n234 ) ;
 assign n289 = ( (~ i_22_)  &  (~ n29) ) | ( (~ i_23_)  &  (~ n29) ) | ( (~ i_22_)  &  n290 ) | ( (~ i_23_)  &  n290 ) ;
 assign n293 = ( (~ i_38_)  &  (~ n17) ) | ( (~ n17)  &  n152 ) | ( (~ i_38_)  &  (~ n299) ) | ( n152  &  (~ n299) ) ;
 assign n299 = ( (~ i_31_)  &  n394 ) ;
 assign n296 = ( (~ i_29_)  &  n299  &  (~ n1057) ) ;
 assign n300 = ( i_8_ ) | ( (~ n11) ) | ( (~ n288) ) | ( (~ n299) ) ;
 assign n304 = ( (~ i_28_)  &  n288 ) ;
 assign n301 = ( n296  &  n304 ) | ( (~ n190)  &  n304  &  (~ n994) ) ;
 assign n308 = ( (~ i_24_)  &  n350 ) ;
 assign n307 = ( (~ i_31_)  &  n402  &  (~ n1057) ) ;
 assign n306 = ( (~ i_30_)  &  n402 ) ;
 assign n305 = ( n308  &  n307 ) | ( (~ n190)  &  n308  &  n306 ) ;
 assign n313 = ( (~ i_25_)  &  n350 ) ;
 assign n311 = ( n33  &  i_9_ ) ;
 assign n309 = ( (~ n293)  &  n313 ) | ( (~ n196)  &  n313  &  n311 ) ;
 assign n315 = ( i_29_ ) | ( n995 ) ;
 assign n314 = ( (~ n35) ) | ( n315 ) ;
 assign n317 = ( i_38_  &  n284 ) | ( i_38_  &  n287 ) | ( i_38_  &  (~ n1081) ) ;
 assign n319 = ( n86  &  n139 ) | ( n139  &  n293 ) | ( n86  &  (~ n414) ) | ( n293  &  (~ n414) ) ;
 assign n322 = ( (~ i_33_)  &  i_38_ ) ;
 assign n320 = ( (~ i_7_)  &  (~ n163)  &  n322 ) ;
 assign n324 = ( (~ i_25_)  &  (~ n163) ) ;
 assign n323 = ( (~ i_32_)  &  n320 ) | ( (~ i_32_)  &  n299  &  n324 ) ;
 assign n326 = ( i_33_ ) | ( (~ n299) ) ;
 assign n325 = ( i_8_  &  (~ n323) ) | ( n163  &  (~ n323) ) | ( (~ n323)  &  n326 ) ;
 assign n328 = ( (~ i_25_)  &  (~ n996) ) | ( (~ i_25_)  &  n11  &  n229 ) ;
 assign n331 = ( (~ n69)  &  (~ n70) ) | ( (~ i_32_)  &  (~ n66)  &  (~ n69) ) ;
 assign n335 = ( (~ n367)  &  n1065 ) | ( (~ n324)  &  (~ n349)  &  n1065 ) ;
 assign n336 = ( (~ n308)  &  n1066 ) | ( n376  &  n1066 ) ;
 assign n334 = ( i_32_ ) | ( (~ n253) ) ;
 assign n332 = ( (~ n313)  &  n335  &  n336 ) | ( n335  &  n336  &  n334 ) ;
 assign n337 = ( (~ n95)  &  (~ n195) ) | ( (~ i_7_)  &  (~ n195)  &  n234 ) ;
 assign n341 = ( n66 ) | ( (~ n350) ) | ( n716 ) ;
 assign n340 = ( i_34_ ) | ( i_33_ ) | ( i_29_ ) ;
 assign n339 = ( n341  &  i_28_ ) | ( n341  &  n70 ) | ( n341  &  n340 ) ;
 assign n342 = ( n101  &  (~ n304) ) | ( (~ n121)  &  (~ n304) ) | ( n101  &  (~ n832) ) | ( (~ n121)  &  (~ n832) ) ;
 assign n345 = ( i_33_ ) | ( n978 ) ;
 assign n346 = ( i_24_ ) | ( i_28_ ) ;
 assign n347 = ( i_33_ ) | ( (~ n350) ) ;
 assign n344 = ( n345  &  n163 ) | ( n346  &  n163 ) | ( n345  &  n347 ) | ( n346  &  n347 ) ;
 assign n349 = ( (~ i_33_)  &  n253 ) ;
 assign n350 = ( (~ i_28_)  &  (~ i_29_) ) ;
 assign n348 = ( (~ n95)  &  (~ n344) ) | ( (~ n95)  &  n349  &  n350 ) ;
 assign n352 = ( (~ n283)  &  (~ n1062) ) | ( (~ n283)  &  n324  &  n350 ) ;
 assign n356 = ( n350  &  i_34_ ) ;
 assign n355 = ( n288  &  (~ n1063) ) | ( (~ n95)  &  n288  &  n356 ) ;
 assign n358 = ( n253  &  n328 ) | ( n253  &  (~ n1067) ) | ( n253  &  (~ n1069) ) ;
 assign n362 = ( (~ i_27_)  &  n350 ) ;
 assign n363 = ( n15  &  i_14_ ) ;
 assign n364 = ( (~ i_16_)  &  n833 ) ;
 assign n361 = ( n362  &  n363  &  n364 ) ;
 assign n367 = ( (~ i_32_)  &  n350 ) ;
 assign n365 = ( (~ n146)  &  (~ n163)  &  n367 ) ;
 assign n368 = ( (~ n17)  &  (~ n290) ) | ( n170  &  (~ n290) ) | ( (~ n17)  &  (~ n308) ) | ( n170  &  (~ n308) ) ;
 assign n371 = ( i_5_ ) | ( n961 ) ;
 assign n372 = ( i_12_ ) | ( i_6_ ) ;
 assign n373 = ( i_5_ ) | ( i_6_ ) ;
 assign n374 = ( i_1_ ) | ( n961 ) ;
 assign n370 = ( n371  &  n373 ) | ( n372  &  n373 ) | ( n371  &  n374 ) | ( n372  &  n374 ) ;
 assign n376 = ( (~ i_34_) ) | ( n970 ) ;
 assign n375 = ( n190  &  (~ n311) ) | ( (~ n311)  &  (~ n324) ) | ( n190  &  n376 ) | ( (~ n324)  &  n376 ) ;
 assign n377 = ( i_29_  &  n192 ) | ( n140  &  n192 ) | ( i_29_  &  (~ n311) ) | ( n140  &  (~ n311) ) ;
 assign n378 = ( (~ i_24_)  &  (~ n370)  &  (~ n1045) ) | ( (~ i_24_)  &  (~ n370)  &  (~ n1046) ) ;
 assign n382 = ( (~ n86)  &  n227 ) | ( n227  &  (~ n1258) ) ;
 assign n385 = ( (~ n1047)  &  (~ n1049) ) | ( (~ n1048)  &  (~ n1049) ) | ( (~ n1047)  &  (~ n1051) ) | ( (~ n1048)  &  (~ n1051) ) ;
 assign n394 = ( (~ i_35_)  &  i_38_ ) ;
 assign n390 = ( n394  &  (~ n1053) ) | ( n394  &  (~ n1055) ) | ( n394  &  (~ n1058) ) ;
 assign n395 = ( (~ n185)  &  n307 ) | ( (~ n185)  &  (~ n283)  &  n322 ) ;
 assign n397 = ( (~ n181)  &  n268 ) | ( i_12_  &  (~ n181)  &  n256 ) ;
 assign n402 = ( (~ i_33_)  &  n394 ) ;
 assign n399 = ( n365  &  n402 ) | ( (~ n138)  &  (~ n186)  &  n402 ) ;
 assign n404 = ( n362  &  (~ n608) ) ;
 assign n403 = ( n245  &  n361 ) | ( (~ n216)  &  n245  &  n404 ) ;
 assign n407 = ( n350  &  n290  &  n246 ) ;
 assign n406 = ( i_14_  &  n407 ) | ( i_14_  &  n121  &  i_33_ ) ;
 assign n408 = ( i_9_  &  (~ n1089) ) | ( i_9_  &  (~ n1091) ) | ( i_9_  &  (~ n1093) ) ;
 assign n413 = ( i_10_  &  n267 ) | ( i_10_  &  n282  &  n279 ) ;
 assign n414 = ( (~ i_24_)  &  n229 ) ;
 assign n412 = ( (~ n136)  &  n269 ) | ( (~ n136)  &  n413  &  n414 ) ;
 assign n415 = ( (~ i_28_)  &  n250 ) | ( (~ i_28_)  &  n252 ) | ( (~ i_28_)  &  (~ n1263) ) ;
 assign n418 = ( i_10_  &  (~ n1102) ) | ( i_10_  &  i_12_  &  (~ n225) ) ;
 assign n421 = ( n48  &  (~ n1106) ) | ( n48  &  (~ n127)  &  (~ n997) ) ;
 assign n425 = ( n213  &  (~ n1108) ) | ( n121  &  n213  &  (~ n234) ) ;
 assign n429 = ( (~ i_22_)  &  n33 ) ;
 assign n428 = ( (~ n371)  &  (~ n1113) ) | ( (~ n85)  &  (~ n371)  &  n429 ) ;
 assign n436 = ( (~ i_27_)  &  (~ n390) ) | ( n179  &  (~ n390) ) | ( (~ n390)  &  (~ n531) ) ;
 assign n437 = ( n1141  &  n49 ) | ( n1141  &  n222 ) | ( n1141  &  n969 ) ;
 assign n438 = ( (~ n35)  &  n1139 ) | ( n234  &  n1139 ) | ( (~ n356)  &  n1139 ) ;
 assign n439 = ( (~ n11)  &  (~ n406)  &  n1146 ) | ( n325  &  (~ n406)  &  n1146 ) ;
 assign n440 = ( n124  &  (~ n399)  &  n1143 ) | ( n368  &  (~ n399)  &  n1143 ) ;
 assign n441 = ( (~ n418)  &  (~ n421)  &  n1149  &  n1152  &  n1153  &  n1157  &  n1159  &  n1160 ) ;
 assign n433 = ( (~ n395)  &  (~ n397)  &  n436  &  n437  &  n438  &  n439  &  n440  &  n441 ) ;
 assign n443 = ( (~ i_34_) ) | ( (~ i_37_) ) ;
 assign n444 = ( i_29_ ) | ( n649 ) ;
 assign n446 = ( (~ i_37_) ) | ( (~ n253) ) ;
 assign n442 = ( (~ n362)  &  n443 ) | ( (~ n362)  &  n444 ) | ( n443  &  n446 ) | ( n444  &  n446 ) ;
 assign n449 = ( i_29_ ) | ( (~ n543) ) | ( n664 ) ;
 assign n448 = ( (~ i_34_) ) | ( (~ n543) ) ;
 assign n447 = ( (~ n362)  &  n449 ) | ( n449  &  n448 ) ;
 assign n451 = ( (~ i_37_) ) | ( (~ n362) ) | ( (~ n832) ) ;
 assign n450 = ( n451  &  i_32_ ) | ( n451  &  n449 ) ;
 assign n455 = ( n371 ) | ( n453 ) | ( n1020 ) ;
 assign n453 = ( i_17_ ) | ( n735 ) ;
 assign n454 = ( i_10_ ) | ( n989 ) ;
 assign n452 = ( n455  &  n371 ) | ( n455  &  n453 ) | ( n455  &  n454 ) ;
 assign n459 = ( n1015 ) | ( n454 ) | ( n522 ) | ( n501 ) ;
 assign n457 = ( (~ i_37_) ) | ( n595 ) | ( n622 ) ;
 assign n458 = ( (~ n543) ) | ( n1015 ) | ( n1114 ) ;
 assign n456 = ( n459  &  n453 ) | ( n459  &  n457  &  n458 ) ;
 assign n462 = ( (~ n494) ) | ( n992 ) | ( n1015 ) ;
 assign n461 = ( i_7_ ) | ( i_0_ ) | ( n1005 ) ;
 assign n460 = ( n462  &  i_12_ ) | ( n462  &  n461 ) ;
 assign n467 = ( (~ i_23_)  &  (~ n163) ) ;
 assign n463 = ( n467  &  (~ n1194) ) | ( (~ n460)  &  n467  &  (~ n629) ) ;
 assign n471 = ( n639 ) | ( n1009 ) | ( n587 ) ;
 assign n469 = ( i_11_ ) | ( n735 ) ;
 assign n470 = ( n81 ) | ( n1015 ) | ( n746 ) ;
 assign n468 = ( (~ n463)  &  n471  &  n469 ) | ( (~ n463)  &  n471  &  n470 ) ;
 assign n474 = ( i_14_ ) | ( (~ n543) ) ;
 assign n473 = ( (~ i_21_)  &  (~ n11) ) | ( (~ i_21_)  &  n474 ) | ( (~ n11)  &  (~ n692) ) | ( n474  &  (~ n692) ) ;
 assign n479 = ( n953  &  n453 ) ;
 assign n477 = ( i_33_  &  n479 ) | ( n479  &  (~ n688) ) ;
 assign n482 = ( n66 ) | ( n763 ) ;
 assign n481 = ( i_10_ ) | ( n735 ) ;
 assign n480 = ( n482  &  n66 ) | ( n482  &  n481 ) ;
 assign n485 = ( (~ i_31_) ) | ( (~ n11) ) | ( n477 ) | ( n572 ) ;
 assign n483 = ( (~ n404)  &  n485 ) | ( n480  &  n485 ) ;
 assign n487 = ( (~ i_29_) ) | ( n456 ) | ( n664 ) | ( n1027 ) ;
 assign n488 = ( n884 ) | ( n561 ) | ( n1023 ) | ( i_29_ ) ;
 assign n489 = ( (~ i_37_)  &  n443 ) | ( n443  &  n468 ) | ( (~ i_37_)  &  n483 ) | ( n468  &  n483 ) ;
 assign n490 = ( n1196  &  i_31_ ) | ( n1196  &  n473 ) | ( n1196  &  n684 ) ;
 assign n486 = ( n487  &  n488  &  n489  &  n490 ) ;
 assign n494 = ( (~ i_27_)  &  n531 ) ;
 assign n495 = ( n833  &  i_22_ ) ;
 assign n491 = ( (~ n479)  &  n494  &  n495 ) | ( n494  &  n495  &  (~ n1011) ) ;
 assign n497 = ( (~ i_33_) ) | ( n685 ) ;
 assign n498 = ( (~ i_25_) ) | ( (~ n833) ) ;
 assign n496 = ( (~ n11)  &  (~ n491) ) | ( (~ n491)  &  n497 ) | ( (~ n491)  &  n498 ) ;
 assign n501 = ( i_33_ ) | ( (~ n543) ) ;
 assign n500 = ( n474  &  i_13_ ) | ( n474  &  n501 ) ;
 assign n503 = ( n481  &  n763 ) ;
 assign n505 = ( i_10_ ) | ( n734 ) ;
 assign n502 = ( n501  &  n503 ) | ( n503  &  n505 ) | ( n501  &  (~ n543) ) | ( n505  &  (~ n543) ) ;
 assign n506 = ( (~ n457)  &  (~ n620) ) | ( (~ i_33_)  &  (~ n457)  &  (~ n609) ) ;
 assign n512 = ( i_20_ ) | ( (~ n1003) ) ;
 assign n513 = ( i_20_ ) | ( n960 ) ;
 assign n511 = ( i_12_  &  i_16_ ) | ( n512  &  i_16_ ) | ( i_12_  &  n513 ) | ( n512  &  n513 ) ;
 assign n516 = ( n1169  &  n990 ) | ( n1169  &  n639 ) | ( n1169  &  n1013 ) ;
 assign n515 = ( i_19_ ) | ( n960 ) ;
 assign n514 = ( n516  &  n59 ) | ( n516  &  n515 ) | ( n516  &  n469 ) ;
 assign n519 = ( n990 ) | ( n640 ) | ( n1013 ) ;
 assign n518 = ( i_11_ ) | ( n734 ) ;
 assign n517 = ( n519  &  n59 ) | ( n519  &  n515 ) | ( n519  &  n518 ) ;
 assign n520 = ( n503  &  i_33_ ) | ( n503  &  n505 ) ;
 assign n522 = ( i_17_ ) | ( n734 ) ;
 assign n521 = ( n453  &  n501 ) | ( n453  &  n522 ) | ( n501  &  (~ n543) ) | ( n522  &  (~ n543) ) ;
 assign n524 = ( n1192  &  i_19_ ) | ( n1192  &  n991 ) | ( n1192  &  n526 ) ;
 assign n523 = ( n524  &  n500 ) | ( n524  &  n372 ) | ( n524  &  n512 ) ;
 assign n526 = ( i_23_ ) | ( i_20_ ) | ( n521 ) ;
 assign n527 = ( (~ i_3_) ) | ( n1007 ) ;
 assign n528 = ( i_9_ ) | ( n373 ) ;
 assign n525 = ( n526 ) | ( n527 ) | ( n528 ) | ( i_18_ ) ;
 assign n531 = ( (~ i_28_)  &  i_29_ ) ;
 assign n529 = ( n506  &  (~ n513)  &  n531 ) | ( (~ n513)  &  n531  &  (~ n1190) ) ;
 assign n534 = ( i_13_ ) | ( n1014 ) | ( n556 ) ;
 assign n533 = ( (~ n367) ) | ( n501 ) | ( n534 ) ;
 assign n539 = ( (~ i_32_)  &  n531 ) ;
 assign n535 = ( (~ n525)  &  n539 ) | ( (~ n523)  &  n539  &  (~ n1015) ) ;
 assign n543 = ( (~ i_35_)  &  i_37_ ) ;
 assign n540 = ( n543  &  (~ n1193) ) | ( n367  &  n543  &  (~ n704) ) ;
 assign n545 = ( n1163  &  n984 ) | ( n1163  &  n640 ) | ( n1163  &  n1013 ) ;
 assign n544 = ( n545  &  n66 ) | ( n545  &  n515 ) | ( n545  &  n518 ) ;
 assign n547 = ( i_18_ ) | ( (~ n833) ) ;
 assign n548 = ( i_19_ ) | ( (~ n833) ) ;
 assign n546 = ( n93  &  n94 ) | ( n547  &  n94 ) | ( n93  &  n548 ) | ( n547  &  n548 ) ;
 assign n550 = ( (~ i_37_) ) | ( n970 ) ;
 assign n549 = ( i_30_ ) | ( (~ i_31_) ) | ( n550 ) | ( (~ n688) ) ;
 assign n554 = ( n371 ) | ( n522 ) | ( n454 ) ;
 assign n552 = ( (~ i_37_) ) | ( n101 ) | ( n554 ) ;
 assign n556 = ( i_16_ ) | ( n960 ) ;
 assign n557 = ( i_13_ ) | ( (~ n229) ) ;
 assign n558 = ( i_23_ ) | ( n734 ) ;
 assign n559 = ( i_12_ ) | ( (~ n229) ) ;
 assign n555 = ( n556  &  n558 ) | ( n557  &  n558 ) | ( n556  &  n559 ) | ( n557  &  n559 ) ;
 assign n562 = ( (~ i_34_) ) | ( (~ n364) ) | ( n501 ) | ( n607 ) ;
 assign n561 = ( i_34_ ) | ( n717 ) ;
 assign n560 = ( n562  &  i_33_ ) | ( n562  &  n555 ) | ( n562  &  n561 ) ;
 assign n563 = ( n467  &  (~ n549) ) | ( n467  &  (~ n552) ) | ( n467  &  (~ n1187) ) ;
 assign n569 = ( n1188  &  n544 ) | ( n1188  &  n716 ) | ( n1188  &  n717 ) ;
 assign n567 = ( i_30_  &  (~ n563)  &  n569 ) | ( n560  &  (~ n563)  &  n569 ) ;
 assign n573 = ( (~ n841) ) | ( n884 ) ;
 assign n572 = ( i_27_ ) | ( (~ n833) ) ;
 assign n570 = ( (~ n356)  &  n573 ) | ( n573  &  n572 ) ;
 assign n576 = ( i_8_ ) | ( n985 ) | ( n586 ) ;
 assign n575 = ( i_11_ ) | ( n1010 ) ;
 assign n574 = ( n576  &  n70 ) | ( n576  &  n575 ) ;
 assign n578 = ( n243 ) | ( n334 ) | ( i_7_ ) | ( i_28_ ) ;
 assign n579 = ( i_9_ ) | ( n69 ) | ( n631 ) | ( (~ n681) ) | ( n1016 ) ;
 assign n577 = ( n578  &  n579  &  n570 ) | ( n578  &  n579  &  n574 ) ;
 assign n580 = ( i_10_  &  i_30_ ) | ( i_30_  &  n70 ) | ( i_10_  &  (~ n229) ) | ( n70  &  (~ n229) ) ;
 assign n583 = ( n442 ) | ( n580 ) | ( n556 ) ;
 assign n584 = ( (~ n543)  &  n1186 ) | ( n973  &  n1186 ) | ( n993  &  n1186 ) ;
 assign n582 = ( (~ i_37_)  &  n583  &  n584 ) | ( n577  &  n583  &  n584 ) ;
 assign n586 = ( i_18_ ) | ( n1006 ) ;
 assign n587 = ( n595 ) | ( n527 ) ;
 assign n585 = ( n586 ) | ( i_8_ ) | ( n587 ) ;
 assign n590 = ( (~ i_9_)  &  (~ n585) ) | ( (~ i_9_)  &  (~ n575)  &  (~ n1016) ) ;
 assign n588 = ( (~ i_14_)  &  n590 ) | ( (~ i_13_)  &  (~ i_33_)  &  n590 ) ;
 assign n591 = ( (~ n953)  &  (~ n1016) ) | ( (~ i_33_)  &  (~ n1011)  &  (~ n1016) ) ;
 assign n595 = ( i_7_ ) | ( n373 ) ;
 assign n594 = ( n522 ) | ( n595 ) | ( n550 ) ;
 assign n596 = ( (~ n594)  &  (~ n622) ) | ( (~ n521)  &  (~ n622)  &  (~ n965) ) ;
 assign n601 = ( (~ i_37_)  &  (~ n596) ) | ( (~ n588)  &  (~ n591)  &  (~ n596) ) ;
 assign n607 = ( i_8_ ) | ( (~ n15) ) ;
 assign n608 = ( i_17_ ) | ( (~ n833) ) ;
 assign n609 = ( i_8_ ) | ( n734 ) ;
 assign n605 = ( (~ n364)  &  n608 ) | ( n607  &  n608 ) | ( (~ n364)  &  n609 ) | ( n607  &  n609 ) ;
 assign n611 = ( i_33_ ) | ( n974 ) ;
 assign n612 = ( n789  &  n1259 ) ;
 assign n610 = ( n605  &  n612 ) | ( n611  &  n612 ) | ( n605  &  n241 ) | ( n611  &  n241 ) ;
 assign n614 = ( (~ n689) ) | ( n953 ) ;
 assign n615 = ( (~ i_29_)  &  n1256 ) | ( n601  &  n1256 ) | ( n1027  &  n1256 ) ;
 assign n613 = ( (~ n543)  &  n614  &  n615 ) | ( n610  &  n614  &  n615 ) ;
 assign n617 = ( (~ i_25_) ) | ( i_28_ ) | ( n497 ) | ( n1026 ) ;
 assign n616 = ( (~ n404)  &  n617 ) | ( n501  &  n617 ) | ( n609  &  n617 ) ;
 assign n619 = ( i_8_ ) | ( n1030 ) ;
 assign n620 = ( i_8_ ) | ( n735 ) ;
 assign n618 = ( (~ n364)  &  n608 ) | ( n608  &  n619 ) | ( (~ n364)  &  n620 ) | ( n619  &  n620 ) ;
 assign n623 = ( i_10_ ) | ( n1016 ) | ( i_33_ ) | ( i_9_ ) ;
 assign n622 = ( i_1_ ) | ( n1007 ) ;
 assign n621 = ( n623  &  n373 ) | ( n623  &  n101 ) | ( n623  &  n622 ) ;
 assign n626 = ( n461 ) | ( (~ n467) ) | ( n550 ) ;
 assign n624 = ( (~ i_37_)  &  n626 ) | ( n621  &  n626 ) | ( n626  &  (~ n681) ) ;
 assign n628 = ( i_20_ ) | ( n734 ) ;
 assign n629 = ( i_20_ ) | ( n735 ) ;
 assign n627 = ( n501  &  (~ n543) ) | ( (~ n543)  &  n628 ) | ( n501  &  n629 ) | ( n628  &  n629 ) ;
 assign n631 = ( i_20_ ) | ( n1006 ) ;
 assign n630 = ( i_12_  &  n500 ) | ( n627  &  n500 ) | ( i_12_  &  n631 ) | ( n627  &  n631 ) ;
 assign n632 = ( (~ i_7_)  &  i_37_  &  n349 ) ;
 assign n633 = ( n350  &  n632 ) | ( n350  &  i_25_  &  n246 ) ;
 assign n634 = ( (~ n253)  &  (~ n633) ) | ( (~ n531)  &  (~ n633) ) | ( (~ n633)  &  (~ n954) ) ;
 assign n639 = ( i_9_ ) | ( n735 ) ;
 assign n640 = ( i_9_ ) | ( n734 ) ;
 assign n638 = ( n501  &  (~ n543) ) | ( n501  &  n639 ) | ( (~ n543)  &  n640 ) | ( n639  &  n640 ) ;
 assign n641 = ( n544  &  n448 ) | ( n443  &  n448 ) | ( n544  &  n534 ) | ( n443  &  n534 ) ;
 assign n644 = ( n986 ) | ( n1011 ) ;
 assign n643 = ( i_11_ ) | ( n70 ) | ( n1010 ) ;
 assign n642 = ( n644  &  i_13_ ) | ( n644  &  n643  &  n576 ) ;
 assign n646 = ( n63 ) | ( n522 ) ;
 assign n645 = ( n642  &  n448 ) | ( n443  &  n448 ) | ( n642  &  n646 ) | ( n443  &  n646 ) ;
 assign n648 = ( i_32_ ) | ( n978 ) ;
 assign n649 = ( i_24_ ) | ( n1004 ) ;
 assign n647 = ( n334  &  n648 ) | ( (~ n362)  &  n648 ) | ( n334  &  n649 ) | ( (~ n362)  &  n649 ) ;
 assign n651 = ( n1179  &  n984 ) | ( n1179  &  n639 ) | ( n1179  &  n1013 ) ;
 assign n650 = ( n651  &  n66 ) | ( n651  &  n515 ) | ( n651  &  n469 ) ;
 assign n653 = ( (~ n367) ) | ( n572 ) ;
 assign n654 = ( n59 ) | ( n505 ) ;
 assign n652 = ( (~ n404)  &  n554 ) | ( (~ n404)  &  n653 ) | ( n554  &  n654 ) | ( n653  &  n654 ) ;
 assign n657 = ( n215 ) | ( (~ n367) ) ;
 assign n655 = ( (~ n349)  &  n376 ) | ( (~ n349)  &  (~ n404) ) | ( n376  &  n657 ) | ( (~ n404)  &  n657 ) ;
 assign n660 = ( n652  &  n647 ) | ( n988  &  n647 ) | ( n652  &  n650 ) | ( n988  &  n650 ) ;
 assign n661 = ( n1180  &  n1181  &  n655 ) | ( n1180  &  n1181  &  n1029 ) ;
 assign n659 = ( n986 ) | ( n953 ) ;
 assign n658 = ( n660  &  n661  &  n570 ) | ( n660  &  n661  &  n659 ) ;
 assign n664 = ( i_26_ ) | ( n1004 ) ;
 assign n662 = ( (~ i_33_)  &  (~ n245) ) | ( (~ i_33_)  &  (~ n362) ) | ( (~ n245)  &  n664 ) | ( (~ n362)  &  n664 ) ;
 assign n665 = ( i_20_  &  (~ i_23_)  &  i_25_  &  (~ n849) ) ;
 assign n670 = ( (~ i_34_)  &  n531 ) ;
 assign n668 = ( (~ i_27_)  &  n891 ) ;
 assign n669 = ( i_22_  &  n1024 ) ;
 assign n667 = ( i_35_  &  n670  &  n668 ) | ( i_35_  &  n670  &  n669 ) ;
 assign n672 = ( i_25_  &  n1024 ) ;
 assign n673 = ( n350  &  i_33_ ) ;
 assign n671 = ( n253  &  n665 ) | ( n253  &  n672  &  n673 ) ;
 assign n676 = ( (~ i_34_)  &  n1175 ) | ( (~ n494)  &  n1175 ) | ( (~ n880)  &  n1175 ) ;
 assign n674 = ( n498  &  (~ n671)  &  n676 ) | ( n662  &  (~ n671)  &  n676 ) ;
 assign n677 = ( i_34_  &  n494  &  (~ n522) ) ;
 assign n680 = ( (~ i_20_)  &  (~ i_21_) ) ;
 assign n681 = ( n467  &  n494 ) ;
 assign n682 = ( (~ n953) ) | ( (~ n1011) ) ;
 assign n679 = ( n680  &  i_2_  &  n681  &  n682 ) ;
 assign n684 = ( i_34_ ) | ( n163 ) ;
 assign n685 = ( i_31_ ) | ( i_32_ ) ;
 assign n683 = ( (~ i_22_) ) | ( n684 ) | ( n685 ) | ( (~ n692) ) ;
 assign n689 = ( i_29_  &  n495 ) ;
 assign n688 = ( (~ n522) ) | ( (~ n1011) ) ;
 assign n686 = ( (~ n453)  &  (~ n664)  &  n689 ) | ( (~ n664)  &  n689  &  n688 ) ;
 assign n692 = ( (~ i_30_)  &  n531 ) ;
 assign n691 = ( n495  &  n677 ) | ( n495  &  n692  &  (~ n973) ) ;
 assign n695 = ( n96 ) | ( n522 ) ;
 assign n696 = ( n96 ) | ( n609 ) ;
 assign n694 = ( (~ n404)  &  n653 ) | ( (~ n404)  &  n695 ) | ( n653  &  n696 ) | ( n695  &  n696 ) ;
 assign n698 = ( n1174  &  n555 ) | ( n1174  &  n611 ) | ( n1174  &  n649 ) ;
 assign n699 = ( (~ n404)  &  n653 ) | ( n653  &  n1021 ) | ( (~ n404)  &  n1023 ) | ( n1021  &  n1023 ) ;
 assign n697 = ( n698  &  n699  &  i_33_ ) | ( n698  &  n699  &  n694 ) ;
 assign n700 = ( i_28_ ) | ( n376 ) | ( (~ n833) ) ;
 assign n703 = ( n1260  &  n517 ) ;
 assign n704 = ( i_14_ ) | ( n1014 ) | ( n556 ) ;
 assign n702 = ( n703  &  n648 ) | ( n345  &  n648 ) | ( n703  &  n704 ) | ( n345  &  n704 ) ;
 assign n705 = ( (~ n243)  &  (~ n700) ) | ( n121  &  (~ n243)  &  (~ n716) ) ;
 assign n710 = ( (~ n356) ) | ( n572 ) | ( n1022 ) ;
 assign n709 = ( n649  &  (~ n705)  &  n710 ) | ( n702  &  (~ n705)  &  n710 ) ;
 assign n712 = ( n347  &  (~ n367) ) | ( n347  &  n480 ) | ( (~ n367)  &  n696 ) | ( n480  &  n696 ) ;
 assign n714 = ( (~ n350) ) | ( n561 ) | ( n1021 ) ;
 assign n713 = ( n714  &  n712 ) | ( n714  &  n446 ) ;
 assign n718 = ( (~ i_37_) ) | ( n334 ) | ( n479 ) ;
 assign n716 = ( i_34_ ) | ( n970 ) ;
 assign n717 = ( (~ i_35_) ) | ( (~ i_37_) ) ;
 assign n715 = ( (~ n688)  &  n718 ) | ( n718  &  n716 ) | ( n718  &  n717 ) ;
 assign n720 = ( n460 ) | ( (~ n467) ) | ( n628 ) ;
 assign n721 = ( n640 ) | ( n1009 ) | ( n587 ) ;
 assign n719 = ( n720  &  n721  &  n518 ) | ( n720  &  n721  &  n470 ) ;
 assign n723 = ( i_27_ ) | ( n995 ) ;
 assign n724 = ( (~ i_31_) ) | ( (~ i_34_) ) ;
 assign n722 = ( (~ n253)  &  n649 ) | ( n649  &  n723 ) | ( (~ n253)  &  n724 ) | ( n723  &  n724 ) ;
 assign n725 = ( (~ i_31_)  &  (~ n362) ) | ( (~ n362)  &  n664 ) | ( (~ i_31_)  &  n724 ) | ( n664  &  n724 ) ;
 assign n727 = ( n215 ) | ( (~ n253) ) | ( n315 ) ;
 assign n728 = ( (~ i_20_) ) | ( n722 ) | ( n960 ) ;
 assign n726 = ( n727  &  n728  &  n725 ) | ( n727  &  n728  &  n608 ) ;
 assign n729 = ( n364  &  (~ n725) ) ;
 assign n731 = ( n15  &  n729 ) | ( n729  &  (~ n1030) ) | ( n15  &  (~ n1170) ) | ( (~ n1030)  &  (~ n1170) ) ;
 assign n734 = ( i_16_ ) | ( i_13_ ) ;
 assign n735 = ( i_16_ ) | ( i_14_ ) ;
 assign n733 = ( n726  &  (~ n731) ) | ( (~ n731)  &  n734  &  n735 ) ;
 assign n739 = ( n138 ) | ( n497 ) | ( i_34_ ) | ( i_24_ ) ;
 assign n737 = ( i_28_  &  n739 ) | ( (~ n246)  &  n739 ) | ( (~ n290)  &  n739 ) ;
 assign n741 = ( (~ n11) ) | ( n684 ) ;
 assign n740 = ( (~ i_20_)  &  n497 ) | ( n497  &  n737 ) | ( (~ i_20_)  &  n741 ) | ( n737  &  n741 ) ;
 assign n743 = ( n514  &  n452 ) | ( n444  &  n452 ) | ( n514  &  n653 ) | ( n444  &  n653 ) ;
 assign n744 = ( n469  &  n501 ) | ( n469  &  n518 ) | ( n501  &  (~ n543) ) | ( n518  &  (~ n543) ) ;
 assign n747 = ( n627 ) | ( (~ n681) ) | ( n975 ) ;
 assign n746 = ( i_19_ ) | ( n1008 ) ;
 assign n745 = ( n747  &  n744 ) | ( n747  &  n84 ) | ( n747  &  n746 ) ;
 assign n749 = ( i_14_ ) | ( n40 ) | ( (~ n364) ) ;
 assign n748 = ( n749  &  n546 ) | ( n749  &  n453 ) ;
 assign n750 = ( (~ i_30_)  &  (~ n1182) ) | ( (~ i_30_)  &  i_34_  &  (~ n616) ) ;
 assign n754 = ( n1009 ) | ( n527 ) | ( n638 ) | ( n965 ) ;
 assign n755 = ( n630 ) | ( n907 ) | ( i_0_ ) | ( i_8_ ) ;
 assign n756 = ( n1198  &  n641 ) | ( n1198  &  n241 ) | ( n1198  &  n649 ) ;
 assign n757 = ( n608  &  n1199  &  n1201 ) | ( (~ n1164)  &  n1199  &  n1201 ) ;
 assign n758 = ( (~ i_25_)  &  n448 ) | ( n448  &  n740 ) | ( (~ i_25_)  &  n743 ) | ( n740  &  n743 ) ;
 assign n759 = ( n450  &  n745 ) | ( n748  &  n745 ) | ( n450  &  n1015 ) | ( n748  &  n1015 ) ;
 assign n760 = ( n1202  &  n884 ) | ( n1202  &  n1172  &  n1203 ) ;
 assign n761 = ( (~ n750)  &  (~ n1033)  &  n1204  &  n1205  &  n1206  &  n1207  &  n1208  &  n1210 ) ;
 assign n753 = ( n754  &  n755  &  n756  &  n757  &  n758  &  n759  &  n760  &  n761 ) ;
 assign n763 = ( (~ i_13_) ) | ( n735 ) ;
 assign n762 = ( i_12_  &  (~ i_13_) ) | ( i_12_  &  n453 ) | ( (~ i_13_)  &  n763 ) | ( n453  &  n763 ) ;
 assign n764 = ( n522  &  n453 ) ;
 assign n765 = ( i_10_  &  (~ i_13_) ) | ( i_10_  &  n453 ) | ( (~ i_13_)  &  n522 ) | ( n453  &  n522 ) ;
 assign n767 = ( (~ i_3_) ) | ( i_4_ ) | ( i_5_ ) ;
 assign n766 = ( n586 ) | ( i_6_ ) | ( n767 ) ;
 assign n769 = ( i_4_ ) | ( n373 ) ;
 assign n768 = ( (~ i_2_)  &  i_8_ ) | ( (~ i_2_)  &  n769 ) | ( (~ i_2_)  &  (~ n951) ) ;
 assign n771 = ( (~ i_7_)  &  (~ i_32_)  &  i_36_  &  (~ n769) ) ;
 assign n773 = ( (~ n765)  &  (~ n768) ) | ( (~ n765)  &  n771 ) ;
 assign n777 = ( (~ i_13_)  &  (~ n766) ) | ( (~ i_13_)  &  (~ n575)  &  (~ n769) ) ;
 assign n778 = ( (~ i_32_)  &  n951 ) ;
 assign n776 = ( (~ i_9_)  &  n773 ) | ( (~ i_9_)  &  n777  &  n778 ) ;
 assign n782 = ( (~ n290)  &  n1242 ) | ( (~ n951)  &  n1242 ) | ( n1242  &  n1241 ) ;
 assign n781 = ( i_31_ ) | ( n769 ) | ( (~ n778) ) | ( n1241 ) ;
 assign n779 = ( (~ i_29_)  &  n782 ) | ( (~ n776)  &  n782  &  n781 ) ;
 assign n784 = ( n1261  &  n654 ) ;
 assign n785 = ( n1021  &  n696 ) ;
 assign n783 = ( (~ i_36_)  &  n784 ) | ( n784  &  n785 ) | ( (~ i_36_)  &  (~ n951) ) | ( n785  &  (~ n951) ) ;
 assign n789 = ( n546 ) | ( n522 ) ;
 assign n787 = ( n608  &  (~ n778) ) | ( (~ n778)  &  n783 ) | ( n608  &  n789 ) | ( n783  &  n789 ) ;
 assign n790 = ( n620  &  n609 ) ;
 assign n792 = ( n607  &  n619 ) ;
 assign n791 = ( (~ n364)  &  n608 ) | ( (~ n364)  &  n790 ) | ( n608  &  n792 ) | ( n790  &  n792 ) ;
 assign n794 = ( n1259  &  n749 ) ;
 assign n793 = ( n794  &  n791 ) | ( n174  &  n791 ) | ( n794  &  n243 ) | ( n174  &  n243 ) ;
 assign n795 = ( n539  &  (~ n769) ) ;
 assign n797 = ( i_9_ ) | ( n769 ) ;
 assign n798 = ( n505  &  n763 ) ;
 assign n796 = ( (~ n229) ) | ( (~ n531) ) | ( n797 ) | ( n798 ) ;
 assign n801 = ( (~ i_21_)  &  n1003 ) ;
 assign n800 = ( (~ i_28_)  &  n234 ) ;
 assign n799 = ( n13  &  n801  &  n795 ) | ( n13  &  n801  &  n800 ) ;
 assign n802 = ( (~ n796)  &  (~ n1040) ) | ( (~ i_28_)  &  (~ n785)  &  (~ n1040) ) ;
 assign n806 = ( n367  &  (~ n1163) ) | ( n367  &  (~ n1179) ) ;
 assign n809 = ( i_19_ ) | ( (~ n229) ) | ( n518 ) | ( n797 ) ;
 assign n810 = ( n767 ) | ( n640 ) | ( n98 ) | ( i_18_ ) ;
 assign n813 = ( (~ n362) ) | ( (~ n467) ) ;
 assign n812 = ( i_21_ ) | ( (~ n833) ) ;
 assign n811 = ( n813  &  n664 ) | ( n813  &  n812 ) ;
 assign n814 = ( (~ n573)  &  (~ n824) ) | ( (~ n811)  &  (~ n824) ) ;
 assign n818 = ( n467  &  (~ n644) ) | ( n467  &  (~ n659) ) ;
 assign n821 = ( n404  &  (~ n785) ) | ( (~ i_32_)  &  n404  &  (~ n1272) ) ;
 assign n826 = ( n828 ) | ( n556 ) | ( n444 ) ;
 assign n824 = ( n1023  &  n695 ) ;
 assign n823 = ( n653  &  (~ n821)  &  n826 ) | ( (~ n821)  &  n826  &  n824 ) ;
 assign n829 = ( n215 ) | ( (~ n367) ) | ( n1272 ) ;
 assign n828 = ( n1017  &  n1028 ) ;
 assign n827 = ( (~ n362)  &  n829 ) | ( n556  &  n829 ) | ( n829  &  n828 ) ;
 assign n830 = ( i_7_  &  n215 ) | ( n215  &  (~ n290) ) | ( i_7_  &  n785 ) | ( (~ n290)  &  n785 ) ;
 assign n832 = ( (~ i_32_)  &  i_34_  &  (~ i_35_) ) ;
 assign n833 = ( (~ i_23_)  &  (~ i_24_) ) ;
 assign n831 = ( (~ n243)  &  n832  &  n833 ) ;
 assign n834 = ( (~ n544)  &  (~ n647) ) | ( (~ n647)  &  (~ n1179) ) ;
 assign n837 = ( (~ n570)  &  (~ n642) ) | ( (~ n570)  &  (~ n659) ) ;
 assign n841 = ( (~ i_29_)  &  n253 ) ;
 assign n840 = ( (~ i_28_)  &  n831 ) | ( (~ i_28_)  &  (~ n830)  &  n841 ) ;
 assign n843 = ( n362  &  n818 ) | ( n362  &  (~ n789)  &  n832 ) ;
 assign n845 = ( (~ i_32_)  &  n814 ) | ( (~ i_7_)  &  (~ i_32_)  &  (~ n1043) ) ;
 assign n847 = ( n10  &  n799 ) | ( n10  &  n802 ) | ( n10  &  n806 ) ;
 assign n849 = ( (~ i_33_) ) | ( n1004 ) ;
 assign n848 = ( (~ n245)  &  (~ n253) ) | ( (~ n253)  &  n649 ) | ( (~ n245)  &  n849 ) | ( n649  &  n849 ) ;
 assign n851 = ( n1260  &  n1169 ) ;
 assign n850 = ( n517  &  i_31_ ) | ( n517  &  n851 ) ;
 assign n853 = ( n1231  &  n868 ) | ( n1231  &  n174 ) | ( n1231  &  n649 ) ;
 assign n854 = ( (~ n404)  &  n653 ) | ( n653  &  n784 ) | ( (~ n404)  &  n1228 ) | ( n784  &  n1228 ) ;
 assign n852 = ( n853  &  n854  &  n850 ) | ( n853  &  n854  &  n444 ) ;
 assign n855 = ( i_31_  &  n135 ) | ( n135  &  (~ n531) ) | ( n135  &  n769 ) ;
 assign n856 = ( (~ i_8_)  &  (~ n1043) ) ;
 assign n857 = ( n362  &  (~ n794)  &  (~ n973) ) ;
 assign n859 = ( (~ i_31_)  &  n856 ) | ( (~ i_31_)  &  (~ n811)  &  (~ n1276) ) ;
 assign n861 = ( n10  &  (~ n1229) ) | ( n10  &  n350  &  (~ n517) ) ;
 assign n866 = ( i_31_ ) | ( n31 ) | ( (~ n467) ) | ( n1004 ) | ( n1014 ) ;
 assign n864 = ( (~ n681)  &  n866 ) | ( n797  &  n866 ) | ( n866  &  (~ n1044) ) ;
 assign n868 = ( n534  &  n704 ) ;
 assign n867 = ( (~ n10) ) | ( n170 ) | ( n868 ) ;
 assign n870 = ( (~ i_34_)  &  n121  &  (~ n243) ) ;
 assign n872 = ( (~ i_14_)  &  (~ i_25_) ) ;
 assign n871 = ( n497 ) | ( n872 ) | ( i_28_ ) | ( i_30_ ) ;
 assign n875 = ( i_24_ ) | ( (~ n290) ) | ( (~ n531) ) ;
 assign n874 = ( n479  &  (~ n688) ) ;
 assign n873 = ( (~ i_29_)  &  n875 ) | ( n649  &  n875 ) | ( n875  &  n874 ) ;
 assign n880 = ( n833  &  i_21_ ) ;
 assign n876 = ( (~ n871)  &  n880 ) | ( (~ n723)  &  n880  &  (~ n1038) ) ;
 assign n882 = ( (~ n10)  &  n238 ) | ( (~ n10)  &  n649 ) | ( n238  &  n995 ) | ( n649  &  n995 ) ;
 assign n881 = ( n211  &  n882 ) | ( (~ n362)  &  n882 ) ;
 assign n884 = ( i_23_ ) | ( n1004 ) ;
 assign n883 = ( n884  &  n572 ) | ( n211  &  n572 ) | ( n884  &  n236 ) | ( n211  &  n236 ) ;
 assign n886 = ( (~ i_21_) ) | ( n883 ) | ( n1006 ) ;
 assign n885 = ( n886  &  n881 ) | ( n886  &  n556 ) ;
 assign n888 = ( i_11_ ) | ( n1036 ) ;
 assign n889 = ( (~ i_3_) ) | ( n1036 ) ;
 assign n887 = ( i_19_  &  i_18_ ) | ( n888  &  i_18_ ) | ( i_19_  &  n889 ) | ( n888  &  n889 ) ;
 assign n891 = ( i_21_  &  (~ i_23_) ) ;
 assign n890 = ( i_25_  &  (~ n849)  &  n891 ) ;
 assign n892 = ( n290  &  n531  &  i_22_ ) ;
 assign n893 = ( (~ n479)  &  n890 ) | ( (~ n479)  &  n672  &  n673 ) ;
 assign n895 = ( i_18_ ) | ( n81 ) | ( n767 ) ;
 assign n894 = ( i_7_  &  n895 ) | ( (~ n19)  &  n895 ) | ( n797  &  n895 ) ;
 assign n897 = ( (~ i_2_) ) | ( (~ i_3_) ) | ( i_9_ ) ;
 assign n896 = ( n84  &  n897 ) | ( n767  &  n897 ) | ( n897  &  (~ n951) ) ;
 assign n898 = ( (~ i_9_)  &  n19  &  (~ n768) ) ;
 assign n899 = ( n531  &  n898 ) | ( (~ i_18_)  &  n531  &  (~ n896) ) ;
 assign n901 = ( (~ i_36_)  &  (~ n899) ) | ( (~ n539)  &  (~ n899) ) | ( n894  &  (~ n899) ) ;
 assign n904 = ( i_31_  &  (~ n1279) ) | ( n334  &  (~ n1279) ) | ( (~ n692)  &  (~ n1279) ) ;
 assign n907 = ( (~ n467) ) | ( n1005 ) ;
 assign n906 = ( (~ n681)  &  n907 ) | ( n769  &  n907 ) ;
 assign n909 = ( n192 ) | ( n608 ) | ( n664 ) ;
 assign n908 = ( (~ n11)  &  n909 ) | ( n215  &  n909 ) | ( n334  &  n909 ) ;
 assign n911 = ( (~ i_34_) ) | ( (~ i_36_) ) | ( (~ n234) ) ;
 assign n910 = ( (~ i_36_)  &  (~ n404) ) | ( (~ n404)  &  n908 ) | ( (~ i_36_)  &  n911 ) | ( n908  &  n911 ) ;
 assign n912 = ( i_2_ ) | ( n135 ) | ( (~ n778) ) ;
 assign n916 = ( (~ n9)  &  (~ n1281) ) | ( (~ n229)  &  (~ n1281) ) | ( n556  &  (~ n1281) ) ;
 assign n914 = ( i_7_  &  n1040 ) | ( n910  &  n1040 ) | ( i_7_  &  (~ n1216) ) | ( n910  &  (~ n1216) ) ;
 assign n915 = ( (~ i_21_)  &  n1257 ) | ( n883  &  n1257 ) | ( n931  &  n1257 ) ;
 assign n913 = ( n916  &  i_16_ ) | ( n916  &  n914  &  n915 ) ;
 assign n917 = ( n548  &  n547 ) | ( n888  &  n547 ) | ( n548  &  n889 ) | ( n888  &  n889 ) ;
 assign n919 = ( n722 ) | ( n887 ) | ( (~ n891) ) ;
 assign n918 = ( n919  &  n725 ) | ( n919  &  n917 ) ;
 assign n920 = ( i_16_  &  i_17_ ) | ( i_16_  &  n216 ) | ( i_17_  &  (~ n363) ) | ( n216  &  (~ n363) ) ;
 assign n922 = ( n497 ) | ( n741 ) ;
 assign n921 = ( (~ i_21_)  &  (~ n407)  &  n922 ) | ( (~ n407)  &  n737  &  n922 ) ;
 assign n926 = ( n791 ) | ( n1039 ) | ( i_31_ ) | ( i_30_ ) ;
 assign n924 = ( (~ n13)  &  n926 ) | ( (~ n364)  &  n926 ) | ( n911  &  n926 ) ;
 assign n927 = ( (~ i_31_)  &  (~ n467) ) | ( (~ n467)  &  n573 ) | ( (~ i_31_)  &  n723 ) | ( n573  &  n723 ) ;
 assign n931 = ( i_12_ ) | ( n1035 ) ;
 assign n929 = ( (~ n9)  &  n881 ) | ( n559  &  n881 ) | ( (~ n9)  &  n931 ) | ( n559  &  n931 ) ;
 assign n939 = ( (~ i_21_)  &  (~ n1280) ) | ( i_20_  &  (~ i_21_)  &  (~ n904) ) ;
 assign n942 = ( n253  &  n892 ) | ( n253  &  n893 ) | ( n253  &  (~ n1223) ) ;
 assign n944 = ( i_34_  &  (~ n496) ) | ( i_34_  &  n876 ) | ( i_34_  &  (~ n1224) ) ;
 assign n947 = ( n778  &  (~ n867) ) | ( n778  &  n870 ) | ( n778  &  (~ n1227) ) ;
 assign n951 = ( (~ i_35_)  &  i_36_ ) ;
 assign n950 = ( n951  &  n857 ) | ( n951  &  n859 ) | ( n951  &  n861 ) ;
 assign n953 = ( i_12_ ) | ( n735 ) ;
 assign n954 = ( i_21_ ) | ( i_22_ ) ;
 assign n957 = ( (~ i_16_)  &  (~ i_27_) ) ;
 assign n960 = ( i_23_ ) | ( i_17_ ) ;
 assign n961 = ( i_2_ ) | ( i_4_ ) ;
 assign n962 = ( (~ i_9_) ) | ( n373 ) ;
 assign n963 = ( i_28_ ) | ( i_26_ ) ;
 assign n964 = ( i_8_ ) | ( (~ i_9_) ) ;
 assign n965 = ( i_8_ ) | ( n373 ) ;
 assign n966 = ( i_2_ ) | ( i_3_ ) ;
 assign n968 = ( i_33_ ) | ( (~ n234) ) ;
 assign n969 = ( (~ i_9_) ) | ( n966 ) ;
 assign n970 = ( i_33_ ) | ( i_32_ ) ;
 assign n972 = ( i_31_ ) | ( n970 ) ;
 assign n973 = ( (~ i_34_) ) | ( n685 ) ;
 assign n974 = ( i_30_ ) | ( i_29_ ) ;
 assign n975 = ( i_8_ ) | ( n372 ) ;
 assign n977 = ( i_4_ ) | ( n966 ) ;
 assign n978 = ( i_29_ ) | ( (~ i_34_) ) ;
 assign n979 = ( (~ i_9_) ) | ( (~ n23) ) ;
 assign n983 = ( (~ i_3_) ) | ( n961 ) ;
 assign n984 = ( n983 ) | ( n595 ) ;
 assign n985 = ( i_9_ ) | ( n984 ) ;
 assign n986 = ( n371 ) | ( n98 ) ;
 assign n987 = ( i_3_ ) | ( i_7_ ) | ( (~ i_10_) ) ;
 assign n988 = ( i_33_ ) | ( (~ i_34_) ) | ( i_35_ ) ;
 assign n989 = ( i_9_ ) | ( i_6_ ) ;
 assign n990 = ( n965 ) | ( n983 ) ;
 assign n991 = ( i_11_ ) | ( n989 ) ;
 assign n992 = ( i_7_ ) | ( n372 ) ;
 assign n993 = ( (~ n11) ) | ( (~ n833) ) ;
 assign n994 = ( (~ n394) ) | ( n974 ) ;
 assign n995 = ( i_28_ ) | ( (~ i_31_) ) ;
 assign n996 = ( i_7_ ) | ( i_28_ ) | ( n192 ) ;
 assign n997 = ( i_8_ ) | ( n966 ) ;
 assign n998 = ( i_22_ ) | ( (~ n531) ) | ( n874 ) | ( (~ n891) ) ;
 assign n1000 = ( i_12_ ) | ( n962 ) | ( n977 ) ;
 assign n1001 = ( i_2_ ) | ( i_7_ ) | ( (~ i_38_) ) ;
 assign n1002 = ( n30 ) | ( n31 ) ;
 assign n1003 = ( (~ i_16_)  &  (~ i_23_) ) ;
 assign n1004 = ( i_27_ ) | ( i_28_ ) ;
 assign n1005 = ( i_30_ ) | ( n1004 ) ;
 assign n1006 = ( i_16_ ) | ( i_17_ ) ;
 assign n1007 = ( i_0_ ) | ( i_4_ ) ;
 assign n1008 = ( i_17_ ) | ( i_20_ ) | ( (~ n681) ) ;
 assign n1009 = ( i_18_ ) | ( n1008 ) ;
 assign n1010 = ( i_19_ ) | ( n1006 ) ;
 assign n1011 = ( i_12_ ) | ( n734 ) ;
 assign n1012 = ( n371 ) | ( n992 ) ;
 assign n1013 = ( i_18_ ) | ( n960 ) ;
 assign n1014 = ( n373 ) | ( n374 ) ;
 assign n1015 = ( i_5_ ) | ( n1007 ) ;
 assign n1016 = ( n98 ) | ( n1015 ) ;
 assign n1017 = ( (~ i_13_) ) | ( i_14_ ) | ( n70 ) ;
 assign n1018 = ( n371 ) | ( n975 ) ;
 assign n1019 = ( i_23_ ) | ( n735 ) ;
 assign n1020 = ( (~ i_13_) ) | ( n989 ) ;
 assign n1021 = ( n96 ) | ( n620 ) ;
 assign n1022 = ( n63 ) | ( n453 ) ;
 assign n1023 = ( n96 ) | ( n453 ) ;
 assign n1024 = ( (~ i_23_)  &  (~ i_27_) ) ;
 assign n1025 = ( (~ i_25_) ) | ( n1004 ) ;
 assign n1026 = ( (~ i_20_) ) | ( (~ n833) ) ;
 assign n1027 = ( i_20_ ) | ( (~ n833) ) ;
 assign n1028 = ( i_13_ ) | ( i_10_ ) | ( n70 ) ;
 assign n1029 = ( n66 ) | ( n505 ) ;
 assign n1030 = ( i_14_ ) | ( i_12_ ) ;
 assign n1033 = ( n679 ) | ( (~ n683) ) | ( n686 ) | ( n691 ) ;
 assign n1035 = ( (~ i_7_) ) | ( i_9_ ) ;
 assign n1036 = ( (~ i_7_) ) | ( (~ i_10_) ) ;
 assign n1038 = ( n762 ) | ( n1036 ) ;
 assign n1039 = ( (~ i_34_) ) | ( (~ n951) ) ;
 assign n1040 = ( i_21_ ) | ( n960 ) ;
 assign n1041 = ( (~ i_20_) ) | ( i_21_ ) | ( i_23_ ) ;
 assign n1042 = ( i_21_ ) | ( n1006 ) ;
 assign n1043 = ( n907 ) | ( n1042 ) | ( i_2_ ) | ( n31 ) ;
 assign n1044 = ( (~ i_10_)  &  (~ i_13_) ) | ( (~ i_10_)  &  (~ i_14_) ) | ( i_13_  &  (~ i_14_) ) ;
 assign n1045 = ( n170  &  n86 ) | ( n376  &  n86 ) | ( n170  &  n174 ) | ( n376  &  n174 ) ;
 assign n1046 = ( n195  &  (~ n313) ) | ( (~ n313)  &  n972 ) | ( n195  &  n973 ) | ( n972  &  n973 ) ;
 assign n1047 = ( (~ n15)  &  n38 ) | ( n38  &  n72 ) | ( (~ n15)  &  n261 ) | ( n72  &  n261 ) ;
 assign n1048 = ( (~ n23)  &  n63 ) | ( n64  &  n63 ) | ( (~ n23)  &  n979 ) | ( n64  &  n979 ) ;
 assign n1050 = ( (~ i_19_) ) | ( n163 ) | ( n347 ) ;
 assign n1049 = ( n1050  &  i_28_ ) | ( n1050  &  n345 ) | ( n1050  &  n199 ) ;
 assign n1051 = ( n200  &  (~ n382) ) | ( n195  &  (~ n356)  &  (~ n382) ) ;
 assign n1053 = ( (~ n121)  &  (~ n378) ) | ( n190  &  (~ n378) ) | ( (~ n378)  &  n611 ) ;
 assign n1055 = ( (~ n11)  &  n86 ) | ( n86  &  n375 ) | ( (~ n11)  &  n377 ) | ( n375  &  n377 ) ;
 assign n1057 = ( n1018  &  n63 ) ;
 assign n1056 = ( n143  &  n168 ) | ( n168  &  (~ n356) ) | ( n143  &  n1057 ) | ( (~ n356)  &  n1057 ) ;
 assign n1058 = ( n78  &  (~ n385)  &  n1056 ) | ( n344  &  (~ n385)  &  n1056 ) ;
 assign n1060 = ( (~ n95)  &  n841 ) | ( n331  &  n841 ) ;
 assign n1062 = ( n130  &  (~ n304) ) | ( (~ n304)  &  n963 ) | ( n130  &  n978 ) | ( n963  &  n978 ) ;
 assign n1063 = ( n92  &  (~ n337) ) | ( n170  &  (~ n337) ) | ( (~ n337)  &  (~ n832) ) ;
 assign n1065 = ( n91 ) | ( n130 ) ;
 assign n1066 = ( (~ n121)  &  (~ n304) ) | ( n241  &  (~ n304) ) | ( (~ n121)  &  n648 ) | ( n241  &  n648 ) ;
 assign n1068 = ( i_28_ ) | ( (~ n229) ) | ( n611 ) ;
 assign n1067 = ( i_7_  &  n1068 ) | ( (~ n350)  &  n1068 ) | ( n968  &  n1068 ) ;
 assign n1070 = ( (~ n313)  &  n347 ) ;
 assign n1069 = ( n1070  &  n65 ) | ( n283  &  n65 ) | ( n1070  &  n240 ) | ( n283  &  n240 ) ;
 assign n1072 = ( n170 ) | ( n101 ) | ( n92 ) | ( n163 ) ;
 assign n1071 = ( i_25_  &  n1072 ) | ( i_28_  &  n1072 ) | ( (~ n1060)  &  n1072 ) ;
 assign n1073 = ( (~ i_35_)  &  n1071 ) | ( n69  &  n1071 ) | ( n339  &  n1071 ) ;
 assign n1074 = ( n243  &  (~ n348)  &  n1073 ) | ( n342  &  (~ n348)  &  n1073 ) ;
 assign n1076 = ( n133  &  (~ n352)  &  (~ n355) ) | ( n249  &  (~ n352)  &  (~ n355) ) ;
 assign n1079 = ( n248  &  (~ n358)  &  n1076 ) | ( n332  &  (~ n358)  &  n1076 ) ;
 assign n1082 = ( i_30_ ) | ( (~ n313) ) | ( (~ n414) ) ;
 assign n1081 = ( (~ n32)  &  n1082 ) | ( n347  &  n1082 ) ;
 assign n1083 = ( i_24_  &  (~ n26) ) | ( i_24_  &  (~ n367) ) | ( (~ n26)  &  n996 ) | ( (~ n367)  &  n996 ) ;
 assign n1084 = ( (~ n11)  &  n283 ) | ( (~ n11)  &  (~ n308) ) | ( n283  &  (~ n414) ) | ( (~ n308)  &  (~ n414) ) ;
 assign n1085 = ( (~ n317)  &  (~ n322) ) | ( (~ n317)  &  n1083  &  n1084 ) ;
 assign n1087 = ( i_13_ ) | ( i_24_ ) ;
 assign n1088 = ( n191  &  n194 ) | ( n1087  &  n194 ) | ( n191  &  n145 ) | ( n1087  &  n145 ) ;
 assign n1089 = ( n127  &  (~ n274) ) | ( (~ n256)  &  (~ n274) ) | ( (~ n274)  &  n997 ) ;
 assign n1092 = ( i_2_ ) | ( (~ n22) ) | ( n49 ) ;
 assign n1091 = ( n1092  &  i_13_ ) | ( n1092  &  i_3_ ) | ( n1092  &  n198 ) ;
 assign n1094 = ( n136 ) | ( n189 ) | ( (~ n229) ) ;
 assign n1093 = ( (~ i_12_)  &  (~ n278)  &  n1094 ) | ( n273  &  (~ n278)  &  n1094 ) ;
 assign n1097 = ( i_26_  &  (~ n841) ) | ( (~ n35)  &  (~ n841) ) | ( i_26_  &  (~ n1002) ) | ( (~ n35)  &  (~ n1002) ) ;
 assign n1100 = ( n146 ) | ( n240 ) | ( n162 ) ;
 assign n1099 = ( n1100  &  i_28_ ) | ( n1100  &  n242 ) | ( n1100  &  n124 ) ;
 assign n1101 = ( (~ i_23_)  &  n237 ) | ( n237  &  (~ n356) ) | ( (~ i_23_)  &  n957 ) | ( (~ n356)  &  n957 ) ;
 assign n1102 = ( n53  &  (~ n230) ) | ( (~ n230)  &  (~ n282) ) | ( (~ n230)  &  (~ n279) ) ;
 assign n1107 = ( (~ i_18_) ) | ( i_24_ ) | ( n191 ) ;
 assign n1106 = ( n1107  &  n194 ) | ( n1107  &  n144 ) ;
 assign n1108 = ( n163  &  n207 ) | ( n163  &  (~ n350) ) | ( n207  &  n995 ) | ( (~ n350)  &  n995 ) ;
 assign n1109 = ( (~ i_9_)  &  (~ n41)  &  (~ n45) ) | ( n36  &  (~ n41)  &  (~ n45) ) ;
 assign n1112 = ( n39  &  (~ n256) ) | ( n147  &  (~ n256) ) | ( n39  &  n1000 ) | ( n147  &  n1000 ) ;
 assign n1114 = ( n1020  &  n454 ) ;
 assign n1113 = ( n1114  &  n69 ) | ( n173  &  n69 ) | ( n1114  &  n164 ) | ( n173  &  n164 ) ;
 assign n1115 = ( n140  &  n143 ) | ( n140  &  (~ n394) ) | ( n143  &  (~ n402) ) | ( (~ n394)  &  (~ n402) ) ;
 assign n1116 = ( i_31_ ) | ( n1127 ) | ( n90 ) ;
 assign n1117 = ( i_2_ ) | ( i_8_ ) | ( n135 ) | ( (~ n394) ) ;
 assign n1120 = ( (~ i_34_) ) | ( (~ n531) ) | ( n680 ) ;
 assign n1118 = ( n78  &  n1120 ) | ( (~ n107)  &  n1120 ) | ( (~ n394)  &  n1120 ) ;
 assign n1122 = ( n89 ) | ( n97 ) | ( n148 ) ;
 assign n1121 = ( (~ i_13_)  &  n1122 ) | ( n85  &  n1122 ) | ( n371  &  n1122 ) ;
 assign n1124 = ( i_2_ ) | ( n972 ) | ( n131 ) ;
 assign n1123 = ( n86  &  (~ n105)  &  n1124 ) | ( n102  &  (~ n105)  &  n1124 ) ;
 assign n1128 = ( i_2_ ) | ( i_8_ ) | ( i_31_ ) | ( (~ n306) ) ;
 assign n1127 = ( n1014  &  n40 ) ;
 assign n1126 = ( (~ n394)  &  n1128 ) | ( n972  &  n1128 ) | ( n1128  &  n1127 ) ;
 assign n1130 = ( i_10_ ) | ( n61 ) | ( (~ n402) ) ;
 assign n1129 = ( (~ i_29_)  &  n1130 ) | ( (~ n1002)  &  n1003  &  n1130 ) ;
 assign n1131 = ( n968  &  n57 ) | ( n1001  &  n57 ) | ( n968  &  n326 ) | ( n1001  &  n326 ) ;
 assign n1132 = ( n68  &  n1131 ) | ( (~ n322)  &  n1131 ) ;
 assign n1134 = ( (~ n253) ) | ( (~ n531) ) | ( n680 ) ;
 assign n1133 = ( (~ n44)  &  n1134 ) | ( n49  &  n1134 ) | ( n969  &  n1134 ) ;
 assign n1135 = ( (~ i_9_)  &  n1133 ) | ( (~ i_12_)  &  n1133 ) | ( n53  &  n1133 ) ;
 assign n1136 = ( n109  &  (~ n113)  &  (~ n117) ) | ( (~ n113)  &  (~ n117)  &  (~ n324) ) ;
 assign n1140 = ( n89 ) | ( n147 ) | ( (~ n429) ) ;
 assign n1139 = ( n1140  &  n140 ) | ( n1140  &  n1070 ) | ( n1140  &  n162 ) ;
 assign n1141 = ( i_35_ ) | ( n186 ) | ( n139 ) ;
 assign n1143 = ( (~ i_38_)  &  (~ n403) ) | ( (~ n403)  &  n1074  &  n1079 ) ;
 assign n1147 = ( n300  &  (~ n301)  &  (~ n305)  &  (~ n309)  &  n314  &  n1085  &  n1226  &  n1264 ) ;
 assign n1146 = ( i_29_  &  (~ i_34_) ) | ( (~ i_34_)  &  n319 ) | ( i_29_  &  n1147 ) | ( n319  &  n1147 ) ;
 assign n1149 = ( (~ n10)  &  (~ n408)  &  (~ n412) ) | ( (~ n408)  &  (~ n412)  &  n998 ) ;
 assign n1152 = ( n127  &  n122 ) | ( n264  &  n122 ) | ( n127  &  n260 ) | ( n264  &  n260 ) ;
 assign n1153 = ( i_24_  &  (~ n415) ) | ( (~ n415)  &  n1099  &  n1101 ) ;
 assign n1155 = ( n205  &  (~ n425) ) | ( (~ n425)  &  n1109  &  n1112 ) ;
 assign n1157 = ( n198  &  (~ n428)  &  n1155 ) | ( (~ n428)  &  n979  &  n1155 ) ;
 assign n1159 = ( n157  &  n132 ) | ( n195  &  n132 ) | ( n157  &  n265 ) | ( n195  &  n265 ) ;
 assign n1160 = ( n217  &  i_22_ ) | ( n217  &  n1136  &  n1135 ) ;
 assign n1163 = ( n1012 ) | ( n558 ) ;
 assign n1164 = ( (~ n447)  &  (~ n1261) ) | ( (~ n59)  &  (~ n447)  &  (~ n481) ) ;
 assign n1169 = ( n1018 ) | ( n1019 ) ;
 assign n1171 = ( n213 ) | ( (~ n253) ) | ( n315 ) ;
 assign n1170 = ( (~ i_20_)  &  n1171 ) | ( n722  &  n1171 ) | ( (~ n1003)  &  n1171 ) ;
 assign n1173 = ( (~ i_31_) ) | ( n715 ) | ( n974 ) ;
 assign n1172 = ( n1173  &  n642 ) | ( n1173  &  n340 ) | ( n1173  &  n717 ) ;
 assign n1174 = ( i_7_ ) | ( n972 ) | ( n993 ) ;
 assign n1175 = ( (~ n245)  &  (~ n667) ) | ( (~ n667)  &  n1025 ) | ( (~ n667)  &  n1026 ) ;
 assign n1179 = ( n1012 ) | ( n1019 ) ;
 assign n1180 = ( n649 ) | ( n1028 ) | ( n345 ) | ( n556 ) ;
 assign n1181 = ( i_0_ ) | ( i_30_ ) | ( (~ n229) ) | ( n477 ) | ( n664 ) | ( n1027 ) ;
 assign n1183 = ( n442 ) | ( n1019 ) | ( n559 ) ;
 assign n1182 = ( n1183  &  n447 ) | ( n1183  &  n618 ) ;
 assign n1186 = ( i_7_ ) | ( i_23_ ) | ( (~ n290) ) | ( (~ n308) ) | ( n443 ) ;
 assign n1187 = ( n501  &  (~ n543) ) | ( (~ n543)  &  n646 ) | ( n501  &  n1022 ) | ( n646  &  n1022 ) ;
 assign n1189 = ( (~ i_37_) ) | ( (~ n349) ) | ( n556 ) | ( n1028 ) ;
 assign n1188 = ( n376  &  n1189 ) | ( (~ n543)  &  n1189 ) | ( n612  &  n1189 ) ;
 assign n1191 = ( (~ i_2_) ) | ( i_16_ ) | ( n31 ) ;
 assign n1190 = ( n1191  &  n502 ) | ( n1191  &  n84 ) | ( n1191  &  n1015 ) ;
 assign n1192 = ( (~ i_37_) ) | ( n81 ) | ( n513 ) | ( n520 ) ;
 assign n1193 = ( n347  &  (~ n350) ) | ( n347  &  n514 ) | ( (~ n350)  &  n703 ) | ( n514  &  n703 ) ;
 assign n1195 = ( i_30_ ) | ( (~ i_31_) ) | ( (~ n362) ) | ( n479 ) ;
 assign n1194 = ( n1195  &  i_14_ ) | ( n1195  &  n631 ) | ( n1195  &  n461 ) ;
 assign n1197 = ( n373 ) | ( n474 ) | ( n622 ) | ( n631 ) | ( (~ n681) ) ;
 assign n1196 = ( n452  &  n1197 ) | ( (~ n543)  &  n1197 ) | ( n813  &  n1197 ) ;
 assign n1198 = ( n645 ) | ( n347 ) | ( n572 ) ;
 assign n1200 = ( (~ n692) ) | ( (~ n880) ) | ( n973 ) ;
 assign n1199 = ( n1200  &  n442 ) | ( n1200  &  n556 ) | ( n1200  &  n1017 ) ;
 assign n1201 = ( i_13_ ) | ( n624 ) | ( n631 ) ;
 assign n1202 = ( (~ i_7_)  &  n550 ) | ( (~ i_7_)  &  n719 ) | ( n550  &  n733 ) | ( n719  &  n733 ) ;
 assign n1203 = ( n241 ) | ( n446 ) | ( n695 ) ;
 assign n1204 = ( n215  &  (~ n543) ) | ( n215  &  n709 ) | ( (~ n543)  &  n713 ) | ( n709  &  n713 ) ;
 assign n1205 = ( n697  &  n874 ) | ( n443  &  n874 ) | ( n697  &  n674 ) | ( n443  &  n674 ) ;
 assign n1206 = ( (~ i_37_)  &  (~ n290) ) | ( (~ i_37_)  &  n634 ) | ( (~ n290)  &  n658 ) | ( n634  &  n658 ) ;
 assign n1207 = ( n613  &  i_14_ ) | ( n664  &  i_14_ ) | ( n613  &  n582 ) | ( n664  &  n582 ) ;
 assign n1209 = ( (~ n529)  &  n533  &  (~ n535)  &  (~ n540)  &  n998  &  n1268 ) ;
 assign n1208 = ( (~ n10)  &  (~ n362) ) | ( (~ n10)  &  n567 ) | ( (~ n362)  &  n1209 ) | ( n567  &  n1209 ) ;
 assign n1210 = ( i_32_  &  (~ i_34_) ) | ( (~ i_34_)  &  n486 ) | ( i_32_  &  n496 ) | ( n486  &  n496 ) ;
 assign n1214 = ( (~ i_34_) ) | ( n649 ) | ( n974 ) ;
 assign n1213 = ( i_30_  &  n1214 ) | ( (~ n253)  &  n1214 ) | ( (~ n362)  &  n1214 ) ;
 assign n1215 = ( (~ n363)  &  n479 ) | ( (~ n364)  &  n479 ) | ( (~ n363)  &  n498 ) | ( (~ n364)  &  n498 ) ;
 assign n1216 = ( n10  &  (~ n912) ) | ( i_0_  &  n10  &  n531 ) ;
 assign n1222 = ( n315 ) | ( (~ n688) ) | ( n887 ) | ( (~ n1024) ) ;
 assign n1220 = ( (~ n668)  &  n1222 ) | ( n995  &  n1222 ) | ( n1038  &  n1222 ) ;
 assign n1223 = ( (~ n494)  &  n1220 ) | ( n874  &  n1220 ) | ( n1041  &  n1220 ) ;
 assign n1225 = ( n315 ) | ( n572 ) | ( n1038 ) ;
 assign n1226 = ( (~ i_14_) ) | ( n497 ) | ( n993 ) ;
 assign n1224 = ( n1225  &  n1226  &  n873 ) | ( n1225  &  n1226  &  n1041 ) ;
 assign n1228 = ( n455  &  n554 ) ;
 assign n1227 = ( n864  &  n1228 ) | ( n1042  &  n1228 ) | ( n864  &  n813 ) | ( n1042  &  n813 ) ;
 assign n1230 = ( n792 ) | ( (~ n801) ) | ( n855 ) ;
 assign n1229 = ( n1230  &  n851 ) | ( n1230  &  n170 ) ;
 assign n1231 = ( n1276 ) | ( n170 ) | ( n572 ) ;
 assign n1232 = ( n681  &  (~ n809) ) | ( n681  &  (~ n810) ) ;
 assign n1237 = ( (~ n11) ) | ( (~ n13) ) | ( n213 ) | ( n334 ) ;
 assign n1236 = ( i_17_  &  n1237 ) | ( i_21_  &  n1237 ) | ( (~ n1232)  &  n1237 ) ;
 assign n1238 = ( n1236  &  i_7_ ) | ( n1236  &  n973 ) | ( n1236  &  n993 ) ;
 assign n1239 = ( (~ i_34_)  &  (~ n253) ) | ( (~ n253)  &  n823 ) | ( (~ i_34_)  &  n827 ) | ( n823  &  n827 ) ;
 assign n1242 = ( i_30_ ) | ( (~ i_36_) ) | ( n249 ) | ( n764 ) ;
 assign n1241 = ( n953  &  n1011 ) ;
 assign n1244 = ( (~ i_36_) ) | ( (~ n13) ) | ( n192 ) | ( (~ n364) ) ;
 assign n1243 = ( n614  &  n793  &  n1244 ) | ( n614  &  (~ n951)  &  n1244 ) ;
 assign n1245 = ( i_29_  &  n779 ) | ( n787  &  n779 ) | ( i_29_  &  n812 ) | ( n787  &  n812 ) ;
 assign n1247 = ( n848 ) | ( (~ n891) ) | ( n920 ) ;
 assign n1246 = ( n1247  &  n929 ) | ( n1247  &  n558  &  n1019 ) ;
 assign n1248 = ( n1246  &  n927 ) | ( n1246  &  n1038 ) ;
 assign n1249 = ( (~ n362)  &  n872 ) | ( (~ n362)  &  n921 ) | ( n872  &  n924 ) | ( n921  &  n924 ) ;
 assign n1250 = ( n31  &  (~ n688) ) | ( (~ n688)  &  n913 ) | ( n31  &  n918 ) | ( n913  &  n918 ) ;
 assign n1251 = ( (~ i_36_)  &  n852 ) | ( (~ i_36_)  &  n1039 ) | ( n852  &  (~ n1273) ) | ( n1039  &  (~ n1273) ) ;
 assign n1253 = ( n1251  &  n664 ) | ( n1251  &  n1245  &  n1243 ) ;
 assign n1256 = ( n608 ) | ( n501 ) | ( n654 ) | ( i_29_ ) ;
 assign n1257 = ( i_21_ ) | ( (~ i_36_) ) | ( n559 ) | ( n906 ) ;
 assign n1258 = ( i_33_ ) | ( n963 ) ;
 assign n1259 = ( i_13_ ) | ( n40 ) | ( (~ n364) ) ;
 assign n1260 = ( n558 ) | ( n1018 ) ;
 assign n1261 = ( n59 ) | ( n763 ) ;
 assign n1263 = ( n179 ) | ( n247 ) | ( (~ n322) ) ;
 assign n1264 = ( i_24_ ) | ( i_28_ ) | ( n289 ) ;
 assign n1268 = ( i_0_ ) | ( n500 ) | ( n511 ) | ( (~ n800) ) ;
 assign n1272 = ( n482  &  n1029 ) ;
 assign n1273 = ( n834 ) | ( n837 ) | ( n840 ) | ( n843 ) | ( n845 ) | ( n847 ) | ( (~ n1238) ) | ( (~ n1239) ) ;
 assign n1276 = ( n646  &  n1022 ) ;
 assign n1279 = ( (~ n163)  &  n290  &  n670 ) ;
 assign n1280 = ( i_23_ ) | ( (~ n10) ) | ( n522 ) | ( n901 ) ;
 assign n1281 = ( i_0_  &  (~ i_12_)  &  n10  &  n531  &  n801 ) ;


endmodule

