// sk = 0110011010011000111001010100010111001101
`timescale 10ns/1ns
module alu4_orig (/* input clk, */ input [39:0] sk, input n, input j, input k, input l, input i, input a, input e, input m, input b, input f, input c, input g, input d, input houtput wire o, output wire p, output wire q, output wire r, output wire s, output wire t, output wire u, output wire v);

//reg [13:0] inputs;
//reg [7:0] outputs;
//reg [39:0] sk_reg;
//always @(posedge clk) inputs = {n, j, k, l, i, a, e, m, b, f, c, g, d, h};
//always @(posedge clk) outputs = {o, p, q, r, s, t, u, v};
//always @(posedge clk) sk_reg = {o, p, q, r, s, t, u, v};

	wire g163, g121, g179, g182, g1, g8, g11, g9, g10, g12, g7;
	wire g13, g15, g17, g14, g16, g18, g19, g20, g22, g23, g27;
	wire g28, g26, g29, g21, g24, g25, g30, g33, g34, g35, g32;
	wire g36, g2, g3, g4, g41, g42, g38, g39, g40, g43, g44;
	wire g45, g46, g47, g50, g51, g54, g55, g48, g49, g52, g206;
	wire g62, g63, g64, g65, g67, g68, g69, g60, g61, g66, g70;
	wire g71, g58, g59, g72, g76, g74, g75, g77, g31, g73, g78;
	wire g81, g83, g84, g85, g86, g82, g87, g88, g89, g90, g53;
	wire g57, g92, g93, g95, g96, g91, g94, g97, g99, g100, g102;
	wire g103, g104, g106, g111, g108, g109, g110, g112, g98, g101, g105;
	wire g107, g113, g114, g118, g122, g123, g125, g126, g129, g130, g127;
	wire g128, g131, g124, g132, g133, g134, g120, g135, g136, g138, g139;
	wire g141, g147, g148, g149, g144, g145, g146, g150, g152, g153, g154;
	wire g137, g140, g142, g143, g151, g155, g159, g157, g158, g160, g80;
	wire g115, g156, g161, g168, g171, g183, g173, g169, g170, g172, g174;
	wire g165, g166, g167, g175, g164, g176, g178, g180, g181, g184, g185;
	wire g186, g189, g187, g188, g190, g191, g192, g194, g195, g196, g199;
	wire g197, g198, g202, g203, g200, g201, g204, g205, g119, g116, g117;
	wire g207, g208, g209, g212, g210, g211, g215, g216, g213, g214, g217;
	wire g218, g56, g220, g221, g222, g225, g223, g224, g228, g229, g226;
	wire g227, g230, g231, g37, g5, g6;


	assign g93 = (((!g82) & (sk[0]) & (g87)) + ((g82) & (!sk[0]) & (!g87)) + ((g82) & (!sk[0]) & (g87)));
	assign g7 = (((!n) & (!i) & (!sk[0]) & (j) & (!g1)) + ((!n) & (!i) & (!sk[0]) & (j) & (g1)) + ((!n) & (i) & (!sk[0]) & (j) & (!g1)) + ((!n) & (i) & (!sk[0]) & (j) & (g1)) + ((n) & (!i) & (!sk[0]) & (!j) & (g1)) + ((n) & (!i) & (!sk[0]) & (j) & (!g1)) + ((n) & (!i) & (!sk[0]) & (j) & (g1)) + ((n) & (i) & (!sk[0]) & (!j) & (g1)) + ((n) & (i) & (!sk[0]) & (j) & (!g1)) + ((n) & (i) & (!sk[0]) & (j) & (g1)) + ((n) & (i) & (sk[0]) & (!j) & (g1)));
	assign g44 = (((!a) & (!g11) & (!g38) & (!g39) & (!g40) & (g43)) + ((!a) & (!g11) & (!g38) & (!g39) & (g40) & (!g43)) + ((!a) & (!g11) & (!g38) & (!g39) & (g40) & (g43)) + ((!a) & (!g11) & (!g38) & (g39) & (!g40) & (g43)) + ((!a) & (!g11) & (!g38) & (g39) & (g40) & (!g43)) + ((!a) & (!g11) & (!g38) & (g39) & (g40) & (g43)) + ((!a) & (!g11) & (g38) & (!g39) & (!g40) & (g43)) + ((!a) & (!g11) & (g38) & (!g39) & (g40) & (!g43)) + ((!a) & (!g11) & (g38) & (!g39) & (g40) & (g43)) + ((!a) & (!g11) & (g38) & (g39) & (!g40) & (g43)) + ((!a) & (!g11) & (g38) & (g39) & (g40) & (!g43)) + ((!a) & (!g11) & (g38) & (g39) & (g40) & (g43)) + ((!a) & (g11) & (!g38) & (!g39) & (!g40) & (g43)) + ((!a) & (g11) & (!g38) & (!g39) & (g40) & (!g43)) + ((!a) & (g11) & (!g38) & (!g39) & (g40) & (g43)) + ((!a) & (g11) & (!g38) & (g39) & (!g40) & (!g43)) + ((!a) & (g11) & (!g38) & (g39) & (!g40) & (g43)) + ((!a) & (g11) & (!g38) & (g39) & (g40) & (!g43)) + ((!a) & (g11) & (!g38) & (g39) & (g40) & (g43)) + ((!a) & (g11) & (g38) & (!g39) & (!g40) & (g43)) + ((!a) & (g11) & (g38) & (!g39) & (g40) & (!g43)) + ((!a) & (g11) & (g38) & (!g39) & (g40) & (g43)) + ((!a) & (g11) & (g38) & (g39) & (!g40) & (!g43)) + ((!a) & (g11) & (g38) & (g39) & (!g40) & (g43)) + ((!a) & (g11) & (g38) & (g39) & (g40) & (!g43)) + ((!a) & (g11) & (g38) & (g39) & (g40) & (g43)) + ((a) & (!g11) & (!g38) & (!g39) & (!g40) & (g43)) + ((a) & (!g11) & (!g38) & (!g39) & (g40) & (!g43)) + ((a) & (!g11) & (!g38) & (!g39) & (g40) & (g43)) + ((a) & (!g11) & (!g38) & (g39) & (!g40) & (g43)) + ((a) & (!g11) & (!g38) & (g39) & (g40) & (!g43)) + ((a) & (!g11) & (!g38) & (g39) & (g40) & (g43)) + ((a) & (!g11) & (g38) & (!g39) & (!g40) & (!g43)) + ((a) & (!g11) & (g38) & (!g39) & (!g40) & (g43)) + ((a) & (!g11) & (g38) & (!g39) & (g40) & (!g43)) + ((a) & (!g11) & (g38) & (!g39) & (g40) & (g43)) + ((a) & (!g11) & (g38) & (g39) & (!g40) & (!g43)) + ((a) & (!g11) & (g38) & (g39) & (!g40) & (g43)) + ((a) & (!g11) & (g38) & (g39) & (g40) & (!g43)) + ((a) & (!g11) & (g38) & (g39) & (g40) & (g43)) + ((a) & (g11) & (!g38) & (!g39) & (!g40) & (g43)) + ((a) & (g11) & (!g38) & (!g39) & (g40) & (!g43)) + ((a) & (g11) & (!g38) & (!g39) & (g40) & (g43)) + ((a) & (g11) & (!g38) & (g39) & (!g40) & (!g43)) + ((a) & (g11) & (!g38) & (g39) & (!g40) & (g43)) + ((a) & (g11) & (!g38) & (g39) & (g40) & (!g43)) + ((a) & (g11) & (!g38) & (g39) & (g40) & (g43)) + ((a) & (g11) & (g38) & (!g39) & (!g40) & (!g43)) + ((a) & (g11) & (g38) & (!g39) & (!g40) & (g43)) + ((a) & (g11) & (g38) & (!g39) & (g40) & (!g43)) + ((a) & (g11) & (g38) & (!g39) & (g40) & (g43)) + ((a) & (g11) & (g38) & (g39) & (!g40) & (!g43)) + ((a) & (g11) & (g38) & (g39) & (!g40) & (g43)) + ((a) & (g11) & (g38) & (g39) & (g40) & (!g43)) + ((a) & (g11) & (g38) & (g39) & (g40) & (g43)));
	assign g182 = (((!sk[0]) & (!g180) & (!g181) & (i)) + ((!sk[0]) & (!g180) & (g181) & (i)) + ((!sk[0]) & (g180) & (!g181) & (i)) + ((!sk[0]) & (g180) & (g181) & (i)) + ((sk[0]) & (!g180) & (g181) & (i)) + ((sk[0]) & (g180) & (!g181) & (!i)) + ((sk[0]) & (g180) & (g181) & (!i)) + ((sk[0]) & (g180) & (g181) & (i)));
	assign g141 = (((!sk[0]) & (!g124) & (g132)) + ((!sk[0]) & (g124) & (g132)) + ((sk[0]) & (!g124) & (g132)));
	assign g46 = (((!g9) & (!g10) & (!g12) & (!b) & (!g44) & (!g45)) + ((!g9) & (!g10) & (!g12) & (!b) & (!g44) & (g45)) + ((!g9) & (!g10) & (!g12) & (!b) & (g44) & (!g45)) + ((!g9) & (!g10) & (!g12) & (!b) & (g44) & (g45)) + ((!g9) & (!g10) & (!g12) & (b) & (!g44) & (!g45)) + ((!g9) & (!g10) & (!g12) & (b) & (g44) & (!g45)) + ((!g9) & (!g10) & (g12) & (!b) & (!g44) & (!g45)) + ((!g9) & (!g10) & (g12) & (!b) & (!g44) & (g45)) + ((!g9) & (g10) & (!g12) & (!b) & (g44) & (!g45)) + ((!g9) & (g10) & (!g12) & (!b) & (g44) & (g45)) + ((!g9) & (g10) & (!g12) & (b) & (g44) & (!g45)) + ((g9) & (!g10) & (!g12) & (!b) & (!g44) & (!g45)) + ((g9) & (!g10) & (!g12) & (!b) & (!g44) & (g45)) + ((g9) & (!g10) & (!g12) & (!b) & (g44) & (!g45)) + ((g9) & (!g10) & (!g12) & (!b) & (g44) & (g45)) + ((g9) & (!g10) & (!g12) & (b) & (!g44) & (!g45)) + ((g9) & (!g10) & (g12) & (!b) & (!g44) & (!g45)) + ((g9) & (!g10) & (g12) & (!b) & (!g44) & (g45)) + ((g9) & (g10) & (!g12) & (!b) & (g44) & (!g45)) + ((g9) & (g10) & (!g12) & (!b) & (g44) & (g45)));
	assign g1 = (((k) & (!sk[1]) & (!l)) + ((k) & (sk[1]) & (!l)) + ((k) & (sk[1]) & (l)));
	assign g14 = (((!a) & (!sk[2]) & (!e) & (!g7) & (g13)) + ((!a) & (!sk[2]) & (!e) & (g7) & (g13)) + ((!a) & (!sk[2]) & (e) & (!g7) & (!g13)) + ((!a) & (!sk[2]) & (e) & (!g7) & (g13)) + ((!a) & (!sk[2]) & (e) & (g7) & (!g13)) + ((!a) & (!sk[2]) & (e) & (g7) & (g13)) + ((!a) & (sk[2]) & (!e) & (!g7) & (g13)) + ((!a) & (sk[2]) & (!e) & (g7) & (g13)) + ((!a) & (sk[2]) & (e) & (!g7) & (g13)) + ((!a) & (sk[2]) & (e) & (g7) & (g13)) + ((a) & (!sk[2]) & (!e) & (!g7) & (g13)) + ((a) & (!sk[2]) & (!e) & (g7) & (g13)) + ((a) & (!sk[2]) & (e) & (!g7) & (!g13)) + ((a) & (!sk[2]) & (e) & (!g7) & (g13)) + ((a) & (!sk[2]) & (e) & (g7) & (!g13)) + ((a) & (!sk[2]) & (e) & (g7) & (g13)) + ((a) & (sk[2]) & (!e) & (!g7) & (g13)) + ((a) & (sk[2]) & (!e) & (g7) & (g13)) + ((a) & (sk[2]) & (e) & (!g7) & (g13)));
	assign g12 = (((!sk[3]) & (l) & (!g11)) + ((!sk[3]) & (l) & (g11)) + ((sk[3]) & (l) & (g11)));
	assign g90 = (((!g10) & (!sk[0]) & (!g82) & (!g87) & (g88) & (!g89)) + ((!g10) & (!sk[0]) & (!g82) & (!g87) & (g88) & (g89)) + ((!g10) & (!sk[0]) & (!g82) & (g87) & (g88) & (!g89)) + ((!g10) & (!sk[0]) & (!g82) & (g87) & (g88) & (g89)) + ((!g10) & (!sk[0]) & (g82) & (!g87) & (!g88) & (!g89)) + ((!g10) & (!sk[0]) & (g82) & (!g87) & (!g88) & (g89)) + ((!g10) & (!sk[0]) & (g82) & (!g87) & (g88) & (!g89)) + ((!g10) & (!sk[0]) & (g82) & (!g87) & (g88) & (g89)) + ((!g10) & (!sk[0]) & (g82) & (g87) & (!g88) & (!g89)) + ((!g10) & (!sk[0]) & (g82) & (g87) & (!g88) & (g89)) + ((!g10) & (!sk[0]) & (g82) & (g87) & (g88) & (!g89)) + ((!g10) & (!sk[0]) & (g82) & (g87) & (g88) & (g89)) + ((!g10) & (sk[0]) & (!g82) & (!g87) & (g88) & (!g89)) + ((!g10) & (sk[0]) & (!g82) & (g87) & (!g88) & (!g89)) + ((!g10) & (sk[0]) & (!g82) & (g87) & (g88) & (!g89)) + ((!g10) & (sk[0]) & (g82) & (!g87) & (g88) & (!g89)) + ((!g10) & (sk[0]) & (g82) & (g87) & (g88) & (!g89)) + ((g10) & (!sk[0]) & (!g82) & (!g87) & (g88) & (!g89)) + ((g10) & (!sk[0]) & (!g82) & (!g87) & (g88) & (g89)) + ((g10) & (!sk[0]) & (!g82) & (g87) & (g88) & (!g89)) + ((g10) & (!sk[0]) & (!g82) & (g87) & (g88) & (g89)) + ((g10) & (!sk[0]) & (g82) & (!g87) & (!g88) & (!g89)) + ((g10) & (!sk[0]) & (g82) & (!g87) & (!g88) & (g89)) + ((g10) & (!sk[0]) & (g82) & (!g87) & (g88) & (!g89)) + ((g10) & (!sk[0]) & (g82) & (!g87) & (g88) & (g89)) + ((g10) & (!sk[0]) & (g82) & (g87) & (!g88) & (!g89)) + ((g10) & (!sk[0]) & (g82) & (g87) & (!g88) & (g89)) + ((g10) & (!sk[0]) & (g82) & (g87) & (g88) & (!g89)) + ((g10) & (!sk[0]) & (g82) & (g87) & (g88) & (g89)) + ((g10) & (sk[0]) & (!g82) & (!g87) & (g88) & (!g89)) + ((g10) & (sk[0]) & (g82) & (!g87) & (g88) & (!g89)) + ((g10) & (sk[0]) & (g82) & (g87) & (g88) & (!g89)));
	assign g135 = (((!sk[4]) & (!g10) & (!g124) & (!g132) & (g133) & (!g134)) + ((!sk[4]) & (!g10) & (!g124) & (g132) & (!g133) & (!g134)) + ((!sk[4]) & (!g10) & (!g124) & (g132) & (g133) & (!g134)) + ((!sk[4]) & (!g10) & (g124) & (!g132) & (g133) & (!g134)) + ((!sk[4]) & (!g10) & (g124) & (g132) & (g133) & (!g134)) + ((!sk[4]) & (g10) & (!g124) & (!g132) & (g133) & (!g134)) + ((!sk[4]) & (g10) & (g124) & (!g132) & (g133) & (!g134)) + ((!sk[4]) & (g10) & (g124) & (g132) & (g133) & (!g134)) + ((sk[4]) & (!g10) & (!g124) & (!g132) & (!g133) & (g134)) + ((sk[4]) & (!g10) & (!g124) & (!g132) & (g133) & (!g134)) + ((sk[4]) & (!g10) & (!g124) & (!g132) & (g133) & (g134)) + ((sk[4]) & (!g10) & (!g124) & (g132) & (!g133) & (g134)) + ((sk[4]) & (!g10) & (!g124) & (g132) & (g133) & (!g134)) + ((sk[4]) & (!g10) & (!g124) & (g132) & (g133) & (g134)) + ((sk[4]) & (!g10) & (g124) & (!g132) & (!g133) & (g134)) + ((sk[4]) & (!g10) & (g124) & (!g132) & (g133) & (!g134)) + ((sk[4]) & (!g10) & (g124) & (!g132) & (g133) & (g134)) + ((sk[4]) & (!g10) & (g124) & (g132) & (!g133) & (g134)) + ((sk[4]) & (!g10) & (g124) & (g132) & (g133) & (!g134)) + ((sk[4]) & (!g10) & (g124) & (g132) & (g133) & (g134)) + ((sk[4]) & (g10) & (!g124) & (!g132) & (!g133) & (!g134)) + ((sk[4]) & (g10) & (!g124) & (!g132) & (!g133) & (g134)) + ((sk[4]) & (g10) & (!g124) & (!g132) & (g133) & (!g134)) + ((sk[4]) & (g10) & (!g124) & (!g132) & (g133) & (g134)) + ((sk[4]) & (g10) & (!g124) & (g132) & (!g133) & (!g134)) + ((sk[4]) & (g10) & (!g124) & (g132) & (!g133) & (g134)) + ((sk[4]) & (g10) & (!g124) & (g132) & (g133) & (!g134)) + ((sk[4]) & (g10) & (!g124) & (g132) & (g133) & (g134)) + ((sk[4]) & (g10) & (g124) & (!g132) & (!g133) & (!g134)) + ((sk[4]) & (g10) & (g124) & (!g132) & (!g133) & (g134)) + ((sk[4]) & (g10) & (g124) & (!g132) & (g133) & (!g134)) + ((sk[4]) & (g10) & (g124) & (!g132) & (g133) & (g134)) + ((sk[4]) & (g10) & (g124) & (g132) & (!g133) & (!g134)) + ((sk[4]) & (g10) & (g124) & (g132) & (!g133) & (g134)) + ((sk[4]) & (g10) & (g124) & (g132) & (g133) & (!g134)) + ((sk[4]) & (g10) & (g124) & (g132) & (g133) & (g134)));
	assign g8 = (((!sk[4]) & (i) & (j)) + ((sk[4]) & (!i) & (j)) + ((sk[4]) & (i) & (j)));
	assign g15 = (((!k) & (!sk[4]) & (g12)) + ((!k) & (sk[4]) & (g12)) + ((k) & (sk[4]) & (g12)));
	assign g92 = (((!g50) & (!b) & (sk[4]) & (g44)) + ((!g50) & (b) & (!sk[4]) & (g44)) + ((!g50) & (b) & (sk[4]) & (g44)) + ((g50) & (!b) & (!sk[4]) & (g44)) + ((g50) & (!b) & (sk[4]) & (g44)) + ((g50) & (b) & (!sk[4]) & (!g44)) + ((g50) & (b) & (!sk[4]) & (g44)) + ((g50) & (b) & (sk[4]) & (g44)));
	assign g103 = (((!g7) & (!sk[5]) & (!g90) & (!g102)) + ((!g7) & (!sk[5]) & (g90) & (!g102)) + ((g7) & (!sk[5]) & (!g90) & (!g102)));
	assign g11 = (((!sk[6]) & (n) & (!i) & (!j)) + ((!sk[6]) & (n) & (!i) & (j)) + ((!sk[6]) & (n) & (i) & (!j)) + ((!sk[6]) & (n) & (i) & (j)) + ((sk[6]) & (n) & (!i) & (j)));
	assign g47 = (((!g15) & (!sk[7]) & (!f) & (b)) + ((!g15) & (!sk[7]) & (f) & (b)) + ((g15) & (!sk[7]) & (!f) & (!b)) + ((g15) & (!sk[7]) & (!f) & (b)) + ((g15) & (!sk[7]) & (f) & (!b)) + ((g15) & (!sk[7]) & (f) & (b)) + ((g15) & (sk[7]) & (f) & (b)));
	assign g51 = (((!k) & (!l) & (sk[1]) & (!i) & (j)) + ((!k) & (!l) & (sk[1]) & (i) & (j)) + ((!k) & (l) & (!sk[1]) & (!i) & (!j)) + ((!k) & (l) & (sk[1]) & (!i) & (j)) + ((!k) & (l) & (sk[1]) & (i) & (j)) + ((k) & (!l) & (sk[1]) & (!i) & (j)) + ((k) & (!l) & (sk[1]) & (i) & (j)) + ((k) & (l) & (!sk[1]) & (!i) & (!j)) + ((k) & (l) & (!sk[1]) & (!i) & (j)) + ((k) & (l) & (!sk[1]) & (i) & (!j)) + ((k) & (l) & (sk[1]) & (!i) & (!j)) + ((k) & (l) & (sk[1]) & (!i) & (j)) + ((k) & (l) & (sk[1]) & (i) & (!j)) + ((k) & (l) & (sk[1]) & (i) & (j)));
	assign g53 = (((!sk[1]) & (!k) & (!l) & (!i) & (!j)) + ((!sk[1]) & (!k) & (l) & (!i) & (!j)) + ((!sk[1]) & (k) & (l) & (!i) & (!j)) + ((!sk[1]) & (k) & (l) & (!i) & (j)) + ((!sk[1]) & (k) & (l) & (i) & (!j)));
	assign g60 = (((!k) & (!sk[8]) & (n) & (!g8)) + ((!k) & (!sk[8]) & (n) & (g8)) + ((k) & (!sk[8]) & (!n) & (g8)) + ((k) & (!sk[8]) & (n) & (!g8)) + ((k) & (!sk[8]) & (n) & (g8)) + ((k) & (sk[8]) & (n) & (g8)));
	assign g121 = (((!d) & (sk[9]) & (h)) + ((d) & (!sk[9]) & (h)) + ((d) & (sk[9]) & (h)));
	assign g138 = (((!g7) & (!g15) & (sk[5]) & (g121) & (!g135)) + ((!g7) & (!g15) & (sk[5]) & (g121) & (g135)) + ((!g7) & (g15) & (!sk[5]) & (g121) & (!g135)) + ((!g7) & (g15) & (!sk[5]) & (g121) & (g135)) + ((!g7) & (g15) & (sk[5]) & (g121) & (!g135)) + ((!g7) & (g15) & (sk[5]) & (g121) & (g135)) + ((g7) & (!g15) & (!sk[5]) & (!g121) & (g135)) + ((g7) & (!g15) & (!sk[5]) & (g121) & (g135)) + ((g7) & (!g15) & (sk[5]) & (!g121) & (g135)) + ((g7) & (!g15) & (sk[5]) & (g121) & (!g135)) + ((g7) & (!g15) & (sk[5]) & (g121) & (g135)) + ((g7) & (g15) & (!sk[5]) & (!g121) & (g135)) + ((g7) & (g15) & (!sk[5]) & (g121) & (!g135)) + ((g7) & (g15) & (!sk[5]) & (g121) & (g135)) + ((g7) & (g15) & (sk[5]) & (!g121) & (g135)) + ((g7) & (g15) & (sk[5]) & (g121) & (!g135)) + ((g7) & (g15) & (sk[5]) & (g121) & (g135)));
	assign g9 = (((!n) & (!g8) & (!sk[8]) & (g1)) + ((!n) & (g8) & (!sk[8]) & (g1)) + ((n) & (!g8) & (!sk[8]) & (g1)) + ((n) & (g8) & (!sk[8]) & (g1)) + ((n) & (g8) & (sk[8]) & (g1)));
	assign g10 = (((!n) & (!i) & (!sk[6]) & (j) & (!g1)) + ((!n) & (!i) & (!sk[6]) & (j) & (g1)) + ((!n) & (i) & (!sk[6]) & (!j) & (!g1)) + ((!n) & (i) & (!sk[6]) & (!j) & (g1)) + ((!n) & (i) & (!sk[6]) & (j) & (!g1)) + ((!n) & (i) & (!sk[6]) & (j) & (g1)) + ((n) & (!i) & (!sk[6]) & (!j) & (!g1)) + ((n) & (!i) & (!sk[6]) & (!j) & (g1)) + ((n) & (!i) & (!sk[6]) & (j) & (!g1)) + ((n) & (!i) & (!sk[6]) & (j) & (g1)) + ((n) & (!i) & (sk[6]) & (!j) & (g1)) + ((n) & (i) & (!sk[6]) & (!j) & (!g1)) + ((n) & (i) & (!sk[6]) & (!j) & (g1)) + ((n) & (i) & (!sk[6]) & (j) & (!g1)) + ((n) & (i) & (!sk[6]) & (j) & (g1)));
	assign g16 = (((!a) & (!e) & (!g7) & (!sk[2]) & (!g13) & (g15)) + ((!a) & (!e) & (!g7) & (!sk[2]) & (g13) & (g15)) + ((!a) & (!e) & (g7) & (!sk[2]) & (!g13) & (g15)) + ((!a) & (!e) & (g7) & (!sk[2]) & (g13) & (g15)) + ((!a) & (!e) & (g7) & (sk[2]) & (g13) & (!g15)) + ((!a) & (!e) & (g7) & (sk[2]) & (g13) & (g15)) + ((!a) & (e) & (!g7) & (!sk[2]) & (!g13) & (!g15)) + ((!a) & (e) & (!g7) & (!sk[2]) & (!g13) & (g15)) + ((!a) & (e) & (!g7) & (!sk[2]) & (g13) & (!g15)) + ((!a) & (e) & (!g7) & (!sk[2]) & (g13) & (g15)) + ((!a) & (e) & (g7) & (!sk[2]) & (!g13) & (!g15)) + ((!a) & (e) & (g7) & (!sk[2]) & (!g13) & (g15)) + ((!a) & (e) & (g7) & (!sk[2]) & (g13) & (!g15)) + ((!a) & (e) & (g7) & (!sk[2]) & (g13) & (g15)) + ((!a) & (e) & (g7) & (sk[2]) & (g13) & (!g15)) + ((!a) & (e) & (g7) & (sk[2]) & (g13) & (g15)) + ((a) & (!e) & (!g7) & (!sk[2]) & (!g13) & (g15)) + ((a) & (!e) & (!g7) & (!sk[2]) & (g13) & (g15)) + ((a) & (!e) & (g7) & (!sk[2]) & (!g13) & (g15)) + ((a) & (!e) & (g7) & (!sk[2]) & (g13) & (g15)) + ((a) & (!e) & (g7) & (sk[2]) & (g13) & (!g15)) + ((a) & (!e) & (g7) & (sk[2]) & (g13) & (g15)) + ((a) & (e) & (!g7) & (!sk[2]) & (!g13) & (!g15)) + ((a) & (e) & (!g7) & (!sk[2]) & (!g13) & (g15)) + ((a) & (e) & (!g7) & (!sk[2]) & (g13) & (!g15)) + ((a) & (e) & (!g7) & (!sk[2]) & (g13) & (g15)) + ((a) & (e) & (!g7) & (sk[2]) & (!g13) & (g15)) + ((a) & (e) & (!g7) & (sk[2]) & (g13) & (g15)) + ((a) & (e) & (g7) & (!sk[2]) & (!g13) & (!g15)) + ((a) & (e) & (g7) & (!sk[2]) & (!g13) & (g15)) + ((a) & (e) & (g7) & (!sk[2]) & (g13) & (!g15)) + ((a) & (e) & (g7) & (!sk[2]) & (g13) & (g15)) + ((a) & (e) & (g7) & (sk[2]) & (!g13) & (g15)) + ((a) & (e) & (g7) & (sk[2]) & (g13) & (g15)));
	assign g22 = (((!l) & (!n) & (!sk[3]) & (j)) + ((!l) & (n) & (!sk[3]) & (j)) + ((!l) & (n) & (sk[3]) & (!j)) + ((l) & (!n) & (!sk[3]) & (!j)) + ((l) & (!n) & (!sk[3]) & (j)) + ((l) & (n) & (!sk[3]) & (!j)) + ((l) & (n) & (!sk[3]) & (j)));
	assign g26 = (((!sk[10]) & (i) & (!g22)) + ((!sk[10]) & (i) & (g22)) + ((sk[10]) & (!i) & (g22)));
	assign g31 = (((!n) & (!g21) & (!g24) & (!sk[11]) & (!g25) & (!g30)) + ((!n) & (!g21) & (!g24) & (!sk[11]) & (g25) & (!g30)) + ((!n) & (!g21) & (!g24) & (!sk[11]) & (g25) & (g30)) + ((!n) & (!g21) & (g24) & (!sk[11]) & (!g25) & (!g30)) + ((!n) & (!g21) & (g24) & (!sk[11]) & (!g25) & (g30)) + ((!n) & (!g21) & (g24) & (!sk[11]) & (g25) & (!g30)) + ((!n) & (!g21) & (g24) & (!sk[11]) & (g25) & (g30)) + ((!n) & (g21) & (!g24) & (!sk[11]) & (!g25) & (!g30)) + ((!n) & (g21) & (!g24) & (!sk[11]) & (g25) & (!g30)) + ((!n) & (g21) & (!g24) & (!sk[11]) & (g25) & (g30)) + ((!n) & (g21) & (g24) & (!sk[11]) & (!g25) & (!g30)) + ((!n) & (g21) & (g24) & (!sk[11]) & (!g25) & (g30)) + ((!n) & (g21) & (g24) & (!sk[11]) & (g25) & (!g30)) + ((!n) & (g21) & (g24) & (!sk[11]) & (g25) & (g30)) + ((n) & (!g21) & (!g24) & (!sk[11]) & (!g25) & (!g30)) + ((n) & (!g21) & (!g24) & (!sk[11]) & (!g25) & (g30)) + ((n) & (!g21) & (!g24) & (!sk[11]) & (g25) & (!g30)) + ((n) & (!g21) & (!g24) & (!sk[11]) & (g25) & (g30)) + ((n) & (!g21) & (g24) & (!sk[11]) & (!g25) & (!g30)) + ((n) & (!g21) & (g24) & (!sk[11]) & (!g25) & (g30)) + ((n) & (!g21) & (g24) & (!sk[11]) & (g25) & (!g30)) + ((n) & (!g21) & (g24) & (!sk[11]) & (g25) & (g30)) + ((n) & (g21) & (!g24) & (!sk[11]) & (!g25) & (!g30)) + ((n) & (g21) & (!g24) & (!sk[11]) & (g25) & (!g30)) + ((n) & (g21) & (!g24) & (!sk[11]) & (g25) & (g30)) + ((n) & (g21) & (g24) & (!sk[11]) & (!g25) & (!g30)) + ((n) & (g21) & (g24) & (!sk[11]) & (!g25) & (g30)) + ((n) & (g21) & (g24) & (!sk[11]) & (g25) & (!g30)) + ((n) & (g21) & (g24) & (!sk[11]) & (g25) & (g30)));
	assign g32 = (((!k) & (!sk[8]) & (n) & (!i)) + ((!k) & (!sk[8]) & (n) & (i)) + ((!k) & (sk[8]) & (!n) & (!i)) + ((k) & (!sk[8]) & (!n) & (!i)) + ((k) & (!sk[8]) & (!n) & (i)) + ((k) & (!sk[8]) & (n) & (!i)) + ((k) & (!sk[8]) & (n) & (i)));
	assign g33 = (((!k) & (!l) & (!n) & (sk[1]) & (!i) & (j)) + ((!k) & (!l) & (!n) & (sk[1]) & (i) & (j)) + ((!k) & (!l) & (n) & (!sk[1]) & (i) & (j)) + ((!k) & (!l) & (n) & (sk[1]) & (!i) & (!j)) + ((!k) & (!l) & (n) & (sk[1]) & (!i) & (j)) + ((!k) & (!l) & (n) & (sk[1]) & (i) & (!j)) + ((!k) & (!l) & (n) & (sk[1]) & (i) & (j)) + ((!k) & (l) & (!n) & (sk[1]) & (!i) & (j)) + ((!k) & (l) & (!n) & (sk[1]) & (i) & (j)) + ((!k) & (l) & (n) & (sk[1]) & (!i) & (!j)) + ((!k) & (l) & (n) & (sk[1]) & (!i) & (j)) + ((!k) & (l) & (n) & (sk[1]) & (i) & (!j)) + ((!k) & (l) & (n) & (sk[1]) & (i) & (j)) + ((k) & (!l) & (!n) & (sk[1]) & (!i) & (j)) + ((k) & (!l) & (!n) & (sk[1]) & (i) & (j)) + ((k) & (!l) & (n) & (sk[1]) & (!i) & (!j)) + ((k) & (!l) & (n) & (sk[1]) & (!i) & (j)) + ((k) & (!l) & (n) & (sk[1]) & (i) & (!j)) + ((k) & (!l) & (n) & (sk[1]) & (i) & (j)) + ((k) & (l) & (!n) & (!sk[1]) & (!i) & (!j)) + ((k) & (l) & (!n) & (sk[1]) & (!i) & (j)) + ((k) & (l) & (!n) & (sk[1]) & (i) & (j)) + ((k) & (l) & (n) & (sk[1]) & (!i) & (!j)) + ((k) & (l) & (n) & (sk[1]) & (!i) & (j)) + ((k) & (l) & (n) & (sk[1]) & (i) & (!j)) + ((k) & (l) & (n) & (sk[1]) & (i) & (j)));
	assign g34 = (((!sk[1]) & (!k) & (l) & (!n) & (!i) & (j)) + ((!sk[1]) & (!k) & (l) & (!n) & (i) & (j)) + ((!sk[1]) & (k) & (!l) & (!n) & (!i) & (j)) + ((!sk[1]) & (k) & (l) & (!n) & (!i) & (j)) + ((!sk[1]) & (k) & (l) & (!n) & (i) & (j)) + ((sk[1]) & (!k) & (!l) & (!n) & (i) & (!j)) + ((sk[1]) & (!k) & (!l) & (!n) & (i) & (j)) + ((sk[1]) & (!k) & (!l) & (n) & (!i) & (!j)) + ((sk[1]) & (!k) & (!l) & (n) & (!i) & (j)) + ((sk[1]) & (!k) & (!l) & (n) & (i) & (!j)) + ((sk[1]) & (!k) & (!l) & (n) & (i) & (j)) + ((sk[1]) & (!k) & (l) & (!n) & (!i) & (j)) + ((sk[1]) & (!k) & (l) & (!n) & (i) & (!j)) + ((sk[1]) & (!k) & (l) & (!n) & (i) & (j)) + ((sk[1]) & (!k) & (l) & (n) & (!i) & (!j)) + ((sk[1]) & (!k) & (l) & (n) & (!i) & (j)) + ((sk[1]) & (!k) & (l) & (n) & (i) & (!j)) + ((sk[1]) & (!k) & (l) & (n) & (i) & (j)) + ((sk[1]) & (k) & (!l) & (!n) & (i) & (!j)) + ((sk[1]) & (k) & (!l) & (!n) & (i) & (j)) + ((sk[1]) & (k) & (!l) & (n) & (!i) & (!j)) + ((sk[1]) & (k) & (!l) & (n) & (!i) & (j)) + ((sk[1]) & (k) & (!l) & (n) & (i) & (!j)) + ((sk[1]) & (k) & (!l) & (n) & (i) & (j)) + ((sk[1]) & (k) & (l) & (!n) & (!i) & (!j)) + ((sk[1]) & (k) & (l) & (!n) & (!i) & (j)) + ((sk[1]) & (k) & (l) & (!n) & (i) & (!j)) + ((sk[1]) & (k) & (l) & (!n) & (i) & (j)) + ((sk[1]) & (k) & (l) & (n) & (!i) & (!j)) + ((sk[1]) & (k) & (l) & (n) & (!i) & (j)) + ((sk[1]) & (k) & (l) & (n) & (i) & (!j)) + ((sk[1]) & (k) & (l) & (n) & (i) & (j)));
	assign g35 = (((!sk[3]) & (!k) & (!l) & (!n) & (i) & (!j)) + ((!sk[3]) & (!k) & (!l) & (!n) & (i) & (j)) + ((!sk[3]) & (!k) & (!l) & (n) & (!i) & (!j)) + ((!sk[3]) & (!k) & (!l) & (n) & (!i) & (j)) + ((!sk[3]) & (!k) & (!l) & (n) & (i) & (!j)) + ((!sk[3]) & (!k) & (!l) & (n) & (i) & (j)) + ((!sk[3]) & (!k) & (l) & (!n) & (!i) & (!j)) + ((!sk[3]) & (!k) & (l) & (!n) & (!i) & (j)) + ((!sk[3]) & (!k) & (l) & (!n) & (i) & (!j)) + ((!sk[3]) & (!k) & (l) & (!n) & (i) & (j)) + ((!sk[3]) & (!k) & (l) & (n) & (!i) & (!j)) + ((!sk[3]) & (!k) & (l) & (n) & (!i) & (j)) + ((!sk[3]) & (!k) & (l) & (n) & (i) & (!j)) + ((!sk[3]) & (!k) & (l) & (n) & (i) & (j)) + ((!sk[3]) & (k) & (!l) & (!n) & (i) & (!j)) + ((!sk[3]) & (k) & (!l) & (!n) & (i) & (j)) + ((!sk[3]) & (k) & (!l) & (n) & (!i) & (!j)) + ((!sk[3]) & (k) & (!l) & (n) & (!i) & (j)) + ((!sk[3]) & (k) & (!l) & (n) & (i) & (!j)) + ((!sk[3]) & (k) & (!l) & (n) & (i) & (j)) + ((!sk[3]) & (k) & (l) & (!n) & (!i) & (!j)) + ((!sk[3]) & (k) & (l) & (!n) & (!i) & (j)) + ((!sk[3]) & (k) & (l) & (!n) & (i) & (!j)) + ((!sk[3]) & (k) & (l) & (!n) & (i) & (j)) + ((!sk[3]) & (k) & (l) & (n) & (!i) & (!j)) + ((!sk[3]) & (k) & (l) & (n) & (!i) & (j)) + ((!sk[3]) & (k) & (l) & (n) & (i) & (!j)) + ((!sk[3]) & (k) & (l) & (n) & (i) & (j)) + ((sk[3]) & (!k) & (l) & (!n) & (!i) & (!j)) + ((sk[3]) & (k) & (l) & (!n) & (!i) & (!j)) + ((sk[3]) & (k) & (l) & (!n) & (!i) & (j)) + ((sk[3]) & (k) & (l) & (!n) & (i) & (!j)) + ((sk[3]) & (k) & (l) & (!n) & (i) & (j)));
	assign g37 = (((!e) & (!g32) & (!sk[12]) & (!g182) & (!g36)) + ((!e) & (!g32) & (!sk[12]) & (g182) & (!g36)) + ((!e) & (g32) & (!sk[12]) & (!g182) & (!g36)) + ((!e) & (g32) & (!sk[12]) & (g182) & (!g36)) + ((e) & (!g32) & (!sk[12]) & (!g182) & (!g36)) + ((e) & (!g32) & (!sk[12]) & (g182) & (!g36)) + ((e) & (g32) & (!sk[12]) & (!g182) & (!g36)) + ((e) & (g32) & (!sk[12]) & (g182) & (!g36)) + ((e) & (g32) & (!sk[12]) & (g182) & (g36)));
	assign g50 = (((a) & (!sk[12]) & (g182)) + ((a) & (sk[12]) & (!g182)) + ((a) & (sk[12]) & (g182)));
	assign g56 = (((!sk[12]) & (!g182) & (g54) & (!g55)) + ((!sk[12]) & (!g182) & (g54) & (g55)) + ((!sk[12]) & (g182) & (!g54) & (g55)) + ((!sk[12]) & (g182) & (g54) & (!g55)) + ((!sk[12]) & (g182) & (g54) & (g55)) + ((sk[12]) & (!g182) & (!g54) & (g55)) + ((sk[12]) & (!g182) & (g54) & (g55)) + ((sk[12]) & (g182) & (!g54) & (!g55)) + ((sk[12]) & (g182) & (!g54) & (g55)) + ((sk[12]) & (g182) & (g54) & (!g55)) + ((sk[12]) & (g182) & (g54) & (g55)));
	assign g57 = (((!k) & (sk[3]) & (!l) & (!g8)) + ((k) & (!sk[3]) & (!l) & (!g8)) + ((k) & (!sk[3]) & (!l) & (g8)) + ((k) & (!sk[3]) & (l) & (!g8)) + ((k) & (!sk[3]) & (l) & (g8)));
	assign g62 = (((!sk[12]) & (!g182) & (!g44)));
	assign g65 = (((!k) & (!sk[6]) & (n) & (!i) & (!j)) + ((!k) & (!sk[6]) & (n) & (!i) & (j)) + ((!k) & (!sk[6]) & (n) & (i) & (!j)) + ((!k) & (!sk[6]) & (n) & (i) & (j)) + ((!k) & (sk[6]) & (n) & (i) & (!j)) + ((k) & (!sk[6]) & (!n) & (!i) & (!j)) + ((k) & (!sk[6]) & (!n) & (!i) & (j)) + ((k) & (!sk[6]) & (!n) & (i) & (!j)) + ((k) & (!sk[6]) & (!n) & (i) & (j)) + ((k) & (!sk[6]) & (n) & (!i) & (!j)) + ((k) & (!sk[6]) & (n) & (!i) & (j)) + ((k) & (!sk[6]) & (n) & (i) & (!j)) + ((k) & (!sk[6]) & (n) & (i) & (j)));
	assign g80 = (((!m) & (!sk[13]) & (!g31) & (!g58) & (!g59) & (!g72)) + ((!m) & (!sk[13]) & (!g31) & (!g58) & (!g59) & (g72)) + ((!m) & (!sk[13]) & (!g31) & (!g58) & (g59) & (!g72)) + ((!m) & (!sk[13]) & (!g31) & (!g58) & (g59) & (g72)) + ((!m) & (!sk[13]) & (!g31) & (g58) & (!g59) & (!g72)) + ((!m) & (!sk[13]) & (!g31) & (g58) & (!g59) & (g72)) + ((!m) & (!sk[13]) & (!g31) & (g58) & (g59) & (!g72)) + ((!m) & (!sk[13]) & (!g31) & (g58) & (g59) & (g72)) + ((!m) & (!sk[13]) & (g31) & (!g58) & (!g59) & (g72)) + ((m) & (!sk[13]) & (!g31) & (!g58) & (!g59) & (!g72)) + ((m) & (!sk[13]) & (!g31) & (!g58) & (!g59) & (g72)) + ((m) & (!sk[13]) & (!g31) & (!g58) & (g59) & (!g72)) + ((m) & (!sk[13]) & (!g31) & (!g58) & (g59) & (g72)) + ((m) & (!sk[13]) & (!g31) & (g58) & (!g59) & (!g72)) + ((m) & (!sk[13]) & (!g31) & (g58) & (!g59) & (g72)) + ((m) & (!sk[13]) & (!g31) & (g58) & (g59) & (!g72)) + ((m) & (!sk[13]) & (!g31) & (g58) & (g59) & (g72)) + ((m) & (!sk[13]) & (g31) & (!g58) & (!g59) & (!g72)) + ((m) & (!sk[13]) & (g31) & (!g58) & (!g59) & (g72)) + ((m) & (!sk[13]) & (g31) & (!g58) & (g59) & (!g72)) + ((m) & (!sk[13]) & (g31) & (!g58) & (g59) & (g72)) + ((m) & (!sk[13]) & (g31) & (g58) & (!g59) & (!g72)) + ((m) & (!sk[13]) & (g31) & (g58) & (!g59) & (g72)) + ((m) & (!sk[13]) & (g31) & (g58) & (g59) & (!g72)) + ((m) & (!sk[13]) & (g31) & (g58) & (g59) & (g72)));
	assign g104 = (((!g182) & (!g7) & (!g16) & (g44) & (!g46) & (g47)) + ((!g182) & (!g7) & (!g16) & (g44) & (g46) & (g47)) + ((!g182) & (!g7) & (g16) & (g44) & (!g46) & (g47)) + ((!g182) & (!g7) & (g16) & (g44) & (g46) & (g47)) + ((!g182) & (g7) & (!g16) & (g44) & (!g46) & (g47)) + ((!g182) & (g7) & (!g16) & (g44) & (g46) & (!g47)) + ((!g182) & (g7) & (!g16) & (g44) & (g46) & (g47)) + ((!g182) & (g7) & (g16) & (g44) & (!g46) & (g47)) + ((!g182) & (g7) & (g16) & (g44) & (g46) & (!g47)) + ((!g182) & (g7) & (g16) & (g44) & (g46) & (g47)) + ((g182) & (!g7) & (!g16) & (g44) & (!g46) & (g47)) + ((g182) & (!g7) & (!g16) & (g44) & (g46) & (g47)) + ((g182) & (!g7) & (g16) & (!g44) & (!g46) & (g47)) + ((g182) & (!g7) & (g16) & (!g44) & (g46) & (g47)) + ((g182) & (!g7) & (g16) & (g44) & (!g46) & (!g47)) + ((g182) & (!g7) & (g16) & (g44) & (!g46) & (g47)) + ((g182) & (!g7) & (g16) & (g44) & (g46) & (!g47)) + ((g182) & (!g7) & (g16) & (g44) & (g46) & (g47)) + ((g182) & (g7) & (!g16) & (g44) & (!g46) & (g47)) + ((g182) & (g7) & (!g16) & (g44) & (g46) & (!g47)) + ((g182) & (g7) & (!g16) & (g44) & (g46) & (g47)) + ((g182) & (g7) & (g16) & (!g44) & (!g46) & (g47)) + ((g182) & (g7) & (g16) & (!g44) & (g46) & (!g47)) + ((g182) & (g7) & (g16) & (!g44) & (g46) & (g47)) + ((g182) & (g7) & (g16) & (g44) & (!g46) & (!g47)) + ((g182) & (g7) & (g16) & (g44) & (!g46) & (g47)) + ((g182) & (g7) & (g16) & (g44) & (g46) & (!g47)) + ((g182) & (g7) & (g16) & (g44) & (g46) & (g47)));
	assign g115 = (((!g98) & (!g101) & (!g105) & (!g107) & (!g113) & (!g114)) + ((!g98) & (!g101) & (!g105) & (!g107) & (!g113) & (g114)) + ((!g98) & (!g101) & (!g105) & (!g107) & (g113) & (g114)) + ((!g98) & (!g101) & (!g105) & (g107) & (!g113) & (!g114)) + ((!g98) & (!g101) & (!g105) & (g107) & (!g113) & (g114)) + ((!g98) & (!g101) & (!g105) & (g107) & (g113) & (!g114)) + ((!g98) & (!g101) & (!g105) & (g107) & (g113) & (g114)) + ((!g98) & (!g101) & (g105) & (!g107) & (!g113) & (!g114)) + ((!g98) & (!g101) & (g105) & (!g107) & (!g113) & (g114)) + ((!g98) & (!g101) & (g105) & (!g107) & (g113) & (!g114)) + ((!g98) & (!g101) & (g105) & (!g107) & (g113) & (g114)) + ((!g98) & (!g101) & (g105) & (g107) & (!g113) & (!g114)) + ((!g98) & (!g101) & (g105) & (g107) & (!g113) & (g114)) + ((!g98) & (!g101) & (g105) & (g107) & (g113) & (!g114)) + ((!g98) & (!g101) & (g105) & (g107) & (g113) & (g114)) + ((!g98) & (g101) & (!g105) & (!g107) & (!g113) & (!g114)) + ((!g98) & (g101) & (!g105) & (!g107) & (!g113) & (g114)) + ((!g98) & (g101) & (!g105) & (!g107) & (g113) & (!g114)) + ((!g98) & (g101) & (!g105) & (!g107) & (g113) & (g114)) + ((!g98) & (g101) & (!g105) & (g107) & (!g113) & (!g114)) + ((!g98) & (g101) & (!g105) & (g107) & (!g113) & (g114)) + ((!g98) & (g101) & (!g105) & (g107) & (g113) & (!g114)) + ((!g98) & (g101) & (!g105) & (g107) & (g113) & (g114)) + ((!g98) & (g101) & (g105) & (!g107) & (!g113) & (!g114)) + ((!g98) & (g101) & (g105) & (!g107) & (!g113) & (g114)) + ((!g98) & (g101) & (g105) & (!g107) & (g113) & (!g114)) + ((!g98) & (g101) & (g105) & (!g107) & (g113) & (g114)) + ((!g98) & (g101) & (g105) & (g107) & (!g113) & (!g114)) + ((!g98) & (g101) & (g105) & (g107) & (!g113) & (g114)) + ((!g98) & (g101) & (g105) & (g107) & (g113) & (!g114)) + ((!g98) & (g101) & (g105) & (g107) & (g113) & (g114)) + ((g98) & (!g101) & (!g105) & (!g107) & (!g113) & (!g114)) + ((g98) & (!g101) & (!g105) & (!g107) & (!g113) & (g114)) + ((g98) & (!g101) & (!g105) & (!g107) & (g113) & (!g114)) + ((g98) & (!g101) & (!g105) & (!g107) & (g113) & (g114)) + ((g98) & (!g101) & (!g105) & (g107) & (!g113) & (!g114)) + ((g98) & (!g101) & (!g105) & (g107) & (!g113) & (g114)) + ((g98) & (!g101) & (!g105) & (g107) & (g113) & (!g114)) + ((g98) & (!g101) & (!g105) & (g107) & (g113) & (g114)) + ((g98) & (!g101) & (g105) & (!g107) & (!g113) & (!g114)) + ((g98) & (!g101) & (g105) & (!g107) & (!g113) & (g114)) + ((g98) & (!g101) & (g105) & (!g107) & (g113) & (!g114)) + ((g98) & (!g101) & (g105) & (!g107) & (g113) & (g114)) + ((g98) & (!g101) & (g105) & (g107) & (!g113) & (!g114)) + ((g98) & (!g101) & (g105) & (g107) & (!g113) & (g114)) + ((g98) & (!g101) & (g105) & (g107) & (g113) & (!g114)) + ((g98) & (!g101) & (g105) & (g107) & (g113) & (g114)) + ((g98) & (g101) & (!g105) & (!g107) & (!g113) & (!g114)) + ((g98) & (g101) & (!g105) & (!g107) & (!g113) & (g114)) + ((g98) & (g101) & (!g105) & (!g107) & (g113) & (!g114)) + ((g98) & (g101) & (!g105) & (!g107) & (g113) & (g114)) + ((g98) & (g101) & (!g105) & (g107) & (!g113) & (!g114)) + ((g98) & (g101) & (!g105) & (g107) & (!g113) & (g114)) + ((g98) & (g101) & (!g105) & (g107) & (g113) & (!g114)) + ((g98) & (g101) & (!g105) & (g107) & (g113) & (g114)) + ((g98) & (g101) & (g105) & (!g107) & (!g113) & (!g114)) + ((g98) & (g101) & (g105) & (!g107) & (!g113) & (g114)) + ((g98) & (g101) & (g105) & (!g107) & (g113) & (!g114)) + ((g98) & (g101) & (g105) & (!g107) & (g113) & (g114)) + ((g98) & (g101) & (g105) & (g107) & (!g113) & (!g114)) + ((g98) & (g101) & (g105) & (g107) & (!g113) & (g114)) + ((g98) & (g101) & (g105) & (g107) & (g113) & (!g114)) + ((g98) & (g101) & (g105) & (g107) & (g113) & (g114)));
	assign g119 = (((!g33) & (!sk[14]) & (!g35) & (c) & (!g) & (!g118)) + ((!g33) & (!sk[14]) & (!g35) & (c) & (!g) & (g118)) + ((!g33) & (!sk[14]) & (!g35) & (c) & (g) & (!g118)) + ((!g33) & (!sk[14]) & (!g35) & (c) & (g) & (g118)) + ((!g33) & (!sk[14]) & (g35) & (!c) & (!g) & (!g118)) + ((!g33) & (!sk[14]) & (g35) & (!c) & (!g) & (g118)) + ((!g33) & (!sk[14]) & (g35) & (!c) & (g) & (!g118)) + ((!g33) & (!sk[14]) & (g35) & (!c) & (g) & (g118)) + ((!g33) & (!sk[14]) & (g35) & (c) & (!g) & (!g118)) + ((!g33) & (!sk[14]) & (g35) & (c) & (!g) & (g118)) + ((!g33) & (!sk[14]) & (g35) & (c) & (g) & (!g118)) + ((!g33) & (!sk[14]) & (g35) & (c) & (g) & (g118)) + ((!g33) & (sk[14]) & (!g35) & (!c) & (g) & (g118)) + ((!g33) & (sk[14]) & (!g35) & (c) & (g) & (g118)) + ((!g33) & (sk[14]) & (g35) & (!c) & (g) & (g118)) + ((!g33) & (sk[14]) & (g35) & (c) & (!g) & (!g118)) + ((!g33) & (sk[14]) & (g35) & (c) & (!g) & (g118)) + ((!g33) & (sk[14]) & (g35) & (c) & (g) & (!g118)) + ((!g33) & (sk[14]) & (g35) & (c) & (g) & (g118)) + ((g33) & (!sk[14]) & (!g35) & (c) & (!g) & (!g118)) + ((g33) & (!sk[14]) & (!g35) & (c) & (!g) & (g118)) + ((g33) & (!sk[14]) & (!g35) & (c) & (g) & (!g118)) + ((g33) & (!sk[14]) & (!g35) & (c) & (g) & (g118)) + ((g33) & (!sk[14]) & (g35) & (!c) & (!g) & (!g118)) + ((g33) & (!sk[14]) & (g35) & (!c) & (!g) & (g118)) + ((g33) & (!sk[14]) & (g35) & (!c) & (g) & (!g118)) + ((g33) & (!sk[14]) & (g35) & (!c) & (g) & (g118)) + ((g33) & (!sk[14]) & (g35) & (c) & (!g) & (!g118)) + ((g33) & (!sk[14]) & (g35) & (c) & (!g) & (g118)) + ((g33) & (!sk[14]) & (g35) & (c) & (g) & (!g118)) + ((g33) & (!sk[14]) & (g35) & (c) & (g) & (g118)) + ((g33) & (sk[14]) & (!g35) & (!c) & (!g) & (!g118)) + ((g33) & (sk[14]) & (!g35) & (!c) & (!g) & (g118)) + ((g33) & (sk[14]) & (!g35) & (!c) & (g) & (!g118)) + ((g33) & (sk[14]) & (!g35) & (!c) & (g) & (g118)) + ((g33) & (sk[14]) & (!g35) & (c) & (!g) & (!g118)) + ((g33) & (sk[14]) & (!g35) & (c) & (!g) & (g118)) + ((g33) & (sk[14]) & (!g35) & (c) & (g) & (!g118)) + ((g33) & (sk[14]) & (!g35) & (c) & (g) & (g118)) + ((g33) & (sk[14]) & (g35) & (!c) & (!g) & (!g118)) + ((g33) & (sk[14]) & (g35) & (!c) & (!g) & (g118)) + ((g33) & (sk[14]) & (g35) & (!c) & (g) & (!g118)) + ((g33) & (sk[14]) & (g35) & (!c) & (g) & (g118)) + ((g33) & (sk[14]) & (g35) & (c) & (!g) & (!g118)) + ((g33) & (sk[14]) & (g35) & (c) & (!g) & (g118)) + ((g33) & (sk[14]) & (g35) & (c) & (g) & (!g118)) + ((g33) & (sk[14]) & (g35) & (c) & (g) & (g118)));
	assign g2 = (((!k) & (!l) & (!n) & (i) & (!sk[6]) & (!j)) + ((!k) & (!l) & (!n) & (i) & (!sk[6]) & (j)) + ((!k) & (!l) & (n) & (!i) & (!sk[6]) & (!j)) + ((!k) & (!l) & (n) & (!i) & (!sk[6]) & (j)) + ((!k) & (!l) & (n) & (!i) & (sk[6]) & (j)) + ((!k) & (!l) & (n) & (i) & (!sk[6]) & (!j)) + ((!k) & (!l) & (n) & (i) & (!sk[6]) & (j)) + ((!k) & (l) & (!n) & (i) & (!sk[6]) & (!j)) + ((!k) & (l) & (!n) & (i) & (!sk[6]) & (j)) + ((!k) & (l) & (n) & (!i) & (!sk[6]) & (!j)) + ((!k) & (l) & (n) & (!i) & (!sk[6]) & (j)) + ((!k) & (l) & (n) & (!i) & (sk[6]) & (j)) + ((!k) & (l) & (n) & (i) & (!sk[6]) & (!j)) + ((!k) & (l) & (n) & (i) & (!sk[6]) & (j)) + ((k) & (!l) & (!n) & (!i) & (!sk[6]) & (j)) + ((k) & (!l) & (!n) & (i) & (!sk[6]) & (!j)) + ((k) & (!l) & (!n) & (i) & (!sk[6]) & (j)) + ((k) & (!l) & (!n) & (i) & (sk[6]) & (j)) + ((k) & (!l) & (n) & (!i) & (!sk[6]) & (!j)) + ((k) & (!l) & (n) & (!i) & (!sk[6]) & (j)) + ((k) & (!l) & (n) & (i) & (!sk[6]) & (!j)) + ((k) & (!l) & (n) & (i) & (!sk[6]) & (j)) + ((k) & (!l) & (n) & (i) & (sk[6]) & (j)) + ((k) & (l) & (!n) & (!i) & (!sk[6]) & (j)) + ((k) & (l) & (!n) & (i) & (!sk[6]) & (!j)) + ((k) & (l) & (!n) & (i) & (!sk[6]) & (j)) + ((k) & (l) & (!n) & (i) & (sk[6]) & (!j)) + ((k) & (l) & (n) & (!i) & (!sk[6]) & (!j)) + ((k) & (l) & (n) & (!i) & (!sk[6]) & (j)) + ((k) & (l) & (n) & (!i) & (sk[6]) & (j)) + ((k) & (l) & (n) & (i) & (!sk[6]) & (!j)) + ((k) & (l) & (n) & (i) & (!sk[6]) & (j)));
	assign g4 = (((!k) & (!l) & (!sk[6]) & (!n) & (i) & (!j)) + ((!k) & (!l) & (!sk[6]) & (!n) & (i) & (j)) + ((!k) & (!l) & (!sk[6]) & (n) & (!i) & (!j)) + ((!k) & (!l) & (!sk[6]) & (n) & (!i) & (j)) + ((!k) & (!l) & (!sk[6]) & (n) & (i) & (!j)) + ((!k) & (!l) & (!sk[6]) & (n) & (i) & (j)) + ((!k) & (!l) & (sk[6]) & (!n) & (i) & (!j)) + ((!k) & (l) & (!sk[6]) & (!n) & (i) & (!j)) + ((!k) & (l) & (!sk[6]) & (!n) & (i) & (j)) + ((!k) & (l) & (!sk[6]) & (n) & (!i) & (!j)) + ((!k) & (l) & (!sk[6]) & (n) & (!i) & (j)) + ((!k) & (l) & (!sk[6]) & (n) & (i) & (!j)) + ((!k) & (l) & (!sk[6]) & (n) & (i) & (j)) + ((k) & (!l) & (!sk[6]) & (!n) & (i) & (!j)) + ((k) & (!l) & (!sk[6]) & (!n) & (i) & (j)) + ((k) & (!l) & (!sk[6]) & (n) & (!i) & (!j)) + ((k) & (!l) & (!sk[6]) & (n) & (!i) & (j)) + ((k) & (!l) & (!sk[6]) & (n) & (i) & (!j)) + ((k) & (!l) & (!sk[6]) & (n) & (i) & (j)) + ((k) & (!l) & (sk[6]) & (n) & (i) & (!j)) + ((k) & (l) & (!sk[6]) & (!n) & (i) & (!j)) + ((k) & (l) & (!sk[6]) & (!n) & (i) & (j)) + ((k) & (l) & (!sk[6]) & (n) & (!i) & (!j)) + ((k) & (l) & (!sk[6]) & (n) & (!i) & (j)) + ((k) & (l) & (!sk[6]) & (n) & (i) & (!j)) + ((k) & (l) & (!sk[6]) & (n) & (i) & (j)) + ((k) & (l) & (sk[6]) & (n) & (i) & (!j)));
	assign g17 = (((!sk[10]) & (!k) & (i) & (!j)) + ((!sk[10]) & (!k) & (i) & (j)) + ((!sk[10]) & (k) & (i) & (!j)) + ((!sk[10]) & (k) & (i) & (j)) + ((sk[10]) & (!k) & (!i) & (j)));
	assign g27 = (((!sk[8]) & (!k) & (!l) & (!n) & (i) & (!j)) + ((!sk[8]) & (!k) & (!l) & (!n) & (i) & (j)) + ((!sk[8]) & (!k) & (!l) & (n) & (i) & (!j)) + ((!sk[8]) & (!k) & (!l) & (n) & (i) & (j)) + ((!sk[8]) & (!k) & (l) & (!n) & (!i) & (!j)) + ((!sk[8]) & (!k) & (l) & (!n) & (!i) & (j)) + ((!sk[8]) & (!k) & (l) & (!n) & (i) & (!j)) + ((!sk[8]) & (!k) & (l) & (!n) & (i) & (j)) + ((!sk[8]) & (!k) & (l) & (n) & (!i) & (!j)) + ((!sk[8]) & (!k) & (l) & (n) & (!i) & (j)) + ((!sk[8]) & (!k) & (l) & (n) & (i) & (!j)) + ((!sk[8]) & (!k) & (l) & (n) & (i) & (j)) + ((!sk[8]) & (k) & (!l) & (!n) & (i) & (!j)) + ((!sk[8]) & (k) & (!l) & (!n) & (i) & (j)) + ((!sk[8]) & (k) & (!l) & (n) & (i) & (!j)) + ((!sk[8]) & (k) & (!l) & (n) & (i) & (j)) + ((!sk[8]) & (k) & (l) & (!n) & (!i) & (!j)) + ((!sk[8]) & (k) & (l) & (!n) & (!i) & (j)) + ((!sk[8]) & (k) & (l) & (!n) & (i) & (!j)) + ((!sk[8]) & (k) & (l) & (!n) & (i) & (j)) + ((!sk[8]) & (k) & (l) & (n) & (!i) & (!j)) + ((!sk[8]) & (k) & (l) & (n) & (!i) & (j)) + ((!sk[8]) & (k) & (l) & (n) & (i) & (!j)) + ((!sk[8]) & (k) & (l) & (n) & (i) & (j)) + ((sk[8]) & (!k) & (l) & (n) & (i) & (j)) + ((sk[8]) & (k) & (!l) & (n) & (!i) & (j)));
	assign g54 = (((!l) & (!sk[15]) & (g17)) + ((l) & (sk[15]) & (!g17)) + ((l) & (sk[15]) & (g17)));
	assign g55 = (((!sk[15]) & (!k) & (!l) & (!i) & (j)) + ((!sk[15]) & (!k) & (l) & (i) & (j)) + ((!sk[15]) & (k) & (!l) & (!i) & (j)) + ((sk[15]) & (!k) & (!l) & (!i) & (j)) + ((sk[15]) & (!k) & (!l) & (i) & (!j)) + ((sk[15]) & (!k) & (!l) & (i) & (j)) + ((sk[15]) & (!k) & (l) & (!i) & (j)) + ((sk[15]) & (!k) & (l) & (i) & (!j)) + ((sk[15]) & (!k) & (l) & (i) & (j)) + ((sk[15]) & (k) & (!l) & (!i) & (!j)) + ((sk[15]) & (k) & (!l) & (!i) & (j)) + ((sk[15]) & (k) & (!l) & (i) & (!j)) + ((sk[15]) & (k) & (!l) & (i) & (j)) + ((sk[15]) & (k) & (l) & (!i) & (!j)) + ((sk[15]) & (k) & (l) & (!i) & (j)) + ((sk[15]) & (k) & (l) & (i) & (!j)) + ((sk[15]) & (k) & (l) & (i) & (j)));
	assign g67 = (((!a) & (!e) & (!sk[2]) & (g15)) + ((!a) & (e) & (!sk[2]) & (g15)) + ((a) & (!e) & (!sk[2]) & (g15)) + ((a) & (e) & (!sk[2]) & (!g15)) + ((a) & (e) & (!sk[2]) & (g15)) + ((a) & (e) & (sk[2]) & (g15)));
	assign g68 = (((!k) & (!sk[3]) & (!l) & (g11)) + ((!k) & (!sk[3]) & (l) & (g11)) + ((!k) & (sk[3]) & (l) & (g11)) + ((k) & (!sk[3]) & (!l) & (!g11)) + ((k) & (!sk[3]) & (!l) & (g11)) + ((k) & (!sk[3]) & (l) & (!g11)) + ((k) & (!sk[3]) & (l) & (g11)));
	assign g81 = (((!a) & (!e) & (f) & (!sk[2]) & (!b)) + ((!a) & (!e) & (f) & (!sk[2]) & (b)) + ((!a) & (!e) & (f) & (sk[2]) & (!b)) + ((!a) & (e) & (!f) & (sk[2]) & (!b)) + ((!a) & (e) & (f) & (!sk[2]) & (!b)) + ((!a) & (e) & (f) & (!sk[2]) & (b)) + ((!a) & (e) & (f) & (sk[2]) & (!b)) + ((!a) & (e) & (f) & (sk[2]) & (b)) + ((a) & (!e) & (!f) & (!sk[2]) & (!b)) + ((a) & (!e) & (!f) & (!sk[2]) & (b)) + ((a) & (!e) & (f) & (!sk[2]) & (!b)) + ((a) & (!e) & (f) & (!sk[2]) & (b)) + ((a) & (!e) & (f) & (sk[2]) & (!b)) + ((a) & (e) & (!f) & (!sk[2]) & (!b)) + ((a) & (e) & (!f) & (!sk[2]) & (b)) + ((a) & (e) & (f) & (!sk[2]) & (!b)) + ((a) & (e) & (f) & (!sk[2]) & (b)) + ((a) & (e) & (f) & (sk[2]) & (!b)));
	assign g96 = (((!sk[2]) & (!a) & (!e) & (f) & (!b)) + ((!sk[2]) & (!a) & (!e) & (f) & (b)) + ((!sk[2]) & (!a) & (e) & (!f) & (!b)) + ((!sk[2]) & (!a) & (e) & (!f) & (b)) + ((!sk[2]) & (!a) & (e) & (f) & (!b)) + ((!sk[2]) & (!a) & (e) & (f) & (b)) + ((!sk[2]) & (a) & (!e) & (!f) & (!b)) + ((!sk[2]) & (a) & (!e) & (!f) & (b)) + ((!sk[2]) & (a) & (!e) & (f) & (!b)) + ((!sk[2]) & (a) & (!e) & (f) & (b)) + ((!sk[2]) & (a) & (e) & (!f) & (!b)) + ((!sk[2]) & (a) & (e) & (!f) & (b)) + ((!sk[2]) & (a) & (e) & (f) & (!b)) + ((!sk[2]) & (a) & (e) & (f) & (b)) + ((sk[2]) & (!a) & (!e) & (f) & (b)) + ((sk[2]) & (!a) & (e) & (f) & (b)) + ((sk[2]) & (a) & (!e) & (f) & (b)) + ((sk[2]) & (a) & (e) & (!f) & (b)) + ((sk[2]) & (a) & (e) & (f) & (!b)) + ((sk[2]) & (a) & (e) & (f) & (b)));
	assign g122 = (((!sk[14]) & (!c) & (!g) & (g81)) + ((!sk[14]) & (!c) & (g) & (g81)) + ((!sk[14]) & (c) & (!g) & (!g81)) + ((!sk[14]) & (c) & (!g) & (g81)) + ((!sk[14]) & (c) & (g) & (!g81)) + ((!sk[14]) & (c) & (g) & (g81)) + ((sk[14]) & (!c) & (!g) & (g81)) + ((sk[14]) & (!c) & (g) & (!g81)) + ((sk[14]) & (!c) & (g) & (g81)) + ((sk[14]) & (c) & (g) & (g81)));
	assign g147 = (((!c) & (!g) & (!sk[14]) & (g96)) + ((!c) & (g) & (!sk[14]) & (g96)) + ((!c) & (g) & (sk[14]) & (g96)) + ((c) & (!g) & (!sk[14]) & (g96)) + ((c) & (!g) & (sk[14]) & (g96)) + ((c) & (g) & (!sk[14]) & (g96)) + ((c) & (g) & (sk[14]) & (!g96)) + ((c) & (g) & (sk[14]) & (g96)));
	assign g152 = (((!a) & (!g14) & (!b) & (!g46) & (c) & (!g90)) + ((!a) & (!g14) & (!b) & (g46) & (c) & (!g90)) + ((!a) & (!g14) & (b) & (!g46) & (!c) & (!g90)) + ((!a) & (!g14) & (b) & (!g46) & (c) & (!g90)) + ((!a) & (!g14) & (b) & (!g46) & (c) & (g90)) + ((!a) & (!g14) & (b) & (g46) & (c) & (!g90)) + ((!a) & (g14) & (!b) & (!g46) & (c) & (!g90)) + ((!a) & (g14) & (!b) & (g46) & (c) & (!g90)) + ((!a) & (g14) & (b) & (!g46) & (!c) & (!g90)) + ((!a) & (g14) & (b) & (!g46) & (c) & (!g90)) + ((!a) & (g14) & (b) & (!g46) & (c) & (g90)) + ((!a) & (g14) & (b) & (g46) & (c) & (!g90)) + ((a) & (!g14) & (!b) & (!g46) & (!c) & (!g90)) + ((a) & (!g14) & (!b) & (!g46) & (c) & (!g90)) + ((a) & (!g14) & (!b) & (!g46) & (c) & (g90)) + ((a) & (!g14) & (!b) & (g46) & (c) & (!g90)) + ((a) & (!g14) & (b) & (!g46) & (!c) & (!g90)) + ((a) & (!g14) & (b) & (!g46) & (c) & (!g90)) + ((a) & (!g14) & (b) & (!g46) & (c) & (g90)) + ((a) & (!g14) & (b) & (g46) & (!c) & (!g90)) + ((a) & (!g14) & (b) & (g46) & (c) & (!g90)) + ((a) & (!g14) & (b) & (g46) & (c) & (g90)) + ((a) & (g14) & (!b) & (!g46) & (c) & (!g90)) + ((a) & (g14) & (!b) & (g46) & (c) & (!g90)) + ((a) & (g14) & (b) & (!g46) & (!c) & (!g90)) + ((a) & (g14) & (b) & (!g46) & (c) & (!g90)) + ((a) & (g14) & (b) & (!g46) & (c) & (g90)) + ((a) & (g14) & (b) & (g46) & (c) & (!g90)));
	assign g3 = (((!k) & (!l) & (!sk[8]) & (n) & (!i) & (!j)) + ((!k) & (!l) & (!sk[8]) & (n) & (!i) & (j)) + ((!k) & (!l) & (!sk[8]) & (n) & (i) & (!j)) + ((!k) & (!l) & (!sk[8]) & (n) & (i) & (j)) + ((!k) & (!l) & (sk[8]) & (!n) & (!i) & (!j)) + ((!k) & (!l) & (sk[8]) & (!n) & (!i) & (j)) + ((!k) & (l) & (!sk[8]) & (n) & (!i) & (!j)) + ((!k) & (l) & (!sk[8]) & (n) & (!i) & (j)) + ((!k) & (l) & (!sk[8]) & (n) & (i) & (!j)) + ((!k) & (l) & (!sk[8]) & (n) & (i) & (j)) + ((!k) & (l) & (sk[8]) & (!n) & (!i) & (!j)) + ((k) & (!l) & (!sk[8]) & (!n) & (i) & (!j)) + ((k) & (!l) & (!sk[8]) & (!n) & (i) & (j)) + ((k) & (!l) & (!sk[8]) & (n) & (!i) & (!j)) + ((k) & (!l) & (!sk[8]) & (n) & (!i) & (j)) + ((k) & (!l) & (!sk[8]) & (n) & (i) & (!j)) + ((k) & (!l) & (!sk[8]) & (n) & (i) & (j)) + ((k) & (l) & (!sk[8]) & (!n) & (i) & (!j)) + ((k) & (l) & (!sk[8]) & (!n) & (i) & (j)) + ((k) & (l) & (!sk[8]) & (n) & (!i) & (!j)) + ((k) & (l) & (!sk[8]) & (n) & (!i) & (j)) + ((k) & (l) & (!sk[8]) & (n) & (i) & (!j)) + ((k) & (l) & (!sk[8]) & (n) & (i) & (j)));
	assign g13 = (((!a) & (!g182) & (!g9) & (!sk[4]) & (!g10) & (!g12)) + ((!a) & (!g182) & (!g9) & (!sk[4]) & (!g10) & (g12)) + ((!a) & (!g182) & (g9) & (!sk[4]) & (!g10) & (!g12)) + ((!a) & (!g182) & (g9) & (!sk[4]) & (!g10) & (g12)) + ((!a) & (g182) & (!g9) & (!sk[4]) & (!g10) & (!g12)) + ((!a) & (g182) & (!g9) & (!sk[4]) & (g10) & (!g12)) + ((!a) & (g182) & (g9) & (!sk[4]) & (!g10) & (!g12)) + ((!a) & (g182) & (g9) & (!sk[4]) & (g10) & (!g12)) + ((a) & (!g182) & (!g9) & (!sk[4]) & (!g10) & (!g12)) + ((a) & (!g182) & (g9) & (!sk[4]) & (!g10) & (!g12)) + ((a) & (g182) & (!g9) & (!sk[4]) & (!g10) & (!g12)) + ((a) & (g182) & (!g9) & (!sk[4]) & (g10) & (!g12)));
	assign g18 = (((!sk[15]) & (l) & (g17)) + ((sk[15]) & (l) & (!g17)) + ((sk[15]) & (l) & (g17)));
	assign g23 = (((!sk[10]) & (!k) & (i) & (!g22)) + ((!sk[10]) & (!k) & (i) & (g22)) + ((!sk[10]) & (k) & (i) & (!g22)) + ((!sk[10]) & (k) & (i) & (g22)) + ((sk[10]) & (k) & (i) & (g22)));
	assign g28 = (((!sk[10]) & (i) & (!g22)) + ((!sk[10]) & (i) & (g22)) + ((sk[10]) & (i) & (g22)));
	assign g38 = (((!sk[11]) & (k) & (l) & (n) & (!i) & (!j)) + ((sk[11]) & (!k) & (!l) & (!n) & (i) & (!j)) + ((sk[11]) & (!k) & (!l) & (!n) & (i) & (j)) + ((sk[11]) & (!k) & (!l) & (n) & (i) & (!j)) + ((sk[11]) & (!k) & (!l) & (n) & (i) & (j)) + ((sk[11]) & (!k) & (l) & (!n) & (i) & (!j)) + ((sk[11]) & (!k) & (l) & (!n) & (i) & (j)) + ((sk[11]) & (!k) & (l) & (n) & (i) & (!j)) + ((sk[11]) & (!k) & (l) & (n) & (i) & (j)) + ((sk[11]) & (k) & (!l) & (!n) & (i) & (!j)) + ((sk[11]) & (k) & (!l) & (!n) & (i) & (j)) + ((sk[11]) & (k) & (!l) & (n) & (i) & (!j)) + ((sk[11]) & (k) & (!l) & (n) & (i) & (j)) + ((sk[11]) & (k) & (l) & (!n) & (i) & (!j)) + ((sk[11]) & (k) & (l) & (!n) & (i) & (j)) + ((sk[11]) & (k) & (l) & (n) & (i) & (!j)) + ((sk[11]) & (k) & (l) & (n) & (i) & (j)));
	assign g41 = (((!k) & (!sk[11]) & (l) & (n) & (!i) & (!j)) + ((!k) & (!sk[11]) & (l) & (n) & (i) & (j)) + ((!k) & (sk[11]) & (l) & (!n) & (!i) & (!j)) + ((!k) & (sk[11]) & (l) & (!n) & (!i) & (j)) + ((!k) & (sk[11]) & (l) & (!n) & (i) & (!j)) + ((!k) & (sk[11]) & (l) & (!n) & (i) & (j)) + ((!k) & (sk[11]) & (l) & (n) & (!i) & (!j)) + ((!k) & (sk[11]) & (l) & (n) & (!i) & (j)) + ((!k) & (sk[11]) & (l) & (n) & (i) & (!j)) + ((!k) & (sk[11]) & (l) & (n) & (i) & (j)) + ((k) & (!sk[11]) & (!l) & (!n) & (!i) & (!j)) + ((k) & (!sk[11]) & (!l) & (n) & (!i) & (!j)) + ((k) & (!sk[11]) & (!l) & (n) & (i) & (!j)) + ((k) & (sk[11]) & (!l) & (!n) & (!i) & (!j)) + ((k) & (sk[11]) & (!l) & (!n) & (!i) & (j)) + ((k) & (sk[11]) & (!l) & (!n) & (i) & (!j)) + ((k) & (sk[11]) & (!l) & (!n) & (i) & (j)) + ((k) & (sk[11]) & (!l) & (n) & (!i) & (!j)) + ((k) & (sk[11]) & (!l) & (n) & (!i) & (j)) + ((k) & (sk[11]) & (!l) & (n) & (i) & (!j)) + ((k) & (sk[11]) & (!l) & (n) & (i) & (j)) + ((k) & (sk[11]) & (l) & (!n) & (!i) & (!j)) + ((k) & (sk[11]) & (l) & (!n) & (!i) & (j)) + ((k) & (sk[11]) & (l) & (!n) & (i) & (!j)) + ((k) & (sk[11]) & (l) & (!n) & (i) & (j)) + ((k) & (sk[11]) & (l) & (n) & (!i) & (!j)) + ((k) & (sk[11]) & (l) & (n) & (!i) & (j)) + ((k) & (sk[11]) & (l) & (n) & (i) & (!j)) + ((k) & (sk[11]) & (l) & (n) & (i) & (j)));
	assign g48 = (((!g7) & (!g46) & (!sk[5]) & (!g47)) + ((!g7) & (g46) & (!sk[5]) & (!g47)) + ((g7) & (!g46) & (!sk[5]) & (!g47)));
	assign g58 = (((n) & (!g46) & (!g48) & (!g49) & (!g52) & (g206)) + ((n) & (!g46) & (!g48) & (!g49) & (g52) & (!g206)) + ((n) & (!g46) & (!g48) & (!g49) & (g52) & (g206)) + ((n) & (!g46) & (!g48) & (g49) & (!g52) & (g206)) + ((n) & (!g46) & (!g48) & (g49) & (g52) & (!g206)) + ((n) & (!g46) & (!g48) & (g49) & (g52) & (g206)) + ((n) & (!g46) & (g48) & (!g49) & (!g52) & (g206)) + ((n) & (!g46) & (g48) & (!g49) & (g52) & (!g206)) + ((n) & (!g46) & (g48) & (!g49) & (g52) & (g206)) + ((n) & (!g46) & (g48) & (g49) & (!g52) & (g206)) + ((n) & (!g46) & (g48) & (g49) & (g52) & (!g206)) + ((n) & (!g46) & (g48) & (g49) & (g52) & (g206)) + ((n) & (g46) & (!g48) & (!g49) & (!g52) & (g206)) + ((n) & (g46) & (!g48) & (!g49) & (g52) & (!g206)) + ((n) & (g46) & (!g48) & (!g49) & (g52) & (g206)) + ((n) & (g46) & (!g48) & (g49) & (!g52) & (g206)) + ((n) & (g46) & (!g48) & (g49) & (g52) & (!g206)) + ((n) & (g46) & (!g48) & (g49) & (g52) & (g206)) + ((n) & (g46) & (g48) & (!g49) & (!g52) & (g206)) + ((n) & (g46) & (g48) & (!g49) & (g52) & (!g206)) + ((n) & (g46) & (g48) & (!g49) & (g52) & (g206)) + ((n) & (g46) & (g48) & (g49) & (!g52) & (!g206)) + ((n) & (g46) & (g48) & (g49) & (!g52) & (g206)) + ((n) & (g46) & (g48) & (g49) & (g52) & (!g206)) + ((n) & (g46) & (g48) & (g49) & (g52) & (g206)));
	assign g59 = (((!g182) & (!g16) & (!g23) & (g44) & (!sk[16]) & (!g48)) + ((!g182) & (!g16) & (!g23) & (g44) & (!sk[16]) & (g48)) + ((!g182) & (!g16) & (g23) & (!g44) & (sk[16]) & (!g48)) + ((!g182) & (!g16) & (g23) & (g44) & (!sk[16]) & (!g48)) + ((!g182) & (!g16) & (g23) & (g44) & (!sk[16]) & (g48)) + ((!g182) & (!g16) & (g23) & (g44) & (sk[16]) & (g48)) + ((!g182) & (g16) & (!g23) & (g44) & (!sk[16]) & (!g48)) + ((!g182) & (g16) & (!g23) & (g44) & (!sk[16]) & (g48)) + ((!g182) & (g16) & (g23) & (!g44) & (sk[16]) & (!g48)) + ((!g182) & (g16) & (g23) & (g44) & (!sk[16]) & (!g48)) + ((!g182) & (g16) & (g23) & (g44) & (!sk[16]) & (g48)) + ((!g182) & (g16) & (g23) & (g44) & (sk[16]) & (g48)) + ((g182) & (!g16) & (!g23) & (g44) & (!sk[16]) & (!g48)) + ((g182) & (!g16) & (!g23) & (g44) & (!sk[16]) & (g48)) + ((g182) & (!g16) & (g23) & (!g44) & (sk[16]) & (!g48)) + ((g182) & (!g16) & (g23) & (g44) & (!sk[16]) & (!g48)) + ((g182) & (!g16) & (g23) & (g44) & (!sk[16]) & (g48)) + ((g182) & (!g16) & (g23) & (g44) & (sk[16]) & (g48)) + ((g182) & (g16) & (!g23) & (g44) & (!sk[16]) & (!g48)) + ((g182) & (g16) & (!g23) & (g44) & (!sk[16]) & (g48)) + ((g182) & (g16) & (g23) & (!g44) & (!sk[16]) & (!g48)) + ((g182) & (g16) & (g23) & (!g44) & (!sk[16]) & (g48)) + ((g182) & (g16) & (g23) & (!g44) & (sk[16]) & (g48)) + ((g182) & (g16) & (g23) & (g44) & (!sk[16]) & (!g48)) + ((g182) & (g16) & (g23) & (g44) & (!sk[16]) & (g48)) + ((g182) & (g16) & (g23) & (g44) & (sk[16]) & (!g48)));
	assign g72 = (((!g60) & (!g61) & (g66) & (!sk[17]) & (!g70) & (!g71)) + ((!g60) & (!g61) & (g66) & (sk[17]) & (!g70) & (!g71)) + ((!g60) & (!g61) & (g66) & (sk[17]) & (!g70) & (g71)) + ((!g60) & (!g61) & (g66) & (sk[17]) & (g70) & (!g71)) + ((!g60) & (!g61) & (g66) & (sk[17]) & (g70) & (g71)) + ((!g60) & (g61) & (!g66) & (sk[17]) & (!g70) & (!g71)) + ((!g60) & (g61) & (!g66) & (sk[17]) & (!g70) & (g71)) + ((!g60) & (g61) & (!g66) & (sk[17]) & (g70) & (!g71)) + ((!g60) & (g61) & (!g66) & (sk[17]) & (g70) & (g71)) + ((!g60) & (g61) & (g66) & (!sk[17]) & (!g70) & (!g71)) + ((!g60) & (g61) & (g66) & (sk[17]) & (!g70) & (!g71)) + ((!g60) & (g61) & (g66) & (sk[17]) & (!g70) & (g71)) + ((!g60) & (g61) & (g66) & (sk[17]) & (g70) & (!g71)) + ((!g60) & (g61) & (g66) & (sk[17]) & (g70) & (g71)) + ((g60) & (!g61) & (g66) & (!sk[17]) & (!g70) & (!g71)) + ((g60) & (!g61) & (g66) & (sk[17]) & (!g70) & (!g71)) + ((g60) & (!g61) & (g66) & (sk[17]) & (!g70) & (g71)) + ((g60) & (!g61) & (g66) & (sk[17]) & (g70) & (!g71)) + ((g60) & (!g61) & (g66) & (sk[17]) & (g70) & (g71)) + ((g60) & (g61) & (!g66) & (sk[17]) & (!g70) & (!g71)) + ((g60) & (g61) & (!g66) & (sk[17]) & (!g70) & (g71)) + ((g60) & (g61) & (!g66) & (sk[17]) & (g70) & (!g71)) + ((g60) & (g61) & (!g66) & (sk[17]) & (g70) & (g71)) + ((g60) & (g61) & (g66) & (sk[17]) & (!g70) & (!g71)) + ((g60) & (g61) & (g66) & (sk[17]) & (!g70) & (g71)) + ((g60) & (g61) & (g66) & (sk[17]) & (g70) & (!g71)) + ((g60) & (g61) & (g66) & (sk[17]) & (g70) & (g71)));
	assign g82 = (((!sk[14]) & (!g1) & (!g11) & (!c) & (!g) & (g81)) + ((!sk[14]) & (!g1) & (!g11) & (!c) & (g) & (g81)) + ((!sk[14]) & (!g1) & (!g11) & (c) & (!g) & (g81)) + ((!sk[14]) & (!g1) & (!g11) & (c) & (g) & (g81)) + ((!sk[14]) & (!g1) & (g11) & (!c) & (!g) & (g81)) + ((!sk[14]) & (!g1) & (g11) & (!c) & (g) & (g81)) + ((!sk[14]) & (!g1) & (g11) & (c) & (!g) & (!g81)) + ((!sk[14]) & (!g1) & (g11) & (c) & (!g) & (g81)) + ((!sk[14]) & (!g1) & (g11) & (c) & (g) & (!g81)) + ((!sk[14]) & (!g1) & (g11) & (c) & (g) & (g81)) + ((!sk[14]) & (g1) & (!g11) & (!c) & (!g) & (!g81)) + ((!sk[14]) & (g1) & (!g11) & (!c) & (!g) & (g81)) + ((!sk[14]) & (g1) & (!g11) & (!c) & (g) & (!g81)) + ((!sk[14]) & (g1) & (!g11) & (!c) & (g) & (g81)) + ((!sk[14]) & (g1) & (!g11) & (c) & (!g) & (!g81)) + ((!sk[14]) & (g1) & (!g11) & (c) & (!g) & (g81)) + ((!sk[14]) & (g1) & (!g11) & (c) & (g) & (!g81)) + ((!sk[14]) & (g1) & (!g11) & (c) & (g) & (g81)) + ((!sk[14]) & (g1) & (g11) & (!c) & (!g) & (!g81)) + ((!sk[14]) & (g1) & (g11) & (!c) & (!g) & (g81)) + ((!sk[14]) & (g1) & (g11) & (!c) & (g) & (!g81)) + ((!sk[14]) & (g1) & (g11) & (!c) & (g) & (g81)) + ((!sk[14]) & (g1) & (g11) & (c) & (!g) & (!g81)) + ((!sk[14]) & (g1) & (g11) & (c) & (!g) & (g81)) + ((!sk[14]) & (g1) & (g11) & (c) & (g) & (!g81)) + ((!sk[14]) & (g1) & (g11) & (c) & (g) & (g81)) + ((sk[14]) & (!g1) & (g11) & (c) & (!g) & (!g81)) + ((sk[14]) & (g1) & (g11) & (!c) & (g) & (!g81)) + ((sk[14]) & (g1) & (g11) & (c) & (!g) & (!g81)));
	assign g87 = (((!b) & (!sk[18]) & (g38) & (!g84) & (!g85) & (!g86)) + ((!b) & (!sk[18]) & (g38) & (!g84) & (!g85) & (g86)) + ((!b) & (!sk[18]) & (g38) & (!g84) & (g85) & (!g86)) + ((!b) & (!sk[18]) & (g38) & (!g84) & (g85) & (g86)) + ((!b) & (!sk[18]) & (g38) & (g84) & (!g85) & (!g86)) + ((!b) & (!sk[18]) & (g38) & (g84) & (!g85) & (g86)) + ((!b) & (!sk[18]) & (g38) & (g84) & (g85) & (!g86)) + ((!b) & (!sk[18]) & (g38) & (g84) & (g85) & (g86)) + ((!b) & (sk[18]) & (!g38) & (!g84) & (!g85) & (!g86)) + ((!b) & (sk[18]) & (g38) & (!g84) & (!g85) & (!g86)) + ((b) & (!sk[18]) & (g38) & (!g84) & (!g85) & (!g86)) + ((b) & (!sk[18]) & (g38) & (!g84) & (!g85) & (g86)) + ((b) & (!sk[18]) & (g38) & (!g84) & (g85) & (!g86)) + ((b) & (!sk[18]) & (g38) & (!g84) & (g85) & (g86)) + ((b) & (!sk[18]) & (g38) & (g84) & (!g85) & (!g86)) + ((b) & (!sk[18]) & (g38) & (g84) & (!g85) & (g86)) + ((b) & (!sk[18]) & (g38) & (g84) & (g85) & (!g86)) + ((b) & (!sk[18]) & (g38) & (g84) & (g85) & (g86)) + ((b) & (sk[18]) & (!g38) & (!g84) & (!g85) & (!g86)));
	assign g91 = (((!a) & (!g14) & (!b) & (!sk[5]) & (!g46) & (!g90)) + ((!a) & (!g14) & (!b) & (!sk[5]) & (g46) & (!g90)) + ((!a) & (!g14) & (b) & (!sk[5]) & (!g46) & (g90)) + ((!a) & (!g14) & (b) & (!sk[5]) & (g46) & (!g90)) + ((!a) & (g14) & (!b) & (!sk[5]) & (!g46) & (!g90)) + ((!a) & (g14) & (!b) & (!sk[5]) & (g46) & (!g90)) + ((!a) & (g14) & (b) & (!sk[5]) & (!g46) & (g90)) + ((!a) & (g14) & (b) & (!sk[5]) & (g46) & (!g90)) + ((a) & (!g14) & (!b) & (!sk[5]) & (!g46) & (g90)) + ((a) & (!g14) & (!b) & (!sk[5]) & (g46) & (!g90)) + ((a) & (!g14) & (b) & (!sk[5]) & (!g46) & (g90)) + ((a) & (!g14) & (b) & (!sk[5]) & (g46) & (g90)) + ((a) & (g14) & (!b) & (!sk[5]) & (!g46) & (!g90)) + ((a) & (g14) & (!b) & (!sk[5]) & (g46) & (!g90)) + ((a) & (g14) & (b) & (!sk[5]) & (!g46) & (g90)) + ((a) & (g14) & (b) & (!sk[5]) & (g46) & (!g90)));
	assign g102 = (((!g15) & (!sk[14]) & (!c) & (g)) + ((!g15) & (!sk[14]) & (c) & (!g)) + ((!g15) & (!sk[14]) & (c) & (g)) + ((g15) & (!sk[14]) & (!c) & (g)) + ((g15) & (!sk[14]) & (c) & (!g)) + ((g15) & (!sk[14]) & (c) & (g)) + ((g15) & (sk[14]) & (c) & (g)));
	assign g106 = (((!g7) & (!sk[5]) & (!g67) & (!g46) & (!g47)) + ((!g7) & (!sk[5]) & (!g67) & (g46) & (!g47)) + ((!g7) & (!sk[5]) & (!g67) & (g46) & (g47)) + ((!g7) & (!sk[5]) & (g67) & (g46) & (!g47)) + ((g7) & (!sk[5]) & (!g67) & (!g46) & (!g47)) + ((g7) & (!sk[5]) & (!g67) & (g46) & (!g47)) + ((g7) & (!sk[5]) & (!g67) & (g46) & (g47)));
	assign g109 = (((!g27) & (sk[19]) & (g62) & (!g93)) + ((!g27) & (sk[19]) & (g62) & (g93)) + ((g27) & (!sk[19]) & (g62) & (g93)) + ((g27) & (sk[19]) & (g62) & (!g93)) + ((g27) & (sk[19]) & (g62) & (g93)));
	assign g120 = (((g14) & (!sk[20]) & (g46) & (g90)) + ((g14) & (sk[20]) & (!g46) & (g90)) + ((g14) & (sk[20]) & (g46) & (g90)));
	assign g124 = (((!sk[11]) & (n) & (g121) & (g123)) + ((sk[11]) & (!n) & (g121) & (!g123)) + ((sk[11]) & (!n) & (g121) & (g123)) + ((sk[11]) & (n) & (g121) & (!g123)) + ((sk[11]) & (n) & (g121) & (g123)));
	assign g132 = (((!g11) & (!sk[20]) & (!g122) & (!g127) & (!g128) & (g131)) + ((!g11) & (!sk[20]) & (!g122) & (!g127) & (g128) & (g131)) + ((!g11) & (!sk[20]) & (g122) & (!g127) & (!g128) & (g131)) + ((!g11) & (!sk[20]) & (g122) & (!g127) & (g128) & (g131)) + ((!g11) & (sk[20]) & (!g122) & (!g127) & (!g128) & (g131)) + ((!g11) & (sk[20]) & (!g122) & (!g127) & (g128) & (g131)) + ((!g11) & (sk[20]) & (!g122) & (g127) & (!g128) & (g131)) + ((!g11) & (sk[20]) & (!g122) & (g127) & (g128) & (!g131)) + ((!g11) & (sk[20]) & (!g122) & (g127) & (g128) & (g131)) + ((!g11) & (sk[20]) & (g122) & (!g127) & (!g128) & (g131)) + ((!g11) & (sk[20]) & (g122) & (!g127) & (g128) & (g131)) + ((!g11) & (sk[20]) & (g122) & (g127) & (!g128) & (!g131)) + ((!g11) & (sk[20]) & (g122) & (g127) & (!g128) & (g131)) + ((!g11) & (sk[20]) & (g122) & (g127) & (g128) & (!g131)) + ((!g11) & (sk[20]) & (g122) & (g127) & (g128) & (g131)) + ((g11) & (!sk[20]) & (!g122) & (!g127) & (!g128) & (g131)) + ((g11) & (!sk[20]) & (g122) & (!g127) & (!g128) & (g131)) + ((g11) & (!sk[20]) & (g122) & (!g127) & (g128) & (g131)) + ((g11) & (sk[20]) & (!g122) & (!g127) & (!g128) & (g131)) + ((g11) & (sk[20]) & (!g122) & (!g127) & (g128) & (g131)) + ((g11) & (sk[20]) & (!g122) & (g127) & (!g128) & (g131)) + ((g11) & (sk[20]) & (!g122) & (g127) & (g128) & (!g131)) + ((g11) & (sk[20]) & (!g122) & (g127) & (g128) & (g131)) + ((g11) & (sk[20]) & (g122) & (!g127) & (!g128) & (g131)) + ((g11) & (sk[20]) & (g122) & (!g127) & (g128) & (g131)) + ((g11) & (sk[20]) & (g122) & (g127) & (!g128) & (!g131)) + ((g11) & (sk[20]) & (g122) & (g127) & (!g128) & (g131)) + ((g11) & (sk[20]) & (g122) & (g127) & (g128) & (!g131)) + ((g11) & (sk[20]) & (g122) & (g127) & (g128) & (g131)));
	assign g139 = (((!g7) & (!g67) & (!g46) & (!g47) & (!g90) & (!g102)) + ((!g7) & (!g67) & (!g46) & (!g47) & (g90) & (!g102)) + ((!g7) & (!g67) & (!g46) & (!g47) & (g90) & (g102)) + ((!g7) & (!g67) & (!g46) & (g47) & (g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (!g47) & (!g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (!g47) & (g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (!g47) & (g90) & (g102)) + ((!g7) & (!g67) & (g46) & (g47) & (!g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (g47) & (g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (g47) & (g90) & (g102)) + ((!g7) & (g67) & (!g46) & (!g47) & (g90) & (!g102)) + ((!g7) & (g67) & (!g46) & (g47) & (g90) & (!g102)) + ((!g7) & (g67) & (g46) & (!g47) & (!g90) & (!g102)) + ((!g7) & (g67) & (g46) & (!g47) & (g90) & (!g102)) + ((!g7) & (g67) & (g46) & (!g47) & (g90) & (g102)) + ((!g7) & (g67) & (g46) & (g47) & (g90) & (!g102)) + ((g7) & (!g67) & (!g46) & (!g47) & (!g90) & (!g102)) + ((g7) & (!g67) & (!g46) & (!g47) & (g90) & (!g102)) + ((g7) & (!g67) & (!g46) & (!g47) & (g90) & (g102)) + ((g7) & (!g67) & (g46) & (!g47) & (!g90) & (!g102)) + ((g7) & (!g67) & (g46) & (!g47) & (g90) & (!g102)) + ((g7) & (!g67) & (g46) & (!g47) & (g90) & (g102)) + ((g7) & (!g67) & (g46) & (g47) & (!g90) & (!g102)) + ((g7) & (!g67) & (g46) & (g47) & (g90) & (!g102)) + ((g7) & (!g67) & (g46) & (g47) & (g90) & (g102)));
	assign g156 = (((!g137) & (!g140) & (!g142) & (!g143) & (g151) & (!g155)));
	assign g163 = (((!d) & (!sk[9]) & (h)) + ((d) & (!sk[9]) & (!h)) + ((d) & (sk[9]) & (!h)) + ((d) & (sk[9]) & (h)));
	assign g5 = (((!k) & (!l) & (!i) & (!a) & (!e) & (g182)) + ((!k) & (!l) & (!i) & (!a) & (e) & (g182)) + ((!k) & (!l) & (!i) & (a) & (!e) & (g182)) + ((!k) & (!l) & (!i) & (a) & (e) & (g182)) + ((!k) & (!l) & (i) & (!a) & (!e) & (!g182)) + ((!k) & (!l) & (i) & (!a) & (e) & (!g182)) + ((!k) & (!l) & (i) & (a) & (!e) & (!g182)) + ((!k) & (!l) & (i) & (a) & (e) & (!g182)) + ((!k) & (l) & (!i) & (!a) & (!e) & (g182)) + ((!k) & (l) & (!i) & (!a) & (e) & (g182)) + ((!k) & (l) & (!i) & (a) & (!e) & (!g182)) + ((!k) & (l) & (!i) & (a) & (!e) & (g182)) + ((!k) & (l) & (!i) & (a) & (e) & (g182)) + ((!k) & (l) & (i) & (!a) & (e) & (!g182)) + ((!k) & (l) & (i) & (!a) & (e) & (g182)) + ((!k) & (l) & (i) & (a) & (!e) & (!g182)) + ((!k) & (l) & (i) & (a) & (!e) & (g182)) + ((k) & (!l) & (!i) & (!a) & (!e) & (!g182)) + ((k) & (!l) & (!i) & (!a) & (e) & (!g182)) + ((k) & (!l) & (!i) & (a) & (!e) & (!g182)) + ((k) & (!l) & (!i) & (a) & (e) & (!g182)) + ((k) & (!l) & (i) & (!a) & (!e) & (!g182)) + ((k) & (!l) & (i) & (!a) & (!e) & (g182)) + ((k) & (!l) & (i) & (a) & (!e) & (!g182)) + ((k) & (!l) & (i) & (a) & (!e) & (g182)) + ((k) & (l) & (!i) & (!a) & (!e) & (!g182)) + ((k) & (l) & (!i) & (!a) & (!e) & (g182)) + ((k) & (l) & (!i) & (!a) & (e) & (!g182)) + ((k) & (l) & (!i) & (!a) & (e) & (g182)) + ((k) & (l) & (!i) & (a) & (!e) & (!g182)) + ((k) & (l) & (!i) & (a) & (!e) & (g182)) + ((k) & (l) & (!i) & (a) & (e) & (!g182)) + ((k) & (l) & (!i) & (a) & (e) & (g182)) + ((k) & (l) & (i) & (!a) & (!e) & (g182)) + ((k) & (l) & (i) & (!a) & (e) & (g182)) + ((k) & (l) & (i) & (a) & (!e) & (!g182)) + ((k) & (l) & (i) & (a) & (!e) & (g182)) + ((k) & (l) & (i) & (a) & (e) & (g182)));
	assign g6 = (((!k) & (l) & (!i) & (!a) & (e) & (!g182)) + ((!k) & (l) & (!i) & (!a) & (e) & (g182)) + ((!k) & (l) & (!i) & (a) & (e) & (!g182)) + ((!k) & (l) & (!i) & (a) & (e) & (g182)) + ((k) & (!l) & (!i) & (!a) & (!e) & (!g182)) + ((k) & (!l) & (!i) & (!a) & (!e) & (g182)) + ((k) & (!l) & (i) & (a) & (!e) & (g182)) + ((k) & (!l) & (i) & (a) & (e) & (g182)) + ((k) & (l) & (!i) & (!a) & (e) & (!g182)) + ((k) & (l) & (!i) & (!a) & (e) & (g182)) + ((k) & (l) & (!i) & (a) & (e) & (!g182)) + ((k) & (l) & (!i) & (a) & (e) & (g182)) + ((k) & (l) & (i) & (a) & (!e) & (g182)) + ((k) & (l) & (i) & (a) & (e) & (g182)));
	assign g19 = (((!l) & (!i) & (!j) & (a) & (!e) & (!g182)) + ((!l) & (!i) & (!j) & (a) & (!e) & (g182)) + ((!l) & (!i) & (!j) & (a) & (e) & (!g182)) + ((!l) & (!i) & (!j) & (a) & (e) & (g182)) + ((!l) & (!i) & (j) & (!a) & (!e) & (g182)) + ((!l) & (!i) & (j) & (!a) & (e) & (g182)) + ((!l) & (!i) & (j) & (a) & (!e) & (!g182)) + ((!l) & (!i) & (j) & (a) & (!e) & (g182)) + ((!l) & (!i) & (j) & (a) & (e) & (!g182)) + ((!l) & (!i) & (j) & (a) & (e) & (g182)) + ((!l) & (i) & (!j) & (!a) & (e) & (!g182)) + ((!l) & (i) & (!j) & (!a) & (e) & (g182)) + ((!l) & (i) & (!j) & (a) & (!e) & (!g182)) + ((!l) & (i) & (!j) & (a) & (!e) & (g182)) + ((l) & (!i) & (!j) & (a) & (!e) & (!g182)) + ((l) & (!i) & (!j) & (a) & (e) & (!g182)) + ((l) & (i) & (!j) & (!a) & (e) & (!g182)) + ((l) & (i) & (!j) & (!a) & (e) & (g182)) + ((l) & (i) & (!j) & (a) & (!e) & (!g182)) + ((l) & (i) & (!j) & (a) & (!e) & (g182)));
	assign g20 = (((!k) & (l) & (!i) & (!j) & (!a) & (g182)) + ((k) & (l) & (!i) & (!j) & (!a) & (g182)) + ((k) & (l) & (!i) & (!j) & (a) & (!g182)) + ((k) & (l) & (!i) & (j) & (!a) & (g182)) + ((k) & (l) & (!i) & (j) & (a) & (!g182)) + ((k) & (l) & (i) & (!j) & (!a) & (g182)) + ((k) & (l) & (i) & (!j) & (a) & (!g182)) + ((k) & (l) & (i) & (j) & (!a) & (g182)));
	assign g21 = (((!k) & (!g14) & (!g16) & (!g18) & (!g19) & (!g20)) + ((!k) & (!g14) & (g16) & (!g18) & (!g19) & (!g20)) + ((!k) & (!g14) & (g16) & (g18) & (!g19) & (!g20)) + ((!k) & (g14) & (!g16) & (!g18) & (!g19) & (!g20)) + ((!k) & (g14) & (!g16) & (g18) & (!g19) & (!g20)) + ((!k) & (g14) & (g16) & (!g18) & (!g19) & (!g20)) + ((k) & (!g14) & (!g16) & (!g18) & (!g19) & (!g20)) + ((k) & (!g14) & (!g16) & (!g18) & (g19) & (!g20)) + ((k) & (!g14) & (g16) & (!g18) & (!g19) & (!g20)) + ((k) & (!g14) & (g16) & (!g18) & (g19) & (!g20)) + ((k) & (!g14) & (g16) & (g18) & (!g19) & (!g20)) + ((k) & (!g14) & (g16) & (g18) & (g19) & (!g20)) + ((k) & (g14) & (!g16) & (!g18) & (!g19) & (!g20)) + ((k) & (g14) & (!g16) & (!g18) & (g19) & (!g20)) + ((k) & (g14) & (!g16) & (g18) & (!g19) & (!g20)) + ((k) & (g14) & (!g16) & (g18) & (g19) & (!g20)) + ((k) & (g14) & (g16) & (!g18) & (!g19) & (!g20)) + ((k) & (g14) & (g16) & (!g18) & (g19) & (!g20)));
	assign g24 = (((!g182) & (!g16) & (!sk[16]) & (g23)) + ((!g182) & (g16) & (!sk[16]) & (g23)) + ((!g182) & (g16) & (sk[16]) & (g23)) + ((g182) & (!g16) & (!sk[16]) & (!g23)) + ((g182) & (!g16) & (!sk[16]) & (g23)) + ((g182) & (!g16) & (sk[16]) & (g23)) + ((g182) & (g16) & (!sk[16]) & (!g23)) + ((g182) & (g16) & (!sk[16]) & (g23)));
	assign g25 = (((k) & (!l) & (n) & (g8) & (!a) & (g14)) + ((k) & (!l) & (n) & (g8) & (a) & (g14)) + ((k) & (l) & (n) & (g8) & (!a) & (!g14)) + ((k) & (l) & (n) & (g8) & (!a) & (g14)));
	assign g29 = (((!k) & (!e) & (!g182) & (g27) & (!sk[12]) & (!g28)) + ((!k) & (!e) & (!g182) & (g27) & (!sk[12]) & (g28)) + ((!k) & (!e) & (!g182) & (g27) & (sk[12]) & (!g28)) + ((!k) & (!e) & (!g182) & (g27) & (sk[12]) & (g28)) + ((!k) & (!e) & (g182) & (!g27) & (sk[12]) & (!g28)) + ((!k) & (!e) & (g182) & (!g27) & (sk[12]) & (g28)) + ((!k) & (!e) & (g182) & (g27) & (sk[12]) & (!g28)) + ((!k) & (!e) & (g182) & (g27) & (sk[12]) & (g28)) + ((!k) & (e) & (!g182) & (!g27) & (!sk[12]) & (g28)) + ((!k) & (e) & (!g182) & (!g27) & (sk[12]) & (!g28)) + ((!k) & (e) & (!g182) & (!g27) & (sk[12]) & (g28)) + ((!k) & (e) & (!g182) & (g27) & (!sk[12]) & (!g28)) + ((!k) & (e) & (!g182) & (g27) & (!sk[12]) & (g28)) + ((!k) & (e) & (!g182) & (g27) & (sk[12]) & (!g28)) + ((!k) & (e) & (!g182) & (g27) & (sk[12]) & (g28)) + ((!k) & (e) & (g182) & (!g27) & (!sk[12]) & (g28)) + ((!k) & (e) & (g182) & (!g27) & (sk[12]) & (!g28)) + ((!k) & (e) & (g182) & (!g27) & (sk[12]) & (g28)) + ((!k) & (e) & (g182) & (g27) & (!sk[12]) & (g28)) + ((!k) & (e) & (g182) & (g27) & (sk[12]) & (!g28)) + ((!k) & (e) & (g182) & (g27) & (sk[12]) & (g28)) + ((k) & (!e) & (!g182) & (!g27) & (sk[12]) & (!g28)) + ((k) & (!e) & (!g182) & (!g27) & (sk[12]) & (g28)) + ((k) & (!e) & (!g182) & (g27) & (!sk[12]) & (!g28)) + ((k) & (!e) & (!g182) & (g27) & (!sk[12]) & (g28)) + ((k) & (!e) & (!g182) & (g27) & (sk[12]) & (!g28)) + ((k) & (!e) & (!g182) & (g27) & (sk[12]) & (g28)) + ((k) & (!e) & (g182) & (!g27) & (sk[12]) & (!g28)) + ((k) & (!e) & (g182) & (!g27) & (sk[12]) & (g28)) + ((k) & (!e) & (g182) & (g27) & (sk[12]) & (!g28)) + ((k) & (!e) & (g182) & (g27) & (sk[12]) & (g28)) + ((k) & (e) & (!g182) & (!g27) & (sk[12]) & (!g28)) + ((k) & (e) & (!g182) & (!g27) & (sk[12]) & (g28)) + ((k) & (e) & (!g182) & (g27) & (!sk[12]) & (!g28)) + ((k) & (e) & (!g182) & (g27) & (!sk[12]) & (g28)) + ((k) & (e) & (!g182) & (g27) & (sk[12]) & (!g28)) + ((k) & (e) & (!g182) & (g27) & (sk[12]) & (g28)) + ((k) & (e) & (g182) & (!g27) & (sk[12]) & (!g28)) + ((k) & (e) & (g182) & (!g27) & (sk[12]) & (g28)) + ((k) & (e) & (g182) & (g27) & (sk[12]) & (!g28)) + ((k) & (e) & (g182) & (g27) & (sk[12]) & (g28)));
	assign g30 = (((!sk[20]) & (!k) & (!a) & (!g14) & (!g26) & (!g29)) + ((!sk[20]) & (!k) & (!a) & (!g14) & (g26) & (!g29)) + ((!sk[20]) & (!k) & (!a) & (g14) & (!g26) & (!g29)) + ((!sk[20]) & (!k) & (!a) & (g14) & (g26) & (!g29)) + ((!sk[20]) & (!k) & (a) & (!g14) & (!g26) & (!g29)) + ((!sk[20]) & (!k) & (a) & (!g14) & (g26) & (!g29)) + ((!sk[20]) & (!k) & (a) & (g14) & (!g26) & (!g29)) + ((!sk[20]) & (k) & (!a) & (!g14) & (!g26) & (!g29)) + ((!sk[20]) & (k) & (!a) & (g14) & (!g26) & (!g29)) + ((!sk[20]) & (k) & (!a) & (g14) & (g26) & (!g29)) + ((!sk[20]) & (k) & (a) & (!g14) & (!g26) & (!g29)) + ((!sk[20]) & (k) & (a) & (!g14) & (g26) & (!g29)) + ((!sk[20]) & (k) & (a) & (g14) & (!g26) & (!g29)));
	assign g36 = (((!g33) & (!a) & (!sk[21]) & (!e) & (!g34) & (g35)) + ((!g33) & (!a) & (!sk[21]) & (!e) & (g34) & (!g35)) + ((!g33) & (!a) & (!sk[21]) & (!e) & (g34) & (g35)) + ((!g33) & (!a) & (!sk[21]) & (e) & (!g34) & (g35)) + ((!g33) & (!a) & (!sk[21]) & (e) & (g34) & (!g35)) + ((!g33) & (!a) & (!sk[21]) & (e) & (g34) & (g35)) + ((!g33) & (!a) & (sk[21]) & (!e) & (!g34) & (!g35)) + ((!g33) & (!a) & (sk[21]) & (!e) & (!g34) & (g35)) + ((!g33) & (!a) & (sk[21]) & (!e) & (g34) & (!g35)) + ((!g33) & (!a) & (sk[21]) & (!e) & (g34) & (g35)) + ((!g33) & (!a) & (sk[21]) & (e) & (!g34) & (!g35)) + ((!g33) & (!a) & (sk[21]) & (e) & (!g34) & (g35)) + ((!g33) & (!a) & (sk[21]) & (e) & (g34) & (!g35)) + ((!g33) & (!a) & (sk[21]) & (e) & (g34) & (g35)) + ((!g33) & (a) & (!sk[21]) & (!e) & (!g34) & (!g35)) + ((!g33) & (a) & (!sk[21]) & (!e) & (!g34) & (g35)) + ((!g33) & (a) & (!sk[21]) & (!e) & (g34) & (!g35)) + ((!g33) & (a) & (!sk[21]) & (!e) & (g34) & (g35)) + ((!g33) & (a) & (!sk[21]) & (e) & (!g34) & (!g35)) + ((!g33) & (a) & (!sk[21]) & (e) & (!g34) & (g35)) + ((!g33) & (a) & (!sk[21]) & (e) & (g34) & (!g35)) + ((!g33) & (a) & (!sk[21]) & (e) & (g34) & (g35)) + ((!g33) & (a) & (sk[21]) & (!e) & (!g34) & (!g35)) + ((!g33) & (a) & (sk[21]) & (!e) & (g34) & (!g35)) + ((!g33) & (a) & (sk[21]) & (e) & (!g34) & (!g35)) + ((g33) & (!a) & (!sk[21]) & (!e) & (!g34) & (!g35)) + ((g33) & (!a) & (!sk[21]) & (!e) & (!g34) & (g35)) + ((g33) & (!a) & (!sk[21]) & (!e) & (g34) & (!g35)) + ((g33) & (!a) & (!sk[21]) & (!e) & (g34) & (g35)) + ((g33) & (!a) & (!sk[21]) & (e) & (!g34) & (!g35)) + ((g33) & (!a) & (!sk[21]) & (e) & (!g34) & (g35)) + ((g33) & (!a) & (!sk[21]) & (e) & (g34) & (!g35)) + ((g33) & (!a) & (!sk[21]) & (e) & (g34) & (g35)) + ((g33) & (a) & (!sk[21]) & (!e) & (!g34) & (!g35)) + ((g33) & (a) & (!sk[21]) & (!e) & (!g34) & (g35)) + ((g33) & (a) & (!sk[21]) & (!e) & (g34) & (!g35)) + ((g33) & (a) & (!sk[21]) & (!e) & (g34) & (g35)) + ((g33) & (a) & (!sk[21]) & (e) & (!g34) & (!g35)) + ((g33) & (a) & (!sk[21]) & (e) & (!g34) & (g35)) + ((g33) & (a) & (!sk[21]) & (e) & (g34) & (!g35)) + ((g33) & (a) & (!sk[21]) & (e) & (g34) & (g35)));
	assign g39 = (((!a) & (!e) & (!g1) & (!sk[7]) & (!f) & (b)) + ((!a) & (!e) & (!g1) & (!sk[7]) & (f) & (!b)) + ((!a) & (!e) & (!g1) & (!sk[7]) & (f) & (b)) + ((!a) & (!e) & (!g1) & (sk[7]) & (!f) & (b)) + ((!a) & (!e) & (g1) & (!sk[7]) & (!f) & (b)) + ((!a) & (!e) & (g1) & (!sk[7]) & (f) & (!b)) + ((!a) & (!e) & (g1) & (!sk[7]) & (f) & (b)) + ((!a) & (!e) & (g1) & (sk[7]) & (!f) & (b)) + ((!a) & (!e) & (g1) & (sk[7]) & (f) & (!b)) + ((!a) & (e) & (!g1) & (!sk[7]) & (!f) & (b)) + ((!a) & (e) & (!g1) & (!sk[7]) & (f) & (!b)) + ((!a) & (e) & (!g1) & (!sk[7]) & (f) & (b)) + ((!a) & (e) & (!g1) & (sk[7]) & (!f) & (!b)) + ((!a) & (e) & (g1) & (!sk[7]) & (!f) & (b)) + ((!a) & (e) & (g1) & (!sk[7]) & (f) & (!b)) + ((!a) & (e) & (g1) & (!sk[7]) & (f) & (b)) + ((!a) & (e) & (g1) & (sk[7]) & (!f) & (!b)) + ((a) & (!e) & (!g1) & (!sk[7]) & (!f) & (!b)) + ((a) & (!e) & (!g1) & (!sk[7]) & (!f) & (b)) + ((a) & (!e) & (!g1) & (!sk[7]) & (f) & (!b)) + ((a) & (!e) & (!g1) & (!sk[7]) & (f) & (b)) + ((a) & (!e) & (!g1) & (sk[7]) & (!f) & (b)) + ((a) & (!e) & (g1) & (!sk[7]) & (!f) & (!b)) + ((a) & (!e) & (g1) & (!sk[7]) & (!f) & (b)) + ((a) & (!e) & (g1) & (!sk[7]) & (f) & (!b)) + ((a) & (!e) & (g1) & (!sk[7]) & (f) & (b)) + ((a) & (!e) & (g1) & (sk[7]) & (!f) & (b)) + ((a) & (!e) & (g1) & (sk[7]) & (f) & (!b)) + ((a) & (e) & (!g1) & (!sk[7]) & (!f) & (!b)) + ((a) & (e) & (!g1) & (!sk[7]) & (!f) & (b)) + ((a) & (e) & (!g1) & (!sk[7]) & (f) & (!b)) + ((a) & (e) & (!g1) & (!sk[7]) & (f) & (b)) + ((a) & (e) & (!g1) & (sk[7]) & (!f) & (b)) + ((a) & (e) & (g1) & (!sk[7]) & (!f) & (!b)) + ((a) & (e) & (g1) & (!sk[7]) & (!f) & (b)) + ((a) & (e) & (g1) & (!sk[7]) & (f) & (!b)) + ((a) & (e) & (g1) & (!sk[7]) & (f) & (b)) + ((a) & (e) & (g1) & (sk[7]) & (!f) & (b)) + ((a) & (e) & (g1) & (sk[7]) & (f) & (!b)));
	assign g40 = (((!g2) & (sk[7]) & (g3) & (!f) & (!b)) + ((!g2) & (sk[7]) & (g3) & (f) & (!b)) + ((g2) & (!sk[7]) & (!g3) & (f) & (!b)) + ((g2) & (!sk[7]) & (!g3) & (f) & (b)) + ((g2) & (!sk[7]) & (g3) & (!f) & (!b)) + ((g2) & (!sk[7]) & (g3) & (!f) & (b)) + ((g2) & (!sk[7]) & (g3) & (f) & (!b)) + ((g2) & (!sk[7]) & (g3) & (f) & (b)) + ((g2) & (sk[7]) & (!g3) & (!f) & (!b)) + ((g2) & (sk[7]) & (!g3) & (!f) & (b)) + ((g2) & (sk[7]) & (g3) & (!f) & (!b)) + ((g2) & (sk[7]) & (g3) & (!f) & (b)) + ((g2) & (sk[7]) & (g3) & (f) & (!b)));
	assign g42 = (((!n) & (!i) & (sk[11]) & (!a) & (!e) & (g1)) + ((!n) & (!i) & (sk[11]) & (!a) & (e) & (!g1)) + ((!n) & (!i) & (sk[11]) & (!a) & (e) & (g1)) + ((!n) & (!i) & (sk[11]) & (a) & (!e) & (!g1)) + ((!n) & (!i) & (sk[11]) & (a) & (!e) & (g1)) + ((!n) & (!i) & (sk[11]) & (a) & (e) & (!g1)) + ((!n) & (!i) & (sk[11]) & (a) & (e) & (g1)) + ((!n) & (i) & (sk[11]) & (!a) & (!e) & (g1)) + ((!n) & (i) & (sk[11]) & (!a) & (e) & (!g1)) + ((!n) & (i) & (sk[11]) & (!a) & (e) & (g1)) + ((!n) & (i) & (sk[11]) & (a) & (!e) & (!g1)) + ((!n) & (i) & (sk[11]) & (a) & (!e) & (g1)) + ((!n) & (i) & (sk[11]) & (a) & (e) & (!g1)) + ((!n) & (i) & (sk[11]) & (a) & (e) & (g1)) + ((n) & (!i) & (!sk[11]) & (!a) & (e) & (g1)) + ((n) & (!i) & (sk[11]) & (!a) & (!e) & (g1)) + ((n) & (!i) & (sk[11]) & (!a) & (e) & (!g1)) + ((n) & (!i) & (sk[11]) & (!a) & (e) & (g1)) + ((n) & (!i) & (sk[11]) & (a) & (!e) & (!g1)) + ((n) & (!i) & (sk[11]) & (a) & (!e) & (g1)) + ((n) & (!i) & (sk[11]) & (a) & (e) & (!g1)) + ((n) & (!i) & (sk[11]) & (a) & (e) & (g1)) + ((n) & (i) & (sk[11]) & (!a) & (!e) & (g1)) + ((n) & (i) & (sk[11]) & (!a) & (e) & (!g1)) + ((n) & (i) & (sk[11]) & (!a) & (e) & (g1)) + ((n) & (i) & (sk[11]) & (a) & (!e) & (!g1)) + ((n) & (i) & (sk[11]) & (a) & (!e) & (g1)) + ((n) & (i) & (sk[11]) & (a) & (e) & (!g1)) + ((n) & (i) & (sk[11]) & (a) & (e) & (g1)));
	assign g43 = (((!g4) & (!f) & (!b) & (g41) & (!sk[7]) & (!g42)) + ((!g4) & (!f) & (!b) & (g41) & (!sk[7]) & (g42)) + ((!g4) & (!f) & (b) & (!g41) & (!sk[7]) & (g42)) + ((!g4) & (!f) & (b) & (g41) & (!sk[7]) & (!g42)) + ((!g4) & (!f) & (b) & (g41) & (!sk[7]) & (g42)) + ((!g4) & (f) & (!b) & (g41) & (!sk[7]) & (!g42)) + ((!g4) & (f) & (!b) & (g41) & (!sk[7]) & (g42)) + ((!g4) & (f) & (b) & (!g41) & (!sk[7]) & (!g42)) + ((!g4) & (f) & (b) & (!g41) & (!sk[7]) & (g42)) + ((!g4) & (f) & (b) & (!g41) & (sk[7]) & (g42)) + ((!g4) & (f) & (b) & (g41) & (!sk[7]) & (!g42)) + ((!g4) & (f) & (b) & (g41) & (!sk[7]) & (g42)) + ((!g4) & (f) & (b) & (g41) & (sk[7]) & (!g42)) + ((!g4) & (f) & (b) & (g41) & (sk[7]) & (g42)) + ((g4) & (!f) & (!b) & (g41) & (!sk[7]) & (!g42)) + ((g4) & (!f) & (!b) & (g41) & (!sk[7]) & (g42)) + ((g4) & (!f) & (b) & (!g41) & (!sk[7]) & (g42)) + ((g4) & (!f) & (b) & (!g41) & (sk[7]) & (!g42)) + ((g4) & (!f) & (b) & (!g41) & (sk[7]) & (g42)) + ((g4) & (!f) & (b) & (g41) & (!sk[7]) & (!g42)) + ((g4) & (!f) & (b) & (g41) & (!sk[7]) & (g42)) + ((g4) & (!f) & (b) & (g41) & (sk[7]) & (!g42)) + ((g4) & (!f) & (b) & (g41) & (sk[7]) & (g42)) + ((g4) & (f) & (!b) & (!g41) & (sk[7]) & (!g42)) + ((g4) & (f) & (!b) & (!g41) & (sk[7]) & (g42)) + ((g4) & (f) & (!b) & (g41) & (!sk[7]) & (!g42)) + ((g4) & (f) & (!b) & (g41) & (!sk[7]) & (g42)) + ((g4) & (f) & (!b) & (g41) & (sk[7]) & (!g42)) + ((g4) & (f) & (!b) & (g41) & (sk[7]) & (g42)) + ((g4) & (f) & (b) & (!g41) & (!sk[7]) & (!g42)) + ((g4) & (f) & (b) & (!g41) & (!sk[7]) & (g42)) + ((g4) & (f) & (b) & (!g41) & (sk[7]) & (!g42)) + ((g4) & (f) & (b) & (!g41) & (sk[7]) & (g42)) + ((g4) & (f) & (b) & (g41) & (!sk[7]) & (!g42)) + ((g4) & (f) & (b) & (g41) & (!sk[7]) & (g42)) + ((g4) & (f) & (b) & (g41) & (sk[7]) & (!g42)) + ((g4) & (f) & (b) & (g41) & (sk[7]) & (g42)));
	assign g45 = (((!sk[21]) & (!g7) & (f)) + ((!sk[21]) & (g7) & (f)) + ((sk[21]) & (g7) & (f)));
	assign g49 = (((!k) & (l) & (!i) & (j) & (a) & (e)));
	assign g52 = (((!g50) & (!sk[16]) & (!b) & (!g44) & (g51)) + ((!g50) & (!sk[16]) & (!b) & (g44) & (!g51)) + ((!g50) & (!sk[16]) & (!b) & (g44) & (g51)) + ((!g50) & (!sk[16]) & (b) & (!g44) & (g51)) + ((!g50) & (!sk[16]) & (b) & (g44) & (!g51)) + ((!g50) & (!sk[16]) & (b) & (g44) & (g51)) + ((g50) & (!sk[16]) & (!b) & (!g44) & (!g51)) + ((g50) & (!sk[16]) & (!b) & (!g44) & (g51)) + ((g50) & (!sk[16]) & (!b) & (g44) & (!g51)) + ((g50) & (!sk[16]) & (!b) & (g44) & (g51)) + ((g50) & (!sk[16]) & (b) & (!g44) & (!g51)) + ((g50) & (!sk[16]) & (b) & (!g44) & (g51)) + ((g50) & (!sk[16]) & (b) & (g44) & (!g51)) + ((g50) & (!sk[16]) & (b) & (g44) & (g51)) + ((g50) & (sk[16]) & (!b) & (!g44) & (g51)));
	assign g61 = (((!l) & (!a) & (!sk[15]) & (!g14) & (!b) & (!g46)) + ((!l) & (!a) & (!sk[15]) & (!g14) & (b) & (!g46)) + ((!l) & (!a) & (!sk[15]) & (g14) & (!b) & (g46)) + ((!l) & (!a) & (!sk[15]) & (g14) & (b) & (g46)) + ((!l) & (a) & (!sk[15]) & (!g14) & (!b) & (!g46)) + ((!l) & (a) & (!sk[15]) & (!g14) & (b) & (!g46)) + ((!l) & (a) & (!sk[15]) & (g14) & (!b) & (g46)) + ((!l) & (a) & (!sk[15]) & (g14) & (b) & (g46)) + ((l) & (!a) & (!sk[15]) & (!g14) & (!b) & (!g46)) + ((l) & (!a) & (!sk[15]) & (!g14) & (!b) & (g46)) + ((l) & (!a) & (!sk[15]) & (g14) & (!b) & (!g46)) + ((l) & (!a) & (!sk[15]) & (g14) & (!b) & (g46)) + ((l) & (a) & (!sk[15]) & (!g14) & (b) & (!g46)) + ((l) & (a) & (!sk[15]) & (!g14) & (b) & (g46)) + ((l) & (a) & (!sk[15]) & (g14) & (b) & (!g46)) + ((l) & (a) & (!sk[15]) & (g14) & (b) & (g46)));
	assign g63 = (((!k) & (!i) & (!sk[10]) & (g22) & (!f)) + ((!k) & (!i) & (!sk[10]) & (g22) & (f)) + ((!k) & (i) & (!sk[10]) & (g22) & (!f)) + ((!k) & (i) & (!sk[10]) & (g22) & (f)) + ((!k) & (i) & (sk[10]) & (g22) & (f)) + ((k) & (!i) & (!sk[10]) & (!g22) & (!f)) + ((k) & (!i) & (!sk[10]) & (!g22) & (f)) + ((k) & (!i) & (!sk[10]) & (g22) & (!f)) + ((k) & (!i) & (!sk[10]) & (g22) & (f)) + ((k) & (i) & (!sk[10]) & (!g22) & (!f)) + ((k) & (i) & (!sk[10]) & (!g22) & (f)) + ((k) & (i) & (!sk[10]) & (g22) & (!f)) + ((k) & (i) & (!sk[10]) & (g22) & (f)));
	assign g64 = (((!l) & (!a) & (!e) & (sk[7]) & (!f) & (b)) + ((!l) & (!a) & (!e) & (sk[7]) & (f) & (!b)) + ((!l) & (!a) & (e) & (sk[7]) & (!f) & (b)) + ((!l) & (!a) & (e) & (sk[7]) & (f) & (!b)) + ((!l) & (a) & (!e) & (!sk[7]) & (!f) & (!b)) + ((!l) & (a) & (!e) & (!sk[7]) & (!f) & (b)) + ((!l) & (a) & (!e) & (!sk[7]) & (f) & (!b)) + ((!l) & (a) & (!e) & (!sk[7]) & (f) & (b)) + ((!l) & (a) & (!e) & (sk[7]) & (!f) & (b)) + ((!l) & (a) & (!e) & (sk[7]) & (f) & (!b)) + ((!l) & (a) & (e) & (!sk[7]) & (!f) & (!b)) + ((!l) & (a) & (e) & (!sk[7]) & (!f) & (b)) + ((!l) & (a) & (e) & (!sk[7]) & (f) & (!b)) + ((!l) & (a) & (e) & (!sk[7]) & (f) & (b)) + ((!l) & (a) & (e) & (sk[7]) & (f) & (b)) + ((l) & (!a) & (!e) & (!sk[7]) & (!f) & (!b)) + ((l) & (!a) & (!e) & (!sk[7]) & (!f) & (b)) + ((l) & (!a) & (!e) & (!sk[7]) & (f) & (!b)) + ((l) & (!a) & (!e) & (!sk[7]) & (f) & (b)) + ((l) & (!a) & (!e) & (sk[7]) & (!f) & (b)) + ((l) & (!a) & (!e) & (sk[7]) & (f) & (!b)) + ((l) & (!a) & (e) & (!sk[7]) & (!f) & (!b)) + ((l) & (!a) & (e) & (!sk[7]) & (!f) & (b)) + ((l) & (!a) & (e) & (!sk[7]) & (f) & (!b)) + ((l) & (!a) & (e) & (!sk[7]) & (f) & (b)) + ((l) & (!a) & (e) & (sk[7]) & (!f) & (b)) + ((l) & (!a) & (e) & (sk[7]) & (f) & (!b)) + ((l) & (a) & (!e) & (!sk[7]) & (!f) & (!b)) + ((l) & (a) & (!e) & (!sk[7]) & (!f) & (b)) + ((l) & (a) & (!e) & (!sk[7]) & (f) & (!b)) + ((l) & (a) & (!e) & (!sk[7]) & (f) & (b)) + ((l) & (a) & (!e) & (sk[7]) & (!f) & (b)) + ((l) & (a) & (!e) & (sk[7]) & (f) & (!b)) + ((l) & (a) & (e) & (!sk[7]) & (!f) & (!b)) + ((l) & (a) & (e) & (!sk[7]) & (!f) & (b)) + ((l) & (a) & (e) & (!sk[7]) & (f) & (!b)) + ((l) & (a) & (e) & (!sk[7]) & (f) & (b)) + ((l) & (a) & (e) & (sk[7]) & (!f) & (!b)) + ((l) & (a) & (e) & (sk[7]) & (f) & (b)));
	assign g66 = (((!sk[19]) & (!g27) & (!g62) & (!g63) & (!g64) & (!g65)) + ((!sk[19]) & (!g27) & (!g62) & (!g63) & (!g64) & (g65)) + ((!sk[19]) & (!g27) & (!g62) & (!g63) & (g64) & (!g65)) + ((!sk[19]) & (!g27) & (g62) & (!g63) & (!g64) & (!g65)) + ((!sk[19]) & (!g27) & (g62) & (!g63) & (!g64) & (g65)) + ((!sk[19]) & (!g27) & (g62) & (!g63) & (g64) & (!g65)) + ((!sk[19]) & (g27) & (!g62) & (!g63) & (!g64) & (!g65)) + ((!sk[19]) & (g27) & (!g62) & (!g63) & (!g64) & (g65)) + ((!sk[19]) & (g27) & (!g62) & (!g63) & (g64) & (!g65)));
	assign g69 = (((!sk[15]) & (l) & (!i) & (a) & (e)) + ((sk[15]) & (!l) & (!i) & (!a) & (e)) + ((sk[15]) & (!l) & (!i) & (a) & (e)) + ((sk[15]) & (!l) & (i) & (!a) & (e)) + ((sk[15]) & (!l) & (i) & (a) & (e)) + ((sk[15]) & (l) & (!i) & (!a) & (e)) + ((sk[15]) & (l) & (!i) & (a) & (!e)) + ((sk[15]) & (l) & (!i) & (a) & (e)) + ((sk[15]) & (l) & (i) & (!a) & (e)) + ((sk[15]) & (l) & (i) & (a) & (!e)) + ((sk[15]) & (l) & (i) & (a) & (e)));
	assign g70 = (((!g7) & (!g67) & (!g46) & (!g47) & (g68) & (!g69)) + ((!g7) & (!g67) & (!g46) & (!g47) & (g68) & (g69)) + ((!g7) & (!g67) & (!g46) & (g47) & (!g68) & (g69)) + ((!g7) & (!g67) & (!g46) & (g47) & (g68) & (g69)) + ((!g7) & (!g67) & (g46) & (g47) & (g68) & (!g69)) + ((!g7) & (!g67) & (g46) & (g47) & (g68) & (g69)) + ((!g7) & (g67) & (!g46) & (g47) & (!g68) & (g69)) + ((!g7) & (g67) & (!g46) & (g47) & (g68) & (g69)) + ((g7) & (!g67) & (!g46) & (!g47) & (g68) & (!g69)) + ((g7) & (!g67) & (!g46) & (!g47) & (g68) & (g69)) + ((g7) & (!g67) & (!g46) & (g47) & (!g68) & (g69)) + ((g7) & (!g67) & (!g46) & (g47) & (g68) & (g69)) + ((g7) & (!g67) & (g46) & (!g47) & (g68) & (!g69)) + ((g7) & (!g67) & (g46) & (!g47) & (g68) & (g69)) + ((g7) & (!g67) & (g46) & (g47) & (g68) & (!g69)) + ((g7) & (!g67) & (g46) & (g47) & (g68) & (g69)) + ((g7) & (g67) & (!g46) & (g47) & (!g68) & (g69)) + ((g7) & (g67) & (!g46) & (g47) & (g68) & (g69)));
	assign g71 = (((!k) & (!a) & (!g14) & (g26) & (b) & (g46)) + ((!k) & (!a) & (g14) & (g26) & (b) & (g46)) + ((!k) & (a) & (!g14) & (g26) & (b) & (!g46)) + ((!k) & (a) & (g14) & (g26) & (b) & (g46)) + ((k) & (!a) & (!g14) & (g26) & (!b) & (!g46)) + ((k) & (!a) & (!g14) & (g26) & (b) & (g46)) + ((k) & (!a) & (g14) & (g26) & (!b) & (!g46)) + ((k) & (!a) & (g14) & (g26) & (b) & (g46)) + ((k) & (a) & (!g14) & (g26) & (!b) & (g46)) + ((k) & (a) & (!g14) & (g26) & (b) & (!g46)) + ((k) & (a) & (g14) & (g26) & (!b) & (!g46)) + ((k) & (a) & (g14) & (g26) & (b) & (g46)));
	assign g73 = (((!sk[13]) & (!g58) & (!g59) & (g72)) + ((sk[13]) & (g58) & (!g59) & (!g72)) + ((sk[13]) & (g58) & (!g59) & (g72)) + ((sk[13]) & (g58) & (g59) & (!g72)) + ((sk[13]) & (g58) & (g59) & (g72)));
	assign g74 = (((!k) & (!l) & (!i) & (!f) & (!b) & (!g44)) + ((!k) & (!l) & (!i) & (!f) & (b) & (!g44)) + ((!k) & (!l) & (!i) & (f) & (!b) & (!g44)) + ((!k) & (!l) & (!i) & (f) & (b) & (!g44)) + ((!k) & (!l) & (i) & (!f) & (!b) & (g44)) + ((!k) & (!l) & (i) & (!f) & (b) & (g44)) + ((!k) & (!l) & (i) & (f) & (!b) & (g44)) + ((!k) & (!l) & (i) & (f) & (b) & (g44)) + ((!k) & (l) & (!i) & (!f) & (!b) & (!g44)) + ((!k) & (l) & (!i) & (f) & (!b) & (!g44)) + ((!k) & (l) & (!i) & (f) & (b) & (!g44)) + ((!k) & (l) & (i) & (!f) & (!b) & (!g44)) + ((!k) & (l) & (i) & (!f) & (!b) & (g44)) + ((!k) & (l) & (i) & (f) & (b) & (!g44)) + ((!k) & (l) & (i) & (f) & (b) & (g44)) + ((k) & (!l) & (!i) & (!f) & (!b) & (g44)) + ((k) & (!l) & (!i) & (!f) & (b) & (g44)) + ((k) & (!l) & (!i) & (f) & (!b) & (g44)) + ((k) & (!l) & (!i) & (f) & (b) & (g44)) + ((k) & (!l) & (i) & (f) & (!b) & (!g44)) + ((k) & (!l) & (i) & (f) & (!b) & (g44)) + ((k) & (!l) & (i) & (f) & (b) & (!g44)) + ((k) & (!l) & (i) & (f) & (b) & (g44)) + ((k) & (l) & (i) & (!f) & (!b) & (!g44)) + ((k) & (l) & (i) & (f) & (!b) & (!g44)) + ((k) & (l) & (i) & (f) & (b) & (!g44)));
	assign g75 = (((!k) & (l) & (!i) & (f) & (!b) & (!g44)) + ((!k) & (l) & (!i) & (f) & (!b) & (g44)) + ((!k) & (l) & (!i) & (f) & (b) & (!g44)) + ((!k) & (l) & (!i) & (f) & (b) & (g44)) + ((k) & (!l) & (!i) & (!f) & (!b) & (!g44)) + ((k) & (!l) & (!i) & (!f) & (!b) & (g44)) + ((k) & (!l) & (i) & (!f) & (b) & (g44)) + ((k) & (!l) & (i) & (f) & (b) & (g44)) + ((k) & (l) & (!i) & (f) & (!b) & (!g44)) + ((k) & (l) & (!i) & (f) & (!b) & (g44)) + ((k) & (l) & (!i) & (f) & (b) & (!g44)) + ((k) & (l) & (!i) & (f) & (b) & (g44)) + ((k) & (l) & (i) & (!f) & (b) & (g44)) + ((k) & (l) & (i) & (f) & (b) & (g44)));
	assign g76 = (((!g34) & (!sk[18]) & (!g35) & (!f) & (b)) + ((!g34) & (!sk[18]) & (!g35) & (f) & (b)) + ((!g34) & (!sk[18]) & (g35) & (!f) & (!b)) + ((!g34) & (!sk[18]) & (g35) & (!f) & (b)) + ((!g34) & (!sk[18]) & (g35) & (f) & (!b)) + ((!g34) & (!sk[18]) & (g35) & (f) & (b)) + ((!g34) & (sk[18]) & (g35) & (!f) & (b)) + ((!g34) & (sk[18]) & (g35) & (f) & (b)) + ((g34) & (!sk[18]) & (!g35) & (!f) & (!b)) + ((g34) & (!sk[18]) & (!g35) & (!f) & (b)) + ((g34) & (!sk[18]) & (!g35) & (f) & (!b)) + ((g34) & (!sk[18]) & (!g35) & (f) & (b)) + ((g34) & (!sk[18]) & (g35) & (!f) & (!b)) + ((g34) & (!sk[18]) & (g35) & (!f) & (b)) + ((g34) & (!sk[18]) & (g35) & (f) & (!b)) + ((g34) & (!sk[18]) & (g35) & (f) & (b)) + ((g34) & (sk[18]) & (!g35) & (f) & (b)) + ((g34) & (sk[18]) & (g35) & (!f) & (b)) + ((g34) & (sk[18]) & (g35) & (f) & (b)));
	assign g77 = (((!g33) & (!sk[16]) & (!g32) & (f) & (!g44) & (!g76)) + ((!g33) & (!sk[16]) & (!g32) & (f) & (!g44) & (g76)) + ((!g33) & (!sk[16]) & (!g32) & (f) & (g44) & (!g76)) + ((!g33) & (!sk[16]) & (!g32) & (f) & (g44) & (g76)) + ((!g33) & (!sk[16]) & (g32) & (f) & (!g44) & (!g76)) + ((!g33) & (!sk[16]) & (g32) & (f) & (!g44) & (g76)) + ((!g33) & (!sk[16]) & (g32) & (f) & (g44) & (!g76)) + ((!g33) & (!sk[16]) & (g32) & (f) & (g44) & (g76)) + ((!g33) & (sk[16]) & (!g32) & (!f) & (!g44) & (!g76)) + ((!g33) & (sk[16]) & (!g32) & (!f) & (g44) & (!g76)) + ((!g33) & (sk[16]) & (!g32) & (f) & (!g44) & (!g76)) + ((!g33) & (sk[16]) & (!g32) & (f) & (g44) & (!g76)) + ((!g33) & (sk[16]) & (g32) & (!f) & (!g44) & (!g76)) + ((!g33) & (sk[16]) & (g32) & (!f) & (g44) & (!g76)) + ((!g33) & (sk[16]) & (g32) & (f) & (!g44) & (!g76)) + ((g33) & (!sk[16]) & (!g32) & (!f) & (!g44) & (!g76)) + ((g33) & (!sk[16]) & (!g32) & (!f) & (!g44) & (g76)) + ((g33) & (!sk[16]) & (!g32) & (!f) & (g44) & (!g76)) + ((g33) & (!sk[16]) & (!g32) & (!f) & (g44) & (g76)) + ((g33) & (!sk[16]) & (!g32) & (f) & (!g44) & (!g76)) + ((g33) & (!sk[16]) & (!g32) & (f) & (!g44) & (g76)) + ((g33) & (!sk[16]) & (!g32) & (f) & (g44) & (!g76)) + ((g33) & (!sk[16]) & (!g32) & (f) & (g44) & (g76)) + ((g33) & (!sk[16]) & (g32) & (!f) & (!g44) & (!g76)) + ((g33) & (!sk[16]) & (g32) & (!f) & (!g44) & (g76)) + ((g33) & (!sk[16]) & (g32) & (!f) & (g44) & (!g76)) + ((g33) & (!sk[16]) & (g32) & (!f) & (g44) & (g76)) + ((g33) & (!sk[16]) & (g32) & (f) & (!g44) & (!g76)) + ((g33) & (!sk[16]) & (g32) & (f) & (!g44) & (g76)) + ((g33) & (!sk[16]) & (g32) & (f) & (g44) & (!g76)) + ((g33) & (!sk[16]) & (g32) & (f) & (g44) & (g76)));
	assign g78 = (((!n) & (!j) & (!g74) & (!g75) & (!sk[22]) & (g77)) + ((!n) & (!j) & (!g74) & (g75) & (!sk[22]) & (g77)) + ((!n) & (!j) & (g74) & (!g75) & (!sk[22]) & (!g77)) + ((!n) & (!j) & (g74) & (!g75) & (!sk[22]) & (g77)) + ((!n) & (!j) & (g74) & (!g75) & (sk[22]) & (g77)) + ((!n) & (!j) & (g74) & (g75) & (!sk[22]) & (!g77)) + ((!n) & (!j) & (g74) & (g75) & (!sk[22]) & (g77)) + ((!n) & (!j) & (g74) & (g75) & (sk[22]) & (g77)) + ((!n) & (j) & (!g74) & (!g75) & (!sk[22]) & (g77)) + ((!n) & (j) & (!g74) & (!g75) & (sk[22]) & (g77)) + ((!n) & (j) & (!g74) & (g75) & (!sk[22]) & (g77)) + ((!n) & (j) & (g74) & (!g75) & (!sk[22]) & (!g77)) + ((!n) & (j) & (g74) & (!g75) & (!sk[22]) & (g77)) + ((!n) & (j) & (g74) & (!g75) & (sk[22]) & (g77)) + ((!n) & (j) & (g74) & (g75) & (!sk[22]) & (!g77)) + ((!n) & (j) & (g74) & (g75) & (!sk[22]) & (g77)) + ((n) & (!j) & (!g74) & (!g75) & (!sk[22]) & (g77)) + ((n) & (!j) & (!g74) & (!g75) & (sk[22]) & (g77)) + ((n) & (!j) & (!g74) & (g75) & (!sk[22]) & (g77)) + ((n) & (!j) & (!g74) & (g75) & (sk[22]) & (g77)) + ((n) & (!j) & (g74) & (!g75) & (!sk[22]) & (!g77)) + ((n) & (!j) & (g74) & (!g75) & (!sk[22]) & (g77)) + ((n) & (!j) & (g74) & (!g75) & (sk[22]) & (g77)) + ((n) & (!j) & (g74) & (g75) & (!sk[22]) & (!g77)) + ((n) & (!j) & (g74) & (g75) & (!sk[22]) & (g77)) + ((n) & (!j) & (g74) & (g75) & (sk[22]) & (g77)) + ((n) & (j) & (!g74) & (!g75) & (!sk[22]) & (g77)) + ((n) & (j) & (!g74) & (!g75) & (sk[22]) & (g77)) + ((n) & (j) & (!g74) & (g75) & (!sk[22]) & (g77)) + ((n) & (j) & (!g74) & (g75) & (sk[22]) & (g77)) + ((n) & (j) & (g74) & (!g75) & (!sk[22]) & (!g77)) + ((n) & (j) & (g74) & (!g75) & (!sk[22]) & (g77)) + ((n) & (j) & (g74) & (!g75) & (sk[22]) & (g77)) + ((n) & (j) & (g74) & (g75) & (!sk[22]) & (!g77)) + ((n) & (j) & (g74) & (g75) & (!sk[22]) & (g77)) + ((n) & (j) & (g74) & (g75) & (sk[22]) & (g77)));
	assign g83 = (((!j) & (!g1) & (!c) & (!sk[22]) & (g)) + ((!j) & (!g1) & (c) & (!sk[22]) & (g)) + ((!j) & (g1) & (!c) & (!sk[22]) & (g)) + ((!j) & (g1) & (c) & (!sk[22]) & (g)) + ((!j) & (g1) & (c) & (sk[22]) & (g)) + ((j) & (!g1) & (!c) & (!sk[22]) & (g)) + ((j) & (!g1) & (!c) & (sk[22]) & (!g)) + ((j) & (!g1) & (c) & (!sk[22]) & (!g)) + ((j) & (!g1) & (c) & (!sk[22]) & (g)) + ((j) & (g1) & (!c) & (!sk[22]) & (g)) + ((j) & (g1) & (!c) & (sk[22]) & (!g)) + ((j) & (g1) & (c) & (!sk[22]) & (!g)) + ((j) & (g1) & (c) & (!sk[22]) & (g)) + ((j) & (g1) & (c) & (sk[22]) & (g)));
	assign g84 = (((!n) & (!sk[23]) & (!i) & (!g81) & (g83)) + ((!n) & (!sk[23]) & (!i) & (g81) & (!g83)) + ((!n) & (!sk[23]) & (!i) & (g81) & (g83)) + ((!n) & (!sk[23]) & (i) & (!g81) & (g83)) + ((!n) & (!sk[23]) & (i) & (g81) & (!g83)) + ((!n) & (!sk[23]) & (i) & (g81) & (g83)) + ((n) & (!sk[23]) & (!i) & (!g81) & (g83)) + ((n) & (!sk[23]) & (!i) & (g81) & (!g83)) + ((n) & (!sk[23]) & (!i) & (g81) & (g83)) + ((n) & (!sk[23]) & (i) & (!g81) & (g83)) + ((n) & (!sk[23]) & (i) & (g81) & (!g83)) + ((n) & (!sk[23]) & (i) & (g81) & (g83)) + ((n) & (sk[23]) & (!i) & (g81) & (g83)));
	assign g85 = (((!g2) & (!g3) & (sk[24]) & (!c) & (g)) + ((!g2) & (!g3) & (sk[24]) & (c) & (g)) + ((!g2) & (g3) & (!sk[24]) & (!c) & (!g)) + ((!g2) & (g3) & (!sk[24]) & (!c) & (g)) + ((!g2) & (g3) & (sk[24]) & (!c) & (g)) + ((!g2) & (g3) & (sk[24]) & (c) & (g)) + ((g2) & (!g3) & (!sk[24]) & (!c) & (!g)) + ((g2) & (!g3) & (!sk[24]) & (c) & (!g)) + ((g2) & (!g3) & (sk[24]) & (!c) & (!g)) + ((g2) & (!g3) & (sk[24]) & (!c) & (g)) + ((g2) & (!g3) & (sk[24]) & (c) & (!g)) + ((g2) & (!g3) & (sk[24]) & (c) & (g)) + ((g2) & (g3) & (!sk[24]) & (!c) & (!g)) + ((g2) & (g3) & (!sk[24]) & (!c) & (g)) + ((g2) & (g3) & (!sk[24]) & (c) & (!g)) + ((g2) & (g3) & (sk[24]) & (!c) & (!g)) + ((g2) & (g3) & (sk[24]) & (!c) & (g)) + ((g2) & (g3) & (sk[24]) & (c) & (!g)) + ((g2) & (g3) & (sk[24]) & (c) & (g)));
	assign g86 = (((!g4) & (!sk[24]) & (g41) & (c) & (g)) + ((!g4) & (sk[24]) & (!g41) & (c) & (!g)) + ((!g4) & (sk[24]) & (!g41) & (c) & (g)) + ((!g4) & (sk[24]) & (g41) & (c) & (!g)) + ((!g4) & (sk[24]) & (g41) & (c) & (g)) + ((g4) & (!sk[24]) & (!g41) & (!c) & (g)) + ((g4) & (!sk[24]) & (!g41) & (c) & (!g)) + ((g4) & (!sk[24]) & (!g41) & (c) & (g)) + ((g4) & (!sk[24]) & (g41) & (!c) & (g)) + ((g4) & (!sk[24]) & (g41) & (c) & (!g)) + ((g4) & (!sk[24]) & (g41) & (c) & (g)) + ((g4) & (sk[24]) & (!g41) & (c) & (!g)) + ((g4) & (sk[24]) & (!g41) & (c) & (g)) + ((g4) & (sk[24]) & (g41) & (c) & (!g)) + ((g4) & (sk[24]) & (g41) & (c) & (g)));
	assign g88 = (((!g9) & (!sk[24]) & (!g12) & (!c)) + ((!g9) & (!sk[24]) & (!g12) & (c)) + ((g9) & (!sk[24]) & (!g12) & (!c)));
	assign g89 = (((!g7) & (!g12) & (c) & (sk[24]) & (g)) + ((!g7) & (g12) & (c) & (!sk[24]) & (!g)) + ((!g7) & (g12) & (c) & (!sk[24]) & (g)) + ((!g7) & (g12) & (c) & (sk[24]) & (g)) + ((g7) & (!g12) & (!c) & (sk[24]) & (!g)) + ((g7) & (!g12) & (!c) & (sk[24]) & (g)) + ((g7) & (!g12) & (c) & (!sk[24]) & (g)) + ((g7) & (!g12) & (c) & (sk[24]) & (!g)) + ((g7) & (!g12) & (c) & (sk[24]) & (g)) + ((g7) & (g12) & (!c) & (sk[24]) & (!g)) + ((g7) & (g12) & (!c) & (sk[24]) & (g)) + ((g7) & (g12) & (c) & (!sk[24]) & (!g)) + ((g7) & (g12) & (c) & (!sk[24]) & (g)) + ((g7) & (g12) & (c) & (sk[24]) & (!g)) + ((g7) & (g12) & (c) & (sk[24]) & (g)));
	assign g94 = (((!n) & (!g53) & (!g57) & (sk[19]) & (!g92) & (g93)) + ((!n) & (!g53) & (!g57) & (sk[19]) & (g92) & (g93)) + ((!n) & (!g53) & (g57) & (sk[19]) & (!g92) & (!g93)) + ((!n) & (!g53) & (g57) & (sk[19]) & (!g92) & (g93)) + ((!n) & (!g53) & (g57) & (sk[19]) & (g92) & (!g93)) + ((!n) & (!g53) & (g57) & (sk[19]) & (g92) & (g93)) + ((!n) & (g53) & (!g57) & (sk[19]) & (!g92) & (!g93)) + ((!n) & (g53) & (!g57) & (sk[19]) & (!g92) & (g93)) + ((!n) & (g53) & (!g57) & (sk[19]) & (g92) & (!g93)) + ((!n) & (g53) & (!g57) & (sk[19]) & (g92) & (g93)) + ((!n) & (g53) & (g57) & (sk[19]) & (!g92) & (!g93)) + ((!n) & (g53) & (g57) & (sk[19]) & (!g92) & (g93)) + ((!n) & (g53) & (g57) & (sk[19]) & (g92) & (!g93)) + ((!n) & (g53) & (g57) & (sk[19]) & (g92) & (g93)) + ((n) & (!g53) & (!g57) & (sk[19]) & (!g92) & (g93)) + ((n) & (!g53) & (!g57) & (sk[19]) & (g92) & (g93)) + ((n) & (!g53) & (g57) & (!sk[19]) & (!g92) & (!g93)) + ((n) & (!g53) & (g57) & (!sk[19]) & (!g92) & (g93)) + ((n) & (!g53) & (g57) & (!sk[19]) & (g92) & (!g93)) + ((n) & (!g53) & (g57) & (!sk[19]) & (g92) & (g93)) + ((n) & (!g53) & (g57) & (sk[19]) & (!g92) & (!g93)) + ((n) & (!g53) & (g57) & (sk[19]) & (!g92) & (g93)) + ((n) & (!g53) & (g57) & (sk[19]) & (g92) & (!g93)) + ((n) & (!g53) & (g57) & (sk[19]) & (g92) & (g93)) + ((n) & (g53) & (!g57) & (!sk[19]) & (!g92) & (g93)) + ((n) & (g53) & (!g57) & (sk[19]) & (!g92) & (!g93)) + ((n) & (g53) & (!g57) & (sk[19]) & (!g92) & (g93)) + ((n) & (g53) & (!g57) & (sk[19]) & (g92) & (!g93)) + ((n) & (g53) & (!g57) & (sk[19]) & (g92) & (g93)) + ((n) & (g53) & (g57) & (!sk[19]) & (!g92) & (!g93)) + ((n) & (g53) & (g57) & (!sk[19]) & (!g92) & (g93)) + ((n) & (g53) & (g57) & (!sk[19]) & (g92) & (!g93)) + ((n) & (g53) & (g57) & (!sk[19]) & (g92) & (g93)) + ((n) & (g53) & (g57) & (sk[19]) & (!g92) & (!g93)) + ((n) & (g53) & (g57) & (sk[19]) & (!g92) & (g93)) + ((n) & (g53) & (g57) & (sk[19]) & (g92) & (!g93)) + ((n) & (g53) & (g57) & (sk[19]) & (g92) & (g93)));
	assign g95 = (((!sk[17]) & (l) & (!a) & (b) & (g60)) + ((!sk[17]) & (l) & (a) & (!b) & (g60)) + ((!sk[17]) & (l) & (a) & (b) & (g60)) + ((sk[17]) & (!l) & (!a) & (b) & (!g60)) + ((sk[17]) & (!l) & (!a) & (b) & (g60)) + ((sk[17]) & (!l) & (a) & (!b) & (!g60)) + ((sk[17]) & (!l) & (a) & (!b) & (g60)) + ((sk[17]) & (!l) & (a) & (b) & (!g60)) + ((sk[17]) & (!l) & (a) & (b) & (g60)) + ((sk[17]) & (l) & (!a) & (!b) & (!g60)) + ((sk[17]) & (l) & (!a) & (!b) & (g60)) + ((sk[17]) & (l) & (!a) & (b) & (!g60)) + ((sk[17]) & (l) & (!a) & (b) & (g60)) + ((sk[17]) & (l) & (a) & (!b) & (!g60)) + ((sk[17]) & (l) & (a) & (!b) & (g60)) + ((sk[17]) & (l) & (a) & (b) & (!g60)) + ((sk[17]) & (l) & (a) & (b) & (g60)));
	assign g97 = (((!sk[24]) & (!g65) & (!g) & (!g95) & (!g96)) + ((!sk[24]) & (!g65) & (!g) & (!g95) & (g96)) + ((!sk[24]) & (!g65) & (g) & (!g95) & (!g96)) + ((!sk[24]) & (!g65) & (g) & (!g95) & (g96)) + ((!sk[24]) & (g65) & (!g) & (!g95) & (g96)) + ((!sk[24]) & (g65) & (g) & (!g95) & (!g96)));
	assign g98 = (((!g26) & (!sk[25]) & (c) & (!g91) & (!g94) & (!g97)) + ((!g26) & (!sk[25]) & (c) & (!g91) & (g94) & (!g97)) + ((!g26) & (!sk[25]) & (c) & (!g91) & (g94) & (g97)) + ((!g26) & (!sk[25]) & (c) & (g91) & (!g94) & (!g97)) + ((!g26) & (!sk[25]) & (c) & (g91) & (g94) & (!g97)) + ((!g26) & (!sk[25]) & (c) & (g91) & (g94) & (g97)) + ((!g26) & (sk[25]) & (!c) & (!g91) & (!g94) & (g97)) + ((!g26) & (sk[25]) & (!c) & (!g91) & (g94) & (g97)) + ((!g26) & (sk[25]) & (!c) & (g91) & (!g94) & (g97)) + ((!g26) & (sk[25]) & (!c) & (g91) & (g94) & (g97)) + ((!g26) & (sk[25]) & (c) & (!g91) & (!g94) & (!g97)) + ((!g26) & (sk[25]) & (c) & (!g91) & (!g94) & (g97)) + ((!g26) & (sk[25]) & (c) & (!g91) & (g94) & (!g97)) + ((!g26) & (sk[25]) & (c) & (!g91) & (g94) & (g97)) + ((!g26) & (sk[25]) & (c) & (g91) & (!g94) & (!g97)) + ((!g26) & (sk[25]) & (c) & (g91) & (!g94) & (g97)) + ((!g26) & (sk[25]) & (c) & (g91) & (g94) & (!g97)) + ((!g26) & (sk[25]) & (c) & (g91) & (g94) & (g97)) + ((g26) & (!sk[25]) & (c) & (!g91) & (!g94) & (!g97)) + ((g26) & (!sk[25]) & (c) & (!g91) & (!g94) & (g97)) + ((g26) & (!sk[25]) & (c) & (!g91) & (g94) & (!g97)) + ((g26) & (!sk[25]) & (c) & (!g91) & (g94) & (g97)) + ((g26) & (!sk[25]) & (c) & (g91) & (!g94) & (!g97)) + ((g26) & (!sk[25]) & (c) & (g91) & (g94) & (!g97)) + ((g26) & (!sk[25]) & (c) & (g91) & (g94) & (g97)) + ((g26) & (sk[25]) & (!c) & (!g91) & (!g94) & (g97)) + ((g26) & (sk[25]) & (!c) & (!g91) & (g94) & (g97)) + ((g26) & (sk[25]) & (!c) & (g91) & (!g94) & (!g97)) + ((g26) & (sk[25]) & (!c) & (g91) & (!g94) & (g97)) + ((g26) & (sk[25]) & (!c) & (g91) & (g94) & (!g97)) + ((g26) & (sk[25]) & (!c) & (g91) & (g94) & (g97)) + ((g26) & (sk[25]) & (c) & (!g91) & (!g94) & (!g97)) + ((g26) & (sk[25]) & (c) & (!g91) & (!g94) & (g97)) + ((g26) & (sk[25]) & (c) & (!g91) & (g94) & (!g97)) + ((g26) & (sk[25]) & (c) & (!g91) & (g94) & (g97)) + ((g26) & (sk[25]) & (c) & (g91) & (!g94) & (!g97)) + ((g26) & (sk[25]) & (c) & (g91) & (!g94) & (g97)) + ((g26) & (sk[25]) & (c) & (g91) & (g94) & (!g97)) + ((g26) & (sk[25]) & (c) & (g91) & (g94) & (g97)));
	assign g99 = (((!sk[25]) & (!l) & (g65) & (g) & (!g96)) + ((!sk[25]) & (l) & (g65) & (!g) & (g96)) + ((!sk[25]) & (l) & (g65) & (g) & (!g96)) + ((sk[25]) & (l) & (!g65) & (!g) & (!g96)) + ((sk[25]) & (l) & (!g65) & (!g) & (g96)) + ((sk[25]) & (l) & (!g65) & (g) & (!g96)) + ((sk[25]) & (l) & (!g65) & (g) & (g96)) + ((sk[25]) & (l) & (g65) & (!g) & (!g96)) + ((sk[25]) & (l) & (g65) & (!g) & (g96)) + ((sk[25]) & (l) & (g65) & (g) & (!g96)) + ((sk[25]) & (l) & (g65) & (g) & (g96)));
	assign g100 = (((!n) & (!sk[19]) & (!g51) & (!g92) & (!g93) & (!g99)) + ((!n) & (!sk[19]) & (!g51) & (!g92) & (g93) & (!g99)) + ((!n) & (!sk[19]) & (!g51) & (g92) & (!g93) & (!g99)) + ((!n) & (!sk[19]) & (!g51) & (g92) & (g93) & (!g99)) + ((!n) & (!sk[19]) & (g51) & (!g92) & (!g93) & (!g99)) + ((!n) & (!sk[19]) & (g51) & (!g92) & (g93) & (!g99)) + ((!n) & (!sk[19]) & (g51) & (g92) & (!g93) & (!g99)) + ((!n) & (!sk[19]) & (g51) & (g92) & (g93) & (!g99)) + ((n) & (!sk[19]) & (!g51) & (!g92) & (!g93) & (!g99)) + ((n) & (!sk[19]) & (!g51) & (!g92) & (g93) & (!g99)) + ((n) & (!sk[19]) & (!g51) & (g92) & (!g93) & (!g99)) + ((n) & (!sk[19]) & (!g51) & (g92) & (g93) & (!g99)) + ((n) & (!sk[19]) & (g51) & (!g92) & (!g93) & (!g99)) + ((n) & (!sk[19]) & (g51) & (!g92) & (g93) & (!g99)) + ((n) & (!sk[19]) & (g51) & (g92) & (!g93) & (!g99)));
	assign g101 = (((!k) & (!g26) & (!sk[25]) & (!c) & (!g91) & (!g100)) + ((!k) & (!g26) & (!sk[25]) & (!c) & (g91) & (!g100)) + ((!k) & (g26) & (!sk[25]) & (!c) & (!g91) & (!g100)) + ((!k) & (g26) & (!sk[25]) & (!c) & (g91) & (!g100)) + ((k) & (!g26) & (!sk[25]) & (!c) & (!g91) & (!g100)) + ((k) & (!g26) & (!sk[25]) & (!c) & (g91) & (!g100)) + ((k) & (g26) & (!sk[25]) & (!c) & (!g91) & (!g100)) + ((k) & (g26) & (!sk[25]) & (!c) & (g91) & (!g100)) + ((k) & (g26) & (!sk[25]) & (!c) & (g91) & (g100)));
	assign g105 = (((!k) & (g28) & (g) & (!g93) & (!g103) & (!g104)) + ((!k) & (g28) & (g) & (!g93) & (!g103) & (g104)) + ((!k) & (g28) & (g) & (!g93) & (g103) & (!g104)) + ((!k) & (g28) & (g) & (!g93) & (g103) & (g104)) + ((!k) & (g28) & (g) & (g93) & (!g103) & (!g104)) + ((!k) & (g28) & (g) & (g93) & (!g103) & (g104)) + ((!k) & (g28) & (g) & (g93) & (g103) & (!g104)) + ((!k) & (g28) & (g) & (g93) & (g103) & (g104)) + ((k) & (g28) & (!g) & (!g93) & (!g103) & (g104)) + ((k) & (g28) & (!g) & (!g93) & (g103) & (!g104)) + ((k) & (g28) & (!g) & (g93) & (!g103) & (!g104)) + ((k) & (g28) & (!g) & (g93) & (g103) & (g104)) + ((k) & (g28) & (g) & (!g93) & (!g103) & (g104)) + ((k) & (g28) & (g) & (!g93) & (g103) & (!g104)) + ((k) & (g28) & (g) & (g93) & (!g103) & (!g104)) + ((k) & (g28) & (g) & (g93) & (g103) & (g104)));
	assign g107 = (((!g68) & (sk[20]) & (!g90) & (!g103) & (g106)) + ((!g68) & (sk[20]) & (!g90) & (g103) & (g106)) + ((!g68) & (sk[20]) & (g90) & (!g103) & (g106)) + ((!g68) & (sk[20]) & (g90) & (g103) & (g106)) + ((g68) & (!sk[20]) & (!g90) & (!g103) & (!g106)) + ((g68) & (!sk[20]) & (g90) & (!g103) & (g106)) + ((g68) & (sk[20]) & (!g90) & (!g103) & (!g106)) + ((g68) & (sk[20]) & (!g90) & (!g103) & (g106)) + ((g68) & (sk[20]) & (!g90) & (g103) & (!g106)) + ((g68) & (sk[20]) & (!g90) & (g103) & (g106)) + ((g68) & (sk[20]) & (g90) & (!g103) & (!g106)) + ((g68) & (sk[20]) & (g90) & (!g103) & (g106)) + ((g68) & (sk[20]) & (g90) & (g103) & (!g106)) + ((g68) & (sk[20]) & (g90) & (g103) & (g106)));
	assign g108 = (((!l) & (!a) & (!b) & (sk[17]) & (g60) & (!c)) + ((!l) & (!a) & (!b) & (sk[17]) & (g60) & (c)) + ((!l) & (!a) & (b) & (sk[17]) & (g60) & (!c)) + ((!l) & (!a) & (b) & (sk[17]) & (g60) & (c)) + ((!l) & (a) & (!b) & (sk[17]) & (g60) & (!c)) + ((!l) & (a) & (!b) & (sk[17]) & (g60) & (c)) + ((!l) & (a) & (b) & (sk[17]) & (g60) & (!c)) + ((!l) & (a) & (b) & (sk[17]) & (g60) & (c)) + ((l) & (!a) & (!b) & (!sk[17]) & (g60) & (!c)) + ((l) & (!a) & (!b) & (sk[17]) & (g60) & (!c)) + ((l) & (!a) & (!b) & (sk[17]) & (g60) & (c)) + ((l) & (!a) & (b) & (sk[17]) & (g60) & (!c)) + ((l) & (!a) & (b) & (sk[17]) & (g60) & (c)) + ((l) & (a) & (!b) & (sk[17]) & (!g60) & (!c)) + ((l) & (a) & (!b) & (sk[17]) & (!g60) & (c)) + ((l) & (a) & (!b) & (sk[17]) & (g60) & (!c)) + ((l) & (a) & (!b) & (sk[17]) & (g60) & (c)) + ((l) & (a) & (b) & (sk[17]) & (!g60) & (!c)) + ((l) & (a) & (b) & (sk[17]) & (!g60) & (c)) + ((l) & (a) & (b) & (sk[17]) & (g60) & (!c)) + ((l) & (a) & (b) & (sk[17]) & (g60) & (c)));
	assign g110 = (((!l) & (!g14) & (!g46) & (!g60) & (sk[17]) & (g90)) + ((!l) & (!g14) & (!g46) & (g60) & (!sk[17]) & (!g90)) + ((!l) & (!g14) & (!g46) & (g60) & (sk[17]) & (!g90)) + ((!l) & (!g14) & (!g46) & (g60) & (sk[17]) & (g90)) + ((!l) & (!g14) & (g46) & (!g60) & (sk[17]) & (!g90)) + ((!l) & (!g14) & (g46) & (!g60) & (sk[17]) & (g90)) + ((!l) & (!g14) & (g46) & (g60) & (!sk[17]) & (!g90)) + ((!l) & (!g14) & (g46) & (g60) & (sk[17]) & (!g90)) + ((!l) & (!g14) & (g46) & (g60) & (sk[17]) & (g90)) + ((!l) & (g14) & (!g46) & (!g60) & (sk[17]) & (g90)) + ((!l) & (g14) & (!g46) & (g60) & (!sk[17]) & (!g90)) + ((!l) & (g14) & (!g46) & (g60) & (sk[17]) & (!g90)) + ((!l) & (g14) & (!g46) & (g60) & (sk[17]) & (g90)) + ((!l) & (g14) & (g46) & (!g60) & (sk[17]) & (!g90)) + ((!l) & (g14) & (g46) & (!g60) & (sk[17]) & (g90)) + ((!l) & (g14) & (g46) & (g60) & (!sk[17]) & (g90)) + ((!l) & (g14) & (g46) & (g60) & (sk[17]) & (!g90)) + ((!l) & (g14) & (g46) & (g60) & (sk[17]) & (g90)) + ((l) & (!g14) & (!g46) & (!g60) & (sk[17]) & (g90)) + ((l) & (!g14) & (!g46) & (g60) & (sk[17]) & (!g90)) + ((l) & (!g14) & (!g46) & (g60) & (sk[17]) & (g90)) + ((l) & (!g14) & (g46) & (!g60) & (sk[17]) & (!g90)) + ((l) & (!g14) & (g46) & (!g60) & (sk[17]) & (g90)) + ((l) & (!g14) & (g46) & (g60) & (sk[17]) & (!g90)) + ((l) & (!g14) & (g46) & (g60) & (sk[17]) & (g90)) + ((l) & (g14) & (!g46) & (!g60) & (sk[17]) & (g90)) + ((l) & (g14) & (!g46) & (g60) & (sk[17]) & (!g90)) + ((l) & (g14) & (!g46) & (g60) & (sk[17]) & (g90)) + ((l) & (g14) & (g46) & (!g60) & (sk[17]) & (!g90)) + ((l) & (g14) & (g46) & (!g60) & (sk[17]) & (g90)) + ((l) & (g14) & (g46) & (g60) & (sk[17]) & (!g90)) + ((l) & (g14) & (g46) & (g60) & (sk[17]) & (g90)));
	assign g111 = (((!sk[16]) & (!g182) & (!g44) & (!g54) & (g55)) + ((!sk[16]) & (!g182) & (!g44) & (g54) & (g55)) + ((!sk[16]) & (!g182) & (g44) & (!g54) & (!g55)) + ((!sk[16]) & (!g182) & (g44) & (!g54) & (g55)) + ((!sk[16]) & (!g182) & (g44) & (g54) & (!g55)) + ((!sk[16]) & (!g182) & (g44) & (g54) & (g55)) + ((!sk[16]) & (g182) & (!g44) & (!g54) & (g55)) + ((!sk[16]) & (g182) & (!g44) & (g54) & (g55)) + ((!sk[16]) & (g182) & (g44) & (!g54) & (!g55)) + ((!sk[16]) & (g182) & (g44) & (!g54) & (g55)) + ((!sk[16]) & (g182) & (g44) & (g54) & (!g55)) + ((!sk[16]) & (g182) & (g44) & (g54) & (g55)) + ((sk[16]) & (!g182) & (!g44) & (!g54) & (!g55)) + ((sk[16]) & (!g182) & (!g44) & (!g54) & (g55)) + ((sk[16]) & (!g182) & (g44) & (!g54) & (!g55)) + ((sk[16]) & (g182) & (!g44) & (!g54) & (!g55)) + ((sk[16]) & (g182) & (g44) & (!g54) & (!g55)));
	assign g112 = (((!g51) & (!g53) & (!c) & (!g92) & (!sk[25]) & (g111)) + ((!g51) & (!g53) & (!c) & (g92) & (!sk[25]) & (g111)) + ((!g51) & (!g53) & (c) & (!g92) & (!sk[25]) & (g111)) + ((!g51) & (!g53) & (c) & (g92) & (!sk[25]) & (g111)) + ((!g51) & (!g53) & (c) & (g92) & (sk[25]) & (!g111)) + ((!g51) & (!g53) & (c) & (g92) & (sk[25]) & (g111)) + ((!g51) & (g53) & (!c) & (!g92) & (!sk[25]) & (g111)) + ((!g51) & (g53) & (!c) & (g92) & (!sk[25]) & (g111)) + ((!g51) & (g53) & (c) & (!g92) & (!sk[25]) & (g111)) + ((!g51) & (g53) & (c) & (g92) & (sk[25]) & (!g111)) + ((!g51) & (g53) & (c) & (g92) & (sk[25]) & (g111)) + ((g51) & (!g53) & (!c) & (!g92) & (sk[25]) & (!g111)) + ((g51) & (!g53) & (!c) & (!g92) & (sk[25]) & (g111)) + ((g51) & (!g53) & (!c) & (g92) & (!sk[25]) & (g111)) + ((g51) & (!g53) & (!c) & (g92) & (sk[25]) & (!g111)) + ((g51) & (!g53) & (!c) & (g92) & (sk[25]) & (g111)) + ((g51) & (!g53) & (c) & (!g92) & (!sk[25]) & (g111)) + ((g51) & (!g53) & (c) & (!g92) & (sk[25]) & (!g111)) + ((g51) & (!g53) & (c) & (!g92) & (sk[25]) & (g111)) + ((g51) & (!g53) & (c) & (g92) & (!sk[25]) & (g111)) + ((g51) & (!g53) & (c) & (g92) & (sk[25]) & (!g111)) + ((g51) & (!g53) & (c) & (g92) & (sk[25]) & (g111)) + ((g51) & (g53) & (!c) & (!g92) & (sk[25]) & (!g111)) + ((g51) & (g53) & (!c) & (!g92) & (sk[25]) & (g111)) + ((g51) & (g53) & (!c) & (g92) & (!sk[25]) & (g111)) + ((g51) & (g53) & (!c) & (g92) & (sk[25]) & (!g111)) + ((g51) & (g53) & (!c) & (g92) & (sk[25]) & (g111)) + ((g51) & (g53) & (c) & (!g92) & (!sk[25]) & (g111)) + ((g51) & (g53) & (c) & (!g92) & (sk[25]) & (!g111)) + ((g51) & (g53) & (c) & (!g92) & (sk[25]) & (g111)) + ((g51) & (g53) & (c) & (g92) & (sk[25]) & (!g111)) + ((g51) & (g53) & (c) & (g92) & (sk[25]) & (g111)));
	assign g113 = (((!n) & (!g93) & (!g108) & (!g109) & (!g110) & (!g112)) + ((!n) & (!g93) & (!g108) & (!g109) & (!g110) & (g112)) + ((!n) & (g93) & (!g108) & (!g109) & (!g110) & (!g112)) + ((!n) & (g93) & (!g108) & (!g109) & (!g110) & (g112)) + ((n) & (!g93) & (!g108) & (!g109) & (!g110) & (g112)) + ((n) & (g93) & (!g108) & (!g109) & (!g110) & (!g112)) + ((n) & (g93) & (!g108) & (!g109) & (!g110) & (g112)));
	assign g114 = (((!g68) & (g90) & (sk[20]) & (!g103) & (!g106)) + ((!g68) & (g90) & (sk[20]) & (!g103) & (g106)) + ((!g68) & (g90) & (sk[20]) & (g103) & (!g106)) + ((!g68) & (g90) & (sk[20]) & (g103) & (g106)) + ((g68) & (!g90) & (!sk[20]) & (g103) & (g106)) + ((g68) & (!g90) & (sk[20]) & (!g103) & (!g106)) + ((g68) & (!g90) & (sk[20]) & (!g103) & (g106)) + ((g68) & (!g90) & (sk[20]) & (g103) & (!g106)) + ((g68) & (!g90) & (sk[20]) & (g103) & (g106)) + ((g68) & (g90) & (!sk[20]) & (g103) & (!g106)) + ((g68) & (g90) & (sk[20]) & (!g103) & (!g106)) + ((g68) & (g90) & (sk[20]) & (!g103) & (g106)) + ((g68) & (g90) & (sk[20]) & (g103) & (!g106)) + ((g68) & (g90) & (sk[20]) & (g103) & (g106)));
	assign g116 = (((!k) & (!l) & (!i) & (!c) & (!g) & (!g93)) + ((!k) & (!l) & (!i) & (!c) & (g) & (!g93)) + ((!k) & (!l) & (!i) & (c) & (!g) & (!g93)) + ((!k) & (!l) & (!i) & (c) & (g) & (!g93)) + ((!k) & (!l) & (i) & (!c) & (!g) & (g93)) + ((!k) & (!l) & (i) & (!c) & (g) & (g93)) + ((!k) & (!l) & (i) & (c) & (!g) & (g93)) + ((!k) & (!l) & (i) & (c) & (g) & (g93)) + ((!k) & (l) & (!i) & (!c) & (!g) & (!g93)) + ((!k) & (l) & (!i) & (!c) & (g) & (!g93)) + ((!k) & (l) & (!i) & (c) & (!g) & (!g93)) + ((!k) & (l) & (!i) & (c) & (!g) & (g93)) + ((!k) & (l) & (!i) & (c) & (g) & (!g93)) + ((!k) & (l) & (i) & (!c) & (g) & (!g93)) + ((!k) & (l) & (i) & (!c) & (g) & (g93)) + ((!k) & (l) & (i) & (c) & (!g) & (!g93)) + ((!k) & (l) & (i) & (c) & (!g) & (g93)) + ((k) & (!l) & (!i) & (!c) & (!g) & (g93)) + ((k) & (!l) & (!i) & (!c) & (g) & (g93)) + ((k) & (!l) & (!i) & (c) & (!g) & (g93)) + ((k) & (!l) & (!i) & (c) & (g) & (g93)) + ((k) & (!l) & (i) & (!c) & (!g) & (!g93)) + ((k) & (!l) & (i) & (!c) & (!g) & (g93)) + ((k) & (!l) & (i) & (c) & (!g) & (!g93)) + ((k) & (!l) & (i) & (c) & (!g) & (g93)) + ((k) & (l) & (!i) & (!c) & (!g) & (!g93)) + ((k) & (l) & (!i) & (!c) & (!g) & (g93)) + ((k) & (l) & (!i) & (!c) & (g) & (!g93)) + ((k) & (l) & (!i) & (!c) & (g) & (g93)) + ((k) & (l) & (!i) & (c) & (!g) & (!g93)) + ((k) & (l) & (!i) & (c) & (!g) & (g93)) + ((k) & (l) & (!i) & (c) & (g) & (!g93)) + ((k) & (l) & (!i) & (c) & (g) & (g93)) + ((k) & (l) & (i) & (!c) & (!g) & (!g93)) + ((k) & (l) & (i) & (!c) & (g) & (!g93)) + ((k) & (l) & (i) & (c) & (!g) & (!g93)) + ((k) & (l) & (i) & (c) & (!g) & (g93)) + ((k) & (l) & (i) & (c) & (g) & (!g93)));
	assign g117 = (((!k) & (l) & (!i) & (!c) & (g) & (!g93)) + ((!k) & (l) & (!i) & (!c) & (g) & (g93)) + ((!k) & (l) & (!i) & (c) & (g) & (!g93)) + ((!k) & (l) & (!i) & (c) & (g) & (g93)) + ((k) & (!l) & (!i) & (!c) & (!g) & (!g93)) + ((k) & (!l) & (!i) & (!c) & (!g) & (g93)) + ((k) & (!l) & (i) & (c) & (!g) & (!g93)) + ((k) & (!l) & (i) & (c) & (g) & (!g93)) + ((k) & (l) & (!i) & (!c) & (g) & (!g93)) + ((k) & (l) & (!i) & (!c) & (g) & (g93)) + ((k) & (l) & (!i) & (c) & (g) & (!g93)) + ((k) & (l) & (!i) & (c) & (g) & (g93)) + ((k) & (l) & (i) & (c) & (!g) & (!g93)) + ((k) & (l) & (i) & (c) & (g) & (!g93)));
	assign g118 = (((!g34) & (g32) & (!sk[21]) & (!c) & (!g93)) + ((!g34) & (g32) & (!sk[21]) & (!c) & (g93)) + ((!g34) & (g32) & (!sk[21]) & (c) & (!g93)) + ((!g34) & (g32) & (!sk[21]) & (c) & (g93)) + ((!g34) & (g32) & (sk[21]) & (!c) & (!g93)) + ((!g34) & (g32) & (sk[21]) & (c) & (!g93)) + ((g34) & (!g32) & (!sk[21]) & (!c) & (!g93)) + ((g34) & (!g32) & (!sk[21]) & (!c) & (g93)) + ((g34) & (!g32) & (!sk[21]) & (c) & (!g93)) + ((g34) & (!g32) & (!sk[21]) & (c) & (g93)) + ((g34) & (!g32) & (sk[21]) & (c) & (!g93)) + ((g34) & (!g32) & (sk[21]) & (c) & (g93)) + ((g34) & (g32) & (!sk[21]) & (!c) & (!g93)) + ((g34) & (g32) & (!sk[21]) & (!c) & (g93)) + ((g34) & (g32) & (!sk[21]) & (c) & (!g93)) + ((g34) & (g32) & (!sk[21]) & (c) & (g93)) + ((g34) & (g32) & (sk[21]) & (!c) & (!g93)) + ((g34) & (g32) & (sk[21]) & (c) & (!g93)) + ((g34) & (g32) & (sk[21]) & (c) & (g93)));
	assign g123 = (((!k) & (!l) & (!i) & (!sk[23]) & (j) & (!g122)) + ((!k) & (!l) & (!i) & (!sk[23]) & (j) & (g122)) + ((!k) & (!l) & (i) & (!sk[23]) & (j) & (!g122)) + ((!k) & (!l) & (i) & (!sk[23]) & (j) & (g122)) + ((!k) & (l) & (!i) & (!sk[23]) & (!j) & (!g122)) + ((!k) & (l) & (!i) & (!sk[23]) & (!j) & (g122)) + ((!k) & (l) & (!i) & (!sk[23]) & (j) & (!g122)) + ((!k) & (l) & (!i) & (!sk[23]) & (j) & (g122)) + ((!k) & (l) & (!i) & (sk[23]) & (!j) & (!g122)) + ((!k) & (l) & (!i) & (sk[23]) & (!j) & (g122)) + ((!k) & (l) & (i) & (!sk[23]) & (!j) & (!g122)) + ((!k) & (l) & (i) & (!sk[23]) & (!j) & (g122)) + ((!k) & (l) & (i) & (!sk[23]) & (j) & (!g122)) + ((!k) & (l) & (i) & (!sk[23]) & (j) & (g122)) + ((!k) & (l) & (i) & (sk[23]) & (j) & (!g122)) + ((!k) & (l) & (i) & (sk[23]) & (j) & (g122)) + ((k) & (!l) & (!i) & (!sk[23]) & (!j) & (g122)) + ((k) & (!l) & (!i) & (!sk[23]) & (j) & (!g122)) + ((k) & (!l) & (!i) & (!sk[23]) & (j) & (g122)) + ((k) & (!l) & (!i) & (sk[23]) & (!j) & (!g122)) + ((k) & (!l) & (!i) & (sk[23]) & (!j) & (g122)) + ((k) & (!l) & (!i) & (sk[23]) & (j) & (g122)) + ((k) & (!l) & (i) & (!sk[23]) & (!j) & (g122)) + ((k) & (!l) & (i) & (!sk[23]) & (j) & (!g122)) + ((k) & (!l) & (i) & (!sk[23]) & (j) & (g122)) + ((k) & (!l) & (i) & (sk[23]) & (!j) & (!g122)) + ((k) & (!l) & (i) & (sk[23]) & (!j) & (g122)) + ((k) & (l) & (!i) & (!sk[23]) & (!j) & (!g122)) + ((k) & (l) & (!i) & (!sk[23]) & (!j) & (g122)) + ((k) & (l) & (!i) & (!sk[23]) & (j) & (!g122)) + ((k) & (l) & (!i) & (!sk[23]) & (j) & (g122)) + ((k) & (l) & (i) & (!sk[23]) & (!j) & (!g122)) + ((k) & (l) & (i) & (!sk[23]) & (!j) & (g122)) + ((k) & (l) & (i) & (!sk[23]) & (j) & (!g122)) + ((k) & (l) & (i) & (!sk[23]) & (j) & (g122)));
	assign g125 = (((!sk[22]) & (!n) & (!j) & (h)) + ((!sk[22]) & (!n) & (j) & (h)) + ((!sk[22]) & (n) & (!j) & (h)) + ((!sk[22]) & (n) & (j) & (h)) + ((sk[22]) & (n) & (j) & (!h)));
	assign g126 = (((!sk[22]) & (!k) & (!l) & (n) & (!j)) + ((!sk[22]) & (!k) & (!l) & (n) & (j)) + ((!sk[22]) & (!k) & (l) & (n) & (!j)) + ((!sk[22]) & (!k) & (l) & (n) & (j)) + ((!sk[22]) & (k) & (!l) & (n) & (!j)) + ((!sk[22]) & (k) & (!l) & (n) & (j)) + ((!sk[22]) & (k) & (l) & (n) & (!j)) + ((!sk[22]) & (k) & (l) & (n) & (j)) + ((sk[22]) & (!k) & (!l) & (!n) & (!j)) + ((sk[22]) & (!k) & (!l) & (!n) & (j)) + ((sk[22]) & (!k) & (l) & (!n) & (!j)));
	assign g127 = (((!i) & (!sk[23]) & (!d) & (!g122) & (!g125) & (g126)) + ((!i) & (!sk[23]) & (!d) & (!g122) & (g125) & (g126)) + ((!i) & (!sk[23]) & (!d) & (g122) & (!g125) & (!g126)) + ((!i) & (!sk[23]) & (!d) & (g122) & (!g125) & (g126)) + ((!i) & (!sk[23]) & (!d) & (g122) & (g125) & (!g126)) + ((!i) & (!sk[23]) & (!d) & (g122) & (g125) & (g126)) + ((!i) & (!sk[23]) & (d) & (!g122) & (!g125) & (g126)) + ((!i) & (!sk[23]) & (d) & (!g122) & (g125) & (!g126)) + ((!i) & (!sk[23]) & (d) & (!g122) & (g125) & (g126)) + ((!i) & (!sk[23]) & (d) & (g122) & (!g125) & (!g126)) + ((!i) & (!sk[23]) & (d) & (g122) & (!g125) & (g126)) + ((!i) & (!sk[23]) & (d) & (g122) & (g125) & (!g126)) + ((!i) & (!sk[23]) & (d) & (g122) & (g125) & (g126)) + ((!i) & (sk[23]) & (!d) & (!g122) & (!g125) & (g126)) + ((!i) & (sk[23]) & (!d) & (!g122) & (g125) & (g126)) + ((!i) & (sk[23]) & (!d) & (g122) & (!g125) & (g126)) + ((!i) & (sk[23]) & (!d) & (g122) & (g125) & (!g126)) + ((!i) & (sk[23]) & (!d) & (g122) & (g125) & (g126)) + ((i) & (!sk[23]) & (!d) & (!g122) & (!g125) & (g126)) + ((i) & (!sk[23]) & (!d) & (!g122) & (g125) & (g126)) + ((i) & (!sk[23]) & (!d) & (g122) & (!g125) & (!g126)) + ((i) & (!sk[23]) & (!d) & (g122) & (!g125) & (g126)) + ((i) & (!sk[23]) & (!d) & (g122) & (g125) & (!g126)) + ((i) & (!sk[23]) & (!d) & (g122) & (g125) & (g126)) + ((i) & (!sk[23]) & (d) & (!g122) & (!g125) & (g126)) + ((i) & (!sk[23]) & (d) & (!g122) & (g125) & (!g126)) + ((i) & (!sk[23]) & (d) & (!g122) & (g125) & (g126)) + ((i) & (!sk[23]) & (d) & (g122) & (!g125) & (!g126)) + ((i) & (!sk[23]) & (d) & (g122) & (!g125) & (g126)) + ((i) & (!sk[23]) & (d) & (g122) & (g125) & (!g126)) + ((i) & (!sk[23]) & (d) & (g122) & (g125) & (g126)));
	assign g128 = (((!g1) & (!d) & (sk[9]) & (h)) + ((!g1) & (d) & (!sk[9]) & (!h)) + ((!g1) & (d) & (sk[9]) & (h)) + ((g1) & (!d) & (!sk[9]) & (h)) + ((g1) & (!d) & (sk[9]) & (!h)) + ((g1) & (!d) & (sk[9]) & (h)) + ((g1) & (d) & (!sk[9]) & (!h)) + ((g1) & (d) & (sk[9]) & (!h)) + ((g1) & (d) & (sk[9]) & (h)));
	assign g129 = (((!k) & (!sk[23]) & (!l) & (n) & (!c) & (!g121)) + ((!k) & (!sk[23]) & (!l) & (n) & (!c) & (g121)) + ((!k) & (!sk[23]) & (!l) & (n) & (c) & (!g121)) + ((!k) & (!sk[23]) & (!l) & (n) & (c) & (g121)) + ((!k) & (!sk[23]) & (l) & (n) & (!c) & (!g121)) + ((!k) & (!sk[23]) & (l) & (n) & (!c) & (g121)) + ((!k) & (!sk[23]) & (l) & (n) & (c) & (!g121)) + ((!k) & (!sk[23]) & (l) & (n) & (c) & (g121)) + ((k) & (!sk[23]) & (!l) & (n) & (!c) & (!g121)) + ((k) & (!sk[23]) & (!l) & (n) & (!c) & (g121)) + ((k) & (!sk[23]) & (!l) & (n) & (c) & (!g121)) + ((k) & (!sk[23]) & (!l) & (n) & (c) & (g121)) + ((k) & (!sk[23]) & (l) & (n) & (!c) & (!g121)) + ((k) & (!sk[23]) & (l) & (n) & (!c) & (g121)) + ((k) & (!sk[23]) & (l) & (n) & (c) & (!g121)) + ((k) & (!sk[23]) & (l) & (n) & (c) & (g121)) + ((k) & (sk[23]) & (!l) & (!n) & (!c) & (g121)) + ((k) & (sk[23]) & (!l) & (!n) & (c) & (g121)) + ((k) & (sk[23]) & (!l) & (n) & (!c) & (g121)) + ((k) & (sk[23]) & (!l) & (n) & (c) & (g121)) + ((k) & (sk[23]) & (l) & (n) & (c) & (!g121)) + ((k) & (sk[23]) & (l) & (n) & (c) & (g121)));
	assign g130 = (((!g2) & (!g4) & (!sk[9]) & (!d) & (!h)) + ((!g2) & (!g4) & (!sk[9]) & (!d) & (h)) + ((!g2) & (!g4) & (!sk[9]) & (d) & (!h)) + ((!g2) & (!g4) & (!sk[9]) & (d) & (h)) + ((!g2) & (g4) & (!sk[9]) & (!d) & (!h)) + ((g2) & (!g4) & (!sk[9]) & (!d) & (h)) + ((g2) & (!g4) & (!sk[9]) & (d) & (h)));
	assign g131 = (((!sk[23]) & (i) & (!j) & (!g129) & (!g130)) + ((!sk[23]) & (i) & (!j) & (!g129) & (g130)) + ((!sk[23]) & (i) & (!j) & (g129) & (!g130)) + ((!sk[23]) & (i) & (!j) & (g129) & (g130)) + ((!sk[23]) & (i) & (j) & (!g129) & (!g130)) + ((!sk[23]) & (i) & (j) & (!g129) & (g130)) + ((!sk[23]) & (i) & (j) & (g129) & (!g130)) + ((!sk[23]) & (i) & (j) & (g129) & (g130)) + ((sk[23]) & (!i) & (!j) & (!g129) & (g130)) + ((sk[23]) & (!i) & (j) & (!g129) & (g130)) + ((sk[23]) & (!i) & (j) & (g129) & (g130)) + ((sk[23]) & (i) & (!j) & (!g129) & (g130)) + ((sk[23]) & (i) & (!j) & (g129) & (g130)) + ((sk[23]) & (i) & (j) & (!g129) & (g130)) + ((sk[23]) & (i) & (j) & (g129) & (g130)));
	assign g133 = (((!g9) & (!g12) & (!sk[25]) & (!d)) + ((!g9) & (!g12) & (!sk[25]) & (d)) + ((g9) & (!g12) & (!sk[25]) & (!d)));
	assign g134 = (((!g7) & (!g12) & (!d) & (sk[9]) & (h)) + ((!g7) & (!g12) & (d) & (sk[9]) & (!h)) + ((!g7) & (!g12) & (d) & (sk[9]) & (h)) + ((!g7) & (g12) & (!d) & (sk[9]) & (!h)) + ((!g7) & (g12) & (!d) & (sk[9]) & (h)) + ((!g7) & (g12) & (d) & (!sk[9]) & (!h)) + ((!g7) & (g12) & (d) & (!sk[9]) & (h)) + ((!g7) & (g12) & (d) & (sk[9]) & (!h)) + ((!g7) & (g12) & (d) & (sk[9]) & (h)) + ((g7) & (!g12) & (!d) & (sk[9]) & (h)) + ((g7) & (!g12) & (d) & (!sk[9]) & (h)) + ((g7) & (!g12) & (d) & (sk[9]) & (!h)) + ((g7) & (!g12) & (d) & (sk[9]) & (h)) + ((g7) & (g12) & (!d) & (sk[9]) & (!h)) + ((g7) & (g12) & (!d) & (sk[9]) & (h)) + ((g7) & (g12) & (d) & (!sk[9]) & (!h)) + ((g7) & (g12) & (d) & (!sk[9]) & (h)) + ((g7) & (g12) & (d) & (sk[9]) & (!h)) + ((g7) & (g12) & (d) & (sk[9]) & (h)));
	assign g136 = (((!a) & (!sk[18]) & (!b) & (!c) & (d)) + ((!a) & (!sk[18]) & (!b) & (c) & (!d)) + ((!a) & (!sk[18]) & (!b) & (c) & (d)) + ((!a) & (!sk[18]) & (b) & (!c) & (d)) + ((!a) & (!sk[18]) & (b) & (c) & (!d)) + ((!a) & (!sk[18]) & (b) & (c) & (d)) + ((!a) & (sk[18]) & (!b) & (!c) & (!d)) + ((!a) & (sk[18]) & (!b) & (c) & (d)) + ((!a) & (sk[18]) & (b) & (!c) & (d)) + ((!a) & (sk[18]) & (b) & (c) & (d)) + ((a) & (!sk[18]) & (!b) & (!c) & (d)) + ((a) & (!sk[18]) & (!b) & (c) & (!d)) + ((a) & (!sk[18]) & (!b) & (c) & (d)) + ((a) & (!sk[18]) & (b) & (!c) & (d)) + ((a) & (!sk[18]) & (b) & (c) & (!d)) + ((a) & (!sk[18]) & (b) & (c) & (d)) + ((a) & (sk[18]) & (!b) & (!c) & (d)) + ((a) & (sk[18]) & (!b) & (c) & (d)) + ((a) & (sk[18]) & (b) & (!c) & (d)) + ((a) & (sk[18]) & (b) & (c) & (d)));
	assign g137 = (((!l) & (!g60) & (!g120) & (sk[17]) & (g135) & (g136)) + ((!l) & (!g60) & (g120) & (sk[17]) & (g135) & (g136)) + ((!l) & (g60) & (!g120) & (!sk[17]) & (!g135) & (!g136)) + ((!l) & (g60) & (!g120) & (!sk[17]) & (!g135) & (g136)) + ((!l) & (g60) & (!g120) & (sk[17]) & (!g135) & (!g136)) + ((!l) & (g60) & (!g120) & (sk[17]) & (!g135) & (g136)) + ((!l) & (g60) & (!g120) & (sk[17]) & (g135) & (!g136)) + ((!l) & (g60) & (!g120) & (sk[17]) & (g135) & (g136)) + ((!l) & (g60) & (g120) & (!sk[17]) & (g135) & (!g136)) + ((!l) & (g60) & (g120) & (!sk[17]) & (g135) & (g136)) + ((!l) & (g60) & (g120) & (sk[17]) & (!g135) & (!g136)) + ((!l) & (g60) & (g120) & (sk[17]) & (!g135) & (g136)) + ((!l) & (g60) & (g120) & (sk[17]) & (g135) & (!g136)) + ((!l) & (g60) & (g120) & (sk[17]) & (g135) & (g136)) + ((l) & (!g60) & (!g120) & (sk[17]) & (g135) & (g136)) + ((l) & (!g60) & (g120) & (sk[17]) & (g135) & (g136)) + ((l) & (g60) & (!g120) & (!sk[17]) & (!g135) & (g136)) + ((l) & (g60) & (!g120) & (!sk[17]) & (g135) & (g136)) + ((l) & (g60) & (!g120) & (sk[17]) & (!g135) & (!g136)) + ((l) & (g60) & (!g120) & (sk[17]) & (!g135) & (g136)) + ((l) & (g60) & (!g120) & (sk[17]) & (g135) & (!g136)) + ((l) & (g60) & (!g120) & (sk[17]) & (g135) & (g136)) + ((l) & (g60) & (g120) & (!sk[17]) & (!g135) & (g136)) + ((l) & (g60) & (g120) & (!sk[17]) & (g135) & (g136)) + ((l) & (g60) & (g120) & (sk[17]) & (!g135) & (!g136)) + ((l) & (g60) & (g120) & (sk[17]) & (!g135) & (g136)) + ((l) & (g60) & (g120) & (sk[17]) & (g135) & (!g136)) + ((l) & (g60) & (g120) & (sk[17]) & (g135) & (g136)));
	assign g140 = (((!n) & (sk[26]) & (!g18) & (!g135) & (g138) & (!g139)) + ((!n) & (sk[26]) & (!g18) & (!g135) & (g138) & (g139)) + ((!n) & (sk[26]) & (!g18) & (g135) & (!g138) & (!g139)) + ((!n) & (sk[26]) & (!g18) & (g135) & (!g138) & (g139)) + ((!n) & (sk[26]) & (!g18) & (g135) & (g138) & (!g139)) + ((!n) & (sk[26]) & (!g18) & (g135) & (g138) & (g139)) + ((!n) & (sk[26]) & (g18) & (!g135) & (!g138) & (g139)) + ((!n) & (sk[26]) & (g18) & (!g135) & (g138) & (!g139)) + ((!n) & (sk[26]) & (g18) & (!g135) & (g138) & (g139)) + ((!n) & (sk[26]) & (g18) & (g135) & (!g138) & (!g139)) + ((!n) & (sk[26]) & (g18) & (g135) & (!g138) & (g139)) + ((!n) & (sk[26]) & (g18) & (g135) & (g138) & (!g139)) + ((!n) & (sk[26]) & (g18) & (g135) & (g138) & (g139)) + ((n) & (!sk[26]) & (g18) & (!g135) & (!g138) & (g139)) + ((n) & (!sk[26]) & (g18) & (!g135) & (g138) & (!g139)) + ((n) & (!sk[26]) & (g18) & (g135) & (!g138) & (!g139)) + ((n) & (!sk[26]) & (g18) & (g135) & (g138) & (g139)) + ((n) & (sk[26]) & (!g18) & (!g135) & (g138) & (!g139)) + ((n) & (sk[26]) & (!g18) & (!g135) & (g138) & (g139)) + ((n) & (sk[26]) & (!g18) & (g135) & (!g138) & (!g139)) + ((n) & (sk[26]) & (!g18) & (g135) & (!g138) & (g139)) + ((n) & (sk[26]) & (!g18) & (g135) & (g138) & (!g139)) + ((n) & (sk[26]) & (!g18) & (g135) & (g138) & (g139)) + ((n) & (sk[26]) & (g18) & (!g135) & (!g138) & (g139)) + ((n) & (sk[26]) & (g18) & (!g135) & (g138) & (!g139)) + ((n) & (sk[26]) & (g18) & (!g135) & (g138) & (g139)) + ((n) & (sk[26]) & (g18) & (g135) & (!g138) & (!g139)) + ((n) & (sk[26]) & (g18) & (g135) & (!g138) & (g139)) + ((n) & (sk[26]) & (g18) & (g135) & (g138) & (!g139)) + ((n) & (sk[26]) & (g18) & (g135) & (g138) & (g139)));
	assign g142 = (((g7) & (!g93) & (g103) & (!g104) & (!g141) & (!g138)) + ((g7) & (!g93) & (g103) & (!g104) & (g141) & (g138)) + ((g7) & (g93) & (!g103) & (!g104) & (!g141) & (!g138)) + ((g7) & (g93) & (!g103) & (!g104) & (g141) & (g138)) + ((g7) & (g93) & (g103) & (!g104) & (!g141) & (!g138)) + ((g7) & (g93) & (g103) & (!g104) & (g141) & (g138)) + ((g7) & (g93) & (g103) & (g104) & (!g141) & (!g138)) + ((g7) & (g93) & (g103) & (g104) & (g141) & (g138)));
	assign g143 = (((g7) & (!g93) & (!g103) & (!g104) & (!g141) & (g138)) + ((g7) & (!g93) & (!g103) & (!g104) & (g141) & (!g138)) + ((g7) & (!g93) & (!g103) & (g104) & (!g141) & (g138)) + ((g7) & (!g93) & (!g103) & (g104) & (g141) & (!g138)) + ((g7) & (!g93) & (g103) & (g104) & (!g141) & (g138)) + ((g7) & (!g93) & (g103) & (g104) & (g141) & (!g138)) + ((g7) & (g93) & (!g103) & (g104) & (!g141) & (g138)) + ((g7) & (g93) & (!g103) & (g104) & (g141) & (!g138)));
	assign g144 = (((!g53) & (!g57) & (!c) & (!g92) & (!g93) & (!g141)) + ((!g53) & (!g57) & (!c) & (!g92) & (!g93) & (g141)) + ((!g53) & (!g57) & (!c) & (!g92) & (g93) & (!g141)) + ((!g53) & (!g57) & (!c) & (!g92) & (g93) & (g141)) + ((!g53) & (!g57) & (!c) & (g92) & (!g93) & (!g141)) + ((!g53) & (!g57) & (!c) & (g92) & (!g93) & (g141)) + ((!g53) & (!g57) & (!c) & (g92) & (g93) & (!g141)) + ((!g53) & (!g57) & (!c) & (g92) & (g93) & (g141)) + ((!g53) & (!g57) & (c) & (!g92) & (!g93) & (!g141)) + ((!g53) & (!g57) & (c) & (!g92) & (!g93) & (g141)) + ((!g53) & (!g57) & (c) & (!g92) & (g93) & (!g141)) + ((!g53) & (!g57) & (c) & (!g92) & (g93) & (g141)) + ((!g53) & (!g57) & (c) & (g92) & (!g93) & (!g141)) + ((!g53) & (!g57) & (c) & (g92) & (!g93) & (g141)) + ((!g53) & (!g57) & (c) & (g92) & (g93) & (!g141)) + ((!g53) & (!g57) & (c) & (g92) & (g93) & (g141)) + ((g53) & (!g57) & (!c) & (!g92) & (!g93) & (!g141)) + ((g53) & (!g57) & (!c) & (!g92) & (g93) & (!g141)) + ((g53) & (!g57) & (!c) & (g92) & (!g93) & (g141)) + ((g53) & (!g57) & (!c) & (g92) & (g93) & (!g141)) + ((g53) & (!g57) & (c) & (!g92) & (!g93) & (g141)) + ((g53) & (!g57) & (c) & (!g92) & (g93) & (!g141)) + ((g53) & (!g57) & (c) & (g92) & (!g93) & (g141)) + ((g53) & (!g57) & (c) & (g92) & (g93) & (g141)));
	assign g145 = (((n) & (!sk[26]) & (d)) + ((n) & (sk[26]) & (!d)) + ((n) & (sk[26]) & (d)));
	assign g146 = (((n) & (!g62) & (!g54) & (g55) & (!g93) & (!g141)) + ((n) & (!g62) & (!g54) & (g55) & (g93) & (!g141)) + ((n) & (!g62) & (g54) & (!g55) & (!g93) & (!g141)) + ((n) & (!g62) & (g54) & (!g55) & (g93) & (!g141)) + ((n) & (!g62) & (g54) & (g55) & (!g93) & (!g141)) + ((n) & (!g62) & (g54) & (g55) & (g93) & (!g141)) + ((n) & (g62) & (!g54) & (g55) & (!g93) & (!g141)) + ((n) & (g62) & (g54) & (!g55) & (!g93) & (!g141)) + ((n) & (g62) & (g54) & (!g55) & (g93) & (!g141)) + ((n) & (g62) & (g54) & (g55) & (!g93) & (!g141)) + ((n) & (g62) & (g54) & (g55) & (g93) & (!g141)));
	assign g148 = (((!l) & (!g65) & (!d) & (!sk[27]) & (h) & (!g147)) + ((!l) & (!g65) & (!d) & (!sk[27]) & (h) & (g147)) + ((!l) & (!g65) & (d) & (!sk[27]) & (h) & (!g147)) + ((!l) & (!g65) & (d) & (!sk[27]) & (h) & (g147)) + ((!l) & (g65) & (!d) & (!sk[27]) & (!h) & (!g147)) + ((!l) & (g65) & (!d) & (!sk[27]) & (!h) & (g147)) + ((!l) & (g65) & (!d) & (!sk[27]) & (h) & (!g147)) + ((!l) & (g65) & (!d) & (!sk[27]) & (h) & (g147)) + ((!l) & (g65) & (!d) & (sk[27]) & (h) & (!g147)) + ((!l) & (g65) & (!d) & (sk[27]) & (h) & (g147)) + ((!l) & (g65) & (d) & (!sk[27]) & (!h) & (!g147)) + ((!l) & (g65) & (d) & (!sk[27]) & (!h) & (g147)) + ((!l) & (g65) & (d) & (!sk[27]) & (h) & (!g147)) + ((!l) & (g65) & (d) & (!sk[27]) & (h) & (g147)) + ((!l) & (g65) & (d) & (sk[27]) & (!h) & (!g147)) + ((!l) & (g65) & (d) & (sk[27]) & (h) & (!g147)) + ((!l) & (g65) & (d) & (sk[27]) & (h) & (g147)) + ((l) & (!g65) & (!d) & (!sk[27]) & (h) & (!g147)) + ((l) & (!g65) & (!d) & (!sk[27]) & (h) & (g147)) + ((l) & (!g65) & (d) & (!sk[27]) & (h) & (!g147)) + ((l) & (!g65) & (d) & (!sk[27]) & (h) & (g147)) + ((l) & (g65) & (!d) & (!sk[27]) & (!h) & (!g147)) + ((l) & (g65) & (!d) & (!sk[27]) & (!h) & (g147)) + ((l) & (g65) & (!d) & (!sk[27]) & (h) & (!g147)) + ((l) & (g65) & (!d) & (!sk[27]) & (h) & (g147)) + ((l) & (g65) & (!d) & (sk[27]) & (!h) & (g147)) + ((l) & (g65) & (!d) & (sk[27]) & (h) & (!g147)) + ((l) & (g65) & (d) & (!sk[27]) & (!h) & (!g147)) + ((l) & (g65) & (d) & (!sk[27]) & (!h) & (g147)) + ((l) & (g65) & (d) & (!sk[27]) & (h) & (!g147)) + ((l) & (g65) & (d) & (!sk[27]) & (h) & (g147)) + ((l) & (g65) & (d) & (sk[27]) & (!h) & (!g147)) + ((l) & (g65) & (d) & (sk[27]) & (h) & (g147)));
	assign g149 = (((!n) & (sk[26]) & (g51) & (!d)) + ((!n) & (sk[26]) & (g51) & (d)) + ((n) & (!sk[26]) & (g51) & (!d)) + ((n) & (sk[26]) & (g51) & (!d)) + ((n) & (sk[26]) & (g51) & (d)));
	assign g150 = (((!c) & (!g92) & (!g93) & (!g141) & (!g148) & (!g149)) + ((!c) & (!g92) & (!g93) & (g141) & (!g148) & (!g149)) + ((!c) & (!g92) & (!g93) & (g141) & (!g148) & (g149)) + ((!c) & (!g92) & (g93) & (!g141) & (!g148) & (!g149)) + ((!c) & (!g92) & (g93) & (g141) & (!g148) & (!g149)) + ((!c) & (!g92) & (g93) & (g141) & (!g148) & (g149)) + ((!c) & (g92) & (!g93) & (!g141) & (!g148) & (!g149)) + ((!c) & (g92) & (!g93) & (!g141) & (!g148) & (g149)) + ((!c) & (g92) & (!g93) & (g141) & (!g148) & (!g149)) + ((!c) & (g92) & (g93) & (!g141) & (!g148) & (!g149)) + ((!c) & (g92) & (g93) & (g141) & (!g148) & (!g149)) + ((!c) & (g92) & (g93) & (g141) & (!g148) & (g149)) + ((c) & (!g92) & (!g93) & (!g141) & (!g148) & (!g149)) + ((c) & (!g92) & (!g93) & (!g141) & (!g148) & (g149)) + ((c) & (!g92) & (!g93) & (g141) & (!g148) & (!g149)) + ((c) & (!g92) & (g93) & (!g141) & (!g148) & (!g149)) + ((c) & (!g92) & (g93) & (g141) & (!g148) & (!g149)) + ((c) & (!g92) & (g93) & (g141) & (!g148) & (g149)) + ((c) & (g92) & (!g93) & (!g141) & (!g148) & (!g149)) + ((c) & (g92) & (!g93) & (!g141) & (!g148) & (g149)) + ((c) & (g92) & (!g93) & (g141) & (!g148) & (!g149)) + ((c) & (g92) & (g93) & (!g141) & (!g148) & (!g149)) + ((c) & (g92) & (g93) & (!g141) & (!g148) & (g149)) + ((c) & (g92) & (g93) & (g141) & (!g148) & (!g149)));
	assign g151 = (((!g109) & (!g141) & (!g144) & (!g145) & (!g146) & (g150)) + ((!g109) & (!g141) & (g144) & (!g145) & (!g146) & (g150)) + ((!g109) & (!g141) & (g144) & (g145) & (!g146) & (g150)) + ((!g109) & (g141) & (!g144) & (!g145) & (!g146) & (g150)) + ((!g109) & (g141) & (g144) & (!g145) & (!g146) & (g150)) + ((!g109) & (g141) & (g144) & (g145) & (!g146) & (g150)) + ((g109) & (!g141) & (!g144) & (!g145) & (!g146) & (g150)) + ((g109) & (!g141) & (g144) & (!g145) & (!g146) & (g150)) + ((g109) & (!g141) & (g144) & (g145) & (!g146) & (g150)));
	assign g153 = (((!sk[27]) & (!l) & (!i) & (j) & (!d)) + ((!sk[27]) & (!l) & (!i) & (j) & (d)) + ((!sk[27]) & (!l) & (i) & (!j) & (d)) + ((!sk[27]) & (!l) & (i) & (j) & (!d)) + ((!sk[27]) & (!l) & (i) & (j) & (d)) + ((!sk[27]) & (l) & (!i) & (j) & (!d)) + ((!sk[27]) & (l) & (!i) & (j) & (d)) + ((!sk[27]) & (l) & (i) & (!j) & (d)) + ((!sk[27]) & (l) & (i) & (j) & (!d)) + ((!sk[27]) & (l) & (i) & (j) & (d)) + ((sk[27]) & (!l) & (!i) & (!j) & (d)));
	assign g154 = (((!sk[28]) & (!i) & (!j) & (!g1) & (d)) + ((!sk[28]) & (!i) & (!j) & (g1) & (d)) + ((!sk[28]) & (!i) & (j) & (!g1) & (d)) + ((!sk[28]) & (!i) & (j) & (g1) & (d)) + ((!sk[28]) & (i) & (!j) & (!g1) & (!d)) + ((!sk[28]) & (i) & (!j) & (!g1) & (d)) + ((!sk[28]) & (i) & (!j) & (g1) & (!d)) + ((!sk[28]) & (i) & (!j) & (g1) & (d)) + ((!sk[28]) & (i) & (j) & (!g1) & (!d)) + ((!sk[28]) & (i) & (j) & (!g1) & (d)) + ((!sk[28]) & (i) & (j) & (g1) & (!d)) + ((!sk[28]) & (i) & (j) & (g1) & (d)) + ((sk[28]) & (!i) & (!j) & (g1) & (!d)));
	assign g155 = (((!n) & (!g135) & (!g152) & (sk[26]) & (!g153) & (g154)) + ((!n) & (!g135) & (!g152) & (sk[26]) & (g153) & (g154)) + ((!n) & (!g135) & (g152) & (sk[26]) & (!g153) & (g154)) + ((!n) & (!g135) & (g152) & (sk[26]) & (g153) & (g154)) + ((!n) & (g135) & (!g152) & (sk[26]) & (!g153) & (g154)) + ((!n) & (g135) & (!g152) & (sk[26]) & (g153) & (g154)) + ((!n) & (g135) & (g152) & (sk[26]) & (!g153) & (!g154)) + ((!n) & (g135) & (g152) & (sk[26]) & (!g153) & (g154)) + ((!n) & (g135) & (g152) & (sk[26]) & (g153) & (!g154)) + ((!n) & (g135) & (g152) & (sk[26]) & (g153) & (g154)) + ((n) & (!g135) & (!g152) & (!sk[26]) & (!g153) & (g154)) + ((n) & (!g135) & (!g152) & (!sk[26]) & (g153) & (g154)) + ((n) & (!g135) & (!g152) & (sk[26]) & (!g153) & (!g154)) + ((n) & (!g135) & (!g152) & (sk[26]) & (!g153) & (g154)) + ((n) & (!g135) & (!g152) & (sk[26]) & (g153) & (!g154)) + ((n) & (!g135) & (!g152) & (sk[26]) & (g153) & (g154)) + ((n) & (!g135) & (g152) & (!sk[26]) & (g153) & (!g154)) + ((n) & (!g135) & (g152) & (!sk[26]) & (g153) & (g154)) + ((n) & (!g135) & (g152) & (sk[26]) & (!g153) & (!g154)) + ((n) & (!g135) & (g152) & (sk[26]) & (!g153) & (g154)) + ((n) & (!g135) & (g152) & (sk[26]) & (g153) & (!g154)) + ((n) & (!g135) & (g152) & (sk[26]) & (g153) & (g154)) + ((n) & (g135) & (!g152) & (!sk[26]) & (g153) & (!g154)) + ((n) & (g135) & (!g152) & (!sk[26]) & (g153) & (g154)) + ((n) & (g135) & (!g152) & (sk[26]) & (!g153) & (!g154)) + ((n) & (g135) & (!g152) & (sk[26]) & (!g153) & (g154)) + ((n) & (g135) & (!g152) & (sk[26]) & (g153) & (!g154)) + ((n) & (g135) & (!g152) & (sk[26]) & (g153) & (g154)) + ((n) & (g135) & (g152) & (!sk[26]) & (!g153) & (g154)) + ((n) & (g135) & (g152) & (!sk[26]) & (g153) & (g154)) + ((n) & (g135) & (g152) & (sk[26]) & (!g153) & (!g154)) + ((n) & (g135) & (g152) & (sk[26]) & (!g153) & (g154)) + ((n) & (g135) & (g152) & (sk[26]) & (g153) & (!g154)) + ((n) & (g135) & (g152) & (sk[26]) & (g153) & (g154)));
	assign g157 = (((!k) & (!l) & (!i) & (!d) & (!h) & (g141)) + ((!k) & (!l) & (!i) & (!d) & (h) & (g141)) + ((!k) & (!l) & (!i) & (d) & (!h) & (g141)) + ((!k) & (!l) & (!i) & (d) & (h) & (g141)) + ((!k) & (!l) & (i) & (!d) & (!h) & (!g141)) + ((!k) & (!l) & (i) & (!d) & (h) & (!g141)) + ((!k) & (!l) & (i) & (d) & (!h) & (!g141)) + ((!k) & (!l) & (i) & (d) & (h) & (!g141)) + ((!k) & (l) & (!i) & (!d) & (!h) & (g141)) + ((!k) & (l) & (!i) & (!d) & (h) & (g141)) + ((!k) & (l) & (!i) & (d) & (h) & (g141)) + ((!k) & (l) & (i) & (!d) & (!h) & (!g141)) + ((!k) & (l) & (i) & (!d) & (!h) & (g141)) + ((!k) & (l) & (i) & (d) & (h) & (!g141)) + ((!k) & (l) & (i) & (d) & (h) & (g141)) + ((k) & (!l) & (!i) & (!d) & (!h) & (!g141)) + ((k) & (!l) & (!i) & (!d) & (h) & (!g141)) + ((k) & (!l) & (!i) & (d) & (!h) & (!g141)) + ((k) & (!l) & (!i) & (d) & (h) & (!g141)) + ((k) & (!l) & (i) & (!d) & (h) & (!g141)) + ((k) & (!l) & (i) & (!d) & (h) & (g141)) + ((k) & (!l) & (i) & (d) & (h) & (!g141)) + ((k) & (!l) & (i) & (d) & (h) & (g141)) + ((k) & (l) & (i) & (!d) & (!h) & (g141)) + ((k) & (l) & (i) & (!d) & (h) & (g141)) + ((k) & (l) & (i) & (d) & (h) & (g141)));
	assign g158 = (((!k) & (l) & (!i) & (!d) & (h) & (!g141)) + ((!k) & (l) & (!i) & (!d) & (h) & (g141)) + ((!k) & (l) & (!i) & (d) & (h) & (!g141)) + ((!k) & (l) & (!i) & (d) & (h) & (g141)) + ((k) & (!l) & (!i) & (!d) & (!h) & (!g141)) + ((k) & (!l) & (!i) & (!d) & (!h) & (g141)) + ((k) & (!l) & (i) & (d) & (!h) & (!g141)) + ((k) & (!l) & (i) & (d) & (h) & (!g141)) + ((k) & (l) & (!i) & (!d) & (h) & (!g141)) + ((k) & (l) & (!i) & (!d) & (h) & (g141)) + ((k) & (l) & (!i) & (d) & (h) & (!g141)) + ((k) & (l) & (!i) & (d) & (h) & (g141)) + ((k) & (l) & (i) & (d) & (!h) & (!g141)) + ((k) & (l) & (i) & (d) & (h) & (!g141)));
	assign g159 = (((!g33) & (!g34) & (!g35) & (!sk[21]) & (!d) & (h)) + ((!g33) & (!g34) & (!g35) & (!sk[21]) & (d) & (h)) + ((!g33) & (!g34) & (!g35) & (sk[21]) & (!d) & (!h)) + ((!g33) & (!g34) & (!g35) & (sk[21]) & (!d) & (h)) + ((!g33) & (!g34) & (!g35) & (sk[21]) & (d) & (!h)) + ((!g33) & (!g34) & (!g35) & (sk[21]) & (d) & (h)) + ((!g33) & (!g34) & (g35) & (!sk[21]) & (!d) & (h)) + ((!g33) & (!g34) & (g35) & (!sk[21]) & (d) & (h)) + ((!g33) & (!g34) & (g35) & (sk[21]) & (!d) & (!h)) + ((!g33) & (!g34) & (g35) & (sk[21]) & (!d) & (h)) + ((!g33) & (g34) & (!g35) & (!sk[21]) & (!d) & (!h)) + ((!g33) & (g34) & (!g35) & (!sk[21]) & (!d) & (h)) + ((!g33) & (g34) & (!g35) & (!sk[21]) & (d) & (!h)) + ((!g33) & (g34) & (!g35) & (!sk[21]) & (d) & (h)) + ((!g33) & (g34) & (!g35) & (sk[21]) & (!d) & (!h)) + ((!g33) & (g34) & (!g35) & (sk[21]) & (!d) & (h)) + ((!g33) & (g34) & (!g35) & (sk[21]) & (d) & (!h)) + ((!g33) & (g34) & (g35) & (!sk[21]) & (!d) & (!h)) + ((!g33) & (g34) & (g35) & (!sk[21]) & (!d) & (h)) + ((!g33) & (g34) & (g35) & (!sk[21]) & (d) & (!h)) + ((!g33) & (g34) & (g35) & (!sk[21]) & (d) & (h)) + ((!g33) & (g34) & (g35) & (sk[21]) & (!d) & (!h)) + ((!g33) & (g34) & (g35) & (sk[21]) & (!d) & (h)) + ((g33) & (!g34) & (!g35) & (!sk[21]) & (!d) & (!h)) + ((g33) & (!g34) & (!g35) & (!sk[21]) & (!d) & (h)) + ((g33) & (!g34) & (!g35) & (!sk[21]) & (d) & (!h)) + ((g33) & (!g34) & (!g35) & (!sk[21]) & (d) & (h)) + ((g33) & (!g34) & (g35) & (!sk[21]) & (!d) & (!h)) + ((g33) & (!g34) & (g35) & (!sk[21]) & (!d) & (h)) + ((g33) & (!g34) & (g35) & (!sk[21]) & (d) & (!h)) + ((g33) & (!g34) & (g35) & (!sk[21]) & (d) & (h)) + ((g33) & (g34) & (!g35) & (!sk[21]) & (!d) & (!h)) + ((g33) & (g34) & (!g35) & (!sk[21]) & (!d) & (h)) + ((g33) & (g34) & (!g35) & (!sk[21]) & (d) & (!h)) + ((g33) & (g34) & (!g35) & (!sk[21]) & (d) & (h)) + ((g33) & (g34) & (g35) & (!sk[21]) & (!d) & (!h)) + ((g33) & (g34) & (g35) & (!sk[21]) & (!d) & (h)) + ((g33) & (g34) & (g35) & (!sk[21]) & (d) & (!h)) + ((g33) & (g34) & (g35) & (!sk[21]) & (d) & (h)));
	assign g160 = (((!g32) & (!h) & (!g141) & (!sk[29]) & (g159)) + ((!g32) & (!h) & (!g141) & (sk[29]) & (g159)) + ((!g32) & (!h) & (g141) & (!sk[29]) & (g159)) + ((!g32) & (!h) & (g141) & (sk[29]) & (g159)) + ((!g32) & (h) & (!g141) & (!sk[29]) & (g159)) + ((!g32) & (h) & (!g141) & (sk[29]) & (!g159)) + ((!g32) & (h) & (!g141) & (sk[29]) & (g159)) + ((!g32) & (h) & (g141) & (!sk[29]) & (g159)) + ((!g32) & (h) & (g141) & (sk[29]) & (!g159)) + ((!g32) & (h) & (g141) & (sk[29]) & (g159)) + ((g32) & (!h) & (!g141) & (!sk[29]) & (g159)) + ((g32) & (!h) & (!g141) & (sk[29]) & (g159)) + ((g32) & (!h) & (g141) & (!sk[29]) & (g159)) + ((g32) & (!h) & (g141) & (sk[29]) & (g159)) + ((g32) & (h) & (!g141) & (sk[29]) & (!g159)) + ((g32) & (h) & (!g141) & (sk[29]) & (g159)) + ((g32) & (h) & (g141) & (!sk[29]) & (g159)) + ((g32) & (h) & (g141) & (sk[29]) & (!g159)) + ((g32) & (h) & (g141) & (sk[29]) & (g159)));
	assign g161 = (((!n) & (!j) & (g157) & (!sk[22]) & (g158) & (g160)) + ((!n) & (!j) & (g157) & (sk[22]) & (!g158) & (g160)) + ((!n) & (!j) & (g157) & (sk[22]) & (g158) & (g160)) + ((!n) & (j) & (!g157) & (!sk[22]) & (!g158) & (!g160)) + ((!n) & (j) & (!g157) & (!sk[22]) & (!g158) & (g160)) + ((!n) & (j) & (!g157) & (!sk[22]) & (g158) & (!g160)) + ((!n) & (j) & (!g157) & (!sk[22]) & (g158) & (g160)) + ((!n) & (j) & (!g157) & (sk[22]) & (!g158) & (g160)) + ((!n) & (j) & (g157) & (!sk[22]) & (!g158) & (!g160)) + ((!n) & (j) & (g157) & (!sk[22]) & (!g158) & (g160)) + ((!n) & (j) & (g157) & (!sk[22]) & (g158) & (!g160)) + ((!n) & (j) & (g157) & (!sk[22]) & (g158) & (g160)) + ((!n) & (j) & (g157) & (sk[22]) & (!g158) & (g160)) + ((n) & (!j) & (!g157) & (sk[22]) & (!g158) & (g160)) + ((n) & (!j) & (!g157) & (sk[22]) & (g158) & (g160)) + ((n) & (!j) & (g157) & (!sk[22]) & (!g158) & (!g160)) + ((n) & (!j) & (g157) & (!sk[22]) & (!g158) & (g160)) + ((n) & (!j) & (g157) & (!sk[22]) & (g158) & (!g160)) + ((n) & (!j) & (g157) & (!sk[22]) & (g158) & (g160)) + ((n) & (!j) & (g157) & (sk[22]) & (!g158) & (g160)) + ((n) & (!j) & (g157) & (sk[22]) & (g158) & (g160)) + ((n) & (j) & (!g157) & (!sk[22]) & (!g158) & (!g160)) + ((n) & (j) & (!g157) & (!sk[22]) & (!g158) & (g160)) + ((n) & (j) & (!g157) & (!sk[22]) & (g158) & (!g160)) + ((n) & (j) & (!g157) & (!sk[22]) & (g158) & (g160)) + ((n) & (j) & (!g157) & (sk[22]) & (!g158) & (g160)) + ((n) & (j) & (!g157) & (sk[22]) & (g158) & (g160)) + ((n) & (j) & (g157) & (!sk[22]) & (!g158) & (!g160)) + ((n) & (j) & (g157) & (!sk[22]) & (!g158) & (g160)) + ((n) & (j) & (g157) & (!sk[22]) & (g158) & (!g160)) + ((n) & (j) & (g157) & (!sk[22]) & (g158) & (g160)) + ((n) & (j) & (g157) & (sk[22]) & (!g158) & (g160)) + ((n) & (j) & (g157) & (sk[22]) & (g158) & (g160)));
	assign g164 = (((!k) & (!l) & (!g8) & (sk[29]) & (!g120) & (g135)) + ((!k) & (!l) & (!g8) & (sk[29]) & (g120) & (!g135)) + ((!k) & (!l) & (!g8) & (sk[29]) & (g120) & (g135)) + ((!k) & (!l) & (g8) & (!sk[29]) & (!g120) & (!g135)) + ((!k) & (!l) & (g8) & (!sk[29]) & (!g120) & (g135)) + ((!k) & (!l) & (g8) & (!sk[29]) & (g120) & (!g135)) + ((!k) & (!l) & (g8) & (!sk[29]) & (g120) & (g135)) + ((!k) & (!l) & (g8) & (sk[29]) & (!g120) & (g135)) + ((!k) & (!l) & (g8) & (sk[29]) & (g120) & (!g135)) + ((!k) & (!l) & (g8) & (sk[29]) & (g120) & (g135)) + ((!k) & (l) & (!g8) & (sk[29]) & (!g120) & (!g135)) + ((!k) & (l) & (!g8) & (sk[29]) & (!g120) & (g135)) + ((!k) & (l) & (!g8) & (sk[29]) & (g120) & (!g135)) + ((!k) & (l) & (!g8) & (sk[29]) & (g120) & (g135)) + ((!k) & (l) & (g8) & (sk[29]) & (!g120) & (!g135)) + ((!k) & (l) & (g8) & (sk[29]) & (!g120) & (g135)) + ((!k) & (l) & (g8) & (sk[29]) & (g120) & (!g135)) + ((!k) & (l) & (g8) & (sk[29]) & (g120) & (g135)) + ((k) & (!l) & (!g8) & (sk[29]) & (!g120) & (g135)) + ((k) & (!l) & (!g8) & (sk[29]) & (g120) & (!g135)) + ((k) & (!l) & (!g8) & (sk[29]) & (g120) & (g135)) + ((k) & (!l) & (g8) & (!sk[29]) & (g120) & (g135)) + ((k) & (!l) & (g8) & (sk[29]) & (!g120) & (g135)) + ((k) & (!l) & (g8) & (sk[29]) & (g120) & (!g135)) + ((k) & (!l) & (g8) & (sk[29]) & (g120) & (g135)) + ((k) & (l) & (!g8) & (sk[29]) & (!g120) & (!g135)) + ((k) & (l) & (!g8) & (sk[29]) & (!g120) & (g135)) + ((k) & (l) & (!g8) & (sk[29]) & (g120) & (!g135)) + ((k) & (l) & (!g8) & (sk[29]) & (g120) & (g135)) + ((k) & (l) & (g8) & (sk[29]) & (!g120) & (!g135)) + ((k) & (l) & (g8) & (sk[29]) & (!g120) & (g135)) + ((k) & (l) & (g8) & (sk[29]) & (g120) & (!g135)) + ((k) & (l) & (g8) & (sk[29]) & (g120) & (g135)));
	assign g165 = (((!sk[28]) & (!i) & (d) & (!g135) & (!g152)) + ((!sk[28]) & (!i) & (d) & (!g135) & (g152)) + ((!sk[28]) & (!i) & (d) & (g135) & (!g152)) + ((!sk[28]) & (!i) & (d) & (g135) & (g152)) + ((!sk[28]) & (i) & (!d) & (g135) & (!g152)) + ((!sk[28]) & (i) & (!d) & (g135) & (g152)) + ((!sk[28]) & (i) & (d) & (!g135) & (!g152)) + ((!sk[28]) & (i) & (d) & (!g135) & (g152)) + ((!sk[28]) & (i) & (d) & (g135) & (!g152)) + ((!sk[28]) & (i) & (d) & (g135) & (g152)) + ((sk[28]) & (!i) & (d) & (!g135) & (!g152)) + ((sk[28]) & (!i) & (d) & (!g135) & (g152)) + ((sk[28]) & (!i) & (d) & (g135) & (g152)));
	assign g166 = (((i) & (!g93) & (!g103) & (!g104) & (!g141) & (!g138)) + ((i) & (!g93) & (!g103) & (!g104) & (!g141) & (g138)) + ((i) & (!g93) & (!g103) & (!g104) & (g141) & (g138)) + ((i) & (!g93) & (!g103) & (g104) & (!g141) & (!g138)) + ((i) & (!g93) & (!g103) & (g104) & (!g141) & (g138)) + ((i) & (!g93) & (!g103) & (g104) & (g141) & (g138)) + ((i) & (!g93) & (g103) & (g104) & (!g141) & (!g138)) + ((i) & (!g93) & (g103) & (g104) & (!g141) & (g138)) + ((i) & (!g93) & (g103) & (g104) & (g141) & (g138)) + ((i) & (g93) & (!g103) & (g104) & (!g141) & (!g138)) + ((i) & (g93) & (!g103) & (g104) & (!g141) & (g138)) + ((i) & (g93) & (!g103) & (g104) & (g141) & (g138)));
	assign g167 = (((!sk[26]) & (!i) & (!g141) & (!g135) & (!g138) & (g152)) + ((!sk[26]) & (!i) & (!g141) & (!g135) & (g138) & (g152)) + ((!sk[26]) & (!i) & (g141) & (!g135) & (!g138) & (g152)) + ((!sk[26]) & (!i) & (g141) & (!g135) & (g138) & (g152)) + ((!sk[26]) & (i) & (!g141) & (!g135) & (g138) & (!g152)) + ((!sk[26]) & (i) & (!g141) & (!g135) & (g138) & (g152)) + ((!sk[26]) & (i) & (!g141) & (g135) & (g138) & (!g152)) + ((!sk[26]) & (i) & (!g141) & (g135) & (g138) & (g152)) + ((sk[26]) & (!i) & (!g141) & (!g135) & (g138) & (!g152)) + ((sk[26]) & (!i) & (!g141) & (!g135) & (g138) & (g152)) + ((sk[26]) & (!i) & (!g141) & (g135) & (g138) & (!g152)) + ((sk[26]) & (!i) & (!g141) & (g135) & (g138) & (g152)) + ((sk[26]) & (!i) & (g141) & (!g135) & (!g138) & (!g152)) + ((sk[26]) & (!i) & (g141) & (!g135) & (!g138) & (g152)) + ((sk[26]) & (!i) & (g141) & (!g135) & (g138) & (!g152)) + ((sk[26]) & (!i) & (g141) & (!g135) & (g138) & (g152)) + ((sk[26]) & (!i) & (g141) & (g135) & (!g138) & (!g152)) + ((sk[26]) & (!i) & (g141) & (g135) & (!g138) & (g152)) + ((sk[26]) & (!i) & (g141) & (g135) & (g138) & (!g152)) + ((sk[26]) & (!i) & (g141) & (g135) & (g138) & (g152)) + ((sk[26]) & (i) & (!g141) & (!g135) & (!g138) & (g152)) + ((sk[26]) & (i) & (!g141) & (!g135) & (g138) & (!g152)) + ((sk[26]) & (i) & (!g141) & (!g135) & (g138) & (g152)) + ((sk[26]) & (i) & (!g141) & (g135) & (!g138) & (g152)) + ((sk[26]) & (i) & (!g141) & (g135) & (g138) & (!g152)) + ((sk[26]) & (i) & (!g141) & (g135) & (g138) & (g152)) + ((sk[26]) & (i) & (g141) & (!g135) & (!g138) & (!g152)) + ((sk[26]) & (i) & (g141) & (!g135) & (!g138) & (g152)) + ((sk[26]) & (i) & (g141) & (!g135) & (g138) & (!g152)) + ((sk[26]) & (i) & (g141) & (!g135) & (g138) & (g152)) + ((sk[26]) & (i) & (g141) & (g135) & (!g138) & (!g152)) + ((sk[26]) & (i) & (g141) & (g135) & (!g138) & (g152)) + ((sk[26]) & (i) & (g141) & (g135) & (g138) & (!g152)) + ((sk[26]) & (i) & (g141) & (g135) & (g138) & (g152)));
	assign g168 = (((!k) & (!i) & (!sk[28]) & (j)) + ((!k) & (!i) & (sk[28]) & (!j)) + ((!k) & (i) & (!sk[28]) & (j)) + ((k) & (!i) & (!sk[28]) & (j)) + ((k) & (!i) & (sk[28]) & (!j)) + ((k) & (!i) & (sk[28]) & (j)) + ((k) & (i) & (!sk[28]) & (j)) + ((k) & (i) & (sk[28]) & (!j)));
	assign g169 = (((!c) & (!g92) & (!g93) & (d) & (!g141) & (g168)) + ((!c) & (!g92) & (g93) & (d) & (!g141) & (g168)) + ((!c) & (g92) & (!g93) & (!d) & (!g141) & (g168)) + ((!c) & (g92) & (!g93) & (d) & (!g141) & (g168)) + ((!c) & (g92) & (!g93) & (d) & (g141) & (g168)) + ((!c) & (g92) & (g93) & (d) & (!g141) & (g168)) + ((c) & (!g92) & (!g93) & (!d) & (!g141) & (g168)) + ((c) & (!g92) & (!g93) & (d) & (!g141) & (g168)) + ((c) & (!g92) & (!g93) & (d) & (g141) & (g168)) + ((c) & (!g92) & (g93) & (d) & (!g141) & (g168)) + ((c) & (g92) & (!g93) & (!d) & (!g141) & (g168)) + ((c) & (g92) & (!g93) & (d) & (!g141) & (g168)) + ((c) & (g92) & (!g93) & (d) & (g141) & (g168)) + ((c) & (g92) & (g93) & (!d) & (!g141) & (g168)) + ((c) & (g92) & (g93) & (d) & (!g141) & (g168)) + ((c) & (g92) & (g93) & (d) & (g141) & (g168)));
	assign g170 = (((!g7) & (!g15) & (!sk[29]) & (g17) & (!g121) & (!g135)) + ((!g7) & (!g15) & (!sk[29]) & (g17) & (g121) & (!g135)) + ((!g7) & (!g15) & (sk[29]) & (g17) & (!g121) & (!g135)) + ((!g7) & (!g15) & (sk[29]) & (g17) & (!g121) & (g135)) + ((!g7) & (!g15) & (sk[29]) & (g17) & (g121) & (!g135)) + ((!g7) & (!g15) & (sk[29]) & (g17) & (g121) & (g135)) + ((!g7) & (g15) & (!sk[29]) & (g17) & (!g121) & (!g135)) + ((!g7) & (g15) & (!sk[29]) & (g17) & (g121) & (!g135)) + ((!g7) & (g15) & (!sk[29]) & (g17) & (g121) & (g135)) + ((!g7) & (g15) & (sk[29]) & (!g17) & (!g121) & (!g135)) + ((!g7) & (g15) & (sk[29]) & (!g17) & (!g121) & (g135)) + ((!g7) & (g15) & (sk[29]) & (!g17) & (g121) & (!g135)) + ((!g7) & (g15) & (sk[29]) & (!g17) & (g121) & (g135)) + ((!g7) & (g15) & (sk[29]) & (g17) & (!g121) & (!g135)) + ((!g7) & (g15) & (sk[29]) & (g17) & (!g121) & (g135)) + ((!g7) & (g15) & (sk[29]) & (g17) & (g121) & (!g135)) + ((!g7) & (g15) & (sk[29]) & (g17) & (g121) & (g135)) + ((g7) & (!g15) & (!sk[29]) & (g17) & (!g121) & (!g135)) + ((g7) & (!g15) & (!sk[29]) & (g17) & (!g121) & (g135)) + ((g7) & (!g15) & (!sk[29]) & (g17) & (g121) & (!g135)) + ((g7) & (!g15) & (!sk[29]) & (g17) & (g121) & (g135)) + ((g7) & (!g15) & (sk[29]) & (g17) & (!g121) & (!g135)) + ((g7) & (!g15) & (sk[29]) & (g17) & (!g121) & (g135)) + ((g7) & (!g15) & (sk[29]) & (g17) & (g121) & (!g135)) + ((g7) & (!g15) & (sk[29]) & (g17) & (g121) & (g135)) + ((g7) & (g15) & (!sk[29]) & (g17) & (!g121) & (!g135)) + ((g7) & (g15) & (!sk[29]) & (g17) & (!g121) & (g135)) + ((g7) & (g15) & (!sk[29]) & (g17) & (g121) & (!g135)) + ((g7) & (g15) & (!sk[29]) & (g17) & (g121) & (g135)) + ((g7) & (g15) & (sk[29]) & (!g17) & (!g121) & (!g135)) + ((g7) & (g15) & (sk[29]) & (!g17) & (!g121) & (g135)) + ((g7) & (g15) & (sk[29]) & (!g17) & (g121) & (!g135)) + ((g7) & (g15) & (sk[29]) & (!g17) & (g121) & (g135)) + ((g7) & (g15) & (sk[29]) & (g17) & (!g121) & (!g135)) + ((g7) & (g15) & (sk[29]) & (g17) & (!g121) & (g135)) + ((g7) & (g15) & (sk[29]) & (g17) & (g121) & (!g135)) + ((g7) & (g15) & (sk[29]) & (g17) & (g121) & (g135)));
	assign g171 = (((!a) & (!sk[18]) & (!b) & (!c) & (d)) + ((!a) & (!sk[18]) & (!b) & (c) & (d)) + ((!a) & (!sk[18]) & (b) & (!c) & (!d)) + ((!a) & (!sk[18]) & (b) & (!c) & (d)) + ((!a) & (!sk[18]) & (b) & (c) & (!d)) + ((!a) & (!sk[18]) & (b) & (c) & (d)) + ((!a) & (sk[18]) & (!b) & (!c) & (!d)) + ((a) & (!sk[18]) & (!b) & (!c) & (!d)) + ((a) & (!sk[18]) & (!b) & (!c) & (d)) + ((a) & (!sk[18]) & (!b) & (c) & (!d)) + ((a) & (!sk[18]) & (!b) & (c) & (d)) + ((a) & (!sk[18]) & (b) & (!c) & (!d)) + ((a) & (!sk[18]) & (b) & (!c) & (d)) + ((a) & (!sk[18]) & (b) & (c) & (!d)) + ((a) & (!sk[18]) & (b) & (c) & (d)));
	assign g172 = (((!k) & (!g8) & (!g171) & (!sk[29]) & (g183)) + ((!k) & (!g8) & (g171) & (!sk[29]) & (g183)) + ((!k) & (!g8) & (g171) & (sk[29]) & (!g183)) + ((!k) & (!g8) & (g171) & (sk[29]) & (g183)) + ((!k) & (g8) & (!g171) & (!sk[29]) & (g183)) + ((!k) & (g8) & (g171) & (!sk[29]) & (g183)) + ((!k) & (g8) & (g171) & (sk[29]) & (!g183)) + ((!k) & (g8) & (g171) & (sk[29]) & (g183)) + ((k) & (!g8) & (g171) & (sk[29]) & (!g183)) + ((k) & (!g8) & (g171) & (sk[29]) & (g183)) + ((k) & (g8) & (g171) & (!sk[29]) & (!g183)) + ((k) & (g8) & (g171) & (!sk[29]) & (g183)) + ((k) & (g8) & (g171) & (sk[29]) & (!g183)) + ((k) & (g8) & (g171) & (sk[29]) & (g183)));
	assign g173 = (((!k) & (!l) & (i) & (sk[28]) & (j)) + ((!k) & (l) & (!i) & (!sk[28]) & (j)) + ((!k) & (l) & (i) & (!sk[28]) & (j)) + ((!k) & (l) & (i) & (sk[28]) & (j)) + ((k) & (!l) & (!i) & (!sk[28]) & (j)) + ((k) & (!l) & (!i) & (sk[28]) & (j)) + ((k) & (!l) & (i) & (!sk[28]) & (j)) + ((k) & (l) & (!i) & (!sk[28]) & (j)) + ((k) & (l) & (i) & (!sk[28]) & (j)));
	assign g174 = (((!sk[19]) & (g62) & (g93) & (g141) & (g173)) + ((sk[19]) & (!g62) & (!g93) & (g141) & (g173)) + ((sk[19]) & (!g62) & (g93) & (!g141) & (!g173)) + ((sk[19]) & (!g62) & (g93) & (!g141) & (g173)) + ((sk[19]) & (!g62) & (g93) & (g141) & (!g173)) + ((sk[19]) & (!g62) & (g93) & (g141) & (g173)) + ((sk[19]) & (g62) & (!g93) & (!g141) & (!g173)) + ((sk[19]) & (g62) & (!g93) & (!g141) & (g173)) + ((sk[19]) & (g62) & (!g93) & (g141) & (!g173)) + ((sk[19]) & (g62) & (!g93) & (g141) & (g173)) + ((sk[19]) & (g62) & (g93) & (!g141) & (!g173)) + ((sk[19]) & (g62) & (g93) & (!g141) & (g173)) + ((sk[19]) & (g62) & (g93) & (g141) & (!g173)) + ((sk[19]) & (g62) & (g93) & (g141) & (g173)));
	assign g175 = (((!l) & (!g139) & (!g169) & (!g170) & (!g172) & (!g174)) + ((!l) & (!g139) & (!g169) & (!g170) & (g172) & (!g174)) + ((!l) & (!g139) & (!g169) & (g170) & (!g172) & (!g174)) + ((!l) & (!g139) & (!g169) & (g170) & (g172) & (!g174)) + ((!l) & (!g139) & (g169) & (!g170) & (!g172) & (!g174)) + ((!l) & (!g139) & (g169) & (!g170) & (g172) & (!g174)) + ((!l) & (!g139) & (g169) & (g170) & (!g172) & (!g174)) + ((!l) & (!g139) & (g169) & (g170) & (g172) & (!g174)) + ((!l) & (g139) & (!g169) & (!g170) & (!g172) & (!g174)) + ((!l) & (g139) & (!g169) & (!g170) & (g172) & (!g174)) + ((!l) & (g139) & (!g169) & (g170) & (!g172) & (!g174)) + ((!l) & (g139) & (!g169) & (g170) & (g172) & (!g174)) + ((!l) & (g139) & (g169) & (!g170) & (!g172) & (!g174)) + ((!l) & (g139) & (g169) & (!g170) & (g172) & (!g174)) + ((!l) & (g139) & (g169) & (g170) & (!g172) & (!g174)) + ((!l) & (g139) & (g169) & (g170) & (g172) & (!g174)) + ((l) & (!g139) & (!g169) & (!g170) & (!g172) & (!g174)) + ((l) & (g139) & (!g169) & (!g170) & (!g172) & (!g174)) + ((l) & (g139) & (!g169) & (g170) & (!g172) & (!g174)));
	assign g176 = (((!j) & (!g1) & (!g165) & (!g166) & (!g167) & (g175)) + ((!j) & (!g1) & (!g165) & (!g166) & (g167) & (g175)) + ((!j) & (!g1) & (!g165) & (g166) & (!g167) & (g175)) + ((!j) & (!g1) & (!g165) & (g166) & (g167) & (g175)) + ((!j) & (!g1) & (g165) & (!g166) & (!g167) & (g175)) + ((!j) & (!g1) & (g165) & (!g166) & (g167) & (g175)) + ((!j) & (!g1) & (g165) & (g166) & (!g167) & (g175)) + ((!j) & (!g1) & (g165) & (g166) & (g167) & (g175)) + ((!j) & (g1) & (!g165) & (!g166) & (!g167) & (g175)) + ((j) & (!g1) & (!g165) & (!g166) & (!g167) & (g175)) + ((j) & (!g1) & (!g165) & (!g166) & (g167) & (g175)) + ((j) & (!g1) & (!g165) & (g166) & (!g167) & (g175)) + ((j) & (!g1) & (!g165) & (g166) & (g167) & (g175)) + ((j) & (!g1) & (g165) & (!g166) & (!g167) & (g175)) + ((j) & (!g1) & (g165) & (!g166) & (g167) & (g175)) + ((j) & (!g1) & (g165) & (g166) & (!g167) & (g175)) + ((j) & (!g1) & (g165) & (g166) & (g167) & (g175)) + ((j) & (g1) & (!g165) & (!g166) & (!g167) & (g175)) + ((j) & (g1) & (!g165) & (!g166) & (g167) & (g175)) + ((j) & (g1) & (!g165) & (g166) & (!g167) & (g175)) + ((j) & (g1) & (!g165) & (g166) & (g167) & (g175)) + ((j) & (g1) & (g165) & (!g166) & (!g167) & (g175)) + ((j) & (g1) & (g165) & (!g166) & (g167) & (g175)) + ((j) & (g1) & (g165) & (g166) & (!g167) & (g175)) + ((j) & (g1) & (g165) & (g166) & (g167) & (g175)));
	assign g178 = (((!a) & (!e) & (sk[21]) & (!g163)) + ((!a) & (e) & (!sk[21]) & (!g163)) + ((!a) & (e) & (!sk[21]) & (g163)) + ((a) & (!e) & (!sk[21]) & (g163)) + ((a) & (e) & (!sk[21]) & (!g163)) + ((a) & (e) & (!sk[21]) & (g163)) + ((a) & (e) & (sk[21]) & (!g163)));
	assign g179 = (((!f) & (!b) & (!c) & (!g) & (sk[18]) & (!g178)) + ((!f) & (!b) & (!c) & (g) & (!sk[18]) & (!g178)) + ((!f) & (!b) & (!c) & (g) & (!sk[18]) & (g178)) + ((!f) & (!b) & (!c) & (g) & (sk[18]) & (!g178)) + ((!f) & (!b) & (!c) & (g) & (sk[18]) & (g178)) + ((!f) & (!b) & (c) & (!g) & (!sk[18]) & (!g178)) + ((!f) & (!b) & (c) & (!g) & (!sk[18]) & (g178)) + ((!f) & (!b) & (c) & (!g) & (sk[18]) & (!g178)) + ((!f) & (!b) & (c) & (!g) & (sk[18]) & (g178)) + ((!f) & (!b) & (c) & (g) & (!sk[18]) & (!g178)) + ((!f) & (!b) & (c) & (g) & (!sk[18]) & (g178)) + ((!f) & (!b) & (c) & (g) & (sk[18]) & (!g178)) + ((!f) & (b) & (!c) & (!g) & (sk[18]) & (!g178)) + ((!f) & (b) & (!c) & (!g) & (sk[18]) & (g178)) + ((!f) & (b) & (!c) & (g) & (!sk[18]) & (!g178)) + ((!f) & (b) & (!c) & (g) & (!sk[18]) & (g178)) + ((!f) & (b) & (!c) & (g) & (sk[18]) & (!g178)) + ((!f) & (b) & (!c) & (g) & (sk[18]) & (g178)) + ((!f) & (b) & (c) & (!g) & (!sk[18]) & (!g178)) + ((!f) & (b) & (c) & (!g) & (!sk[18]) & (g178)) + ((!f) & (b) & (c) & (!g) & (sk[18]) & (!g178)) + ((!f) & (b) & (c) & (!g) & (sk[18]) & (g178)) + ((!f) & (b) & (c) & (g) & (!sk[18]) & (!g178)) + ((!f) & (b) & (c) & (g) & (!sk[18]) & (g178)) + ((!f) & (b) & (c) & (g) & (sk[18]) & (!g178)) + ((!f) & (b) & (c) & (g) & (sk[18]) & (g178)) + ((f) & (!b) & (!c) & (!g) & (!sk[18]) & (!g178)) + ((f) & (!b) & (!c) & (!g) & (!sk[18]) & (g178)) + ((f) & (!b) & (!c) & (!g) & (sk[18]) & (!g178)) + ((f) & (!b) & (!c) & (!g) & (sk[18]) & (g178)) + ((f) & (!b) & (!c) & (g) & (!sk[18]) & (!g178)) + ((f) & (!b) & (!c) & (g) & (!sk[18]) & (g178)) + ((f) & (!b) & (!c) & (g) & (sk[18]) & (!g178)) + ((f) & (!b) & (!c) & (g) & (sk[18]) & (g178)) + ((f) & (!b) & (c) & (!g) & (!sk[18]) & (!g178)) + ((f) & (!b) & (c) & (!g) & (!sk[18]) & (g178)) + ((f) & (!b) & (c) & (!g) & (sk[18]) & (!g178)) + ((f) & (!b) & (c) & (!g) & (sk[18]) & (g178)) + ((f) & (!b) & (c) & (g) & (!sk[18]) & (!g178)) + ((f) & (!b) & (c) & (g) & (!sk[18]) & (g178)) + ((f) & (!b) & (c) & (g) & (sk[18]) & (!g178)) + ((f) & (!b) & (c) & (g) & (sk[18]) & (g178)) + ((f) & (b) & (!c) & (!g) & (!sk[18]) & (!g178)) + ((f) & (b) & (!c) & (!g) & (!sk[18]) & (g178)) + ((f) & (b) & (!c) & (!g) & (sk[18]) & (!g178)) + ((f) & (b) & (!c) & (g) & (!sk[18]) & (!g178)) + ((f) & (b) & (!c) & (g) & (!sk[18]) & (g178)) + ((f) & (b) & (!c) & (g) & (sk[18]) & (!g178)) + ((f) & (b) & (!c) & (g) & (sk[18]) & (g178)) + ((f) & (b) & (c) & (!g) & (!sk[18]) & (!g178)) + ((f) & (b) & (c) & (!g) & (!sk[18]) & (g178)) + ((f) & (b) & (c) & (!g) & (sk[18]) & (!g178)) + ((f) & (b) & (c) & (!g) & (sk[18]) & (g178)) + ((f) & (b) & (c) & (g) & (!sk[18]) & (!g178)) + ((f) & (b) & (c) & (g) & (!sk[18]) & (g178)) + ((f) & (b) & (c) & (g) & (sk[18]) & (!g178)));
	assign g180 = (((!l) & (!k) & (!e) & (!a) & (!j) & (!n)) + ((!l) & (!k) & (!e) & (!a) & (j) & (!n)) + ((!l) & (!k) & (!e) & (!a) & (j) & (n)) + ((!l) & (!k) & (!e) & (a) & (j) & (n)) + ((!l) & (!k) & (e) & (!a) & (!j) & (!n)) + ((!l) & (!k) & (e) & (!a) & (j) & (!n)) + ((!l) & (k) & (!e) & (a) & (j) & (n)) + ((!l) & (k) & (e) & (!a) & (j) & (n)) + ((!l) & (k) & (e) & (a) & (!j) & (!n)) + ((!l) & (k) & (e) & (a) & (!j) & (n)) + ((l) & (!k) & (!e) & (!a) & (!j) & (!n)) + ((l) & (!k) & (!e) & (!a) & (j) & (n)) + ((l) & (!k) & (!e) & (a) & (j) & (n)) + ((l) & (!k) & (e) & (!a) & (!j) & (!n)) + ((l) & (!k) & (e) & (a) & (!j) & (n)) + ((l) & (k) & (!e) & (!a) & (j) & (n)) + ((l) & (k) & (!e) & (a) & (j) & (n)));
	assign g181 = (((!l) & (!k) & (!e) & (a) & (!j) & (!n)) + ((!l) & (!k) & (e) & (!a) & (!j) & (!n)) + ((!l) & (!k) & (e) & (a) & (!j) & (!n)) + ((!l) & (k) & (!e) & (!a) & (j) & (!n)) + ((!l) & (k) & (!e) & (!a) & (j) & (n)) + ((!l) & (k) & (!e) & (a) & (!j) & (n)) + ((!l) & (k) & (!e) & (a) & (j) & (!n)) + ((!l) & (k) & (!e) & (a) & (j) & (n)) + ((!l) & (k) & (e) & (!a) & (!j) & (n)) + ((!l) & (k) & (e) & (a) & (!j) & (n)) + ((l) & (!k) & (e) & (a) & (j) & (n)) + ((l) & (k) & (!e) & (!a) & (!j) & (!n)) + ((l) & (k) & (!e) & (a) & (!j) & (!n)) + ((l) & (k) & (!e) & (a) & (!j) & (n)) + ((l) & (k) & (e) & (!a) & (!j) & (n)) + ((l) & (k) & (e) & (a) & (!j) & (n)));
	assign g183 = (((!sk[29]) & (!g184) & (!g185)));
	assign g184 = (((!sk[30]) & (!k) & (g186)) + ((sk[30]) & (k) & (!g186)) + ((sk[30]) & (k) & (g186)));
	assign g185 = (((!sk[30]) & (k) & (g189)) + ((sk[30]) & (!k) & (g189)) + ((sk[30]) & (k) & (g189)));
	assign g186 = (((!sk[30]) & (!g187) & (!g188)));
	assign g187 = (((!sk[28]) & (j) & (!g190)) + ((!sk[28]) & (j) & (g190)) + ((sk[28]) & (!j) & (g190)));
	assign g188 = (((!sk[30]) & (j) & (g191)) + ((sk[30]) & (j) & (!g191)) + ((sk[30]) & (j) & (g191)));
	assign g189 = (((!sk[30]) & (!j) & (g192)) + ((sk[30]) & (j) & (!g192)) + ((sk[30]) & (j) & (g192)));
	assign g190 = (((!h) & (!d) & (!g147) & (!sk[27]) & (i)) + ((!h) & (!d) & (g147) & (!sk[27]) & (!i)) + ((!h) & (!d) & (g147) & (!sk[27]) & (i)) + ((!h) & (d) & (!g147) & (!sk[27]) & (!i)) + ((!h) & (d) & (!g147) & (!sk[27]) & (i)) + ((!h) & (d) & (g147) & (!sk[27]) & (!i)) + ((!h) & (d) & (g147) & (!sk[27]) & (i)) + ((!h) & (d) & (g147) & (sk[27]) & (i)) + ((h) & (!d) & (!g147) & (!sk[27]) & (i)) + ((h) & (!d) & (g147) & (!sk[27]) & (!i)) + ((h) & (!d) & (g147) & (!sk[27]) & (i)) + ((h) & (!d) & (g147) & (sk[27]) & (i)) + ((h) & (d) & (!g147) & (!sk[27]) & (!i)) + ((h) & (d) & (!g147) & (!sk[27]) & (i)) + ((h) & (d) & (!g147) & (sk[27]) & (i)) + ((h) & (d) & (g147) & (!sk[27]) & (!i)) + ((h) & (d) & (g147) & (!sk[27]) & (i)) + ((h) & (d) & (g147) & (sk[27]) & (i)));
	assign g191 = (((!h) & (!d) & (!sk[27]) & (!g12) & (i)) + ((!h) & (!d) & (!sk[27]) & (g12) & (!i)) + ((!h) & (!d) & (!sk[27]) & (g12) & (i)) + ((!h) & (d) & (!sk[27]) & (!g12) & (i)) + ((!h) & (d) & (!sk[27]) & (g12) & (!i)) + ((!h) & (d) & (!sk[27]) & (g12) & (i)) + ((h) & (!d) & (!sk[27]) & (!g12) & (!i)) + ((h) & (!d) & (!sk[27]) & (!g12) & (i)) + ((h) & (!d) & (!sk[27]) & (g12) & (!i)) + ((h) & (!d) & (!sk[27]) & (g12) & (i)) + ((h) & (d) & (!sk[27]) & (!g12) & (!i)) + ((h) & (d) & (!sk[27]) & (!g12) & (i)) + ((h) & (d) & (!sk[27]) & (g12) & (!i)) + ((h) & (d) & (!sk[27]) & (g12) & (i)) + ((h) & (d) & (sk[27]) & (g12) & (!i)));
	assign g192 = (((!h) & (!d) & (!sk[27]) & (g147) & (!i)) + ((!h) & (!d) & (!sk[27]) & (g147) & (i)) + ((!h) & (d) & (!sk[27]) & (!g147) & (!i)) + ((!h) & (d) & (!sk[27]) & (!g147) & (i)) + ((!h) & (d) & (!sk[27]) & (g147) & (!i)) + ((!h) & (d) & (!sk[27]) & (g147) & (i)) + ((!h) & (d) & (sk[27]) & (g147) & (i)) + ((h) & (!d) & (!sk[27]) & (!g147) & (i)) + ((h) & (!d) & (!sk[27]) & (g147) & (!i)) + ((h) & (!d) & (!sk[27]) & (g147) & (i)) + ((h) & (!d) & (sk[27]) & (g147) & (i)) + ((h) & (d) & (!sk[27]) & (!g147) & (!i)) + ((h) & (d) & (!sk[27]) & (!g147) & (i)) + ((h) & (d) & (!sk[27]) & (g147) & (!i)) + ((h) & (d) & (!sk[27]) & (g147) & (i)) + ((h) & (d) & (sk[27]) & (!g147) & (i)) + ((h) & (d) & (sk[27]) & (g147) & (i)));
	assign g194 = (((!sk[31]) & (!n) & (g196)) + ((!sk[31]) & (n) & (g196)) + ((sk[31]) & (!n) & (g196)));
	assign g195 = (((!sk[31]) & (n) & (!g199)) + ((!sk[31]) & (n) & (g199)) + ((sk[31]) & (n) & (g199)));
	assign g196 = (((!sk[32]) & (!g197) & (!g198)));
	assign g197 = (((!j) & (!sk[32]) & (g202)) + ((!j) & (sk[32]) & (g202)) + ((j) & (sk[32]) & (g202)));
	assign g198 = (((!j) & (sk[32]) & (g203)) + ((j) & (!sk[32]) & (g203)) + ((j) & (sk[32]) & (g203)));
	assign g199 = (((!sk[32]) & (!g200) & (!g201)));
	assign g200 = (((!j) & (!sk[32]) & (g204)) + ((j) & (sk[32]) & (g204)));
	assign g201 = (((!j) & (!sk[33]) & (g205)) + ((j) & (!sk[33]) & (g205)) + ((j) & (sk[33]) & (g205)));
	assign g202 = (((!sk[34]) & (g119) & (!g116)) + ((!sk[34]) & (g119) & (g116)) + ((sk[34]) & (!g119) & (g116)) + ((sk[34]) & (g119) & (!g116)) + ((sk[34]) & (g119) & (g116)));
	assign g203 = (((!g119) & (!sk[34]) & (g117)) + ((!g119) & (sk[34]) & (g117)) + ((g119) & (!sk[34]) & (g117)) + ((g119) & (sk[34]) & (!g117)) + ((g119) & (sk[34]) & (g117)));
	assign g204 = (((!sk[34]) & (!g119) & (!g115) & (g80)) + ((!sk[34]) & (!g119) & (g115) & (!g80)) + ((!sk[34]) & (!g119) & (g115) & (g80)) + ((!sk[34]) & (g119) & (!g115) & (g80)) + ((!sk[34]) & (g119) & (g115) & (!g80)) + ((!sk[34]) & (g119) & (g115) & (g80)) + ((sk[34]) & (!g119) & (!g115) & (!g80)) + ((sk[34]) & (!g119) & (g115) & (g80)) + ((sk[34]) & (g119) & (!g115) & (!g80)) + ((sk[34]) & (g119) & (!g115) & (g80)) + ((sk[34]) & (g119) & (g115) & (!g80)) + ((sk[34]) & (g119) & (g115) & (g80)));
	assign g205 = (((!g119) & (sk[34]) & (!g115) & (!g80)) + ((!g119) & (sk[34]) & (g115) & (g80)) + ((g119) & (!sk[34]) & (!g115) & (!g80)) + ((g119) & (!sk[34]) & (!g115) & (g80)) + ((g119) & (!sk[34]) & (g115) & (!g80)) + ((g119) & (!sk[34]) & (g115) & (g80)) + ((g119) & (sk[34]) & (!g115) & (!g80)) + ((g119) & (sk[34]) & (!g115) & (g80)) + ((g119) & (sk[34]) & (g115) & (!g80)) + ((g119) & (sk[34]) & (g115) & (g80)));
	assign g206 = (((!g207) & (sk[34]) & (!g208)) + ((g207) & (!sk[34]) & (!g208)) + ((g207) & (!sk[34]) & (g208)));
	assign g207 = (((!g50) & (!sk[35]) & (g209)) + ((!g50) & (sk[35]) & (g209)) + ((g50) & (sk[35]) & (g209)));
	assign g208 = (((!g50) & (sk[35]) & (g212)) + ((g50) & (!sk[35]) & (g212)) + ((g50) & (sk[35]) & (g212)));
	assign g209 = (((!sk[35]) & (!g210) & (!g211)));
	assign g210 = (((!b) & (!sk[35]) & (g215)) + ((!b) & (sk[35]) & (g215)) + ((b) & (sk[35]) & (g215)));
	assign g211 = (((b) & (!sk[35]) & (g216)) + ((b) & (sk[35]) & (!g216)) + ((b) & (sk[35]) & (g216)));
	assign g212 = (((!sk[36]) & (!g213) & (!g214)));
	assign g213 = (((!b) & (!sk[36]) & (g217)) + ((!b) & (sk[36]) & (g217)) + ((b) & (sk[36]) & (g217)));
	assign g214 = (((!sk[36]) & (b) & (g218)) + ((sk[36]) & (!b) & (g218)) + ((sk[36]) & (b) & (g218)));
	assign g215 = (((!g56) & (!sk[36]) & (g51) & (g44)) + ((!g56) & (sk[36]) & (g51) & (!g44)) + ((!g56) & (sk[36]) & (g51) & (g44)) + ((g56) & (!sk[36]) & (!g51) & (g44)) + ((g56) & (!sk[36]) & (g51) & (g44)) + ((g56) & (sk[36]) & (g51) & (!g44)) + ((g56) & (sk[36]) & (g51) & (g44)));
	assign g216 = (((!g56) & (!g57) & (g53) & (!sk[36]) & (!g44)) + ((!g56) & (g57) & (!g53) & (!sk[36]) & (!g44)) + ((!g56) & (g57) & (!g53) & (!sk[36]) & (g44)) + ((!g56) & (g57) & (!g53) & (sk[36]) & (!g44)) + ((!g56) & (g57) & (!g53) & (sk[36]) & (g44)) + ((!g56) & (g57) & (g53) & (!sk[36]) & (!g44)) + ((!g56) & (g57) & (g53) & (!sk[36]) & (g44)) + ((!g56) & (g57) & (g53) & (sk[36]) & (!g44)) + ((!g56) & (g57) & (g53) & (sk[36]) & (g44)) + ((g56) & (!g57) & (!g53) & (!sk[36]) & (g44)) + ((g56) & (!g57) & (!g53) & (sk[36]) & (!g44)) + ((g56) & (!g57) & (!g53) & (sk[36]) & (g44)) + ((g56) & (!g57) & (g53) & (!sk[36]) & (!g44)) + ((g56) & (!g57) & (g53) & (!sk[36]) & (g44)) + ((g56) & (!g57) & (g53) & (sk[36]) & (!g44)) + ((g56) & (!g57) & (g53) & (sk[36]) & (g44)) + ((g56) & (g57) & (!g53) & (!sk[36]) & (!g44)) + ((g56) & (g57) & (!g53) & (!sk[36]) & (g44)) + ((g56) & (g57) & (!g53) & (sk[36]) & (!g44)) + ((g56) & (g57) & (!g53) & (sk[36]) & (g44)) + ((g56) & (g57) & (g53) & (!sk[36]) & (!g44)) + ((g56) & (g57) & (g53) & (!sk[36]) & (g44)) + ((g56) & (g57) & (g53) & (sk[36]) & (!g44)) + ((g56) & (g57) & (g53) & (sk[36]) & (g44)));
	assign g217 = (((!sk[37]) & (!g56) & (g44)) + ((!sk[37]) & (g56) & (g44)) + ((sk[37]) & (g56) & (g44)));
	assign g218 = (((!g56) & (!g57) & (!sk[37]) & (!g53) & (g44)) + ((!g56) & (!g57) & (!sk[37]) & (g53) & (g44)) + ((!g56) & (!g57) & (sk[37]) & (g53) & (g44)) + ((!g56) & (g57) & (!sk[37]) & (!g53) & (g44)) + ((!g56) & (g57) & (!sk[37]) & (g53) & (!g44)) + ((!g56) & (g57) & (!sk[37]) & (g53) & (g44)) + ((!g56) & (g57) & (sk[37]) & (!g53) & (!g44)) + ((!g56) & (g57) & (sk[37]) & (!g53) & (g44)) + ((!g56) & (g57) & (sk[37]) & (g53) & (!g44)) + ((!g56) & (g57) & (sk[37]) & (g53) & (g44)) + ((g56) & (!g57) & (!sk[37]) & (!g53) & (!g44)) + ((g56) & (!g57) & (!sk[37]) & (!g53) & (g44)) + ((g56) & (!g57) & (!sk[37]) & (g53) & (!g44)) + ((g56) & (!g57) & (!sk[37]) & (g53) & (g44)) + ((g56) & (!g57) & (sk[37]) & (!g53) & (g44)) + ((g56) & (!g57) & (sk[37]) & (g53) & (g44)) + ((g56) & (g57) & (!sk[37]) & (!g53) & (!g44)) + ((g56) & (g57) & (!sk[37]) & (!g53) & (g44)) + ((g56) & (g57) & (!sk[37]) & (g53) & (!g44)) + ((g56) & (g57) & (!sk[37]) & (g53) & (g44)) + ((g56) & (g57) & (sk[37]) & (!g53) & (!g44)) + ((g56) & (g57) & (sk[37]) & (!g53) & (g44)) + ((g56) & (g57) & (sk[37]) & (g53) & (!g44)) + ((g56) & (g57) & (sk[37]) & (g53) & (g44)));
	assign g220 = (((!sk[31]) & (!n) & (g222)) + ((!sk[31]) & (n) & (g222)) + ((sk[31]) & (!n) & (g222)));
	assign g221 = (((!sk[31]) & (n) & (!g225)) + ((!sk[31]) & (n) & (g225)) + ((sk[31]) & (n) & (g225)));
	assign g222 = (((!sk[37]) & (g223) & (!g224)) + ((!sk[37]) & (g223) & (g224)) + ((sk[37]) & (!g223) & (!g224)));
	assign g223 = (((!sk[33]) & (!j) & (g228)) + ((!sk[33]) & (j) & (g228)) + ((sk[33]) & (!j) & (g228)));
	assign g224 = (((j) & (!sk[33]) & (!g229)) + ((j) & (!sk[33]) & (g229)) + ((j) & (sk[33]) & (g229)));
	assign g225 = (((!sk[37]) & (!g226) & (g227)) + ((!sk[37]) & (g226) & (g227)) + ((sk[37]) & (!g226) & (!g227)));
	assign g226 = (((!j) & (sk[33]) & (g230)) + ((j) & (!sk[33]) & (!g230)) + ((j) & (!sk[33]) & (g230)));
	assign g227 = (((j) & (!sk[33]) & (!g231)) + ((j) & (!sk[33]) & (g231)) + ((j) & (sk[33]) & (g231)));
	assign g228 = (((!g37) & (sk[37]) & (g5)) + ((g37) & (!sk[37]) & (!g5)) + ((g37) & (!sk[37]) & (g5)) + ((g37) & (sk[37]) & (!g5)) + ((g37) & (sk[37]) & (g5)));
	assign g229 = (((!g37) & (sk[38]) & (g6)) + ((g37) & (!sk[38]) & (!g6)) + ((g37) & (!sk[38]) & (g6)) + ((g37) & (sk[38]) & (!g6)) + ((g37) & (sk[38]) & (g6)));
	assign g230 = (((!g37) & (!g31) & (!sk[13]) & (!m)) + ((!g37) & (g31) & (!sk[13]) & (m)) + ((g37) & (!g31) & (!sk[13]) & (!m)) + ((g37) & (!g31) & (!sk[13]) & (m)) + ((g37) & (g31) & (!sk[13]) & (!m)) + ((g37) & (g31) & (!sk[13]) & (m)));
	assign g231 = (((!g37) & (!g31) & (!sk[13]) & (!m)) + ((!g37) & (g31) & (!sk[13]) & (m)) + ((g37) & (!g31) & (!sk[13]) & (!m)) + ((g37) & (!g31) & (!sk[13]) & (m)) + ((g37) & (g31) & (!sk[13]) & (!m)) + ((g37) & (g31) & (!sk[13]) & (m)));
	assign s = (((sk[38]) & (!g163)));
	assign t = (((sk[38]) & (g121)));
	assign v = (((sk[38]) & (!g179)));
	assign p = (((!n) & (!m) & (!g31) & (!g73) & (!sk[13]) & (!g78)) + ((!n) & (!m) & (!g31) & (g73) & (!sk[13]) & (!g78)) + ((!n) & (!m) & (g31) & (!g73) & (!sk[13]) & (!g78)) + ((!n) & (!m) & (g31) & (g73) & (!sk[13]) & (!g78)) + ((!n) & (m) & (!g31) & (!g73) & (!sk[13]) & (!g78)) + ((!n) & (m) & (!g31) & (g73) & (!sk[13]) & (!g78)) + ((!n) & (m) & (g31) & (!g73) & (!sk[13]) & (!g78)) + ((!n) & (m) & (g31) & (g73) & (!sk[13]) & (!g78)) + ((n) & (!m) & (!g31) & (!g73) & (!sk[13]) & (!g78)) + ((n) & (!m) & (!g31) & (!g73) & (!sk[13]) & (g78)) + ((n) & (!m) & (!g31) & (g73) & (!sk[13]) & (!g78)) + ((n) & (!m) & (g31) & (!g73) & (!sk[13]) & (!g78)) + ((n) & (!m) & (g31) & (g73) & (!sk[13]) & (!g78)) + ((n) & (!m) & (g31) & (g73) & (!sk[13]) & (g78)) + ((n) & (m) & (!g31) & (!g73) & (!sk[13]) & (!g78)) + ((n) & (m) & (!g31) & (!g73) & (!sk[13]) & (g78)) + ((n) & (m) & (!g31) & (g73) & (!sk[13]) & (!g78)) + ((n) & (m) & (g31) & (!g73) & (!sk[13]) & (!g78)) + ((n) & (m) & (g31) & (!g73) & (!sk[13]) & (g78)) + ((n) & (m) & (g31) & (g73) & (!sk[13]) & (!g78)));
	assign r = (((!sk[31]) & (!n) & (g80) & (!g115) & (!g156) & (!g161)) + ((!sk[31]) & (!n) & (g80) & (!g115) & (!g156) & (g161)) + ((!sk[31]) & (!n) & (g80) & (!g115) & (g156) & (!g161)) + ((!sk[31]) & (!n) & (g80) & (!g115) & (g156) & (g161)) + ((!sk[31]) & (!n) & (g80) & (g115) & (!g156) & (!g161)) + ((!sk[31]) & (!n) & (g80) & (g115) & (!g156) & (g161)) + ((!sk[31]) & (!n) & (g80) & (g115) & (g156) & (!g161)) + ((!sk[31]) & (!n) & (g80) & (g115) & (g156) & (g161)) + ((!sk[31]) & (n) & (!g80) & (!g115) & (g156) & (!g161)) + ((!sk[31]) & (n) & (!g80) & (!g115) & (g156) & (g161)) + ((!sk[31]) & (n) & (!g80) & (g115) & (g156) & (!g161)) + ((!sk[31]) & (n) & (!g80) & (g115) & (g156) & (g161)) + ((!sk[31]) & (n) & (g80) & (!g115) & (!g156) & (!g161)) + ((!sk[31]) & (n) & (g80) & (!g115) & (!g156) & (g161)) + ((!sk[31]) & (n) & (g80) & (!g115) & (g156) & (!g161)) + ((!sk[31]) & (n) & (g80) & (!g115) & (g156) & (g161)) + ((!sk[31]) & (n) & (g80) & (g115) & (!g156) & (!g161)) + ((!sk[31]) & (n) & (g80) & (g115) & (!g156) & (g161)) + ((!sk[31]) & (n) & (g80) & (g115) & (g156) & (!g161)) + ((!sk[31]) & (n) & (g80) & (g115) & (g156) & (g161)) + ((sk[31]) & (!n) & (!g80) & (!g115) & (!g156) & (!g161)) + ((sk[31]) & (!n) & (!g80) & (!g115) & (g156) & (!g161)) + ((sk[31]) & (!n) & (!g80) & (g115) & (!g156) & (!g161)) + ((sk[31]) & (!n) & (!g80) & (g115) & (g156) & (!g161)) + ((sk[31]) & (!n) & (g80) & (!g115) & (!g156) & (!g161)) + ((sk[31]) & (!n) & (g80) & (!g115) & (g156) & (!g161)) + ((sk[31]) & (!n) & (g80) & (g115) & (!g156) & (!g161)) + ((sk[31]) & (!n) & (g80) & (g115) & (g156) & (!g161)) + ((sk[31]) & (n) & (!g80) & (!g115) & (!g156) & (!g161)) + ((sk[31]) & (n) & (!g80) & (!g115) & (!g156) & (g161)) + ((sk[31]) & (n) & (!g80) & (!g115) & (g156) & (!g161)) + ((sk[31]) & (n) & (!g80) & (g115) & (!g156) & (!g161)) + ((sk[31]) & (n) & (!g80) & (g115) & (g156) & (!g161)) + ((sk[31]) & (n) & (!g80) & (g115) & (g156) & (g161)) + ((sk[31]) & (n) & (g80) & (!g115) & (!g156) & (!g161)) + ((sk[31]) & (n) & (g80) & (!g115) & (!g156) & (g161)) + ((sk[31]) & (n) & (g80) & (!g115) & (g156) & (!g161)) + ((sk[31]) & (n) & (g80) & (g115) & (!g156) & (!g161)) + ((sk[31]) & (n) & (g80) & (g115) & (!g156) & (g161)) + ((sk[31]) & (n) & (g80) & (g115) & (g156) & (!g161)));
	assign u = (((n) & (!g80) & (!g115) & (!g156) & (!g164) & (!g176)) + ((n) & (!g80) & (!g115) & (!g156) & (g164) & (!g176)) + ((n) & (!g80) & (!g115) & (!g156) & (g164) & (g176)) + ((n) & (!g80) & (!g115) & (g156) & (!g164) & (!g176)) + ((n) & (!g80) & (!g115) & (g156) & (g164) & (!g176)) + ((n) & (!g80) & (!g115) & (g156) & (g164) & (g176)) + ((n) & (!g80) & (g115) & (!g156) & (!g164) & (!g176)) + ((n) & (!g80) & (g115) & (!g156) & (!g164) & (g176)) + ((n) & (!g80) & (g115) & (!g156) & (g164) & (!g176)) + ((n) & (!g80) & (g115) & (!g156) & (g164) & (g176)) + ((n) & (!g80) & (g115) & (g156) & (!g164) & (!g176)) + ((n) & (!g80) & (g115) & (g156) & (g164) & (!g176)) + ((n) & (!g80) & (g115) & (g156) & (g164) & (g176)) + ((n) & (g80) & (!g115) & (!g156) & (!g164) & (!g176)) + ((n) & (g80) & (!g115) & (!g156) & (g164) & (!g176)) + ((n) & (g80) & (!g115) & (!g156) & (g164) & (g176)) + ((n) & (g80) & (!g115) & (g156) & (!g164) & (!g176)) + ((n) & (g80) & (!g115) & (g156) & (g164) & (!g176)) + ((n) & (g80) & (!g115) & (g156) & (g164) & (g176)) + ((n) & (g80) & (g115) & (!g156) & (!g164) & (!g176)) + ((n) & (g80) & (g115) & (!g156) & (g164) & (!g176)) + ((n) & (g80) & (g115) & (!g156) & (g164) & (g176)) + ((n) & (g80) & (g115) & (g156) & (!g164) & (!g176)) + ((n) & (g80) & (g115) & (g156) & (g164) & (!g176)) + ((n) & (g80) & (g115) & (g156) & (g164) & (g176)));
	assign q = (((!g194) & (sk[38]) & (!g195)) + ((g194) & (!sk[38]) & (!g195)) + ((g194) & (!sk[38]) & (g195)));
	assign o = (((!g220) & (!sk[39]) & (!g221)));
endmodule
