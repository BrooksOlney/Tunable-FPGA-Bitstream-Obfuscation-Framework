module ks_ex1010_qmap_map (sk, i_9_, i_2_, i_0_, i_1_, i_8_, i_6_, i_7_, i_5_, i_3_, i_4_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_);

	input i_9_;
	input i_2_;
	input i_0_;
	input i_1_;
	input i_8_;
	input i_6_;
	input i_7_;
	input i_5_;
	input i_3_;
	input i_4_;
	output o_0_;
	output o_1_;
	output o_2_;
	output o_3_;
	output o_4_;
	output o_5_;
	output o_6_;
	output o_7_;
	output o_8_;
	output o_9_;

	input [127 : 0] sk /* synthesis noprune */;


	wire g217, g298, g364, g431, g486, g542, g585, g627, g662, g689, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11;
	wire g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32;
	wire g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g52, g53;
	wire g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73, g74;
	wire g75, g76, g77, g78, g79, g80, g81, g82, g83, g84, g85, g86, g765, g87, g88, g787, g774, g89, g90, g91, g92;
	wire g93, g94, g95, g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113;
	wire g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134;
	wire g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155;
	wire g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g170, g171, g172, g747, g173, g174, g175;
	wire g176, g177, g178, g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195, g196;
	wire g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207, g208, g209, g210, g211, g212, g213, g214, g215, g216, g758;
	wire g218, g219, g220, g221, g222, g223, g224, g225, g226, g227, g228, g229, g230, g231, g232, g233, g234, g235, g236, g237, g238;
	wire g239, g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250, g251, g252, g253, g254, g255, g256, g257, g258, g259;
	wire g260, g261, g262, g263, g264, g265, g266, g267, g268, g269, g270, g271, g272, g273, g274, g275, g276, g277, g278, g279, g280;
	wire g281, g282, g283, g284, g285, g286, g287, g288, g289, g729, g290, g291, g292, g293, g294, g295, g296, g722, g297, g735, g299;
	wire g300, g301, g302, g303, g304, g305, g306, g307, g308, g309, g310, g311, g312, g313, g314, g315, g316, g317, g318, g319, g320;
	wire g321, g322, g323, g324, g325, g326, g327, g328, g329, g330, g331, g332, g333, g334, g335, g336, g337, g338, g339, g340, g341;
	wire g342, g343, g344, g345, g346, g347, g348, g349, g350, g351, g352, g353, g354, g355, g356, g357, g358, g359, g360, g711, g361;
	wire g362, g363, g365, g366, g367, g368, g369, g370, g371, g372, g373, g374, g375, g376, g377, g378, g379, g380, g381, g382, g383;
	wire g384, g385, g386, g387, g388, g389, g390, g391, g392, g393, g394, g395, g396, g397, g398, g399, g400, g401, g402, g403, g404;
	wire g405, g406, g407, g408, g409, g410, g411, g412, g413, g414, g415, g416, g417, g418, g419, g420, g421, g422, g423, g424, g425;
	wire g426, g427, g428, g429, g430, g432, g433, g434, g435, g436, g437, g438, g439, g440, g441, g442, g443, g444, g445, g446, g447;
	wire g448, g449, g450, g451, g452, g453, g454, g455, g456, g457, g458, g459, g460, g461, g462, g463, g464, g465, g466, g467, g468;
	wire g469, g470, g471, g472, g473, g474, g475, g476, g477, g478, g479, g480, g481, g482, g483, g704, g484, g485, g487, g488, g489;
	wire g490, g491, g492, g493, g494, g495, g496, g497, g498, g499, g500, g501, g502, g503, g504, g505, g506, g507, g508, g509, g510;
	wire g511, g512, g513, g514, g515, g516, g517, g518, g519, g520, g521, g522, g523, g524, g525, g526, g527, g528, g529, g530, g531;
	wire g532, g533, g534, g535, g536, g537, g538, g697, g539, g540, g541, g543, g544, g545, g546, g690, g547, g548, g549, g550, g551;
	wire g552, g553, g554, g555, g556, g557, g558, g559, g560, g561, g562, g563, g564, g565, g566, g567, g568, g569, g570, g571, g572;
	wire g573, g574, g575, g576, g577, g578, g579, g580, g581, g582, g583, g584, g586, g587, g588, g589, g590, g591, g592, g593, g594;
	wire g595, g596, g597, g598, g599, g600, g601, g602, g603, g604, g605, g606, g607, g608, g609, g610, g611, g612, g613, g614, g615;
	wire g616, g617, g618, g619, g620, g621, g622, g623, g624, g625, g626, g628, g629, g630, g631, g632, g633, g634, g635, g636, g637;
	wire g638, g639, g640, g641, g642, g643, g644, g645, g646, g647, g648, g649, g650, g651, g652, g653, g654, g655, g656, g657, g658;
	wire g659, g660, g661, g663, g664, g665, g666, g667, g668, g669, g670, g671, g672, g673, g674, g675, g676, g677, g678, g679, g680;
	wire g681, g682, g683, g684, g685, g686, g687, g688, g691, g692, g693, g694, g695, g696, g698, g699, g700, g701, g702, g703, g705;
	wire g706, g707, g708, g709, g710, g712, g713, g714, g717, g715, g716, g719, g720, g718, g721, g723, g724, g725, g726, g727, g728;
	wire g730, g731, g732, g733, g734, g736, g737, g738, g741, g739, g740, g744, g745, g742, g743, g746, g748, g749, g750, g753, g751;
	wire g752, g755, g756, g754, g757, g759, g760, g761, g762, g763, g764, g766, g767, g768, g770, g769, g772, g771, g773, g775, g776;
	wire g777, g780, g778, g779, g783, g784, g781, g782, g785, g786, g788, g789, g790, g793, g791, g792, g796, g797, g794, g795, g798;
	wire g799;

	assign o_0_ = (((sk[0]) & (!g217)));
	assign o_1_ = (((sk[1]) & (!g298)));
	assign o_2_ = (((sk[2]) & (!g364)));
	assign o_3_ = (((sk[3]) & (!g431)));
	assign o_4_ = (((sk[4]) & (!g486)));
	assign o_5_ = (((sk[5]) & (!g542)));
	assign o_6_ = (((sk[6]) & (!g585)));
	assign o_7_ = (((sk[7]) & (!g627)));
	assign o_8_ = (((sk[8]) & (!g662)));
	assign o_9_ = (((sk[9]) & (!g689)));
	assign g1 = (((!sk[10]) & (!i_2_) & (!i_0_) & (i_1_)) + ((sk[10]) & (i_2_) & (!i_0_) & (!i_1_)) + ((sk[10]) & (!i_2_) & (i_0_) & (!i_1_)) + ((!sk[10]) & (i_2_) & (i_0_) & (!i_1_)));
	assign g2 = (((i_9_) & (!sk[11]) & (g1)) + ((!i_9_) & (sk[11]) & (!g1)));
	assign g3 = (((!i_8_) & (!sk[12]) & (!i_6_) & (i_7_)) + ((!i_8_) & (sk[12]) & (!i_6_) & (!i_7_)) + ((i_8_) & (!sk[12]) & (i_6_) & (!i_7_)));
	assign g4 = (((i_5_) & (!sk[13]) & (i_3_) & (!i_4_)) + ((!i_5_) & (!sk[13]) & (!i_3_) & (i_4_)) + ((!i_5_) & (sk[13]) & (!i_3_) & (!i_4_)) + ((!i_5_) & (!sk[13]) & (!i_3_) & (i_4_)));
	assign g5 = (((g3) & (!sk[14]) & (g4)) + ((!g3) & (sk[14]) & (!g4)));
	assign g6 = (((!sk[15]) & (!i_2_) & (!i_0_) & (i_1_)) + ((sk[15]) & (!i_2_) & (!i_0_) & (!i_1_)) + ((!sk[15]) & (i_2_) & (i_0_) & (!i_1_)));
	assign g7 = (((!sk[16]) & (!i_5_) & (!i_3_) & (i_4_)) + ((!sk[16]) & (i_5_) & (i_3_) & (!i_4_)) + ((sk[16]) & (!i_5_) & (i_3_) & (!i_4_)));
	assign g8 = (((!sk[17]) & (!i_8_) & (!i_6_) & (i_7_)) + ((!sk[17]) & (i_8_) & (i_6_) & (!i_7_)) + ((sk[17]) & (!i_8_) & (i_6_) & (!i_7_)));
	assign g9 = (((g7) & (!sk[18]) & (g8)));
	assign g10 = (((!i_5_) & (!i_3_) & (!sk[19]) & (i_4_)) + ((i_5_) & (i_3_) & (!sk[19]) & (!i_4_)) + ((i_5_) & (!i_3_) & (sk[19]) & (!i_4_)) + ((!i_5_) & (i_3_) & (sk[19]) & (!i_4_)));
	assign g11 = (((!sk[20]) & (!i_2_) & (!i_0_) & (i_1_)) + ((!sk[20]) & (i_2_) & (i_0_) & (!i_1_)) + ((!sk[20]) & (i_2_) & (!i_0_) & (i_1_)));
	assign g12 = (((!sk[21]) & (g10) & (g11)) + ((sk[21]) & (!g10) & (!g11)));
	assign g13 = (((i_2_) & (i_0_) & (!sk[22]) & (!i_1_) & (!i_9_)) + ((!i_2_) & (!i_0_) & (sk[22]) & (!i_1_) & (!i_9_)) + ((!i_2_) & (!i_0_) & (sk[22]) & (!i_1_) & (!i_9_)) + ((i_2_) & (!i_0_) & (!sk[22]) & (!i_1_) & (i_9_)) + ((!i_2_) & (!i_0_) & (sk[22]) & (!i_1_) & (i_9_)));
	assign g14 = (((sk[23]) & (!i_5_) & (!i_3_) & (!i_4_)) + ((sk[23]) & (!i_5_) & (!i_3_) & (!i_4_)) + ((!sk[23]) & (!i_5_) & (!i_3_) & (i_4_)) + ((!sk[23]) & (i_5_) & (i_3_) & (!i_4_)));
	assign g15 = (((!sk[24]) & (g3) & (g14)) + ((sk[24]) & (!g3) & (!g14)));
	assign g16 = (((!i_8_) & (!i_6_) & (!sk[25]) & (i_7_)) + ((i_8_) & (i_6_) & (!sk[25]) & (!i_7_)) + ((!i_8_) & (!i_6_) & (!sk[25]) & (i_7_)));
	assign g17 = (((g16) & (!sk[26]) & (g4)) + ((g16) & (sk[26]) & (!g4)));
	assign g18 = (((!i_8_) & (!sk[27]) & (!i_6_) & (i_7_)) + ((i_8_) & (!sk[27]) & (i_6_) & (!i_7_)) + ((!i_8_) & (sk[27]) & (!i_6_) & (!i_7_)));
	assign g19 = (((!sk[28]) & (g7) & (g18)));
	assign g20 = (((i_9_) & (i_8_) & (!i_6_) & (!sk[29]) & (!i_7_)) + ((i_9_) & (!i_8_) & (!i_6_) & (!sk[29]) & (i_7_)) + ((i_9_) & (i_8_) & (!i_6_) & (!sk[29]) & (i_7_)));
	assign g21 = (((!i_2_) & (!i_0_) & (sk[30]) & (!i_1_) & (!i_9_)) + ((!i_2_) & (!i_0_) & (sk[30]) & (!i_1_) & (!i_9_)) + ((i_2_) & (!i_0_) & (!sk[30]) & (!i_1_) & (i_9_)) + ((i_2_) & (i_0_) & (!sk[30]) & (!i_1_) & (!i_9_)) + ((i_2_) & (i_0_) & (!sk[30]) & (i_1_) & (!i_9_)));
	assign g22 = (((!i_2_) & (!sk[31]) & (!i_0_) & (i_1_)) + ((i_2_) & (!sk[31]) & (i_0_) & (!i_1_)) + ((i_2_) & (!sk[31]) & (i_0_) & (i_1_)));
	assign g23 = (((g22) & (!sk[32]) & (g14)) + ((g22) & (sk[32]) & (!g14)));
	assign g24 = (((!sk[33]) & (g20) & (!g21) & (!g19) & (g23)) + ((!sk[33]) & (g20) & (g21) & (!g19) & (!g23)) + ((sk[33]) & (!g20) & (!g21) & (g19) & (!g23)));
	assign g25 = (((!sk[34]) & (!i_2_) & (!i_0_) & (i_1_)) + ((!sk[34]) & (i_2_) & (i_0_) & (!i_1_)));
	assign g26 = (((g25) & (!sk[35]) & (g14)) + ((g25) & (sk[35]) & (!g14)));
	assign g27 = (((!sk[36]) & (i_9_) & (i_8_) & (!i_6_) & (!i_7_)) + ((!sk[36]) & (i_9_) & (!i_8_) & (!i_6_) & (i_7_)) + ((!sk[36]) & (i_9_) & (i_8_) & (i_6_) & (!i_7_)));
	assign g28 = (((i_5_) & (i_3_) & (!sk[37]) & (!i_4_)) + ((!i_5_) & (!i_3_) & (!sk[37]) & (i_4_)) + ((!i_5_) & (!i_3_) & (sk[37]) & (!i_4_)) + ((i_5_) & (!i_3_) & (!sk[37]) & (i_4_)) + ((!i_5_) & (i_3_) & (!sk[37]) & (i_4_)));
	assign g29 = (((g28) & (!sk[38]) & (g6)) + ((!g28) & (sk[38]) & (!g6)));
	assign g30 = (((!i_5_) & (!sk[39]) & (!i_3_) & (i_4_)) + ((i_5_) & (!sk[39]) & (i_3_) & (!i_4_)) + ((i_5_) & (sk[39]) & (!i_3_) & (!i_4_)));
	assign g31 = (((g16) & (!sk[40]) & (g30)));
	assign g32 = (((g8) & (!sk[41]) & (g10)) + ((g8) & (sk[41]) & (!g10)));
	assign g33 = (((i_2_) & (!i_0_) & (i_1_) & (!i_9_) & (g31) & (!g32)) + ((!i_2_) & (i_0_) & (!i_1_) & (!i_9_) & (!g31) & (g32)));
	assign g34 = (((g20) & (!g26) & (!sk[43]) & (!g27) & (!g29) & (!g33)) + ((!g20) & (g26) & (!sk[43]) & (g27) & (!g29) & (!g33)) + ((!g20) & (!g26) & (!sk[43]) & (!g27) & (g29) & (g33)) + ((!g20) & (!g26) & (sk[43]) & (!g27) & (!g29) & (!g33)) + ((!g20) & (!g26) & (sk[43]) & (!g27) & (!g29) & (!g33)) + ((!g20) & (!g26) & (sk[43]) & (!g27) & (!g29) & (!g33)) + ((!g20) & (!g26) & (sk[43]) & (!g27) & (!g29) & (!g33)));
	assign g35 = (((i_2_) & (i_0_) & (!sk[44]) & (!i_1_) & (!i_9_)) + ((i_2_) & (!i_0_) & (!sk[44]) & (!i_1_) & (i_9_)) + ((!i_2_) & (!i_0_) & (sk[44]) & (i_1_) & (!i_9_)));
	assign g36 = (((!sk[45]) & (!i_5_) & (!i_3_) & (i_4_)) + ((!sk[45]) & (i_5_) & (i_3_) & (!i_4_)) + ((!sk[45]) & (i_5_) & (!i_3_) & (i_4_)));
	assign g37 = (((!g36) & (sk[46]) & (!g16)) + ((!g36) & (sk[46]) & (!g16)) + ((g36) & (!sk[46]) & (g16)));
	assign g38 = (((i_9_) & (i_8_) & (!sk[47]) & (!i_6_) & (!i_7_)) + ((!i_9_) & (!i_8_) & (sk[47]) & (!i_6_) & (!i_7_)) + ((!i_9_) & (!i_8_) & (sk[47]) & (!i_6_) & (!i_7_)) + ((i_9_) & (!i_8_) & (!sk[47]) & (!i_6_) & (i_7_)));
	assign g39 = (((!i_2_) & (!sk[48]) & (!i_0_) & (i_1_)) + ((i_2_) & (!sk[48]) & (i_0_) & (!i_1_)) + ((!i_2_) & (!sk[48]) & (!i_0_) & (i_1_)));
	assign g40 = (((!sk[49]) & (i_9_) & (i_8_) & (!i_6_) & (!i_7_)) + ((!sk[49]) & (i_9_) & (!i_8_) & (!i_6_) & (i_7_)) + ((sk[49]) & (i_9_) & (!i_8_) & (!i_6_) & (!i_7_)));
	assign g41 = (((g38) & (!sk[50]) & (!g39) & (!g25) & (!g10) & (!g40)) + ((!g38) & (!sk[50]) & (g39) & (g25) & (!g10) & (!g40)) + ((!g38) & (!sk[50]) & (!g39) & (!g25) & (g10) & (g40)) + ((!g38) & (sk[50]) & (!g39) & (g25) & (!g10) & (!g40)) + ((!g38) & (sk[50]) & (g39) & (!g25) & (!g10) & (g40)));
	assign g42 = (((i_2_) & (i_0_) & (!sk[51]) & (!i_1_) & (!i_9_)) + ((i_2_) & (!i_0_) & (!sk[51]) & (!i_1_) & (i_9_)) + ((i_2_) & (!i_0_) & (sk[51]) & (!i_1_) & (!i_9_)));
	assign g43 = (((!sk[52]) & (i_9_) & (g11)) + ((sk[52]) & (!i_9_) & (!g11)));
	assign g44 = (((!sk[53]) & (g28) & (g3)) + ((sk[53]) & (!g28) & (!g3)));
	assign g45 = (((!i_8_) & (!i_6_) & (!sk[54]) & (i_7_)) + ((!i_8_) & (!i_6_) & (sk[54]) & (!i_7_)) + ((!i_8_) & (!i_6_) & (sk[54]) & (!i_7_)) + ((i_8_) & (i_6_) & (!sk[54]) & (!i_7_)));
	assign g46 = (((g28) & (!sk[55]) & (g45)) + ((!g28) & (sk[55]) & (!g45)));
	assign g47 = (((g42) & (!g43) & (!g44) & (!sk[56]) & (g46)) + ((!g42) & (!g43) & (g44) & (sk[56]) & (!g46)) + ((g42) & (g43) & (!g44) & (!sk[56]) & (!g46)));
	assign g48 = (((g20) & (!g28) & (!sk[57]) & (!g1) & (g47)) + ((!g20) & (!g28) & (sk[57]) & (!g1) & (!g47)) + ((!g20) & (!g28) & (sk[57]) & (g1) & (!g47)) + ((g20) & (g28) & (!sk[57]) & (!g1) & (!g47)));
	assign g49 = (((i_2_) & (i_0_) & (!i_1_) & (!sk[58]) & (!i_9_)) + ((i_2_) & (!i_0_) & (!i_1_) & (!sk[58]) & (i_9_)) + ((i_2_) & (i_0_) & (i_1_) & (!sk[58]) & (!i_9_)));
	assign g50 = (((i_8_) & (i_6_) & (!sk[59]) & (!i_7_)) + ((!i_8_) & (!i_6_) & (!sk[59]) & (i_7_)) + ((!i_8_) & (!i_6_) & (sk[59]) & (!i_7_)) + ((!i_8_) & (!i_6_) & (!sk[59]) & (i_7_)));
	assign g51 = (((!sk[60]) & (g50) & (g14)) + ((sk[60]) & (!g50) & (!g14)));
	assign g52 = (((!sk[61]) & (g39) & (g14)) + ((sk[61]) & (g39) & (!g14)));
	assign g53 = (((i_9_) & (!sk[62]) & (g50)) + ((i_9_) & (sk[62]) & (!g50)));
	assign g54 = (((!sk[63]) & (i_8_) & (i_6_) & (!i_7_)) + ((!sk[63]) & (!i_8_) & (!i_6_) & (i_7_)) + ((sk[63]) & (!i_8_) & (!i_6_) & (!i_7_)) + ((!sk[63]) & (!i_8_) & (!i_6_) & (i_7_)));
	assign g55 = (((!sk[64]) & (g54) & (g30)) + ((sk[64]) & (!g54) & (g30)));
	assign g56 = (((g49) & (!sk[65]) & (!g52) & (!g53) & (g55)) + ((g49) & (!sk[65]) & (g52) & (!g53) & (!g55)) + ((!g49) & (sk[65]) & (g52) & (g53) & (!g55)));
	assign g57 = (((g6) & (!sk[66]) & (g4)) + ((!g6) & (sk[66]) & (!g4)));
	assign g58 = (((sk[67]) & (!i_9_) & (!i_8_) & (!i_6_) & (!i_7_)) + ((sk[67]) & (!i_9_) & (!i_8_) & (!i_6_) & (!i_7_)) + ((!sk[67]) & (i_9_) & (i_8_) & (!i_6_) & (!i_7_)) + ((!sk[67]) & (i_9_) & (!i_8_) & (!i_6_) & (i_7_)) + ((!sk[67]) & (i_9_) & (i_8_) & (!i_6_) & (!i_7_)));
	assign g59 = (((!i_2_) & (!sk[68]) & (!i_0_) & (i_1_)) + ((i_2_) & (!sk[68]) & (i_0_) & (!i_1_)) + ((!i_2_) & (!sk[68]) & (i_0_) & (i_1_)));
	assign g60 = (((!sk[69]) & (g7) & (g59)));
	assign g61 = (((!sk[70]) & (g39) & (!g30) & (!g57) & (!g58) & (!g60)) + ((!sk[70]) & (!g39) & (g30) & (g57) & (!g58) & (!g60)) + ((!sk[70]) & (g39) & (g30) & (!g57) & (!g58) & (!g60)) + ((sk[70]) & (!g39) & (!g30) & (g57) & (!g58) & (!g60)) + ((!sk[70]) & (!g39) & (!g30) & (!g57) & (g58) & (g60)) + ((sk[70]) & (!g39) & (!g30) & (!g57) & (!g58) & (g60)));
	assign g62 = (((!sk[71]) & (g59) & (g4)) + ((sk[71]) & (g59) & (!g4)));
	assign g63 = (((!sk[72]) & (!i_2_) & (!i_0_) & (i_1_)) + ((!sk[72]) & (i_2_) & (i_0_) & (!i_1_)) + ((sk[72]) & (!i_2_) & (i_0_) & (!i_1_)));
	assign g64 = (((g63) & (!sk[73]) & (g14)) + ((g63) & (sk[73]) & (!g14)));
	assign g65 = (((!sk[74]) & (g62) & (g53) & (!g64)) + ((!sk[74]) & (!g62) & (!g53) & (g64)) + ((!sk[74]) & (!g62) & (g53) & (g64)));
	assign g66 = (((g49) & (!g51) & (!g56) & (!g61) & (!sk[75]) & (!g65)) + ((!g49) & (g51) & (g56) & (!g61) & (!sk[75]) & (!g65)) + ((!g49) & (!g51) & (!g56) & (g61) & (!sk[75]) & (g65)) + ((!g49) & (!g51) & (!g56) & (!g61) & (sk[75]) & (!g65)) + ((!g49) & (!g51) & (!g56) & (!g61) & (sk[75]) & (!g65)));
	assign g67 = (((g35) & (!g37) & (!sk[76]) & (!g41) & (!g48) & (!g66)) + ((!g35) & (g37) & (!sk[76]) & (g41) & (!g48) & (!g66)) + ((!g35) & (!g37) & (!sk[76]) & (!g41) & (g48) & (g66)) + ((!g35) & (!g37) & (!sk[76]) & (!g41) & (g48) & (g66)) + ((!g35) & (g37) & (!sk[76]) & (!g41) & (g48) & (g66)));
	assign g68 = (((!i_6_) & (sk[77]) & (i_7_)) + ((i_6_) & (!sk[77]) & (i_7_)));
	assign g69 = (((!sk[78]) & (i_9_) & (g68)));
	assign g70 = (((g22) & (!g36) & (!g20) & (!sk[79]) & (!g58) & (!g12)) + ((g22) & (g36) & (g20) & (!sk[79]) & (!g58) & (!g12)) + ((!g22) & (g36) & (g20) & (!sk[79]) & (!g58) & (!g12)) + ((!g22) & (!g36) & (!g20) & (!sk[79]) & (g58) & (g12)) + ((!g22) & (!g36) & (!g20) & (sk[79]) & (!g58) & (!g12)));
	assign g71 = (((!sk[80]) & (g6) & (g14)) + ((sk[80]) & (!g6) & (!g14)));
	assign g72 = (((!sk[81]) & (i_8_) & (g28) & (!g59) & (!g71)) + ((!sk[81]) & (i_8_) & (!g28) & (!g59) & (g71)) + ((sk[81]) & (!i_8_) & (!g28) & (!g59) & (g71)) + ((sk[81]) & (i_8_) & (!g28) & (g59) & (!g71)));
	assign g73 = (((!sk[82]) & (i_9_) & (i_8_) & (!i_6_) & (!i_7_)) + ((!sk[82]) & (i_9_) & (!i_8_) & (!i_6_) & (i_7_)) + ((!sk[82]) & (i_9_) & (i_8_) & (!i_6_) & (!i_7_)));
	assign g74 = (((g4) & (sk[83]) & (!g1)) + ((g4) & (!sk[83]) & (g1)) + ((!g4) & (sk[83]) & (g1)));
	assign g75 = (((!sk[84]) & (i_0_) & (i_1_)) + ((sk[84]) & (i_0_) & (!i_1_)));
	assign g76 = (((!sk[85]) & (!i_5_) & (!i_3_) & (i_4_)) + ((sk[85]) & (!i_5_) & (!i_3_) & (!i_4_)) + ((sk[85]) & (!i_5_) & (!i_3_) & (!i_4_)) + ((!sk[85]) & (i_5_) & (i_3_) & (!i_4_)));
	assign g77 = (((!sk[86]) & (g76) & (g45)) + ((sk[86]) & (!g76) & (!g45)));
	assign g78 = (((!sk[87]) & (i_0_) & (i_1_)));
	assign g79 = (((!i_2_) & (!g78) & (!sk[88]) & (i_9_)) + ((!i_2_) & (!g78) & (sk[88]) & (!i_9_)) + ((i_2_) & (g78) & (!sk[88]) & (!i_9_)));
	assign g80 = (((i_2_) & (g7) & (!g75) & (g16) & (!g77) & (g79)) + ((!i_2_) & (!g7) & (g75) & (!g16) & (g77) & (g79)));
	assign g81 = (((i_6_) & (!sk[90]) & (i_7_)) + ((i_6_) & (sk[90]) & (!i_7_)));
	assign g82 = (((!sk[91]) & (g63) & (g4)) + ((sk[91]) & (g63) & (!g4)));
	assign g83 = (((!sk[92]) & (i_6_) & (i_7_)));
	assign g84 = (((!sk[93]) & (g76) & (g63)) + ((sk[93]) & (!g76) & (g63)));
	assign g85 = (((!sk[94]) & (g54) & (g14)) + ((sk[94]) & (!g54) & (!g14)));
	assign g86 = (((!sk[95]) & (g35) & (!g20) & (!g84) & (g85)) + ((!sk[95]) & (g35) & (g20) & (!g84) & (!g85)) + ((sk[95]) & (!g35) & (g20) & (g84) & (!g85)));
	assign g87 = (((g73) & (!sk[96]) & (!g74) & (!g80) & (!g765) & (!g86)) + ((!g73) & (!sk[96]) & (g74) & (g80) & (!g765) & (!g86)) + ((!g73) & (!sk[96]) & (!g74) & (!g80) & (g765) & (g86)) + ((!g73) & (sk[96]) & (!g74) & (!g80) & (g765) & (!g86)) + ((!g73) & (sk[96]) & (g74) & (!g80) & (g765) & (!g86)));
	assign g88 = (((!sk[97]) & (g69) & (g70) & (!g72) & (!g87)) + ((!sk[97]) & (g69) & (!g70) & (!g72) & (g87)) + ((sk[97]) & (!g69) & (!g70) & (!g72) & (g87)) + ((!sk[97]) & (g69) & (!g70) & (!g72) & (g87)));
	assign g89 = (((g787) & (g774) & (!g24) & (g34) & (g67) & (g88)));
	assign g90 = (((g36) & (!sk[99]) & (g63)));
	assign g91 = (((g22) & (!sk[100]) & (!g28) & (!g73) & (!g27) & (!g90)) + ((!g22) & (!sk[100]) & (!g28) & (!g73) & (g27) & (g90)) + ((!g22) & (!sk[100]) & (g28) & (g73) & (!g27) & (!g90)) + ((g22) & (!sk[100]) & (!g28) & (g73) & (!g27) & (!g90)));
	assign g92 = (((!sk[101]) & (i_3_) & (i_4_)));
	assign g93 = (((g22) & (!i_9_) & (!g50) & (!i_5_) & (g92) & (!g18)) + ((g22) & (i_9_) & (!g50) & (i_5_) & (g92) & (g18)));
	assign g94 = (((g39) & (!sk[103]) & (g4)) + ((g39) & (sk[103]) & (!g4)));
	assign g95 = (((i_6_) & (i_7_) & (!sk[104]) & (!g6) & (!g10)) + ((i_6_) & (!i_7_) & (sk[104]) & (!g6) & (!g10)) + ((!i_6_) & (i_7_) & (sk[104]) & (!g6) & (!g10)) + ((!i_6_) & (!i_7_) & (sk[104]) & (g6) & (!g10)) + ((i_6_) & (!i_7_) & (!sk[104]) & (!g6) & (g10)) + ((!i_6_) & (!i_7_) & (sk[104]) & (!g6) & (g10)));
	assign g96 = (((i_9_) & (!sk[105]) & (!i_8_) & (!g83) & (!g94) & (!g95)) + ((!i_9_) & (!sk[105]) & (i_8_) & (g83) & (!g94) & (!g95)) + ((!i_9_) & (!sk[105]) & (!i_8_) & (!g83) & (g94) & (g95)) + ((i_9_) & (!sk[105]) & (i_8_) & (!g83) & (!g94) & (!g95)) + ((i_9_) & (!sk[105]) & (!i_8_) & (g83) & (g94) & (!g95)));
	assign g97 = (((!sk[106]) & (g50) & (g10)) + ((sk[106]) & (!g50) & (!g10)));
	assign g98 = (((g42) & (!g13) & (g85) & (sk[107]) & (!g97)) + ((g42) & (g13) & (!g85) & (!sk[107]) & (!g97)) + ((!g42) & (!g13) & (!g85) & (sk[107]) & (g97)) + ((g42) & (!g13) & (!g85) & (!sk[107]) & (g97)));
	assign g99 = (((!sk[108]) & (g63) & (g30)));
	assign g100 = (((g99) & (!sk[109]) & (g40) & (!g12)) + ((!g99) & (!sk[109]) & (!g40) & (g12)) + ((!g99) & (sk[109]) & (g40) & (!g12)));
	assign g101 = (((!g50) & (sk[110]) & (g36)) + ((g50) & (!sk[110]) & (g36)));
	assign g102 = (((!i_2_) & (!i_9_) & (!g7) & (g101) & (g75) & (!g3)) + ((!i_2_) & (i_9_) & (g7) & (!g101) & (g75) & (!g3)));
	assign g103 = (((!sk[112]) & (!g20) & (!g25) & (g4)) + ((!sk[112]) & (g20) & (g25) & (!g4)));
	assign g104 = (((g36) & (!g20) & (!g59) & (!g53) & (!sk[113]) & (!g103)) + ((!g36) & (g20) & (g59) & (!g53) & (!sk[113]) & (!g103)) + ((!g36) & (!g20) & (!g59) & (g53) & (!sk[113]) & (g103)) + ((!g36) & (!g20) & (!g59) & (!g53) & (sk[113]) & (!g103)) + ((!g36) & (!g20) & (!g59) & (!g53) & (sk[113]) & (!g103)) + ((!g36) & (!g20) & (!g59) & (!g53) & (sk[113]) & (!g103)));
	assign g105 = (((g22) & (!sk[114]) & (!g50) & (!g38) & (!g35) & (!g76)) + ((!g22) & (!sk[114]) & (g50) & (g38) & (!g35) & (!g76)) + ((!g22) & (!sk[114]) & (!g50) & (!g38) & (g35) & (g76)) + ((g22) & (!sk[114]) & (!g50) & (!g38) & (!g35) & (!g76)) + ((!g22) & (sk[114]) & (!g50) & (!g38) & (g35) & (!g76)));
	assign g106 = (((!sk[115]) & (g7) & (!g1) & (!g14) & (!g53) & (!g27)) + ((!sk[115]) & (!g7) & (g1) & (g14) & (!g53) & (!g27)) + ((!sk[115]) & (g7) & (!g1) & (!g14) & (g53) & (!g27)) + ((!sk[115]) & (!g7) & (!g1) & (!g14) & (g53) & (g27)) + ((sk[115]) & (!g7) & (!g1) & (!g14) & (!g53) & (g27)));
	assign g107 = (((g100) & (!sk[116]) & (!g102) & (!g104) & (!g105) & (!g106)) + ((!g100) & (!sk[116]) & (g102) & (g104) & (!g105) & (!g106)) + ((!g100) & (!sk[116]) & (!g102) & (!g104) & (g105) & (g106)) + ((!g100) & (sk[116]) & (!g102) & (g104) & (!g105) & (!g106)));
	assign g108 = (((g91) & (!sk[117]) & (!g93) & (!g96) & (!g98) & (!g107)) + ((!g91) & (!sk[117]) & (g93) & (g96) & (!g98) & (!g107)) + ((!g91) & (!sk[117]) & (!g93) & (!g96) & (g98) & (g107)) + ((!g91) & (sk[117]) & (!g93) & (!g96) & (!g98) & (g107)));
	assign g109 = (((!i_9_) & (sk[118]) & (g3) & (!g63) & (!g30)) + ((i_9_) & (!sk[118]) & (g3) & (!g63) & (!g30)) + ((!i_9_) & (sk[118]) & (!g3) & (!g63) & (!g30)) + ((i_9_) & (!sk[118]) & (!g3) & (!g63) & (g30)) + ((!i_9_) & (sk[118]) & (!g3) & (!g63) & (!g30)));
	assign g110 = (((!sk[119]) & (i_9_) & (g7) & (!g39) & (!g16)) + ((!sk[119]) & (i_9_) & (g7) & (!g39) & (!g16)) + ((!sk[119]) & (i_9_) & (!g7) & (!g39) & (g16)) + ((sk[119]) & (i_9_) & (!g7) & (!g39) & (!g16)));
	assign g111 = (((!sk[120]) & (i_9_) & (!i_8_) & (!g81) & (!g84) & (!g62)) + ((!sk[120]) & (!i_9_) & (i_8_) & (g81) & (!g84) & (!g62)) + ((!sk[120]) & (!i_9_) & (!i_8_) & (!g81) & (g84) & (g62)) + ((!sk[120]) & (i_9_) & (i_8_) & (g81) & (!g84) & (g62)) + ((sk[120]) & (!i_9_) & (!i_8_) & (g81) & (g84) & (!g62)));
	assign g112 = (((!sk[121]) & (g36) & (g1)) + ((sk[121]) & (g36) & (!g1)));
	assign g113 = (((g20) & (!g73) & (!g30) & (!g11) & (!sk[122]) & (!g112)) + ((g20) & (!g73) & (g30) & (g11) & (!sk[122]) & (!g112)) + ((!g20) & (g73) & (g30) & (!g11) & (!sk[122]) & (!g112)) + ((!g20) & (g73) & (!g30) & (!g11) & (sk[122]) & (g112)) + ((!g20) & (!g73) & (!g30) & (g11) & (!sk[122]) & (g112)));
	assign g114 = (((!sk[123]) & (g109) & (g110) & (!g111) & (!g113)) + ((!sk[123]) & (g109) & (!g110) & (!g111) & (g113)) + ((sk[123]) & (g109) & (!g110) & (!g111) & (!g113)) + ((sk[123]) & (!g109) & (g110) & (!g111) & (!g113)));
	assign g115 = (((!sk[124]) & (g38) & (g57) & (!g53) & (!g90)) + ((sk[124]) & (!g38) & (g57) & (g53) & (!g90)) + ((!sk[124]) & (g38) & (!g57) & (!g53) & (g90)) + ((sk[124]) & (!g38) & (!g57) & (!g53) & (g90)));
	assign g116 = (((!sk[125]) & (g76) & (g16)) + ((sk[125]) & (!g76) & (g16)));
	assign g117 = (((!sk[126]) & (g10) & (g45)) + ((sk[126]) & (!g10) & (!g45)));
	assign g118 = (((g20) & (!g13) & (g57) & (sk[127]) & (!g117)) + ((g20) & (g13) & (!g57) & (!sk[127]) & (!g117)) + ((!g20) & (!g13) & (!g57) & (sk[127]) & (g117)) + ((g20) & (!g13) & (!g57) & (!sk[127]) & (g117)));
	assign g119 = (((i_0_) & (sk[0]) & (!i_1_)) + ((i_0_) & (!sk[0]) & (i_1_)) + ((!i_0_) & (sk[0]) & (i_1_)));
	assign g120 = (((g54) & (!sk[1]) & (g76)) + ((!g54) & (sk[1]) & (!g76)));
	assign g121 = (((i_2_) & (!i_9_) & (!g119) & (!g120) & (!sk[2]) & (!g9)) + ((!i_2_) & (i_9_) & (g119) & (!g120) & (!sk[2]) & (!g9)) + ((!i_2_) & (!i_9_) & (!g119) & (g120) & (!sk[2]) & (g9)) + ((i_2_) & (!i_9_) & (!g119) & (g120) & (!sk[2]) & (!g9)) + ((!i_2_) & (i_9_) & (!g119) & (!g120) & (sk[2]) & (g9)));
	assign g122 = (((g50) & (!sk[3]) & (g28)) + ((!g50) & (sk[3]) & (!g28)));
	assign g123 = (((i_2_) & (!sk[4]) & (!g78) & (!i_9_) & (!g122) & (!g17)) + ((!i_2_) & (!sk[4]) & (g78) & (i_9_) & (!g122) & (!g17)) + ((!i_2_) & (!sk[4]) & (!g78) & (!i_9_) & (g122) & (g17)) + ((i_2_) & (!sk[4]) & (g78) & (i_9_) & (!g122) & (g17)) + ((!i_2_) & (sk[4]) & (g78) & (!i_9_) & (g122) & (!g17)));
	assign g124 = (((g39) & (!sk[5]) & (g76)) + ((g39) & (sk[5]) & (!g76)));
	assign g125 = (((!g50) & (sk[6]) & (g30)) + ((g50) & (!sk[6]) & (g30)));
	assign g126 = (((!g101) & (!g35) & (!g20) & (!g124) & (!g125) & (!g13)) + ((!g101) & (!g35) & (!g20) & (!g124) & (!g125) & (!g13)) + ((!g101) & (!g35) & (!g20) & (!g124) & (!g125) & (!g13)) + ((!g101) & (!g35) & (!g20) & (!g124) & (!g125) & (!g13)) + ((!g101) & (!g35) & (!g20) & (!g124) & (!g125) & (g13)) + ((!g101) & (!g35) & (!g20) & (!g124) & (!g125) & (g13)) + ((!g101) & (!g35) & (!g20) & (!g124) & (!g125) & (g13)) + ((!g101) & (!g35) & (!g20) & (!g124) & (!g125) & (g13)));
	assign g127 = (((g20) & (!g28) & (!sk[8]) & (!g25) & (g99)) + ((g20) & (g28) & (!sk[8]) & (!g25) & (!g99)) + ((g20) & (!g28) & (sk[8]) & (g25) & (!g99)));
	assign g128 = (((g73) & (!g84) & (!g123) & (!sk[9]) & (!g126) & (!g127)) + ((!g73) & (g84) & (g123) & (!sk[9]) & (!g126) & (!g127)) + ((!g73) & (!g84) & (!g123) & (!sk[9]) & (g126) & (g127)) + ((!g73) & (!g84) & (!g123) & (sk[9]) & (g126) & (!g127)) + ((!g73) & (!g84) & (!g123) & (sk[9]) & (g126) & (!g127)));
	assign g129 = (((!sk[10]) & (g42) & (!g116) & (!g118) & (!g121) & (!g128)) + ((!sk[10]) & (!g42) & (g116) & (g118) & (!g121) & (!g128)) + ((!sk[10]) & (!g42) & (!g116) & (!g118) & (g121) & (g128)) + ((sk[10]) & (!g42) & (!g116) & (!g118) & (!g121) & (g128)) + ((!sk[10]) & (g42) & (!g116) & (!g118) & (!g121) & (g128)));
	assign g130 = (((i_9_) & (i_8_) & (g81) & (!g36) & (g57) & (!g11)) + ((!i_9_) & (!i_8_) & (g81) & (g36) & (!g57) & (g11)));
	assign g131 = (((!sk[12]) & (!i_2_) & (!i_0_) & (i_9_)) + ((!sk[12]) & (i_2_) & (i_0_) & (!i_9_)) + ((sk[12]) & (!i_2_) & (!i_0_) & (!i_9_)));
	assign g132 = (((!g50) & (g35) & (!g10) & (!g2) & (!g14) & (g131)) + ((!g50) & (!g35) & (!g10) & (!g2) & (!g14) & (g131)) + ((!g50) & (!g35) & (!g10) & (g2) & (!g14) & (g131)));
	assign g133 = (((i_9_) & (!sk[14]) & (g63)) + ((!i_9_) & (sk[14]) & (!g63)));
	assign g134 = (((g8) & (!sk[15]) & (g28)) + ((g8) & (sk[15]) & (!g28)));
	assign g135 = (((g8) & (!sk[16]) & (g14)) + ((g8) & (sk[16]) & (!g14)));
	assign g136 = (((!g49) & (g13) & (g133) & (!g134) & (!g32) & (!g135)) + ((!g49) & (g13) & (g133) & (!g134) & (!g32) & (!g135)) + ((!g49) & (!g13) & (g133) & (!g134) & (!g32) & (!g135)) + ((!g49) & (!g13) & (g133) & (!g134) & (!g32) & (!g135)) + ((!g49) & (g13) & (!g133) & (!g134) & (!g32) & (!g135)) + ((!g49) & (g13) & (!g133) & (!g134) & (!g32) & (!g135)) + ((!g49) & (!g13) & (!g133) & (!g134) & (!g32) & (!g135)) + ((!g49) & (!g13) & (!g133) & (!g134) & (!g32) & (!g135)));
	assign g137 = (((i_9_) & (!sk[18]) & (g16)));
	assign g138 = (((!sk[19]) & (!i_8_) & (!i_6_) & (i_7_)) + ((!sk[19]) & (i_8_) & (i_6_) & (!i_7_)) + ((!sk[19]) & (i_8_) & (i_6_) & (i_7_)));
	assign g139 = (((!sk[20]) & (g138) & (g14)) + ((sk[20]) & (g138) & (!g14)));
	assign g140 = (((g7) & (!g43) & (!sk[21]) & (!g137) & (!g1) & (!g139)) + ((!g7) & (g43) & (!sk[21]) & (g137) & (!g1) & (!g139)) + ((g7) & (!g43) & (!sk[21]) & (g137) & (!g1) & (!g139)) + ((!g7) & (!g43) & (sk[21]) & (!g137) & (!g1) & (g139)) + ((!g7) & (!g43) & (!sk[21]) & (!g137) & (g1) & (g139)));
	assign g141 = (((!sk[22]) & (g76) & (g138)) + ((sk[22]) & (!g76) & (g138)));
	assign g142 = (((sk[23]) & (!g36) & (!g25)) + ((sk[23]) & (!g36) & (!g25)) + ((!sk[23]) & (g36) & (g25)));
	assign g143 = (((g76) & (!sk[24]) & (g11) & (!g40) & (!g142)) + ((g76) & (!sk[24]) & (!g11) & (!g40) & (g142)) + ((!g76) & (sk[24]) & (!g11) & (g40) & (!g142)) + ((!g76) & (sk[24]) & (g11) & (g40) & (!g142)));
	assign g144 = (((!sk[25]) & (g25) & (g30)));
	assign g145 = (((g38) & (!g42) & (!g77) & (!g27) & (!g29) & (!g144)) + ((g38) & (!g42) & (!g77) & (!g27) & (!g29) & (!g144)) + ((g38) & (!g42) & (!g77) & (!g27) & (!g29) & (!g144)) + ((g38) & (!g42) & (!g77) & (!g27) & (!g29) & (!g144)) + ((!g38) & (!g42) & (!g77) & (!g27) & (!g29) & (!g144)) + ((!g38) & (!g42) & (!g77) & (!g27) & (!g29) & (!g144)));
	assign g146 = (((g21) & (!g15) & (!g141) & (!g143) & (!sk[27]) & (!g145)) + ((!g21) & (g15) & (g141) & (!g143) & (!sk[27]) & (!g145)) + ((g21) & (!g15) & (!g141) & (!g143) & (!sk[27]) & (g145)) + ((!g21) & (!g15) & (!g141) & (g143) & (!sk[27]) & (g145)) + ((!g21) & (!g15) & (!g141) & (!g143) & (sk[27]) & (g145)));
	assign g147 = (((g130) & (!g132) & (!g136) & (!g140) & (!sk[28]) & (!g146)) + ((!g130) & (g132) & (g136) & (!g140) & (!sk[28]) & (!g146)) + ((!g130) & (!g132) & (!g136) & (g140) & (!sk[28]) & (g146)) + ((!g130) & (!g132) & (g136) & (!g140) & (sk[28]) & (g146)));
	assign g148 = (((g54) & (!sk[29]) & (g28)) + ((!g54) & (sk[29]) & (!g28)));
	assign g149 = (((!i_9_) & (!g36) & (!g39) & (!g45) & (!g1) & (g148)) + ((i_9_) & (g36) & (g39) & (!g45) & (!g1) & (!g148)));
	assign g150 = (((g36) & (!g20) & (!g18) & (!g21) & (!sk[31]) & (!g144)) + ((g36) & (!g20) & (g18) & (!g21) & (!sk[31]) & (!g144)) + ((!g36) & (g20) & (g18) & (!g21) & (!sk[31]) & (!g144)) + ((!g36) & (g20) & (!g18) & (!g21) & (sk[31]) & (g144)) + ((!g36) & (!g20) & (!g18) & (g21) & (!sk[31]) & (g144)));
	assign g151 = (((!sk[32]) & (!i_2_) & (!i_9_) & (g75)) + ((!sk[32]) & (!i_2_) & (!i_9_) & (g75)) + ((!sk[32]) & (i_2_) & (i_9_) & (!g75)) + ((sk[32]) & (!i_2_) & (!i_9_) & (!g75)));
	assign g152 = (((!sk[33]) & (!g78) & (!g3) & (g30)) + ((!sk[33]) & (g78) & (g3) & (!g30)) + ((!sk[33]) & (g78) & (!g3) & (g30)));
	assign g153 = (((i_2_) & (!g76) & (!g16) & (!g151) & (!sk[34]) & (!g152)) + ((!i_2_) & (g76) & (g16) & (!g151) & (!sk[34]) & (!g152)) + ((!i_2_) & (!g76) & (!g16) & (g151) & (!sk[34]) & (g152)) + ((i_2_) & (!g76) & (g16) & (g151) & (!sk[34]) & (!g152)));
	assign g154 = (((i_8_) & (i_6_) & (!i_7_) & (g36) & (!g133) & (!g43)) + ((!i_8_) & (!i_6_) & (!i_7_) & (g36) & (!g133) & (!g43)));
	assign g155 = (((!sk[36]) & (g149) & (g150) & (!g153) & (!g154)) + ((!sk[36]) & (g149) & (!g150) & (!g153) & (g154)) + ((sk[36]) & (!g149) & (!g150) & (!g153) & (!g154)));
	assign g156 = (((g54) & (!sk[37]) & (g4)) + ((!g54) & (sk[37]) & (!g4)));
	assign g157 = (((!sk[38]) & (g8) & (g4)) + ((sk[38]) & (g8) & (!g4)));
	assign g158 = (((!sk[39]) & (g8) & (g30)));
	assign g159 = (((g42) & (!sk[40]) & (g156) & (!g157) & (!g158)) + ((g42) & (!sk[40]) & (!g156) & (!g157) & (g158)) + ((g42) & (sk[40]) & (!g156) & (g157) & (!g158)));
	assign g160 = (((i_9_) & (!sk[41]) & (i_8_) & (!i_6_) & (!g36)) + ((i_9_) & (!sk[41]) & (!i_8_) & (!i_6_) & (g36)) + ((i_9_) & (!sk[41]) & (!i_8_) & (!i_6_) & (g36)) + ((!i_9_) & (sk[41]) & (!i_8_) & (i_6_) & (g36)));
	assign g161 = (((!sk[42]) & (g36) & (g54)) + ((sk[42]) & (g36) & (!g54)));
	assign g162 = (((i_9_) & (!sk[43]) & (!g25) & (!g3) & (!g10) & (!g161)) + ((!i_9_) & (!sk[43]) & (g25) & (g3) & (!g10) & (!g161)) + ((!i_9_) & (!sk[43]) & (!g25) & (!g3) & (g10) & (g161)) + ((i_9_) & (!sk[43]) & (g25) & (!g3) & (!g10) & (!g161)) + ((!i_9_) & (sk[43]) & (g25) & (!g3) & (!g10) & (g161)));
	assign g163 = (((i_7_) & (!g6) & (!sk[44]) & (!g160) & (g162)) + ((i_7_) & (!g6) & (sk[44]) & (!g160) & (!g162)) + ((!i_7_) & (g6) & (sk[44]) & (!g160) & (!g162)) + ((!i_7_) & (!g6) & (sk[44]) & (!g160) & (!g162)) + ((i_7_) & (g6) & (!sk[44]) & (!g160) & (!g162)));
	assign g164 = (((g28) & (g25) & (!sk[45]) & (!g84) & (!g53)) + ((g28) & (!g25) & (!sk[45]) & (!g84) & (g53)) + ((!g28) & (!g25) & (sk[45]) & (g84) & (g53)) + ((!g28) & (g25) & (sk[45]) & (!g84) & (g53)));
	assign g165 = (((!sk[46]) & (g18) & (g14)) + ((sk[46]) & (g18) & (!g14)));
	assign g166 = (((!sk[47]) & (g49) & (!g50) & (!g7) & (g165)) + ((!sk[47]) & (g49) & (g50) & (!g7) & (!g165)) + ((sk[47]) & (g49) & (!g50) & (g7) & (!g165)));
	assign g167 = (((!g38) & (g36) & (g39) & (!g28) & (!g137) & (!g40)) + ((!g38) & (!g36) & (g39) & (!g28) & (g137) & (!g40)) + ((!g38) & (g36) & (g39) & (!g28) & (!g137) & (g40)));
	assign g168 = (((g7) & (!sk[49]) & (g45)) + ((g7) & (sk[49]) & (!g45)));
	assign g169 = (((!sk[50]) & (g28) & (g16)) + ((sk[50]) & (!g28) & (g16)));
	assign g170 = (((!sk[51]) & (g7) & (g54)) + ((sk[51]) & (g7) & (!g54)));
	assign g171 = (((!sk[52]) & (g7) & (g138)));
	assign g172 = (((g99) & (!g134) & (!sk[53]) & (!g43) & (!g58) & (!g171)) + ((!g99) & (!g134) & (sk[53]) & (g43) & (!g58) & (!g171)) + ((!g99) & (!g134) & (!sk[53]) & (!g43) & (g58) & (g171)) + ((!g99) & (!g134) & (sk[53]) & (!g43) & (!g58) & (!g171)) + ((!g99) & (g134) & (!sk[53]) & (g43) & (!g58) & (!g171)) + ((!g99) & (!g134) & (sk[53]) & (g43) & (g58) & (!g171)) + ((!g99) & (!g134) & (sk[53]) & (!g43) & (g58) & (!g171)));
	assign g173 = (((g164) & (!sk[54]) & (!g166) & (!g167) & (!g747) & (!g172)) + ((!g164) & (!sk[54]) & (g166) & (g167) & (!g747) & (!g172)) + ((!g164) & (!sk[54]) & (!g166) & (!g167) & (g747) & (g172)) + ((!g164) & (!sk[54]) & (!g166) & (!g167) & (g747) & (g172)));
	assign g174 = (((g2) & (!sk[55]) & (!g46) & (!g159) & (!g163) & (!g173)) + ((!g2) & (!sk[55]) & (g46) & (g159) & (!g163) & (!g173)) + ((!g2) & (!sk[55]) & (!g46) & (!g159) & (g163) & (g173)) + ((!g2) & (!sk[55]) & (!g46) & (!g159) & (g163) & (g173)) + ((!g2) & (!sk[55]) & (!g46) & (!g159) & (g163) & (g173)));
	assign g175 = (((!g38) & (!sk[56]) & (!g6) & (g30)) + ((g38) & (!sk[56]) & (g6) & (!g30)) + ((!g38) & (!sk[56]) & (!g6) & (g30)));
	assign g176 = (((g39) & (g20) & (!g10) & (!sk[57]) & (!g175)) + ((g39) & (!g20) & (!g10) & (!sk[57]) & (g175)) + ((!g39) & (!g20) & (!g10) & (sk[57]) & (!g175)) + ((!g39) & (!g20) & (!g10) & (sk[57]) & (!g175)) + ((g39) & (g20) & (g10) & (!sk[57]) & (!g175)));
	assign g177 = (((g3) & (!sk[58]) & (g10)) + ((!g3) & (sk[58]) & (!g10)));
	assign g178 = (((g22) & (!i_9_) & (!g101) & (!sk[59]) & (!g16) & (!g26)) + ((g22) & (!i_9_) & (g101) & (!sk[59]) & (!g16) & (!g26)) + ((!g22) & (i_9_) & (g101) & (!sk[59]) & (!g16) & (!g26)) + ((!g22) & (i_9_) & (!g101) & (!sk[59]) & (g16) & (g26)) + ((!g22) & (!i_9_) & (!g101) & (!sk[59]) & (g16) & (g26)));
	assign g179 = (((!sk[60]) & (g16) & (g10)) + ((sk[60]) & (g16) & (!g10)));
	assign g180 = (((!sk[61]) & (g36) & (g138)));
	assign g181 = (((g35) & (!sk[62]) & (g179) & (!g21) & (!g180)) + ((g35) & (!sk[62]) & (!g179) & (!g21) & (g180)) + ((!g35) & (sk[62]) & (!g179) & (!g21) & (g180)));
	assign g182 = (((g30) & (!sk[63]) & (g138)));
	assign g183 = (((!g4) & (sk[64]) & (g18)) + ((g4) & (!sk[64]) & (g18)));
	assign g184 = (((g42) & (!g2) & (!g182) & (!g183) & (!sk[65]) & (!g44)) + ((!g42) & (!g2) & (!g182) & (!g183) & (sk[65]) & (!g44)) + ((!g42) & (g2) & (g182) & (!g183) & (!sk[65]) & (!g44)) + ((!g42) & (!g2) & (!g182) & (g183) & (!sk[65]) & (g44)) + ((!g42) & (!g2) & (!g182) & (!g183) & (sk[65]) & (!g44)) + ((!g42) & (!g2) & (!g182) & (!g183) & (sk[65]) & (!g44)) + ((!g42) & (!g2) & (!g182) & (!g183) & (sk[65]) & (!g44)));
	assign g185 = (((!sk[66]) & (g49) & (!g177) & (!g178) & (!g181) & (!g184)) + ((!sk[66]) & (!g49) & (g177) & (g178) & (!g181) & (!g184)) + ((!sk[66]) & (!g49) & (!g177) & (!g178) & (g181) & (g184)) + ((sk[66]) & (!g49) & (!g177) & (!g178) & (!g181) & (g184)) + ((!sk[66]) & (g49) & (!g177) & (!g178) & (!g181) & (g184)));
	assign g186 = (((!sk[67]) & (g45) & (g14)) + ((sk[67]) & (!g45) & (!g14)));
	assign g187 = (((!i_2_) & (i_0_) & (!i_1_) & (!i_9_) & (g179) & (!g186)) + ((i_2_) & (!i_0_) & (i_1_) & (!i_9_) & (!g179) & (g186)));
	assign g188 = (((g7) & (!g36) & (!g35) & (!sk[69]) & (!g42) & (!g16)) + ((!g7) & (g36) & (g35) & (!sk[69]) & (!g42) & (!g16)) + ((g7) & (!g36) & (g35) & (!sk[69]) & (!g42) & (g16)) + ((!g7) & (g36) & (!g35) & (!sk[69]) & (g42) & (g16)) + ((!g7) & (!g36) & (!g35) & (!sk[69]) & (g42) & (g16)));
	assign g189 = (((g38) & (!g11) & (!sk[70]) & (!g14) & (g188)) + ((!g38) & (!g11) & (sk[70]) & (!g14) & (!g188)) + ((!g38) & (!g11) & (sk[70]) & (g14) & (!g188)) + ((g38) & (g11) & (!sk[70]) & (!g14) & (!g188)));
	assign g190 = (((g176) & (g185) & (!g187) & (!sk[71]) & (!g189)) + ((g176) & (!g185) & (!g187) & (!sk[71]) & (g189)) + ((g176) & (g185) & (!g187) & (!sk[71]) & (g189)));
	assign g191 = (((!g115) & (g129) & (g147) & (g155) & (g174) & (g190)));
	assign g192 = (((!i_9_) & (!sk[73]) & (!i_8_) & (i_6_)) + ((i_9_) & (!sk[73]) & (i_8_) & (!i_6_)) + ((i_9_) & (!sk[73]) & (!i_8_) & (i_6_)));
	assign g193 = (((!sk[74]) & (g36) & (g45)) + ((sk[74]) & (g36) & (!g45)));
	assign g194 = (((i_9_) & (!g7) & (!g3) & (!sk[75]) & (!g11) & (!g193)) + ((!i_9_) & (g7) & (g3) & (!sk[75]) & (!g11) & (!g193)) + ((i_9_) & (!g7) & (!g3) & (!sk[75]) & (g11) & (g193)) + ((!i_9_) & (!g7) & (!g3) & (!sk[75]) & (g11) & (g193)) + ((!i_9_) & (g7) & (!g3) & (sk[75]) & (g11) & (!g193)));
	assign g195 = (((!sk[76]) & (g36) & (g11)));
	assign g196 = (((g7) & (!g38) & (!sk[77]) & (!g63) & (!g53) & (!g195)) + ((!g7) & (!g38) & (!sk[77]) & (!g63) & (g53) & (g195)) + ((g7) & (!g38) & (!sk[77]) & (g63) & (!g53) & (!g195)) + ((!g7) & (g38) & (!sk[77]) & (g63) & (!g53) & (!g195)) + ((g7) & (!g38) & (!sk[77]) & (g63) & (!g53) & (g195)));
	assign g197 = (((i_9_) & (!i_8_) & (!sk[78]) & (!i_6_) & (!i_7_) & (!g25)) + ((!i_9_) & (i_8_) & (!sk[78]) & (i_6_) & (!i_7_) & (!g25)) + ((!i_9_) & (!i_8_) & (!sk[78]) & (!i_6_) & (i_7_) & (g25)) + ((!i_9_) & (!i_8_) & (sk[78]) & (!i_6_) & (!i_7_) & (!g25)) + ((!i_9_) & (i_8_) & (sk[78]) & (!i_6_) & (!i_7_) & (g25)));
	assign g198 = (((i_9_) & (!i_8_) & (!sk[79]) & (!g30) & (!g82) & (!g197)) + ((!i_9_) & (i_8_) & (!sk[79]) & (g30) & (!g82) & (!g197)) + ((i_9_) & (!i_8_) & (!sk[79]) & (g30) & (!g82) & (g197)) + ((!i_9_) & (!i_8_) & (!sk[79]) & (!g30) & (g82) & (g197)) + ((!i_9_) & (!i_8_) & (!sk[79]) & (!g30) & (g82) & (g197)));
	assign g199 = (((i_2_) & (!g78) & (!g122) & (!sk[80]) & (!g139) & (!g151)) + ((!i_2_) & (g78) & (g122) & (!sk[80]) & (!g139) & (!g151)) + ((i_2_) & (!g78) & (g122) & (!sk[80]) & (!g139) & (g151)) + ((!i_2_) & (!g78) & (!g122) & (!sk[80]) & (g139) & (g151)) + ((!i_2_) & (g78) & (!g122) & (!sk[80]) & (g139) & (g151)));
	assign g200 = (((!g50) & (!g6) & (!sk[81]) & (g30)) + ((g50) & (g6) & (!sk[81]) & (!g30)) + ((!g50) & (!g6) & (!sk[81]) & (g30)));
	assign g201 = (((!g28) & (sk[82]) & (g138)) + ((g28) & (!sk[82]) & (g138)));
	assign g202 = (((!i_9_) & (!g25) & (g59) & (g183) & (!g141) & (!g201)) + ((!i_9_) & (!g25) & (g59) & (!g183) & (g141) & (!g201)) + ((i_9_) & (g25) & (!g59) & (!g183) & (!g141) & (g201)));
	assign g203 = (((g21) & (!g5) & (!g198) & (!g199) & (!g200) & (!g202)) + ((!g21) & (!g5) & (!g198) & (!g199) & (!g200) & (!g202)));
	assign g204 = (((!sk[85]) & (i_9_) & (!i_8_) & (!i_7_) & (!g59) & (!g14)) + ((!sk[85]) & (!i_9_) & (i_8_) & (i_7_) & (!g59) & (!g14)) + ((!sk[85]) & (!i_9_) & (!i_8_) & (!i_7_) & (g59) & (g14)) + ((!sk[85]) & (i_9_) & (!i_8_) & (i_7_) & (g59) & (!g14)));
	assign g205 = (((i_2_) & (!i_9_) & (!g50) & (!g8) & (!sk[86]) & (!g119)) + ((!i_2_) & (i_9_) & (g50) & (!g8) & (!sk[86]) & (!g119)) + ((!i_2_) & (!i_9_) & (!g50) & (g8) & (!sk[86]) & (g119)) + ((i_2_) & (i_9_) & (!g50) & (g8) & (!sk[86]) & (!g119)) + ((!i_2_) & (!i_9_) & (!g50) & (!g8) & (sk[86]) & (!g119)));
	assign g206 = (((!i_8_) & (sk[87]) & (i_7_)) + ((i_8_) & (!sk[87]) & (i_7_)) + ((i_8_) & (sk[87]) & (!i_7_)));
	assign g207 = (((!i_9_) & (!i_6_) & (!sk[88]) & (g206)) + ((i_9_) & (i_6_) & (!sk[88]) & (!g206)) + ((i_9_) & (!i_6_) & (sk[88]) & (!g206)));
	assign g208 = (((!g28) & (sk[89]) & (g11)) + ((g28) & (!sk[89]) & (g11)));
	assign g209 = (((!g4) & (sk[90]) & (g138)) + ((g4) & (!sk[90]) & (g138)));
	assign g210 = (((i_9_) & (!sk[91]) & (!g25) & (!g18) & (!g208) & (!g209)) + ((!i_9_) & (!sk[91]) & (g25) & (g18) & (!g208) & (!g209)) + ((i_9_) & (!sk[91]) & (!g25) & (g18) & (g208) & (!g209)) + ((!i_9_) & (!sk[91]) & (!g25) & (!g18) & (g208) & (g209)) + ((!i_9_) & (sk[91]) & (g25) & (!g18) & (!g208) & (g209)));
	assign g211 = (((g36) & (!sk[92]) & (g3)) + ((g36) & (sk[92]) & (!g3)));
	assign g212 = (((i_9_) & (!g25) & (!g45) & (!g52) & (!sk[93]) & (!g211)) + ((i_9_) & (!g25) & (!g45) & (g52) & (!sk[93]) & (!g211)) + ((!i_9_) & (g25) & (g45) & (!g52) & (!sk[93]) & (!g211)) + ((!i_9_) & (!g25) & (!g45) & (g52) & (!sk[93]) & (g211)) + ((!i_9_) & (g25) & (!g45) & (!g52) & (sk[93]) & (g211)));
	assign g213 = (((i_5_) & (!g39) & (!sk[94]) & (!g20) & (!g92) & (!g40)) + ((!i_5_) & (g39) & (!sk[94]) & (g20) & (!g92) & (!g40)) + ((!i_5_) & (!g39) & (!sk[94]) & (!g20) & (g92) & (g40)) + ((!i_5_) & (g39) & (!sk[94]) & (g20) & (g92) & (!g40)) + ((i_5_) & (g39) & (!sk[94]) & (!g20) & (g92) & (g40)));
	assign g214 = (((!sk[95]) & (g207) & (g210) & (!g212) & (!g213)) + ((!sk[95]) & (g207) & (!g210) & (!g212) & (g213)) + ((sk[95]) & (!g207) & (!g210) & (!g212) & (!g213)) + ((sk[95]) & (!g207) & (!g210) & (!g212) & (!g213)));
	assign g215 = (((g7) & (!sk[96]) & (g204) & (!g205) & (!g214)) + ((g7) & (!sk[96]) & (!g204) & (!g205) & (g214)) + ((!g7) & (sk[96]) & (!g204) & (!g205) & (g214)) + ((!g7) & (sk[96]) & (!g204) & (!g205) & (g214)));
	assign g216 = (((!sk[97]) & (g192) & (!g194) & (!g196) & (!g203) & (!g215)) + ((!sk[97]) & (!g192) & (g194) & (g196) & (!g203) & (!g215)) + ((!sk[97]) & (!g192) & (!g194) & (!g196) & (g203) & (g215)) + ((!sk[97]) & (!g192) & (!g194) & (!g196) & (g203) & (g215)) + ((!sk[97]) & (!g192) & (!g194) & (!g196) & (g203) & (g215)));
	assign g217 = (((g89) & (g108) & (g758) & (g114) & (g191) & (g216)));
	assign g218 = (((i_9_) & (i_8_) & (!i_6_) & (!i_7_) & (g29) & (!g142)) + ((i_9_) & (i_8_) & (i_6_) & (i_7_) & (!g29) & (!g142)));
	assign g219 = (((g10) & (!sk[100]) & (!g1) & (!g58) & (g218)) + ((g10) & (sk[100]) & (!g1) & (!g58) & (!g218)) + ((!g10) & (sk[100]) & (g1) & (!g58) & (!g218)) + ((!g10) & (sk[100]) & (!g1) & (g58) & (!g218)) + ((g10) & (!sk[100]) & (g1) & (!g58) & (!g218)));
	assign g220 = (((i_9_) & (!g50) & (g124) & (!g59) & (!g134) & (!g77)) + ((!i_9_) & (!g50) & (!g124) & (g59) & (g134) & (!g77)) + ((i_9_) & (!g50) & (!g124) & (g59) & (!g134) & (g77)));
	assign g221 = (((!sk[102]) & (g39) & (g28)) + ((sk[102]) & (g39) & (!g28)));
	assign g222 = (((g76) & (!sk[103]) & (g1)) + ((!g76) & (sk[103]) & (!g1)));
	assign g223 = (((g20) & (!g42) & (!g221) & (!g135) & (!sk[104]) & (!g222)) + ((!g20) & (!g42) & (!g221) & (!g135) & (sk[104]) & (!g222)) + ((!g20) & (!g42) & (!g221) & (!g135) & (sk[104]) & (!g222)) + ((!g20) & (g42) & (g221) & (!g135) & (!sk[104]) & (!g222)) + ((!g20) & (!g42) & (!g221) & (g135) & (!sk[104]) & (g222)) + ((!g20) & (!g42) & (!g221) & (!g135) & (sk[104]) & (!g222)) + ((!g20) & (!g42) & (!g221) & (!g135) & (sk[104]) & (!g222)));
	assign g224 = (((!sk[105]) & (g4) & (g11)) + ((sk[105]) & (!g4) & (g11)));
	assign g225 = (((!sk[106]) & (g50) & (g4)) + ((sk[106]) & (!g50) & (!g4)));
	assign g226 = (((g21) & (g27) & (!sk[107]) & (!g224) & (!g225)) + ((!g21) & (g27) & (sk[107]) & (g224) & (!g225)) + ((!g21) & (!g27) & (sk[107]) & (!g224) & (g225)) + ((g21) & (!g27) & (!sk[107]) & (!g224) & (g225)));
	assign g227 = (((!sk[108]) & (g219) & (g220) & (!g223) & (!g226)) + ((!sk[108]) & (g219) & (!g220) & (!g223) & (g226)) + ((sk[108]) & (g219) & (!g220) & (g223) & (!g226)));
	assign g228 = (((!sk[109]) & (g30) & (g45)) + ((sk[109]) & (g30) & (!g45)));
	assign g229 = (((!g35) & (sk[110]) & (g133) & (!g165) & (!g228)) + ((g35) & (!sk[110]) & (g133) & (!g165) & (!g228)) + ((g35) & (!sk[110]) & (!g133) & (!g165) & (g228)) + ((!g35) & (sk[110]) & (!g133) & (!g165) & (!g228)) + ((!g35) & (sk[110]) & (!g133) & (!g165) & (!g228)) + ((!g35) & (sk[110]) & (g133) & (!g165) & (!g228)));
	assign g230 = (((g8) & (!sk[111]) & (g76)) + ((g8) & (sk[111]) & (!g76)));
	assign g231 = (((g84) & (!g1) & (!g14) & (g40) & (!sk[112]) & (!g142)) + ((g84) & (!g1) & (!g14) & (!g40) & (!sk[112]) & (!g142)) + ((!g84) & (g1) & (g14) & (!g40) & (!sk[112]) & (!g142)) + ((!g84) & (!g1) & (!g14) & (g40) & (!sk[112]) & (g142)) + ((!g84) & (!g1) & (!g14) & (g40) & (sk[112]) & (!g142)) + ((!g84) & (!g1) & (!g14) & (g40) & (!sk[112]) & (g142)));
	assign g232 = (((!sk[113]) & (g42) & (!g2) & (!g186) & (!g230) & (!g231)) + ((!sk[113]) & (!g42) & (g2) & (g186) & (!g230) & (!g231)) + ((!sk[113]) & (!g42) & (!g2) & (!g186) & (g230) & (g231)) + ((sk[113]) & (!g42) & (!g2) & (!g186) & (!g230) & (!g231)) + ((sk[113]) & (!g42) & (!g2) & (!g186) & (!g230) & (!g231)) + ((!sk[113]) & (g42) & (!g2) & (!g186) & (!g230) & (!g231)) + ((!sk[113]) & (g42) & (!g2) & (!g186) & (!g230) & (!g231)));
	assign g233 = (((g30) & (!sk[114]) & (g18)));
	assign g234 = (((!sk[115]) & (g35) & (!g28) & (!g1) & (!g40) & (!g233)) + ((!sk[115]) & (g35) & (!g28) & (!g1) & (!g40) & (g233)) + ((!sk[115]) & (!g35) & (g28) & (g1) & (!g40) & (!g233)) + ((!sk[115]) & (!g35) & (!g28) & (!g1) & (g40) & (g233)) + ((sk[115]) & (!g35) & (!g28) & (!g1) & (g40) & (!g233)));
	assign g235 = (((i_2_) & (i_0_) & (!i_1_) & (!sk[116]) & (!g186)) + ((i_2_) & (!i_0_) & (!i_1_) & (!sk[116]) & (g186)) + ((!i_2_) & (!i_0_) & (i_1_) & (sk[116]) & (!g186)) + ((i_2_) & (!i_0_) & (!i_1_) & (!sk[116]) & (g186)));
	assign g236 = (((!g7) & (!g6) & (g16) & (!g4) & (!g133) & (!g53)) + ((g7) & (!g6) & (!g16) & (!g4) & (!g133) & (g53)));
	assign g237 = (((!i_2_) & (i_9_) & (!g125) & (!g234) & (!g235) & (!g236)) + ((!i_2_) & (!i_9_) & (!g125) & (!g234) & (!g235) & (!g236)) + ((!i_2_) & (!i_9_) & (!g125) & (!g234) & (!g235) & (!g236)));
	assign g238 = (((i_9_) & (!g50) & (!g25) & (!g60) & (!sk[119]) & (!g230)) + ((i_9_) & (!g50) & (!g25) & (g60) & (!sk[119]) & (!g230)) + ((!i_9_) & (g50) & (g25) & (!g60) & (!sk[119]) & (!g230)) + ((!i_9_) & (!g50) & (!g25) & (g60) & (!sk[119]) & (g230)) + ((!i_9_) & (!g50) & (g25) & (!g60) & (sk[119]) & (g230)));
	assign g239 = (((!sk[120]) & (g49) & (g38) & (!g182) & (!g142)) + ((!sk[120]) & (g49) & (!g38) & (!g182) & (g142)) + ((sk[120]) & (!g49) & (!g38) & (!g182) & (!g142)) + ((sk[120]) & (g49) & (!g38) & (g182) & (!g142)));
	assign g240 = (((!sk[121]) & (g22) & (g30)));
	assign g241 = (((i_9_) & (i_8_) & (!i_6_) & (i_7_) & (g26) & (!g240)) + ((i_9_) & (!i_8_) & (i_6_) & (i_7_) & (!g26) & (g240)));
	assign g242 = (((!g42) & (!g233) & (!sk[123]) & (g241)) + ((g42) & (g233) & (!sk[123]) & (!g241)) + ((!g42) & (!g233) & (sk[123]) & (!g241)) + ((!g42) & (!g233) & (sk[123]) & (!g241)));
	assign g243 = (((g20) & (!g28) & (!g25) & (!g137) & (!sk[124]) & (!g74)) + ((g20) & (!g28) & (!g25) & (!g137) & (!sk[124]) & (!g74)) + ((!g20) & (g28) & (g25) & (!g137) & (!sk[124]) & (!g74)) + ((!g20) & (!g28) & (!g25) & (g137) & (!sk[124]) & (g74)) + ((!g20) & (!g28) & (g25) & (g137) & (sk[124]) & (!g74)));
	assign g244 = (((!g10) & (sk[125]) & (g18)) + ((g10) & (!sk[125]) & (g18)));
	assign g245 = (((!sk[126]) & (g22) & (!g38) & (!g73) & (!g4) & (!g10)) + ((!sk[126]) & (!g22) & (g38) & (g73) & (!g4) & (!g10)) + ((!sk[126]) & (g22) & (!g38) & (g73) & (!g4) & (!g10)) + ((!sk[126]) & (!g22) & (!g38) & (!g73) & (g4) & (g10)) + ((!sk[126]) & (g22) & (!g38) & (!g73) & (!g4) & (!g10)));
	assign g246 = (((!g133) & (!g244) & (!sk[127]) & (g245)) + ((!g133) & (!g244) & (sk[127]) & (!g245)) + ((g133) & (g244) & (!sk[127]) & (!g245)));
	assign g247 = (((!g35) & (!g42) & (!g2) & (!g161) & (!g141) & (!g244)) + ((!g35) & (!g42) & (!g2) & (!g161) & (!g141) & (!g244)) + ((!g35) & (!g42) & (!g2) & (!g161) & (!g141) & (!g244)) + ((!g35) & (!g42) & (!g2) & (!g161) & (!g141) & (!g244)) + ((!g35) & (!g42) & (!g2) & (!g161) & (!g141) & (!g244)) + ((!g35) & (!g42) & (!g2) & (!g161) & (!g141) & (!g244)) + ((!g35) & (!g42) & (!g2) & (!g161) & (!g141) & (!g244)) + ((!g35) & (!g42) & (!g2) & (!g161) & (!g141) & (!g244)));
	assign g248 = (((g239) & (!g242) & (!g243) & (!g246) & (!sk[1]) & (!g247)) + ((!g239) & (g242) & (g243) & (!g246) & (!sk[1]) & (!g247)) + ((!g239) & (!g242) & (!g243) & (g246) & (!sk[1]) & (g247)) + ((!g239) & (g242) & (!g243) & (g246) & (!sk[1]) & (g247)));
	assign g249 = (((!sk[2]) & (i_9_) & (!g25) & (!g3) & (!g125) & (!g62)) + ((!sk[2]) & (!i_9_) & (g25) & (g3) & (!g125) & (!g62)) + ((!sk[2]) & (i_9_) & (!g25) & (!g3) & (!g125) & (g62)) + ((!sk[2]) & (!i_9_) & (!g25) & (!g3) & (g125) & (g62)) + ((sk[2]) & (!i_9_) & (g25) & (!g3) & (g125) & (!g62)));
	assign g250 = (((!sk[3]) & (g22) & (!i_9_) & (!g54) & (!g122) & (!g10)) + ((!sk[3]) & (!g22) & (i_9_) & (g54) & (!g122) & (!g10)) + ((!sk[3]) & (g22) & (i_9_) & (!g54) & (g122) & (!g10)) + ((!sk[3]) & (!g22) & (!i_9_) & (!g54) & (g122) & (g10)) + ((!sk[3]) & (g22) & (!i_9_) & (!g54) & (!g122) & (!g10)));
	assign g251 = (((!g76) & (sk[4]) & (g18)) + ((g76) & (!sk[4]) & (g18)));
	assign g252 = (((!g42) & (g13) & (g43) & (!g19) & (!g165) & (!g251)) + ((!g42) & (g13) & (!g43) & (!g19) & (!g165) & (!g251)) + ((!g42) & (!g13) & (g43) & (!g19) & (!g165) & (!g251)) + ((!g42) & (!g13) & (!g43) & (!g19) & (!g165) & (!g251)) + ((!g42) & (g13) & (g43) & (!g19) & (!g165) & (!g251)) + ((!g42) & (g13) & (!g43) & (!g19) & (!g165) & (!g251)) + ((!g42) & (!g13) & (g43) & (!g19) & (!g165) & (!g251)) + ((!g42) & (!g13) & (!g43) & (!g19) & (!g165) & (!g251)));
	assign g253 = (((!g117) & (g133) & (g21) & (!g161) & (!sk[6]) & (!g55)) + ((g117) & (!g133) & (!g21) & (!g161) & (!sk[6]) & (!g55)) + ((!g117) & (g133) & (!g21) & (!g161) & (sk[6]) & (!g55)) + ((!g117) & (!g133) & (!g21) & (g161) & (!sk[6]) & (g55)) + ((!g117) & (!g133) & (g21) & (!g161) & (sk[6]) & (!g55)) + ((!g117) & (!g133) & (!g21) & (!g161) & (sk[6]) & (!g55)));
	assign g254 = (((!g38) & (g73) & (g57) & (!sk[7]) & (!g1) & (!g14)) + ((g38) & (!g73) & (!g57) & (!sk[7]) & (!g1) & (!g14)) + ((!g38) & (!g73) & (!g57) & (!sk[7]) & (g1) & (g14)) + ((!g38) & (!g73) & (!g57) & (sk[7]) & (!g1) & (!g14)));
	assign g255 = (((g249) & (!sk[8]) & (!g250) & (!g252) & (!g253) & (!g254)) + ((!g249) & (!sk[8]) & (g250) & (g252) & (!g253) & (!g254)) + ((!g249) & (!sk[8]) & (!g250) & (!g252) & (g253) & (g254)) + ((!g249) & (sk[8]) & (!g250) & (g252) & (g253) & (!g254)));
	assign g256 = (((!i_2_) & (!i_0_) & (i_1_) & (!g38) & (g30) & (!g40)) + ((!i_2_) & (i_0_) & (i_1_) & (!g38) & (g30) & (g40)) + ((!i_2_) & (!i_0_) & (!i_1_) & (!g38) & (g30) & (g40)));
	assign g257 = (((i_2_) & (g119) & (!g30) & (!sk[10]) & (!g10)) + ((i_2_) & (!g119) & (!g30) & (!sk[10]) & (g10)) + ((!i_2_) & (!g119) & (g30) & (sk[10]) & (!g10)) + ((i_2_) & (!g119) & (!g30) & (sk[10]) & (!g10)));
	assign g258 = (((g21) & (!sk[11]) & (!g58) & (!g85) & (!g141) & (!g257)) + ((g21) & (!sk[11]) & (g58) & (!g85) & (!g141) & (!g257)) + ((g21) & (!sk[11]) & (!g58) & (!g85) & (!g141) & (!g257)) + ((!g21) & (!sk[11]) & (g58) & (g85) & (!g141) & (!g257)) + ((!g21) & (!sk[11]) & (!g58) & (!g85) & (g141) & (g257)) + ((!g21) & (sk[11]) & (g58) & (!g85) & (!g141) & (!g257)) + ((!g21) & (sk[11]) & (!g58) & (!g85) & (!g141) & (!g257)));
	assign g259 = (((g16) & (!sk[12]) & (g14)) + ((g16) & (sk[12]) & (!g14)));
	assign g260 = (((g49) & (!sk[13]) & (g77) & (!g259)) + ((g49) & (!sk[13]) & (!g77) & (g259)) + ((!g49) & (!sk[13]) & (!g77) & (g259)));
	assign g261 = (((g22) & (!g38) & (!g6) & (!g76) & (!sk[14]) & (!g260)) + ((!g22) & (g38) & (g6) & (!g76) & (!sk[14]) & (!g260)) + ((!g22) & (!g38) & (!g6) & (g76) & (!sk[14]) & (g260)) + ((!g22) & (g38) & (!g6) & (!g76) & (sk[14]) & (!g260)) + ((!g22) & (!g38) & (!g6) & (g76) & (sk[14]) & (!g260)) + ((!g22) & (!g38) & (g6) & (!g76) & (sk[14]) & (!g260)));
	assign g262 = (((g133) & (g43) & (!sk[15]) & (!g169) & (!g135) & (!g211)) + ((g133) & (!g43) & (!sk[15]) & (!g169) & (!g135) & (!g211)) + ((!g133) & (g43) & (!sk[15]) & (g169) & (!g135) & (!g211)) + ((g133) & (!g43) & (!sk[15]) & (!g169) & (!g135) & (!g211)) + ((!g133) & (!g43) & (!sk[15]) & (!g169) & (g135) & (g211)) + ((!g133) & (!g43) & (sk[15]) & (!g169) & (!g135) & (!g211)) + ((!g133) & (g43) & (!sk[15]) & (g169) & (!g135) & (!g211)));
	assign g263 = (((!g10) & (sk[16]) & (g27)) + ((g10) & (!sk[16]) & (g27)));
	assign g264 = (((!sk[17]) & (i_9_) & (!g25) & (!g77) & (!g209) & (!g263)) + ((!sk[17]) & (!i_9_) & (g25) & (g77) & (!g209) & (!g263)) + ((!sk[17]) & (i_9_) & (g25) & (!g77) & (g209) & (!g263)) + ((sk[17]) & (!i_9_) & (g25) & (!g77) & (!g209) & (g263)) + ((!sk[17]) & (!i_9_) & (!g25) & (!g77) & (g209) & (g263)));
	assign g265 = (((!i_9_) & (g39) & (g182) & (!g44) & (!g161) & (!g251)) + ((i_9_) & (g39) & (!g182) & (g44) & (!g161) & (!g251)) + ((i_9_) & (g39) & (!g182) & (!g44) & (g161) & (!g251)) + ((!i_9_) & (g39) & (!g182) & (!g44) & (!g161) & (g251)));
	assign g266 = (((g258) & (!sk[19]) & (!g261) & (!g262) & (!g264) & (!g265)) + ((!g258) & (!sk[19]) & (g261) & (g262) & (!g264) & (!g265)) + ((!g258) & (!sk[19]) & (!g261) & (!g262) & (g264) & (g265)) + ((g258) & (!sk[19]) & (g261) & (g262) & (!g264) & (!g265)));
	assign g267 = (((!sk[20]) & (!i_2_) & (!g78) & (g180)) + ((!sk[20]) & (i_2_) & (g78) & (!g180)) + ((sk[20]) & (!i_2_) & (!g78) & (!g180)) + ((!sk[20]) & (!i_2_) & (!g78) & (g180)));
	assign g268 = (((g22) & (!g42) & (!g76) & (!g27) & (!sk[21]) & (!g201)) + ((g22) & (!g42) & (!g76) & (g27) & (!sk[21]) & (!g201)) + ((!g22) & (g42) & (g76) & (!g27) & (!sk[21]) & (!g201)) + ((!g22) & (g42) & (!g76) & (!g27) & (sk[21]) & (g201)) + ((!g22) & (!g42) & (!g76) & (g27) & (!sk[21]) & (g201)));
	assign g269 = (((i_2_) & (!i_9_) & (!g8) & (!g119) & (!sk[22]) & (!g10)) + ((!i_2_) & (!i_9_) & (!g8) & (!g119) & (sk[22]) & (!g10)) + ((!i_2_) & (i_9_) & (g8) & (!g119) & (!sk[22]) & (!g10)) + ((!i_2_) & (!i_9_) & (!g8) & (g119) & (!sk[22]) & (g10)) + ((!i_2_) & (!i_9_) & (g8) & (!g119) & (sk[22]) & (!g10)));
	assign g270 = (((g42) & (!g124) & (!sk[23]) & (!g40) & (g15)) + ((g42) & (g124) & (!sk[23]) & (!g40) & (!g15)) + ((!g42) & (g124) & (sk[23]) & (g40) & (!g15)));
	assign g271 = (((g22) & (!sk[24]) & (!i_9_) & (!g36) & (!g10) & (!g18)) + ((!g22) & (!sk[24]) & (i_9_) & (g36) & (!g10) & (!g18)) + ((!g22) & (!sk[24]) & (!i_9_) & (!g36) & (g10) & (g18)) + ((g22) & (!sk[24]) & (i_9_) & (g36) & (!g10) & (g18)) + ((g22) & (!sk[24]) & (!i_9_) & (!g36) & (!g10) & (g18)));
	assign g272 = (((!i_0_) & (sk[25]) & (i_1_)) + ((i_0_) & (!sk[25]) & (i_1_)));
	assign g273 = (((i_2_) & (!i_9_) & (!g272) & (!sk[26]) & (!g32) & (!g141)) + ((!i_2_) & (i_9_) & (g272) & (!sk[26]) & (!g32) & (!g141)) + ((!i_2_) & (!i_9_) & (!g272) & (!sk[26]) & (g32) & (g141)) + ((!i_2_) & (i_9_) & (g272) & (!sk[26]) & (g32) & (!g141)) + ((i_2_) & (!i_9_) & (g272) & (!sk[26]) & (!g32) & (g141)));
	assign g274 = (((!sk[27]) & (i_2_) & (!i_9_) & (!g119) & (!g31) & (!g139)) + ((!sk[27]) & (!i_2_) & (i_9_) & (g119) & (!g31) & (!g139)) + ((!sk[27]) & (!i_2_) & (!i_9_) & (!g119) & (g31) & (g139)) + ((!sk[27]) & (i_2_) & (i_9_) & (!g119) & (g31) & (!g139)) + ((sk[27]) & (!i_2_) & (!i_9_) & (!g119) & (!g31) & (g139)));
	assign g275 = (((!sk[28]) & (i_5_) & (!g92) & (!g11) & (!g137) & (!g1)) + ((!sk[28]) & (!i_5_) & (g92) & (g11) & (!g137) & (!g1)) + ((!sk[28]) & (!i_5_) & (g92) & (g11) & (g137) & (!g1)) + ((!sk[28]) & (!i_5_) & (!g92) & (!g11) & (g137) & (g1)) + ((!sk[28]) & (i_5_) & (g92) & (!g11) & (g137) & (!g1)));
	assign g276 = (((g271) & (g273) & (!g274) & (!sk[29]) & (!g275)) + ((g271) & (!g273) & (!g274) & (!sk[29]) & (g275)) + ((!g271) & (!g273) & (!g274) & (sk[29]) & (!g275)));
	assign g277 = (((!sk[30]) & (g267) & (!g268) & (!g269) & (!g270) & (!g276)) + ((!sk[30]) & (!g267) & (g268) & (g269) & (!g270) & (!g276)) + ((!sk[30]) & (!g267) & (!g268) & (!g269) & (g270) & (g276)) + ((!sk[30]) & (g267) & (!g268) & (!g269) & (!g270) & (g276)) + ((sk[30]) & (!g267) & (!g268) & (!g269) & (!g270) & (g276)));
	assign g278 = (((!g238) & (g248) & (g255) & (!g256) & (g266) & (g277)));
	assign g279 = (((!sk[32]) & (g43) & (g21) & (!g51) & (!g157)) + ((sk[32]) & (!g43) & (!g21) & (g51) & (!g157)) + ((!sk[32]) & (g43) & (!g21) & (!g51) & (g157)) + ((sk[32]) & (!g43) & (!g21) & (!g51) & (g157)));
	assign g280 = (((g20) & (!g122) & (!g43) & (!g179) & (!sk[33]) & (!g60)) + ((!g20) & (!g122) & (!g43) & (g179) & (!sk[33]) & (g60)) + ((!g20) & (!g122) & (!g43) & (!g179) & (sk[33]) & (!g60)) + ((!g20) & (g122) & (g43) & (!g179) & (!sk[33]) & (!g60)) + ((!g20) & (!g122) & (g43) & (!g179) & (sk[33]) & (!g60)) + ((!g20) & (!g122) & (g43) & (!g179) & (sk[33]) & (!g60)) + ((!g20) & (!g122) & (!g43) & (!g179) & (sk[33]) & (!g60)));
	assign g281 = (((g57) & (!sk[34]) & (g137) & (!g2) & (!g201)) + ((g57) & (!sk[34]) & (!g137) & (!g2) & (g201)) + ((!g57) & (sk[34]) & (!g137) & (g2) & (g201)));
	assign g282 = (((!g38) & (!sk[35]) & (!g175) & (g26)) + ((g38) & (!sk[35]) & (g175) & (!g26)) + ((!g38) & (sk[35]) & (!g175) & (!g26)) + ((g38) & (!sk[35]) & (!g175) & (g26)));
	assign g283 = (((g73) & (!sk[36]) & (!g43) & (!g64) & (!g85) & (!g240)) + ((!g73) & (sk[36]) & (!g43) & (!g64) & (!g85) & (!g240)) + ((!g73) & (!sk[36]) & (!g43) & (!g64) & (g85) & (g240)) + ((!g73) & (sk[36]) & (g43) & (!g64) & (!g85) & (!g240)) + ((!g73) & (!sk[36]) & (g43) & (g64) & (!g85) & (!g240)) + ((!g73) & (sk[36]) & (g43) & (!g64) & (!g85) & (!g240)) + ((!g73) & (sk[36]) & (!g43) & (!g64) & (!g85) & (!g240)));
	assign g284 = (((!sk[37]) & (i_9_) & (!g50) & (!g28) & (!g63) & (!g45)) + ((!sk[37]) & (!i_9_) & (g50) & (g28) & (!g63) & (!g45)) + ((!sk[37]) & (!i_9_) & (!g50) & (!g28) & (g63) & (g45)) + ((!sk[37]) & (i_9_) & (!g50) & (!g28) & (g63) & (!g45)) + ((sk[37]) & (!i_9_) & (!g50) & (!g28) & (g63) & (!g45)));
	assign g285 = (((i_2_) & (i_0_) & (i_1_) & (g7) & (!g36) & (g40)) + ((i_2_) & (!i_0_) & (!i_1_) & (g7) & (!g36) & (g40)) + ((!i_2_) & (i_0_) & (i_1_) & (!g7) & (g36) & (g40)));
	assign g286 = (((g54) & (!sk[39]) & (!g10) & (!g133) & (!g284) & (!g285)) + ((!g54) & (!sk[39]) & (g10) & (g133) & (!g284) & (!g285)) + ((!g54) & (!sk[39]) & (!g10) & (!g133) & (g284) & (g285)) + ((g54) & (!sk[39]) & (!g10) & (!g133) & (!g284) & (!g285)) + ((!g54) & (sk[39]) & (g10) & (!g133) & (!g284) & (!g285)) + ((!g54) & (sk[39]) & (!g10) & (g133) & (!g284) & (!g285)));
	assign g287 = (((!sk[40]) & (g21) & (!g158) & (!g282) & (!g283) & (!g286)) + ((!sk[40]) & (!g21) & (g158) & (g282) & (!g283) & (!g286)) + ((!sk[40]) & (!g21) & (!g158) & (!g282) & (g283) & (g286)) + ((!sk[40]) & (g21) & (!g158) & (g282) & (g283) & (g286)) + ((!sk[40]) & (!g21) & (!g158) & (g282) & (g283) & (g286)));
	assign g288 = (((i_2_) & (!sk[41]) & (!g78) & (!i_9_) & (!g117) & (!g230)) + ((!i_2_) & (!sk[41]) & (g78) & (i_9_) & (!g117) & (!g230)) + ((!i_2_) & (!sk[41]) & (!g78) & (!i_9_) & (g117) & (g230)) + ((i_2_) & (!sk[41]) & (g78) & (!i_9_) & (g117) & (!g230)) + ((!i_2_) & (sk[41]) & (g78) & (!i_9_) & (!g117) & (g230)));
	assign g289 = (((g76) & (!sk[42]) & (!g1) & (!g40) & (!g150) & (!g288)) + ((!g76) & (!sk[42]) & (g1) & (g40) & (!g150) & (!g288)) + ((!g76) & (!sk[42]) & (!g1) & (!g40) & (g150) & (g288)) + ((g76) & (!sk[42]) & (!g1) & (!g40) & (!g150) & (!g288)) + ((!g76) & (sk[42]) & (!g1) & (!g40) & (!g150) & (!g288)) + ((!g76) & (!sk[42]) & (g1) & (g40) & (!g150) & (!g288)));
	assign g290 = (((g279) & (!g729) & (!g281) & (!g287) & (!sk[43]) & (!g289)) + ((!g279) & (g729) & (g281) & (!g287) & (!sk[43]) & (!g289)) + ((!g279) & (!g729) & (!g281) & (g287) & (!sk[43]) & (g289)) + ((!g279) & (g729) & (!g281) & (g287) & (!sk[43]) & (g289)));
	assign g291 = (((i_9_) & (!i_5_) & (i_3_) & (!i_4_) & (!g3) & (!g45)) + ((!i_9_) & (i_5_) & (i_3_) & (!i_4_) & (!g3) & (!g45)));
	assign g292 = (((!sk[45]) & (i_0_) & (i_1_) & (!g9) & (!g46)) + ((!sk[45]) & (i_0_) & (!i_1_) & (!g9) & (g46)) + ((sk[45]) & (!i_0_) & (i_1_) & (g9) & (!g46)));
	assign g293 = (((i_2_) & (!i_9_) & (!g119) & (!g125) & (!g117) & (g292)) + ((!i_2_) & (!i_9_) & (!g119) & (g125) & (!g117) & (!g292)) + ((i_2_) & (!i_9_) & (!g119) & (!g125) & (g117) & (!g292)));
	assign g294 = (((!g73) & (!sk[47]) & (!g23) & (g293)) + ((g73) & (!sk[47]) & (g23) & (!g293)) + ((!g73) & (sk[47]) & (!g23) & (!g293)) + ((!g73) & (sk[47]) & (!g23) & (!g293)));
	assign g295 = (((!sk[48]) & (g35) & (!g28) & (!g2) & (!g18) & (!g225)) + ((!sk[48]) & (!g35) & (g28) & (g2) & (!g18) & (!g225)) + ((!sk[48]) & (g35) & (!g28) & (!g2) & (g18) & (!g225)) + ((sk[48]) & (!g35) & (!g28) & (g2) & (!g18) & (g225)) + ((!sk[48]) & (!g35) & (!g28) & (!g2) & (g18) & (g225)));
	assign g296 = (((g181) & (g70) & (!sk[49]) & (!g295) & (!g189)) + ((g181) & (!g70) & (!sk[49]) & (!g295) & (g189)) + ((!g181) & (!g70) & (sk[49]) & (!g295) & (g189)));
	assign g297 = (((!g59) & (g290) & (g722) & (!g291) & (g294) & (g296)) + ((!g59) & (g290) & (g722) & (!g291) & (g294) & (g296)));
	assign g298 = (((g227) & (g735) & (g232) & (g237) & (g278) & (g297)));
	assign g299 = (((g22) & (!i_9_) & (!sk[52]) & (!g25) & (!g134) & (!g171)) + ((!g22) & (i_9_) & (!sk[52]) & (g25) & (!g134) & (!g171)) + ((g22) & (i_9_) & (!sk[52]) & (!g25) & (!g134) & (g171)) + ((!g22) & (!i_9_) & (!sk[52]) & (!g25) & (g134) & (g171)) + ((!g22) & (!i_9_) & (sk[52]) & (g25) & (g134) & (!g171)));
	assign g300 = (((!sk[53]) & (g22) & (!g73) & (!g30) & (!g11) & (!g137)) + ((!sk[53]) & (!g22) & (g73) & (g30) & (!g11) & (!g137)) + ((!sk[53]) & (g22) & (g73) & (g30) & (!g11) & (!g137)) + ((!sk[53]) & (!g22) & (!g73) & (!g30) & (g11) & (g137)) + ((!sk[53]) & (!g22) & (!g73) & (g30) & (g11) & (g137)));
	assign g301 = (((!sk[54]) & (g20) & (!g6) & (!g10) & (g300)) + ((sk[54]) & (!g20) & (!g6) & (!g10) & (!g300)) + ((sk[54]) & (!g20) & (!g6) & (g10) & (!g300)) + ((!sk[54]) & (g20) & (g6) & (!g10) & (!g300)));
	assign g302 = (((!sk[55]) & (g6) & (g76)) + ((sk[55]) & (!g6) & (!g76)));
	assign g303 = (((g28) & (!sk[56]) & (!g42) & (!g63) & (!g40) & (!g139)) + ((!g28) & (!sk[56]) & (g42) & (g63) & (!g40) & (!g139)) + ((!g28) & (sk[56]) & (g42) & (!g63) & (!g40) & (g139)) + ((!g28) & (!sk[56]) & (!g42) & (!g63) & (g40) & (g139)) + ((!g28) & (sk[56]) & (!g42) & (g63) & (g40) & (!g139)));
	assign g304 = (((!sk[57]) & (!g27) & (!g302) & (g303)) + ((!sk[57]) & (g27) & (g302) & (!g303)) + ((sk[57]) & (!g27) & (!g302) & (!g303)) + ((sk[57]) & (!g27) & (!g302) & (!g303)));
	assign g305 = (((!sk[58]) & (i_9_) & (!g50) & (!g7) & (!g6) & (!g62)) + ((!sk[58]) & (!i_9_) & (g50) & (g7) & (!g6) & (!g62)) + ((!sk[58]) & (i_9_) & (!g50) & (!g7) & (!g6) & (g62)) + ((!sk[58]) & (!i_9_) & (!g50) & (!g7) & (g6) & (g62)) + ((sk[58]) & (!i_9_) & (!g50) & (g7) & (!g6) & (!g62)));
	assign g306 = (((!g49) & (!g28) & (!sk[59]) & (g18)) + ((g49) & (g28) & (!sk[59]) & (!g18)) + ((g49) & (!g28) & (!sk[59]) & (g18)));
	assign g307 = (((!g76) & (sk[60]) & (g59)) + ((g76) & (!sk[60]) & (g59)));
	assign g308 = (((g22) & (!g10) & (!g53) & (!g306) & (!sk[61]) & (!g307)) + ((!g22) & (!g10) & (!g53) & (!g306) & (sk[61]) & (!g307)) + ((!g22) & (g10) & (g53) & (!g306) & (!sk[61]) & (!g307)) + ((!g22) & (!g10) & (!g53) & (g306) & (!sk[61]) & (g307)) + ((!g22) & (!g10) & (!g53) & (!g306) & (sk[61]) & (!g307)) + ((!g22) & (g10) & (!g53) & (!g306) & (sk[61]) & (!g307)));
	assign g309 = (((!sk[62]) & (g49) & (!g1) & (!g183) & (!g14) & (!g40)) + ((!sk[62]) & (g49) & (!g1) & (g183) & (!g14) & (!g40)) + ((!sk[62]) & (!g49) & (g1) & (g183) & (!g14) & (!g40)) + ((!sk[62]) & (!g49) & (!g1) & (!g183) & (g14) & (g40)) + ((sk[62]) & (!g49) & (!g1) & (!g183) & (!g14) & (g40)));
	assign g310 = (((g22) & (!g38) & (!g36) & (!sk[63]) & (!g39) & (!g58)) + ((!g22) & (g38) & (g36) & (!sk[63]) & (!g39) & (!g58)) + ((!g22) & (!g38) & (!g36) & (!sk[63]) & (g39) & (g58)) + ((g22) & (!g38) & (g36) & (!sk[63]) & (!g39) & (!g58)) + ((!g22) & (!g38) & (g36) & (sk[63]) & (g39) & (!g58)));
	assign g311 = (((!g35) & (!sk[64]) & (!g170) & (g310)) + ((g35) & (!sk[64]) & (g170) & (!g310)) + ((!g35) & (sk[64]) & (!g170) & (!g310)) + ((!g35) & (sk[64]) & (!g170) & (!g310)));
	assign g312 = (((g49) & (!g141) & (!g308) & (!g309) & (!sk[65]) & (!g311)) + ((!g49) & (g141) & (g308) & (!g309) & (!sk[65]) & (!g311)) + ((!g49) & (!g141) & (!g308) & (g309) & (!sk[65]) & (g311)) + ((!g49) & (!g141) & (g308) & (!g309) & (sk[65]) & (g311)) + ((!g49) & (!g141) & (g308) & (!g309) & (sk[65]) & (g311)));
	assign g313 = (((g76) & (!sk[66]) & (!g3) & (!g13) & (!g305) & (!g312)) + ((!g76) & (!sk[66]) & (g3) & (g13) & (!g305) & (!g312)) + ((!g76) & (!sk[66]) & (!g3) & (!g13) & (g305) & (g312)) + ((g76) & (!sk[66]) & (!g3) & (!g13) & (!g305) & (g312)) + ((!g76) & (sk[66]) & (g3) & (!g13) & (!g305) & (g312)) + ((!g76) & (sk[66]) & (!g3) & (g13) & (!g305) & (g312)));
	assign g314 = (((g234) & (!g299) & (!g301) & (!g304) & (!sk[67]) & (!g313)) + ((!g234) & (g299) & (g301) & (!g304) & (!sk[67]) & (!g313)) + ((!g234) & (!g299) & (!g301) & (g304) & (!sk[67]) & (g313)) + ((!g234) & (!g299) & (g301) & (g304) & (!sk[67]) & (g313)));
	assign g315 = (((i_9_) & (!g39) & (!sk[68]) & (!g3) & (!g55) & (!g302)) + ((!i_9_) & (g39) & (!sk[68]) & (g3) & (!g55) & (!g302)) + ((i_9_) & (!g39) & (!sk[68]) & (!g3) & (!g55) & (g302)) + ((!i_9_) & (!g39) & (!sk[68]) & (!g3) & (g55) & (g302)) + ((!i_9_) & (g39) & (sk[68]) & (!g3) & (g55) & (!g302)));
	assign g316 = (((!sk[69]) & (g73) & (!g133) & (!g64) & (!g19) & (!g208)) + ((sk[69]) & (!g73) & (!g133) & (!g64) & (!g19) & (!g208)) + ((!sk[69]) & (!g73) & (!g133) & (!g64) & (g19) & (g208)) + ((sk[69]) & (!g73) & (g133) & (!g64) & (!g19) & (!g208)) + ((!sk[69]) & (!g73) & (g133) & (g64) & (!g19) & (!g208)) + ((sk[69]) & (!g73) & (g133) & (!g64) & (!g19) & (!g208)) + ((!sk[69]) & (g73) & (!g133) & (!g64) & (!g19) & (!g208)));
	assign g317 = (((g2) & (g251) & (!sk[70]) & (!g315) & (!g316)) + ((g2) & (!g251) & (!sk[70]) & (!g315) & (g316)) + ((!g2) & (!g251) & (sk[70]) & (!g315) & (g316)) + ((!g2) & (!g251) & (sk[70]) & (!g315) & (g316)));
	assign g318 = (((!sk[71]) & (g38) & (g94) & (!g58) & (!g23)) + ((sk[71]) & (!g38) & (g94) & (!g58) & (!g23)) + ((!sk[71]) & (g38) & (!g94) & (!g58) & (g23)) + ((sk[71]) & (!g38) & (!g94) & (!g58) & (g23)));
	assign g319 = (((g28) & (!g73) & (!g63) & (!g13) & (!sk[72]) & (!g18)) + ((!g28) & (g73) & (g63) & (!g13) & (!sk[72]) & (!g18)) + ((!g28) & (!g73) & (!g63) & (g13) & (!sk[72]) & (g18)) + ((!g28) & (!g73) & (!g63) & (!g13) & (sk[72]) & (g18)));
	assign g320 = (((g73) & (g26) & (!g318) & (!sk[73]) & (!g319)) + ((g73) & (!g26) & (!g318) & (!sk[73]) & (g319)) + ((!g73) & (!g26) & (!g318) & (sk[73]) & (!g319)) + ((!g73) & (!g26) & (!g318) & (sk[73]) & (!g319)));
	assign g321 = (((g7) & (g20) & (!sk[74]) & (!g6) & (!g320)) + ((!g7) & (!g20) & (sk[74]) & (!g6) & (g320)) + ((g7) & (!g20) & (!sk[74]) & (!g6) & (g320)) + ((!g7) & (!g20) & (sk[74]) & (g6) & (g320)));
	assign g322 = (((!sk[75]) & (i_9_) & (!g6) & (!g45) & (!g94) & (!g171)) + ((!sk[75]) & (!i_9_) & (g6) & (g45) & (!g94) & (!g171)) + ((!sk[75]) & (i_9_) & (!g6) & (!g45) & (g94) & (!g171)) + ((!sk[75]) & (!i_9_) & (!g6) & (!g45) & (g94) & (g171)) + ((sk[75]) & (!i_9_) & (!g6) & (!g45) & (!g94) & (g171)));
	assign g323 = (((!g73) & (!g57) & (!g94) & (!g58) & (!g82) & (!g195)) + ((!g73) & (!g57) & (!g94) & (g58) & (!g82) & (!g195)) + ((!g73) & (!g57) & (!g94) & (!g58) & (!g82) & (!g195)) + ((!g73) & (!g57) & (!g94) & (g58) & (!g82) & (!g195)));
	assign g324 = (((g49) & (!g35) & (g170) & (sk[77]) & (!g228)) + ((g49) & (g35) & (!g170) & (!sk[77]) & (!g228)) + ((!g49) & (g35) & (!g170) & (sk[77]) & (g228)) + ((g49) & (!g35) & (!g170) & (!sk[77]) & (g228)));
	assign g325 = (((!sk[78]) & (g53) & (!g112) & (!g322) & (!g323) & (!g324)) + ((!sk[78]) & (!g53) & (g112) & (g322) & (!g323) & (!g324)) + ((!sk[78]) & (!g53) & (!g112) & (!g322) & (g323) & (g324)) + ((sk[78]) & (!g53) & (!g112) & (!g322) & (g323) & (!g324)) + ((!sk[78]) & (g53) & (!g112) & (!g322) & (g323) & (!g324)));
	assign g326 = (((g7) & (!g35) & (!sk[79]) & (!g16) & (!g2) & (!g225)) + ((!g7) & (g35) & (!sk[79]) & (g16) & (!g2) & (!g225)) + ((g7) & (!g35) & (!sk[79]) & (g16) & (g2) & (!g225)) + ((!g7) & (g35) & (sk[79]) & (!g16) & (!g2) & (g225)) + ((g7) & (!g35) & (!sk[79]) & (g16) & (!g2) & (g225)) + ((!g7) & (!g35) & (!sk[79]) & (!g16) & (g2) & (g225)));
	assign g327 = (((i_9_) & (!g50) & (!g7) & (!sk[80]) & (g31)) + ((i_9_) & (g50) & (!g7) & (!sk[80]) & (!g31)) + ((!i_9_) & (!g50) & (g7) & (sk[80]) & (!g31)));
	assign g328 = (((g59) & (!g131) & (!g325) & (!g326) & (!sk[81]) & (!g327)) + ((!g59) & (g131) & (g325) & (!g326) & (!sk[81]) & (!g327)) + ((!g59) & (!g131) & (!g325) & (g326) & (!sk[81]) & (g327)) + ((!g59) & (!g131) & (g325) & (!g326) & (sk[81]) & (!g327)) + ((!g59) & (!g131) & (g325) & (!g326) & (sk[81]) & (!g327)) + ((!g59) & (!g131) & (g325) & (!g326) & (sk[81]) & (!g327)) + ((!g59) & (!g131) & (g325) & (!g326) & (sk[81]) & (!g327)));
	assign g329 = (((g22) & (!i_5_) & (!i_3_) & (!i_4_) & (!g20) & (g207)) + ((g22) & (!i_5_) & (!i_3_) & (!i_4_) & (g20) & (g207)));
	assign g330 = (((!sk[83]) & (i_2_) & (!g272) & (!g168) & (!g79) & (!g97)) + ((!sk[83]) & (!i_2_) & (g272) & (g168) & (!g79) & (!g97)) + ((!sk[83]) & (!i_2_) & (!g272) & (!g168) & (g79) & (g97)) + ((!sk[83]) & (i_2_) & (!g272) & (!g168) & (g79) & (g97)) + ((!sk[83]) & (!i_2_) & (g272) & (g168) & (g79) & (!g97)));
	assign g331 = (((i_9_) & (i_8_) & (!sk[84]) & (!i_6_) & (!i_7_)) + ((i_9_) & (!i_8_) & (!sk[84]) & (!i_6_) & (i_7_)) + ((i_9_) & (!i_8_) & (!sk[84]) & (!i_6_) & (i_7_)) + ((i_9_) & (!i_8_) & (sk[84]) & (i_6_) & (!i_7_)));
	assign g332 = (((g38) & (!sk[85]) & (!g137) & (!g64) & (!g195) & (!g331)) + ((!g38) & (!sk[85]) & (g137) & (g64) & (!g195) & (!g331)) + ((!g38) & (!sk[85]) & (g137) & (g64) & (!g195) & (g331)) + ((!g38) & (!sk[85]) & (!g137) & (!g64) & (g195) & (g331)) + ((!g38) & (!sk[85]) & (!g137) & (g64) & (g195) & (g331)));
	assign g333 = (((i_9_) & (!g50) & (!sk[86]) & (!g36) & (!g6) & (!g170)) + ((!i_9_) & (g50) & (!sk[86]) & (g36) & (!g6) & (!g170)) + ((!i_9_) & (!g50) & (!sk[86]) & (!g36) & (g6) & (g170)) + ((i_9_) & (!g50) & (!sk[86]) & (g36) & (!g6) & (!g170)) + ((!i_9_) & (!g50) & (sk[86]) & (!g36) & (!g6) & (g170)));
	assign g334 = (((g21) & (g60) & (!sk[87]) & (!g27) & (!g171)) + ((!g21) & (g60) & (sk[87]) & (g27) & (!g171)) + ((!g21) & (!g60) & (sk[87]) & (!g27) & (g171)) + ((g21) & (!g60) & (!sk[87]) & (!g27) & (g171)));
	assign g335 = (((g40) & (!sk[88]) & (!g195) & (!g332) & (!g333) & (!g334)) + ((!g40) & (!sk[88]) & (g195) & (g332) & (!g333) & (!g334)) + ((!g40) & (!sk[88]) & (!g195) & (!g332) & (g333) & (g334)) + ((!g40) & (sk[88]) & (!g195) & (!g332) & (!g333) & (!g334)) + ((!g40) & (sk[88]) & (!g195) & (!g332) & (!g333) & (!g334)));
	assign g336 = (((g28) & (!g40) & (!g329) & (!sk[89]) & (!g330) & (!g335)) + ((!g28) & (g40) & (g329) & (!sk[89]) & (!g330) & (!g335)) + ((!g28) & (!g40) & (!g329) & (!sk[89]) & (g330) & (g335)) + ((g28) & (!g40) & (!g329) & (!sk[89]) & (!g330) & (g335)) + ((!g28) & (!g40) & (!g329) & (sk[89]) & (!g330) & (g335)));
	assign g337 = (((i_9_) & (!g39) & (!g30) & (!g44) & (!sk[90]) & (!g58)) + ((!i_9_) & (g39) & (g30) & (!g44) & (!sk[90]) & (!g58)) + ((!i_9_) & (!g39) & (!g30) & (g44) & (!sk[90]) & (g58)) + ((!i_9_) & (g39) & (g30) & (!g44) & (!sk[90]) & (!g58)) + ((!i_9_) & (g39) & (!g30) & (g44) & (sk[90]) & (!g58)));
	assign g338 = (((!g49) & (!g53) & (!g82) & (!g19) & (!g230) & (!g337)) + ((!g49) & (!g53) & (!g82) & (!g19) & (!g230) & (!g337)) + ((!g49) & (!g53) & (!g82) & (!g19) & (!g230) & (!g337)) + ((!g49) & (!g53) & (!g82) & (!g19) & (!g230) & (!g337)));
	assign g339 = (((!g22) & (i_9_) & (!g28) & (g84) & (!g45) & (!g177)) + ((g22) & (i_9_) & (!g28) & (!g84) & (!g45) & (g177)) + ((g22) & (!i_9_) & (!g28) & (!g84) & (!g45) & (!g177)));
	assign g340 = (((!g30) & (!g11) & (!sk[93]) & (g58)) + ((g30) & (g11) & (!sk[93]) & (!g58)));
	assign g341 = (((g39) & (!g10) & (!sk[94]) & (!g53) & (!g144) & (!g340)) + ((!g39) & (g10) & (!sk[94]) & (g53) & (!g144) & (!g340)) + ((!g39) & (!g10) & (!sk[94]) & (!g53) & (g144) & (g340)) + ((!g39) & (!g10) & (sk[94]) & (!g53) & (!g144) & (!g340)) + ((!g39) & (!g10) & (sk[94]) & (!g53) & (!g144) & (!g340)) + ((!g39) & (g10) & (!sk[94]) & (g53) & (!g144) & (!g340)));
	assign g342 = (((g116) & (g59) & (!g10) & (!g43) & (!g137) & (!g259)) + ((!g116) & (!g59) & (!g10) & (!g43) & (!g137) & (g259)) + ((!g116) & (g59) & (!g10) & (!g43) & (g137) & (!g259)));
	assign g343 = (((!g49) & (!i_6_) & (g36) & (g39) & (g73) & (!g206)) + ((g49) & (i_6_) & (g36) & (!g39) & (!g73) & (!g206)));
	assign g344 = (((i_9_) & (!i_8_) & (!i_6_) & (!i_7_) & (!sk[97]) & (!i_5_)) + ((!i_9_) & (i_8_) & (i_6_) & (!i_7_) & (!sk[97]) & (!i_5_)) + ((!i_9_) & (!i_8_) & (!i_6_) & (i_7_) & (!sk[97]) & (i_5_)) + ((i_9_) & (i_8_) & (i_6_) & (!i_7_) & (!sk[97]) & (i_5_)) + ((i_9_) & (!i_8_) & (!i_6_) & (!i_7_) & (!sk[97]) & (!i_5_)));
	assign g345 = (((!sk[98]) & (i_3_) & (i_4_) & (!g63) & (!g344)) + ((!sk[98]) & (i_3_) & (!i_4_) & (!g63) & (g344)) + ((sk[98]) & (!i_3_) & (!i_4_) & (g63) & (g344)));
	assign g346 = (((!sk[99]) & (i_6_) & (!g76) & (!g9) & (!g133) & (!g206)) + ((!sk[99]) & (!i_6_) & (g76) & (g9) & (!g133) & (!g206)) + ((sk[99]) & (!i_6_) & (!g76) & (g9) & (!g133) & (!g206)) + ((!sk[99]) & (!i_6_) & (!g76) & (!g9) & (g133) & (g206)) + ((sk[99]) & (!i_6_) & (!g76) & (!g9) & (!g133) & (!g206)));
	assign g347 = (((g38) & (g28) & (!sk[100]) & (!g10) & (!g1)) + ((g38) & (!g28) & (!sk[100]) & (!g10) & (g1)) + ((!g38) & (!g28) & (sk[100]) & (!g10) & (!g1)) + ((!g38) & (!g28) & (sk[100]) & (!g10) & (!g1)));
	assign g348 = (((g35) & (!g169) & (!sk[101]) & (!g345) & (!g346) & (!g347)) + ((!g35) & (g169) & (!sk[101]) & (g345) & (!g346) & (!g347)) + ((!g35) & (!g169) & (!sk[101]) & (!g345) & (g346) & (g347)) + ((!g35) & (!g169) & (sk[101]) & (!g345) & (!g346) & (!g347)) + ((!g35) & (!g169) & (sk[101]) & (!g345) & (!g346) & (!g347)));
	assign g349 = (((!sk[102]) & (g339) & (!g341) & (!g342) & (!g343) & (!g348)) + ((!sk[102]) & (!g339) & (g341) & (g342) & (!g343) & (!g348)) + ((!sk[102]) & (!g339) & (!g341) & (!g342) & (g343) & (g348)) + ((sk[102]) & (!g339) & (g341) & (!g342) & (!g343) & (g348)));
	assign g350 = (((i_6_) & (i_7_) & (!sk[103]) & (!i_5_) & (!i_3_)) + ((i_6_) & (!i_7_) & (!sk[103]) & (!i_5_) & (i_3_)) + ((!i_6_) & (!i_7_) & (sk[103]) & (!i_5_) & (i_3_)));
	assign g351 = (((g22) & (!i_9_) & (!i_8_) & (!i_4_) & (!sk[104]) & (!g350)) + ((!g22) & (i_9_) & (i_8_) & (!i_4_) & (!sk[104]) & (!g350)) + ((!g22) & (!i_9_) & (!i_8_) & (i_4_) & (!sk[104]) & (g350)) + ((g22) & (i_9_) & (!i_8_) & (i_4_) & (!sk[104]) & (g350)) + ((g22) & (i_9_) & (i_8_) & (!i_4_) & (!sk[104]) & (g350)));
	assign g352 = (((!sk[105]) & (i_2_) & (i_9_) & (!i_7_) & (!g272)) + ((!sk[105]) & (i_2_) & (!i_9_) & (!i_7_) & (g272)) + ((!sk[105]) & (i_2_) & (!i_9_) & (!i_7_) & (g272)) + ((sk[105]) & (!i_2_) & (!i_9_) & (i_7_) & (g272)));
	assign g353 = (((i_8_) & (i_6_) & (!g4) & (!sk[106]) & (!g352)) + ((i_8_) & (!i_6_) & (!g4) & (!sk[106]) & (g352)) + ((i_8_) & (i_6_) & (!g4) & (!sk[106]) & (g352)));
	assign g354 = (((!sk[107]) & (g7) & (g25)));
	assign g355 = (((i_9_) & (!i_8_) & (!sk[108]) & (!g83) & (!g82) & (!g354)) + ((!i_9_) & (i_8_) & (!sk[108]) & (g83) & (!g82) & (!g354)) + ((!i_9_) & (!i_8_) & (!sk[108]) & (!g83) & (g82) & (g354)) + ((i_9_) & (i_8_) & (!sk[108]) & (g83) & (g82) & (!g354)) + ((i_9_) & (!i_8_) & (!sk[108]) & (g83) & (!g82) & (g354)));
	assign g356 = (((!sk[109]) & (g10) & (g138)) + ((sk[109]) & (!g10) & (g138)));
	assign g357 = (((i_2_) & (!g119) & (!g157) & (!g151) & (!sk[110]) & (!g356)) + ((i_2_) & (!g119) & (g157) & (g151) & (!sk[110]) & (!g356)) + ((!i_2_) & (g119) & (g157) & (!g151) & (!sk[110]) & (!g356)) + ((!i_2_) & (!g119) & (!g157) & (g151) & (!sk[110]) & (g356)) + ((!i_2_) & (!g119) & (!g157) & (g151) & (!sk[110]) & (g356)));
	assign g358 = (((!i_2_) & (!i_9_) & (!i_8_) & (!i_6_) & (sk[111]) & (!i_7_)) + ((!i_2_) & (i_9_) & (i_8_) & (!i_6_) & (!sk[111]) & (!i_7_)) + ((i_2_) & (!i_9_) & (i_8_) & (!i_6_) & (!sk[111]) & (!i_7_)) + ((!i_2_) & (!i_9_) & (!i_8_) & (!i_6_) & (sk[111]) & (!i_7_)) + ((i_2_) & (!i_9_) & (!i_8_) & (!i_6_) & (!sk[111]) & (!i_7_)) + ((!i_2_) & (!i_9_) & (!i_8_) & (i_6_) & (!sk[111]) & (i_7_)) + ((!i_2_) & (!i_9_) & (!i_8_) & (!i_6_) & (sk[111]) & (!i_7_)));
	assign g359 = (((!g38) & (!sk[112]) & (!g28) & (g59)) + ((g38) & (!sk[112]) & (g28) & (!g59)) + ((!g38) & (!sk[112]) & (!g28) & (g59)));
	assign g360 = (((g40) & (!g27) & (!g142) & (!sk[113]) & (!g90) & (!g359)) + ((!g40) & (g27) & (g142) & (!sk[113]) & (!g90) & (!g359)) + ((!g40) & (!g27) & (!g142) & (!sk[113]) & (g90) & (g359)) + ((!g40) & (!g27) & (!g142) & (sk[113]) & (!g90) & (!g359)) + ((!g40) & (!g27) & (g142) & (sk[113]) & (!g90) & (!g359)) + ((!g40) & (!g27) & (!g142) & (sk[113]) & (!g90) & (!g359)) + ((!g40) & (!g27) & (g142) & (sk[113]) & (!g90) & (!g359)));
	assign g361 = (((g20) & (!g307) & (!sk[114]) & (!g357) & (!g711) & (!g360)) + ((!g20) & (g307) & (!sk[114]) & (g357) & (!g711) & (!g360)) + ((!g20) & (!g307) & (!sk[114]) & (!g357) & (g711) & (g360)) + ((!g20) & (!g307) & (!sk[114]) & (!g357) & (g711) & (g360)) + ((!g20) & (!g307) & (!sk[114]) & (!g357) & (g711) & (g360)));
	assign g362 = (((!sk[115]) & (g56) & (!g351) & (!g353) & (!g355) & (!g361)) + ((!sk[115]) & (!g56) & (g351) & (g353) & (!g355) & (!g361)) + ((!sk[115]) & (!g56) & (!g351) & (!g353) & (g355) & (g361)) + ((sk[115]) & (!g56) & (!g351) & (!g353) & (!g355) & (g361)));
	assign g363 = (((g729) & (g248) & (g336) & (g338) & (g349) & (g362)));
	assign g364 = (((g108) & (g314) & (g317) & (g321) & (g328) & (g363)));
	assign g365 = (((g35) & (!g76) & (!sk[118]) & (!g1) & (!g40) & (!g201)) + ((g35) & (!g76) & (!sk[118]) & (!g1) & (!g40) & (g201)) + ((!g35) & (g76) & (!sk[118]) & (g1) & (!g40) & (!g201)) + ((!g35) & (!g76) & (!sk[118]) & (!g1) & (g40) & (g201)) + ((!g35) & (!g76) & (sk[118]) & (!g1) & (g40) & (!g201)));
	assign g366 = (((!sk[119]) & (i_9_) & (g116) & (!g63) & (!g161)) + ((!sk[119]) & (i_9_) & (g116) & (g63) & (!g161)) + ((!sk[119]) & (i_9_) & (!g116) & (!g63) & (g161)) + ((sk[119]) & (!i_9_) & (!g116) & (g63) & (g161)));
	assign g367 = (((g133) & (g64) & (!sk[120]) & (!g27) & (!g165)) + ((!g133) & (g64) & (sk[120]) & (g27) & (!g165)) + ((!g133) & (!g64) & (sk[120]) & (!g27) & (g165)) + ((g133) & (!g64) & (!sk[120]) & (!g27) & (g165)));
	assign g368 = (((!sk[121]) & (g38) & (!g307) & (!g354) & (g367)) + ((sk[121]) & (g38) & (!g307) & (!g354) & (!g367)) + ((sk[121]) & (!g38) & (!g307) & (!g354) & (!g367)) + ((!sk[121]) & (g38) & (g307) & (!g354) & (!g367)));
	assign g369 = (((!g35) & (g43) & (!g169) & (g58) & (!g71) & (!g171)) + ((!g35) & (!g43) & (!g169) & (g58) & (!g71) & (!g171)) + ((!g35) & (g43) & (!g169) & (!g58) & (!g71) & (!g171)) + ((!g35) & (!g43) & (!g169) & (!g58) & (!g71) & (!g171)) + ((!g35) & (g43) & (!g169) & (g58) & (!g71) & (!g171)) + ((!g35) & (!g43) & (!g169) & (g58) & (!g71) & (!g171)) + ((!g35) & (g43) & (!g169) & (!g58) & (!g71) & (!g171)) + ((!g35) & (!g43) & (!g169) & (!g58) & (!g71) & (!g171)));
	assign g370 = (((g8) & (!g36) & (!g42) & (!g13) & (!sk[123]) & (!g183)) + ((g8) & (g36) & (!g42) & (!g13) & (!sk[123]) & (!g183)) + ((!g8) & (g36) & (g42) & (!g13) & (!sk[123]) & (!g183)) + ((!g8) & (!g36) & (g42) & (!g13) & (sk[123]) & (g183)) + ((!g8) & (!g36) & (!g42) & (g13) & (!sk[123]) & (g183)));
	assign g371 = (((g365) & (!g366) & (!g368) & (!sk[124]) & (!g369) & (!g370)) + ((!g365) & (g366) & (g368) & (!sk[124]) & (!g369) & (!g370)) + ((!g365) & (!g366) & (!g368) & (!sk[124]) & (g369) & (g370)) + ((!g365) & (!g366) & (g368) & (sk[124]) & (g369) & (!g370)));
	assign g372 = (((!sk[125]) & (g59) & (g10) & (!g58) & (!g371)) + ((!sk[125]) & (g59) & (!g10) & (!g58) & (g371)) + ((sk[125]) & (!g59) & (!g10) & (!g58) & (g371)) + ((!sk[125]) & (g59) & (g10) & (!g58) & (g371)) + ((!sk[125]) & (g59) & (!g10) & (g58) & (g371)));
	assign g373 = (((g49) & (!g7) & (!g3) & (!g21) & (!sk[126]) & (!g156)) + ((g49) & (g7) & (!g3) & (!g21) & (!sk[126]) & (!g156)) + ((!g49) & (g7) & (g3) & (!g21) & (!sk[126]) & (!g156)) + ((!g49) & (!g7) & (!g3) & (!g21) & (sk[126]) & (g156)) + ((!g49) & (!g7) & (!g3) & (g21) & (!sk[126]) & (g156)) + ((!g49) & (g7) & (!g3) & (!g21) & (sk[126]) & (g156)));
	assign g374 = (((!sk[127]) & (i_9_) & (g39) & (!g101) & (!g31)) + ((!sk[127]) & (i_9_) & (g39) & (g101) & (!g31)) + ((!sk[127]) & (i_9_) & (!g39) & (!g101) & (g31)) + ((sk[127]) & (!i_9_) & (g39) & (!g101) & (g31)));
	assign g375 = (((!g43) & (!g37) & (!sk[0]) & (g55)) + ((!g43) & (!g37) & (!sk[0]) & (g55)) + ((!g43) & (!g37) & (sk[0]) & (!g55)) + ((g43) & (g37) & (!sk[0]) & (!g55)));
	assign g376 = (((g76) & (!g73) & (!g11) & (!sk[1]) & (!g90) & (!g375)) + ((!g76) & (g73) & (g11) & (!sk[1]) & (!g90) & (!g375)) + ((!g76) & (!g73) & (!g11) & (!sk[1]) & (g90) & (g375)) + ((!g76) & (!g73) & (!g11) & (sk[1]) & (!g90) & (!g375)) + ((g76) & (!g73) & (!g11) & (!sk[1]) & (!g90) & (!g375)) + ((!g76) & (!g73) & (!g11) & (sk[1]) & (!g90) & (!g375)));
	assign g377 = (((g20) & (!g28) & (!g25) & (!sk[2]) & (!g10) & (!g137)) + ((g20) & (!g28) & (g25) & (!sk[2]) & (!g10) & (!g137)) + ((!g20) & (g28) & (g25) & (!sk[2]) & (!g10) & (!g137)) + ((!g20) & (!g28) & (!g25) & (!sk[2]) & (g10) & (g137)) + ((!g20) & (!g28) & (g25) & (sk[2]) & (!g10) & (g137)));
	assign g378 = (((!g35) & (!g165) & (!sk[3]) & (g377)) + ((g35) & (g165) & (!sk[3]) & (!g377)) + ((!g35) & (!g165) & (sk[3]) & (!g377)) + ((!g35) & (!g165) & (sk[3]) & (!g377)));
	assign g379 = (((!g2) & (!sk[4]) & (!g77) & (g115)) + ((g2) & (!sk[4]) & (g77) & (!g115)) + ((!g2) & (sk[4]) & (!g77) & (!g115)) + ((!g2) & (sk[4]) & (!g77) & (!g115)));
	assign g380 = (((g24) & (!g374) & (!g376) & (!sk[5]) & (!g378) & (!g379)) + ((!g24) & (g374) & (g376) & (!sk[5]) & (!g378) & (!g379)) + ((!g24) & (!g374) & (!g376) & (!sk[5]) & (g378) & (g379)) + ((!g24) & (!g374) & (g376) & (!sk[5]) & (g378) & (g379)));
	assign g381 = (((i_2_) & (!i_0_) & (!i_9_) & (!sk[6]) & (!g373) & (!g380)) + ((!i_2_) & (i_0_) & (i_9_) & (!sk[6]) & (!g373) & (!g380)) + ((!i_2_) & (!i_0_) & (!i_9_) & (sk[6]) & (!g373) & (g380)) + ((!i_2_) & (!i_0_) & (i_9_) & (sk[6]) & (!g373) & (g380)) + ((!i_2_) & (!i_0_) & (!i_9_) & (!sk[6]) & (g373) & (g380)) + ((!i_2_) & (!i_0_) & (!i_9_) & (sk[6]) & (!g373) & (g380)));
	assign g382 = (((i_9_) & (!g7) & (!g25) & (!g16) & (!sk[7]) & (!g157)) + ((!i_9_) & (g7) & (g25) & (!g16) & (!sk[7]) & (!g157)) + ((i_9_) & (!g7) & (g25) & (!g16) & (!sk[7]) & (g157)) + ((!i_9_) & (!g7) & (!g25) & (g16) & (!sk[7]) & (g157)) + ((!i_9_) & (g7) & (g25) & (g16) & (!sk[7]) & (!g157)));
	assign g383 = (((g42) & (!g21) & (!g32) & (!g135) & (!sk[8]) & (!g244)) + ((!g42) & (!g21) & (!g32) & (!g135) & (sk[8]) & (!g244)) + ((!g42) & (!g21) & (!g32) & (g135) & (!sk[8]) & (g244)) + ((!g42) & (g21) & (g32) & (!g135) & (!sk[8]) & (!g244)) + ((!g42) & (g21) & (!g32) & (!g135) & (sk[8]) & (!g244)) + ((!g42) & (!g21) & (!g32) & (!g135) & (sk[8]) & (!g244)));
	assign g384 = (((i_9_) & (g16) & (g124) & (!g59) & (!g1) & (!g14)) + ((!i_9_) & (g16) & (!g124) & (g59) & (!g1) & (!g14)) + ((i_9_) & (g16) & (!g124) & (!g59) & (!g1) & (!g14)));
	assign g385 = (((g22) & (!g7) & (!sk[10]) & (!g221) & (!g14) & (!g53)) + ((!g22) & (g7) & (!sk[10]) & (g221) & (!g14) & (!g53)) + ((g22) & (g7) & (!sk[10]) & (!g221) & (!g14) & (g53)) + ((!g22) & (!g7) & (sk[10]) & (g221) & (!g14) & (g53)) + ((!g22) & (!g7) & (!sk[10]) & (!g221) & (g14) & (g53)) + ((g22) & (!g7) & (!sk[10]) & (!g221) & (!g14) & (g53)));
	assign g386 = (((i_9_) & (!sk[11]) & (!i_8_) & (!g68) & (!g28) & (!g63)) + ((!i_9_) & (!sk[11]) & (i_8_) & (g68) & (!g28) & (!g63)) + ((!i_9_) & (!sk[11]) & (!i_8_) & (!g68) & (g28) & (g63)) + ((i_9_) & (!sk[11]) & (i_8_) & (g68) & (!g28) & (g63)) + ((!i_9_) & (sk[11]) & (!i_8_) & (g68) & (!g28) & (g63)));
	assign g387 = (((g20) & (g84) & (!g62) & (!sk[12]) & (!g386)) + ((g20) & (!g84) & (!g62) & (!sk[12]) & (g386)) + ((!g20) & (!g84) & (!g62) & (sk[12]) & (!g386)) + ((!g20) & (!g84) & (!g62) & (sk[12]) & (!g386)));
	assign g388 = (((!g49) & (!g117) & (!g134) & (!g2) & (!g179) & (!g171)) + ((!g49) & (!g117) & (!g134) & (!g2) & (!g179) & (!g171)) + ((!g49) & (!g117) & (!g134) & (!g2) & (!g179) & (!g171)) + ((!g49) & (!g117) & (!g134) & (!g2) & (!g179) & (!g171)));
	assign g389 = (((g22) & (!sk[14]) & (!g20) & (!g10) & (!g40) & (!g307)) + ((!g22) & (!sk[14]) & (!g20) & (!g10) & (g40) & (g307)) + ((!g22) & (!sk[14]) & (g20) & (g10) & (!g40) & (!g307)) + ((g22) & (!sk[14]) & (g20) & (!g10) & (!g40) & (!g307)));
	assign g390 = (((!sk[15]) & (!g40) & (!g144) & (g389)) + ((!sk[15]) & (g40) & (g144) & (!g389)) + ((sk[15]) & (!g40) & (!g144) & (!g389)) + ((sk[15]) & (!g40) & (!g144) & (!g389)));
	assign g391 = (((g383) & (!g384) & (!g385) & (g387) & (g388) & (g390)));
	assign g392 = (((!g133) & (!sk[17]) & (!g5) & (g80)) + ((!g133) & (sk[17]) & (!g5) & (!g80)) + ((g133) & (!sk[17]) & (g5) & (!g80)));
	assign g393 = (((i_2_) & (!i_0_) & (!i_1_) & (!g4) & (!sk[18]) & (!g137)) + ((!i_2_) & (i_0_) & (i_1_) & (!g4) & (!sk[18]) & (!g137)) + ((!i_2_) & (!i_0_) & (!i_1_) & (g4) & (!sk[18]) & (g137)) + ((!i_2_) & (!i_0_) & (!i_1_) & (!g4) & (sk[18]) & (!g137)) + ((i_2_) & (i_0_) & (!i_1_) & (!g4) & (!sk[18]) & (g137)));
	assign g394 = (((i_9_) & (!sk[19]) & (i_8_) & (!i_6_) & (!g393)) + ((i_9_) & (!sk[19]) & (!i_8_) & (!i_6_) & (g393)) + ((i_9_) & (!sk[19]) & (!i_8_) & (!i_6_) & (g393)));
	assign g395 = (((g7) & (!g38) & (!g39) & (!sk[20]) & (!g43) & (!g156)) + ((g7) & (!g38) & (g39) & (!sk[20]) & (!g43) & (!g156)) + ((!g7) & (g38) & (g39) & (!sk[20]) & (!g43) & (!g156)) + ((!g7) & (!g38) & (!g39) & (!sk[20]) & (g43) & (g156)) + ((!g7) & (!g38) & (!g39) & (sk[20]) & (!g43) & (g156)));
	assign g396 = (((g28) & (!g2) & (!sk[21]) & (!g18) & (g395)) + ((!g28) & (!g2) & (sk[21]) & (!g18) & (!g395)) + ((!g28) & (!g2) & (sk[21]) & (!g18) & (!g395)) + ((g28) & (g2) & (!sk[21]) & (!g18) & (!g395)));
	assign g397 = (((g25) & (!sk[22]) & (g40) & (!g394) & (!g396)) + ((g25) & (!sk[22]) & (!g40) & (!g394) & (g396)) + ((!g25) & (sk[22]) & (!g40) & (!g394) & (g396)) + ((!g25) & (sk[22]) & (!g40) & (!g394) & (g396)));
	assign g398 = (((i_9_) & (!g54) & (!sk[23]) & (!g45) & (!g60) & (!g240)) + ((!i_9_) & (g54) & (!sk[23]) & (g45) & (!g60) & (!g240)) + ((i_9_) & (!g54) & (!sk[23]) & (!g45) & (!g60) & (g240)) + ((!i_9_) & (!g54) & (!sk[23]) & (!g45) & (g60) & (g240)) + ((!i_9_) & (!g54) & (sk[23]) & (!g45) & (g60) & (!g240)));
	assign g399 = (((g22) & (!i_9_) & (!g50) & (!g76) & (!sk[24]) & (!g156)) + ((!g22) & (i_9_) & (g50) & (!g76) & (!sk[24]) & (!g156)) + ((g22) & (!i_9_) & (!g50) & (!g76) & (!sk[24]) & (g156)) + ((!g22) & (!i_9_) & (!g50) & (g76) & (!sk[24]) & (g156)) + ((g22) & (i_9_) & (!g50) & (!g76) & (!sk[24]) & (!g156)));
	assign g400 = (((i_9_) & (!g6) & (!g3) & (!sk[25]) & (!g30) & (!g179)) + ((!i_9_) & (g6) & (g3) & (!sk[25]) & (!g30) & (!g179)) + ((!i_9_) & (!g6) & (!g3) & (!sk[25]) & (g30) & (g179)) + ((i_9_) & (!g6) & (!g3) & (!sk[25]) & (g30) & (!g179)) + ((!i_9_) & (!g6) & (!g3) & (sk[25]) & (!g30) & (g179)));
	assign g401 = (((i_2_) & (!sk[26]) & (i_9_) & (!g7) & (!g16)) + ((!i_2_) & (sk[26]) & (!i_9_) & (!g7) & (g16)) + ((i_2_) & (!sk[26]) & (!i_9_) & (g7) & (g16)) + ((i_2_) & (!sk[26]) & (!i_9_) & (!g7) & (g16)));
	assign g402 = (((i_2_) & (!i_9_) & (!g119) & (!g10) & (!sk[27]) & (!g401)) + ((!i_2_) & (i_9_) & (g119) & (!g10) & (!sk[27]) & (!g401)) + ((!i_2_) & (!i_9_) & (!g119) & (g10) & (!sk[27]) & (g401)) + ((!i_2_) & (!i_9_) & (!g119) & (!g10) & (sk[27]) & (g401)) + ((!i_2_) & (i_9_) & (!g119) & (!g10) & (sk[27]) & (g401)));
	assign g403 = (((!g28) & (!sk[28]) & (!g18) & (g21)) + ((g28) & (!sk[28]) & (g18) & (!g21)) + ((!g28) & (sk[28]) & (g18) & (!g21)));
	assign g404 = (((!sk[29]) & (g133) & (!g53) & (!g46) & (!g224) & (!g403)) + ((!sk[29]) & (!g133) & (g53) & (g46) & (!g224) & (!g403)) + ((!sk[29]) & (!g133) & (!g53) & (!g46) & (g224) & (g403)) + ((!sk[29]) & (g133) & (!g53) & (!g46) & (!g224) & (!g403)) + ((!sk[29]) & (g133) & (!g53) & (!g46) & (!g224) & (!g403)) + ((sk[29]) & (!g133) & (!g53) & (!g46) & (!g224) & (!g403)) + ((sk[29]) & (!g133) & (!g53) & (!g46) & (!g224) & (!g403)));
	assign g405 = (((g398) & (!sk[30]) & (!g399) & (!g400) & (!g402) & (!g404)) + ((!g398) & (!sk[30]) & (g399) & (g400) & (!g402) & (!g404)) + ((!g398) & (!sk[30]) & (!g399) & (!g400) & (g402) & (g404)) + ((!g398) & (sk[30]) & (!g399) & (!g400) & (!g402) & (g404)));
	assign g406 = (((i_9_) & (!g25) & (!g5) & (!g148) & (!sk[31]) & (!g405)) + ((!i_9_) & (g25) & (g5) & (!g148) & (!sk[31]) & (!g405)) + ((i_9_) & (!g25) & (!g5) & (!g148) & (!sk[31]) & (g405)) + ((!i_9_) & (!g25) & (!g5) & (g148) & (!sk[31]) & (g405)) + ((!i_9_) & (!g25) & (!g5) & (!g148) & (sk[31]) & (g405)) + ((!i_9_) & (!g25) & (!g5) & (!g148) & (sk[31]) & (g405)));
	assign g407 = (((!sk[32]) & (i_9_) & (g59) & (!g37) & (!g19)) + ((!sk[32]) & (i_9_) & (!g59) & (!g37) & (g19)) + ((!sk[32]) & (i_9_) & (g59) & (!g37) & (g19)) + ((sk[32]) & (!i_9_) & (g59) & (!g37) & (!g19)));
	assign g408 = (((i_9_) & (!g39) & (!g76) & (!g3) & (!sk[33]) & (!g209)) + ((!i_9_) & (g39) & (g76) & (!g3) & (!sk[33]) & (!g209)) + ((i_9_) & (g39) & (!g76) & (!g3) & (!sk[33]) & (g209)) + ((!i_9_) & (!g39) & (!g76) & (g3) & (!sk[33]) & (g209)) + ((!i_9_) & (g39) & (!g76) & (!g3) & (sk[33]) & (!g209)));
	assign g409 = (((!sk[34]) & (i_9_) & (!i_5_) & (!g6) & (!g45) & (!g11)) + ((!sk[34]) & (!i_9_) & (i_5_) & (g6) & (!g45) & (!g11)) + ((!sk[34]) & (!i_9_) & (!i_5_) & (!g6) & (g45) & (g11)) + ((!sk[34]) & (i_9_) & (i_5_) & (!g6) & (!g45) & (g11)) + ((sk[34]) & (!i_9_) & (!i_5_) & (!g6) & (!g45) & (!g11)));
	assign g410 = (((i_3_) & (!sk[35]) & (!i_4_) & (!g407) & (!g408) & (!g409)) + ((!i_3_) & (!sk[35]) & (i_4_) & (g407) & (!g408) & (!g409)) + ((!i_3_) & (!sk[35]) & (!i_4_) & (!g407) & (g408) & (g409)) + ((!i_3_) & (sk[35]) & (!i_4_) & (!g407) & (!g408) & (!g409)) + ((!i_3_) & (sk[35]) & (i_4_) & (!g407) & (!g408) & (!g409)) + ((!i_3_) & (sk[35]) & (!i_4_) & (!g407) & (!g408) & (!g409)));
	assign g411 = (((i_2_) & (!sk[36]) & (!i_9_) & (!g119) & (!g233) & (!g259)) + ((!i_2_) & (!sk[36]) & (i_9_) & (g119) & (!g233) & (!g259)) + ((!i_2_) & (!sk[36]) & (!i_9_) & (!g119) & (g233) & (g259)) + ((i_2_) & (!sk[36]) & (i_9_) & (!g119) & (g233) & (!g259)) + ((!i_2_) & (sk[36]) & (!i_9_) & (!g119) & (!g233) & (g259)));
	assign g412 = (((g7) & (!g63) & (!g13) & (!g27) & (!sk[37]) & (!g193)) + ((g7) & (g63) & (!g13) & (g27) & (!sk[37]) & (!g193)) + ((!g7) & (g63) & (g13) & (!g27) & (!sk[37]) & (!g193)) + ((!g7) & (!g63) & (!g13) & (!g27) & (sk[37]) & (g193)) + ((!g7) & (!g63) & (!g13) & (g27) & (!sk[37]) & (g193)));
	assign g413 = (((g22) & (!g28) & (!sk[38]) & (!g2) & (!g177) & (!g58)) + ((!g22) & (g28) & (!sk[38]) & (g2) & (!g177) & (!g58)) + ((!g22) & (!g28) & (sk[38]) & (g2) & (g177) & (!g58)) + ((!g22) & (!g28) & (!sk[38]) & (!g2) & (g177) & (g58)) + ((g22) & (!g28) & (!sk[38]) & (!g2) & (!g177) & (!g58)));
	assign g414 = (((g35) & (!sk[39]) & (!g85) & (!g411) & (!g412) & (!g413)) + ((!g35) & (!sk[39]) & (g85) & (g411) & (!g412) & (!g413)) + ((!g35) & (!sk[39]) & (!g85) & (!g411) & (g412) & (g413)) + ((!g35) & (sk[39]) & (!g85) & (!g411) & (!g412) & (!g413)) + ((!g35) & (sk[39]) & (!g85) & (!g411) & (!g412) & (!g413)));
	assign g415 = (((i_8_) & (!g7) & (!sk[40]) & (!g36) & (!g63) & (!g69)) + ((!i_8_) & (g7) & (!sk[40]) & (g36) & (!g63) & (!g69)) + ((!i_8_) & (!g7) & (!sk[40]) & (!g36) & (g63) & (g69)) + ((!i_8_) & (g7) & (!sk[40]) & (!g36) & (g63) & (g69)) + ((i_8_) & (!g7) & (!sk[40]) & (g36) & (g63) & (g69)));
	assign g416 = (((i_9_) & (!g39) & (!g76) & (!g16) & (!sk[41]) & (!g4)) + ((!i_9_) & (g39) & (g76) & (!g16) & (!sk[41]) & (!g4)) + ((!i_9_) & (!g39) & (!g76) & (g16) & (!sk[41]) & (g4)) + ((i_9_) & (g39) & (!g76) & (g16) & (!sk[41]) & (!g4)) + ((!i_9_) & (g39) & (!g76) & (g16) & (sk[41]) & (!g4)));
	assign g417 = (((g42) & (!sk[42]) & (g193) & (!g415) & (!g416)) + ((g42) & (!sk[42]) & (!g193) & (!g415) & (g416)) + ((!g42) & (sk[42]) & (!g193) & (!g415) & (!g416)) + ((!g42) & (sk[42]) & (!g193) & (!g415) & (!g416)));
	assign g418 = (((!g22) & (!i_9_) & (!g3) & (g63) & (!g10) & (!g31)) + ((g22) & (!i_9_) & (!g3) & (!g63) & (!g10) & (g31)));
	assign g419 = (((i_9_) & (!sk[44]) & (!i_6_) & (!g39) & (!g30) & (!g206)) + ((!i_9_) & (!sk[44]) & (i_6_) & (g39) & (!g30) & (!g206)) + ((!i_9_) & (!sk[44]) & (!i_6_) & (!g39) & (g30) & (g206)) + ((i_9_) & (!sk[44]) & (i_6_) & (g39) & (g30) & (g206)));
	assign g420 = (((!sk[45]) & (g20) & (!g13) & (!g161) & (!g112) & (!g208)) + ((sk[45]) & (!g20) & (!g13) & (!g161) & (!g112) & (!g208)) + ((!sk[45]) & (!g20) & (!g13) & (!g161) & (g112) & (g208)) + ((!sk[45]) & (!g20) & (g13) & (g161) & (!g112) & (!g208)) + ((!sk[45]) & (g20) & (g13) & (!g161) & (!g112) & (!g208)) + ((!sk[45]) & (g20) & (!g13) & (!g161) & (!g112) & (!g208)));
	assign g421 = (((g38) & (!g35) & (!g120) & (!g9) & (!sk[46]) & (!g57)) + ((g38) & (!g35) & (!g120) & (!g9) & (!sk[46]) & (!g57)) + ((g38) & (!g35) & (!g120) & (!g9) & (!sk[46]) & (!g57)) + ((!g38) & (g35) & (g120) & (!g9) & (!sk[46]) & (!g57)) + ((!g38) & (!g35) & (!g120) & (g9) & (!sk[46]) & (g57)) + ((!g38) & (!g35) & (!g120) & (!g9) & (sk[46]) & (!g57)) + ((!g38) & (!g35) & (!g120) & (!g9) & (sk[46]) & (!g57)));
	assign g422 = (((!sk[47]) & (g76) & (g3) & (!g4) & (!g45)) + ((sk[47]) & (!g76) & (!g3) & (!g4) & (!g45)) + ((!sk[47]) & (g76) & (!g3) & (!g4) & (g45)) + ((sk[47]) & (!g76) & (!g3) & (!g4) & (!g45)));
	assign g423 = (((!sk[48]) & (g122) & (g2) & (!g15) & (!g422)) + ((sk[48]) & (!g122) & (g2) & (g15) & (!g422)) + ((!sk[48]) & (g122) & (!g2) & (!g15) & (g422)) + ((sk[48]) & (!g122) & (g2) & (!g15) & (g422)));
	assign g424 = (((!sk[49]) & (!i_9_) & (!i_8_) & (i_7_)) + ((!sk[49]) & (i_9_) & (i_8_) & (!i_7_)) + ((!sk[49]) & (i_9_) & (i_8_) & (i_7_)));
	assign g425 = (((i_6_) & (i_5_) & (!i_3_) & (!i_4_) & (g25) & (g424)) + ((!i_6_) & (!i_5_) & (!i_3_) & (!i_4_) & (g25) & (g424)));
	assign g426 = (((!i_5_) & (!i_3_) & (!i_4_) & (g39) & (!g59) & (g40)) + ((i_5_) & (!i_3_) & (i_4_) & (!g39) & (g59) & (g40)));
	assign g427 = (((!sk[52]) & (g26) & (!g27) & (!g354) & (!g425) & (!g426)) + ((!sk[52]) & (!g26) & (g27) & (g354) & (!g425) & (!g426)) + ((!sk[52]) & (!g26) & (!g27) & (!g354) & (g425) & (g426)) + ((sk[52]) & (!g26) & (!g27) & (!g354) & (!g425) & (!g426)) + ((sk[52]) & (!g26) & (!g27) & (!g354) & (!g425) & (!g426)));
	assign g428 = (((g419) & (!g420) & (!g421) & (!g423) & (!sk[53]) & (!g427)) + ((!g419) & (g420) & (g421) & (!g423) & (!sk[53]) & (!g427)) + ((!g419) & (!g420) & (!g421) & (g423) & (!sk[53]) & (g427)) + ((!g419) & (g420) & (g421) & (!g423) & (!sk[53]) & (g427)));
	assign g429 = (((g255) & (!sk[54]) & (!g414) & (!g417) & (!g418) & (!g428)) + ((!g255) & (!sk[54]) & (g414) & (g417) & (!g418) & (!g428)) + ((!g255) & (!sk[54]) & (!g414) & (!g417) & (g418) & (g428)) + ((g255) & (!sk[54]) & (g414) & (g417) & (!g418) & (g428)));
	assign g430 = (((g392) & (g203) & (g397) & (g406) & (g410) & (g429)));
	assign g431 = (((g314) & (g372) & (g381) & (!g382) & (g391) & (g430)));
	assign g432 = (((i_2_) & (!sk[57]) & (!i_9_) & (!g272) & (!g157) & (!g233)) + ((!i_2_) & (!sk[57]) & (i_9_) & (g272) & (!g157) & (!g233)) + ((!i_2_) & (!sk[57]) & (!i_9_) & (!g272) & (g157) & (g233)) + ((i_2_) & (!sk[57]) & (i_9_) & (g272) & (!g157) & (g233)) + ((!i_2_) & (sk[57]) & (!i_9_) & (g272) & (g157) & (!g233)));
	assign g433 = (((i_9_) & (!g50) & (!sk[58]) & (!g7) & (!g6) & (!g221)) + ((!i_9_) & (g50) & (!sk[58]) & (g7) & (!g6) & (!g221)) + ((i_9_) & (!g50) & (!sk[58]) & (!g7) & (!g6) & (g221)) + ((!i_9_) & (!g50) & (!sk[58]) & (!g7) & (g6) & (g221)) + ((!i_9_) & (!g50) & (sk[58]) & (g7) & (!g6) & (!g221)));
	assign g434 = (((!sk[59]) & (g20) & (g240) & (!g432) & (!g433)) + ((!sk[59]) & (g20) & (!g240) & (!g432) & (g433)) + ((sk[59]) & (!g20) & (!g240) & (!g432) & (!g433)) + ((sk[59]) & (!g20) & (!g240) & (!g432) & (!g433)));
	assign g435 = (((i_9_) & (g8) & (!g28) & (!g63) & (g11) & (!g138)) + ((!i_9_) & (!g8) & (!g28) & (g63) & (!g11) & (g138)));
	assign g436 = (((i_2_) & (!g78) & (!g156) & (!sk[61]) & (!g31) & (!g151)) + ((!i_2_) & (g78) & (g156) & (!sk[61]) & (!g31) & (!g151)) + ((i_2_) & (!g78) & (!g156) & (!sk[61]) & (g31) & (g151)) + ((!i_2_) & (!g78) & (!g156) & (!sk[61]) & (g31) & (g151)) + ((!i_2_) & (g78) & (g156) & (!sk[61]) & (!g31) & (g151)));
	assign g437 = (((g22) & (!i_9_) & (g9) & (!g11) & (!g165) & (!g193)) + ((!g22) & (i_9_) & (!g9) & (g11) & (g165) & (!g193)) + ((g22) & (i_9_) & (!g9) & (!g11) & (!g165) & (g193)) + ((!g22) & (!i_9_) & (!g9) & (g11) & (!g165) & (g193)));
	assign g438 = (((i_9_) & (g25) & (!sk[63]) & (!g44) & (!g31)) + ((i_9_) & (g25) & (!sk[63]) & (!g44) & (g31)) + ((i_9_) & (!g25) & (!sk[63]) & (!g44) & (g31)) + ((!i_9_) & (g25) & (sk[63]) & (g44) & (!g31)));
	assign g439 = (((i_9_) & (!g54) & (!g59) & (!sk[64]) & (!g10) & (!g31)) + ((!i_9_) & (g54) & (g59) & (!sk[64]) & (!g10) & (!g31)) + ((!i_9_) & (!g54) & (!g59) & (!sk[64]) & (g10) & (g31)) + ((i_9_) & (!g54) & (g59) & (!sk[64]) & (!g10) & (!g31)) + ((!i_9_) & (!g54) & (g59) & (sk[64]) & (!g10) & (g31)));
	assign g440 = (((g25) & (!sk[65]) & (g76)) + ((g25) & (sk[65]) & (!g76)));
	assign g441 = (((!g20) & (!g53) & (!g27) & (!g12) & (!g208) & (!g440)) + ((!g20) & (!g53) & (!g27) & (g12) & (!g208) & (!g440)) + ((!g20) & (!g53) & (!g27) & (g12) & (!g208) & (!g440)) + ((!g20) & (!g53) & (!g27) & (g12) & (!g208) & (!g440)) + ((!g20) & (!g53) & (!g27) & (!g12) & (!g208) & (!g440)));
	assign g442 = (((g7) & (g42) & (!g3) & (!sk[67]) & (!g356)) + ((g7) & (g42) & (!g3) & (!sk[67]) & (!g356)) + ((!g7) & (g42) & (!g3) & (sk[67]) & (g356)) + ((g7) & (!g42) & (!g3) & (!sk[67]) & (g356)));
	assign g443 = (((!g120) & (!sk[68]) & (!g4) & (g45)) + ((!g120) & (!sk[68]) & (!g4) & (g45)) + ((!g120) & (sk[68]) & (g4) & (!g45)) + ((g120) & (!sk[68]) & (g4) & (!g45)));
	assign g444 = (((!sk[69]) & (g13) & (!g161) & (!g51) & (!g442) & (!g443)) + ((!sk[69]) & (g13) & (!g161) & (!g51) & (!g442) & (!g443)) + ((!sk[69]) & (!g13) & (g161) & (g51) & (!g442) & (!g443)) + ((!sk[69]) & (!g13) & (!g161) & (!g51) & (g442) & (g443)) + ((sk[69]) & (!g13) & (!g161) & (!g51) & (!g442) & (g443)));
	assign g445 = (((!sk[70]) & (g49) & (!i_5_) & (!i_3_) & (!i_4_) & (!g3)) + ((!sk[70]) & (!g49) & (i_5_) & (i_3_) & (!i_4_) & (!g3)) + ((!sk[70]) & (!g49) & (!i_5_) & (!i_3_) & (i_4_) & (g3)) + ((!sk[70]) & (g49) & (!i_5_) & (!i_3_) & (i_4_) & (!g3)) + ((!sk[70]) & (g49) & (i_5_) & (!i_3_) & (!i_4_) & (!g3)));
	assign g446 = (((g35) & (!sk[71]) & (g5) & (!g230) & (!g445)) + ((g35) & (!sk[71]) & (!g5) & (!g230) & (g445)) + ((!g35) & (sk[71]) & (!g5) & (!g230) & (!g445)) + ((!g35) & (sk[71]) & (!g5) & (!g230) & (!g445)));
	assign g447 = (((i_5_) & (!i_4_) & (!sk[72]) & (!g8) & (!g117) & (!g133)) + ((!i_5_) & (i_4_) & (!sk[72]) & (g8) & (!g117) & (!g133)) + ((!i_5_) & (!i_4_) & (!sk[72]) & (!g8) & (g117) & (g133)) + ((!i_5_) & (!i_4_) & (sk[72]) & (!g8) & (g117) & (!g133)) + ((!i_5_) & (i_4_) & (!sk[72]) & (g8) & (!g117) & (!g133)));
	assign g448 = (((g22) & (!g28) & (!g73) & (!g27) & (!sk[73]) & (!g90)) + ((!g22) & (!g28) & (!g73) & (g27) & (!sk[73]) & (g90)) + ((g22) & (!g28) & (g73) & (!g27) & (!sk[73]) & (!g90)) + ((!g22) & (g28) & (g73) & (!g27) & (!sk[73]) & (!g90)) + ((!g22) & (!g28) & (g73) & (!g27) & (sk[73]) & (g90)));
	assign g449 = (((g63) & (!g263) & (!g446) & (!sk[74]) & (!g447) & (!g448)) + ((!g63) & (g263) & (g446) & (!sk[74]) & (!g447) & (!g448)) + ((!g63) & (!g263) & (!g446) & (!sk[74]) & (g447) & (g448)) + ((!g63) & (!g263) & (g446) & (sk[74]) & (!g447) & (!g448)) + ((!g63) & (!g263) & (g446) & (sk[74]) & (!g447) & (!g448)));
	assign g450 = (((g438) & (!g439) & (!g441) & (!sk[75]) & (!g444) & (!g449)) + ((!g438) & (g439) & (g441) & (!sk[75]) & (!g444) & (!g449)) + ((!g438) & (!g439) & (!g441) & (!sk[75]) & (g444) & (g449)) + ((!g438) & (!g439) & (g441) & (!sk[75]) & (g444) & (g449)));
	assign g451 = (((!sk[76]) & (i_9_) & (i_3_) & (!i_4_) & (!g1)) + ((!sk[76]) & (i_9_) & (!i_3_) & (!i_4_) & (g1)) + ((sk[76]) & (!i_9_) & (i_3_) & (i_4_) & (!g1)) + ((sk[76]) & (i_9_) & (!i_3_) & (!i_4_) & (!g1)));
	assign g452 = (((i_9_) & (!g63) & (!sk[77]) & (!g11) & (!g51) & (!g32)) + ((!i_9_) & (g63) & (!sk[77]) & (g11) & (!g51) & (!g32)) + ((i_9_) & (g63) & (!sk[77]) & (!g11) & (!g51) & (g32)) + ((!i_9_) & (!g63) & (!sk[77]) & (!g11) & (g51) & (g32)) + ((!i_9_) & (!g63) & (sk[77]) & (g11) & (g51) & (!g32)));
	assign g453 = (((!g2) & (g21) & (!g40) & (!g64) & (!g15) & (!g165)) + ((!g2) & (g21) & (!g40) & (!g64) & (!g15) & (!g165)) + ((!g2) & (!g21) & (!g40) & (!g64) & (!g15) & (!g165)) + ((!g2) & (!g21) & (!g40) & (!g64) & (!g15) & (!g165)) + ((!g2) & (g21) & (!g40) & (!g64) & (!g15) & (!g165)) + ((!g2) & (g21) & (!g40) & (!g64) & (!g15) & (!g165)) + ((!g2) & (!g21) & (!g40) & (!g64) & (!g15) & (!g165)) + ((!g2) & (!g21) & (!g40) & (!g64) & (!g15) & (!g165)));
	assign g454 = (((g7) & (!g39) & (!g42) & (!g58) & (!sk[79]) & (!g209)) + ((g7) & (g39) & (!g42) & (!g58) & (!sk[79]) & (!g209)) + ((!g7) & (g39) & (g42) & (!g58) & (!sk[79]) & (!g209)) + ((!g7) & (!g39) & (g42) & (!g58) & (sk[79]) & (g209)) + ((!g7) & (!g39) & (!g42) & (g58) & (!sk[79]) & (g209)));
	assign g455 = (((g137) & (!sk[80]) & (!g302) & (!g452) & (!g453) & (!g454)) + ((!g137) & (!sk[80]) & (g302) & (g452) & (!g453) & (!g454)) + ((!g137) & (!sk[80]) & (!g302) & (!g452) & (g453) & (g454)) + ((!g137) & (sk[80]) & (!g302) & (!g452) & (g453) & (!g454)) + ((!g137) & (sk[80]) & (!g302) & (!g452) & (g453) & (!g454)));
	assign g456 = (((i_5_) & (!g54) & (g308) & (!g389) & (!g451) & (g455)) + ((!i_5_) & (g54) & (g308) & (!g389) & (!g451) & (g455)) + ((!i_5_) & (!g54) & (g308) & (!g389) & (!g451) & (g455)));
	assign g457 = (((!sk[82]) & (g73) & (g124) & (!g133) & (!g97)) + ((!sk[82]) & (g73) & (!g124) & (!g133) & (g97)) + ((sk[82]) & (!g73) & (!g124) & (!g133) & (g97)));
	assign g458 = (((i_9_) & (i_8_) & (!sk[83]) & (!i_6_) & (!i_7_)) + ((i_9_) & (!i_8_) & (!sk[83]) & (!i_6_) & (i_7_)) + ((i_9_) & (!i_8_) & (!sk[83]) & (i_6_) & (i_7_)) + ((i_9_) & (!i_8_) & (sk[83]) & (!i_6_) & (!i_7_)));
	assign g459 = (((i_5_) & (!i_3_) & (!i_4_) & (!g11) & (!sk[84]) & (!g40)) + ((!i_5_) & (i_3_) & (i_4_) & (!g11) & (!sk[84]) & (!g40)) + ((!i_5_) & (!i_3_) & (!i_4_) & (g11) & (!sk[84]) & (g40)) + ((!i_5_) & (!i_3_) & (!i_4_) & (g11) & (sk[84]) & (!g40)) + ((!i_5_) & (i_3_) & (i_4_) & (g11) & (!sk[84]) & (g40)));
	assign g460 = (((g4) & (g53) & (!g458) & (!sk[85]) & (!g459)) + ((g4) & (!g53) & (!g458) & (!sk[85]) & (g459)) + ((!g4) & (!g53) & (g458) & (sk[85]) & (g459)) + ((!g4) & (g53) & (g458) & (sk[85]) & (g459)));
	assign g461 = (((!sk[86]) & (g9) & (g21) & (!g169) & (!g32)) + ((sk[86]) & (g9) & (!g21) & (!g169) & (!g32)) + ((sk[86]) & (!g9) & (!g21) & (g169) & (!g32)) + ((sk[86]) & (!g9) & (!g21) & (!g169) & (g32)) + ((!sk[86]) & (g9) & (!g21) & (!g169) & (g32)));
	assign g462 = (((!g35) & (!g120) & (!g43) & (!g2) & (!g85) & (!g186)) + ((!g35) & (!g120) & (g43) & (!g2) & (!g85) & (!g186)) + ((!g35) & (!g120) & (!g43) & (!g2) & (!g85) & (!g186)) + ((!g35) & (!g120) & (g43) & (!g2) & (!g85) & (!g186)) + ((!g35) & (!g120) & (!g43) & (!g2) & (!g85) & (!g186)) + ((!g35) & (!g120) & (g43) & (!g2) & (!g85) & (!g186)) + ((!g35) & (!g120) & (!g43) & (!g2) & (!g85) & (!g186)) + ((!g35) & (!g120) & (g43) & (!g2) & (!g85) & (!g186)));
	assign g463 = (((!g49) & (!g38) & (!g76) & (!g3) & (!g138) & (g112)) + ((g49) & (!g38) & (!g76) & (!g3) & (!g138) & (!g112)) + ((g49) & (!g38) & (!g76) & (!g3) & (g138) & (!g112)));
	assign g464 = (((!sk[89]) & (g73) & (!g440) & (!g461) & (!g462) & (!g463)) + ((!sk[89]) & (!g73) & (g440) & (g461) & (!g462) & (!g463)) + ((!sk[89]) & (!g73) & (!g440) & (!g461) & (g462) & (g463)) + ((sk[89]) & (!g73) & (!g440) & (!g461) & (g462) & (!g463)) + ((!sk[89]) & (g73) & (!g440) & (!g461) & (g462) & (!g463)));
	assign g465 = (((i_9_) & (!i_8_) & (!sk[90]) & (!i_6_) & (!i_7_) & (!g76)) + ((!i_9_) & (i_8_) & (!sk[90]) & (i_6_) & (!i_7_) & (!g76)) + ((!i_9_) & (!i_8_) & (!sk[90]) & (!i_6_) & (i_7_) & (g76)) + ((i_9_) & (i_8_) & (!sk[90]) & (!i_6_) & (!i_7_) & (!g76)) + ((i_9_) & (i_8_) & (!sk[90]) & (i_6_) & (i_7_) & (!g76)));
	assign g466 = (((!sk[91]) & (i_5_) & (i_4_) & (!g11) & (!g465)) + ((!sk[91]) & (i_5_) & (!i_4_) & (!g11) & (g465)) + ((!sk[91]) & (i_5_) & (!i_4_) & (g11) & (g465)));
	assign g467 = (((!g30) & (!g58) & (!g457) & (!g460) & (g464) & (!g466)) + ((!g30) & (g58) & (!g457) & (!g460) & (g464) & (!g466)));
	assign g468 = (((g129) & (!g436) & (!g437) & (g450) & (g456) & (g467)));
	assign g469 = (((g20) & (!g73) & (!sk[94]) & (!g63) & (!g10) & (!g307)) + ((!g20) & (g73) & (!sk[94]) & (g63) & (!g10) & (!g307)) + ((g20) & (!g73) & (!sk[94]) & (g63) & (!g10) & (!g307)) + ((!g20) & (g73) & (sk[94]) & (!g63) & (!g10) & (g307)) + ((!g20) & (!g73) & (!sk[94]) & (!g63) & (g10) & (g307)) + ((!g20) & (!g73) & (sk[94]) & (g63) & (!g10) & (g307)));
	assign g470 = (((!i_2_) & (!i_9_) & (!g36) & (!g54) & (g75) & (g51)) + ((i_2_) & (i_9_) & (g36) & (!g54) & (g75) & (!g51)));
	assign g471 = (((!sk[96]) & (g117) & (g133) & (!g21) & (!g31)) + ((sk[96]) & (g117) & (!g133) & (!g21) & (!g31)) + ((sk[96]) & (!g117) & (!g133) & (!g21) & (g31)) + ((!sk[96]) & (g117) & (!g133) & (!g21) & (g31)));
	assign g472 = (((g49) & (g42) & (!sk[97]) & (!g211) & (!g225)) + ((g49) & (!g42) & (sk[97]) & (g211) & (!g225)) + ((!g49) & (g42) & (sk[97]) & (!g211) & (g225)) + ((g49) & (!g42) & (!sk[97]) & (!g211) & (g225)));
	assign g473 = (((g20) & (!sk[98]) & (!g208) & (!g470) & (!g471) & (!g472)) + ((!g20) & (!sk[98]) & (g208) & (g470) & (!g471) & (!g472)) + ((!g20) & (!sk[98]) & (!g208) & (!g470) & (g471) & (g472)) + ((!g20) & (sk[98]) & (!g208) & (!g470) & (!g471) & (!g472)) + ((!g20) & (sk[98]) & (!g208) & (!g470) & (!g471) & (!g472)));
	assign g474 = (((i_9_) & (!sk[99]) & (!i_8_) & (!i_6_) & (!g469) & (!g473)) + ((!i_9_) & (!sk[99]) & (i_8_) & (i_6_) & (!g469) & (!g473)) + ((!i_9_) & (sk[99]) & (!i_8_) & (!i_6_) & (!g469) & (g473)) + ((!i_9_) & (!sk[99]) & (i_8_) & (i_6_) & (!g469) & (g473)) + ((!i_9_) & (!sk[99]) & (!i_8_) & (!i_6_) & (g469) & (g473)) + ((!i_9_) & (sk[99]) & (!i_8_) & (!i_6_) & (!g469) & (g473)));
	assign g475 = (((!sk[100]) & (!g28) & (!g1) & (g40)) + ((!sk[100]) & (!g28) & (!g1) & (g40)) + ((!sk[100]) & (g28) & (g1) & (!g40)) + ((sk[100]) & (!g28) & (!g1) & (!g40)));
	assign g476 = (((g22) & (!g1) & (!sk[101]) & (!g53) & (g458)) + ((g22) & (g1) & (!sk[101]) & (!g53) & (!g458)) + ((!g22) & (!g1) & (sk[101]) & (g53) & (g458)));
	assign g477 = (((i_9_) & (!g28) & (!g63) & (!sk[102]) & (!g45) & (!g94)) + ((!i_9_) & (g28) & (g63) & (!sk[102]) & (!g45) & (!g94)) + ((!i_9_) & (!g28) & (!g63) & (!sk[102]) & (g45) & (g94)) + ((i_9_) & (!g28) & (g63) & (!sk[102]) & (!g45) & (!g94)) + ((!i_9_) & (!g28) & (!g63) & (sk[102]) & (!g45) & (g94)));
	assign g478 = (((g20) & (!g30) & (!g59) & (!sk[103]) & (!g120) & (!g2)) + ((!g20) & (!g30) & (!g59) & (!sk[103]) & (g120) & (g2)) + ((g20) & (g30) & (g59) & (!sk[103]) & (!g120) & (!g2)) + ((!g20) & (g30) & (g59) & (!sk[103]) & (!g120) & (!g2)));
	assign g479 = (((g475) & (g476) & (!sk[104]) & (!g477) & (!g478)) + ((g475) & (!g476) & (!sk[104]) & (!g477) & (g478)) + ((!g475) & (!g476) & (sk[104]) & (!g477) & (!g478)) + ((!g475) & (!g476) & (sk[104]) & (!g477) & (!g478)));
	assign g480 = (((i_2_) & (i_0_) & (!i_1_) & (!sk[105]) & (!i_9_)) + ((!i_2_) & (!i_0_) & (!i_1_) & (sk[105]) & (!i_9_)) + ((i_2_) & (!i_0_) & (!i_1_) & (!sk[105]) & (i_9_)) + ((!i_2_) & (!i_0_) & (!i_1_) & (sk[105]) & (i_9_)) + ((!i_2_) & (!i_0_) & (!i_1_) & (sk[105]) & (!i_9_)));
	assign g481 = (((i_2_) & (!g78) & (!i_9_) & (!sk[106]) & (!g201) & (!g228)) + ((!i_2_) & (g78) & (i_9_) & (!sk[106]) & (!g201) & (!g228)) + ((!i_2_) & (!g78) & (!i_9_) & (!sk[106]) & (g201) & (g228)) + ((i_2_) & (g78) & (!i_9_) & (!sk[106]) & (!g201) & (g228)) + ((!i_2_) & (g78) & (!i_9_) & (sk[106]) & (g201) & (!g228)));
	assign g482 = (((!sk[107]) & (g22) & (i_9_) & (!g15) & (!g251)) + ((!sk[107]) & (g22) & (!i_9_) & (!g15) & (g251)) + ((!sk[107]) & (g22) & (i_9_) & (!g15) & (g251)) + ((sk[107]) & (g22) & (!i_9_) & (g15) & (!g251)));
	assign g483 = (((g42) & (!sk[108]) & (!g73) & (!g74) & (g77)) + ((g42) & (!sk[108]) & (g73) & (!g74) & (!g77)) + ((!g42) & (sk[108]) & (g73) & (!g74) & (!g77)));
	assign g484 = (((g704) & (g481) & (!g482) & (!sk[109]) & (!g483)) + ((g704) & (!g481) & (!g482) & (!sk[109]) & (g483)) + ((g704) & (!g481) & (!g482) & (sk[109]) & (!g483)));
	assign g485 = (((g290) & (!sk[110]) & (g474) & (!g479) & (!g484)) + ((g290) & (!sk[110]) & (!g474) & (!g479) & (g484)) + ((g290) & (!sk[110]) & (g474) & (g479) & (g484)));
	assign g486 = (((g34) & (g336) & (g434) & (!g435) & (g468) & (g485)));
	assign g487 = (((i_2_) & (g36) & (!sk[112]) & (!g18) & (!g209)) + ((i_2_) & (g36) & (!sk[112]) & (g18) & (!g209)) + ((!i_2_) & (!g36) & (sk[112]) & (!g18) & (g209)) + ((i_2_) & (!g36) & (!sk[112]) & (!g18) & (g209)));
	assign g488 = (((!sk[113]) & (g78) & (!i_9_) & (!g16) & (!g29) & (!g487)) + ((!sk[113]) & (!g78) & (i_9_) & (g16) & (!g29) & (!g487)) + ((!sk[113]) & (!g78) & (i_9_) & (g16) & (g29) & (!g487)) + ((!sk[113]) & (g78) & (!i_9_) & (!g16) & (!g29) & (g487)) + ((!sk[113]) & (!g78) & (!i_9_) & (!g16) & (g29) & (g487)));
	assign g489 = (((g22) & (!g7) & (!g35) & (!g18) & (!sk[114]) & (!g53)) + ((!g22) & (g7) & (g35) & (g18) & (!sk[114]) & (!g53)) + ((!g22) & (g7) & (g35) & (!g18) & (!sk[114]) & (!g53)) + ((g22) & (g7) & (!g35) & (!g18) & (!sk[114]) & (g53)) + ((!g22) & (!g7) & (!g35) & (g18) & (!sk[114]) & (g53)));
	assign g490 = (((!sk[115]) & (g49) & (g134) & (!g5) & (!g306)) + ((!sk[115]) & (g49) & (!g134) & (!g5) & (g306)) + ((sk[115]) & (!g49) & (!g134) & (!g5) & (!g306)) + ((sk[115]) & (!g49) & (!g134) & (!g5) & (!g306)));
	assign g491 = (((g38) & (!sk[116]) & (!g36) & (!g59) & (!g1) & (!g58)) + ((!g38) & (!sk[116]) & (!g36) & (!g59) & (g1) & (g58)) + ((!g38) & (!sk[116]) & (g36) & (g59) & (!g1) & (!g58)) + ((!g38) & (sk[116]) & (g36) & (!g59) & (!g1) & (!g58)) + ((!g38) & (!sk[116]) & (g36) & (g59) & (!g1) & (!g58)));
	assign g492 = (((!g25) & (g73) & (!g10) & (!g43) & (g82) & (!g211)) + ((!g25) & (!g73) & (!g10) & (!g43) & (!g82) & (g211)) + ((g25) & (g73) & (!g10) & (!g43) & (!g82) & (!g211)));
	assign g493 = (((g73) & (!g240) & (!sk[118]) & (!g490) & (!g491) & (!g492)) + ((!g73) & (g240) & (!sk[118]) & (g490) & (!g491) & (!g492)) + ((!g73) & (!g240) & (!sk[118]) & (!g490) & (g491) & (g492)) + ((!g73) & (!g240) & (sk[118]) & (g490) & (!g491) & (!g492)) + ((!g73) & (!g240) & (sk[118]) & (g490) & (!g491) & (!g492)));
	assign g494 = (((i_9_) & (g25) & (!g30) & (g120) & (!g138) & (!g208)) + ((i_9_) & (!g25) & (!g30) & (!g120) & (g138) & (g208)) + ((!i_9_) & (g25) & (g30) & (!g120) & (g138) & (!g208)));
	assign g495 = (((!sk[120]) & (g43) & (g58) & (!g148) & (!g222)) + ((sk[120]) & (!g43) & (!g58) & (g148) & (!g222)) + ((sk[120]) & (!g43) & (!g58) & (!g148) & (g222)) + ((!sk[120]) & (g43) & (!g58) & (!g148) & (g222)));
	assign g496 = (((g20) & (!g28) & (!sk[121]) & (!g1) & (!g40) & (!g62)) + ((!g20) & (!g28) & (!sk[121]) & (!g1) & (g40) & (g62)) + ((!g20) & (g28) & (!sk[121]) & (g1) & (!g40) & (!g62)) + ((g20) & (!g28) & (!sk[121]) & (!g1) & (!g40) & (!g62)));
	assign g497 = (((g118) & (!sk[122]) & (!g392) & (!g494) & (!g495) & (!g496)) + ((!g118) & (!sk[122]) & (g392) & (g494) & (!g495) & (!g496)) + ((!g118) & (!sk[122]) & (!g392) & (!g494) & (g495) & (g496)) + ((!g118) & (sk[122]) & (g392) & (!g494) & (!g495) & (!g496)));
	assign g498 = (((g295) & (!g488) & (!g489) & (!sk[123]) & (!g493) & (!g497)) + ((!g295) & (g488) & (g489) & (!sk[123]) & (!g493) & (!g497)) + ((!g295) & (!g488) & (!g489) & (!sk[123]) & (g493) & (g497)) + ((!g295) & (!g488) & (!g489) & (!sk[123]) & (g493) & (g497)));
	assign g499 = (((!i_9_) & (g59) & (!g45) & (!g11) & (g44) & (!g14)) + ((i_9_) & (!g59) & (!g45) & (g11) & (!g44) & (!g14)));
	assign g500 = (((!sk[125]) & (!g36) & (!g119) & (g18)) + ((!sk[125]) & (g36) & (g119) & (!g18)) + ((!sk[125]) & (g36) & (!g119) & (g18)));
	assign g501 = (((i_2_) & (!g7) & (!sk[126]) & (!g3) & (!g151) & (!g500)) + ((!i_2_) & (g7) & (!sk[126]) & (g3) & (!g151) & (!g500)) + ((!i_2_) & (!g7) & (!sk[126]) & (!g3) & (g151) & (g500)) + ((i_2_) & (g7) & (!sk[126]) & (!g3) & (g151) & (!g500)));
	assign g502 = (((g30) & (!g168) & (!g11) & (!sk[127]) & (!g2) & (!g53)) + ((!g30) & (g168) & (g11) & (!sk[127]) & (!g2) & (!g53)) + ((!g30) & (g168) & (!g11) & (sk[127]) & (g2) & (!g53)) + ((g30) & (!g168) & (g11) & (!sk[127]) & (!g2) & (g53)) + ((!g30) & (!g168) & (!g11) & (!sk[127]) & (g2) & (g53)));
	assign g503 = (((!sk[0]) & (g279) & (g499) & (!g501) & (!g502)) + ((!sk[0]) & (g279) & (!g499) & (!g501) & (g502)) + ((sk[0]) & (!g279) & (!g499) & (!g501) & (!g502)));
	assign g504 = (((i_9_) & (!i_8_) & (!sk[1]) & (!g81) & (!g23) & (!g440)) + ((!i_9_) & (i_8_) & (!sk[1]) & (g81) & (!g23) & (!g440)) + ((!i_9_) & (!i_8_) & (!sk[1]) & (!g81) & (g23) & (g440)) + ((i_9_) & (i_8_) & (!sk[1]) & (g81) & (g23) & (!g440)) + ((i_9_) & (!i_8_) & (!sk[1]) & (g81) & (!g23) & (g440)));
	assign g505 = (((g42) & (g133) & (!sk[2]) & (!g141) & (!g171)) + ((g42) & (!g133) & (sk[2]) & (g141) & (!g171)) + ((!g42) & (!g133) & (sk[2]) & (!g141) & (g171)) + ((g42) & (!g133) & (!sk[2]) & (!g141) & (g171)));
	assign g506 = (((i_9_) & (!sk[3]) & (!g50) & (!g28) & (!g11) & (!g14)) + ((!i_9_) & (!sk[3]) & (g50) & (g28) & (!g11) & (!g14)) + ((!i_9_) & (!sk[3]) & (!g50) & (!g28) & (g11) & (g14)) + ((i_9_) & (!sk[3]) & (!g50) & (!g28) & (g11) & (!g14)) + ((!i_9_) & (sk[3]) & (!g50) & (!g28) & (g11) & (!g14)));
	assign g507 = (((g58) & (!g90) & (!g504) & (!g505) & (!sk[4]) & (!g506)) + ((!g58) & (g90) & (g504) & (!g505) & (!sk[4]) & (!g506)) + ((!g58) & (!g90) & (!g504) & (g505) & (!sk[4]) & (g506)) + ((g58) & (!g90) & (!g504) & (!g505) & (!sk[4]) & (!g506)) + ((!g58) & (!g90) & (!g504) & (!g505) & (sk[4]) & (!g506)));
	assign g508 = (((i_9_) & (!g50) & (!sk[5]) & (!g7) & (!g75) & (!g74)) + ((!i_9_) & (g50) & (!sk[5]) & (g7) & (!g75) & (!g74)) + ((!i_9_) & (!g50) & (!sk[5]) & (!g7) & (g75) & (g74)) + ((i_9_) & (!g50) & (!sk[5]) & (!g7) & (!g75) & (!g74)) + ((!i_9_) & (!g50) & (sk[5]) & (g7) & (g75) & (!g74)));
	assign g509 = (((g1) & (!sk[6]) & (!g14) & (!g27) & (g508)) + ((g1) & (sk[6]) & (!g14) & (!g27) & (!g508)) + ((!g1) & (sk[6]) & (g14) & (!g27) & (!g508)) + ((!g1) & (sk[6]) & (!g14) & (!g27) & (!g508)) + ((g1) & (!sk[6]) & (g14) & (!g27) & (!g508)));
	assign g510 = (((g28) & (!sk[7]) & (!g25) & (!g73) & (g509)) + ((g28) & (!sk[7]) & (g25) & (!g73) & (!g509)) + ((!g28) & (sk[7]) & (!g25) & (!g73) & (g509)) + ((!g28) & (sk[7]) & (!g25) & (!g73) & (g509)));
	assign g511 = (((!i_9_) & (!i_6_) & (!sk[8]) & (g206)) + ((i_9_) & (i_6_) & (!sk[8]) & (!g206)));
	assign g512 = (((i_2_) & (i_0_) & (!i_1_) & (g7) & (!g38) & (g511)) + ((!i_2_) & (i_0_) & (i_1_) & (g7) & (!g38) & (g511)));
	assign g513 = (((!sk[10]) & (i_2_) & (!i_9_) & (!g272) & (!g141) & (!g244)) + ((!sk[10]) & (!i_2_) & (i_9_) & (g272) & (!g141) & (!g244)) + ((!sk[10]) & (!i_2_) & (!i_9_) & (!g272) & (g141) & (g244)) + ((!sk[10]) & (i_2_) & (!i_9_) & (g272) & (!g141) & (g244)) + ((sk[10]) & (!i_2_) & (!i_9_) & (g272) & (g141) & (!g244)));
	assign g514 = (((i_9_) & (!g39) & (!sk[11]) & (!g6) & (!g122) & (!g55)) + ((!i_9_) & (g39) & (!sk[11]) & (g6) & (!g122) & (!g55)) + ((i_9_) & (!g39) & (!sk[11]) & (!g6) & (!g122) & (g55)) + ((!i_9_) & (!g39) & (!sk[11]) & (!g6) & (g122) & (g55)) + ((!i_9_) & (g39) & (sk[11]) & (!g6) & (g122) & (!g55)));
	assign g515 = (((!sk[12]) & (!g25) & (!g4) & (g45)) + ((!sk[12]) & (g25) & (g4) & (!g45)) + ((sk[12]) & (g25) & (!g4) & (!g45)));
	assign g516 = (((i_9_) & (!g54) & (!g59) & (!g14) & (!sk[13]) & (!g515)) + ((!i_9_) & (g54) & (g59) & (!g14) & (!sk[13]) & (!g515)) + ((!i_9_) & (!g54) & (!g59) & (!g14) & (sk[13]) & (g515)) + ((i_9_) & (!g54) & (g59) & (!g14) & (!sk[13]) & (!g515)) + ((!i_9_) & (!g54) & (!g59) & (g14) & (!sk[13]) & (g515)));
	assign g517 = (((i_5_) & (!i_3_) & (!i_4_) & (!g8) & (!sk[14]) & (!g54)) + ((!i_5_) & (i_3_) & (i_4_) & (!g8) & (!sk[14]) & (!g54)) + ((!i_5_) & (!i_3_) & (!i_4_) & (g8) & (!sk[14]) & (g54)) + ((i_5_) & (!i_3_) & (i_4_) & (g8) & (!sk[14]) & (!g54)) + ((i_5_) & (i_3_) & (!i_4_) & (g8) & (!sk[14]) & (!g54)) + ((i_5_) & (!i_3_) & (i_4_) & (!g8) & (!sk[14]) & (!g54)) + ((i_5_) & (i_3_) & (!i_4_) & (!g8) & (!sk[14]) & (!g54)));
	assign g518 = (((g22) & (!i_9_) & (!sk[15]) & (!g36) & (!g20) & (!g517)) + ((!g22) & (i_9_) & (!sk[15]) & (g36) & (!g20) & (!g517)) + ((!g22) & (!i_9_) & (!sk[15]) & (!g36) & (g20) & (g517)) + ((g22) & (i_9_) & (!sk[15]) & (g36) & (!g20) & (g517)) + ((g22) & (i_9_) & (!sk[15]) & (!g36) & (g20) & (g517)));
	assign g519 = (((g38) & (!g76) & (!g514) & (!g516) & (!sk[16]) & (!g518)) + ((!g38) & (g76) & (g514) & (!g516) & (!sk[16]) & (!g518)) + ((!g38) & (!g76) & (!g514) & (g516) & (!sk[16]) & (g518)) + ((g38) & (g76) & (!g514) & (!g516) & (!sk[16]) & (!g518)) + ((!g38) & (!g76) & (!g514) & (!g516) & (sk[16]) & (!g518)));
	assign g520 = (((g59) & (!sk[17]) & (!g58) & (!g512) & (!g513) & (!g519)) + ((!g59) & (!sk[17]) & (g58) & (g512) & (!g513) & (!g519)) + ((!g59) & (!sk[17]) & (!g58) & (!g512) & (g513) & (g519)) + ((!g59) & (sk[17]) & (!g58) & (!g512) & (!g513) & (g519)) + ((!g59) & (!sk[17]) & (g58) & (g512) & (!g513) & (g519)));
	assign g521 = (((!sk[18]) & (g49) & (i_3_) & (!i_4_) & (!g13)) + ((!sk[18]) & (g49) & (!i_3_) & (!i_4_) & (g13)) + ((sk[18]) & (g49) & (!i_3_) & (!i_4_) & (!g13)) + ((sk[18]) & (!g49) & (i_3_) & (i_4_) & (!g13)));
	assign g522 = (((g50) & (!g76) & (!sk[19]) & (!g13) & (!g46) & (!g157)) + ((!g50) & (g76) & (!sk[19]) & (g13) & (!g46) & (!g157)) + ((!g50) & (!g76) & (sk[19]) & (!g13) & (g46) & (!g157)) + ((!g50) & (!g76) & (sk[19]) & (!g13) & (!g46) & (g157)) + ((!g50) & (!g76) & (!sk[19]) & (!g13) & (g46) & (g157)) + ((!g50) & (!g76) & (sk[19]) & (!g13) & (!g46) & (!g157)));
	assign g523 = (((i_5_) & (g8) & (!g521) & (!sk[20]) & (!g522)) + ((i_5_) & (!g8) & (!g521) & (!sk[20]) & (g522)) + ((!i_5_) & (!g8) & (!g521) & (sk[20]) & (!g522)) + ((!i_5_) & (!g8) & (!g521) & (sk[20]) & (!g522)) + ((i_5_) & (g8) & (!g521) & (!sk[20]) & (!g522)));
	assign g524 = (((g22) & (!i_9_) & (i_5_) & (i_3_) & (i_4_) & (g138)) + ((g22) & (i_9_) & (i_5_) & (i_3_) & (!i_4_) & (g138)));
	assign g525 = (((g35) & (!sk[22]) & (g183) & (!g148) & (!g524)) + ((g35) & (!sk[22]) & (!g183) & (!g148) & (g524)) + ((!g35) & (sk[22]) & (!g183) & (!g148) & (!g524)) + ((!g35) & (sk[22]) & (!g183) & (!g148) & (!g524)));
	assign g526 = (((g22) & (!sk[23]) & (!i_9_) & (!g28) & (!g16) & (!g45)) + ((!g22) & (!sk[23]) & (i_9_) & (g28) & (!g16) & (!g45)) + ((!g22) & (!sk[23]) & (!i_9_) & (!g28) & (g16) & (g45)) + ((g22) & (!sk[23]) & (!i_9_) & (!g28) & (g16) & (!g45)) + ((g22) & (!sk[23]) & (i_9_) & (!g28) & (!g16) & (!g45)));
	assign g527 = (((!g120) & (g43) & (!g161) & (!g251) & (!g228) & (!g526)) + ((!g120) & (!g43) & (!g161) & (!g251) & (!g228) & (!g526)));
	assign g528 = (((!sk[25]) & (g168) & (!g21) & (!g55) & (!g356) & (!g103)) + ((!sk[25]) & (!g168) & (g21) & (g55) & (!g356) & (!g103)) + ((!sk[25]) & (!g168) & (!g21) & (!g55) & (g356) & (g103)) + ((sk[25]) & (!g168) & (g21) & (!g55) & (!g356) & (!g103)) + ((sk[25]) & (!g168) & (!g21) & (!g55) & (!g356) & (!g103)));
	assign g529 = (((i_9_) & (!sk[26]) & (!g59) & (!g1) & (!g244) & (!g263)) + ((!i_9_) & (!sk[26]) & (g59) & (g1) & (!g244) & (!g263)) + ((!i_9_) & (sk[26]) & (!g59) & (!g1) & (!g244) & (g263)) + ((!i_9_) & (!sk[26]) & (!g59) & (!g1) & (g244) & (g263)) + ((!i_9_) & (sk[26]) & (!g59) & (!g1) & (g244) & (!g263)) + ((!i_9_) & (!sk[26]) & (g59) & (g1) & (!g244) & (g263)));
	assign g530 = (((g16) & (!sk[27]) & (!g30) & (!g133) & (!g139) & (!g90)) + ((g16) & (!sk[27]) & (!g30) & (!g133) & (!g139) & (g90)) + ((!g16) & (!sk[27]) & (g30) & (g133) & (!g139) & (!g90)) + ((g16) & (!sk[27]) & (g30) & (!g133) & (!g139) & (!g90)) + ((!g16) & (sk[27]) & (!g30) & (!g133) & (g139) & (!g90)) + ((!g16) & (!sk[27]) & (!g30) & (!g133) & (g139) & (g90)));
	assign g531 = (((!g20) & (!g99) & (g527) & (g528) & (!g529) & (!g530)) + ((!g20) & (!g99) & (g527) & (g528) & (!g529) & (!g530)));
	assign g532 = (((i_9_) & (!i_8_) & (!i_6_) & (!g59) & (!sk[29]) & (!g14)) + ((!i_9_) & (i_8_) & (i_6_) & (!g59) & (!sk[29]) & (!g14)) + ((!i_9_) & (!i_8_) & (!i_6_) & (g59) & (!sk[29]) & (g14)) + ((i_9_) & (i_8_) & (i_6_) & (g59) & (!sk[29]) & (!g14)));
	assign g533 = (((g20) & (!g137) & (!g52) & (!g71) & (!sk[30]) & (!g532)) + ((!g20) & (g137) & (g52) & (!g71) & (!sk[30]) & (!g532)) + ((!g20) & (!g137) & (!g52) & (g71) & (!sk[30]) & (g532)) + ((!g20) & (!g137) & (!g52) & (!g71) & (sk[30]) & (!g532)) + ((!g20) & (!g137) & (!g52) & (!g71) & (sk[30]) & (!g532)) + ((!g20) & (!g137) & (!g52) & (!g71) & (sk[30]) & (!g532)) + ((!g20) & (!g137) & (!g52) & (!g71) & (sk[30]) & (!g532)));
	assign g534 = (((g22) & (!i_7_) & (!i_5_) & (!g92) & (!sk[31]) & (!g192)) + ((!g22) & (i_7_) & (i_5_) & (!g92) & (!sk[31]) & (!g192)) + ((!g22) & (!i_7_) & (!i_5_) & (g92) & (!sk[31]) & (g192)) + ((g22) & (!i_7_) & (i_5_) & (g92) & (!sk[31]) & (g192)) + ((g22) & (i_7_) & (!i_5_) & (g92) & (!sk[31]) & (g192)));
	assign g535 = (((!sk[32]) & (i_9_) & (!g6) & (!g165) & (!g193) & (!g534)) + ((!sk[32]) & (!i_9_) & (g6) & (g165) & (!g193) & (!g534)) + ((!sk[32]) & (!i_9_) & (!g6) & (!g165) & (g193) & (g534)) + ((!sk[32]) & (i_9_) & (!g6) & (!g165) & (!g193) & (!g534)) + ((sk[32]) & (!i_9_) & (!g6) & (!g165) & (!g193) & (!g534)) + ((sk[32]) & (!i_9_) & (g6) & (!g165) & (!g193) & (!g534)));
	assign g536 = (((!sk[33]) & (i_9_) & (!i_8_) & (!i_6_) & (!i_7_) & (!g119)) + ((!sk[33]) & (!i_9_) & (i_8_) & (i_6_) & (!i_7_) & (!g119)) + ((!sk[33]) & (!i_9_) & (!i_8_) & (!i_6_) & (i_7_) & (g119)) + ((!sk[33]) & (i_9_) & (i_8_) & (i_6_) & (!i_7_) & (!g119)) + ((!sk[33]) & (i_9_) & (!i_8_) & (!i_6_) & (!i_7_) & (!g119)));
	assign g537 = (((i_2_) & (g7) & (g75) & (g73) & (!g14) & (!g40)) + ((!i_2_) & (!g7) & (g75) & (g73) & (!g14) & (!g40)) + ((!i_2_) & (g7) & (g75) & (!g73) & (!g14) & (g40)));
	assign g538 = (((g27) & (!g29) & (!sk[35]) & (!g475) & (!g536) & (!g537)) + ((!g27) & (g29) & (!sk[35]) & (g475) & (!g536) & (!g537)) + ((!g27) & (!g29) & (!sk[35]) & (!g475) & (g536) & (g537)) + ((!g27) & (!g29) & (sk[35]) & (!g475) & (!g536) & (!g537)) + ((!g27) & (!g29) & (sk[35]) & (!g475) & (!g536) & (!g537)) + ((!g27) & (!g29) & (sk[35]) & (!g475) & (!g536) & (!g537)));
	assign g539 = (((g303) & (!g697) & (!g533) & (!g535) & (!sk[36]) & (!g538)) + ((!g303) & (g697) & (g533) & (!g535) & (!sk[36]) & (!g538)) + ((!g303) & (!g697) & (!g533) & (g535) & (!sk[36]) & (g538)) + ((!g303) & (g697) & (g533) & (g535) & (!sk[36]) & (g538)));
	assign g540 = (((g774) & (g114) & (g523) & (g525) & (g531) & (g539)));
	assign g541 = (((g227) & (g338) & (g434) & (g510) & (g520) & (g540)));
	assign g542 = (((g381) & (!sk[39]) & (!g498) & (!g503) & (!g507) & (!g541)) + ((!g381) & (!sk[39]) & (g498) & (g503) & (!g507) & (!g541)) + ((!g381) & (!sk[39]) & (!g498) & (!g503) & (g507) & (g541)) + ((g381) & (!sk[39]) & (g498) & (g503) & (g507) & (g541)));
	assign g543 = (((!sk[40]) & (g20) & (g52) & (!g58) & (!g302)) + ((sk[40]) & (!g20) & (!g52) & (!g58) & (!g302)) + ((!sk[40]) & (g20) & (!g52) & (!g58) & (g302)) + ((sk[40]) & (!g20) & (!g52) & (!g58) & (!g302)) + ((sk[40]) & (!g20) & (!g52) & (g58) & (!g302)));
	assign g544 = (((i_9_) & (!g6) & (!g46) & (!sk[41]) & (!g19) & (!g488)) + ((!i_9_) & (g6) & (g46) & (!sk[41]) & (!g19) & (!g488)) + ((!i_9_) & (!g6) & (!g46) & (!sk[41]) & (g19) & (g488)) + ((i_9_) & (!g6) & (!g46) & (!sk[41]) & (!g19) & (!g488)) + ((!i_9_) & (g6) & (!g46) & (sk[41]) & (!g19) & (!g488)) + ((!i_9_) & (!g6) & (!g46) & (sk[41]) & (!g19) & (!g488)));
	assign g545 = (((g220) & (!g339) & (!g424) & (!g543) & (!sk[42]) & (!g544)) + ((!g220) & (g339) & (g424) & (!g543) & (!sk[42]) & (!g544)) + ((!g220) & (!g339) & (!g424) & (g543) & (!sk[42]) & (g544)) + ((!g220) & (!g339) & (!g424) & (g543) & (!sk[42]) & (g544)) + ((!g220) & (!g339) & (!g424) & (!g543) & (sk[42]) & (g544)));
	assign g546 = (((i_0_) & (!sk[43]) & (i_1_) & (!g135) & (!g251)) + ((i_0_) & (!sk[43]) & (!i_1_) & (!g135) & (g251)) + ((i_0_) & (!sk[43]) & (i_1_) & (!g135) & (g251)) + ((!i_0_) & (sk[43]) & (i_1_) & (g135) & (!g251)));
	assign g547 = (((i_2_) & (!sk[44]) & (!i_9_) & (!g546) & (g690)) + ((i_2_) & (!sk[44]) & (i_9_) & (!g546) & (!g690)) + ((!i_2_) & (sk[44]) & (i_9_) & (!g546) & (g690)) + ((!i_2_) & (sk[44]) & (!i_9_) & (!g546) & (g690)));
	assign g548 = (((!sk[45]) & (i_8_) & (g36) & (!g68) & (!g59)) + ((sk[45]) & (!i_8_) & (!g36) & (!g68) & (!g59)) + ((sk[45]) & (!i_8_) & (!g36) & (!g68) & (!g59)) + ((!sk[45]) & (i_8_) & (!g36) & (!g68) & (g59)) + ((sk[45]) & (!i_8_) & (!g36) & (!g68) & (!g59)));
	assign g549 = (((g22) & (!i_9_) & (!i_8_) & (!g83) & (!sk[46]) & (!g10)) + ((!g22) & (i_9_) & (!i_8_) & (!g83) & (sk[46]) & (!g10)) + ((!g22) & (i_9_) & (i_8_) & (!g83) & (!sk[46]) & (!g10)) + ((!g22) & (!i_9_) & (!i_8_) & (g83) & (!sk[46]) & (g10)) + ((g22) & (i_9_) & (!i_8_) & (g83) & (!sk[46]) & (!g10)));
	assign g550 = (((!i_9_) & (!sk[47]) & (!i_6_) & (i_7_)) + ((i_9_) & (!sk[47]) & (i_6_) & (!i_7_)) + ((i_9_) & (sk[47]) & (!i_6_) & (!i_7_)));
	assign g551 = (((!sk[48]) & (i_8_) & (!g39) & (!g30) & (!g71) & (!g550)) + ((!sk[48]) & (!i_8_) & (g39) & (g30) & (!g71) & (!g550)) + ((!sk[48]) & (!i_8_) & (!g39) & (!g30) & (g71) & (g550)) + ((!sk[48]) & (i_8_) & (!g39) & (!g30) & (g71) & (g550)) + ((!sk[48]) & (!i_8_) & (g39) & (g30) & (!g71) & (g550)));
	assign g552 = (((!i_9_) & (!g38) & (!g30) & (!g59) & (g94) & (!g46)) + ((!i_9_) & (!g38) & (g30) & (g59) & (!g94) & (!g46)) + ((!i_9_) & (!g38) & (!g30) & (g59) & (!g94) & (g46)));
	assign g553 = (((g49) & (!g35) & (!g116) & (!g135) & (!sk[50]) & (!g259)) + ((!g49) & (!g35) & (!g116) & (!g135) & (sk[50]) & (!g259)) + ((!g49) & (g35) & (g116) & (!g135) & (!sk[50]) & (!g259)) + ((!g49) & (!g35) & (!g116) & (g135) & (!sk[50]) & (g259)) + ((!g49) & (!g35) & (!g116) & (!g135) & (sk[50]) & (!g259)) + ((!g49) & (!g35) & (!g116) & (!g135) & (sk[50]) & (!g259)) + ((!g49) & (!g35) & (!g116) & (!g135) & (sk[50]) & (!g259)));
	assign g554 = (((!i_9_) & (!g50) & (!g28) & (!g63) & (g11) & (g182)) + ((i_9_) & (!g50) & (!g28) & (g63) & (!g11) & (!g182)) + ((i_9_) & (!g50) & (!g28) & (!g63) & (g11) & (!g182)));
	assign g555 = (((g101) & (g42) & (!g209) & (!sk[52]) & (!g148)) + ((!g101) & (g42) & (g209) & (sk[52]) & (!g148)) + ((!g101) & (g42) & (!g209) & (sk[52]) & (g148)) + ((g101) & (!g42) & (!g209) & (!sk[52]) & (g148)));
	assign g556 = (((g268) & (!sk[53]) & (g553) & (!g554) & (!g555)) + ((g268) & (!sk[53]) & (!g553) & (!g554) & (g555)) + ((!g268) & (sk[53]) & (g553) & (!g554) & (!g555)));
	assign g557 = (((g548) & (!g549) & (!g551) & (!g552) & (!sk[54]) & (!g556)) + ((!g548) & (g549) & (g551) & (!g552) & (!sk[54]) & (!g556)) + ((!g548) & (!g549) & (!g551) & (g552) & (!sk[54]) & (g556)) + ((g548) & (!g549) & (!g551) & (!g552) & (!sk[54]) & (g556)) + ((!g548) & (!g549) & (!g551) & (!g552) & (sk[54]) & (g556)));
	assign g558 = (((i_9_) & (!sk[55]) & (!g50) & (!g7) & (!g45) & (!g11)) + ((!i_9_) & (!sk[55]) & (g50) & (g7) & (!g45) & (!g11)) + ((!i_9_) & (!sk[55]) & (!g50) & (!g7) & (g45) & (g11)) + ((i_9_) & (!sk[55]) & (!g50) & (g7) & (!g45) & (g11)) + ((!i_9_) & (sk[55]) & (!g50) & (g7) & (!g45) & (g11)));
	assign g559 = (((g43) & (!g37) & (!g230) & (!sk[56]) & (!g225) & (!g558)) + ((g43) & (!g37) & (!g230) & (!sk[56]) & (!g225) & (!g558)) + ((!g43) & (g37) & (g230) & (!sk[56]) & (!g225) & (!g558)) + ((!g43) & (!g37) & (!g230) & (!sk[56]) & (g225) & (g558)) + ((!g43) & (g37) & (!g230) & (sk[56]) & (!g225) & (!g558)));
	assign g560 = (((i_9_) & (g16) & (!sk[57]) & (!g138) & (!g112)) + ((i_9_) & (g16) & (!sk[57]) & (!g138) & (g112)) + ((i_9_) & (!g16) & (!sk[57]) & (!g138) & (g112)) + ((!i_9_) & (!g16) & (sk[57]) & (g138) & (g112)));
	assign g561 = (((g13) & (!g158) & (!g259) & (!sk[58]) & (g560)) + ((g13) & (!g158) & (!g259) & (sk[58]) & (!g560)) + ((!g13) & (!g158) & (!g259) & (sk[58]) & (!g560)) + ((g13) & (g158) & (!g259) & (!sk[58]) & (!g560)));
	assign g562 = (((i_2_) & (i_9_) & (g36) & (!sk[59]) & (!g76)) + ((i_2_) & (i_9_) & (!g36) & (!sk[59]) & (!g76)) + ((i_2_) & (!i_9_) & (!g36) & (!sk[59]) & (g76)) + ((!i_2_) & (!i_9_) & (!g36) & (sk[59]) & (!g76)));
	assign g563 = (((g54) & (!g10) & (!sk[60]) & (!g133) & (!g18) & (!g141)) + ((!g54) & (g10) & (!sk[60]) & (g133) & (!g18) & (!g141)) + ((!g54) & (!g10) & (sk[60]) & (!g133) & (!g18) & (g141)) + ((!g54) & (!g10) & (!sk[60]) & (!g133) & (g18) & (g141)) + ((!g54) & (!g10) & (sk[60]) & (!g133) & (!g18) & (!g141)) + ((!g54) & (!g10) & (sk[60]) & (!g133) & (g18) & (!g141)));
	assign g564 = (((g50) & (!g75) & (!sk[61]) & (!g562) & (g563)) + ((!g50) & (!g75) & (sk[61]) & (!g562) & (!g563)) + ((!g50) & (!g75) & (sk[61]) & (!g562) & (!g563)) + ((g50) & (g75) & (!sk[61]) & (!g562) & (!g563)));
	assign g565 = (((!g81) & (!g35) & (!g10) & (g2) & (g233) & (!g228)) + ((!g81) & (g35) & (!g10) & (!g2) & (!g233) & (g228)) + ((g81) & (!g35) & (!g10) & (g2) & (!g233) & (!g228)));
	assign g566 = (((i_9_) & (!i_8_) & (!sk[63]) & (!i_5_) & (!i_3_) & (!i_4_)) + ((!i_9_) & (i_8_) & (!sk[63]) & (i_5_) & (!i_3_) & (!i_4_)) + ((!i_9_) & (!i_8_) & (!sk[63]) & (!i_5_) & (i_3_) & (i_4_)) + ((i_9_) & (i_8_) & (!sk[63]) & (i_5_) & (i_3_) & (i_4_)) + ((i_9_) & (i_8_) & (!sk[63]) & (!i_5_) & (i_3_) & (!i_4_)));
	assign g567 = (((i_7_) & (!sk[64]) & (!g6) & (!g73) & (!g14) & (!g566)) + ((!i_7_) & (!sk[64]) & (g6) & (g73) & (!g14) & (!g566)) + ((!i_7_) & (!sk[64]) & (!g6) & (!g73) & (g14) & (g566)) + ((!i_7_) & (sk[64]) & (!g6) & (!g73) & (!g14) & (g566)) + ((!i_7_) & (!sk[64]) & (!g6) & (g73) & (g14) & (g566)));
	assign g568 = (((!i_2_) & (i_0_) & (!i_1_) & (!g28) & (g73) & (!g40)) + ((!i_2_) & (i_0_) & (i_1_) & (!g28) & (!g73) & (g40)) + ((!i_2_) & (!i_0_) & (!i_1_) & (!g28) & (!g73) & (g40)));
	assign g569 = (((g7) & (g27) & (!g567) & (!sk[66]) & (!g568)) + ((g7) & (!g27) & (!g567) & (!sk[66]) & (g568)) + ((!g7) & (!g27) & (!g567) & (sk[66]) & (!g568)) + ((!g7) & (!g27) & (!g567) & (sk[66]) & (!g568)));
	assign g570 = (((g559) & (!g561) & (!sk[67]) & (!g564) & (!g565) & (!g569)) + ((!g559) & (g561) & (!sk[67]) & (g564) & (!g565) & (!g569)) + ((!g559) & (!g561) & (!sk[67]) & (!g564) & (g565) & (g569)) + ((g559) & (g561) & (!sk[67]) & (g564) & (!g565) & (g569)));
	assign g571 = (((i_9_) & (!sk[68]) & (i_8_) & (!g81) & (!g124)) + ((i_9_) & (!sk[68]) & (!i_8_) & (!g81) & (g124)) + ((i_9_) & (!sk[68]) & (!i_8_) & (g81) & (g124)) + ((!i_9_) & (sk[68]) & (i_8_) & (g81) & (g124)));
	assign g572 = (((g39) & (g20) & (!g10) & (!g14) & (!g58) & (g424)) + ((g39) & (!g20) & (!g10) & (!g14) & (!g58) & (g424)) + ((g39) & (!g20) & (!g10) & (!g14) & (!g58) & (g424)));
	assign g573 = (((g49) & (g32) & (!g157) & (!sk[70]) & (!g251)) + ((g49) & (!g32) & (!g157) & (!sk[70]) & (g251)) + ((g49) & (!g32) & (g157) & (sk[70]) & (!g251)));
	assign g574 = (((g460) & (!g464) & (!g571) & (!g572) & (!sk[71]) & (!g573)) + ((!g460) & (g464) & (g571) & (!g572) & (!sk[71]) & (!g573)) + ((!g460) & (!g464) & (!g571) & (g572) & (!sk[71]) & (g573)) + ((!g460) & (g464) & (!g571) & (!g572) & (sk[71]) & (!g573)));
	assign g575 = (((i_2_) & (i_9_) & (!g28) & (!g119) & (!g16) & (g180)) + ((!i_2_) & (i_9_) & (!g28) & (!g119) & (g16) & (!g180)) + ((i_2_) & (!i_9_) & (!g28) & (!g119) & (g16) & (!g180)));
	assign g576 = (((i_9_) & (!g7) & (g36) & (g16) & (!g45) & (g11)) + ((i_9_) & (g7) & (!g36) & (!g16) & (!g45) & (g11)));
	assign g577 = (((i_9_) & (!g7) & (!sk[74]) & (!g3) & (g125)) + ((i_9_) & (g7) & (!sk[74]) & (!g3) & (!g125)) + ((!i_9_) & (g7) & (sk[74]) & (!g3) & (!g125)));
	assign g578 = (((i_9_) & (!sk[75]) & (i_3_) & (!i_4_) & (!g25)) + ((i_9_) & (!sk[75]) & (!i_3_) & (!i_4_) & (g25)) + ((i_9_) & (!sk[75]) & (i_3_) & (!i_4_) & (g25)) + ((!i_9_) & (sk[75]) & (!i_3_) & (!i_4_) & (g25)));
	assign g579 = (((i_5_) & (!sk[76]) & (!g54) & (!g63) & (!g577) & (!g578)) + ((!i_5_) & (!sk[76]) & (g54) & (g63) & (!g577) & (!g578)) + ((!i_5_) & (sk[76]) & (!g54) & (g63) & (g577) & (!g578)) + ((!i_5_) & (!sk[76]) & (!g54) & (!g63) & (g577) & (g578)) + ((!i_5_) & (sk[76]) & (!g54) & (!g63) & (!g577) & (g578)));
	assign g580 = (((!i_9_) & (g39) & (!g3) & (!g92) & (g117) & (!g224)) + ((i_9_) & (!g39) & (!g3) & (!g92) & (!g117) & (g224)) + ((i_9_) & (g39) & (!g3) & (g92) & (!g117) & (!g224)));
	assign g581 = (((g26) & (g58) & (!sk[78]) & (!g53) & (!g440)) + ((g26) & (!g58) & (sk[78]) & (g53) & (!g440)) + ((!g26) & (!g58) & (sk[78]) & (!g53) & (g440)) + ((g26) & (!g58) & (!sk[78]) & (!g53) & (g440)));
	assign g582 = (((!i_9_) & (!g25) & (!g120) & (!g183) & (!g179) & (!g581)) + ((i_9_) & (!g25) & (!g120) & (!g183) & (!g179) & (!g581)) + ((!i_9_) & (!g25) & (!g120) & (!g183) & (!g179) & (!g581)));
	assign g583 = (((g575) & (!g576) & (!g579) & (!sk[80]) & (!g580) & (!g582)) + ((!g575) & (g576) & (g579) & (!sk[80]) & (!g580) & (!g582)) + ((!g575) & (!g576) & (!g579) & (!sk[80]) & (g580) & (g582)) + ((!g575) & (!g576) & (!g579) & (sk[80]) & (!g580) & (g582)));
	assign g584 = (((g547) & (g735) & (g557) & (g570) & (g574) & (g583)));
	assign g585 = (((g89) & (!g372) & (!sk[82]) & (!g507) & (!g545) & (!g584)) + ((!g89) & (g372) & (!sk[82]) & (g507) & (!g545) & (!g584)) + ((!g89) & (!g372) & (!sk[82]) & (!g507) & (g545) & (g584)) + ((g89) & (g372) & (!sk[82]) & (g507) & (g545) & (g584)));
	assign g586 = (((i_9_) & (g101) & (!g59) & (!sk[83]) & (!g141)) + ((i_9_) & (!g101) & (g59) & (!sk[83]) & (g141)) + ((i_9_) & (!g101) & (!g59) & (!sk[83]) & (g141)) + ((!i_9_) & (g101) & (g59) & (sk[83]) & (!g141)));
	assign g587 = (((g22) & (g36) & (!g26) & (!sk[84]) & (!g53)) + ((g22) & (g36) & (!g26) & (!sk[84]) & (g53)) + ((!g22) & (!g36) & (g26) & (sk[84]) & (g53)) + ((g22) & (!g36) & (!g26) & (!sk[84]) & (g53)));
	assign g588 = (((!sk[85]) & (g50) & (!g35) & (!g76) & (g587)) + ((sk[85]) & (!g50) & (!g35) & (!g76) & (!g587)) + ((sk[85]) & (!g50) & (!g35) & (g76) & (!g587)) + ((!sk[85]) & (g50) & (g35) & (!g76) & (!g587)));
	assign g589 = (((g124) & (g137) & (!sk[86]) & (!g2) & (!g46)) + ((g124) & (!g137) & (!sk[86]) & (!g2) & (g46)) + ((!g124) & (!g137) & (sk[86]) & (g2) & (g46)));
	assign g590 = (((g22) & (!g36) & (!sk[87]) & (!g6) & (!g73) & (!g4)) + ((!g22) & (g36) & (!sk[87]) & (g6) & (!g73) & (!g4)) + ((!g22) & (!g36) & (!sk[87]) & (!g6) & (g73) & (g4)) + ((g22) & (!g36) & (!sk[87]) & (!g6) & (g73) & (!g4)) + ((!g22) & (g36) & (sk[87]) & (!g6) & (g73) & (!g4)));
	assign g591 = (((g39) & (g20) & (g30) & (!sk[88]) & (!g59)) + ((g39) & (g20) & (!g30) & (!sk[88]) & (!g59)) + ((g39) & (!g20) & (!g30) & (!sk[88]) & (g59)) + ((!g39) & (g20) & (g30) & (sk[88]) & (g59)));
	assign g592 = (((!sk[89]) & (g42) & (!g116) & (!g340) & (!g590) & (!g591)) + ((!sk[89]) & (!g42) & (g116) & (g340) & (!g590) & (!g591)) + ((!sk[89]) & (!g42) & (!g116) & (!g340) & (g590) & (g591)) + ((sk[89]) & (!g42) & (!g116) & (!g340) & (!g590) & (!g591)) + ((!sk[89]) & (g42) & (!g116) & (!g340) & (!g590) & (!g591)));
	assign g593 = (((g404) & (!g586) & (!g588) & (!sk[90]) & (!g589) & (!g592)) + ((!g404) & (g586) & (g588) & (!sk[90]) & (!g589) & (!g592)) + ((!g404) & (!g586) & (!g588) & (!sk[90]) & (g589) & (g592)) + ((g404) & (!g586) & (g588) & (!sk[90]) & (!g589) & (g592)));
	assign g594 = (((g62) & (!sk[91]) & (g27) & (!g192) & (!g224)) + ((g62) & (sk[91]) & (!g27) & (g192) & (!g224)) + ((g62) & (!sk[91]) & (!g27) & (!g192) & (g224)) + ((!g62) & (sk[91]) & (g27) & (!g192) & (g224)));
	assign g595 = (((g49) & (!sk[92]) & (g17) & (!g193) & (!g594)) + ((g49) & (!sk[92]) & (!g17) & (!g193) & (g594)) + ((!g49) & (sk[92]) & (!g17) & (!g193) & (!g594)) + ((!g49) & (sk[92]) & (!g17) & (!g193) & (!g594)));
	assign g596 = (((g125) & (!sk[93]) & (g13) & (!g2) & (!g161)) + ((g125) & (sk[93]) & (!g13) & (!g2) & (!g161)) + ((!g125) & (sk[93]) & (!g13) & (g2) & (g161)) + ((g125) & (!sk[93]) & (!g13) & (!g2) & (g161)));
	assign g597 = (((!sk[94]) & (g495) & (g325) & (!g595) & (!g596)) + ((!sk[94]) & (g495) & (!g325) & (!g595) & (g596)) + ((sk[94]) & (!g495) & (g325) & (g595) & (!g596)));
	assign g598 = (((i_9_) & (!g39) & (!g45) & (!g139) & (!sk[95]) & (!g208)) + ((!i_9_) & (g39) & (g45) & (!g139) & (!sk[95]) & (!g208)) + ((i_9_) & (!g39) & (!g45) & (!g139) & (!sk[95]) & (g208)) + ((!i_9_) & (!g39) & (!g45) & (g139) & (!sk[95]) & (g208)) + ((!i_9_) & (g39) & (!g45) & (g139) & (sk[95]) & (!g208)));
	assign g599 = (((i_9_) & (!sk[96]) & (g120) & (!g11) & (!g5)) + ((i_9_) & (!sk[96]) & (g120) & (g11) & (!g5)) + ((i_9_) & (!sk[96]) & (!g120) & (!g11) & (g5)) + ((!i_9_) & (sk[96]) & (!g120) & (g11) & (g5)));
	assign g600 = (((i_9_) & (g63) & (!sk[97]) & (!g179) & (!g158)) + ((i_9_) & (g63) & (!sk[97]) & (g179) & (!g158)) + ((i_9_) & (!g63) & (!sk[97]) & (!g179) & (g158)) + ((!i_9_) & (g63) & (sk[97]) & (!g179) & (g158)));
	assign g601 = (((!sk[98]) & (g22) & (!i_9_) & (!g10) & (!g45) & (!g148)) + ((!sk[98]) & (!g22) & (i_9_) & (g10) & (!g45) & (!g148)) + ((!sk[98]) & (g22) & (!i_9_) & (!g10) & (!g45) & (g148)) + ((!sk[98]) & (!g22) & (!i_9_) & (!g10) & (g45) & (g148)) + ((!sk[98]) & (g22) & (i_9_) & (!g10) & (!g45) & (!g148)));
	assign g602 = (((g365) & (!sk[99]) & (!g598) & (!g599) & (!g600) & (!g601)) + ((!g365) & (!sk[99]) & (g598) & (g599) & (!g600) & (!g601)) + ((!g365) & (!sk[99]) & (!g598) & (!g599) & (g600) & (g601)) + ((!g365) & (sk[99]) & (!g598) & (!g599) & (!g600) & (!g601)));
	assign g603 = (((i_9_) & (!sk[100]) & (!g59) & (!g177) & (!g55) & (!g602)) + ((!i_9_) & (!sk[100]) & (g59) & (g177) & (!g55) & (!g602)) + ((i_9_) & (!sk[100]) & (!g59) & (!g177) & (!g55) & (g602)) + ((!i_9_) & (!sk[100]) & (!g59) & (!g177) & (g55) & (g602)) + ((!i_9_) & (sk[100]) & (!g59) & (!g177) & (!g55) & (g602)) + ((!i_9_) & (sk[100]) & (!g59) & (!g177) & (!g55) & (g602)));
	assign g604 = (((!sk[101]) & (i_2_) & (!i_9_) & (!g272) & (!g156) & (!g169)) + ((!sk[101]) & (!i_2_) & (i_9_) & (g272) & (!g156) & (!g169)) + ((!sk[101]) & (!i_2_) & (!i_9_) & (!g272) & (g156) & (g169)) + ((!sk[101]) & (i_2_) & (i_9_) & (g272) & (!g156) & (g169)) + ((sk[101]) & (!i_2_) & (!i_9_) & (g272) & (g156) & (!g169)));
	assign g605 = (((!sk[102]) & (!g28) & (!g3) & (g1)) + ((!sk[102]) & (g28) & (g3) & (!g1)) + ((sk[102]) & (!g28) & (!g3) & (!g1)));
	assign g606 = (((g7) & (!sk[103]) & (!g20) & (!g16) & (!g63) & (!g13)) + ((!g7) & (!sk[103]) & (g20) & (g16) & (!g63) & (!g13)) + ((g7) & (!sk[103]) & (g20) & (!g16) & (g63) & (!g13)) + ((!g7) & (!sk[103]) & (!g20) & (!g16) & (g63) & (g13)) + ((g7) & (!sk[103]) & (!g20) & (g16) & (!g63) & (!g13)));
	assign g607 = (((!g133) & (!sk[104]) & (!g139) & (g606)) + ((!g133) & (sk[104]) & (!g139) & (!g606)) + ((g133) & (!sk[104]) & (g139) & (!g606)));
	assign g608 = (((g101) & (g42) & (!sk[105]) & (!g43) & (!g180)) + ((g101) & (!g42) & (sk[105]) & (!g43) & (!g180)) + ((!g101) & (g42) & (sk[105]) & (!g43) & (g180)) + ((g101) & (!g42) & (!sk[105]) & (!g43) & (g180)));
	assign g609 = (((g57) & (!g40) & (!g457) & (!g607) & (!sk[106]) & (!g608)) + ((!g57) & (g40) & (g457) & (!g607) & (!sk[106]) & (!g608)) + ((!g57) & (!g40) & (!g457) & (g607) & (!sk[106]) & (g608)) + ((!g57) & (!g40) & (!g457) & (g607) & (sk[106]) & (!g608)) + ((!g57) & (!g40) & (!g457) & (g607) & (sk[106]) & (!g608)));
	assign g610 = (((!i_9_) & (!g39) & (!g239) & (!g356) & (!g605) & (g609)) + ((!i_9_) & (!g39) & (!g239) & (!g356) & (!g605) & (g609)) + ((i_9_) & (!g39) & (!g239) & (!g356) & (!g605) & (g609)));
	assign g611 = (((!i_5_) & (!i_3_) & (i_4_) & (g63) & (g137) & (!g58)) + ((i_5_) & (i_3_) & (i_4_) & (g63) & (!g137) & (!g58)));
	assign g612 = (((g7) & (!g28) & (!sk[109]) & (!g73) & (!g59) & (!g1)) + ((!g7) & (g28) & (!sk[109]) & (g73) & (!g59) & (!g1)) + ((!g7) & (!g28) & (!sk[109]) & (!g73) & (g59) & (g1)) + ((g7) & (!g28) & (!sk[109]) & (g73) & (!g59) & (!g1)) + ((!g7) & (!g28) & (sk[109]) & (g73) & (g59) & (!g1)));
	assign g613 = (((i_9_) & (!g50) & (i_5_) & (!g6) & (g92) & (!g45)) + ((!i_9_) & (!g50) & (!i_5_) & (!g6) & (g92) & (!g45)));
	assign g614 = (((g38) & (!g1) & (!g14) & (!sk[111]) & (g613)) + ((g38) & (!g1) & (!g14) & (sk[111]) & (!g613)) + ((!g38) & (g1) & (!g14) & (sk[111]) & (!g613)) + ((!g38) & (!g1) & (g14) & (sk[111]) & (!g613)) + ((g38) & (g1) & (!g14) & (!sk[111]) & (!g613)));
	assign g615 = (((g7) & (!g28) & (!sk[112]) & (!g25) & (!g6) & (!g40)) + ((!g7) & (g28) & (!sk[112]) & (g25) & (!g6) & (!g40)) + ((g7) & (!g28) & (!sk[112]) & (g25) & (!g6) & (g40)) + ((!g7) & (!g28) & (!sk[112]) & (!g25) & (g6) & (g40)) + ((g7) & (!g28) & (!sk[112]) & (!g25) & (!g6) & (g40)) + ((!g7) & (!g28) & (sk[112]) & (g25) & (!g6) & (g40)));
	assign g616 = (((g38) & (!g42) & (!g122) & (!g17) & (!g46) & (!g29)) + ((!g38) & (!g42) & (!g122) & (!g17) & (!g46) & (!g29)) + ((g38) & (!g42) & (!g122) & (!g17) & (!g46) & (!g29)) + ((!g38) & (!g42) & (!g122) & (!g17) & (!g46) & (!g29)));
	assign g617 = (((g101) & (!sk[114]) & (!g21) & (!g53) & (!g23) & (!g97)) + ((!g101) & (!sk[114]) & (g21) & (g53) & (!g23) & (!g97)) + ((!g101) & (!sk[114]) & (!g21) & (!g53) & (g23) & (g97)) + ((!g101) & (sk[114]) & (!g21) & (!g53) & (!g23) & (!g97)) + ((!g101) & (sk[114]) & (!g21) & (!g53) & (!g23) & (!g97)) + ((!g101) & (sk[114]) & (g21) & (!g53) & (!g23) & (!g97)) + ((!g101) & (sk[114]) & (g21) & (!g53) & (!g23) & (!g97)));
	assign g618 = (((g21) & (!sk[115]) & (!g165) & (!g615) & (!g616) & (!g617)) + ((!g21) & (!sk[115]) & (g165) & (g615) & (!g616) & (!g617)) + ((!g21) & (!sk[115]) & (!g165) & (!g615) & (g616) & (g617)) + ((g21) & (!sk[115]) & (!g165) & (!g615) & (g616) & (g617)) + ((!g21) & (!sk[115]) & (!g165) & (!g615) & (g616) & (g617)));
	assign g619 = (((!sk[116]) & (g13) & (!g177) & (!g612) & (!g614) & (!g618)) + ((!sk[116]) & (!g13) & (g177) & (g612) & (!g614) & (!g618)) + ((!sk[116]) & (!g13) & (!g177) & (!g612) & (g614) & (g618)) + ((!sk[116]) & (g13) & (!g177) & (!g612) & (g614) & (g618)) + ((!sk[116]) & (!g13) & (!g177) & (!g612) & (g614) & (g618)));
	assign g620 = (((g8) & (!g36) & (!g122) & (!sk[117]) & (g133)) + ((g8) & (g36) & (!g122) & (!sk[117]) & (!g133)) + ((!g8) & (!g36) & (g122) & (sk[117]) & (!g133)));
	assign g621 = (((!sk[118]) & (g35) & (!g43) & (!g165) & (g244)) + ((!sk[118]) & (g35) & (g43) & (!g165) & (!g244)) + ((sk[118]) & (!g35) & (!g43) & (g165) & (!g244)));
	assign g622 = (((g7) & (!sk[119]) & (!g39) & (!g16) & (!g133) & (!g53)) + ((!g7) & (!sk[119]) & (g39) & (g16) & (!g133) & (!g53)) + ((g7) & (!sk[119]) & (!g39) & (g16) & (!g133) & (!g53)) + ((g7) & (!sk[119]) & (g39) & (!g16) & (!g133) & (g53)) + ((!g7) & (!sk[119]) & (!g39) & (!g16) & (g133) & (g53)));
	assign g623 = (((g620) & (!g176) & (!g185) & (!sk[120]) & (!g621) & (!g622)) + ((!g620) & (g176) & (g185) & (!sk[120]) & (!g621) & (!g622)) + ((!g620) & (!g176) & (!g185) & (!sk[120]) & (g621) & (g622)) + ((!g620) & (g176) & (g185) & (!sk[120]) & (!g621) & (!g622)));
	assign g624 = (((g604) & (!g610) & (!g611) & (!g619) & (!sk[121]) & (!g623)) + ((!g604) & (g610) & (g611) & (!g619) & (!sk[121]) & (!g623)) + ((!g604) & (!g610) & (!g611) & (g619) & (!sk[121]) & (g623)) + ((!g604) & (g610) & (!g611) & (g619) & (!sk[121]) & (g623)));
	assign g625 = (((i_9_) & (i_8_) & (!i_6_) & (!i_7_) & (g99) & (!g195)) + ((i_9_) & (i_8_) & (!i_6_) & (i_7_) & (!g99) & (g195)));
	assign g626 = (((g547) & (!sk[123]) & (!g397) & (!g474) & (!g503) & (!g625)) + ((!g547) & (!sk[123]) & (g397) & (g474) & (!g503) & (!g625)) + ((!g547) & (!sk[123]) & (!g397) & (!g474) & (g503) & (g625)) + ((g547) & (!sk[123]) & (g397) & (g474) & (g503) & (!g625)));
	assign g627 = (((g237) & (g593) & (g597) & (g603) & (g624) & (g626)));
	assign g628 = (((g22) & (i_9_) & (!sk[125]) & (!g182) & (!g186)) + ((g22) & (i_9_) & (!sk[125]) & (g182) & (!g186)) + ((g22) & (!i_9_) & (!sk[125]) & (!g182) & (g186)));
	assign g629 = (((!sk[126]) & (g20) & (!g137) & (!g60) & (g307)) + ((!sk[126]) & (g20) & (g137) & (!g60) & (!g307)) + ((sk[126]) & (!g20) & (g137) & (g60) & (!g307)));
	assign g630 = (((g38) & (!sk[127]) & (!g137) & (!g52) & (!g222) & (!g331)) + ((!g38) & (!sk[127]) & (g137) & (g52) & (!g222) & (!g331)) + ((!g38) & (!sk[127]) & (!g137) & (!g52) & (g222) & (g331)) + ((!g38) & (!sk[127]) & (g137) & (!g52) & (g222) & (g331)) + ((!g38) & (!sk[127]) & (!g137) & (g52) & (g222) & (g331)) + ((!g38) & (sk[127]) & (!g137) & (g52) & (!g222) & (g331)));
	assign g631 = (((!sk[0]) & (g76) & (!g3) & (!g21) & (!g171) & (!g193)) + ((!sk[0]) & (!g76) & (g3) & (g21) & (!g171) & (!g193)) + ((sk[0]) & (!g76) & (!g3) & (!g21) & (g171) & (!g193)) + ((sk[0]) & (!g76) & (!g3) & (!g21) & (!g171) & (g193)) + ((!sk[0]) & (!g76) & (!g3) & (!g21) & (g171) & (g193)) + ((sk[0]) & (!g76) & (!g3) & (!g21) & (!g171) & (!g193)));
	assign g632 = (((g53) & (!sk[1]) & (g440) & (!g630) & (!g631)) + ((g53) & (!sk[1]) & (!g440) & (!g630) & (g631)) + ((!g53) & (sk[1]) & (!g440) & (!g630) & (!g631)) + ((!g53) & (sk[1]) & (!g440) & (!g630) & (!g631)));
	assign g633 = (((g43) & (!g209) & (!g628) & (!g629) & (!sk[2]) & (!g632)) + ((!g43) & (g209) & (g628) & (!g629) & (!sk[2]) & (!g632)) + ((!g43) & (!g209) & (!g628) & (g629) & (!sk[2]) & (g632)) + ((g43) & (!g209) & (!g628) & (!g629) & (!sk[2]) & (g632)) + ((!g43) & (!g209) & (!g628) & (!g629) & (sk[2]) & (g632)));
	assign g634 = (((!sk[3]) & (i_5_) & (!i_3_) & (!i_4_) & (!g25) & (!g137)) + ((!sk[3]) & (!i_5_) & (i_3_) & (i_4_) & (!g25) & (!g137)) + ((!sk[3]) & (!i_5_) & (!i_3_) & (!i_4_) & (g25) & (g137)) + ((!sk[3]) & (i_5_) & (i_3_) & (i_4_) & (g25) & (!g137)) + ((!sk[3]) & (i_5_) & (i_3_) & (!i_4_) & (g25) & (g137)));
	assign g635 = (((!sk[4]) & (i_9_) & (i_8_) & (!i_6_) & (!g634)) + ((!sk[4]) & (i_9_) & (!i_8_) & (!i_6_) & (g634)) + ((!sk[4]) & (i_9_) & (!i_8_) & (!i_6_) & (g634)));
	assign g636 = (((g40) & (!g243) & (!sk[5]) & (!g440) & (!g633) & (!g635)) + ((!g40) & (g243) & (!sk[5]) & (g440) & (!g633) & (!g635)) + ((!g40) & (!g243) & (!sk[5]) & (!g440) & (g633) & (g635)) + ((!g40) & (!g243) & (sk[5]) & (!g440) & (g633) & (!g635)) + ((!g40) & (!g243) & (!sk[5]) & (!g440) & (g633) & (g635)));
	assign g637 = (((i_9_) & (!sk[6]) & (!g6) & (!g30) & (!g134) & (!g138)) + ((!i_9_) & (!sk[6]) & (g6) & (g30) & (!g134) & (!g138)) + ((!i_9_) & (!sk[6]) & (!g6) & (!g30) & (g134) & (g138)) + ((!i_9_) & (sk[6]) & (!g6) & (!g30) & (g134) & (!g138)) + ((i_9_) & (!sk[6]) & (!g6) & (g30) & (!g134) & (g138)));
	assign g638 = (((i_9_) & (!g7) & (!sk[7]) & (!g63) & (!g30) & (!g138)) + ((!i_9_) & (g7) & (!sk[7]) & (g63) & (!g30) & (!g138)) + ((!i_9_) & (!g7) & (!sk[7]) & (!g63) & (g30) & (g138)) + ((i_9_) & (g7) & (!sk[7]) & (g63) & (!g30) & (g138)) + ((!i_9_) & (!g7) & (!sk[7]) & (g63) & (g30) & (g138)));
	assign g639 = (((i_9_) & (!i_8_) & (!i_6_) & (!sk[8]) & (!i_7_) & (!i_5_)) + ((!i_9_) & (i_8_) & (i_6_) & (!sk[8]) & (!i_7_) & (!i_5_)) + ((!i_9_) & (!i_8_) & (!i_6_) & (!sk[8]) & (i_7_) & (i_5_)) + ((i_9_) & (i_8_) & (!i_6_) & (!sk[8]) & (!i_7_) & (i_5_)) + ((i_9_) & (i_8_) & (i_6_) & (!sk[8]) & (i_7_) & (!i_5_)));
	assign g640 = (((i_3_) & (!sk[9]) & (i_4_) & (!g1) & (!g639)) + ((i_3_) & (!sk[9]) & (!i_4_) & (!g1) & (g639)) + ((i_3_) & (!sk[9]) & (!i_4_) & (!g1) & (g639)));
	assign g641 = (((g13) & (!sk[10]) & (g85) & (!g638) & (!g640)) + ((g13) & (!sk[10]) & (!g85) & (!g638) & (g640)) + ((!g13) & (sk[10]) & (!g85) & (!g638) & (!g640)) + ((g13) & (!sk[10]) & (g85) & (!g638) & (!g640)));
	assign g642 = (((!sk[11]) & (g36) & (!g54) & (!g28) & (!g6) & (!g58)) + ((!sk[11]) & (!g36) & (g54) & (g28) & (!g6) & (!g58)) + ((!sk[11]) & (g36) & (!g54) & (!g28) & (!g6) & (!g58)) + ((!sk[11]) & (!g36) & (!g54) & (!g28) & (g6) & (g58)) + ((sk[11]) & (!g36) & (!g54) & (!g28) & (!g6) & (!g58)));
	assign g643 = (((!i_2_) & (g78) & (i_9_) & (g122) & (!g168) & (!g85)) + ((i_2_) & (g78) & (i_9_) & (!g122) & (g168) & (!g85)) + ((!i_2_) & (g78) & (!i_9_) & (!g122) & (g168) & (!g85)) + ((i_2_) & (g78) & (!i_9_) & (!g122) & (!g168) & (g85)));
	assign g644 = (((i_9_) & (g39) & (!g1) & (!g37) & (!g32) & (!g228)) + ((!i_9_) & (!g39) & (!g1) & (!g37) & (!g32) & (!g228)) + ((!i_9_) & (g39) & (!g1) & (!g37) & (g32) & (!g228)) + ((i_9_) & (!g39) & (!g1) & (!g37) & (!g32) & (g228)));
	assign g645 = (((!i_9_) & (i_5_) & (!i_3_) & (!i_4_) & (!g3) & (g11)) + ((i_9_) & (i_5_) & (i_3_) & (i_4_) & (!g3) & (g11)));
	assign g646 = (((g35) & (!g42) & (!g3) & (!g10) & (!g18) & (!g21)) + ((!g35) & (g42) & (!g3) & (!g10) & (!g18) & (!g21)) + ((!g35) & (!g42) & (!g3) & (!g10) & (g18) & (!g21)));
	assign g647 = (((g7) & (!g16) & (!g43) & (!g645) & (!sk[16]) & (!g646)) + ((!g7) & (g16) & (g43) & (!g645) & (!sk[16]) & (!g646)) + ((!g7) & (!g16) & (!g43) & (g645) & (!sk[16]) & (g646)) + ((!g7) & (!g16) & (!g43) & (!g645) & (sk[16]) & (!g646)) + ((!g7) & (!g16) & (!g43) & (!g645) & (sk[16]) & (!g646)) + ((!g7) & (!g16) & (g43) & (!g645) & (sk[16]) & (!g646)));
	assign g648 = (((g641) & (!g642) & (!g643) & (!sk[17]) & (!g644) & (!g647)) + ((!g641) & (g642) & (g643) & (!sk[17]) & (!g644) & (!g647)) + ((!g641) & (!g642) & (!g643) & (!sk[17]) & (g644) & (g647)) + ((g641) & (!g642) & (!g643) & (!sk[17]) & (!g644) & (g647)));
	assign g649 = (((!g78) & (!sk[18]) & (!g54) & (g10)) + ((g78) & (!sk[18]) & (g54) & (!g10)) + ((g78) & (sk[18]) & (!g54) & (!g10)));
	assign g650 = (((i_2_) & (!sk[19]) & (!g16) & (!g14) & (!g151) & (!g649)) + ((!i_2_) & (!sk[19]) & (g16) & (g14) & (!g151) & (!g649)) + ((!i_2_) & (!sk[19]) & (!g16) & (!g14) & (g151) & (g649)) + ((i_2_) & (!sk[19]) & (g16) & (!g14) & (g151) & (!g649)));
	assign g651 = (((g22) & (!sk[20]) & (!i_9_) & (!g1) & (!g44) & (!g156)) + ((!g22) & (!sk[20]) & (i_9_) & (g1) & (!g44) & (!g156)) + ((g22) & (!sk[20]) & (i_9_) & (!g1) & (!g44) & (g156)) + ((!g22) & (!sk[20]) & (!i_9_) & (!g1) & (g44) & (g156)) + ((!g22) & (sk[20]) & (!i_9_) & (!g1) & (g44) & (!g156)));
	assign g652 = (((!sk[21]) & (i_9_) & (!g16) & (!g63) & (!g156) & (!g354)) + ((!sk[21]) & (!i_9_) & (g16) & (g63) & (!g156) & (!g354)) + ((!sk[21]) & (i_9_) & (g16) & (!g63) & (!g156) & (g354)) + ((!sk[21]) & (!i_9_) & (!g16) & (!g63) & (g156) & (g354)) + ((sk[21]) & (!i_9_) & (!g16) & (g63) & (g156) & (!g354)));
	assign g653 = (((g22) & (!sk[22]) & (!i_9_) & (!g7) & (!g40) & (!g356)) + ((!g22) & (!sk[22]) & (i_9_) & (g7) & (!g40) & (!g356)) + ((g22) & (!sk[22]) & (!i_9_) & (g7) & (g40) & (!g356)) + ((g22) & (!sk[22]) & (!i_9_) & (!g7) & (!g40) & (g356)) + ((!g22) & (!sk[22]) & (!i_9_) & (!g7) & (g40) & (g356)));
	assign g654 = (((!sk[23]) & (g133) & (!g422) & (!g651) & (!g652) & (!g653)) + ((!sk[23]) & (!g133) & (g422) & (g651) & (!g652) & (!g653)) + ((!sk[23]) & (!g133) & (!g422) & (!g651) & (g652) & (g653)) + ((!sk[23]) & (g133) & (!g422) & (!g651) & (!g652) & (!g653)) + ((sk[23]) & (!g133) & (!g422) & (!g651) & (!g652) & (!g653)));
	assign g655 = (((g219) & (g494) & (!sk[24]) & (!g650) & (!g654)) + ((g219) & (!g494) & (!sk[24]) & (!g650) & (g654)) + ((g219) & (!g494) & (!sk[24]) & (!g650) & (g654)));
	assign g656 = (((g147) & (!g610) & (!sk[25]) & (!g637) & (!g648) & (!g655)) + ((!g147) & (g610) & (!sk[25]) & (g637) & (!g648) & (!g655)) + ((!g147) & (!g610) & (!sk[25]) & (!g637) & (g648) & (g655)) + ((g147) & (g610) & (!sk[25]) & (!g637) & (g648) & (g655)));
	assign g657 = (((i_9_) & (!g39) & (!g3) & (!g30) & (!sk[26]) & (!g77)) + ((!i_9_) & (g39) & (g3) & (!g30) & (!sk[26]) & (!g77)) + ((i_9_) & (g39) & (!g3) & (!g30) & (!sk[26]) & (g77)) + ((!i_9_) & (!g39) & (!g3) & (g30) & (!sk[26]) & (g77)) + ((!i_9_) & (g39) & (!g3) & (g30) & (sk[26]) & (!g77)));
	assign g658 = (((!sk[27]) & (i_9_) & (g25) & (!g17) & (!g139)) + ((!sk[27]) & (i_9_) & (!g25) & (!g17) & (g139)) + ((!sk[27]) & (i_9_) & (g25) & (!g17) & (g139)) + ((sk[27]) & (!i_9_) & (g25) & (g17) & (!g139)));
	assign g659 = (((i_2_) & (!sk[28]) & (g78) & (!i_9_) & (!g4)) + ((!i_2_) & (sk[28]) & (g78) & (i_9_) & (!g4)) + ((i_2_) & (!sk[28]) & (!g78) & (!i_9_) & (g4)) + ((!i_2_) & (sk[28]) & (g78) & (!i_9_) & (!g4)));
	assign g660 = (((g787) & (!sk[29]) & (!g401) & (!g657) & (!g658) & (!g659)) + ((!g787) & (!sk[29]) & (g401) & (g657) & (!g658) & (!g659)) + ((!g787) & (!sk[29]) & (!g401) & (!g657) & (g658) & (g659)) + ((g787) & (!sk[29]) & (!g401) & (!g657) & (!g658) & (!g659)) + ((g787) & (!sk[29]) & (!g401) & (!g657) & (!g658) & (!g659)));
	assign g661 = (((g294) & (!sk[30]) & (!g382) & (!g391) & (!g510) & (!g660)) + ((!g294) & (!sk[30]) & (g382) & (g391) & (!g510) & (!g660)) + ((!g294) & (!sk[30]) & (!g382) & (!g391) & (g510) & (g660)) + ((g294) & (!sk[30]) & (!g382) & (g391) & (g510) & (g660)));
	assign g662 = (((g317) & (g479) & (g557) & (g636) & (g656) & (g661)));
	assign g663 = (((i_9_) & (!g45) & (!g221) & (!g138) & (!sk[32]) & (!g302)) + ((!i_9_) & (g45) & (g221) & (!g138) & (!sk[32]) & (!g302)) + ((i_9_) & (!g45) & (!g221) & (g138) & (!sk[32]) & (g302)) + ((!i_9_) & (!g45) & (!g221) & (g138) & (!sk[32]) & (g302)) + ((!i_9_) & (!g45) & (g221) & (!g138) & (sk[32]) & (!g302)));
	assign g664 = (((!sk[33]) & (i_9_) & (!i_8_) & (!i_6_) & (!i_7_) & (!i_5_)) + ((!sk[33]) & (!i_9_) & (i_8_) & (i_6_) & (!i_7_) & (!i_5_)) + ((!sk[33]) & (!i_9_) & (!i_8_) & (!i_6_) & (i_7_) & (i_5_)) + ((!sk[33]) & (i_9_) & (i_8_) & (!i_6_) & (!i_7_) & (i_5_)) + ((!sk[33]) & (i_9_) & (!i_8_) & (!i_6_) & (i_7_) & (!i_5_)));
	assign g665 = (((g22) & (!i_3_) & (!sk[34]) & (!i_4_) & (!g206) & (!g664)) + ((!g22) & (i_3_) & (!sk[34]) & (i_4_) & (!g206) & (!g664)) + ((!g22) & (!i_3_) & (!sk[34]) & (!i_4_) & (g206) & (g664)) + ((g22) & (!i_3_) & (!sk[34]) & (i_4_) & (g206) & (g664)));
	assign g666 = (((i_9_) & (!sk[35]) & (!g8) & (!g59) & (!g10) & (!g142)) + ((!i_9_) & (!sk[35]) & (g8) & (g59) & (!g10) & (!g142)) + ((!i_9_) & (!sk[35]) & (!g8) & (!g59) & (g10) & (g142)) + ((i_9_) & (!sk[35]) & (g8) & (g59) & (!g10) & (!g142)) + ((!i_9_) & (sk[35]) & (g8) & (!g59) & (!g10) & (!g142)));
	assign g667 = (((g35) & (!g116) & (!sk[36]) & (!g43) & (!g158) & (!g193)) + ((!g35) & (!g116) & (!sk[36]) & (!g43) & (g158) & (g193)) + ((!g35) & (!g116) & (sk[36]) & (!g43) & (!g158) & (!g193)) + ((!g35) & (g116) & (!sk[36]) & (g43) & (!g158) & (!g193)) + ((!g35) & (!g116) & (sk[36]) & (g43) & (!g158) & (!g193)) + ((!g35) & (!g116) & (sk[36]) & (g43) & (!g158) & (!g193)) + ((!g35) & (!g116) & (sk[36]) & (!g43) & (!g158) & (!g193)));
	assign g668 = (((!sk[37]) & (g13) & (!g141) & (!g225) & (g667)) + ((!sk[37]) & (g13) & (g141) & (!g225) & (!g667)) + ((sk[37]) & (!g13) & (!g141) & (!g225) & (g667)));
	assign g669 = (((!sk[38]) & (i_9_) & (i_8_) & (!i_6_) & (!g221)) + ((!sk[38]) & (i_9_) & (!i_8_) & (!i_6_) & (g221)) + ((!sk[38]) & (i_9_) & (i_8_) & (i_6_) & (g221)));
	assign g670 = (((i_9_) & (i_5_) & (g16) & (!sk[39]) & (!g138)) + ((i_9_) & (i_5_) & (!g16) & (!sk[39]) & (!g138)) + ((i_9_) & (!i_5_) & (!g16) & (!sk[39]) & (g138)));
	assign g671 = (((i_3_) & (!i_4_) & (!g63) & (!sk[40]) & (!g669) & (!g670)) + ((i_3_) & (!i_4_) & (!g63) & (!sk[40]) & (!g669) & (!g670)) + ((!i_3_) & (i_4_) & (g63) & (!sk[40]) & (!g669) & (!g670)) + ((!i_3_) & (!i_4_) & (!g63) & (sk[40]) & (!g669) & (!g670)) + ((!i_3_) & (!i_4_) & (!g63) & (!sk[40]) & (g669) & (g670)) + ((!i_3_) & (!i_4_) & (!g63) & (sk[40]) & (!g669) & (!g670)) + ((!i_3_) & (i_4_) & (!g63) & (sk[40]) & (!g669) & (!g670)));
	assign g672 = (((g663) & (!sk[41]) & (!g665) & (!g666) & (!g668) & (!g671)) + ((!g663) & (!sk[41]) & (g665) & (g666) & (!g668) & (!g671)) + ((!g663) & (!sk[41]) & (!g665) & (!g666) & (g668) & (g671)) + ((!g663) & (!sk[41]) & (!g665) & (!g666) & (g668) & (g671)));
	assign g673 = (((g22) & (!i_9_) & (!sk[42]) & (!i_3_) & (!i_4_) & (!g68)) + ((!g22) & (i_9_) & (!sk[42]) & (i_3_) & (!i_4_) & (!g68)) + ((!g22) & (!i_9_) & (!sk[42]) & (!i_3_) & (i_4_) & (g68)) + ((g22) & (i_9_) & (!sk[42]) & (i_3_) & (!i_4_) & (g68)));
	assign g674 = (((g7) & (!g20) & (!g76) & (!sk[43]) & (!g137) & (!g673)) + ((!g7) & (g20) & (g76) & (!sk[43]) & (!g137) & (!g673)) + ((g7) & (g20) & (!g76) & (!sk[43]) & (!g137) & (g673)) + ((g7) & (!g20) & (!g76) & (!sk[43]) & (!g137) & (g673)) + ((!g7) & (g20) & (!g76) & (!sk[43]) & (g137) & (g673)) + ((!g7) & (!g20) & (!g76) & (!sk[43]) & (g137) & (g673)) + ((!g7) & (!g20) & (!g76) & (!sk[43]) & (g137) & (g673)));
	assign g675 = (((!sk[44]) & (g242) & (g232)));
	assign g676 = (((!sk[45]) & (g16) & (g45) & (!g133) & (!g14)) + ((!sk[45]) & (g16) & (!g45) & (!g133) & (g14)) + ((sk[45]) & (!g16) & (!g45) & (!g133) & (!g14)) + ((!sk[45]) & (g16) & (g45) & (!g133) & (!g14)));
	assign g677 = (((g7) & (!g1) & (!sk[46]) & (!g27) & (g676)) + ((!g7) & (!g1) & (sk[46]) & (!g27) & (!g676)) + ((!g7) & (!g1) & (sk[46]) & (!g27) & (!g676)) + ((g7) & (g1) & (!sk[46]) & (!g27) & (!g676)));
	assign g678 = (((i_2_) & (!i_9_) & (!g119) & (g182) & (!g55) & (!g97)) + ((!i_2_) & (i_9_) & (!g119) & (!g182) & (g55) & (!g97)) + ((i_2_) & (i_9_) & (!g119) & (!g182) & (!g55) & (g97)) + ((!i_2_) & (!i_9_) & (!g119) & (!g182) & (!g55) & (g97)));
	assign g679 = (((i_9_) & (!g30) & (!g59) & (!g45) & (!sk[48]) & (!g18)) + ((!i_9_) & (g30) & (g59) & (!g45) & (!sk[48]) & (!g18)) + ((!i_9_) & (!g30) & (!g59) & (g45) & (!sk[48]) & (g18)) + ((i_9_) & (g30) & (g59) & (!g45) & (!sk[48]) & (!g18)) + ((!i_9_) & (g30) & (g59) & (!g45) & (!sk[48]) & (g18)));
	assign g680 = (((g21) & (!g40) & (!g112) & (!g233) & (!sk[49]) & (!g679)) + ((!g21) & (g40) & (g112) & (!g233) & (!sk[49]) & (!g679)) + ((!g21) & (!g40) & (!g112) & (g233) & (!sk[49]) & (g679)) + ((g21) & (!g40) & (!g112) & (!g233) & (!sk[49]) & (!g679)) + ((g21) & (!g40) & (!g112) & (!g233) & (!sk[49]) & (!g679)) + ((!g21) & (!g40) & (!g112) & (!g233) & (sk[49]) & (!g679)) + ((!g21) & (!g40) & (!g112) & (!g233) & (sk[49]) & (!g679)));
	assign g681 = (((g38) & (!g25) & (!g4) & (!g10) & (!sk[50]) & (!g11)) + ((!g38) & (g25) & (g4) & (!g10) & (!sk[50]) & (!g11)) + ((!g38) & (!g25) & (!g4) & (g10) & (!sk[50]) & (g11)) + ((!g38) & (g25) & (!g4) & (!g10) & (sk[50]) & (!g11)) + ((!g38) & (!g25) & (!g4) & (!g10) & (sk[50]) & (g11)));
	assign g682 = (((!sk[51]) & (g2) & (g158) & (!g201) & (!g681)) + ((!sk[51]) & (g2) & (!g158) & (!g201) & (g681)) + ((sk[51]) & (!g2) & (!g158) & (!g201) & (!g681)) + ((sk[51]) & (!g2) & (!g158) & (!g201) & (!g681)));
	assign g683 = (((!g28) & (g42) & (!g59) & (!g10) & (g18) & (!g58)) + ((!g28) & (!g42) & (g59) & (!g10) & (!g18) & (!g58)) + ((!g28) & (!g42) & (g59) & (!g10) & (!g18) & (!g58)));
	assign g684 = (((!sk[53]) & (i_8_) & (!g7) & (!g35) & (!g68) & (!g42)) + ((!sk[53]) & (!i_8_) & (g7) & (g35) & (!g68) & (!g42)) + ((!sk[53]) & (!i_8_) & (!g7) & (!g35) & (g68) & (g42)) + ((!sk[53]) & (!i_8_) & (g7) & (!g35) & (g68) & (g42)) + ((!sk[53]) & (i_8_) & (g7) & (g35) & (g68) & (!g42)));
	assign g685 = (((g35) & (!sk[54]) & (g180) & (!g259) & (!g684)) + ((g35) & (!sk[54]) & (!g180) & (!g259) & (g684)) + ((!g35) & (sk[54]) & (!g180) & (!g259) & (!g684)) + ((!g35) & (sk[54]) & (!g180) & (!g259) & (!g684)));
	assign g686 = (((g680) & (g682) & (!g683) & (!sk[55]) & (!g685)) + ((g680) & (!g682) & (!g683) & (!sk[55]) & (g685)) + ((g680) & (g682) & (!g683) & (!sk[55]) & (g685)));
	assign g687 = (((g155) & (g677) & (!sk[56]) & (!g678) & (!g686)) + ((g155) & (!g677) & (!sk[56]) & (!g678) & (g686)) + ((g155) & (g677) & (!sk[56]) & (!g678) & (g686)));
	assign g688 = (((!g575) & (g593) & (g633) & (!g674) & (g675) & (g687)));
	assign g689 = (((g321) & (g414) & (g484) & (g498) & (g672) & (g688)));
	assign g690 = (((g4) & (!sk[59]) & (g691)) + ((!g4) & (sk[59]) & (!g691)));
	assign g691 = (((!sk[60]) & (g4) & (g692)) + ((sk[60]) & (!g4) & (g692)));
	assign g692 = (((!sk[61]) & (g693) & (g694)) + ((sk[61]) & (!g693) & (!g694)));
	assign g693 = (((!sk[62]) & (i_1_) & (g695)) + ((sk[62]) & (!i_1_) & (g695)));
	assign g694 = (((i_1_) & (!sk[63]) & (g696)));
	assign g695 = (((g511) & (i_0_) & (!sk[64]) & (!g38) & (!i_2_)) + ((!g511) & (!i_0_) & (sk[64]) & (!g38) & (!i_2_)) + ((!g511) & (!i_0_) & (sk[64]) & (g38) & (!i_2_)) + ((g511) & (!i_0_) & (!sk[64]) & (!g38) & (i_2_)));
	assign g696 = (((!g511) & (!i_0_) & (sk[65]) & (!g58) & (!i_2_)) + ((!g511) & (!i_0_) & (sk[65]) & (!g58) & (!i_2_)) + ((g511) & (!i_0_) & (!sk[65]) & (!g58) & (i_2_)) + ((g511) & (i_0_) & (!sk[65]) & (!g58) & (!i_2_)) + ((g511) & (i_0_) & (!sk[65]) & (g58) & (!i_2_)));
	assign g697 = (((i_9_) & (!sk[66]) & (g698)) + ((i_9_) & (sk[66]) & (!g698)));
	assign g698 = (((i_9_) & (!sk[67]) & (g699)));
	assign g699 = (((g700) & (!sk[68]) & (g701)) + ((!g700) & (sk[68]) & (!g701)));
	assign g700 = (((!sk[69]) & (i_7_) & (g702)) + ((sk[69]) & (!i_7_) & (g702)));
	assign g701 = (((!sk[70]) & (i_7_) & (g703)));
	assign g702 = (((g6) & (!sk[71]) & (i_6_) & (!g7) & (!i_8_)) + ((!g6) & (sk[71]) & (!i_6_) & (!g7) & (!i_8_)) + ((!g6) & (sk[71]) & (!i_6_) & (!g7) & (!i_8_)) + ((g6) & (!sk[71]) & (!i_6_) & (!g7) & (i_8_)) + ((!g6) & (sk[71]) & (!i_6_) & (!g7) & (!i_8_)));
	assign g703 = (((!sk[72]) & (!i_6_) & (!g74) & (i_8_)) + ((sk[72]) & (i_6_) & (!g74) & (!i_8_)) + ((sk[72]) & (!i_6_) & (g74) & (!i_8_)) + ((!sk[72]) & (i_6_) & (g74) & (!i_8_)));
	assign g704 = (((!sk[73]) & (i_5_) & (g705)) + ((sk[73]) & (!i_5_) & (!g705)));
	assign g705 = (((!i_5_) & (sk[74]) & (g706)) + ((i_5_) & (!sk[74]) & (g706)));
	assign g706 = (((g707) & (!sk[75]) & (g708)) + ((!g707) & (sk[75]) & (!g708)));
	assign g707 = (((!i_4_) & (sk[76]) & (g709)) + ((i_4_) & (!sk[76]) & (g709)));
	assign g708 = (((i_4_) & (!sk[77]) & (g710)));
	assign g709 = (((g480) & (g138) & (!g13) & (!sk[78]) & (!i_3_)) + ((!g480) & (!g138) & (!g13) & (sk[78]) & (!i_3_)) + ((!g480) & (!g138) & (g13) & (sk[78]) & (!i_3_)) + ((g480) & (!g138) & (!g13) & (!sk[78]) & (i_3_)) + ((!g480) & (!g138) & (!g13) & (sk[78]) & (i_3_)));
	assign g710 = (((g480) & (g138) & (!g43) & (!sk[79]) & (!i_3_)) + ((!g480) & (!g138) & (!g43) & (sk[79]) & (!i_3_)) + ((!g480) & (!g138) & (g43) & (sk[79]) & (!i_3_)) + ((g480) & (!g138) & (!g43) & (!sk[79]) & (i_3_)) + ((!g480) & (!g138) & (!g43) & (sk[79]) & (i_3_)));
	assign g711 = (((g712) & (!sk[80]) & (g713)) + ((!g712) & (sk[80]) & (!g713)));
	assign g712 = (((!sk[81]) & (g358) & (g714)) + ((sk[81]) & (!g358) & (g714)));
	assign g713 = (((g358) & (!sk[82]) & (g717)));
	assign g714 = (((g715) & (!sk[83]) & (g716)) + ((!g715) & (sk[83]) & (!g716)));
	assign g715 = (((!sk[84]) & (i_4_) & (g719)) + ((sk[84]) & (!i_4_) & (g719)));
	assign g716 = (((i_4_) & (!sk[85]) & (g720)));
	assign g717 = (((i_4_) & (!sk[86]) & (g718)) + ((i_4_) & (sk[86]) & (!g718)));
	assign g718 = (((!sk[87]) & (i_4_) & (g721)));
	assign g719 = (((!sk[88]) & (i_3_) & (g119) & (!i_5_)) + ((!sk[88]) & (!i_3_) & (!g119) & (i_5_)) + ((sk[88]) & (!i_3_) & (!g119) & (!i_5_)) + ((!sk[88]) & (!i_3_) & (!g119) & (i_5_)));
	assign g720 = (((g21) & (sk[89]) & (!i_3_) & (!g138) & (!i_5_)) + ((g21) & (!sk[89]) & (i_3_) & (!g138) & (!i_5_)) + ((!g21) & (sk[89]) & (!i_3_) & (!g138) & (!i_5_)) + ((g21) & (!sk[89]) & (!i_3_) & (!g138) & (i_5_)) + ((!g21) & (sk[89]) & (!i_3_) & (!g138) & (i_5_)) + ((!g21) & (sk[89]) & (i_3_) & (!g138) & (!i_5_)));
	assign g721 = (((g21) & (i_3_) & (!g138) & (!sk[90]) & (!i_5_)) + ((g21) & (!i_3_) & (!g138) & (sk[90]) & (!i_5_)) + ((!g21) & (!i_3_) & (!g138) & (sk[90]) & (!i_5_)) + ((g21) & (!i_3_) & (!g138) & (!sk[90]) & (i_5_)) + ((!g21) & (!i_3_) & (!g138) & (sk[90]) & (i_5_)) + ((!g21) & (i_3_) & (!g138) & (sk[90]) & (!i_5_)));
	assign g722 = (((!sk[91]) & (i_9_) & (g723)) + ((sk[91]) & (i_9_) & (!g723)));
	assign g723 = (((i_9_) & (!sk[92]) & (g724)));
	assign g724 = (((g725) & (!sk[93]) & (g726)) + ((!g725) & (sk[93]) & (!g726)));
	assign g725 = (((!sk[94]) & (i_7_) & (g727)) + ((sk[94]) & (!i_7_) & (g727)));
	assign g726 = (((!sk[95]) & (i_7_) & (g728)));
	assign g727 = (((!sk[96]) & (i_6_) & (g142) & (!i_8_)) + ((!sk[96]) & (!i_6_) & (!g142) & (i_8_)) + ((sk[96]) & (!i_6_) & (!g142) & (!i_8_)) + ((!sk[96]) & (i_6_) & (!g142) & (i_8_)) + ((!sk[96]) & (!i_6_) & (g142) & (i_8_)));
	assign g728 = (((!g11) & (sk[97]) & (!i_6_) & (!g14) & (!i_8_)) + ((g11) & (!sk[97]) & (i_6_) & (!g14) & (!i_8_)) + ((!g11) & (sk[97]) & (!i_6_) & (!g14) & (!i_8_)) + ((g11) & (!sk[97]) & (!i_6_) & (!g14) & (i_8_)) + ((g11) & (!sk[97]) & (!i_6_) & (g14) & (i_8_)));
	assign g729 = (((!sk[98]) & (g280) & (g730)));
	assign g730 = (((!sk[99]) & (g731) & (g732)) + ((sk[99]) & (!g731) & (!g732)));
	assign g731 = (((!i_8_) & (sk[100]) & (g733)) + ((i_8_) & (!sk[100]) & (g733)));
	assign g732 = (((i_8_) & (!sk[101]) & (g734)));
	assign g733 = (((!sk[102]) & (g95) & (i_9_)) + ((sk[102]) & (!g95) & (!i_9_)));
	assign g734 = (((!sk[103]) & (g1) & (g68) & (!g14) & (!i_9_)) + ((sk[103]) & (!g1) & (!g68) & (!g14) & (!i_9_)) + ((sk[103]) & (!g1) & (!g68) & (g14) & (!i_9_)) + ((!sk[103]) & (g1) & (!g68) & (!g14) & (i_9_)) + ((sk[103]) & (!g1) & (!g68) & (!g14) & (!i_9_)));
	assign g735 = (((g736) & (!sk[104]) & (g737)) + ((!g736) & (sk[104]) & (!g737)));
	assign g736 = (((!sk[105]) & (g45) & (g738)) + ((sk[105]) & (!g45) & (g738)));
	assign g737 = (((g45) & (!sk[106]) & (g741)));
	assign g738 = (((g739) & (!sk[107]) & (g740)) + ((!g739) & (sk[107]) & (!g740)));
	assign g739 = (((!sk[108]) & (i_9_) & (g744)) + ((sk[108]) & (!i_9_) & (g744)));
	assign g740 = (((!sk[109]) & (i_9_) & (g745)));
	assign g741 = (((!sk[110]) & (g742) & (g743)) + ((sk[110]) & (!g742) & (!g743)));
	assign g742 = (((!i_9_) & (sk[111]) & (g746)) + ((i_9_) & (!sk[111]) & (g746)));
	assign g743 = (((!sk[112]) & (i_9_) & (g229)));
	assign g744 = (((g10) & (!g54) & (!sk[113]) & (!g1) & (g229)) + ((g10) & (g54) & (!sk[113]) & (!g1) & (!g229)) + ((!g10) & (g54) & (sk[113]) & (!g1) & (g229)) + ((!g10) & (!g54) & (sk[113]) & (g1) & (g229)));
	assign g745 = (((g10) & (!g39) & (!sk[114]) & (g229)) + ((!g10) & (!g39) & (!sk[114]) & (g229)) + ((!g10) & (!g39) & (!sk[114]) & (g229)) + ((g10) & (g39) & (!sk[114]) & (!g229)));
	assign g746 = (((g10) & (!g54) & (!g1) & (!sk[115]) & (g229)) + ((g10) & (g54) & (!g1) & (!sk[115]) & (!g229)) + ((!g10) & (g54) & (!g1) & (sk[115]) & (g229)) + ((!g10) & (!g54) & (g1) & (sk[115]) & (g229)));
	assign g747 = (((!sk[116]) & (g748) & (g749)) + ((sk[116]) & (!g748) & (!g749)));
	assign g748 = (((!sk[117]) & (g133) & (g750)) + ((sk[117]) & (!g133) & (g750)));
	assign g749 = (((g133) & (!sk[118]) & (g753)));
	assign g750 = (((!sk[119]) & (g751) & (g752)) + ((sk[119]) & (!g751) & (!g752)));
	assign g751 = (((!i_8_) & (sk[120]) & (g755)) + ((i_8_) & (!sk[120]) & (g755)));
	assign g752 = (((!sk[121]) & (i_8_) & (g756)));
	assign g753 = (((i_8_) & (!sk[122]) & (g754)) + ((!i_8_) & (sk[122]) & (!g754)));
	assign g754 = (((!sk[123]) & (i_8_) & (g757)) + ((sk[123]) & (!i_8_) & (g757)));
	assign g755 = (((!i_7_) & (!sk[124]) & (!i_6_) & (g28)) + ((!i_7_) & (sk[124]) & (!i_6_) & (!g28)) + ((i_7_) & (!sk[124]) & (i_6_) & (!g28)));
	assign g756 = (((!sk[125]) & (i_7_) & (i_6_) & (!g7) & (!g28)) + ((sk[125]) & (!i_7_) & (!i_6_) & (!g7) & (!g28)) + ((!sk[125]) & (i_7_) & (!i_6_) & (!g7) & (g28)) + ((sk[125]) & (!i_7_) & (i_6_) & (!g7) & (!g28)) + ((!sk[125]) & (i_7_) & (!i_6_) & (!g7) & (g28)));
	assign g757 = (((i_7_) & (i_6_) & (!sk[126]) & (!g13) & (!g28)) + ((!i_7_) & (!i_6_) & (sk[126]) & (!g13) & (!g28)) + ((!i_7_) & (!i_6_) & (sk[126]) & (g13) & (!g28)) + ((i_7_) & (!i_6_) & (!sk[126]) & (!g13) & (g28)));
	assign g758 = (((!sk[127]) & (i_2_) & (g759)) + ((sk[127]) & (i_2_) & (!g759)));
	assign g759 = (((!sk[0]) & (i_2_) & (g760)));
	assign g760 = (((g761) & (!sk[1]) & (g762)) + ((!g761) & (sk[1]) & (!g762)));
	assign g761 = (((!i_1_) & (sk[2]) & (g763)) + ((i_1_) & (!sk[2]) & (g763)));
	assign g762 = (((!sk[3]) & (i_1_) & (g764)));
	assign g763 = (((i_9_) & (!sk[4]) & (g37) & (!i_0_)) + ((!i_9_) & (!sk[4]) & (!g37) & (i_0_)) + ((!i_9_) & (sk[4]) & (!g37) & (!i_0_)) + ((i_9_) & (!sk[4]) & (!g37) & (i_0_)) + ((!i_9_) & (!sk[4]) & (g37) & (i_0_)));
	assign g764 = (((g50) & (i_9_) & (!sk[5]) & (!g76) & (!i_0_)) + ((!g50) & (i_9_) & (sk[5]) & (!g76) & (!i_0_)) + ((!g50) & (!i_9_) & (sk[5]) & (g76) & (!i_0_)) + ((g50) & (!i_9_) & (!sk[5]) & (!g76) & (i_0_)) + ((!g50) & (!i_9_) & (sk[5]) & (!g76) & (!i_0_)));
	assign g765 = (((!sk[6]) & (g766) & (g767)) + ((sk[6]) & (!g766) & (!g767)));
	assign g766 = (((!sk[7]) & (i_8_) & (g768)) + ((sk[7]) & (!i_8_) & (g768)));
	assign g767 = (((!sk[8]) & (i_8_) & (g770)));
	assign g768 = (((i_7_) & (!sk[9]) & (g769)) + ((!i_7_) & (sk[9]) & (!g769)));
	assign g769 = (((!sk[10]) & (i_7_) & (g772)) + ((sk[10]) & (!i_7_) & (g772)));
	assign g770 = (((i_7_) & (!sk[11]) & (g771)) + ((i_7_) & (sk[11]) & (!g771)));
	assign g771 = (((i_7_) & (!sk[12]) & (g773)));
	assign g772 = (((sk[13]) & (!i_9_) & (!g82) & (!i_6_)) + ((sk[13]) & (!i_9_) & (!g82) & (!i_6_)) + ((!sk[13]) & (!i_9_) & (!g82) & (i_6_)) + ((!sk[13]) & (i_9_) & (g82) & (!i_6_)));
	assign g773 = (((sk[14]) & (!g11) & (!i_9_) & (!g7) & (!i_6_)) + ((sk[14]) & (!g11) & (!i_9_) & (!g7) & (!i_6_)) + ((!sk[14]) & (g11) & (i_9_) & (!g7) & (!i_6_)) + ((!sk[14]) & (g11) & (!i_9_) & (!g7) & (i_6_)) + ((!sk[14]) & (g11) & (i_9_) & (!g7) & (!i_6_)));
	assign g774 = (((!sk[15]) & (g775) & (g776)) + ((sk[15]) & (!g775) & (!g776)));
	assign g775 = (((!sk[16]) & (g15) & (g777)) + ((sk[16]) & (!g15) & (g777)));
	assign g776 = (((g15) & (!sk[17]) & (g780)));
	assign g777 = (((!sk[18]) & (g778) & (g779)) + ((sk[18]) & (!g778) & (!g779)));
	assign g778 = (((!i_9_) & (sk[19]) & (g783)) + ((i_9_) & (!sk[19]) & (g783)));
	assign g779 = (((!sk[20]) & (i_9_) & (g784)));
	assign g780 = (((!sk[21]) & (g781) & (g782)) + ((sk[21]) & (!g781) & (!g782)));
	assign g781 = (((!i_9_) & (sk[22]) & (g785)) + ((i_9_) & (!sk[22]) & (g785)));
	assign g782 = (((i_9_) & (!sk[23]) & (g786)));
	assign g783 = (((i_1_) & (i_0_) & (!g17) & (!sk[24]) & (!i_2_)) + ((i_1_) & (!i_0_) & (!g17) & (sk[24]) & (!i_2_)) + ((!i_1_) & (i_0_) & (!g17) & (sk[24]) & (!i_2_)) + ((!i_1_) & (!i_0_) & (!g17) & (sk[24]) & (!i_2_)) + ((i_1_) & (!i_0_) & (!g17) & (!sk[24]) & (i_2_)) + ((!i_1_) & (!i_0_) & (!g17) & (sk[24]) & (i_2_)));
	assign g784 = (((sk[25]) & (!i_1_) & (!i_0_) & (!g19) & (!i_2_)) + ((!sk[25]) & (i_1_) & (i_0_) & (!g19) & (!i_2_)) + ((sk[25]) & (!i_1_) & (!i_0_) & (!g19) & (!i_2_)) + ((!sk[25]) & (i_1_) & (!i_0_) & (!g19) & (i_2_)) + ((!sk[25]) & (i_1_) & (!i_0_) & (!g19) & (i_2_)));
	assign g785 = (((i_1_) & (!sk[26]) & (!i_0_) & (!g17) & (i_2_)) + ((!i_1_) & (sk[26]) & (!i_0_) & (!g17) & (i_2_)) + ((!i_1_) & (sk[26]) & (i_0_) & (!g17) & (!i_2_)) + ((i_1_) & (!sk[26]) & (i_0_) & (!g17) & (!i_2_)) + ((i_1_) & (sk[26]) & (!i_0_) & (!g17) & (!i_2_)) + ((!i_1_) & (sk[26]) & (!i_0_) & (!g17) & (!i_2_)));
	assign g786 = (((sk[27]) & (!i_1_) & (!i_0_) & (!g19) & (!i_2_)) + ((!sk[27]) & (i_1_) & (i_0_) & (!g19) & (!i_2_)) + ((sk[27]) & (!i_1_) & (!i_0_) & (!g19) & (!i_2_)) + ((!sk[27]) & (i_1_) & (!i_0_) & (!g19) & (i_2_)) + ((!sk[27]) & (i_1_) & (!i_0_) & (!g19) & (i_2_)));
	assign g787 = (((!sk[28]) & (g788) & (g789)) + ((sk[28]) & (!g788) & (!g789)));
	assign g788 = (((!g1) & (sk[29]) & (g790)) + ((g1) & (!sk[29]) & (g790)));
	assign g789 = (((g1) & (!sk[30]) & (g793)));
	assign g790 = (((g791) & (!sk[31]) & (g792)) + ((!g791) & (sk[31]) & (!g792)));
	assign g791 = (((!sk[32]) & (i_9_) & (g796)) + ((sk[32]) & (!i_9_) & (g796)));
	assign g792 = (((!sk[33]) & (i_9_) & (g797)));
	assign g793 = (((g794) & (!sk[34]) & (g795)) + ((!g794) & (sk[34]) & (!g795)));
	assign g794 = (((!sk[35]) & (i_9_) & (g798)) + ((sk[35]) & (!i_9_) & (g798)));
	assign g795 = (((!sk[36]) & (i_9_) & (g799)));
	assign g796 = (((!sk[37]) & (g6) & (g4) & (!g9) & (!g3)) + ((!sk[37]) & (g6) & (!g4) & (!g9) & (g3)) + ((sk[37]) & (!g6) & (g4) & (!g9) & (!g3)) + ((sk[37]) & (!g6) & (!g4) & (!g9) & (g3)));
	assign g797 = (((sk[38]) & (g12) & (!g3)) + ((sk[38]) & (!g12) & (g3)) + ((!sk[38]) & (g12) & (g3)));
	assign g798 = (((!sk[39]) & (g6) & (g9)) + ((sk[39]) & (!g6) & (!g9)));
	assign g799 = (((sk[40]) & (g12) & (!g3)) + ((sk[40]) & (!g12) & (g3)) + ((!sk[40]) & (g12) & (g3)));

endmodule