module ks__aes_cipher_top_qmap_map (sk, ld, clk, rst, keyx0x, keyx1x, keyx2x, keyx3x, keyx4x, keyx5x, keyx6x, keyx7x, keyx8x, keyx9x, keyx10x, keyx11x, keyx12x, keyx13x, keyx14x, keyx15x, keyx16x, keyx17x, keyx18x, keyx19x, keyx20x, keyx21x, keyx22x, keyx23x, keyx24x, keyx25x, keyx26x, keyx27x, keyx28x, keyx29x, keyx30x, keyx31x, keyx32x, keyx33x, keyx34x, keyx35x, keyx36x, keyx37x, keyx38x, keyx39x, keyx40x, keyx41x, keyx42x, keyx43x, keyx44x, keyx45x, keyx46x, keyx47x, keyx48x, keyx49x, keyx50x, keyx51x, keyx52x, keyx53x, keyx54x, keyx55x, keyx56x, keyx57x, keyx58x, keyx59x, keyx60x, keyx61x, keyx62x, keyx63x, keyx64x, keyx65x, keyx66x, keyx67x, keyx68x, keyx69x, keyx70x, keyx71x, keyx72x, keyx73x, keyx74x, keyx75x, keyx76x, keyx77x, keyx78x, keyx79x, keyx80x, keyx81x, keyx82x, keyx83x, keyx84x, keyx85x, keyx86x, keyx87x, keyx88x, keyx89x, keyx90x, keyx91x, keyx92x, keyx93x, keyx94x, keyx95x, keyx96x, keyx97x, keyx98x, keyx99x, keyx100x, keyx101x, keyx102x, keyx103x, keyx104x, keyx105x, keyx106x, keyx107x, keyx108x, keyx109x, keyx110x, keyx111x, keyx112x, keyx113x, keyx114x, keyx115x, keyx116x, keyx117x, keyx118x, keyx119x, keyx120x, keyx121x, keyx122x, keyx123x, keyx124x, keyx125x, keyx126x, keyx127x, text_inx32x, text_inx33x, text_inx34x, text_inx35x, text_inx38x, text_inx37x, text_inx36x, text_inx39x, text_inx72x, text_inx73x, text_inx74x, text_inx75x, text_inx78x, text_inx77x, text_inx76x, text_inx79x, text_inx112x, text_inx113x, text_inx114x, text_inx115x, text_inx118x, text_inx117x, text_inx116x, text_inx119x, text_inx24x, text_inx25x, text_inx26x, text_inx27x, text_inx30x, text_inx29x, text_inx28x, text_inx31x, text_inx64x, text_inx65x, text_inx66x, text_inx67x, text_inx70x, text_inx69x, text_inx68x, text_inx71x, text_inx104x, text_inx105x, text_inx106x, text_inx107x, text_inx110x, text_inx109x, text_inx108x, text_inx111x, text_inx16x, text_inx17x, text_inx18x, text_inx19x, text_inx22x, text_inx21x, text_inx20x, text_inx23x, text_inx56x, text_inx57x, text_inx58x, text_inx59x, text_inx62x, text_inx61x, text_inx60x, text_inx63x, text_inx96x, text_inx97x, text_inx98x, text_inx99x, text_inx102x, text_inx101x, text_inx100x, text_inx103x, text_inx8x, text_inx9x, text_inx10x, text_inx11x, text_inx14x, text_inx13x, text_inx12x, text_inx15x, text_inx48x, text_inx49x, text_inx50x, text_inx51x, text_inx54x, text_inx53x, text_inx52x, text_inx55x, text_inx88x, text_inx89x, text_inx90x, text_inx91x, text_inx94x, text_inx93x, text_inx92x, text_inx95x, text_inx0x, text_inx1x, text_inx2x, text_inx3x, text_inx6x, text_inx5x, text_inx4x, text_inx7x, text_inx40x, text_inx41x, text_inx42x, text_inx43x, text_inx46x, text_inx45x, text_inx44x, text_inx47x, text_inx80x, text_inx81x, text_inx82x, text_inx83x, text_inx86x, text_inx85x, text_inx84x, text_inx87x, text_inx120x, text_inx121x, text_inx122x, text_inx123x, text_inx126x, text_inx125x, text_inx124x, text_inx127x, done, text_outx0x, text_outx1x, text_outx2x, text_outx3x, text_outx4x, text_outx5x, text_outx6x, text_outx7x, text_outx8x, text_outx9x, text_outx10x, text_outx11x, text_outx12x, text_outx13x, text_outx14x, text_outx15x, text_outx16x, text_outx17x, text_outx18x, text_outx19x, text_outx20x, text_outx21x, text_outx22x, text_outx23x, text_outx24x, text_outx25x, text_outx26x, text_outx27x, text_outx28x, text_outx29x, text_outx30x, text_outx31x, text_outx32x, text_outx33x, text_outx34x, text_outx35x, text_outx36x, text_outx37x, text_outx38x, text_outx39x, text_outx40x, text_outx41x, text_outx42x, text_outx43x, text_outx44x, text_outx45x, text_outx46x, text_outx47x, text_outx48x, text_outx49x, text_outx50x, text_outx51x, text_outx52x, text_outx53x, text_outx54x, text_outx55x, text_outx56x, text_outx57x, text_outx58x, text_outx59x, text_outx60x, text_outx61x, text_outx62x, text_outx63x, text_outx64x, text_outx65x, text_outx66x, text_outx67x, text_outx68x, text_outx69x, text_outx70x, text_outx71x, text_outx72x, text_outx73x, text_outx74x, text_outx75x, text_outx76x, text_outx77x, text_outx78x, text_outx79x, text_outx80x, text_outx81x, text_outx82x, text_outx83x, text_outx84x, text_outx85x, text_outx86x, text_outx87x, text_outx88x, text_outx89x, text_outx90x, text_outx91x, text_outx92x, text_outx93x, text_outx94x, text_outx95x, text_outx96x, text_outx97x, text_outx98x, text_outx99x, text_outx100x, text_outx101x, text_outx102x, text_outx103x, text_outx104x, text_outx105x, text_outx106x, text_outx107x, text_outx108x, text_outx109x, text_outx110x, text_outx111x, text_outx112x, text_outx113x, text_outx114x, text_outx115x, text_outx116x, text_outx117x, text_outx118x, text_outx119x, text_outx120x, text_outx121x, text_outx122x, text_outx123x, text_outx124x, text_outx125x, text_outx126x, text_outx127x);

	input ld;
	input clk;
	input rst;
	input keyx0x;
	input keyx1x;
	input keyx2x;
	input keyx3x;
	input keyx4x;
	input keyx5x;
	input keyx6x;
	input keyx7x;
	input keyx8x;
	input keyx9x;
	input keyx10x;
	input keyx11x;
	input keyx12x;
	input keyx13x;
	input keyx14x;
	input keyx15x;
	input keyx16x;
	input keyx17x;
	input keyx18x;
	input keyx19x;
	input keyx20x;
	input keyx21x;
	input keyx22x;
	input keyx23x;
	input keyx24x;
	input keyx25x;
	input keyx26x;
	input keyx27x;
	input keyx28x;
	input keyx29x;
	input keyx30x;
	input keyx31x;
	input keyx32x;
	input keyx33x;
	input keyx34x;
	input keyx35x;
	input keyx36x;
	input keyx37x;
	input keyx38x;
	input keyx39x;
	input keyx40x;
	input keyx41x;
	input keyx42x;
	input keyx43x;
	input keyx44x;
	input keyx45x;
	input keyx46x;
	input keyx47x;
	input keyx48x;
	input keyx49x;
	input keyx50x;
	input keyx51x;
	input keyx52x;
	input keyx53x;
	input keyx54x;
	input keyx55x;
	input keyx56x;
	input keyx57x;
	input keyx58x;
	input keyx59x;
	input keyx60x;
	input keyx61x;
	input keyx62x;
	input keyx63x;
	input keyx64x;
	input keyx65x;
	input keyx66x;
	input keyx67x;
	input keyx68x;
	input keyx69x;
	input keyx70x;
	input keyx71x;
	input keyx72x;
	input keyx73x;
	input keyx74x;
	input keyx75x;
	input keyx76x;
	input keyx77x;
	input keyx78x;
	input keyx79x;
	input keyx80x;
	input keyx81x;
	input keyx82x;
	input keyx83x;
	input keyx84x;
	input keyx85x;
	input keyx86x;
	input keyx87x;
	input keyx88x;
	input keyx89x;
	input keyx90x;
	input keyx91x;
	input keyx92x;
	input keyx93x;
	input keyx94x;
	input keyx95x;
	input keyx96x;
	input keyx97x;
	input keyx98x;
	input keyx99x;
	input keyx100x;
	input keyx101x;
	input keyx102x;
	input keyx103x;
	input keyx104x;
	input keyx105x;
	input keyx106x;
	input keyx107x;
	input keyx108x;
	input keyx109x;
	input keyx110x;
	input keyx111x;
	input keyx112x;
	input keyx113x;
	input keyx114x;
	input keyx115x;
	input keyx116x;
	input keyx117x;
	input keyx118x;
	input keyx119x;
	input keyx120x;
	input keyx121x;
	input keyx122x;
	input keyx123x;
	input keyx124x;
	input keyx125x;
	input keyx126x;
	input keyx127x;
	input text_inx32x;
	input text_inx33x;
	input text_inx34x;
	input text_inx35x;
	input text_inx38x;
	input text_inx37x;
	input text_inx36x;
	input text_inx39x;
	input text_inx72x;
	input text_inx73x;
	input text_inx74x;
	input text_inx75x;
	input text_inx78x;
	input text_inx77x;
	input text_inx76x;
	input text_inx79x;
	input text_inx112x;
	input text_inx113x;
	input text_inx114x;
	input text_inx115x;
	input text_inx118x;
	input text_inx117x;
	input text_inx116x;
	input text_inx119x;
	input text_inx24x;
	input text_inx25x;
	input text_inx26x;
	input text_inx27x;
	input text_inx30x;
	input text_inx29x;
	input text_inx28x;
	input text_inx31x;
	input text_inx64x;
	input text_inx65x;
	input text_inx66x;
	input text_inx67x;
	input text_inx70x;
	input text_inx69x;
	input text_inx68x;
	input text_inx71x;
	input text_inx104x;
	input text_inx105x;
	input text_inx106x;
	input text_inx107x;
	input text_inx110x;
	input text_inx109x;
	input text_inx108x;
	input text_inx111x;
	input text_inx16x;
	input text_inx17x;
	input text_inx18x;
	input text_inx19x;
	input text_inx22x;
	input text_inx21x;
	input text_inx20x;
	input text_inx23x;
	input text_inx56x;
	input text_inx57x;
	input text_inx58x;
	input text_inx59x;
	input text_inx62x;
	input text_inx61x;
	input text_inx60x;
	input text_inx63x;
	input text_inx96x;
	input text_inx97x;
	input text_inx98x;
	input text_inx99x;
	input text_inx102x;
	input text_inx101x;
	input text_inx100x;
	input text_inx103x;
	input text_inx8x;
	input text_inx9x;
	input text_inx10x;
	input text_inx11x;
	input text_inx14x;
	input text_inx13x;
	input text_inx12x;
	input text_inx15x;
	input text_inx48x;
	input text_inx49x;
	input text_inx50x;
	input text_inx51x;
	input text_inx54x;
	input text_inx53x;
	input text_inx52x;
	input text_inx55x;
	input text_inx88x;
	input text_inx89x;
	input text_inx90x;
	input text_inx91x;
	input text_inx94x;
	input text_inx93x;
	input text_inx92x;
	input text_inx95x;
	input text_inx0x;
	input text_inx1x;
	input text_inx2x;
	input text_inx3x;
	input text_inx6x;
	input text_inx5x;
	input text_inx4x;
	input text_inx7x;
	input text_inx40x;
	input text_inx41x;
	input text_inx42x;
	input text_inx43x;
	input text_inx46x;
	input text_inx45x;
	input text_inx44x;
	input text_inx47x;
	input text_inx80x;
	input text_inx81x;
	input text_inx82x;
	input text_inx83x;
	input text_inx86x;
	input text_inx85x;
	input text_inx84x;
	input text_inx87x;
	input text_inx120x;
	input text_inx121x;
	input text_inx122x;
	input text_inx123x;
	input text_inx126x;
	input text_inx125x;
	input text_inx124x;
	input text_inx127x;
	output done;
	output text_outx0x;
	output text_outx1x;
	output text_outx2x;
	output text_outx3x;
	output text_outx4x;
	output text_outx5x;
	output text_outx6x;
	output text_outx7x;
	output text_outx8x;
	output text_outx9x;
	output text_outx10x;
	output text_outx11x;
	output text_outx12x;
	output text_outx13x;
	output text_outx14x;
	output text_outx15x;
	output text_outx16x;
	output text_outx17x;
	output text_outx18x;
	output text_outx19x;
	output text_outx20x;
	output text_outx21x;
	output text_outx22x;
	output text_outx23x;
	output text_outx24x;
	output text_outx25x;
	output text_outx26x;
	output text_outx27x;
	output text_outx28x;
	output text_outx29x;
	output text_outx30x;
	output text_outx31x;
	output text_outx32x;
	output text_outx33x;
	output text_outx34x;
	output text_outx35x;
	output text_outx36x;
	output text_outx37x;
	output text_outx38x;
	output text_outx39x;
	output text_outx40x;
	output text_outx41x;
	output text_outx42x;
	output text_outx43x;
	output text_outx44x;
	output text_outx45x;
	output text_outx46x;
	output text_outx47x;
	output text_outx48x;
	output text_outx49x;
	output text_outx50x;
	output text_outx51x;
	output text_outx52x;
	output text_outx53x;
	output text_outx54x;
	output text_outx55x;
	output text_outx56x;
	output text_outx57x;
	output text_outx58x;
	output text_outx59x;
	output text_outx60x;
	output text_outx61x;
	output text_outx62x;
	output text_outx63x;
	output text_outx64x;
	output text_outx65x;
	output text_outx66x;
	output text_outx67x;
	output text_outx68x;
	output text_outx69x;
	output text_outx70x;
	output text_outx71x;
	output text_outx72x;
	output text_outx73x;
	output text_outx74x;
	output text_outx75x;
	output text_outx76x;
	output text_outx77x;
	output text_outx78x;
	output text_outx79x;
	output text_outx80x;
	output text_outx81x;
	output text_outx82x;
	output text_outx83x;
	output text_outx84x;
	output text_outx85x;
	output text_outx86x;
	output text_outx87x;
	output text_outx88x;
	output text_outx89x;
	output text_outx90x;
	output text_outx91x;
	output text_outx92x;
	output text_outx93x;
	output text_outx94x;
	output text_outx95x;
	output text_outx96x;
	output text_outx97x;
	output text_outx98x;
	output text_outx99x;
	output text_outx100x;
	output text_outx101x;
	output text_outx102x;
	output text_outx103x;
	output text_outx104x;
	output text_outx105x;
	output text_outx106x;
	output text_outx107x;
	output text_outx108x;
	output text_outx109x;
	output text_outx110x;
	output text_outx111x;
	output text_outx112x;
	output text_outx113x;
	output text_outx114x;
	output text_outx115x;
	output text_outx116x;
	output text_outx117x;
	output text_outx118x;
	output text_outx119x;
	output text_outx120x;
	output text_outx121x;
	output text_outx122x;
	output text_outx123x;
	output text_outx124x;
	output text_outx125x;
	output text_outx126x;
	output text_outx127x;

	input [127 : 0] sk /* synthesis noprune */;


	wire g134, g141, g142, g143, g144, g147, g149, g150, g151, g152, g153;
	wire g154, g156, g157, g158, g159, g160, g161, g163, g164, g165, g166;
	wire g167, g168, g170, g171, g172, g173, g174, g175, g177, g178, g179;
	wire g180, g181, g182, g184, g185, g186, g187, g188, g189, g191, g192;
	wire g193, g194, g195, g196, g198, g205, g206, g207, g208, g211, g213;
	wire g214, g215, g216, g217, g218, g220, g221, g222, g223, g224, g225;
	wire g227, g228, g229, g230, g231, g232, g234, g235, g236, g237, g238;
	wire g239, g241, g242, g243, g244, g245, g246, g248, g249, g250, g251;
	wire g252, g253, g255, g256, g257, g258, g259, g260, g262, g269, g270;
	wire g271, g272, g275, g277, g278, g279, g280, g281, g282, g284, g285;
	wire g286, g287, g288, g289, g291, g292, g293, g294, g295, g296, g298;
	wire g299, g300, g301, g302, g303, g305, g306, g307, g308, g309, g310;
	wire g312, g313, g314, g315, g316, g317, g319, g320, g321, g322, g323;
	wire g324, g326, g333, g334, g335, g336, g339, g341, g342, g343, g344;
	wire g345, g346, g348, g349, g350, g351, g352, g353, g355, g356, g357;
	wire g358, g359, g360, g362, g363, g364, g365, g366, g367, g369, g370;
	wire g371, g372, g373, g374, g376, g377, g378, g379, g380, g381, g383;
	wire g384, g385, g386, g387, g388, g390, g397, g398, g399, g400, g403;
	wire g405, g406, g407, g408, g409, g410, g412, g413, g414, g415, g416;
	wire g417, g419, g420, g421, g422, g423, g424, g426, g427, g428, g429;
	wire g430, g431, g433, g434, g435, g436, g437, g438, g440, g441, g442;
	wire g443, g444, g445, g447, g448, g449, g450, g451, g452, g454, g461;
	wire g462, g463, g464, g467, g469, g470, g471, g472, g473, g474, g476;
	wire g477, g478, g479, g480, g481, g483, g484, g485, g486, g487, g488;
	wire g490, g491, g492, g493, g494, g495, g497, g498, g499, g500, g501;
	wire g502, g504, g505, g506, g507, g508, g509, g511, g512, g513, g514;
	wire g515, g516, g518, g525, g526, g527, g528, g531, g533, g534, g535;
	wire g536, g537, g538, g540, g541, g542, g543, g544, g545, g547, g548;
	wire g549, g550, g551, g552, g554, g555, g556, g557, g558, g559, g561;
	wire g562, g563, g564, g565, g566, g568, g569, g570, g571, g572, g573;
	wire g575, g576, g577, g578, g579, g580, g582, g589, g590, g591, g592;
	wire g595, g597, g598, g599, g600, g601, g602, g604, g605, g606, g607;
	wire g608, g609, g611, g612, g613, g614, g615, g616, g618, g619, g620;
	wire g621, g622, g623, g625, g626, g627, g628, g629, g630, g632, g633;
	wire g634, g635, g636, g637, g639, g640, g641, g642, g643, g644, g646;
	wire g653, g654, g655, g656, g659, g661, g662, g663, g664, g665, g666;
	wire g668, g669, g670, g671, g672, g673, g675, g676, g677, g678, g679;
	wire g680, g682, g683, g684, g685, g686, g687, g689, g690, g691, g692;
	wire g693, g694, g696, g697, g698, g699, g700, g701, g703, g704, g705;
	wire g706, g707, g708, g710, g717, g718, g719, g720, g723, g725, g726;
	wire g727, g728, g729, g730, g732, g733, g734, g735, g736, g737, g739;
	wire g740, g741, g742, g743, g744, g746, g747, g748, g749, g750, g751;
	wire g753, g754, g755, g756, g757, g758, g760, g761, g762, g763, g764;
	wire g765, g767, g768, g769, g770, g771, g772, g774, g781, g782, g783;
	wire g784, g787, g789, g790, g791, g792, g793, g794, g796, g797, g798;
	wire g799, g800, g801, g803, g804, g805, g806, g807, g808, g810, g811;
	wire g812, g813, g814, g815, g817, g818, g819, g820, g821, g822, g824;
	wire g825, g826, g827, g828, g829, g831, g832, g833, g834, g835, g836;
	wire g838, g845, g846, g847, g848, g851, g853, g854, g855, g856, g857;
	wire g858, g860, g861, g862, g863, g864, g865, g867, g868, g869, g870;
	wire g871, g872, g874, g875, g876, g877, g878, g879, g881, g882, g883;
	wire g884, g885, g886, g888, g889, g890, g891, g892, g893, g895, g896;
	wire g897, g898, g899, g900, g902, g909, g910, g911, g912, g915, g917;
	wire g918, g919, g920, g921, g922, g924, g925, g926, g927, g928, g929;
	wire g931, g932, g933, g934, g935, g936, g938, g939, g940, g941, g942;
	wire g943, g945, g946, g947, g948, g949, g950, g952, g953, g954, g955;
	wire g956, g957, g959, g960, g961, g962, g963, g964, g966, g973, g974;
	wire g975, g976, g979, g981, g982, g983, g984, g985, g986, g988, g989;
	wire g990, g991, g992, g993, g995, g996, g997, g998, g999, g1000, g1002;
	wire g1003, g1004, g1005, g1006, g1007, g1009, g1010, g1011, g1012, g1013, g1014;
	wire g1016, g1017, g1018, g1019, g1020, g1021, g1023, g1024, g1025, g1026, g1027;
	wire g1028, g1030, g1037, g1038, g1039, g1040, g1043, g1045, g1046, g1047, g1048;
	wire g1049, g1050, g1052, g1053, g1054, g1055, g1056, g1057, g1059, g1060, g1061;
	wire g1062, g1063, g1064, g1066, g1067, g1068, g1069, g1070, g1071, g1073, g1074;
	wire g1075, g1076, g1077, g1078, g1080, g1081, g1082, g1083, g1084, g1085, g1087;
	wire g1088, g1089, g1090, g1091, g1092, g1094, g1101, g1102, g1103, g1104, g1107;
	wire g1109, g1110, g1111, g1112, g1113, g1114, g1116, g1117, g1118, g1119, g1120;
	wire g1121, g1123, g1124, g1125, g1126, g1127, g1128, g1130, g1131, g1132, g1133;
	wire g1134, g1135, g1137, g1138, g1139, g1140, g1141, g1142, g1144, g1145, g1146;
	wire g1147, g1148, g1149, g1151, g1152, g1153, g1154, g1155, g1156, g1158, g1159;
	wire g1160, g1161, g1162, g2082, g1165, g1166, g2083, g1168, g1169, g1170, g2084;
	wire g1172, g1173, g2085, g1175, g2086, g1177, g1178, g2087, g1180, g1181, g2088;
	wire g1183, g1184, g1185, g2089, g1187, g1188, g1189, g1190, g1191, g1192, g1193;
	wire g1194, g1195, g1196, g1197, g1198, g1199, g1200, g1201, g1202, g1203, g1204;
	wire g1205, g1206, g1207, g1208, g1209, g1210, g1211, g1212, g1213, g1214, g1215;
	wire g1216, g1217, g1218, g1219, g1220, g1221, g1222, g1223, g1224, g1225, g1226;
	wire g1227, g1228, g1229, g1230, g1231, g1232, g1233, g1234, g1235, g1236, g1237;
	wire g1238, g1239, g1240, g1241, g1242, g1243, g1244, g2090, g1246, g1247, g1248;
	wire g2091, g1250, g1251, g1252, g2092, g1254, g1255, g2093, g1257, g1258, g2094;
	wire g1260, g1261, g2095, g1263, g1264, g2096, g1266, g1267, g2097, g1269, g1270;
	wire g1271, g1272, g1273, g1274, g1275, g1276, g1277, g1278, g1279, g1280, g1281;
	wire g1282, g1283, g1284, g1285, g1286, g1287, g1288, g1289, g1290, g1291, g1292;
	wire g1293, g1294, g1295, g1296, g1297, g1298, g1299, g1300, g1301, g1302, g1303;
	wire g1304, g1305, g1306, g1307, g1308, g1309, g1310, g1311, g1312, g1313, g1314;
	wire g1315, g1316, g1317, g1318, g1319, g1320, g1321, g1322, g1323, g1324, g1325;
	wire g1326, g1327, g2098, g1329, g1330, g1331, g2099, g1333, g1334, g1335, g2100;
	wire g1337, g1338, g2101, g1340, g2102, g1342, g1343, g2103, g1345, g1346, g2104;
	wire g1348, g1349, g1350, g2105, g1352, g1353, g1354, g1355, g1356, g1357, g1358;
	wire g1359, g1360, g1361, g1362, g1363, g1364, g1365, g1366, g1367, g1368, g1369;
	wire g1370, g1371, g1372, g1373, g1374, g1375, g1376, g1377, g1378, g1379, g1380;
	wire g1381, g1382, g1383, g1384, g1385, g1386, g1387, g1388, g1389, g1390, g1391;
	wire g1392, g1393, g1394, g1395, g1396, g1397, g1398, g1399, g1400, g1401, g1402;
	wire g1403, g1404, g1405, g1406, g1407, g1408, g1409, g2106, g1411, g1412, g1413;
	wire g2107, g1415, g2108, g1417, g1418, g2109, g1420, g1421, g2110, g1423, g1424;
	wire g2111, g1426, g1427, g2112, g1429, g2113, g1431, g1432, g1433, g1434, g1435;
	wire g1436, g1437, g1438, g1440, g1441, g1442, g1443, g1444, g1445, g1446, g1447;
	wire g1449, g1450, g1451, g1452, g1453, g1454, g1455, g1456, g1458, g1459, g1460;
	wire g1461, g1462, g1463, g1464, g1465, g1467, g1468, g1469, g1470, g1471, g1472;
	wire g1473, g1474, g1476, g1477, g1478, g1479, g1480, g1481, g1482, g1483, g1485;
	wire g1486, g1487, g1488, g1489, g1490, g1491, g1492, g1494, g1495, g1496, g1497;
	wire g1498, g1499, g1500, g1501, g1503, g1504, g1505, g2114, g1507, g2115, g1509;
	wire g1510, g2116, g1512, g2117, g1514, g2118, g1516, g2119, g1518, g2120, g1520;
	wire g1521, g2121, g1523, g1524, g1525, g1526, g1527, g1528, g1529, g1530, g1531;
	wire g1532, g2122, g1534, g1535, g2123, g1537, g1538, g1539, g2124, g1541, g1542;
	wire g2125, g1544, g1545, g1546, g2126, g1548, g1549, g2127, g1551, g1552, g2128;
	wire g1554, g2129, g1556, g1557, g1558, g1559, g1560, g1561, g1562, g1563, g1564;
	wire g2130, g1566, g1567, g2131, g2132, g1570, g2133, g1572, g1573, g2134, g1575;
	wire g2135, g1577, g2136, g2137, g1580, g1581, g1582, g1583, g1584, g1585, g1586;
	wire g1587, g2138, g1589, g1590, g2139, g1592, g2140, g1594, g1595, g2141, g2142;
	wire g1598, g1599, g2143, g1601, g1602, g2144, g1604, g1605, g1606, g2145, g1608;
	wire g1609, g1610, g1611, g1612, g1613, g1614, g1615, g1616, g1617, g1618, g2146;
	wire g1620, g2147, g1622, g1623, g1624, g2148, g1626, g2149, g1628, g1629, g2150;
	wire g1631, g2151, g1633, g2152, g1635, g2153, g1637, g1638, g1639, g1640, g1641;
	wire g1642, g1643, g1644, g2154, g2155, g1647, g1648, g1649, g2156, g1651, g1652;
	wire g2157, g1654, g1655, g1656, g2158, g1658, g1659, g2159, g1661, g1662, g2160;
	wire g1664, g1665, g1666, g2161, g1668, g1669, g1670, g1671, g1672, g1673, g1674;
	wire g1675, g1676, g1677, g2162, g1679, g1680, g2163, g1682, g2164, g1684, g2165;
	wire g1686, g1687, g1688, g2166, g1690, g2167, g1692, g2168, g1694, g1695, g2169;
	wire g1697, g1698, g1699, g1700, g1701, g1702, g1703, g1704, g1705, g2170, g1707;
	wire g1708, g2171, g1710, g1711, g2172, g1713, g1714, g2173, g1716, g1717, g2174;
	wire g1719, g1720, g2175, g1722, g1723, g2176, g1725, g1726, g1727, g1728, g2177;
	wire g1730, g1731, g1732, g1733, g1734, g1735, g1736, g1737, g1738, g2178, g1740;
	wire g1741, g2179, g1743, g2180, g1745, g2181, g1747, g1748, g2182, g1750, g2183;
	wire g1752, g2184, g1754, g1755, g2185, g1757, g1758, g1759, g1760, g1761, g1762;
	wire g1763, g1764, g2186, g1766, g1767, g2187, g2188, g1770, g2189, g1772, g1773;
	wire g2190, g1775, g2191, g1777, g2192, g1779, g1780, g2193, g1782, g1783, g1784;
	wire g1785, g1786, g1787, g1788, g1789, g1790, g2194, g1792, g1793, g2195, g1795;
	wire g1796, g2196, g1798, g2197, g1800, g1801, g2198, g1803, g2199, g1805, g2200;
	wire g1807, g1808, g2201, g1810, g1811, g1812, g1813, g1814, g1815, g1816, g1817;
	wire g2202, g1819, g1820, g2203, g1822, g2204, g1824, g2205, g2206, g1827, g2207;
	wire g1829, g2208, g1831, g2209, g1833, g1834, g1835, g1836, g1837, g1838, g1839;
	wire g1840, g1841, g1845, g1847, g1848, g1849, g1850, g1851, g1852, g1853, g1854;
	wire g1855, g1856, g1857, g1859, g1860, g1858, g1861, g1864, g1862, g1863, g1867;
	wire g1868, g1865, g1866, g1869, g1870, g1872, g1873, g1871, g1874, g1877, g1875;
	wire g1876, g1880, g1881, g1878, g1879, g1882, g1883, g1885, g1886, g1884, g1887;
	wire g1890, g1888, g1889, g1893, g1891, g1892, g1894, g1896, g1897, g1895, g1898;
	wire g1901, g1899, g1900, g1904, g1905, g1902, g1903, g1906, g1907, g1909, g1910;
	wire g1908, g1911, g1914, g1912, g1913, g1917, g1915, g1916, g1918, g1920, g1921;
	wire g1919, g1922, g1925, g1923, g1924, g1928, g1929, g1926, g1927, g1930, g1931;
	wire g1933, g1934, g1932, g1935, g1938, g1936, g1937, g1941, g1939, g1940, g1942;
	wire g1944, g1945, g1943, g1946, g1949, g1947, g1948, g1952, g1950, g1951, g1953;
	wire g1955, g1956, g1954, g1957, g1960, g1958, g1959, g1963, g1964, g1961, g1962;
	wire g1965, g1966, g1968, g1969, g1967, g1970, g1973, g1971, g1972, g1976, g1977;
	wire g1974, g1975, g1978, g1979, g1981, g1982, g1980, g1983, g1986, g1984, g1985;
	wire g1989, g1987, g1988, g1990, g1992, g1993, g1991, g1994, g1997, g1995, g1996;
	wire g2000, g2001, g1998, g1999, g2002, g2003, g2005, g2006, g2004, g2007, g2010;
	wire g2008, g2009, g2013, g2014, g2011, g2012, g2015, g2016, g2018, g2019, g2017;
	wire g2020, g2023, g2021, g2022, g2026, g2027, g2024, g2025, g2028, g2029, g2031;
	wire g2032, g2030, g2033, g2036, g2034, g2035, g2039, g2040, g2037, g2038, g2041;
	wire g2042, g2044, g2045, g2043, g2046, g2049, g2047, g2048, g2052, g2053, g2050;
	wire g2051, g2054, g2055, g2057, g2058, g2056, g2059, g2062, g2060, g2061, g2065;
	wire g2066, g2063, g2064, g2067, g2068, g2070, g2071, g2069, g2072, g2075, g2073;
	wire g2074, g2078, g2079, g2076, g2077, g2080, g2081;


	reg done, text_outx0x, text_outx1x, text_outx2x, text_outx3x, text_outx4x, text_outx5x, text_outx6x, text_outx7x;
	reg text_outx8x, text_outx9x, text_outx10x, text_outx11x, text_outx12x, text_outx13x, text_outx14x, text_outx15x, text_outx16x;
	reg text_outx17x, text_outx18x, text_outx19x, text_outx20x, text_outx21x, text_outx22x, text_outx23x, text_outx24x, text_outx25x;
	reg text_outx26x, text_outx27x, text_outx28x, text_outx29x, text_outx30x, text_outx31x, text_outx32x, text_outx33x, text_outx34x;
	reg text_outx35x, text_outx36x, text_outx37x, text_outx38x, text_outx39x, text_outx40x, text_outx41x, text_outx42x, text_outx43x;
	reg text_outx44x, text_outx45x, text_outx46x, text_outx47x, text_outx48x, text_outx49x, text_outx50x, text_outx51x, text_outx52x;
	reg text_outx53x, text_outx54x, text_outx55x, text_outx56x, text_outx57x, text_outx58x, text_outx59x, text_outx60x, text_outx61x;
	reg text_outx62x, text_outx63x, text_outx64x, text_outx65x, text_outx66x, text_outx67x, text_outx68x, text_outx69x, text_outx70x;
	reg text_outx71x, text_outx72x, text_outx73x, text_outx74x, text_outx75x, text_outx76x, text_outx77x, text_outx78x, text_outx79x;
	reg text_outx80x, text_outx81x, text_outx82x, text_outx83x, text_outx84x, text_outx85x, text_outx86x, text_outx87x, text_outx88x;
	reg text_outx89x, text_outx90x, text_outx91x, text_outx92x, text_outx93x, text_outx94x, text_outx95x, text_outx96x, text_outx97x;
	reg text_outx98x, text_outx99x, text_outx100x, text_outx101x, text_outx102x, text_outx103x, text_outx104x, text_outx105x, text_outx106x;
	reg text_outx107x, text_outx108x, text_outx109x, text_outx110x, text_outx111x, text_outx112x, text_outx113x, text_outx114x, text_outx115x;
	reg text_outx116x, text_outx117x, text_outx118x, text_outx119x, text_outx120x, text_outx121x, text_outx122x, text_outx123x, text_outx124x;
	reg text_outx125x, text_outx126x, text_outx127x, g130, g131, g132, g133, g135, g136;
	reg g137, g138, g139, g140, g145, g146, g148, g155, g162;
	reg g169, g176, g183, g190, g197, g199, g200, g201, g202;
	reg g203, g204, g209, g210, g212, g219, g226, g233, g240;
	reg g247, g254, g261, g263, g264, g265, g266, g267, g268;
	reg g273, g274, g276, g283, g290, g297, g304, g311, g318;
	reg g325, g327, g328, g329, g330, g331, g332, g337, g338;
	reg g340, g347, g354, g361, g368, g375, g382, g389, g391;
	reg g392, g393, g394, g395, g396, g401, g402, g404, g411;
	reg g418, g425, g432, g439, g446, g453, g455, g456, g457;
	reg g458, g459, g460, g465, g466, g468, g475, g482, g489;
	reg g496, g503, g510, g517, g519, g520, g521, g522, g523;
	reg g524, g529, g530, g532, g539, g546, g553, g560, g567;
	reg g574, g581, g583, g584, g585, g586, g587, g588, g593;
	reg g594, g596, g603, g610, g617, g624, g631, g638, g645;
	reg g647, g648, g649, g650, g651, g652, g657, g658, g660;
	reg g667, g674, g681, g688, g695, g702, g709, g711, g712;
	reg g713, g714, g715, g716, g721, g722, g724, g731, g738;
	reg g745, g752, g759, g766, g773, g775, g776, g777, g778;
	reg g779, g780, g785, g786, g788, g795, g802, g809, g816;
	reg g823, g830, g837, g839, g840, g841, g842, g843, g844;
	reg g849, g850, g852, g859, g866, g873, g880, g887, g894;
	reg g901, g903, g904, g905, g906, g907, g908, g913, g914;
	reg g916, g923, g930, g937, g944, g951, g958, g965, g967;
	reg g968, g969, g970, g971, g972, g977, g978, g980, g987;
	reg g994, g1001, g1008, g1015, g1022, g1029, g1031, g1032, g1033;
	reg g1034, g1035, g1036, g1041, g1042, g1044, g1051, g1058, g1065;
	reg g1072, g1079, g1086, g1093, g1095, g1096, g1097, g1098, g1099;
	reg g1100, g1105, g1106, g1108, g1115, g1122, g1129, g1136, g1143;
	reg g1150, g1157, g1163, g1164, g1167, g1171, g1174, g1176, g1179;
	reg g1182, g1186, g1245, g1249, g1253, g1256, g1259, g1262, g1265;
	reg g1268, g1328, g1332, g1336, g1339, g1341, g1344, g1347, g1351;
	reg g1410, g1414, g1416, g1419, g1422, g1425, g1428, g1430, g1439;
	reg g1448, g1457, g1466, g1475, g1484, g1493, g1502, g1506, g1508;
	reg g1511, g1513, g1515, g1517, g1519, g1522, g1533, g1536, g1540;
	reg g1543, g1547, g1550, g1553, g1555, g1565, g1568, g1569, g1571;
	reg g1574, g1576, g1578, g1579, g1588, g1591, g1593, g1596, g1597;
	reg g1600, g1603, g1607, g1619, g1621, g1625, g1627, g1630, g1632;
	reg g1634, g1636, g1645, g1646, g1650, g1653, g1657, g1660, g1663;
	reg g1667, g1678, g1681, g1683, g1685, g1689, g1691, g1693, g1696;
	reg g1706, g1709, g1712, g1715, g1718, g1721, g1724, g1729, g1739;
	reg g1742, g1744, g1746, g1749, g1751, g1753, g1756, g1765, g1768;
	reg g1769, g1771, g1774, g1776, g1778, g1781, g1791, g1794, g1797;
	reg g1799, g1802, g1804, g1806, g1809, g1818, g1821, g1823, g1825;
	reg g1826, g1828, g1830, g1832, g1842, g1843, g1844, g1846;

	always @ (posedge clk) begin done <= g134; end
	always @ (posedge clk) begin text_outx0x <= g149; end
	always @ (posedge clk) begin text_outx1x <= g156; end
	always @ (posedge clk) begin text_outx2x <= g163; end
	always @ (posedge clk) begin text_outx3x <= g170; end
	always @ (posedge clk) begin text_outx4x <= g177; end
	always @ (posedge clk) begin text_outx5x <= g184; end
	always @ (posedge clk) begin text_outx6x <= g191; end
	always @ (posedge clk) begin text_outx7x <= g198; end
	always @ (posedge clk) begin text_outx8x <= g213; end
	always @ (posedge clk) begin text_outx9x <= g220; end
	always @ (posedge clk) begin text_outx10x <= g227; end
	always @ (posedge clk) begin text_outx11x <= g234; end
	always @ (posedge clk) begin text_outx12x <= g241; end
	always @ (posedge clk) begin text_outx13x <= g248; end
	always @ (posedge clk) begin text_outx14x <= g255; end
	always @ (posedge clk) begin text_outx15x <= g262; end
	always @ (posedge clk) begin text_outx16x <= g277; end
	always @ (posedge clk) begin text_outx17x <= g284; end
	always @ (posedge clk) begin text_outx18x <= g291; end
	always @ (posedge clk) begin text_outx19x <= g298; end
	always @ (posedge clk) begin text_outx20x <= g305; end
	always @ (posedge clk) begin text_outx21x <= g312; end
	always @ (posedge clk) begin text_outx22x <= g319; end
	always @ (posedge clk) begin text_outx23x <= g326; end
	always @ (posedge clk) begin text_outx24x <= g341; end
	always @ (posedge clk) begin text_outx25x <= g348; end
	always @ (posedge clk) begin text_outx26x <= g355; end
	always @ (posedge clk) begin text_outx27x <= g362; end
	always @ (posedge clk) begin text_outx28x <= g369; end
	always @ (posedge clk) begin text_outx29x <= g376; end
	always @ (posedge clk) begin text_outx30x <= g383; end
	always @ (posedge clk) begin text_outx31x <= g390; end
	always @ (posedge clk) begin text_outx32x <= g405; end
	always @ (posedge clk) begin text_outx33x <= g412; end
	always @ (posedge clk) begin text_outx34x <= g419; end
	always @ (posedge clk) begin text_outx35x <= g426; end
	always @ (posedge clk) begin text_outx36x <= g433; end
	always @ (posedge clk) begin text_outx37x <= g440; end
	always @ (posedge clk) begin text_outx38x <= g447; end
	always @ (posedge clk) begin text_outx39x <= g454; end
	always @ (posedge clk) begin text_outx40x <= g469; end
	always @ (posedge clk) begin text_outx41x <= g476; end
	always @ (posedge clk) begin text_outx42x <= g483; end
	always @ (posedge clk) begin text_outx43x <= g490; end
	always @ (posedge clk) begin text_outx44x <= g497; end
	always @ (posedge clk) begin text_outx45x <= g504; end
	always @ (posedge clk) begin text_outx46x <= g511; end
	always @ (posedge clk) begin text_outx47x <= g518; end
	always @ (posedge clk) begin text_outx48x <= g533; end
	always @ (posedge clk) begin text_outx49x <= g540; end
	always @ (posedge clk) begin text_outx50x <= g547; end
	always @ (posedge clk) begin text_outx51x <= g554; end
	always @ (posedge clk) begin text_outx52x <= g561; end
	always @ (posedge clk) begin text_outx53x <= g568; end
	always @ (posedge clk) begin text_outx54x <= g575; end
	always @ (posedge clk) begin text_outx55x <= g582; end
	always @ (posedge clk) begin text_outx56x <= g597; end
	always @ (posedge clk) begin text_outx57x <= g604; end
	always @ (posedge clk) begin text_outx58x <= g611; end
	always @ (posedge clk) begin text_outx59x <= g618; end
	always @ (posedge clk) begin text_outx60x <= g625; end
	always @ (posedge clk) begin text_outx61x <= g632; end
	always @ (posedge clk) begin text_outx62x <= g639; end
	always @ (posedge clk) begin text_outx63x <= g646; end
	always @ (posedge clk) begin text_outx64x <= g661; end
	always @ (posedge clk) begin text_outx65x <= g668; end
	always @ (posedge clk) begin text_outx66x <= g675; end
	always @ (posedge clk) begin text_outx67x <= g682; end
	always @ (posedge clk) begin text_outx68x <= g689; end
	always @ (posedge clk) begin text_outx69x <= g696; end
	always @ (posedge clk) begin text_outx70x <= g703; end
	always @ (posedge clk) begin text_outx71x <= g710; end
	always @ (posedge clk) begin text_outx72x <= g725; end
	always @ (posedge clk) begin text_outx73x <= g732; end
	always @ (posedge clk) begin text_outx74x <= g739; end
	always @ (posedge clk) begin text_outx75x <= g746; end
	always @ (posedge clk) begin text_outx76x <= g753; end
	always @ (posedge clk) begin text_outx77x <= g760; end
	always @ (posedge clk) begin text_outx78x <= g767; end
	always @ (posedge clk) begin text_outx79x <= g774; end
	always @ (posedge clk) begin text_outx80x <= g789; end
	always @ (posedge clk) begin text_outx81x <= g796; end
	always @ (posedge clk) begin text_outx82x <= g803; end
	always @ (posedge clk) begin text_outx83x <= g810; end
	always @ (posedge clk) begin text_outx84x <= g817; end
	always @ (posedge clk) begin text_outx85x <= g824; end
	always @ (posedge clk) begin text_outx86x <= g831; end
	always @ (posedge clk) begin text_outx87x <= g838; end
	always @ (posedge clk) begin text_outx88x <= g853; end
	always @ (posedge clk) begin text_outx89x <= g860; end
	always @ (posedge clk) begin text_outx90x <= g867; end
	always @ (posedge clk) begin text_outx91x <= g874; end
	always @ (posedge clk) begin text_outx92x <= g881; end
	always @ (posedge clk) begin text_outx93x <= g888; end
	always @ (posedge clk) begin text_outx94x <= g895; end
	always @ (posedge clk) begin text_outx95x <= g902; end
	always @ (posedge clk) begin text_outx96x <= g917; end
	always @ (posedge clk) begin text_outx97x <= g924; end
	always @ (posedge clk) begin text_outx98x <= g931; end
	always @ (posedge clk) begin text_outx99x <= g938; end
	always @ (posedge clk) begin text_outx100x <= g945; end
	always @ (posedge clk) begin text_outx101x <= g952; end
	always @ (posedge clk) begin text_outx102x <= g959; end
	always @ (posedge clk) begin text_outx103x <= g966; end
	always @ (posedge clk) begin text_outx104x <= g981; end
	always @ (posedge clk) begin text_outx105x <= g988; end
	always @ (posedge clk) begin text_outx106x <= g995; end
	always @ (posedge clk) begin text_outx107x <= g1002; end
	always @ (posedge clk) begin text_outx108x <= g1009; end
	always @ (posedge clk) begin text_outx109x <= g1016; end
	always @ (posedge clk) begin text_outx110x <= g1023; end
	always @ (posedge clk) begin text_outx111x <= g1030; end
	always @ (posedge clk) begin text_outx112x <= g1045; end
	always @ (posedge clk) begin text_outx113x <= g1052; end
	always @ (posedge clk) begin text_outx114x <= g1059; end
	always @ (posedge clk) begin text_outx115x <= g1066; end
	always @ (posedge clk) begin text_outx116x <= g1073; end
	always @ (posedge clk) begin text_outx117x <= g1080; end
	always @ (posedge clk) begin text_outx118x <= g1087; end
	always @ (posedge clk) begin text_outx119x <= g1094; end
	always @ (posedge clk) begin text_outx120x <= g1109; end
	always @ (posedge clk) begin text_outx121x <= g1116; end
	always @ (posedge clk) begin text_outx122x <= g1123; end
	always @ (posedge clk) begin text_outx123x <= g1130; end
	always @ (posedge clk) begin text_outx124x <= g1137; end
	always @ (posedge clk) begin text_outx125x <= g1144; end
	always @ (posedge clk) begin text_outx126x <= g1151; end
	always @ (posedge clk) begin text_outx127x <= g1158; end
	always @ (posedge clk) begin g130 <= g1159; end
	always @ (posedge clk) begin g131 <= g1160; end
	always @ (posedge clk) begin g132 <= g1161; end
	always @ (posedge clk) begin g133 <= g1162; end
	always @ (posedge clk) begin g135 <= g1166; end
	always @ (posedge clk) begin g136 <= g1170; end
	always @ (posedge clk) begin g137 <= g1173; end
	always @ (posedge clk) begin g138 <= g2069; end
	always @ (posedge clk) begin g139 <= g1178; end
	always @ (posedge clk) begin g140 <= g1181; end
	always @ (posedge clk) begin g145 <= g1185; end
	always @ (posedge clk) begin g146 <= g1188; end
	always @ (posedge clk) begin g148 <= g1195; end
	always @ (posedge clk) begin g155 <= g1202; end
	always @ (posedge clk) begin g162 <= g1209; end
	always @ (posedge clk) begin g169 <= g1216; end
	always @ (posedge clk) begin g176 <= g1223; end
	always @ (posedge clk) begin g183 <= g1230; end
	always @ (posedge clk) begin g190 <= g1237; end
	always @ (posedge clk) begin g197 <= g1244; end
	always @ (posedge clk) begin g199 <= g1248; end
	always @ (posedge clk) begin g200 <= g1252; end
	always @ (posedge clk) begin g201 <= g1255; end
	always @ (posedge clk) begin g202 <= g1258; end
	always @ (posedge clk) begin g203 <= g1261; end
	always @ (posedge clk) begin g204 <= g1264; end
	always @ (posedge clk) begin g209 <= g1267; end
	always @ (posedge clk) begin g210 <= g1271; end
	always @ (posedge clk) begin g212 <= g1278; end
	always @ (posedge clk) begin g219 <= g1285; end
	always @ (posedge clk) begin g226 <= g1292; end
	always @ (posedge clk) begin g233 <= g1299; end
	always @ (posedge clk) begin g240 <= g1306; end
	always @ (posedge clk) begin g247 <= g1313; end
	always @ (posedge clk) begin g254 <= g1320; end
	always @ (posedge clk) begin g261 <= g1327; end
	always @ (posedge clk) begin g263 <= g1331; end
	always @ (posedge clk) begin g264 <= g1335; end
	always @ (posedge clk) begin g265 <= g1338; end
	always @ (posedge clk) begin g266 <= g2056; end
	always @ (posedge clk) begin g267 <= g1343; end
	always @ (posedge clk) begin g268 <= g1346; end
	always @ (posedge clk) begin g273 <= g1350; end
	always @ (posedge clk) begin g274 <= g1353; end
	always @ (posedge clk) begin g276 <= g1360; end
	always @ (posedge clk) begin g283 <= g1367; end
	always @ (posedge clk) begin g290 <= g1374; end
	always @ (posedge clk) begin g297 <= g1381; end
	always @ (posedge clk) begin g304 <= g1388; end
	always @ (posedge clk) begin g311 <= g1395; end
	always @ (posedge clk) begin g318 <= g1402; end
	always @ (posedge clk) begin g325 <= g1409; end
	always @ (posedge clk) begin g327 <= g1413; end
	always @ (posedge clk) begin g328 <= g2043; end
	always @ (posedge clk) begin g329 <= g1418; end
	always @ (posedge clk) begin g330 <= g1421; end
	always @ (posedge clk) begin g331 <= g1424; end
	always @ (posedge clk) begin g332 <= g1427; end
	always @ (posedge clk) begin g337 <= g2030; end
	always @ (posedge clk) begin g338 <= g1433; end
	always @ (posedge clk) begin g340 <= g1442; end
	always @ (posedge clk) begin g347 <= g1451; end
	always @ (posedge clk) begin g354 <= g1460; end
	always @ (posedge clk) begin g361 <= g1469; end
	always @ (posedge clk) begin g368 <= g1478; end
	always @ (posedge clk) begin g375 <= g1487; end
	always @ (posedge clk) begin g382 <= g1496; end
	always @ (posedge clk) begin g389 <= g1505; end
	always @ (posedge clk) begin g391 <= g1507; end
	always @ (posedge clk) begin g392 <= g1510; end
	always @ (posedge clk) begin g393 <= g1512; end
	always @ (posedge clk) begin g394 <= g2017; end
	always @ (posedge clk) begin g395 <= g1516; end
	always @ (posedge clk) begin g396 <= g1518; end
	always @ (posedge clk) begin g401 <= g1521; end
	always @ (posedge clk) begin g402 <= g1524; end
	always @ (posedge clk) begin g404 <= g1525; end
	always @ (posedge clk) begin g411 <= g1526; end
	always @ (posedge clk) begin g418 <= g1527; end
	always @ (posedge clk) begin g425 <= g1528; end
	always @ (posedge clk) begin g432 <= g1529; end
	always @ (posedge clk) begin g439 <= g1530; end
	always @ (posedge clk) begin g446 <= g1531; end
	always @ (posedge clk) begin g453 <= g1532; end
	always @ (posedge clk) begin g455 <= g1535; end
	always @ (posedge clk) begin g456 <= g1539; end
	always @ (posedge clk) begin g457 <= g1542; end
	always @ (posedge clk) begin g458 <= g1546; end
	always @ (posedge clk) begin g459 <= g1549; end
	always @ (posedge clk) begin g460 <= g1552; end
	always @ (posedge clk) begin g465 <= g1554; end
	always @ (posedge clk) begin g466 <= g1556; end
	always @ (posedge clk) begin g468 <= g1557; end
	always @ (posedge clk) begin g475 <= g1558; end
	always @ (posedge clk) begin g482 <= g1559; end
	always @ (posedge clk) begin g489 <= g1560; end
	always @ (posedge clk) begin g496 <= g1561; end
	always @ (posedge clk) begin g503 <= g1562; end
	always @ (posedge clk) begin g510 <= g1563; end
	always @ (posedge clk) begin g517 <= g1564; end
	always @ (posedge clk) begin g519 <= g1567; end
	always @ (posedge clk) begin g520 <= g2004; end
	always @ (posedge clk) begin g521 <= g1570; end
	always @ (posedge clk) begin g522 <= g1573; end
	always @ (posedge clk) begin g523 <= g1575; end
	always @ (posedge clk) begin g524 <= g1577; end
	always @ (posedge clk) begin g529 <= g1991; end
	always @ (posedge clk) begin g530 <= g1980; end
	always @ (posedge clk) begin g532 <= g1580; end
	always @ (posedge clk) begin g539 <= g1581; end
	always @ (posedge clk) begin g546 <= g1582; end
	always @ (posedge clk) begin g553 <= g1583; end
	always @ (posedge clk) begin g560 <= g1584; end
	always @ (posedge clk) begin g567 <= g1585; end
	always @ (posedge clk) begin g574 <= g1586; end
	always @ (posedge clk) begin g581 <= g1587; end
	always @ (posedge clk) begin g583 <= g1590; end
	always @ (posedge clk) begin g584 <= g1592; end
	always @ (posedge clk) begin g585 <= g1595; end
	always @ (posedge clk) begin g586 <= g1967; end
	always @ (posedge clk) begin g587 <= g1599; end
	always @ (posedge clk) begin g588 <= g1602; end
	always @ (posedge clk) begin g593 <= g1606; end
	always @ (posedge clk) begin g594 <= g1609; end
	always @ (posedge clk) begin g596 <= g1610; end
	always @ (posedge clk) begin g603 <= g1611; end
	always @ (posedge clk) begin g610 <= g1612; end
	always @ (posedge clk) begin g617 <= g1613; end
	always @ (posedge clk) begin g624 <= g1614; end
	always @ (posedge clk) begin g631 <= g1615; end
	always @ (posedge clk) begin g638 <= g1616; end
	always @ (posedge clk) begin g645 <= g1617; end
	always @ (posedge clk) begin g647 <= g1620; end
	always @ (posedge clk) begin g648 <= g1624; end
	always @ (posedge clk) begin g649 <= g1626; end
	always @ (posedge clk) begin g650 <= g1629; end
	always @ (posedge clk) begin g651 <= g1631; end
	always @ (posedge clk) begin g652 <= g1633; end
	always @ (posedge clk) begin g657 <= g1954; end
	always @ (posedge clk) begin g658 <= g1943; end
	always @ (posedge clk) begin g660 <= g1637; end
	always @ (posedge clk) begin g667 <= g1638; end
	always @ (posedge clk) begin g674 <= g1639; end
	always @ (posedge clk) begin g681 <= g1640; end
	always @ (posedge clk) begin g688 <= g1641; end
	always @ (posedge clk) begin g695 <= g1642; end
	always @ (posedge clk) begin g702 <= g1643; end
	always @ (posedge clk) begin g709 <= g1644; end
	always @ (posedge clk) begin g711 <= g1932; end
	always @ (posedge clk) begin g712 <= g1649; end
	always @ (posedge clk) begin g713 <= g1652; end
	always @ (posedge clk) begin g714 <= g1656; end
	always @ (posedge clk) begin g715 <= g1659; end
	always @ (posedge clk) begin g716 <= g1662; end
	always @ (posedge clk) begin g721 <= g1666; end
	always @ (posedge clk) begin g722 <= g1669; end
	always @ (posedge clk) begin g724 <= g1670; end
	always @ (posedge clk) begin g731 <= g1671; end
	always @ (posedge clk) begin g738 <= g1672; end
	always @ (posedge clk) begin g745 <= g1673; end
	always @ (posedge clk) begin g752 <= g1674; end
	always @ (posedge clk) begin g759 <= g1675; end
	always @ (posedge clk) begin g766 <= g1676; end
	always @ (posedge clk) begin g773 <= g1677; end
	always @ (posedge clk) begin g775 <= g1680; end
	always @ (posedge clk) begin g776 <= g1919; end
	always @ (posedge clk) begin g777 <= g1684; end
	always @ (posedge clk) begin g778 <= g1688; end
	always @ (posedge clk) begin g779 <= g1690; end
	always @ (posedge clk) begin g780 <= g1692; end
	always @ (posedge clk) begin g785 <= g1695; end
	always @ (posedge clk) begin g786 <= g1697; end
	always @ (posedge clk) begin g788 <= g1698; end
	always @ (posedge clk) begin g795 <= g1699; end
	always @ (posedge clk) begin g802 <= g1700; end
	always @ (posedge clk) begin g809 <= g1701; end
	always @ (posedge clk) begin g816 <= g1702; end
	always @ (posedge clk) begin g823 <= g1703; end
	always @ (posedge clk) begin g830 <= g1704; end
	always @ (posedge clk) begin g837 <= g1705; end
	always @ (posedge clk) begin g839 <= g1708; end
	always @ (posedge clk) begin g840 <= g1711; end
	always @ (posedge clk) begin g841 <= g1714; end
	always @ (posedge clk) begin g842 <= g1717; end
	always @ (posedge clk) begin g843 <= g1720; end
	always @ (posedge clk) begin g844 <= g1723; end
	always @ (posedge clk) begin g849 <= g1727; end
	always @ (posedge clk) begin g850 <= g1730; end
	always @ (posedge clk) begin g852 <= g1731; end
	always @ (posedge clk) begin g859 <= g1732; end
	always @ (posedge clk) begin g866 <= g1733; end
	always @ (posedge clk) begin g873 <= g1734; end
	always @ (posedge clk) begin g880 <= g1735; end
	always @ (posedge clk) begin g887 <= g1736; end
	always @ (posedge clk) begin g894 <= g1737; end
	always @ (posedge clk) begin g901 <= g1738; end
	always @ (posedge clk) begin g903 <= g1741; end
	always @ (posedge clk) begin g904 <= g1743; end
	always @ (posedge clk) begin g905 <= g1745; end
	always @ (posedge clk) begin g906 <= g1748; end
	always @ (posedge clk) begin g907 <= g1750; end
	always @ (posedge clk) begin g908 <= g1752; end
	always @ (posedge clk) begin g913 <= g1755; end
	always @ (posedge clk) begin g914 <= g1908; end
	always @ (posedge clk) begin g916 <= g1757; end
	always @ (posedge clk) begin g923 <= g1758; end
	always @ (posedge clk) begin g930 <= g1759; end
	always @ (posedge clk) begin g937 <= g1760; end
	always @ (posedge clk) begin g944 <= g1761; end
	always @ (posedge clk) begin g951 <= g1762; end
	always @ (posedge clk) begin g958 <= g1763; end
	always @ (posedge clk) begin g965 <= g1764; end
	always @ (posedge clk) begin g967 <= g1767; end
	always @ (posedge clk) begin g968 <= g1895; end
	always @ (posedge clk) begin g969 <= g1770; end
	always @ (posedge clk) begin g970 <= g1773; end
	always @ (posedge clk) begin g971 <= g1775; end
	always @ (posedge clk) begin g972 <= g1777; end
	always @ (posedge clk) begin g977 <= g1780; end
	always @ (posedge clk) begin g978 <= g1782; end
	always @ (posedge clk) begin g980 <= g1783; end
	always @ (posedge clk) begin g987 <= g1784; end
	always @ (posedge clk) begin g994 <= g1785; end
	always @ (posedge clk) begin g1001 <= g1786; end
	always @ (posedge clk) begin g1008 <= g1787; end
	always @ (posedge clk) begin g1015 <= g1788; end
	always @ (posedge clk) begin g1022 <= g1789; end
	always @ (posedge clk) begin g1029 <= g1790; end
	always @ (posedge clk) begin g1031 <= g1793; end
	always @ (posedge clk) begin g1032 <= g1796; end
	always @ (posedge clk) begin g1033 <= g1798; end
	always @ (posedge clk) begin g1034 <= g1801; end
	always @ (posedge clk) begin g1035 <= g1803; end
	always @ (posedge clk) begin g1036 <= g1805; end
	always @ (posedge clk) begin g1041 <= g1808; end
	always @ (posedge clk) begin g1042 <= g1884; end
	always @ (posedge clk) begin g1044 <= g1810; end
	always @ (posedge clk) begin g1051 <= g1811; end
	always @ (posedge clk) begin g1058 <= g1812; end
	always @ (posedge clk) begin g1065 <= g1813; end
	always @ (posedge clk) begin g1072 <= g1814; end
	always @ (posedge clk) begin g1079 <= g1815; end
	always @ (posedge clk) begin g1086 <= g1816; end
	always @ (posedge clk) begin g1093 <= g1817; end
	always @ (posedge clk) begin g1095 <= g1820; end
	always @ (posedge clk) begin g1096 <= g1822; end
	always @ (posedge clk) begin g1097 <= g1824; end
	always @ (posedge clk) begin g1098 <= g1871; end
	always @ (posedge clk) begin g1099 <= g1827; end
	always @ (posedge clk) begin g1100 <= g1829; end
	always @ (posedge clk) begin g1105 <= g1858; end
	always @ (posedge clk) begin g1106 <= g1833; end
	always @ (posedge clk) begin g1108 <= g1834; end
	always @ (posedge clk) begin g1115 <= g1835; end
	always @ (posedge clk) begin g1122 <= g1836; end
	always @ (posedge clk) begin g1129 <= g1837; end
	always @ (posedge clk) begin g1136 <= g1838; end
	always @ (posedge clk) begin g1143 <= g1839; end
	always @ (posedge clk) begin g1150 <= g1840; end
	always @ (posedge clk) begin g1157 <= g1841; end
	always @ (posedge clk) begin g1163 <= ld; end
	always @ (posedge clk) begin g1164 <= g2082; end
	always @ (posedge clk) begin g1167 <= g2083; end
	always @ (posedge clk) begin g1171 <= g2084; end
	always @ (posedge clk) begin g1174 <= g2085; end
	always @ (posedge clk) begin g1176 <= g2086; end
	always @ (posedge clk) begin g1179 <= g2087; end
	always @ (posedge clk) begin g1182 <= g2088; end
	always @ (posedge clk) begin g1186 <= g2089; end
	always @ (posedge clk) begin g1245 <= g2090; end
	always @ (posedge clk) begin g1249 <= g2091; end
	always @ (posedge clk) begin g1253 <= g2092; end
	always @ (posedge clk) begin g1256 <= g2093; end
	always @ (posedge clk) begin g1259 <= g2094; end
	always @ (posedge clk) begin g1262 <= g2095; end
	always @ (posedge clk) begin g1265 <= g2096; end
	always @ (posedge clk) begin g1268 <= g2097; end
	always @ (posedge clk) begin g1328 <= g2098; end
	always @ (posedge clk) begin g1332 <= g2099; end
	always @ (posedge clk) begin g1336 <= g2100; end
	always @ (posedge clk) begin g1339 <= g2101; end
	always @ (posedge clk) begin g1341 <= g2102; end
	always @ (posedge clk) begin g1344 <= g2103; end
	always @ (posedge clk) begin g1347 <= g2104; end
	always @ (posedge clk) begin g1351 <= g2105; end
	always @ (posedge clk) begin g1410 <= g2106; end
	always @ (posedge clk) begin g1414 <= g2107; end
	always @ (posedge clk) begin g1416 <= g2108; end
	always @ (posedge clk) begin g1419 <= g2109; end
	always @ (posedge clk) begin g1422 <= g2110; end
	always @ (posedge clk) begin g1425 <= g2111; end
	always @ (posedge clk) begin g1428 <= g2112; end
	always @ (posedge clk) begin g1430 <= g2113; end
	always @ (posedge clk) begin g1439 <= g1845; end
	always @ (posedge clk) begin g1448 <= g1857; end
	always @ (posedge clk) begin g1457 <= g1856; end
	always @ (posedge clk) begin g1466 <= g1855; end
	always @ (posedge clk) begin g1475 <= g1854; end
	always @ (posedge clk) begin g1484 <= g1853; end
	always @ (posedge clk) begin g1493 <= g1847; end
	always @ (posedge clk) begin g1502 <= g1848; end
	always @ (posedge clk) begin g1506 <= g2114; end
	always @ (posedge clk) begin g1508 <= g2115; end
	always @ (posedge clk) begin g1511 <= g2116; end
	always @ (posedge clk) begin g1513 <= g2117; end
	always @ (posedge clk) begin g1515 <= g2118; end
	always @ (posedge clk) begin g1517 <= g2119; end
	always @ (posedge clk) begin g1519 <= g2120; end
	always @ (posedge clk) begin g1522 <= g2121; end
	always @ (posedge clk) begin g1533 <= g2122; end
	always @ (posedge clk) begin g1536 <= g2123; end
	always @ (posedge clk) begin g1540 <= g2124; end
	always @ (posedge clk) begin g1543 <= g2125; end
	always @ (posedge clk) begin g1547 <= g2126; end
	always @ (posedge clk) begin g1550 <= g2127; end
	always @ (posedge clk) begin g1553 <= g2128; end
	always @ (posedge clk) begin g1555 <= g2129; end
	always @ (posedge clk) begin g1565 <= g2130; end
	always @ (posedge clk) begin g1568 <= g2131; end
	always @ (posedge clk) begin g1569 <= g2132; end
	always @ (posedge clk) begin g1571 <= g2133; end
	always @ (posedge clk) begin g1574 <= g2134; end
	always @ (posedge clk) begin g1576 <= g2135; end
	always @ (posedge clk) begin g1578 <= g2136; end
	always @ (posedge clk) begin g1579 <= g2137; end
	always @ (posedge clk) begin g1588 <= g2138; end
	always @ (posedge clk) begin g1591 <= g2139; end
	always @ (posedge clk) begin g1593 <= g2140; end
	always @ (posedge clk) begin g1596 <= g2141; end
	always @ (posedge clk) begin g1597 <= g2142; end
	always @ (posedge clk) begin g1600 <= g2143; end
	always @ (posedge clk) begin g1603 <= g2144; end
	always @ (posedge clk) begin g1607 <= g2145; end
	always @ (posedge clk) begin g1619 <= g2146; end
	always @ (posedge clk) begin g1621 <= g2147; end
	always @ (posedge clk) begin g1625 <= g2148; end
	always @ (posedge clk) begin g1627 <= g2149; end
	always @ (posedge clk) begin g1630 <= g2150; end
	always @ (posedge clk) begin g1632 <= g2151; end
	always @ (posedge clk) begin g1634 <= g2152; end
	always @ (posedge clk) begin g1636 <= g2153; end
	always @ (posedge clk) begin g1645 <= g2154; end
	always @ (posedge clk) begin g1646 <= g2155; end
	always @ (posedge clk) begin g1650 <= g2156; end
	always @ (posedge clk) begin g1653 <= g2157; end
	always @ (posedge clk) begin g1657 <= g2158; end
	always @ (posedge clk) begin g1660 <= g2159; end
	always @ (posedge clk) begin g1663 <= g2160; end
	always @ (posedge clk) begin g1667 <= g2161; end
	always @ (posedge clk) begin g1678 <= g2162; end
	always @ (posedge clk) begin g1681 <= g2163; end
	always @ (posedge clk) begin g1683 <= g2164; end
	always @ (posedge clk) begin g1685 <= g2165; end
	always @ (posedge clk) begin g1689 <= g2166; end
	always @ (posedge clk) begin g1691 <= g2167; end
	always @ (posedge clk) begin g1693 <= g2168; end
	always @ (posedge clk) begin g1696 <= g2169; end
	always @ (posedge clk) begin g1706 <= g2170; end
	always @ (posedge clk) begin g1709 <= g2171; end
	always @ (posedge clk) begin g1712 <= g2172; end
	always @ (posedge clk) begin g1715 <= g2173; end
	always @ (posedge clk) begin g1718 <= g2174; end
	always @ (posedge clk) begin g1721 <= g2175; end
	always @ (posedge clk) begin g1724 <= g2176; end
	always @ (posedge clk) begin g1729 <= g2177; end
	always @ (posedge clk) begin g1739 <= g2178; end
	always @ (posedge clk) begin g1742 <= g2179; end
	always @ (posedge clk) begin g1744 <= g2180; end
	always @ (posedge clk) begin g1746 <= g2181; end
	always @ (posedge clk) begin g1749 <= g2182; end
	always @ (posedge clk) begin g1751 <= g2183; end
	always @ (posedge clk) begin g1753 <= g2184; end
	always @ (posedge clk) begin g1756 <= g2185; end
	always @ (posedge clk) begin g1765 <= g2186; end
	always @ (posedge clk) begin g1768 <= g2187; end
	always @ (posedge clk) begin g1769 <= g2188; end
	always @ (posedge clk) begin g1771 <= g2189; end
	always @ (posedge clk) begin g1774 <= g2190; end
	always @ (posedge clk) begin g1776 <= g2191; end
	always @ (posedge clk) begin g1778 <= g2192; end
	always @ (posedge clk) begin g1781 <= g2193; end
	always @ (posedge clk) begin g1791 <= g2194; end
	always @ (posedge clk) begin g1794 <= g2195; end
	always @ (posedge clk) begin g1797 <= g2196; end
	always @ (posedge clk) begin g1799 <= g2197; end
	always @ (posedge clk) begin g1802 <= g2198; end
	always @ (posedge clk) begin g1804 <= g2199; end
	always @ (posedge clk) begin g1806 <= g2200; end
	always @ (posedge clk) begin g1809 <= g2201; end
	always @ (posedge clk) begin g1818 <= g2202; end
	always @ (posedge clk) begin g1821 <= g2203; end
	always @ (posedge clk) begin g1823 <= g2204; end
	always @ (posedge clk) begin g1825 <= g2205; end
	always @ (posedge clk) begin g1826 <= g2206; end
	always @ (posedge clk) begin g1828 <= g2207; end
	always @ (posedge clk) begin g1830 <= g2208; end
	always @ (posedge clk) begin g1832 <= g2209; end
	always @ (posedge clk) begin g1842 <= g1849; end
	always @ (posedge clk) begin g1843 <= g1850; end
	always @ (posedge clk) begin g1844 <= g1851; end
	always @ (posedge clk) begin g1846 <= g1852; end

	assign g134 = (((!g130) & (!g131) & (!sk[0]) & (!g132) & (!g133) & (ld)) + ((!g130) & (!g131) & (!sk[0]) & (!g132) & (g133) & (ld)) + ((!g130) & (!g131) & (!sk[0]) & (g132) & (!g133) & (ld)) + ((!g130) & (!g131) & (!sk[0]) & (g132) & (g133) & (ld)) + ((!g130) & (g131) & (!sk[0]) & (!g132) & (!g133) & (!ld)) + ((!g130) & (g131) & (!sk[0]) & (!g132) & (!g133) & (ld)) + ((!g130) & (g131) & (!sk[0]) & (!g132) & (g133) & (!ld)) + ((!g130) & (g131) & (!sk[0]) & (!g132) & (g133) & (ld)) + ((!g130) & (g131) & (!sk[0]) & (g132) & (!g133) & (!ld)) + ((!g130) & (g131) & (!sk[0]) & (g132) & (!g133) & (ld)) + ((!g130) & (g131) & (!sk[0]) & (g132) & (g133) & (!ld)) + ((!g130) & (g131) & (!sk[0]) & (g132) & (g133) & (ld)) + ((g130) & (!g131) & (!sk[0]) & (!g132) & (!g133) & (ld)) + ((g130) & (!g131) & (!sk[0]) & (!g132) & (g133) & (!ld)) + ((g130) & (!g131) & (!sk[0]) & (!g132) & (g133) & (ld)) + ((g130) & (!g131) & (!sk[0]) & (g132) & (!g133) & (ld)) + ((g130) & (!g131) & (!sk[0]) & (g132) & (g133) & (!ld)) + ((g130) & (!g131) & (!sk[0]) & (g132) & (g133) & (ld)) + ((g130) & (!g131) & (sk[0]) & (!g132) & (!g133) & (!ld)) + ((g130) & (g131) & (!sk[0]) & (!g132) & (!g133) & (!ld)) + ((g130) & (g131) & (!sk[0]) & (!g132) & (!g133) & (ld)) + ((g130) & (g131) & (!sk[0]) & (!g132) & (g133) & (!ld)) + ((g130) & (g131) & (!sk[0]) & (!g132) & (g133) & (ld)) + ((g130) & (g131) & (!sk[0]) & (g132) & (!g133) & (!ld)) + ((g130) & (g131) & (!sk[0]) & (g132) & (!g133) & (ld)) + ((g130) & (g131) & (!sk[0]) & (g132) & (g133) & (!ld)) + ((g130) & (g131) & (!sk[0]) & (g132) & (g133) & (ld)));
	assign g141 = (((!g135) & (!g136) & (!g137) & (!g138) & (g139) & (g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g139) & (!g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g139) & (g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (g139) & (!g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (!g139) & (!g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (!g139) & (g140)) + ((!g135) & (!g136) & (g137) & (g138) & (!g139) & (!g140)) + ((!g135) & (!g136) & (g137) & (g138) & (g139) & (g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (g139) & (!g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (g139) & (g140)) + ((!g135) & (g136) & (!g137) & (g138) & (g139) & (!g140)) + ((!g135) & (g136) & (!g137) & (g138) & (g139) & (g140)) + ((!g135) & (g136) & (g137) & (!g138) & (g139) & (!g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (!g139) & (!g140)) + ((g135) & (!g136) & (g137) & (!g138) & (g139) & (!g140)) + ((g135) & (!g136) & (g137) & (g138) & (!g139) & (g140)) + ((g135) & (!g136) & (g137) & (g138) & (g139) & (g140)) + ((g135) & (g136) & (!g137) & (!g138) & (!g139) & (g140)) + ((g135) & (g136) & (!g137) & (!g138) & (g139) & (!g140)) + ((g135) & (g136) & (g137) & (!g138) & (!g139) & (g140)) + ((g135) & (g136) & (g137) & (!g138) & (g139) & (!g140)) + ((g135) & (g136) & (g137) & (g138) & (!g139) & (!g140)) + ((g135) & (g136) & (g137) & (g138) & (g139) & (!g140)) + ((g135) & (g136) & (g137) & (g138) & (g139) & (g140)));
	assign g142 = (((!g135) & (!g136) & (!g137) & (!g138) & (g139) & (!g140)) + ((!g135) & (!g136) & (!g137) & (!g138) & (g139) & (g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g139) & (!g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g139) & (g140)) + ((!g135) & (!g136) & (g137) & (g138) & (!g139) & (g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (!g139) & (!g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (!g139) & (g140)) + ((!g135) & (g136) & (g137) & (!g138) & (!g139) & (!g140)) + ((!g135) & (g136) & (g137) & (!g138) & (!g139) & (g140)) + ((!g135) & (g136) & (g137) & (!g138) & (g139) & (!g140)) + ((!g135) & (g136) & (g137) & (g138) & (g139) & (g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (!g139) & (g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (g139) & (!g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (g139) & (g140)) + ((g135) & (!g136) & (!g137) & (g138) & (g139) & (!g140)) + ((g135) & (!g136) & (g137) & (!g138) & (!g139) & (!g140)) + ((g135) & (!g136) & (g137) & (!g138) & (g139) & (g140)) + ((g135) & (!g136) & (g137) & (g138) & (!g139) & (g140)) + ((g135) & (!g136) & (g137) & (g138) & (g139) & (g140)) + ((g135) & (g136) & (!g137) & (!g138) & (!g139) & (!g140)) + ((g135) & (g136) & (!g137) & (!g138) & (!g139) & (g140)) + ((g135) & (g136) & (!g137) & (!g138) & (g139) & (!g140)) + ((g135) & (g136) & (!g137) & (!g138) & (g139) & (g140)) + ((g135) & (g136) & (!g137) & (g138) & (!g139) & (!g140)) + ((g135) & (g136) & (!g137) & (g138) & (g139) & (!g140)) + ((g135) & (g136) & (!g137) & (g138) & (g139) & (g140)) + ((g135) & (g136) & (g137) & (!g138) & (g139) & (!g140)) + ((g135) & (g136) & (g137) & (!g138) & (g139) & (g140)) + ((g135) & (g136) & (g137) & (g138) & (!g139) & (g140)) + ((g135) & (g136) & (g137) & (g138) & (g139) & (!g140)));
	assign g143 = (((!g135) & (!g136) & (!g137) & (!g138) & (!g139) & (!g140)) + ((!g135) & (!g136) & (!g137) & (!g138) & (g139) & (g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (g139) & (g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (!g139) & (!g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (!g139) & (g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (g139) & (g140)) + ((!g135) & (!g136) & (g137) & (g138) & (!g139) & (g140)) + ((!g135) & (!g136) & (g137) & (g138) & (g139) & (!g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (!g139) & (!g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (g139) & (!g140)) + ((!g135) & (g136) & (!g137) & (g138) & (g139) & (g140)) + ((!g135) & (g136) & (g137) & (g138) & (!g139) & (!g140)) + ((!g135) & (g136) & (g137) & (g138) & (g139) & (!g140)) + ((g135) & (!g136) & (!g137) & (g138) & (!g139) & (!g140)) + ((g135) & (!g136) & (!g137) & (g138) & (!g139) & (g140)) + ((g135) & (!g136) & (!g137) & (g138) & (g139) & (!g140)) + ((g135) & (!g136) & (g137) & (!g138) & (!g139) & (!g140)) + ((g135) & (!g136) & (g137) & (!g138) & (g139) & (g140)) + ((g135) & (!g136) & (g137) & (g138) & (!g139) & (!g140)) + ((g135) & (!g136) & (g137) & (g138) & (!g139) & (g140)) + ((g135) & (!g136) & (g137) & (g138) & (g139) & (!g140)) + ((g135) & (!g136) & (g137) & (g138) & (g139) & (g140)) + ((g135) & (g136) & (!g137) & (!g138) & (g139) & (g140)) + ((g135) & (g136) & (!g137) & (g138) & (!g139) & (!g140)) + ((g135) & (g136) & (!g137) & (g138) & (g139) & (!g140)) + ((g135) & (g136) & (!g137) & (g138) & (g139) & (g140)) + ((g135) & (g136) & (g137) & (!g138) & (!g139) & (!g140)) + ((g135) & (g136) & (g137) & (g138) & (!g139) & (!g140)) + ((g135) & (g136) & (g137) & (g138) & (!g139) & (g140)) + ((g135) & (g136) & (g137) & (g138) & (g139) & (g140)));
	assign g144 = (((!g135) & (!g136) & (!g137) & (!g138) & (!g139) & (g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (g139) & (!g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (g139) & (g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (!g139) & (g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (g139) & (g140)) + ((!g135) & (!g136) & (g137) & (g138) & (!g139) & (g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (!g139) & (!g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (!g139) & (g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (g139) & (!g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (g139) & (g140)) + ((!g135) & (g136) & (!g137) & (g138) & (g139) & (!g140)) + ((!g135) & (g136) & (!g137) & (g138) & (g139) & (g140)) + ((!g135) & (g136) & (g137) & (g138) & (!g139) & (!g140)) + ((!g135) & (g136) & (g137) & (g138) & (g139) & (!g140)) + ((!g135) & (g136) & (g137) & (g138) & (g139) & (g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (!g139) & (!g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (g139) & (g140)) + ((g135) & (!g136) & (!g137) & (g138) & (g139) & (!g140)) + ((g135) & (!g136) & (!g137) & (g138) & (g139) & (g140)) + ((g135) & (!g136) & (g137) & (!g138) & (!g139) & (g140)) + ((g135) & (!g136) & (g137) & (!g138) & (g139) & (!g140)) + ((g135) & (!g136) & (g137) & (g138) & (g139) & (!g140)) + ((g135) & (g136) & (!g137) & (!g138) & (!g139) & (g140)) + ((g135) & (g136) & (!g137) & (!g138) & (g139) & (g140)) + ((g135) & (g136) & (!g137) & (g138) & (g139) & (!g140)) + ((g135) & (g136) & (!g137) & (g138) & (g139) & (g140)) + ((g135) & (g136) & (g137) & (!g138) & (!g139) & (g140)) + ((g135) & (g136) & (g137) & (g138) & (!g139) & (!g140)));
	assign g147 = (((!g141) & (!g142) & (!g143) & (!g144) & (!g145) & (!g146)) + ((!g141) & (!g142) & (!g143) & (g144) & (!g145) & (!g146)) + ((!g141) & (!g142) & (!g143) & (g144) & (g145) & (g146)) + ((!g141) & (!g142) & (g143) & (!g144) & (!g145) & (!g146)) + ((!g141) & (!g142) & (g143) & (!g144) & (!g145) & (g146)) + ((!g141) & (!g142) & (g143) & (g144) & (!g145) & (!g146)) + ((!g141) & (!g142) & (g143) & (g144) & (!g145) & (g146)) + ((!g141) & (!g142) & (g143) & (g144) & (g145) & (g146)) + ((!g141) & (g142) & (!g143) & (!g144) & (!g145) & (!g146)) + ((!g141) & (g142) & (!g143) & (!g144) & (g145) & (!g146)) + ((!g141) & (g142) & (!g143) & (g144) & (!g145) & (!g146)) + ((!g141) & (g142) & (!g143) & (g144) & (g145) & (!g146)) + ((!g141) & (g142) & (!g143) & (g144) & (g145) & (g146)) + ((!g141) & (g142) & (g143) & (!g144) & (!g145) & (!g146)) + ((!g141) & (g142) & (g143) & (!g144) & (!g145) & (g146)) + ((!g141) & (g142) & (g143) & (!g144) & (g145) & (!g146)) + ((!g141) & (g142) & (g143) & (g144) & (!g145) & (!g146)) + ((!g141) & (g142) & (g143) & (g144) & (!g145) & (g146)) + ((!g141) & (g142) & (g143) & (g144) & (g145) & (!g146)) + ((!g141) & (g142) & (g143) & (g144) & (g145) & (g146)) + ((g141) & (!g142) & (!g143) & (g144) & (g145) & (g146)) + ((g141) & (!g142) & (g143) & (!g144) & (!g145) & (g146)) + ((g141) & (!g142) & (g143) & (g144) & (!g145) & (g146)) + ((g141) & (!g142) & (g143) & (g144) & (g145) & (g146)) + ((g141) & (g142) & (!g143) & (!g144) & (g145) & (!g146)) + ((g141) & (g142) & (!g143) & (g144) & (g145) & (!g146)) + ((g141) & (g142) & (!g143) & (g144) & (g145) & (g146)) + ((g141) & (g142) & (g143) & (!g144) & (!g145) & (g146)) + ((g141) & (g142) & (g143) & (!g144) & (g145) & (!g146)) + ((g141) & (g142) & (g143) & (g144) & (!g145) & (g146)) + ((g141) & (g142) & (g143) & (g144) & (g145) & (!g146)) + ((g141) & (g142) & (g143) & (g144) & (g145) & (g146)));
	assign g149 = (((!g147) & (sk[6]) & (g148)) + ((g147) & (!sk[6]) & (!g148)) + ((g147) & (!sk[6]) & (g148)) + ((g147) & (sk[6]) & (!g148)));
	assign g150 = (((!g135) & (!g136) & (!g137) & (!g138) & (!g145) & (g139)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g145) & (!g139)) + ((!g135) & (!g136) & (!g137) & (g138) & (g145) & (!g139)) + ((!g135) & (!g136) & (g137) & (!g138) & (g145) & (g139)) + ((!g135) & (!g136) & (g137) & (g138) & (!g145) & (g139)) + ((!g135) & (!g136) & (g137) & (g138) & (g145) & (!g139)) + ((!g135) & (g136) & (!g137) & (!g138) & (!g145) & (g139)) + ((!g135) & (g136) & (!g137) & (!g138) & (g145) & (!g139)) + ((!g135) & (g136) & (!g137) & (!g138) & (g145) & (g139)) + ((!g135) & (g136) & (g137) & (!g138) & (g145) & (g139)) + ((!g135) & (g136) & (g137) & (g138) & (g145) & (g139)) + ((g135) & (!g136) & (!g137) & (!g138) & (!g145) & (!g139)) + ((g135) & (!g136) & (!g137) & (!g138) & (g145) & (g139)) + ((g135) & (!g136) & (!g137) & (g138) & (!g145) & (!g139)) + ((g135) & (!g136) & (!g137) & (g138) & (g145) & (!g139)) + ((g135) & (!g136) & (g137) & (!g138) & (g145) & (!g139)) + ((g135) & (!g136) & (g137) & (!g138) & (g145) & (g139)) + ((g135) & (!g136) & (g137) & (g138) & (g145) & (!g139)) + ((g135) & (!g136) & (g137) & (g138) & (g145) & (g139)) + ((g135) & (g136) & (!g137) & (!g138) & (g145) & (!g139)) + ((g135) & (g136) & (!g137) & (!g138) & (g145) & (g139)) + ((g135) & (g136) & (!g137) & (g138) & (g145) & (g139)) + ((g135) & (g136) & (g137) & (!g138) & (!g145) & (!g139)) + ((g135) & (g136) & (g137) & (!g138) & (!g145) & (g139)) + ((g135) & (g136) & (g137) & (!g138) & (g145) & (!g139)) + ((g135) & (g136) & (g137) & (g138) & (!g145) & (g139)) + ((g135) & (g136) & (g137) & (g138) & (g145) & (!g139)));
	assign g151 = (((!g135) & (!g136) & (!g137) & (!g138) & (!g145) & (g139)) + ((!g135) & (!g136) & (!g137) & (!g138) & (g145) & (!g139)) + ((!g135) & (!g136) & (!g137) & (!g138) & (g145) & (g139)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g145) & (!g139)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g145) & (g139)) + ((!g135) & (!g136) & (!g137) & (g138) & (g145) & (g139)) + ((!g135) & (!g136) & (g137) & (!g138) & (g145) & (!g139)) + ((!g135) & (!g136) & (g137) & (g138) & (!g145) & (!g139)) + ((!g135) & (!g136) & (g137) & (g138) & (!g145) & (g139)) + ((!g135) & (!g136) & (g137) & (g138) & (g145) & (g139)) + ((!g135) & (g136) & (!g137) & (!g138) & (g145) & (g139)) + ((!g135) & (g136) & (!g137) & (g138) & (!g145) & (!g139)) + ((!g135) & (g136) & (!g137) & (g138) & (g145) & (!g139)) + ((!g135) & (g136) & (g137) & (!g138) & (g145) & (!g139)) + ((!g135) & (g136) & (g137) & (!g138) & (g145) & (g139)) + ((!g135) & (g136) & (g137) & (g138) & (!g145) & (!g139)) + ((g135) & (!g136) & (!g137) & (!g138) & (!g145) & (!g139)) + ((g135) & (!g136) & (!g137) & (g138) & (!g145) & (!g139)) + ((g135) & (!g136) & (!g137) & (g138) & (!g145) & (g139)) + ((g135) & (!g136) & (g137) & (!g138) & (!g145) & (g139)) + ((g135) & (!g136) & (g137) & (!g138) & (g145) & (g139)) + ((g135) & (!g136) & (g137) & (g138) & (!g145) & (!g139)) + ((g135) & (!g136) & (g137) & (g138) & (!g145) & (g139)) + ((g135) & (g136) & (!g137) & (g138) & (!g145) & (!g139)) + ((g135) & (g136) & (!g137) & (g138) & (g145) & (g139)) + ((g135) & (g136) & (g137) & (!g138) & (!g145) & (!g139)) + ((g135) & (g136) & (g137) & (!g138) & (!g145) & (g139)) + ((g135) & (g136) & (g137) & (!g138) & (g145) & (g139)) + ((g135) & (g136) & (g137) & (g138) & (!g145) & (!g139)) + ((g135) & (g136) & (g137) & (g138) & (!g145) & (g139)) + ((g135) & (g136) & (g137) & (g138) & (g145) & (!g139)));
	assign g152 = (((!g135) & (!g136) & (!g137) & (!g138) & (!g145) & (g139)) + ((!g135) & (!g136) & (!g137) & (g138) & (g145) & (!g139)) + ((!g135) & (!g136) & (g137) & (!g138) & (!g145) & (!g139)) + ((!g135) & (!g136) & (g137) & (!g138) & (g145) & (!g139)) + ((!g135) & (!g136) & (g137) & (g138) & (!g145) & (g139)) + ((!g135) & (!g136) & (g137) & (g138) & (g145) & (!g139)) + ((!g135) & (!g136) & (g137) & (g138) & (g145) & (g139)) + ((!g135) & (g136) & (!g137) & (!g138) & (!g145) & (!g139)) + ((!g135) & (g136) & (!g137) & (!g138) & (g145) & (!g139)) + ((!g135) & (g136) & (!g137) & (g138) & (!g145) & (!g139)) + ((!g135) & (g136) & (!g137) & (g138) & (g145) & (g139)) + ((!g135) & (g136) & (g137) & (!g138) & (g145) & (g139)) + ((!g135) & (g136) & (g137) & (g138) & (!g145) & (g139)) + ((!g135) & (g136) & (g137) & (g138) & (g145) & (!g139)) + ((g135) & (!g136) & (!g137) & (!g138) & (g145) & (g139)) + ((g135) & (!g136) & (!g137) & (g138) & (!g145) & (!g139)) + ((g135) & (!g136) & (!g137) & (g138) & (g145) & (!g139)) + ((g135) & (!g136) & (g137) & (!g138) & (!g145) & (!g139)) + ((g135) & (!g136) & (g137) & (!g138) & (!g145) & (g139)) + ((g135) & (!g136) & (g137) & (!g138) & (g145) & (!g139)) + ((g135) & (!g136) & (g137) & (!g138) & (g145) & (g139)) + ((g135) & (!g136) & (g137) & (g138) & (g145) & (!g139)) + ((g135) & (g136) & (!g137) & (!g138) & (!g145) & (g139)) + ((g135) & (g136) & (!g137) & (!g138) & (g145) & (g139)) + ((g135) & (g136) & (!g137) & (g138) & (!g145) & (g139)) + ((g135) & (g136) & (g137) & (!g138) & (!g145) & (!g139)) + ((g135) & (g136) & (g137) & (!g138) & (!g145) & (g139)) + ((g135) & (g136) & (g137) & (!g138) & (g145) & (g139)) + ((g135) & (g136) & (g137) & (g138) & (!g145) & (!g139)) + ((g135) & (g136) & (g137) & (g138) & (!g145) & (g139)) + ((g135) & (g136) & (g137) & (g138) & (g145) & (!g139)) + ((g135) & (g136) & (g137) & (g138) & (g145) & (g139)));
	assign g153 = (((!g135) & (!g136) & (!g137) & (!g138) & (g145) & (!g139)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g145) & (!g139)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g145) & (g139)) + ((!g135) & (!g136) & (g137) & (!g138) & (g145) & (g139)) + ((!g135) & (!g136) & (g137) & (g138) & (!g145) & (g139)) + ((!g135) & (g136) & (!g137) & (!g138) & (!g145) & (!g139)) + ((!g135) & (g136) & (!g137) & (!g138) & (g145) & (!g139)) + ((!g135) & (g136) & (!g137) & (g138) & (!g145) & (g139)) + ((!g135) & (g136) & (g137) & (!g138) & (!g145) & (g139)) + ((!g135) & (g136) & (g137) & (!g138) & (g145) & (!g139)) + ((!g135) & (g136) & (g137) & (!g138) & (g145) & (g139)) + ((!g135) & (g136) & (g137) & (g138) & (g145) & (!g139)) + ((!g135) & (g136) & (g137) & (g138) & (g145) & (g139)) + ((g135) & (!g136) & (!g137) & (!g138) & (!g145) & (!g139)) + ((g135) & (!g136) & (!g137) & (g138) & (!g145) & (!g139)) + ((g135) & (!g136) & (!g137) & (g138) & (!g145) & (g139)) + ((g135) & (!g136) & (!g137) & (g138) & (g145) & (!g139)) + ((g135) & (!g136) & (g137) & (!g138) & (!g145) & (!g139)) + ((g135) & (!g136) & (g137) & (!g138) & (g145) & (g139)) + ((g135) & (!g136) & (g137) & (g138) & (g145) & (!g139)) + ((g135) & (g136) & (!g137) & (!g138) & (!g145) & (!g139)) + ((g135) & (g136) & (!g137) & (g138) & (!g145) & (!g139)) + ((g135) & (g136) & (!g137) & (g138) & (g145) & (!g139)) + ((g135) & (g136) & (!g137) & (g138) & (g145) & (g139)) + ((g135) & (g136) & (g137) & (g138) & (!g145) & (g139)) + ((g135) & (g136) & (g137) & (g138) & (g145) & (g139)));
	assign g154 = (((!g150) & (!g151) & (!g152) & (!g153) & (!g140) & (!g146)) + ((!g150) & (!g151) & (!g152) & (!g153) & (g140) & (!g146)) + ((!g150) & (!g151) & (!g152) & (g153) & (!g140) & (!g146)) + ((!g150) & (!g151) & (!g152) & (g153) & (g140) & (!g146)) + ((!g150) & (!g151) & (!g152) & (g153) & (g140) & (g146)) + ((!g150) & (!g151) & (g152) & (!g153) & (!g140) & (!g146)) + ((!g150) & (!g151) & (g152) & (!g153) & (!g140) & (g146)) + ((!g150) & (!g151) & (g152) & (!g153) & (g140) & (!g146)) + ((!g150) & (!g151) & (g152) & (g153) & (!g140) & (!g146)) + ((!g150) & (!g151) & (g152) & (g153) & (!g140) & (g146)) + ((!g150) & (!g151) & (g152) & (g153) & (g140) & (!g146)) + ((!g150) & (!g151) & (g152) & (g153) & (g140) & (g146)) + ((!g150) & (g151) & (!g152) & (!g153) & (!g140) & (!g146)) + ((!g150) & (g151) & (!g152) & (g153) & (!g140) & (!g146)) + ((!g150) & (g151) & (!g152) & (g153) & (g140) & (g146)) + ((!g150) & (g151) & (g152) & (!g153) & (!g140) & (!g146)) + ((!g150) & (g151) & (g152) & (!g153) & (!g140) & (g146)) + ((!g150) & (g151) & (g152) & (g153) & (!g140) & (!g146)) + ((!g150) & (g151) & (g152) & (g153) & (!g140) & (g146)) + ((!g150) & (g151) & (g152) & (g153) & (g140) & (g146)) + ((g150) & (!g151) & (!g152) & (!g153) & (g140) & (!g146)) + ((g150) & (!g151) & (!g152) & (g153) & (g140) & (!g146)) + ((g150) & (!g151) & (!g152) & (g153) & (g140) & (g146)) + ((g150) & (!g151) & (g152) & (!g153) & (!g140) & (g146)) + ((g150) & (!g151) & (g152) & (!g153) & (g140) & (!g146)) + ((g150) & (!g151) & (g152) & (g153) & (!g140) & (g146)) + ((g150) & (!g151) & (g152) & (g153) & (g140) & (!g146)) + ((g150) & (!g151) & (g152) & (g153) & (g140) & (g146)) + ((g150) & (g151) & (!g152) & (g153) & (g140) & (g146)) + ((g150) & (g151) & (g152) & (!g153) & (!g140) & (g146)) + ((g150) & (g151) & (g152) & (g153) & (!g140) & (g146)) + ((g150) & (g151) & (g152) & (g153) & (g140) & (g146)));
	assign g156 = (((!sk[12]) & (g154) & (!g155)) + ((!sk[12]) & (g154) & (g155)) + ((sk[12]) & (!g154) & (g155)) + ((sk[12]) & (g154) & (!g155)));
	assign g157 = (((!g139) & (!g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((!g139) & (!g136) & (!g137) & (!g138) & (g145) & (g140)) + ((!g139) & (!g136) & (!g137) & (g138) & (!g145) & (g140)) + ((!g139) & (!g136) & (!g137) & (g138) & (g145) & (!g140)) + ((!g139) & (!g136) & (!g137) & (g138) & (g145) & (g140)) + ((!g139) & (!g136) & (g137) & (!g138) & (!g145) & (g140)) + ((!g139) & (!g136) & (g137) & (g138) & (!g145) & (!g140)) + ((!g139) & (!g136) & (g137) & (g138) & (g145) & (!g140)) + ((!g139) & (g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((!g139) & (g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((!g139) & (g136) & (!g137) & (g138) & (!g145) & (g140)) + ((!g139) & (g136) & (g137) & (!g138) & (!g145) & (!g140)) + ((!g139) & (g136) & (g137) & (!g138) & (!g145) & (g140)) + ((!g139) & (g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g139) & (g136) & (g137) & (!g138) & (g145) & (g140)) + ((g139) & (!g136) & (!g137) & (g138) & (!g145) & (g140)) + ((g139) & (!g136) & (!g137) & (g138) & (g145) & (g140)) + ((g139) & (g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((g139) & (g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((g139) & (g136) & (!g137) & (g138) & (g145) & (!g140)) + ((g139) & (g136) & (g137) & (g138) & (!g145) & (!g140)) + ((g139) & (g136) & (g137) & (g138) & (!g145) & (g140)));
	assign g158 = (((!g139) & (!g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((!g139) & (!g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((!g139) & (!g136) & (!g137) & (g138) & (g145) & (g140)) + ((!g139) & (!g136) & (g137) & (!g138) & (!g145) & (!g140)) + ((!g139) & (!g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g139) & (!g136) & (g137) & (g138) & (!g145) & (g140)) + ((!g139) & (g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((!g139) & (g136) & (!g137) & (!g138) & (g145) & (g140)) + ((!g139) & (g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((!g139) & (g136) & (!g137) & (g138) & (!g145) & (g140)) + ((!g139) & (g136) & (!g137) & (g138) & (g145) & (g140)) + ((!g139) & (g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g139) & (g136) & (g137) & (!g138) & (g145) & (g140)) + ((!g139) & (g136) & (g137) & (g138) & (g145) & (!g140)) + ((g139) & (!g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((g139) & (!g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((g139) & (!g136) & (!g137) & (!g138) & (g145) & (g140)) + ((g139) & (!g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((g139) & (!g136) & (!g137) & (g138) & (!g145) & (g140)) + ((g139) & (!g136) & (!g137) & (g138) & (g145) & (!g140)) + ((g139) & (!g136) & (g137) & (g138) & (!g145) & (!g140)) + ((g139) & (g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((g139) & (g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((g139) & (g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((g139) & (g136) & (!g137) & (g138) & (g145) & (!g140)) + ((g139) & (g136) & (!g137) & (g138) & (g145) & (g140)) + ((g139) & (g136) & (g137) & (!g138) & (!g145) & (!g140)) + ((g139) & (g136) & (g137) & (!g138) & (g145) & (!g140)) + ((g139) & (g136) & (g137) & (g138) & (!g145) & (g140)) + ((g139) & (g136) & (g137) & (g138) & (g145) & (g140)));
	assign g159 = (((!g139) & (!g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((!g139) & (!g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((!g139) & (!g136) & (!g137) & (g138) & (!g145) & (g140)) + ((!g139) & (!g136) & (g137) & (!g138) & (!g145) & (g140)) + ((!g139) & (!g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g139) & (!g136) & (g137) & (g138) & (!g145) & (g140)) + ((!g139) & (g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((!g139) & (g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((!g139) & (g136) & (!g137) & (g138) & (g145) & (!g140)) + ((!g139) & (g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g139) & (g136) & (g137) & (g138) & (!g145) & (!g140)) + ((!g139) & (g136) & (g137) & (g138) & (g145) & (!g140)) + ((g139) & (!g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((g139) & (!g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((g139) & (!g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((g139) & (!g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((g139) & (!g136) & (!g137) & (g138) & (!g145) & (g140)) + ((g139) & (!g136) & (!g137) & (g138) & (g145) & (!g140)) + ((g139) & (!g136) & (!g137) & (g138) & (g145) & (g140)) + ((g139) & (!g136) & (g137) & (!g138) & (!g145) & (g140)) + ((g139) & (!g136) & (g137) & (!g138) & (g145) & (!g140)) + ((g139) & (!g136) & (g137) & (g138) & (!g145) & (!g140)) + ((g139) & (!g136) & (g137) & (g138) & (g145) & (g140)) + ((g139) & (g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((g139) & (g136) & (!g137) & (!g138) & (g145) & (g140)) + ((g139) & (g136) & (g137) & (!g138) & (g145) & (g140)) + ((g139) & (g136) & (g137) & (g138) & (!g145) & (!g140)) + ((g139) & (g136) & (g137) & (g138) & (!g145) & (g140)) + ((g139) & (g136) & (g137) & (g138) & (g145) & (g140)));
	assign g160 = (((!g139) & (!g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((!g139) & (!g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((!g139) & (!g136) & (!g137) & (!g138) & (g145) & (g140)) + ((!g139) & (!g136) & (!g137) & (g138) & (!g145) & (g140)) + ((!g139) & (!g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g139) & (!g136) & (g137) & (g138) & (g145) & (g140)) + ((!g139) & (g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((!g139) & (g136) & (!g137) & (g138) & (!g145) & (g140)) + ((!g139) & (g136) & (!g137) & (g138) & (g145) & (g140)) + ((!g139) & (g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g139) & (g136) & (g137) & (!g138) & (g145) & (g140)) + ((!g139) & (g136) & (g137) & (g138) & (!g145) & (!g140)) + ((!g139) & (g136) & (g137) & (g138) & (!g145) & (g140)) + ((!g139) & (g136) & (g137) & (g138) & (g145) & (!g140)) + ((!g139) & (g136) & (g137) & (g138) & (g145) & (g140)) + ((g139) & (!g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((g139) & (!g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((g139) & (!g136) & (!g137) & (!g138) & (g145) & (g140)) + ((g139) & (!g136) & (!g137) & (g138) & (g145) & (g140)) + ((g139) & (!g136) & (g137) & (!g138) & (!g145) & (g140)) + ((g139) & (!g136) & (g137) & (!g138) & (g145) & (!g140)) + ((g139) & (!g136) & (g137) & (g138) & (g145) & (!g140)) + ((g139) & (g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((g139) & (g136) & (!g137) & (g138) & (!g145) & (g140)) + ((g139) & (g136) & (!g137) & (g138) & (g145) & (!g140)) + ((g139) & (g136) & (g137) & (!g138) & (g145) & (g140)) + ((g139) & (g136) & (g137) & (g138) & (!g145) & (!g140)));
	assign g161 = (((!g157) & (!g158) & (!g159) & (!g160) & (!g135) & (g146)) + ((!g157) & (!g158) & (!g159) & (!g160) & (g135) & (!g146)) + ((!g157) & (!g158) & (!g159) & (!g160) & (g135) & (g146)) + ((!g157) & (!g158) & (!g159) & (g160) & (!g135) & (g146)) + ((!g157) & (!g158) & (!g159) & (g160) & (g135) & (!g146)) + ((!g157) & (!g158) & (g159) & (!g160) & (g135) & (!g146)) + ((!g157) & (!g158) & (g159) & (!g160) & (g135) & (g146)) + ((!g157) & (!g158) & (g159) & (g160) & (g135) & (!g146)) + ((!g157) & (g158) & (!g159) & (!g160) & (!g135) & (g146)) + ((!g157) & (g158) & (!g159) & (!g160) & (g135) & (g146)) + ((!g157) & (g158) & (!g159) & (g160) & (!g135) & (g146)) + ((!g157) & (g158) & (g159) & (!g160) & (g135) & (g146)) + ((g157) & (!g158) & (!g159) & (!g160) & (!g135) & (!g146)) + ((g157) & (!g158) & (!g159) & (!g160) & (!g135) & (g146)) + ((g157) & (!g158) & (!g159) & (!g160) & (g135) & (!g146)) + ((g157) & (!g158) & (!g159) & (!g160) & (g135) & (g146)) + ((g157) & (!g158) & (!g159) & (g160) & (!g135) & (!g146)) + ((g157) & (!g158) & (!g159) & (g160) & (!g135) & (g146)) + ((g157) & (!g158) & (!g159) & (g160) & (g135) & (!g146)) + ((g157) & (!g158) & (g159) & (!g160) & (!g135) & (!g146)) + ((g157) & (!g158) & (g159) & (!g160) & (g135) & (!g146)) + ((g157) & (!g158) & (g159) & (!g160) & (g135) & (g146)) + ((g157) & (!g158) & (g159) & (g160) & (!g135) & (!g146)) + ((g157) & (!g158) & (g159) & (g160) & (g135) & (!g146)) + ((g157) & (g158) & (!g159) & (!g160) & (!g135) & (!g146)) + ((g157) & (g158) & (!g159) & (!g160) & (!g135) & (g146)) + ((g157) & (g158) & (!g159) & (!g160) & (g135) & (g146)) + ((g157) & (g158) & (!g159) & (g160) & (!g135) & (!g146)) + ((g157) & (g158) & (!g159) & (g160) & (!g135) & (g146)) + ((g157) & (g158) & (g159) & (!g160) & (!g135) & (!g146)) + ((g157) & (g158) & (g159) & (!g160) & (g135) & (g146)) + ((g157) & (g158) & (g159) & (g160) & (!g135) & (!g146)));
	assign g163 = (((!g161) & (sk[18]) & (g162)) + ((g161) & (!sk[18]) & (!g162)) + ((g161) & (!sk[18]) & (g162)) + ((g161) & (sk[18]) & (!g162)));
	assign g164 = (((!g135) & (!g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (g145) & (g140)) + ((!g135) & (!g136) & (g137) & (g138) & (!g145) & (!g140)) + ((!g135) & (!g136) & (g137) & (g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (g137) & (g138) & (g145) & (g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (g136) & (g137) & (!g138) & (!g145) & (!g140)) + ((!g135) & (g136) & (g137) & (g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((g135) & (!g136) & (g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (g137) & (!g138) & (!g145) & (g140)) + ((g135) & (!g136) & (g137) & (!g138) & (g145) & (!g140)) + ((g135) & (!g136) & (g137) & (g138) & (!g145) & (g140)) + ((g135) & (g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((g135) & (g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((g135) & (g136) & (!g137) & (g138) & (g145) & (!g140)) + ((g135) & (g136) & (g137) & (!g138) & (!g145) & (g140)) + ((g135) & (g136) & (g137) & (!g138) & (g145) & (g140)));
	assign g165 = (((!g135) & (!g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (!g137) & (!g138) & (g145) & (g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (g137) & (g138) & (!g145) & (!g140)) + ((!g135) & (!g136) & (g137) & (g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (g137) & (g138) & (g145) & (g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (g145) & (g140)) + ((!g135) & (g136) & (!g137) & (g138) & (g145) & (g140)) + ((!g135) & (g136) & (g137) & (!g138) & (!g145) & (!g140)) + ((!g135) & (g136) & (g137) & (!g138) & (!g145) & (g140)) + ((!g135) & (g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (g136) & (g137) & (g138) & (!g145) & (g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((g135) & (!g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (!g137) & (g138) & (!g145) & (g140)) + ((g135) & (!g136) & (!g137) & (g138) & (g145) & (g140)) + ((g135) & (!g136) & (g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (g137) & (!g138) & (!g145) & (g140)) + ((g135) & (!g136) & (g137) & (!g138) & (g145) & (g140)) + ((g135) & (!g136) & (g137) & (g138) & (!g145) & (g140)) + ((g135) & (g136) & (!g137) & (g138) & (!g145) & (g140)) + ((g135) & (g136) & (!g137) & (g138) & (g145) & (!g140)) + ((g135) & (g136) & (g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (g136) & (g137) & (g138) & (!g145) & (!g140)));
	assign g166 = (((!g135) & (!g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (!g137) & (!g138) & (g145) & (g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (g137) & (!g138) & (g145) & (g140)) + ((!g135) & (!g136) & (g137) & (g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (g137) & (g138) & (g145) & (g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (g145) & (g140)) + ((!g135) & (g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((!g135) & (g136) & (!g137) & (g138) & (!g145) & (g140)) + ((!g135) & (g136) & (g137) & (!g138) & (!g145) & (g140)) + ((!g135) & (g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (g136) & (g137) & (g138) & (g145) & (g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (g145) & (g140)) + ((g135) & (!g136) & (!g137) & (g138) & (g145) & (g140)) + ((g135) & (!g136) & (g137) & (g138) & (!g145) & (!g140)) + ((g135) & (g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((g135) & (g136) & (!g137) & (g138) & (g145) & (g140)) + ((g135) & (g136) & (g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (g136) & (g137) & (!g138) & (!g145) & (g140)) + ((g135) & (g136) & (g137) & (!g138) & (g145) & (g140)) + ((g135) & (g136) & (g137) & (g138) & (!g145) & (!g140)) + ((g135) & (g136) & (g137) & (g138) & (g145) & (g140)));
	assign g167 = (((!g135) & (!g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (!g137) & (g138) & (g145) & (g140)) + ((!g135) & (!g136) & (g137) & (g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (g137) & (g138) & (g145) & (g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (!g145) & (!g140)) + ((!g135) & (g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (g136) & (!g137) & (g138) & (!g145) & (!g140)) + ((!g135) & (g136) & (!g137) & (g138) & (!g145) & (g140)) + ((!g135) & (g136) & (!g137) & (g138) & (g145) & (!g140)) + ((!g135) & (g136) & (g137) & (!g138) & (!g145) & (!g140)) + ((!g135) & (g136) & (g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (g136) & (g137) & (!g138) & (g145) & (g140)) + ((g135) & (!g136) & (!g137) & (!g138) & (g145) & (g140)) + ((g135) & (!g136) & (!g137) & (g138) & (g145) & (!g140)) + ((g135) & (!g136) & (g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (g137) & (!g138) & (g145) & (!g140)) + ((g135) & (!g136) & (g137) & (!g138) & (g145) & (g140)) + ((g135) & (!g136) & (g137) & (g138) & (!g145) & (g140)) + ((g135) & (!g136) & (g137) & (g138) & (g145) & (!g140)) + ((g135) & (!g136) & (g137) & (g138) & (g145) & (g140)) + ((g135) & (g136) & (!g137) & (!g138) & (!g145) & (g140)) + ((g135) & (g136) & (!g137) & (!g138) & (g145) & (!g140)) + ((g135) & (g136) & (g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (g136) & (g137) & (!g138) & (!g145) & (g140)) + ((g135) & (g136) & (g137) & (g138) & (g145) & (g140)));
	assign g168 = (((!g164) & (!g165) & (!g166) & (!g167) & (!g146) & (g139)) + ((!g164) & (!g165) & (!g166) & (!g167) & (g146) & (!g139)) + ((!g164) & (!g165) & (!g166) & (!g167) & (g146) & (g139)) + ((!g164) & (!g165) & (!g166) & (g167) & (!g146) & (g139)) + ((!g164) & (!g165) & (!g166) & (g167) & (g146) & (!g139)) + ((!g164) & (!g165) & (g166) & (!g167) & (g146) & (!g139)) + ((!g164) & (!g165) & (g166) & (!g167) & (g146) & (g139)) + ((!g164) & (!g165) & (g166) & (g167) & (g146) & (!g139)) + ((!g164) & (g165) & (!g166) & (!g167) & (!g146) & (g139)) + ((!g164) & (g165) & (!g166) & (!g167) & (g146) & (g139)) + ((!g164) & (g165) & (!g166) & (g167) & (!g146) & (g139)) + ((!g164) & (g165) & (g166) & (!g167) & (g146) & (g139)) + ((g164) & (!g165) & (!g166) & (!g167) & (!g146) & (!g139)) + ((g164) & (!g165) & (!g166) & (!g167) & (!g146) & (g139)) + ((g164) & (!g165) & (!g166) & (!g167) & (g146) & (!g139)) + ((g164) & (!g165) & (!g166) & (!g167) & (g146) & (g139)) + ((g164) & (!g165) & (!g166) & (g167) & (!g146) & (!g139)) + ((g164) & (!g165) & (!g166) & (g167) & (!g146) & (g139)) + ((g164) & (!g165) & (!g166) & (g167) & (g146) & (!g139)) + ((g164) & (!g165) & (g166) & (!g167) & (!g146) & (!g139)) + ((g164) & (!g165) & (g166) & (!g167) & (g146) & (!g139)) + ((g164) & (!g165) & (g166) & (!g167) & (g146) & (g139)) + ((g164) & (!g165) & (g166) & (g167) & (!g146) & (!g139)) + ((g164) & (!g165) & (g166) & (g167) & (g146) & (!g139)) + ((g164) & (g165) & (!g166) & (!g167) & (!g146) & (!g139)) + ((g164) & (g165) & (!g166) & (!g167) & (!g146) & (g139)) + ((g164) & (g165) & (!g166) & (!g167) & (g146) & (g139)) + ((g164) & (g165) & (!g166) & (g167) & (!g146) & (!g139)) + ((g164) & (g165) & (!g166) & (g167) & (!g146) & (g139)) + ((g164) & (g165) & (g166) & (!g167) & (!g146) & (!g139)) + ((g164) & (g165) & (g166) & (!g167) & (g146) & (g139)) + ((g164) & (g165) & (g166) & (g167) & (!g146) & (!g139)));
	assign g170 = (((!g168) & (sk[24]) & (g169)) + ((g168) & (!sk[24]) & (!g169)) + ((g168) & (!sk[24]) & (g169)) + ((g168) & (sk[24]) & (!g169)));
	assign g171 = (((!g135) & (!g136) & (!g139) & (!g146) & (!g145) & (g140)) + ((!g135) & (!g136) & (g139) & (!g146) & (!g145) & (g140)) + ((!g135) & (!g136) & (g139) & (!g146) & (g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (!g146) & (g145) & (g140)) + ((!g135) & (!g136) & (g139) & (g146) & (!g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (g146) & (g145) & (!g140)) + ((!g135) & (g136) & (!g139) & (!g146) & (!g145) & (!g140)) + ((!g135) & (g136) & (!g139) & (!g146) & (!g145) & (g140)) + ((!g135) & (g136) & (!g139) & (g146) & (!g145) & (!g140)) + ((!g135) & (g136) & (!g139) & (g146) & (!g145) & (g140)) + ((!g135) & (g136) & (!g139) & (g146) & (g145) & (g140)) + ((!g135) & (g136) & (g139) & (g146) & (!g145) & (g140)) + ((!g135) & (g136) & (g139) & (g146) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g146) & (!g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g146) & (!g145) & (g140)) + ((g135) & (!g136) & (!g139) & (g146) & (!g145) & (g140)) + ((g135) & (!g136) & (g139) & (!g146) & (g145) & (!g140)) + ((g135) & (!g136) & (g139) & (g146) & (!g145) & (!g140)) + ((g135) & (!g136) & (g139) & (g146) & (!g145) & (g140)) + ((g135) & (!g136) & (g139) & (g146) & (g145) & (!g140)) + ((g135) & (g136) & (!g139) & (!g146) & (!g145) & (!g140)) + ((g135) & (g136) & (!g139) & (!g146) & (g145) & (!g140)) + ((g135) & (g136) & (!g139) & (g146) & (g145) & (!g140)) + ((g135) & (g136) & (g139) & (!g146) & (!g145) & (!g140)) + ((g135) & (g136) & (g139) & (!g146) & (!g145) & (g140)) + ((g135) & (g136) & (g139) & (g146) & (!g145) & (g140)));
	assign g172 = (((!g135) & (!g136) & (!g139) & (!g146) & (!g145) & (!g140)) + ((!g135) & (!g136) & (!g139) & (!g146) & (!g145) & (g140)) + ((!g135) & (!g136) & (!g139) & (!g146) & (g145) & (!g140)) + ((!g135) & (!g136) & (!g139) & (!g146) & (g145) & (g140)) + ((!g135) & (!g136) & (!g139) & (g146) & (!g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (!g146) & (!g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (!g146) & (g145) & (g140)) + ((!g135) & (!g136) & (g139) & (g146) & (!g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (g146) & (g145) & (g140)) + ((!g135) & (g136) & (!g139) & (!g146) & (!g145) & (g140)) + ((!g135) & (g136) & (!g139) & (g146) & (g145) & (!g140)) + ((!g135) & (g136) & (g139) & (!g146) & (!g145) & (!g140)) + ((!g135) & (g136) & (g139) & (!g146) & (!g145) & (g140)) + ((!g135) & (g136) & (g139) & (!g146) & (g145) & (!g140)) + ((!g135) & (g136) & (g139) & (!g146) & (g145) & (g140)) + ((!g135) & (g136) & (g139) & (g146) & (!g145) & (!g140)) + ((!g135) & (g136) & (g139) & (g146) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g146) & (!g145) & (g140)) + ((g135) & (!g136) & (!g139) & (!g146) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g146) & (g145) & (g140)) + ((g135) & (!g136) & (!g139) & (g146) & (!g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (g146) & (g145) & (g140)) + ((g135) & (!g136) & (g139) & (!g146) & (g145) & (!g140)) + ((g135) & (!g136) & (g139) & (!g146) & (g145) & (g140)) + ((g135) & (!g136) & (g139) & (g146) & (!g145) & (g140)) + ((g135) & (g136) & (!g139) & (!g146) & (g145) & (!g140)) + ((g135) & (g136) & (!g139) & (!g146) & (g145) & (g140)) + ((g135) & (g136) & (!g139) & (g146) & (!g145) & (!g140)) + ((g135) & (g136) & (!g139) & (g146) & (!g145) & (g140)) + ((g135) & (g136) & (g139) & (!g146) & (g145) & (!g140)) + ((g135) & (g136) & (g139) & (!g146) & (g145) & (g140)) + ((g135) & (g136) & (g139) & (g146) & (!g145) & (g140)));
	assign g173 = (((!g135) & (!g136) & (!g139) & (!g146) & (!g145) & (!g140)) + ((!g135) & (!g136) & (!g139) & (!g146) & (!g145) & (g140)) + ((!g135) & (!g136) & (g139) & (!g146) & (!g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (!g146) & (g145) & (g140)) + ((!g135) & (!g136) & (g139) & (g146) & (!g145) & (g140)) + ((!g135) & (g136) & (!g139) & (g146) & (!g145) & (!g140)) + ((!g135) & (g136) & (!g139) & (g146) & (g145) & (!g140)) + ((!g135) & (g136) & (!g139) & (g146) & (g145) & (g140)) + ((!g135) & (g136) & (g139) & (!g146) & (!g145) & (!g140)) + ((!g135) & (g136) & (g139) & (!g146) & (g145) & (!g140)) + ((!g135) & (g136) & (g139) & (!g146) & (g145) & (g140)) + ((!g135) & (g136) & (g139) & (g146) & (!g145) & (!g140)) + ((!g135) & (g136) & (g139) & (g146) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g146) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g146) & (g145) & (g140)) + ((g135) & (!g136) & (!g139) & (g146) & (!g145) & (g140)) + ((g135) & (!g136) & (!g139) & (g146) & (g145) & (g140)) + ((g135) & (!g136) & (g139) & (!g146) & (!g145) & (!g140)) + ((g135) & (!g136) & (g139) & (!g146) & (!g145) & (g140)) + ((g135) & (!g136) & (g139) & (!g146) & (g145) & (g140)) + ((g135) & (!g136) & (g139) & (g146) & (!g145) & (!g140)) + ((g135) & (!g136) & (g139) & (g146) & (!g145) & (g140)) + ((g135) & (!g136) & (g139) & (g146) & (g145) & (!g140)) + ((g135) & (!g136) & (g139) & (g146) & (g145) & (g140)) + ((g135) & (g136) & (!g139) & (!g146) & (!g145) & (g140)) + ((g135) & (g136) & (!g139) & (g146) & (!g145) & (!g140)) + ((g135) & (g136) & (!g139) & (g146) & (g145) & (!g140)) + ((g135) & (g136) & (g139) & (!g146) & (!g145) & (!g140)) + ((g135) & (g136) & (g139) & (!g146) & (!g145) & (g140)) + ((g135) & (g136) & (g139) & (!g146) & (g145) & (!g140)) + ((g135) & (g136) & (g139) & (g146) & (!g145) & (!g140)) + ((g135) & (g136) & (g139) & (g146) & (g145) & (!g140)));
	assign g174 = (((!g135) & (!g136) & (!g139) & (!g146) & (g145) & (g140)) + ((!g135) & (!g136) & (!g139) & (g146) & (!g145) & (!g140)) + ((!g135) & (!g136) & (!g139) & (g146) & (g145) & (g140)) + ((!g135) & (!g136) & (g139) & (!g146) & (!g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (!g146) & (g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (g146) & (!g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (g146) & (!g145) & (g140)) + ((!g135) & (!g136) & (g139) & (g146) & (g145) & (!g140)) + ((!g135) & (g136) & (!g139) & (!g146) & (!g145) & (!g140)) + ((!g135) & (g136) & (!g139) & (g146) & (!g145) & (g140)) + ((!g135) & (g136) & (!g139) & (g146) & (g145) & (!g140)) + ((!g135) & (g136) & (!g139) & (g146) & (g145) & (g140)) + ((!g135) & (g136) & (g139) & (!g146) & (!g145) & (!g140)) + ((!g135) & (g136) & (g139) & (g146) & (!g145) & (!g140)) + ((!g135) & (g136) & (g139) & (g146) & (!g145) & (g140)) + ((g135) & (!g136) & (!g139) & (!g146) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g146) & (g145) & (g140)) + ((g135) & (!g136) & (g139) & (!g146) & (!g145) & (!g140)) + ((g135) & (!g136) & (g139) & (!g146) & (g145) & (!g140)) + ((g135) & (!g136) & (g139) & (g146) & (g145) & (!g140)) + ((g135) & (g136) & (!g139) & (!g146) & (g145) & (!g140)) + ((g135) & (g136) & (!g139) & (g146) & (g145) & (g140)) + ((g135) & (g136) & (g139) & (!g146) & (!g145) & (!g140)) + ((g135) & (g136) & (g139) & (!g146) & (!g145) & (g140)) + ((g135) & (g136) & (g139) & (!g146) & (g145) & (!g140)) + ((g135) & (g136) & (g139) & (g146) & (!g145) & (!g140)));
	assign g175 = (((!g171) & (!g172) & (!g173) & (!g174) & (g137) & (g138)) + ((!g171) & (!g172) & (g173) & (!g174) & (!g137) & (g138)) + ((!g171) & (!g172) & (g173) & (!g174) & (g137) & (g138)) + ((!g171) & (!g172) & (g173) & (g174) & (!g137) & (g138)) + ((!g171) & (g172) & (!g173) & (!g174) & (g137) & (!g138)) + ((!g171) & (g172) & (!g173) & (!g174) & (g137) & (g138)) + ((!g171) & (g172) & (!g173) & (g174) & (g137) & (!g138)) + ((!g171) & (g172) & (g173) & (!g174) & (!g137) & (g138)) + ((!g171) & (g172) & (g173) & (!g174) & (g137) & (!g138)) + ((!g171) & (g172) & (g173) & (!g174) & (g137) & (g138)) + ((!g171) & (g172) & (g173) & (g174) & (!g137) & (g138)) + ((!g171) & (g172) & (g173) & (g174) & (g137) & (!g138)) + ((g171) & (!g172) & (!g173) & (!g174) & (!g137) & (!g138)) + ((g171) & (!g172) & (!g173) & (!g174) & (g137) & (g138)) + ((g171) & (!g172) & (!g173) & (g174) & (!g137) & (!g138)) + ((g171) & (!g172) & (g173) & (!g174) & (!g137) & (!g138)) + ((g171) & (!g172) & (g173) & (!g174) & (!g137) & (g138)) + ((g171) & (!g172) & (g173) & (!g174) & (g137) & (g138)) + ((g171) & (!g172) & (g173) & (g174) & (!g137) & (!g138)) + ((g171) & (!g172) & (g173) & (g174) & (!g137) & (g138)) + ((g171) & (g172) & (!g173) & (!g174) & (!g137) & (!g138)) + ((g171) & (g172) & (!g173) & (!g174) & (g137) & (!g138)) + ((g171) & (g172) & (!g173) & (!g174) & (g137) & (g138)) + ((g171) & (g172) & (!g173) & (g174) & (!g137) & (!g138)) + ((g171) & (g172) & (!g173) & (g174) & (g137) & (!g138)) + ((g171) & (g172) & (g173) & (!g174) & (!g137) & (!g138)) + ((g171) & (g172) & (g173) & (!g174) & (!g137) & (g138)) + ((g171) & (g172) & (g173) & (!g174) & (g137) & (!g138)) + ((g171) & (g172) & (g173) & (!g174) & (g137) & (g138)) + ((g171) & (g172) & (g173) & (g174) & (!g137) & (!g138)) + ((g171) & (g172) & (g173) & (g174) & (!g137) & (g138)) + ((g171) & (g172) & (g173) & (g174) & (g137) & (!g138)));
	assign g177 = (((!g175) & (sk[30]) & (g176)) + ((g175) & (!sk[30]) & (!g176)) + ((g175) & (!sk[30]) & (g176)) + ((g175) & (sk[30]) & (!g176)));
	assign g178 = (((!g135) & (!g136) & (!g139) & (!g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (!g139) & (!g138) & (g145) & (g140)) + ((!g135) & (!g136) & (!g139) & (g138) & (g145) & (g140)) + ((!g135) & (!g136) & (g139) & (!g138) & (!g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (!g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (g139) & (!g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (!g138) & (g145) & (g140)) + ((!g135) & (!g136) & (g139) & (g138) & (!g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (g138) & (!g145) & (g140)) + ((!g135) & (g136) & (!g139) & (!g138) & (!g145) & (g140)) + ((!g135) & (g136) & (!g139) & (!g138) & (g145) & (!g140)) + ((!g135) & (g136) & (!g139) & (g138) & (g145) & (g140)) + ((!g135) & (g136) & (g139) & (!g138) & (g145) & (!g140)) + ((!g135) & (g136) & (g139) & (!g138) & (g145) & (g140)) + ((!g135) & (g136) & (g139) & (g138) & (!g145) & (!g140)) + ((!g135) & (g136) & (g139) & (g138) & (!g145) & (g140)) + ((!g135) & (g136) & (g139) & (g138) & (g145) & (g140)) + ((g135) & (!g136) & (!g139) & (!g138) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g138) & (g145) & (g140)) + ((g135) & (!g136) & (!g139) & (g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (g138) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (g138) & (g145) & (g140)) + ((g135) & (!g136) & (g139) & (!g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (g139) & (!g138) & (g145) & (!g140)) + ((g135) & (!g136) & (g139) & (g138) & (g145) & (!g140)) + ((g135) & (g136) & (!g139) & (!g138) & (g145) & (g140)) + ((g135) & (g136) & (g139) & (!g138) & (!g145) & (!g140)) + ((g135) & (g136) & (g139) & (!g138) & (g145) & (g140)));
	assign g179 = (((!g135) & (!g136) & (!g139) & (!g138) & (!g145) & (!g140)) + ((!g135) & (!g136) & (!g139) & (g138) & (!g145) & (!g140)) + ((!g135) & (!g136) & (!g139) & (g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (!g139) & (g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (!g138) & (g145) & (g140)) + ((!g135) & (!g136) & (g139) & (g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (g139) & (g138) & (g145) & (g140)) + ((!g135) & (g136) & (!g139) & (!g138) & (!g145) & (!g140)) + ((!g135) & (g136) & (!g139) & (!g138) & (g145) & (!g140)) + ((!g135) & (g136) & (g139) & (!g138) & (!g145) & (g140)) + ((!g135) & (g136) & (g139) & (!g138) & (g145) & (g140)) + ((!g135) & (g136) & (g139) & (g138) & (!g145) & (g140)) + ((!g135) & (g136) & (g139) & (g138) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g138) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g138) & (g145) & (g140)) + ((g135) & (!g136) & (!g139) & (g138) & (!g145) & (g140)) + ((g135) & (!g136) & (!g139) & (g138) & (g145) & (g140)) + ((g135) & (!g136) & (g139) & (g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (g139) & (g138) & (!g145) & (g140)) + ((g135) & (!g136) & (g139) & (g138) & (g145) & (g140)) + ((g135) & (g136) & (!g139) & (!g138) & (!g145) & (g140)) + ((g135) & (g136) & (!g139) & (!g138) & (g145) & (!g140)) + ((g135) & (g136) & (!g139) & (g138) & (g145) & (!g140)) + ((g135) & (g136) & (g139) & (!g138) & (!g145) & (g140)) + ((g135) & (g136) & (g139) & (!g138) & (g145) & (g140)) + ((g135) & (g136) & (g139) & (g138) & (!g145) & (!g140)) + ((g135) & (g136) & (g139) & (g138) & (g145) & (g140)));
	assign g180 = (((!g135) & (!g136) & (!g139) & (!g138) & (g145) & (g140)) + ((!g135) & (!g136) & (!g139) & (g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (!g138) & (!g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (!g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (g139) & (!g138) & (g145) & (g140)) + ((!g135) & (!g136) & (g139) & (g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (g139) & (g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (g139) & (g138) & (g145) & (g140)) + ((!g135) & (g136) & (!g139) & (!g138) & (g145) & (!g140)) + ((!g135) & (g136) & (!g139) & (!g138) & (g145) & (g140)) + ((!g135) & (g136) & (g139) & (!g138) & (!g145) & (!g140)) + ((!g135) & (g136) & (g139) & (g138) & (!g145) & (g140)) + ((!g135) & (g136) & (g139) & (g138) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g138) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (!g138) & (g145) & (g140)) + ((g135) & (!g136) & (!g139) & (g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (g138) & (!g145) & (g140)) + ((g135) & (!g136) & (g139) & (!g138) & (!g145) & (g140)) + ((g135) & (!g136) & (g139) & (!g138) & (g145) & (g140)) + ((g135) & (!g136) & (g139) & (g138) & (g145) & (!g140)) + ((g135) & (g136) & (!g139) & (!g138) & (!g145) & (!g140)) + ((g135) & (g136) & (!g139) & (!g138) & (!g145) & (g140)) + ((g135) & (g136) & (!g139) & (!g138) & (g145) & (g140)) + ((g135) & (g136) & (!g139) & (g138) & (!g145) & (g140)) + ((g135) & (g136) & (!g139) & (g138) & (g145) & (!g140)) + ((g135) & (g136) & (g139) & (!g138) & (!g145) & (g140)) + ((g135) & (g136) & (g139) & (!g138) & (g145) & (!g140)) + ((g135) & (g136) & (g139) & (g138) & (!g145) & (!g140)) + ((g135) & (g136) & (g139) & (g138) & (g145) & (!g140)) + ((g135) & (g136) & (g139) & (g138) & (g145) & (g140)));
	assign g181 = (((!g135) & (!g136) & (!g139) & (!g138) & (g145) & (!g140)) + ((!g135) & (!g136) & (!g139) & (g138) & (!g145) & (!g140)) + ((!g135) & (!g136) & (!g139) & (g138) & (g145) & (g140)) + ((!g135) & (!g136) & (g139) & (!g138) & (!g145) & (g140)) + ((!g135) & (!g136) & (g139) & (!g138) & (g145) & (g140)) + ((!g135) & (!g136) & (g139) & (g138) & (g145) & (g140)) + ((!g135) & (g136) & (!g139) & (!g138) & (!g145) & (g140)) + ((!g135) & (g136) & (!g139) & (g138) & (!g145) & (g140)) + ((!g135) & (g136) & (!g139) & (g138) & (g145) & (g140)) + ((!g135) & (g136) & (g139) & (!g138) & (!g145) & (!g140)) + ((!g135) & (g136) & (g139) & (!g138) & (g145) & (!g140)) + ((!g135) & (g136) & (g139) & (g138) & (!g145) & (g140)) + ((!g135) & (g136) & (g139) & (g138) & (g145) & (g140)) + ((g135) & (!g136) & (!g139) & (!g138) & (g145) & (!g140)) + ((g135) & (!g136) & (!g139) & (g138) & (g145) & (g140)) + ((g135) & (!g136) & (g139) & (!g138) & (!g145) & (!g140)) + ((g135) & (!g136) & (g139) & (!g138) & (g145) & (g140)) + ((g135) & (!g136) & (g139) & (g138) & (!g145) & (!g140)) + ((g135) & (g136) & (!g139) & (!g138) & (g145) & (g140)) + ((g135) & (g136) & (!g139) & (g138) & (!g145) & (!g140)) + ((g135) & (g136) & (!g139) & (g138) & (!g145) & (g140)) + ((g135) & (g136) & (g139) & (!g138) & (g145) & (g140)));
	assign g182 = (((!g178) & (!g179) & (!g180) & (!g181) & (!g146) & (!g137)) + ((!g178) & (!g179) & (!g180) & (!g181) & (!g146) & (g137)) + ((!g178) & (!g179) & (!g180) & (!g181) & (g146) & (!g137)) + ((!g178) & (!g179) & (!g180) & (g181) & (!g146) & (!g137)) + ((!g178) & (!g179) & (!g180) & (g181) & (!g146) & (g137)) + ((!g178) & (!g179) & (!g180) & (g181) & (g146) & (!g137)) + ((!g178) & (!g179) & (!g180) & (g181) & (g146) & (g137)) + ((!g178) & (!g179) & (g180) & (!g181) & (!g146) & (!g137)) + ((!g178) & (!g179) & (g180) & (!g181) & (g146) & (!g137)) + ((!g178) & (!g179) & (g180) & (g181) & (!g146) & (!g137)) + ((!g178) & (!g179) & (g180) & (g181) & (g146) & (!g137)) + ((!g178) & (!g179) & (g180) & (g181) & (g146) & (g137)) + ((!g178) & (g179) & (!g180) & (!g181) & (!g146) & (!g137)) + ((!g178) & (g179) & (!g180) & (!g181) & (!g146) & (g137)) + ((!g178) & (g179) & (!g180) & (g181) & (!g146) & (!g137)) + ((!g178) & (g179) & (!g180) & (g181) & (!g146) & (g137)) + ((!g178) & (g179) & (!g180) & (g181) & (g146) & (g137)) + ((!g178) & (g179) & (g180) & (!g181) & (!g146) & (!g137)) + ((!g178) & (g179) & (g180) & (g181) & (!g146) & (!g137)) + ((!g178) & (g179) & (g180) & (g181) & (g146) & (g137)) + ((g178) & (!g179) & (!g180) & (!g181) & (!g146) & (g137)) + ((g178) & (!g179) & (!g180) & (!g181) & (g146) & (!g137)) + ((g178) & (!g179) & (!g180) & (g181) & (!g146) & (g137)) + ((g178) & (!g179) & (!g180) & (g181) & (g146) & (!g137)) + ((g178) & (!g179) & (!g180) & (g181) & (g146) & (g137)) + ((g178) & (!g179) & (g180) & (!g181) & (g146) & (!g137)) + ((g178) & (!g179) & (g180) & (g181) & (g146) & (!g137)) + ((g178) & (!g179) & (g180) & (g181) & (g146) & (g137)) + ((g178) & (g179) & (!g180) & (!g181) & (!g146) & (g137)) + ((g178) & (g179) & (!g180) & (g181) & (!g146) & (g137)) + ((g178) & (g179) & (!g180) & (g181) & (g146) & (g137)) + ((g178) & (g179) & (g180) & (g181) & (g146) & (g137)));
	assign g184 = (((!sk[36]) & (g182) & (!g183)) + ((!sk[36]) & (g182) & (g183)) + ((sk[36]) & (!g182) & (g183)) + ((sk[36]) & (g182) & (!g183)));
	assign g185 = (((!g135) & (!g146) & (!g137) & (!g138) & (!g145) & (g140)) + ((!g135) & (!g146) & (!g137) & (!g138) & (g145) & (g140)) + ((!g135) & (!g146) & (!g137) & (g138) & (!g145) & (!g140)) + ((!g135) & (!g146) & (!g137) & (g138) & (!g145) & (g140)) + ((!g135) & (!g146) & (!g137) & (g138) & (g145) & (!g140)) + ((!g135) & (!g146) & (!g137) & (g138) & (g145) & (g140)) + ((!g135) & (!g146) & (g137) & (!g138) & (!g145) & (g140)) + ((!g135) & (!g146) & (g137) & (!g138) & (g145) & (g140)) + ((!g135) & (!g146) & (g137) & (g138) & (g145) & (!g140)) + ((!g135) & (g146) & (g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (g146) & (g137) & (!g138) & (g145) & (g140)) + ((!g135) & (g146) & (g137) & (g138) & (!g145) & (g140)) + ((g135) & (!g146) & (!g137) & (!g138) & (g145) & (!g140)) + ((g135) & (!g146) & (!g137) & (g138) & (!g145) & (!g140)) + ((g135) & (!g146) & (!g137) & (g138) & (!g145) & (g140)) + ((g135) & (!g146) & (!g137) & (g138) & (g145) & (g140)) + ((g135) & (!g146) & (g137) & (!g138) & (!g145) & (g140)) + ((g135) & (!g146) & (g137) & (!g138) & (g145) & (g140)) + ((g135) & (!g146) & (g137) & (g138) & (g145) & (!g140)) + ((g135) & (!g146) & (g137) & (g138) & (g145) & (g140)) + ((g135) & (g146) & (!g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (g146) & (!g137) & (!g138) & (!g145) & (g140)) + ((g135) & (g146) & (!g137) & (!g138) & (g145) & (!g140)) + ((g135) & (g146) & (!g137) & (g138) & (!g145) & (!g140)) + ((g135) & (g146) & (g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (g146) & (g137) & (!g138) & (!g145) & (g140)) + ((g135) & (g146) & (g137) & (!g138) & (g145) & (!g140)) + ((g135) & (g146) & (g137) & (g138) & (!g145) & (g140)));
	assign g186 = (((!g135) & (!g146) & (!g137) & (!g138) & (!g145) & (!g140)) + ((!g135) & (!g146) & (!g137) & (g138) & (g145) & (g140)) + ((!g135) & (!g146) & (g137) & (!g138) & (!g145) & (!g140)) + ((!g135) & (!g146) & (g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (!g146) & (g137) & (!g138) & (g145) & (g140)) + ((!g135) & (!g146) & (g137) & (g138) & (!g145) & (!g140)) + ((!g135) & (!g146) & (g137) & (g138) & (g145) & (g140)) + ((!g135) & (g146) & (!g137) & (!g138) & (!g145) & (!g140)) + ((!g135) & (g146) & (!g137) & (!g138) & (g145) & (g140)) + ((!g135) & (g146) & (!g137) & (g138) & (!g145) & (g140)) + ((!g135) & (g146) & (g137) & (!g138) & (!g145) & (!g140)) + ((!g135) & (g146) & (g137) & (!g138) & (g145) & (g140)) + ((!g135) & (g146) & (g137) & (g138) & (g145) & (!g140)) + ((!g135) & (g146) & (g137) & (g138) & (g145) & (g140)) + ((g135) & (!g146) & (!g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (!g146) & (!g137) & (!g138) & (g145) & (g140)) + ((g135) & (!g146) & (!g137) & (g138) & (!g145) & (!g140)) + ((g135) & (!g146) & (!g137) & (g138) & (g145) & (g140)) + ((g135) & (!g146) & (g137) & (!g138) & (g145) & (g140)) + ((g135) & (!g146) & (g137) & (g138) & (!g145) & (g140)) + ((g135) & (g146) & (!g137) & (!g138) & (g145) & (!g140)) + ((g135) & (g146) & (!g137) & (!g138) & (g145) & (g140)) + ((g135) & (g146) & (!g137) & (g138) & (!g145) & (g140)) + ((g135) & (g146) & (!g137) & (g138) & (g145) & (!g140)) + ((g135) & (g146) & (!g137) & (g138) & (g145) & (g140)) + ((g135) & (g146) & (g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (g146) & (g137) & (!g138) & (g145) & (!g140)) + ((g135) & (g146) & (g137) & (g138) & (!g145) & (!g140)));
	assign g187 = (((!g135) & (!g146) & (!g137) & (!g138) & (!g145) & (g140)) + ((!g135) & (!g146) & (!g137) & (!g138) & (g145) & (g140)) + ((!g135) & (!g146) & (!g137) & (g138) & (g145) & (!g140)) + ((!g135) & (!g146) & (!g137) & (g138) & (g145) & (g140)) + ((!g135) & (!g146) & (g137) & (!g138) & (g145) & (g140)) + ((!g135) & (!g146) & (g137) & (g138) & (!g145) & (!g140)) + ((!g135) & (!g146) & (g137) & (g138) & (!g145) & (g140)) + ((!g135) & (!g146) & (g137) & (g138) & (g145) & (g140)) + ((!g135) & (g146) & (!g137) & (!g138) & (!g145) & (!g140)) + ((!g135) & (g146) & (!g137) & (!g138) & (!g145) & (g140)) + ((!g135) & (g146) & (!g137) & (!g138) & (g145) & (g140)) + ((!g135) & (g146) & (!g137) & (g138) & (!g145) & (g140)) + ((!g135) & (g146) & (!g137) & (g138) & (g145) & (!g140)) + ((!g135) & (g146) & (g137) & (!g138) & (!g145) & (g140)) + ((!g135) & (g146) & (g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (g146) & (g137) & (g138) & (!g145) & (!g140)) + ((!g135) & (g146) & (g137) & (g138) & (g145) & (!g140)) + ((!g135) & (g146) & (g137) & (g138) & (g145) & (g140)) + ((g135) & (!g146) & (!g137) & (!g138) & (!g145) & (g140)) + ((g135) & (!g146) & (!g137) & (g138) & (!g145) & (!g140)) + ((g135) & (!g146) & (!g137) & (g138) & (g145) & (!g140)) + ((g135) & (!g146) & (g137) & (!g138) & (g145) & (g140)) + ((g135) & (!g146) & (g137) & (g138) & (!g145) & (g140)) + ((g135) & (g146) & (!g137) & (!g138) & (!g145) & (g140)) + ((g135) & (g146) & (!g137) & (g138) & (!g145) & (!g140)) + ((g135) & (g146) & (!g137) & (g138) & (g145) & (!g140)) + ((g135) & (g146) & (g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (g146) & (g137) & (!g138) & (g145) & (!g140)) + ((g135) & (g146) & (g137) & (!g138) & (g145) & (g140)) + ((g135) & (g146) & (g137) & (g138) & (g145) & (g140)));
	assign g188 = (((!g135) & (!g146) & (!g137) & (!g138) & (g145) & (g140)) + ((!g135) & (!g146) & (!g137) & (g138) & (!g145) & (!g140)) + ((!g135) & (!g146) & (!g137) & (g138) & (g145) & (g140)) + ((!g135) & (!g146) & (g137) & (!g138) & (!g145) & (!g140)) + ((!g135) & (!g146) & (g137) & (g138) & (g145) & (!g140)) + ((!g135) & (!g146) & (g137) & (g138) & (g145) & (g140)) + ((!g135) & (g146) & (!g137) & (g138) & (!g145) & (!g140)) + ((!g135) & (g146) & (!g137) & (g138) & (g145) & (!g140)) + ((!g135) & (g146) & (g137) & (!g138) & (g145) & (!g140)) + ((!g135) & (g146) & (g137) & (!g138) & (g145) & (g140)) + ((g135) & (!g146) & (!g137) & (!g138) & (!g145) & (g140)) + ((g135) & (!g146) & (!g137) & (!g138) & (g145) & (!g140)) + ((g135) & (!g146) & (!g137) & (g138) & (!g145) & (g140)) + ((g135) & (!g146) & (g137) & (!g138) & (g145) & (!g140)) + ((g135) & (!g146) & (g137) & (!g138) & (g145) & (g140)) + ((g135) & (!g146) & (g137) & (g138) & (g145) & (!g140)) + ((g135) & (!g146) & (g137) & (g138) & (g145) & (g140)) + ((g135) & (g146) & (!g137) & (!g138) & (g145) & (!g140)) + ((g135) & (g146) & (!g137) & (g138) & (!g145) & (g140)) + ((g135) & (g146) & (g137) & (!g138) & (!g145) & (!g140)) + ((g135) & (g146) & (g137) & (!g138) & (g145) & (g140)) + ((g135) & (g146) & (g137) & (g138) & (!g145) & (g140)));
	assign g189 = (((!g185) & (!g186) & (!g187) & (!g188) & (!g139) & (!g136)) + ((!g185) & (!g186) & (!g187) & (!g188) & (!g139) & (g136)) + ((!g185) & (!g186) & (!g187) & (!g188) & (g139) & (!g136)) + ((!g185) & (!g186) & (!g187) & (g188) & (!g139) & (!g136)) + ((!g185) & (!g186) & (!g187) & (g188) & (!g139) & (g136)) + ((!g185) & (!g186) & (!g187) & (g188) & (g139) & (!g136)) + ((!g185) & (!g186) & (!g187) & (g188) & (g139) & (g136)) + ((!g185) & (!g186) & (g187) & (!g188) & (!g139) & (!g136)) + ((!g185) & (!g186) & (g187) & (!g188) & (g139) & (!g136)) + ((!g185) & (!g186) & (g187) & (g188) & (!g139) & (!g136)) + ((!g185) & (!g186) & (g187) & (g188) & (g139) & (!g136)) + ((!g185) & (!g186) & (g187) & (g188) & (g139) & (g136)) + ((!g185) & (g186) & (!g187) & (!g188) & (!g139) & (!g136)) + ((!g185) & (g186) & (!g187) & (!g188) & (!g139) & (g136)) + ((!g185) & (g186) & (!g187) & (g188) & (!g139) & (!g136)) + ((!g185) & (g186) & (!g187) & (g188) & (!g139) & (g136)) + ((!g185) & (g186) & (!g187) & (g188) & (g139) & (g136)) + ((!g185) & (g186) & (g187) & (!g188) & (!g139) & (!g136)) + ((!g185) & (g186) & (g187) & (g188) & (!g139) & (!g136)) + ((!g185) & (g186) & (g187) & (g188) & (g139) & (g136)) + ((g185) & (!g186) & (!g187) & (!g188) & (!g139) & (g136)) + ((g185) & (!g186) & (!g187) & (!g188) & (g139) & (!g136)) + ((g185) & (!g186) & (!g187) & (g188) & (!g139) & (g136)) + ((g185) & (!g186) & (!g187) & (g188) & (g139) & (!g136)) + ((g185) & (!g186) & (!g187) & (g188) & (g139) & (g136)) + ((g185) & (!g186) & (g187) & (!g188) & (g139) & (!g136)) + ((g185) & (!g186) & (g187) & (g188) & (g139) & (!g136)) + ((g185) & (!g186) & (g187) & (g188) & (g139) & (g136)) + ((g185) & (g186) & (!g187) & (!g188) & (!g139) & (g136)) + ((g185) & (g186) & (!g187) & (g188) & (!g139) & (g136)) + ((g185) & (g186) & (!g187) & (g188) & (g139) & (g136)) + ((g185) & (g186) & (g187) & (g188) & (g139) & (g136)));
	assign g191 = (((!sk[42]) & (g189) & (!g190)) + ((!sk[42]) & (g189) & (g190)) + ((sk[42]) & (!g189) & (g190)) + ((sk[42]) & (g189) & (!g190)));
	assign g192 = (((!g139) & (!g136) & (!g137) & (!g138) & (!g145) & (g146)) + ((!g139) & (!g136) & (!g137) & (!g138) & (g145) & (!g146)) + ((!g139) & (!g136) & (!g137) & (g138) & (!g145) & (g146)) + ((!g139) & (!g136) & (!g137) & (g138) & (g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (!g138) & (!g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (!g138) & (g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (g138) & (!g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (g138) & (g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (g138) & (g145) & (g146)) + ((!g139) & (g136) & (!g137) & (!g138) & (g145) & (!g146)) + ((!g139) & (g136) & (!g137) & (g138) & (g145) & (!g146)) + ((!g139) & (g136) & (!g137) & (g138) & (g145) & (g146)) + ((!g139) & (g136) & (g137) & (!g138) & (g145) & (g146)) + ((!g139) & (g136) & (g137) & (g138) & (!g145) & (!g146)) + ((g139) & (!g136) & (!g137) & (!g138) & (!g145) & (g146)) + ((g139) & (!g136) & (!g137) & (g138) & (!g145) & (g146)) + ((g139) & (!g136) & (g137) & (g138) & (g145) & (g146)) + ((g139) & (g136) & (!g137) & (!g138) & (g145) & (g146)) + ((g139) & (g136) & (!g137) & (g138) & (!g145) & (!g146)) + ((g139) & (g136) & (!g137) & (g138) & (g145) & (!g146)) + ((g139) & (g136) & (g137) & (!g138) & (!g145) & (g146)) + ((g139) & (g136) & (g137) & (!g138) & (g145) & (!g146)) + ((g139) & (g136) & (g137) & (!g138) & (g145) & (g146)) + ((g139) & (g136) & (g137) & (g138) & (!g145) & (g146)));
	assign g193 = (((!g139) & (!g136) & (!g137) & (!g138) & (!g145) & (!g146)) + ((!g139) & (!g136) & (!g137) & (!g138) & (!g145) & (g146)) + ((!g139) & (!g136) & (!g137) & (g138) & (!g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (!g138) & (!g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (!g138) & (g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (!g138) & (g145) & (g146)) + ((!g139) & (!g136) & (g137) & (g138) & (!g145) & (g146)) + ((!g139) & (!g136) & (g137) & (g138) & (g145) & (g146)) + ((!g139) & (g136) & (!g137) & (!g138) & (!g145) & (!g146)) + ((!g139) & (g136) & (!g137) & (!g138) & (g145) & (!g146)) + ((!g139) & (g136) & (!g137) & (g138) & (!g145) & (!g146)) + ((!g139) & (g136) & (!g137) & (g138) & (!g145) & (g146)) + ((!g139) & (g136) & (!g137) & (g138) & (g145) & (g146)) + ((!g139) & (g136) & (g137) & (!g138) & (!g145) & (g146)) + ((!g139) & (g136) & (g137) & (g138) & (!g145) & (!g146)) + ((!g139) & (g136) & (g137) & (g138) & (!g145) & (g146)) + ((g139) & (!g136) & (!g137) & (!g138) & (!g145) & (g146)) + ((g139) & (!g136) & (!g137) & (!g138) & (g145) & (g146)) + ((g139) & (!g136) & (!g137) & (g138) & (!g145) & (!g146)) + ((g139) & (!g136) & (!g137) & (g138) & (g145) & (g146)) + ((g139) & (!g136) & (g137) & (!g138) & (!g145) & (!g146)) + ((g139) & (!g136) & (g137) & (!g138) & (g145) & (g146)) + ((g139) & (!g136) & (g137) & (g138) & (g145) & (!g146)) + ((g139) & (g136) & (!g137) & (!g138) & (!g145) & (!g146)) + ((g139) & (g136) & (!g137) & (!g138) & (!g145) & (g146)) + ((g139) & (g136) & (!g137) & (!g138) & (g145) & (g146)) + ((g139) & (g136) & (!g137) & (g138) & (!g145) & (g146)) + ((g139) & (g136) & (!g137) & (g138) & (g145) & (!g146)) + ((g139) & (g136) & (g137) & (!g138) & (g145) & (!g146)) + ((g139) & (g136) & (g137) & (!g138) & (g145) & (g146)));
	assign g194 = (((!g139) & (!g136) & (!g137) & (!g138) & (g145) & (!g146)) + ((!g139) & (!g136) & (!g137) & (g138) & (!g145) & (!g146)) + ((!g139) & (!g136) & (!g137) & (g138) & (g145) & (!g146)) + ((!g139) & (!g136) & (!g137) & (g138) & (g145) & (g146)) + ((!g139) & (!g136) & (g137) & (!g138) & (!g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (!g138) & (!g145) & (g146)) + ((!g139) & (!g136) & (g137) & (!g138) & (g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (g138) & (!g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (g138) & (g145) & (g146)) + ((!g139) & (g136) & (!g137) & (!g138) & (!g145) & (g146)) + ((!g139) & (g136) & (!g137) & (!g138) & (g145) & (!g146)) + ((!g139) & (g136) & (!g137) & (!g138) & (g145) & (g146)) + ((!g139) & (g136) & (g137) & (!g138) & (!g145) & (g146)) + ((!g139) & (g136) & (g137) & (!g138) & (g145) & (!g146)) + ((!g139) & (g136) & (g137) & (!g138) & (g145) & (g146)) + ((!g139) & (g136) & (g137) & (g138) & (!g145) & (!g146)) + ((g139) & (!g136) & (!g137) & (!g138) & (g145) & (!g146)) + ((g139) & (!g136) & (!g137) & (g138) & (!g145) & (!g146)) + ((g139) & (!g136) & (!g137) & (g138) & (g145) & (g146)) + ((g139) & (!g136) & (g137) & (!g138) & (!g145) & (!g146)) + ((g139) & (!g136) & (g137) & (!g138) & (!g145) & (g146)) + ((g139) & (!g136) & (g137) & (g138) & (!g145) & (!g146)) + ((g139) & (!g136) & (g137) & (g138) & (g145) & (!g146)) + ((g139) & (g136) & (!g137) & (!g138) & (g145) & (!g146)) + ((g139) & (g136) & (!g137) & (g138) & (!g145) & (!g146)) + ((g139) & (g136) & (!g137) & (g138) & (g145) & (g146)) + ((g139) & (g136) & (g137) & (!g138) & (!g145) & (!g146)) + ((g139) & (g136) & (g137) & (!g138) & (g145) & (!g146)) + ((g139) & (g136) & (g137) & (!g138) & (g145) & (g146)) + ((g139) & (g136) & (g137) & (g138) & (!g145) & (g146)));
	assign g195 = (((!g139) & (!g136) & (!g137) & (!g138) & (!g145) & (g146)) + ((!g139) & (!g136) & (!g137) & (g138) & (g145) & (!g146)) + ((!g139) & (!g136) & (!g137) & (g138) & (g145) & (g146)) + ((!g139) & (!g136) & (g137) & (!g138) & (!g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (!g138) & (!g145) & (g146)) + ((!g139) & (!g136) & (g137) & (g138) & (g145) & (!g146)) + ((!g139) & (!g136) & (g137) & (g138) & (g145) & (g146)) + ((!g139) & (g136) & (!g137) & (!g138) & (!g145) & (!g146)) + ((!g139) & (g136) & (!g137) & (!g138) & (!g145) & (g146)) + ((!g139) & (g136) & (!g137) & (!g138) & (g145) & (g146)) + ((!g139) & (g136) & (!g137) & (g138) & (!g145) & (g146)) + ((!g139) & (g136) & (g137) & (!g138) & (!g145) & (g146)) + ((!g139) & (g136) & (g137) & (g138) & (!g145) & (!g146)) + ((!g139) & (g136) & (g137) & (g138) & (!g145) & (g146)) + ((!g139) & (g136) & (g137) & (g138) & (g145) & (!g146)) + ((!g139) & (g136) & (g137) & (g138) & (g145) & (g146)) + ((g139) & (!g136) & (!g137) & (g138) & (!g145) & (g146)) + ((g139) & (!g136) & (g137) & (!g138) & (!g145) & (!g146)) + ((g139) & (!g136) & (g137) & (g138) & (!g145) & (!g146)) + ((g139) & (!g136) & (g137) & (g138) & (!g145) & (g146)) + ((g139) & (!g136) & (g137) & (g138) & (g145) & (g146)) + ((g139) & (g136) & (!g137) & (!g138) & (!g145) & (g146)) + ((g139) & (g136) & (!g137) & (!g138) & (g145) & (g146)) + ((g139) & (g136) & (!g137) & (g138) & (!g145) & (!g146)) + ((g139) & (g136) & (!g137) & (g138) & (g145) & (!g146)) + ((g139) & (g136) & (!g137) & (g138) & (g145) & (g146)) + ((g139) & (g136) & (g137) & (!g138) & (g145) & (g146)) + ((g139) & (g136) & (g137) & (g138) & (g145) & (g146)));
	assign g196 = (((!g192) & (!g193) & (!g194) & (!g195) & (!g135) & (g140)) + ((!g192) & (!g193) & (!g194) & (!g195) & (g135) & (!g140)) + ((!g192) & (!g193) & (!g194) & (!g195) & (g135) & (g140)) + ((!g192) & (!g193) & (!g194) & (g195) & (!g135) & (g140)) + ((!g192) & (!g193) & (!g194) & (g195) & (g135) & (!g140)) + ((!g192) & (!g193) & (g194) & (!g195) & (g135) & (!g140)) + ((!g192) & (!g193) & (g194) & (!g195) & (g135) & (g140)) + ((!g192) & (!g193) & (g194) & (g195) & (g135) & (!g140)) + ((!g192) & (g193) & (!g194) & (!g195) & (!g135) & (g140)) + ((!g192) & (g193) & (!g194) & (!g195) & (g135) & (g140)) + ((!g192) & (g193) & (!g194) & (g195) & (!g135) & (g140)) + ((!g192) & (g193) & (g194) & (!g195) & (g135) & (g140)) + ((g192) & (!g193) & (!g194) & (!g195) & (!g135) & (!g140)) + ((g192) & (!g193) & (!g194) & (!g195) & (!g135) & (g140)) + ((g192) & (!g193) & (!g194) & (!g195) & (g135) & (!g140)) + ((g192) & (!g193) & (!g194) & (!g195) & (g135) & (g140)) + ((g192) & (!g193) & (!g194) & (g195) & (!g135) & (!g140)) + ((g192) & (!g193) & (!g194) & (g195) & (!g135) & (g140)) + ((g192) & (!g193) & (!g194) & (g195) & (g135) & (!g140)) + ((g192) & (!g193) & (g194) & (!g195) & (!g135) & (!g140)) + ((g192) & (!g193) & (g194) & (!g195) & (g135) & (!g140)) + ((g192) & (!g193) & (g194) & (!g195) & (g135) & (g140)) + ((g192) & (!g193) & (g194) & (g195) & (!g135) & (!g140)) + ((g192) & (!g193) & (g194) & (g195) & (g135) & (!g140)) + ((g192) & (g193) & (!g194) & (!g195) & (!g135) & (!g140)) + ((g192) & (g193) & (!g194) & (!g195) & (!g135) & (g140)) + ((g192) & (g193) & (!g194) & (!g195) & (g135) & (g140)) + ((g192) & (g193) & (!g194) & (g195) & (!g135) & (!g140)) + ((g192) & (g193) & (!g194) & (g195) & (!g135) & (g140)) + ((g192) & (g193) & (g194) & (!g195) & (!g135) & (!g140)) + ((g192) & (g193) & (g194) & (!g195) & (g135) & (g140)) + ((g192) & (g193) & (g194) & (g195) & (!g135) & (!g140)));
	assign g198 = (((!g196) & (sk[48]) & (g197)) + ((g196) & (!sk[48]) & (!g197)) + ((g196) & (!sk[48]) & (g197)) + ((g196) & (sk[48]) & (!g197)));
	assign g205 = (((!g199) & (!g200) & (!g201) & (!g202) & (g203) & (g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g203) & (!g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g203) & (g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (g203) & (!g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (!g203) & (!g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (!g203) & (g204)) + ((!g199) & (!g200) & (g201) & (g202) & (!g203) & (!g204)) + ((!g199) & (!g200) & (g201) & (g202) & (g203) & (g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (g203) & (!g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (g203) & (g204)) + ((!g199) & (g200) & (!g201) & (g202) & (g203) & (!g204)) + ((!g199) & (g200) & (!g201) & (g202) & (g203) & (g204)) + ((!g199) & (g200) & (g201) & (!g202) & (g203) & (!g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (!g203) & (!g204)) + ((g199) & (!g200) & (g201) & (!g202) & (g203) & (!g204)) + ((g199) & (!g200) & (g201) & (g202) & (!g203) & (g204)) + ((g199) & (!g200) & (g201) & (g202) & (g203) & (g204)) + ((g199) & (g200) & (!g201) & (!g202) & (!g203) & (g204)) + ((g199) & (g200) & (!g201) & (!g202) & (g203) & (!g204)) + ((g199) & (g200) & (g201) & (!g202) & (!g203) & (g204)) + ((g199) & (g200) & (g201) & (!g202) & (g203) & (!g204)) + ((g199) & (g200) & (g201) & (g202) & (!g203) & (!g204)) + ((g199) & (g200) & (g201) & (g202) & (g203) & (!g204)) + ((g199) & (g200) & (g201) & (g202) & (g203) & (g204)));
	assign g206 = (((!g199) & (!g200) & (!g201) & (!g202) & (g203) & (!g204)) + ((!g199) & (!g200) & (!g201) & (!g202) & (g203) & (g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g203) & (!g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g203) & (g204)) + ((!g199) & (!g200) & (g201) & (g202) & (!g203) & (g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (!g203) & (!g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (!g203) & (g204)) + ((!g199) & (g200) & (g201) & (!g202) & (!g203) & (!g204)) + ((!g199) & (g200) & (g201) & (!g202) & (!g203) & (g204)) + ((!g199) & (g200) & (g201) & (!g202) & (g203) & (!g204)) + ((!g199) & (g200) & (g201) & (g202) & (g203) & (g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (!g203) & (g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (g203) & (!g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (g203) & (g204)) + ((g199) & (!g200) & (!g201) & (g202) & (g203) & (!g204)) + ((g199) & (!g200) & (g201) & (!g202) & (!g203) & (!g204)) + ((g199) & (!g200) & (g201) & (!g202) & (g203) & (g204)) + ((g199) & (!g200) & (g201) & (g202) & (!g203) & (g204)) + ((g199) & (!g200) & (g201) & (g202) & (g203) & (g204)) + ((g199) & (g200) & (!g201) & (!g202) & (!g203) & (!g204)) + ((g199) & (g200) & (!g201) & (!g202) & (!g203) & (g204)) + ((g199) & (g200) & (!g201) & (!g202) & (g203) & (!g204)) + ((g199) & (g200) & (!g201) & (!g202) & (g203) & (g204)) + ((g199) & (g200) & (!g201) & (g202) & (!g203) & (!g204)) + ((g199) & (g200) & (!g201) & (g202) & (g203) & (!g204)) + ((g199) & (g200) & (!g201) & (g202) & (g203) & (g204)) + ((g199) & (g200) & (g201) & (!g202) & (g203) & (!g204)) + ((g199) & (g200) & (g201) & (!g202) & (g203) & (g204)) + ((g199) & (g200) & (g201) & (g202) & (!g203) & (g204)) + ((g199) & (g200) & (g201) & (g202) & (g203) & (!g204)));
	assign g207 = (((!g199) & (!g200) & (!g201) & (!g202) & (!g203) & (!g204)) + ((!g199) & (!g200) & (!g201) & (!g202) & (g203) & (g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (g203) & (g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (!g203) & (!g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (!g203) & (g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (g203) & (g204)) + ((!g199) & (!g200) & (g201) & (g202) & (!g203) & (g204)) + ((!g199) & (!g200) & (g201) & (g202) & (g203) & (!g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (!g203) & (!g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (g203) & (!g204)) + ((!g199) & (g200) & (!g201) & (g202) & (g203) & (g204)) + ((!g199) & (g200) & (g201) & (g202) & (!g203) & (!g204)) + ((!g199) & (g200) & (g201) & (g202) & (g203) & (!g204)) + ((g199) & (!g200) & (!g201) & (g202) & (!g203) & (!g204)) + ((g199) & (!g200) & (!g201) & (g202) & (!g203) & (g204)) + ((g199) & (!g200) & (!g201) & (g202) & (g203) & (!g204)) + ((g199) & (!g200) & (g201) & (!g202) & (!g203) & (!g204)) + ((g199) & (!g200) & (g201) & (!g202) & (g203) & (g204)) + ((g199) & (!g200) & (g201) & (g202) & (!g203) & (!g204)) + ((g199) & (!g200) & (g201) & (g202) & (!g203) & (g204)) + ((g199) & (!g200) & (g201) & (g202) & (g203) & (!g204)) + ((g199) & (!g200) & (g201) & (g202) & (g203) & (g204)) + ((g199) & (g200) & (!g201) & (!g202) & (g203) & (g204)) + ((g199) & (g200) & (!g201) & (g202) & (!g203) & (!g204)) + ((g199) & (g200) & (!g201) & (g202) & (g203) & (!g204)) + ((g199) & (g200) & (!g201) & (g202) & (g203) & (g204)) + ((g199) & (g200) & (g201) & (!g202) & (!g203) & (!g204)) + ((g199) & (g200) & (g201) & (g202) & (!g203) & (!g204)) + ((g199) & (g200) & (g201) & (g202) & (!g203) & (g204)) + ((g199) & (g200) & (g201) & (g202) & (g203) & (g204)));
	assign g208 = (((!g199) & (!g200) & (!g201) & (!g202) & (!g203) & (g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (g203) & (!g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (g203) & (g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (!g203) & (g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (g203) & (g204)) + ((!g199) & (!g200) & (g201) & (g202) & (!g203) & (g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (!g203) & (!g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (!g203) & (g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (g203) & (!g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (g203) & (g204)) + ((!g199) & (g200) & (!g201) & (g202) & (g203) & (!g204)) + ((!g199) & (g200) & (!g201) & (g202) & (g203) & (g204)) + ((!g199) & (g200) & (g201) & (g202) & (!g203) & (!g204)) + ((!g199) & (g200) & (g201) & (g202) & (g203) & (!g204)) + ((!g199) & (g200) & (g201) & (g202) & (g203) & (g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (!g203) & (!g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (g203) & (g204)) + ((g199) & (!g200) & (!g201) & (g202) & (g203) & (!g204)) + ((g199) & (!g200) & (!g201) & (g202) & (g203) & (g204)) + ((g199) & (!g200) & (g201) & (!g202) & (!g203) & (g204)) + ((g199) & (!g200) & (g201) & (!g202) & (g203) & (!g204)) + ((g199) & (!g200) & (g201) & (g202) & (g203) & (!g204)) + ((g199) & (g200) & (!g201) & (!g202) & (!g203) & (g204)) + ((g199) & (g200) & (!g201) & (!g202) & (g203) & (g204)) + ((g199) & (g200) & (!g201) & (g202) & (g203) & (!g204)) + ((g199) & (g200) & (!g201) & (g202) & (g203) & (g204)) + ((g199) & (g200) & (g201) & (!g202) & (!g203) & (g204)) + ((g199) & (g200) & (g201) & (g202) & (!g203) & (!g204)));
	assign g211 = (((!g205) & (!g206) & (!g207) & (!g208) & (!g209) & (!g210)) + ((!g205) & (!g206) & (!g207) & (g208) & (!g209) & (!g210)) + ((!g205) & (!g206) & (!g207) & (g208) & (g209) & (g210)) + ((!g205) & (!g206) & (g207) & (!g208) & (!g209) & (!g210)) + ((!g205) & (!g206) & (g207) & (!g208) & (!g209) & (g210)) + ((!g205) & (!g206) & (g207) & (g208) & (!g209) & (!g210)) + ((!g205) & (!g206) & (g207) & (g208) & (!g209) & (g210)) + ((!g205) & (!g206) & (g207) & (g208) & (g209) & (g210)) + ((!g205) & (g206) & (!g207) & (!g208) & (!g209) & (!g210)) + ((!g205) & (g206) & (!g207) & (!g208) & (g209) & (!g210)) + ((!g205) & (g206) & (!g207) & (g208) & (!g209) & (!g210)) + ((!g205) & (g206) & (!g207) & (g208) & (g209) & (!g210)) + ((!g205) & (g206) & (!g207) & (g208) & (g209) & (g210)) + ((!g205) & (g206) & (g207) & (!g208) & (!g209) & (!g210)) + ((!g205) & (g206) & (g207) & (!g208) & (!g209) & (g210)) + ((!g205) & (g206) & (g207) & (!g208) & (g209) & (!g210)) + ((!g205) & (g206) & (g207) & (g208) & (!g209) & (!g210)) + ((!g205) & (g206) & (g207) & (g208) & (!g209) & (g210)) + ((!g205) & (g206) & (g207) & (g208) & (g209) & (!g210)) + ((!g205) & (g206) & (g207) & (g208) & (g209) & (g210)) + ((g205) & (!g206) & (!g207) & (g208) & (g209) & (g210)) + ((g205) & (!g206) & (g207) & (!g208) & (!g209) & (g210)) + ((g205) & (!g206) & (g207) & (g208) & (!g209) & (g210)) + ((g205) & (!g206) & (g207) & (g208) & (g209) & (g210)) + ((g205) & (g206) & (!g207) & (!g208) & (g209) & (!g210)) + ((g205) & (g206) & (!g207) & (g208) & (g209) & (!g210)) + ((g205) & (g206) & (!g207) & (g208) & (g209) & (g210)) + ((g205) & (g206) & (g207) & (!g208) & (!g209) & (g210)) + ((g205) & (g206) & (g207) & (!g208) & (g209) & (!g210)) + ((g205) & (g206) & (g207) & (g208) & (!g209) & (g210)) + ((g205) & (g206) & (g207) & (g208) & (g209) & (!g210)) + ((g205) & (g206) & (g207) & (g208) & (g209) & (g210)));
	assign g213 = (((!sk[54]) & (g211) & (!g212)) + ((!sk[54]) & (g211) & (g212)) + ((sk[54]) & (!g211) & (g212)) + ((sk[54]) & (g211) & (!g212)));
	assign g214 = (((!g199) & (!g200) & (!g201) & (!g202) & (!g209) & (g203)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g209) & (!g203)) + ((!g199) & (!g200) & (!g201) & (g202) & (g209) & (!g203)) + ((!g199) & (!g200) & (g201) & (!g202) & (g209) & (g203)) + ((!g199) & (!g200) & (g201) & (g202) & (!g209) & (g203)) + ((!g199) & (!g200) & (g201) & (g202) & (g209) & (!g203)) + ((!g199) & (g200) & (!g201) & (!g202) & (!g209) & (g203)) + ((!g199) & (g200) & (!g201) & (!g202) & (g209) & (!g203)) + ((!g199) & (g200) & (!g201) & (!g202) & (g209) & (g203)) + ((!g199) & (g200) & (g201) & (!g202) & (g209) & (g203)) + ((!g199) & (g200) & (g201) & (g202) & (g209) & (g203)) + ((g199) & (!g200) & (!g201) & (!g202) & (!g209) & (!g203)) + ((g199) & (!g200) & (!g201) & (!g202) & (g209) & (g203)) + ((g199) & (!g200) & (!g201) & (g202) & (!g209) & (!g203)) + ((g199) & (!g200) & (!g201) & (g202) & (g209) & (!g203)) + ((g199) & (!g200) & (g201) & (!g202) & (g209) & (!g203)) + ((g199) & (!g200) & (g201) & (!g202) & (g209) & (g203)) + ((g199) & (!g200) & (g201) & (g202) & (g209) & (!g203)) + ((g199) & (!g200) & (g201) & (g202) & (g209) & (g203)) + ((g199) & (g200) & (!g201) & (!g202) & (g209) & (!g203)) + ((g199) & (g200) & (!g201) & (!g202) & (g209) & (g203)) + ((g199) & (g200) & (!g201) & (g202) & (g209) & (g203)) + ((g199) & (g200) & (g201) & (!g202) & (!g209) & (!g203)) + ((g199) & (g200) & (g201) & (!g202) & (!g209) & (g203)) + ((g199) & (g200) & (g201) & (!g202) & (g209) & (!g203)) + ((g199) & (g200) & (g201) & (g202) & (!g209) & (g203)) + ((g199) & (g200) & (g201) & (g202) & (g209) & (!g203)));
	assign g215 = (((!g199) & (!g200) & (!g201) & (!g202) & (!g209) & (g203)) + ((!g199) & (!g200) & (!g201) & (!g202) & (g209) & (!g203)) + ((!g199) & (!g200) & (!g201) & (!g202) & (g209) & (g203)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g209) & (!g203)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g209) & (g203)) + ((!g199) & (!g200) & (!g201) & (g202) & (g209) & (g203)) + ((!g199) & (!g200) & (g201) & (!g202) & (g209) & (!g203)) + ((!g199) & (!g200) & (g201) & (g202) & (!g209) & (!g203)) + ((!g199) & (!g200) & (g201) & (g202) & (!g209) & (g203)) + ((!g199) & (!g200) & (g201) & (g202) & (g209) & (g203)) + ((!g199) & (g200) & (!g201) & (!g202) & (g209) & (g203)) + ((!g199) & (g200) & (!g201) & (g202) & (!g209) & (!g203)) + ((!g199) & (g200) & (!g201) & (g202) & (g209) & (!g203)) + ((!g199) & (g200) & (g201) & (!g202) & (g209) & (!g203)) + ((!g199) & (g200) & (g201) & (!g202) & (g209) & (g203)) + ((!g199) & (g200) & (g201) & (g202) & (!g209) & (!g203)) + ((g199) & (!g200) & (!g201) & (!g202) & (!g209) & (!g203)) + ((g199) & (!g200) & (!g201) & (g202) & (!g209) & (!g203)) + ((g199) & (!g200) & (!g201) & (g202) & (!g209) & (g203)) + ((g199) & (!g200) & (g201) & (!g202) & (!g209) & (g203)) + ((g199) & (!g200) & (g201) & (!g202) & (g209) & (g203)) + ((g199) & (!g200) & (g201) & (g202) & (!g209) & (!g203)) + ((g199) & (!g200) & (g201) & (g202) & (!g209) & (g203)) + ((g199) & (g200) & (!g201) & (g202) & (!g209) & (!g203)) + ((g199) & (g200) & (!g201) & (g202) & (g209) & (g203)) + ((g199) & (g200) & (g201) & (!g202) & (!g209) & (!g203)) + ((g199) & (g200) & (g201) & (!g202) & (!g209) & (g203)) + ((g199) & (g200) & (g201) & (!g202) & (g209) & (g203)) + ((g199) & (g200) & (g201) & (g202) & (!g209) & (!g203)) + ((g199) & (g200) & (g201) & (g202) & (!g209) & (g203)) + ((g199) & (g200) & (g201) & (g202) & (g209) & (!g203)));
	assign g216 = (((!g199) & (!g200) & (!g201) & (!g202) & (!g209) & (g203)) + ((!g199) & (!g200) & (!g201) & (g202) & (g209) & (!g203)) + ((!g199) & (!g200) & (g201) & (!g202) & (!g209) & (!g203)) + ((!g199) & (!g200) & (g201) & (!g202) & (g209) & (!g203)) + ((!g199) & (!g200) & (g201) & (g202) & (!g209) & (g203)) + ((!g199) & (!g200) & (g201) & (g202) & (g209) & (!g203)) + ((!g199) & (!g200) & (g201) & (g202) & (g209) & (g203)) + ((!g199) & (g200) & (!g201) & (!g202) & (!g209) & (!g203)) + ((!g199) & (g200) & (!g201) & (!g202) & (g209) & (!g203)) + ((!g199) & (g200) & (!g201) & (g202) & (!g209) & (!g203)) + ((!g199) & (g200) & (!g201) & (g202) & (g209) & (g203)) + ((!g199) & (g200) & (g201) & (!g202) & (g209) & (g203)) + ((!g199) & (g200) & (g201) & (g202) & (!g209) & (g203)) + ((!g199) & (g200) & (g201) & (g202) & (g209) & (!g203)) + ((g199) & (!g200) & (!g201) & (!g202) & (g209) & (g203)) + ((g199) & (!g200) & (!g201) & (g202) & (!g209) & (!g203)) + ((g199) & (!g200) & (!g201) & (g202) & (g209) & (!g203)) + ((g199) & (!g200) & (g201) & (!g202) & (!g209) & (!g203)) + ((g199) & (!g200) & (g201) & (!g202) & (!g209) & (g203)) + ((g199) & (!g200) & (g201) & (!g202) & (g209) & (!g203)) + ((g199) & (!g200) & (g201) & (!g202) & (g209) & (g203)) + ((g199) & (!g200) & (g201) & (g202) & (g209) & (!g203)) + ((g199) & (g200) & (!g201) & (!g202) & (!g209) & (g203)) + ((g199) & (g200) & (!g201) & (!g202) & (g209) & (g203)) + ((g199) & (g200) & (!g201) & (g202) & (!g209) & (g203)) + ((g199) & (g200) & (g201) & (!g202) & (!g209) & (!g203)) + ((g199) & (g200) & (g201) & (!g202) & (!g209) & (g203)) + ((g199) & (g200) & (g201) & (!g202) & (g209) & (g203)) + ((g199) & (g200) & (g201) & (g202) & (!g209) & (!g203)) + ((g199) & (g200) & (g201) & (g202) & (!g209) & (g203)) + ((g199) & (g200) & (g201) & (g202) & (g209) & (!g203)) + ((g199) & (g200) & (g201) & (g202) & (g209) & (g203)));
	assign g217 = (((!g199) & (!g200) & (!g201) & (!g202) & (g209) & (!g203)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g209) & (!g203)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g209) & (g203)) + ((!g199) & (!g200) & (g201) & (!g202) & (g209) & (g203)) + ((!g199) & (!g200) & (g201) & (g202) & (!g209) & (g203)) + ((!g199) & (g200) & (!g201) & (!g202) & (!g209) & (!g203)) + ((!g199) & (g200) & (!g201) & (!g202) & (g209) & (!g203)) + ((!g199) & (g200) & (!g201) & (g202) & (!g209) & (g203)) + ((!g199) & (g200) & (g201) & (!g202) & (!g209) & (g203)) + ((!g199) & (g200) & (g201) & (!g202) & (g209) & (!g203)) + ((!g199) & (g200) & (g201) & (!g202) & (g209) & (g203)) + ((!g199) & (g200) & (g201) & (g202) & (g209) & (!g203)) + ((!g199) & (g200) & (g201) & (g202) & (g209) & (g203)) + ((g199) & (!g200) & (!g201) & (!g202) & (!g209) & (!g203)) + ((g199) & (!g200) & (!g201) & (g202) & (!g209) & (!g203)) + ((g199) & (!g200) & (!g201) & (g202) & (!g209) & (g203)) + ((g199) & (!g200) & (!g201) & (g202) & (g209) & (!g203)) + ((g199) & (!g200) & (g201) & (!g202) & (!g209) & (!g203)) + ((g199) & (!g200) & (g201) & (!g202) & (g209) & (g203)) + ((g199) & (!g200) & (g201) & (g202) & (g209) & (!g203)) + ((g199) & (g200) & (!g201) & (!g202) & (!g209) & (!g203)) + ((g199) & (g200) & (!g201) & (g202) & (!g209) & (!g203)) + ((g199) & (g200) & (!g201) & (g202) & (g209) & (!g203)) + ((g199) & (g200) & (!g201) & (g202) & (g209) & (g203)) + ((g199) & (g200) & (g201) & (g202) & (!g209) & (g203)) + ((g199) & (g200) & (g201) & (g202) & (g209) & (g203)));
	assign g218 = (((!g214) & (!g215) & (!g216) & (!g217) & (!g204) & (!g210)) + ((!g214) & (!g215) & (!g216) & (!g217) & (g204) & (!g210)) + ((!g214) & (!g215) & (!g216) & (g217) & (!g204) & (!g210)) + ((!g214) & (!g215) & (!g216) & (g217) & (g204) & (!g210)) + ((!g214) & (!g215) & (!g216) & (g217) & (g204) & (g210)) + ((!g214) & (!g215) & (g216) & (!g217) & (!g204) & (!g210)) + ((!g214) & (!g215) & (g216) & (!g217) & (!g204) & (g210)) + ((!g214) & (!g215) & (g216) & (!g217) & (g204) & (!g210)) + ((!g214) & (!g215) & (g216) & (g217) & (!g204) & (!g210)) + ((!g214) & (!g215) & (g216) & (g217) & (!g204) & (g210)) + ((!g214) & (!g215) & (g216) & (g217) & (g204) & (!g210)) + ((!g214) & (!g215) & (g216) & (g217) & (g204) & (g210)) + ((!g214) & (g215) & (!g216) & (!g217) & (!g204) & (!g210)) + ((!g214) & (g215) & (!g216) & (g217) & (!g204) & (!g210)) + ((!g214) & (g215) & (!g216) & (g217) & (g204) & (g210)) + ((!g214) & (g215) & (g216) & (!g217) & (!g204) & (!g210)) + ((!g214) & (g215) & (g216) & (!g217) & (!g204) & (g210)) + ((!g214) & (g215) & (g216) & (g217) & (!g204) & (!g210)) + ((!g214) & (g215) & (g216) & (g217) & (!g204) & (g210)) + ((!g214) & (g215) & (g216) & (g217) & (g204) & (g210)) + ((g214) & (!g215) & (!g216) & (!g217) & (g204) & (!g210)) + ((g214) & (!g215) & (!g216) & (g217) & (g204) & (!g210)) + ((g214) & (!g215) & (!g216) & (g217) & (g204) & (g210)) + ((g214) & (!g215) & (g216) & (!g217) & (!g204) & (g210)) + ((g214) & (!g215) & (g216) & (!g217) & (g204) & (!g210)) + ((g214) & (!g215) & (g216) & (g217) & (!g204) & (g210)) + ((g214) & (!g215) & (g216) & (g217) & (g204) & (!g210)) + ((g214) & (!g215) & (g216) & (g217) & (g204) & (g210)) + ((g214) & (g215) & (!g216) & (g217) & (g204) & (g210)) + ((g214) & (g215) & (g216) & (!g217) & (!g204) & (g210)) + ((g214) & (g215) & (g216) & (g217) & (!g204) & (g210)) + ((g214) & (g215) & (g216) & (g217) & (g204) & (g210)));
	assign g220 = (((!sk[60]) & (g218) & (!g219)) + ((!sk[60]) & (g218) & (g219)) + ((sk[60]) & (!g218) & (g219)) + ((sk[60]) & (g218) & (!g219)));
	assign g221 = (((!g203) & (!g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((!g203) & (!g200) & (!g201) & (!g202) & (g209) & (g204)) + ((!g203) & (!g200) & (!g201) & (g202) & (!g209) & (g204)) + ((!g203) & (!g200) & (!g201) & (g202) & (g209) & (!g204)) + ((!g203) & (!g200) & (!g201) & (g202) & (g209) & (g204)) + ((!g203) & (!g200) & (g201) & (!g202) & (!g209) & (g204)) + ((!g203) & (!g200) & (g201) & (g202) & (!g209) & (!g204)) + ((!g203) & (!g200) & (g201) & (g202) & (g209) & (!g204)) + ((!g203) & (g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((!g203) & (g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((!g203) & (g200) & (!g201) & (g202) & (!g209) & (g204)) + ((!g203) & (g200) & (g201) & (!g202) & (!g209) & (!g204)) + ((!g203) & (g200) & (g201) & (!g202) & (!g209) & (g204)) + ((!g203) & (g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g203) & (g200) & (g201) & (!g202) & (g209) & (g204)) + ((g203) & (!g200) & (!g201) & (g202) & (!g209) & (g204)) + ((g203) & (!g200) & (!g201) & (g202) & (g209) & (g204)) + ((g203) & (g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((g203) & (g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((g203) & (g200) & (!g201) & (g202) & (g209) & (!g204)) + ((g203) & (g200) & (g201) & (g202) & (!g209) & (!g204)) + ((g203) & (g200) & (g201) & (g202) & (!g209) & (g204)));
	assign g222 = (((!g203) & (!g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((!g203) & (!g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((!g203) & (!g200) & (!g201) & (g202) & (g209) & (g204)) + ((!g203) & (!g200) & (g201) & (!g202) & (!g209) & (!g204)) + ((!g203) & (!g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g203) & (!g200) & (g201) & (g202) & (!g209) & (g204)) + ((!g203) & (g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((!g203) & (g200) & (!g201) & (!g202) & (g209) & (g204)) + ((!g203) & (g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((!g203) & (g200) & (!g201) & (g202) & (!g209) & (g204)) + ((!g203) & (g200) & (!g201) & (g202) & (g209) & (g204)) + ((!g203) & (g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g203) & (g200) & (g201) & (!g202) & (g209) & (g204)) + ((!g203) & (g200) & (g201) & (g202) & (g209) & (!g204)) + ((g203) & (!g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((g203) & (!g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((g203) & (!g200) & (!g201) & (!g202) & (g209) & (g204)) + ((g203) & (!g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((g203) & (!g200) & (!g201) & (g202) & (!g209) & (g204)) + ((g203) & (!g200) & (!g201) & (g202) & (g209) & (!g204)) + ((g203) & (!g200) & (g201) & (g202) & (!g209) & (!g204)) + ((g203) & (g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((g203) & (g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((g203) & (g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((g203) & (g200) & (!g201) & (g202) & (g209) & (!g204)) + ((g203) & (g200) & (!g201) & (g202) & (g209) & (g204)) + ((g203) & (g200) & (g201) & (!g202) & (!g209) & (!g204)) + ((g203) & (g200) & (g201) & (!g202) & (g209) & (!g204)) + ((g203) & (g200) & (g201) & (g202) & (!g209) & (g204)) + ((g203) & (g200) & (g201) & (g202) & (g209) & (g204)));
	assign g223 = (((!g203) & (!g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((!g203) & (!g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((!g203) & (!g200) & (!g201) & (g202) & (!g209) & (g204)) + ((!g203) & (!g200) & (g201) & (!g202) & (!g209) & (g204)) + ((!g203) & (!g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g203) & (!g200) & (g201) & (g202) & (!g209) & (g204)) + ((!g203) & (g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((!g203) & (g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((!g203) & (g200) & (!g201) & (g202) & (g209) & (!g204)) + ((!g203) & (g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g203) & (g200) & (g201) & (g202) & (!g209) & (!g204)) + ((!g203) & (g200) & (g201) & (g202) & (g209) & (!g204)) + ((g203) & (!g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((g203) & (!g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((g203) & (!g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((g203) & (!g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((g203) & (!g200) & (!g201) & (g202) & (!g209) & (g204)) + ((g203) & (!g200) & (!g201) & (g202) & (g209) & (!g204)) + ((g203) & (!g200) & (!g201) & (g202) & (g209) & (g204)) + ((g203) & (!g200) & (g201) & (!g202) & (!g209) & (g204)) + ((g203) & (!g200) & (g201) & (!g202) & (g209) & (!g204)) + ((g203) & (!g200) & (g201) & (g202) & (!g209) & (!g204)) + ((g203) & (!g200) & (g201) & (g202) & (g209) & (g204)) + ((g203) & (g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((g203) & (g200) & (!g201) & (!g202) & (g209) & (g204)) + ((g203) & (g200) & (g201) & (!g202) & (g209) & (g204)) + ((g203) & (g200) & (g201) & (g202) & (!g209) & (!g204)) + ((g203) & (g200) & (g201) & (g202) & (!g209) & (g204)) + ((g203) & (g200) & (g201) & (g202) & (g209) & (g204)));
	assign g224 = (((!g203) & (!g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((!g203) & (!g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((!g203) & (!g200) & (!g201) & (!g202) & (g209) & (g204)) + ((!g203) & (!g200) & (!g201) & (g202) & (!g209) & (g204)) + ((!g203) & (!g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g203) & (!g200) & (g201) & (g202) & (g209) & (g204)) + ((!g203) & (g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((!g203) & (g200) & (!g201) & (g202) & (!g209) & (g204)) + ((!g203) & (g200) & (!g201) & (g202) & (g209) & (g204)) + ((!g203) & (g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g203) & (g200) & (g201) & (!g202) & (g209) & (g204)) + ((!g203) & (g200) & (g201) & (g202) & (!g209) & (!g204)) + ((!g203) & (g200) & (g201) & (g202) & (!g209) & (g204)) + ((!g203) & (g200) & (g201) & (g202) & (g209) & (!g204)) + ((!g203) & (g200) & (g201) & (g202) & (g209) & (g204)) + ((g203) & (!g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((g203) & (!g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((g203) & (!g200) & (!g201) & (!g202) & (g209) & (g204)) + ((g203) & (!g200) & (!g201) & (g202) & (g209) & (g204)) + ((g203) & (!g200) & (g201) & (!g202) & (!g209) & (g204)) + ((g203) & (!g200) & (g201) & (!g202) & (g209) & (!g204)) + ((g203) & (!g200) & (g201) & (g202) & (g209) & (!g204)) + ((g203) & (g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((g203) & (g200) & (!g201) & (g202) & (!g209) & (g204)) + ((g203) & (g200) & (!g201) & (g202) & (g209) & (!g204)) + ((g203) & (g200) & (g201) & (!g202) & (g209) & (g204)) + ((g203) & (g200) & (g201) & (g202) & (!g209) & (!g204)));
	assign g225 = (((!g221) & (!g222) & (!g223) & (!g224) & (!g199) & (g210)) + ((!g221) & (!g222) & (!g223) & (!g224) & (g199) & (!g210)) + ((!g221) & (!g222) & (!g223) & (!g224) & (g199) & (g210)) + ((!g221) & (!g222) & (!g223) & (g224) & (!g199) & (g210)) + ((!g221) & (!g222) & (!g223) & (g224) & (g199) & (!g210)) + ((!g221) & (!g222) & (g223) & (!g224) & (g199) & (!g210)) + ((!g221) & (!g222) & (g223) & (!g224) & (g199) & (g210)) + ((!g221) & (!g222) & (g223) & (g224) & (g199) & (!g210)) + ((!g221) & (g222) & (!g223) & (!g224) & (!g199) & (g210)) + ((!g221) & (g222) & (!g223) & (!g224) & (g199) & (g210)) + ((!g221) & (g222) & (!g223) & (g224) & (!g199) & (g210)) + ((!g221) & (g222) & (g223) & (!g224) & (g199) & (g210)) + ((g221) & (!g222) & (!g223) & (!g224) & (!g199) & (!g210)) + ((g221) & (!g222) & (!g223) & (!g224) & (!g199) & (g210)) + ((g221) & (!g222) & (!g223) & (!g224) & (g199) & (!g210)) + ((g221) & (!g222) & (!g223) & (!g224) & (g199) & (g210)) + ((g221) & (!g222) & (!g223) & (g224) & (!g199) & (!g210)) + ((g221) & (!g222) & (!g223) & (g224) & (!g199) & (g210)) + ((g221) & (!g222) & (!g223) & (g224) & (g199) & (!g210)) + ((g221) & (!g222) & (g223) & (!g224) & (!g199) & (!g210)) + ((g221) & (!g222) & (g223) & (!g224) & (g199) & (!g210)) + ((g221) & (!g222) & (g223) & (!g224) & (g199) & (g210)) + ((g221) & (!g222) & (g223) & (g224) & (!g199) & (!g210)) + ((g221) & (!g222) & (g223) & (g224) & (g199) & (!g210)) + ((g221) & (g222) & (!g223) & (!g224) & (!g199) & (!g210)) + ((g221) & (g222) & (!g223) & (!g224) & (!g199) & (g210)) + ((g221) & (g222) & (!g223) & (!g224) & (g199) & (g210)) + ((g221) & (g222) & (!g223) & (g224) & (!g199) & (!g210)) + ((g221) & (g222) & (!g223) & (g224) & (!g199) & (g210)) + ((g221) & (g222) & (g223) & (!g224) & (!g199) & (!g210)) + ((g221) & (g222) & (g223) & (!g224) & (g199) & (g210)) + ((g221) & (g222) & (g223) & (g224) & (!g199) & (!g210)));
	assign g227 = (((!g225) & (sk[66]) & (g226)) + ((g225) & (!sk[66]) & (!g226)) + ((g225) & (!sk[66]) & (g226)) + ((g225) & (sk[66]) & (!g226)));
	assign g228 = (((!g199) & (!g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (g209) & (g204)) + ((!g199) & (!g200) & (g201) & (g202) & (!g209) & (!g204)) + ((!g199) & (!g200) & (g201) & (g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (g201) & (g202) & (g209) & (g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (g200) & (g201) & (!g202) & (!g209) & (!g204)) + ((!g199) & (g200) & (g201) & (g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((g199) & (!g200) & (g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (g201) & (!g202) & (!g209) & (g204)) + ((g199) & (!g200) & (g201) & (!g202) & (g209) & (!g204)) + ((g199) & (!g200) & (g201) & (g202) & (!g209) & (g204)) + ((g199) & (g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((g199) & (g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((g199) & (g200) & (!g201) & (g202) & (g209) & (!g204)) + ((g199) & (g200) & (g201) & (!g202) & (!g209) & (g204)) + ((g199) & (g200) & (g201) & (!g202) & (g209) & (g204)));
	assign g229 = (((!g199) & (!g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (!g201) & (!g202) & (g209) & (g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (g201) & (g202) & (!g209) & (!g204)) + ((!g199) & (!g200) & (g201) & (g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (g201) & (g202) & (g209) & (g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (g209) & (g204)) + ((!g199) & (g200) & (!g201) & (g202) & (g209) & (g204)) + ((!g199) & (g200) & (g201) & (!g202) & (!g209) & (!g204)) + ((!g199) & (g200) & (g201) & (!g202) & (!g209) & (g204)) + ((!g199) & (g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (g200) & (g201) & (g202) & (!g209) & (g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((g199) & (!g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (!g201) & (g202) & (!g209) & (g204)) + ((g199) & (!g200) & (!g201) & (g202) & (g209) & (g204)) + ((g199) & (!g200) & (g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (g201) & (!g202) & (!g209) & (g204)) + ((g199) & (!g200) & (g201) & (!g202) & (g209) & (g204)) + ((g199) & (!g200) & (g201) & (g202) & (!g209) & (g204)) + ((g199) & (g200) & (!g201) & (g202) & (!g209) & (g204)) + ((g199) & (g200) & (!g201) & (g202) & (g209) & (!g204)) + ((g199) & (g200) & (g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (g200) & (g201) & (g202) & (!g209) & (!g204)));
	assign g230 = (((!g199) & (!g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (!g201) & (!g202) & (g209) & (g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (g201) & (!g202) & (g209) & (g204)) + ((!g199) & (!g200) & (g201) & (g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (g201) & (g202) & (g209) & (g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (g209) & (g204)) + ((!g199) & (g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((!g199) & (g200) & (!g201) & (g202) & (!g209) & (g204)) + ((!g199) & (g200) & (g201) & (!g202) & (!g209) & (g204)) + ((!g199) & (g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (g200) & (g201) & (g202) & (g209) & (g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (g209) & (g204)) + ((g199) & (!g200) & (!g201) & (g202) & (g209) & (g204)) + ((g199) & (!g200) & (g201) & (g202) & (!g209) & (!g204)) + ((g199) & (g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((g199) & (g200) & (!g201) & (g202) & (g209) & (g204)) + ((g199) & (g200) & (g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (g200) & (g201) & (!g202) & (!g209) & (g204)) + ((g199) & (g200) & (g201) & (!g202) & (g209) & (g204)) + ((g199) & (g200) & (g201) & (g202) & (!g209) & (!g204)) + ((g199) & (g200) & (g201) & (g202) & (g209) & (g204)));
	assign g231 = (((!g199) & (!g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (!g201) & (g202) & (g209) & (g204)) + ((!g199) & (!g200) & (g201) & (g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (g201) & (g202) & (g209) & (g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (!g209) & (!g204)) + ((!g199) & (g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (g200) & (!g201) & (g202) & (!g209) & (!g204)) + ((!g199) & (g200) & (!g201) & (g202) & (!g209) & (g204)) + ((!g199) & (g200) & (!g201) & (g202) & (g209) & (!g204)) + ((!g199) & (g200) & (g201) & (!g202) & (!g209) & (!g204)) + ((!g199) & (g200) & (g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (g200) & (g201) & (!g202) & (g209) & (g204)) + ((g199) & (!g200) & (!g201) & (!g202) & (g209) & (g204)) + ((g199) & (!g200) & (!g201) & (g202) & (g209) & (!g204)) + ((g199) & (!g200) & (g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (g201) & (!g202) & (g209) & (!g204)) + ((g199) & (!g200) & (g201) & (!g202) & (g209) & (g204)) + ((g199) & (!g200) & (g201) & (g202) & (!g209) & (g204)) + ((g199) & (!g200) & (g201) & (g202) & (g209) & (!g204)) + ((g199) & (!g200) & (g201) & (g202) & (g209) & (g204)) + ((g199) & (g200) & (!g201) & (!g202) & (!g209) & (g204)) + ((g199) & (g200) & (!g201) & (!g202) & (g209) & (!g204)) + ((g199) & (g200) & (g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (g200) & (g201) & (!g202) & (!g209) & (g204)) + ((g199) & (g200) & (g201) & (g202) & (g209) & (g204)));
	assign g232 = (((!g228) & (!g229) & (!g230) & (!g231) & (!g210) & (g203)) + ((!g228) & (!g229) & (!g230) & (!g231) & (g210) & (!g203)) + ((!g228) & (!g229) & (!g230) & (!g231) & (g210) & (g203)) + ((!g228) & (!g229) & (!g230) & (g231) & (!g210) & (g203)) + ((!g228) & (!g229) & (!g230) & (g231) & (g210) & (!g203)) + ((!g228) & (!g229) & (g230) & (!g231) & (g210) & (!g203)) + ((!g228) & (!g229) & (g230) & (!g231) & (g210) & (g203)) + ((!g228) & (!g229) & (g230) & (g231) & (g210) & (!g203)) + ((!g228) & (g229) & (!g230) & (!g231) & (!g210) & (g203)) + ((!g228) & (g229) & (!g230) & (!g231) & (g210) & (g203)) + ((!g228) & (g229) & (!g230) & (g231) & (!g210) & (g203)) + ((!g228) & (g229) & (g230) & (!g231) & (g210) & (g203)) + ((g228) & (!g229) & (!g230) & (!g231) & (!g210) & (!g203)) + ((g228) & (!g229) & (!g230) & (!g231) & (!g210) & (g203)) + ((g228) & (!g229) & (!g230) & (!g231) & (g210) & (!g203)) + ((g228) & (!g229) & (!g230) & (!g231) & (g210) & (g203)) + ((g228) & (!g229) & (!g230) & (g231) & (!g210) & (!g203)) + ((g228) & (!g229) & (!g230) & (g231) & (!g210) & (g203)) + ((g228) & (!g229) & (!g230) & (g231) & (g210) & (!g203)) + ((g228) & (!g229) & (g230) & (!g231) & (!g210) & (!g203)) + ((g228) & (!g229) & (g230) & (!g231) & (g210) & (!g203)) + ((g228) & (!g229) & (g230) & (!g231) & (g210) & (g203)) + ((g228) & (!g229) & (g230) & (g231) & (!g210) & (!g203)) + ((g228) & (!g229) & (g230) & (g231) & (g210) & (!g203)) + ((g228) & (g229) & (!g230) & (!g231) & (!g210) & (!g203)) + ((g228) & (g229) & (!g230) & (!g231) & (!g210) & (g203)) + ((g228) & (g229) & (!g230) & (!g231) & (g210) & (g203)) + ((g228) & (g229) & (!g230) & (g231) & (!g210) & (!g203)) + ((g228) & (g229) & (!g230) & (g231) & (!g210) & (g203)) + ((g228) & (g229) & (g230) & (!g231) & (!g210) & (!g203)) + ((g228) & (g229) & (g230) & (!g231) & (g210) & (g203)) + ((g228) & (g229) & (g230) & (g231) & (!g210) & (!g203)));
	assign g234 = (((!g232) & (sk[72]) & (g233)) + ((g232) & (!sk[72]) & (!g233)) + ((g232) & (!sk[72]) & (g233)) + ((g232) & (sk[72]) & (!g233)));
	assign g235 = (((!g199) & (!g200) & (!g203) & (!g210) & (!g209) & (g204)) + ((!g199) & (!g200) & (g203) & (!g210) & (!g209) & (g204)) + ((!g199) & (!g200) & (g203) & (!g210) & (g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (!g210) & (g209) & (g204)) + ((!g199) & (!g200) & (g203) & (g210) & (!g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (g210) & (g209) & (!g204)) + ((!g199) & (g200) & (!g203) & (!g210) & (!g209) & (!g204)) + ((!g199) & (g200) & (!g203) & (!g210) & (!g209) & (g204)) + ((!g199) & (g200) & (!g203) & (g210) & (!g209) & (!g204)) + ((!g199) & (g200) & (!g203) & (g210) & (!g209) & (g204)) + ((!g199) & (g200) & (!g203) & (g210) & (g209) & (g204)) + ((!g199) & (g200) & (g203) & (g210) & (!g209) & (g204)) + ((!g199) & (g200) & (g203) & (g210) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g210) & (!g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g210) & (!g209) & (g204)) + ((g199) & (!g200) & (!g203) & (g210) & (!g209) & (g204)) + ((g199) & (!g200) & (g203) & (!g210) & (g209) & (!g204)) + ((g199) & (!g200) & (g203) & (g210) & (!g209) & (!g204)) + ((g199) & (!g200) & (g203) & (g210) & (!g209) & (g204)) + ((g199) & (!g200) & (g203) & (g210) & (g209) & (!g204)) + ((g199) & (g200) & (!g203) & (!g210) & (!g209) & (!g204)) + ((g199) & (g200) & (!g203) & (!g210) & (g209) & (!g204)) + ((g199) & (g200) & (!g203) & (g210) & (g209) & (!g204)) + ((g199) & (g200) & (g203) & (!g210) & (!g209) & (!g204)) + ((g199) & (g200) & (g203) & (!g210) & (!g209) & (g204)) + ((g199) & (g200) & (g203) & (g210) & (!g209) & (g204)));
	assign g236 = (((!g199) & (!g200) & (!g203) & (!g210) & (!g209) & (!g204)) + ((!g199) & (!g200) & (!g203) & (!g210) & (!g209) & (g204)) + ((!g199) & (!g200) & (!g203) & (!g210) & (g209) & (!g204)) + ((!g199) & (!g200) & (!g203) & (!g210) & (g209) & (g204)) + ((!g199) & (!g200) & (!g203) & (g210) & (!g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (!g210) & (!g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (!g210) & (g209) & (g204)) + ((!g199) & (!g200) & (g203) & (g210) & (!g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (g210) & (g209) & (g204)) + ((!g199) & (g200) & (!g203) & (!g210) & (!g209) & (g204)) + ((!g199) & (g200) & (!g203) & (g210) & (g209) & (!g204)) + ((!g199) & (g200) & (g203) & (!g210) & (!g209) & (!g204)) + ((!g199) & (g200) & (g203) & (!g210) & (!g209) & (g204)) + ((!g199) & (g200) & (g203) & (!g210) & (g209) & (!g204)) + ((!g199) & (g200) & (g203) & (!g210) & (g209) & (g204)) + ((!g199) & (g200) & (g203) & (g210) & (!g209) & (!g204)) + ((!g199) & (g200) & (g203) & (g210) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g210) & (!g209) & (g204)) + ((g199) & (!g200) & (!g203) & (!g210) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g210) & (g209) & (g204)) + ((g199) & (!g200) & (!g203) & (g210) & (!g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (g210) & (g209) & (g204)) + ((g199) & (!g200) & (g203) & (!g210) & (g209) & (!g204)) + ((g199) & (!g200) & (g203) & (!g210) & (g209) & (g204)) + ((g199) & (!g200) & (g203) & (g210) & (!g209) & (g204)) + ((g199) & (g200) & (!g203) & (!g210) & (g209) & (!g204)) + ((g199) & (g200) & (!g203) & (!g210) & (g209) & (g204)) + ((g199) & (g200) & (!g203) & (g210) & (!g209) & (!g204)) + ((g199) & (g200) & (!g203) & (g210) & (!g209) & (g204)) + ((g199) & (g200) & (g203) & (!g210) & (g209) & (!g204)) + ((g199) & (g200) & (g203) & (!g210) & (g209) & (g204)) + ((g199) & (g200) & (g203) & (g210) & (!g209) & (g204)));
	assign g237 = (((!g199) & (!g200) & (!g203) & (!g210) & (!g209) & (!g204)) + ((!g199) & (!g200) & (!g203) & (!g210) & (!g209) & (g204)) + ((!g199) & (!g200) & (g203) & (!g210) & (!g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (!g210) & (g209) & (g204)) + ((!g199) & (!g200) & (g203) & (g210) & (!g209) & (g204)) + ((!g199) & (g200) & (!g203) & (g210) & (!g209) & (!g204)) + ((!g199) & (g200) & (!g203) & (g210) & (g209) & (!g204)) + ((!g199) & (g200) & (!g203) & (g210) & (g209) & (g204)) + ((!g199) & (g200) & (g203) & (!g210) & (!g209) & (!g204)) + ((!g199) & (g200) & (g203) & (!g210) & (g209) & (!g204)) + ((!g199) & (g200) & (g203) & (!g210) & (g209) & (g204)) + ((!g199) & (g200) & (g203) & (g210) & (!g209) & (!g204)) + ((!g199) & (g200) & (g203) & (g210) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g210) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g210) & (g209) & (g204)) + ((g199) & (!g200) & (!g203) & (g210) & (!g209) & (g204)) + ((g199) & (!g200) & (!g203) & (g210) & (g209) & (g204)) + ((g199) & (!g200) & (g203) & (!g210) & (!g209) & (!g204)) + ((g199) & (!g200) & (g203) & (!g210) & (!g209) & (g204)) + ((g199) & (!g200) & (g203) & (!g210) & (g209) & (g204)) + ((g199) & (!g200) & (g203) & (g210) & (!g209) & (!g204)) + ((g199) & (!g200) & (g203) & (g210) & (!g209) & (g204)) + ((g199) & (!g200) & (g203) & (g210) & (g209) & (!g204)) + ((g199) & (!g200) & (g203) & (g210) & (g209) & (g204)) + ((g199) & (g200) & (!g203) & (!g210) & (!g209) & (g204)) + ((g199) & (g200) & (!g203) & (g210) & (!g209) & (!g204)) + ((g199) & (g200) & (!g203) & (g210) & (g209) & (!g204)) + ((g199) & (g200) & (g203) & (!g210) & (!g209) & (!g204)) + ((g199) & (g200) & (g203) & (!g210) & (!g209) & (g204)) + ((g199) & (g200) & (g203) & (!g210) & (g209) & (!g204)) + ((g199) & (g200) & (g203) & (g210) & (!g209) & (!g204)) + ((g199) & (g200) & (g203) & (g210) & (g209) & (!g204)));
	assign g238 = (((!g199) & (!g200) & (!g203) & (!g210) & (g209) & (g204)) + ((!g199) & (!g200) & (!g203) & (g210) & (!g209) & (!g204)) + ((!g199) & (!g200) & (!g203) & (g210) & (g209) & (g204)) + ((!g199) & (!g200) & (g203) & (!g210) & (!g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (!g210) & (g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (g210) & (!g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (g210) & (!g209) & (g204)) + ((!g199) & (!g200) & (g203) & (g210) & (g209) & (!g204)) + ((!g199) & (g200) & (!g203) & (!g210) & (!g209) & (!g204)) + ((!g199) & (g200) & (!g203) & (g210) & (!g209) & (g204)) + ((!g199) & (g200) & (!g203) & (g210) & (g209) & (!g204)) + ((!g199) & (g200) & (!g203) & (g210) & (g209) & (g204)) + ((!g199) & (g200) & (g203) & (!g210) & (!g209) & (!g204)) + ((!g199) & (g200) & (g203) & (g210) & (!g209) & (!g204)) + ((!g199) & (g200) & (g203) & (g210) & (!g209) & (g204)) + ((g199) & (!g200) & (!g203) & (!g210) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g210) & (g209) & (g204)) + ((g199) & (!g200) & (g203) & (!g210) & (!g209) & (!g204)) + ((g199) & (!g200) & (g203) & (!g210) & (g209) & (!g204)) + ((g199) & (!g200) & (g203) & (g210) & (g209) & (!g204)) + ((g199) & (g200) & (!g203) & (!g210) & (g209) & (!g204)) + ((g199) & (g200) & (!g203) & (g210) & (g209) & (g204)) + ((g199) & (g200) & (g203) & (!g210) & (!g209) & (!g204)) + ((g199) & (g200) & (g203) & (!g210) & (!g209) & (g204)) + ((g199) & (g200) & (g203) & (!g210) & (g209) & (!g204)) + ((g199) & (g200) & (g203) & (g210) & (!g209) & (!g204)));
	assign g239 = (((!g235) & (!g236) & (!g237) & (!g238) & (g201) & (g202)) + ((!g235) & (!g236) & (g237) & (!g238) & (!g201) & (g202)) + ((!g235) & (!g236) & (g237) & (!g238) & (g201) & (g202)) + ((!g235) & (!g236) & (g237) & (g238) & (!g201) & (g202)) + ((!g235) & (g236) & (!g237) & (!g238) & (g201) & (!g202)) + ((!g235) & (g236) & (!g237) & (!g238) & (g201) & (g202)) + ((!g235) & (g236) & (!g237) & (g238) & (g201) & (!g202)) + ((!g235) & (g236) & (g237) & (!g238) & (!g201) & (g202)) + ((!g235) & (g236) & (g237) & (!g238) & (g201) & (!g202)) + ((!g235) & (g236) & (g237) & (!g238) & (g201) & (g202)) + ((!g235) & (g236) & (g237) & (g238) & (!g201) & (g202)) + ((!g235) & (g236) & (g237) & (g238) & (g201) & (!g202)) + ((g235) & (!g236) & (!g237) & (!g238) & (!g201) & (!g202)) + ((g235) & (!g236) & (!g237) & (!g238) & (g201) & (g202)) + ((g235) & (!g236) & (!g237) & (g238) & (!g201) & (!g202)) + ((g235) & (!g236) & (g237) & (!g238) & (!g201) & (!g202)) + ((g235) & (!g236) & (g237) & (!g238) & (!g201) & (g202)) + ((g235) & (!g236) & (g237) & (!g238) & (g201) & (g202)) + ((g235) & (!g236) & (g237) & (g238) & (!g201) & (!g202)) + ((g235) & (!g236) & (g237) & (g238) & (!g201) & (g202)) + ((g235) & (g236) & (!g237) & (!g238) & (!g201) & (!g202)) + ((g235) & (g236) & (!g237) & (!g238) & (g201) & (!g202)) + ((g235) & (g236) & (!g237) & (!g238) & (g201) & (g202)) + ((g235) & (g236) & (!g237) & (g238) & (!g201) & (!g202)) + ((g235) & (g236) & (!g237) & (g238) & (g201) & (!g202)) + ((g235) & (g236) & (g237) & (!g238) & (!g201) & (!g202)) + ((g235) & (g236) & (g237) & (!g238) & (!g201) & (g202)) + ((g235) & (g236) & (g237) & (!g238) & (g201) & (!g202)) + ((g235) & (g236) & (g237) & (!g238) & (g201) & (g202)) + ((g235) & (g236) & (g237) & (g238) & (!g201) & (!g202)) + ((g235) & (g236) & (g237) & (g238) & (!g201) & (g202)) + ((g235) & (g236) & (g237) & (g238) & (g201) & (!g202)));
	assign g241 = (((!sk[78]) & (g239) & (!g240)) + ((!sk[78]) & (g239) & (g240)) + ((sk[78]) & (!g239) & (g240)) + ((sk[78]) & (g239) & (!g240)));
	assign g242 = (((!g199) & (!g200) & (!g203) & (!g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (!g203) & (!g202) & (g209) & (g204)) + ((!g199) & (!g200) & (!g203) & (g202) & (g209) & (g204)) + ((!g199) & (!g200) & (g203) & (!g202) & (!g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (!g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (g203) & (!g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (!g202) & (g209) & (g204)) + ((!g199) & (!g200) & (g203) & (g202) & (!g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (g202) & (!g209) & (g204)) + ((!g199) & (g200) & (!g203) & (!g202) & (!g209) & (g204)) + ((!g199) & (g200) & (!g203) & (!g202) & (g209) & (!g204)) + ((!g199) & (g200) & (!g203) & (g202) & (g209) & (g204)) + ((!g199) & (g200) & (g203) & (!g202) & (g209) & (!g204)) + ((!g199) & (g200) & (g203) & (!g202) & (g209) & (g204)) + ((!g199) & (g200) & (g203) & (g202) & (!g209) & (!g204)) + ((!g199) & (g200) & (g203) & (g202) & (!g209) & (g204)) + ((!g199) & (g200) & (g203) & (g202) & (g209) & (g204)) + ((g199) & (!g200) & (!g203) & (!g202) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g202) & (g209) & (g204)) + ((g199) & (!g200) & (!g203) & (g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (g202) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (g202) & (g209) & (g204)) + ((g199) & (!g200) & (g203) & (!g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (g203) & (!g202) & (g209) & (!g204)) + ((g199) & (!g200) & (g203) & (g202) & (g209) & (!g204)) + ((g199) & (g200) & (!g203) & (!g202) & (g209) & (g204)) + ((g199) & (g200) & (g203) & (!g202) & (!g209) & (!g204)) + ((g199) & (g200) & (g203) & (!g202) & (g209) & (g204)));
	assign g243 = (((!g199) & (!g200) & (!g203) & (!g202) & (!g209) & (!g204)) + ((!g199) & (!g200) & (!g203) & (g202) & (!g209) & (!g204)) + ((!g199) & (!g200) & (!g203) & (g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (!g203) & (g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (!g202) & (g209) & (g204)) + ((!g199) & (!g200) & (g203) & (g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (g203) & (g202) & (g209) & (g204)) + ((!g199) & (g200) & (!g203) & (!g202) & (!g209) & (!g204)) + ((!g199) & (g200) & (!g203) & (!g202) & (g209) & (!g204)) + ((!g199) & (g200) & (g203) & (!g202) & (!g209) & (g204)) + ((!g199) & (g200) & (g203) & (!g202) & (g209) & (g204)) + ((!g199) & (g200) & (g203) & (g202) & (!g209) & (g204)) + ((!g199) & (g200) & (g203) & (g202) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g202) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g202) & (g209) & (g204)) + ((g199) & (!g200) & (!g203) & (g202) & (!g209) & (g204)) + ((g199) & (!g200) & (!g203) & (g202) & (g209) & (g204)) + ((g199) & (!g200) & (g203) & (g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (g203) & (g202) & (!g209) & (g204)) + ((g199) & (!g200) & (g203) & (g202) & (g209) & (g204)) + ((g199) & (g200) & (!g203) & (!g202) & (!g209) & (g204)) + ((g199) & (g200) & (!g203) & (!g202) & (g209) & (!g204)) + ((g199) & (g200) & (!g203) & (g202) & (g209) & (!g204)) + ((g199) & (g200) & (g203) & (!g202) & (!g209) & (g204)) + ((g199) & (g200) & (g203) & (!g202) & (g209) & (g204)) + ((g199) & (g200) & (g203) & (g202) & (!g209) & (!g204)) + ((g199) & (g200) & (g203) & (g202) & (g209) & (g204)));
	assign g244 = (((!g199) & (!g200) & (!g203) & (!g202) & (g209) & (g204)) + ((!g199) & (!g200) & (!g203) & (g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (!g202) & (!g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (!g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (g203) & (!g202) & (g209) & (g204)) + ((!g199) & (!g200) & (g203) & (g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (g203) & (g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (g203) & (g202) & (g209) & (g204)) + ((!g199) & (g200) & (!g203) & (!g202) & (g209) & (!g204)) + ((!g199) & (g200) & (!g203) & (!g202) & (g209) & (g204)) + ((!g199) & (g200) & (g203) & (!g202) & (!g209) & (!g204)) + ((!g199) & (g200) & (g203) & (g202) & (!g209) & (g204)) + ((!g199) & (g200) & (g203) & (g202) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g202) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (!g202) & (g209) & (g204)) + ((g199) & (!g200) & (!g203) & (g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (g202) & (!g209) & (g204)) + ((g199) & (!g200) & (g203) & (!g202) & (!g209) & (g204)) + ((g199) & (!g200) & (g203) & (!g202) & (g209) & (g204)) + ((g199) & (!g200) & (g203) & (g202) & (g209) & (!g204)) + ((g199) & (g200) & (!g203) & (!g202) & (!g209) & (!g204)) + ((g199) & (g200) & (!g203) & (!g202) & (!g209) & (g204)) + ((g199) & (g200) & (!g203) & (!g202) & (g209) & (g204)) + ((g199) & (g200) & (!g203) & (g202) & (!g209) & (g204)) + ((g199) & (g200) & (!g203) & (g202) & (g209) & (!g204)) + ((g199) & (g200) & (g203) & (!g202) & (!g209) & (g204)) + ((g199) & (g200) & (g203) & (!g202) & (g209) & (!g204)) + ((g199) & (g200) & (g203) & (g202) & (!g209) & (!g204)) + ((g199) & (g200) & (g203) & (g202) & (g209) & (!g204)) + ((g199) & (g200) & (g203) & (g202) & (g209) & (g204)));
	assign g245 = (((!g199) & (!g200) & (!g203) & (!g202) & (g209) & (!g204)) + ((!g199) & (!g200) & (!g203) & (g202) & (!g209) & (!g204)) + ((!g199) & (!g200) & (!g203) & (g202) & (g209) & (g204)) + ((!g199) & (!g200) & (g203) & (!g202) & (!g209) & (g204)) + ((!g199) & (!g200) & (g203) & (!g202) & (g209) & (g204)) + ((!g199) & (!g200) & (g203) & (g202) & (g209) & (g204)) + ((!g199) & (g200) & (!g203) & (!g202) & (!g209) & (g204)) + ((!g199) & (g200) & (!g203) & (g202) & (!g209) & (g204)) + ((!g199) & (g200) & (!g203) & (g202) & (g209) & (g204)) + ((!g199) & (g200) & (g203) & (!g202) & (!g209) & (!g204)) + ((!g199) & (g200) & (g203) & (!g202) & (g209) & (!g204)) + ((!g199) & (g200) & (g203) & (g202) & (!g209) & (g204)) + ((!g199) & (g200) & (g203) & (g202) & (g209) & (g204)) + ((g199) & (!g200) & (!g203) & (!g202) & (g209) & (!g204)) + ((g199) & (!g200) & (!g203) & (g202) & (g209) & (g204)) + ((g199) & (!g200) & (g203) & (!g202) & (!g209) & (!g204)) + ((g199) & (!g200) & (g203) & (!g202) & (g209) & (g204)) + ((g199) & (!g200) & (g203) & (g202) & (!g209) & (!g204)) + ((g199) & (g200) & (!g203) & (!g202) & (g209) & (g204)) + ((g199) & (g200) & (!g203) & (g202) & (!g209) & (!g204)) + ((g199) & (g200) & (!g203) & (g202) & (!g209) & (g204)) + ((g199) & (g200) & (g203) & (!g202) & (g209) & (g204)));
	assign g246 = (((!g242) & (!g243) & (!g244) & (!g245) & (!g210) & (!g201)) + ((!g242) & (!g243) & (!g244) & (!g245) & (!g210) & (g201)) + ((!g242) & (!g243) & (!g244) & (!g245) & (g210) & (!g201)) + ((!g242) & (!g243) & (!g244) & (g245) & (!g210) & (!g201)) + ((!g242) & (!g243) & (!g244) & (g245) & (!g210) & (g201)) + ((!g242) & (!g243) & (!g244) & (g245) & (g210) & (!g201)) + ((!g242) & (!g243) & (!g244) & (g245) & (g210) & (g201)) + ((!g242) & (!g243) & (g244) & (!g245) & (!g210) & (!g201)) + ((!g242) & (!g243) & (g244) & (!g245) & (g210) & (!g201)) + ((!g242) & (!g243) & (g244) & (g245) & (!g210) & (!g201)) + ((!g242) & (!g243) & (g244) & (g245) & (g210) & (!g201)) + ((!g242) & (!g243) & (g244) & (g245) & (g210) & (g201)) + ((!g242) & (g243) & (!g244) & (!g245) & (!g210) & (!g201)) + ((!g242) & (g243) & (!g244) & (!g245) & (!g210) & (g201)) + ((!g242) & (g243) & (!g244) & (g245) & (!g210) & (!g201)) + ((!g242) & (g243) & (!g244) & (g245) & (!g210) & (g201)) + ((!g242) & (g243) & (!g244) & (g245) & (g210) & (g201)) + ((!g242) & (g243) & (g244) & (!g245) & (!g210) & (!g201)) + ((!g242) & (g243) & (g244) & (g245) & (!g210) & (!g201)) + ((!g242) & (g243) & (g244) & (g245) & (g210) & (g201)) + ((g242) & (!g243) & (!g244) & (!g245) & (!g210) & (g201)) + ((g242) & (!g243) & (!g244) & (!g245) & (g210) & (!g201)) + ((g242) & (!g243) & (!g244) & (g245) & (!g210) & (g201)) + ((g242) & (!g243) & (!g244) & (g245) & (g210) & (!g201)) + ((g242) & (!g243) & (!g244) & (g245) & (g210) & (g201)) + ((g242) & (!g243) & (g244) & (!g245) & (g210) & (!g201)) + ((g242) & (!g243) & (g244) & (g245) & (g210) & (!g201)) + ((g242) & (!g243) & (g244) & (g245) & (g210) & (g201)) + ((g242) & (g243) & (!g244) & (!g245) & (!g210) & (g201)) + ((g242) & (g243) & (!g244) & (g245) & (!g210) & (g201)) + ((g242) & (g243) & (!g244) & (g245) & (g210) & (g201)) + ((g242) & (g243) & (g244) & (g245) & (g210) & (g201)));
	assign g248 = (((!g246) & (sk[84]) & (g247)) + ((g246) & (!sk[84]) & (!g247)) + ((g246) & (!sk[84]) & (g247)) + ((g246) & (sk[84]) & (!g247)));
	assign g249 = (((!g199) & (!g210) & (!g201) & (!g202) & (!g209) & (g204)) + ((!g199) & (!g210) & (!g201) & (!g202) & (g209) & (g204)) + ((!g199) & (!g210) & (!g201) & (g202) & (!g209) & (!g204)) + ((!g199) & (!g210) & (!g201) & (g202) & (!g209) & (g204)) + ((!g199) & (!g210) & (!g201) & (g202) & (g209) & (!g204)) + ((!g199) & (!g210) & (!g201) & (g202) & (g209) & (g204)) + ((!g199) & (!g210) & (g201) & (!g202) & (!g209) & (g204)) + ((!g199) & (!g210) & (g201) & (!g202) & (g209) & (g204)) + ((!g199) & (!g210) & (g201) & (g202) & (g209) & (!g204)) + ((!g199) & (g210) & (g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (g210) & (g201) & (!g202) & (g209) & (g204)) + ((!g199) & (g210) & (g201) & (g202) & (!g209) & (g204)) + ((g199) & (!g210) & (!g201) & (!g202) & (g209) & (!g204)) + ((g199) & (!g210) & (!g201) & (g202) & (!g209) & (!g204)) + ((g199) & (!g210) & (!g201) & (g202) & (!g209) & (g204)) + ((g199) & (!g210) & (!g201) & (g202) & (g209) & (g204)) + ((g199) & (!g210) & (g201) & (!g202) & (!g209) & (g204)) + ((g199) & (!g210) & (g201) & (!g202) & (g209) & (g204)) + ((g199) & (!g210) & (g201) & (g202) & (g209) & (!g204)) + ((g199) & (!g210) & (g201) & (g202) & (g209) & (g204)) + ((g199) & (g210) & (!g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (g210) & (!g201) & (!g202) & (!g209) & (g204)) + ((g199) & (g210) & (!g201) & (!g202) & (g209) & (!g204)) + ((g199) & (g210) & (!g201) & (g202) & (!g209) & (!g204)) + ((g199) & (g210) & (g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (g210) & (g201) & (!g202) & (!g209) & (g204)) + ((g199) & (g210) & (g201) & (!g202) & (g209) & (!g204)) + ((g199) & (g210) & (g201) & (g202) & (!g209) & (g204)));
	assign g250 = (((!g199) & (!g210) & (!g201) & (!g202) & (!g209) & (!g204)) + ((!g199) & (!g210) & (!g201) & (g202) & (g209) & (g204)) + ((!g199) & (!g210) & (g201) & (!g202) & (!g209) & (!g204)) + ((!g199) & (!g210) & (g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (!g210) & (g201) & (!g202) & (g209) & (g204)) + ((!g199) & (!g210) & (g201) & (g202) & (!g209) & (!g204)) + ((!g199) & (!g210) & (g201) & (g202) & (g209) & (g204)) + ((!g199) & (g210) & (!g201) & (!g202) & (!g209) & (!g204)) + ((!g199) & (g210) & (!g201) & (!g202) & (g209) & (g204)) + ((!g199) & (g210) & (!g201) & (g202) & (!g209) & (g204)) + ((!g199) & (g210) & (g201) & (!g202) & (!g209) & (!g204)) + ((!g199) & (g210) & (g201) & (!g202) & (g209) & (g204)) + ((!g199) & (g210) & (g201) & (g202) & (g209) & (!g204)) + ((!g199) & (g210) & (g201) & (g202) & (g209) & (g204)) + ((g199) & (!g210) & (!g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (!g210) & (!g201) & (!g202) & (g209) & (g204)) + ((g199) & (!g210) & (!g201) & (g202) & (!g209) & (!g204)) + ((g199) & (!g210) & (!g201) & (g202) & (g209) & (g204)) + ((g199) & (!g210) & (g201) & (!g202) & (g209) & (g204)) + ((g199) & (!g210) & (g201) & (g202) & (!g209) & (g204)) + ((g199) & (g210) & (!g201) & (!g202) & (g209) & (!g204)) + ((g199) & (g210) & (!g201) & (!g202) & (g209) & (g204)) + ((g199) & (g210) & (!g201) & (g202) & (!g209) & (g204)) + ((g199) & (g210) & (!g201) & (g202) & (g209) & (!g204)) + ((g199) & (g210) & (!g201) & (g202) & (g209) & (g204)) + ((g199) & (g210) & (g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (g210) & (g201) & (!g202) & (g209) & (!g204)) + ((g199) & (g210) & (g201) & (g202) & (!g209) & (!g204)));
	assign g251 = (((!g199) & (!g210) & (!g201) & (!g202) & (!g209) & (g204)) + ((!g199) & (!g210) & (!g201) & (!g202) & (g209) & (g204)) + ((!g199) & (!g210) & (!g201) & (g202) & (g209) & (!g204)) + ((!g199) & (!g210) & (!g201) & (g202) & (g209) & (g204)) + ((!g199) & (!g210) & (g201) & (!g202) & (g209) & (g204)) + ((!g199) & (!g210) & (g201) & (g202) & (!g209) & (!g204)) + ((!g199) & (!g210) & (g201) & (g202) & (!g209) & (g204)) + ((!g199) & (!g210) & (g201) & (g202) & (g209) & (g204)) + ((!g199) & (g210) & (!g201) & (!g202) & (!g209) & (!g204)) + ((!g199) & (g210) & (!g201) & (!g202) & (!g209) & (g204)) + ((!g199) & (g210) & (!g201) & (!g202) & (g209) & (g204)) + ((!g199) & (g210) & (!g201) & (g202) & (!g209) & (g204)) + ((!g199) & (g210) & (!g201) & (g202) & (g209) & (!g204)) + ((!g199) & (g210) & (g201) & (!g202) & (!g209) & (g204)) + ((!g199) & (g210) & (g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (g210) & (g201) & (g202) & (!g209) & (!g204)) + ((!g199) & (g210) & (g201) & (g202) & (g209) & (!g204)) + ((!g199) & (g210) & (g201) & (g202) & (g209) & (g204)) + ((g199) & (!g210) & (!g201) & (!g202) & (!g209) & (g204)) + ((g199) & (!g210) & (!g201) & (g202) & (!g209) & (!g204)) + ((g199) & (!g210) & (!g201) & (g202) & (g209) & (!g204)) + ((g199) & (!g210) & (g201) & (!g202) & (g209) & (g204)) + ((g199) & (!g210) & (g201) & (g202) & (!g209) & (g204)) + ((g199) & (g210) & (!g201) & (!g202) & (!g209) & (g204)) + ((g199) & (g210) & (!g201) & (g202) & (!g209) & (!g204)) + ((g199) & (g210) & (!g201) & (g202) & (g209) & (!g204)) + ((g199) & (g210) & (g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (g210) & (g201) & (!g202) & (g209) & (!g204)) + ((g199) & (g210) & (g201) & (!g202) & (g209) & (g204)) + ((g199) & (g210) & (g201) & (g202) & (g209) & (g204)));
	assign g252 = (((!g199) & (!g210) & (!g201) & (!g202) & (g209) & (g204)) + ((!g199) & (!g210) & (!g201) & (g202) & (!g209) & (!g204)) + ((!g199) & (!g210) & (!g201) & (g202) & (g209) & (g204)) + ((!g199) & (!g210) & (g201) & (!g202) & (!g209) & (!g204)) + ((!g199) & (!g210) & (g201) & (g202) & (g209) & (!g204)) + ((!g199) & (!g210) & (g201) & (g202) & (g209) & (g204)) + ((!g199) & (g210) & (!g201) & (g202) & (!g209) & (!g204)) + ((!g199) & (g210) & (!g201) & (g202) & (g209) & (!g204)) + ((!g199) & (g210) & (g201) & (!g202) & (g209) & (!g204)) + ((!g199) & (g210) & (g201) & (!g202) & (g209) & (g204)) + ((g199) & (!g210) & (!g201) & (!g202) & (!g209) & (g204)) + ((g199) & (!g210) & (!g201) & (!g202) & (g209) & (!g204)) + ((g199) & (!g210) & (!g201) & (g202) & (!g209) & (g204)) + ((g199) & (!g210) & (g201) & (!g202) & (g209) & (!g204)) + ((g199) & (!g210) & (g201) & (!g202) & (g209) & (g204)) + ((g199) & (!g210) & (g201) & (g202) & (g209) & (!g204)) + ((g199) & (!g210) & (g201) & (g202) & (g209) & (g204)) + ((g199) & (g210) & (!g201) & (!g202) & (g209) & (!g204)) + ((g199) & (g210) & (!g201) & (g202) & (!g209) & (g204)) + ((g199) & (g210) & (g201) & (!g202) & (!g209) & (!g204)) + ((g199) & (g210) & (g201) & (!g202) & (g209) & (g204)) + ((g199) & (g210) & (g201) & (g202) & (!g209) & (g204)));
	assign g253 = (((!g249) & (!g250) & (!g251) & (!g252) & (!g203) & (!g200)) + ((!g249) & (!g250) & (!g251) & (!g252) & (!g203) & (g200)) + ((!g249) & (!g250) & (!g251) & (!g252) & (g203) & (!g200)) + ((!g249) & (!g250) & (!g251) & (g252) & (!g203) & (!g200)) + ((!g249) & (!g250) & (!g251) & (g252) & (!g203) & (g200)) + ((!g249) & (!g250) & (!g251) & (g252) & (g203) & (!g200)) + ((!g249) & (!g250) & (!g251) & (g252) & (g203) & (g200)) + ((!g249) & (!g250) & (g251) & (!g252) & (!g203) & (!g200)) + ((!g249) & (!g250) & (g251) & (!g252) & (g203) & (!g200)) + ((!g249) & (!g250) & (g251) & (g252) & (!g203) & (!g200)) + ((!g249) & (!g250) & (g251) & (g252) & (g203) & (!g200)) + ((!g249) & (!g250) & (g251) & (g252) & (g203) & (g200)) + ((!g249) & (g250) & (!g251) & (!g252) & (!g203) & (!g200)) + ((!g249) & (g250) & (!g251) & (!g252) & (!g203) & (g200)) + ((!g249) & (g250) & (!g251) & (g252) & (!g203) & (!g200)) + ((!g249) & (g250) & (!g251) & (g252) & (!g203) & (g200)) + ((!g249) & (g250) & (!g251) & (g252) & (g203) & (g200)) + ((!g249) & (g250) & (g251) & (!g252) & (!g203) & (!g200)) + ((!g249) & (g250) & (g251) & (g252) & (!g203) & (!g200)) + ((!g249) & (g250) & (g251) & (g252) & (g203) & (g200)) + ((g249) & (!g250) & (!g251) & (!g252) & (!g203) & (g200)) + ((g249) & (!g250) & (!g251) & (!g252) & (g203) & (!g200)) + ((g249) & (!g250) & (!g251) & (g252) & (!g203) & (g200)) + ((g249) & (!g250) & (!g251) & (g252) & (g203) & (!g200)) + ((g249) & (!g250) & (!g251) & (g252) & (g203) & (g200)) + ((g249) & (!g250) & (g251) & (!g252) & (g203) & (!g200)) + ((g249) & (!g250) & (g251) & (g252) & (g203) & (!g200)) + ((g249) & (!g250) & (g251) & (g252) & (g203) & (g200)) + ((g249) & (g250) & (!g251) & (!g252) & (!g203) & (g200)) + ((g249) & (g250) & (!g251) & (g252) & (!g203) & (g200)) + ((g249) & (g250) & (!g251) & (g252) & (g203) & (g200)) + ((g249) & (g250) & (g251) & (g252) & (g203) & (g200)));
	assign g255 = (((!g253) & (sk[90]) & (g254)) + ((g253) & (!sk[90]) & (!g254)) + ((g253) & (!sk[90]) & (g254)) + ((g253) & (sk[90]) & (!g254)));
	assign g256 = (((!g203) & (!g200) & (!g201) & (!g202) & (!g209) & (g210)) + ((!g203) & (!g200) & (!g201) & (!g202) & (g209) & (!g210)) + ((!g203) & (!g200) & (!g201) & (g202) & (!g209) & (g210)) + ((!g203) & (!g200) & (!g201) & (g202) & (g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (!g202) & (!g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (!g202) & (g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (g202) & (!g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (g202) & (g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (g202) & (g209) & (g210)) + ((!g203) & (g200) & (!g201) & (!g202) & (g209) & (!g210)) + ((!g203) & (g200) & (!g201) & (g202) & (g209) & (!g210)) + ((!g203) & (g200) & (!g201) & (g202) & (g209) & (g210)) + ((!g203) & (g200) & (g201) & (!g202) & (g209) & (g210)) + ((!g203) & (g200) & (g201) & (g202) & (!g209) & (!g210)) + ((g203) & (!g200) & (!g201) & (!g202) & (!g209) & (g210)) + ((g203) & (!g200) & (!g201) & (g202) & (!g209) & (g210)) + ((g203) & (!g200) & (g201) & (g202) & (g209) & (g210)) + ((g203) & (g200) & (!g201) & (!g202) & (g209) & (g210)) + ((g203) & (g200) & (!g201) & (g202) & (!g209) & (!g210)) + ((g203) & (g200) & (!g201) & (g202) & (g209) & (!g210)) + ((g203) & (g200) & (g201) & (!g202) & (!g209) & (g210)) + ((g203) & (g200) & (g201) & (!g202) & (g209) & (!g210)) + ((g203) & (g200) & (g201) & (!g202) & (g209) & (g210)) + ((g203) & (g200) & (g201) & (g202) & (!g209) & (g210)));
	assign g257 = (((!g203) & (!g200) & (!g201) & (!g202) & (!g209) & (!g210)) + ((!g203) & (!g200) & (!g201) & (!g202) & (!g209) & (g210)) + ((!g203) & (!g200) & (!g201) & (g202) & (!g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (!g202) & (!g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (!g202) & (g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (!g202) & (g209) & (g210)) + ((!g203) & (!g200) & (g201) & (g202) & (!g209) & (g210)) + ((!g203) & (!g200) & (g201) & (g202) & (g209) & (g210)) + ((!g203) & (g200) & (!g201) & (!g202) & (!g209) & (!g210)) + ((!g203) & (g200) & (!g201) & (!g202) & (g209) & (!g210)) + ((!g203) & (g200) & (!g201) & (g202) & (!g209) & (!g210)) + ((!g203) & (g200) & (!g201) & (g202) & (!g209) & (g210)) + ((!g203) & (g200) & (!g201) & (g202) & (g209) & (g210)) + ((!g203) & (g200) & (g201) & (!g202) & (!g209) & (g210)) + ((!g203) & (g200) & (g201) & (g202) & (!g209) & (!g210)) + ((!g203) & (g200) & (g201) & (g202) & (!g209) & (g210)) + ((g203) & (!g200) & (!g201) & (!g202) & (!g209) & (g210)) + ((g203) & (!g200) & (!g201) & (!g202) & (g209) & (g210)) + ((g203) & (!g200) & (!g201) & (g202) & (!g209) & (!g210)) + ((g203) & (!g200) & (!g201) & (g202) & (g209) & (g210)) + ((g203) & (!g200) & (g201) & (!g202) & (!g209) & (!g210)) + ((g203) & (!g200) & (g201) & (!g202) & (g209) & (g210)) + ((g203) & (!g200) & (g201) & (g202) & (g209) & (!g210)) + ((g203) & (g200) & (!g201) & (!g202) & (!g209) & (!g210)) + ((g203) & (g200) & (!g201) & (!g202) & (!g209) & (g210)) + ((g203) & (g200) & (!g201) & (!g202) & (g209) & (g210)) + ((g203) & (g200) & (!g201) & (g202) & (!g209) & (g210)) + ((g203) & (g200) & (!g201) & (g202) & (g209) & (!g210)) + ((g203) & (g200) & (g201) & (!g202) & (g209) & (!g210)) + ((g203) & (g200) & (g201) & (!g202) & (g209) & (g210)));
	assign g258 = (((!g203) & (!g200) & (!g201) & (!g202) & (g209) & (!g210)) + ((!g203) & (!g200) & (!g201) & (g202) & (!g209) & (!g210)) + ((!g203) & (!g200) & (!g201) & (g202) & (g209) & (!g210)) + ((!g203) & (!g200) & (!g201) & (g202) & (g209) & (g210)) + ((!g203) & (!g200) & (g201) & (!g202) & (!g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (!g202) & (!g209) & (g210)) + ((!g203) & (!g200) & (g201) & (!g202) & (g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (g202) & (!g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (g202) & (g209) & (g210)) + ((!g203) & (g200) & (!g201) & (!g202) & (!g209) & (g210)) + ((!g203) & (g200) & (!g201) & (!g202) & (g209) & (!g210)) + ((!g203) & (g200) & (!g201) & (!g202) & (g209) & (g210)) + ((!g203) & (g200) & (g201) & (!g202) & (!g209) & (g210)) + ((!g203) & (g200) & (g201) & (!g202) & (g209) & (!g210)) + ((!g203) & (g200) & (g201) & (!g202) & (g209) & (g210)) + ((!g203) & (g200) & (g201) & (g202) & (!g209) & (!g210)) + ((g203) & (!g200) & (!g201) & (!g202) & (g209) & (!g210)) + ((g203) & (!g200) & (!g201) & (g202) & (!g209) & (!g210)) + ((g203) & (!g200) & (!g201) & (g202) & (g209) & (g210)) + ((g203) & (!g200) & (g201) & (!g202) & (!g209) & (!g210)) + ((g203) & (!g200) & (g201) & (!g202) & (!g209) & (g210)) + ((g203) & (!g200) & (g201) & (g202) & (!g209) & (!g210)) + ((g203) & (!g200) & (g201) & (g202) & (g209) & (!g210)) + ((g203) & (g200) & (!g201) & (!g202) & (g209) & (!g210)) + ((g203) & (g200) & (!g201) & (g202) & (!g209) & (!g210)) + ((g203) & (g200) & (!g201) & (g202) & (g209) & (g210)) + ((g203) & (g200) & (g201) & (!g202) & (!g209) & (!g210)) + ((g203) & (g200) & (g201) & (!g202) & (g209) & (!g210)) + ((g203) & (g200) & (g201) & (!g202) & (g209) & (g210)) + ((g203) & (g200) & (g201) & (g202) & (!g209) & (g210)));
	assign g259 = (((!g203) & (!g200) & (!g201) & (!g202) & (!g209) & (g210)) + ((!g203) & (!g200) & (!g201) & (g202) & (g209) & (!g210)) + ((!g203) & (!g200) & (!g201) & (g202) & (g209) & (g210)) + ((!g203) & (!g200) & (g201) & (!g202) & (!g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (!g202) & (!g209) & (g210)) + ((!g203) & (!g200) & (g201) & (g202) & (g209) & (!g210)) + ((!g203) & (!g200) & (g201) & (g202) & (g209) & (g210)) + ((!g203) & (g200) & (!g201) & (!g202) & (!g209) & (!g210)) + ((!g203) & (g200) & (!g201) & (!g202) & (!g209) & (g210)) + ((!g203) & (g200) & (!g201) & (!g202) & (g209) & (g210)) + ((!g203) & (g200) & (!g201) & (g202) & (!g209) & (g210)) + ((!g203) & (g200) & (g201) & (!g202) & (!g209) & (g210)) + ((!g203) & (g200) & (g201) & (g202) & (!g209) & (!g210)) + ((!g203) & (g200) & (g201) & (g202) & (!g209) & (g210)) + ((!g203) & (g200) & (g201) & (g202) & (g209) & (!g210)) + ((!g203) & (g200) & (g201) & (g202) & (g209) & (g210)) + ((g203) & (!g200) & (!g201) & (g202) & (!g209) & (g210)) + ((g203) & (!g200) & (g201) & (!g202) & (!g209) & (!g210)) + ((g203) & (!g200) & (g201) & (g202) & (!g209) & (!g210)) + ((g203) & (!g200) & (g201) & (g202) & (!g209) & (g210)) + ((g203) & (!g200) & (g201) & (g202) & (g209) & (g210)) + ((g203) & (g200) & (!g201) & (!g202) & (!g209) & (g210)) + ((g203) & (g200) & (!g201) & (!g202) & (g209) & (g210)) + ((g203) & (g200) & (!g201) & (g202) & (!g209) & (!g210)) + ((g203) & (g200) & (!g201) & (g202) & (g209) & (!g210)) + ((g203) & (g200) & (!g201) & (g202) & (g209) & (g210)) + ((g203) & (g200) & (g201) & (!g202) & (g209) & (g210)) + ((g203) & (g200) & (g201) & (g202) & (g209) & (g210)));
	assign g260 = (((!g256) & (!g257) & (!g258) & (!g259) & (!g199) & (g204)) + ((!g256) & (!g257) & (!g258) & (!g259) & (g199) & (!g204)) + ((!g256) & (!g257) & (!g258) & (!g259) & (g199) & (g204)) + ((!g256) & (!g257) & (!g258) & (g259) & (!g199) & (g204)) + ((!g256) & (!g257) & (!g258) & (g259) & (g199) & (!g204)) + ((!g256) & (!g257) & (g258) & (!g259) & (g199) & (!g204)) + ((!g256) & (!g257) & (g258) & (!g259) & (g199) & (g204)) + ((!g256) & (!g257) & (g258) & (g259) & (g199) & (!g204)) + ((!g256) & (g257) & (!g258) & (!g259) & (!g199) & (g204)) + ((!g256) & (g257) & (!g258) & (!g259) & (g199) & (g204)) + ((!g256) & (g257) & (!g258) & (g259) & (!g199) & (g204)) + ((!g256) & (g257) & (g258) & (!g259) & (g199) & (g204)) + ((g256) & (!g257) & (!g258) & (!g259) & (!g199) & (!g204)) + ((g256) & (!g257) & (!g258) & (!g259) & (!g199) & (g204)) + ((g256) & (!g257) & (!g258) & (!g259) & (g199) & (!g204)) + ((g256) & (!g257) & (!g258) & (!g259) & (g199) & (g204)) + ((g256) & (!g257) & (!g258) & (g259) & (!g199) & (!g204)) + ((g256) & (!g257) & (!g258) & (g259) & (!g199) & (g204)) + ((g256) & (!g257) & (!g258) & (g259) & (g199) & (!g204)) + ((g256) & (!g257) & (g258) & (!g259) & (!g199) & (!g204)) + ((g256) & (!g257) & (g258) & (!g259) & (g199) & (!g204)) + ((g256) & (!g257) & (g258) & (!g259) & (g199) & (g204)) + ((g256) & (!g257) & (g258) & (g259) & (!g199) & (!g204)) + ((g256) & (!g257) & (g258) & (g259) & (g199) & (!g204)) + ((g256) & (g257) & (!g258) & (!g259) & (!g199) & (!g204)) + ((g256) & (g257) & (!g258) & (!g259) & (!g199) & (g204)) + ((g256) & (g257) & (!g258) & (!g259) & (g199) & (g204)) + ((g256) & (g257) & (!g258) & (g259) & (!g199) & (!g204)) + ((g256) & (g257) & (!g258) & (g259) & (!g199) & (g204)) + ((g256) & (g257) & (g258) & (!g259) & (!g199) & (!g204)) + ((g256) & (g257) & (g258) & (!g259) & (g199) & (g204)) + ((g256) & (g257) & (g258) & (g259) & (!g199) & (!g204)));
	assign g262 = (((!g260) & (sk[96]) & (g261)) + ((g260) & (!sk[96]) & (!g261)) + ((g260) & (!sk[96]) & (g261)) + ((g260) & (sk[96]) & (!g261)));
	assign g269 = (((!g263) & (!g264) & (!g265) & (!g266) & (g267) & (g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g267) & (!g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g267) & (g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (g267) & (!g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (!g267) & (!g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (!g267) & (g268)) + ((!g263) & (!g264) & (g265) & (g266) & (!g267) & (!g268)) + ((!g263) & (!g264) & (g265) & (g266) & (g267) & (g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (g267) & (!g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (g267) & (g268)) + ((!g263) & (g264) & (!g265) & (g266) & (g267) & (!g268)) + ((!g263) & (g264) & (!g265) & (g266) & (g267) & (g268)) + ((!g263) & (g264) & (g265) & (!g266) & (g267) & (!g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (!g267) & (!g268)) + ((g263) & (!g264) & (g265) & (!g266) & (g267) & (!g268)) + ((g263) & (!g264) & (g265) & (g266) & (!g267) & (g268)) + ((g263) & (!g264) & (g265) & (g266) & (g267) & (g268)) + ((g263) & (g264) & (!g265) & (!g266) & (!g267) & (g268)) + ((g263) & (g264) & (!g265) & (!g266) & (g267) & (!g268)) + ((g263) & (g264) & (g265) & (!g266) & (!g267) & (g268)) + ((g263) & (g264) & (g265) & (!g266) & (g267) & (!g268)) + ((g263) & (g264) & (g265) & (g266) & (!g267) & (!g268)) + ((g263) & (g264) & (g265) & (g266) & (g267) & (!g268)) + ((g263) & (g264) & (g265) & (g266) & (g267) & (g268)));
	assign g270 = (((!g263) & (!g264) & (!g265) & (!g266) & (g267) & (!g268)) + ((!g263) & (!g264) & (!g265) & (!g266) & (g267) & (g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g267) & (!g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g267) & (g268)) + ((!g263) & (!g264) & (g265) & (g266) & (!g267) & (g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (!g267) & (!g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (!g267) & (g268)) + ((!g263) & (g264) & (g265) & (!g266) & (!g267) & (!g268)) + ((!g263) & (g264) & (g265) & (!g266) & (!g267) & (g268)) + ((!g263) & (g264) & (g265) & (!g266) & (g267) & (!g268)) + ((!g263) & (g264) & (g265) & (g266) & (g267) & (g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (!g267) & (g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (g267) & (!g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (g267) & (g268)) + ((g263) & (!g264) & (!g265) & (g266) & (g267) & (!g268)) + ((g263) & (!g264) & (g265) & (!g266) & (!g267) & (!g268)) + ((g263) & (!g264) & (g265) & (!g266) & (g267) & (g268)) + ((g263) & (!g264) & (g265) & (g266) & (!g267) & (g268)) + ((g263) & (!g264) & (g265) & (g266) & (g267) & (g268)) + ((g263) & (g264) & (!g265) & (!g266) & (!g267) & (!g268)) + ((g263) & (g264) & (!g265) & (!g266) & (!g267) & (g268)) + ((g263) & (g264) & (!g265) & (!g266) & (g267) & (!g268)) + ((g263) & (g264) & (!g265) & (!g266) & (g267) & (g268)) + ((g263) & (g264) & (!g265) & (g266) & (!g267) & (!g268)) + ((g263) & (g264) & (!g265) & (g266) & (g267) & (!g268)) + ((g263) & (g264) & (!g265) & (g266) & (g267) & (g268)) + ((g263) & (g264) & (g265) & (!g266) & (g267) & (!g268)) + ((g263) & (g264) & (g265) & (!g266) & (g267) & (g268)) + ((g263) & (g264) & (g265) & (g266) & (!g267) & (g268)) + ((g263) & (g264) & (g265) & (g266) & (g267) & (!g268)));
	assign g271 = (((!g263) & (!g264) & (!g265) & (!g266) & (!g267) & (!g268)) + ((!g263) & (!g264) & (!g265) & (!g266) & (g267) & (g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (g267) & (g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (!g267) & (!g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (!g267) & (g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (g267) & (g268)) + ((!g263) & (!g264) & (g265) & (g266) & (!g267) & (g268)) + ((!g263) & (!g264) & (g265) & (g266) & (g267) & (!g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (!g267) & (!g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (g267) & (!g268)) + ((!g263) & (g264) & (!g265) & (g266) & (g267) & (g268)) + ((!g263) & (g264) & (g265) & (g266) & (!g267) & (!g268)) + ((!g263) & (g264) & (g265) & (g266) & (g267) & (!g268)) + ((g263) & (!g264) & (!g265) & (g266) & (!g267) & (!g268)) + ((g263) & (!g264) & (!g265) & (g266) & (!g267) & (g268)) + ((g263) & (!g264) & (!g265) & (g266) & (g267) & (!g268)) + ((g263) & (!g264) & (g265) & (!g266) & (!g267) & (!g268)) + ((g263) & (!g264) & (g265) & (!g266) & (g267) & (g268)) + ((g263) & (!g264) & (g265) & (g266) & (!g267) & (!g268)) + ((g263) & (!g264) & (g265) & (g266) & (!g267) & (g268)) + ((g263) & (!g264) & (g265) & (g266) & (g267) & (!g268)) + ((g263) & (!g264) & (g265) & (g266) & (g267) & (g268)) + ((g263) & (g264) & (!g265) & (!g266) & (g267) & (g268)) + ((g263) & (g264) & (!g265) & (g266) & (!g267) & (!g268)) + ((g263) & (g264) & (!g265) & (g266) & (g267) & (!g268)) + ((g263) & (g264) & (!g265) & (g266) & (g267) & (g268)) + ((g263) & (g264) & (g265) & (!g266) & (!g267) & (!g268)) + ((g263) & (g264) & (g265) & (g266) & (!g267) & (!g268)) + ((g263) & (g264) & (g265) & (g266) & (!g267) & (g268)) + ((g263) & (g264) & (g265) & (g266) & (g267) & (g268)));
	assign g272 = (((!g263) & (!g264) & (!g265) & (!g266) & (!g267) & (g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (g267) & (!g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (g267) & (g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (!g267) & (g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (g267) & (g268)) + ((!g263) & (!g264) & (g265) & (g266) & (!g267) & (g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (!g267) & (!g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (!g267) & (g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (g267) & (!g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (g267) & (g268)) + ((!g263) & (g264) & (!g265) & (g266) & (g267) & (!g268)) + ((!g263) & (g264) & (!g265) & (g266) & (g267) & (g268)) + ((!g263) & (g264) & (g265) & (g266) & (!g267) & (!g268)) + ((!g263) & (g264) & (g265) & (g266) & (g267) & (!g268)) + ((!g263) & (g264) & (g265) & (g266) & (g267) & (g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (!g267) & (!g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (g267) & (g268)) + ((g263) & (!g264) & (!g265) & (g266) & (g267) & (!g268)) + ((g263) & (!g264) & (!g265) & (g266) & (g267) & (g268)) + ((g263) & (!g264) & (g265) & (!g266) & (!g267) & (g268)) + ((g263) & (!g264) & (g265) & (!g266) & (g267) & (!g268)) + ((g263) & (!g264) & (g265) & (g266) & (g267) & (!g268)) + ((g263) & (g264) & (!g265) & (!g266) & (!g267) & (g268)) + ((g263) & (g264) & (!g265) & (!g266) & (g267) & (g268)) + ((g263) & (g264) & (!g265) & (g266) & (g267) & (!g268)) + ((g263) & (g264) & (!g265) & (g266) & (g267) & (g268)) + ((g263) & (g264) & (g265) & (!g266) & (!g267) & (g268)) + ((g263) & (g264) & (g265) & (g266) & (!g267) & (!g268)));
	assign g275 = (((!g269) & (!g270) & (!g271) & (!g272) & (!g273) & (!g274)) + ((!g269) & (!g270) & (!g271) & (g272) & (!g273) & (!g274)) + ((!g269) & (!g270) & (!g271) & (g272) & (g273) & (g274)) + ((!g269) & (!g270) & (g271) & (!g272) & (!g273) & (!g274)) + ((!g269) & (!g270) & (g271) & (!g272) & (!g273) & (g274)) + ((!g269) & (!g270) & (g271) & (g272) & (!g273) & (!g274)) + ((!g269) & (!g270) & (g271) & (g272) & (!g273) & (g274)) + ((!g269) & (!g270) & (g271) & (g272) & (g273) & (g274)) + ((!g269) & (g270) & (!g271) & (!g272) & (!g273) & (!g274)) + ((!g269) & (g270) & (!g271) & (!g272) & (g273) & (!g274)) + ((!g269) & (g270) & (!g271) & (g272) & (!g273) & (!g274)) + ((!g269) & (g270) & (!g271) & (g272) & (g273) & (!g274)) + ((!g269) & (g270) & (!g271) & (g272) & (g273) & (g274)) + ((!g269) & (g270) & (g271) & (!g272) & (!g273) & (!g274)) + ((!g269) & (g270) & (g271) & (!g272) & (!g273) & (g274)) + ((!g269) & (g270) & (g271) & (!g272) & (g273) & (!g274)) + ((!g269) & (g270) & (g271) & (g272) & (!g273) & (!g274)) + ((!g269) & (g270) & (g271) & (g272) & (!g273) & (g274)) + ((!g269) & (g270) & (g271) & (g272) & (g273) & (!g274)) + ((!g269) & (g270) & (g271) & (g272) & (g273) & (g274)) + ((g269) & (!g270) & (!g271) & (g272) & (g273) & (g274)) + ((g269) & (!g270) & (g271) & (!g272) & (!g273) & (g274)) + ((g269) & (!g270) & (g271) & (g272) & (!g273) & (g274)) + ((g269) & (!g270) & (g271) & (g272) & (g273) & (g274)) + ((g269) & (g270) & (!g271) & (!g272) & (g273) & (!g274)) + ((g269) & (g270) & (!g271) & (g272) & (g273) & (!g274)) + ((g269) & (g270) & (!g271) & (g272) & (g273) & (g274)) + ((g269) & (g270) & (g271) & (!g272) & (!g273) & (g274)) + ((g269) & (g270) & (g271) & (!g272) & (g273) & (!g274)) + ((g269) & (g270) & (g271) & (g272) & (!g273) & (g274)) + ((g269) & (g270) & (g271) & (g272) & (g273) & (!g274)) + ((g269) & (g270) & (g271) & (g272) & (g273) & (g274)));
	assign g277 = (((!sk[102]) & (g275) & (!g276)) + ((!sk[102]) & (g275) & (g276)) + ((sk[102]) & (!g275) & (g276)) + ((sk[102]) & (g275) & (!g276)));
	assign g278 = (((!g263) & (!g264) & (!g265) & (!g266) & (!g273) & (g267)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g273) & (!g267)) + ((!g263) & (!g264) & (!g265) & (g266) & (g273) & (!g267)) + ((!g263) & (!g264) & (g265) & (!g266) & (g273) & (g267)) + ((!g263) & (!g264) & (g265) & (g266) & (!g273) & (g267)) + ((!g263) & (!g264) & (g265) & (g266) & (g273) & (!g267)) + ((!g263) & (g264) & (!g265) & (!g266) & (!g273) & (g267)) + ((!g263) & (g264) & (!g265) & (!g266) & (g273) & (!g267)) + ((!g263) & (g264) & (!g265) & (!g266) & (g273) & (g267)) + ((!g263) & (g264) & (g265) & (!g266) & (g273) & (g267)) + ((!g263) & (g264) & (g265) & (g266) & (g273) & (g267)) + ((g263) & (!g264) & (!g265) & (!g266) & (!g273) & (!g267)) + ((g263) & (!g264) & (!g265) & (!g266) & (g273) & (g267)) + ((g263) & (!g264) & (!g265) & (g266) & (!g273) & (!g267)) + ((g263) & (!g264) & (!g265) & (g266) & (g273) & (!g267)) + ((g263) & (!g264) & (g265) & (!g266) & (g273) & (!g267)) + ((g263) & (!g264) & (g265) & (!g266) & (g273) & (g267)) + ((g263) & (!g264) & (g265) & (g266) & (g273) & (!g267)) + ((g263) & (!g264) & (g265) & (g266) & (g273) & (g267)) + ((g263) & (g264) & (!g265) & (!g266) & (g273) & (!g267)) + ((g263) & (g264) & (!g265) & (!g266) & (g273) & (g267)) + ((g263) & (g264) & (!g265) & (g266) & (g273) & (g267)) + ((g263) & (g264) & (g265) & (!g266) & (!g273) & (!g267)) + ((g263) & (g264) & (g265) & (!g266) & (!g273) & (g267)) + ((g263) & (g264) & (g265) & (!g266) & (g273) & (!g267)) + ((g263) & (g264) & (g265) & (g266) & (!g273) & (g267)) + ((g263) & (g264) & (g265) & (g266) & (g273) & (!g267)));
	assign g279 = (((!g263) & (!g264) & (!g265) & (!g266) & (!g273) & (g267)) + ((!g263) & (!g264) & (!g265) & (!g266) & (g273) & (!g267)) + ((!g263) & (!g264) & (!g265) & (!g266) & (g273) & (g267)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g273) & (!g267)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g273) & (g267)) + ((!g263) & (!g264) & (!g265) & (g266) & (g273) & (g267)) + ((!g263) & (!g264) & (g265) & (!g266) & (g273) & (!g267)) + ((!g263) & (!g264) & (g265) & (g266) & (!g273) & (!g267)) + ((!g263) & (!g264) & (g265) & (g266) & (!g273) & (g267)) + ((!g263) & (!g264) & (g265) & (g266) & (g273) & (g267)) + ((!g263) & (g264) & (!g265) & (!g266) & (g273) & (g267)) + ((!g263) & (g264) & (!g265) & (g266) & (!g273) & (!g267)) + ((!g263) & (g264) & (!g265) & (g266) & (g273) & (!g267)) + ((!g263) & (g264) & (g265) & (!g266) & (g273) & (!g267)) + ((!g263) & (g264) & (g265) & (!g266) & (g273) & (g267)) + ((!g263) & (g264) & (g265) & (g266) & (!g273) & (!g267)) + ((g263) & (!g264) & (!g265) & (!g266) & (!g273) & (!g267)) + ((g263) & (!g264) & (!g265) & (g266) & (!g273) & (!g267)) + ((g263) & (!g264) & (!g265) & (g266) & (!g273) & (g267)) + ((g263) & (!g264) & (g265) & (!g266) & (!g273) & (g267)) + ((g263) & (!g264) & (g265) & (!g266) & (g273) & (g267)) + ((g263) & (!g264) & (g265) & (g266) & (!g273) & (!g267)) + ((g263) & (!g264) & (g265) & (g266) & (!g273) & (g267)) + ((g263) & (g264) & (!g265) & (g266) & (!g273) & (!g267)) + ((g263) & (g264) & (!g265) & (g266) & (g273) & (g267)) + ((g263) & (g264) & (g265) & (!g266) & (!g273) & (!g267)) + ((g263) & (g264) & (g265) & (!g266) & (!g273) & (g267)) + ((g263) & (g264) & (g265) & (!g266) & (g273) & (g267)) + ((g263) & (g264) & (g265) & (g266) & (!g273) & (!g267)) + ((g263) & (g264) & (g265) & (g266) & (!g273) & (g267)) + ((g263) & (g264) & (g265) & (g266) & (g273) & (!g267)));
	assign g280 = (((!g263) & (!g264) & (!g265) & (!g266) & (!g273) & (g267)) + ((!g263) & (!g264) & (!g265) & (g266) & (g273) & (!g267)) + ((!g263) & (!g264) & (g265) & (!g266) & (!g273) & (!g267)) + ((!g263) & (!g264) & (g265) & (!g266) & (g273) & (!g267)) + ((!g263) & (!g264) & (g265) & (g266) & (!g273) & (g267)) + ((!g263) & (!g264) & (g265) & (g266) & (g273) & (!g267)) + ((!g263) & (!g264) & (g265) & (g266) & (g273) & (g267)) + ((!g263) & (g264) & (!g265) & (!g266) & (!g273) & (!g267)) + ((!g263) & (g264) & (!g265) & (!g266) & (g273) & (!g267)) + ((!g263) & (g264) & (!g265) & (g266) & (!g273) & (!g267)) + ((!g263) & (g264) & (!g265) & (g266) & (g273) & (g267)) + ((!g263) & (g264) & (g265) & (!g266) & (g273) & (g267)) + ((!g263) & (g264) & (g265) & (g266) & (!g273) & (g267)) + ((!g263) & (g264) & (g265) & (g266) & (g273) & (!g267)) + ((g263) & (!g264) & (!g265) & (!g266) & (g273) & (g267)) + ((g263) & (!g264) & (!g265) & (g266) & (!g273) & (!g267)) + ((g263) & (!g264) & (!g265) & (g266) & (g273) & (!g267)) + ((g263) & (!g264) & (g265) & (!g266) & (!g273) & (!g267)) + ((g263) & (!g264) & (g265) & (!g266) & (!g273) & (g267)) + ((g263) & (!g264) & (g265) & (!g266) & (g273) & (!g267)) + ((g263) & (!g264) & (g265) & (!g266) & (g273) & (g267)) + ((g263) & (!g264) & (g265) & (g266) & (g273) & (!g267)) + ((g263) & (g264) & (!g265) & (!g266) & (!g273) & (g267)) + ((g263) & (g264) & (!g265) & (!g266) & (g273) & (g267)) + ((g263) & (g264) & (!g265) & (g266) & (!g273) & (g267)) + ((g263) & (g264) & (g265) & (!g266) & (!g273) & (!g267)) + ((g263) & (g264) & (g265) & (!g266) & (!g273) & (g267)) + ((g263) & (g264) & (g265) & (!g266) & (g273) & (g267)) + ((g263) & (g264) & (g265) & (g266) & (!g273) & (!g267)) + ((g263) & (g264) & (g265) & (g266) & (!g273) & (g267)) + ((g263) & (g264) & (g265) & (g266) & (g273) & (!g267)) + ((g263) & (g264) & (g265) & (g266) & (g273) & (g267)));
	assign g281 = (((!g263) & (!g264) & (!g265) & (!g266) & (g273) & (!g267)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g273) & (!g267)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g273) & (g267)) + ((!g263) & (!g264) & (g265) & (!g266) & (g273) & (g267)) + ((!g263) & (!g264) & (g265) & (g266) & (!g273) & (g267)) + ((!g263) & (g264) & (!g265) & (!g266) & (!g273) & (!g267)) + ((!g263) & (g264) & (!g265) & (!g266) & (g273) & (!g267)) + ((!g263) & (g264) & (!g265) & (g266) & (!g273) & (g267)) + ((!g263) & (g264) & (g265) & (!g266) & (!g273) & (g267)) + ((!g263) & (g264) & (g265) & (!g266) & (g273) & (!g267)) + ((!g263) & (g264) & (g265) & (!g266) & (g273) & (g267)) + ((!g263) & (g264) & (g265) & (g266) & (g273) & (!g267)) + ((!g263) & (g264) & (g265) & (g266) & (g273) & (g267)) + ((g263) & (!g264) & (!g265) & (!g266) & (!g273) & (!g267)) + ((g263) & (!g264) & (!g265) & (g266) & (!g273) & (!g267)) + ((g263) & (!g264) & (!g265) & (g266) & (!g273) & (g267)) + ((g263) & (!g264) & (!g265) & (g266) & (g273) & (!g267)) + ((g263) & (!g264) & (g265) & (!g266) & (!g273) & (!g267)) + ((g263) & (!g264) & (g265) & (!g266) & (g273) & (g267)) + ((g263) & (!g264) & (g265) & (g266) & (g273) & (!g267)) + ((g263) & (g264) & (!g265) & (!g266) & (!g273) & (!g267)) + ((g263) & (g264) & (!g265) & (g266) & (!g273) & (!g267)) + ((g263) & (g264) & (!g265) & (g266) & (g273) & (!g267)) + ((g263) & (g264) & (!g265) & (g266) & (g273) & (g267)) + ((g263) & (g264) & (g265) & (g266) & (!g273) & (g267)) + ((g263) & (g264) & (g265) & (g266) & (g273) & (g267)));
	assign g282 = (((!g278) & (!g279) & (!g280) & (!g281) & (!g268) & (!g274)) + ((!g278) & (!g279) & (!g280) & (!g281) & (g268) & (!g274)) + ((!g278) & (!g279) & (!g280) & (g281) & (!g268) & (!g274)) + ((!g278) & (!g279) & (!g280) & (g281) & (g268) & (!g274)) + ((!g278) & (!g279) & (!g280) & (g281) & (g268) & (g274)) + ((!g278) & (!g279) & (g280) & (!g281) & (!g268) & (!g274)) + ((!g278) & (!g279) & (g280) & (!g281) & (!g268) & (g274)) + ((!g278) & (!g279) & (g280) & (!g281) & (g268) & (!g274)) + ((!g278) & (!g279) & (g280) & (g281) & (!g268) & (!g274)) + ((!g278) & (!g279) & (g280) & (g281) & (!g268) & (g274)) + ((!g278) & (!g279) & (g280) & (g281) & (g268) & (!g274)) + ((!g278) & (!g279) & (g280) & (g281) & (g268) & (g274)) + ((!g278) & (g279) & (!g280) & (!g281) & (!g268) & (!g274)) + ((!g278) & (g279) & (!g280) & (g281) & (!g268) & (!g274)) + ((!g278) & (g279) & (!g280) & (g281) & (g268) & (g274)) + ((!g278) & (g279) & (g280) & (!g281) & (!g268) & (!g274)) + ((!g278) & (g279) & (g280) & (!g281) & (!g268) & (g274)) + ((!g278) & (g279) & (g280) & (g281) & (!g268) & (!g274)) + ((!g278) & (g279) & (g280) & (g281) & (!g268) & (g274)) + ((!g278) & (g279) & (g280) & (g281) & (g268) & (g274)) + ((g278) & (!g279) & (!g280) & (!g281) & (g268) & (!g274)) + ((g278) & (!g279) & (!g280) & (g281) & (g268) & (!g274)) + ((g278) & (!g279) & (!g280) & (g281) & (g268) & (g274)) + ((g278) & (!g279) & (g280) & (!g281) & (!g268) & (g274)) + ((g278) & (!g279) & (g280) & (!g281) & (g268) & (!g274)) + ((g278) & (!g279) & (g280) & (g281) & (!g268) & (g274)) + ((g278) & (!g279) & (g280) & (g281) & (g268) & (!g274)) + ((g278) & (!g279) & (g280) & (g281) & (g268) & (g274)) + ((g278) & (g279) & (!g280) & (g281) & (g268) & (g274)) + ((g278) & (g279) & (g280) & (!g281) & (!g268) & (g274)) + ((g278) & (g279) & (g280) & (g281) & (!g268) & (g274)) + ((g278) & (g279) & (g280) & (g281) & (g268) & (g274)));
	assign g284 = (((!sk[108]) & (g282) & (!g283)) + ((!sk[108]) & (g282) & (g283)) + ((sk[108]) & (!g282) & (g283)) + ((sk[108]) & (g282) & (!g283)));
	assign g285 = (((!g267) & (!g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((!g267) & (!g264) & (!g265) & (!g266) & (g273) & (g268)) + ((!g267) & (!g264) & (!g265) & (g266) & (!g273) & (g268)) + ((!g267) & (!g264) & (!g265) & (g266) & (g273) & (!g268)) + ((!g267) & (!g264) & (!g265) & (g266) & (g273) & (g268)) + ((!g267) & (!g264) & (g265) & (!g266) & (!g273) & (g268)) + ((!g267) & (!g264) & (g265) & (g266) & (!g273) & (!g268)) + ((!g267) & (!g264) & (g265) & (g266) & (g273) & (!g268)) + ((!g267) & (g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((!g267) & (g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((!g267) & (g264) & (!g265) & (g266) & (!g273) & (g268)) + ((!g267) & (g264) & (g265) & (!g266) & (!g273) & (!g268)) + ((!g267) & (g264) & (g265) & (!g266) & (!g273) & (g268)) + ((!g267) & (g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g267) & (g264) & (g265) & (!g266) & (g273) & (g268)) + ((g267) & (!g264) & (!g265) & (g266) & (!g273) & (g268)) + ((g267) & (!g264) & (!g265) & (g266) & (g273) & (g268)) + ((g267) & (g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((g267) & (g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((g267) & (g264) & (!g265) & (g266) & (g273) & (!g268)) + ((g267) & (g264) & (g265) & (g266) & (!g273) & (!g268)) + ((g267) & (g264) & (g265) & (g266) & (!g273) & (g268)));
	assign g286 = (((!g267) & (!g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((!g267) & (!g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((!g267) & (!g264) & (!g265) & (g266) & (g273) & (g268)) + ((!g267) & (!g264) & (g265) & (!g266) & (!g273) & (!g268)) + ((!g267) & (!g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g267) & (!g264) & (g265) & (g266) & (!g273) & (g268)) + ((!g267) & (g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((!g267) & (g264) & (!g265) & (!g266) & (g273) & (g268)) + ((!g267) & (g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((!g267) & (g264) & (!g265) & (g266) & (!g273) & (g268)) + ((!g267) & (g264) & (!g265) & (g266) & (g273) & (g268)) + ((!g267) & (g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g267) & (g264) & (g265) & (!g266) & (g273) & (g268)) + ((!g267) & (g264) & (g265) & (g266) & (g273) & (!g268)) + ((g267) & (!g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((g267) & (!g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((g267) & (!g264) & (!g265) & (!g266) & (g273) & (g268)) + ((g267) & (!g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((g267) & (!g264) & (!g265) & (g266) & (!g273) & (g268)) + ((g267) & (!g264) & (!g265) & (g266) & (g273) & (!g268)) + ((g267) & (!g264) & (g265) & (g266) & (!g273) & (!g268)) + ((g267) & (g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((g267) & (g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((g267) & (g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((g267) & (g264) & (!g265) & (g266) & (g273) & (!g268)) + ((g267) & (g264) & (!g265) & (g266) & (g273) & (g268)) + ((g267) & (g264) & (g265) & (!g266) & (!g273) & (!g268)) + ((g267) & (g264) & (g265) & (!g266) & (g273) & (!g268)) + ((g267) & (g264) & (g265) & (g266) & (!g273) & (g268)) + ((g267) & (g264) & (g265) & (g266) & (g273) & (g268)));
	assign g287 = (((!g267) & (!g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((!g267) & (!g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((!g267) & (!g264) & (!g265) & (g266) & (!g273) & (g268)) + ((!g267) & (!g264) & (g265) & (!g266) & (!g273) & (g268)) + ((!g267) & (!g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g267) & (!g264) & (g265) & (g266) & (!g273) & (g268)) + ((!g267) & (g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((!g267) & (g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((!g267) & (g264) & (!g265) & (g266) & (g273) & (!g268)) + ((!g267) & (g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g267) & (g264) & (g265) & (g266) & (!g273) & (!g268)) + ((!g267) & (g264) & (g265) & (g266) & (g273) & (!g268)) + ((g267) & (!g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((g267) & (!g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((g267) & (!g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((g267) & (!g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((g267) & (!g264) & (!g265) & (g266) & (!g273) & (g268)) + ((g267) & (!g264) & (!g265) & (g266) & (g273) & (!g268)) + ((g267) & (!g264) & (!g265) & (g266) & (g273) & (g268)) + ((g267) & (!g264) & (g265) & (!g266) & (!g273) & (g268)) + ((g267) & (!g264) & (g265) & (!g266) & (g273) & (!g268)) + ((g267) & (!g264) & (g265) & (g266) & (!g273) & (!g268)) + ((g267) & (!g264) & (g265) & (g266) & (g273) & (g268)) + ((g267) & (g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((g267) & (g264) & (!g265) & (!g266) & (g273) & (g268)) + ((g267) & (g264) & (g265) & (!g266) & (g273) & (g268)) + ((g267) & (g264) & (g265) & (g266) & (!g273) & (!g268)) + ((g267) & (g264) & (g265) & (g266) & (!g273) & (g268)) + ((g267) & (g264) & (g265) & (g266) & (g273) & (g268)));
	assign g288 = (((!g267) & (!g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((!g267) & (!g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((!g267) & (!g264) & (!g265) & (!g266) & (g273) & (g268)) + ((!g267) & (!g264) & (!g265) & (g266) & (!g273) & (g268)) + ((!g267) & (!g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g267) & (!g264) & (g265) & (g266) & (g273) & (g268)) + ((!g267) & (g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((!g267) & (g264) & (!g265) & (g266) & (!g273) & (g268)) + ((!g267) & (g264) & (!g265) & (g266) & (g273) & (g268)) + ((!g267) & (g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g267) & (g264) & (g265) & (!g266) & (g273) & (g268)) + ((!g267) & (g264) & (g265) & (g266) & (!g273) & (!g268)) + ((!g267) & (g264) & (g265) & (g266) & (!g273) & (g268)) + ((!g267) & (g264) & (g265) & (g266) & (g273) & (!g268)) + ((!g267) & (g264) & (g265) & (g266) & (g273) & (g268)) + ((g267) & (!g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((g267) & (!g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((g267) & (!g264) & (!g265) & (!g266) & (g273) & (g268)) + ((g267) & (!g264) & (!g265) & (g266) & (g273) & (g268)) + ((g267) & (!g264) & (g265) & (!g266) & (!g273) & (g268)) + ((g267) & (!g264) & (g265) & (!g266) & (g273) & (!g268)) + ((g267) & (!g264) & (g265) & (g266) & (g273) & (!g268)) + ((g267) & (g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((g267) & (g264) & (!g265) & (g266) & (!g273) & (g268)) + ((g267) & (g264) & (!g265) & (g266) & (g273) & (!g268)) + ((g267) & (g264) & (g265) & (!g266) & (g273) & (g268)) + ((g267) & (g264) & (g265) & (g266) & (!g273) & (!g268)));
	assign g289 = (((!g285) & (!g286) & (!g287) & (!g288) & (!g263) & (g274)) + ((!g285) & (!g286) & (!g287) & (!g288) & (g263) & (!g274)) + ((!g285) & (!g286) & (!g287) & (!g288) & (g263) & (g274)) + ((!g285) & (!g286) & (!g287) & (g288) & (!g263) & (g274)) + ((!g285) & (!g286) & (!g287) & (g288) & (g263) & (!g274)) + ((!g285) & (!g286) & (g287) & (!g288) & (g263) & (!g274)) + ((!g285) & (!g286) & (g287) & (!g288) & (g263) & (g274)) + ((!g285) & (!g286) & (g287) & (g288) & (g263) & (!g274)) + ((!g285) & (g286) & (!g287) & (!g288) & (!g263) & (g274)) + ((!g285) & (g286) & (!g287) & (!g288) & (g263) & (g274)) + ((!g285) & (g286) & (!g287) & (g288) & (!g263) & (g274)) + ((!g285) & (g286) & (g287) & (!g288) & (g263) & (g274)) + ((g285) & (!g286) & (!g287) & (!g288) & (!g263) & (!g274)) + ((g285) & (!g286) & (!g287) & (!g288) & (!g263) & (g274)) + ((g285) & (!g286) & (!g287) & (!g288) & (g263) & (!g274)) + ((g285) & (!g286) & (!g287) & (!g288) & (g263) & (g274)) + ((g285) & (!g286) & (!g287) & (g288) & (!g263) & (!g274)) + ((g285) & (!g286) & (!g287) & (g288) & (!g263) & (g274)) + ((g285) & (!g286) & (!g287) & (g288) & (g263) & (!g274)) + ((g285) & (!g286) & (g287) & (!g288) & (!g263) & (!g274)) + ((g285) & (!g286) & (g287) & (!g288) & (g263) & (!g274)) + ((g285) & (!g286) & (g287) & (!g288) & (g263) & (g274)) + ((g285) & (!g286) & (g287) & (g288) & (!g263) & (!g274)) + ((g285) & (!g286) & (g287) & (g288) & (g263) & (!g274)) + ((g285) & (g286) & (!g287) & (!g288) & (!g263) & (!g274)) + ((g285) & (g286) & (!g287) & (!g288) & (!g263) & (g274)) + ((g285) & (g286) & (!g287) & (!g288) & (g263) & (g274)) + ((g285) & (g286) & (!g287) & (g288) & (!g263) & (!g274)) + ((g285) & (g286) & (!g287) & (g288) & (!g263) & (g274)) + ((g285) & (g286) & (g287) & (!g288) & (!g263) & (!g274)) + ((g285) & (g286) & (g287) & (!g288) & (g263) & (g274)) + ((g285) & (g286) & (g287) & (g288) & (!g263) & (!g274)));
	assign g291 = (((!sk[114]) & (g289) & (!g290)) + ((!sk[114]) & (g289) & (g290)) + ((sk[114]) & (!g289) & (g290)) + ((sk[114]) & (g289) & (!g290)));
	assign g292 = (((!g263) & (!g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (g273) & (g268)) + ((!g263) & (!g264) & (g265) & (g266) & (!g273) & (!g268)) + ((!g263) & (!g264) & (g265) & (g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (g265) & (g266) & (g273) & (g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (g264) & (g265) & (!g266) & (!g273) & (!g268)) + ((!g263) & (g264) & (g265) & (g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((g263) & (!g264) & (g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (g265) & (!g266) & (!g273) & (g268)) + ((g263) & (!g264) & (g265) & (!g266) & (g273) & (!g268)) + ((g263) & (!g264) & (g265) & (g266) & (!g273) & (g268)) + ((g263) & (g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((g263) & (g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((g263) & (g264) & (!g265) & (g266) & (g273) & (!g268)) + ((g263) & (g264) & (g265) & (!g266) & (!g273) & (g268)) + ((g263) & (g264) & (g265) & (!g266) & (g273) & (g268)));
	assign g293 = (((!g263) & (!g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (!g265) & (!g266) & (g273) & (g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (g265) & (g266) & (!g273) & (!g268)) + ((!g263) & (!g264) & (g265) & (g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (g265) & (g266) & (g273) & (g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (g273) & (g268)) + ((!g263) & (g264) & (!g265) & (g266) & (g273) & (g268)) + ((!g263) & (g264) & (g265) & (!g266) & (!g273) & (!g268)) + ((!g263) & (g264) & (g265) & (!g266) & (!g273) & (g268)) + ((!g263) & (g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (g264) & (g265) & (g266) & (!g273) & (g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((g263) & (!g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (!g265) & (g266) & (!g273) & (g268)) + ((g263) & (!g264) & (!g265) & (g266) & (g273) & (g268)) + ((g263) & (!g264) & (g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (g265) & (!g266) & (!g273) & (g268)) + ((g263) & (!g264) & (g265) & (!g266) & (g273) & (g268)) + ((g263) & (!g264) & (g265) & (g266) & (!g273) & (g268)) + ((g263) & (g264) & (!g265) & (g266) & (!g273) & (g268)) + ((g263) & (g264) & (!g265) & (g266) & (g273) & (!g268)) + ((g263) & (g264) & (g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (g264) & (g265) & (g266) & (!g273) & (!g268)));
	assign g294 = (((!g263) & (!g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (!g265) & (!g266) & (g273) & (g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (g265) & (!g266) & (g273) & (g268)) + ((!g263) & (!g264) & (g265) & (g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (g265) & (g266) & (g273) & (g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (g273) & (g268)) + ((!g263) & (g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((!g263) & (g264) & (!g265) & (g266) & (!g273) & (g268)) + ((!g263) & (g264) & (g265) & (!g266) & (!g273) & (g268)) + ((!g263) & (g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (g264) & (g265) & (g266) & (g273) & (g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (g273) & (g268)) + ((g263) & (!g264) & (!g265) & (g266) & (g273) & (g268)) + ((g263) & (!g264) & (g265) & (g266) & (!g273) & (!g268)) + ((g263) & (g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((g263) & (g264) & (!g265) & (g266) & (g273) & (g268)) + ((g263) & (g264) & (g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (g264) & (g265) & (!g266) & (!g273) & (g268)) + ((g263) & (g264) & (g265) & (!g266) & (g273) & (g268)) + ((g263) & (g264) & (g265) & (g266) & (!g273) & (!g268)) + ((g263) & (g264) & (g265) & (g266) & (g273) & (g268)));
	assign g295 = (((!g263) & (!g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (!g265) & (g266) & (g273) & (g268)) + ((!g263) & (!g264) & (g265) & (g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (g265) & (g266) & (g273) & (g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (!g273) & (!g268)) + ((!g263) & (g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (g264) & (!g265) & (g266) & (!g273) & (!g268)) + ((!g263) & (g264) & (!g265) & (g266) & (!g273) & (g268)) + ((!g263) & (g264) & (!g265) & (g266) & (g273) & (!g268)) + ((!g263) & (g264) & (g265) & (!g266) & (!g273) & (!g268)) + ((!g263) & (g264) & (g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (g264) & (g265) & (!g266) & (g273) & (g268)) + ((g263) & (!g264) & (!g265) & (!g266) & (g273) & (g268)) + ((g263) & (!g264) & (!g265) & (g266) & (g273) & (!g268)) + ((g263) & (!g264) & (g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (g265) & (!g266) & (g273) & (!g268)) + ((g263) & (!g264) & (g265) & (!g266) & (g273) & (g268)) + ((g263) & (!g264) & (g265) & (g266) & (!g273) & (g268)) + ((g263) & (!g264) & (g265) & (g266) & (g273) & (!g268)) + ((g263) & (!g264) & (g265) & (g266) & (g273) & (g268)) + ((g263) & (g264) & (!g265) & (!g266) & (!g273) & (g268)) + ((g263) & (g264) & (!g265) & (!g266) & (g273) & (!g268)) + ((g263) & (g264) & (g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (g264) & (g265) & (!g266) & (!g273) & (g268)) + ((g263) & (g264) & (g265) & (g266) & (g273) & (g268)));
	assign g296 = (((!g292) & (!g293) & (!g294) & (!g295) & (!g274) & (g267)) + ((!g292) & (!g293) & (!g294) & (!g295) & (g274) & (!g267)) + ((!g292) & (!g293) & (!g294) & (!g295) & (g274) & (g267)) + ((!g292) & (!g293) & (!g294) & (g295) & (!g274) & (g267)) + ((!g292) & (!g293) & (!g294) & (g295) & (g274) & (!g267)) + ((!g292) & (!g293) & (g294) & (!g295) & (g274) & (!g267)) + ((!g292) & (!g293) & (g294) & (!g295) & (g274) & (g267)) + ((!g292) & (!g293) & (g294) & (g295) & (g274) & (!g267)) + ((!g292) & (g293) & (!g294) & (!g295) & (!g274) & (g267)) + ((!g292) & (g293) & (!g294) & (!g295) & (g274) & (g267)) + ((!g292) & (g293) & (!g294) & (g295) & (!g274) & (g267)) + ((!g292) & (g293) & (g294) & (!g295) & (g274) & (g267)) + ((g292) & (!g293) & (!g294) & (!g295) & (!g274) & (!g267)) + ((g292) & (!g293) & (!g294) & (!g295) & (!g274) & (g267)) + ((g292) & (!g293) & (!g294) & (!g295) & (g274) & (!g267)) + ((g292) & (!g293) & (!g294) & (!g295) & (g274) & (g267)) + ((g292) & (!g293) & (!g294) & (g295) & (!g274) & (!g267)) + ((g292) & (!g293) & (!g294) & (g295) & (!g274) & (g267)) + ((g292) & (!g293) & (!g294) & (g295) & (g274) & (!g267)) + ((g292) & (!g293) & (g294) & (!g295) & (!g274) & (!g267)) + ((g292) & (!g293) & (g294) & (!g295) & (g274) & (!g267)) + ((g292) & (!g293) & (g294) & (!g295) & (g274) & (g267)) + ((g292) & (!g293) & (g294) & (g295) & (!g274) & (!g267)) + ((g292) & (!g293) & (g294) & (g295) & (g274) & (!g267)) + ((g292) & (g293) & (!g294) & (!g295) & (!g274) & (!g267)) + ((g292) & (g293) & (!g294) & (!g295) & (!g274) & (g267)) + ((g292) & (g293) & (!g294) & (!g295) & (g274) & (g267)) + ((g292) & (g293) & (!g294) & (g295) & (!g274) & (!g267)) + ((g292) & (g293) & (!g294) & (g295) & (!g274) & (g267)) + ((g292) & (g293) & (g294) & (!g295) & (!g274) & (!g267)) + ((g292) & (g293) & (g294) & (!g295) & (g274) & (g267)) + ((g292) & (g293) & (g294) & (g295) & (!g274) & (!g267)));
	assign g298 = (((!sk[120]) & (g296) & (!g297)) + ((!sk[120]) & (g296) & (g297)) + ((sk[120]) & (!g296) & (g297)) + ((sk[120]) & (g296) & (!g297)));
	assign g299 = (((!g263) & (!g264) & (!g267) & (!g274) & (!g273) & (g268)) + ((!g263) & (!g264) & (g267) & (!g274) & (!g273) & (g268)) + ((!g263) & (!g264) & (g267) & (!g274) & (g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (!g274) & (g273) & (g268)) + ((!g263) & (!g264) & (g267) & (g274) & (!g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (g274) & (g273) & (!g268)) + ((!g263) & (g264) & (!g267) & (!g274) & (!g273) & (!g268)) + ((!g263) & (g264) & (!g267) & (!g274) & (!g273) & (g268)) + ((!g263) & (g264) & (!g267) & (g274) & (!g273) & (!g268)) + ((!g263) & (g264) & (!g267) & (g274) & (!g273) & (g268)) + ((!g263) & (g264) & (!g267) & (g274) & (g273) & (g268)) + ((!g263) & (g264) & (g267) & (g274) & (!g273) & (g268)) + ((!g263) & (g264) & (g267) & (g274) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g274) & (!g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g274) & (!g273) & (g268)) + ((g263) & (!g264) & (!g267) & (g274) & (!g273) & (g268)) + ((g263) & (!g264) & (g267) & (!g274) & (g273) & (!g268)) + ((g263) & (!g264) & (g267) & (g274) & (!g273) & (!g268)) + ((g263) & (!g264) & (g267) & (g274) & (!g273) & (g268)) + ((g263) & (!g264) & (g267) & (g274) & (g273) & (!g268)) + ((g263) & (g264) & (!g267) & (!g274) & (!g273) & (!g268)) + ((g263) & (g264) & (!g267) & (!g274) & (g273) & (!g268)) + ((g263) & (g264) & (!g267) & (g274) & (g273) & (!g268)) + ((g263) & (g264) & (g267) & (!g274) & (!g273) & (!g268)) + ((g263) & (g264) & (g267) & (!g274) & (!g273) & (g268)) + ((g263) & (g264) & (g267) & (g274) & (!g273) & (g268)));
	assign g300 = (((!g263) & (!g264) & (!g267) & (!g274) & (!g273) & (!g268)) + ((!g263) & (!g264) & (!g267) & (!g274) & (!g273) & (g268)) + ((!g263) & (!g264) & (!g267) & (!g274) & (g273) & (!g268)) + ((!g263) & (!g264) & (!g267) & (!g274) & (g273) & (g268)) + ((!g263) & (!g264) & (!g267) & (g274) & (!g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (!g274) & (!g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (!g274) & (g273) & (g268)) + ((!g263) & (!g264) & (g267) & (g274) & (!g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (g274) & (g273) & (g268)) + ((!g263) & (g264) & (!g267) & (!g274) & (!g273) & (g268)) + ((!g263) & (g264) & (!g267) & (g274) & (g273) & (!g268)) + ((!g263) & (g264) & (g267) & (!g274) & (!g273) & (!g268)) + ((!g263) & (g264) & (g267) & (!g274) & (!g273) & (g268)) + ((!g263) & (g264) & (g267) & (!g274) & (g273) & (!g268)) + ((!g263) & (g264) & (g267) & (!g274) & (g273) & (g268)) + ((!g263) & (g264) & (g267) & (g274) & (!g273) & (!g268)) + ((!g263) & (g264) & (g267) & (g274) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g274) & (!g273) & (g268)) + ((g263) & (!g264) & (!g267) & (!g274) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g274) & (g273) & (g268)) + ((g263) & (!g264) & (!g267) & (g274) & (!g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (g274) & (g273) & (g268)) + ((g263) & (!g264) & (g267) & (!g274) & (g273) & (!g268)) + ((g263) & (!g264) & (g267) & (!g274) & (g273) & (g268)) + ((g263) & (!g264) & (g267) & (g274) & (!g273) & (g268)) + ((g263) & (g264) & (!g267) & (!g274) & (g273) & (!g268)) + ((g263) & (g264) & (!g267) & (!g274) & (g273) & (g268)) + ((g263) & (g264) & (!g267) & (g274) & (!g273) & (!g268)) + ((g263) & (g264) & (!g267) & (g274) & (!g273) & (g268)) + ((g263) & (g264) & (g267) & (!g274) & (g273) & (!g268)) + ((g263) & (g264) & (g267) & (!g274) & (g273) & (g268)) + ((g263) & (g264) & (g267) & (g274) & (!g273) & (g268)));
	assign g301 = (((!g263) & (!g264) & (!g267) & (!g274) & (!g273) & (!g268)) + ((!g263) & (!g264) & (!g267) & (!g274) & (!g273) & (g268)) + ((!g263) & (!g264) & (g267) & (!g274) & (!g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (!g274) & (g273) & (g268)) + ((!g263) & (!g264) & (g267) & (g274) & (!g273) & (g268)) + ((!g263) & (g264) & (!g267) & (g274) & (!g273) & (!g268)) + ((!g263) & (g264) & (!g267) & (g274) & (g273) & (!g268)) + ((!g263) & (g264) & (!g267) & (g274) & (g273) & (g268)) + ((!g263) & (g264) & (g267) & (!g274) & (!g273) & (!g268)) + ((!g263) & (g264) & (g267) & (!g274) & (g273) & (!g268)) + ((!g263) & (g264) & (g267) & (!g274) & (g273) & (g268)) + ((!g263) & (g264) & (g267) & (g274) & (!g273) & (!g268)) + ((!g263) & (g264) & (g267) & (g274) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g274) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g274) & (g273) & (g268)) + ((g263) & (!g264) & (!g267) & (g274) & (!g273) & (g268)) + ((g263) & (!g264) & (!g267) & (g274) & (g273) & (g268)) + ((g263) & (!g264) & (g267) & (!g274) & (!g273) & (!g268)) + ((g263) & (!g264) & (g267) & (!g274) & (!g273) & (g268)) + ((g263) & (!g264) & (g267) & (!g274) & (g273) & (g268)) + ((g263) & (!g264) & (g267) & (g274) & (!g273) & (!g268)) + ((g263) & (!g264) & (g267) & (g274) & (!g273) & (g268)) + ((g263) & (!g264) & (g267) & (g274) & (g273) & (!g268)) + ((g263) & (!g264) & (g267) & (g274) & (g273) & (g268)) + ((g263) & (g264) & (!g267) & (!g274) & (!g273) & (g268)) + ((g263) & (g264) & (!g267) & (g274) & (!g273) & (!g268)) + ((g263) & (g264) & (!g267) & (g274) & (g273) & (!g268)) + ((g263) & (g264) & (g267) & (!g274) & (!g273) & (!g268)) + ((g263) & (g264) & (g267) & (!g274) & (!g273) & (g268)) + ((g263) & (g264) & (g267) & (!g274) & (g273) & (!g268)) + ((g263) & (g264) & (g267) & (g274) & (!g273) & (!g268)) + ((g263) & (g264) & (g267) & (g274) & (g273) & (!g268)));
	assign g302 = (((!g263) & (!g264) & (!g267) & (!g274) & (g273) & (g268)) + ((!g263) & (!g264) & (!g267) & (g274) & (!g273) & (!g268)) + ((!g263) & (!g264) & (!g267) & (g274) & (g273) & (g268)) + ((!g263) & (!g264) & (g267) & (!g274) & (!g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (!g274) & (g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (g274) & (!g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (g274) & (!g273) & (g268)) + ((!g263) & (!g264) & (g267) & (g274) & (g273) & (!g268)) + ((!g263) & (g264) & (!g267) & (!g274) & (!g273) & (!g268)) + ((!g263) & (g264) & (!g267) & (g274) & (!g273) & (g268)) + ((!g263) & (g264) & (!g267) & (g274) & (g273) & (!g268)) + ((!g263) & (g264) & (!g267) & (g274) & (g273) & (g268)) + ((!g263) & (g264) & (g267) & (!g274) & (!g273) & (!g268)) + ((!g263) & (g264) & (g267) & (g274) & (!g273) & (!g268)) + ((!g263) & (g264) & (g267) & (g274) & (!g273) & (g268)) + ((g263) & (!g264) & (!g267) & (!g274) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g274) & (g273) & (g268)) + ((g263) & (!g264) & (g267) & (!g274) & (!g273) & (!g268)) + ((g263) & (!g264) & (g267) & (!g274) & (g273) & (!g268)) + ((g263) & (!g264) & (g267) & (g274) & (g273) & (!g268)) + ((g263) & (g264) & (!g267) & (!g274) & (g273) & (!g268)) + ((g263) & (g264) & (!g267) & (g274) & (g273) & (g268)) + ((g263) & (g264) & (g267) & (!g274) & (!g273) & (!g268)) + ((g263) & (g264) & (g267) & (!g274) & (!g273) & (g268)) + ((g263) & (g264) & (g267) & (!g274) & (g273) & (!g268)) + ((g263) & (g264) & (g267) & (g274) & (!g273) & (!g268)));
	assign g303 = (((!g299) & (!g300) & (!g301) & (!g302) & (g265) & (g266)) + ((!g299) & (!g300) & (g301) & (!g302) & (!g265) & (g266)) + ((!g299) & (!g300) & (g301) & (!g302) & (g265) & (g266)) + ((!g299) & (!g300) & (g301) & (g302) & (!g265) & (g266)) + ((!g299) & (g300) & (!g301) & (!g302) & (g265) & (!g266)) + ((!g299) & (g300) & (!g301) & (!g302) & (g265) & (g266)) + ((!g299) & (g300) & (!g301) & (g302) & (g265) & (!g266)) + ((!g299) & (g300) & (g301) & (!g302) & (!g265) & (g266)) + ((!g299) & (g300) & (g301) & (!g302) & (g265) & (!g266)) + ((!g299) & (g300) & (g301) & (!g302) & (g265) & (g266)) + ((!g299) & (g300) & (g301) & (g302) & (!g265) & (g266)) + ((!g299) & (g300) & (g301) & (g302) & (g265) & (!g266)) + ((g299) & (!g300) & (!g301) & (!g302) & (!g265) & (!g266)) + ((g299) & (!g300) & (!g301) & (!g302) & (g265) & (g266)) + ((g299) & (!g300) & (!g301) & (g302) & (!g265) & (!g266)) + ((g299) & (!g300) & (g301) & (!g302) & (!g265) & (!g266)) + ((g299) & (!g300) & (g301) & (!g302) & (!g265) & (g266)) + ((g299) & (!g300) & (g301) & (!g302) & (g265) & (g266)) + ((g299) & (!g300) & (g301) & (g302) & (!g265) & (!g266)) + ((g299) & (!g300) & (g301) & (g302) & (!g265) & (g266)) + ((g299) & (g300) & (!g301) & (!g302) & (!g265) & (!g266)) + ((g299) & (g300) & (!g301) & (!g302) & (g265) & (!g266)) + ((g299) & (g300) & (!g301) & (!g302) & (g265) & (g266)) + ((g299) & (g300) & (!g301) & (g302) & (!g265) & (!g266)) + ((g299) & (g300) & (!g301) & (g302) & (g265) & (!g266)) + ((g299) & (g300) & (g301) & (!g302) & (!g265) & (!g266)) + ((g299) & (g300) & (g301) & (!g302) & (!g265) & (g266)) + ((g299) & (g300) & (g301) & (!g302) & (g265) & (!g266)) + ((g299) & (g300) & (g301) & (!g302) & (g265) & (g266)) + ((g299) & (g300) & (g301) & (g302) & (!g265) & (!g266)) + ((g299) & (g300) & (g301) & (g302) & (!g265) & (g266)) + ((g299) & (g300) & (g301) & (g302) & (g265) & (!g266)));
	assign g305 = (((!sk[126]) & (g303) & (!g304)) + ((!sk[126]) & (g303) & (g304)) + ((sk[126]) & (!g303) & (g304)) + ((sk[126]) & (g303) & (!g304)));
	assign g306 = (((!g263) & (!g264) & (!g267) & (!g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (!g267) & (!g266) & (g273) & (g268)) + ((!g263) & (!g264) & (!g267) & (g266) & (g273) & (g268)) + ((!g263) & (!g264) & (g267) & (!g266) & (!g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (!g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (g267) & (!g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (!g266) & (g273) & (g268)) + ((!g263) & (!g264) & (g267) & (g266) & (!g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (g266) & (!g273) & (g268)) + ((!g263) & (g264) & (!g267) & (!g266) & (!g273) & (g268)) + ((!g263) & (g264) & (!g267) & (!g266) & (g273) & (!g268)) + ((!g263) & (g264) & (!g267) & (g266) & (g273) & (g268)) + ((!g263) & (g264) & (g267) & (!g266) & (g273) & (!g268)) + ((!g263) & (g264) & (g267) & (!g266) & (g273) & (g268)) + ((!g263) & (g264) & (g267) & (g266) & (!g273) & (!g268)) + ((!g263) & (g264) & (g267) & (g266) & (!g273) & (g268)) + ((!g263) & (g264) & (g267) & (g266) & (g273) & (g268)) + ((g263) & (!g264) & (!g267) & (!g266) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g266) & (g273) & (g268)) + ((g263) & (!g264) & (!g267) & (g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (g266) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (g266) & (g273) & (g268)) + ((g263) & (!g264) & (g267) & (!g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (g267) & (!g266) & (g273) & (!g268)) + ((g263) & (!g264) & (g267) & (g266) & (g273) & (!g268)) + ((g263) & (g264) & (!g267) & (!g266) & (g273) & (g268)) + ((g263) & (g264) & (g267) & (!g266) & (!g273) & (!g268)) + ((g263) & (g264) & (g267) & (!g266) & (g273) & (g268)));
	assign g307 = (((!g263) & (!g264) & (!g267) & (!g266) & (!g273) & (!g268)) + ((!g263) & (!g264) & (!g267) & (g266) & (!g273) & (!g268)) + ((!g263) & (!g264) & (!g267) & (g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (!g267) & (g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (!g266) & (g273) & (g268)) + ((!g263) & (!g264) & (g267) & (g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (g267) & (g266) & (g273) & (g268)) + ((!g263) & (g264) & (!g267) & (!g266) & (!g273) & (!g268)) + ((!g263) & (g264) & (!g267) & (!g266) & (g273) & (!g268)) + ((!g263) & (g264) & (g267) & (!g266) & (!g273) & (g268)) + ((!g263) & (g264) & (g267) & (!g266) & (g273) & (g268)) + ((!g263) & (g264) & (g267) & (g266) & (!g273) & (g268)) + ((!g263) & (g264) & (g267) & (g266) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g266) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g266) & (g273) & (g268)) + ((g263) & (!g264) & (!g267) & (g266) & (!g273) & (g268)) + ((g263) & (!g264) & (!g267) & (g266) & (g273) & (g268)) + ((g263) & (!g264) & (g267) & (g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (g267) & (g266) & (!g273) & (g268)) + ((g263) & (!g264) & (g267) & (g266) & (g273) & (g268)) + ((g263) & (g264) & (!g267) & (!g266) & (!g273) & (g268)) + ((g263) & (g264) & (!g267) & (!g266) & (g273) & (!g268)) + ((g263) & (g264) & (!g267) & (g266) & (g273) & (!g268)) + ((g263) & (g264) & (g267) & (!g266) & (!g273) & (g268)) + ((g263) & (g264) & (g267) & (!g266) & (g273) & (g268)) + ((g263) & (g264) & (g267) & (g266) & (!g273) & (!g268)) + ((g263) & (g264) & (g267) & (g266) & (g273) & (g268)));
	assign g308 = (((!g263) & (!g264) & (!g267) & (!g266) & (g273) & (g268)) + ((!g263) & (!g264) & (!g267) & (g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (!g266) & (!g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (!g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (g267) & (!g266) & (g273) & (g268)) + ((!g263) & (!g264) & (g267) & (g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (g267) & (g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (g267) & (g266) & (g273) & (g268)) + ((!g263) & (g264) & (!g267) & (!g266) & (g273) & (!g268)) + ((!g263) & (g264) & (!g267) & (!g266) & (g273) & (g268)) + ((!g263) & (g264) & (g267) & (!g266) & (!g273) & (!g268)) + ((!g263) & (g264) & (g267) & (g266) & (!g273) & (g268)) + ((!g263) & (g264) & (g267) & (g266) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g266) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (!g266) & (g273) & (g268)) + ((g263) & (!g264) & (!g267) & (g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (g266) & (!g273) & (g268)) + ((g263) & (!g264) & (g267) & (!g266) & (!g273) & (g268)) + ((g263) & (!g264) & (g267) & (!g266) & (g273) & (g268)) + ((g263) & (!g264) & (g267) & (g266) & (g273) & (!g268)) + ((g263) & (g264) & (!g267) & (!g266) & (!g273) & (!g268)) + ((g263) & (g264) & (!g267) & (!g266) & (!g273) & (g268)) + ((g263) & (g264) & (!g267) & (!g266) & (g273) & (g268)) + ((g263) & (g264) & (!g267) & (g266) & (!g273) & (g268)) + ((g263) & (g264) & (!g267) & (g266) & (g273) & (!g268)) + ((g263) & (g264) & (g267) & (!g266) & (!g273) & (g268)) + ((g263) & (g264) & (g267) & (!g266) & (g273) & (!g268)) + ((g263) & (g264) & (g267) & (g266) & (!g273) & (!g268)) + ((g263) & (g264) & (g267) & (g266) & (g273) & (!g268)) + ((g263) & (g264) & (g267) & (g266) & (g273) & (g268)));
	assign g309 = (((!g263) & (!g264) & (!g267) & (!g266) & (g273) & (!g268)) + ((!g263) & (!g264) & (!g267) & (g266) & (!g273) & (!g268)) + ((!g263) & (!g264) & (!g267) & (g266) & (g273) & (g268)) + ((!g263) & (!g264) & (g267) & (!g266) & (!g273) & (g268)) + ((!g263) & (!g264) & (g267) & (!g266) & (g273) & (g268)) + ((!g263) & (!g264) & (g267) & (g266) & (g273) & (g268)) + ((!g263) & (g264) & (!g267) & (!g266) & (!g273) & (g268)) + ((!g263) & (g264) & (!g267) & (g266) & (!g273) & (g268)) + ((!g263) & (g264) & (!g267) & (g266) & (g273) & (g268)) + ((!g263) & (g264) & (g267) & (!g266) & (!g273) & (!g268)) + ((!g263) & (g264) & (g267) & (!g266) & (g273) & (!g268)) + ((!g263) & (g264) & (g267) & (g266) & (!g273) & (g268)) + ((!g263) & (g264) & (g267) & (g266) & (g273) & (g268)) + ((g263) & (!g264) & (!g267) & (!g266) & (g273) & (!g268)) + ((g263) & (!g264) & (!g267) & (g266) & (g273) & (g268)) + ((g263) & (!g264) & (g267) & (!g266) & (!g273) & (!g268)) + ((g263) & (!g264) & (g267) & (!g266) & (g273) & (g268)) + ((g263) & (!g264) & (g267) & (g266) & (!g273) & (!g268)) + ((g263) & (g264) & (!g267) & (!g266) & (g273) & (g268)) + ((g263) & (g264) & (!g267) & (g266) & (!g273) & (!g268)) + ((g263) & (g264) & (!g267) & (g266) & (!g273) & (g268)) + ((g263) & (g264) & (g267) & (!g266) & (g273) & (g268)));
	assign g310 = (((!g306) & (!g307) & (!g308) & (!g309) & (!g274) & (!g265)) + ((!g306) & (!g307) & (!g308) & (!g309) & (!g274) & (g265)) + ((!g306) & (!g307) & (!g308) & (!g309) & (g274) & (!g265)) + ((!g306) & (!g307) & (!g308) & (g309) & (!g274) & (!g265)) + ((!g306) & (!g307) & (!g308) & (g309) & (!g274) & (g265)) + ((!g306) & (!g307) & (!g308) & (g309) & (g274) & (!g265)) + ((!g306) & (!g307) & (!g308) & (g309) & (g274) & (g265)) + ((!g306) & (!g307) & (g308) & (!g309) & (!g274) & (!g265)) + ((!g306) & (!g307) & (g308) & (!g309) & (g274) & (!g265)) + ((!g306) & (!g307) & (g308) & (g309) & (!g274) & (!g265)) + ((!g306) & (!g307) & (g308) & (g309) & (g274) & (!g265)) + ((!g306) & (!g307) & (g308) & (g309) & (g274) & (g265)) + ((!g306) & (g307) & (!g308) & (!g309) & (!g274) & (!g265)) + ((!g306) & (g307) & (!g308) & (!g309) & (!g274) & (g265)) + ((!g306) & (g307) & (!g308) & (g309) & (!g274) & (!g265)) + ((!g306) & (g307) & (!g308) & (g309) & (!g274) & (g265)) + ((!g306) & (g307) & (!g308) & (g309) & (g274) & (g265)) + ((!g306) & (g307) & (g308) & (!g309) & (!g274) & (!g265)) + ((!g306) & (g307) & (g308) & (g309) & (!g274) & (!g265)) + ((!g306) & (g307) & (g308) & (g309) & (g274) & (g265)) + ((g306) & (!g307) & (!g308) & (!g309) & (!g274) & (g265)) + ((g306) & (!g307) & (!g308) & (!g309) & (g274) & (!g265)) + ((g306) & (!g307) & (!g308) & (g309) & (!g274) & (g265)) + ((g306) & (!g307) & (!g308) & (g309) & (g274) & (!g265)) + ((g306) & (!g307) & (!g308) & (g309) & (g274) & (g265)) + ((g306) & (!g307) & (g308) & (!g309) & (g274) & (!g265)) + ((g306) & (!g307) & (g308) & (g309) & (g274) & (!g265)) + ((g306) & (!g307) & (g308) & (g309) & (g274) & (g265)) + ((g306) & (g307) & (!g308) & (!g309) & (!g274) & (g265)) + ((g306) & (g307) & (!g308) & (g309) & (!g274) & (g265)) + ((g306) & (g307) & (!g308) & (g309) & (g274) & (g265)) + ((g306) & (g307) & (g308) & (g309) & (g274) & (g265)));
	assign g312 = (((!g310) & (sk[4]) & (g311)) + ((g310) & (!sk[4]) & (!g311)) + ((g310) & (!sk[4]) & (g311)) + ((g310) & (sk[4]) & (!g311)));
	assign g313 = (((!g263) & (!g274) & (!g265) & (!g266) & (!g273) & (g268)) + ((!g263) & (!g274) & (!g265) & (!g266) & (g273) & (g268)) + ((!g263) & (!g274) & (!g265) & (g266) & (!g273) & (!g268)) + ((!g263) & (!g274) & (!g265) & (g266) & (!g273) & (g268)) + ((!g263) & (!g274) & (!g265) & (g266) & (g273) & (!g268)) + ((!g263) & (!g274) & (!g265) & (g266) & (g273) & (g268)) + ((!g263) & (!g274) & (g265) & (!g266) & (!g273) & (g268)) + ((!g263) & (!g274) & (g265) & (!g266) & (g273) & (g268)) + ((!g263) & (!g274) & (g265) & (g266) & (g273) & (!g268)) + ((!g263) & (g274) & (g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (g274) & (g265) & (!g266) & (g273) & (g268)) + ((!g263) & (g274) & (g265) & (g266) & (!g273) & (g268)) + ((g263) & (!g274) & (!g265) & (!g266) & (g273) & (!g268)) + ((g263) & (!g274) & (!g265) & (g266) & (!g273) & (!g268)) + ((g263) & (!g274) & (!g265) & (g266) & (!g273) & (g268)) + ((g263) & (!g274) & (!g265) & (g266) & (g273) & (g268)) + ((g263) & (!g274) & (g265) & (!g266) & (!g273) & (g268)) + ((g263) & (!g274) & (g265) & (!g266) & (g273) & (g268)) + ((g263) & (!g274) & (g265) & (g266) & (g273) & (!g268)) + ((g263) & (!g274) & (g265) & (g266) & (g273) & (g268)) + ((g263) & (g274) & (!g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (g274) & (!g265) & (!g266) & (!g273) & (g268)) + ((g263) & (g274) & (!g265) & (!g266) & (g273) & (!g268)) + ((g263) & (g274) & (!g265) & (g266) & (!g273) & (!g268)) + ((g263) & (g274) & (g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (g274) & (g265) & (!g266) & (!g273) & (g268)) + ((g263) & (g274) & (g265) & (!g266) & (g273) & (!g268)) + ((g263) & (g274) & (g265) & (g266) & (!g273) & (g268)));
	assign g314 = (((!g263) & (!g274) & (!g265) & (!g266) & (!g273) & (!g268)) + ((!g263) & (!g274) & (!g265) & (g266) & (g273) & (g268)) + ((!g263) & (!g274) & (g265) & (!g266) & (!g273) & (!g268)) + ((!g263) & (!g274) & (g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (!g274) & (g265) & (!g266) & (g273) & (g268)) + ((!g263) & (!g274) & (g265) & (g266) & (!g273) & (!g268)) + ((!g263) & (!g274) & (g265) & (g266) & (g273) & (g268)) + ((!g263) & (g274) & (!g265) & (!g266) & (!g273) & (!g268)) + ((!g263) & (g274) & (!g265) & (!g266) & (g273) & (g268)) + ((!g263) & (g274) & (!g265) & (g266) & (!g273) & (g268)) + ((!g263) & (g274) & (g265) & (!g266) & (!g273) & (!g268)) + ((!g263) & (g274) & (g265) & (!g266) & (g273) & (g268)) + ((!g263) & (g274) & (g265) & (g266) & (g273) & (!g268)) + ((!g263) & (g274) & (g265) & (g266) & (g273) & (g268)) + ((g263) & (!g274) & (!g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (!g274) & (!g265) & (!g266) & (g273) & (g268)) + ((g263) & (!g274) & (!g265) & (g266) & (!g273) & (!g268)) + ((g263) & (!g274) & (!g265) & (g266) & (g273) & (g268)) + ((g263) & (!g274) & (g265) & (!g266) & (g273) & (g268)) + ((g263) & (!g274) & (g265) & (g266) & (!g273) & (g268)) + ((g263) & (g274) & (!g265) & (!g266) & (g273) & (!g268)) + ((g263) & (g274) & (!g265) & (!g266) & (g273) & (g268)) + ((g263) & (g274) & (!g265) & (g266) & (!g273) & (g268)) + ((g263) & (g274) & (!g265) & (g266) & (g273) & (!g268)) + ((g263) & (g274) & (!g265) & (g266) & (g273) & (g268)) + ((g263) & (g274) & (g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (g274) & (g265) & (!g266) & (g273) & (!g268)) + ((g263) & (g274) & (g265) & (g266) & (!g273) & (!g268)));
	assign g315 = (((!g263) & (!g274) & (!g265) & (!g266) & (!g273) & (g268)) + ((!g263) & (!g274) & (!g265) & (!g266) & (g273) & (g268)) + ((!g263) & (!g274) & (!g265) & (g266) & (g273) & (!g268)) + ((!g263) & (!g274) & (!g265) & (g266) & (g273) & (g268)) + ((!g263) & (!g274) & (g265) & (!g266) & (g273) & (g268)) + ((!g263) & (!g274) & (g265) & (g266) & (!g273) & (!g268)) + ((!g263) & (!g274) & (g265) & (g266) & (!g273) & (g268)) + ((!g263) & (!g274) & (g265) & (g266) & (g273) & (g268)) + ((!g263) & (g274) & (!g265) & (!g266) & (!g273) & (!g268)) + ((!g263) & (g274) & (!g265) & (!g266) & (!g273) & (g268)) + ((!g263) & (g274) & (!g265) & (!g266) & (g273) & (g268)) + ((!g263) & (g274) & (!g265) & (g266) & (!g273) & (g268)) + ((!g263) & (g274) & (!g265) & (g266) & (g273) & (!g268)) + ((!g263) & (g274) & (g265) & (!g266) & (!g273) & (g268)) + ((!g263) & (g274) & (g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (g274) & (g265) & (g266) & (!g273) & (!g268)) + ((!g263) & (g274) & (g265) & (g266) & (g273) & (!g268)) + ((!g263) & (g274) & (g265) & (g266) & (g273) & (g268)) + ((g263) & (!g274) & (!g265) & (!g266) & (!g273) & (g268)) + ((g263) & (!g274) & (!g265) & (g266) & (!g273) & (!g268)) + ((g263) & (!g274) & (!g265) & (g266) & (g273) & (!g268)) + ((g263) & (!g274) & (g265) & (!g266) & (g273) & (g268)) + ((g263) & (!g274) & (g265) & (g266) & (!g273) & (g268)) + ((g263) & (g274) & (!g265) & (!g266) & (!g273) & (g268)) + ((g263) & (g274) & (!g265) & (g266) & (!g273) & (!g268)) + ((g263) & (g274) & (!g265) & (g266) & (g273) & (!g268)) + ((g263) & (g274) & (g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (g274) & (g265) & (!g266) & (g273) & (!g268)) + ((g263) & (g274) & (g265) & (!g266) & (g273) & (g268)) + ((g263) & (g274) & (g265) & (g266) & (g273) & (g268)));
	assign g316 = (((!g263) & (!g274) & (!g265) & (!g266) & (g273) & (g268)) + ((!g263) & (!g274) & (!g265) & (g266) & (!g273) & (!g268)) + ((!g263) & (!g274) & (!g265) & (g266) & (g273) & (g268)) + ((!g263) & (!g274) & (g265) & (!g266) & (!g273) & (!g268)) + ((!g263) & (!g274) & (g265) & (g266) & (g273) & (!g268)) + ((!g263) & (!g274) & (g265) & (g266) & (g273) & (g268)) + ((!g263) & (g274) & (!g265) & (g266) & (!g273) & (!g268)) + ((!g263) & (g274) & (!g265) & (g266) & (g273) & (!g268)) + ((!g263) & (g274) & (g265) & (!g266) & (g273) & (!g268)) + ((!g263) & (g274) & (g265) & (!g266) & (g273) & (g268)) + ((g263) & (!g274) & (!g265) & (!g266) & (!g273) & (g268)) + ((g263) & (!g274) & (!g265) & (!g266) & (g273) & (!g268)) + ((g263) & (!g274) & (!g265) & (g266) & (!g273) & (g268)) + ((g263) & (!g274) & (g265) & (!g266) & (g273) & (!g268)) + ((g263) & (!g274) & (g265) & (!g266) & (g273) & (g268)) + ((g263) & (!g274) & (g265) & (g266) & (g273) & (!g268)) + ((g263) & (!g274) & (g265) & (g266) & (g273) & (g268)) + ((g263) & (g274) & (!g265) & (!g266) & (g273) & (!g268)) + ((g263) & (g274) & (!g265) & (g266) & (!g273) & (g268)) + ((g263) & (g274) & (g265) & (!g266) & (!g273) & (!g268)) + ((g263) & (g274) & (g265) & (!g266) & (g273) & (g268)) + ((g263) & (g274) & (g265) & (g266) & (!g273) & (g268)));
	assign g317 = (((!g313) & (!g314) & (!g315) & (!g316) & (!g267) & (!g264)) + ((!g313) & (!g314) & (!g315) & (!g316) & (!g267) & (g264)) + ((!g313) & (!g314) & (!g315) & (!g316) & (g267) & (!g264)) + ((!g313) & (!g314) & (!g315) & (g316) & (!g267) & (!g264)) + ((!g313) & (!g314) & (!g315) & (g316) & (!g267) & (g264)) + ((!g313) & (!g314) & (!g315) & (g316) & (g267) & (!g264)) + ((!g313) & (!g314) & (!g315) & (g316) & (g267) & (g264)) + ((!g313) & (!g314) & (g315) & (!g316) & (!g267) & (!g264)) + ((!g313) & (!g314) & (g315) & (!g316) & (g267) & (!g264)) + ((!g313) & (!g314) & (g315) & (g316) & (!g267) & (!g264)) + ((!g313) & (!g314) & (g315) & (g316) & (g267) & (!g264)) + ((!g313) & (!g314) & (g315) & (g316) & (g267) & (g264)) + ((!g313) & (g314) & (!g315) & (!g316) & (!g267) & (!g264)) + ((!g313) & (g314) & (!g315) & (!g316) & (!g267) & (g264)) + ((!g313) & (g314) & (!g315) & (g316) & (!g267) & (!g264)) + ((!g313) & (g314) & (!g315) & (g316) & (!g267) & (g264)) + ((!g313) & (g314) & (!g315) & (g316) & (g267) & (g264)) + ((!g313) & (g314) & (g315) & (!g316) & (!g267) & (!g264)) + ((!g313) & (g314) & (g315) & (g316) & (!g267) & (!g264)) + ((!g313) & (g314) & (g315) & (g316) & (g267) & (g264)) + ((g313) & (!g314) & (!g315) & (!g316) & (!g267) & (g264)) + ((g313) & (!g314) & (!g315) & (!g316) & (g267) & (!g264)) + ((g313) & (!g314) & (!g315) & (g316) & (!g267) & (g264)) + ((g313) & (!g314) & (!g315) & (g316) & (g267) & (!g264)) + ((g313) & (!g314) & (!g315) & (g316) & (g267) & (g264)) + ((g313) & (!g314) & (g315) & (!g316) & (g267) & (!g264)) + ((g313) & (!g314) & (g315) & (g316) & (g267) & (!g264)) + ((g313) & (!g314) & (g315) & (g316) & (g267) & (g264)) + ((g313) & (g314) & (!g315) & (!g316) & (!g267) & (g264)) + ((g313) & (g314) & (!g315) & (g316) & (!g267) & (g264)) + ((g313) & (g314) & (!g315) & (g316) & (g267) & (g264)) + ((g313) & (g314) & (g315) & (g316) & (g267) & (g264)));
	assign g319 = (((!sk[10]) & (g317) & (!g318)) + ((!sk[10]) & (g317) & (g318)) + ((sk[10]) & (!g317) & (g318)) + ((sk[10]) & (g317) & (!g318)));
	assign g320 = (((!g267) & (!g264) & (!g265) & (!g266) & (!g273) & (g274)) + ((!g267) & (!g264) & (!g265) & (!g266) & (g273) & (!g274)) + ((!g267) & (!g264) & (!g265) & (g266) & (!g273) & (g274)) + ((!g267) & (!g264) & (!g265) & (g266) & (g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (!g266) & (!g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (!g266) & (g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (g266) & (!g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (g266) & (g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (g266) & (g273) & (g274)) + ((!g267) & (g264) & (!g265) & (!g266) & (g273) & (!g274)) + ((!g267) & (g264) & (!g265) & (g266) & (g273) & (!g274)) + ((!g267) & (g264) & (!g265) & (g266) & (g273) & (g274)) + ((!g267) & (g264) & (g265) & (!g266) & (g273) & (g274)) + ((!g267) & (g264) & (g265) & (g266) & (!g273) & (!g274)) + ((g267) & (!g264) & (!g265) & (!g266) & (!g273) & (g274)) + ((g267) & (!g264) & (!g265) & (g266) & (!g273) & (g274)) + ((g267) & (!g264) & (g265) & (g266) & (g273) & (g274)) + ((g267) & (g264) & (!g265) & (!g266) & (g273) & (g274)) + ((g267) & (g264) & (!g265) & (g266) & (!g273) & (!g274)) + ((g267) & (g264) & (!g265) & (g266) & (g273) & (!g274)) + ((g267) & (g264) & (g265) & (!g266) & (!g273) & (g274)) + ((g267) & (g264) & (g265) & (!g266) & (g273) & (!g274)) + ((g267) & (g264) & (g265) & (!g266) & (g273) & (g274)) + ((g267) & (g264) & (g265) & (g266) & (!g273) & (g274)));
	assign g321 = (((!g267) & (!g264) & (!g265) & (!g266) & (!g273) & (!g274)) + ((!g267) & (!g264) & (!g265) & (!g266) & (!g273) & (g274)) + ((!g267) & (!g264) & (!g265) & (g266) & (!g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (!g266) & (!g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (!g266) & (g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (!g266) & (g273) & (g274)) + ((!g267) & (!g264) & (g265) & (g266) & (!g273) & (g274)) + ((!g267) & (!g264) & (g265) & (g266) & (g273) & (g274)) + ((!g267) & (g264) & (!g265) & (!g266) & (!g273) & (!g274)) + ((!g267) & (g264) & (!g265) & (!g266) & (g273) & (!g274)) + ((!g267) & (g264) & (!g265) & (g266) & (!g273) & (!g274)) + ((!g267) & (g264) & (!g265) & (g266) & (!g273) & (g274)) + ((!g267) & (g264) & (!g265) & (g266) & (g273) & (g274)) + ((!g267) & (g264) & (g265) & (!g266) & (!g273) & (g274)) + ((!g267) & (g264) & (g265) & (g266) & (!g273) & (!g274)) + ((!g267) & (g264) & (g265) & (g266) & (!g273) & (g274)) + ((g267) & (!g264) & (!g265) & (!g266) & (!g273) & (g274)) + ((g267) & (!g264) & (!g265) & (!g266) & (g273) & (g274)) + ((g267) & (!g264) & (!g265) & (g266) & (!g273) & (!g274)) + ((g267) & (!g264) & (!g265) & (g266) & (g273) & (g274)) + ((g267) & (!g264) & (g265) & (!g266) & (!g273) & (!g274)) + ((g267) & (!g264) & (g265) & (!g266) & (g273) & (g274)) + ((g267) & (!g264) & (g265) & (g266) & (g273) & (!g274)) + ((g267) & (g264) & (!g265) & (!g266) & (!g273) & (!g274)) + ((g267) & (g264) & (!g265) & (!g266) & (!g273) & (g274)) + ((g267) & (g264) & (!g265) & (!g266) & (g273) & (g274)) + ((g267) & (g264) & (!g265) & (g266) & (!g273) & (g274)) + ((g267) & (g264) & (!g265) & (g266) & (g273) & (!g274)) + ((g267) & (g264) & (g265) & (!g266) & (g273) & (!g274)) + ((g267) & (g264) & (g265) & (!g266) & (g273) & (g274)));
	assign g322 = (((!g267) & (!g264) & (!g265) & (!g266) & (g273) & (!g274)) + ((!g267) & (!g264) & (!g265) & (g266) & (!g273) & (!g274)) + ((!g267) & (!g264) & (!g265) & (g266) & (g273) & (!g274)) + ((!g267) & (!g264) & (!g265) & (g266) & (g273) & (g274)) + ((!g267) & (!g264) & (g265) & (!g266) & (!g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (!g266) & (!g273) & (g274)) + ((!g267) & (!g264) & (g265) & (!g266) & (g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (g266) & (!g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (g266) & (g273) & (g274)) + ((!g267) & (g264) & (!g265) & (!g266) & (!g273) & (g274)) + ((!g267) & (g264) & (!g265) & (!g266) & (g273) & (!g274)) + ((!g267) & (g264) & (!g265) & (!g266) & (g273) & (g274)) + ((!g267) & (g264) & (g265) & (!g266) & (!g273) & (g274)) + ((!g267) & (g264) & (g265) & (!g266) & (g273) & (!g274)) + ((!g267) & (g264) & (g265) & (!g266) & (g273) & (g274)) + ((!g267) & (g264) & (g265) & (g266) & (!g273) & (!g274)) + ((g267) & (!g264) & (!g265) & (!g266) & (g273) & (!g274)) + ((g267) & (!g264) & (!g265) & (g266) & (!g273) & (!g274)) + ((g267) & (!g264) & (!g265) & (g266) & (g273) & (g274)) + ((g267) & (!g264) & (g265) & (!g266) & (!g273) & (!g274)) + ((g267) & (!g264) & (g265) & (!g266) & (!g273) & (g274)) + ((g267) & (!g264) & (g265) & (g266) & (!g273) & (!g274)) + ((g267) & (!g264) & (g265) & (g266) & (g273) & (!g274)) + ((g267) & (g264) & (!g265) & (!g266) & (g273) & (!g274)) + ((g267) & (g264) & (!g265) & (g266) & (!g273) & (!g274)) + ((g267) & (g264) & (!g265) & (g266) & (g273) & (g274)) + ((g267) & (g264) & (g265) & (!g266) & (!g273) & (!g274)) + ((g267) & (g264) & (g265) & (!g266) & (g273) & (!g274)) + ((g267) & (g264) & (g265) & (!g266) & (g273) & (g274)) + ((g267) & (g264) & (g265) & (g266) & (!g273) & (g274)));
	assign g323 = (((!g267) & (!g264) & (!g265) & (!g266) & (!g273) & (g274)) + ((!g267) & (!g264) & (!g265) & (g266) & (g273) & (!g274)) + ((!g267) & (!g264) & (!g265) & (g266) & (g273) & (g274)) + ((!g267) & (!g264) & (g265) & (!g266) & (!g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (!g266) & (!g273) & (g274)) + ((!g267) & (!g264) & (g265) & (g266) & (g273) & (!g274)) + ((!g267) & (!g264) & (g265) & (g266) & (g273) & (g274)) + ((!g267) & (g264) & (!g265) & (!g266) & (!g273) & (!g274)) + ((!g267) & (g264) & (!g265) & (!g266) & (!g273) & (g274)) + ((!g267) & (g264) & (!g265) & (!g266) & (g273) & (g274)) + ((!g267) & (g264) & (!g265) & (g266) & (!g273) & (g274)) + ((!g267) & (g264) & (g265) & (!g266) & (!g273) & (g274)) + ((!g267) & (g264) & (g265) & (g266) & (!g273) & (!g274)) + ((!g267) & (g264) & (g265) & (g266) & (!g273) & (g274)) + ((!g267) & (g264) & (g265) & (g266) & (g273) & (!g274)) + ((!g267) & (g264) & (g265) & (g266) & (g273) & (g274)) + ((g267) & (!g264) & (!g265) & (g266) & (!g273) & (g274)) + ((g267) & (!g264) & (g265) & (!g266) & (!g273) & (!g274)) + ((g267) & (!g264) & (g265) & (g266) & (!g273) & (!g274)) + ((g267) & (!g264) & (g265) & (g266) & (!g273) & (g274)) + ((g267) & (!g264) & (g265) & (g266) & (g273) & (g274)) + ((g267) & (g264) & (!g265) & (!g266) & (!g273) & (g274)) + ((g267) & (g264) & (!g265) & (!g266) & (g273) & (g274)) + ((g267) & (g264) & (!g265) & (g266) & (!g273) & (!g274)) + ((g267) & (g264) & (!g265) & (g266) & (g273) & (!g274)) + ((g267) & (g264) & (!g265) & (g266) & (g273) & (g274)) + ((g267) & (g264) & (g265) & (!g266) & (g273) & (g274)) + ((g267) & (g264) & (g265) & (g266) & (g273) & (g274)));
	assign g324 = (((!g320) & (!g321) & (!g322) & (!g323) & (!g263) & (g268)) + ((!g320) & (!g321) & (!g322) & (!g323) & (g263) & (!g268)) + ((!g320) & (!g321) & (!g322) & (!g323) & (g263) & (g268)) + ((!g320) & (!g321) & (!g322) & (g323) & (!g263) & (g268)) + ((!g320) & (!g321) & (!g322) & (g323) & (g263) & (!g268)) + ((!g320) & (!g321) & (g322) & (!g323) & (g263) & (!g268)) + ((!g320) & (!g321) & (g322) & (!g323) & (g263) & (g268)) + ((!g320) & (!g321) & (g322) & (g323) & (g263) & (!g268)) + ((!g320) & (g321) & (!g322) & (!g323) & (!g263) & (g268)) + ((!g320) & (g321) & (!g322) & (!g323) & (g263) & (g268)) + ((!g320) & (g321) & (!g322) & (g323) & (!g263) & (g268)) + ((!g320) & (g321) & (g322) & (!g323) & (g263) & (g268)) + ((g320) & (!g321) & (!g322) & (!g323) & (!g263) & (!g268)) + ((g320) & (!g321) & (!g322) & (!g323) & (!g263) & (g268)) + ((g320) & (!g321) & (!g322) & (!g323) & (g263) & (!g268)) + ((g320) & (!g321) & (!g322) & (!g323) & (g263) & (g268)) + ((g320) & (!g321) & (!g322) & (g323) & (!g263) & (!g268)) + ((g320) & (!g321) & (!g322) & (g323) & (!g263) & (g268)) + ((g320) & (!g321) & (!g322) & (g323) & (g263) & (!g268)) + ((g320) & (!g321) & (g322) & (!g323) & (!g263) & (!g268)) + ((g320) & (!g321) & (g322) & (!g323) & (g263) & (!g268)) + ((g320) & (!g321) & (g322) & (!g323) & (g263) & (g268)) + ((g320) & (!g321) & (g322) & (g323) & (!g263) & (!g268)) + ((g320) & (!g321) & (g322) & (g323) & (g263) & (!g268)) + ((g320) & (g321) & (!g322) & (!g323) & (!g263) & (!g268)) + ((g320) & (g321) & (!g322) & (!g323) & (!g263) & (g268)) + ((g320) & (g321) & (!g322) & (!g323) & (g263) & (g268)) + ((g320) & (g321) & (!g322) & (g323) & (!g263) & (!g268)) + ((g320) & (g321) & (!g322) & (g323) & (!g263) & (g268)) + ((g320) & (g321) & (g322) & (!g323) & (!g263) & (!g268)) + ((g320) & (g321) & (g322) & (!g323) & (g263) & (g268)) + ((g320) & (g321) & (g322) & (g323) & (!g263) & (!g268)));
	assign g326 = (((!sk[16]) & (g324) & (!g325)) + ((!sk[16]) & (g324) & (g325)) + ((sk[16]) & (!g324) & (g325)) + ((sk[16]) & (g324) & (!g325)));
	assign g333 = (((!g327) & (!g328) & (!g329) & (!g330) & (g331) & (g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g331) & (!g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g331) & (g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (g331) & (!g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (!g331) & (!g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (!g331) & (g332)) + ((!g327) & (!g328) & (g329) & (g330) & (!g331) & (!g332)) + ((!g327) & (!g328) & (g329) & (g330) & (g331) & (g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (g331) & (!g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (g331) & (g332)) + ((!g327) & (g328) & (!g329) & (g330) & (g331) & (!g332)) + ((!g327) & (g328) & (!g329) & (g330) & (g331) & (g332)) + ((!g327) & (g328) & (g329) & (!g330) & (g331) & (!g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (!g331) & (!g332)) + ((g327) & (!g328) & (g329) & (!g330) & (g331) & (!g332)) + ((g327) & (!g328) & (g329) & (g330) & (!g331) & (g332)) + ((g327) & (!g328) & (g329) & (g330) & (g331) & (g332)) + ((g327) & (g328) & (!g329) & (!g330) & (!g331) & (g332)) + ((g327) & (g328) & (!g329) & (!g330) & (g331) & (!g332)) + ((g327) & (g328) & (g329) & (!g330) & (!g331) & (g332)) + ((g327) & (g328) & (g329) & (!g330) & (g331) & (!g332)) + ((g327) & (g328) & (g329) & (g330) & (!g331) & (!g332)) + ((g327) & (g328) & (g329) & (g330) & (g331) & (!g332)) + ((g327) & (g328) & (g329) & (g330) & (g331) & (g332)));
	assign g334 = (((!g327) & (!g328) & (!g329) & (!g330) & (g331) & (!g332)) + ((!g327) & (!g328) & (!g329) & (!g330) & (g331) & (g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g331) & (!g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g331) & (g332)) + ((!g327) & (!g328) & (g329) & (g330) & (!g331) & (g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (!g331) & (!g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (!g331) & (g332)) + ((!g327) & (g328) & (g329) & (!g330) & (!g331) & (!g332)) + ((!g327) & (g328) & (g329) & (!g330) & (!g331) & (g332)) + ((!g327) & (g328) & (g329) & (!g330) & (g331) & (!g332)) + ((!g327) & (g328) & (g329) & (g330) & (g331) & (g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (!g331) & (g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (g331) & (!g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (g331) & (g332)) + ((g327) & (!g328) & (!g329) & (g330) & (g331) & (!g332)) + ((g327) & (!g328) & (g329) & (!g330) & (!g331) & (!g332)) + ((g327) & (!g328) & (g329) & (!g330) & (g331) & (g332)) + ((g327) & (!g328) & (g329) & (g330) & (!g331) & (g332)) + ((g327) & (!g328) & (g329) & (g330) & (g331) & (g332)) + ((g327) & (g328) & (!g329) & (!g330) & (!g331) & (!g332)) + ((g327) & (g328) & (!g329) & (!g330) & (!g331) & (g332)) + ((g327) & (g328) & (!g329) & (!g330) & (g331) & (!g332)) + ((g327) & (g328) & (!g329) & (!g330) & (g331) & (g332)) + ((g327) & (g328) & (!g329) & (g330) & (!g331) & (!g332)) + ((g327) & (g328) & (!g329) & (g330) & (g331) & (!g332)) + ((g327) & (g328) & (!g329) & (g330) & (g331) & (g332)) + ((g327) & (g328) & (g329) & (!g330) & (g331) & (!g332)) + ((g327) & (g328) & (g329) & (!g330) & (g331) & (g332)) + ((g327) & (g328) & (g329) & (g330) & (!g331) & (g332)) + ((g327) & (g328) & (g329) & (g330) & (g331) & (!g332)));
	assign g335 = (((!g327) & (!g328) & (!g329) & (!g330) & (!g331) & (!g332)) + ((!g327) & (!g328) & (!g329) & (!g330) & (g331) & (g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (g331) & (g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (!g331) & (!g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (!g331) & (g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (g331) & (g332)) + ((!g327) & (!g328) & (g329) & (g330) & (!g331) & (g332)) + ((!g327) & (!g328) & (g329) & (g330) & (g331) & (!g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (!g331) & (!g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (g331) & (!g332)) + ((!g327) & (g328) & (!g329) & (g330) & (g331) & (g332)) + ((!g327) & (g328) & (g329) & (g330) & (!g331) & (!g332)) + ((!g327) & (g328) & (g329) & (g330) & (g331) & (!g332)) + ((g327) & (!g328) & (!g329) & (g330) & (!g331) & (!g332)) + ((g327) & (!g328) & (!g329) & (g330) & (!g331) & (g332)) + ((g327) & (!g328) & (!g329) & (g330) & (g331) & (!g332)) + ((g327) & (!g328) & (g329) & (!g330) & (!g331) & (!g332)) + ((g327) & (!g328) & (g329) & (!g330) & (g331) & (g332)) + ((g327) & (!g328) & (g329) & (g330) & (!g331) & (!g332)) + ((g327) & (!g328) & (g329) & (g330) & (!g331) & (g332)) + ((g327) & (!g328) & (g329) & (g330) & (g331) & (!g332)) + ((g327) & (!g328) & (g329) & (g330) & (g331) & (g332)) + ((g327) & (g328) & (!g329) & (!g330) & (g331) & (g332)) + ((g327) & (g328) & (!g329) & (g330) & (!g331) & (!g332)) + ((g327) & (g328) & (!g329) & (g330) & (g331) & (!g332)) + ((g327) & (g328) & (!g329) & (g330) & (g331) & (g332)) + ((g327) & (g328) & (g329) & (!g330) & (!g331) & (!g332)) + ((g327) & (g328) & (g329) & (g330) & (!g331) & (!g332)) + ((g327) & (g328) & (g329) & (g330) & (!g331) & (g332)) + ((g327) & (g328) & (g329) & (g330) & (g331) & (g332)));
	assign g336 = (((!g327) & (!g328) & (!g329) & (!g330) & (!g331) & (g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (g331) & (!g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (g331) & (g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (!g331) & (g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (g331) & (g332)) + ((!g327) & (!g328) & (g329) & (g330) & (!g331) & (g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (!g331) & (!g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (!g331) & (g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (g331) & (!g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (g331) & (g332)) + ((!g327) & (g328) & (!g329) & (g330) & (g331) & (!g332)) + ((!g327) & (g328) & (!g329) & (g330) & (g331) & (g332)) + ((!g327) & (g328) & (g329) & (g330) & (!g331) & (!g332)) + ((!g327) & (g328) & (g329) & (g330) & (g331) & (!g332)) + ((!g327) & (g328) & (g329) & (g330) & (g331) & (g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (!g331) & (!g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (g331) & (g332)) + ((g327) & (!g328) & (!g329) & (g330) & (g331) & (!g332)) + ((g327) & (!g328) & (!g329) & (g330) & (g331) & (g332)) + ((g327) & (!g328) & (g329) & (!g330) & (!g331) & (g332)) + ((g327) & (!g328) & (g329) & (!g330) & (g331) & (!g332)) + ((g327) & (!g328) & (g329) & (g330) & (g331) & (!g332)) + ((g327) & (g328) & (!g329) & (!g330) & (!g331) & (g332)) + ((g327) & (g328) & (!g329) & (!g330) & (g331) & (g332)) + ((g327) & (g328) & (!g329) & (g330) & (g331) & (!g332)) + ((g327) & (g328) & (!g329) & (g330) & (g331) & (g332)) + ((g327) & (g328) & (g329) & (!g330) & (!g331) & (g332)) + ((g327) & (g328) & (g329) & (g330) & (!g331) & (!g332)));
	assign g339 = (((!g333) & (!g334) & (!g335) & (!g336) & (!g337) & (!g338)) + ((!g333) & (!g334) & (!g335) & (g336) & (!g337) & (!g338)) + ((!g333) & (!g334) & (!g335) & (g336) & (g337) & (g338)) + ((!g333) & (!g334) & (g335) & (!g336) & (!g337) & (!g338)) + ((!g333) & (!g334) & (g335) & (!g336) & (!g337) & (g338)) + ((!g333) & (!g334) & (g335) & (g336) & (!g337) & (!g338)) + ((!g333) & (!g334) & (g335) & (g336) & (!g337) & (g338)) + ((!g333) & (!g334) & (g335) & (g336) & (g337) & (g338)) + ((!g333) & (g334) & (!g335) & (!g336) & (!g337) & (!g338)) + ((!g333) & (g334) & (!g335) & (!g336) & (g337) & (!g338)) + ((!g333) & (g334) & (!g335) & (g336) & (!g337) & (!g338)) + ((!g333) & (g334) & (!g335) & (g336) & (g337) & (!g338)) + ((!g333) & (g334) & (!g335) & (g336) & (g337) & (g338)) + ((!g333) & (g334) & (g335) & (!g336) & (!g337) & (!g338)) + ((!g333) & (g334) & (g335) & (!g336) & (!g337) & (g338)) + ((!g333) & (g334) & (g335) & (!g336) & (g337) & (!g338)) + ((!g333) & (g334) & (g335) & (g336) & (!g337) & (!g338)) + ((!g333) & (g334) & (g335) & (g336) & (!g337) & (g338)) + ((!g333) & (g334) & (g335) & (g336) & (g337) & (!g338)) + ((!g333) & (g334) & (g335) & (g336) & (g337) & (g338)) + ((g333) & (!g334) & (!g335) & (g336) & (g337) & (g338)) + ((g333) & (!g334) & (g335) & (!g336) & (!g337) & (g338)) + ((g333) & (!g334) & (g335) & (g336) & (!g337) & (g338)) + ((g333) & (!g334) & (g335) & (g336) & (g337) & (g338)) + ((g333) & (g334) & (!g335) & (!g336) & (g337) & (!g338)) + ((g333) & (g334) & (!g335) & (g336) & (g337) & (!g338)) + ((g333) & (g334) & (!g335) & (g336) & (g337) & (g338)) + ((g333) & (g334) & (g335) & (!g336) & (!g337) & (g338)) + ((g333) & (g334) & (g335) & (!g336) & (g337) & (!g338)) + ((g333) & (g334) & (g335) & (g336) & (!g337) & (g338)) + ((g333) & (g334) & (g335) & (g336) & (g337) & (!g338)) + ((g333) & (g334) & (g335) & (g336) & (g337) & (g338)));
	assign g341 = (((!g339) & (sk[22]) & (g340)) + ((g339) & (!sk[22]) & (!g340)) + ((g339) & (!sk[22]) & (g340)) + ((g339) & (sk[22]) & (!g340)));
	assign g342 = (((!g327) & (!g328) & (!g329) & (!g330) & (!g337) & (g331)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g337) & (!g331)) + ((!g327) & (!g328) & (!g329) & (g330) & (g337) & (!g331)) + ((!g327) & (!g328) & (g329) & (!g330) & (g337) & (g331)) + ((!g327) & (!g328) & (g329) & (g330) & (!g337) & (g331)) + ((!g327) & (!g328) & (g329) & (g330) & (g337) & (!g331)) + ((!g327) & (g328) & (!g329) & (!g330) & (!g337) & (g331)) + ((!g327) & (g328) & (!g329) & (!g330) & (g337) & (!g331)) + ((!g327) & (g328) & (!g329) & (!g330) & (g337) & (g331)) + ((!g327) & (g328) & (g329) & (!g330) & (g337) & (g331)) + ((!g327) & (g328) & (g329) & (g330) & (g337) & (g331)) + ((g327) & (!g328) & (!g329) & (!g330) & (!g337) & (!g331)) + ((g327) & (!g328) & (!g329) & (!g330) & (g337) & (g331)) + ((g327) & (!g328) & (!g329) & (g330) & (!g337) & (!g331)) + ((g327) & (!g328) & (!g329) & (g330) & (g337) & (!g331)) + ((g327) & (!g328) & (g329) & (!g330) & (g337) & (!g331)) + ((g327) & (!g328) & (g329) & (!g330) & (g337) & (g331)) + ((g327) & (!g328) & (g329) & (g330) & (g337) & (!g331)) + ((g327) & (!g328) & (g329) & (g330) & (g337) & (g331)) + ((g327) & (g328) & (!g329) & (!g330) & (g337) & (!g331)) + ((g327) & (g328) & (!g329) & (!g330) & (g337) & (g331)) + ((g327) & (g328) & (!g329) & (g330) & (g337) & (g331)) + ((g327) & (g328) & (g329) & (!g330) & (!g337) & (!g331)) + ((g327) & (g328) & (g329) & (!g330) & (!g337) & (g331)) + ((g327) & (g328) & (g329) & (!g330) & (g337) & (!g331)) + ((g327) & (g328) & (g329) & (g330) & (!g337) & (g331)) + ((g327) & (g328) & (g329) & (g330) & (g337) & (!g331)));
	assign g343 = (((!g327) & (!g328) & (!g329) & (!g330) & (!g337) & (g331)) + ((!g327) & (!g328) & (!g329) & (!g330) & (g337) & (!g331)) + ((!g327) & (!g328) & (!g329) & (!g330) & (g337) & (g331)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g337) & (!g331)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g337) & (g331)) + ((!g327) & (!g328) & (!g329) & (g330) & (g337) & (g331)) + ((!g327) & (!g328) & (g329) & (!g330) & (g337) & (!g331)) + ((!g327) & (!g328) & (g329) & (g330) & (!g337) & (!g331)) + ((!g327) & (!g328) & (g329) & (g330) & (!g337) & (g331)) + ((!g327) & (!g328) & (g329) & (g330) & (g337) & (g331)) + ((!g327) & (g328) & (!g329) & (!g330) & (g337) & (g331)) + ((!g327) & (g328) & (!g329) & (g330) & (!g337) & (!g331)) + ((!g327) & (g328) & (!g329) & (g330) & (g337) & (!g331)) + ((!g327) & (g328) & (g329) & (!g330) & (g337) & (!g331)) + ((!g327) & (g328) & (g329) & (!g330) & (g337) & (g331)) + ((!g327) & (g328) & (g329) & (g330) & (!g337) & (!g331)) + ((g327) & (!g328) & (!g329) & (!g330) & (!g337) & (!g331)) + ((g327) & (!g328) & (!g329) & (g330) & (!g337) & (!g331)) + ((g327) & (!g328) & (!g329) & (g330) & (!g337) & (g331)) + ((g327) & (!g328) & (g329) & (!g330) & (!g337) & (g331)) + ((g327) & (!g328) & (g329) & (!g330) & (g337) & (g331)) + ((g327) & (!g328) & (g329) & (g330) & (!g337) & (!g331)) + ((g327) & (!g328) & (g329) & (g330) & (!g337) & (g331)) + ((g327) & (g328) & (!g329) & (g330) & (!g337) & (!g331)) + ((g327) & (g328) & (!g329) & (g330) & (g337) & (g331)) + ((g327) & (g328) & (g329) & (!g330) & (!g337) & (!g331)) + ((g327) & (g328) & (g329) & (!g330) & (!g337) & (g331)) + ((g327) & (g328) & (g329) & (!g330) & (g337) & (g331)) + ((g327) & (g328) & (g329) & (g330) & (!g337) & (!g331)) + ((g327) & (g328) & (g329) & (g330) & (!g337) & (g331)) + ((g327) & (g328) & (g329) & (g330) & (g337) & (!g331)));
	assign g344 = (((!g327) & (!g328) & (!g329) & (!g330) & (!g337) & (g331)) + ((!g327) & (!g328) & (!g329) & (g330) & (g337) & (!g331)) + ((!g327) & (!g328) & (g329) & (!g330) & (!g337) & (!g331)) + ((!g327) & (!g328) & (g329) & (!g330) & (g337) & (!g331)) + ((!g327) & (!g328) & (g329) & (g330) & (!g337) & (g331)) + ((!g327) & (!g328) & (g329) & (g330) & (g337) & (!g331)) + ((!g327) & (!g328) & (g329) & (g330) & (g337) & (g331)) + ((!g327) & (g328) & (!g329) & (!g330) & (!g337) & (!g331)) + ((!g327) & (g328) & (!g329) & (!g330) & (g337) & (!g331)) + ((!g327) & (g328) & (!g329) & (g330) & (!g337) & (!g331)) + ((!g327) & (g328) & (!g329) & (g330) & (g337) & (g331)) + ((!g327) & (g328) & (g329) & (!g330) & (g337) & (g331)) + ((!g327) & (g328) & (g329) & (g330) & (!g337) & (g331)) + ((!g327) & (g328) & (g329) & (g330) & (g337) & (!g331)) + ((g327) & (!g328) & (!g329) & (!g330) & (g337) & (g331)) + ((g327) & (!g328) & (!g329) & (g330) & (!g337) & (!g331)) + ((g327) & (!g328) & (!g329) & (g330) & (g337) & (!g331)) + ((g327) & (!g328) & (g329) & (!g330) & (!g337) & (!g331)) + ((g327) & (!g328) & (g329) & (!g330) & (!g337) & (g331)) + ((g327) & (!g328) & (g329) & (!g330) & (g337) & (!g331)) + ((g327) & (!g328) & (g329) & (!g330) & (g337) & (g331)) + ((g327) & (!g328) & (g329) & (g330) & (g337) & (!g331)) + ((g327) & (g328) & (!g329) & (!g330) & (!g337) & (g331)) + ((g327) & (g328) & (!g329) & (!g330) & (g337) & (g331)) + ((g327) & (g328) & (!g329) & (g330) & (!g337) & (g331)) + ((g327) & (g328) & (g329) & (!g330) & (!g337) & (!g331)) + ((g327) & (g328) & (g329) & (!g330) & (!g337) & (g331)) + ((g327) & (g328) & (g329) & (!g330) & (g337) & (g331)) + ((g327) & (g328) & (g329) & (g330) & (!g337) & (!g331)) + ((g327) & (g328) & (g329) & (g330) & (!g337) & (g331)) + ((g327) & (g328) & (g329) & (g330) & (g337) & (!g331)) + ((g327) & (g328) & (g329) & (g330) & (g337) & (g331)));
	assign g345 = (((!g327) & (!g328) & (!g329) & (!g330) & (g337) & (!g331)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g337) & (!g331)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g337) & (g331)) + ((!g327) & (!g328) & (g329) & (!g330) & (g337) & (g331)) + ((!g327) & (!g328) & (g329) & (g330) & (!g337) & (g331)) + ((!g327) & (g328) & (!g329) & (!g330) & (!g337) & (!g331)) + ((!g327) & (g328) & (!g329) & (!g330) & (g337) & (!g331)) + ((!g327) & (g328) & (!g329) & (g330) & (!g337) & (g331)) + ((!g327) & (g328) & (g329) & (!g330) & (!g337) & (g331)) + ((!g327) & (g328) & (g329) & (!g330) & (g337) & (!g331)) + ((!g327) & (g328) & (g329) & (!g330) & (g337) & (g331)) + ((!g327) & (g328) & (g329) & (g330) & (g337) & (!g331)) + ((!g327) & (g328) & (g329) & (g330) & (g337) & (g331)) + ((g327) & (!g328) & (!g329) & (!g330) & (!g337) & (!g331)) + ((g327) & (!g328) & (!g329) & (g330) & (!g337) & (!g331)) + ((g327) & (!g328) & (!g329) & (g330) & (!g337) & (g331)) + ((g327) & (!g328) & (!g329) & (g330) & (g337) & (!g331)) + ((g327) & (!g328) & (g329) & (!g330) & (!g337) & (!g331)) + ((g327) & (!g328) & (g329) & (!g330) & (g337) & (g331)) + ((g327) & (!g328) & (g329) & (g330) & (g337) & (!g331)) + ((g327) & (g328) & (!g329) & (!g330) & (!g337) & (!g331)) + ((g327) & (g328) & (!g329) & (g330) & (!g337) & (!g331)) + ((g327) & (g328) & (!g329) & (g330) & (g337) & (!g331)) + ((g327) & (g328) & (!g329) & (g330) & (g337) & (g331)) + ((g327) & (g328) & (g329) & (g330) & (!g337) & (g331)) + ((g327) & (g328) & (g329) & (g330) & (g337) & (g331)));
	assign g346 = (((!g342) & (!g343) & (!g344) & (!g345) & (!g332) & (!g338)) + ((!g342) & (!g343) & (!g344) & (!g345) & (g332) & (!g338)) + ((!g342) & (!g343) & (!g344) & (g345) & (!g332) & (!g338)) + ((!g342) & (!g343) & (!g344) & (g345) & (g332) & (!g338)) + ((!g342) & (!g343) & (!g344) & (g345) & (g332) & (g338)) + ((!g342) & (!g343) & (g344) & (!g345) & (!g332) & (!g338)) + ((!g342) & (!g343) & (g344) & (!g345) & (!g332) & (g338)) + ((!g342) & (!g343) & (g344) & (!g345) & (g332) & (!g338)) + ((!g342) & (!g343) & (g344) & (g345) & (!g332) & (!g338)) + ((!g342) & (!g343) & (g344) & (g345) & (!g332) & (g338)) + ((!g342) & (!g343) & (g344) & (g345) & (g332) & (!g338)) + ((!g342) & (!g343) & (g344) & (g345) & (g332) & (g338)) + ((!g342) & (g343) & (!g344) & (!g345) & (!g332) & (!g338)) + ((!g342) & (g343) & (!g344) & (g345) & (!g332) & (!g338)) + ((!g342) & (g343) & (!g344) & (g345) & (g332) & (g338)) + ((!g342) & (g343) & (g344) & (!g345) & (!g332) & (!g338)) + ((!g342) & (g343) & (g344) & (!g345) & (!g332) & (g338)) + ((!g342) & (g343) & (g344) & (g345) & (!g332) & (!g338)) + ((!g342) & (g343) & (g344) & (g345) & (!g332) & (g338)) + ((!g342) & (g343) & (g344) & (g345) & (g332) & (g338)) + ((g342) & (!g343) & (!g344) & (!g345) & (g332) & (!g338)) + ((g342) & (!g343) & (!g344) & (g345) & (g332) & (!g338)) + ((g342) & (!g343) & (!g344) & (g345) & (g332) & (g338)) + ((g342) & (!g343) & (g344) & (!g345) & (!g332) & (g338)) + ((g342) & (!g343) & (g344) & (!g345) & (g332) & (!g338)) + ((g342) & (!g343) & (g344) & (g345) & (!g332) & (g338)) + ((g342) & (!g343) & (g344) & (g345) & (g332) & (!g338)) + ((g342) & (!g343) & (g344) & (g345) & (g332) & (g338)) + ((g342) & (g343) & (!g344) & (g345) & (g332) & (g338)) + ((g342) & (g343) & (g344) & (!g345) & (!g332) & (g338)) + ((g342) & (g343) & (g344) & (g345) & (!g332) & (g338)) + ((g342) & (g343) & (g344) & (g345) & (g332) & (g338)));
	assign g348 = (((!sk[28]) & (g346) & (!g347)) + ((!sk[28]) & (g346) & (g347)) + ((sk[28]) & (!g346) & (g347)) + ((sk[28]) & (g346) & (!g347)));
	assign g349 = (((!g331) & (!g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((!g331) & (!g328) & (!g329) & (!g330) & (g337) & (g332)) + ((!g331) & (!g328) & (!g329) & (g330) & (!g337) & (g332)) + ((!g331) & (!g328) & (!g329) & (g330) & (g337) & (!g332)) + ((!g331) & (!g328) & (!g329) & (g330) & (g337) & (g332)) + ((!g331) & (!g328) & (g329) & (!g330) & (!g337) & (g332)) + ((!g331) & (!g328) & (g329) & (g330) & (!g337) & (!g332)) + ((!g331) & (!g328) & (g329) & (g330) & (g337) & (!g332)) + ((!g331) & (g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((!g331) & (g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((!g331) & (g328) & (!g329) & (g330) & (!g337) & (g332)) + ((!g331) & (g328) & (g329) & (!g330) & (!g337) & (!g332)) + ((!g331) & (g328) & (g329) & (!g330) & (!g337) & (g332)) + ((!g331) & (g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g331) & (g328) & (g329) & (!g330) & (g337) & (g332)) + ((g331) & (!g328) & (!g329) & (g330) & (!g337) & (g332)) + ((g331) & (!g328) & (!g329) & (g330) & (g337) & (g332)) + ((g331) & (g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((g331) & (g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((g331) & (g328) & (!g329) & (g330) & (g337) & (!g332)) + ((g331) & (g328) & (g329) & (g330) & (!g337) & (!g332)) + ((g331) & (g328) & (g329) & (g330) & (!g337) & (g332)));
	assign g350 = (((!g331) & (!g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((!g331) & (!g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((!g331) & (!g328) & (!g329) & (g330) & (g337) & (g332)) + ((!g331) & (!g328) & (g329) & (!g330) & (!g337) & (!g332)) + ((!g331) & (!g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g331) & (!g328) & (g329) & (g330) & (!g337) & (g332)) + ((!g331) & (g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((!g331) & (g328) & (!g329) & (!g330) & (g337) & (g332)) + ((!g331) & (g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((!g331) & (g328) & (!g329) & (g330) & (!g337) & (g332)) + ((!g331) & (g328) & (!g329) & (g330) & (g337) & (g332)) + ((!g331) & (g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g331) & (g328) & (g329) & (!g330) & (g337) & (g332)) + ((!g331) & (g328) & (g329) & (g330) & (g337) & (!g332)) + ((g331) & (!g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((g331) & (!g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((g331) & (!g328) & (!g329) & (!g330) & (g337) & (g332)) + ((g331) & (!g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((g331) & (!g328) & (!g329) & (g330) & (!g337) & (g332)) + ((g331) & (!g328) & (!g329) & (g330) & (g337) & (!g332)) + ((g331) & (!g328) & (g329) & (g330) & (!g337) & (!g332)) + ((g331) & (g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((g331) & (g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((g331) & (g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((g331) & (g328) & (!g329) & (g330) & (g337) & (!g332)) + ((g331) & (g328) & (!g329) & (g330) & (g337) & (g332)) + ((g331) & (g328) & (g329) & (!g330) & (!g337) & (!g332)) + ((g331) & (g328) & (g329) & (!g330) & (g337) & (!g332)) + ((g331) & (g328) & (g329) & (g330) & (!g337) & (g332)) + ((g331) & (g328) & (g329) & (g330) & (g337) & (g332)));
	assign g351 = (((!g331) & (!g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((!g331) & (!g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((!g331) & (!g328) & (!g329) & (g330) & (!g337) & (g332)) + ((!g331) & (!g328) & (g329) & (!g330) & (!g337) & (g332)) + ((!g331) & (!g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g331) & (!g328) & (g329) & (g330) & (!g337) & (g332)) + ((!g331) & (g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((!g331) & (g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((!g331) & (g328) & (!g329) & (g330) & (g337) & (!g332)) + ((!g331) & (g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g331) & (g328) & (g329) & (g330) & (!g337) & (!g332)) + ((!g331) & (g328) & (g329) & (g330) & (g337) & (!g332)) + ((g331) & (!g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((g331) & (!g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((g331) & (!g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((g331) & (!g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((g331) & (!g328) & (!g329) & (g330) & (!g337) & (g332)) + ((g331) & (!g328) & (!g329) & (g330) & (g337) & (!g332)) + ((g331) & (!g328) & (!g329) & (g330) & (g337) & (g332)) + ((g331) & (!g328) & (g329) & (!g330) & (!g337) & (g332)) + ((g331) & (!g328) & (g329) & (!g330) & (g337) & (!g332)) + ((g331) & (!g328) & (g329) & (g330) & (!g337) & (!g332)) + ((g331) & (!g328) & (g329) & (g330) & (g337) & (g332)) + ((g331) & (g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((g331) & (g328) & (!g329) & (!g330) & (g337) & (g332)) + ((g331) & (g328) & (g329) & (!g330) & (g337) & (g332)) + ((g331) & (g328) & (g329) & (g330) & (!g337) & (!g332)) + ((g331) & (g328) & (g329) & (g330) & (!g337) & (g332)) + ((g331) & (g328) & (g329) & (g330) & (g337) & (g332)));
	assign g352 = (((!g331) & (!g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((!g331) & (!g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((!g331) & (!g328) & (!g329) & (!g330) & (g337) & (g332)) + ((!g331) & (!g328) & (!g329) & (g330) & (!g337) & (g332)) + ((!g331) & (!g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g331) & (!g328) & (g329) & (g330) & (g337) & (g332)) + ((!g331) & (g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((!g331) & (g328) & (!g329) & (g330) & (!g337) & (g332)) + ((!g331) & (g328) & (!g329) & (g330) & (g337) & (g332)) + ((!g331) & (g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g331) & (g328) & (g329) & (!g330) & (g337) & (g332)) + ((!g331) & (g328) & (g329) & (g330) & (!g337) & (!g332)) + ((!g331) & (g328) & (g329) & (g330) & (!g337) & (g332)) + ((!g331) & (g328) & (g329) & (g330) & (g337) & (!g332)) + ((!g331) & (g328) & (g329) & (g330) & (g337) & (g332)) + ((g331) & (!g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((g331) & (!g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((g331) & (!g328) & (!g329) & (!g330) & (g337) & (g332)) + ((g331) & (!g328) & (!g329) & (g330) & (g337) & (g332)) + ((g331) & (!g328) & (g329) & (!g330) & (!g337) & (g332)) + ((g331) & (!g328) & (g329) & (!g330) & (g337) & (!g332)) + ((g331) & (!g328) & (g329) & (g330) & (g337) & (!g332)) + ((g331) & (g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((g331) & (g328) & (!g329) & (g330) & (!g337) & (g332)) + ((g331) & (g328) & (!g329) & (g330) & (g337) & (!g332)) + ((g331) & (g328) & (g329) & (!g330) & (g337) & (g332)) + ((g331) & (g328) & (g329) & (g330) & (!g337) & (!g332)));
	assign g353 = (((!g349) & (!g350) & (!g351) & (!g352) & (!g327) & (g338)) + ((!g349) & (!g350) & (!g351) & (!g352) & (g327) & (!g338)) + ((!g349) & (!g350) & (!g351) & (!g352) & (g327) & (g338)) + ((!g349) & (!g350) & (!g351) & (g352) & (!g327) & (g338)) + ((!g349) & (!g350) & (!g351) & (g352) & (g327) & (!g338)) + ((!g349) & (!g350) & (g351) & (!g352) & (g327) & (!g338)) + ((!g349) & (!g350) & (g351) & (!g352) & (g327) & (g338)) + ((!g349) & (!g350) & (g351) & (g352) & (g327) & (!g338)) + ((!g349) & (g350) & (!g351) & (!g352) & (!g327) & (g338)) + ((!g349) & (g350) & (!g351) & (!g352) & (g327) & (g338)) + ((!g349) & (g350) & (!g351) & (g352) & (!g327) & (g338)) + ((!g349) & (g350) & (g351) & (!g352) & (g327) & (g338)) + ((g349) & (!g350) & (!g351) & (!g352) & (!g327) & (!g338)) + ((g349) & (!g350) & (!g351) & (!g352) & (!g327) & (g338)) + ((g349) & (!g350) & (!g351) & (!g352) & (g327) & (!g338)) + ((g349) & (!g350) & (!g351) & (!g352) & (g327) & (g338)) + ((g349) & (!g350) & (!g351) & (g352) & (!g327) & (!g338)) + ((g349) & (!g350) & (!g351) & (g352) & (!g327) & (g338)) + ((g349) & (!g350) & (!g351) & (g352) & (g327) & (!g338)) + ((g349) & (!g350) & (g351) & (!g352) & (!g327) & (!g338)) + ((g349) & (!g350) & (g351) & (!g352) & (g327) & (!g338)) + ((g349) & (!g350) & (g351) & (!g352) & (g327) & (g338)) + ((g349) & (!g350) & (g351) & (g352) & (!g327) & (!g338)) + ((g349) & (!g350) & (g351) & (g352) & (g327) & (!g338)) + ((g349) & (g350) & (!g351) & (!g352) & (!g327) & (!g338)) + ((g349) & (g350) & (!g351) & (!g352) & (!g327) & (g338)) + ((g349) & (g350) & (!g351) & (!g352) & (g327) & (g338)) + ((g349) & (g350) & (!g351) & (g352) & (!g327) & (!g338)) + ((g349) & (g350) & (!g351) & (g352) & (!g327) & (g338)) + ((g349) & (g350) & (g351) & (!g352) & (!g327) & (!g338)) + ((g349) & (g350) & (g351) & (!g352) & (g327) & (g338)) + ((g349) & (g350) & (g351) & (g352) & (!g327) & (!g338)));
	assign g355 = (((!sk[34]) & (g353) & (!g354)) + ((!sk[34]) & (g353) & (g354)) + ((sk[34]) & (!g353) & (g354)) + ((sk[34]) & (g353) & (!g354)));
	assign g356 = (((!g327) & (!g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (g337) & (g332)) + ((!g327) & (!g328) & (g329) & (g330) & (!g337) & (!g332)) + ((!g327) & (!g328) & (g329) & (g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (g329) & (g330) & (g337) & (g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (g328) & (g329) & (!g330) & (!g337) & (!g332)) + ((!g327) & (g328) & (g329) & (g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((g327) & (!g328) & (g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (g329) & (!g330) & (!g337) & (g332)) + ((g327) & (!g328) & (g329) & (!g330) & (g337) & (!g332)) + ((g327) & (!g328) & (g329) & (g330) & (!g337) & (g332)) + ((g327) & (g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((g327) & (g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((g327) & (g328) & (!g329) & (g330) & (g337) & (!g332)) + ((g327) & (g328) & (g329) & (!g330) & (!g337) & (g332)) + ((g327) & (g328) & (g329) & (!g330) & (g337) & (g332)));
	assign g357 = (((!g327) & (!g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (!g329) & (!g330) & (g337) & (g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (g329) & (g330) & (!g337) & (!g332)) + ((!g327) & (!g328) & (g329) & (g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (g329) & (g330) & (g337) & (g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (g337) & (g332)) + ((!g327) & (g328) & (!g329) & (g330) & (g337) & (g332)) + ((!g327) & (g328) & (g329) & (!g330) & (!g337) & (!g332)) + ((!g327) & (g328) & (g329) & (!g330) & (!g337) & (g332)) + ((!g327) & (g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (g328) & (g329) & (g330) & (!g337) & (g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((g327) & (!g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (!g329) & (g330) & (!g337) & (g332)) + ((g327) & (!g328) & (!g329) & (g330) & (g337) & (g332)) + ((g327) & (!g328) & (g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (g329) & (!g330) & (!g337) & (g332)) + ((g327) & (!g328) & (g329) & (!g330) & (g337) & (g332)) + ((g327) & (!g328) & (g329) & (g330) & (!g337) & (g332)) + ((g327) & (g328) & (!g329) & (g330) & (!g337) & (g332)) + ((g327) & (g328) & (!g329) & (g330) & (g337) & (!g332)) + ((g327) & (g328) & (g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (g328) & (g329) & (g330) & (!g337) & (!g332)));
	assign g358 = (((!g327) & (!g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (!g329) & (!g330) & (g337) & (g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (g329) & (!g330) & (g337) & (g332)) + ((!g327) & (!g328) & (g329) & (g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (g329) & (g330) & (g337) & (g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (g337) & (g332)) + ((!g327) & (g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((!g327) & (g328) & (!g329) & (g330) & (!g337) & (g332)) + ((!g327) & (g328) & (g329) & (!g330) & (!g337) & (g332)) + ((!g327) & (g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (g328) & (g329) & (g330) & (g337) & (g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (g337) & (g332)) + ((g327) & (!g328) & (!g329) & (g330) & (g337) & (g332)) + ((g327) & (!g328) & (g329) & (g330) & (!g337) & (!g332)) + ((g327) & (g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((g327) & (g328) & (!g329) & (g330) & (g337) & (g332)) + ((g327) & (g328) & (g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (g328) & (g329) & (!g330) & (!g337) & (g332)) + ((g327) & (g328) & (g329) & (!g330) & (g337) & (g332)) + ((g327) & (g328) & (g329) & (g330) & (!g337) & (!g332)) + ((g327) & (g328) & (g329) & (g330) & (g337) & (g332)));
	assign g359 = (((!g327) & (!g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (!g329) & (g330) & (g337) & (g332)) + ((!g327) & (!g328) & (g329) & (g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (g329) & (g330) & (g337) & (g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (!g337) & (!g332)) + ((!g327) & (g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (g328) & (!g329) & (g330) & (!g337) & (!g332)) + ((!g327) & (g328) & (!g329) & (g330) & (!g337) & (g332)) + ((!g327) & (g328) & (!g329) & (g330) & (g337) & (!g332)) + ((!g327) & (g328) & (g329) & (!g330) & (!g337) & (!g332)) + ((!g327) & (g328) & (g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (g328) & (g329) & (!g330) & (g337) & (g332)) + ((g327) & (!g328) & (!g329) & (!g330) & (g337) & (g332)) + ((g327) & (!g328) & (!g329) & (g330) & (g337) & (!g332)) + ((g327) & (!g328) & (g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (g329) & (!g330) & (g337) & (!g332)) + ((g327) & (!g328) & (g329) & (!g330) & (g337) & (g332)) + ((g327) & (!g328) & (g329) & (g330) & (!g337) & (g332)) + ((g327) & (!g328) & (g329) & (g330) & (g337) & (!g332)) + ((g327) & (!g328) & (g329) & (g330) & (g337) & (g332)) + ((g327) & (g328) & (!g329) & (!g330) & (!g337) & (g332)) + ((g327) & (g328) & (!g329) & (!g330) & (g337) & (!g332)) + ((g327) & (g328) & (g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (g328) & (g329) & (!g330) & (!g337) & (g332)) + ((g327) & (g328) & (g329) & (g330) & (g337) & (g332)));
	assign g360 = (((!g356) & (!g357) & (!g358) & (!g359) & (!g338) & (g331)) + ((!g356) & (!g357) & (!g358) & (!g359) & (g338) & (!g331)) + ((!g356) & (!g357) & (!g358) & (!g359) & (g338) & (g331)) + ((!g356) & (!g357) & (!g358) & (g359) & (!g338) & (g331)) + ((!g356) & (!g357) & (!g358) & (g359) & (g338) & (!g331)) + ((!g356) & (!g357) & (g358) & (!g359) & (g338) & (!g331)) + ((!g356) & (!g357) & (g358) & (!g359) & (g338) & (g331)) + ((!g356) & (!g357) & (g358) & (g359) & (g338) & (!g331)) + ((!g356) & (g357) & (!g358) & (!g359) & (!g338) & (g331)) + ((!g356) & (g357) & (!g358) & (!g359) & (g338) & (g331)) + ((!g356) & (g357) & (!g358) & (g359) & (!g338) & (g331)) + ((!g356) & (g357) & (g358) & (!g359) & (g338) & (g331)) + ((g356) & (!g357) & (!g358) & (!g359) & (!g338) & (!g331)) + ((g356) & (!g357) & (!g358) & (!g359) & (!g338) & (g331)) + ((g356) & (!g357) & (!g358) & (!g359) & (g338) & (!g331)) + ((g356) & (!g357) & (!g358) & (!g359) & (g338) & (g331)) + ((g356) & (!g357) & (!g358) & (g359) & (!g338) & (!g331)) + ((g356) & (!g357) & (!g358) & (g359) & (!g338) & (g331)) + ((g356) & (!g357) & (!g358) & (g359) & (g338) & (!g331)) + ((g356) & (!g357) & (g358) & (!g359) & (!g338) & (!g331)) + ((g356) & (!g357) & (g358) & (!g359) & (g338) & (!g331)) + ((g356) & (!g357) & (g358) & (!g359) & (g338) & (g331)) + ((g356) & (!g357) & (g358) & (g359) & (!g338) & (!g331)) + ((g356) & (!g357) & (g358) & (g359) & (g338) & (!g331)) + ((g356) & (g357) & (!g358) & (!g359) & (!g338) & (!g331)) + ((g356) & (g357) & (!g358) & (!g359) & (!g338) & (g331)) + ((g356) & (g357) & (!g358) & (!g359) & (g338) & (g331)) + ((g356) & (g357) & (!g358) & (g359) & (!g338) & (!g331)) + ((g356) & (g357) & (!g358) & (g359) & (!g338) & (g331)) + ((g356) & (g357) & (g358) & (!g359) & (!g338) & (!g331)) + ((g356) & (g357) & (g358) & (!g359) & (g338) & (g331)) + ((g356) & (g357) & (g358) & (g359) & (!g338) & (!g331)));
	assign g362 = (((!g360) & (sk[40]) & (g361)) + ((g360) & (!sk[40]) & (!g361)) + ((g360) & (!sk[40]) & (g361)) + ((g360) & (sk[40]) & (!g361)));
	assign g363 = (((!g327) & (!g328) & (!g331) & (!g338) & (!g337) & (g332)) + ((!g327) & (!g328) & (g331) & (!g338) & (!g337) & (g332)) + ((!g327) & (!g328) & (g331) & (!g338) & (g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (!g338) & (g337) & (g332)) + ((!g327) & (!g328) & (g331) & (g338) & (!g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (g338) & (g337) & (!g332)) + ((!g327) & (g328) & (!g331) & (!g338) & (!g337) & (!g332)) + ((!g327) & (g328) & (!g331) & (!g338) & (!g337) & (g332)) + ((!g327) & (g328) & (!g331) & (g338) & (!g337) & (!g332)) + ((!g327) & (g328) & (!g331) & (g338) & (!g337) & (g332)) + ((!g327) & (g328) & (!g331) & (g338) & (g337) & (g332)) + ((!g327) & (g328) & (g331) & (g338) & (!g337) & (g332)) + ((!g327) & (g328) & (g331) & (g338) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g338) & (!g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g338) & (!g337) & (g332)) + ((g327) & (!g328) & (!g331) & (g338) & (!g337) & (g332)) + ((g327) & (!g328) & (g331) & (!g338) & (g337) & (!g332)) + ((g327) & (!g328) & (g331) & (g338) & (!g337) & (!g332)) + ((g327) & (!g328) & (g331) & (g338) & (!g337) & (g332)) + ((g327) & (!g328) & (g331) & (g338) & (g337) & (!g332)) + ((g327) & (g328) & (!g331) & (!g338) & (!g337) & (!g332)) + ((g327) & (g328) & (!g331) & (!g338) & (g337) & (!g332)) + ((g327) & (g328) & (!g331) & (g338) & (g337) & (!g332)) + ((g327) & (g328) & (g331) & (!g338) & (!g337) & (!g332)) + ((g327) & (g328) & (g331) & (!g338) & (!g337) & (g332)) + ((g327) & (g328) & (g331) & (g338) & (!g337) & (g332)));
	assign g364 = (((!g327) & (!g328) & (!g331) & (!g338) & (!g337) & (!g332)) + ((!g327) & (!g328) & (!g331) & (!g338) & (!g337) & (g332)) + ((!g327) & (!g328) & (!g331) & (!g338) & (g337) & (!g332)) + ((!g327) & (!g328) & (!g331) & (!g338) & (g337) & (g332)) + ((!g327) & (!g328) & (!g331) & (g338) & (!g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (!g338) & (!g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (!g338) & (g337) & (g332)) + ((!g327) & (!g328) & (g331) & (g338) & (!g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (g338) & (g337) & (g332)) + ((!g327) & (g328) & (!g331) & (!g338) & (!g337) & (g332)) + ((!g327) & (g328) & (!g331) & (g338) & (g337) & (!g332)) + ((!g327) & (g328) & (g331) & (!g338) & (!g337) & (!g332)) + ((!g327) & (g328) & (g331) & (!g338) & (!g337) & (g332)) + ((!g327) & (g328) & (g331) & (!g338) & (g337) & (!g332)) + ((!g327) & (g328) & (g331) & (!g338) & (g337) & (g332)) + ((!g327) & (g328) & (g331) & (g338) & (!g337) & (!g332)) + ((!g327) & (g328) & (g331) & (g338) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g338) & (!g337) & (g332)) + ((g327) & (!g328) & (!g331) & (!g338) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g338) & (g337) & (g332)) + ((g327) & (!g328) & (!g331) & (g338) & (!g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (g338) & (g337) & (g332)) + ((g327) & (!g328) & (g331) & (!g338) & (g337) & (!g332)) + ((g327) & (!g328) & (g331) & (!g338) & (g337) & (g332)) + ((g327) & (!g328) & (g331) & (g338) & (!g337) & (g332)) + ((g327) & (g328) & (!g331) & (!g338) & (g337) & (!g332)) + ((g327) & (g328) & (!g331) & (!g338) & (g337) & (g332)) + ((g327) & (g328) & (!g331) & (g338) & (!g337) & (!g332)) + ((g327) & (g328) & (!g331) & (g338) & (!g337) & (g332)) + ((g327) & (g328) & (g331) & (!g338) & (g337) & (!g332)) + ((g327) & (g328) & (g331) & (!g338) & (g337) & (g332)) + ((g327) & (g328) & (g331) & (g338) & (!g337) & (g332)));
	assign g365 = (((!g327) & (!g328) & (!g331) & (!g338) & (!g337) & (!g332)) + ((!g327) & (!g328) & (!g331) & (!g338) & (!g337) & (g332)) + ((!g327) & (!g328) & (g331) & (!g338) & (!g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (!g338) & (g337) & (g332)) + ((!g327) & (!g328) & (g331) & (g338) & (!g337) & (g332)) + ((!g327) & (g328) & (!g331) & (g338) & (!g337) & (!g332)) + ((!g327) & (g328) & (!g331) & (g338) & (g337) & (!g332)) + ((!g327) & (g328) & (!g331) & (g338) & (g337) & (g332)) + ((!g327) & (g328) & (g331) & (!g338) & (!g337) & (!g332)) + ((!g327) & (g328) & (g331) & (!g338) & (g337) & (!g332)) + ((!g327) & (g328) & (g331) & (!g338) & (g337) & (g332)) + ((!g327) & (g328) & (g331) & (g338) & (!g337) & (!g332)) + ((!g327) & (g328) & (g331) & (g338) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g338) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g338) & (g337) & (g332)) + ((g327) & (!g328) & (!g331) & (g338) & (!g337) & (g332)) + ((g327) & (!g328) & (!g331) & (g338) & (g337) & (g332)) + ((g327) & (!g328) & (g331) & (!g338) & (!g337) & (!g332)) + ((g327) & (!g328) & (g331) & (!g338) & (!g337) & (g332)) + ((g327) & (!g328) & (g331) & (!g338) & (g337) & (g332)) + ((g327) & (!g328) & (g331) & (g338) & (!g337) & (!g332)) + ((g327) & (!g328) & (g331) & (g338) & (!g337) & (g332)) + ((g327) & (!g328) & (g331) & (g338) & (g337) & (!g332)) + ((g327) & (!g328) & (g331) & (g338) & (g337) & (g332)) + ((g327) & (g328) & (!g331) & (!g338) & (!g337) & (g332)) + ((g327) & (g328) & (!g331) & (g338) & (!g337) & (!g332)) + ((g327) & (g328) & (!g331) & (g338) & (g337) & (!g332)) + ((g327) & (g328) & (g331) & (!g338) & (!g337) & (!g332)) + ((g327) & (g328) & (g331) & (!g338) & (!g337) & (g332)) + ((g327) & (g328) & (g331) & (!g338) & (g337) & (!g332)) + ((g327) & (g328) & (g331) & (g338) & (!g337) & (!g332)) + ((g327) & (g328) & (g331) & (g338) & (g337) & (!g332)));
	assign g366 = (((!g327) & (!g328) & (!g331) & (!g338) & (g337) & (g332)) + ((!g327) & (!g328) & (!g331) & (g338) & (!g337) & (!g332)) + ((!g327) & (!g328) & (!g331) & (g338) & (g337) & (g332)) + ((!g327) & (!g328) & (g331) & (!g338) & (!g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (!g338) & (g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (g338) & (!g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (g338) & (!g337) & (g332)) + ((!g327) & (!g328) & (g331) & (g338) & (g337) & (!g332)) + ((!g327) & (g328) & (!g331) & (!g338) & (!g337) & (!g332)) + ((!g327) & (g328) & (!g331) & (g338) & (!g337) & (g332)) + ((!g327) & (g328) & (!g331) & (g338) & (g337) & (!g332)) + ((!g327) & (g328) & (!g331) & (g338) & (g337) & (g332)) + ((!g327) & (g328) & (g331) & (!g338) & (!g337) & (!g332)) + ((!g327) & (g328) & (g331) & (g338) & (!g337) & (!g332)) + ((!g327) & (g328) & (g331) & (g338) & (!g337) & (g332)) + ((g327) & (!g328) & (!g331) & (!g338) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g338) & (g337) & (g332)) + ((g327) & (!g328) & (g331) & (!g338) & (!g337) & (!g332)) + ((g327) & (!g328) & (g331) & (!g338) & (g337) & (!g332)) + ((g327) & (!g328) & (g331) & (g338) & (g337) & (!g332)) + ((g327) & (g328) & (!g331) & (!g338) & (g337) & (!g332)) + ((g327) & (g328) & (!g331) & (g338) & (g337) & (g332)) + ((g327) & (g328) & (g331) & (!g338) & (!g337) & (!g332)) + ((g327) & (g328) & (g331) & (!g338) & (!g337) & (g332)) + ((g327) & (g328) & (g331) & (!g338) & (g337) & (!g332)) + ((g327) & (g328) & (g331) & (g338) & (!g337) & (!g332)));
	assign g367 = (((!g363) & (!g364) & (!g365) & (!g366) & (g329) & (g330)) + ((!g363) & (!g364) & (g365) & (!g366) & (!g329) & (g330)) + ((!g363) & (!g364) & (g365) & (!g366) & (g329) & (g330)) + ((!g363) & (!g364) & (g365) & (g366) & (!g329) & (g330)) + ((!g363) & (g364) & (!g365) & (!g366) & (g329) & (!g330)) + ((!g363) & (g364) & (!g365) & (!g366) & (g329) & (g330)) + ((!g363) & (g364) & (!g365) & (g366) & (g329) & (!g330)) + ((!g363) & (g364) & (g365) & (!g366) & (!g329) & (g330)) + ((!g363) & (g364) & (g365) & (!g366) & (g329) & (!g330)) + ((!g363) & (g364) & (g365) & (!g366) & (g329) & (g330)) + ((!g363) & (g364) & (g365) & (g366) & (!g329) & (g330)) + ((!g363) & (g364) & (g365) & (g366) & (g329) & (!g330)) + ((g363) & (!g364) & (!g365) & (!g366) & (!g329) & (!g330)) + ((g363) & (!g364) & (!g365) & (!g366) & (g329) & (g330)) + ((g363) & (!g364) & (!g365) & (g366) & (!g329) & (!g330)) + ((g363) & (!g364) & (g365) & (!g366) & (!g329) & (!g330)) + ((g363) & (!g364) & (g365) & (!g366) & (!g329) & (g330)) + ((g363) & (!g364) & (g365) & (!g366) & (g329) & (g330)) + ((g363) & (!g364) & (g365) & (g366) & (!g329) & (!g330)) + ((g363) & (!g364) & (g365) & (g366) & (!g329) & (g330)) + ((g363) & (g364) & (!g365) & (!g366) & (!g329) & (!g330)) + ((g363) & (g364) & (!g365) & (!g366) & (g329) & (!g330)) + ((g363) & (g364) & (!g365) & (!g366) & (g329) & (g330)) + ((g363) & (g364) & (!g365) & (g366) & (!g329) & (!g330)) + ((g363) & (g364) & (!g365) & (g366) & (g329) & (!g330)) + ((g363) & (g364) & (g365) & (!g366) & (!g329) & (!g330)) + ((g363) & (g364) & (g365) & (!g366) & (!g329) & (g330)) + ((g363) & (g364) & (g365) & (!g366) & (g329) & (!g330)) + ((g363) & (g364) & (g365) & (!g366) & (g329) & (g330)) + ((g363) & (g364) & (g365) & (g366) & (!g329) & (!g330)) + ((g363) & (g364) & (g365) & (g366) & (!g329) & (g330)) + ((g363) & (g364) & (g365) & (g366) & (g329) & (!g330)));
	assign g369 = (((!g367) & (sk[46]) & (g368)) + ((g367) & (!sk[46]) & (!g368)) + ((g367) & (!sk[46]) & (g368)) + ((g367) & (sk[46]) & (!g368)));
	assign g370 = (((!g327) & (!g328) & (!g331) & (!g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (!g331) & (!g330) & (g337) & (g332)) + ((!g327) & (!g328) & (!g331) & (g330) & (g337) & (g332)) + ((!g327) & (!g328) & (g331) & (!g330) & (!g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (!g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (g331) & (!g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (!g330) & (g337) & (g332)) + ((!g327) & (!g328) & (g331) & (g330) & (!g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (g330) & (!g337) & (g332)) + ((!g327) & (g328) & (!g331) & (!g330) & (!g337) & (g332)) + ((!g327) & (g328) & (!g331) & (!g330) & (g337) & (!g332)) + ((!g327) & (g328) & (!g331) & (g330) & (g337) & (g332)) + ((!g327) & (g328) & (g331) & (!g330) & (g337) & (!g332)) + ((!g327) & (g328) & (g331) & (!g330) & (g337) & (g332)) + ((!g327) & (g328) & (g331) & (g330) & (!g337) & (!g332)) + ((!g327) & (g328) & (g331) & (g330) & (!g337) & (g332)) + ((!g327) & (g328) & (g331) & (g330) & (g337) & (g332)) + ((g327) & (!g328) & (!g331) & (!g330) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g330) & (g337) & (g332)) + ((g327) & (!g328) & (!g331) & (g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (g330) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (g330) & (g337) & (g332)) + ((g327) & (!g328) & (g331) & (!g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (g331) & (!g330) & (g337) & (!g332)) + ((g327) & (!g328) & (g331) & (g330) & (g337) & (!g332)) + ((g327) & (g328) & (!g331) & (!g330) & (g337) & (g332)) + ((g327) & (g328) & (g331) & (!g330) & (!g337) & (!g332)) + ((g327) & (g328) & (g331) & (!g330) & (g337) & (g332)));
	assign g371 = (((!g327) & (!g328) & (!g331) & (!g330) & (!g337) & (!g332)) + ((!g327) & (!g328) & (!g331) & (g330) & (!g337) & (!g332)) + ((!g327) & (!g328) & (!g331) & (g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (!g331) & (g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (!g330) & (g337) & (g332)) + ((!g327) & (!g328) & (g331) & (g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (g331) & (g330) & (g337) & (g332)) + ((!g327) & (g328) & (!g331) & (!g330) & (!g337) & (!g332)) + ((!g327) & (g328) & (!g331) & (!g330) & (g337) & (!g332)) + ((!g327) & (g328) & (g331) & (!g330) & (!g337) & (g332)) + ((!g327) & (g328) & (g331) & (!g330) & (g337) & (g332)) + ((!g327) & (g328) & (g331) & (g330) & (!g337) & (g332)) + ((!g327) & (g328) & (g331) & (g330) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g330) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g330) & (g337) & (g332)) + ((g327) & (!g328) & (!g331) & (g330) & (!g337) & (g332)) + ((g327) & (!g328) & (!g331) & (g330) & (g337) & (g332)) + ((g327) & (!g328) & (g331) & (g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (g331) & (g330) & (!g337) & (g332)) + ((g327) & (!g328) & (g331) & (g330) & (g337) & (g332)) + ((g327) & (g328) & (!g331) & (!g330) & (!g337) & (g332)) + ((g327) & (g328) & (!g331) & (!g330) & (g337) & (!g332)) + ((g327) & (g328) & (!g331) & (g330) & (g337) & (!g332)) + ((g327) & (g328) & (g331) & (!g330) & (!g337) & (g332)) + ((g327) & (g328) & (g331) & (!g330) & (g337) & (g332)) + ((g327) & (g328) & (g331) & (g330) & (!g337) & (!g332)) + ((g327) & (g328) & (g331) & (g330) & (g337) & (g332)));
	assign g372 = (((!g327) & (!g328) & (!g331) & (!g330) & (g337) & (g332)) + ((!g327) & (!g328) & (!g331) & (g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (!g330) & (!g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (!g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (g331) & (!g330) & (g337) & (g332)) + ((!g327) & (!g328) & (g331) & (g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (g331) & (g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (g331) & (g330) & (g337) & (g332)) + ((!g327) & (g328) & (!g331) & (!g330) & (g337) & (!g332)) + ((!g327) & (g328) & (!g331) & (!g330) & (g337) & (g332)) + ((!g327) & (g328) & (g331) & (!g330) & (!g337) & (!g332)) + ((!g327) & (g328) & (g331) & (g330) & (!g337) & (g332)) + ((!g327) & (g328) & (g331) & (g330) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g330) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (!g330) & (g337) & (g332)) + ((g327) & (!g328) & (!g331) & (g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (g330) & (!g337) & (g332)) + ((g327) & (!g328) & (g331) & (!g330) & (!g337) & (g332)) + ((g327) & (!g328) & (g331) & (!g330) & (g337) & (g332)) + ((g327) & (!g328) & (g331) & (g330) & (g337) & (!g332)) + ((g327) & (g328) & (!g331) & (!g330) & (!g337) & (!g332)) + ((g327) & (g328) & (!g331) & (!g330) & (!g337) & (g332)) + ((g327) & (g328) & (!g331) & (!g330) & (g337) & (g332)) + ((g327) & (g328) & (!g331) & (g330) & (!g337) & (g332)) + ((g327) & (g328) & (!g331) & (g330) & (g337) & (!g332)) + ((g327) & (g328) & (g331) & (!g330) & (!g337) & (g332)) + ((g327) & (g328) & (g331) & (!g330) & (g337) & (!g332)) + ((g327) & (g328) & (g331) & (g330) & (!g337) & (!g332)) + ((g327) & (g328) & (g331) & (g330) & (g337) & (!g332)) + ((g327) & (g328) & (g331) & (g330) & (g337) & (g332)));
	assign g373 = (((!g327) & (!g328) & (!g331) & (!g330) & (g337) & (!g332)) + ((!g327) & (!g328) & (!g331) & (g330) & (!g337) & (!g332)) + ((!g327) & (!g328) & (!g331) & (g330) & (g337) & (g332)) + ((!g327) & (!g328) & (g331) & (!g330) & (!g337) & (g332)) + ((!g327) & (!g328) & (g331) & (!g330) & (g337) & (g332)) + ((!g327) & (!g328) & (g331) & (g330) & (g337) & (g332)) + ((!g327) & (g328) & (!g331) & (!g330) & (!g337) & (g332)) + ((!g327) & (g328) & (!g331) & (g330) & (!g337) & (g332)) + ((!g327) & (g328) & (!g331) & (g330) & (g337) & (g332)) + ((!g327) & (g328) & (g331) & (!g330) & (!g337) & (!g332)) + ((!g327) & (g328) & (g331) & (!g330) & (g337) & (!g332)) + ((!g327) & (g328) & (g331) & (g330) & (!g337) & (g332)) + ((!g327) & (g328) & (g331) & (g330) & (g337) & (g332)) + ((g327) & (!g328) & (!g331) & (!g330) & (g337) & (!g332)) + ((g327) & (!g328) & (!g331) & (g330) & (g337) & (g332)) + ((g327) & (!g328) & (g331) & (!g330) & (!g337) & (!g332)) + ((g327) & (!g328) & (g331) & (!g330) & (g337) & (g332)) + ((g327) & (!g328) & (g331) & (g330) & (!g337) & (!g332)) + ((g327) & (g328) & (!g331) & (!g330) & (g337) & (g332)) + ((g327) & (g328) & (!g331) & (g330) & (!g337) & (!g332)) + ((g327) & (g328) & (!g331) & (g330) & (!g337) & (g332)) + ((g327) & (g328) & (g331) & (!g330) & (g337) & (g332)));
	assign g374 = (((!g370) & (!g371) & (!g372) & (!g373) & (!g338) & (!g329)) + ((!g370) & (!g371) & (!g372) & (!g373) & (!g338) & (g329)) + ((!g370) & (!g371) & (!g372) & (!g373) & (g338) & (!g329)) + ((!g370) & (!g371) & (!g372) & (g373) & (!g338) & (!g329)) + ((!g370) & (!g371) & (!g372) & (g373) & (!g338) & (g329)) + ((!g370) & (!g371) & (!g372) & (g373) & (g338) & (!g329)) + ((!g370) & (!g371) & (!g372) & (g373) & (g338) & (g329)) + ((!g370) & (!g371) & (g372) & (!g373) & (!g338) & (!g329)) + ((!g370) & (!g371) & (g372) & (!g373) & (g338) & (!g329)) + ((!g370) & (!g371) & (g372) & (g373) & (!g338) & (!g329)) + ((!g370) & (!g371) & (g372) & (g373) & (g338) & (!g329)) + ((!g370) & (!g371) & (g372) & (g373) & (g338) & (g329)) + ((!g370) & (g371) & (!g372) & (!g373) & (!g338) & (!g329)) + ((!g370) & (g371) & (!g372) & (!g373) & (!g338) & (g329)) + ((!g370) & (g371) & (!g372) & (g373) & (!g338) & (!g329)) + ((!g370) & (g371) & (!g372) & (g373) & (!g338) & (g329)) + ((!g370) & (g371) & (!g372) & (g373) & (g338) & (g329)) + ((!g370) & (g371) & (g372) & (!g373) & (!g338) & (!g329)) + ((!g370) & (g371) & (g372) & (g373) & (!g338) & (!g329)) + ((!g370) & (g371) & (g372) & (g373) & (g338) & (g329)) + ((g370) & (!g371) & (!g372) & (!g373) & (!g338) & (g329)) + ((g370) & (!g371) & (!g372) & (!g373) & (g338) & (!g329)) + ((g370) & (!g371) & (!g372) & (g373) & (!g338) & (g329)) + ((g370) & (!g371) & (!g372) & (g373) & (g338) & (!g329)) + ((g370) & (!g371) & (!g372) & (g373) & (g338) & (g329)) + ((g370) & (!g371) & (g372) & (!g373) & (g338) & (!g329)) + ((g370) & (!g371) & (g372) & (g373) & (g338) & (!g329)) + ((g370) & (!g371) & (g372) & (g373) & (g338) & (g329)) + ((g370) & (g371) & (!g372) & (!g373) & (!g338) & (g329)) + ((g370) & (g371) & (!g372) & (g373) & (!g338) & (g329)) + ((g370) & (g371) & (!g372) & (g373) & (g338) & (g329)) + ((g370) & (g371) & (g372) & (g373) & (g338) & (g329)));
	assign g376 = (((!g374) & (sk[52]) & (g375)) + ((g374) & (!sk[52]) & (!g375)) + ((g374) & (!sk[52]) & (g375)) + ((g374) & (sk[52]) & (!g375)));
	assign g377 = (((!g327) & (!g338) & (!g329) & (!g330) & (!g337) & (g332)) + ((!g327) & (!g338) & (!g329) & (!g330) & (g337) & (g332)) + ((!g327) & (!g338) & (!g329) & (g330) & (!g337) & (!g332)) + ((!g327) & (!g338) & (!g329) & (g330) & (!g337) & (g332)) + ((!g327) & (!g338) & (!g329) & (g330) & (g337) & (!g332)) + ((!g327) & (!g338) & (!g329) & (g330) & (g337) & (g332)) + ((!g327) & (!g338) & (g329) & (!g330) & (!g337) & (g332)) + ((!g327) & (!g338) & (g329) & (!g330) & (g337) & (g332)) + ((!g327) & (!g338) & (g329) & (g330) & (g337) & (!g332)) + ((!g327) & (g338) & (g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (g338) & (g329) & (!g330) & (g337) & (g332)) + ((!g327) & (g338) & (g329) & (g330) & (!g337) & (g332)) + ((g327) & (!g338) & (!g329) & (!g330) & (g337) & (!g332)) + ((g327) & (!g338) & (!g329) & (g330) & (!g337) & (!g332)) + ((g327) & (!g338) & (!g329) & (g330) & (!g337) & (g332)) + ((g327) & (!g338) & (!g329) & (g330) & (g337) & (g332)) + ((g327) & (!g338) & (g329) & (!g330) & (!g337) & (g332)) + ((g327) & (!g338) & (g329) & (!g330) & (g337) & (g332)) + ((g327) & (!g338) & (g329) & (g330) & (g337) & (!g332)) + ((g327) & (!g338) & (g329) & (g330) & (g337) & (g332)) + ((g327) & (g338) & (!g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (g338) & (!g329) & (!g330) & (!g337) & (g332)) + ((g327) & (g338) & (!g329) & (!g330) & (g337) & (!g332)) + ((g327) & (g338) & (!g329) & (g330) & (!g337) & (!g332)) + ((g327) & (g338) & (g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (g338) & (g329) & (!g330) & (!g337) & (g332)) + ((g327) & (g338) & (g329) & (!g330) & (g337) & (!g332)) + ((g327) & (g338) & (g329) & (g330) & (!g337) & (g332)));
	assign g378 = (((!g327) & (!g338) & (!g329) & (!g330) & (!g337) & (!g332)) + ((!g327) & (!g338) & (!g329) & (g330) & (g337) & (g332)) + ((!g327) & (!g338) & (g329) & (!g330) & (!g337) & (!g332)) + ((!g327) & (!g338) & (g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (!g338) & (g329) & (!g330) & (g337) & (g332)) + ((!g327) & (!g338) & (g329) & (g330) & (!g337) & (!g332)) + ((!g327) & (!g338) & (g329) & (g330) & (g337) & (g332)) + ((!g327) & (g338) & (!g329) & (!g330) & (!g337) & (!g332)) + ((!g327) & (g338) & (!g329) & (!g330) & (g337) & (g332)) + ((!g327) & (g338) & (!g329) & (g330) & (!g337) & (g332)) + ((!g327) & (g338) & (g329) & (!g330) & (!g337) & (!g332)) + ((!g327) & (g338) & (g329) & (!g330) & (g337) & (g332)) + ((!g327) & (g338) & (g329) & (g330) & (g337) & (!g332)) + ((!g327) & (g338) & (g329) & (g330) & (g337) & (g332)) + ((g327) & (!g338) & (!g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (!g338) & (!g329) & (!g330) & (g337) & (g332)) + ((g327) & (!g338) & (!g329) & (g330) & (!g337) & (!g332)) + ((g327) & (!g338) & (!g329) & (g330) & (g337) & (g332)) + ((g327) & (!g338) & (g329) & (!g330) & (g337) & (g332)) + ((g327) & (!g338) & (g329) & (g330) & (!g337) & (g332)) + ((g327) & (g338) & (!g329) & (!g330) & (g337) & (!g332)) + ((g327) & (g338) & (!g329) & (!g330) & (g337) & (g332)) + ((g327) & (g338) & (!g329) & (g330) & (!g337) & (g332)) + ((g327) & (g338) & (!g329) & (g330) & (g337) & (!g332)) + ((g327) & (g338) & (!g329) & (g330) & (g337) & (g332)) + ((g327) & (g338) & (g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (g338) & (g329) & (!g330) & (g337) & (!g332)) + ((g327) & (g338) & (g329) & (g330) & (!g337) & (!g332)));
	assign g379 = (((!g327) & (!g338) & (!g329) & (!g330) & (!g337) & (g332)) + ((!g327) & (!g338) & (!g329) & (!g330) & (g337) & (g332)) + ((!g327) & (!g338) & (!g329) & (g330) & (g337) & (!g332)) + ((!g327) & (!g338) & (!g329) & (g330) & (g337) & (g332)) + ((!g327) & (!g338) & (g329) & (!g330) & (g337) & (g332)) + ((!g327) & (!g338) & (g329) & (g330) & (!g337) & (!g332)) + ((!g327) & (!g338) & (g329) & (g330) & (!g337) & (g332)) + ((!g327) & (!g338) & (g329) & (g330) & (g337) & (g332)) + ((!g327) & (g338) & (!g329) & (!g330) & (!g337) & (!g332)) + ((!g327) & (g338) & (!g329) & (!g330) & (!g337) & (g332)) + ((!g327) & (g338) & (!g329) & (!g330) & (g337) & (g332)) + ((!g327) & (g338) & (!g329) & (g330) & (!g337) & (g332)) + ((!g327) & (g338) & (!g329) & (g330) & (g337) & (!g332)) + ((!g327) & (g338) & (g329) & (!g330) & (!g337) & (g332)) + ((!g327) & (g338) & (g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (g338) & (g329) & (g330) & (!g337) & (!g332)) + ((!g327) & (g338) & (g329) & (g330) & (g337) & (!g332)) + ((!g327) & (g338) & (g329) & (g330) & (g337) & (g332)) + ((g327) & (!g338) & (!g329) & (!g330) & (!g337) & (g332)) + ((g327) & (!g338) & (!g329) & (g330) & (!g337) & (!g332)) + ((g327) & (!g338) & (!g329) & (g330) & (g337) & (!g332)) + ((g327) & (!g338) & (g329) & (!g330) & (g337) & (g332)) + ((g327) & (!g338) & (g329) & (g330) & (!g337) & (g332)) + ((g327) & (g338) & (!g329) & (!g330) & (!g337) & (g332)) + ((g327) & (g338) & (!g329) & (g330) & (!g337) & (!g332)) + ((g327) & (g338) & (!g329) & (g330) & (g337) & (!g332)) + ((g327) & (g338) & (g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (g338) & (g329) & (!g330) & (g337) & (!g332)) + ((g327) & (g338) & (g329) & (!g330) & (g337) & (g332)) + ((g327) & (g338) & (g329) & (g330) & (g337) & (g332)));
	assign g380 = (((!g327) & (!g338) & (!g329) & (!g330) & (g337) & (g332)) + ((!g327) & (!g338) & (!g329) & (g330) & (!g337) & (!g332)) + ((!g327) & (!g338) & (!g329) & (g330) & (g337) & (g332)) + ((!g327) & (!g338) & (g329) & (!g330) & (!g337) & (!g332)) + ((!g327) & (!g338) & (g329) & (g330) & (g337) & (!g332)) + ((!g327) & (!g338) & (g329) & (g330) & (g337) & (g332)) + ((!g327) & (g338) & (!g329) & (g330) & (!g337) & (!g332)) + ((!g327) & (g338) & (!g329) & (g330) & (g337) & (!g332)) + ((!g327) & (g338) & (g329) & (!g330) & (g337) & (!g332)) + ((!g327) & (g338) & (g329) & (!g330) & (g337) & (g332)) + ((g327) & (!g338) & (!g329) & (!g330) & (!g337) & (g332)) + ((g327) & (!g338) & (!g329) & (!g330) & (g337) & (!g332)) + ((g327) & (!g338) & (!g329) & (g330) & (!g337) & (g332)) + ((g327) & (!g338) & (g329) & (!g330) & (g337) & (!g332)) + ((g327) & (!g338) & (g329) & (!g330) & (g337) & (g332)) + ((g327) & (!g338) & (g329) & (g330) & (g337) & (!g332)) + ((g327) & (!g338) & (g329) & (g330) & (g337) & (g332)) + ((g327) & (g338) & (!g329) & (!g330) & (g337) & (!g332)) + ((g327) & (g338) & (!g329) & (g330) & (!g337) & (g332)) + ((g327) & (g338) & (g329) & (!g330) & (!g337) & (!g332)) + ((g327) & (g338) & (g329) & (!g330) & (g337) & (g332)) + ((g327) & (g338) & (g329) & (g330) & (!g337) & (g332)));
	assign g381 = (((!g377) & (!g378) & (!g379) & (!g380) & (!g331) & (!g328)) + ((!g377) & (!g378) & (!g379) & (!g380) & (!g331) & (g328)) + ((!g377) & (!g378) & (!g379) & (!g380) & (g331) & (!g328)) + ((!g377) & (!g378) & (!g379) & (g380) & (!g331) & (!g328)) + ((!g377) & (!g378) & (!g379) & (g380) & (!g331) & (g328)) + ((!g377) & (!g378) & (!g379) & (g380) & (g331) & (!g328)) + ((!g377) & (!g378) & (!g379) & (g380) & (g331) & (g328)) + ((!g377) & (!g378) & (g379) & (!g380) & (!g331) & (!g328)) + ((!g377) & (!g378) & (g379) & (!g380) & (g331) & (!g328)) + ((!g377) & (!g378) & (g379) & (g380) & (!g331) & (!g328)) + ((!g377) & (!g378) & (g379) & (g380) & (g331) & (!g328)) + ((!g377) & (!g378) & (g379) & (g380) & (g331) & (g328)) + ((!g377) & (g378) & (!g379) & (!g380) & (!g331) & (!g328)) + ((!g377) & (g378) & (!g379) & (!g380) & (!g331) & (g328)) + ((!g377) & (g378) & (!g379) & (g380) & (!g331) & (!g328)) + ((!g377) & (g378) & (!g379) & (g380) & (!g331) & (g328)) + ((!g377) & (g378) & (!g379) & (g380) & (g331) & (g328)) + ((!g377) & (g378) & (g379) & (!g380) & (!g331) & (!g328)) + ((!g377) & (g378) & (g379) & (g380) & (!g331) & (!g328)) + ((!g377) & (g378) & (g379) & (g380) & (g331) & (g328)) + ((g377) & (!g378) & (!g379) & (!g380) & (!g331) & (g328)) + ((g377) & (!g378) & (!g379) & (!g380) & (g331) & (!g328)) + ((g377) & (!g378) & (!g379) & (g380) & (!g331) & (g328)) + ((g377) & (!g378) & (!g379) & (g380) & (g331) & (!g328)) + ((g377) & (!g378) & (!g379) & (g380) & (g331) & (g328)) + ((g377) & (!g378) & (g379) & (!g380) & (g331) & (!g328)) + ((g377) & (!g378) & (g379) & (g380) & (g331) & (!g328)) + ((g377) & (!g378) & (g379) & (g380) & (g331) & (g328)) + ((g377) & (g378) & (!g379) & (!g380) & (!g331) & (g328)) + ((g377) & (g378) & (!g379) & (g380) & (!g331) & (g328)) + ((g377) & (g378) & (!g379) & (g380) & (g331) & (g328)) + ((g377) & (g378) & (g379) & (g380) & (g331) & (g328)));
	assign g383 = (((!g381) & (sk[58]) & (g382)) + ((g381) & (!sk[58]) & (!g382)) + ((g381) & (!sk[58]) & (g382)) + ((g381) & (sk[58]) & (!g382)));
	assign g384 = (((!g331) & (!g328) & (!g329) & (!g330) & (!g337) & (g338)) + ((!g331) & (!g328) & (!g329) & (!g330) & (g337) & (!g338)) + ((!g331) & (!g328) & (!g329) & (g330) & (!g337) & (g338)) + ((!g331) & (!g328) & (!g329) & (g330) & (g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (!g330) & (!g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (!g330) & (g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (g330) & (!g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (g330) & (g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (g330) & (g337) & (g338)) + ((!g331) & (g328) & (!g329) & (!g330) & (g337) & (!g338)) + ((!g331) & (g328) & (!g329) & (g330) & (g337) & (!g338)) + ((!g331) & (g328) & (!g329) & (g330) & (g337) & (g338)) + ((!g331) & (g328) & (g329) & (!g330) & (g337) & (g338)) + ((!g331) & (g328) & (g329) & (g330) & (!g337) & (!g338)) + ((g331) & (!g328) & (!g329) & (!g330) & (!g337) & (g338)) + ((g331) & (!g328) & (!g329) & (g330) & (!g337) & (g338)) + ((g331) & (!g328) & (g329) & (g330) & (g337) & (g338)) + ((g331) & (g328) & (!g329) & (!g330) & (g337) & (g338)) + ((g331) & (g328) & (!g329) & (g330) & (!g337) & (!g338)) + ((g331) & (g328) & (!g329) & (g330) & (g337) & (!g338)) + ((g331) & (g328) & (g329) & (!g330) & (!g337) & (g338)) + ((g331) & (g328) & (g329) & (!g330) & (g337) & (!g338)) + ((g331) & (g328) & (g329) & (!g330) & (g337) & (g338)) + ((g331) & (g328) & (g329) & (g330) & (!g337) & (g338)));
	assign g385 = (((!g331) & (!g328) & (!g329) & (!g330) & (!g337) & (!g338)) + ((!g331) & (!g328) & (!g329) & (!g330) & (!g337) & (g338)) + ((!g331) & (!g328) & (!g329) & (g330) & (!g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (!g330) & (!g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (!g330) & (g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (!g330) & (g337) & (g338)) + ((!g331) & (!g328) & (g329) & (g330) & (!g337) & (g338)) + ((!g331) & (!g328) & (g329) & (g330) & (g337) & (g338)) + ((!g331) & (g328) & (!g329) & (!g330) & (!g337) & (!g338)) + ((!g331) & (g328) & (!g329) & (!g330) & (g337) & (!g338)) + ((!g331) & (g328) & (!g329) & (g330) & (!g337) & (!g338)) + ((!g331) & (g328) & (!g329) & (g330) & (!g337) & (g338)) + ((!g331) & (g328) & (!g329) & (g330) & (g337) & (g338)) + ((!g331) & (g328) & (g329) & (!g330) & (!g337) & (g338)) + ((!g331) & (g328) & (g329) & (g330) & (!g337) & (!g338)) + ((!g331) & (g328) & (g329) & (g330) & (!g337) & (g338)) + ((g331) & (!g328) & (!g329) & (!g330) & (!g337) & (g338)) + ((g331) & (!g328) & (!g329) & (!g330) & (g337) & (g338)) + ((g331) & (!g328) & (!g329) & (g330) & (!g337) & (!g338)) + ((g331) & (!g328) & (!g329) & (g330) & (g337) & (g338)) + ((g331) & (!g328) & (g329) & (!g330) & (!g337) & (!g338)) + ((g331) & (!g328) & (g329) & (!g330) & (g337) & (g338)) + ((g331) & (!g328) & (g329) & (g330) & (g337) & (!g338)) + ((g331) & (g328) & (!g329) & (!g330) & (!g337) & (!g338)) + ((g331) & (g328) & (!g329) & (!g330) & (!g337) & (g338)) + ((g331) & (g328) & (!g329) & (!g330) & (g337) & (g338)) + ((g331) & (g328) & (!g329) & (g330) & (!g337) & (g338)) + ((g331) & (g328) & (!g329) & (g330) & (g337) & (!g338)) + ((g331) & (g328) & (g329) & (!g330) & (g337) & (!g338)) + ((g331) & (g328) & (g329) & (!g330) & (g337) & (g338)));
	assign g386 = (((!g331) & (!g328) & (!g329) & (!g330) & (g337) & (!g338)) + ((!g331) & (!g328) & (!g329) & (g330) & (!g337) & (!g338)) + ((!g331) & (!g328) & (!g329) & (g330) & (g337) & (!g338)) + ((!g331) & (!g328) & (!g329) & (g330) & (g337) & (g338)) + ((!g331) & (!g328) & (g329) & (!g330) & (!g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (!g330) & (!g337) & (g338)) + ((!g331) & (!g328) & (g329) & (!g330) & (g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (g330) & (!g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (g330) & (g337) & (g338)) + ((!g331) & (g328) & (!g329) & (!g330) & (!g337) & (g338)) + ((!g331) & (g328) & (!g329) & (!g330) & (g337) & (!g338)) + ((!g331) & (g328) & (!g329) & (!g330) & (g337) & (g338)) + ((!g331) & (g328) & (g329) & (!g330) & (!g337) & (g338)) + ((!g331) & (g328) & (g329) & (!g330) & (g337) & (!g338)) + ((!g331) & (g328) & (g329) & (!g330) & (g337) & (g338)) + ((!g331) & (g328) & (g329) & (g330) & (!g337) & (!g338)) + ((g331) & (!g328) & (!g329) & (!g330) & (g337) & (!g338)) + ((g331) & (!g328) & (!g329) & (g330) & (!g337) & (!g338)) + ((g331) & (!g328) & (!g329) & (g330) & (g337) & (g338)) + ((g331) & (!g328) & (g329) & (!g330) & (!g337) & (!g338)) + ((g331) & (!g328) & (g329) & (!g330) & (!g337) & (g338)) + ((g331) & (!g328) & (g329) & (g330) & (!g337) & (!g338)) + ((g331) & (!g328) & (g329) & (g330) & (g337) & (!g338)) + ((g331) & (g328) & (!g329) & (!g330) & (g337) & (!g338)) + ((g331) & (g328) & (!g329) & (g330) & (!g337) & (!g338)) + ((g331) & (g328) & (!g329) & (g330) & (g337) & (g338)) + ((g331) & (g328) & (g329) & (!g330) & (!g337) & (!g338)) + ((g331) & (g328) & (g329) & (!g330) & (g337) & (!g338)) + ((g331) & (g328) & (g329) & (!g330) & (g337) & (g338)) + ((g331) & (g328) & (g329) & (g330) & (!g337) & (g338)));
	assign g387 = (((!g331) & (!g328) & (!g329) & (!g330) & (!g337) & (g338)) + ((!g331) & (!g328) & (!g329) & (g330) & (g337) & (!g338)) + ((!g331) & (!g328) & (!g329) & (g330) & (g337) & (g338)) + ((!g331) & (!g328) & (g329) & (!g330) & (!g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (!g330) & (!g337) & (g338)) + ((!g331) & (!g328) & (g329) & (g330) & (g337) & (!g338)) + ((!g331) & (!g328) & (g329) & (g330) & (g337) & (g338)) + ((!g331) & (g328) & (!g329) & (!g330) & (!g337) & (!g338)) + ((!g331) & (g328) & (!g329) & (!g330) & (!g337) & (g338)) + ((!g331) & (g328) & (!g329) & (!g330) & (g337) & (g338)) + ((!g331) & (g328) & (!g329) & (g330) & (!g337) & (g338)) + ((!g331) & (g328) & (g329) & (!g330) & (!g337) & (g338)) + ((!g331) & (g328) & (g329) & (g330) & (!g337) & (!g338)) + ((!g331) & (g328) & (g329) & (g330) & (!g337) & (g338)) + ((!g331) & (g328) & (g329) & (g330) & (g337) & (!g338)) + ((!g331) & (g328) & (g329) & (g330) & (g337) & (g338)) + ((g331) & (!g328) & (!g329) & (g330) & (!g337) & (g338)) + ((g331) & (!g328) & (g329) & (!g330) & (!g337) & (!g338)) + ((g331) & (!g328) & (g329) & (g330) & (!g337) & (!g338)) + ((g331) & (!g328) & (g329) & (g330) & (!g337) & (g338)) + ((g331) & (!g328) & (g329) & (g330) & (g337) & (g338)) + ((g331) & (g328) & (!g329) & (!g330) & (!g337) & (g338)) + ((g331) & (g328) & (!g329) & (!g330) & (g337) & (g338)) + ((g331) & (g328) & (!g329) & (g330) & (!g337) & (!g338)) + ((g331) & (g328) & (!g329) & (g330) & (g337) & (!g338)) + ((g331) & (g328) & (!g329) & (g330) & (g337) & (g338)) + ((g331) & (g328) & (g329) & (!g330) & (g337) & (g338)) + ((g331) & (g328) & (g329) & (g330) & (g337) & (g338)));
	assign g388 = (((!g384) & (!g385) & (!g386) & (!g387) & (!g327) & (g332)) + ((!g384) & (!g385) & (!g386) & (!g387) & (g327) & (!g332)) + ((!g384) & (!g385) & (!g386) & (!g387) & (g327) & (g332)) + ((!g384) & (!g385) & (!g386) & (g387) & (!g327) & (g332)) + ((!g384) & (!g385) & (!g386) & (g387) & (g327) & (!g332)) + ((!g384) & (!g385) & (g386) & (!g387) & (g327) & (!g332)) + ((!g384) & (!g385) & (g386) & (!g387) & (g327) & (g332)) + ((!g384) & (!g385) & (g386) & (g387) & (g327) & (!g332)) + ((!g384) & (g385) & (!g386) & (!g387) & (!g327) & (g332)) + ((!g384) & (g385) & (!g386) & (!g387) & (g327) & (g332)) + ((!g384) & (g385) & (!g386) & (g387) & (!g327) & (g332)) + ((!g384) & (g385) & (g386) & (!g387) & (g327) & (g332)) + ((g384) & (!g385) & (!g386) & (!g387) & (!g327) & (!g332)) + ((g384) & (!g385) & (!g386) & (!g387) & (!g327) & (g332)) + ((g384) & (!g385) & (!g386) & (!g387) & (g327) & (!g332)) + ((g384) & (!g385) & (!g386) & (!g387) & (g327) & (g332)) + ((g384) & (!g385) & (!g386) & (g387) & (!g327) & (!g332)) + ((g384) & (!g385) & (!g386) & (g387) & (!g327) & (g332)) + ((g384) & (!g385) & (!g386) & (g387) & (g327) & (!g332)) + ((g384) & (!g385) & (g386) & (!g387) & (!g327) & (!g332)) + ((g384) & (!g385) & (g386) & (!g387) & (g327) & (!g332)) + ((g384) & (!g385) & (g386) & (!g387) & (g327) & (g332)) + ((g384) & (!g385) & (g386) & (g387) & (!g327) & (!g332)) + ((g384) & (!g385) & (g386) & (g387) & (g327) & (!g332)) + ((g384) & (g385) & (!g386) & (!g387) & (!g327) & (!g332)) + ((g384) & (g385) & (!g386) & (!g387) & (!g327) & (g332)) + ((g384) & (g385) & (!g386) & (!g387) & (g327) & (g332)) + ((g384) & (g385) & (!g386) & (g387) & (!g327) & (!g332)) + ((g384) & (g385) & (!g386) & (g387) & (!g327) & (g332)) + ((g384) & (g385) & (g386) & (!g387) & (!g327) & (!g332)) + ((g384) & (g385) & (g386) & (!g387) & (g327) & (g332)) + ((g384) & (g385) & (g386) & (g387) & (!g327) & (!g332)));
	assign g390 = (((!g388) & (sk[64]) & (g389)) + ((g388) & (!sk[64]) & (!g389)) + ((g388) & (!sk[64]) & (g389)) + ((g388) & (sk[64]) & (!g389)));
	assign g397 = (((!g391) & (!g392) & (!g393) & (!g394) & (g395) & (g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g395) & (!g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g395) & (g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (g395) & (!g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (!g395) & (!g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (!g395) & (g396)) + ((!g391) & (!g392) & (g393) & (g394) & (!g395) & (!g396)) + ((!g391) & (!g392) & (g393) & (g394) & (g395) & (g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (g395) & (!g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (g395) & (g396)) + ((!g391) & (g392) & (!g393) & (g394) & (g395) & (!g396)) + ((!g391) & (g392) & (!g393) & (g394) & (g395) & (g396)) + ((!g391) & (g392) & (g393) & (!g394) & (g395) & (!g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (!g395) & (!g396)) + ((g391) & (!g392) & (g393) & (!g394) & (g395) & (!g396)) + ((g391) & (!g392) & (g393) & (g394) & (!g395) & (g396)) + ((g391) & (!g392) & (g393) & (g394) & (g395) & (g396)) + ((g391) & (g392) & (!g393) & (!g394) & (!g395) & (g396)) + ((g391) & (g392) & (!g393) & (!g394) & (g395) & (!g396)) + ((g391) & (g392) & (g393) & (!g394) & (!g395) & (g396)) + ((g391) & (g392) & (g393) & (!g394) & (g395) & (!g396)) + ((g391) & (g392) & (g393) & (g394) & (!g395) & (!g396)) + ((g391) & (g392) & (g393) & (g394) & (g395) & (!g396)) + ((g391) & (g392) & (g393) & (g394) & (g395) & (g396)));
	assign g398 = (((!g391) & (!g392) & (!g393) & (!g394) & (g395) & (!g396)) + ((!g391) & (!g392) & (!g393) & (!g394) & (g395) & (g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g395) & (!g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g395) & (g396)) + ((!g391) & (!g392) & (g393) & (g394) & (!g395) & (g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (!g395) & (!g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (!g395) & (g396)) + ((!g391) & (g392) & (g393) & (!g394) & (!g395) & (!g396)) + ((!g391) & (g392) & (g393) & (!g394) & (!g395) & (g396)) + ((!g391) & (g392) & (g393) & (!g394) & (g395) & (!g396)) + ((!g391) & (g392) & (g393) & (g394) & (g395) & (g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (!g395) & (g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (g395) & (!g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (g395) & (g396)) + ((g391) & (!g392) & (!g393) & (g394) & (g395) & (!g396)) + ((g391) & (!g392) & (g393) & (!g394) & (!g395) & (!g396)) + ((g391) & (!g392) & (g393) & (!g394) & (g395) & (g396)) + ((g391) & (!g392) & (g393) & (g394) & (!g395) & (g396)) + ((g391) & (!g392) & (g393) & (g394) & (g395) & (g396)) + ((g391) & (g392) & (!g393) & (!g394) & (!g395) & (!g396)) + ((g391) & (g392) & (!g393) & (!g394) & (!g395) & (g396)) + ((g391) & (g392) & (!g393) & (!g394) & (g395) & (!g396)) + ((g391) & (g392) & (!g393) & (!g394) & (g395) & (g396)) + ((g391) & (g392) & (!g393) & (g394) & (!g395) & (!g396)) + ((g391) & (g392) & (!g393) & (g394) & (g395) & (!g396)) + ((g391) & (g392) & (!g393) & (g394) & (g395) & (g396)) + ((g391) & (g392) & (g393) & (!g394) & (g395) & (!g396)) + ((g391) & (g392) & (g393) & (!g394) & (g395) & (g396)) + ((g391) & (g392) & (g393) & (g394) & (!g395) & (g396)) + ((g391) & (g392) & (g393) & (g394) & (g395) & (!g396)));
	assign g399 = (((!g391) & (!g392) & (!g393) & (!g394) & (!g395) & (!g396)) + ((!g391) & (!g392) & (!g393) & (!g394) & (g395) & (g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (g395) & (g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (!g395) & (!g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (!g395) & (g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (g395) & (g396)) + ((!g391) & (!g392) & (g393) & (g394) & (!g395) & (g396)) + ((!g391) & (!g392) & (g393) & (g394) & (g395) & (!g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (!g395) & (!g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (g395) & (!g396)) + ((!g391) & (g392) & (!g393) & (g394) & (g395) & (g396)) + ((!g391) & (g392) & (g393) & (g394) & (!g395) & (!g396)) + ((!g391) & (g392) & (g393) & (g394) & (g395) & (!g396)) + ((g391) & (!g392) & (!g393) & (g394) & (!g395) & (!g396)) + ((g391) & (!g392) & (!g393) & (g394) & (!g395) & (g396)) + ((g391) & (!g392) & (!g393) & (g394) & (g395) & (!g396)) + ((g391) & (!g392) & (g393) & (!g394) & (!g395) & (!g396)) + ((g391) & (!g392) & (g393) & (!g394) & (g395) & (g396)) + ((g391) & (!g392) & (g393) & (g394) & (!g395) & (!g396)) + ((g391) & (!g392) & (g393) & (g394) & (!g395) & (g396)) + ((g391) & (!g392) & (g393) & (g394) & (g395) & (!g396)) + ((g391) & (!g392) & (g393) & (g394) & (g395) & (g396)) + ((g391) & (g392) & (!g393) & (!g394) & (g395) & (g396)) + ((g391) & (g392) & (!g393) & (g394) & (!g395) & (!g396)) + ((g391) & (g392) & (!g393) & (g394) & (g395) & (!g396)) + ((g391) & (g392) & (!g393) & (g394) & (g395) & (g396)) + ((g391) & (g392) & (g393) & (!g394) & (!g395) & (!g396)) + ((g391) & (g392) & (g393) & (g394) & (!g395) & (!g396)) + ((g391) & (g392) & (g393) & (g394) & (!g395) & (g396)) + ((g391) & (g392) & (g393) & (g394) & (g395) & (g396)));
	assign g400 = (((!g391) & (!g392) & (!g393) & (!g394) & (!g395) & (g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (g395) & (!g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (g395) & (g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (!g395) & (g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (g395) & (g396)) + ((!g391) & (!g392) & (g393) & (g394) & (!g395) & (g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (!g395) & (!g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (!g395) & (g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (g395) & (!g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (g395) & (g396)) + ((!g391) & (g392) & (!g393) & (g394) & (g395) & (!g396)) + ((!g391) & (g392) & (!g393) & (g394) & (g395) & (g396)) + ((!g391) & (g392) & (g393) & (g394) & (!g395) & (!g396)) + ((!g391) & (g392) & (g393) & (g394) & (g395) & (!g396)) + ((!g391) & (g392) & (g393) & (g394) & (g395) & (g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (!g395) & (!g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (g395) & (g396)) + ((g391) & (!g392) & (!g393) & (g394) & (g395) & (!g396)) + ((g391) & (!g392) & (!g393) & (g394) & (g395) & (g396)) + ((g391) & (!g392) & (g393) & (!g394) & (!g395) & (g396)) + ((g391) & (!g392) & (g393) & (!g394) & (g395) & (!g396)) + ((g391) & (!g392) & (g393) & (g394) & (g395) & (!g396)) + ((g391) & (g392) & (!g393) & (!g394) & (!g395) & (g396)) + ((g391) & (g392) & (!g393) & (!g394) & (g395) & (g396)) + ((g391) & (g392) & (!g393) & (g394) & (g395) & (!g396)) + ((g391) & (g392) & (!g393) & (g394) & (g395) & (g396)) + ((g391) & (g392) & (g393) & (!g394) & (!g395) & (g396)) + ((g391) & (g392) & (g393) & (g394) & (!g395) & (!g396)));
	assign g403 = (((!g397) & (!g398) & (!g399) & (!g400) & (!g401) & (!g402)) + ((!g397) & (!g398) & (!g399) & (g400) & (!g401) & (!g402)) + ((!g397) & (!g398) & (!g399) & (g400) & (g401) & (g402)) + ((!g397) & (!g398) & (g399) & (!g400) & (!g401) & (!g402)) + ((!g397) & (!g398) & (g399) & (!g400) & (!g401) & (g402)) + ((!g397) & (!g398) & (g399) & (g400) & (!g401) & (!g402)) + ((!g397) & (!g398) & (g399) & (g400) & (!g401) & (g402)) + ((!g397) & (!g398) & (g399) & (g400) & (g401) & (g402)) + ((!g397) & (g398) & (!g399) & (!g400) & (!g401) & (!g402)) + ((!g397) & (g398) & (!g399) & (!g400) & (g401) & (!g402)) + ((!g397) & (g398) & (!g399) & (g400) & (!g401) & (!g402)) + ((!g397) & (g398) & (!g399) & (g400) & (g401) & (!g402)) + ((!g397) & (g398) & (!g399) & (g400) & (g401) & (g402)) + ((!g397) & (g398) & (g399) & (!g400) & (!g401) & (!g402)) + ((!g397) & (g398) & (g399) & (!g400) & (!g401) & (g402)) + ((!g397) & (g398) & (g399) & (!g400) & (g401) & (!g402)) + ((!g397) & (g398) & (g399) & (g400) & (!g401) & (!g402)) + ((!g397) & (g398) & (g399) & (g400) & (!g401) & (g402)) + ((!g397) & (g398) & (g399) & (g400) & (g401) & (!g402)) + ((!g397) & (g398) & (g399) & (g400) & (g401) & (g402)) + ((g397) & (!g398) & (!g399) & (g400) & (g401) & (g402)) + ((g397) & (!g398) & (g399) & (!g400) & (!g401) & (g402)) + ((g397) & (!g398) & (g399) & (g400) & (!g401) & (g402)) + ((g397) & (!g398) & (g399) & (g400) & (g401) & (g402)) + ((g397) & (g398) & (!g399) & (!g400) & (g401) & (!g402)) + ((g397) & (g398) & (!g399) & (g400) & (g401) & (!g402)) + ((g397) & (g398) & (!g399) & (g400) & (g401) & (g402)) + ((g397) & (g398) & (g399) & (!g400) & (!g401) & (g402)) + ((g397) & (g398) & (g399) & (!g400) & (g401) & (!g402)) + ((g397) & (g398) & (g399) & (g400) & (!g401) & (g402)) + ((g397) & (g398) & (g399) & (g400) & (g401) & (!g402)) + ((g397) & (g398) & (g399) & (g400) & (g401) & (g402)));
	assign g405 = (((!sk[70]) & (g403) & (!g404)) + ((!sk[70]) & (g403) & (g404)) + ((sk[70]) & (!g403) & (g404)) + ((sk[70]) & (g403) & (!g404)));
	assign g406 = (((!g391) & (!g392) & (!g393) & (!g394) & (!g401) & (g395)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g401) & (!g395)) + ((!g391) & (!g392) & (!g393) & (g394) & (g401) & (!g395)) + ((!g391) & (!g392) & (g393) & (!g394) & (g401) & (g395)) + ((!g391) & (!g392) & (g393) & (g394) & (!g401) & (g395)) + ((!g391) & (!g392) & (g393) & (g394) & (g401) & (!g395)) + ((!g391) & (g392) & (!g393) & (!g394) & (!g401) & (g395)) + ((!g391) & (g392) & (!g393) & (!g394) & (g401) & (!g395)) + ((!g391) & (g392) & (!g393) & (!g394) & (g401) & (g395)) + ((!g391) & (g392) & (g393) & (!g394) & (g401) & (g395)) + ((!g391) & (g392) & (g393) & (g394) & (g401) & (g395)) + ((g391) & (!g392) & (!g393) & (!g394) & (!g401) & (!g395)) + ((g391) & (!g392) & (!g393) & (!g394) & (g401) & (g395)) + ((g391) & (!g392) & (!g393) & (g394) & (!g401) & (!g395)) + ((g391) & (!g392) & (!g393) & (g394) & (g401) & (!g395)) + ((g391) & (!g392) & (g393) & (!g394) & (g401) & (!g395)) + ((g391) & (!g392) & (g393) & (!g394) & (g401) & (g395)) + ((g391) & (!g392) & (g393) & (g394) & (g401) & (!g395)) + ((g391) & (!g392) & (g393) & (g394) & (g401) & (g395)) + ((g391) & (g392) & (!g393) & (!g394) & (g401) & (!g395)) + ((g391) & (g392) & (!g393) & (!g394) & (g401) & (g395)) + ((g391) & (g392) & (!g393) & (g394) & (g401) & (g395)) + ((g391) & (g392) & (g393) & (!g394) & (!g401) & (!g395)) + ((g391) & (g392) & (g393) & (!g394) & (!g401) & (g395)) + ((g391) & (g392) & (g393) & (!g394) & (g401) & (!g395)) + ((g391) & (g392) & (g393) & (g394) & (!g401) & (g395)) + ((g391) & (g392) & (g393) & (g394) & (g401) & (!g395)));
	assign g407 = (((!g391) & (!g392) & (!g393) & (!g394) & (!g401) & (g395)) + ((!g391) & (!g392) & (!g393) & (!g394) & (g401) & (!g395)) + ((!g391) & (!g392) & (!g393) & (!g394) & (g401) & (g395)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g401) & (!g395)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g401) & (g395)) + ((!g391) & (!g392) & (!g393) & (g394) & (g401) & (g395)) + ((!g391) & (!g392) & (g393) & (!g394) & (g401) & (!g395)) + ((!g391) & (!g392) & (g393) & (g394) & (!g401) & (!g395)) + ((!g391) & (!g392) & (g393) & (g394) & (!g401) & (g395)) + ((!g391) & (!g392) & (g393) & (g394) & (g401) & (g395)) + ((!g391) & (g392) & (!g393) & (!g394) & (g401) & (g395)) + ((!g391) & (g392) & (!g393) & (g394) & (!g401) & (!g395)) + ((!g391) & (g392) & (!g393) & (g394) & (g401) & (!g395)) + ((!g391) & (g392) & (g393) & (!g394) & (g401) & (!g395)) + ((!g391) & (g392) & (g393) & (!g394) & (g401) & (g395)) + ((!g391) & (g392) & (g393) & (g394) & (!g401) & (!g395)) + ((g391) & (!g392) & (!g393) & (!g394) & (!g401) & (!g395)) + ((g391) & (!g392) & (!g393) & (g394) & (!g401) & (!g395)) + ((g391) & (!g392) & (!g393) & (g394) & (!g401) & (g395)) + ((g391) & (!g392) & (g393) & (!g394) & (!g401) & (g395)) + ((g391) & (!g392) & (g393) & (!g394) & (g401) & (g395)) + ((g391) & (!g392) & (g393) & (g394) & (!g401) & (!g395)) + ((g391) & (!g392) & (g393) & (g394) & (!g401) & (g395)) + ((g391) & (g392) & (!g393) & (g394) & (!g401) & (!g395)) + ((g391) & (g392) & (!g393) & (g394) & (g401) & (g395)) + ((g391) & (g392) & (g393) & (!g394) & (!g401) & (!g395)) + ((g391) & (g392) & (g393) & (!g394) & (!g401) & (g395)) + ((g391) & (g392) & (g393) & (!g394) & (g401) & (g395)) + ((g391) & (g392) & (g393) & (g394) & (!g401) & (!g395)) + ((g391) & (g392) & (g393) & (g394) & (!g401) & (g395)) + ((g391) & (g392) & (g393) & (g394) & (g401) & (!g395)));
	assign g408 = (((!g391) & (!g392) & (!g393) & (!g394) & (!g401) & (g395)) + ((!g391) & (!g392) & (!g393) & (g394) & (g401) & (!g395)) + ((!g391) & (!g392) & (g393) & (!g394) & (!g401) & (!g395)) + ((!g391) & (!g392) & (g393) & (!g394) & (g401) & (!g395)) + ((!g391) & (!g392) & (g393) & (g394) & (!g401) & (g395)) + ((!g391) & (!g392) & (g393) & (g394) & (g401) & (!g395)) + ((!g391) & (!g392) & (g393) & (g394) & (g401) & (g395)) + ((!g391) & (g392) & (!g393) & (!g394) & (!g401) & (!g395)) + ((!g391) & (g392) & (!g393) & (!g394) & (g401) & (!g395)) + ((!g391) & (g392) & (!g393) & (g394) & (!g401) & (!g395)) + ((!g391) & (g392) & (!g393) & (g394) & (g401) & (g395)) + ((!g391) & (g392) & (g393) & (!g394) & (g401) & (g395)) + ((!g391) & (g392) & (g393) & (g394) & (!g401) & (g395)) + ((!g391) & (g392) & (g393) & (g394) & (g401) & (!g395)) + ((g391) & (!g392) & (!g393) & (!g394) & (g401) & (g395)) + ((g391) & (!g392) & (!g393) & (g394) & (!g401) & (!g395)) + ((g391) & (!g392) & (!g393) & (g394) & (g401) & (!g395)) + ((g391) & (!g392) & (g393) & (!g394) & (!g401) & (!g395)) + ((g391) & (!g392) & (g393) & (!g394) & (!g401) & (g395)) + ((g391) & (!g392) & (g393) & (!g394) & (g401) & (!g395)) + ((g391) & (!g392) & (g393) & (!g394) & (g401) & (g395)) + ((g391) & (!g392) & (g393) & (g394) & (g401) & (!g395)) + ((g391) & (g392) & (!g393) & (!g394) & (!g401) & (g395)) + ((g391) & (g392) & (!g393) & (!g394) & (g401) & (g395)) + ((g391) & (g392) & (!g393) & (g394) & (!g401) & (g395)) + ((g391) & (g392) & (g393) & (!g394) & (!g401) & (!g395)) + ((g391) & (g392) & (g393) & (!g394) & (!g401) & (g395)) + ((g391) & (g392) & (g393) & (!g394) & (g401) & (g395)) + ((g391) & (g392) & (g393) & (g394) & (!g401) & (!g395)) + ((g391) & (g392) & (g393) & (g394) & (!g401) & (g395)) + ((g391) & (g392) & (g393) & (g394) & (g401) & (!g395)) + ((g391) & (g392) & (g393) & (g394) & (g401) & (g395)));
	assign g409 = (((!g391) & (!g392) & (!g393) & (!g394) & (g401) & (!g395)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g401) & (!g395)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g401) & (g395)) + ((!g391) & (!g392) & (g393) & (!g394) & (g401) & (g395)) + ((!g391) & (!g392) & (g393) & (g394) & (!g401) & (g395)) + ((!g391) & (g392) & (!g393) & (!g394) & (!g401) & (!g395)) + ((!g391) & (g392) & (!g393) & (!g394) & (g401) & (!g395)) + ((!g391) & (g392) & (!g393) & (g394) & (!g401) & (g395)) + ((!g391) & (g392) & (g393) & (!g394) & (!g401) & (g395)) + ((!g391) & (g392) & (g393) & (!g394) & (g401) & (!g395)) + ((!g391) & (g392) & (g393) & (!g394) & (g401) & (g395)) + ((!g391) & (g392) & (g393) & (g394) & (g401) & (!g395)) + ((!g391) & (g392) & (g393) & (g394) & (g401) & (g395)) + ((g391) & (!g392) & (!g393) & (!g394) & (!g401) & (!g395)) + ((g391) & (!g392) & (!g393) & (g394) & (!g401) & (!g395)) + ((g391) & (!g392) & (!g393) & (g394) & (!g401) & (g395)) + ((g391) & (!g392) & (!g393) & (g394) & (g401) & (!g395)) + ((g391) & (!g392) & (g393) & (!g394) & (!g401) & (!g395)) + ((g391) & (!g392) & (g393) & (!g394) & (g401) & (g395)) + ((g391) & (!g392) & (g393) & (g394) & (g401) & (!g395)) + ((g391) & (g392) & (!g393) & (!g394) & (!g401) & (!g395)) + ((g391) & (g392) & (!g393) & (g394) & (!g401) & (!g395)) + ((g391) & (g392) & (!g393) & (g394) & (g401) & (!g395)) + ((g391) & (g392) & (!g393) & (g394) & (g401) & (g395)) + ((g391) & (g392) & (g393) & (g394) & (!g401) & (g395)) + ((g391) & (g392) & (g393) & (g394) & (g401) & (g395)));
	assign g410 = (((!g406) & (!g407) & (!g408) & (!g409) & (!g396) & (!g402)) + ((!g406) & (!g407) & (!g408) & (!g409) & (g396) & (!g402)) + ((!g406) & (!g407) & (!g408) & (g409) & (!g396) & (!g402)) + ((!g406) & (!g407) & (!g408) & (g409) & (g396) & (!g402)) + ((!g406) & (!g407) & (!g408) & (g409) & (g396) & (g402)) + ((!g406) & (!g407) & (g408) & (!g409) & (!g396) & (!g402)) + ((!g406) & (!g407) & (g408) & (!g409) & (!g396) & (g402)) + ((!g406) & (!g407) & (g408) & (!g409) & (g396) & (!g402)) + ((!g406) & (!g407) & (g408) & (g409) & (!g396) & (!g402)) + ((!g406) & (!g407) & (g408) & (g409) & (!g396) & (g402)) + ((!g406) & (!g407) & (g408) & (g409) & (g396) & (!g402)) + ((!g406) & (!g407) & (g408) & (g409) & (g396) & (g402)) + ((!g406) & (g407) & (!g408) & (!g409) & (!g396) & (!g402)) + ((!g406) & (g407) & (!g408) & (g409) & (!g396) & (!g402)) + ((!g406) & (g407) & (!g408) & (g409) & (g396) & (g402)) + ((!g406) & (g407) & (g408) & (!g409) & (!g396) & (!g402)) + ((!g406) & (g407) & (g408) & (!g409) & (!g396) & (g402)) + ((!g406) & (g407) & (g408) & (g409) & (!g396) & (!g402)) + ((!g406) & (g407) & (g408) & (g409) & (!g396) & (g402)) + ((!g406) & (g407) & (g408) & (g409) & (g396) & (g402)) + ((g406) & (!g407) & (!g408) & (!g409) & (g396) & (!g402)) + ((g406) & (!g407) & (!g408) & (g409) & (g396) & (!g402)) + ((g406) & (!g407) & (!g408) & (g409) & (g396) & (g402)) + ((g406) & (!g407) & (g408) & (!g409) & (!g396) & (g402)) + ((g406) & (!g407) & (g408) & (!g409) & (g396) & (!g402)) + ((g406) & (!g407) & (g408) & (g409) & (!g396) & (g402)) + ((g406) & (!g407) & (g408) & (g409) & (g396) & (!g402)) + ((g406) & (!g407) & (g408) & (g409) & (g396) & (g402)) + ((g406) & (g407) & (!g408) & (g409) & (g396) & (g402)) + ((g406) & (g407) & (g408) & (!g409) & (!g396) & (g402)) + ((g406) & (g407) & (g408) & (g409) & (!g396) & (g402)) + ((g406) & (g407) & (g408) & (g409) & (g396) & (g402)));
	assign g412 = (((!g410) & (sk[76]) & (g411)) + ((g410) & (!sk[76]) & (!g411)) + ((g410) & (!sk[76]) & (g411)) + ((g410) & (sk[76]) & (!g411)));
	assign g413 = (((!g395) & (!g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((!g395) & (!g392) & (!g393) & (!g394) & (g401) & (g396)) + ((!g395) & (!g392) & (!g393) & (g394) & (!g401) & (g396)) + ((!g395) & (!g392) & (!g393) & (g394) & (g401) & (!g396)) + ((!g395) & (!g392) & (!g393) & (g394) & (g401) & (g396)) + ((!g395) & (!g392) & (g393) & (!g394) & (!g401) & (g396)) + ((!g395) & (!g392) & (g393) & (g394) & (!g401) & (!g396)) + ((!g395) & (!g392) & (g393) & (g394) & (g401) & (!g396)) + ((!g395) & (g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((!g395) & (g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((!g395) & (g392) & (!g393) & (g394) & (!g401) & (g396)) + ((!g395) & (g392) & (g393) & (!g394) & (!g401) & (!g396)) + ((!g395) & (g392) & (g393) & (!g394) & (!g401) & (g396)) + ((!g395) & (g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g395) & (g392) & (g393) & (!g394) & (g401) & (g396)) + ((g395) & (!g392) & (!g393) & (g394) & (!g401) & (g396)) + ((g395) & (!g392) & (!g393) & (g394) & (g401) & (g396)) + ((g395) & (g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((g395) & (g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((g395) & (g392) & (!g393) & (g394) & (g401) & (!g396)) + ((g395) & (g392) & (g393) & (g394) & (!g401) & (!g396)) + ((g395) & (g392) & (g393) & (g394) & (!g401) & (g396)));
	assign g414 = (((!g395) & (!g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((!g395) & (!g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((!g395) & (!g392) & (!g393) & (g394) & (g401) & (g396)) + ((!g395) & (!g392) & (g393) & (!g394) & (!g401) & (!g396)) + ((!g395) & (!g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g395) & (!g392) & (g393) & (g394) & (!g401) & (g396)) + ((!g395) & (g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((!g395) & (g392) & (!g393) & (!g394) & (g401) & (g396)) + ((!g395) & (g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((!g395) & (g392) & (!g393) & (g394) & (!g401) & (g396)) + ((!g395) & (g392) & (!g393) & (g394) & (g401) & (g396)) + ((!g395) & (g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g395) & (g392) & (g393) & (!g394) & (g401) & (g396)) + ((!g395) & (g392) & (g393) & (g394) & (g401) & (!g396)) + ((g395) & (!g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((g395) & (!g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((g395) & (!g392) & (!g393) & (!g394) & (g401) & (g396)) + ((g395) & (!g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((g395) & (!g392) & (!g393) & (g394) & (!g401) & (g396)) + ((g395) & (!g392) & (!g393) & (g394) & (g401) & (!g396)) + ((g395) & (!g392) & (g393) & (g394) & (!g401) & (!g396)) + ((g395) & (g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((g395) & (g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((g395) & (g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((g395) & (g392) & (!g393) & (g394) & (g401) & (!g396)) + ((g395) & (g392) & (!g393) & (g394) & (g401) & (g396)) + ((g395) & (g392) & (g393) & (!g394) & (!g401) & (!g396)) + ((g395) & (g392) & (g393) & (!g394) & (g401) & (!g396)) + ((g395) & (g392) & (g393) & (g394) & (!g401) & (g396)) + ((g395) & (g392) & (g393) & (g394) & (g401) & (g396)));
	assign g415 = (((!g395) & (!g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((!g395) & (!g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((!g395) & (!g392) & (!g393) & (g394) & (!g401) & (g396)) + ((!g395) & (!g392) & (g393) & (!g394) & (!g401) & (g396)) + ((!g395) & (!g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g395) & (!g392) & (g393) & (g394) & (!g401) & (g396)) + ((!g395) & (g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((!g395) & (g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((!g395) & (g392) & (!g393) & (g394) & (g401) & (!g396)) + ((!g395) & (g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g395) & (g392) & (g393) & (g394) & (!g401) & (!g396)) + ((!g395) & (g392) & (g393) & (g394) & (g401) & (!g396)) + ((g395) & (!g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((g395) & (!g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((g395) & (!g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((g395) & (!g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((g395) & (!g392) & (!g393) & (g394) & (!g401) & (g396)) + ((g395) & (!g392) & (!g393) & (g394) & (g401) & (!g396)) + ((g395) & (!g392) & (!g393) & (g394) & (g401) & (g396)) + ((g395) & (!g392) & (g393) & (!g394) & (!g401) & (g396)) + ((g395) & (!g392) & (g393) & (!g394) & (g401) & (!g396)) + ((g395) & (!g392) & (g393) & (g394) & (!g401) & (!g396)) + ((g395) & (!g392) & (g393) & (g394) & (g401) & (g396)) + ((g395) & (g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((g395) & (g392) & (!g393) & (!g394) & (g401) & (g396)) + ((g395) & (g392) & (g393) & (!g394) & (g401) & (g396)) + ((g395) & (g392) & (g393) & (g394) & (!g401) & (!g396)) + ((g395) & (g392) & (g393) & (g394) & (!g401) & (g396)) + ((g395) & (g392) & (g393) & (g394) & (g401) & (g396)));
	assign g416 = (((!g395) & (!g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((!g395) & (!g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((!g395) & (!g392) & (!g393) & (!g394) & (g401) & (g396)) + ((!g395) & (!g392) & (!g393) & (g394) & (!g401) & (g396)) + ((!g395) & (!g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g395) & (!g392) & (g393) & (g394) & (g401) & (g396)) + ((!g395) & (g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((!g395) & (g392) & (!g393) & (g394) & (!g401) & (g396)) + ((!g395) & (g392) & (!g393) & (g394) & (g401) & (g396)) + ((!g395) & (g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g395) & (g392) & (g393) & (!g394) & (g401) & (g396)) + ((!g395) & (g392) & (g393) & (g394) & (!g401) & (!g396)) + ((!g395) & (g392) & (g393) & (g394) & (!g401) & (g396)) + ((!g395) & (g392) & (g393) & (g394) & (g401) & (!g396)) + ((!g395) & (g392) & (g393) & (g394) & (g401) & (g396)) + ((g395) & (!g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((g395) & (!g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((g395) & (!g392) & (!g393) & (!g394) & (g401) & (g396)) + ((g395) & (!g392) & (!g393) & (g394) & (g401) & (g396)) + ((g395) & (!g392) & (g393) & (!g394) & (!g401) & (g396)) + ((g395) & (!g392) & (g393) & (!g394) & (g401) & (!g396)) + ((g395) & (!g392) & (g393) & (g394) & (g401) & (!g396)) + ((g395) & (g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((g395) & (g392) & (!g393) & (g394) & (!g401) & (g396)) + ((g395) & (g392) & (!g393) & (g394) & (g401) & (!g396)) + ((g395) & (g392) & (g393) & (!g394) & (g401) & (g396)) + ((g395) & (g392) & (g393) & (g394) & (!g401) & (!g396)));
	assign g417 = (((!g413) & (!g414) & (!g415) & (!g416) & (!g391) & (g402)) + ((!g413) & (!g414) & (!g415) & (!g416) & (g391) & (!g402)) + ((!g413) & (!g414) & (!g415) & (!g416) & (g391) & (g402)) + ((!g413) & (!g414) & (!g415) & (g416) & (!g391) & (g402)) + ((!g413) & (!g414) & (!g415) & (g416) & (g391) & (!g402)) + ((!g413) & (!g414) & (g415) & (!g416) & (g391) & (!g402)) + ((!g413) & (!g414) & (g415) & (!g416) & (g391) & (g402)) + ((!g413) & (!g414) & (g415) & (g416) & (g391) & (!g402)) + ((!g413) & (g414) & (!g415) & (!g416) & (!g391) & (g402)) + ((!g413) & (g414) & (!g415) & (!g416) & (g391) & (g402)) + ((!g413) & (g414) & (!g415) & (g416) & (!g391) & (g402)) + ((!g413) & (g414) & (g415) & (!g416) & (g391) & (g402)) + ((g413) & (!g414) & (!g415) & (!g416) & (!g391) & (!g402)) + ((g413) & (!g414) & (!g415) & (!g416) & (!g391) & (g402)) + ((g413) & (!g414) & (!g415) & (!g416) & (g391) & (!g402)) + ((g413) & (!g414) & (!g415) & (!g416) & (g391) & (g402)) + ((g413) & (!g414) & (!g415) & (g416) & (!g391) & (!g402)) + ((g413) & (!g414) & (!g415) & (g416) & (!g391) & (g402)) + ((g413) & (!g414) & (!g415) & (g416) & (g391) & (!g402)) + ((g413) & (!g414) & (g415) & (!g416) & (!g391) & (!g402)) + ((g413) & (!g414) & (g415) & (!g416) & (g391) & (!g402)) + ((g413) & (!g414) & (g415) & (!g416) & (g391) & (g402)) + ((g413) & (!g414) & (g415) & (g416) & (!g391) & (!g402)) + ((g413) & (!g414) & (g415) & (g416) & (g391) & (!g402)) + ((g413) & (g414) & (!g415) & (!g416) & (!g391) & (!g402)) + ((g413) & (g414) & (!g415) & (!g416) & (!g391) & (g402)) + ((g413) & (g414) & (!g415) & (!g416) & (g391) & (g402)) + ((g413) & (g414) & (!g415) & (g416) & (!g391) & (!g402)) + ((g413) & (g414) & (!g415) & (g416) & (!g391) & (g402)) + ((g413) & (g414) & (g415) & (!g416) & (!g391) & (!g402)) + ((g413) & (g414) & (g415) & (!g416) & (g391) & (g402)) + ((g413) & (g414) & (g415) & (g416) & (!g391) & (!g402)));
	assign g419 = (((!sk[82]) & (g417) & (!g418)) + ((!sk[82]) & (g417) & (g418)) + ((sk[82]) & (!g417) & (g418)) + ((sk[82]) & (g417) & (!g418)));
	assign g420 = (((!g391) & (!g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (g401) & (g396)) + ((!g391) & (!g392) & (g393) & (g394) & (!g401) & (!g396)) + ((!g391) & (!g392) & (g393) & (g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (g393) & (g394) & (g401) & (g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (g392) & (g393) & (!g394) & (!g401) & (!g396)) + ((!g391) & (g392) & (g393) & (g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((g391) & (!g392) & (g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (g393) & (!g394) & (!g401) & (g396)) + ((g391) & (!g392) & (g393) & (!g394) & (g401) & (!g396)) + ((g391) & (!g392) & (g393) & (g394) & (!g401) & (g396)) + ((g391) & (g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((g391) & (g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((g391) & (g392) & (!g393) & (g394) & (g401) & (!g396)) + ((g391) & (g392) & (g393) & (!g394) & (!g401) & (g396)) + ((g391) & (g392) & (g393) & (!g394) & (g401) & (g396)));
	assign g421 = (((!g391) & (!g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (!g393) & (!g394) & (g401) & (g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (g393) & (g394) & (!g401) & (!g396)) + ((!g391) & (!g392) & (g393) & (g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (g393) & (g394) & (g401) & (g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (g401) & (g396)) + ((!g391) & (g392) & (!g393) & (g394) & (g401) & (g396)) + ((!g391) & (g392) & (g393) & (!g394) & (!g401) & (!g396)) + ((!g391) & (g392) & (g393) & (!g394) & (!g401) & (g396)) + ((!g391) & (g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (g392) & (g393) & (g394) & (!g401) & (g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((g391) & (!g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (!g393) & (g394) & (!g401) & (g396)) + ((g391) & (!g392) & (!g393) & (g394) & (g401) & (g396)) + ((g391) & (!g392) & (g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (g393) & (!g394) & (!g401) & (g396)) + ((g391) & (!g392) & (g393) & (!g394) & (g401) & (g396)) + ((g391) & (!g392) & (g393) & (g394) & (!g401) & (g396)) + ((g391) & (g392) & (!g393) & (g394) & (!g401) & (g396)) + ((g391) & (g392) & (!g393) & (g394) & (g401) & (!g396)) + ((g391) & (g392) & (g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (g392) & (g393) & (g394) & (!g401) & (!g396)));
	assign g422 = (((!g391) & (!g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (!g393) & (!g394) & (g401) & (g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (g393) & (!g394) & (g401) & (g396)) + ((!g391) & (!g392) & (g393) & (g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (g393) & (g394) & (g401) & (g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (g401) & (g396)) + ((!g391) & (g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((!g391) & (g392) & (!g393) & (g394) & (!g401) & (g396)) + ((!g391) & (g392) & (g393) & (!g394) & (!g401) & (g396)) + ((!g391) & (g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (g392) & (g393) & (g394) & (g401) & (g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (g401) & (g396)) + ((g391) & (!g392) & (!g393) & (g394) & (g401) & (g396)) + ((g391) & (!g392) & (g393) & (g394) & (!g401) & (!g396)) + ((g391) & (g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((g391) & (g392) & (!g393) & (g394) & (g401) & (g396)) + ((g391) & (g392) & (g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (g392) & (g393) & (!g394) & (!g401) & (g396)) + ((g391) & (g392) & (g393) & (!g394) & (g401) & (g396)) + ((g391) & (g392) & (g393) & (g394) & (!g401) & (!g396)) + ((g391) & (g392) & (g393) & (g394) & (g401) & (g396)));
	assign g423 = (((!g391) & (!g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (!g393) & (g394) & (g401) & (g396)) + ((!g391) & (!g392) & (g393) & (g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (g393) & (g394) & (g401) & (g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (!g401) & (!g396)) + ((!g391) & (g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (g392) & (!g393) & (g394) & (!g401) & (!g396)) + ((!g391) & (g392) & (!g393) & (g394) & (!g401) & (g396)) + ((!g391) & (g392) & (!g393) & (g394) & (g401) & (!g396)) + ((!g391) & (g392) & (g393) & (!g394) & (!g401) & (!g396)) + ((!g391) & (g392) & (g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (g392) & (g393) & (!g394) & (g401) & (g396)) + ((g391) & (!g392) & (!g393) & (!g394) & (g401) & (g396)) + ((g391) & (!g392) & (!g393) & (g394) & (g401) & (!g396)) + ((g391) & (!g392) & (g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (g393) & (!g394) & (g401) & (!g396)) + ((g391) & (!g392) & (g393) & (!g394) & (g401) & (g396)) + ((g391) & (!g392) & (g393) & (g394) & (!g401) & (g396)) + ((g391) & (!g392) & (g393) & (g394) & (g401) & (!g396)) + ((g391) & (!g392) & (g393) & (g394) & (g401) & (g396)) + ((g391) & (g392) & (!g393) & (!g394) & (!g401) & (g396)) + ((g391) & (g392) & (!g393) & (!g394) & (g401) & (!g396)) + ((g391) & (g392) & (g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (g392) & (g393) & (!g394) & (!g401) & (g396)) + ((g391) & (g392) & (g393) & (g394) & (g401) & (g396)));
	assign g424 = (((!g420) & (!g421) & (!g422) & (!g423) & (!g402) & (g395)) + ((!g420) & (!g421) & (!g422) & (!g423) & (g402) & (!g395)) + ((!g420) & (!g421) & (!g422) & (!g423) & (g402) & (g395)) + ((!g420) & (!g421) & (!g422) & (g423) & (!g402) & (g395)) + ((!g420) & (!g421) & (!g422) & (g423) & (g402) & (!g395)) + ((!g420) & (!g421) & (g422) & (!g423) & (g402) & (!g395)) + ((!g420) & (!g421) & (g422) & (!g423) & (g402) & (g395)) + ((!g420) & (!g421) & (g422) & (g423) & (g402) & (!g395)) + ((!g420) & (g421) & (!g422) & (!g423) & (!g402) & (g395)) + ((!g420) & (g421) & (!g422) & (!g423) & (g402) & (g395)) + ((!g420) & (g421) & (!g422) & (g423) & (!g402) & (g395)) + ((!g420) & (g421) & (g422) & (!g423) & (g402) & (g395)) + ((g420) & (!g421) & (!g422) & (!g423) & (!g402) & (!g395)) + ((g420) & (!g421) & (!g422) & (!g423) & (!g402) & (g395)) + ((g420) & (!g421) & (!g422) & (!g423) & (g402) & (!g395)) + ((g420) & (!g421) & (!g422) & (!g423) & (g402) & (g395)) + ((g420) & (!g421) & (!g422) & (g423) & (!g402) & (!g395)) + ((g420) & (!g421) & (!g422) & (g423) & (!g402) & (g395)) + ((g420) & (!g421) & (!g422) & (g423) & (g402) & (!g395)) + ((g420) & (!g421) & (g422) & (!g423) & (!g402) & (!g395)) + ((g420) & (!g421) & (g422) & (!g423) & (g402) & (!g395)) + ((g420) & (!g421) & (g422) & (!g423) & (g402) & (g395)) + ((g420) & (!g421) & (g422) & (g423) & (!g402) & (!g395)) + ((g420) & (!g421) & (g422) & (g423) & (g402) & (!g395)) + ((g420) & (g421) & (!g422) & (!g423) & (!g402) & (!g395)) + ((g420) & (g421) & (!g422) & (!g423) & (!g402) & (g395)) + ((g420) & (g421) & (!g422) & (!g423) & (g402) & (g395)) + ((g420) & (g421) & (!g422) & (g423) & (!g402) & (!g395)) + ((g420) & (g421) & (!g422) & (g423) & (!g402) & (g395)) + ((g420) & (g421) & (g422) & (!g423) & (!g402) & (!g395)) + ((g420) & (g421) & (g422) & (!g423) & (g402) & (g395)) + ((g420) & (g421) & (g422) & (g423) & (!g402) & (!g395)));
	assign g426 = (((!g424) & (sk[88]) & (g425)) + ((g424) & (!sk[88]) & (!g425)) + ((g424) & (!sk[88]) & (g425)) + ((g424) & (sk[88]) & (!g425)));
	assign g427 = (((!g391) & (!g392) & (!g395) & (!g402) & (!g401) & (g396)) + ((!g391) & (!g392) & (g395) & (!g402) & (!g401) & (g396)) + ((!g391) & (!g392) & (g395) & (!g402) & (g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (!g402) & (g401) & (g396)) + ((!g391) & (!g392) & (g395) & (g402) & (!g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (g402) & (g401) & (!g396)) + ((!g391) & (g392) & (!g395) & (!g402) & (!g401) & (!g396)) + ((!g391) & (g392) & (!g395) & (!g402) & (!g401) & (g396)) + ((!g391) & (g392) & (!g395) & (g402) & (!g401) & (!g396)) + ((!g391) & (g392) & (!g395) & (g402) & (!g401) & (g396)) + ((!g391) & (g392) & (!g395) & (g402) & (g401) & (g396)) + ((!g391) & (g392) & (g395) & (g402) & (!g401) & (g396)) + ((!g391) & (g392) & (g395) & (g402) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g402) & (!g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g402) & (!g401) & (g396)) + ((g391) & (!g392) & (!g395) & (g402) & (!g401) & (g396)) + ((g391) & (!g392) & (g395) & (!g402) & (g401) & (!g396)) + ((g391) & (!g392) & (g395) & (g402) & (!g401) & (!g396)) + ((g391) & (!g392) & (g395) & (g402) & (!g401) & (g396)) + ((g391) & (!g392) & (g395) & (g402) & (g401) & (!g396)) + ((g391) & (g392) & (!g395) & (!g402) & (!g401) & (!g396)) + ((g391) & (g392) & (!g395) & (!g402) & (g401) & (!g396)) + ((g391) & (g392) & (!g395) & (g402) & (g401) & (!g396)) + ((g391) & (g392) & (g395) & (!g402) & (!g401) & (!g396)) + ((g391) & (g392) & (g395) & (!g402) & (!g401) & (g396)) + ((g391) & (g392) & (g395) & (g402) & (!g401) & (g396)));
	assign g428 = (((!g391) & (!g392) & (!g395) & (!g402) & (!g401) & (!g396)) + ((!g391) & (!g392) & (!g395) & (!g402) & (!g401) & (g396)) + ((!g391) & (!g392) & (!g395) & (!g402) & (g401) & (!g396)) + ((!g391) & (!g392) & (!g395) & (!g402) & (g401) & (g396)) + ((!g391) & (!g392) & (!g395) & (g402) & (!g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (!g402) & (!g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (!g402) & (g401) & (g396)) + ((!g391) & (!g392) & (g395) & (g402) & (!g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (g402) & (g401) & (g396)) + ((!g391) & (g392) & (!g395) & (!g402) & (!g401) & (g396)) + ((!g391) & (g392) & (!g395) & (g402) & (g401) & (!g396)) + ((!g391) & (g392) & (g395) & (!g402) & (!g401) & (!g396)) + ((!g391) & (g392) & (g395) & (!g402) & (!g401) & (g396)) + ((!g391) & (g392) & (g395) & (!g402) & (g401) & (!g396)) + ((!g391) & (g392) & (g395) & (!g402) & (g401) & (g396)) + ((!g391) & (g392) & (g395) & (g402) & (!g401) & (!g396)) + ((!g391) & (g392) & (g395) & (g402) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g402) & (!g401) & (g396)) + ((g391) & (!g392) & (!g395) & (!g402) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g402) & (g401) & (g396)) + ((g391) & (!g392) & (!g395) & (g402) & (!g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (g402) & (g401) & (g396)) + ((g391) & (!g392) & (g395) & (!g402) & (g401) & (!g396)) + ((g391) & (!g392) & (g395) & (!g402) & (g401) & (g396)) + ((g391) & (!g392) & (g395) & (g402) & (!g401) & (g396)) + ((g391) & (g392) & (!g395) & (!g402) & (g401) & (!g396)) + ((g391) & (g392) & (!g395) & (!g402) & (g401) & (g396)) + ((g391) & (g392) & (!g395) & (g402) & (!g401) & (!g396)) + ((g391) & (g392) & (!g395) & (g402) & (!g401) & (g396)) + ((g391) & (g392) & (g395) & (!g402) & (g401) & (!g396)) + ((g391) & (g392) & (g395) & (!g402) & (g401) & (g396)) + ((g391) & (g392) & (g395) & (g402) & (!g401) & (g396)));
	assign g429 = (((!g391) & (!g392) & (!g395) & (!g402) & (!g401) & (!g396)) + ((!g391) & (!g392) & (!g395) & (!g402) & (!g401) & (g396)) + ((!g391) & (!g392) & (g395) & (!g402) & (!g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (!g402) & (g401) & (g396)) + ((!g391) & (!g392) & (g395) & (g402) & (!g401) & (g396)) + ((!g391) & (g392) & (!g395) & (g402) & (!g401) & (!g396)) + ((!g391) & (g392) & (!g395) & (g402) & (g401) & (!g396)) + ((!g391) & (g392) & (!g395) & (g402) & (g401) & (g396)) + ((!g391) & (g392) & (g395) & (!g402) & (!g401) & (!g396)) + ((!g391) & (g392) & (g395) & (!g402) & (g401) & (!g396)) + ((!g391) & (g392) & (g395) & (!g402) & (g401) & (g396)) + ((!g391) & (g392) & (g395) & (g402) & (!g401) & (!g396)) + ((!g391) & (g392) & (g395) & (g402) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g402) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g402) & (g401) & (g396)) + ((g391) & (!g392) & (!g395) & (g402) & (!g401) & (g396)) + ((g391) & (!g392) & (!g395) & (g402) & (g401) & (g396)) + ((g391) & (!g392) & (g395) & (!g402) & (!g401) & (!g396)) + ((g391) & (!g392) & (g395) & (!g402) & (!g401) & (g396)) + ((g391) & (!g392) & (g395) & (!g402) & (g401) & (g396)) + ((g391) & (!g392) & (g395) & (g402) & (!g401) & (!g396)) + ((g391) & (!g392) & (g395) & (g402) & (!g401) & (g396)) + ((g391) & (!g392) & (g395) & (g402) & (g401) & (!g396)) + ((g391) & (!g392) & (g395) & (g402) & (g401) & (g396)) + ((g391) & (g392) & (!g395) & (!g402) & (!g401) & (g396)) + ((g391) & (g392) & (!g395) & (g402) & (!g401) & (!g396)) + ((g391) & (g392) & (!g395) & (g402) & (g401) & (!g396)) + ((g391) & (g392) & (g395) & (!g402) & (!g401) & (!g396)) + ((g391) & (g392) & (g395) & (!g402) & (!g401) & (g396)) + ((g391) & (g392) & (g395) & (!g402) & (g401) & (!g396)) + ((g391) & (g392) & (g395) & (g402) & (!g401) & (!g396)) + ((g391) & (g392) & (g395) & (g402) & (g401) & (!g396)));
	assign g430 = (((!g391) & (!g392) & (!g395) & (!g402) & (g401) & (g396)) + ((!g391) & (!g392) & (!g395) & (g402) & (!g401) & (!g396)) + ((!g391) & (!g392) & (!g395) & (g402) & (g401) & (g396)) + ((!g391) & (!g392) & (g395) & (!g402) & (!g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (!g402) & (g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (g402) & (!g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (g402) & (!g401) & (g396)) + ((!g391) & (!g392) & (g395) & (g402) & (g401) & (!g396)) + ((!g391) & (g392) & (!g395) & (!g402) & (!g401) & (!g396)) + ((!g391) & (g392) & (!g395) & (g402) & (!g401) & (g396)) + ((!g391) & (g392) & (!g395) & (g402) & (g401) & (!g396)) + ((!g391) & (g392) & (!g395) & (g402) & (g401) & (g396)) + ((!g391) & (g392) & (g395) & (!g402) & (!g401) & (!g396)) + ((!g391) & (g392) & (g395) & (g402) & (!g401) & (!g396)) + ((!g391) & (g392) & (g395) & (g402) & (!g401) & (g396)) + ((g391) & (!g392) & (!g395) & (!g402) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g402) & (g401) & (g396)) + ((g391) & (!g392) & (g395) & (!g402) & (!g401) & (!g396)) + ((g391) & (!g392) & (g395) & (!g402) & (g401) & (!g396)) + ((g391) & (!g392) & (g395) & (g402) & (g401) & (!g396)) + ((g391) & (g392) & (!g395) & (!g402) & (g401) & (!g396)) + ((g391) & (g392) & (!g395) & (g402) & (g401) & (g396)) + ((g391) & (g392) & (g395) & (!g402) & (!g401) & (!g396)) + ((g391) & (g392) & (g395) & (!g402) & (!g401) & (g396)) + ((g391) & (g392) & (g395) & (!g402) & (g401) & (!g396)) + ((g391) & (g392) & (g395) & (g402) & (!g401) & (!g396)));
	assign g431 = (((!g427) & (!g428) & (!g429) & (!g430) & (g393) & (g394)) + ((!g427) & (!g428) & (g429) & (!g430) & (!g393) & (g394)) + ((!g427) & (!g428) & (g429) & (!g430) & (g393) & (g394)) + ((!g427) & (!g428) & (g429) & (g430) & (!g393) & (g394)) + ((!g427) & (g428) & (!g429) & (!g430) & (g393) & (!g394)) + ((!g427) & (g428) & (!g429) & (!g430) & (g393) & (g394)) + ((!g427) & (g428) & (!g429) & (g430) & (g393) & (!g394)) + ((!g427) & (g428) & (g429) & (!g430) & (!g393) & (g394)) + ((!g427) & (g428) & (g429) & (!g430) & (g393) & (!g394)) + ((!g427) & (g428) & (g429) & (!g430) & (g393) & (g394)) + ((!g427) & (g428) & (g429) & (g430) & (!g393) & (g394)) + ((!g427) & (g428) & (g429) & (g430) & (g393) & (!g394)) + ((g427) & (!g428) & (!g429) & (!g430) & (!g393) & (!g394)) + ((g427) & (!g428) & (!g429) & (!g430) & (g393) & (g394)) + ((g427) & (!g428) & (!g429) & (g430) & (!g393) & (!g394)) + ((g427) & (!g428) & (g429) & (!g430) & (!g393) & (!g394)) + ((g427) & (!g428) & (g429) & (!g430) & (!g393) & (g394)) + ((g427) & (!g428) & (g429) & (!g430) & (g393) & (g394)) + ((g427) & (!g428) & (g429) & (g430) & (!g393) & (!g394)) + ((g427) & (!g428) & (g429) & (g430) & (!g393) & (g394)) + ((g427) & (g428) & (!g429) & (!g430) & (!g393) & (!g394)) + ((g427) & (g428) & (!g429) & (!g430) & (g393) & (!g394)) + ((g427) & (g428) & (!g429) & (!g430) & (g393) & (g394)) + ((g427) & (g428) & (!g429) & (g430) & (!g393) & (!g394)) + ((g427) & (g428) & (!g429) & (g430) & (g393) & (!g394)) + ((g427) & (g428) & (g429) & (!g430) & (!g393) & (!g394)) + ((g427) & (g428) & (g429) & (!g430) & (!g393) & (g394)) + ((g427) & (g428) & (g429) & (!g430) & (g393) & (!g394)) + ((g427) & (g428) & (g429) & (!g430) & (g393) & (g394)) + ((g427) & (g428) & (g429) & (g430) & (!g393) & (!g394)) + ((g427) & (g428) & (g429) & (g430) & (!g393) & (g394)) + ((g427) & (g428) & (g429) & (g430) & (g393) & (!g394)));
	assign g433 = (((!sk[94]) & (g431) & (!g432)) + ((!sk[94]) & (g431) & (g432)) + ((sk[94]) & (!g431) & (g432)) + ((sk[94]) & (g431) & (!g432)));
	assign g434 = (((!g391) & (!g392) & (!g395) & (!g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (!g395) & (!g394) & (g401) & (g396)) + ((!g391) & (!g392) & (!g395) & (g394) & (g401) & (g396)) + ((!g391) & (!g392) & (g395) & (!g394) & (!g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (!g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (g395) & (!g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (!g394) & (g401) & (g396)) + ((!g391) & (!g392) & (g395) & (g394) & (!g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (g394) & (!g401) & (g396)) + ((!g391) & (g392) & (!g395) & (!g394) & (!g401) & (g396)) + ((!g391) & (g392) & (!g395) & (!g394) & (g401) & (!g396)) + ((!g391) & (g392) & (!g395) & (g394) & (g401) & (g396)) + ((!g391) & (g392) & (g395) & (!g394) & (g401) & (!g396)) + ((!g391) & (g392) & (g395) & (!g394) & (g401) & (g396)) + ((!g391) & (g392) & (g395) & (g394) & (!g401) & (!g396)) + ((!g391) & (g392) & (g395) & (g394) & (!g401) & (g396)) + ((!g391) & (g392) & (g395) & (g394) & (g401) & (g396)) + ((g391) & (!g392) & (!g395) & (!g394) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g394) & (g401) & (g396)) + ((g391) & (!g392) & (!g395) & (g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (g394) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (g394) & (g401) & (g396)) + ((g391) & (!g392) & (g395) & (!g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (g395) & (!g394) & (g401) & (!g396)) + ((g391) & (!g392) & (g395) & (g394) & (g401) & (!g396)) + ((g391) & (g392) & (!g395) & (!g394) & (g401) & (g396)) + ((g391) & (g392) & (g395) & (!g394) & (!g401) & (!g396)) + ((g391) & (g392) & (g395) & (!g394) & (g401) & (g396)));
	assign g435 = (((!g391) & (!g392) & (!g395) & (!g394) & (!g401) & (!g396)) + ((!g391) & (!g392) & (!g395) & (g394) & (!g401) & (!g396)) + ((!g391) & (!g392) & (!g395) & (g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (!g395) & (g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (!g394) & (g401) & (g396)) + ((!g391) & (!g392) & (g395) & (g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (g395) & (g394) & (g401) & (g396)) + ((!g391) & (g392) & (!g395) & (!g394) & (!g401) & (!g396)) + ((!g391) & (g392) & (!g395) & (!g394) & (g401) & (!g396)) + ((!g391) & (g392) & (g395) & (!g394) & (!g401) & (g396)) + ((!g391) & (g392) & (g395) & (!g394) & (g401) & (g396)) + ((!g391) & (g392) & (g395) & (g394) & (!g401) & (g396)) + ((!g391) & (g392) & (g395) & (g394) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g394) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g394) & (g401) & (g396)) + ((g391) & (!g392) & (!g395) & (g394) & (!g401) & (g396)) + ((g391) & (!g392) & (!g395) & (g394) & (g401) & (g396)) + ((g391) & (!g392) & (g395) & (g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (g395) & (g394) & (!g401) & (g396)) + ((g391) & (!g392) & (g395) & (g394) & (g401) & (g396)) + ((g391) & (g392) & (!g395) & (!g394) & (!g401) & (g396)) + ((g391) & (g392) & (!g395) & (!g394) & (g401) & (!g396)) + ((g391) & (g392) & (!g395) & (g394) & (g401) & (!g396)) + ((g391) & (g392) & (g395) & (!g394) & (!g401) & (g396)) + ((g391) & (g392) & (g395) & (!g394) & (g401) & (g396)) + ((g391) & (g392) & (g395) & (g394) & (!g401) & (!g396)) + ((g391) & (g392) & (g395) & (g394) & (g401) & (g396)));
	assign g436 = (((!g391) & (!g392) & (!g395) & (!g394) & (g401) & (g396)) + ((!g391) & (!g392) & (!g395) & (g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (!g394) & (!g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (!g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (g395) & (!g394) & (g401) & (g396)) + ((!g391) & (!g392) & (g395) & (g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (g395) & (g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (g395) & (g394) & (g401) & (g396)) + ((!g391) & (g392) & (!g395) & (!g394) & (g401) & (!g396)) + ((!g391) & (g392) & (!g395) & (!g394) & (g401) & (g396)) + ((!g391) & (g392) & (g395) & (!g394) & (!g401) & (!g396)) + ((!g391) & (g392) & (g395) & (g394) & (!g401) & (g396)) + ((!g391) & (g392) & (g395) & (g394) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g394) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (!g394) & (g401) & (g396)) + ((g391) & (!g392) & (!g395) & (g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (g394) & (!g401) & (g396)) + ((g391) & (!g392) & (g395) & (!g394) & (!g401) & (g396)) + ((g391) & (!g392) & (g395) & (!g394) & (g401) & (g396)) + ((g391) & (!g392) & (g395) & (g394) & (g401) & (!g396)) + ((g391) & (g392) & (!g395) & (!g394) & (!g401) & (!g396)) + ((g391) & (g392) & (!g395) & (!g394) & (!g401) & (g396)) + ((g391) & (g392) & (!g395) & (!g394) & (g401) & (g396)) + ((g391) & (g392) & (!g395) & (g394) & (!g401) & (g396)) + ((g391) & (g392) & (!g395) & (g394) & (g401) & (!g396)) + ((g391) & (g392) & (g395) & (!g394) & (!g401) & (g396)) + ((g391) & (g392) & (g395) & (!g394) & (g401) & (!g396)) + ((g391) & (g392) & (g395) & (g394) & (!g401) & (!g396)) + ((g391) & (g392) & (g395) & (g394) & (g401) & (!g396)) + ((g391) & (g392) & (g395) & (g394) & (g401) & (g396)));
	assign g437 = (((!g391) & (!g392) & (!g395) & (!g394) & (g401) & (!g396)) + ((!g391) & (!g392) & (!g395) & (g394) & (!g401) & (!g396)) + ((!g391) & (!g392) & (!g395) & (g394) & (g401) & (g396)) + ((!g391) & (!g392) & (g395) & (!g394) & (!g401) & (g396)) + ((!g391) & (!g392) & (g395) & (!g394) & (g401) & (g396)) + ((!g391) & (!g392) & (g395) & (g394) & (g401) & (g396)) + ((!g391) & (g392) & (!g395) & (!g394) & (!g401) & (g396)) + ((!g391) & (g392) & (!g395) & (g394) & (!g401) & (g396)) + ((!g391) & (g392) & (!g395) & (g394) & (g401) & (g396)) + ((!g391) & (g392) & (g395) & (!g394) & (!g401) & (!g396)) + ((!g391) & (g392) & (g395) & (!g394) & (g401) & (!g396)) + ((!g391) & (g392) & (g395) & (g394) & (!g401) & (g396)) + ((!g391) & (g392) & (g395) & (g394) & (g401) & (g396)) + ((g391) & (!g392) & (!g395) & (!g394) & (g401) & (!g396)) + ((g391) & (!g392) & (!g395) & (g394) & (g401) & (g396)) + ((g391) & (!g392) & (g395) & (!g394) & (!g401) & (!g396)) + ((g391) & (!g392) & (g395) & (!g394) & (g401) & (g396)) + ((g391) & (!g392) & (g395) & (g394) & (!g401) & (!g396)) + ((g391) & (g392) & (!g395) & (!g394) & (g401) & (g396)) + ((g391) & (g392) & (!g395) & (g394) & (!g401) & (!g396)) + ((g391) & (g392) & (!g395) & (g394) & (!g401) & (g396)) + ((g391) & (g392) & (g395) & (!g394) & (g401) & (g396)));
	assign g438 = (((!g434) & (!g435) & (!g436) & (!g437) & (!g402) & (!g393)) + ((!g434) & (!g435) & (!g436) & (!g437) & (!g402) & (g393)) + ((!g434) & (!g435) & (!g436) & (!g437) & (g402) & (!g393)) + ((!g434) & (!g435) & (!g436) & (g437) & (!g402) & (!g393)) + ((!g434) & (!g435) & (!g436) & (g437) & (!g402) & (g393)) + ((!g434) & (!g435) & (!g436) & (g437) & (g402) & (!g393)) + ((!g434) & (!g435) & (!g436) & (g437) & (g402) & (g393)) + ((!g434) & (!g435) & (g436) & (!g437) & (!g402) & (!g393)) + ((!g434) & (!g435) & (g436) & (!g437) & (g402) & (!g393)) + ((!g434) & (!g435) & (g436) & (g437) & (!g402) & (!g393)) + ((!g434) & (!g435) & (g436) & (g437) & (g402) & (!g393)) + ((!g434) & (!g435) & (g436) & (g437) & (g402) & (g393)) + ((!g434) & (g435) & (!g436) & (!g437) & (!g402) & (!g393)) + ((!g434) & (g435) & (!g436) & (!g437) & (!g402) & (g393)) + ((!g434) & (g435) & (!g436) & (g437) & (!g402) & (!g393)) + ((!g434) & (g435) & (!g436) & (g437) & (!g402) & (g393)) + ((!g434) & (g435) & (!g436) & (g437) & (g402) & (g393)) + ((!g434) & (g435) & (g436) & (!g437) & (!g402) & (!g393)) + ((!g434) & (g435) & (g436) & (g437) & (!g402) & (!g393)) + ((!g434) & (g435) & (g436) & (g437) & (g402) & (g393)) + ((g434) & (!g435) & (!g436) & (!g437) & (!g402) & (g393)) + ((g434) & (!g435) & (!g436) & (!g437) & (g402) & (!g393)) + ((g434) & (!g435) & (!g436) & (g437) & (!g402) & (g393)) + ((g434) & (!g435) & (!g436) & (g437) & (g402) & (!g393)) + ((g434) & (!g435) & (!g436) & (g437) & (g402) & (g393)) + ((g434) & (!g435) & (g436) & (!g437) & (g402) & (!g393)) + ((g434) & (!g435) & (g436) & (g437) & (g402) & (!g393)) + ((g434) & (!g435) & (g436) & (g437) & (g402) & (g393)) + ((g434) & (g435) & (!g436) & (!g437) & (!g402) & (g393)) + ((g434) & (g435) & (!g436) & (g437) & (!g402) & (g393)) + ((g434) & (g435) & (!g436) & (g437) & (g402) & (g393)) + ((g434) & (g435) & (g436) & (g437) & (g402) & (g393)));
	assign g440 = (((!sk[100]) & (g438) & (!g439)) + ((!sk[100]) & (g438) & (g439)) + ((sk[100]) & (!g438) & (g439)) + ((sk[100]) & (g438) & (!g439)));
	assign g441 = (((!g391) & (!g402) & (!g393) & (!g394) & (!g401) & (g396)) + ((!g391) & (!g402) & (!g393) & (!g394) & (g401) & (g396)) + ((!g391) & (!g402) & (!g393) & (g394) & (!g401) & (!g396)) + ((!g391) & (!g402) & (!g393) & (g394) & (!g401) & (g396)) + ((!g391) & (!g402) & (!g393) & (g394) & (g401) & (!g396)) + ((!g391) & (!g402) & (!g393) & (g394) & (g401) & (g396)) + ((!g391) & (!g402) & (g393) & (!g394) & (!g401) & (g396)) + ((!g391) & (!g402) & (g393) & (!g394) & (g401) & (g396)) + ((!g391) & (!g402) & (g393) & (g394) & (g401) & (!g396)) + ((!g391) & (g402) & (g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (g402) & (g393) & (!g394) & (g401) & (g396)) + ((!g391) & (g402) & (g393) & (g394) & (!g401) & (g396)) + ((g391) & (!g402) & (!g393) & (!g394) & (g401) & (!g396)) + ((g391) & (!g402) & (!g393) & (g394) & (!g401) & (!g396)) + ((g391) & (!g402) & (!g393) & (g394) & (!g401) & (g396)) + ((g391) & (!g402) & (!g393) & (g394) & (g401) & (g396)) + ((g391) & (!g402) & (g393) & (!g394) & (!g401) & (g396)) + ((g391) & (!g402) & (g393) & (!g394) & (g401) & (g396)) + ((g391) & (!g402) & (g393) & (g394) & (g401) & (!g396)) + ((g391) & (!g402) & (g393) & (g394) & (g401) & (g396)) + ((g391) & (g402) & (!g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (g402) & (!g393) & (!g394) & (!g401) & (g396)) + ((g391) & (g402) & (!g393) & (!g394) & (g401) & (!g396)) + ((g391) & (g402) & (!g393) & (g394) & (!g401) & (!g396)) + ((g391) & (g402) & (g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (g402) & (g393) & (!g394) & (!g401) & (g396)) + ((g391) & (g402) & (g393) & (!g394) & (g401) & (!g396)) + ((g391) & (g402) & (g393) & (g394) & (!g401) & (g396)));
	assign g442 = (((!g391) & (!g402) & (!g393) & (!g394) & (!g401) & (!g396)) + ((!g391) & (!g402) & (!g393) & (g394) & (g401) & (g396)) + ((!g391) & (!g402) & (g393) & (!g394) & (!g401) & (!g396)) + ((!g391) & (!g402) & (g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (!g402) & (g393) & (!g394) & (g401) & (g396)) + ((!g391) & (!g402) & (g393) & (g394) & (!g401) & (!g396)) + ((!g391) & (!g402) & (g393) & (g394) & (g401) & (g396)) + ((!g391) & (g402) & (!g393) & (!g394) & (!g401) & (!g396)) + ((!g391) & (g402) & (!g393) & (!g394) & (g401) & (g396)) + ((!g391) & (g402) & (!g393) & (g394) & (!g401) & (g396)) + ((!g391) & (g402) & (g393) & (!g394) & (!g401) & (!g396)) + ((!g391) & (g402) & (g393) & (!g394) & (g401) & (g396)) + ((!g391) & (g402) & (g393) & (g394) & (g401) & (!g396)) + ((!g391) & (g402) & (g393) & (g394) & (g401) & (g396)) + ((g391) & (!g402) & (!g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (!g402) & (!g393) & (!g394) & (g401) & (g396)) + ((g391) & (!g402) & (!g393) & (g394) & (!g401) & (!g396)) + ((g391) & (!g402) & (!g393) & (g394) & (g401) & (g396)) + ((g391) & (!g402) & (g393) & (!g394) & (g401) & (g396)) + ((g391) & (!g402) & (g393) & (g394) & (!g401) & (g396)) + ((g391) & (g402) & (!g393) & (!g394) & (g401) & (!g396)) + ((g391) & (g402) & (!g393) & (!g394) & (g401) & (g396)) + ((g391) & (g402) & (!g393) & (g394) & (!g401) & (g396)) + ((g391) & (g402) & (!g393) & (g394) & (g401) & (!g396)) + ((g391) & (g402) & (!g393) & (g394) & (g401) & (g396)) + ((g391) & (g402) & (g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (g402) & (g393) & (!g394) & (g401) & (!g396)) + ((g391) & (g402) & (g393) & (g394) & (!g401) & (!g396)));
	assign g443 = (((!g391) & (!g402) & (!g393) & (!g394) & (!g401) & (g396)) + ((!g391) & (!g402) & (!g393) & (!g394) & (g401) & (g396)) + ((!g391) & (!g402) & (!g393) & (g394) & (g401) & (!g396)) + ((!g391) & (!g402) & (!g393) & (g394) & (g401) & (g396)) + ((!g391) & (!g402) & (g393) & (!g394) & (g401) & (g396)) + ((!g391) & (!g402) & (g393) & (g394) & (!g401) & (!g396)) + ((!g391) & (!g402) & (g393) & (g394) & (!g401) & (g396)) + ((!g391) & (!g402) & (g393) & (g394) & (g401) & (g396)) + ((!g391) & (g402) & (!g393) & (!g394) & (!g401) & (!g396)) + ((!g391) & (g402) & (!g393) & (!g394) & (!g401) & (g396)) + ((!g391) & (g402) & (!g393) & (!g394) & (g401) & (g396)) + ((!g391) & (g402) & (!g393) & (g394) & (!g401) & (g396)) + ((!g391) & (g402) & (!g393) & (g394) & (g401) & (!g396)) + ((!g391) & (g402) & (g393) & (!g394) & (!g401) & (g396)) + ((!g391) & (g402) & (g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (g402) & (g393) & (g394) & (!g401) & (!g396)) + ((!g391) & (g402) & (g393) & (g394) & (g401) & (!g396)) + ((!g391) & (g402) & (g393) & (g394) & (g401) & (g396)) + ((g391) & (!g402) & (!g393) & (!g394) & (!g401) & (g396)) + ((g391) & (!g402) & (!g393) & (g394) & (!g401) & (!g396)) + ((g391) & (!g402) & (!g393) & (g394) & (g401) & (!g396)) + ((g391) & (!g402) & (g393) & (!g394) & (g401) & (g396)) + ((g391) & (!g402) & (g393) & (g394) & (!g401) & (g396)) + ((g391) & (g402) & (!g393) & (!g394) & (!g401) & (g396)) + ((g391) & (g402) & (!g393) & (g394) & (!g401) & (!g396)) + ((g391) & (g402) & (!g393) & (g394) & (g401) & (!g396)) + ((g391) & (g402) & (g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (g402) & (g393) & (!g394) & (g401) & (!g396)) + ((g391) & (g402) & (g393) & (!g394) & (g401) & (g396)) + ((g391) & (g402) & (g393) & (g394) & (g401) & (g396)));
	assign g444 = (((!g391) & (!g402) & (!g393) & (!g394) & (g401) & (g396)) + ((!g391) & (!g402) & (!g393) & (g394) & (!g401) & (!g396)) + ((!g391) & (!g402) & (!g393) & (g394) & (g401) & (g396)) + ((!g391) & (!g402) & (g393) & (!g394) & (!g401) & (!g396)) + ((!g391) & (!g402) & (g393) & (g394) & (g401) & (!g396)) + ((!g391) & (!g402) & (g393) & (g394) & (g401) & (g396)) + ((!g391) & (g402) & (!g393) & (g394) & (!g401) & (!g396)) + ((!g391) & (g402) & (!g393) & (g394) & (g401) & (!g396)) + ((!g391) & (g402) & (g393) & (!g394) & (g401) & (!g396)) + ((!g391) & (g402) & (g393) & (!g394) & (g401) & (g396)) + ((g391) & (!g402) & (!g393) & (!g394) & (!g401) & (g396)) + ((g391) & (!g402) & (!g393) & (!g394) & (g401) & (!g396)) + ((g391) & (!g402) & (!g393) & (g394) & (!g401) & (g396)) + ((g391) & (!g402) & (g393) & (!g394) & (g401) & (!g396)) + ((g391) & (!g402) & (g393) & (!g394) & (g401) & (g396)) + ((g391) & (!g402) & (g393) & (g394) & (g401) & (!g396)) + ((g391) & (!g402) & (g393) & (g394) & (g401) & (g396)) + ((g391) & (g402) & (!g393) & (!g394) & (g401) & (!g396)) + ((g391) & (g402) & (!g393) & (g394) & (!g401) & (g396)) + ((g391) & (g402) & (g393) & (!g394) & (!g401) & (!g396)) + ((g391) & (g402) & (g393) & (!g394) & (g401) & (g396)) + ((g391) & (g402) & (g393) & (g394) & (!g401) & (g396)));
	assign g445 = (((!g441) & (!g442) & (!g443) & (!g444) & (!g395) & (!g392)) + ((!g441) & (!g442) & (!g443) & (!g444) & (!g395) & (g392)) + ((!g441) & (!g442) & (!g443) & (!g444) & (g395) & (!g392)) + ((!g441) & (!g442) & (!g443) & (g444) & (!g395) & (!g392)) + ((!g441) & (!g442) & (!g443) & (g444) & (!g395) & (g392)) + ((!g441) & (!g442) & (!g443) & (g444) & (g395) & (!g392)) + ((!g441) & (!g442) & (!g443) & (g444) & (g395) & (g392)) + ((!g441) & (!g442) & (g443) & (!g444) & (!g395) & (!g392)) + ((!g441) & (!g442) & (g443) & (!g444) & (g395) & (!g392)) + ((!g441) & (!g442) & (g443) & (g444) & (!g395) & (!g392)) + ((!g441) & (!g442) & (g443) & (g444) & (g395) & (!g392)) + ((!g441) & (!g442) & (g443) & (g444) & (g395) & (g392)) + ((!g441) & (g442) & (!g443) & (!g444) & (!g395) & (!g392)) + ((!g441) & (g442) & (!g443) & (!g444) & (!g395) & (g392)) + ((!g441) & (g442) & (!g443) & (g444) & (!g395) & (!g392)) + ((!g441) & (g442) & (!g443) & (g444) & (!g395) & (g392)) + ((!g441) & (g442) & (!g443) & (g444) & (g395) & (g392)) + ((!g441) & (g442) & (g443) & (!g444) & (!g395) & (!g392)) + ((!g441) & (g442) & (g443) & (g444) & (!g395) & (!g392)) + ((!g441) & (g442) & (g443) & (g444) & (g395) & (g392)) + ((g441) & (!g442) & (!g443) & (!g444) & (!g395) & (g392)) + ((g441) & (!g442) & (!g443) & (!g444) & (g395) & (!g392)) + ((g441) & (!g442) & (!g443) & (g444) & (!g395) & (g392)) + ((g441) & (!g442) & (!g443) & (g444) & (g395) & (!g392)) + ((g441) & (!g442) & (!g443) & (g444) & (g395) & (g392)) + ((g441) & (!g442) & (g443) & (!g444) & (g395) & (!g392)) + ((g441) & (!g442) & (g443) & (g444) & (g395) & (!g392)) + ((g441) & (!g442) & (g443) & (g444) & (g395) & (g392)) + ((g441) & (g442) & (!g443) & (!g444) & (!g395) & (g392)) + ((g441) & (g442) & (!g443) & (g444) & (!g395) & (g392)) + ((g441) & (g442) & (!g443) & (g444) & (g395) & (g392)) + ((g441) & (g442) & (g443) & (g444) & (g395) & (g392)));
	assign g447 = (((!sk[106]) & (g445) & (!g446)) + ((!sk[106]) & (g445) & (g446)) + ((sk[106]) & (!g445) & (g446)) + ((sk[106]) & (g445) & (!g446)));
	assign g448 = (((!g395) & (!g392) & (!g393) & (!g394) & (!g401) & (g402)) + ((!g395) & (!g392) & (!g393) & (!g394) & (g401) & (!g402)) + ((!g395) & (!g392) & (!g393) & (g394) & (!g401) & (g402)) + ((!g395) & (!g392) & (!g393) & (g394) & (g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (!g394) & (!g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (!g394) & (g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (g394) & (!g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (g394) & (g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (g394) & (g401) & (g402)) + ((!g395) & (g392) & (!g393) & (!g394) & (g401) & (!g402)) + ((!g395) & (g392) & (!g393) & (g394) & (g401) & (!g402)) + ((!g395) & (g392) & (!g393) & (g394) & (g401) & (g402)) + ((!g395) & (g392) & (g393) & (!g394) & (g401) & (g402)) + ((!g395) & (g392) & (g393) & (g394) & (!g401) & (!g402)) + ((g395) & (!g392) & (!g393) & (!g394) & (!g401) & (g402)) + ((g395) & (!g392) & (!g393) & (g394) & (!g401) & (g402)) + ((g395) & (!g392) & (g393) & (g394) & (g401) & (g402)) + ((g395) & (g392) & (!g393) & (!g394) & (g401) & (g402)) + ((g395) & (g392) & (!g393) & (g394) & (!g401) & (!g402)) + ((g395) & (g392) & (!g393) & (g394) & (g401) & (!g402)) + ((g395) & (g392) & (g393) & (!g394) & (!g401) & (g402)) + ((g395) & (g392) & (g393) & (!g394) & (g401) & (!g402)) + ((g395) & (g392) & (g393) & (!g394) & (g401) & (g402)) + ((g395) & (g392) & (g393) & (g394) & (!g401) & (g402)));
	assign g449 = (((!g395) & (!g392) & (!g393) & (!g394) & (!g401) & (!g402)) + ((!g395) & (!g392) & (!g393) & (!g394) & (!g401) & (g402)) + ((!g395) & (!g392) & (!g393) & (g394) & (!g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (!g394) & (!g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (!g394) & (g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (!g394) & (g401) & (g402)) + ((!g395) & (!g392) & (g393) & (g394) & (!g401) & (g402)) + ((!g395) & (!g392) & (g393) & (g394) & (g401) & (g402)) + ((!g395) & (g392) & (!g393) & (!g394) & (!g401) & (!g402)) + ((!g395) & (g392) & (!g393) & (!g394) & (g401) & (!g402)) + ((!g395) & (g392) & (!g393) & (g394) & (!g401) & (!g402)) + ((!g395) & (g392) & (!g393) & (g394) & (!g401) & (g402)) + ((!g395) & (g392) & (!g393) & (g394) & (g401) & (g402)) + ((!g395) & (g392) & (g393) & (!g394) & (!g401) & (g402)) + ((!g395) & (g392) & (g393) & (g394) & (!g401) & (!g402)) + ((!g395) & (g392) & (g393) & (g394) & (!g401) & (g402)) + ((g395) & (!g392) & (!g393) & (!g394) & (!g401) & (g402)) + ((g395) & (!g392) & (!g393) & (!g394) & (g401) & (g402)) + ((g395) & (!g392) & (!g393) & (g394) & (!g401) & (!g402)) + ((g395) & (!g392) & (!g393) & (g394) & (g401) & (g402)) + ((g395) & (!g392) & (g393) & (!g394) & (!g401) & (!g402)) + ((g395) & (!g392) & (g393) & (!g394) & (g401) & (g402)) + ((g395) & (!g392) & (g393) & (g394) & (g401) & (!g402)) + ((g395) & (g392) & (!g393) & (!g394) & (!g401) & (!g402)) + ((g395) & (g392) & (!g393) & (!g394) & (!g401) & (g402)) + ((g395) & (g392) & (!g393) & (!g394) & (g401) & (g402)) + ((g395) & (g392) & (!g393) & (g394) & (!g401) & (g402)) + ((g395) & (g392) & (!g393) & (g394) & (g401) & (!g402)) + ((g395) & (g392) & (g393) & (!g394) & (g401) & (!g402)) + ((g395) & (g392) & (g393) & (!g394) & (g401) & (g402)));
	assign g450 = (((!g395) & (!g392) & (!g393) & (!g394) & (g401) & (!g402)) + ((!g395) & (!g392) & (!g393) & (g394) & (!g401) & (!g402)) + ((!g395) & (!g392) & (!g393) & (g394) & (g401) & (!g402)) + ((!g395) & (!g392) & (!g393) & (g394) & (g401) & (g402)) + ((!g395) & (!g392) & (g393) & (!g394) & (!g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (!g394) & (!g401) & (g402)) + ((!g395) & (!g392) & (g393) & (!g394) & (g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (g394) & (!g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (g394) & (g401) & (g402)) + ((!g395) & (g392) & (!g393) & (!g394) & (!g401) & (g402)) + ((!g395) & (g392) & (!g393) & (!g394) & (g401) & (!g402)) + ((!g395) & (g392) & (!g393) & (!g394) & (g401) & (g402)) + ((!g395) & (g392) & (g393) & (!g394) & (!g401) & (g402)) + ((!g395) & (g392) & (g393) & (!g394) & (g401) & (!g402)) + ((!g395) & (g392) & (g393) & (!g394) & (g401) & (g402)) + ((!g395) & (g392) & (g393) & (g394) & (!g401) & (!g402)) + ((g395) & (!g392) & (!g393) & (!g394) & (g401) & (!g402)) + ((g395) & (!g392) & (!g393) & (g394) & (!g401) & (!g402)) + ((g395) & (!g392) & (!g393) & (g394) & (g401) & (g402)) + ((g395) & (!g392) & (g393) & (!g394) & (!g401) & (!g402)) + ((g395) & (!g392) & (g393) & (!g394) & (!g401) & (g402)) + ((g395) & (!g392) & (g393) & (g394) & (!g401) & (!g402)) + ((g395) & (!g392) & (g393) & (g394) & (g401) & (!g402)) + ((g395) & (g392) & (!g393) & (!g394) & (g401) & (!g402)) + ((g395) & (g392) & (!g393) & (g394) & (!g401) & (!g402)) + ((g395) & (g392) & (!g393) & (g394) & (g401) & (g402)) + ((g395) & (g392) & (g393) & (!g394) & (!g401) & (!g402)) + ((g395) & (g392) & (g393) & (!g394) & (g401) & (!g402)) + ((g395) & (g392) & (g393) & (!g394) & (g401) & (g402)) + ((g395) & (g392) & (g393) & (g394) & (!g401) & (g402)));
	assign g451 = (((!g395) & (!g392) & (!g393) & (!g394) & (!g401) & (g402)) + ((!g395) & (!g392) & (!g393) & (g394) & (g401) & (!g402)) + ((!g395) & (!g392) & (!g393) & (g394) & (g401) & (g402)) + ((!g395) & (!g392) & (g393) & (!g394) & (!g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (!g394) & (!g401) & (g402)) + ((!g395) & (!g392) & (g393) & (g394) & (g401) & (!g402)) + ((!g395) & (!g392) & (g393) & (g394) & (g401) & (g402)) + ((!g395) & (g392) & (!g393) & (!g394) & (!g401) & (!g402)) + ((!g395) & (g392) & (!g393) & (!g394) & (!g401) & (g402)) + ((!g395) & (g392) & (!g393) & (!g394) & (g401) & (g402)) + ((!g395) & (g392) & (!g393) & (g394) & (!g401) & (g402)) + ((!g395) & (g392) & (g393) & (!g394) & (!g401) & (g402)) + ((!g395) & (g392) & (g393) & (g394) & (!g401) & (!g402)) + ((!g395) & (g392) & (g393) & (g394) & (!g401) & (g402)) + ((!g395) & (g392) & (g393) & (g394) & (g401) & (!g402)) + ((!g395) & (g392) & (g393) & (g394) & (g401) & (g402)) + ((g395) & (!g392) & (!g393) & (g394) & (!g401) & (g402)) + ((g395) & (!g392) & (g393) & (!g394) & (!g401) & (!g402)) + ((g395) & (!g392) & (g393) & (g394) & (!g401) & (!g402)) + ((g395) & (!g392) & (g393) & (g394) & (!g401) & (g402)) + ((g395) & (!g392) & (g393) & (g394) & (g401) & (g402)) + ((g395) & (g392) & (!g393) & (!g394) & (!g401) & (g402)) + ((g395) & (g392) & (!g393) & (!g394) & (g401) & (g402)) + ((g395) & (g392) & (!g393) & (g394) & (!g401) & (!g402)) + ((g395) & (g392) & (!g393) & (g394) & (g401) & (!g402)) + ((g395) & (g392) & (!g393) & (g394) & (g401) & (g402)) + ((g395) & (g392) & (g393) & (!g394) & (g401) & (g402)) + ((g395) & (g392) & (g393) & (g394) & (g401) & (g402)));
	assign g452 = (((!g448) & (!g449) & (!g450) & (!g451) & (!g391) & (g396)) + ((!g448) & (!g449) & (!g450) & (!g451) & (g391) & (!g396)) + ((!g448) & (!g449) & (!g450) & (!g451) & (g391) & (g396)) + ((!g448) & (!g449) & (!g450) & (g451) & (!g391) & (g396)) + ((!g448) & (!g449) & (!g450) & (g451) & (g391) & (!g396)) + ((!g448) & (!g449) & (g450) & (!g451) & (g391) & (!g396)) + ((!g448) & (!g449) & (g450) & (!g451) & (g391) & (g396)) + ((!g448) & (!g449) & (g450) & (g451) & (g391) & (!g396)) + ((!g448) & (g449) & (!g450) & (!g451) & (!g391) & (g396)) + ((!g448) & (g449) & (!g450) & (!g451) & (g391) & (g396)) + ((!g448) & (g449) & (!g450) & (g451) & (!g391) & (g396)) + ((!g448) & (g449) & (g450) & (!g451) & (g391) & (g396)) + ((g448) & (!g449) & (!g450) & (!g451) & (!g391) & (!g396)) + ((g448) & (!g449) & (!g450) & (!g451) & (!g391) & (g396)) + ((g448) & (!g449) & (!g450) & (!g451) & (g391) & (!g396)) + ((g448) & (!g449) & (!g450) & (!g451) & (g391) & (g396)) + ((g448) & (!g449) & (!g450) & (g451) & (!g391) & (!g396)) + ((g448) & (!g449) & (!g450) & (g451) & (!g391) & (g396)) + ((g448) & (!g449) & (!g450) & (g451) & (g391) & (!g396)) + ((g448) & (!g449) & (g450) & (!g451) & (!g391) & (!g396)) + ((g448) & (!g449) & (g450) & (!g451) & (g391) & (!g396)) + ((g448) & (!g449) & (g450) & (!g451) & (g391) & (g396)) + ((g448) & (!g449) & (g450) & (g451) & (!g391) & (!g396)) + ((g448) & (!g449) & (g450) & (g451) & (g391) & (!g396)) + ((g448) & (g449) & (!g450) & (!g451) & (!g391) & (!g396)) + ((g448) & (g449) & (!g450) & (!g451) & (!g391) & (g396)) + ((g448) & (g449) & (!g450) & (!g451) & (g391) & (g396)) + ((g448) & (g449) & (!g450) & (g451) & (!g391) & (!g396)) + ((g448) & (g449) & (!g450) & (g451) & (!g391) & (g396)) + ((g448) & (g449) & (g450) & (!g451) & (!g391) & (!g396)) + ((g448) & (g449) & (g450) & (!g451) & (g391) & (g396)) + ((g448) & (g449) & (g450) & (g451) & (!g391) & (!g396)));
	assign g454 = (((!sk[112]) & (g452) & (!g453)) + ((!sk[112]) & (g452) & (g453)) + ((sk[112]) & (!g452) & (g453)) + ((sk[112]) & (g452) & (!g453)));
	assign g461 = (((!g455) & (!g456) & (!g457) & (!g458) & (g459) & (g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g459) & (!g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g459) & (g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (g459) & (!g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (!g459) & (!g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (!g459) & (g460)) + ((!g455) & (!g456) & (g457) & (g458) & (!g459) & (!g460)) + ((!g455) & (!g456) & (g457) & (g458) & (g459) & (g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (g459) & (!g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (g459) & (g460)) + ((!g455) & (g456) & (!g457) & (g458) & (g459) & (!g460)) + ((!g455) & (g456) & (!g457) & (g458) & (g459) & (g460)) + ((!g455) & (g456) & (g457) & (!g458) & (g459) & (!g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (!g459) & (!g460)) + ((g455) & (!g456) & (g457) & (!g458) & (g459) & (!g460)) + ((g455) & (!g456) & (g457) & (g458) & (!g459) & (g460)) + ((g455) & (!g456) & (g457) & (g458) & (g459) & (g460)) + ((g455) & (g456) & (!g457) & (!g458) & (!g459) & (g460)) + ((g455) & (g456) & (!g457) & (!g458) & (g459) & (!g460)) + ((g455) & (g456) & (g457) & (!g458) & (!g459) & (g460)) + ((g455) & (g456) & (g457) & (!g458) & (g459) & (!g460)) + ((g455) & (g456) & (g457) & (g458) & (!g459) & (!g460)) + ((g455) & (g456) & (g457) & (g458) & (g459) & (!g460)) + ((g455) & (g456) & (g457) & (g458) & (g459) & (g460)));
	assign g462 = (((!g455) & (!g456) & (!g457) & (!g458) & (g459) & (!g460)) + ((!g455) & (!g456) & (!g457) & (!g458) & (g459) & (g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g459) & (!g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g459) & (g460)) + ((!g455) & (!g456) & (g457) & (g458) & (!g459) & (g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (!g459) & (!g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (!g459) & (g460)) + ((!g455) & (g456) & (g457) & (!g458) & (!g459) & (!g460)) + ((!g455) & (g456) & (g457) & (!g458) & (!g459) & (g460)) + ((!g455) & (g456) & (g457) & (!g458) & (g459) & (!g460)) + ((!g455) & (g456) & (g457) & (g458) & (g459) & (g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (!g459) & (g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (g459) & (!g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (g459) & (g460)) + ((g455) & (!g456) & (!g457) & (g458) & (g459) & (!g460)) + ((g455) & (!g456) & (g457) & (!g458) & (!g459) & (!g460)) + ((g455) & (!g456) & (g457) & (!g458) & (g459) & (g460)) + ((g455) & (!g456) & (g457) & (g458) & (!g459) & (g460)) + ((g455) & (!g456) & (g457) & (g458) & (g459) & (g460)) + ((g455) & (g456) & (!g457) & (!g458) & (!g459) & (!g460)) + ((g455) & (g456) & (!g457) & (!g458) & (!g459) & (g460)) + ((g455) & (g456) & (!g457) & (!g458) & (g459) & (!g460)) + ((g455) & (g456) & (!g457) & (!g458) & (g459) & (g460)) + ((g455) & (g456) & (!g457) & (g458) & (!g459) & (!g460)) + ((g455) & (g456) & (!g457) & (g458) & (g459) & (!g460)) + ((g455) & (g456) & (!g457) & (g458) & (g459) & (g460)) + ((g455) & (g456) & (g457) & (!g458) & (g459) & (!g460)) + ((g455) & (g456) & (g457) & (!g458) & (g459) & (g460)) + ((g455) & (g456) & (g457) & (g458) & (!g459) & (g460)) + ((g455) & (g456) & (g457) & (g458) & (g459) & (!g460)));
	assign g463 = (((!g455) & (!g456) & (!g457) & (!g458) & (!g459) & (!g460)) + ((!g455) & (!g456) & (!g457) & (!g458) & (g459) & (g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (g459) & (g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (!g459) & (!g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (!g459) & (g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (g459) & (g460)) + ((!g455) & (!g456) & (g457) & (g458) & (!g459) & (g460)) + ((!g455) & (!g456) & (g457) & (g458) & (g459) & (!g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (!g459) & (!g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (g459) & (!g460)) + ((!g455) & (g456) & (!g457) & (g458) & (g459) & (g460)) + ((!g455) & (g456) & (g457) & (g458) & (!g459) & (!g460)) + ((!g455) & (g456) & (g457) & (g458) & (g459) & (!g460)) + ((g455) & (!g456) & (!g457) & (g458) & (!g459) & (!g460)) + ((g455) & (!g456) & (!g457) & (g458) & (!g459) & (g460)) + ((g455) & (!g456) & (!g457) & (g458) & (g459) & (!g460)) + ((g455) & (!g456) & (g457) & (!g458) & (!g459) & (!g460)) + ((g455) & (!g456) & (g457) & (!g458) & (g459) & (g460)) + ((g455) & (!g456) & (g457) & (g458) & (!g459) & (!g460)) + ((g455) & (!g456) & (g457) & (g458) & (!g459) & (g460)) + ((g455) & (!g456) & (g457) & (g458) & (g459) & (!g460)) + ((g455) & (!g456) & (g457) & (g458) & (g459) & (g460)) + ((g455) & (g456) & (!g457) & (!g458) & (g459) & (g460)) + ((g455) & (g456) & (!g457) & (g458) & (!g459) & (!g460)) + ((g455) & (g456) & (!g457) & (g458) & (g459) & (!g460)) + ((g455) & (g456) & (!g457) & (g458) & (g459) & (g460)) + ((g455) & (g456) & (g457) & (!g458) & (!g459) & (!g460)) + ((g455) & (g456) & (g457) & (g458) & (!g459) & (!g460)) + ((g455) & (g456) & (g457) & (g458) & (!g459) & (g460)) + ((g455) & (g456) & (g457) & (g458) & (g459) & (g460)));
	assign g464 = (((!g455) & (!g456) & (!g457) & (!g458) & (!g459) & (g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (g459) & (!g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (g459) & (g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (!g459) & (g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (g459) & (g460)) + ((!g455) & (!g456) & (g457) & (g458) & (!g459) & (g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (!g459) & (!g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (!g459) & (g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (g459) & (!g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (g459) & (g460)) + ((!g455) & (g456) & (!g457) & (g458) & (g459) & (!g460)) + ((!g455) & (g456) & (!g457) & (g458) & (g459) & (g460)) + ((!g455) & (g456) & (g457) & (g458) & (!g459) & (!g460)) + ((!g455) & (g456) & (g457) & (g458) & (g459) & (!g460)) + ((!g455) & (g456) & (g457) & (g458) & (g459) & (g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (!g459) & (!g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (g459) & (g460)) + ((g455) & (!g456) & (!g457) & (g458) & (g459) & (!g460)) + ((g455) & (!g456) & (!g457) & (g458) & (g459) & (g460)) + ((g455) & (!g456) & (g457) & (!g458) & (!g459) & (g460)) + ((g455) & (!g456) & (g457) & (!g458) & (g459) & (!g460)) + ((g455) & (!g456) & (g457) & (g458) & (g459) & (!g460)) + ((g455) & (g456) & (!g457) & (!g458) & (!g459) & (g460)) + ((g455) & (g456) & (!g457) & (!g458) & (g459) & (g460)) + ((g455) & (g456) & (!g457) & (g458) & (g459) & (!g460)) + ((g455) & (g456) & (!g457) & (g458) & (g459) & (g460)) + ((g455) & (g456) & (g457) & (!g458) & (!g459) & (g460)) + ((g455) & (g456) & (g457) & (g458) & (!g459) & (!g460)));
	assign g467 = (((!g461) & (!g462) & (!g463) & (!g464) & (!g465) & (!g466)) + ((!g461) & (!g462) & (!g463) & (g464) & (!g465) & (!g466)) + ((!g461) & (!g462) & (!g463) & (g464) & (g465) & (g466)) + ((!g461) & (!g462) & (g463) & (!g464) & (!g465) & (!g466)) + ((!g461) & (!g462) & (g463) & (!g464) & (!g465) & (g466)) + ((!g461) & (!g462) & (g463) & (g464) & (!g465) & (!g466)) + ((!g461) & (!g462) & (g463) & (g464) & (!g465) & (g466)) + ((!g461) & (!g462) & (g463) & (g464) & (g465) & (g466)) + ((!g461) & (g462) & (!g463) & (!g464) & (!g465) & (!g466)) + ((!g461) & (g462) & (!g463) & (!g464) & (g465) & (!g466)) + ((!g461) & (g462) & (!g463) & (g464) & (!g465) & (!g466)) + ((!g461) & (g462) & (!g463) & (g464) & (g465) & (!g466)) + ((!g461) & (g462) & (!g463) & (g464) & (g465) & (g466)) + ((!g461) & (g462) & (g463) & (!g464) & (!g465) & (!g466)) + ((!g461) & (g462) & (g463) & (!g464) & (!g465) & (g466)) + ((!g461) & (g462) & (g463) & (!g464) & (g465) & (!g466)) + ((!g461) & (g462) & (g463) & (g464) & (!g465) & (!g466)) + ((!g461) & (g462) & (g463) & (g464) & (!g465) & (g466)) + ((!g461) & (g462) & (g463) & (g464) & (g465) & (!g466)) + ((!g461) & (g462) & (g463) & (g464) & (g465) & (g466)) + ((g461) & (!g462) & (!g463) & (g464) & (g465) & (g466)) + ((g461) & (!g462) & (g463) & (!g464) & (!g465) & (g466)) + ((g461) & (!g462) & (g463) & (g464) & (!g465) & (g466)) + ((g461) & (!g462) & (g463) & (g464) & (g465) & (g466)) + ((g461) & (g462) & (!g463) & (!g464) & (g465) & (!g466)) + ((g461) & (g462) & (!g463) & (g464) & (g465) & (!g466)) + ((g461) & (g462) & (!g463) & (g464) & (g465) & (g466)) + ((g461) & (g462) & (g463) & (!g464) & (!g465) & (g466)) + ((g461) & (g462) & (g463) & (!g464) & (g465) & (!g466)) + ((g461) & (g462) & (g463) & (g464) & (!g465) & (g466)) + ((g461) & (g462) & (g463) & (g464) & (g465) & (!g466)) + ((g461) & (g462) & (g463) & (g464) & (g465) & (g466)));
	assign g469 = (((!g467) & (sk[118]) & (g468)) + ((g467) & (!sk[118]) & (!g468)) + ((g467) & (!sk[118]) & (g468)) + ((g467) & (sk[118]) & (!g468)));
	assign g470 = (((!g455) & (!g456) & (!g457) & (!g458) & (!g465) & (g459)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g465) & (!g459)) + ((!g455) & (!g456) & (!g457) & (g458) & (g465) & (!g459)) + ((!g455) & (!g456) & (g457) & (!g458) & (g465) & (g459)) + ((!g455) & (!g456) & (g457) & (g458) & (!g465) & (g459)) + ((!g455) & (!g456) & (g457) & (g458) & (g465) & (!g459)) + ((!g455) & (g456) & (!g457) & (!g458) & (!g465) & (g459)) + ((!g455) & (g456) & (!g457) & (!g458) & (g465) & (!g459)) + ((!g455) & (g456) & (!g457) & (!g458) & (g465) & (g459)) + ((!g455) & (g456) & (g457) & (!g458) & (g465) & (g459)) + ((!g455) & (g456) & (g457) & (g458) & (g465) & (g459)) + ((g455) & (!g456) & (!g457) & (!g458) & (!g465) & (!g459)) + ((g455) & (!g456) & (!g457) & (!g458) & (g465) & (g459)) + ((g455) & (!g456) & (!g457) & (g458) & (!g465) & (!g459)) + ((g455) & (!g456) & (!g457) & (g458) & (g465) & (!g459)) + ((g455) & (!g456) & (g457) & (!g458) & (g465) & (!g459)) + ((g455) & (!g456) & (g457) & (!g458) & (g465) & (g459)) + ((g455) & (!g456) & (g457) & (g458) & (g465) & (!g459)) + ((g455) & (!g456) & (g457) & (g458) & (g465) & (g459)) + ((g455) & (g456) & (!g457) & (!g458) & (g465) & (!g459)) + ((g455) & (g456) & (!g457) & (!g458) & (g465) & (g459)) + ((g455) & (g456) & (!g457) & (g458) & (g465) & (g459)) + ((g455) & (g456) & (g457) & (!g458) & (!g465) & (!g459)) + ((g455) & (g456) & (g457) & (!g458) & (!g465) & (g459)) + ((g455) & (g456) & (g457) & (!g458) & (g465) & (!g459)) + ((g455) & (g456) & (g457) & (g458) & (!g465) & (g459)) + ((g455) & (g456) & (g457) & (g458) & (g465) & (!g459)));
	assign g471 = (((!g455) & (!g456) & (!g457) & (!g458) & (!g465) & (g459)) + ((!g455) & (!g456) & (!g457) & (!g458) & (g465) & (!g459)) + ((!g455) & (!g456) & (!g457) & (!g458) & (g465) & (g459)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g465) & (!g459)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g465) & (g459)) + ((!g455) & (!g456) & (!g457) & (g458) & (g465) & (g459)) + ((!g455) & (!g456) & (g457) & (!g458) & (g465) & (!g459)) + ((!g455) & (!g456) & (g457) & (g458) & (!g465) & (!g459)) + ((!g455) & (!g456) & (g457) & (g458) & (!g465) & (g459)) + ((!g455) & (!g456) & (g457) & (g458) & (g465) & (g459)) + ((!g455) & (g456) & (!g457) & (!g458) & (g465) & (g459)) + ((!g455) & (g456) & (!g457) & (g458) & (!g465) & (!g459)) + ((!g455) & (g456) & (!g457) & (g458) & (g465) & (!g459)) + ((!g455) & (g456) & (g457) & (!g458) & (g465) & (!g459)) + ((!g455) & (g456) & (g457) & (!g458) & (g465) & (g459)) + ((!g455) & (g456) & (g457) & (g458) & (!g465) & (!g459)) + ((g455) & (!g456) & (!g457) & (!g458) & (!g465) & (!g459)) + ((g455) & (!g456) & (!g457) & (g458) & (!g465) & (!g459)) + ((g455) & (!g456) & (!g457) & (g458) & (!g465) & (g459)) + ((g455) & (!g456) & (g457) & (!g458) & (!g465) & (g459)) + ((g455) & (!g456) & (g457) & (!g458) & (g465) & (g459)) + ((g455) & (!g456) & (g457) & (g458) & (!g465) & (!g459)) + ((g455) & (!g456) & (g457) & (g458) & (!g465) & (g459)) + ((g455) & (g456) & (!g457) & (g458) & (!g465) & (!g459)) + ((g455) & (g456) & (!g457) & (g458) & (g465) & (g459)) + ((g455) & (g456) & (g457) & (!g458) & (!g465) & (!g459)) + ((g455) & (g456) & (g457) & (!g458) & (!g465) & (g459)) + ((g455) & (g456) & (g457) & (!g458) & (g465) & (g459)) + ((g455) & (g456) & (g457) & (g458) & (!g465) & (!g459)) + ((g455) & (g456) & (g457) & (g458) & (!g465) & (g459)) + ((g455) & (g456) & (g457) & (g458) & (g465) & (!g459)));
	assign g472 = (((!g455) & (!g456) & (!g457) & (!g458) & (!g465) & (g459)) + ((!g455) & (!g456) & (!g457) & (g458) & (g465) & (!g459)) + ((!g455) & (!g456) & (g457) & (!g458) & (!g465) & (!g459)) + ((!g455) & (!g456) & (g457) & (!g458) & (g465) & (!g459)) + ((!g455) & (!g456) & (g457) & (g458) & (!g465) & (g459)) + ((!g455) & (!g456) & (g457) & (g458) & (g465) & (!g459)) + ((!g455) & (!g456) & (g457) & (g458) & (g465) & (g459)) + ((!g455) & (g456) & (!g457) & (!g458) & (!g465) & (!g459)) + ((!g455) & (g456) & (!g457) & (!g458) & (g465) & (!g459)) + ((!g455) & (g456) & (!g457) & (g458) & (!g465) & (!g459)) + ((!g455) & (g456) & (!g457) & (g458) & (g465) & (g459)) + ((!g455) & (g456) & (g457) & (!g458) & (g465) & (g459)) + ((!g455) & (g456) & (g457) & (g458) & (!g465) & (g459)) + ((!g455) & (g456) & (g457) & (g458) & (g465) & (!g459)) + ((g455) & (!g456) & (!g457) & (!g458) & (g465) & (g459)) + ((g455) & (!g456) & (!g457) & (g458) & (!g465) & (!g459)) + ((g455) & (!g456) & (!g457) & (g458) & (g465) & (!g459)) + ((g455) & (!g456) & (g457) & (!g458) & (!g465) & (!g459)) + ((g455) & (!g456) & (g457) & (!g458) & (!g465) & (g459)) + ((g455) & (!g456) & (g457) & (!g458) & (g465) & (!g459)) + ((g455) & (!g456) & (g457) & (!g458) & (g465) & (g459)) + ((g455) & (!g456) & (g457) & (g458) & (g465) & (!g459)) + ((g455) & (g456) & (!g457) & (!g458) & (!g465) & (g459)) + ((g455) & (g456) & (!g457) & (!g458) & (g465) & (g459)) + ((g455) & (g456) & (!g457) & (g458) & (!g465) & (g459)) + ((g455) & (g456) & (g457) & (!g458) & (!g465) & (!g459)) + ((g455) & (g456) & (g457) & (!g458) & (!g465) & (g459)) + ((g455) & (g456) & (g457) & (!g458) & (g465) & (g459)) + ((g455) & (g456) & (g457) & (g458) & (!g465) & (!g459)) + ((g455) & (g456) & (g457) & (g458) & (!g465) & (g459)) + ((g455) & (g456) & (g457) & (g458) & (g465) & (!g459)) + ((g455) & (g456) & (g457) & (g458) & (g465) & (g459)));
	assign g473 = (((!g455) & (!g456) & (!g457) & (!g458) & (g465) & (!g459)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g465) & (!g459)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g465) & (g459)) + ((!g455) & (!g456) & (g457) & (!g458) & (g465) & (g459)) + ((!g455) & (!g456) & (g457) & (g458) & (!g465) & (g459)) + ((!g455) & (g456) & (!g457) & (!g458) & (!g465) & (!g459)) + ((!g455) & (g456) & (!g457) & (!g458) & (g465) & (!g459)) + ((!g455) & (g456) & (!g457) & (g458) & (!g465) & (g459)) + ((!g455) & (g456) & (g457) & (!g458) & (!g465) & (g459)) + ((!g455) & (g456) & (g457) & (!g458) & (g465) & (!g459)) + ((!g455) & (g456) & (g457) & (!g458) & (g465) & (g459)) + ((!g455) & (g456) & (g457) & (g458) & (g465) & (!g459)) + ((!g455) & (g456) & (g457) & (g458) & (g465) & (g459)) + ((g455) & (!g456) & (!g457) & (!g458) & (!g465) & (!g459)) + ((g455) & (!g456) & (!g457) & (g458) & (!g465) & (!g459)) + ((g455) & (!g456) & (!g457) & (g458) & (!g465) & (g459)) + ((g455) & (!g456) & (!g457) & (g458) & (g465) & (!g459)) + ((g455) & (!g456) & (g457) & (!g458) & (!g465) & (!g459)) + ((g455) & (!g456) & (g457) & (!g458) & (g465) & (g459)) + ((g455) & (!g456) & (g457) & (g458) & (g465) & (!g459)) + ((g455) & (g456) & (!g457) & (!g458) & (!g465) & (!g459)) + ((g455) & (g456) & (!g457) & (g458) & (!g465) & (!g459)) + ((g455) & (g456) & (!g457) & (g458) & (g465) & (!g459)) + ((g455) & (g456) & (!g457) & (g458) & (g465) & (g459)) + ((g455) & (g456) & (g457) & (g458) & (!g465) & (g459)) + ((g455) & (g456) & (g457) & (g458) & (g465) & (g459)));
	assign g474 = (((!g470) & (!g471) & (!g472) & (!g473) & (!g460) & (!g466)) + ((!g470) & (!g471) & (!g472) & (!g473) & (g460) & (!g466)) + ((!g470) & (!g471) & (!g472) & (g473) & (!g460) & (!g466)) + ((!g470) & (!g471) & (!g472) & (g473) & (g460) & (!g466)) + ((!g470) & (!g471) & (!g472) & (g473) & (g460) & (g466)) + ((!g470) & (!g471) & (g472) & (!g473) & (!g460) & (!g466)) + ((!g470) & (!g471) & (g472) & (!g473) & (!g460) & (g466)) + ((!g470) & (!g471) & (g472) & (!g473) & (g460) & (!g466)) + ((!g470) & (!g471) & (g472) & (g473) & (!g460) & (!g466)) + ((!g470) & (!g471) & (g472) & (g473) & (!g460) & (g466)) + ((!g470) & (!g471) & (g472) & (g473) & (g460) & (!g466)) + ((!g470) & (!g471) & (g472) & (g473) & (g460) & (g466)) + ((!g470) & (g471) & (!g472) & (!g473) & (!g460) & (!g466)) + ((!g470) & (g471) & (!g472) & (g473) & (!g460) & (!g466)) + ((!g470) & (g471) & (!g472) & (g473) & (g460) & (g466)) + ((!g470) & (g471) & (g472) & (!g473) & (!g460) & (!g466)) + ((!g470) & (g471) & (g472) & (!g473) & (!g460) & (g466)) + ((!g470) & (g471) & (g472) & (g473) & (!g460) & (!g466)) + ((!g470) & (g471) & (g472) & (g473) & (!g460) & (g466)) + ((!g470) & (g471) & (g472) & (g473) & (g460) & (g466)) + ((g470) & (!g471) & (!g472) & (!g473) & (g460) & (!g466)) + ((g470) & (!g471) & (!g472) & (g473) & (g460) & (!g466)) + ((g470) & (!g471) & (!g472) & (g473) & (g460) & (g466)) + ((g470) & (!g471) & (g472) & (!g473) & (!g460) & (g466)) + ((g470) & (!g471) & (g472) & (!g473) & (g460) & (!g466)) + ((g470) & (!g471) & (g472) & (g473) & (!g460) & (g466)) + ((g470) & (!g471) & (g472) & (g473) & (g460) & (!g466)) + ((g470) & (!g471) & (g472) & (g473) & (g460) & (g466)) + ((g470) & (g471) & (!g472) & (g473) & (g460) & (g466)) + ((g470) & (g471) & (g472) & (!g473) & (!g460) & (g466)) + ((g470) & (g471) & (g472) & (g473) & (!g460) & (g466)) + ((g470) & (g471) & (g472) & (g473) & (g460) & (g466)));
	assign g476 = (((!g474) & (sk[124]) & (g475)) + ((g474) & (!sk[124]) & (!g475)) + ((g474) & (!sk[124]) & (g475)) + ((g474) & (sk[124]) & (!g475)));
	assign g477 = (((!g459) & (!g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((!g459) & (!g456) & (!g457) & (!g458) & (g465) & (g460)) + ((!g459) & (!g456) & (!g457) & (g458) & (!g465) & (g460)) + ((!g459) & (!g456) & (!g457) & (g458) & (g465) & (!g460)) + ((!g459) & (!g456) & (!g457) & (g458) & (g465) & (g460)) + ((!g459) & (!g456) & (g457) & (!g458) & (!g465) & (g460)) + ((!g459) & (!g456) & (g457) & (g458) & (!g465) & (!g460)) + ((!g459) & (!g456) & (g457) & (g458) & (g465) & (!g460)) + ((!g459) & (g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((!g459) & (g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((!g459) & (g456) & (!g457) & (g458) & (!g465) & (g460)) + ((!g459) & (g456) & (g457) & (!g458) & (!g465) & (!g460)) + ((!g459) & (g456) & (g457) & (!g458) & (!g465) & (g460)) + ((!g459) & (g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g459) & (g456) & (g457) & (!g458) & (g465) & (g460)) + ((g459) & (!g456) & (!g457) & (g458) & (!g465) & (g460)) + ((g459) & (!g456) & (!g457) & (g458) & (g465) & (g460)) + ((g459) & (g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((g459) & (g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((g459) & (g456) & (!g457) & (g458) & (g465) & (!g460)) + ((g459) & (g456) & (g457) & (g458) & (!g465) & (!g460)) + ((g459) & (g456) & (g457) & (g458) & (!g465) & (g460)));
	assign g478 = (((!g459) & (!g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((!g459) & (!g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((!g459) & (!g456) & (!g457) & (g458) & (g465) & (g460)) + ((!g459) & (!g456) & (g457) & (!g458) & (!g465) & (!g460)) + ((!g459) & (!g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g459) & (!g456) & (g457) & (g458) & (!g465) & (g460)) + ((!g459) & (g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((!g459) & (g456) & (!g457) & (!g458) & (g465) & (g460)) + ((!g459) & (g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((!g459) & (g456) & (!g457) & (g458) & (!g465) & (g460)) + ((!g459) & (g456) & (!g457) & (g458) & (g465) & (g460)) + ((!g459) & (g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g459) & (g456) & (g457) & (!g458) & (g465) & (g460)) + ((!g459) & (g456) & (g457) & (g458) & (g465) & (!g460)) + ((g459) & (!g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((g459) & (!g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((g459) & (!g456) & (!g457) & (!g458) & (g465) & (g460)) + ((g459) & (!g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((g459) & (!g456) & (!g457) & (g458) & (!g465) & (g460)) + ((g459) & (!g456) & (!g457) & (g458) & (g465) & (!g460)) + ((g459) & (!g456) & (g457) & (g458) & (!g465) & (!g460)) + ((g459) & (g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((g459) & (g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((g459) & (g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((g459) & (g456) & (!g457) & (g458) & (g465) & (!g460)) + ((g459) & (g456) & (!g457) & (g458) & (g465) & (g460)) + ((g459) & (g456) & (g457) & (!g458) & (!g465) & (!g460)) + ((g459) & (g456) & (g457) & (!g458) & (g465) & (!g460)) + ((g459) & (g456) & (g457) & (g458) & (!g465) & (g460)) + ((g459) & (g456) & (g457) & (g458) & (g465) & (g460)));
	assign g479 = (((!g459) & (!g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((!g459) & (!g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((!g459) & (!g456) & (!g457) & (g458) & (!g465) & (g460)) + ((!g459) & (!g456) & (g457) & (!g458) & (!g465) & (g460)) + ((!g459) & (!g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g459) & (!g456) & (g457) & (g458) & (!g465) & (g460)) + ((!g459) & (g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((!g459) & (g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((!g459) & (g456) & (!g457) & (g458) & (g465) & (!g460)) + ((!g459) & (g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g459) & (g456) & (g457) & (g458) & (!g465) & (!g460)) + ((!g459) & (g456) & (g457) & (g458) & (g465) & (!g460)) + ((g459) & (!g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((g459) & (!g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((g459) & (!g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((g459) & (!g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((g459) & (!g456) & (!g457) & (g458) & (!g465) & (g460)) + ((g459) & (!g456) & (!g457) & (g458) & (g465) & (!g460)) + ((g459) & (!g456) & (!g457) & (g458) & (g465) & (g460)) + ((g459) & (!g456) & (g457) & (!g458) & (!g465) & (g460)) + ((g459) & (!g456) & (g457) & (!g458) & (g465) & (!g460)) + ((g459) & (!g456) & (g457) & (g458) & (!g465) & (!g460)) + ((g459) & (!g456) & (g457) & (g458) & (g465) & (g460)) + ((g459) & (g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((g459) & (g456) & (!g457) & (!g458) & (g465) & (g460)) + ((g459) & (g456) & (g457) & (!g458) & (g465) & (g460)) + ((g459) & (g456) & (g457) & (g458) & (!g465) & (!g460)) + ((g459) & (g456) & (g457) & (g458) & (!g465) & (g460)) + ((g459) & (g456) & (g457) & (g458) & (g465) & (g460)));
	assign g480 = (((!g459) & (!g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((!g459) & (!g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((!g459) & (!g456) & (!g457) & (!g458) & (g465) & (g460)) + ((!g459) & (!g456) & (!g457) & (g458) & (!g465) & (g460)) + ((!g459) & (!g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g459) & (!g456) & (g457) & (g458) & (g465) & (g460)) + ((!g459) & (g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((!g459) & (g456) & (!g457) & (g458) & (!g465) & (g460)) + ((!g459) & (g456) & (!g457) & (g458) & (g465) & (g460)) + ((!g459) & (g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g459) & (g456) & (g457) & (!g458) & (g465) & (g460)) + ((!g459) & (g456) & (g457) & (g458) & (!g465) & (!g460)) + ((!g459) & (g456) & (g457) & (g458) & (!g465) & (g460)) + ((!g459) & (g456) & (g457) & (g458) & (g465) & (!g460)) + ((!g459) & (g456) & (g457) & (g458) & (g465) & (g460)) + ((g459) & (!g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((g459) & (!g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((g459) & (!g456) & (!g457) & (!g458) & (g465) & (g460)) + ((g459) & (!g456) & (!g457) & (g458) & (g465) & (g460)) + ((g459) & (!g456) & (g457) & (!g458) & (!g465) & (g460)) + ((g459) & (!g456) & (g457) & (!g458) & (g465) & (!g460)) + ((g459) & (!g456) & (g457) & (g458) & (g465) & (!g460)) + ((g459) & (g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((g459) & (g456) & (!g457) & (g458) & (!g465) & (g460)) + ((g459) & (g456) & (!g457) & (g458) & (g465) & (!g460)) + ((g459) & (g456) & (g457) & (!g458) & (g465) & (g460)) + ((g459) & (g456) & (g457) & (g458) & (!g465) & (!g460)));
	assign g481 = (((!g477) & (!g478) & (!g479) & (!g480) & (!g455) & (g466)) + ((!g477) & (!g478) & (!g479) & (!g480) & (g455) & (!g466)) + ((!g477) & (!g478) & (!g479) & (!g480) & (g455) & (g466)) + ((!g477) & (!g478) & (!g479) & (g480) & (!g455) & (g466)) + ((!g477) & (!g478) & (!g479) & (g480) & (g455) & (!g466)) + ((!g477) & (!g478) & (g479) & (!g480) & (g455) & (!g466)) + ((!g477) & (!g478) & (g479) & (!g480) & (g455) & (g466)) + ((!g477) & (!g478) & (g479) & (g480) & (g455) & (!g466)) + ((!g477) & (g478) & (!g479) & (!g480) & (!g455) & (g466)) + ((!g477) & (g478) & (!g479) & (!g480) & (g455) & (g466)) + ((!g477) & (g478) & (!g479) & (g480) & (!g455) & (g466)) + ((!g477) & (g478) & (g479) & (!g480) & (g455) & (g466)) + ((g477) & (!g478) & (!g479) & (!g480) & (!g455) & (!g466)) + ((g477) & (!g478) & (!g479) & (!g480) & (!g455) & (g466)) + ((g477) & (!g478) & (!g479) & (!g480) & (g455) & (!g466)) + ((g477) & (!g478) & (!g479) & (!g480) & (g455) & (g466)) + ((g477) & (!g478) & (!g479) & (g480) & (!g455) & (!g466)) + ((g477) & (!g478) & (!g479) & (g480) & (!g455) & (g466)) + ((g477) & (!g478) & (!g479) & (g480) & (g455) & (!g466)) + ((g477) & (!g478) & (g479) & (!g480) & (!g455) & (!g466)) + ((g477) & (!g478) & (g479) & (!g480) & (g455) & (!g466)) + ((g477) & (!g478) & (g479) & (!g480) & (g455) & (g466)) + ((g477) & (!g478) & (g479) & (g480) & (!g455) & (!g466)) + ((g477) & (!g478) & (g479) & (g480) & (g455) & (!g466)) + ((g477) & (g478) & (!g479) & (!g480) & (!g455) & (!g466)) + ((g477) & (g478) & (!g479) & (!g480) & (!g455) & (g466)) + ((g477) & (g478) & (!g479) & (!g480) & (g455) & (g466)) + ((g477) & (g478) & (!g479) & (g480) & (!g455) & (!g466)) + ((g477) & (g478) & (!g479) & (g480) & (!g455) & (g466)) + ((g477) & (g478) & (g479) & (!g480) & (!g455) & (!g466)) + ((g477) & (g478) & (g479) & (!g480) & (g455) & (g466)) + ((g477) & (g478) & (g479) & (g480) & (!g455) & (!g466)));
	assign g483 = (((!sk[2]) & (g481) & (!g482)) + ((!sk[2]) & (g481) & (g482)) + ((sk[2]) & (!g481) & (g482)) + ((sk[2]) & (g481) & (!g482)));
	assign g484 = (((!g455) & (!g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (g465) & (g460)) + ((!g455) & (!g456) & (g457) & (g458) & (!g465) & (!g460)) + ((!g455) & (!g456) & (g457) & (g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (g457) & (g458) & (g465) & (g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (g456) & (g457) & (!g458) & (!g465) & (!g460)) + ((!g455) & (g456) & (g457) & (g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((g455) & (!g456) & (g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (g457) & (!g458) & (!g465) & (g460)) + ((g455) & (!g456) & (g457) & (!g458) & (g465) & (!g460)) + ((g455) & (!g456) & (g457) & (g458) & (!g465) & (g460)) + ((g455) & (g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((g455) & (g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((g455) & (g456) & (!g457) & (g458) & (g465) & (!g460)) + ((g455) & (g456) & (g457) & (!g458) & (!g465) & (g460)) + ((g455) & (g456) & (g457) & (!g458) & (g465) & (g460)));
	assign g485 = (((!g455) & (!g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (!g457) & (!g458) & (g465) & (g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (g457) & (g458) & (!g465) & (!g460)) + ((!g455) & (!g456) & (g457) & (g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (g457) & (g458) & (g465) & (g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (g465) & (g460)) + ((!g455) & (g456) & (!g457) & (g458) & (g465) & (g460)) + ((!g455) & (g456) & (g457) & (!g458) & (!g465) & (!g460)) + ((!g455) & (g456) & (g457) & (!g458) & (!g465) & (g460)) + ((!g455) & (g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (g456) & (g457) & (g458) & (!g465) & (g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((g455) & (!g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (!g457) & (g458) & (!g465) & (g460)) + ((g455) & (!g456) & (!g457) & (g458) & (g465) & (g460)) + ((g455) & (!g456) & (g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (g457) & (!g458) & (!g465) & (g460)) + ((g455) & (!g456) & (g457) & (!g458) & (g465) & (g460)) + ((g455) & (!g456) & (g457) & (g458) & (!g465) & (g460)) + ((g455) & (g456) & (!g457) & (g458) & (!g465) & (g460)) + ((g455) & (g456) & (!g457) & (g458) & (g465) & (!g460)) + ((g455) & (g456) & (g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (g456) & (g457) & (g458) & (!g465) & (!g460)));
	assign g486 = (((!g455) & (!g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (!g457) & (!g458) & (g465) & (g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (g457) & (!g458) & (g465) & (g460)) + ((!g455) & (!g456) & (g457) & (g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (g457) & (g458) & (g465) & (g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (g465) & (g460)) + ((!g455) & (g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((!g455) & (g456) & (!g457) & (g458) & (!g465) & (g460)) + ((!g455) & (g456) & (g457) & (!g458) & (!g465) & (g460)) + ((!g455) & (g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (g456) & (g457) & (g458) & (g465) & (g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (g465) & (g460)) + ((g455) & (!g456) & (!g457) & (g458) & (g465) & (g460)) + ((g455) & (!g456) & (g457) & (g458) & (!g465) & (!g460)) + ((g455) & (g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((g455) & (g456) & (!g457) & (g458) & (g465) & (g460)) + ((g455) & (g456) & (g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (g456) & (g457) & (!g458) & (!g465) & (g460)) + ((g455) & (g456) & (g457) & (!g458) & (g465) & (g460)) + ((g455) & (g456) & (g457) & (g458) & (!g465) & (!g460)) + ((g455) & (g456) & (g457) & (g458) & (g465) & (g460)));
	assign g487 = (((!g455) & (!g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (!g457) & (g458) & (g465) & (g460)) + ((!g455) & (!g456) & (g457) & (g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (g457) & (g458) & (g465) & (g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (!g465) & (!g460)) + ((!g455) & (g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (g456) & (!g457) & (g458) & (!g465) & (!g460)) + ((!g455) & (g456) & (!g457) & (g458) & (!g465) & (g460)) + ((!g455) & (g456) & (!g457) & (g458) & (g465) & (!g460)) + ((!g455) & (g456) & (g457) & (!g458) & (!g465) & (!g460)) + ((!g455) & (g456) & (g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (g456) & (g457) & (!g458) & (g465) & (g460)) + ((g455) & (!g456) & (!g457) & (!g458) & (g465) & (g460)) + ((g455) & (!g456) & (!g457) & (g458) & (g465) & (!g460)) + ((g455) & (!g456) & (g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (g457) & (!g458) & (g465) & (!g460)) + ((g455) & (!g456) & (g457) & (!g458) & (g465) & (g460)) + ((g455) & (!g456) & (g457) & (g458) & (!g465) & (g460)) + ((g455) & (!g456) & (g457) & (g458) & (g465) & (!g460)) + ((g455) & (!g456) & (g457) & (g458) & (g465) & (g460)) + ((g455) & (g456) & (!g457) & (!g458) & (!g465) & (g460)) + ((g455) & (g456) & (!g457) & (!g458) & (g465) & (!g460)) + ((g455) & (g456) & (g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (g456) & (g457) & (!g458) & (!g465) & (g460)) + ((g455) & (g456) & (g457) & (g458) & (g465) & (g460)));
	assign g488 = (((!g484) & (!g485) & (!g486) & (!g487) & (!g466) & (g459)) + ((!g484) & (!g485) & (!g486) & (!g487) & (g466) & (!g459)) + ((!g484) & (!g485) & (!g486) & (!g487) & (g466) & (g459)) + ((!g484) & (!g485) & (!g486) & (g487) & (!g466) & (g459)) + ((!g484) & (!g485) & (!g486) & (g487) & (g466) & (!g459)) + ((!g484) & (!g485) & (g486) & (!g487) & (g466) & (!g459)) + ((!g484) & (!g485) & (g486) & (!g487) & (g466) & (g459)) + ((!g484) & (!g485) & (g486) & (g487) & (g466) & (!g459)) + ((!g484) & (g485) & (!g486) & (!g487) & (!g466) & (g459)) + ((!g484) & (g485) & (!g486) & (!g487) & (g466) & (g459)) + ((!g484) & (g485) & (!g486) & (g487) & (!g466) & (g459)) + ((!g484) & (g485) & (g486) & (!g487) & (g466) & (g459)) + ((g484) & (!g485) & (!g486) & (!g487) & (!g466) & (!g459)) + ((g484) & (!g485) & (!g486) & (!g487) & (!g466) & (g459)) + ((g484) & (!g485) & (!g486) & (!g487) & (g466) & (!g459)) + ((g484) & (!g485) & (!g486) & (!g487) & (g466) & (g459)) + ((g484) & (!g485) & (!g486) & (g487) & (!g466) & (!g459)) + ((g484) & (!g485) & (!g486) & (g487) & (!g466) & (g459)) + ((g484) & (!g485) & (!g486) & (g487) & (g466) & (!g459)) + ((g484) & (!g485) & (g486) & (!g487) & (!g466) & (!g459)) + ((g484) & (!g485) & (g486) & (!g487) & (g466) & (!g459)) + ((g484) & (!g485) & (g486) & (!g487) & (g466) & (g459)) + ((g484) & (!g485) & (g486) & (g487) & (!g466) & (!g459)) + ((g484) & (!g485) & (g486) & (g487) & (g466) & (!g459)) + ((g484) & (g485) & (!g486) & (!g487) & (!g466) & (!g459)) + ((g484) & (g485) & (!g486) & (!g487) & (!g466) & (g459)) + ((g484) & (g485) & (!g486) & (!g487) & (g466) & (g459)) + ((g484) & (g485) & (!g486) & (g487) & (!g466) & (!g459)) + ((g484) & (g485) & (!g486) & (g487) & (!g466) & (g459)) + ((g484) & (g485) & (g486) & (!g487) & (!g466) & (!g459)) + ((g484) & (g485) & (g486) & (!g487) & (g466) & (g459)) + ((g484) & (g485) & (g486) & (g487) & (!g466) & (!g459)));
	assign g490 = (((!g488) & (sk[8]) & (g489)) + ((g488) & (!sk[8]) & (!g489)) + ((g488) & (!sk[8]) & (g489)) + ((g488) & (sk[8]) & (!g489)));
	assign g491 = (((!g455) & (!g456) & (!g459) & (!g466) & (!g465) & (g460)) + ((!g455) & (!g456) & (g459) & (!g466) & (!g465) & (g460)) + ((!g455) & (!g456) & (g459) & (!g466) & (g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (!g466) & (g465) & (g460)) + ((!g455) & (!g456) & (g459) & (g466) & (!g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (g466) & (g465) & (!g460)) + ((!g455) & (g456) & (!g459) & (!g466) & (!g465) & (!g460)) + ((!g455) & (g456) & (!g459) & (!g466) & (!g465) & (g460)) + ((!g455) & (g456) & (!g459) & (g466) & (!g465) & (!g460)) + ((!g455) & (g456) & (!g459) & (g466) & (!g465) & (g460)) + ((!g455) & (g456) & (!g459) & (g466) & (g465) & (g460)) + ((!g455) & (g456) & (g459) & (g466) & (!g465) & (g460)) + ((!g455) & (g456) & (g459) & (g466) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g466) & (!g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g466) & (!g465) & (g460)) + ((g455) & (!g456) & (!g459) & (g466) & (!g465) & (g460)) + ((g455) & (!g456) & (g459) & (!g466) & (g465) & (!g460)) + ((g455) & (!g456) & (g459) & (g466) & (!g465) & (!g460)) + ((g455) & (!g456) & (g459) & (g466) & (!g465) & (g460)) + ((g455) & (!g456) & (g459) & (g466) & (g465) & (!g460)) + ((g455) & (g456) & (!g459) & (!g466) & (!g465) & (!g460)) + ((g455) & (g456) & (!g459) & (!g466) & (g465) & (!g460)) + ((g455) & (g456) & (!g459) & (g466) & (g465) & (!g460)) + ((g455) & (g456) & (g459) & (!g466) & (!g465) & (!g460)) + ((g455) & (g456) & (g459) & (!g466) & (!g465) & (g460)) + ((g455) & (g456) & (g459) & (g466) & (!g465) & (g460)));
	assign g492 = (((!g455) & (!g456) & (!g459) & (!g466) & (!g465) & (!g460)) + ((!g455) & (!g456) & (!g459) & (!g466) & (!g465) & (g460)) + ((!g455) & (!g456) & (!g459) & (!g466) & (g465) & (!g460)) + ((!g455) & (!g456) & (!g459) & (!g466) & (g465) & (g460)) + ((!g455) & (!g456) & (!g459) & (g466) & (!g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (!g466) & (!g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (!g466) & (g465) & (g460)) + ((!g455) & (!g456) & (g459) & (g466) & (!g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (g466) & (g465) & (g460)) + ((!g455) & (g456) & (!g459) & (!g466) & (!g465) & (g460)) + ((!g455) & (g456) & (!g459) & (g466) & (g465) & (!g460)) + ((!g455) & (g456) & (g459) & (!g466) & (!g465) & (!g460)) + ((!g455) & (g456) & (g459) & (!g466) & (!g465) & (g460)) + ((!g455) & (g456) & (g459) & (!g466) & (g465) & (!g460)) + ((!g455) & (g456) & (g459) & (!g466) & (g465) & (g460)) + ((!g455) & (g456) & (g459) & (g466) & (!g465) & (!g460)) + ((!g455) & (g456) & (g459) & (g466) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g466) & (!g465) & (g460)) + ((g455) & (!g456) & (!g459) & (!g466) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g466) & (g465) & (g460)) + ((g455) & (!g456) & (!g459) & (g466) & (!g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (g466) & (g465) & (g460)) + ((g455) & (!g456) & (g459) & (!g466) & (g465) & (!g460)) + ((g455) & (!g456) & (g459) & (!g466) & (g465) & (g460)) + ((g455) & (!g456) & (g459) & (g466) & (!g465) & (g460)) + ((g455) & (g456) & (!g459) & (!g466) & (g465) & (!g460)) + ((g455) & (g456) & (!g459) & (!g466) & (g465) & (g460)) + ((g455) & (g456) & (!g459) & (g466) & (!g465) & (!g460)) + ((g455) & (g456) & (!g459) & (g466) & (!g465) & (g460)) + ((g455) & (g456) & (g459) & (!g466) & (g465) & (!g460)) + ((g455) & (g456) & (g459) & (!g466) & (g465) & (g460)) + ((g455) & (g456) & (g459) & (g466) & (!g465) & (g460)));
	assign g493 = (((!g455) & (!g456) & (!g459) & (!g466) & (!g465) & (!g460)) + ((!g455) & (!g456) & (!g459) & (!g466) & (!g465) & (g460)) + ((!g455) & (!g456) & (g459) & (!g466) & (!g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (!g466) & (g465) & (g460)) + ((!g455) & (!g456) & (g459) & (g466) & (!g465) & (g460)) + ((!g455) & (g456) & (!g459) & (g466) & (!g465) & (!g460)) + ((!g455) & (g456) & (!g459) & (g466) & (g465) & (!g460)) + ((!g455) & (g456) & (!g459) & (g466) & (g465) & (g460)) + ((!g455) & (g456) & (g459) & (!g466) & (!g465) & (!g460)) + ((!g455) & (g456) & (g459) & (!g466) & (g465) & (!g460)) + ((!g455) & (g456) & (g459) & (!g466) & (g465) & (g460)) + ((!g455) & (g456) & (g459) & (g466) & (!g465) & (!g460)) + ((!g455) & (g456) & (g459) & (g466) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g466) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g466) & (g465) & (g460)) + ((g455) & (!g456) & (!g459) & (g466) & (!g465) & (g460)) + ((g455) & (!g456) & (!g459) & (g466) & (g465) & (g460)) + ((g455) & (!g456) & (g459) & (!g466) & (!g465) & (!g460)) + ((g455) & (!g456) & (g459) & (!g466) & (!g465) & (g460)) + ((g455) & (!g456) & (g459) & (!g466) & (g465) & (g460)) + ((g455) & (!g456) & (g459) & (g466) & (!g465) & (!g460)) + ((g455) & (!g456) & (g459) & (g466) & (!g465) & (g460)) + ((g455) & (!g456) & (g459) & (g466) & (g465) & (!g460)) + ((g455) & (!g456) & (g459) & (g466) & (g465) & (g460)) + ((g455) & (g456) & (!g459) & (!g466) & (!g465) & (g460)) + ((g455) & (g456) & (!g459) & (g466) & (!g465) & (!g460)) + ((g455) & (g456) & (!g459) & (g466) & (g465) & (!g460)) + ((g455) & (g456) & (g459) & (!g466) & (!g465) & (!g460)) + ((g455) & (g456) & (g459) & (!g466) & (!g465) & (g460)) + ((g455) & (g456) & (g459) & (!g466) & (g465) & (!g460)) + ((g455) & (g456) & (g459) & (g466) & (!g465) & (!g460)) + ((g455) & (g456) & (g459) & (g466) & (g465) & (!g460)));
	assign g494 = (((!g455) & (!g456) & (!g459) & (!g466) & (g465) & (g460)) + ((!g455) & (!g456) & (!g459) & (g466) & (!g465) & (!g460)) + ((!g455) & (!g456) & (!g459) & (g466) & (g465) & (g460)) + ((!g455) & (!g456) & (g459) & (!g466) & (!g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (!g466) & (g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (g466) & (!g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (g466) & (!g465) & (g460)) + ((!g455) & (!g456) & (g459) & (g466) & (g465) & (!g460)) + ((!g455) & (g456) & (!g459) & (!g466) & (!g465) & (!g460)) + ((!g455) & (g456) & (!g459) & (g466) & (!g465) & (g460)) + ((!g455) & (g456) & (!g459) & (g466) & (g465) & (!g460)) + ((!g455) & (g456) & (!g459) & (g466) & (g465) & (g460)) + ((!g455) & (g456) & (g459) & (!g466) & (!g465) & (!g460)) + ((!g455) & (g456) & (g459) & (g466) & (!g465) & (!g460)) + ((!g455) & (g456) & (g459) & (g466) & (!g465) & (g460)) + ((g455) & (!g456) & (!g459) & (!g466) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g466) & (g465) & (g460)) + ((g455) & (!g456) & (g459) & (!g466) & (!g465) & (!g460)) + ((g455) & (!g456) & (g459) & (!g466) & (g465) & (!g460)) + ((g455) & (!g456) & (g459) & (g466) & (g465) & (!g460)) + ((g455) & (g456) & (!g459) & (!g466) & (g465) & (!g460)) + ((g455) & (g456) & (!g459) & (g466) & (g465) & (g460)) + ((g455) & (g456) & (g459) & (!g466) & (!g465) & (!g460)) + ((g455) & (g456) & (g459) & (!g466) & (!g465) & (g460)) + ((g455) & (g456) & (g459) & (!g466) & (g465) & (!g460)) + ((g455) & (g456) & (g459) & (g466) & (!g465) & (!g460)));
	assign g495 = (((!g491) & (!g492) & (!g493) & (!g494) & (g457) & (g458)) + ((!g491) & (!g492) & (g493) & (!g494) & (!g457) & (g458)) + ((!g491) & (!g492) & (g493) & (!g494) & (g457) & (g458)) + ((!g491) & (!g492) & (g493) & (g494) & (!g457) & (g458)) + ((!g491) & (g492) & (!g493) & (!g494) & (g457) & (!g458)) + ((!g491) & (g492) & (!g493) & (!g494) & (g457) & (g458)) + ((!g491) & (g492) & (!g493) & (g494) & (g457) & (!g458)) + ((!g491) & (g492) & (g493) & (!g494) & (!g457) & (g458)) + ((!g491) & (g492) & (g493) & (!g494) & (g457) & (!g458)) + ((!g491) & (g492) & (g493) & (!g494) & (g457) & (g458)) + ((!g491) & (g492) & (g493) & (g494) & (!g457) & (g458)) + ((!g491) & (g492) & (g493) & (g494) & (g457) & (!g458)) + ((g491) & (!g492) & (!g493) & (!g494) & (!g457) & (!g458)) + ((g491) & (!g492) & (!g493) & (!g494) & (g457) & (g458)) + ((g491) & (!g492) & (!g493) & (g494) & (!g457) & (!g458)) + ((g491) & (!g492) & (g493) & (!g494) & (!g457) & (!g458)) + ((g491) & (!g492) & (g493) & (!g494) & (!g457) & (g458)) + ((g491) & (!g492) & (g493) & (!g494) & (g457) & (g458)) + ((g491) & (!g492) & (g493) & (g494) & (!g457) & (!g458)) + ((g491) & (!g492) & (g493) & (g494) & (!g457) & (g458)) + ((g491) & (g492) & (!g493) & (!g494) & (!g457) & (!g458)) + ((g491) & (g492) & (!g493) & (!g494) & (g457) & (!g458)) + ((g491) & (g492) & (!g493) & (!g494) & (g457) & (g458)) + ((g491) & (g492) & (!g493) & (g494) & (!g457) & (!g458)) + ((g491) & (g492) & (!g493) & (g494) & (g457) & (!g458)) + ((g491) & (g492) & (g493) & (!g494) & (!g457) & (!g458)) + ((g491) & (g492) & (g493) & (!g494) & (!g457) & (g458)) + ((g491) & (g492) & (g493) & (!g494) & (g457) & (!g458)) + ((g491) & (g492) & (g493) & (!g494) & (g457) & (g458)) + ((g491) & (g492) & (g493) & (g494) & (!g457) & (!g458)) + ((g491) & (g492) & (g493) & (g494) & (!g457) & (g458)) + ((g491) & (g492) & (g493) & (g494) & (g457) & (!g458)));
	assign g497 = (((!g495) & (sk[14]) & (g496)) + ((g495) & (!sk[14]) & (!g496)) + ((g495) & (!sk[14]) & (g496)) + ((g495) & (sk[14]) & (!g496)));
	assign g498 = (((!g455) & (!g456) & (!g459) & (!g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (!g459) & (!g458) & (g465) & (g460)) + ((!g455) & (!g456) & (!g459) & (g458) & (g465) & (g460)) + ((!g455) & (!g456) & (g459) & (!g458) & (!g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (!g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (g459) & (!g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (!g458) & (g465) & (g460)) + ((!g455) & (!g456) & (g459) & (g458) & (!g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (g458) & (!g465) & (g460)) + ((!g455) & (g456) & (!g459) & (!g458) & (!g465) & (g460)) + ((!g455) & (g456) & (!g459) & (!g458) & (g465) & (!g460)) + ((!g455) & (g456) & (!g459) & (g458) & (g465) & (g460)) + ((!g455) & (g456) & (g459) & (!g458) & (g465) & (!g460)) + ((!g455) & (g456) & (g459) & (!g458) & (g465) & (g460)) + ((!g455) & (g456) & (g459) & (g458) & (!g465) & (!g460)) + ((!g455) & (g456) & (g459) & (g458) & (!g465) & (g460)) + ((!g455) & (g456) & (g459) & (g458) & (g465) & (g460)) + ((g455) & (!g456) & (!g459) & (!g458) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g458) & (g465) & (g460)) + ((g455) & (!g456) & (!g459) & (g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (g458) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (g458) & (g465) & (g460)) + ((g455) & (!g456) & (g459) & (!g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (g459) & (!g458) & (g465) & (!g460)) + ((g455) & (!g456) & (g459) & (g458) & (g465) & (!g460)) + ((g455) & (g456) & (!g459) & (!g458) & (g465) & (g460)) + ((g455) & (g456) & (g459) & (!g458) & (!g465) & (!g460)) + ((g455) & (g456) & (g459) & (!g458) & (g465) & (g460)));
	assign g499 = (((!g455) & (!g456) & (!g459) & (!g458) & (!g465) & (!g460)) + ((!g455) & (!g456) & (!g459) & (g458) & (!g465) & (!g460)) + ((!g455) & (!g456) & (!g459) & (g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (!g459) & (g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (!g458) & (g465) & (g460)) + ((!g455) & (!g456) & (g459) & (g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (g459) & (g458) & (g465) & (g460)) + ((!g455) & (g456) & (!g459) & (!g458) & (!g465) & (!g460)) + ((!g455) & (g456) & (!g459) & (!g458) & (g465) & (!g460)) + ((!g455) & (g456) & (g459) & (!g458) & (!g465) & (g460)) + ((!g455) & (g456) & (g459) & (!g458) & (g465) & (g460)) + ((!g455) & (g456) & (g459) & (g458) & (!g465) & (g460)) + ((!g455) & (g456) & (g459) & (g458) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g458) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g458) & (g465) & (g460)) + ((g455) & (!g456) & (!g459) & (g458) & (!g465) & (g460)) + ((g455) & (!g456) & (!g459) & (g458) & (g465) & (g460)) + ((g455) & (!g456) & (g459) & (g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (g459) & (g458) & (!g465) & (g460)) + ((g455) & (!g456) & (g459) & (g458) & (g465) & (g460)) + ((g455) & (g456) & (!g459) & (!g458) & (!g465) & (g460)) + ((g455) & (g456) & (!g459) & (!g458) & (g465) & (!g460)) + ((g455) & (g456) & (!g459) & (g458) & (g465) & (!g460)) + ((g455) & (g456) & (g459) & (!g458) & (!g465) & (g460)) + ((g455) & (g456) & (g459) & (!g458) & (g465) & (g460)) + ((g455) & (g456) & (g459) & (g458) & (!g465) & (!g460)) + ((g455) & (g456) & (g459) & (g458) & (g465) & (g460)));
	assign g500 = (((!g455) & (!g456) & (!g459) & (!g458) & (g465) & (g460)) + ((!g455) & (!g456) & (!g459) & (g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (!g458) & (!g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (!g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (g459) & (!g458) & (g465) & (g460)) + ((!g455) & (!g456) & (g459) & (g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (g459) & (g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (g459) & (g458) & (g465) & (g460)) + ((!g455) & (g456) & (!g459) & (!g458) & (g465) & (!g460)) + ((!g455) & (g456) & (!g459) & (!g458) & (g465) & (g460)) + ((!g455) & (g456) & (g459) & (!g458) & (!g465) & (!g460)) + ((!g455) & (g456) & (g459) & (g458) & (!g465) & (g460)) + ((!g455) & (g456) & (g459) & (g458) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g458) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (!g458) & (g465) & (g460)) + ((g455) & (!g456) & (!g459) & (g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (g458) & (!g465) & (g460)) + ((g455) & (!g456) & (g459) & (!g458) & (!g465) & (g460)) + ((g455) & (!g456) & (g459) & (!g458) & (g465) & (g460)) + ((g455) & (!g456) & (g459) & (g458) & (g465) & (!g460)) + ((g455) & (g456) & (!g459) & (!g458) & (!g465) & (!g460)) + ((g455) & (g456) & (!g459) & (!g458) & (!g465) & (g460)) + ((g455) & (g456) & (!g459) & (!g458) & (g465) & (g460)) + ((g455) & (g456) & (!g459) & (g458) & (!g465) & (g460)) + ((g455) & (g456) & (!g459) & (g458) & (g465) & (!g460)) + ((g455) & (g456) & (g459) & (!g458) & (!g465) & (g460)) + ((g455) & (g456) & (g459) & (!g458) & (g465) & (!g460)) + ((g455) & (g456) & (g459) & (g458) & (!g465) & (!g460)) + ((g455) & (g456) & (g459) & (g458) & (g465) & (!g460)) + ((g455) & (g456) & (g459) & (g458) & (g465) & (g460)));
	assign g501 = (((!g455) & (!g456) & (!g459) & (!g458) & (g465) & (!g460)) + ((!g455) & (!g456) & (!g459) & (g458) & (!g465) & (!g460)) + ((!g455) & (!g456) & (!g459) & (g458) & (g465) & (g460)) + ((!g455) & (!g456) & (g459) & (!g458) & (!g465) & (g460)) + ((!g455) & (!g456) & (g459) & (!g458) & (g465) & (g460)) + ((!g455) & (!g456) & (g459) & (g458) & (g465) & (g460)) + ((!g455) & (g456) & (!g459) & (!g458) & (!g465) & (g460)) + ((!g455) & (g456) & (!g459) & (g458) & (!g465) & (g460)) + ((!g455) & (g456) & (!g459) & (g458) & (g465) & (g460)) + ((!g455) & (g456) & (g459) & (!g458) & (!g465) & (!g460)) + ((!g455) & (g456) & (g459) & (!g458) & (g465) & (!g460)) + ((!g455) & (g456) & (g459) & (g458) & (!g465) & (g460)) + ((!g455) & (g456) & (g459) & (g458) & (g465) & (g460)) + ((g455) & (!g456) & (!g459) & (!g458) & (g465) & (!g460)) + ((g455) & (!g456) & (!g459) & (g458) & (g465) & (g460)) + ((g455) & (!g456) & (g459) & (!g458) & (!g465) & (!g460)) + ((g455) & (!g456) & (g459) & (!g458) & (g465) & (g460)) + ((g455) & (!g456) & (g459) & (g458) & (!g465) & (!g460)) + ((g455) & (g456) & (!g459) & (!g458) & (g465) & (g460)) + ((g455) & (g456) & (!g459) & (g458) & (!g465) & (!g460)) + ((g455) & (g456) & (!g459) & (g458) & (!g465) & (g460)) + ((g455) & (g456) & (g459) & (!g458) & (g465) & (g460)));
	assign g502 = (((!g498) & (!g499) & (!g500) & (!g501) & (!g466) & (!g457)) + ((!g498) & (!g499) & (!g500) & (!g501) & (!g466) & (g457)) + ((!g498) & (!g499) & (!g500) & (!g501) & (g466) & (!g457)) + ((!g498) & (!g499) & (!g500) & (g501) & (!g466) & (!g457)) + ((!g498) & (!g499) & (!g500) & (g501) & (!g466) & (g457)) + ((!g498) & (!g499) & (!g500) & (g501) & (g466) & (!g457)) + ((!g498) & (!g499) & (!g500) & (g501) & (g466) & (g457)) + ((!g498) & (!g499) & (g500) & (!g501) & (!g466) & (!g457)) + ((!g498) & (!g499) & (g500) & (!g501) & (g466) & (!g457)) + ((!g498) & (!g499) & (g500) & (g501) & (!g466) & (!g457)) + ((!g498) & (!g499) & (g500) & (g501) & (g466) & (!g457)) + ((!g498) & (!g499) & (g500) & (g501) & (g466) & (g457)) + ((!g498) & (g499) & (!g500) & (!g501) & (!g466) & (!g457)) + ((!g498) & (g499) & (!g500) & (!g501) & (!g466) & (g457)) + ((!g498) & (g499) & (!g500) & (g501) & (!g466) & (!g457)) + ((!g498) & (g499) & (!g500) & (g501) & (!g466) & (g457)) + ((!g498) & (g499) & (!g500) & (g501) & (g466) & (g457)) + ((!g498) & (g499) & (g500) & (!g501) & (!g466) & (!g457)) + ((!g498) & (g499) & (g500) & (g501) & (!g466) & (!g457)) + ((!g498) & (g499) & (g500) & (g501) & (g466) & (g457)) + ((g498) & (!g499) & (!g500) & (!g501) & (!g466) & (g457)) + ((g498) & (!g499) & (!g500) & (!g501) & (g466) & (!g457)) + ((g498) & (!g499) & (!g500) & (g501) & (!g466) & (g457)) + ((g498) & (!g499) & (!g500) & (g501) & (g466) & (!g457)) + ((g498) & (!g499) & (!g500) & (g501) & (g466) & (g457)) + ((g498) & (!g499) & (g500) & (!g501) & (g466) & (!g457)) + ((g498) & (!g499) & (g500) & (g501) & (g466) & (!g457)) + ((g498) & (!g499) & (g500) & (g501) & (g466) & (g457)) + ((g498) & (g499) & (!g500) & (!g501) & (!g466) & (g457)) + ((g498) & (g499) & (!g500) & (g501) & (!g466) & (g457)) + ((g498) & (g499) & (!g500) & (g501) & (g466) & (g457)) + ((g498) & (g499) & (g500) & (g501) & (g466) & (g457)));
	assign g504 = (((!sk[20]) & (g502) & (!g503)) + ((!sk[20]) & (g502) & (g503)) + ((sk[20]) & (!g502) & (g503)) + ((sk[20]) & (g502) & (!g503)));
	assign g505 = (((!g455) & (!g466) & (!g457) & (!g458) & (!g465) & (g460)) + ((!g455) & (!g466) & (!g457) & (!g458) & (g465) & (g460)) + ((!g455) & (!g466) & (!g457) & (g458) & (!g465) & (!g460)) + ((!g455) & (!g466) & (!g457) & (g458) & (!g465) & (g460)) + ((!g455) & (!g466) & (!g457) & (g458) & (g465) & (!g460)) + ((!g455) & (!g466) & (!g457) & (g458) & (g465) & (g460)) + ((!g455) & (!g466) & (g457) & (!g458) & (!g465) & (g460)) + ((!g455) & (!g466) & (g457) & (!g458) & (g465) & (g460)) + ((!g455) & (!g466) & (g457) & (g458) & (g465) & (!g460)) + ((!g455) & (g466) & (g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (g466) & (g457) & (!g458) & (g465) & (g460)) + ((!g455) & (g466) & (g457) & (g458) & (!g465) & (g460)) + ((g455) & (!g466) & (!g457) & (!g458) & (g465) & (!g460)) + ((g455) & (!g466) & (!g457) & (g458) & (!g465) & (!g460)) + ((g455) & (!g466) & (!g457) & (g458) & (!g465) & (g460)) + ((g455) & (!g466) & (!g457) & (g458) & (g465) & (g460)) + ((g455) & (!g466) & (g457) & (!g458) & (!g465) & (g460)) + ((g455) & (!g466) & (g457) & (!g458) & (g465) & (g460)) + ((g455) & (!g466) & (g457) & (g458) & (g465) & (!g460)) + ((g455) & (!g466) & (g457) & (g458) & (g465) & (g460)) + ((g455) & (g466) & (!g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (g466) & (!g457) & (!g458) & (!g465) & (g460)) + ((g455) & (g466) & (!g457) & (!g458) & (g465) & (!g460)) + ((g455) & (g466) & (!g457) & (g458) & (!g465) & (!g460)) + ((g455) & (g466) & (g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (g466) & (g457) & (!g458) & (!g465) & (g460)) + ((g455) & (g466) & (g457) & (!g458) & (g465) & (!g460)) + ((g455) & (g466) & (g457) & (g458) & (!g465) & (g460)));
	assign g506 = (((!g455) & (!g466) & (!g457) & (!g458) & (!g465) & (!g460)) + ((!g455) & (!g466) & (!g457) & (g458) & (g465) & (g460)) + ((!g455) & (!g466) & (g457) & (!g458) & (!g465) & (!g460)) + ((!g455) & (!g466) & (g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (!g466) & (g457) & (!g458) & (g465) & (g460)) + ((!g455) & (!g466) & (g457) & (g458) & (!g465) & (!g460)) + ((!g455) & (!g466) & (g457) & (g458) & (g465) & (g460)) + ((!g455) & (g466) & (!g457) & (!g458) & (!g465) & (!g460)) + ((!g455) & (g466) & (!g457) & (!g458) & (g465) & (g460)) + ((!g455) & (g466) & (!g457) & (g458) & (!g465) & (g460)) + ((!g455) & (g466) & (g457) & (!g458) & (!g465) & (!g460)) + ((!g455) & (g466) & (g457) & (!g458) & (g465) & (g460)) + ((!g455) & (g466) & (g457) & (g458) & (g465) & (!g460)) + ((!g455) & (g466) & (g457) & (g458) & (g465) & (g460)) + ((g455) & (!g466) & (!g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (!g466) & (!g457) & (!g458) & (g465) & (g460)) + ((g455) & (!g466) & (!g457) & (g458) & (!g465) & (!g460)) + ((g455) & (!g466) & (!g457) & (g458) & (g465) & (g460)) + ((g455) & (!g466) & (g457) & (!g458) & (g465) & (g460)) + ((g455) & (!g466) & (g457) & (g458) & (!g465) & (g460)) + ((g455) & (g466) & (!g457) & (!g458) & (g465) & (!g460)) + ((g455) & (g466) & (!g457) & (!g458) & (g465) & (g460)) + ((g455) & (g466) & (!g457) & (g458) & (!g465) & (g460)) + ((g455) & (g466) & (!g457) & (g458) & (g465) & (!g460)) + ((g455) & (g466) & (!g457) & (g458) & (g465) & (g460)) + ((g455) & (g466) & (g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (g466) & (g457) & (!g458) & (g465) & (!g460)) + ((g455) & (g466) & (g457) & (g458) & (!g465) & (!g460)));
	assign g507 = (((!g455) & (!g466) & (!g457) & (!g458) & (!g465) & (g460)) + ((!g455) & (!g466) & (!g457) & (!g458) & (g465) & (g460)) + ((!g455) & (!g466) & (!g457) & (g458) & (g465) & (!g460)) + ((!g455) & (!g466) & (!g457) & (g458) & (g465) & (g460)) + ((!g455) & (!g466) & (g457) & (!g458) & (g465) & (g460)) + ((!g455) & (!g466) & (g457) & (g458) & (!g465) & (!g460)) + ((!g455) & (!g466) & (g457) & (g458) & (!g465) & (g460)) + ((!g455) & (!g466) & (g457) & (g458) & (g465) & (g460)) + ((!g455) & (g466) & (!g457) & (!g458) & (!g465) & (!g460)) + ((!g455) & (g466) & (!g457) & (!g458) & (!g465) & (g460)) + ((!g455) & (g466) & (!g457) & (!g458) & (g465) & (g460)) + ((!g455) & (g466) & (!g457) & (g458) & (!g465) & (g460)) + ((!g455) & (g466) & (!g457) & (g458) & (g465) & (!g460)) + ((!g455) & (g466) & (g457) & (!g458) & (!g465) & (g460)) + ((!g455) & (g466) & (g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (g466) & (g457) & (g458) & (!g465) & (!g460)) + ((!g455) & (g466) & (g457) & (g458) & (g465) & (!g460)) + ((!g455) & (g466) & (g457) & (g458) & (g465) & (g460)) + ((g455) & (!g466) & (!g457) & (!g458) & (!g465) & (g460)) + ((g455) & (!g466) & (!g457) & (g458) & (!g465) & (!g460)) + ((g455) & (!g466) & (!g457) & (g458) & (g465) & (!g460)) + ((g455) & (!g466) & (g457) & (!g458) & (g465) & (g460)) + ((g455) & (!g466) & (g457) & (g458) & (!g465) & (g460)) + ((g455) & (g466) & (!g457) & (!g458) & (!g465) & (g460)) + ((g455) & (g466) & (!g457) & (g458) & (!g465) & (!g460)) + ((g455) & (g466) & (!g457) & (g458) & (g465) & (!g460)) + ((g455) & (g466) & (g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (g466) & (g457) & (!g458) & (g465) & (!g460)) + ((g455) & (g466) & (g457) & (!g458) & (g465) & (g460)) + ((g455) & (g466) & (g457) & (g458) & (g465) & (g460)));
	assign g508 = (((!g455) & (!g466) & (!g457) & (!g458) & (g465) & (g460)) + ((!g455) & (!g466) & (!g457) & (g458) & (!g465) & (!g460)) + ((!g455) & (!g466) & (!g457) & (g458) & (g465) & (g460)) + ((!g455) & (!g466) & (g457) & (!g458) & (!g465) & (!g460)) + ((!g455) & (!g466) & (g457) & (g458) & (g465) & (!g460)) + ((!g455) & (!g466) & (g457) & (g458) & (g465) & (g460)) + ((!g455) & (g466) & (!g457) & (g458) & (!g465) & (!g460)) + ((!g455) & (g466) & (!g457) & (g458) & (g465) & (!g460)) + ((!g455) & (g466) & (g457) & (!g458) & (g465) & (!g460)) + ((!g455) & (g466) & (g457) & (!g458) & (g465) & (g460)) + ((g455) & (!g466) & (!g457) & (!g458) & (!g465) & (g460)) + ((g455) & (!g466) & (!g457) & (!g458) & (g465) & (!g460)) + ((g455) & (!g466) & (!g457) & (g458) & (!g465) & (g460)) + ((g455) & (!g466) & (g457) & (!g458) & (g465) & (!g460)) + ((g455) & (!g466) & (g457) & (!g458) & (g465) & (g460)) + ((g455) & (!g466) & (g457) & (g458) & (g465) & (!g460)) + ((g455) & (!g466) & (g457) & (g458) & (g465) & (g460)) + ((g455) & (g466) & (!g457) & (!g458) & (g465) & (!g460)) + ((g455) & (g466) & (!g457) & (g458) & (!g465) & (g460)) + ((g455) & (g466) & (g457) & (!g458) & (!g465) & (!g460)) + ((g455) & (g466) & (g457) & (!g458) & (g465) & (g460)) + ((g455) & (g466) & (g457) & (g458) & (!g465) & (g460)));
	assign g509 = (((!g505) & (!g506) & (!g507) & (!g508) & (!g459) & (!g456)) + ((!g505) & (!g506) & (!g507) & (!g508) & (!g459) & (g456)) + ((!g505) & (!g506) & (!g507) & (!g508) & (g459) & (!g456)) + ((!g505) & (!g506) & (!g507) & (g508) & (!g459) & (!g456)) + ((!g505) & (!g506) & (!g507) & (g508) & (!g459) & (g456)) + ((!g505) & (!g506) & (!g507) & (g508) & (g459) & (!g456)) + ((!g505) & (!g506) & (!g507) & (g508) & (g459) & (g456)) + ((!g505) & (!g506) & (g507) & (!g508) & (!g459) & (!g456)) + ((!g505) & (!g506) & (g507) & (!g508) & (g459) & (!g456)) + ((!g505) & (!g506) & (g507) & (g508) & (!g459) & (!g456)) + ((!g505) & (!g506) & (g507) & (g508) & (g459) & (!g456)) + ((!g505) & (!g506) & (g507) & (g508) & (g459) & (g456)) + ((!g505) & (g506) & (!g507) & (!g508) & (!g459) & (!g456)) + ((!g505) & (g506) & (!g507) & (!g508) & (!g459) & (g456)) + ((!g505) & (g506) & (!g507) & (g508) & (!g459) & (!g456)) + ((!g505) & (g506) & (!g507) & (g508) & (!g459) & (g456)) + ((!g505) & (g506) & (!g507) & (g508) & (g459) & (g456)) + ((!g505) & (g506) & (g507) & (!g508) & (!g459) & (!g456)) + ((!g505) & (g506) & (g507) & (g508) & (!g459) & (!g456)) + ((!g505) & (g506) & (g507) & (g508) & (g459) & (g456)) + ((g505) & (!g506) & (!g507) & (!g508) & (!g459) & (g456)) + ((g505) & (!g506) & (!g507) & (!g508) & (g459) & (!g456)) + ((g505) & (!g506) & (!g507) & (g508) & (!g459) & (g456)) + ((g505) & (!g506) & (!g507) & (g508) & (g459) & (!g456)) + ((g505) & (!g506) & (!g507) & (g508) & (g459) & (g456)) + ((g505) & (!g506) & (g507) & (!g508) & (g459) & (!g456)) + ((g505) & (!g506) & (g507) & (g508) & (g459) & (!g456)) + ((g505) & (!g506) & (g507) & (g508) & (g459) & (g456)) + ((g505) & (g506) & (!g507) & (!g508) & (!g459) & (g456)) + ((g505) & (g506) & (!g507) & (g508) & (!g459) & (g456)) + ((g505) & (g506) & (!g507) & (g508) & (g459) & (g456)) + ((g505) & (g506) & (g507) & (g508) & (g459) & (g456)));
	assign g511 = (((!sk[26]) & (g509) & (!g510)) + ((!sk[26]) & (g509) & (g510)) + ((sk[26]) & (!g509) & (g510)) + ((sk[26]) & (g509) & (!g510)));
	assign g512 = (((!g459) & (!g456) & (!g457) & (!g458) & (!g465) & (g466)) + ((!g459) & (!g456) & (!g457) & (!g458) & (g465) & (!g466)) + ((!g459) & (!g456) & (!g457) & (g458) & (!g465) & (g466)) + ((!g459) & (!g456) & (!g457) & (g458) & (g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (!g458) & (!g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (!g458) & (g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (g458) & (!g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (g458) & (g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (g458) & (g465) & (g466)) + ((!g459) & (g456) & (!g457) & (!g458) & (g465) & (!g466)) + ((!g459) & (g456) & (!g457) & (g458) & (g465) & (!g466)) + ((!g459) & (g456) & (!g457) & (g458) & (g465) & (g466)) + ((!g459) & (g456) & (g457) & (!g458) & (g465) & (g466)) + ((!g459) & (g456) & (g457) & (g458) & (!g465) & (!g466)) + ((g459) & (!g456) & (!g457) & (!g458) & (!g465) & (g466)) + ((g459) & (!g456) & (!g457) & (g458) & (!g465) & (g466)) + ((g459) & (!g456) & (g457) & (g458) & (g465) & (g466)) + ((g459) & (g456) & (!g457) & (!g458) & (g465) & (g466)) + ((g459) & (g456) & (!g457) & (g458) & (!g465) & (!g466)) + ((g459) & (g456) & (!g457) & (g458) & (g465) & (!g466)) + ((g459) & (g456) & (g457) & (!g458) & (!g465) & (g466)) + ((g459) & (g456) & (g457) & (!g458) & (g465) & (!g466)) + ((g459) & (g456) & (g457) & (!g458) & (g465) & (g466)) + ((g459) & (g456) & (g457) & (g458) & (!g465) & (g466)));
	assign g513 = (((!g459) & (!g456) & (!g457) & (!g458) & (!g465) & (!g466)) + ((!g459) & (!g456) & (!g457) & (!g458) & (!g465) & (g466)) + ((!g459) & (!g456) & (!g457) & (g458) & (!g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (!g458) & (!g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (!g458) & (g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (!g458) & (g465) & (g466)) + ((!g459) & (!g456) & (g457) & (g458) & (!g465) & (g466)) + ((!g459) & (!g456) & (g457) & (g458) & (g465) & (g466)) + ((!g459) & (g456) & (!g457) & (!g458) & (!g465) & (!g466)) + ((!g459) & (g456) & (!g457) & (!g458) & (g465) & (!g466)) + ((!g459) & (g456) & (!g457) & (g458) & (!g465) & (!g466)) + ((!g459) & (g456) & (!g457) & (g458) & (!g465) & (g466)) + ((!g459) & (g456) & (!g457) & (g458) & (g465) & (g466)) + ((!g459) & (g456) & (g457) & (!g458) & (!g465) & (g466)) + ((!g459) & (g456) & (g457) & (g458) & (!g465) & (!g466)) + ((!g459) & (g456) & (g457) & (g458) & (!g465) & (g466)) + ((g459) & (!g456) & (!g457) & (!g458) & (!g465) & (g466)) + ((g459) & (!g456) & (!g457) & (!g458) & (g465) & (g466)) + ((g459) & (!g456) & (!g457) & (g458) & (!g465) & (!g466)) + ((g459) & (!g456) & (!g457) & (g458) & (g465) & (g466)) + ((g459) & (!g456) & (g457) & (!g458) & (!g465) & (!g466)) + ((g459) & (!g456) & (g457) & (!g458) & (g465) & (g466)) + ((g459) & (!g456) & (g457) & (g458) & (g465) & (!g466)) + ((g459) & (g456) & (!g457) & (!g458) & (!g465) & (!g466)) + ((g459) & (g456) & (!g457) & (!g458) & (!g465) & (g466)) + ((g459) & (g456) & (!g457) & (!g458) & (g465) & (g466)) + ((g459) & (g456) & (!g457) & (g458) & (!g465) & (g466)) + ((g459) & (g456) & (!g457) & (g458) & (g465) & (!g466)) + ((g459) & (g456) & (g457) & (!g458) & (g465) & (!g466)) + ((g459) & (g456) & (g457) & (!g458) & (g465) & (g466)));
	assign g514 = (((!g459) & (!g456) & (!g457) & (!g458) & (g465) & (!g466)) + ((!g459) & (!g456) & (!g457) & (g458) & (!g465) & (!g466)) + ((!g459) & (!g456) & (!g457) & (g458) & (g465) & (!g466)) + ((!g459) & (!g456) & (!g457) & (g458) & (g465) & (g466)) + ((!g459) & (!g456) & (g457) & (!g458) & (!g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (!g458) & (!g465) & (g466)) + ((!g459) & (!g456) & (g457) & (!g458) & (g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (g458) & (!g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (g458) & (g465) & (g466)) + ((!g459) & (g456) & (!g457) & (!g458) & (!g465) & (g466)) + ((!g459) & (g456) & (!g457) & (!g458) & (g465) & (!g466)) + ((!g459) & (g456) & (!g457) & (!g458) & (g465) & (g466)) + ((!g459) & (g456) & (g457) & (!g458) & (!g465) & (g466)) + ((!g459) & (g456) & (g457) & (!g458) & (g465) & (!g466)) + ((!g459) & (g456) & (g457) & (!g458) & (g465) & (g466)) + ((!g459) & (g456) & (g457) & (g458) & (!g465) & (!g466)) + ((g459) & (!g456) & (!g457) & (!g458) & (g465) & (!g466)) + ((g459) & (!g456) & (!g457) & (g458) & (!g465) & (!g466)) + ((g459) & (!g456) & (!g457) & (g458) & (g465) & (g466)) + ((g459) & (!g456) & (g457) & (!g458) & (!g465) & (!g466)) + ((g459) & (!g456) & (g457) & (!g458) & (!g465) & (g466)) + ((g459) & (!g456) & (g457) & (g458) & (!g465) & (!g466)) + ((g459) & (!g456) & (g457) & (g458) & (g465) & (!g466)) + ((g459) & (g456) & (!g457) & (!g458) & (g465) & (!g466)) + ((g459) & (g456) & (!g457) & (g458) & (!g465) & (!g466)) + ((g459) & (g456) & (!g457) & (g458) & (g465) & (g466)) + ((g459) & (g456) & (g457) & (!g458) & (!g465) & (!g466)) + ((g459) & (g456) & (g457) & (!g458) & (g465) & (!g466)) + ((g459) & (g456) & (g457) & (!g458) & (g465) & (g466)) + ((g459) & (g456) & (g457) & (g458) & (!g465) & (g466)));
	assign g515 = (((!g459) & (!g456) & (!g457) & (!g458) & (!g465) & (g466)) + ((!g459) & (!g456) & (!g457) & (g458) & (g465) & (!g466)) + ((!g459) & (!g456) & (!g457) & (g458) & (g465) & (g466)) + ((!g459) & (!g456) & (g457) & (!g458) & (!g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (!g458) & (!g465) & (g466)) + ((!g459) & (!g456) & (g457) & (g458) & (g465) & (!g466)) + ((!g459) & (!g456) & (g457) & (g458) & (g465) & (g466)) + ((!g459) & (g456) & (!g457) & (!g458) & (!g465) & (!g466)) + ((!g459) & (g456) & (!g457) & (!g458) & (!g465) & (g466)) + ((!g459) & (g456) & (!g457) & (!g458) & (g465) & (g466)) + ((!g459) & (g456) & (!g457) & (g458) & (!g465) & (g466)) + ((!g459) & (g456) & (g457) & (!g458) & (!g465) & (g466)) + ((!g459) & (g456) & (g457) & (g458) & (!g465) & (!g466)) + ((!g459) & (g456) & (g457) & (g458) & (!g465) & (g466)) + ((!g459) & (g456) & (g457) & (g458) & (g465) & (!g466)) + ((!g459) & (g456) & (g457) & (g458) & (g465) & (g466)) + ((g459) & (!g456) & (!g457) & (g458) & (!g465) & (g466)) + ((g459) & (!g456) & (g457) & (!g458) & (!g465) & (!g466)) + ((g459) & (!g456) & (g457) & (g458) & (!g465) & (!g466)) + ((g459) & (!g456) & (g457) & (g458) & (!g465) & (g466)) + ((g459) & (!g456) & (g457) & (g458) & (g465) & (g466)) + ((g459) & (g456) & (!g457) & (!g458) & (!g465) & (g466)) + ((g459) & (g456) & (!g457) & (!g458) & (g465) & (g466)) + ((g459) & (g456) & (!g457) & (g458) & (!g465) & (!g466)) + ((g459) & (g456) & (!g457) & (g458) & (g465) & (!g466)) + ((g459) & (g456) & (!g457) & (g458) & (g465) & (g466)) + ((g459) & (g456) & (g457) & (!g458) & (g465) & (g466)) + ((g459) & (g456) & (g457) & (g458) & (g465) & (g466)));
	assign g516 = (((!g512) & (!g513) & (!g514) & (!g515) & (!g455) & (g460)) + ((!g512) & (!g513) & (!g514) & (!g515) & (g455) & (!g460)) + ((!g512) & (!g513) & (!g514) & (!g515) & (g455) & (g460)) + ((!g512) & (!g513) & (!g514) & (g515) & (!g455) & (g460)) + ((!g512) & (!g513) & (!g514) & (g515) & (g455) & (!g460)) + ((!g512) & (!g513) & (g514) & (!g515) & (g455) & (!g460)) + ((!g512) & (!g513) & (g514) & (!g515) & (g455) & (g460)) + ((!g512) & (!g513) & (g514) & (g515) & (g455) & (!g460)) + ((!g512) & (g513) & (!g514) & (!g515) & (!g455) & (g460)) + ((!g512) & (g513) & (!g514) & (!g515) & (g455) & (g460)) + ((!g512) & (g513) & (!g514) & (g515) & (!g455) & (g460)) + ((!g512) & (g513) & (g514) & (!g515) & (g455) & (g460)) + ((g512) & (!g513) & (!g514) & (!g515) & (!g455) & (!g460)) + ((g512) & (!g513) & (!g514) & (!g515) & (!g455) & (g460)) + ((g512) & (!g513) & (!g514) & (!g515) & (g455) & (!g460)) + ((g512) & (!g513) & (!g514) & (!g515) & (g455) & (g460)) + ((g512) & (!g513) & (!g514) & (g515) & (!g455) & (!g460)) + ((g512) & (!g513) & (!g514) & (g515) & (!g455) & (g460)) + ((g512) & (!g513) & (!g514) & (g515) & (g455) & (!g460)) + ((g512) & (!g513) & (g514) & (!g515) & (!g455) & (!g460)) + ((g512) & (!g513) & (g514) & (!g515) & (g455) & (!g460)) + ((g512) & (!g513) & (g514) & (!g515) & (g455) & (g460)) + ((g512) & (!g513) & (g514) & (g515) & (!g455) & (!g460)) + ((g512) & (!g513) & (g514) & (g515) & (g455) & (!g460)) + ((g512) & (g513) & (!g514) & (!g515) & (!g455) & (!g460)) + ((g512) & (g513) & (!g514) & (!g515) & (!g455) & (g460)) + ((g512) & (g513) & (!g514) & (!g515) & (g455) & (g460)) + ((g512) & (g513) & (!g514) & (g515) & (!g455) & (!g460)) + ((g512) & (g513) & (!g514) & (g515) & (!g455) & (g460)) + ((g512) & (g513) & (g514) & (!g515) & (!g455) & (!g460)) + ((g512) & (g513) & (g514) & (!g515) & (g455) & (g460)) + ((g512) & (g513) & (g514) & (g515) & (!g455) & (!g460)));
	assign g518 = (((!g516) & (sk[32]) & (g517)) + ((g516) & (!sk[32]) & (!g517)) + ((g516) & (!sk[32]) & (g517)) + ((g516) & (sk[32]) & (!g517)));
	assign g525 = (((!g519) & (!g520) & (!g521) & (!g522) & (g523) & (g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g523) & (!g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g523) & (g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (g523) & (!g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (!g523) & (!g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (!g523) & (g524)) + ((!g519) & (!g520) & (g521) & (g522) & (!g523) & (!g524)) + ((!g519) & (!g520) & (g521) & (g522) & (g523) & (g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (g523) & (!g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (g523) & (g524)) + ((!g519) & (g520) & (!g521) & (g522) & (g523) & (!g524)) + ((!g519) & (g520) & (!g521) & (g522) & (g523) & (g524)) + ((!g519) & (g520) & (g521) & (!g522) & (g523) & (!g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (!g523) & (!g524)) + ((g519) & (!g520) & (g521) & (!g522) & (g523) & (!g524)) + ((g519) & (!g520) & (g521) & (g522) & (!g523) & (g524)) + ((g519) & (!g520) & (g521) & (g522) & (g523) & (g524)) + ((g519) & (g520) & (!g521) & (!g522) & (!g523) & (g524)) + ((g519) & (g520) & (!g521) & (!g522) & (g523) & (!g524)) + ((g519) & (g520) & (g521) & (!g522) & (!g523) & (g524)) + ((g519) & (g520) & (g521) & (!g522) & (g523) & (!g524)) + ((g519) & (g520) & (g521) & (g522) & (!g523) & (!g524)) + ((g519) & (g520) & (g521) & (g522) & (g523) & (!g524)) + ((g519) & (g520) & (g521) & (g522) & (g523) & (g524)));
	assign g526 = (((!g519) & (!g520) & (!g521) & (!g522) & (g523) & (!g524)) + ((!g519) & (!g520) & (!g521) & (!g522) & (g523) & (g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g523) & (!g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g523) & (g524)) + ((!g519) & (!g520) & (g521) & (g522) & (!g523) & (g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (!g523) & (!g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (!g523) & (g524)) + ((!g519) & (g520) & (g521) & (!g522) & (!g523) & (!g524)) + ((!g519) & (g520) & (g521) & (!g522) & (!g523) & (g524)) + ((!g519) & (g520) & (g521) & (!g522) & (g523) & (!g524)) + ((!g519) & (g520) & (g521) & (g522) & (g523) & (g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (!g523) & (g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (g523) & (!g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (g523) & (g524)) + ((g519) & (!g520) & (!g521) & (g522) & (g523) & (!g524)) + ((g519) & (!g520) & (g521) & (!g522) & (!g523) & (!g524)) + ((g519) & (!g520) & (g521) & (!g522) & (g523) & (g524)) + ((g519) & (!g520) & (g521) & (g522) & (!g523) & (g524)) + ((g519) & (!g520) & (g521) & (g522) & (g523) & (g524)) + ((g519) & (g520) & (!g521) & (!g522) & (!g523) & (!g524)) + ((g519) & (g520) & (!g521) & (!g522) & (!g523) & (g524)) + ((g519) & (g520) & (!g521) & (!g522) & (g523) & (!g524)) + ((g519) & (g520) & (!g521) & (!g522) & (g523) & (g524)) + ((g519) & (g520) & (!g521) & (g522) & (!g523) & (!g524)) + ((g519) & (g520) & (!g521) & (g522) & (g523) & (!g524)) + ((g519) & (g520) & (!g521) & (g522) & (g523) & (g524)) + ((g519) & (g520) & (g521) & (!g522) & (g523) & (!g524)) + ((g519) & (g520) & (g521) & (!g522) & (g523) & (g524)) + ((g519) & (g520) & (g521) & (g522) & (!g523) & (g524)) + ((g519) & (g520) & (g521) & (g522) & (g523) & (!g524)));
	assign g527 = (((!g519) & (!g520) & (!g521) & (!g522) & (!g523) & (!g524)) + ((!g519) & (!g520) & (!g521) & (!g522) & (g523) & (g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (g523) & (g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (!g523) & (!g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (!g523) & (g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (g523) & (g524)) + ((!g519) & (!g520) & (g521) & (g522) & (!g523) & (g524)) + ((!g519) & (!g520) & (g521) & (g522) & (g523) & (!g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (!g523) & (!g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (g523) & (!g524)) + ((!g519) & (g520) & (!g521) & (g522) & (g523) & (g524)) + ((!g519) & (g520) & (g521) & (g522) & (!g523) & (!g524)) + ((!g519) & (g520) & (g521) & (g522) & (g523) & (!g524)) + ((g519) & (!g520) & (!g521) & (g522) & (!g523) & (!g524)) + ((g519) & (!g520) & (!g521) & (g522) & (!g523) & (g524)) + ((g519) & (!g520) & (!g521) & (g522) & (g523) & (!g524)) + ((g519) & (!g520) & (g521) & (!g522) & (!g523) & (!g524)) + ((g519) & (!g520) & (g521) & (!g522) & (g523) & (g524)) + ((g519) & (!g520) & (g521) & (g522) & (!g523) & (!g524)) + ((g519) & (!g520) & (g521) & (g522) & (!g523) & (g524)) + ((g519) & (!g520) & (g521) & (g522) & (g523) & (!g524)) + ((g519) & (!g520) & (g521) & (g522) & (g523) & (g524)) + ((g519) & (g520) & (!g521) & (!g522) & (g523) & (g524)) + ((g519) & (g520) & (!g521) & (g522) & (!g523) & (!g524)) + ((g519) & (g520) & (!g521) & (g522) & (g523) & (!g524)) + ((g519) & (g520) & (!g521) & (g522) & (g523) & (g524)) + ((g519) & (g520) & (g521) & (!g522) & (!g523) & (!g524)) + ((g519) & (g520) & (g521) & (g522) & (!g523) & (!g524)) + ((g519) & (g520) & (g521) & (g522) & (!g523) & (g524)) + ((g519) & (g520) & (g521) & (g522) & (g523) & (g524)));
	assign g528 = (((!g519) & (!g520) & (!g521) & (!g522) & (!g523) & (g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (g523) & (!g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (g523) & (g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (!g523) & (g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (g523) & (g524)) + ((!g519) & (!g520) & (g521) & (g522) & (!g523) & (g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (!g523) & (!g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (!g523) & (g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (g523) & (!g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (g523) & (g524)) + ((!g519) & (g520) & (!g521) & (g522) & (g523) & (!g524)) + ((!g519) & (g520) & (!g521) & (g522) & (g523) & (g524)) + ((!g519) & (g520) & (g521) & (g522) & (!g523) & (!g524)) + ((!g519) & (g520) & (g521) & (g522) & (g523) & (!g524)) + ((!g519) & (g520) & (g521) & (g522) & (g523) & (g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (!g523) & (!g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (g523) & (g524)) + ((g519) & (!g520) & (!g521) & (g522) & (g523) & (!g524)) + ((g519) & (!g520) & (!g521) & (g522) & (g523) & (g524)) + ((g519) & (!g520) & (g521) & (!g522) & (!g523) & (g524)) + ((g519) & (!g520) & (g521) & (!g522) & (g523) & (!g524)) + ((g519) & (!g520) & (g521) & (g522) & (g523) & (!g524)) + ((g519) & (g520) & (!g521) & (!g522) & (!g523) & (g524)) + ((g519) & (g520) & (!g521) & (!g522) & (g523) & (g524)) + ((g519) & (g520) & (!g521) & (g522) & (g523) & (!g524)) + ((g519) & (g520) & (!g521) & (g522) & (g523) & (g524)) + ((g519) & (g520) & (g521) & (!g522) & (!g523) & (g524)) + ((g519) & (g520) & (g521) & (g522) & (!g523) & (!g524)));
	assign g531 = (((!g525) & (!g526) & (!g527) & (!g528) & (!g529) & (!g530)) + ((!g525) & (!g526) & (!g527) & (g528) & (!g529) & (!g530)) + ((!g525) & (!g526) & (!g527) & (g528) & (g529) & (g530)) + ((!g525) & (!g526) & (g527) & (!g528) & (!g529) & (!g530)) + ((!g525) & (!g526) & (g527) & (!g528) & (!g529) & (g530)) + ((!g525) & (!g526) & (g527) & (g528) & (!g529) & (!g530)) + ((!g525) & (!g526) & (g527) & (g528) & (!g529) & (g530)) + ((!g525) & (!g526) & (g527) & (g528) & (g529) & (g530)) + ((!g525) & (g526) & (!g527) & (!g528) & (!g529) & (!g530)) + ((!g525) & (g526) & (!g527) & (!g528) & (g529) & (!g530)) + ((!g525) & (g526) & (!g527) & (g528) & (!g529) & (!g530)) + ((!g525) & (g526) & (!g527) & (g528) & (g529) & (!g530)) + ((!g525) & (g526) & (!g527) & (g528) & (g529) & (g530)) + ((!g525) & (g526) & (g527) & (!g528) & (!g529) & (!g530)) + ((!g525) & (g526) & (g527) & (!g528) & (!g529) & (g530)) + ((!g525) & (g526) & (g527) & (!g528) & (g529) & (!g530)) + ((!g525) & (g526) & (g527) & (g528) & (!g529) & (!g530)) + ((!g525) & (g526) & (g527) & (g528) & (!g529) & (g530)) + ((!g525) & (g526) & (g527) & (g528) & (g529) & (!g530)) + ((!g525) & (g526) & (g527) & (g528) & (g529) & (g530)) + ((g525) & (!g526) & (!g527) & (g528) & (g529) & (g530)) + ((g525) & (!g526) & (g527) & (!g528) & (!g529) & (g530)) + ((g525) & (!g526) & (g527) & (g528) & (!g529) & (g530)) + ((g525) & (!g526) & (g527) & (g528) & (g529) & (g530)) + ((g525) & (g526) & (!g527) & (!g528) & (g529) & (!g530)) + ((g525) & (g526) & (!g527) & (g528) & (g529) & (!g530)) + ((g525) & (g526) & (!g527) & (g528) & (g529) & (g530)) + ((g525) & (g526) & (g527) & (!g528) & (!g529) & (g530)) + ((g525) & (g526) & (g527) & (!g528) & (g529) & (!g530)) + ((g525) & (g526) & (g527) & (g528) & (!g529) & (g530)) + ((g525) & (g526) & (g527) & (g528) & (g529) & (!g530)) + ((g525) & (g526) & (g527) & (g528) & (g529) & (g530)));
	assign g533 = (((!sk[38]) & (g531) & (!g532)) + ((!sk[38]) & (g531) & (g532)) + ((sk[38]) & (!g531) & (g532)) + ((sk[38]) & (g531) & (!g532)));
	assign g534 = (((!g519) & (!g520) & (!g521) & (!g522) & (!g529) & (g523)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g529) & (!g523)) + ((!g519) & (!g520) & (!g521) & (g522) & (g529) & (!g523)) + ((!g519) & (!g520) & (g521) & (!g522) & (g529) & (g523)) + ((!g519) & (!g520) & (g521) & (g522) & (!g529) & (g523)) + ((!g519) & (!g520) & (g521) & (g522) & (g529) & (!g523)) + ((!g519) & (g520) & (!g521) & (!g522) & (!g529) & (g523)) + ((!g519) & (g520) & (!g521) & (!g522) & (g529) & (!g523)) + ((!g519) & (g520) & (!g521) & (!g522) & (g529) & (g523)) + ((!g519) & (g520) & (g521) & (!g522) & (g529) & (g523)) + ((!g519) & (g520) & (g521) & (g522) & (g529) & (g523)) + ((g519) & (!g520) & (!g521) & (!g522) & (!g529) & (!g523)) + ((g519) & (!g520) & (!g521) & (!g522) & (g529) & (g523)) + ((g519) & (!g520) & (!g521) & (g522) & (!g529) & (!g523)) + ((g519) & (!g520) & (!g521) & (g522) & (g529) & (!g523)) + ((g519) & (!g520) & (g521) & (!g522) & (g529) & (!g523)) + ((g519) & (!g520) & (g521) & (!g522) & (g529) & (g523)) + ((g519) & (!g520) & (g521) & (g522) & (g529) & (!g523)) + ((g519) & (!g520) & (g521) & (g522) & (g529) & (g523)) + ((g519) & (g520) & (!g521) & (!g522) & (g529) & (!g523)) + ((g519) & (g520) & (!g521) & (!g522) & (g529) & (g523)) + ((g519) & (g520) & (!g521) & (g522) & (g529) & (g523)) + ((g519) & (g520) & (g521) & (!g522) & (!g529) & (!g523)) + ((g519) & (g520) & (g521) & (!g522) & (!g529) & (g523)) + ((g519) & (g520) & (g521) & (!g522) & (g529) & (!g523)) + ((g519) & (g520) & (g521) & (g522) & (!g529) & (g523)) + ((g519) & (g520) & (g521) & (g522) & (g529) & (!g523)));
	assign g535 = (((!g519) & (!g520) & (!g521) & (!g522) & (!g529) & (g523)) + ((!g519) & (!g520) & (!g521) & (!g522) & (g529) & (!g523)) + ((!g519) & (!g520) & (!g521) & (!g522) & (g529) & (g523)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g529) & (!g523)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g529) & (g523)) + ((!g519) & (!g520) & (!g521) & (g522) & (g529) & (g523)) + ((!g519) & (!g520) & (g521) & (!g522) & (g529) & (!g523)) + ((!g519) & (!g520) & (g521) & (g522) & (!g529) & (!g523)) + ((!g519) & (!g520) & (g521) & (g522) & (!g529) & (g523)) + ((!g519) & (!g520) & (g521) & (g522) & (g529) & (g523)) + ((!g519) & (g520) & (!g521) & (!g522) & (g529) & (g523)) + ((!g519) & (g520) & (!g521) & (g522) & (!g529) & (!g523)) + ((!g519) & (g520) & (!g521) & (g522) & (g529) & (!g523)) + ((!g519) & (g520) & (g521) & (!g522) & (g529) & (!g523)) + ((!g519) & (g520) & (g521) & (!g522) & (g529) & (g523)) + ((!g519) & (g520) & (g521) & (g522) & (!g529) & (!g523)) + ((g519) & (!g520) & (!g521) & (!g522) & (!g529) & (!g523)) + ((g519) & (!g520) & (!g521) & (g522) & (!g529) & (!g523)) + ((g519) & (!g520) & (!g521) & (g522) & (!g529) & (g523)) + ((g519) & (!g520) & (g521) & (!g522) & (!g529) & (g523)) + ((g519) & (!g520) & (g521) & (!g522) & (g529) & (g523)) + ((g519) & (!g520) & (g521) & (g522) & (!g529) & (!g523)) + ((g519) & (!g520) & (g521) & (g522) & (!g529) & (g523)) + ((g519) & (g520) & (!g521) & (g522) & (!g529) & (!g523)) + ((g519) & (g520) & (!g521) & (g522) & (g529) & (g523)) + ((g519) & (g520) & (g521) & (!g522) & (!g529) & (!g523)) + ((g519) & (g520) & (g521) & (!g522) & (!g529) & (g523)) + ((g519) & (g520) & (g521) & (!g522) & (g529) & (g523)) + ((g519) & (g520) & (g521) & (g522) & (!g529) & (!g523)) + ((g519) & (g520) & (g521) & (g522) & (!g529) & (g523)) + ((g519) & (g520) & (g521) & (g522) & (g529) & (!g523)));
	assign g536 = (((!g519) & (!g520) & (!g521) & (!g522) & (!g529) & (g523)) + ((!g519) & (!g520) & (!g521) & (g522) & (g529) & (!g523)) + ((!g519) & (!g520) & (g521) & (!g522) & (!g529) & (!g523)) + ((!g519) & (!g520) & (g521) & (!g522) & (g529) & (!g523)) + ((!g519) & (!g520) & (g521) & (g522) & (!g529) & (g523)) + ((!g519) & (!g520) & (g521) & (g522) & (g529) & (!g523)) + ((!g519) & (!g520) & (g521) & (g522) & (g529) & (g523)) + ((!g519) & (g520) & (!g521) & (!g522) & (!g529) & (!g523)) + ((!g519) & (g520) & (!g521) & (!g522) & (g529) & (!g523)) + ((!g519) & (g520) & (!g521) & (g522) & (!g529) & (!g523)) + ((!g519) & (g520) & (!g521) & (g522) & (g529) & (g523)) + ((!g519) & (g520) & (g521) & (!g522) & (g529) & (g523)) + ((!g519) & (g520) & (g521) & (g522) & (!g529) & (g523)) + ((!g519) & (g520) & (g521) & (g522) & (g529) & (!g523)) + ((g519) & (!g520) & (!g521) & (!g522) & (g529) & (g523)) + ((g519) & (!g520) & (!g521) & (g522) & (!g529) & (!g523)) + ((g519) & (!g520) & (!g521) & (g522) & (g529) & (!g523)) + ((g519) & (!g520) & (g521) & (!g522) & (!g529) & (!g523)) + ((g519) & (!g520) & (g521) & (!g522) & (!g529) & (g523)) + ((g519) & (!g520) & (g521) & (!g522) & (g529) & (!g523)) + ((g519) & (!g520) & (g521) & (!g522) & (g529) & (g523)) + ((g519) & (!g520) & (g521) & (g522) & (g529) & (!g523)) + ((g519) & (g520) & (!g521) & (!g522) & (!g529) & (g523)) + ((g519) & (g520) & (!g521) & (!g522) & (g529) & (g523)) + ((g519) & (g520) & (!g521) & (g522) & (!g529) & (g523)) + ((g519) & (g520) & (g521) & (!g522) & (!g529) & (!g523)) + ((g519) & (g520) & (g521) & (!g522) & (!g529) & (g523)) + ((g519) & (g520) & (g521) & (!g522) & (g529) & (g523)) + ((g519) & (g520) & (g521) & (g522) & (!g529) & (!g523)) + ((g519) & (g520) & (g521) & (g522) & (!g529) & (g523)) + ((g519) & (g520) & (g521) & (g522) & (g529) & (!g523)) + ((g519) & (g520) & (g521) & (g522) & (g529) & (g523)));
	assign g537 = (((!g519) & (!g520) & (!g521) & (!g522) & (g529) & (!g523)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g529) & (!g523)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g529) & (g523)) + ((!g519) & (!g520) & (g521) & (!g522) & (g529) & (g523)) + ((!g519) & (!g520) & (g521) & (g522) & (!g529) & (g523)) + ((!g519) & (g520) & (!g521) & (!g522) & (!g529) & (!g523)) + ((!g519) & (g520) & (!g521) & (!g522) & (g529) & (!g523)) + ((!g519) & (g520) & (!g521) & (g522) & (!g529) & (g523)) + ((!g519) & (g520) & (g521) & (!g522) & (!g529) & (g523)) + ((!g519) & (g520) & (g521) & (!g522) & (g529) & (!g523)) + ((!g519) & (g520) & (g521) & (!g522) & (g529) & (g523)) + ((!g519) & (g520) & (g521) & (g522) & (g529) & (!g523)) + ((!g519) & (g520) & (g521) & (g522) & (g529) & (g523)) + ((g519) & (!g520) & (!g521) & (!g522) & (!g529) & (!g523)) + ((g519) & (!g520) & (!g521) & (g522) & (!g529) & (!g523)) + ((g519) & (!g520) & (!g521) & (g522) & (!g529) & (g523)) + ((g519) & (!g520) & (!g521) & (g522) & (g529) & (!g523)) + ((g519) & (!g520) & (g521) & (!g522) & (!g529) & (!g523)) + ((g519) & (!g520) & (g521) & (!g522) & (g529) & (g523)) + ((g519) & (!g520) & (g521) & (g522) & (g529) & (!g523)) + ((g519) & (g520) & (!g521) & (!g522) & (!g529) & (!g523)) + ((g519) & (g520) & (!g521) & (g522) & (!g529) & (!g523)) + ((g519) & (g520) & (!g521) & (g522) & (g529) & (!g523)) + ((g519) & (g520) & (!g521) & (g522) & (g529) & (g523)) + ((g519) & (g520) & (g521) & (g522) & (!g529) & (g523)) + ((g519) & (g520) & (g521) & (g522) & (g529) & (g523)));
	assign g538 = (((!g534) & (!g535) & (!g536) & (!g537) & (!g524) & (!g530)) + ((!g534) & (!g535) & (!g536) & (!g537) & (g524) & (!g530)) + ((!g534) & (!g535) & (!g536) & (g537) & (!g524) & (!g530)) + ((!g534) & (!g535) & (!g536) & (g537) & (g524) & (!g530)) + ((!g534) & (!g535) & (!g536) & (g537) & (g524) & (g530)) + ((!g534) & (!g535) & (g536) & (!g537) & (!g524) & (!g530)) + ((!g534) & (!g535) & (g536) & (!g537) & (!g524) & (g530)) + ((!g534) & (!g535) & (g536) & (!g537) & (g524) & (!g530)) + ((!g534) & (!g535) & (g536) & (g537) & (!g524) & (!g530)) + ((!g534) & (!g535) & (g536) & (g537) & (!g524) & (g530)) + ((!g534) & (!g535) & (g536) & (g537) & (g524) & (!g530)) + ((!g534) & (!g535) & (g536) & (g537) & (g524) & (g530)) + ((!g534) & (g535) & (!g536) & (!g537) & (!g524) & (!g530)) + ((!g534) & (g535) & (!g536) & (g537) & (!g524) & (!g530)) + ((!g534) & (g535) & (!g536) & (g537) & (g524) & (g530)) + ((!g534) & (g535) & (g536) & (!g537) & (!g524) & (!g530)) + ((!g534) & (g535) & (g536) & (!g537) & (!g524) & (g530)) + ((!g534) & (g535) & (g536) & (g537) & (!g524) & (!g530)) + ((!g534) & (g535) & (g536) & (g537) & (!g524) & (g530)) + ((!g534) & (g535) & (g536) & (g537) & (g524) & (g530)) + ((g534) & (!g535) & (!g536) & (!g537) & (g524) & (!g530)) + ((g534) & (!g535) & (!g536) & (g537) & (g524) & (!g530)) + ((g534) & (!g535) & (!g536) & (g537) & (g524) & (g530)) + ((g534) & (!g535) & (g536) & (!g537) & (!g524) & (g530)) + ((g534) & (!g535) & (g536) & (!g537) & (g524) & (!g530)) + ((g534) & (!g535) & (g536) & (g537) & (!g524) & (g530)) + ((g534) & (!g535) & (g536) & (g537) & (g524) & (!g530)) + ((g534) & (!g535) & (g536) & (g537) & (g524) & (g530)) + ((g534) & (g535) & (!g536) & (g537) & (g524) & (g530)) + ((g534) & (g535) & (g536) & (!g537) & (!g524) & (g530)) + ((g534) & (g535) & (g536) & (g537) & (!g524) & (g530)) + ((g534) & (g535) & (g536) & (g537) & (g524) & (g530)));
	assign g540 = (((!sk[44]) & (g538) & (!g539)) + ((!sk[44]) & (g538) & (g539)) + ((sk[44]) & (!g538) & (g539)) + ((sk[44]) & (g538) & (!g539)));
	assign g541 = (((!g523) & (!g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((!g523) & (!g520) & (!g521) & (!g522) & (g529) & (g524)) + ((!g523) & (!g520) & (!g521) & (g522) & (!g529) & (g524)) + ((!g523) & (!g520) & (!g521) & (g522) & (g529) & (!g524)) + ((!g523) & (!g520) & (!g521) & (g522) & (g529) & (g524)) + ((!g523) & (!g520) & (g521) & (!g522) & (!g529) & (g524)) + ((!g523) & (!g520) & (g521) & (g522) & (!g529) & (!g524)) + ((!g523) & (!g520) & (g521) & (g522) & (g529) & (!g524)) + ((!g523) & (g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((!g523) & (g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((!g523) & (g520) & (!g521) & (g522) & (!g529) & (g524)) + ((!g523) & (g520) & (g521) & (!g522) & (!g529) & (!g524)) + ((!g523) & (g520) & (g521) & (!g522) & (!g529) & (g524)) + ((!g523) & (g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g523) & (g520) & (g521) & (!g522) & (g529) & (g524)) + ((g523) & (!g520) & (!g521) & (g522) & (!g529) & (g524)) + ((g523) & (!g520) & (!g521) & (g522) & (g529) & (g524)) + ((g523) & (g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((g523) & (g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((g523) & (g520) & (!g521) & (g522) & (g529) & (!g524)) + ((g523) & (g520) & (g521) & (g522) & (!g529) & (!g524)) + ((g523) & (g520) & (g521) & (g522) & (!g529) & (g524)));
	assign g542 = (((!g523) & (!g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((!g523) & (!g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((!g523) & (!g520) & (!g521) & (g522) & (g529) & (g524)) + ((!g523) & (!g520) & (g521) & (!g522) & (!g529) & (!g524)) + ((!g523) & (!g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g523) & (!g520) & (g521) & (g522) & (!g529) & (g524)) + ((!g523) & (g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((!g523) & (g520) & (!g521) & (!g522) & (g529) & (g524)) + ((!g523) & (g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((!g523) & (g520) & (!g521) & (g522) & (!g529) & (g524)) + ((!g523) & (g520) & (!g521) & (g522) & (g529) & (g524)) + ((!g523) & (g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g523) & (g520) & (g521) & (!g522) & (g529) & (g524)) + ((!g523) & (g520) & (g521) & (g522) & (g529) & (!g524)) + ((g523) & (!g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((g523) & (!g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((g523) & (!g520) & (!g521) & (!g522) & (g529) & (g524)) + ((g523) & (!g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((g523) & (!g520) & (!g521) & (g522) & (!g529) & (g524)) + ((g523) & (!g520) & (!g521) & (g522) & (g529) & (!g524)) + ((g523) & (!g520) & (g521) & (g522) & (!g529) & (!g524)) + ((g523) & (g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((g523) & (g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((g523) & (g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((g523) & (g520) & (!g521) & (g522) & (g529) & (!g524)) + ((g523) & (g520) & (!g521) & (g522) & (g529) & (g524)) + ((g523) & (g520) & (g521) & (!g522) & (!g529) & (!g524)) + ((g523) & (g520) & (g521) & (!g522) & (g529) & (!g524)) + ((g523) & (g520) & (g521) & (g522) & (!g529) & (g524)) + ((g523) & (g520) & (g521) & (g522) & (g529) & (g524)));
	assign g543 = (((!g523) & (!g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((!g523) & (!g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((!g523) & (!g520) & (!g521) & (g522) & (!g529) & (g524)) + ((!g523) & (!g520) & (g521) & (!g522) & (!g529) & (g524)) + ((!g523) & (!g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g523) & (!g520) & (g521) & (g522) & (!g529) & (g524)) + ((!g523) & (g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((!g523) & (g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((!g523) & (g520) & (!g521) & (g522) & (g529) & (!g524)) + ((!g523) & (g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g523) & (g520) & (g521) & (g522) & (!g529) & (!g524)) + ((!g523) & (g520) & (g521) & (g522) & (g529) & (!g524)) + ((g523) & (!g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((g523) & (!g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((g523) & (!g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((g523) & (!g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((g523) & (!g520) & (!g521) & (g522) & (!g529) & (g524)) + ((g523) & (!g520) & (!g521) & (g522) & (g529) & (!g524)) + ((g523) & (!g520) & (!g521) & (g522) & (g529) & (g524)) + ((g523) & (!g520) & (g521) & (!g522) & (!g529) & (g524)) + ((g523) & (!g520) & (g521) & (!g522) & (g529) & (!g524)) + ((g523) & (!g520) & (g521) & (g522) & (!g529) & (!g524)) + ((g523) & (!g520) & (g521) & (g522) & (g529) & (g524)) + ((g523) & (g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((g523) & (g520) & (!g521) & (!g522) & (g529) & (g524)) + ((g523) & (g520) & (g521) & (!g522) & (g529) & (g524)) + ((g523) & (g520) & (g521) & (g522) & (!g529) & (!g524)) + ((g523) & (g520) & (g521) & (g522) & (!g529) & (g524)) + ((g523) & (g520) & (g521) & (g522) & (g529) & (g524)));
	assign g544 = (((!g523) & (!g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((!g523) & (!g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((!g523) & (!g520) & (!g521) & (!g522) & (g529) & (g524)) + ((!g523) & (!g520) & (!g521) & (g522) & (!g529) & (g524)) + ((!g523) & (!g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g523) & (!g520) & (g521) & (g522) & (g529) & (g524)) + ((!g523) & (g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((!g523) & (g520) & (!g521) & (g522) & (!g529) & (g524)) + ((!g523) & (g520) & (!g521) & (g522) & (g529) & (g524)) + ((!g523) & (g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g523) & (g520) & (g521) & (!g522) & (g529) & (g524)) + ((!g523) & (g520) & (g521) & (g522) & (!g529) & (!g524)) + ((!g523) & (g520) & (g521) & (g522) & (!g529) & (g524)) + ((!g523) & (g520) & (g521) & (g522) & (g529) & (!g524)) + ((!g523) & (g520) & (g521) & (g522) & (g529) & (g524)) + ((g523) & (!g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((g523) & (!g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((g523) & (!g520) & (!g521) & (!g522) & (g529) & (g524)) + ((g523) & (!g520) & (!g521) & (g522) & (g529) & (g524)) + ((g523) & (!g520) & (g521) & (!g522) & (!g529) & (g524)) + ((g523) & (!g520) & (g521) & (!g522) & (g529) & (!g524)) + ((g523) & (!g520) & (g521) & (g522) & (g529) & (!g524)) + ((g523) & (g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((g523) & (g520) & (!g521) & (g522) & (!g529) & (g524)) + ((g523) & (g520) & (!g521) & (g522) & (g529) & (!g524)) + ((g523) & (g520) & (g521) & (!g522) & (g529) & (g524)) + ((g523) & (g520) & (g521) & (g522) & (!g529) & (!g524)));
	assign g545 = (((!g541) & (!g542) & (!g543) & (!g544) & (!g519) & (g530)) + ((!g541) & (!g542) & (!g543) & (!g544) & (g519) & (!g530)) + ((!g541) & (!g542) & (!g543) & (!g544) & (g519) & (g530)) + ((!g541) & (!g542) & (!g543) & (g544) & (!g519) & (g530)) + ((!g541) & (!g542) & (!g543) & (g544) & (g519) & (!g530)) + ((!g541) & (!g542) & (g543) & (!g544) & (g519) & (!g530)) + ((!g541) & (!g542) & (g543) & (!g544) & (g519) & (g530)) + ((!g541) & (!g542) & (g543) & (g544) & (g519) & (!g530)) + ((!g541) & (g542) & (!g543) & (!g544) & (!g519) & (g530)) + ((!g541) & (g542) & (!g543) & (!g544) & (g519) & (g530)) + ((!g541) & (g542) & (!g543) & (g544) & (!g519) & (g530)) + ((!g541) & (g542) & (g543) & (!g544) & (g519) & (g530)) + ((g541) & (!g542) & (!g543) & (!g544) & (!g519) & (!g530)) + ((g541) & (!g542) & (!g543) & (!g544) & (!g519) & (g530)) + ((g541) & (!g542) & (!g543) & (!g544) & (g519) & (!g530)) + ((g541) & (!g542) & (!g543) & (!g544) & (g519) & (g530)) + ((g541) & (!g542) & (!g543) & (g544) & (!g519) & (!g530)) + ((g541) & (!g542) & (!g543) & (g544) & (!g519) & (g530)) + ((g541) & (!g542) & (!g543) & (g544) & (g519) & (!g530)) + ((g541) & (!g542) & (g543) & (!g544) & (!g519) & (!g530)) + ((g541) & (!g542) & (g543) & (!g544) & (g519) & (!g530)) + ((g541) & (!g542) & (g543) & (!g544) & (g519) & (g530)) + ((g541) & (!g542) & (g543) & (g544) & (!g519) & (!g530)) + ((g541) & (!g542) & (g543) & (g544) & (g519) & (!g530)) + ((g541) & (g542) & (!g543) & (!g544) & (!g519) & (!g530)) + ((g541) & (g542) & (!g543) & (!g544) & (!g519) & (g530)) + ((g541) & (g542) & (!g543) & (!g544) & (g519) & (g530)) + ((g541) & (g542) & (!g543) & (g544) & (!g519) & (!g530)) + ((g541) & (g542) & (!g543) & (g544) & (!g519) & (g530)) + ((g541) & (g542) & (g543) & (!g544) & (!g519) & (!g530)) + ((g541) & (g542) & (g543) & (!g544) & (g519) & (g530)) + ((g541) & (g542) & (g543) & (g544) & (!g519) & (!g530)));
	assign g547 = (((!g545) & (sk[50]) & (g546)) + ((g545) & (!sk[50]) & (!g546)) + ((g545) & (!sk[50]) & (g546)) + ((g545) & (sk[50]) & (!g546)));
	assign g548 = (((!g519) & (!g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (g529) & (g524)) + ((!g519) & (!g520) & (g521) & (g522) & (!g529) & (!g524)) + ((!g519) & (!g520) & (g521) & (g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (g521) & (g522) & (g529) & (g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (g520) & (g521) & (!g522) & (!g529) & (!g524)) + ((!g519) & (g520) & (g521) & (g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((g519) & (!g520) & (g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (g521) & (!g522) & (!g529) & (g524)) + ((g519) & (!g520) & (g521) & (!g522) & (g529) & (!g524)) + ((g519) & (!g520) & (g521) & (g522) & (!g529) & (g524)) + ((g519) & (g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((g519) & (g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((g519) & (g520) & (!g521) & (g522) & (g529) & (!g524)) + ((g519) & (g520) & (g521) & (!g522) & (!g529) & (g524)) + ((g519) & (g520) & (g521) & (!g522) & (g529) & (g524)));
	assign g549 = (((!g519) & (!g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (!g521) & (!g522) & (g529) & (g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (g521) & (g522) & (!g529) & (!g524)) + ((!g519) & (!g520) & (g521) & (g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (g521) & (g522) & (g529) & (g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (g529) & (g524)) + ((!g519) & (g520) & (!g521) & (g522) & (g529) & (g524)) + ((!g519) & (g520) & (g521) & (!g522) & (!g529) & (!g524)) + ((!g519) & (g520) & (g521) & (!g522) & (!g529) & (g524)) + ((!g519) & (g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (g520) & (g521) & (g522) & (!g529) & (g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((g519) & (!g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (!g521) & (g522) & (!g529) & (g524)) + ((g519) & (!g520) & (!g521) & (g522) & (g529) & (g524)) + ((g519) & (!g520) & (g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (g521) & (!g522) & (!g529) & (g524)) + ((g519) & (!g520) & (g521) & (!g522) & (g529) & (g524)) + ((g519) & (!g520) & (g521) & (g522) & (!g529) & (g524)) + ((g519) & (g520) & (!g521) & (g522) & (!g529) & (g524)) + ((g519) & (g520) & (!g521) & (g522) & (g529) & (!g524)) + ((g519) & (g520) & (g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (g520) & (g521) & (g522) & (!g529) & (!g524)));
	assign g550 = (((!g519) & (!g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (!g521) & (!g522) & (g529) & (g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (g521) & (!g522) & (g529) & (g524)) + ((!g519) & (!g520) & (g521) & (g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (g521) & (g522) & (g529) & (g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (g529) & (g524)) + ((!g519) & (g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((!g519) & (g520) & (!g521) & (g522) & (!g529) & (g524)) + ((!g519) & (g520) & (g521) & (!g522) & (!g529) & (g524)) + ((!g519) & (g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (g520) & (g521) & (g522) & (g529) & (g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (g529) & (g524)) + ((g519) & (!g520) & (!g521) & (g522) & (g529) & (g524)) + ((g519) & (!g520) & (g521) & (g522) & (!g529) & (!g524)) + ((g519) & (g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((g519) & (g520) & (!g521) & (g522) & (g529) & (g524)) + ((g519) & (g520) & (g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (g520) & (g521) & (!g522) & (!g529) & (g524)) + ((g519) & (g520) & (g521) & (!g522) & (g529) & (g524)) + ((g519) & (g520) & (g521) & (g522) & (!g529) & (!g524)) + ((g519) & (g520) & (g521) & (g522) & (g529) & (g524)));
	assign g551 = (((!g519) & (!g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (!g521) & (g522) & (g529) & (g524)) + ((!g519) & (!g520) & (g521) & (g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (g521) & (g522) & (g529) & (g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (!g529) & (!g524)) + ((!g519) & (g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (g520) & (!g521) & (g522) & (!g529) & (!g524)) + ((!g519) & (g520) & (!g521) & (g522) & (!g529) & (g524)) + ((!g519) & (g520) & (!g521) & (g522) & (g529) & (!g524)) + ((!g519) & (g520) & (g521) & (!g522) & (!g529) & (!g524)) + ((!g519) & (g520) & (g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (g520) & (g521) & (!g522) & (g529) & (g524)) + ((g519) & (!g520) & (!g521) & (!g522) & (g529) & (g524)) + ((g519) & (!g520) & (!g521) & (g522) & (g529) & (!g524)) + ((g519) & (!g520) & (g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (g521) & (!g522) & (g529) & (!g524)) + ((g519) & (!g520) & (g521) & (!g522) & (g529) & (g524)) + ((g519) & (!g520) & (g521) & (g522) & (!g529) & (g524)) + ((g519) & (!g520) & (g521) & (g522) & (g529) & (!g524)) + ((g519) & (!g520) & (g521) & (g522) & (g529) & (g524)) + ((g519) & (g520) & (!g521) & (!g522) & (!g529) & (g524)) + ((g519) & (g520) & (!g521) & (!g522) & (g529) & (!g524)) + ((g519) & (g520) & (g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (g520) & (g521) & (!g522) & (!g529) & (g524)) + ((g519) & (g520) & (g521) & (g522) & (g529) & (g524)));
	assign g552 = (((!g548) & (!g549) & (!g550) & (!g551) & (!g530) & (g523)) + ((!g548) & (!g549) & (!g550) & (!g551) & (g530) & (!g523)) + ((!g548) & (!g549) & (!g550) & (!g551) & (g530) & (g523)) + ((!g548) & (!g549) & (!g550) & (g551) & (!g530) & (g523)) + ((!g548) & (!g549) & (!g550) & (g551) & (g530) & (!g523)) + ((!g548) & (!g549) & (g550) & (!g551) & (g530) & (!g523)) + ((!g548) & (!g549) & (g550) & (!g551) & (g530) & (g523)) + ((!g548) & (!g549) & (g550) & (g551) & (g530) & (!g523)) + ((!g548) & (g549) & (!g550) & (!g551) & (!g530) & (g523)) + ((!g548) & (g549) & (!g550) & (!g551) & (g530) & (g523)) + ((!g548) & (g549) & (!g550) & (g551) & (!g530) & (g523)) + ((!g548) & (g549) & (g550) & (!g551) & (g530) & (g523)) + ((g548) & (!g549) & (!g550) & (!g551) & (!g530) & (!g523)) + ((g548) & (!g549) & (!g550) & (!g551) & (!g530) & (g523)) + ((g548) & (!g549) & (!g550) & (!g551) & (g530) & (!g523)) + ((g548) & (!g549) & (!g550) & (!g551) & (g530) & (g523)) + ((g548) & (!g549) & (!g550) & (g551) & (!g530) & (!g523)) + ((g548) & (!g549) & (!g550) & (g551) & (!g530) & (g523)) + ((g548) & (!g549) & (!g550) & (g551) & (g530) & (!g523)) + ((g548) & (!g549) & (g550) & (!g551) & (!g530) & (!g523)) + ((g548) & (!g549) & (g550) & (!g551) & (g530) & (!g523)) + ((g548) & (!g549) & (g550) & (!g551) & (g530) & (g523)) + ((g548) & (!g549) & (g550) & (g551) & (!g530) & (!g523)) + ((g548) & (!g549) & (g550) & (g551) & (g530) & (!g523)) + ((g548) & (g549) & (!g550) & (!g551) & (!g530) & (!g523)) + ((g548) & (g549) & (!g550) & (!g551) & (!g530) & (g523)) + ((g548) & (g549) & (!g550) & (!g551) & (g530) & (g523)) + ((g548) & (g549) & (!g550) & (g551) & (!g530) & (!g523)) + ((g548) & (g549) & (!g550) & (g551) & (!g530) & (g523)) + ((g548) & (g549) & (g550) & (!g551) & (!g530) & (!g523)) + ((g548) & (g549) & (g550) & (!g551) & (g530) & (g523)) + ((g548) & (g549) & (g550) & (g551) & (!g530) & (!g523)));
	assign g554 = (((!sk[56]) & (g552) & (!g553)) + ((!sk[56]) & (g552) & (g553)) + ((sk[56]) & (!g552) & (g553)) + ((sk[56]) & (g552) & (!g553)));
	assign g555 = (((!g519) & (!g520) & (!g523) & (!g530) & (!g529) & (g524)) + ((!g519) & (!g520) & (g523) & (!g530) & (!g529) & (g524)) + ((!g519) & (!g520) & (g523) & (!g530) & (g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (!g530) & (g529) & (g524)) + ((!g519) & (!g520) & (g523) & (g530) & (!g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (g530) & (g529) & (!g524)) + ((!g519) & (g520) & (!g523) & (!g530) & (!g529) & (!g524)) + ((!g519) & (g520) & (!g523) & (!g530) & (!g529) & (g524)) + ((!g519) & (g520) & (!g523) & (g530) & (!g529) & (!g524)) + ((!g519) & (g520) & (!g523) & (g530) & (!g529) & (g524)) + ((!g519) & (g520) & (!g523) & (g530) & (g529) & (g524)) + ((!g519) & (g520) & (g523) & (g530) & (!g529) & (g524)) + ((!g519) & (g520) & (g523) & (g530) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g530) & (!g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g530) & (!g529) & (g524)) + ((g519) & (!g520) & (!g523) & (g530) & (!g529) & (g524)) + ((g519) & (!g520) & (g523) & (!g530) & (g529) & (!g524)) + ((g519) & (!g520) & (g523) & (g530) & (!g529) & (!g524)) + ((g519) & (!g520) & (g523) & (g530) & (!g529) & (g524)) + ((g519) & (!g520) & (g523) & (g530) & (g529) & (!g524)) + ((g519) & (g520) & (!g523) & (!g530) & (!g529) & (!g524)) + ((g519) & (g520) & (!g523) & (!g530) & (g529) & (!g524)) + ((g519) & (g520) & (!g523) & (g530) & (g529) & (!g524)) + ((g519) & (g520) & (g523) & (!g530) & (!g529) & (!g524)) + ((g519) & (g520) & (g523) & (!g530) & (!g529) & (g524)) + ((g519) & (g520) & (g523) & (g530) & (!g529) & (g524)));
	assign g556 = (((!g519) & (!g520) & (!g523) & (!g530) & (!g529) & (!g524)) + ((!g519) & (!g520) & (!g523) & (!g530) & (!g529) & (g524)) + ((!g519) & (!g520) & (!g523) & (!g530) & (g529) & (!g524)) + ((!g519) & (!g520) & (!g523) & (!g530) & (g529) & (g524)) + ((!g519) & (!g520) & (!g523) & (g530) & (!g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (!g530) & (!g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (!g530) & (g529) & (g524)) + ((!g519) & (!g520) & (g523) & (g530) & (!g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (g530) & (g529) & (g524)) + ((!g519) & (g520) & (!g523) & (!g530) & (!g529) & (g524)) + ((!g519) & (g520) & (!g523) & (g530) & (g529) & (!g524)) + ((!g519) & (g520) & (g523) & (!g530) & (!g529) & (!g524)) + ((!g519) & (g520) & (g523) & (!g530) & (!g529) & (g524)) + ((!g519) & (g520) & (g523) & (!g530) & (g529) & (!g524)) + ((!g519) & (g520) & (g523) & (!g530) & (g529) & (g524)) + ((!g519) & (g520) & (g523) & (g530) & (!g529) & (!g524)) + ((!g519) & (g520) & (g523) & (g530) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g530) & (!g529) & (g524)) + ((g519) & (!g520) & (!g523) & (!g530) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g530) & (g529) & (g524)) + ((g519) & (!g520) & (!g523) & (g530) & (!g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (g530) & (g529) & (g524)) + ((g519) & (!g520) & (g523) & (!g530) & (g529) & (!g524)) + ((g519) & (!g520) & (g523) & (!g530) & (g529) & (g524)) + ((g519) & (!g520) & (g523) & (g530) & (!g529) & (g524)) + ((g519) & (g520) & (!g523) & (!g530) & (g529) & (!g524)) + ((g519) & (g520) & (!g523) & (!g530) & (g529) & (g524)) + ((g519) & (g520) & (!g523) & (g530) & (!g529) & (!g524)) + ((g519) & (g520) & (!g523) & (g530) & (!g529) & (g524)) + ((g519) & (g520) & (g523) & (!g530) & (g529) & (!g524)) + ((g519) & (g520) & (g523) & (!g530) & (g529) & (g524)) + ((g519) & (g520) & (g523) & (g530) & (!g529) & (g524)));
	assign g557 = (((!g519) & (!g520) & (!g523) & (!g530) & (!g529) & (!g524)) + ((!g519) & (!g520) & (!g523) & (!g530) & (!g529) & (g524)) + ((!g519) & (!g520) & (g523) & (!g530) & (!g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (!g530) & (g529) & (g524)) + ((!g519) & (!g520) & (g523) & (g530) & (!g529) & (g524)) + ((!g519) & (g520) & (!g523) & (g530) & (!g529) & (!g524)) + ((!g519) & (g520) & (!g523) & (g530) & (g529) & (!g524)) + ((!g519) & (g520) & (!g523) & (g530) & (g529) & (g524)) + ((!g519) & (g520) & (g523) & (!g530) & (!g529) & (!g524)) + ((!g519) & (g520) & (g523) & (!g530) & (g529) & (!g524)) + ((!g519) & (g520) & (g523) & (!g530) & (g529) & (g524)) + ((!g519) & (g520) & (g523) & (g530) & (!g529) & (!g524)) + ((!g519) & (g520) & (g523) & (g530) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g530) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g530) & (g529) & (g524)) + ((g519) & (!g520) & (!g523) & (g530) & (!g529) & (g524)) + ((g519) & (!g520) & (!g523) & (g530) & (g529) & (g524)) + ((g519) & (!g520) & (g523) & (!g530) & (!g529) & (!g524)) + ((g519) & (!g520) & (g523) & (!g530) & (!g529) & (g524)) + ((g519) & (!g520) & (g523) & (!g530) & (g529) & (g524)) + ((g519) & (!g520) & (g523) & (g530) & (!g529) & (!g524)) + ((g519) & (!g520) & (g523) & (g530) & (!g529) & (g524)) + ((g519) & (!g520) & (g523) & (g530) & (g529) & (!g524)) + ((g519) & (!g520) & (g523) & (g530) & (g529) & (g524)) + ((g519) & (g520) & (!g523) & (!g530) & (!g529) & (g524)) + ((g519) & (g520) & (!g523) & (g530) & (!g529) & (!g524)) + ((g519) & (g520) & (!g523) & (g530) & (g529) & (!g524)) + ((g519) & (g520) & (g523) & (!g530) & (!g529) & (!g524)) + ((g519) & (g520) & (g523) & (!g530) & (!g529) & (g524)) + ((g519) & (g520) & (g523) & (!g530) & (g529) & (!g524)) + ((g519) & (g520) & (g523) & (g530) & (!g529) & (!g524)) + ((g519) & (g520) & (g523) & (g530) & (g529) & (!g524)));
	assign g558 = (((!g519) & (!g520) & (!g523) & (!g530) & (g529) & (g524)) + ((!g519) & (!g520) & (!g523) & (g530) & (!g529) & (!g524)) + ((!g519) & (!g520) & (!g523) & (g530) & (g529) & (g524)) + ((!g519) & (!g520) & (g523) & (!g530) & (!g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (!g530) & (g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (g530) & (!g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (g530) & (!g529) & (g524)) + ((!g519) & (!g520) & (g523) & (g530) & (g529) & (!g524)) + ((!g519) & (g520) & (!g523) & (!g530) & (!g529) & (!g524)) + ((!g519) & (g520) & (!g523) & (g530) & (!g529) & (g524)) + ((!g519) & (g520) & (!g523) & (g530) & (g529) & (!g524)) + ((!g519) & (g520) & (!g523) & (g530) & (g529) & (g524)) + ((!g519) & (g520) & (g523) & (!g530) & (!g529) & (!g524)) + ((!g519) & (g520) & (g523) & (g530) & (!g529) & (!g524)) + ((!g519) & (g520) & (g523) & (g530) & (!g529) & (g524)) + ((g519) & (!g520) & (!g523) & (!g530) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g530) & (g529) & (g524)) + ((g519) & (!g520) & (g523) & (!g530) & (!g529) & (!g524)) + ((g519) & (!g520) & (g523) & (!g530) & (g529) & (!g524)) + ((g519) & (!g520) & (g523) & (g530) & (g529) & (!g524)) + ((g519) & (g520) & (!g523) & (!g530) & (g529) & (!g524)) + ((g519) & (g520) & (!g523) & (g530) & (g529) & (g524)) + ((g519) & (g520) & (g523) & (!g530) & (!g529) & (!g524)) + ((g519) & (g520) & (g523) & (!g530) & (!g529) & (g524)) + ((g519) & (g520) & (g523) & (!g530) & (g529) & (!g524)) + ((g519) & (g520) & (g523) & (g530) & (!g529) & (!g524)));
	assign g559 = (((!g555) & (!g556) & (!g557) & (!g558) & (g521) & (g522)) + ((!g555) & (!g556) & (g557) & (!g558) & (!g521) & (g522)) + ((!g555) & (!g556) & (g557) & (!g558) & (g521) & (g522)) + ((!g555) & (!g556) & (g557) & (g558) & (!g521) & (g522)) + ((!g555) & (g556) & (!g557) & (!g558) & (g521) & (!g522)) + ((!g555) & (g556) & (!g557) & (!g558) & (g521) & (g522)) + ((!g555) & (g556) & (!g557) & (g558) & (g521) & (!g522)) + ((!g555) & (g556) & (g557) & (!g558) & (!g521) & (g522)) + ((!g555) & (g556) & (g557) & (!g558) & (g521) & (!g522)) + ((!g555) & (g556) & (g557) & (!g558) & (g521) & (g522)) + ((!g555) & (g556) & (g557) & (g558) & (!g521) & (g522)) + ((!g555) & (g556) & (g557) & (g558) & (g521) & (!g522)) + ((g555) & (!g556) & (!g557) & (!g558) & (!g521) & (!g522)) + ((g555) & (!g556) & (!g557) & (!g558) & (g521) & (g522)) + ((g555) & (!g556) & (!g557) & (g558) & (!g521) & (!g522)) + ((g555) & (!g556) & (g557) & (!g558) & (!g521) & (!g522)) + ((g555) & (!g556) & (g557) & (!g558) & (!g521) & (g522)) + ((g555) & (!g556) & (g557) & (!g558) & (g521) & (g522)) + ((g555) & (!g556) & (g557) & (g558) & (!g521) & (!g522)) + ((g555) & (!g556) & (g557) & (g558) & (!g521) & (g522)) + ((g555) & (g556) & (!g557) & (!g558) & (!g521) & (!g522)) + ((g555) & (g556) & (!g557) & (!g558) & (g521) & (!g522)) + ((g555) & (g556) & (!g557) & (!g558) & (g521) & (g522)) + ((g555) & (g556) & (!g557) & (g558) & (!g521) & (!g522)) + ((g555) & (g556) & (!g557) & (g558) & (g521) & (!g522)) + ((g555) & (g556) & (g557) & (!g558) & (!g521) & (!g522)) + ((g555) & (g556) & (g557) & (!g558) & (!g521) & (g522)) + ((g555) & (g556) & (g557) & (!g558) & (g521) & (!g522)) + ((g555) & (g556) & (g557) & (!g558) & (g521) & (g522)) + ((g555) & (g556) & (g557) & (g558) & (!g521) & (!g522)) + ((g555) & (g556) & (g557) & (g558) & (!g521) & (g522)) + ((g555) & (g556) & (g557) & (g558) & (g521) & (!g522)));
	assign g561 = (((!sk[62]) & (g559) & (!g560)) + ((!sk[62]) & (g559) & (g560)) + ((sk[62]) & (!g559) & (g560)) + ((sk[62]) & (g559) & (!g560)));
	assign g562 = (((!g519) & (!g520) & (!g523) & (!g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (!g523) & (!g522) & (g529) & (g524)) + ((!g519) & (!g520) & (!g523) & (g522) & (g529) & (g524)) + ((!g519) & (!g520) & (g523) & (!g522) & (!g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (!g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (g523) & (!g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (!g522) & (g529) & (g524)) + ((!g519) & (!g520) & (g523) & (g522) & (!g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (g522) & (!g529) & (g524)) + ((!g519) & (g520) & (!g523) & (!g522) & (!g529) & (g524)) + ((!g519) & (g520) & (!g523) & (!g522) & (g529) & (!g524)) + ((!g519) & (g520) & (!g523) & (g522) & (g529) & (g524)) + ((!g519) & (g520) & (g523) & (!g522) & (g529) & (!g524)) + ((!g519) & (g520) & (g523) & (!g522) & (g529) & (g524)) + ((!g519) & (g520) & (g523) & (g522) & (!g529) & (!g524)) + ((!g519) & (g520) & (g523) & (g522) & (!g529) & (g524)) + ((!g519) & (g520) & (g523) & (g522) & (g529) & (g524)) + ((g519) & (!g520) & (!g523) & (!g522) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g522) & (g529) & (g524)) + ((g519) & (!g520) & (!g523) & (g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (g522) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (g522) & (g529) & (g524)) + ((g519) & (!g520) & (g523) & (!g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (g523) & (!g522) & (g529) & (!g524)) + ((g519) & (!g520) & (g523) & (g522) & (g529) & (!g524)) + ((g519) & (g520) & (!g523) & (!g522) & (g529) & (g524)) + ((g519) & (g520) & (g523) & (!g522) & (!g529) & (!g524)) + ((g519) & (g520) & (g523) & (!g522) & (g529) & (g524)));
	assign g563 = (((!g519) & (!g520) & (!g523) & (!g522) & (!g529) & (!g524)) + ((!g519) & (!g520) & (!g523) & (g522) & (!g529) & (!g524)) + ((!g519) & (!g520) & (!g523) & (g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (!g523) & (g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (!g522) & (g529) & (g524)) + ((!g519) & (!g520) & (g523) & (g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (g523) & (g522) & (g529) & (g524)) + ((!g519) & (g520) & (!g523) & (!g522) & (!g529) & (!g524)) + ((!g519) & (g520) & (!g523) & (!g522) & (g529) & (!g524)) + ((!g519) & (g520) & (g523) & (!g522) & (!g529) & (g524)) + ((!g519) & (g520) & (g523) & (!g522) & (g529) & (g524)) + ((!g519) & (g520) & (g523) & (g522) & (!g529) & (g524)) + ((!g519) & (g520) & (g523) & (g522) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g522) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g522) & (g529) & (g524)) + ((g519) & (!g520) & (!g523) & (g522) & (!g529) & (g524)) + ((g519) & (!g520) & (!g523) & (g522) & (g529) & (g524)) + ((g519) & (!g520) & (g523) & (g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (g523) & (g522) & (!g529) & (g524)) + ((g519) & (!g520) & (g523) & (g522) & (g529) & (g524)) + ((g519) & (g520) & (!g523) & (!g522) & (!g529) & (g524)) + ((g519) & (g520) & (!g523) & (!g522) & (g529) & (!g524)) + ((g519) & (g520) & (!g523) & (g522) & (g529) & (!g524)) + ((g519) & (g520) & (g523) & (!g522) & (!g529) & (g524)) + ((g519) & (g520) & (g523) & (!g522) & (g529) & (g524)) + ((g519) & (g520) & (g523) & (g522) & (!g529) & (!g524)) + ((g519) & (g520) & (g523) & (g522) & (g529) & (g524)));
	assign g564 = (((!g519) & (!g520) & (!g523) & (!g522) & (g529) & (g524)) + ((!g519) & (!g520) & (!g523) & (g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (!g522) & (!g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (!g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (g523) & (!g522) & (g529) & (g524)) + ((!g519) & (!g520) & (g523) & (g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (g523) & (g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (g523) & (g522) & (g529) & (g524)) + ((!g519) & (g520) & (!g523) & (!g522) & (g529) & (!g524)) + ((!g519) & (g520) & (!g523) & (!g522) & (g529) & (g524)) + ((!g519) & (g520) & (g523) & (!g522) & (!g529) & (!g524)) + ((!g519) & (g520) & (g523) & (g522) & (!g529) & (g524)) + ((!g519) & (g520) & (g523) & (g522) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g522) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (!g522) & (g529) & (g524)) + ((g519) & (!g520) & (!g523) & (g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (g522) & (!g529) & (g524)) + ((g519) & (!g520) & (g523) & (!g522) & (!g529) & (g524)) + ((g519) & (!g520) & (g523) & (!g522) & (g529) & (g524)) + ((g519) & (!g520) & (g523) & (g522) & (g529) & (!g524)) + ((g519) & (g520) & (!g523) & (!g522) & (!g529) & (!g524)) + ((g519) & (g520) & (!g523) & (!g522) & (!g529) & (g524)) + ((g519) & (g520) & (!g523) & (!g522) & (g529) & (g524)) + ((g519) & (g520) & (!g523) & (g522) & (!g529) & (g524)) + ((g519) & (g520) & (!g523) & (g522) & (g529) & (!g524)) + ((g519) & (g520) & (g523) & (!g522) & (!g529) & (g524)) + ((g519) & (g520) & (g523) & (!g522) & (g529) & (!g524)) + ((g519) & (g520) & (g523) & (g522) & (!g529) & (!g524)) + ((g519) & (g520) & (g523) & (g522) & (g529) & (!g524)) + ((g519) & (g520) & (g523) & (g522) & (g529) & (g524)));
	assign g565 = (((!g519) & (!g520) & (!g523) & (!g522) & (g529) & (!g524)) + ((!g519) & (!g520) & (!g523) & (g522) & (!g529) & (!g524)) + ((!g519) & (!g520) & (!g523) & (g522) & (g529) & (g524)) + ((!g519) & (!g520) & (g523) & (!g522) & (!g529) & (g524)) + ((!g519) & (!g520) & (g523) & (!g522) & (g529) & (g524)) + ((!g519) & (!g520) & (g523) & (g522) & (g529) & (g524)) + ((!g519) & (g520) & (!g523) & (!g522) & (!g529) & (g524)) + ((!g519) & (g520) & (!g523) & (g522) & (!g529) & (g524)) + ((!g519) & (g520) & (!g523) & (g522) & (g529) & (g524)) + ((!g519) & (g520) & (g523) & (!g522) & (!g529) & (!g524)) + ((!g519) & (g520) & (g523) & (!g522) & (g529) & (!g524)) + ((!g519) & (g520) & (g523) & (g522) & (!g529) & (g524)) + ((!g519) & (g520) & (g523) & (g522) & (g529) & (g524)) + ((g519) & (!g520) & (!g523) & (!g522) & (g529) & (!g524)) + ((g519) & (!g520) & (!g523) & (g522) & (g529) & (g524)) + ((g519) & (!g520) & (g523) & (!g522) & (!g529) & (!g524)) + ((g519) & (!g520) & (g523) & (!g522) & (g529) & (g524)) + ((g519) & (!g520) & (g523) & (g522) & (!g529) & (!g524)) + ((g519) & (g520) & (!g523) & (!g522) & (g529) & (g524)) + ((g519) & (g520) & (!g523) & (g522) & (!g529) & (!g524)) + ((g519) & (g520) & (!g523) & (g522) & (!g529) & (g524)) + ((g519) & (g520) & (g523) & (!g522) & (g529) & (g524)));
	assign g566 = (((!g562) & (!g563) & (!g564) & (!g565) & (!g530) & (!g521)) + ((!g562) & (!g563) & (!g564) & (!g565) & (!g530) & (g521)) + ((!g562) & (!g563) & (!g564) & (!g565) & (g530) & (!g521)) + ((!g562) & (!g563) & (!g564) & (g565) & (!g530) & (!g521)) + ((!g562) & (!g563) & (!g564) & (g565) & (!g530) & (g521)) + ((!g562) & (!g563) & (!g564) & (g565) & (g530) & (!g521)) + ((!g562) & (!g563) & (!g564) & (g565) & (g530) & (g521)) + ((!g562) & (!g563) & (g564) & (!g565) & (!g530) & (!g521)) + ((!g562) & (!g563) & (g564) & (!g565) & (g530) & (!g521)) + ((!g562) & (!g563) & (g564) & (g565) & (!g530) & (!g521)) + ((!g562) & (!g563) & (g564) & (g565) & (g530) & (!g521)) + ((!g562) & (!g563) & (g564) & (g565) & (g530) & (g521)) + ((!g562) & (g563) & (!g564) & (!g565) & (!g530) & (!g521)) + ((!g562) & (g563) & (!g564) & (!g565) & (!g530) & (g521)) + ((!g562) & (g563) & (!g564) & (g565) & (!g530) & (!g521)) + ((!g562) & (g563) & (!g564) & (g565) & (!g530) & (g521)) + ((!g562) & (g563) & (!g564) & (g565) & (g530) & (g521)) + ((!g562) & (g563) & (g564) & (!g565) & (!g530) & (!g521)) + ((!g562) & (g563) & (g564) & (g565) & (!g530) & (!g521)) + ((!g562) & (g563) & (g564) & (g565) & (g530) & (g521)) + ((g562) & (!g563) & (!g564) & (!g565) & (!g530) & (g521)) + ((g562) & (!g563) & (!g564) & (!g565) & (g530) & (!g521)) + ((g562) & (!g563) & (!g564) & (g565) & (!g530) & (g521)) + ((g562) & (!g563) & (!g564) & (g565) & (g530) & (!g521)) + ((g562) & (!g563) & (!g564) & (g565) & (g530) & (g521)) + ((g562) & (!g563) & (g564) & (!g565) & (g530) & (!g521)) + ((g562) & (!g563) & (g564) & (g565) & (g530) & (!g521)) + ((g562) & (!g563) & (g564) & (g565) & (g530) & (g521)) + ((g562) & (g563) & (!g564) & (!g565) & (!g530) & (g521)) + ((g562) & (g563) & (!g564) & (g565) & (!g530) & (g521)) + ((g562) & (g563) & (!g564) & (g565) & (g530) & (g521)) + ((g562) & (g563) & (g564) & (g565) & (g530) & (g521)));
	assign g568 = (((!sk[68]) & (g566) & (!g567)) + ((!sk[68]) & (g566) & (g567)) + ((sk[68]) & (!g566) & (g567)) + ((sk[68]) & (g566) & (!g567)));
	assign g569 = (((!g519) & (!g530) & (!g521) & (!g522) & (!g529) & (g524)) + ((!g519) & (!g530) & (!g521) & (!g522) & (g529) & (g524)) + ((!g519) & (!g530) & (!g521) & (g522) & (!g529) & (!g524)) + ((!g519) & (!g530) & (!g521) & (g522) & (!g529) & (g524)) + ((!g519) & (!g530) & (!g521) & (g522) & (g529) & (!g524)) + ((!g519) & (!g530) & (!g521) & (g522) & (g529) & (g524)) + ((!g519) & (!g530) & (g521) & (!g522) & (!g529) & (g524)) + ((!g519) & (!g530) & (g521) & (!g522) & (g529) & (g524)) + ((!g519) & (!g530) & (g521) & (g522) & (g529) & (!g524)) + ((!g519) & (g530) & (g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (g530) & (g521) & (!g522) & (g529) & (g524)) + ((!g519) & (g530) & (g521) & (g522) & (!g529) & (g524)) + ((g519) & (!g530) & (!g521) & (!g522) & (g529) & (!g524)) + ((g519) & (!g530) & (!g521) & (g522) & (!g529) & (!g524)) + ((g519) & (!g530) & (!g521) & (g522) & (!g529) & (g524)) + ((g519) & (!g530) & (!g521) & (g522) & (g529) & (g524)) + ((g519) & (!g530) & (g521) & (!g522) & (!g529) & (g524)) + ((g519) & (!g530) & (g521) & (!g522) & (g529) & (g524)) + ((g519) & (!g530) & (g521) & (g522) & (g529) & (!g524)) + ((g519) & (!g530) & (g521) & (g522) & (g529) & (g524)) + ((g519) & (g530) & (!g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (g530) & (!g521) & (!g522) & (!g529) & (g524)) + ((g519) & (g530) & (!g521) & (!g522) & (g529) & (!g524)) + ((g519) & (g530) & (!g521) & (g522) & (!g529) & (!g524)) + ((g519) & (g530) & (g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (g530) & (g521) & (!g522) & (!g529) & (g524)) + ((g519) & (g530) & (g521) & (!g522) & (g529) & (!g524)) + ((g519) & (g530) & (g521) & (g522) & (!g529) & (g524)));
	assign g570 = (((!g519) & (!g530) & (!g521) & (!g522) & (!g529) & (!g524)) + ((!g519) & (!g530) & (!g521) & (g522) & (g529) & (g524)) + ((!g519) & (!g530) & (g521) & (!g522) & (!g529) & (!g524)) + ((!g519) & (!g530) & (g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (!g530) & (g521) & (!g522) & (g529) & (g524)) + ((!g519) & (!g530) & (g521) & (g522) & (!g529) & (!g524)) + ((!g519) & (!g530) & (g521) & (g522) & (g529) & (g524)) + ((!g519) & (g530) & (!g521) & (!g522) & (!g529) & (!g524)) + ((!g519) & (g530) & (!g521) & (!g522) & (g529) & (g524)) + ((!g519) & (g530) & (!g521) & (g522) & (!g529) & (g524)) + ((!g519) & (g530) & (g521) & (!g522) & (!g529) & (!g524)) + ((!g519) & (g530) & (g521) & (!g522) & (g529) & (g524)) + ((!g519) & (g530) & (g521) & (g522) & (g529) & (!g524)) + ((!g519) & (g530) & (g521) & (g522) & (g529) & (g524)) + ((g519) & (!g530) & (!g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (!g530) & (!g521) & (!g522) & (g529) & (g524)) + ((g519) & (!g530) & (!g521) & (g522) & (!g529) & (!g524)) + ((g519) & (!g530) & (!g521) & (g522) & (g529) & (g524)) + ((g519) & (!g530) & (g521) & (!g522) & (g529) & (g524)) + ((g519) & (!g530) & (g521) & (g522) & (!g529) & (g524)) + ((g519) & (g530) & (!g521) & (!g522) & (g529) & (!g524)) + ((g519) & (g530) & (!g521) & (!g522) & (g529) & (g524)) + ((g519) & (g530) & (!g521) & (g522) & (!g529) & (g524)) + ((g519) & (g530) & (!g521) & (g522) & (g529) & (!g524)) + ((g519) & (g530) & (!g521) & (g522) & (g529) & (g524)) + ((g519) & (g530) & (g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (g530) & (g521) & (!g522) & (g529) & (!g524)) + ((g519) & (g530) & (g521) & (g522) & (!g529) & (!g524)));
	assign g571 = (((!g519) & (!g530) & (!g521) & (!g522) & (!g529) & (g524)) + ((!g519) & (!g530) & (!g521) & (!g522) & (g529) & (g524)) + ((!g519) & (!g530) & (!g521) & (g522) & (g529) & (!g524)) + ((!g519) & (!g530) & (!g521) & (g522) & (g529) & (g524)) + ((!g519) & (!g530) & (g521) & (!g522) & (g529) & (g524)) + ((!g519) & (!g530) & (g521) & (g522) & (!g529) & (!g524)) + ((!g519) & (!g530) & (g521) & (g522) & (!g529) & (g524)) + ((!g519) & (!g530) & (g521) & (g522) & (g529) & (g524)) + ((!g519) & (g530) & (!g521) & (!g522) & (!g529) & (!g524)) + ((!g519) & (g530) & (!g521) & (!g522) & (!g529) & (g524)) + ((!g519) & (g530) & (!g521) & (!g522) & (g529) & (g524)) + ((!g519) & (g530) & (!g521) & (g522) & (!g529) & (g524)) + ((!g519) & (g530) & (!g521) & (g522) & (g529) & (!g524)) + ((!g519) & (g530) & (g521) & (!g522) & (!g529) & (g524)) + ((!g519) & (g530) & (g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (g530) & (g521) & (g522) & (!g529) & (!g524)) + ((!g519) & (g530) & (g521) & (g522) & (g529) & (!g524)) + ((!g519) & (g530) & (g521) & (g522) & (g529) & (g524)) + ((g519) & (!g530) & (!g521) & (!g522) & (!g529) & (g524)) + ((g519) & (!g530) & (!g521) & (g522) & (!g529) & (!g524)) + ((g519) & (!g530) & (!g521) & (g522) & (g529) & (!g524)) + ((g519) & (!g530) & (g521) & (!g522) & (g529) & (g524)) + ((g519) & (!g530) & (g521) & (g522) & (!g529) & (g524)) + ((g519) & (g530) & (!g521) & (!g522) & (!g529) & (g524)) + ((g519) & (g530) & (!g521) & (g522) & (!g529) & (!g524)) + ((g519) & (g530) & (!g521) & (g522) & (g529) & (!g524)) + ((g519) & (g530) & (g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (g530) & (g521) & (!g522) & (g529) & (!g524)) + ((g519) & (g530) & (g521) & (!g522) & (g529) & (g524)) + ((g519) & (g530) & (g521) & (g522) & (g529) & (g524)));
	assign g572 = (((!g519) & (!g530) & (!g521) & (!g522) & (g529) & (g524)) + ((!g519) & (!g530) & (!g521) & (g522) & (!g529) & (!g524)) + ((!g519) & (!g530) & (!g521) & (g522) & (g529) & (g524)) + ((!g519) & (!g530) & (g521) & (!g522) & (!g529) & (!g524)) + ((!g519) & (!g530) & (g521) & (g522) & (g529) & (!g524)) + ((!g519) & (!g530) & (g521) & (g522) & (g529) & (g524)) + ((!g519) & (g530) & (!g521) & (g522) & (!g529) & (!g524)) + ((!g519) & (g530) & (!g521) & (g522) & (g529) & (!g524)) + ((!g519) & (g530) & (g521) & (!g522) & (g529) & (!g524)) + ((!g519) & (g530) & (g521) & (!g522) & (g529) & (g524)) + ((g519) & (!g530) & (!g521) & (!g522) & (!g529) & (g524)) + ((g519) & (!g530) & (!g521) & (!g522) & (g529) & (!g524)) + ((g519) & (!g530) & (!g521) & (g522) & (!g529) & (g524)) + ((g519) & (!g530) & (g521) & (!g522) & (g529) & (!g524)) + ((g519) & (!g530) & (g521) & (!g522) & (g529) & (g524)) + ((g519) & (!g530) & (g521) & (g522) & (g529) & (!g524)) + ((g519) & (!g530) & (g521) & (g522) & (g529) & (g524)) + ((g519) & (g530) & (!g521) & (!g522) & (g529) & (!g524)) + ((g519) & (g530) & (!g521) & (g522) & (!g529) & (g524)) + ((g519) & (g530) & (g521) & (!g522) & (!g529) & (!g524)) + ((g519) & (g530) & (g521) & (!g522) & (g529) & (g524)) + ((g519) & (g530) & (g521) & (g522) & (!g529) & (g524)));
	assign g573 = (((!g569) & (!g570) & (!g571) & (!g572) & (!g523) & (!g520)) + ((!g569) & (!g570) & (!g571) & (!g572) & (!g523) & (g520)) + ((!g569) & (!g570) & (!g571) & (!g572) & (g523) & (!g520)) + ((!g569) & (!g570) & (!g571) & (g572) & (!g523) & (!g520)) + ((!g569) & (!g570) & (!g571) & (g572) & (!g523) & (g520)) + ((!g569) & (!g570) & (!g571) & (g572) & (g523) & (!g520)) + ((!g569) & (!g570) & (!g571) & (g572) & (g523) & (g520)) + ((!g569) & (!g570) & (g571) & (!g572) & (!g523) & (!g520)) + ((!g569) & (!g570) & (g571) & (!g572) & (g523) & (!g520)) + ((!g569) & (!g570) & (g571) & (g572) & (!g523) & (!g520)) + ((!g569) & (!g570) & (g571) & (g572) & (g523) & (!g520)) + ((!g569) & (!g570) & (g571) & (g572) & (g523) & (g520)) + ((!g569) & (g570) & (!g571) & (!g572) & (!g523) & (!g520)) + ((!g569) & (g570) & (!g571) & (!g572) & (!g523) & (g520)) + ((!g569) & (g570) & (!g571) & (g572) & (!g523) & (!g520)) + ((!g569) & (g570) & (!g571) & (g572) & (!g523) & (g520)) + ((!g569) & (g570) & (!g571) & (g572) & (g523) & (g520)) + ((!g569) & (g570) & (g571) & (!g572) & (!g523) & (!g520)) + ((!g569) & (g570) & (g571) & (g572) & (!g523) & (!g520)) + ((!g569) & (g570) & (g571) & (g572) & (g523) & (g520)) + ((g569) & (!g570) & (!g571) & (!g572) & (!g523) & (g520)) + ((g569) & (!g570) & (!g571) & (!g572) & (g523) & (!g520)) + ((g569) & (!g570) & (!g571) & (g572) & (!g523) & (g520)) + ((g569) & (!g570) & (!g571) & (g572) & (g523) & (!g520)) + ((g569) & (!g570) & (!g571) & (g572) & (g523) & (g520)) + ((g569) & (!g570) & (g571) & (!g572) & (g523) & (!g520)) + ((g569) & (!g570) & (g571) & (g572) & (g523) & (!g520)) + ((g569) & (!g570) & (g571) & (g572) & (g523) & (g520)) + ((g569) & (g570) & (!g571) & (!g572) & (!g523) & (g520)) + ((g569) & (g570) & (!g571) & (g572) & (!g523) & (g520)) + ((g569) & (g570) & (!g571) & (g572) & (g523) & (g520)) + ((g569) & (g570) & (g571) & (g572) & (g523) & (g520)));
	assign g575 = (((!sk[74]) & (g573) & (!g574)) + ((!sk[74]) & (g573) & (g574)) + ((sk[74]) & (!g573) & (g574)) + ((sk[74]) & (g573) & (!g574)));
	assign g576 = (((!g523) & (!g520) & (!g521) & (!g522) & (!g529) & (g530)) + ((!g523) & (!g520) & (!g521) & (!g522) & (g529) & (!g530)) + ((!g523) & (!g520) & (!g521) & (g522) & (!g529) & (g530)) + ((!g523) & (!g520) & (!g521) & (g522) & (g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (!g522) & (!g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (!g522) & (g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (g522) & (!g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (g522) & (g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (g522) & (g529) & (g530)) + ((!g523) & (g520) & (!g521) & (!g522) & (g529) & (!g530)) + ((!g523) & (g520) & (!g521) & (g522) & (g529) & (!g530)) + ((!g523) & (g520) & (!g521) & (g522) & (g529) & (g530)) + ((!g523) & (g520) & (g521) & (!g522) & (g529) & (g530)) + ((!g523) & (g520) & (g521) & (g522) & (!g529) & (!g530)) + ((g523) & (!g520) & (!g521) & (!g522) & (!g529) & (g530)) + ((g523) & (!g520) & (!g521) & (g522) & (!g529) & (g530)) + ((g523) & (!g520) & (g521) & (g522) & (g529) & (g530)) + ((g523) & (g520) & (!g521) & (!g522) & (g529) & (g530)) + ((g523) & (g520) & (!g521) & (g522) & (!g529) & (!g530)) + ((g523) & (g520) & (!g521) & (g522) & (g529) & (!g530)) + ((g523) & (g520) & (g521) & (!g522) & (!g529) & (g530)) + ((g523) & (g520) & (g521) & (!g522) & (g529) & (!g530)) + ((g523) & (g520) & (g521) & (!g522) & (g529) & (g530)) + ((g523) & (g520) & (g521) & (g522) & (!g529) & (g530)));
	assign g577 = (((!g523) & (!g520) & (!g521) & (!g522) & (!g529) & (!g530)) + ((!g523) & (!g520) & (!g521) & (!g522) & (!g529) & (g530)) + ((!g523) & (!g520) & (!g521) & (g522) & (!g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (!g522) & (!g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (!g522) & (g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (!g522) & (g529) & (g530)) + ((!g523) & (!g520) & (g521) & (g522) & (!g529) & (g530)) + ((!g523) & (!g520) & (g521) & (g522) & (g529) & (g530)) + ((!g523) & (g520) & (!g521) & (!g522) & (!g529) & (!g530)) + ((!g523) & (g520) & (!g521) & (!g522) & (g529) & (!g530)) + ((!g523) & (g520) & (!g521) & (g522) & (!g529) & (!g530)) + ((!g523) & (g520) & (!g521) & (g522) & (!g529) & (g530)) + ((!g523) & (g520) & (!g521) & (g522) & (g529) & (g530)) + ((!g523) & (g520) & (g521) & (!g522) & (!g529) & (g530)) + ((!g523) & (g520) & (g521) & (g522) & (!g529) & (!g530)) + ((!g523) & (g520) & (g521) & (g522) & (!g529) & (g530)) + ((g523) & (!g520) & (!g521) & (!g522) & (!g529) & (g530)) + ((g523) & (!g520) & (!g521) & (!g522) & (g529) & (g530)) + ((g523) & (!g520) & (!g521) & (g522) & (!g529) & (!g530)) + ((g523) & (!g520) & (!g521) & (g522) & (g529) & (g530)) + ((g523) & (!g520) & (g521) & (!g522) & (!g529) & (!g530)) + ((g523) & (!g520) & (g521) & (!g522) & (g529) & (g530)) + ((g523) & (!g520) & (g521) & (g522) & (g529) & (!g530)) + ((g523) & (g520) & (!g521) & (!g522) & (!g529) & (!g530)) + ((g523) & (g520) & (!g521) & (!g522) & (!g529) & (g530)) + ((g523) & (g520) & (!g521) & (!g522) & (g529) & (g530)) + ((g523) & (g520) & (!g521) & (g522) & (!g529) & (g530)) + ((g523) & (g520) & (!g521) & (g522) & (g529) & (!g530)) + ((g523) & (g520) & (g521) & (!g522) & (g529) & (!g530)) + ((g523) & (g520) & (g521) & (!g522) & (g529) & (g530)));
	assign g578 = (((!g523) & (!g520) & (!g521) & (!g522) & (g529) & (!g530)) + ((!g523) & (!g520) & (!g521) & (g522) & (!g529) & (!g530)) + ((!g523) & (!g520) & (!g521) & (g522) & (g529) & (!g530)) + ((!g523) & (!g520) & (!g521) & (g522) & (g529) & (g530)) + ((!g523) & (!g520) & (g521) & (!g522) & (!g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (!g522) & (!g529) & (g530)) + ((!g523) & (!g520) & (g521) & (!g522) & (g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (g522) & (!g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (g522) & (g529) & (g530)) + ((!g523) & (g520) & (!g521) & (!g522) & (!g529) & (g530)) + ((!g523) & (g520) & (!g521) & (!g522) & (g529) & (!g530)) + ((!g523) & (g520) & (!g521) & (!g522) & (g529) & (g530)) + ((!g523) & (g520) & (g521) & (!g522) & (!g529) & (g530)) + ((!g523) & (g520) & (g521) & (!g522) & (g529) & (!g530)) + ((!g523) & (g520) & (g521) & (!g522) & (g529) & (g530)) + ((!g523) & (g520) & (g521) & (g522) & (!g529) & (!g530)) + ((g523) & (!g520) & (!g521) & (!g522) & (g529) & (!g530)) + ((g523) & (!g520) & (!g521) & (g522) & (!g529) & (!g530)) + ((g523) & (!g520) & (!g521) & (g522) & (g529) & (g530)) + ((g523) & (!g520) & (g521) & (!g522) & (!g529) & (!g530)) + ((g523) & (!g520) & (g521) & (!g522) & (!g529) & (g530)) + ((g523) & (!g520) & (g521) & (g522) & (!g529) & (!g530)) + ((g523) & (!g520) & (g521) & (g522) & (g529) & (!g530)) + ((g523) & (g520) & (!g521) & (!g522) & (g529) & (!g530)) + ((g523) & (g520) & (!g521) & (g522) & (!g529) & (!g530)) + ((g523) & (g520) & (!g521) & (g522) & (g529) & (g530)) + ((g523) & (g520) & (g521) & (!g522) & (!g529) & (!g530)) + ((g523) & (g520) & (g521) & (!g522) & (g529) & (!g530)) + ((g523) & (g520) & (g521) & (!g522) & (g529) & (g530)) + ((g523) & (g520) & (g521) & (g522) & (!g529) & (g530)));
	assign g579 = (((!g523) & (!g520) & (!g521) & (!g522) & (!g529) & (g530)) + ((!g523) & (!g520) & (!g521) & (g522) & (g529) & (!g530)) + ((!g523) & (!g520) & (!g521) & (g522) & (g529) & (g530)) + ((!g523) & (!g520) & (g521) & (!g522) & (!g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (!g522) & (!g529) & (g530)) + ((!g523) & (!g520) & (g521) & (g522) & (g529) & (!g530)) + ((!g523) & (!g520) & (g521) & (g522) & (g529) & (g530)) + ((!g523) & (g520) & (!g521) & (!g522) & (!g529) & (!g530)) + ((!g523) & (g520) & (!g521) & (!g522) & (!g529) & (g530)) + ((!g523) & (g520) & (!g521) & (!g522) & (g529) & (g530)) + ((!g523) & (g520) & (!g521) & (g522) & (!g529) & (g530)) + ((!g523) & (g520) & (g521) & (!g522) & (!g529) & (g530)) + ((!g523) & (g520) & (g521) & (g522) & (!g529) & (!g530)) + ((!g523) & (g520) & (g521) & (g522) & (!g529) & (g530)) + ((!g523) & (g520) & (g521) & (g522) & (g529) & (!g530)) + ((!g523) & (g520) & (g521) & (g522) & (g529) & (g530)) + ((g523) & (!g520) & (!g521) & (g522) & (!g529) & (g530)) + ((g523) & (!g520) & (g521) & (!g522) & (!g529) & (!g530)) + ((g523) & (!g520) & (g521) & (g522) & (!g529) & (!g530)) + ((g523) & (!g520) & (g521) & (g522) & (!g529) & (g530)) + ((g523) & (!g520) & (g521) & (g522) & (g529) & (g530)) + ((g523) & (g520) & (!g521) & (!g522) & (!g529) & (g530)) + ((g523) & (g520) & (!g521) & (!g522) & (g529) & (g530)) + ((g523) & (g520) & (!g521) & (g522) & (!g529) & (!g530)) + ((g523) & (g520) & (!g521) & (g522) & (g529) & (!g530)) + ((g523) & (g520) & (!g521) & (g522) & (g529) & (g530)) + ((g523) & (g520) & (g521) & (!g522) & (g529) & (g530)) + ((g523) & (g520) & (g521) & (g522) & (g529) & (g530)));
	assign g580 = (((!g576) & (!g577) & (!g578) & (!g579) & (!g519) & (g524)) + ((!g576) & (!g577) & (!g578) & (!g579) & (g519) & (!g524)) + ((!g576) & (!g577) & (!g578) & (!g579) & (g519) & (g524)) + ((!g576) & (!g577) & (!g578) & (g579) & (!g519) & (g524)) + ((!g576) & (!g577) & (!g578) & (g579) & (g519) & (!g524)) + ((!g576) & (!g577) & (g578) & (!g579) & (g519) & (!g524)) + ((!g576) & (!g577) & (g578) & (!g579) & (g519) & (g524)) + ((!g576) & (!g577) & (g578) & (g579) & (g519) & (!g524)) + ((!g576) & (g577) & (!g578) & (!g579) & (!g519) & (g524)) + ((!g576) & (g577) & (!g578) & (!g579) & (g519) & (g524)) + ((!g576) & (g577) & (!g578) & (g579) & (!g519) & (g524)) + ((!g576) & (g577) & (g578) & (!g579) & (g519) & (g524)) + ((g576) & (!g577) & (!g578) & (!g579) & (!g519) & (!g524)) + ((g576) & (!g577) & (!g578) & (!g579) & (!g519) & (g524)) + ((g576) & (!g577) & (!g578) & (!g579) & (g519) & (!g524)) + ((g576) & (!g577) & (!g578) & (!g579) & (g519) & (g524)) + ((g576) & (!g577) & (!g578) & (g579) & (!g519) & (!g524)) + ((g576) & (!g577) & (!g578) & (g579) & (!g519) & (g524)) + ((g576) & (!g577) & (!g578) & (g579) & (g519) & (!g524)) + ((g576) & (!g577) & (g578) & (!g579) & (!g519) & (!g524)) + ((g576) & (!g577) & (g578) & (!g579) & (g519) & (!g524)) + ((g576) & (!g577) & (g578) & (!g579) & (g519) & (g524)) + ((g576) & (!g577) & (g578) & (g579) & (!g519) & (!g524)) + ((g576) & (!g577) & (g578) & (g579) & (g519) & (!g524)) + ((g576) & (g577) & (!g578) & (!g579) & (!g519) & (!g524)) + ((g576) & (g577) & (!g578) & (!g579) & (!g519) & (g524)) + ((g576) & (g577) & (!g578) & (!g579) & (g519) & (g524)) + ((g576) & (g577) & (!g578) & (g579) & (!g519) & (!g524)) + ((g576) & (g577) & (!g578) & (g579) & (!g519) & (g524)) + ((g576) & (g577) & (g578) & (!g579) & (!g519) & (!g524)) + ((g576) & (g577) & (g578) & (!g579) & (g519) & (g524)) + ((g576) & (g577) & (g578) & (g579) & (!g519) & (!g524)));
	assign g582 = (((!g580) & (sk[80]) & (g581)) + ((g580) & (!sk[80]) & (!g581)) + ((g580) & (!sk[80]) & (g581)) + ((g580) & (sk[80]) & (!g581)));
	assign g589 = (((!g583) & (!g584) & (!g585) & (!g586) & (g587) & (g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g587) & (!g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g587) & (g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (g587) & (!g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (!g587) & (!g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (!g587) & (g588)) + ((!g583) & (!g584) & (g585) & (g586) & (!g587) & (!g588)) + ((!g583) & (!g584) & (g585) & (g586) & (g587) & (g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (g587) & (!g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (g587) & (g588)) + ((!g583) & (g584) & (!g585) & (g586) & (g587) & (!g588)) + ((!g583) & (g584) & (!g585) & (g586) & (g587) & (g588)) + ((!g583) & (g584) & (g585) & (!g586) & (g587) & (!g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (!g587) & (!g588)) + ((g583) & (!g584) & (g585) & (!g586) & (g587) & (!g588)) + ((g583) & (!g584) & (g585) & (g586) & (!g587) & (g588)) + ((g583) & (!g584) & (g585) & (g586) & (g587) & (g588)) + ((g583) & (g584) & (!g585) & (!g586) & (!g587) & (g588)) + ((g583) & (g584) & (!g585) & (!g586) & (g587) & (!g588)) + ((g583) & (g584) & (g585) & (!g586) & (!g587) & (g588)) + ((g583) & (g584) & (g585) & (!g586) & (g587) & (!g588)) + ((g583) & (g584) & (g585) & (g586) & (!g587) & (!g588)) + ((g583) & (g584) & (g585) & (g586) & (g587) & (!g588)) + ((g583) & (g584) & (g585) & (g586) & (g587) & (g588)));
	assign g590 = (((!g583) & (!g584) & (!g585) & (!g586) & (g587) & (!g588)) + ((!g583) & (!g584) & (!g585) & (!g586) & (g587) & (g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g587) & (!g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g587) & (g588)) + ((!g583) & (!g584) & (g585) & (g586) & (!g587) & (g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (!g587) & (!g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (!g587) & (g588)) + ((!g583) & (g584) & (g585) & (!g586) & (!g587) & (!g588)) + ((!g583) & (g584) & (g585) & (!g586) & (!g587) & (g588)) + ((!g583) & (g584) & (g585) & (!g586) & (g587) & (!g588)) + ((!g583) & (g584) & (g585) & (g586) & (g587) & (g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (!g587) & (g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (g587) & (!g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (g587) & (g588)) + ((g583) & (!g584) & (!g585) & (g586) & (g587) & (!g588)) + ((g583) & (!g584) & (g585) & (!g586) & (!g587) & (!g588)) + ((g583) & (!g584) & (g585) & (!g586) & (g587) & (g588)) + ((g583) & (!g584) & (g585) & (g586) & (!g587) & (g588)) + ((g583) & (!g584) & (g585) & (g586) & (g587) & (g588)) + ((g583) & (g584) & (!g585) & (!g586) & (!g587) & (!g588)) + ((g583) & (g584) & (!g585) & (!g586) & (!g587) & (g588)) + ((g583) & (g584) & (!g585) & (!g586) & (g587) & (!g588)) + ((g583) & (g584) & (!g585) & (!g586) & (g587) & (g588)) + ((g583) & (g584) & (!g585) & (g586) & (!g587) & (!g588)) + ((g583) & (g584) & (!g585) & (g586) & (g587) & (!g588)) + ((g583) & (g584) & (!g585) & (g586) & (g587) & (g588)) + ((g583) & (g584) & (g585) & (!g586) & (g587) & (!g588)) + ((g583) & (g584) & (g585) & (!g586) & (g587) & (g588)) + ((g583) & (g584) & (g585) & (g586) & (!g587) & (g588)) + ((g583) & (g584) & (g585) & (g586) & (g587) & (!g588)));
	assign g591 = (((!g583) & (!g584) & (!g585) & (!g586) & (!g587) & (!g588)) + ((!g583) & (!g584) & (!g585) & (!g586) & (g587) & (g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (g587) & (g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (!g587) & (!g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (!g587) & (g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (g587) & (g588)) + ((!g583) & (!g584) & (g585) & (g586) & (!g587) & (g588)) + ((!g583) & (!g584) & (g585) & (g586) & (g587) & (!g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (!g587) & (!g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (g587) & (!g588)) + ((!g583) & (g584) & (!g585) & (g586) & (g587) & (g588)) + ((!g583) & (g584) & (g585) & (g586) & (!g587) & (!g588)) + ((!g583) & (g584) & (g585) & (g586) & (g587) & (!g588)) + ((g583) & (!g584) & (!g585) & (g586) & (!g587) & (!g588)) + ((g583) & (!g584) & (!g585) & (g586) & (!g587) & (g588)) + ((g583) & (!g584) & (!g585) & (g586) & (g587) & (!g588)) + ((g583) & (!g584) & (g585) & (!g586) & (!g587) & (!g588)) + ((g583) & (!g584) & (g585) & (!g586) & (g587) & (g588)) + ((g583) & (!g584) & (g585) & (g586) & (!g587) & (!g588)) + ((g583) & (!g584) & (g585) & (g586) & (!g587) & (g588)) + ((g583) & (!g584) & (g585) & (g586) & (g587) & (!g588)) + ((g583) & (!g584) & (g585) & (g586) & (g587) & (g588)) + ((g583) & (g584) & (!g585) & (!g586) & (g587) & (g588)) + ((g583) & (g584) & (!g585) & (g586) & (!g587) & (!g588)) + ((g583) & (g584) & (!g585) & (g586) & (g587) & (!g588)) + ((g583) & (g584) & (!g585) & (g586) & (g587) & (g588)) + ((g583) & (g584) & (g585) & (!g586) & (!g587) & (!g588)) + ((g583) & (g584) & (g585) & (g586) & (!g587) & (!g588)) + ((g583) & (g584) & (g585) & (g586) & (!g587) & (g588)) + ((g583) & (g584) & (g585) & (g586) & (g587) & (g588)));
	assign g592 = (((!g583) & (!g584) & (!g585) & (!g586) & (!g587) & (g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (g587) & (!g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (g587) & (g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (!g587) & (g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (g587) & (g588)) + ((!g583) & (!g584) & (g585) & (g586) & (!g587) & (g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (!g587) & (!g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (!g587) & (g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (g587) & (!g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (g587) & (g588)) + ((!g583) & (g584) & (!g585) & (g586) & (g587) & (!g588)) + ((!g583) & (g584) & (!g585) & (g586) & (g587) & (g588)) + ((!g583) & (g584) & (g585) & (g586) & (!g587) & (!g588)) + ((!g583) & (g584) & (g585) & (g586) & (g587) & (!g588)) + ((!g583) & (g584) & (g585) & (g586) & (g587) & (g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (!g587) & (!g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (g587) & (g588)) + ((g583) & (!g584) & (!g585) & (g586) & (g587) & (!g588)) + ((g583) & (!g584) & (!g585) & (g586) & (g587) & (g588)) + ((g583) & (!g584) & (g585) & (!g586) & (!g587) & (g588)) + ((g583) & (!g584) & (g585) & (!g586) & (g587) & (!g588)) + ((g583) & (!g584) & (g585) & (g586) & (g587) & (!g588)) + ((g583) & (g584) & (!g585) & (!g586) & (!g587) & (g588)) + ((g583) & (g584) & (!g585) & (!g586) & (g587) & (g588)) + ((g583) & (g584) & (!g585) & (g586) & (g587) & (!g588)) + ((g583) & (g584) & (!g585) & (g586) & (g587) & (g588)) + ((g583) & (g584) & (g585) & (!g586) & (!g587) & (g588)) + ((g583) & (g584) & (g585) & (g586) & (!g587) & (!g588)));
	assign g595 = (((!g589) & (!g590) & (!g591) & (!g592) & (!g593) & (!g594)) + ((!g589) & (!g590) & (!g591) & (g592) & (!g593) & (!g594)) + ((!g589) & (!g590) & (!g591) & (g592) & (g593) & (g594)) + ((!g589) & (!g590) & (g591) & (!g592) & (!g593) & (!g594)) + ((!g589) & (!g590) & (g591) & (!g592) & (!g593) & (g594)) + ((!g589) & (!g590) & (g591) & (g592) & (!g593) & (!g594)) + ((!g589) & (!g590) & (g591) & (g592) & (!g593) & (g594)) + ((!g589) & (!g590) & (g591) & (g592) & (g593) & (g594)) + ((!g589) & (g590) & (!g591) & (!g592) & (!g593) & (!g594)) + ((!g589) & (g590) & (!g591) & (!g592) & (g593) & (!g594)) + ((!g589) & (g590) & (!g591) & (g592) & (!g593) & (!g594)) + ((!g589) & (g590) & (!g591) & (g592) & (g593) & (!g594)) + ((!g589) & (g590) & (!g591) & (g592) & (g593) & (g594)) + ((!g589) & (g590) & (g591) & (!g592) & (!g593) & (!g594)) + ((!g589) & (g590) & (g591) & (!g592) & (!g593) & (g594)) + ((!g589) & (g590) & (g591) & (!g592) & (g593) & (!g594)) + ((!g589) & (g590) & (g591) & (g592) & (!g593) & (!g594)) + ((!g589) & (g590) & (g591) & (g592) & (!g593) & (g594)) + ((!g589) & (g590) & (g591) & (g592) & (g593) & (!g594)) + ((!g589) & (g590) & (g591) & (g592) & (g593) & (g594)) + ((g589) & (!g590) & (!g591) & (g592) & (g593) & (g594)) + ((g589) & (!g590) & (g591) & (!g592) & (!g593) & (g594)) + ((g589) & (!g590) & (g591) & (g592) & (!g593) & (g594)) + ((g589) & (!g590) & (g591) & (g592) & (g593) & (g594)) + ((g589) & (g590) & (!g591) & (!g592) & (g593) & (!g594)) + ((g589) & (g590) & (!g591) & (g592) & (g593) & (!g594)) + ((g589) & (g590) & (!g591) & (g592) & (g593) & (g594)) + ((g589) & (g590) & (g591) & (!g592) & (!g593) & (g594)) + ((g589) & (g590) & (g591) & (!g592) & (g593) & (!g594)) + ((g589) & (g590) & (g591) & (g592) & (!g593) & (g594)) + ((g589) & (g590) & (g591) & (g592) & (g593) & (!g594)) + ((g589) & (g590) & (g591) & (g592) & (g593) & (g594)));
	assign g597 = (((!sk[86]) & (g595) & (!g596)) + ((!sk[86]) & (g595) & (g596)) + ((sk[86]) & (!g595) & (g596)) + ((sk[86]) & (g595) & (!g596)));
	assign g598 = (((!g583) & (!g584) & (!g585) & (!g586) & (!g593) & (g587)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g593) & (!g587)) + ((!g583) & (!g584) & (!g585) & (g586) & (g593) & (!g587)) + ((!g583) & (!g584) & (g585) & (!g586) & (g593) & (g587)) + ((!g583) & (!g584) & (g585) & (g586) & (!g593) & (g587)) + ((!g583) & (!g584) & (g585) & (g586) & (g593) & (!g587)) + ((!g583) & (g584) & (!g585) & (!g586) & (!g593) & (g587)) + ((!g583) & (g584) & (!g585) & (!g586) & (g593) & (!g587)) + ((!g583) & (g584) & (!g585) & (!g586) & (g593) & (g587)) + ((!g583) & (g584) & (g585) & (!g586) & (g593) & (g587)) + ((!g583) & (g584) & (g585) & (g586) & (g593) & (g587)) + ((g583) & (!g584) & (!g585) & (!g586) & (!g593) & (!g587)) + ((g583) & (!g584) & (!g585) & (!g586) & (g593) & (g587)) + ((g583) & (!g584) & (!g585) & (g586) & (!g593) & (!g587)) + ((g583) & (!g584) & (!g585) & (g586) & (g593) & (!g587)) + ((g583) & (!g584) & (g585) & (!g586) & (g593) & (!g587)) + ((g583) & (!g584) & (g585) & (!g586) & (g593) & (g587)) + ((g583) & (!g584) & (g585) & (g586) & (g593) & (!g587)) + ((g583) & (!g584) & (g585) & (g586) & (g593) & (g587)) + ((g583) & (g584) & (!g585) & (!g586) & (g593) & (!g587)) + ((g583) & (g584) & (!g585) & (!g586) & (g593) & (g587)) + ((g583) & (g584) & (!g585) & (g586) & (g593) & (g587)) + ((g583) & (g584) & (g585) & (!g586) & (!g593) & (!g587)) + ((g583) & (g584) & (g585) & (!g586) & (!g593) & (g587)) + ((g583) & (g584) & (g585) & (!g586) & (g593) & (!g587)) + ((g583) & (g584) & (g585) & (g586) & (!g593) & (g587)) + ((g583) & (g584) & (g585) & (g586) & (g593) & (!g587)));
	assign g599 = (((!g583) & (!g584) & (!g585) & (!g586) & (!g593) & (g587)) + ((!g583) & (!g584) & (!g585) & (!g586) & (g593) & (!g587)) + ((!g583) & (!g584) & (!g585) & (!g586) & (g593) & (g587)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g593) & (!g587)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g593) & (g587)) + ((!g583) & (!g584) & (!g585) & (g586) & (g593) & (g587)) + ((!g583) & (!g584) & (g585) & (!g586) & (g593) & (!g587)) + ((!g583) & (!g584) & (g585) & (g586) & (!g593) & (!g587)) + ((!g583) & (!g584) & (g585) & (g586) & (!g593) & (g587)) + ((!g583) & (!g584) & (g585) & (g586) & (g593) & (g587)) + ((!g583) & (g584) & (!g585) & (!g586) & (g593) & (g587)) + ((!g583) & (g584) & (!g585) & (g586) & (!g593) & (!g587)) + ((!g583) & (g584) & (!g585) & (g586) & (g593) & (!g587)) + ((!g583) & (g584) & (g585) & (!g586) & (g593) & (!g587)) + ((!g583) & (g584) & (g585) & (!g586) & (g593) & (g587)) + ((!g583) & (g584) & (g585) & (g586) & (!g593) & (!g587)) + ((g583) & (!g584) & (!g585) & (!g586) & (!g593) & (!g587)) + ((g583) & (!g584) & (!g585) & (g586) & (!g593) & (!g587)) + ((g583) & (!g584) & (!g585) & (g586) & (!g593) & (g587)) + ((g583) & (!g584) & (g585) & (!g586) & (!g593) & (g587)) + ((g583) & (!g584) & (g585) & (!g586) & (g593) & (g587)) + ((g583) & (!g584) & (g585) & (g586) & (!g593) & (!g587)) + ((g583) & (!g584) & (g585) & (g586) & (!g593) & (g587)) + ((g583) & (g584) & (!g585) & (g586) & (!g593) & (!g587)) + ((g583) & (g584) & (!g585) & (g586) & (g593) & (g587)) + ((g583) & (g584) & (g585) & (!g586) & (!g593) & (!g587)) + ((g583) & (g584) & (g585) & (!g586) & (!g593) & (g587)) + ((g583) & (g584) & (g585) & (!g586) & (g593) & (g587)) + ((g583) & (g584) & (g585) & (g586) & (!g593) & (!g587)) + ((g583) & (g584) & (g585) & (g586) & (!g593) & (g587)) + ((g583) & (g584) & (g585) & (g586) & (g593) & (!g587)));
	assign g600 = (((!g583) & (!g584) & (!g585) & (!g586) & (!g593) & (g587)) + ((!g583) & (!g584) & (!g585) & (g586) & (g593) & (!g587)) + ((!g583) & (!g584) & (g585) & (!g586) & (!g593) & (!g587)) + ((!g583) & (!g584) & (g585) & (!g586) & (g593) & (!g587)) + ((!g583) & (!g584) & (g585) & (g586) & (!g593) & (g587)) + ((!g583) & (!g584) & (g585) & (g586) & (g593) & (!g587)) + ((!g583) & (!g584) & (g585) & (g586) & (g593) & (g587)) + ((!g583) & (g584) & (!g585) & (!g586) & (!g593) & (!g587)) + ((!g583) & (g584) & (!g585) & (!g586) & (g593) & (!g587)) + ((!g583) & (g584) & (!g585) & (g586) & (!g593) & (!g587)) + ((!g583) & (g584) & (!g585) & (g586) & (g593) & (g587)) + ((!g583) & (g584) & (g585) & (!g586) & (g593) & (g587)) + ((!g583) & (g584) & (g585) & (g586) & (!g593) & (g587)) + ((!g583) & (g584) & (g585) & (g586) & (g593) & (!g587)) + ((g583) & (!g584) & (!g585) & (!g586) & (g593) & (g587)) + ((g583) & (!g584) & (!g585) & (g586) & (!g593) & (!g587)) + ((g583) & (!g584) & (!g585) & (g586) & (g593) & (!g587)) + ((g583) & (!g584) & (g585) & (!g586) & (!g593) & (!g587)) + ((g583) & (!g584) & (g585) & (!g586) & (!g593) & (g587)) + ((g583) & (!g584) & (g585) & (!g586) & (g593) & (!g587)) + ((g583) & (!g584) & (g585) & (!g586) & (g593) & (g587)) + ((g583) & (!g584) & (g585) & (g586) & (g593) & (!g587)) + ((g583) & (g584) & (!g585) & (!g586) & (!g593) & (g587)) + ((g583) & (g584) & (!g585) & (!g586) & (g593) & (g587)) + ((g583) & (g584) & (!g585) & (g586) & (!g593) & (g587)) + ((g583) & (g584) & (g585) & (!g586) & (!g593) & (!g587)) + ((g583) & (g584) & (g585) & (!g586) & (!g593) & (g587)) + ((g583) & (g584) & (g585) & (!g586) & (g593) & (g587)) + ((g583) & (g584) & (g585) & (g586) & (!g593) & (!g587)) + ((g583) & (g584) & (g585) & (g586) & (!g593) & (g587)) + ((g583) & (g584) & (g585) & (g586) & (g593) & (!g587)) + ((g583) & (g584) & (g585) & (g586) & (g593) & (g587)));
	assign g601 = (((!g583) & (!g584) & (!g585) & (!g586) & (g593) & (!g587)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g593) & (!g587)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g593) & (g587)) + ((!g583) & (!g584) & (g585) & (!g586) & (g593) & (g587)) + ((!g583) & (!g584) & (g585) & (g586) & (!g593) & (g587)) + ((!g583) & (g584) & (!g585) & (!g586) & (!g593) & (!g587)) + ((!g583) & (g584) & (!g585) & (!g586) & (g593) & (!g587)) + ((!g583) & (g584) & (!g585) & (g586) & (!g593) & (g587)) + ((!g583) & (g584) & (g585) & (!g586) & (!g593) & (g587)) + ((!g583) & (g584) & (g585) & (!g586) & (g593) & (!g587)) + ((!g583) & (g584) & (g585) & (!g586) & (g593) & (g587)) + ((!g583) & (g584) & (g585) & (g586) & (g593) & (!g587)) + ((!g583) & (g584) & (g585) & (g586) & (g593) & (g587)) + ((g583) & (!g584) & (!g585) & (!g586) & (!g593) & (!g587)) + ((g583) & (!g584) & (!g585) & (g586) & (!g593) & (!g587)) + ((g583) & (!g584) & (!g585) & (g586) & (!g593) & (g587)) + ((g583) & (!g584) & (!g585) & (g586) & (g593) & (!g587)) + ((g583) & (!g584) & (g585) & (!g586) & (!g593) & (!g587)) + ((g583) & (!g584) & (g585) & (!g586) & (g593) & (g587)) + ((g583) & (!g584) & (g585) & (g586) & (g593) & (!g587)) + ((g583) & (g584) & (!g585) & (!g586) & (!g593) & (!g587)) + ((g583) & (g584) & (!g585) & (g586) & (!g593) & (!g587)) + ((g583) & (g584) & (!g585) & (g586) & (g593) & (!g587)) + ((g583) & (g584) & (!g585) & (g586) & (g593) & (g587)) + ((g583) & (g584) & (g585) & (g586) & (!g593) & (g587)) + ((g583) & (g584) & (g585) & (g586) & (g593) & (g587)));
	assign g602 = (((!g598) & (!g599) & (!g600) & (!g601) & (!g588) & (!g594)) + ((!g598) & (!g599) & (!g600) & (!g601) & (g588) & (!g594)) + ((!g598) & (!g599) & (!g600) & (g601) & (!g588) & (!g594)) + ((!g598) & (!g599) & (!g600) & (g601) & (g588) & (!g594)) + ((!g598) & (!g599) & (!g600) & (g601) & (g588) & (g594)) + ((!g598) & (!g599) & (g600) & (!g601) & (!g588) & (!g594)) + ((!g598) & (!g599) & (g600) & (!g601) & (!g588) & (g594)) + ((!g598) & (!g599) & (g600) & (!g601) & (g588) & (!g594)) + ((!g598) & (!g599) & (g600) & (g601) & (!g588) & (!g594)) + ((!g598) & (!g599) & (g600) & (g601) & (!g588) & (g594)) + ((!g598) & (!g599) & (g600) & (g601) & (g588) & (!g594)) + ((!g598) & (!g599) & (g600) & (g601) & (g588) & (g594)) + ((!g598) & (g599) & (!g600) & (!g601) & (!g588) & (!g594)) + ((!g598) & (g599) & (!g600) & (g601) & (!g588) & (!g594)) + ((!g598) & (g599) & (!g600) & (g601) & (g588) & (g594)) + ((!g598) & (g599) & (g600) & (!g601) & (!g588) & (!g594)) + ((!g598) & (g599) & (g600) & (!g601) & (!g588) & (g594)) + ((!g598) & (g599) & (g600) & (g601) & (!g588) & (!g594)) + ((!g598) & (g599) & (g600) & (g601) & (!g588) & (g594)) + ((!g598) & (g599) & (g600) & (g601) & (g588) & (g594)) + ((g598) & (!g599) & (!g600) & (!g601) & (g588) & (!g594)) + ((g598) & (!g599) & (!g600) & (g601) & (g588) & (!g594)) + ((g598) & (!g599) & (!g600) & (g601) & (g588) & (g594)) + ((g598) & (!g599) & (g600) & (!g601) & (!g588) & (g594)) + ((g598) & (!g599) & (g600) & (!g601) & (g588) & (!g594)) + ((g598) & (!g599) & (g600) & (g601) & (!g588) & (g594)) + ((g598) & (!g599) & (g600) & (g601) & (g588) & (!g594)) + ((g598) & (!g599) & (g600) & (g601) & (g588) & (g594)) + ((g598) & (g599) & (!g600) & (g601) & (g588) & (g594)) + ((g598) & (g599) & (g600) & (!g601) & (!g588) & (g594)) + ((g598) & (g599) & (g600) & (g601) & (!g588) & (g594)) + ((g598) & (g599) & (g600) & (g601) & (g588) & (g594)));
	assign g604 = (((!g602) & (sk[92]) & (g603)) + ((g602) & (!sk[92]) & (!g603)) + ((g602) & (!sk[92]) & (g603)) + ((g602) & (sk[92]) & (!g603)));
	assign g605 = (((!g587) & (!g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((!g587) & (!g584) & (!g585) & (!g586) & (g593) & (g588)) + ((!g587) & (!g584) & (!g585) & (g586) & (!g593) & (g588)) + ((!g587) & (!g584) & (!g585) & (g586) & (g593) & (!g588)) + ((!g587) & (!g584) & (!g585) & (g586) & (g593) & (g588)) + ((!g587) & (!g584) & (g585) & (!g586) & (!g593) & (g588)) + ((!g587) & (!g584) & (g585) & (g586) & (!g593) & (!g588)) + ((!g587) & (!g584) & (g585) & (g586) & (g593) & (!g588)) + ((!g587) & (g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((!g587) & (g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((!g587) & (g584) & (!g585) & (g586) & (!g593) & (g588)) + ((!g587) & (g584) & (g585) & (!g586) & (!g593) & (!g588)) + ((!g587) & (g584) & (g585) & (!g586) & (!g593) & (g588)) + ((!g587) & (g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g587) & (g584) & (g585) & (!g586) & (g593) & (g588)) + ((g587) & (!g584) & (!g585) & (g586) & (!g593) & (g588)) + ((g587) & (!g584) & (!g585) & (g586) & (g593) & (g588)) + ((g587) & (g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((g587) & (g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((g587) & (g584) & (!g585) & (g586) & (g593) & (!g588)) + ((g587) & (g584) & (g585) & (g586) & (!g593) & (!g588)) + ((g587) & (g584) & (g585) & (g586) & (!g593) & (g588)));
	assign g606 = (((!g587) & (!g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((!g587) & (!g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((!g587) & (!g584) & (!g585) & (g586) & (g593) & (g588)) + ((!g587) & (!g584) & (g585) & (!g586) & (!g593) & (!g588)) + ((!g587) & (!g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g587) & (!g584) & (g585) & (g586) & (!g593) & (g588)) + ((!g587) & (g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((!g587) & (g584) & (!g585) & (!g586) & (g593) & (g588)) + ((!g587) & (g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((!g587) & (g584) & (!g585) & (g586) & (!g593) & (g588)) + ((!g587) & (g584) & (!g585) & (g586) & (g593) & (g588)) + ((!g587) & (g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g587) & (g584) & (g585) & (!g586) & (g593) & (g588)) + ((!g587) & (g584) & (g585) & (g586) & (g593) & (!g588)) + ((g587) & (!g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((g587) & (!g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((g587) & (!g584) & (!g585) & (!g586) & (g593) & (g588)) + ((g587) & (!g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((g587) & (!g584) & (!g585) & (g586) & (!g593) & (g588)) + ((g587) & (!g584) & (!g585) & (g586) & (g593) & (!g588)) + ((g587) & (!g584) & (g585) & (g586) & (!g593) & (!g588)) + ((g587) & (g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((g587) & (g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((g587) & (g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((g587) & (g584) & (!g585) & (g586) & (g593) & (!g588)) + ((g587) & (g584) & (!g585) & (g586) & (g593) & (g588)) + ((g587) & (g584) & (g585) & (!g586) & (!g593) & (!g588)) + ((g587) & (g584) & (g585) & (!g586) & (g593) & (!g588)) + ((g587) & (g584) & (g585) & (g586) & (!g593) & (g588)) + ((g587) & (g584) & (g585) & (g586) & (g593) & (g588)));
	assign g607 = (((!g587) & (!g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((!g587) & (!g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((!g587) & (!g584) & (!g585) & (g586) & (!g593) & (g588)) + ((!g587) & (!g584) & (g585) & (!g586) & (!g593) & (g588)) + ((!g587) & (!g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g587) & (!g584) & (g585) & (g586) & (!g593) & (g588)) + ((!g587) & (g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((!g587) & (g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((!g587) & (g584) & (!g585) & (g586) & (g593) & (!g588)) + ((!g587) & (g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g587) & (g584) & (g585) & (g586) & (!g593) & (!g588)) + ((!g587) & (g584) & (g585) & (g586) & (g593) & (!g588)) + ((g587) & (!g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((g587) & (!g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((g587) & (!g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((g587) & (!g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((g587) & (!g584) & (!g585) & (g586) & (!g593) & (g588)) + ((g587) & (!g584) & (!g585) & (g586) & (g593) & (!g588)) + ((g587) & (!g584) & (!g585) & (g586) & (g593) & (g588)) + ((g587) & (!g584) & (g585) & (!g586) & (!g593) & (g588)) + ((g587) & (!g584) & (g585) & (!g586) & (g593) & (!g588)) + ((g587) & (!g584) & (g585) & (g586) & (!g593) & (!g588)) + ((g587) & (!g584) & (g585) & (g586) & (g593) & (g588)) + ((g587) & (g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((g587) & (g584) & (!g585) & (!g586) & (g593) & (g588)) + ((g587) & (g584) & (g585) & (!g586) & (g593) & (g588)) + ((g587) & (g584) & (g585) & (g586) & (!g593) & (!g588)) + ((g587) & (g584) & (g585) & (g586) & (!g593) & (g588)) + ((g587) & (g584) & (g585) & (g586) & (g593) & (g588)));
	assign g608 = (((!g587) & (!g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((!g587) & (!g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((!g587) & (!g584) & (!g585) & (!g586) & (g593) & (g588)) + ((!g587) & (!g584) & (!g585) & (g586) & (!g593) & (g588)) + ((!g587) & (!g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g587) & (!g584) & (g585) & (g586) & (g593) & (g588)) + ((!g587) & (g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((!g587) & (g584) & (!g585) & (g586) & (!g593) & (g588)) + ((!g587) & (g584) & (!g585) & (g586) & (g593) & (g588)) + ((!g587) & (g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g587) & (g584) & (g585) & (!g586) & (g593) & (g588)) + ((!g587) & (g584) & (g585) & (g586) & (!g593) & (!g588)) + ((!g587) & (g584) & (g585) & (g586) & (!g593) & (g588)) + ((!g587) & (g584) & (g585) & (g586) & (g593) & (!g588)) + ((!g587) & (g584) & (g585) & (g586) & (g593) & (g588)) + ((g587) & (!g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((g587) & (!g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((g587) & (!g584) & (!g585) & (!g586) & (g593) & (g588)) + ((g587) & (!g584) & (!g585) & (g586) & (g593) & (g588)) + ((g587) & (!g584) & (g585) & (!g586) & (!g593) & (g588)) + ((g587) & (!g584) & (g585) & (!g586) & (g593) & (!g588)) + ((g587) & (!g584) & (g585) & (g586) & (g593) & (!g588)) + ((g587) & (g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((g587) & (g584) & (!g585) & (g586) & (!g593) & (g588)) + ((g587) & (g584) & (!g585) & (g586) & (g593) & (!g588)) + ((g587) & (g584) & (g585) & (!g586) & (g593) & (g588)) + ((g587) & (g584) & (g585) & (g586) & (!g593) & (!g588)));
	assign g609 = (((!g605) & (!g606) & (!g607) & (!g608) & (!g583) & (g594)) + ((!g605) & (!g606) & (!g607) & (!g608) & (g583) & (!g594)) + ((!g605) & (!g606) & (!g607) & (!g608) & (g583) & (g594)) + ((!g605) & (!g606) & (!g607) & (g608) & (!g583) & (g594)) + ((!g605) & (!g606) & (!g607) & (g608) & (g583) & (!g594)) + ((!g605) & (!g606) & (g607) & (!g608) & (g583) & (!g594)) + ((!g605) & (!g606) & (g607) & (!g608) & (g583) & (g594)) + ((!g605) & (!g606) & (g607) & (g608) & (g583) & (!g594)) + ((!g605) & (g606) & (!g607) & (!g608) & (!g583) & (g594)) + ((!g605) & (g606) & (!g607) & (!g608) & (g583) & (g594)) + ((!g605) & (g606) & (!g607) & (g608) & (!g583) & (g594)) + ((!g605) & (g606) & (g607) & (!g608) & (g583) & (g594)) + ((g605) & (!g606) & (!g607) & (!g608) & (!g583) & (!g594)) + ((g605) & (!g606) & (!g607) & (!g608) & (!g583) & (g594)) + ((g605) & (!g606) & (!g607) & (!g608) & (g583) & (!g594)) + ((g605) & (!g606) & (!g607) & (!g608) & (g583) & (g594)) + ((g605) & (!g606) & (!g607) & (g608) & (!g583) & (!g594)) + ((g605) & (!g606) & (!g607) & (g608) & (!g583) & (g594)) + ((g605) & (!g606) & (!g607) & (g608) & (g583) & (!g594)) + ((g605) & (!g606) & (g607) & (!g608) & (!g583) & (!g594)) + ((g605) & (!g606) & (g607) & (!g608) & (g583) & (!g594)) + ((g605) & (!g606) & (g607) & (!g608) & (g583) & (g594)) + ((g605) & (!g606) & (g607) & (g608) & (!g583) & (!g594)) + ((g605) & (!g606) & (g607) & (g608) & (g583) & (!g594)) + ((g605) & (g606) & (!g607) & (!g608) & (!g583) & (!g594)) + ((g605) & (g606) & (!g607) & (!g608) & (!g583) & (g594)) + ((g605) & (g606) & (!g607) & (!g608) & (g583) & (g594)) + ((g605) & (g606) & (!g607) & (g608) & (!g583) & (!g594)) + ((g605) & (g606) & (!g607) & (g608) & (!g583) & (g594)) + ((g605) & (g606) & (g607) & (!g608) & (!g583) & (!g594)) + ((g605) & (g606) & (g607) & (!g608) & (g583) & (g594)) + ((g605) & (g606) & (g607) & (g608) & (!g583) & (!g594)));
	assign g611 = (((!sk[98]) & (g609) & (!g610)) + ((!sk[98]) & (g609) & (g610)) + ((sk[98]) & (!g609) & (g610)) + ((sk[98]) & (g609) & (!g610)));
	assign g612 = (((!g583) & (!g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (g593) & (g588)) + ((!g583) & (!g584) & (g585) & (g586) & (!g593) & (!g588)) + ((!g583) & (!g584) & (g585) & (g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (g585) & (g586) & (g593) & (g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (g584) & (g585) & (!g586) & (!g593) & (!g588)) + ((!g583) & (g584) & (g585) & (g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((g583) & (!g584) & (g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (g585) & (!g586) & (!g593) & (g588)) + ((g583) & (!g584) & (g585) & (!g586) & (g593) & (!g588)) + ((g583) & (!g584) & (g585) & (g586) & (!g593) & (g588)) + ((g583) & (g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((g583) & (g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((g583) & (g584) & (!g585) & (g586) & (g593) & (!g588)) + ((g583) & (g584) & (g585) & (!g586) & (!g593) & (g588)) + ((g583) & (g584) & (g585) & (!g586) & (g593) & (g588)));
	assign g613 = (((!g583) & (!g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (!g585) & (!g586) & (g593) & (g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (g585) & (g586) & (!g593) & (!g588)) + ((!g583) & (!g584) & (g585) & (g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (g585) & (g586) & (g593) & (g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (g593) & (g588)) + ((!g583) & (g584) & (!g585) & (g586) & (g593) & (g588)) + ((!g583) & (g584) & (g585) & (!g586) & (!g593) & (!g588)) + ((!g583) & (g584) & (g585) & (!g586) & (!g593) & (g588)) + ((!g583) & (g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (g584) & (g585) & (g586) & (!g593) & (g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((g583) & (!g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (!g585) & (g586) & (!g593) & (g588)) + ((g583) & (!g584) & (!g585) & (g586) & (g593) & (g588)) + ((g583) & (!g584) & (g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (g585) & (!g586) & (!g593) & (g588)) + ((g583) & (!g584) & (g585) & (!g586) & (g593) & (g588)) + ((g583) & (!g584) & (g585) & (g586) & (!g593) & (g588)) + ((g583) & (g584) & (!g585) & (g586) & (!g593) & (g588)) + ((g583) & (g584) & (!g585) & (g586) & (g593) & (!g588)) + ((g583) & (g584) & (g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (g584) & (g585) & (g586) & (!g593) & (!g588)));
	assign g614 = (((!g583) & (!g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (!g585) & (!g586) & (g593) & (g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (g585) & (!g586) & (g593) & (g588)) + ((!g583) & (!g584) & (g585) & (g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (g585) & (g586) & (g593) & (g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (g593) & (g588)) + ((!g583) & (g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((!g583) & (g584) & (!g585) & (g586) & (!g593) & (g588)) + ((!g583) & (g584) & (g585) & (!g586) & (!g593) & (g588)) + ((!g583) & (g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (g584) & (g585) & (g586) & (g593) & (g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (g593) & (g588)) + ((g583) & (!g584) & (!g585) & (g586) & (g593) & (g588)) + ((g583) & (!g584) & (g585) & (g586) & (!g593) & (!g588)) + ((g583) & (g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((g583) & (g584) & (!g585) & (g586) & (g593) & (g588)) + ((g583) & (g584) & (g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (g584) & (g585) & (!g586) & (!g593) & (g588)) + ((g583) & (g584) & (g585) & (!g586) & (g593) & (g588)) + ((g583) & (g584) & (g585) & (g586) & (!g593) & (!g588)) + ((g583) & (g584) & (g585) & (g586) & (g593) & (g588)));
	assign g615 = (((!g583) & (!g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (!g585) & (g586) & (g593) & (g588)) + ((!g583) & (!g584) & (g585) & (g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (g585) & (g586) & (g593) & (g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (!g593) & (!g588)) + ((!g583) & (g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (g584) & (!g585) & (g586) & (!g593) & (!g588)) + ((!g583) & (g584) & (!g585) & (g586) & (!g593) & (g588)) + ((!g583) & (g584) & (!g585) & (g586) & (g593) & (!g588)) + ((!g583) & (g584) & (g585) & (!g586) & (!g593) & (!g588)) + ((!g583) & (g584) & (g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (g584) & (g585) & (!g586) & (g593) & (g588)) + ((g583) & (!g584) & (!g585) & (!g586) & (g593) & (g588)) + ((g583) & (!g584) & (!g585) & (g586) & (g593) & (!g588)) + ((g583) & (!g584) & (g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (g585) & (!g586) & (g593) & (!g588)) + ((g583) & (!g584) & (g585) & (!g586) & (g593) & (g588)) + ((g583) & (!g584) & (g585) & (g586) & (!g593) & (g588)) + ((g583) & (!g584) & (g585) & (g586) & (g593) & (!g588)) + ((g583) & (!g584) & (g585) & (g586) & (g593) & (g588)) + ((g583) & (g584) & (!g585) & (!g586) & (!g593) & (g588)) + ((g583) & (g584) & (!g585) & (!g586) & (g593) & (!g588)) + ((g583) & (g584) & (g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (g584) & (g585) & (!g586) & (!g593) & (g588)) + ((g583) & (g584) & (g585) & (g586) & (g593) & (g588)));
	assign g616 = (((!g612) & (!g613) & (!g614) & (!g615) & (!g594) & (g587)) + ((!g612) & (!g613) & (!g614) & (!g615) & (g594) & (!g587)) + ((!g612) & (!g613) & (!g614) & (!g615) & (g594) & (g587)) + ((!g612) & (!g613) & (!g614) & (g615) & (!g594) & (g587)) + ((!g612) & (!g613) & (!g614) & (g615) & (g594) & (!g587)) + ((!g612) & (!g613) & (g614) & (!g615) & (g594) & (!g587)) + ((!g612) & (!g613) & (g614) & (!g615) & (g594) & (g587)) + ((!g612) & (!g613) & (g614) & (g615) & (g594) & (!g587)) + ((!g612) & (g613) & (!g614) & (!g615) & (!g594) & (g587)) + ((!g612) & (g613) & (!g614) & (!g615) & (g594) & (g587)) + ((!g612) & (g613) & (!g614) & (g615) & (!g594) & (g587)) + ((!g612) & (g613) & (g614) & (!g615) & (g594) & (g587)) + ((g612) & (!g613) & (!g614) & (!g615) & (!g594) & (!g587)) + ((g612) & (!g613) & (!g614) & (!g615) & (!g594) & (g587)) + ((g612) & (!g613) & (!g614) & (!g615) & (g594) & (!g587)) + ((g612) & (!g613) & (!g614) & (!g615) & (g594) & (g587)) + ((g612) & (!g613) & (!g614) & (g615) & (!g594) & (!g587)) + ((g612) & (!g613) & (!g614) & (g615) & (!g594) & (g587)) + ((g612) & (!g613) & (!g614) & (g615) & (g594) & (!g587)) + ((g612) & (!g613) & (g614) & (!g615) & (!g594) & (!g587)) + ((g612) & (!g613) & (g614) & (!g615) & (g594) & (!g587)) + ((g612) & (!g613) & (g614) & (!g615) & (g594) & (g587)) + ((g612) & (!g613) & (g614) & (g615) & (!g594) & (!g587)) + ((g612) & (!g613) & (g614) & (g615) & (g594) & (!g587)) + ((g612) & (g613) & (!g614) & (!g615) & (!g594) & (!g587)) + ((g612) & (g613) & (!g614) & (!g615) & (!g594) & (g587)) + ((g612) & (g613) & (!g614) & (!g615) & (g594) & (g587)) + ((g612) & (g613) & (!g614) & (g615) & (!g594) & (!g587)) + ((g612) & (g613) & (!g614) & (g615) & (!g594) & (g587)) + ((g612) & (g613) & (g614) & (!g615) & (!g594) & (!g587)) + ((g612) & (g613) & (g614) & (!g615) & (g594) & (g587)) + ((g612) & (g613) & (g614) & (g615) & (!g594) & (!g587)));
	assign g618 = (((!g616) & (sk[104]) & (g617)) + ((g616) & (!sk[104]) & (!g617)) + ((g616) & (!sk[104]) & (g617)) + ((g616) & (sk[104]) & (!g617)));
	assign g619 = (((!g583) & (!g584) & (!g587) & (!g594) & (!g593) & (g588)) + ((!g583) & (!g584) & (g587) & (!g594) & (!g593) & (g588)) + ((!g583) & (!g584) & (g587) & (!g594) & (g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (!g594) & (g593) & (g588)) + ((!g583) & (!g584) & (g587) & (g594) & (!g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (g594) & (g593) & (!g588)) + ((!g583) & (g584) & (!g587) & (!g594) & (!g593) & (!g588)) + ((!g583) & (g584) & (!g587) & (!g594) & (!g593) & (g588)) + ((!g583) & (g584) & (!g587) & (g594) & (!g593) & (!g588)) + ((!g583) & (g584) & (!g587) & (g594) & (!g593) & (g588)) + ((!g583) & (g584) & (!g587) & (g594) & (g593) & (g588)) + ((!g583) & (g584) & (g587) & (g594) & (!g593) & (g588)) + ((!g583) & (g584) & (g587) & (g594) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g594) & (!g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g594) & (!g593) & (g588)) + ((g583) & (!g584) & (!g587) & (g594) & (!g593) & (g588)) + ((g583) & (!g584) & (g587) & (!g594) & (g593) & (!g588)) + ((g583) & (!g584) & (g587) & (g594) & (!g593) & (!g588)) + ((g583) & (!g584) & (g587) & (g594) & (!g593) & (g588)) + ((g583) & (!g584) & (g587) & (g594) & (g593) & (!g588)) + ((g583) & (g584) & (!g587) & (!g594) & (!g593) & (!g588)) + ((g583) & (g584) & (!g587) & (!g594) & (g593) & (!g588)) + ((g583) & (g584) & (!g587) & (g594) & (g593) & (!g588)) + ((g583) & (g584) & (g587) & (!g594) & (!g593) & (!g588)) + ((g583) & (g584) & (g587) & (!g594) & (!g593) & (g588)) + ((g583) & (g584) & (g587) & (g594) & (!g593) & (g588)));
	assign g620 = (((!g583) & (!g584) & (!g587) & (!g594) & (!g593) & (!g588)) + ((!g583) & (!g584) & (!g587) & (!g594) & (!g593) & (g588)) + ((!g583) & (!g584) & (!g587) & (!g594) & (g593) & (!g588)) + ((!g583) & (!g584) & (!g587) & (!g594) & (g593) & (g588)) + ((!g583) & (!g584) & (!g587) & (g594) & (!g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (!g594) & (!g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (!g594) & (g593) & (g588)) + ((!g583) & (!g584) & (g587) & (g594) & (!g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (g594) & (g593) & (g588)) + ((!g583) & (g584) & (!g587) & (!g594) & (!g593) & (g588)) + ((!g583) & (g584) & (!g587) & (g594) & (g593) & (!g588)) + ((!g583) & (g584) & (g587) & (!g594) & (!g593) & (!g588)) + ((!g583) & (g584) & (g587) & (!g594) & (!g593) & (g588)) + ((!g583) & (g584) & (g587) & (!g594) & (g593) & (!g588)) + ((!g583) & (g584) & (g587) & (!g594) & (g593) & (g588)) + ((!g583) & (g584) & (g587) & (g594) & (!g593) & (!g588)) + ((!g583) & (g584) & (g587) & (g594) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g594) & (!g593) & (g588)) + ((g583) & (!g584) & (!g587) & (!g594) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g594) & (g593) & (g588)) + ((g583) & (!g584) & (!g587) & (g594) & (!g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (g594) & (g593) & (g588)) + ((g583) & (!g584) & (g587) & (!g594) & (g593) & (!g588)) + ((g583) & (!g584) & (g587) & (!g594) & (g593) & (g588)) + ((g583) & (!g584) & (g587) & (g594) & (!g593) & (g588)) + ((g583) & (g584) & (!g587) & (!g594) & (g593) & (!g588)) + ((g583) & (g584) & (!g587) & (!g594) & (g593) & (g588)) + ((g583) & (g584) & (!g587) & (g594) & (!g593) & (!g588)) + ((g583) & (g584) & (!g587) & (g594) & (!g593) & (g588)) + ((g583) & (g584) & (g587) & (!g594) & (g593) & (!g588)) + ((g583) & (g584) & (g587) & (!g594) & (g593) & (g588)) + ((g583) & (g584) & (g587) & (g594) & (!g593) & (g588)));
	assign g621 = (((!g583) & (!g584) & (!g587) & (!g594) & (!g593) & (!g588)) + ((!g583) & (!g584) & (!g587) & (!g594) & (!g593) & (g588)) + ((!g583) & (!g584) & (g587) & (!g594) & (!g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (!g594) & (g593) & (g588)) + ((!g583) & (!g584) & (g587) & (g594) & (!g593) & (g588)) + ((!g583) & (g584) & (!g587) & (g594) & (!g593) & (!g588)) + ((!g583) & (g584) & (!g587) & (g594) & (g593) & (!g588)) + ((!g583) & (g584) & (!g587) & (g594) & (g593) & (g588)) + ((!g583) & (g584) & (g587) & (!g594) & (!g593) & (!g588)) + ((!g583) & (g584) & (g587) & (!g594) & (g593) & (!g588)) + ((!g583) & (g584) & (g587) & (!g594) & (g593) & (g588)) + ((!g583) & (g584) & (g587) & (g594) & (!g593) & (!g588)) + ((!g583) & (g584) & (g587) & (g594) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g594) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g594) & (g593) & (g588)) + ((g583) & (!g584) & (!g587) & (g594) & (!g593) & (g588)) + ((g583) & (!g584) & (!g587) & (g594) & (g593) & (g588)) + ((g583) & (!g584) & (g587) & (!g594) & (!g593) & (!g588)) + ((g583) & (!g584) & (g587) & (!g594) & (!g593) & (g588)) + ((g583) & (!g584) & (g587) & (!g594) & (g593) & (g588)) + ((g583) & (!g584) & (g587) & (g594) & (!g593) & (!g588)) + ((g583) & (!g584) & (g587) & (g594) & (!g593) & (g588)) + ((g583) & (!g584) & (g587) & (g594) & (g593) & (!g588)) + ((g583) & (!g584) & (g587) & (g594) & (g593) & (g588)) + ((g583) & (g584) & (!g587) & (!g594) & (!g593) & (g588)) + ((g583) & (g584) & (!g587) & (g594) & (!g593) & (!g588)) + ((g583) & (g584) & (!g587) & (g594) & (g593) & (!g588)) + ((g583) & (g584) & (g587) & (!g594) & (!g593) & (!g588)) + ((g583) & (g584) & (g587) & (!g594) & (!g593) & (g588)) + ((g583) & (g584) & (g587) & (!g594) & (g593) & (!g588)) + ((g583) & (g584) & (g587) & (g594) & (!g593) & (!g588)) + ((g583) & (g584) & (g587) & (g594) & (g593) & (!g588)));
	assign g622 = (((!g583) & (!g584) & (!g587) & (!g594) & (g593) & (g588)) + ((!g583) & (!g584) & (!g587) & (g594) & (!g593) & (!g588)) + ((!g583) & (!g584) & (!g587) & (g594) & (g593) & (g588)) + ((!g583) & (!g584) & (g587) & (!g594) & (!g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (!g594) & (g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (g594) & (!g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (g594) & (!g593) & (g588)) + ((!g583) & (!g584) & (g587) & (g594) & (g593) & (!g588)) + ((!g583) & (g584) & (!g587) & (!g594) & (!g593) & (!g588)) + ((!g583) & (g584) & (!g587) & (g594) & (!g593) & (g588)) + ((!g583) & (g584) & (!g587) & (g594) & (g593) & (!g588)) + ((!g583) & (g584) & (!g587) & (g594) & (g593) & (g588)) + ((!g583) & (g584) & (g587) & (!g594) & (!g593) & (!g588)) + ((!g583) & (g584) & (g587) & (g594) & (!g593) & (!g588)) + ((!g583) & (g584) & (g587) & (g594) & (!g593) & (g588)) + ((g583) & (!g584) & (!g587) & (!g594) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g594) & (g593) & (g588)) + ((g583) & (!g584) & (g587) & (!g594) & (!g593) & (!g588)) + ((g583) & (!g584) & (g587) & (!g594) & (g593) & (!g588)) + ((g583) & (!g584) & (g587) & (g594) & (g593) & (!g588)) + ((g583) & (g584) & (!g587) & (!g594) & (g593) & (!g588)) + ((g583) & (g584) & (!g587) & (g594) & (g593) & (g588)) + ((g583) & (g584) & (g587) & (!g594) & (!g593) & (!g588)) + ((g583) & (g584) & (g587) & (!g594) & (!g593) & (g588)) + ((g583) & (g584) & (g587) & (!g594) & (g593) & (!g588)) + ((g583) & (g584) & (g587) & (g594) & (!g593) & (!g588)));
	assign g623 = (((!g619) & (!g620) & (!g621) & (!g622) & (g585) & (g586)) + ((!g619) & (!g620) & (g621) & (!g622) & (!g585) & (g586)) + ((!g619) & (!g620) & (g621) & (!g622) & (g585) & (g586)) + ((!g619) & (!g620) & (g621) & (g622) & (!g585) & (g586)) + ((!g619) & (g620) & (!g621) & (!g622) & (g585) & (!g586)) + ((!g619) & (g620) & (!g621) & (!g622) & (g585) & (g586)) + ((!g619) & (g620) & (!g621) & (g622) & (g585) & (!g586)) + ((!g619) & (g620) & (g621) & (!g622) & (!g585) & (g586)) + ((!g619) & (g620) & (g621) & (!g622) & (g585) & (!g586)) + ((!g619) & (g620) & (g621) & (!g622) & (g585) & (g586)) + ((!g619) & (g620) & (g621) & (g622) & (!g585) & (g586)) + ((!g619) & (g620) & (g621) & (g622) & (g585) & (!g586)) + ((g619) & (!g620) & (!g621) & (!g622) & (!g585) & (!g586)) + ((g619) & (!g620) & (!g621) & (!g622) & (g585) & (g586)) + ((g619) & (!g620) & (!g621) & (g622) & (!g585) & (!g586)) + ((g619) & (!g620) & (g621) & (!g622) & (!g585) & (!g586)) + ((g619) & (!g620) & (g621) & (!g622) & (!g585) & (g586)) + ((g619) & (!g620) & (g621) & (!g622) & (g585) & (g586)) + ((g619) & (!g620) & (g621) & (g622) & (!g585) & (!g586)) + ((g619) & (!g620) & (g621) & (g622) & (!g585) & (g586)) + ((g619) & (g620) & (!g621) & (!g622) & (!g585) & (!g586)) + ((g619) & (g620) & (!g621) & (!g622) & (g585) & (!g586)) + ((g619) & (g620) & (!g621) & (!g622) & (g585) & (g586)) + ((g619) & (g620) & (!g621) & (g622) & (!g585) & (!g586)) + ((g619) & (g620) & (!g621) & (g622) & (g585) & (!g586)) + ((g619) & (g620) & (g621) & (!g622) & (!g585) & (!g586)) + ((g619) & (g620) & (g621) & (!g622) & (!g585) & (g586)) + ((g619) & (g620) & (g621) & (!g622) & (g585) & (!g586)) + ((g619) & (g620) & (g621) & (!g622) & (g585) & (g586)) + ((g619) & (g620) & (g621) & (g622) & (!g585) & (!g586)) + ((g619) & (g620) & (g621) & (g622) & (!g585) & (g586)) + ((g619) & (g620) & (g621) & (g622) & (g585) & (!g586)));
	assign g625 = (((!sk[110]) & (g623) & (!g624)) + ((!sk[110]) & (g623) & (g624)) + ((sk[110]) & (!g623) & (g624)) + ((sk[110]) & (g623) & (!g624)));
	assign g626 = (((!g583) & (!g584) & (!g587) & (!g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (!g587) & (!g586) & (g593) & (g588)) + ((!g583) & (!g584) & (!g587) & (g586) & (g593) & (g588)) + ((!g583) & (!g584) & (g587) & (!g586) & (!g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (!g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (g587) & (!g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (!g586) & (g593) & (g588)) + ((!g583) & (!g584) & (g587) & (g586) & (!g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (g586) & (!g593) & (g588)) + ((!g583) & (g584) & (!g587) & (!g586) & (!g593) & (g588)) + ((!g583) & (g584) & (!g587) & (!g586) & (g593) & (!g588)) + ((!g583) & (g584) & (!g587) & (g586) & (g593) & (g588)) + ((!g583) & (g584) & (g587) & (!g586) & (g593) & (!g588)) + ((!g583) & (g584) & (g587) & (!g586) & (g593) & (g588)) + ((!g583) & (g584) & (g587) & (g586) & (!g593) & (!g588)) + ((!g583) & (g584) & (g587) & (g586) & (!g593) & (g588)) + ((!g583) & (g584) & (g587) & (g586) & (g593) & (g588)) + ((g583) & (!g584) & (!g587) & (!g586) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g586) & (g593) & (g588)) + ((g583) & (!g584) & (!g587) & (g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (g586) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (g586) & (g593) & (g588)) + ((g583) & (!g584) & (g587) & (!g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (g587) & (!g586) & (g593) & (!g588)) + ((g583) & (!g584) & (g587) & (g586) & (g593) & (!g588)) + ((g583) & (g584) & (!g587) & (!g586) & (g593) & (g588)) + ((g583) & (g584) & (g587) & (!g586) & (!g593) & (!g588)) + ((g583) & (g584) & (g587) & (!g586) & (g593) & (g588)));
	assign g627 = (((!g583) & (!g584) & (!g587) & (!g586) & (!g593) & (!g588)) + ((!g583) & (!g584) & (!g587) & (g586) & (!g593) & (!g588)) + ((!g583) & (!g584) & (!g587) & (g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (!g587) & (g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (!g586) & (g593) & (g588)) + ((!g583) & (!g584) & (g587) & (g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (g587) & (g586) & (g593) & (g588)) + ((!g583) & (g584) & (!g587) & (!g586) & (!g593) & (!g588)) + ((!g583) & (g584) & (!g587) & (!g586) & (g593) & (!g588)) + ((!g583) & (g584) & (g587) & (!g586) & (!g593) & (g588)) + ((!g583) & (g584) & (g587) & (!g586) & (g593) & (g588)) + ((!g583) & (g584) & (g587) & (g586) & (!g593) & (g588)) + ((!g583) & (g584) & (g587) & (g586) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g586) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g586) & (g593) & (g588)) + ((g583) & (!g584) & (!g587) & (g586) & (!g593) & (g588)) + ((g583) & (!g584) & (!g587) & (g586) & (g593) & (g588)) + ((g583) & (!g584) & (g587) & (g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (g587) & (g586) & (!g593) & (g588)) + ((g583) & (!g584) & (g587) & (g586) & (g593) & (g588)) + ((g583) & (g584) & (!g587) & (!g586) & (!g593) & (g588)) + ((g583) & (g584) & (!g587) & (!g586) & (g593) & (!g588)) + ((g583) & (g584) & (!g587) & (g586) & (g593) & (!g588)) + ((g583) & (g584) & (g587) & (!g586) & (!g593) & (g588)) + ((g583) & (g584) & (g587) & (!g586) & (g593) & (g588)) + ((g583) & (g584) & (g587) & (g586) & (!g593) & (!g588)) + ((g583) & (g584) & (g587) & (g586) & (g593) & (g588)));
	assign g628 = (((!g583) & (!g584) & (!g587) & (!g586) & (g593) & (g588)) + ((!g583) & (!g584) & (!g587) & (g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (!g586) & (!g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (!g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (g587) & (!g586) & (g593) & (g588)) + ((!g583) & (!g584) & (g587) & (g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (g587) & (g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (g587) & (g586) & (g593) & (g588)) + ((!g583) & (g584) & (!g587) & (!g586) & (g593) & (!g588)) + ((!g583) & (g584) & (!g587) & (!g586) & (g593) & (g588)) + ((!g583) & (g584) & (g587) & (!g586) & (!g593) & (!g588)) + ((!g583) & (g584) & (g587) & (g586) & (!g593) & (g588)) + ((!g583) & (g584) & (g587) & (g586) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g586) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (!g586) & (g593) & (g588)) + ((g583) & (!g584) & (!g587) & (g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (g586) & (!g593) & (g588)) + ((g583) & (!g584) & (g587) & (!g586) & (!g593) & (g588)) + ((g583) & (!g584) & (g587) & (!g586) & (g593) & (g588)) + ((g583) & (!g584) & (g587) & (g586) & (g593) & (!g588)) + ((g583) & (g584) & (!g587) & (!g586) & (!g593) & (!g588)) + ((g583) & (g584) & (!g587) & (!g586) & (!g593) & (g588)) + ((g583) & (g584) & (!g587) & (!g586) & (g593) & (g588)) + ((g583) & (g584) & (!g587) & (g586) & (!g593) & (g588)) + ((g583) & (g584) & (!g587) & (g586) & (g593) & (!g588)) + ((g583) & (g584) & (g587) & (!g586) & (!g593) & (g588)) + ((g583) & (g584) & (g587) & (!g586) & (g593) & (!g588)) + ((g583) & (g584) & (g587) & (g586) & (!g593) & (!g588)) + ((g583) & (g584) & (g587) & (g586) & (g593) & (!g588)) + ((g583) & (g584) & (g587) & (g586) & (g593) & (g588)));
	assign g629 = (((!g583) & (!g584) & (!g587) & (!g586) & (g593) & (!g588)) + ((!g583) & (!g584) & (!g587) & (g586) & (!g593) & (!g588)) + ((!g583) & (!g584) & (!g587) & (g586) & (g593) & (g588)) + ((!g583) & (!g584) & (g587) & (!g586) & (!g593) & (g588)) + ((!g583) & (!g584) & (g587) & (!g586) & (g593) & (g588)) + ((!g583) & (!g584) & (g587) & (g586) & (g593) & (g588)) + ((!g583) & (g584) & (!g587) & (!g586) & (!g593) & (g588)) + ((!g583) & (g584) & (!g587) & (g586) & (!g593) & (g588)) + ((!g583) & (g584) & (!g587) & (g586) & (g593) & (g588)) + ((!g583) & (g584) & (g587) & (!g586) & (!g593) & (!g588)) + ((!g583) & (g584) & (g587) & (!g586) & (g593) & (!g588)) + ((!g583) & (g584) & (g587) & (g586) & (!g593) & (g588)) + ((!g583) & (g584) & (g587) & (g586) & (g593) & (g588)) + ((g583) & (!g584) & (!g587) & (!g586) & (g593) & (!g588)) + ((g583) & (!g584) & (!g587) & (g586) & (g593) & (g588)) + ((g583) & (!g584) & (g587) & (!g586) & (!g593) & (!g588)) + ((g583) & (!g584) & (g587) & (!g586) & (g593) & (g588)) + ((g583) & (!g584) & (g587) & (g586) & (!g593) & (!g588)) + ((g583) & (g584) & (!g587) & (!g586) & (g593) & (g588)) + ((g583) & (g584) & (!g587) & (g586) & (!g593) & (!g588)) + ((g583) & (g584) & (!g587) & (g586) & (!g593) & (g588)) + ((g583) & (g584) & (g587) & (!g586) & (g593) & (g588)));
	assign g630 = (((!g626) & (!g627) & (!g628) & (!g629) & (!g594) & (!g585)) + ((!g626) & (!g627) & (!g628) & (!g629) & (!g594) & (g585)) + ((!g626) & (!g627) & (!g628) & (!g629) & (g594) & (!g585)) + ((!g626) & (!g627) & (!g628) & (g629) & (!g594) & (!g585)) + ((!g626) & (!g627) & (!g628) & (g629) & (!g594) & (g585)) + ((!g626) & (!g627) & (!g628) & (g629) & (g594) & (!g585)) + ((!g626) & (!g627) & (!g628) & (g629) & (g594) & (g585)) + ((!g626) & (!g627) & (g628) & (!g629) & (!g594) & (!g585)) + ((!g626) & (!g627) & (g628) & (!g629) & (g594) & (!g585)) + ((!g626) & (!g627) & (g628) & (g629) & (!g594) & (!g585)) + ((!g626) & (!g627) & (g628) & (g629) & (g594) & (!g585)) + ((!g626) & (!g627) & (g628) & (g629) & (g594) & (g585)) + ((!g626) & (g627) & (!g628) & (!g629) & (!g594) & (!g585)) + ((!g626) & (g627) & (!g628) & (!g629) & (!g594) & (g585)) + ((!g626) & (g627) & (!g628) & (g629) & (!g594) & (!g585)) + ((!g626) & (g627) & (!g628) & (g629) & (!g594) & (g585)) + ((!g626) & (g627) & (!g628) & (g629) & (g594) & (g585)) + ((!g626) & (g627) & (g628) & (!g629) & (!g594) & (!g585)) + ((!g626) & (g627) & (g628) & (g629) & (!g594) & (!g585)) + ((!g626) & (g627) & (g628) & (g629) & (g594) & (g585)) + ((g626) & (!g627) & (!g628) & (!g629) & (!g594) & (g585)) + ((g626) & (!g627) & (!g628) & (!g629) & (g594) & (!g585)) + ((g626) & (!g627) & (!g628) & (g629) & (!g594) & (g585)) + ((g626) & (!g627) & (!g628) & (g629) & (g594) & (!g585)) + ((g626) & (!g627) & (!g628) & (g629) & (g594) & (g585)) + ((g626) & (!g627) & (g628) & (!g629) & (g594) & (!g585)) + ((g626) & (!g627) & (g628) & (g629) & (g594) & (!g585)) + ((g626) & (!g627) & (g628) & (g629) & (g594) & (g585)) + ((g626) & (g627) & (!g628) & (!g629) & (!g594) & (g585)) + ((g626) & (g627) & (!g628) & (g629) & (!g594) & (g585)) + ((g626) & (g627) & (!g628) & (g629) & (g594) & (g585)) + ((g626) & (g627) & (g628) & (g629) & (g594) & (g585)));
	assign g632 = (((!sk[116]) & (g630) & (!g631)) + ((!sk[116]) & (g630) & (g631)) + ((sk[116]) & (!g630) & (g631)) + ((sk[116]) & (g630) & (!g631)));
	assign g633 = (((!g583) & (!g594) & (!g585) & (!g586) & (!g593) & (g588)) + ((!g583) & (!g594) & (!g585) & (!g586) & (g593) & (g588)) + ((!g583) & (!g594) & (!g585) & (g586) & (!g593) & (!g588)) + ((!g583) & (!g594) & (!g585) & (g586) & (!g593) & (g588)) + ((!g583) & (!g594) & (!g585) & (g586) & (g593) & (!g588)) + ((!g583) & (!g594) & (!g585) & (g586) & (g593) & (g588)) + ((!g583) & (!g594) & (g585) & (!g586) & (!g593) & (g588)) + ((!g583) & (!g594) & (g585) & (!g586) & (g593) & (g588)) + ((!g583) & (!g594) & (g585) & (g586) & (g593) & (!g588)) + ((!g583) & (g594) & (g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (g594) & (g585) & (!g586) & (g593) & (g588)) + ((!g583) & (g594) & (g585) & (g586) & (!g593) & (g588)) + ((g583) & (!g594) & (!g585) & (!g586) & (g593) & (!g588)) + ((g583) & (!g594) & (!g585) & (g586) & (!g593) & (!g588)) + ((g583) & (!g594) & (!g585) & (g586) & (!g593) & (g588)) + ((g583) & (!g594) & (!g585) & (g586) & (g593) & (g588)) + ((g583) & (!g594) & (g585) & (!g586) & (!g593) & (g588)) + ((g583) & (!g594) & (g585) & (!g586) & (g593) & (g588)) + ((g583) & (!g594) & (g585) & (g586) & (g593) & (!g588)) + ((g583) & (!g594) & (g585) & (g586) & (g593) & (g588)) + ((g583) & (g594) & (!g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (g594) & (!g585) & (!g586) & (!g593) & (g588)) + ((g583) & (g594) & (!g585) & (!g586) & (g593) & (!g588)) + ((g583) & (g594) & (!g585) & (g586) & (!g593) & (!g588)) + ((g583) & (g594) & (g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (g594) & (g585) & (!g586) & (!g593) & (g588)) + ((g583) & (g594) & (g585) & (!g586) & (g593) & (!g588)) + ((g583) & (g594) & (g585) & (g586) & (!g593) & (g588)));
	assign g634 = (((!g583) & (!g594) & (!g585) & (!g586) & (!g593) & (!g588)) + ((!g583) & (!g594) & (!g585) & (g586) & (g593) & (g588)) + ((!g583) & (!g594) & (g585) & (!g586) & (!g593) & (!g588)) + ((!g583) & (!g594) & (g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (!g594) & (g585) & (!g586) & (g593) & (g588)) + ((!g583) & (!g594) & (g585) & (g586) & (!g593) & (!g588)) + ((!g583) & (!g594) & (g585) & (g586) & (g593) & (g588)) + ((!g583) & (g594) & (!g585) & (!g586) & (!g593) & (!g588)) + ((!g583) & (g594) & (!g585) & (!g586) & (g593) & (g588)) + ((!g583) & (g594) & (!g585) & (g586) & (!g593) & (g588)) + ((!g583) & (g594) & (g585) & (!g586) & (!g593) & (!g588)) + ((!g583) & (g594) & (g585) & (!g586) & (g593) & (g588)) + ((!g583) & (g594) & (g585) & (g586) & (g593) & (!g588)) + ((!g583) & (g594) & (g585) & (g586) & (g593) & (g588)) + ((g583) & (!g594) & (!g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (!g594) & (!g585) & (!g586) & (g593) & (g588)) + ((g583) & (!g594) & (!g585) & (g586) & (!g593) & (!g588)) + ((g583) & (!g594) & (!g585) & (g586) & (g593) & (g588)) + ((g583) & (!g594) & (g585) & (!g586) & (g593) & (g588)) + ((g583) & (!g594) & (g585) & (g586) & (!g593) & (g588)) + ((g583) & (g594) & (!g585) & (!g586) & (g593) & (!g588)) + ((g583) & (g594) & (!g585) & (!g586) & (g593) & (g588)) + ((g583) & (g594) & (!g585) & (g586) & (!g593) & (g588)) + ((g583) & (g594) & (!g585) & (g586) & (g593) & (!g588)) + ((g583) & (g594) & (!g585) & (g586) & (g593) & (g588)) + ((g583) & (g594) & (g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (g594) & (g585) & (!g586) & (g593) & (!g588)) + ((g583) & (g594) & (g585) & (g586) & (!g593) & (!g588)));
	assign g635 = (((!g583) & (!g594) & (!g585) & (!g586) & (!g593) & (g588)) + ((!g583) & (!g594) & (!g585) & (!g586) & (g593) & (g588)) + ((!g583) & (!g594) & (!g585) & (g586) & (g593) & (!g588)) + ((!g583) & (!g594) & (!g585) & (g586) & (g593) & (g588)) + ((!g583) & (!g594) & (g585) & (!g586) & (g593) & (g588)) + ((!g583) & (!g594) & (g585) & (g586) & (!g593) & (!g588)) + ((!g583) & (!g594) & (g585) & (g586) & (!g593) & (g588)) + ((!g583) & (!g594) & (g585) & (g586) & (g593) & (g588)) + ((!g583) & (g594) & (!g585) & (!g586) & (!g593) & (!g588)) + ((!g583) & (g594) & (!g585) & (!g586) & (!g593) & (g588)) + ((!g583) & (g594) & (!g585) & (!g586) & (g593) & (g588)) + ((!g583) & (g594) & (!g585) & (g586) & (!g593) & (g588)) + ((!g583) & (g594) & (!g585) & (g586) & (g593) & (!g588)) + ((!g583) & (g594) & (g585) & (!g586) & (!g593) & (g588)) + ((!g583) & (g594) & (g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (g594) & (g585) & (g586) & (!g593) & (!g588)) + ((!g583) & (g594) & (g585) & (g586) & (g593) & (!g588)) + ((!g583) & (g594) & (g585) & (g586) & (g593) & (g588)) + ((g583) & (!g594) & (!g585) & (!g586) & (!g593) & (g588)) + ((g583) & (!g594) & (!g585) & (g586) & (!g593) & (!g588)) + ((g583) & (!g594) & (!g585) & (g586) & (g593) & (!g588)) + ((g583) & (!g594) & (g585) & (!g586) & (g593) & (g588)) + ((g583) & (!g594) & (g585) & (g586) & (!g593) & (g588)) + ((g583) & (g594) & (!g585) & (!g586) & (!g593) & (g588)) + ((g583) & (g594) & (!g585) & (g586) & (!g593) & (!g588)) + ((g583) & (g594) & (!g585) & (g586) & (g593) & (!g588)) + ((g583) & (g594) & (g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (g594) & (g585) & (!g586) & (g593) & (!g588)) + ((g583) & (g594) & (g585) & (!g586) & (g593) & (g588)) + ((g583) & (g594) & (g585) & (g586) & (g593) & (g588)));
	assign g636 = (((!g583) & (!g594) & (!g585) & (!g586) & (g593) & (g588)) + ((!g583) & (!g594) & (!g585) & (g586) & (!g593) & (!g588)) + ((!g583) & (!g594) & (!g585) & (g586) & (g593) & (g588)) + ((!g583) & (!g594) & (g585) & (!g586) & (!g593) & (!g588)) + ((!g583) & (!g594) & (g585) & (g586) & (g593) & (!g588)) + ((!g583) & (!g594) & (g585) & (g586) & (g593) & (g588)) + ((!g583) & (g594) & (!g585) & (g586) & (!g593) & (!g588)) + ((!g583) & (g594) & (!g585) & (g586) & (g593) & (!g588)) + ((!g583) & (g594) & (g585) & (!g586) & (g593) & (!g588)) + ((!g583) & (g594) & (g585) & (!g586) & (g593) & (g588)) + ((g583) & (!g594) & (!g585) & (!g586) & (!g593) & (g588)) + ((g583) & (!g594) & (!g585) & (!g586) & (g593) & (!g588)) + ((g583) & (!g594) & (!g585) & (g586) & (!g593) & (g588)) + ((g583) & (!g594) & (g585) & (!g586) & (g593) & (!g588)) + ((g583) & (!g594) & (g585) & (!g586) & (g593) & (g588)) + ((g583) & (!g594) & (g585) & (g586) & (g593) & (!g588)) + ((g583) & (!g594) & (g585) & (g586) & (g593) & (g588)) + ((g583) & (g594) & (!g585) & (!g586) & (g593) & (!g588)) + ((g583) & (g594) & (!g585) & (g586) & (!g593) & (g588)) + ((g583) & (g594) & (g585) & (!g586) & (!g593) & (!g588)) + ((g583) & (g594) & (g585) & (!g586) & (g593) & (g588)) + ((g583) & (g594) & (g585) & (g586) & (!g593) & (g588)));
	assign g637 = (((!g633) & (!g634) & (!g635) & (!g636) & (!g587) & (!g584)) + ((!g633) & (!g634) & (!g635) & (!g636) & (!g587) & (g584)) + ((!g633) & (!g634) & (!g635) & (!g636) & (g587) & (!g584)) + ((!g633) & (!g634) & (!g635) & (g636) & (!g587) & (!g584)) + ((!g633) & (!g634) & (!g635) & (g636) & (!g587) & (g584)) + ((!g633) & (!g634) & (!g635) & (g636) & (g587) & (!g584)) + ((!g633) & (!g634) & (!g635) & (g636) & (g587) & (g584)) + ((!g633) & (!g634) & (g635) & (!g636) & (!g587) & (!g584)) + ((!g633) & (!g634) & (g635) & (!g636) & (g587) & (!g584)) + ((!g633) & (!g634) & (g635) & (g636) & (!g587) & (!g584)) + ((!g633) & (!g634) & (g635) & (g636) & (g587) & (!g584)) + ((!g633) & (!g634) & (g635) & (g636) & (g587) & (g584)) + ((!g633) & (g634) & (!g635) & (!g636) & (!g587) & (!g584)) + ((!g633) & (g634) & (!g635) & (!g636) & (!g587) & (g584)) + ((!g633) & (g634) & (!g635) & (g636) & (!g587) & (!g584)) + ((!g633) & (g634) & (!g635) & (g636) & (!g587) & (g584)) + ((!g633) & (g634) & (!g635) & (g636) & (g587) & (g584)) + ((!g633) & (g634) & (g635) & (!g636) & (!g587) & (!g584)) + ((!g633) & (g634) & (g635) & (g636) & (!g587) & (!g584)) + ((!g633) & (g634) & (g635) & (g636) & (g587) & (g584)) + ((g633) & (!g634) & (!g635) & (!g636) & (!g587) & (g584)) + ((g633) & (!g634) & (!g635) & (!g636) & (g587) & (!g584)) + ((g633) & (!g634) & (!g635) & (g636) & (!g587) & (g584)) + ((g633) & (!g634) & (!g635) & (g636) & (g587) & (!g584)) + ((g633) & (!g634) & (!g635) & (g636) & (g587) & (g584)) + ((g633) & (!g634) & (g635) & (!g636) & (g587) & (!g584)) + ((g633) & (!g634) & (g635) & (g636) & (g587) & (!g584)) + ((g633) & (!g634) & (g635) & (g636) & (g587) & (g584)) + ((g633) & (g634) & (!g635) & (!g636) & (!g587) & (g584)) + ((g633) & (g634) & (!g635) & (g636) & (!g587) & (g584)) + ((g633) & (g634) & (!g635) & (g636) & (g587) & (g584)) + ((g633) & (g634) & (g635) & (g636) & (g587) & (g584)));
	assign g639 = (((!g637) & (sk[122]) & (g638)) + ((g637) & (!sk[122]) & (!g638)) + ((g637) & (!sk[122]) & (g638)) + ((g637) & (sk[122]) & (!g638)));
	assign g640 = (((!g587) & (!g584) & (!g585) & (!g586) & (!g593) & (g594)) + ((!g587) & (!g584) & (!g585) & (!g586) & (g593) & (!g594)) + ((!g587) & (!g584) & (!g585) & (g586) & (!g593) & (g594)) + ((!g587) & (!g584) & (!g585) & (g586) & (g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (!g586) & (!g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (!g586) & (g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (g586) & (!g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (g586) & (g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (g586) & (g593) & (g594)) + ((!g587) & (g584) & (!g585) & (!g586) & (g593) & (!g594)) + ((!g587) & (g584) & (!g585) & (g586) & (g593) & (!g594)) + ((!g587) & (g584) & (!g585) & (g586) & (g593) & (g594)) + ((!g587) & (g584) & (g585) & (!g586) & (g593) & (g594)) + ((!g587) & (g584) & (g585) & (g586) & (!g593) & (!g594)) + ((g587) & (!g584) & (!g585) & (!g586) & (!g593) & (g594)) + ((g587) & (!g584) & (!g585) & (g586) & (!g593) & (g594)) + ((g587) & (!g584) & (g585) & (g586) & (g593) & (g594)) + ((g587) & (g584) & (!g585) & (!g586) & (g593) & (g594)) + ((g587) & (g584) & (!g585) & (g586) & (!g593) & (!g594)) + ((g587) & (g584) & (!g585) & (g586) & (g593) & (!g594)) + ((g587) & (g584) & (g585) & (!g586) & (!g593) & (g594)) + ((g587) & (g584) & (g585) & (!g586) & (g593) & (!g594)) + ((g587) & (g584) & (g585) & (!g586) & (g593) & (g594)) + ((g587) & (g584) & (g585) & (g586) & (!g593) & (g594)));
	assign g641 = (((!g587) & (!g584) & (!g585) & (!g586) & (!g593) & (!g594)) + ((!g587) & (!g584) & (!g585) & (!g586) & (!g593) & (g594)) + ((!g587) & (!g584) & (!g585) & (g586) & (!g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (!g586) & (!g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (!g586) & (g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (!g586) & (g593) & (g594)) + ((!g587) & (!g584) & (g585) & (g586) & (!g593) & (g594)) + ((!g587) & (!g584) & (g585) & (g586) & (g593) & (g594)) + ((!g587) & (g584) & (!g585) & (!g586) & (!g593) & (!g594)) + ((!g587) & (g584) & (!g585) & (!g586) & (g593) & (!g594)) + ((!g587) & (g584) & (!g585) & (g586) & (!g593) & (!g594)) + ((!g587) & (g584) & (!g585) & (g586) & (!g593) & (g594)) + ((!g587) & (g584) & (!g585) & (g586) & (g593) & (g594)) + ((!g587) & (g584) & (g585) & (!g586) & (!g593) & (g594)) + ((!g587) & (g584) & (g585) & (g586) & (!g593) & (!g594)) + ((!g587) & (g584) & (g585) & (g586) & (!g593) & (g594)) + ((g587) & (!g584) & (!g585) & (!g586) & (!g593) & (g594)) + ((g587) & (!g584) & (!g585) & (!g586) & (g593) & (g594)) + ((g587) & (!g584) & (!g585) & (g586) & (!g593) & (!g594)) + ((g587) & (!g584) & (!g585) & (g586) & (g593) & (g594)) + ((g587) & (!g584) & (g585) & (!g586) & (!g593) & (!g594)) + ((g587) & (!g584) & (g585) & (!g586) & (g593) & (g594)) + ((g587) & (!g584) & (g585) & (g586) & (g593) & (!g594)) + ((g587) & (g584) & (!g585) & (!g586) & (!g593) & (!g594)) + ((g587) & (g584) & (!g585) & (!g586) & (!g593) & (g594)) + ((g587) & (g584) & (!g585) & (!g586) & (g593) & (g594)) + ((g587) & (g584) & (!g585) & (g586) & (!g593) & (g594)) + ((g587) & (g584) & (!g585) & (g586) & (g593) & (!g594)) + ((g587) & (g584) & (g585) & (!g586) & (g593) & (!g594)) + ((g587) & (g584) & (g585) & (!g586) & (g593) & (g594)));
	assign g642 = (((!g587) & (!g584) & (!g585) & (!g586) & (g593) & (!g594)) + ((!g587) & (!g584) & (!g585) & (g586) & (!g593) & (!g594)) + ((!g587) & (!g584) & (!g585) & (g586) & (g593) & (!g594)) + ((!g587) & (!g584) & (!g585) & (g586) & (g593) & (g594)) + ((!g587) & (!g584) & (g585) & (!g586) & (!g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (!g586) & (!g593) & (g594)) + ((!g587) & (!g584) & (g585) & (!g586) & (g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (g586) & (!g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (g586) & (g593) & (g594)) + ((!g587) & (g584) & (!g585) & (!g586) & (!g593) & (g594)) + ((!g587) & (g584) & (!g585) & (!g586) & (g593) & (!g594)) + ((!g587) & (g584) & (!g585) & (!g586) & (g593) & (g594)) + ((!g587) & (g584) & (g585) & (!g586) & (!g593) & (g594)) + ((!g587) & (g584) & (g585) & (!g586) & (g593) & (!g594)) + ((!g587) & (g584) & (g585) & (!g586) & (g593) & (g594)) + ((!g587) & (g584) & (g585) & (g586) & (!g593) & (!g594)) + ((g587) & (!g584) & (!g585) & (!g586) & (g593) & (!g594)) + ((g587) & (!g584) & (!g585) & (g586) & (!g593) & (!g594)) + ((g587) & (!g584) & (!g585) & (g586) & (g593) & (g594)) + ((g587) & (!g584) & (g585) & (!g586) & (!g593) & (!g594)) + ((g587) & (!g584) & (g585) & (!g586) & (!g593) & (g594)) + ((g587) & (!g584) & (g585) & (g586) & (!g593) & (!g594)) + ((g587) & (!g584) & (g585) & (g586) & (g593) & (!g594)) + ((g587) & (g584) & (!g585) & (!g586) & (g593) & (!g594)) + ((g587) & (g584) & (!g585) & (g586) & (!g593) & (!g594)) + ((g587) & (g584) & (!g585) & (g586) & (g593) & (g594)) + ((g587) & (g584) & (g585) & (!g586) & (!g593) & (!g594)) + ((g587) & (g584) & (g585) & (!g586) & (g593) & (!g594)) + ((g587) & (g584) & (g585) & (!g586) & (g593) & (g594)) + ((g587) & (g584) & (g585) & (g586) & (!g593) & (g594)));
	assign g643 = (((!g587) & (!g584) & (!g585) & (!g586) & (!g593) & (g594)) + ((!g587) & (!g584) & (!g585) & (g586) & (g593) & (!g594)) + ((!g587) & (!g584) & (!g585) & (g586) & (g593) & (g594)) + ((!g587) & (!g584) & (g585) & (!g586) & (!g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (!g586) & (!g593) & (g594)) + ((!g587) & (!g584) & (g585) & (g586) & (g593) & (!g594)) + ((!g587) & (!g584) & (g585) & (g586) & (g593) & (g594)) + ((!g587) & (g584) & (!g585) & (!g586) & (!g593) & (!g594)) + ((!g587) & (g584) & (!g585) & (!g586) & (!g593) & (g594)) + ((!g587) & (g584) & (!g585) & (!g586) & (g593) & (g594)) + ((!g587) & (g584) & (!g585) & (g586) & (!g593) & (g594)) + ((!g587) & (g584) & (g585) & (!g586) & (!g593) & (g594)) + ((!g587) & (g584) & (g585) & (g586) & (!g593) & (!g594)) + ((!g587) & (g584) & (g585) & (g586) & (!g593) & (g594)) + ((!g587) & (g584) & (g585) & (g586) & (g593) & (!g594)) + ((!g587) & (g584) & (g585) & (g586) & (g593) & (g594)) + ((g587) & (!g584) & (!g585) & (g586) & (!g593) & (g594)) + ((g587) & (!g584) & (g585) & (!g586) & (!g593) & (!g594)) + ((g587) & (!g584) & (g585) & (g586) & (!g593) & (!g594)) + ((g587) & (!g584) & (g585) & (g586) & (!g593) & (g594)) + ((g587) & (!g584) & (g585) & (g586) & (g593) & (g594)) + ((g587) & (g584) & (!g585) & (!g586) & (!g593) & (g594)) + ((g587) & (g584) & (!g585) & (!g586) & (g593) & (g594)) + ((g587) & (g584) & (!g585) & (g586) & (!g593) & (!g594)) + ((g587) & (g584) & (!g585) & (g586) & (g593) & (!g594)) + ((g587) & (g584) & (!g585) & (g586) & (g593) & (g594)) + ((g587) & (g584) & (g585) & (!g586) & (g593) & (g594)) + ((g587) & (g584) & (g585) & (g586) & (g593) & (g594)));
	assign g644 = (((!g640) & (!g641) & (!g642) & (!g643) & (!g583) & (g588)) + ((!g640) & (!g641) & (!g642) & (!g643) & (g583) & (!g588)) + ((!g640) & (!g641) & (!g642) & (!g643) & (g583) & (g588)) + ((!g640) & (!g641) & (!g642) & (g643) & (!g583) & (g588)) + ((!g640) & (!g641) & (!g642) & (g643) & (g583) & (!g588)) + ((!g640) & (!g641) & (g642) & (!g643) & (g583) & (!g588)) + ((!g640) & (!g641) & (g642) & (!g643) & (g583) & (g588)) + ((!g640) & (!g641) & (g642) & (g643) & (g583) & (!g588)) + ((!g640) & (g641) & (!g642) & (!g643) & (!g583) & (g588)) + ((!g640) & (g641) & (!g642) & (!g643) & (g583) & (g588)) + ((!g640) & (g641) & (!g642) & (g643) & (!g583) & (g588)) + ((!g640) & (g641) & (g642) & (!g643) & (g583) & (g588)) + ((g640) & (!g641) & (!g642) & (!g643) & (!g583) & (!g588)) + ((g640) & (!g641) & (!g642) & (!g643) & (!g583) & (g588)) + ((g640) & (!g641) & (!g642) & (!g643) & (g583) & (!g588)) + ((g640) & (!g641) & (!g642) & (!g643) & (g583) & (g588)) + ((g640) & (!g641) & (!g642) & (g643) & (!g583) & (!g588)) + ((g640) & (!g641) & (!g642) & (g643) & (!g583) & (g588)) + ((g640) & (!g641) & (!g642) & (g643) & (g583) & (!g588)) + ((g640) & (!g641) & (g642) & (!g643) & (!g583) & (!g588)) + ((g640) & (!g641) & (g642) & (!g643) & (g583) & (!g588)) + ((g640) & (!g641) & (g642) & (!g643) & (g583) & (g588)) + ((g640) & (!g641) & (g642) & (g643) & (!g583) & (!g588)) + ((g640) & (!g641) & (g642) & (g643) & (g583) & (!g588)) + ((g640) & (g641) & (!g642) & (!g643) & (!g583) & (!g588)) + ((g640) & (g641) & (!g642) & (!g643) & (!g583) & (g588)) + ((g640) & (g641) & (!g642) & (!g643) & (g583) & (g588)) + ((g640) & (g641) & (!g642) & (g643) & (!g583) & (!g588)) + ((g640) & (g641) & (!g642) & (g643) & (!g583) & (g588)) + ((g640) & (g641) & (g642) & (!g643) & (!g583) & (!g588)) + ((g640) & (g641) & (g642) & (!g643) & (g583) & (g588)) + ((g640) & (g641) & (g642) & (g643) & (!g583) & (!g588)));
	assign g646 = (((!g644) & (sk[0]) & (g645)) + ((g644) & (!sk[0]) & (!g645)) + ((g644) & (!sk[0]) & (g645)) + ((g644) & (sk[0]) & (!g645)));
	assign g653 = (((!g647) & (!g648) & (!g649) & (!g650) & (g651) & (g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g651) & (!g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g651) & (g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (g651) & (!g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (!g651) & (!g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (!g651) & (g652)) + ((!g647) & (!g648) & (g649) & (g650) & (!g651) & (!g652)) + ((!g647) & (!g648) & (g649) & (g650) & (g651) & (g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (g651) & (!g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (g651) & (g652)) + ((!g647) & (g648) & (!g649) & (g650) & (g651) & (!g652)) + ((!g647) & (g648) & (!g649) & (g650) & (g651) & (g652)) + ((!g647) & (g648) & (g649) & (!g650) & (g651) & (!g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (!g651) & (!g652)) + ((g647) & (!g648) & (g649) & (!g650) & (g651) & (!g652)) + ((g647) & (!g648) & (g649) & (g650) & (!g651) & (g652)) + ((g647) & (!g648) & (g649) & (g650) & (g651) & (g652)) + ((g647) & (g648) & (!g649) & (!g650) & (!g651) & (g652)) + ((g647) & (g648) & (!g649) & (!g650) & (g651) & (!g652)) + ((g647) & (g648) & (g649) & (!g650) & (!g651) & (g652)) + ((g647) & (g648) & (g649) & (!g650) & (g651) & (!g652)) + ((g647) & (g648) & (g649) & (g650) & (!g651) & (!g652)) + ((g647) & (g648) & (g649) & (g650) & (g651) & (!g652)) + ((g647) & (g648) & (g649) & (g650) & (g651) & (g652)));
	assign g654 = (((!g647) & (!g648) & (!g649) & (!g650) & (g651) & (!g652)) + ((!g647) & (!g648) & (!g649) & (!g650) & (g651) & (g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g651) & (!g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g651) & (g652)) + ((!g647) & (!g648) & (g649) & (g650) & (!g651) & (g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (!g651) & (!g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (!g651) & (g652)) + ((!g647) & (g648) & (g649) & (!g650) & (!g651) & (!g652)) + ((!g647) & (g648) & (g649) & (!g650) & (!g651) & (g652)) + ((!g647) & (g648) & (g649) & (!g650) & (g651) & (!g652)) + ((!g647) & (g648) & (g649) & (g650) & (g651) & (g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (!g651) & (g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (g651) & (!g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (g651) & (g652)) + ((g647) & (!g648) & (!g649) & (g650) & (g651) & (!g652)) + ((g647) & (!g648) & (g649) & (!g650) & (!g651) & (!g652)) + ((g647) & (!g648) & (g649) & (!g650) & (g651) & (g652)) + ((g647) & (!g648) & (g649) & (g650) & (!g651) & (g652)) + ((g647) & (!g648) & (g649) & (g650) & (g651) & (g652)) + ((g647) & (g648) & (!g649) & (!g650) & (!g651) & (!g652)) + ((g647) & (g648) & (!g649) & (!g650) & (!g651) & (g652)) + ((g647) & (g648) & (!g649) & (!g650) & (g651) & (!g652)) + ((g647) & (g648) & (!g649) & (!g650) & (g651) & (g652)) + ((g647) & (g648) & (!g649) & (g650) & (!g651) & (!g652)) + ((g647) & (g648) & (!g649) & (g650) & (g651) & (!g652)) + ((g647) & (g648) & (!g649) & (g650) & (g651) & (g652)) + ((g647) & (g648) & (g649) & (!g650) & (g651) & (!g652)) + ((g647) & (g648) & (g649) & (!g650) & (g651) & (g652)) + ((g647) & (g648) & (g649) & (g650) & (!g651) & (g652)) + ((g647) & (g648) & (g649) & (g650) & (g651) & (!g652)));
	assign g655 = (((!g647) & (!g648) & (!g649) & (!g650) & (!g651) & (!g652)) + ((!g647) & (!g648) & (!g649) & (!g650) & (g651) & (g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (g651) & (g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (!g651) & (!g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (!g651) & (g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (g651) & (g652)) + ((!g647) & (!g648) & (g649) & (g650) & (!g651) & (g652)) + ((!g647) & (!g648) & (g649) & (g650) & (g651) & (!g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (!g651) & (!g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (g651) & (!g652)) + ((!g647) & (g648) & (!g649) & (g650) & (g651) & (g652)) + ((!g647) & (g648) & (g649) & (g650) & (!g651) & (!g652)) + ((!g647) & (g648) & (g649) & (g650) & (g651) & (!g652)) + ((g647) & (!g648) & (!g649) & (g650) & (!g651) & (!g652)) + ((g647) & (!g648) & (!g649) & (g650) & (!g651) & (g652)) + ((g647) & (!g648) & (!g649) & (g650) & (g651) & (!g652)) + ((g647) & (!g648) & (g649) & (!g650) & (!g651) & (!g652)) + ((g647) & (!g648) & (g649) & (!g650) & (g651) & (g652)) + ((g647) & (!g648) & (g649) & (g650) & (!g651) & (!g652)) + ((g647) & (!g648) & (g649) & (g650) & (!g651) & (g652)) + ((g647) & (!g648) & (g649) & (g650) & (g651) & (!g652)) + ((g647) & (!g648) & (g649) & (g650) & (g651) & (g652)) + ((g647) & (g648) & (!g649) & (!g650) & (g651) & (g652)) + ((g647) & (g648) & (!g649) & (g650) & (!g651) & (!g652)) + ((g647) & (g648) & (!g649) & (g650) & (g651) & (!g652)) + ((g647) & (g648) & (!g649) & (g650) & (g651) & (g652)) + ((g647) & (g648) & (g649) & (!g650) & (!g651) & (!g652)) + ((g647) & (g648) & (g649) & (g650) & (!g651) & (!g652)) + ((g647) & (g648) & (g649) & (g650) & (!g651) & (g652)) + ((g647) & (g648) & (g649) & (g650) & (g651) & (g652)));
	assign g656 = (((!g647) & (!g648) & (!g649) & (!g650) & (!g651) & (g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (g651) & (!g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (g651) & (g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (!g651) & (g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (g651) & (g652)) + ((!g647) & (!g648) & (g649) & (g650) & (!g651) & (g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (!g651) & (!g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (!g651) & (g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (g651) & (!g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (g651) & (g652)) + ((!g647) & (g648) & (!g649) & (g650) & (g651) & (!g652)) + ((!g647) & (g648) & (!g649) & (g650) & (g651) & (g652)) + ((!g647) & (g648) & (g649) & (g650) & (!g651) & (!g652)) + ((!g647) & (g648) & (g649) & (g650) & (g651) & (!g652)) + ((!g647) & (g648) & (g649) & (g650) & (g651) & (g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (!g651) & (!g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (g651) & (g652)) + ((g647) & (!g648) & (!g649) & (g650) & (g651) & (!g652)) + ((g647) & (!g648) & (!g649) & (g650) & (g651) & (g652)) + ((g647) & (!g648) & (g649) & (!g650) & (!g651) & (g652)) + ((g647) & (!g648) & (g649) & (!g650) & (g651) & (!g652)) + ((g647) & (!g648) & (g649) & (g650) & (g651) & (!g652)) + ((g647) & (g648) & (!g649) & (!g650) & (!g651) & (g652)) + ((g647) & (g648) & (!g649) & (!g650) & (g651) & (g652)) + ((g647) & (g648) & (!g649) & (g650) & (g651) & (!g652)) + ((g647) & (g648) & (!g649) & (g650) & (g651) & (g652)) + ((g647) & (g648) & (g649) & (!g650) & (!g651) & (g652)) + ((g647) & (g648) & (g649) & (g650) & (!g651) & (!g652)));
	assign g659 = (((!g653) & (!g654) & (!g655) & (!g656) & (!g657) & (!g658)) + ((!g653) & (!g654) & (!g655) & (g656) & (!g657) & (!g658)) + ((!g653) & (!g654) & (!g655) & (g656) & (g657) & (g658)) + ((!g653) & (!g654) & (g655) & (!g656) & (!g657) & (!g658)) + ((!g653) & (!g654) & (g655) & (!g656) & (!g657) & (g658)) + ((!g653) & (!g654) & (g655) & (g656) & (!g657) & (!g658)) + ((!g653) & (!g654) & (g655) & (g656) & (!g657) & (g658)) + ((!g653) & (!g654) & (g655) & (g656) & (g657) & (g658)) + ((!g653) & (g654) & (!g655) & (!g656) & (!g657) & (!g658)) + ((!g653) & (g654) & (!g655) & (!g656) & (g657) & (!g658)) + ((!g653) & (g654) & (!g655) & (g656) & (!g657) & (!g658)) + ((!g653) & (g654) & (!g655) & (g656) & (g657) & (!g658)) + ((!g653) & (g654) & (!g655) & (g656) & (g657) & (g658)) + ((!g653) & (g654) & (g655) & (!g656) & (!g657) & (!g658)) + ((!g653) & (g654) & (g655) & (!g656) & (!g657) & (g658)) + ((!g653) & (g654) & (g655) & (!g656) & (g657) & (!g658)) + ((!g653) & (g654) & (g655) & (g656) & (!g657) & (!g658)) + ((!g653) & (g654) & (g655) & (g656) & (!g657) & (g658)) + ((!g653) & (g654) & (g655) & (g656) & (g657) & (!g658)) + ((!g653) & (g654) & (g655) & (g656) & (g657) & (g658)) + ((g653) & (!g654) & (!g655) & (g656) & (g657) & (g658)) + ((g653) & (!g654) & (g655) & (!g656) & (!g657) & (g658)) + ((g653) & (!g654) & (g655) & (g656) & (!g657) & (g658)) + ((g653) & (!g654) & (g655) & (g656) & (g657) & (g658)) + ((g653) & (g654) & (!g655) & (!g656) & (g657) & (!g658)) + ((g653) & (g654) & (!g655) & (g656) & (g657) & (!g658)) + ((g653) & (g654) & (!g655) & (g656) & (g657) & (g658)) + ((g653) & (g654) & (g655) & (!g656) & (!g657) & (g658)) + ((g653) & (g654) & (g655) & (!g656) & (g657) & (!g658)) + ((g653) & (g654) & (g655) & (g656) & (!g657) & (g658)) + ((g653) & (g654) & (g655) & (g656) & (g657) & (!g658)) + ((g653) & (g654) & (g655) & (g656) & (g657) & (g658)));
	assign g661 = (((!sk[6]) & (g659) & (!g660)) + ((!sk[6]) & (g659) & (g660)) + ((sk[6]) & (!g659) & (g660)) + ((sk[6]) & (g659) & (!g660)));
	assign g662 = (((!g647) & (!g648) & (!g649) & (!g650) & (!g657) & (g651)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g657) & (!g651)) + ((!g647) & (!g648) & (!g649) & (g650) & (g657) & (!g651)) + ((!g647) & (!g648) & (g649) & (!g650) & (g657) & (g651)) + ((!g647) & (!g648) & (g649) & (g650) & (!g657) & (g651)) + ((!g647) & (!g648) & (g649) & (g650) & (g657) & (!g651)) + ((!g647) & (g648) & (!g649) & (!g650) & (!g657) & (g651)) + ((!g647) & (g648) & (!g649) & (!g650) & (g657) & (!g651)) + ((!g647) & (g648) & (!g649) & (!g650) & (g657) & (g651)) + ((!g647) & (g648) & (g649) & (!g650) & (g657) & (g651)) + ((!g647) & (g648) & (g649) & (g650) & (g657) & (g651)) + ((g647) & (!g648) & (!g649) & (!g650) & (!g657) & (!g651)) + ((g647) & (!g648) & (!g649) & (!g650) & (g657) & (g651)) + ((g647) & (!g648) & (!g649) & (g650) & (!g657) & (!g651)) + ((g647) & (!g648) & (!g649) & (g650) & (g657) & (!g651)) + ((g647) & (!g648) & (g649) & (!g650) & (g657) & (!g651)) + ((g647) & (!g648) & (g649) & (!g650) & (g657) & (g651)) + ((g647) & (!g648) & (g649) & (g650) & (g657) & (!g651)) + ((g647) & (!g648) & (g649) & (g650) & (g657) & (g651)) + ((g647) & (g648) & (!g649) & (!g650) & (g657) & (!g651)) + ((g647) & (g648) & (!g649) & (!g650) & (g657) & (g651)) + ((g647) & (g648) & (!g649) & (g650) & (g657) & (g651)) + ((g647) & (g648) & (g649) & (!g650) & (!g657) & (!g651)) + ((g647) & (g648) & (g649) & (!g650) & (!g657) & (g651)) + ((g647) & (g648) & (g649) & (!g650) & (g657) & (!g651)) + ((g647) & (g648) & (g649) & (g650) & (!g657) & (g651)) + ((g647) & (g648) & (g649) & (g650) & (g657) & (!g651)));
	assign g663 = (((!g647) & (!g648) & (!g649) & (!g650) & (!g657) & (g651)) + ((!g647) & (!g648) & (!g649) & (!g650) & (g657) & (!g651)) + ((!g647) & (!g648) & (!g649) & (!g650) & (g657) & (g651)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g657) & (!g651)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g657) & (g651)) + ((!g647) & (!g648) & (!g649) & (g650) & (g657) & (g651)) + ((!g647) & (!g648) & (g649) & (!g650) & (g657) & (!g651)) + ((!g647) & (!g648) & (g649) & (g650) & (!g657) & (!g651)) + ((!g647) & (!g648) & (g649) & (g650) & (!g657) & (g651)) + ((!g647) & (!g648) & (g649) & (g650) & (g657) & (g651)) + ((!g647) & (g648) & (!g649) & (!g650) & (g657) & (g651)) + ((!g647) & (g648) & (!g649) & (g650) & (!g657) & (!g651)) + ((!g647) & (g648) & (!g649) & (g650) & (g657) & (!g651)) + ((!g647) & (g648) & (g649) & (!g650) & (g657) & (!g651)) + ((!g647) & (g648) & (g649) & (!g650) & (g657) & (g651)) + ((!g647) & (g648) & (g649) & (g650) & (!g657) & (!g651)) + ((g647) & (!g648) & (!g649) & (!g650) & (!g657) & (!g651)) + ((g647) & (!g648) & (!g649) & (g650) & (!g657) & (!g651)) + ((g647) & (!g648) & (!g649) & (g650) & (!g657) & (g651)) + ((g647) & (!g648) & (g649) & (!g650) & (!g657) & (g651)) + ((g647) & (!g648) & (g649) & (!g650) & (g657) & (g651)) + ((g647) & (!g648) & (g649) & (g650) & (!g657) & (!g651)) + ((g647) & (!g648) & (g649) & (g650) & (!g657) & (g651)) + ((g647) & (g648) & (!g649) & (g650) & (!g657) & (!g651)) + ((g647) & (g648) & (!g649) & (g650) & (g657) & (g651)) + ((g647) & (g648) & (g649) & (!g650) & (!g657) & (!g651)) + ((g647) & (g648) & (g649) & (!g650) & (!g657) & (g651)) + ((g647) & (g648) & (g649) & (!g650) & (g657) & (g651)) + ((g647) & (g648) & (g649) & (g650) & (!g657) & (!g651)) + ((g647) & (g648) & (g649) & (g650) & (!g657) & (g651)) + ((g647) & (g648) & (g649) & (g650) & (g657) & (!g651)));
	assign g664 = (((!g647) & (!g648) & (!g649) & (!g650) & (!g657) & (g651)) + ((!g647) & (!g648) & (!g649) & (g650) & (g657) & (!g651)) + ((!g647) & (!g648) & (g649) & (!g650) & (!g657) & (!g651)) + ((!g647) & (!g648) & (g649) & (!g650) & (g657) & (!g651)) + ((!g647) & (!g648) & (g649) & (g650) & (!g657) & (g651)) + ((!g647) & (!g648) & (g649) & (g650) & (g657) & (!g651)) + ((!g647) & (!g648) & (g649) & (g650) & (g657) & (g651)) + ((!g647) & (g648) & (!g649) & (!g650) & (!g657) & (!g651)) + ((!g647) & (g648) & (!g649) & (!g650) & (g657) & (!g651)) + ((!g647) & (g648) & (!g649) & (g650) & (!g657) & (!g651)) + ((!g647) & (g648) & (!g649) & (g650) & (g657) & (g651)) + ((!g647) & (g648) & (g649) & (!g650) & (g657) & (g651)) + ((!g647) & (g648) & (g649) & (g650) & (!g657) & (g651)) + ((!g647) & (g648) & (g649) & (g650) & (g657) & (!g651)) + ((g647) & (!g648) & (!g649) & (!g650) & (g657) & (g651)) + ((g647) & (!g648) & (!g649) & (g650) & (!g657) & (!g651)) + ((g647) & (!g648) & (!g649) & (g650) & (g657) & (!g651)) + ((g647) & (!g648) & (g649) & (!g650) & (!g657) & (!g651)) + ((g647) & (!g648) & (g649) & (!g650) & (!g657) & (g651)) + ((g647) & (!g648) & (g649) & (!g650) & (g657) & (!g651)) + ((g647) & (!g648) & (g649) & (!g650) & (g657) & (g651)) + ((g647) & (!g648) & (g649) & (g650) & (g657) & (!g651)) + ((g647) & (g648) & (!g649) & (!g650) & (!g657) & (g651)) + ((g647) & (g648) & (!g649) & (!g650) & (g657) & (g651)) + ((g647) & (g648) & (!g649) & (g650) & (!g657) & (g651)) + ((g647) & (g648) & (g649) & (!g650) & (!g657) & (!g651)) + ((g647) & (g648) & (g649) & (!g650) & (!g657) & (g651)) + ((g647) & (g648) & (g649) & (!g650) & (g657) & (g651)) + ((g647) & (g648) & (g649) & (g650) & (!g657) & (!g651)) + ((g647) & (g648) & (g649) & (g650) & (!g657) & (g651)) + ((g647) & (g648) & (g649) & (g650) & (g657) & (!g651)) + ((g647) & (g648) & (g649) & (g650) & (g657) & (g651)));
	assign g665 = (((!g647) & (!g648) & (!g649) & (!g650) & (g657) & (!g651)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g657) & (!g651)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g657) & (g651)) + ((!g647) & (!g648) & (g649) & (!g650) & (g657) & (g651)) + ((!g647) & (!g648) & (g649) & (g650) & (!g657) & (g651)) + ((!g647) & (g648) & (!g649) & (!g650) & (!g657) & (!g651)) + ((!g647) & (g648) & (!g649) & (!g650) & (g657) & (!g651)) + ((!g647) & (g648) & (!g649) & (g650) & (!g657) & (g651)) + ((!g647) & (g648) & (g649) & (!g650) & (!g657) & (g651)) + ((!g647) & (g648) & (g649) & (!g650) & (g657) & (!g651)) + ((!g647) & (g648) & (g649) & (!g650) & (g657) & (g651)) + ((!g647) & (g648) & (g649) & (g650) & (g657) & (!g651)) + ((!g647) & (g648) & (g649) & (g650) & (g657) & (g651)) + ((g647) & (!g648) & (!g649) & (!g650) & (!g657) & (!g651)) + ((g647) & (!g648) & (!g649) & (g650) & (!g657) & (!g651)) + ((g647) & (!g648) & (!g649) & (g650) & (!g657) & (g651)) + ((g647) & (!g648) & (!g649) & (g650) & (g657) & (!g651)) + ((g647) & (!g648) & (g649) & (!g650) & (!g657) & (!g651)) + ((g647) & (!g648) & (g649) & (!g650) & (g657) & (g651)) + ((g647) & (!g648) & (g649) & (g650) & (g657) & (!g651)) + ((g647) & (g648) & (!g649) & (!g650) & (!g657) & (!g651)) + ((g647) & (g648) & (!g649) & (g650) & (!g657) & (!g651)) + ((g647) & (g648) & (!g649) & (g650) & (g657) & (!g651)) + ((g647) & (g648) & (!g649) & (g650) & (g657) & (g651)) + ((g647) & (g648) & (g649) & (g650) & (!g657) & (g651)) + ((g647) & (g648) & (g649) & (g650) & (g657) & (g651)));
	assign g666 = (((!g662) & (!g663) & (!g664) & (!g665) & (!g652) & (!g658)) + ((!g662) & (!g663) & (!g664) & (!g665) & (g652) & (!g658)) + ((!g662) & (!g663) & (!g664) & (g665) & (!g652) & (!g658)) + ((!g662) & (!g663) & (!g664) & (g665) & (g652) & (!g658)) + ((!g662) & (!g663) & (!g664) & (g665) & (g652) & (g658)) + ((!g662) & (!g663) & (g664) & (!g665) & (!g652) & (!g658)) + ((!g662) & (!g663) & (g664) & (!g665) & (!g652) & (g658)) + ((!g662) & (!g663) & (g664) & (!g665) & (g652) & (!g658)) + ((!g662) & (!g663) & (g664) & (g665) & (!g652) & (!g658)) + ((!g662) & (!g663) & (g664) & (g665) & (!g652) & (g658)) + ((!g662) & (!g663) & (g664) & (g665) & (g652) & (!g658)) + ((!g662) & (!g663) & (g664) & (g665) & (g652) & (g658)) + ((!g662) & (g663) & (!g664) & (!g665) & (!g652) & (!g658)) + ((!g662) & (g663) & (!g664) & (g665) & (!g652) & (!g658)) + ((!g662) & (g663) & (!g664) & (g665) & (g652) & (g658)) + ((!g662) & (g663) & (g664) & (!g665) & (!g652) & (!g658)) + ((!g662) & (g663) & (g664) & (!g665) & (!g652) & (g658)) + ((!g662) & (g663) & (g664) & (g665) & (!g652) & (!g658)) + ((!g662) & (g663) & (g664) & (g665) & (!g652) & (g658)) + ((!g662) & (g663) & (g664) & (g665) & (g652) & (g658)) + ((g662) & (!g663) & (!g664) & (!g665) & (g652) & (!g658)) + ((g662) & (!g663) & (!g664) & (g665) & (g652) & (!g658)) + ((g662) & (!g663) & (!g664) & (g665) & (g652) & (g658)) + ((g662) & (!g663) & (g664) & (!g665) & (!g652) & (g658)) + ((g662) & (!g663) & (g664) & (!g665) & (g652) & (!g658)) + ((g662) & (!g663) & (g664) & (g665) & (!g652) & (g658)) + ((g662) & (!g663) & (g664) & (g665) & (g652) & (!g658)) + ((g662) & (!g663) & (g664) & (g665) & (g652) & (g658)) + ((g662) & (g663) & (!g664) & (g665) & (g652) & (g658)) + ((g662) & (g663) & (g664) & (!g665) & (!g652) & (g658)) + ((g662) & (g663) & (g664) & (g665) & (!g652) & (g658)) + ((g662) & (g663) & (g664) & (g665) & (g652) & (g658)));
	assign g668 = (((!g666) & (sk[12]) & (g667)) + ((g666) & (!sk[12]) & (!g667)) + ((g666) & (!sk[12]) & (g667)) + ((g666) & (sk[12]) & (!g667)));
	assign g669 = (((!g651) & (!g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((!g651) & (!g648) & (!g649) & (!g650) & (g657) & (g652)) + ((!g651) & (!g648) & (!g649) & (g650) & (!g657) & (g652)) + ((!g651) & (!g648) & (!g649) & (g650) & (g657) & (!g652)) + ((!g651) & (!g648) & (!g649) & (g650) & (g657) & (g652)) + ((!g651) & (!g648) & (g649) & (!g650) & (!g657) & (g652)) + ((!g651) & (!g648) & (g649) & (g650) & (!g657) & (!g652)) + ((!g651) & (!g648) & (g649) & (g650) & (g657) & (!g652)) + ((!g651) & (g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((!g651) & (g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((!g651) & (g648) & (!g649) & (g650) & (!g657) & (g652)) + ((!g651) & (g648) & (g649) & (!g650) & (!g657) & (!g652)) + ((!g651) & (g648) & (g649) & (!g650) & (!g657) & (g652)) + ((!g651) & (g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g651) & (g648) & (g649) & (!g650) & (g657) & (g652)) + ((g651) & (!g648) & (!g649) & (g650) & (!g657) & (g652)) + ((g651) & (!g648) & (!g649) & (g650) & (g657) & (g652)) + ((g651) & (g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((g651) & (g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((g651) & (g648) & (!g649) & (g650) & (g657) & (!g652)) + ((g651) & (g648) & (g649) & (g650) & (!g657) & (!g652)) + ((g651) & (g648) & (g649) & (g650) & (!g657) & (g652)));
	assign g670 = (((!g651) & (!g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((!g651) & (!g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((!g651) & (!g648) & (!g649) & (g650) & (g657) & (g652)) + ((!g651) & (!g648) & (g649) & (!g650) & (!g657) & (!g652)) + ((!g651) & (!g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g651) & (!g648) & (g649) & (g650) & (!g657) & (g652)) + ((!g651) & (g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((!g651) & (g648) & (!g649) & (!g650) & (g657) & (g652)) + ((!g651) & (g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((!g651) & (g648) & (!g649) & (g650) & (!g657) & (g652)) + ((!g651) & (g648) & (!g649) & (g650) & (g657) & (g652)) + ((!g651) & (g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g651) & (g648) & (g649) & (!g650) & (g657) & (g652)) + ((!g651) & (g648) & (g649) & (g650) & (g657) & (!g652)) + ((g651) & (!g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((g651) & (!g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((g651) & (!g648) & (!g649) & (!g650) & (g657) & (g652)) + ((g651) & (!g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((g651) & (!g648) & (!g649) & (g650) & (!g657) & (g652)) + ((g651) & (!g648) & (!g649) & (g650) & (g657) & (!g652)) + ((g651) & (!g648) & (g649) & (g650) & (!g657) & (!g652)) + ((g651) & (g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((g651) & (g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((g651) & (g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((g651) & (g648) & (!g649) & (g650) & (g657) & (!g652)) + ((g651) & (g648) & (!g649) & (g650) & (g657) & (g652)) + ((g651) & (g648) & (g649) & (!g650) & (!g657) & (!g652)) + ((g651) & (g648) & (g649) & (!g650) & (g657) & (!g652)) + ((g651) & (g648) & (g649) & (g650) & (!g657) & (g652)) + ((g651) & (g648) & (g649) & (g650) & (g657) & (g652)));
	assign g671 = (((!g651) & (!g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((!g651) & (!g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((!g651) & (!g648) & (!g649) & (g650) & (!g657) & (g652)) + ((!g651) & (!g648) & (g649) & (!g650) & (!g657) & (g652)) + ((!g651) & (!g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g651) & (!g648) & (g649) & (g650) & (!g657) & (g652)) + ((!g651) & (g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((!g651) & (g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((!g651) & (g648) & (!g649) & (g650) & (g657) & (!g652)) + ((!g651) & (g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g651) & (g648) & (g649) & (g650) & (!g657) & (!g652)) + ((!g651) & (g648) & (g649) & (g650) & (g657) & (!g652)) + ((g651) & (!g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((g651) & (!g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((g651) & (!g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((g651) & (!g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((g651) & (!g648) & (!g649) & (g650) & (!g657) & (g652)) + ((g651) & (!g648) & (!g649) & (g650) & (g657) & (!g652)) + ((g651) & (!g648) & (!g649) & (g650) & (g657) & (g652)) + ((g651) & (!g648) & (g649) & (!g650) & (!g657) & (g652)) + ((g651) & (!g648) & (g649) & (!g650) & (g657) & (!g652)) + ((g651) & (!g648) & (g649) & (g650) & (!g657) & (!g652)) + ((g651) & (!g648) & (g649) & (g650) & (g657) & (g652)) + ((g651) & (g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((g651) & (g648) & (!g649) & (!g650) & (g657) & (g652)) + ((g651) & (g648) & (g649) & (!g650) & (g657) & (g652)) + ((g651) & (g648) & (g649) & (g650) & (!g657) & (!g652)) + ((g651) & (g648) & (g649) & (g650) & (!g657) & (g652)) + ((g651) & (g648) & (g649) & (g650) & (g657) & (g652)));
	assign g672 = (((!g651) & (!g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((!g651) & (!g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((!g651) & (!g648) & (!g649) & (!g650) & (g657) & (g652)) + ((!g651) & (!g648) & (!g649) & (g650) & (!g657) & (g652)) + ((!g651) & (!g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g651) & (!g648) & (g649) & (g650) & (g657) & (g652)) + ((!g651) & (g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((!g651) & (g648) & (!g649) & (g650) & (!g657) & (g652)) + ((!g651) & (g648) & (!g649) & (g650) & (g657) & (g652)) + ((!g651) & (g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g651) & (g648) & (g649) & (!g650) & (g657) & (g652)) + ((!g651) & (g648) & (g649) & (g650) & (!g657) & (!g652)) + ((!g651) & (g648) & (g649) & (g650) & (!g657) & (g652)) + ((!g651) & (g648) & (g649) & (g650) & (g657) & (!g652)) + ((!g651) & (g648) & (g649) & (g650) & (g657) & (g652)) + ((g651) & (!g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((g651) & (!g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((g651) & (!g648) & (!g649) & (!g650) & (g657) & (g652)) + ((g651) & (!g648) & (!g649) & (g650) & (g657) & (g652)) + ((g651) & (!g648) & (g649) & (!g650) & (!g657) & (g652)) + ((g651) & (!g648) & (g649) & (!g650) & (g657) & (!g652)) + ((g651) & (!g648) & (g649) & (g650) & (g657) & (!g652)) + ((g651) & (g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((g651) & (g648) & (!g649) & (g650) & (!g657) & (g652)) + ((g651) & (g648) & (!g649) & (g650) & (g657) & (!g652)) + ((g651) & (g648) & (g649) & (!g650) & (g657) & (g652)) + ((g651) & (g648) & (g649) & (g650) & (!g657) & (!g652)));
	assign g673 = (((!g669) & (!g670) & (!g671) & (!g672) & (!g647) & (g658)) + ((!g669) & (!g670) & (!g671) & (!g672) & (g647) & (!g658)) + ((!g669) & (!g670) & (!g671) & (!g672) & (g647) & (g658)) + ((!g669) & (!g670) & (!g671) & (g672) & (!g647) & (g658)) + ((!g669) & (!g670) & (!g671) & (g672) & (g647) & (!g658)) + ((!g669) & (!g670) & (g671) & (!g672) & (g647) & (!g658)) + ((!g669) & (!g670) & (g671) & (!g672) & (g647) & (g658)) + ((!g669) & (!g670) & (g671) & (g672) & (g647) & (!g658)) + ((!g669) & (g670) & (!g671) & (!g672) & (!g647) & (g658)) + ((!g669) & (g670) & (!g671) & (!g672) & (g647) & (g658)) + ((!g669) & (g670) & (!g671) & (g672) & (!g647) & (g658)) + ((!g669) & (g670) & (g671) & (!g672) & (g647) & (g658)) + ((g669) & (!g670) & (!g671) & (!g672) & (!g647) & (!g658)) + ((g669) & (!g670) & (!g671) & (!g672) & (!g647) & (g658)) + ((g669) & (!g670) & (!g671) & (!g672) & (g647) & (!g658)) + ((g669) & (!g670) & (!g671) & (!g672) & (g647) & (g658)) + ((g669) & (!g670) & (!g671) & (g672) & (!g647) & (!g658)) + ((g669) & (!g670) & (!g671) & (g672) & (!g647) & (g658)) + ((g669) & (!g670) & (!g671) & (g672) & (g647) & (!g658)) + ((g669) & (!g670) & (g671) & (!g672) & (!g647) & (!g658)) + ((g669) & (!g670) & (g671) & (!g672) & (g647) & (!g658)) + ((g669) & (!g670) & (g671) & (!g672) & (g647) & (g658)) + ((g669) & (!g670) & (g671) & (g672) & (!g647) & (!g658)) + ((g669) & (!g670) & (g671) & (g672) & (g647) & (!g658)) + ((g669) & (g670) & (!g671) & (!g672) & (!g647) & (!g658)) + ((g669) & (g670) & (!g671) & (!g672) & (!g647) & (g658)) + ((g669) & (g670) & (!g671) & (!g672) & (g647) & (g658)) + ((g669) & (g670) & (!g671) & (g672) & (!g647) & (!g658)) + ((g669) & (g670) & (!g671) & (g672) & (!g647) & (g658)) + ((g669) & (g670) & (g671) & (!g672) & (!g647) & (!g658)) + ((g669) & (g670) & (g671) & (!g672) & (g647) & (g658)) + ((g669) & (g670) & (g671) & (g672) & (!g647) & (!g658)));
	assign g675 = (((!sk[18]) & (g673) & (!g674)) + ((!sk[18]) & (g673) & (g674)) + ((sk[18]) & (!g673) & (g674)) + ((sk[18]) & (g673) & (!g674)));
	assign g676 = (((!g647) & (!g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (g657) & (g652)) + ((!g647) & (!g648) & (g649) & (g650) & (!g657) & (!g652)) + ((!g647) & (!g648) & (g649) & (g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (g649) & (g650) & (g657) & (g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (g648) & (g649) & (!g650) & (!g657) & (!g652)) + ((!g647) & (g648) & (g649) & (g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((g647) & (!g648) & (g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (g649) & (!g650) & (!g657) & (g652)) + ((g647) & (!g648) & (g649) & (!g650) & (g657) & (!g652)) + ((g647) & (!g648) & (g649) & (g650) & (!g657) & (g652)) + ((g647) & (g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((g647) & (g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((g647) & (g648) & (!g649) & (g650) & (g657) & (!g652)) + ((g647) & (g648) & (g649) & (!g650) & (!g657) & (g652)) + ((g647) & (g648) & (g649) & (!g650) & (g657) & (g652)));
	assign g677 = (((!g647) & (!g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (!g649) & (!g650) & (g657) & (g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (g649) & (g650) & (!g657) & (!g652)) + ((!g647) & (!g648) & (g649) & (g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (g649) & (g650) & (g657) & (g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (g657) & (g652)) + ((!g647) & (g648) & (!g649) & (g650) & (g657) & (g652)) + ((!g647) & (g648) & (g649) & (!g650) & (!g657) & (!g652)) + ((!g647) & (g648) & (g649) & (!g650) & (!g657) & (g652)) + ((!g647) & (g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (g648) & (g649) & (g650) & (!g657) & (g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((g647) & (!g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (!g649) & (g650) & (!g657) & (g652)) + ((g647) & (!g648) & (!g649) & (g650) & (g657) & (g652)) + ((g647) & (!g648) & (g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (g649) & (!g650) & (!g657) & (g652)) + ((g647) & (!g648) & (g649) & (!g650) & (g657) & (g652)) + ((g647) & (!g648) & (g649) & (g650) & (!g657) & (g652)) + ((g647) & (g648) & (!g649) & (g650) & (!g657) & (g652)) + ((g647) & (g648) & (!g649) & (g650) & (g657) & (!g652)) + ((g647) & (g648) & (g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (g648) & (g649) & (g650) & (!g657) & (!g652)));
	assign g678 = (((!g647) & (!g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (!g649) & (!g650) & (g657) & (g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (g649) & (!g650) & (g657) & (g652)) + ((!g647) & (!g648) & (g649) & (g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (g649) & (g650) & (g657) & (g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (g657) & (g652)) + ((!g647) & (g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((!g647) & (g648) & (!g649) & (g650) & (!g657) & (g652)) + ((!g647) & (g648) & (g649) & (!g650) & (!g657) & (g652)) + ((!g647) & (g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (g648) & (g649) & (g650) & (g657) & (g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (g657) & (g652)) + ((g647) & (!g648) & (!g649) & (g650) & (g657) & (g652)) + ((g647) & (!g648) & (g649) & (g650) & (!g657) & (!g652)) + ((g647) & (g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((g647) & (g648) & (!g649) & (g650) & (g657) & (g652)) + ((g647) & (g648) & (g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (g648) & (g649) & (!g650) & (!g657) & (g652)) + ((g647) & (g648) & (g649) & (!g650) & (g657) & (g652)) + ((g647) & (g648) & (g649) & (g650) & (!g657) & (!g652)) + ((g647) & (g648) & (g649) & (g650) & (g657) & (g652)));
	assign g679 = (((!g647) & (!g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (!g649) & (g650) & (g657) & (g652)) + ((!g647) & (!g648) & (g649) & (g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (g649) & (g650) & (g657) & (g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (!g657) & (!g652)) + ((!g647) & (g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (g648) & (!g649) & (g650) & (!g657) & (!g652)) + ((!g647) & (g648) & (!g649) & (g650) & (!g657) & (g652)) + ((!g647) & (g648) & (!g649) & (g650) & (g657) & (!g652)) + ((!g647) & (g648) & (g649) & (!g650) & (!g657) & (!g652)) + ((!g647) & (g648) & (g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (g648) & (g649) & (!g650) & (g657) & (g652)) + ((g647) & (!g648) & (!g649) & (!g650) & (g657) & (g652)) + ((g647) & (!g648) & (!g649) & (g650) & (g657) & (!g652)) + ((g647) & (!g648) & (g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (g649) & (!g650) & (g657) & (!g652)) + ((g647) & (!g648) & (g649) & (!g650) & (g657) & (g652)) + ((g647) & (!g648) & (g649) & (g650) & (!g657) & (g652)) + ((g647) & (!g648) & (g649) & (g650) & (g657) & (!g652)) + ((g647) & (!g648) & (g649) & (g650) & (g657) & (g652)) + ((g647) & (g648) & (!g649) & (!g650) & (!g657) & (g652)) + ((g647) & (g648) & (!g649) & (!g650) & (g657) & (!g652)) + ((g647) & (g648) & (g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (g648) & (g649) & (!g650) & (!g657) & (g652)) + ((g647) & (g648) & (g649) & (g650) & (g657) & (g652)));
	assign g680 = (((!g676) & (!g677) & (!g678) & (!g679) & (!g658) & (g651)) + ((!g676) & (!g677) & (!g678) & (!g679) & (g658) & (!g651)) + ((!g676) & (!g677) & (!g678) & (!g679) & (g658) & (g651)) + ((!g676) & (!g677) & (!g678) & (g679) & (!g658) & (g651)) + ((!g676) & (!g677) & (!g678) & (g679) & (g658) & (!g651)) + ((!g676) & (!g677) & (g678) & (!g679) & (g658) & (!g651)) + ((!g676) & (!g677) & (g678) & (!g679) & (g658) & (g651)) + ((!g676) & (!g677) & (g678) & (g679) & (g658) & (!g651)) + ((!g676) & (g677) & (!g678) & (!g679) & (!g658) & (g651)) + ((!g676) & (g677) & (!g678) & (!g679) & (g658) & (g651)) + ((!g676) & (g677) & (!g678) & (g679) & (!g658) & (g651)) + ((!g676) & (g677) & (g678) & (!g679) & (g658) & (g651)) + ((g676) & (!g677) & (!g678) & (!g679) & (!g658) & (!g651)) + ((g676) & (!g677) & (!g678) & (!g679) & (!g658) & (g651)) + ((g676) & (!g677) & (!g678) & (!g679) & (g658) & (!g651)) + ((g676) & (!g677) & (!g678) & (!g679) & (g658) & (g651)) + ((g676) & (!g677) & (!g678) & (g679) & (!g658) & (!g651)) + ((g676) & (!g677) & (!g678) & (g679) & (!g658) & (g651)) + ((g676) & (!g677) & (!g678) & (g679) & (g658) & (!g651)) + ((g676) & (!g677) & (g678) & (!g679) & (!g658) & (!g651)) + ((g676) & (!g677) & (g678) & (!g679) & (g658) & (!g651)) + ((g676) & (!g677) & (g678) & (!g679) & (g658) & (g651)) + ((g676) & (!g677) & (g678) & (g679) & (!g658) & (!g651)) + ((g676) & (!g677) & (g678) & (g679) & (g658) & (!g651)) + ((g676) & (g677) & (!g678) & (!g679) & (!g658) & (!g651)) + ((g676) & (g677) & (!g678) & (!g679) & (!g658) & (g651)) + ((g676) & (g677) & (!g678) & (!g679) & (g658) & (g651)) + ((g676) & (g677) & (!g678) & (g679) & (!g658) & (!g651)) + ((g676) & (g677) & (!g678) & (g679) & (!g658) & (g651)) + ((g676) & (g677) & (g678) & (!g679) & (!g658) & (!g651)) + ((g676) & (g677) & (g678) & (!g679) & (g658) & (g651)) + ((g676) & (g677) & (g678) & (g679) & (!g658) & (!g651)));
	assign g682 = (((!sk[24]) & (g680) & (!g681)) + ((!sk[24]) & (g680) & (g681)) + ((sk[24]) & (!g680) & (g681)) + ((sk[24]) & (g680) & (!g681)));
	assign g683 = (((!g647) & (!g648) & (!g651) & (!g658) & (!g657) & (g652)) + ((!g647) & (!g648) & (g651) & (!g658) & (!g657) & (g652)) + ((!g647) & (!g648) & (g651) & (!g658) & (g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (!g658) & (g657) & (g652)) + ((!g647) & (!g648) & (g651) & (g658) & (!g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (g658) & (g657) & (!g652)) + ((!g647) & (g648) & (!g651) & (!g658) & (!g657) & (!g652)) + ((!g647) & (g648) & (!g651) & (!g658) & (!g657) & (g652)) + ((!g647) & (g648) & (!g651) & (g658) & (!g657) & (!g652)) + ((!g647) & (g648) & (!g651) & (g658) & (!g657) & (g652)) + ((!g647) & (g648) & (!g651) & (g658) & (g657) & (g652)) + ((!g647) & (g648) & (g651) & (g658) & (!g657) & (g652)) + ((!g647) & (g648) & (g651) & (g658) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g658) & (!g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g658) & (!g657) & (g652)) + ((g647) & (!g648) & (!g651) & (g658) & (!g657) & (g652)) + ((g647) & (!g648) & (g651) & (!g658) & (g657) & (!g652)) + ((g647) & (!g648) & (g651) & (g658) & (!g657) & (!g652)) + ((g647) & (!g648) & (g651) & (g658) & (!g657) & (g652)) + ((g647) & (!g648) & (g651) & (g658) & (g657) & (!g652)) + ((g647) & (g648) & (!g651) & (!g658) & (!g657) & (!g652)) + ((g647) & (g648) & (!g651) & (!g658) & (g657) & (!g652)) + ((g647) & (g648) & (!g651) & (g658) & (g657) & (!g652)) + ((g647) & (g648) & (g651) & (!g658) & (!g657) & (!g652)) + ((g647) & (g648) & (g651) & (!g658) & (!g657) & (g652)) + ((g647) & (g648) & (g651) & (g658) & (!g657) & (g652)));
	assign g684 = (((!g647) & (!g648) & (!g651) & (!g658) & (!g657) & (!g652)) + ((!g647) & (!g648) & (!g651) & (!g658) & (!g657) & (g652)) + ((!g647) & (!g648) & (!g651) & (!g658) & (g657) & (!g652)) + ((!g647) & (!g648) & (!g651) & (!g658) & (g657) & (g652)) + ((!g647) & (!g648) & (!g651) & (g658) & (!g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (!g658) & (!g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (!g658) & (g657) & (g652)) + ((!g647) & (!g648) & (g651) & (g658) & (!g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (g658) & (g657) & (g652)) + ((!g647) & (g648) & (!g651) & (!g658) & (!g657) & (g652)) + ((!g647) & (g648) & (!g651) & (g658) & (g657) & (!g652)) + ((!g647) & (g648) & (g651) & (!g658) & (!g657) & (!g652)) + ((!g647) & (g648) & (g651) & (!g658) & (!g657) & (g652)) + ((!g647) & (g648) & (g651) & (!g658) & (g657) & (!g652)) + ((!g647) & (g648) & (g651) & (!g658) & (g657) & (g652)) + ((!g647) & (g648) & (g651) & (g658) & (!g657) & (!g652)) + ((!g647) & (g648) & (g651) & (g658) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g658) & (!g657) & (g652)) + ((g647) & (!g648) & (!g651) & (!g658) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g658) & (g657) & (g652)) + ((g647) & (!g648) & (!g651) & (g658) & (!g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (g658) & (g657) & (g652)) + ((g647) & (!g648) & (g651) & (!g658) & (g657) & (!g652)) + ((g647) & (!g648) & (g651) & (!g658) & (g657) & (g652)) + ((g647) & (!g648) & (g651) & (g658) & (!g657) & (g652)) + ((g647) & (g648) & (!g651) & (!g658) & (g657) & (!g652)) + ((g647) & (g648) & (!g651) & (!g658) & (g657) & (g652)) + ((g647) & (g648) & (!g651) & (g658) & (!g657) & (!g652)) + ((g647) & (g648) & (!g651) & (g658) & (!g657) & (g652)) + ((g647) & (g648) & (g651) & (!g658) & (g657) & (!g652)) + ((g647) & (g648) & (g651) & (!g658) & (g657) & (g652)) + ((g647) & (g648) & (g651) & (g658) & (!g657) & (g652)));
	assign g685 = (((!g647) & (!g648) & (!g651) & (!g658) & (!g657) & (!g652)) + ((!g647) & (!g648) & (!g651) & (!g658) & (!g657) & (g652)) + ((!g647) & (!g648) & (g651) & (!g658) & (!g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (!g658) & (g657) & (g652)) + ((!g647) & (!g648) & (g651) & (g658) & (!g657) & (g652)) + ((!g647) & (g648) & (!g651) & (g658) & (!g657) & (!g652)) + ((!g647) & (g648) & (!g651) & (g658) & (g657) & (!g652)) + ((!g647) & (g648) & (!g651) & (g658) & (g657) & (g652)) + ((!g647) & (g648) & (g651) & (!g658) & (!g657) & (!g652)) + ((!g647) & (g648) & (g651) & (!g658) & (g657) & (!g652)) + ((!g647) & (g648) & (g651) & (!g658) & (g657) & (g652)) + ((!g647) & (g648) & (g651) & (g658) & (!g657) & (!g652)) + ((!g647) & (g648) & (g651) & (g658) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g658) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g658) & (g657) & (g652)) + ((g647) & (!g648) & (!g651) & (g658) & (!g657) & (g652)) + ((g647) & (!g648) & (!g651) & (g658) & (g657) & (g652)) + ((g647) & (!g648) & (g651) & (!g658) & (!g657) & (!g652)) + ((g647) & (!g648) & (g651) & (!g658) & (!g657) & (g652)) + ((g647) & (!g648) & (g651) & (!g658) & (g657) & (g652)) + ((g647) & (!g648) & (g651) & (g658) & (!g657) & (!g652)) + ((g647) & (!g648) & (g651) & (g658) & (!g657) & (g652)) + ((g647) & (!g648) & (g651) & (g658) & (g657) & (!g652)) + ((g647) & (!g648) & (g651) & (g658) & (g657) & (g652)) + ((g647) & (g648) & (!g651) & (!g658) & (!g657) & (g652)) + ((g647) & (g648) & (!g651) & (g658) & (!g657) & (!g652)) + ((g647) & (g648) & (!g651) & (g658) & (g657) & (!g652)) + ((g647) & (g648) & (g651) & (!g658) & (!g657) & (!g652)) + ((g647) & (g648) & (g651) & (!g658) & (!g657) & (g652)) + ((g647) & (g648) & (g651) & (!g658) & (g657) & (!g652)) + ((g647) & (g648) & (g651) & (g658) & (!g657) & (!g652)) + ((g647) & (g648) & (g651) & (g658) & (g657) & (!g652)));
	assign g686 = (((!g647) & (!g648) & (!g651) & (!g658) & (g657) & (g652)) + ((!g647) & (!g648) & (!g651) & (g658) & (!g657) & (!g652)) + ((!g647) & (!g648) & (!g651) & (g658) & (g657) & (g652)) + ((!g647) & (!g648) & (g651) & (!g658) & (!g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (!g658) & (g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (g658) & (!g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (g658) & (!g657) & (g652)) + ((!g647) & (!g648) & (g651) & (g658) & (g657) & (!g652)) + ((!g647) & (g648) & (!g651) & (!g658) & (!g657) & (!g652)) + ((!g647) & (g648) & (!g651) & (g658) & (!g657) & (g652)) + ((!g647) & (g648) & (!g651) & (g658) & (g657) & (!g652)) + ((!g647) & (g648) & (!g651) & (g658) & (g657) & (g652)) + ((!g647) & (g648) & (g651) & (!g658) & (!g657) & (!g652)) + ((!g647) & (g648) & (g651) & (g658) & (!g657) & (!g652)) + ((!g647) & (g648) & (g651) & (g658) & (!g657) & (g652)) + ((g647) & (!g648) & (!g651) & (!g658) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g658) & (g657) & (g652)) + ((g647) & (!g648) & (g651) & (!g658) & (!g657) & (!g652)) + ((g647) & (!g648) & (g651) & (!g658) & (g657) & (!g652)) + ((g647) & (!g648) & (g651) & (g658) & (g657) & (!g652)) + ((g647) & (g648) & (!g651) & (!g658) & (g657) & (!g652)) + ((g647) & (g648) & (!g651) & (g658) & (g657) & (g652)) + ((g647) & (g648) & (g651) & (!g658) & (!g657) & (!g652)) + ((g647) & (g648) & (g651) & (!g658) & (!g657) & (g652)) + ((g647) & (g648) & (g651) & (!g658) & (g657) & (!g652)) + ((g647) & (g648) & (g651) & (g658) & (!g657) & (!g652)));
	assign g687 = (((!g683) & (!g684) & (!g685) & (!g686) & (g649) & (g650)) + ((!g683) & (!g684) & (g685) & (!g686) & (!g649) & (g650)) + ((!g683) & (!g684) & (g685) & (!g686) & (g649) & (g650)) + ((!g683) & (!g684) & (g685) & (g686) & (!g649) & (g650)) + ((!g683) & (g684) & (!g685) & (!g686) & (g649) & (!g650)) + ((!g683) & (g684) & (!g685) & (!g686) & (g649) & (g650)) + ((!g683) & (g684) & (!g685) & (g686) & (g649) & (!g650)) + ((!g683) & (g684) & (g685) & (!g686) & (!g649) & (g650)) + ((!g683) & (g684) & (g685) & (!g686) & (g649) & (!g650)) + ((!g683) & (g684) & (g685) & (!g686) & (g649) & (g650)) + ((!g683) & (g684) & (g685) & (g686) & (!g649) & (g650)) + ((!g683) & (g684) & (g685) & (g686) & (g649) & (!g650)) + ((g683) & (!g684) & (!g685) & (!g686) & (!g649) & (!g650)) + ((g683) & (!g684) & (!g685) & (!g686) & (g649) & (g650)) + ((g683) & (!g684) & (!g685) & (g686) & (!g649) & (!g650)) + ((g683) & (!g684) & (g685) & (!g686) & (!g649) & (!g650)) + ((g683) & (!g684) & (g685) & (!g686) & (!g649) & (g650)) + ((g683) & (!g684) & (g685) & (!g686) & (g649) & (g650)) + ((g683) & (!g684) & (g685) & (g686) & (!g649) & (!g650)) + ((g683) & (!g684) & (g685) & (g686) & (!g649) & (g650)) + ((g683) & (g684) & (!g685) & (!g686) & (!g649) & (!g650)) + ((g683) & (g684) & (!g685) & (!g686) & (g649) & (!g650)) + ((g683) & (g684) & (!g685) & (!g686) & (g649) & (g650)) + ((g683) & (g684) & (!g685) & (g686) & (!g649) & (!g650)) + ((g683) & (g684) & (!g685) & (g686) & (g649) & (!g650)) + ((g683) & (g684) & (g685) & (!g686) & (!g649) & (!g650)) + ((g683) & (g684) & (g685) & (!g686) & (!g649) & (g650)) + ((g683) & (g684) & (g685) & (!g686) & (g649) & (!g650)) + ((g683) & (g684) & (g685) & (!g686) & (g649) & (g650)) + ((g683) & (g684) & (g685) & (g686) & (!g649) & (!g650)) + ((g683) & (g684) & (g685) & (g686) & (!g649) & (g650)) + ((g683) & (g684) & (g685) & (g686) & (g649) & (!g650)));
	assign g689 = (((!g687) & (sk[30]) & (g688)) + ((g687) & (!sk[30]) & (!g688)) + ((g687) & (!sk[30]) & (g688)) + ((g687) & (sk[30]) & (!g688)));
	assign g690 = (((!g647) & (!g648) & (!g651) & (!g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (!g651) & (!g650) & (g657) & (g652)) + ((!g647) & (!g648) & (!g651) & (g650) & (g657) & (g652)) + ((!g647) & (!g648) & (g651) & (!g650) & (!g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (!g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (g651) & (!g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (!g650) & (g657) & (g652)) + ((!g647) & (!g648) & (g651) & (g650) & (!g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (g650) & (!g657) & (g652)) + ((!g647) & (g648) & (!g651) & (!g650) & (!g657) & (g652)) + ((!g647) & (g648) & (!g651) & (!g650) & (g657) & (!g652)) + ((!g647) & (g648) & (!g651) & (g650) & (g657) & (g652)) + ((!g647) & (g648) & (g651) & (!g650) & (g657) & (!g652)) + ((!g647) & (g648) & (g651) & (!g650) & (g657) & (g652)) + ((!g647) & (g648) & (g651) & (g650) & (!g657) & (!g652)) + ((!g647) & (g648) & (g651) & (g650) & (!g657) & (g652)) + ((!g647) & (g648) & (g651) & (g650) & (g657) & (g652)) + ((g647) & (!g648) & (!g651) & (!g650) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g650) & (g657) & (g652)) + ((g647) & (!g648) & (!g651) & (g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (g650) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (g650) & (g657) & (g652)) + ((g647) & (!g648) & (g651) & (!g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (g651) & (!g650) & (g657) & (!g652)) + ((g647) & (!g648) & (g651) & (g650) & (g657) & (!g652)) + ((g647) & (g648) & (!g651) & (!g650) & (g657) & (g652)) + ((g647) & (g648) & (g651) & (!g650) & (!g657) & (!g652)) + ((g647) & (g648) & (g651) & (!g650) & (g657) & (g652)));
	assign g691 = (((!g647) & (!g648) & (!g651) & (!g650) & (!g657) & (!g652)) + ((!g647) & (!g648) & (!g651) & (g650) & (!g657) & (!g652)) + ((!g647) & (!g648) & (!g651) & (g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (!g651) & (g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (!g650) & (g657) & (g652)) + ((!g647) & (!g648) & (g651) & (g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (g651) & (g650) & (g657) & (g652)) + ((!g647) & (g648) & (!g651) & (!g650) & (!g657) & (!g652)) + ((!g647) & (g648) & (!g651) & (!g650) & (g657) & (!g652)) + ((!g647) & (g648) & (g651) & (!g650) & (!g657) & (g652)) + ((!g647) & (g648) & (g651) & (!g650) & (g657) & (g652)) + ((!g647) & (g648) & (g651) & (g650) & (!g657) & (g652)) + ((!g647) & (g648) & (g651) & (g650) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g650) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g650) & (g657) & (g652)) + ((g647) & (!g648) & (!g651) & (g650) & (!g657) & (g652)) + ((g647) & (!g648) & (!g651) & (g650) & (g657) & (g652)) + ((g647) & (!g648) & (g651) & (g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (g651) & (g650) & (!g657) & (g652)) + ((g647) & (!g648) & (g651) & (g650) & (g657) & (g652)) + ((g647) & (g648) & (!g651) & (!g650) & (!g657) & (g652)) + ((g647) & (g648) & (!g651) & (!g650) & (g657) & (!g652)) + ((g647) & (g648) & (!g651) & (g650) & (g657) & (!g652)) + ((g647) & (g648) & (g651) & (!g650) & (!g657) & (g652)) + ((g647) & (g648) & (g651) & (!g650) & (g657) & (g652)) + ((g647) & (g648) & (g651) & (g650) & (!g657) & (!g652)) + ((g647) & (g648) & (g651) & (g650) & (g657) & (g652)));
	assign g692 = (((!g647) & (!g648) & (!g651) & (!g650) & (g657) & (g652)) + ((!g647) & (!g648) & (!g651) & (g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (!g650) & (!g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (!g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (g651) & (!g650) & (g657) & (g652)) + ((!g647) & (!g648) & (g651) & (g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (g651) & (g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (g651) & (g650) & (g657) & (g652)) + ((!g647) & (g648) & (!g651) & (!g650) & (g657) & (!g652)) + ((!g647) & (g648) & (!g651) & (!g650) & (g657) & (g652)) + ((!g647) & (g648) & (g651) & (!g650) & (!g657) & (!g652)) + ((!g647) & (g648) & (g651) & (g650) & (!g657) & (g652)) + ((!g647) & (g648) & (g651) & (g650) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g650) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (!g650) & (g657) & (g652)) + ((g647) & (!g648) & (!g651) & (g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (g650) & (!g657) & (g652)) + ((g647) & (!g648) & (g651) & (!g650) & (!g657) & (g652)) + ((g647) & (!g648) & (g651) & (!g650) & (g657) & (g652)) + ((g647) & (!g648) & (g651) & (g650) & (g657) & (!g652)) + ((g647) & (g648) & (!g651) & (!g650) & (!g657) & (!g652)) + ((g647) & (g648) & (!g651) & (!g650) & (!g657) & (g652)) + ((g647) & (g648) & (!g651) & (!g650) & (g657) & (g652)) + ((g647) & (g648) & (!g651) & (g650) & (!g657) & (g652)) + ((g647) & (g648) & (!g651) & (g650) & (g657) & (!g652)) + ((g647) & (g648) & (g651) & (!g650) & (!g657) & (g652)) + ((g647) & (g648) & (g651) & (!g650) & (g657) & (!g652)) + ((g647) & (g648) & (g651) & (g650) & (!g657) & (!g652)) + ((g647) & (g648) & (g651) & (g650) & (g657) & (!g652)) + ((g647) & (g648) & (g651) & (g650) & (g657) & (g652)));
	assign g693 = (((!g647) & (!g648) & (!g651) & (!g650) & (g657) & (!g652)) + ((!g647) & (!g648) & (!g651) & (g650) & (!g657) & (!g652)) + ((!g647) & (!g648) & (!g651) & (g650) & (g657) & (g652)) + ((!g647) & (!g648) & (g651) & (!g650) & (!g657) & (g652)) + ((!g647) & (!g648) & (g651) & (!g650) & (g657) & (g652)) + ((!g647) & (!g648) & (g651) & (g650) & (g657) & (g652)) + ((!g647) & (g648) & (!g651) & (!g650) & (!g657) & (g652)) + ((!g647) & (g648) & (!g651) & (g650) & (!g657) & (g652)) + ((!g647) & (g648) & (!g651) & (g650) & (g657) & (g652)) + ((!g647) & (g648) & (g651) & (!g650) & (!g657) & (!g652)) + ((!g647) & (g648) & (g651) & (!g650) & (g657) & (!g652)) + ((!g647) & (g648) & (g651) & (g650) & (!g657) & (g652)) + ((!g647) & (g648) & (g651) & (g650) & (g657) & (g652)) + ((g647) & (!g648) & (!g651) & (!g650) & (g657) & (!g652)) + ((g647) & (!g648) & (!g651) & (g650) & (g657) & (g652)) + ((g647) & (!g648) & (g651) & (!g650) & (!g657) & (!g652)) + ((g647) & (!g648) & (g651) & (!g650) & (g657) & (g652)) + ((g647) & (!g648) & (g651) & (g650) & (!g657) & (!g652)) + ((g647) & (g648) & (!g651) & (!g650) & (g657) & (g652)) + ((g647) & (g648) & (!g651) & (g650) & (!g657) & (!g652)) + ((g647) & (g648) & (!g651) & (g650) & (!g657) & (g652)) + ((g647) & (g648) & (g651) & (!g650) & (g657) & (g652)));
	assign g694 = (((!g690) & (!g691) & (!g692) & (!g693) & (!g658) & (!g649)) + ((!g690) & (!g691) & (!g692) & (!g693) & (!g658) & (g649)) + ((!g690) & (!g691) & (!g692) & (!g693) & (g658) & (!g649)) + ((!g690) & (!g691) & (!g692) & (g693) & (!g658) & (!g649)) + ((!g690) & (!g691) & (!g692) & (g693) & (!g658) & (g649)) + ((!g690) & (!g691) & (!g692) & (g693) & (g658) & (!g649)) + ((!g690) & (!g691) & (!g692) & (g693) & (g658) & (g649)) + ((!g690) & (!g691) & (g692) & (!g693) & (!g658) & (!g649)) + ((!g690) & (!g691) & (g692) & (!g693) & (g658) & (!g649)) + ((!g690) & (!g691) & (g692) & (g693) & (!g658) & (!g649)) + ((!g690) & (!g691) & (g692) & (g693) & (g658) & (!g649)) + ((!g690) & (!g691) & (g692) & (g693) & (g658) & (g649)) + ((!g690) & (g691) & (!g692) & (!g693) & (!g658) & (!g649)) + ((!g690) & (g691) & (!g692) & (!g693) & (!g658) & (g649)) + ((!g690) & (g691) & (!g692) & (g693) & (!g658) & (!g649)) + ((!g690) & (g691) & (!g692) & (g693) & (!g658) & (g649)) + ((!g690) & (g691) & (!g692) & (g693) & (g658) & (g649)) + ((!g690) & (g691) & (g692) & (!g693) & (!g658) & (!g649)) + ((!g690) & (g691) & (g692) & (g693) & (!g658) & (!g649)) + ((!g690) & (g691) & (g692) & (g693) & (g658) & (g649)) + ((g690) & (!g691) & (!g692) & (!g693) & (!g658) & (g649)) + ((g690) & (!g691) & (!g692) & (!g693) & (g658) & (!g649)) + ((g690) & (!g691) & (!g692) & (g693) & (!g658) & (g649)) + ((g690) & (!g691) & (!g692) & (g693) & (g658) & (!g649)) + ((g690) & (!g691) & (!g692) & (g693) & (g658) & (g649)) + ((g690) & (!g691) & (g692) & (!g693) & (g658) & (!g649)) + ((g690) & (!g691) & (g692) & (g693) & (g658) & (!g649)) + ((g690) & (!g691) & (g692) & (g693) & (g658) & (g649)) + ((g690) & (g691) & (!g692) & (!g693) & (!g658) & (g649)) + ((g690) & (g691) & (!g692) & (g693) & (!g658) & (g649)) + ((g690) & (g691) & (!g692) & (g693) & (g658) & (g649)) + ((g690) & (g691) & (g692) & (g693) & (g658) & (g649)));
	assign g696 = (((!sk[36]) & (g694) & (!g695)) + ((!sk[36]) & (g694) & (g695)) + ((sk[36]) & (!g694) & (g695)) + ((sk[36]) & (g694) & (!g695)));
	assign g697 = (((!g647) & (!g658) & (!g649) & (!g650) & (!g657) & (g652)) + ((!g647) & (!g658) & (!g649) & (!g650) & (g657) & (g652)) + ((!g647) & (!g658) & (!g649) & (g650) & (!g657) & (!g652)) + ((!g647) & (!g658) & (!g649) & (g650) & (!g657) & (g652)) + ((!g647) & (!g658) & (!g649) & (g650) & (g657) & (!g652)) + ((!g647) & (!g658) & (!g649) & (g650) & (g657) & (g652)) + ((!g647) & (!g658) & (g649) & (!g650) & (!g657) & (g652)) + ((!g647) & (!g658) & (g649) & (!g650) & (g657) & (g652)) + ((!g647) & (!g658) & (g649) & (g650) & (g657) & (!g652)) + ((!g647) & (g658) & (g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (g658) & (g649) & (!g650) & (g657) & (g652)) + ((!g647) & (g658) & (g649) & (g650) & (!g657) & (g652)) + ((g647) & (!g658) & (!g649) & (!g650) & (g657) & (!g652)) + ((g647) & (!g658) & (!g649) & (g650) & (!g657) & (!g652)) + ((g647) & (!g658) & (!g649) & (g650) & (!g657) & (g652)) + ((g647) & (!g658) & (!g649) & (g650) & (g657) & (g652)) + ((g647) & (!g658) & (g649) & (!g650) & (!g657) & (g652)) + ((g647) & (!g658) & (g649) & (!g650) & (g657) & (g652)) + ((g647) & (!g658) & (g649) & (g650) & (g657) & (!g652)) + ((g647) & (!g658) & (g649) & (g650) & (g657) & (g652)) + ((g647) & (g658) & (!g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (g658) & (!g649) & (!g650) & (!g657) & (g652)) + ((g647) & (g658) & (!g649) & (!g650) & (g657) & (!g652)) + ((g647) & (g658) & (!g649) & (g650) & (!g657) & (!g652)) + ((g647) & (g658) & (g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (g658) & (g649) & (!g650) & (!g657) & (g652)) + ((g647) & (g658) & (g649) & (!g650) & (g657) & (!g652)) + ((g647) & (g658) & (g649) & (g650) & (!g657) & (g652)));
	assign g698 = (((!g647) & (!g658) & (!g649) & (!g650) & (!g657) & (!g652)) + ((!g647) & (!g658) & (!g649) & (g650) & (g657) & (g652)) + ((!g647) & (!g658) & (g649) & (!g650) & (!g657) & (!g652)) + ((!g647) & (!g658) & (g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (!g658) & (g649) & (!g650) & (g657) & (g652)) + ((!g647) & (!g658) & (g649) & (g650) & (!g657) & (!g652)) + ((!g647) & (!g658) & (g649) & (g650) & (g657) & (g652)) + ((!g647) & (g658) & (!g649) & (!g650) & (!g657) & (!g652)) + ((!g647) & (g658) & (!g649) & (!g650) & (g657) & (g652)) + ((!g647) & (g658) & (!g649) & (g650) & (!g657) & (g652)) + ((!g647) & (g658) & (g649) & (!g650) & (!g657) & (!g652)) + ((!g647) & (g658) & (g649) & (!g650) & (g657) & (g652)) + ((!g647) & (g658) & (g649) & (g650) & (g657) & (!g652)) + ((!g647) & (g658) & (g649) & (g650) & (g657) & (g652)) + ((g647) & (!g658) & (!g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (!g658) & (!g649) & (!g650) & (g657) & (g652)) + ((g647) & (!g658) & (!g649) & (g650) & (!g657) & (!g652)) + ((g647) & (!g658) & (!g649) & (g650) & (g657) & (g652)) + ((g647) & (!g658) & (g649) & (!g650) & (g657) & (g652)) + ((g647) & (!g658) & (g649) & (g650) & (!g657) & (g652)) + ((g647) & (g658) & (!g649) & (!g650) & (g657) & (!g652)) + ((g647) & (g658) & (!g649) & (!g650) & (g657) & (g652)) + ((g647) & (g658) & (!g649) & (g650) & (!g657) & (g652)) + ((g647) & (g658) & (!g649) & (g650) & (g657) & (!g652)) + ((g647) & (g658) & (!g649) & (g650) & (g657) & (g652)) + ((g647) & (g658) & (g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (g658) & (g649) & (!g650) & (g657) & (!g652)) + ((g647) & (g658) & (g649) & (g650) & (!g657) & (!g652)));
	assign g699 = (((!g647) & (!g658) & (!g649) & (!g650) & (!g657) & (g652)) + ((!g647) & (!g658) & (!g649) & (!g650) & (g657) & (g652)) + ((!g647) & (!g658) & (!g649) & (g650) & (g657) & (!g652)) + ((!g647) & (!g658) & (!g649) & (g650) & (g657) & (g652)) + ((!g647) & (!g658) & (g649) & (!g650) & (g657) & (g652)) + ((!g647) & (!g658) & (g649) & (g650) & (!g657) & (!g652)) + ((!g647) & (!g658) & (g649) & (g650) & (!g657) & (g652)) + ((!g647) & (!g658) & (g649) & (g650) & (g657) & (g652)) + ((!g647) & (g658) & (!g649) & (!g650) & (!g657) & (!g652)) + ((!g647) & (g658) & (!g649) & (!g650) & (!g657) & (g652)) + ((!g647) & (g658) & (!g649) & (!g650) & (g657) & (g652)) + ((!g647) & (g658) & (!g649) & (g650) & (!g657) & (g652)) + ((!g647) & (g658) & (!g649) & (g650) & (g657) & (!g652)) + ((!g647) & (g658) & (g649) & (!g650) & (!g657) & (g652)) + ((!g647) & (g658) & (g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (g658) & (g649) & (g650) & (!g657) & (!g652)) + ((!g647) & (g658) & (g649) & (g650) & (g657) & (!g652)) + ((!g647) & (g658) & (g649) & (g650) & (g657) & (g652)) + ((g647) & (!g658) & (!g649) & (!g650) & (!g657) & (g652)) + ((g647) & (!g658) & (!g649) & (g650) & (!g657) & (!g652)) + ((g647) & (!g658) & (!g649) & (g650) & (g657) & (!g652)) + ((g647) & (!g658) & (g649) & (!g650) & (g657) & (g652)) + ((g647) & (!g658) & (g649) & (g650) & (!g657) & (g652)) + ((g647) & (g658) & (!g649) & (!g650) & (!g657) & (g652)) + ((g647) & (g658) & (!g649) & (g650) & (!g657) & (!g652)) + ((g647) & (g658) & (!g649) & (g650) & (g657) & (!g652)) + ((g647) & (g658) & (g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (g658) & (g649) & (!g650) & (g657) & (!g652)) + ((g647) & (g658) & (g649) & (!g650) & (g657) & (g652)) + ((g647) & (g658) & (g649) & (g650) & (g657) & (g652)));
	assign g700 = (((!g647) & (!g658) & (!g649) & (!g650) & (g657) & (g652)) + ((!g647) & (!g658) & (!g649) & (g650) & (!g657) & (!g652)) + ((!g647) & (!g658) & (!g649) & (g650) & (g657) & (g652)) + ((!g647) & (!g658) & (g649) & (!g650) & (!g657) & (!g652)) + ((!g647) & (!g658) & (g649) & (g650) & (g657) & (!g652)) + ((!g647) & (!g658) & (g649) & (g650) & (g657) & (g652)) + ((!g647) & (g658) & (!g649) & (g650) & (!g657) & (!g652)) + ((!g647) & (g658) & (!g649) & (g650) & (g657) & (!g652)) + ((!g647) & (g658) & (g649) & (!g650) & (g657) & (!g652)) + ((!g647) & (g658) & (g649) & (!g650) & (g657) & (g652)) + ((g647) & (!g658) & (!g649) & (!g650) & (!g657) & (g652)) + ((g647) & (!g658) & (!g649) & (!g650) & (g657) & (!g652)) + ((g647) & (!g658) & (!g649) & (g650) & (!g657) & (g652)) + ((g647) & (!g658) & (g649) & (!g650) & (g657) & (!g652)) + ((g647) & (!g658) & (g649) & (!g650) & (g657) & (g652)) + ((g647) & (!g658) & (g649) & (g650) & (g657) & (!g652)) + ((g647) & (!g658) & (g649) & (g650) & (g657) & (g652)) + ((g647) & (g658) & (!g649) & (!g650) & (g657) & (!g652)) + ((g647) & (g658) & (!g649) & (g650) & (!g657) & (g652)) + ((g647) & (g658) & (g649) & (!g650) & (!g657) & (!g652)) + ((g647) & (g658) & (g649) & (!g650) & (g657) & (g652)) + ((g647) & (g658) & (g649) & (g650) & (!g657) & (g652)));
	assign g701 = (((!g697) & (!g698) & (!g699) & (!g700) & (!g651) & (!g648)) + ((!g697) & (!g698) & (!g699) & (!g700) & (!g651) & (g648)) + ((!g697) & (!g698) & (!g699) & (!g700) & (g651) & (!g648)) + ((!g697) & (!g698) & (!g699) & (g700) & (!g651) & (!g648)) + ((!g697) & (!g698) & (!g699) & (g700) & (!g651) & (g648)) + ((!g697) & (!g698) & (!g699) & (g700) & (g651) & (!g648)) + ((!g697) & (!g698) & (!g699) & (g700) & (g651) & (g648)) + ((!g697) & (!g698) & (g699) & (!g700) & (!g651) & (!g648)) + ((!g697) & (!g698) & (g699) & (!g700) & (g651) & (!g648)) + ((!g697) & (!g698) & (g699) & (g700) & (!g651) & (!g648)) + ((!g697) & (!g698) & (g699) & (g700) & (g651) & (!g648)) + ((!g697) & (!g698) & (g699) & (g700) & (g651) & (g648)) + ((!g697) & (g698) & (!g699) & (!g700) & (!g651) & (!g648)) + ((!g697) & (g698) & (!g699) & (!g700) & (!g651) & (g648)) + ((!g697) & (g698) & (!g699) & (g700) & (!g651) & (!g648)) + ((!g697) & (g698) & (!g699) & (g700) & (!g651) & (g648)) + ((!g697) & (g698) & (!g699) & (g700) & (g651) & (g648)) + ((!g697) & (g698) & (g699) & (!g700) & (!g651) & (!g648)) + ((!g697) & (g698) & (g699) & (g700) & (!g651) & (!g648)) + ((!g697) & (g698) & (g699) & (g700) & (g651) & (g648)) + ((g697) & (!g698) & (!g699) & (!g700) & (!g651) & (g648)) + ((g697) & (!g698) & (!g699) & (!g700) & (g651) & (!g648)) + ((g697) & (!g698) & (!g699) & (g700) & (!g651) & (g648)) + ((g697) & (!g698) & (!g699) & (g700) & (g651) & (!g648)) + ((g697) & (!g698) & (!g699) & (g700) & (g651) & (g648)) + ((g697) & (!g698) & (g699) & (!g700) & (g651) & (!g648)) + ((g697) & (!g698) & (g699) & (g700) & (g651) & (!g648)) + ((g697) & (!g698) & (g699) & (g700) & (g651) & (g648)) + ((g697) & (g698) & (!g699) & (!g700) & (!g651) & (g648)) + ((g697) & (g698) & (!g699) & (g700) & (!g651) & (g648)) + ((g697) & (g698) & (!g699) & (g700) & (g651) & (g648)) + ((g697) & (g698) & (g699) & (g700) & (g651) & (g648)));
	assign g703 = (((!sk[42]) & (g701) & (!g702)) + ((!sk[42]) & (g701) & (g702)) + ((sk[42]) & (!g701) & (g702)) + ((sk[42]) & (g701) & (!g702)));
	assign g704 = (((!g651) & (!g648) & (!g649) & (!g650) & (!g657) & (g658)) + ((!g651) & (!g648) & (!g649) & (!g650) & (g657) & (!g658)) + ((!g651) & (!g648) & (!g649) & (g650) & (!g657) & (g658)) + ((!g651) & (!g648) & (!g649) & (g650) & (g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (!g650) & (!g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (!g650) & (g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (g650) & (!g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (g650) & (g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (g650) & (g657) & (g658)) + ((!g651) & (g648) & (!g649) & (!g650) & (g657) & (!g658)) + ((!g651) & (g648) & (!g649) & (g650) & (g657) & (!g658)) + ((!g651) & (g648) & (!g649) & (g650) & (g657) & (g658)) + ((!g651) & (g648) & (g649) & (!g650) & (g657) & (g658)) + ((!g651) & (g648) & (g649) & (g650) & (!g657) & (!g658)) + ((g651) & (!g648) & (!g649) & (!g650) & (!g657) & (g658)) + ((g651) & (!g648) & (!g649) & (g650) & (!g657) & (g658)) + ((g651) & (!g648) & (g649) & (g650) & (g657) & (g658)) + ((g651) & (g648) & (!g649) & (!g650) & (g657) & (g658)) + ((g651) & (g648) & (!g649) & (g650) & (!g657) & (!g658)) + ((g651) & (g648) & (!g649) & (g650) & (g657) & (!g658)) + ((g651) & (g648) & (g649) & (!g650) & (!g657) & (g658)) + ((g651) & (g648) & (g649) & (!g650) & (g657) & (!g658)) + ((g651) & (g648) & (g649) & (!g650) & (g657) & (g658)) + ((g651) & (g648) & (g649) & (g650) & (!g657) & (g658)));
	assign g705 = (((!g651) & (!g648) & (!g649) & (!g650) & (!g657) & (!g658)) + ((!g651) & (!g648) & (!g649) & (!g650) & (!g657) & (g658)) + ((!g651) & (!g648) & (!g649) & (g650) & (!g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (!g650) & (!g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (!g650) & (g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (!g650) & (g657) & (g658)) + ((!g651) & (!g648) & (g649) & (g650) & (!g657) & (g658)) + ((!g651) & (!g648) & (g649) & (g650) & (g657) & (g658)) + ((!g651) & (g648) & (!g649) & (!g650) & (!g657) & (!g658)) + ((!g651) & (g648) & (!g649) & (!g650) & (g657) & (!g658)) + ((!g651) & (g648) & (!g649) & (g650) & (!g657) & (!g658)) + ((!g651) & (g648) & (!g649) & (g650) & (!g657) & (g658)) + ((!g651) & (g648) & (!g649) & (g650) & (g657) & (g658)) + ((!g651) & (g648) & (g649) & (!g650) & (!g657) & (g658)) + ((!g651) & (g648) & (g649) & (g650) & (!g657) & (!g658)) + ((!g651) & (g648) & (g649) & (g650) & (!g657) & (g658)) + ((g651) & (!g648) & (!g649) & (!g650) & (!g657) & (g658)) + ((g651) & (!g648) & (!g649) & (!g650) & (g657) & (g658)) + ((g651) & (!g648) & (!g649) & (g650) & (!g657) & (!g658)) + ((g651) & (!g648) & (!g649) & (g650) & (g657) & (g658)) + ((g651) & (!g648) & (g649) & (!g650) & (!g657) & (!g658)) + ((g651) & (!g648) & (g649) & (!g650) & (g657) & (g658)) + ((g651) & (!g648) & (g649) & (g650) & (g657) & (!g658)) + ((g651) & (g648) & (!g649) & (!g650) & (!g657) & (!g658)) + ((g651) & (g648) & (!g649) & (!g650) & (!g657) & (g658)) + ((g651) & (g648) & (!g649) & (!g650) & (g657) & (g658)) + ((g651) & (g648) & (!g649) & (g650) & (!g657) & (g658)) + ((g651) & (g648) & (!g649) & (g650) & (g657) & (!g658)) + ((g651) & (g648) & (g649) & (!g650) & (g657) & (!g658)) + ((g651) & (g648) & (g649) & (!g650) & (g657) & (g658)));
	assign g706 = (((!g651) & (!g648) & (!g649) & (!g650) & (g657) & (!g658)) + ((!g651) & (!g648) & (!g649) & (g650) & (!g657) & (!g658)) + ((!g651) & (!g648) & (!g649) & (g650) & (g657) & (!g658)) + ((!g651) & (!g648) & (!g649) & (g650) & (g657) & (g658)) + ((!g651) & (!g648) & (g649) & (!g650) & (!g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (!g650) & (!g657) & (g658)) + ((!g651) & (!g648) & (g649) & (!g650) & (g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (g650) & (!g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (g650) & (g657) & (g658)) + ((!g651) & (g648) & (!g649) & (!g650) & (!g657) & (g658)) + ((!g651) & (g648) & (!g649) & (!g650) & (g657) & (!g658)) + ((!g651) & (g648) & (!g649) & (!g650) & (g657) & (g658)) + ((!g651) & (g648) & (g649) & (!g650) & (!g657) & (g658)) + ((!g651) & (g648) & (g649) & (!g650) & (g657) & (!g658)) + ((!g651) & (g648) & (g649) & (!g650) & (g657) & (g658)) + ((!g651) & (g648) & (g649) & (g650) & (!g657) & (!g658)) + ((g651) & (!g648) & (!g649) & (!g650) & (g657) & (!g658)) + ((g651) & (!g648) & (!g649) & (g650) & (!g657) & (!g658)) + ((g651) & (!g648) & (!g649) & (g650) & (g657) & (g658)) + ((g651) & (!g648) & (g649) & (!g650) & (!g657) & (!g658)) + ((g651) & (!g648) & (g649) & (!g650) & (!g657) & (g658)) + ((g651) & (!g648) & (g649) & (g650) & (!g657) & (!g658)) + ((g651) & (!g648) & (g649) & (g650) & (g657) & (!g658)) + ((g651) & (g648) & (!g649) & (!g650) & (g657) & (!g658)) + ((g651) & (g648) & (!g649) & (g650) & (!g657) & (!g658)) + ((g651) & (g648) & (!g649) & (g650) & (g657) & (g658)) + ((g651) & (g648) & (g649) & (!g650) & (!g657) & (!g658)) + ((g651) & (g648) & (g649) & (!g650) & (g657) & (!g658)) + ((g651) & (g648) & (g649) & (!g650) & (g657) & (g658)) + ((g651) & (g648) & (g649) & (g650) & (!g657) & (g658)));
	assign g707 = (((!g651) & (!g648) & (!g649) & (!g650) & (!g657) & (g658)) + ((!g651) & (!g648) & (!g649) & (g650) & (g657) & (!g658)) + ((!g651) & (!g648) & (!g649) & (g650) & (g657) & (g658)) + ((!g651) & (!g648) & (g649) & (!g650) & (!g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (!g650) & (!g657) & (g658)) + ((!g651) & (!g648) & (g649) & (g650) & (g657) & (!g658)) + ((!g651) & (!g648) & (g649) & (g650) & (g657) & (g658)) + ((!g651) & (g648) & (!g649) & (!g650) & (!g657) & (!g658)) + ((!g651) & (g648) & (!g649) & (!g650) & (!g657) & (g658)) + ((!g651) & (g648) & (!g649) & (!g650) & (g657) & (g658)) + ((!g651) & (g648) & (!g649) & (g650) & (!g657) & (g658)) + ((!g651) & (g648) & (g649) & (!g650) & (!g657) & (g658)) + ((!g651) & (g648) & (g649) & (g650) & (!g657) & (!g658)) + ((!g651) & (g648) & (g649) & (g650) & (!g657) & (g658)) + ((!g651) & (g648) & (g649) & (g650) & (g657) & (!g658)) + ((!g651) & (g648) & (g649) & (g650) & (g657) & (g658)) + ((g651) & (!g648) & (!g649) & (g650) & (!g657) & (g658)) + ((g651) & (!g648) & (g649) & (!g650) & (!g657) & (!g658)) + ((g651) & (!g648) & (g649) & (g650) & (!g657) & (!g658)) + ((g651) & (!g648) & (g649) & (g650) & (!g657) & (g658)) + ((g651) & (!g648) & (g649) & (g650) & (g657) & (g658)) + ((g651) & (g648) & (!g649) & (!g650) & (!g657) & (g658)) + ((g651) & (g648) & (!g649) & (!g650) & (g657) & (g658)) + ((g651) & (g648) & (!g649) & (g650) & (!g657) & (!g658)) + ((g651) & (g648) & (!g649) & (g650) & (g657) & (!g658)) + ((g651) & (g648) & (!g649) & (g650) & (g657) & (g658)) + ((g651) & (g648) & (g649) & (!g650) & (g657) & (g658)) + ((g651) & (g648) & (g649) & (g650) & (g657) & (g658)));
	assign g708 = (((!g704) & (!g705) & (!g706) & (!g707) & (!g647) & (g652)) + ((!g704) & (!g705) & (!g706) & (!g707) & (g647) & (!g652)) + ((!g704) & (!g705) & (!g706) & (!g707) & (g647) & (g652)) + ((!g704) & (!g705) & (!g706) & (g707) & (!g647) & (g652)) + ((!g704) & (!g705) & (!g706) & (g707) & (g647) & (!g652)) + ((!g704) & (!g705) & (g706) & (!g707) & (g647) & (!g652)) + ((!g704) & (!g705) & (g706) & (!g707) & (g647) & (g652)) + ((!g704) & (!g705) & (g706) & (g707) & (g647) & (!g652)) + ((!g704) & (g705) & (!g706) & (!g707) & (!g647) & (g652)) + ((!g704) & (g705) & (!g706) & (!g707) & (g647) & (g652)) + ((!g704) & (g705) & (!g706) & (g707) & (!g647) & (g652)) + ((!g704) & (g705) & (g706) & (!g707) & (g647) & (g652)) + ((g704) & (!g705) & (!g706) & (!g707) & (!g647) & (!g652)) + ((g704) & (!g705) & (!g706) & (!g707) & (!g647) & (g652)) + ((g704) & (!g705) & (!g706) & (!g707) & (g647) & (!g652)) + ((g704) & (!g705) & (!g706) & (!g707) & (g647) & (g652)) + ((g704) & (!g705) & (!g706) & (g707) & (!g647) & (!g652)) + ((g704) & (!g705) & (!g706) & (g707) & (!g647) & (g652)) + ((g704) & (!g705) & (!g706) & (g707) & (g647) & (!g652)) + ((g704) & (!g705) & (g706) & (!g707) & (!g647) & (!g652)) + ((g704) & (!g705) & (g706) & (!g707) & (g647) & (!g652)) + ((g704) & (!g705) & (g706) & (!g707) & (g647) & (g652)) + ((g704) & (!g705) & (g706) & (g707) & (!g647) & (!g652)) + ((g704) & (!g705) & (g706) & (g707) & (g647) & (!g652)) + ((g704) & (g705) & (!g706) & (!g707) & (!g647) & (!g652)) + ((g704) & (g705) & (!g706) & (!g707) & (!g647) & (g652)) + ((g704) & (g705) & (!g706) & (!g707) & (g647) & (g652)) + ((g704) & (g705) & (!g706) & (g707) & (!g647) & (!g652)) + ((g704) & (g705) & (!g706) & (g707) & (!g647) & (g652)) + ((g704) & (g705) & (g706) & (!g707) & (!g647) & (!g652)) + ((g704) & (g705) & (g706) & (!g707) & (g647) & (g652)) + ((g704) & (g705) & (g706) & (g707) & (!g647) & (!g652)));
	assign g710 = (((!sk[48]) & (g708) & (!g709)) + ((!sk[48]) & (g708) & (g709)) + ((sk[48]) & (!g708) & (g709)) + ((sk[48]) & (g708) & (!g709)));
	assign g717 = (((!g711) & (!g712) & (!g713) & (!g714) & (g715) & (g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g715) & (!g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g715) & (g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (g715) & (!g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (!g715) & (!g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (!g715) & (g716)) + ((!g711) & (!g712) & (g713) & (g714) & (!g715) & (!g716)) + ((!g711) & (!g712) & (g713) & (g714) & (g715) & (g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (g715) & (!g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (g715) & (g716)) + ((!g711) & (g712) & (!g713) & (g714) & (g715) & (!g716)) + ((!g711) & (g712) & (!g713) & (g714) & (g715) & (g716)) + ((!g711) & (g712) & (g713) & (!g714) & (g715) & (!g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (!g715) & (!g716)) + ((g711) & (!g712) & (g713) & (!g714) & (g715) & (!g716)) + ((g711) & (!g712) & (g713) & (g714) & (!g715) & (g716)) + ((g711) & (!g712) & (g713) & (g714) & (g715) & (g716)) + ((g711) & (g712) & (!g713) & (!g714) & (!g715) & (g716)) + ((g711) & (g712) & (!g713) & (!g714) & (g715) & (!g716)) + ((g711) & (g712) & (g713) & (!g714) & (!g715) & (g716)) + ((g711) & (g712) & (g713) & (!g714) & (g715) & (!g716)) + ((g711) & (g712) & (g713) & (g714) & (!g715) & (!g716)) + ((g711) & (g712) & (g713) & (g714) & (g715) & (!g716)) + ((g711) & (g712) & (g713) & (g714) & (g715) & (g716)));
	assign g718 = (((!g711) & (!g712) & (!g713) & (!g714) & (g715) & (!g716)) + ((!g711) & (!g712) & (!g713) & (!g714) & (g715) & (g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g715) & (!g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g715) & (g716)) + ((!g711) & (!g712) & (g713) & (g714) & (!g715) & (g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (!g715) & (!g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (!g715) & (g716)) + ((!g711) & (g712) & (g713) & (!g714) & (!g715) & (!g716)) + ((!g711) & (g712) & (g713) & (!g714) & (!g715) & (g716)) + ((!g711) & (g712) & (g713) & (!g714) & (g715) & (!g716)) + ((!g711) & (g712) & (g713) & (g714) & (g715) & (g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (!g715) & (g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (g715) & (!g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (g715) & (g716)) + ((g711) & (!g712) & (!g713) & (g714) & (g715) & (!g716)) + ((g711) & (!g712) & (g713) & (!g714) & (!g715) & (!g716)) + ((g711) & (!g712) & (g713) & (!g714) & (g715) & (g716)) + ((g711) & (!g712) & (g713) & (g714) & (!g715) & (g716)) + ((g711) & (!g712) & (g713) & (g714) & (g715) & (g716)) + ((g711) & (g712) & (!g713) & (!g714) & (!g715) & (!g716)) + ((g711) & (g712) & (!g713) & (!g714) & (!g715) & (g716)) + ((g711) & (g712) & (!g713) & (!g714) & (g715) & (!g716)) + ((g711) & (g712) & (!g713) & (!g714) & (g715) & (g716)) + ((g711) & (g712) & (!g713) & (g714) & (!g715) & (!g716)) + ((g711) & (g712) & (!g713) & (g714) & (g715) & (!g716)) + ((g711) & (g712) & (!g713) & (g714) & (g715) & (g716)) + ((g711) & (g712) & (g713) & (!g714) & (g715) & (!g716)) + ((g711) & (g712) & (g713) & (!g714) & (g715) & (g716)) + ((g711) & (g712) & (g713) & (g714) & (!g715) & (g716)) + ((g711) & (g712) & (g713) & (g714) & (g715) & (!g716)));
	assign g719 = (((!g711) & (!g712) & (!g713) & (!g714) & (!g715) & (!g716)) + ((!g711) & (!g712) & (!g713) & (!g714) & (g715) & (g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (g715) & (g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (!g715) & (!g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (!g715) & (g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (g715) & (g716)) + ((!g711) & (!g712) & (g713) & (g714) & (!g715) & (g716)) + ((!g711) & (!g712) & (g713) & (g714) & (g715) & (!g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (!g715) & (!g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (g715) & (!g716)) + ((!g711) & (g712) & (!g713) & (g714) & (g715) & (g716)) + ((!g711) & (g712) & (g713) & (g714) & (!g715) & (!g716)) + ((!g711) & (g712) & (g713) & (g714) & (g715) & (!g716)) + ((g711) & (!g712) & (!g713) & (g714) & (!g715) & (!g716)) + ((g711) & (!g712) & (!g713) & (g714) & (!g715) & (g716)) + ((g711) & (!g712) & (!g713) & (g714) & (g715) & (!g716)) + ((g711) & (!g712) & (g713) & (!g714) & (!g715) & (!g716)) + ((g711) & (!g712) & (g713) & (!g714) & (g715) & (g716)) + ((g711) & (!g712) & (g713) & (g714) & (!g715) & (!g716)) + ((g711) & (!g712) & (g713) & (g714) & (!g715) & (g716)) + ((g711) & (!g712) & (g713) & (g714) & (g715) & (!g716)) + ((g711) & (!g712) & (g713) & (g714) & (g715) & (g716)) + ((g711) & (g712) & (!g713) & (!g714) & (g715) & (g716)) + ((g711) & (g712) & (!g713) & (g714) & (!g715) & (!g716)) + ((g711) & (g712) & (!g713) & (g714) & (g715) & (!g716)) + ((g711) & (g712) & (!g713) & (g714) & (g715) & (g716)) + ((g711) & (g712) & (g713) & (!g714) & (!g715) & (!g716)) + ((g711) & (g712) & (g713) & (g714) & (!g715) & (!g716)) + ((g711) & (g712) & (g713) & (g714) & (!g715) & (g716)) + ((g711) & (g712) & (g713) & (g714) & (g715) & (g716)));
	assign g720 = (((!g711) & (!g712) & (!g713) & (!g714) & (!g715) & (g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (g715) & (!g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (g715) & (g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (!g715) & (g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (g715) & (g716)) + ((!g711) & (!g712) & (g713) & (g714) & (!g715) & (g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (!g715) & (!g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (!g715) & (g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (g715) & (!g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (g715) & (g716)) + ((!g711) & (g712) & (!g713) & (g714) & (g715) & (!g716)) + ((!g711) & (g712) & (!g713) & (g714) & (g715) & (g716)) + ((!g711) & (g712) & (g713) & (g714) & (!g715) & (!g716)) + ((!g711) & (g712) & (g713) & (g714) & (g715) & (!g716)) + ((!g711) & (g712) & (g713) & (g714) & (g715) & (g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (!g715) & (!g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (g715) & (g716)) + ((g711) & (!g712) & (!g713) & (g714) & (g715) & (!g716)) + ((g711) & (!g712) & (!g713) & (g714) & (g715) & (g716)) + ((g711) & (!g712) & (g713) & (!g714) & (!g715) & (g716)) + ((g711) & (!g712) & (g713) & (!g714) & (g715) & (!g716)) + ((g711) & (!g712) & (g713) & (g714) & (g715) & (!g716)) + ((g711) & (g712) & (!g713) & (!g714) & (!g715) & (g716)) + ((g711) & (g712) & (!g713) & (!g714) & (g715) & (g716)) + ((g711) & (g712) & (!g713) & (g714) & (g715) & (!g716)) + ((g711) & (g712) & (!g713) & (g714) & (g715) & (g716)) + ((g711) & (g712) & (g713) & (!g714) & (!g715) & (g716)) + ((g711) & (g712) & (g713) & (g714) & (!g715) & (!g716)));
	assign g723 = (((!g717) & (!g718) & (!g719) & (!g720) & (!g721) & (!g722)) + ((!g717) & (!g718) & (!g719) & (g720) & (!g721) & (!g722)) + ((!g717) & (!g718) & (!g719) & (g720) & (g721) & (g722)) + ((!g717) & (!g718) & (g719) & (!g720) & (!g721) & (!g722)) + ((!g717) & (!g718) & (g719) & (!g720) & (!g721) & (g722)) + ((!g717) & (!g718) & (g719) & (g720) & (!g721) & (!g722)) + ((!g717) & (!g718) & (g719) & (g720) & (!g721) & (g722)) + ((!g717) & (!g718) & (g719) & (g720) & (g721) & (g722)) + ((!g717) & (g718) & (!g719) & (!g720) & (!g721) & (!g722)) + ((!g717) & (g718) & (!g719) & (!g720) & (g721) & (!g722)) + ((!g717) & (g718) & (!g719) & (g720) & (!g721) & (!g722)) + ((!g717) & (g718) & (!g719) & (g720) & (g721) & (!g722)) + ((!g717) & (g718) & (!g719) & (g720) & (g721) & (g722)) + ((!g717) & (g718) & (g719) & (!g720) & (!g721) & (!g722)) + ((!g717) & (g718) & (g719) & (!g720) & (!g721) & (g722)) + ((!g717) & (g718) & (g719) & (!g720) & (g721) & (!g722)) + ((!g717) & (g718) & (g719) & (g720) & (!g721) & (!g722)) + ((!g717) & (g718) & (g719) & (g720) & (!g721) & (g722)) + ((!g717) & (g718) & (g719) & (g720) & (g721) & (!g722)) + ((!g717) & (g718) & (g719) & (g720) & (g721) & (g722)) + ((g717) & (!g718) & (!g719) & (g720) & (g721) & (g722)) + ((g717) & (!g718) & (g719) & (!g720) & (!g721) & (g722)) + ((g717) & (!g718) & (g719) & (g720) & (!g721) & (g722)) + ((g717) & (!g718) & (g719) & (g720) & (g721) & (g722)) + ((g717) & (g718) & (!g719) & (!g720) & (g721) & (!g722)) + ((g717) & (g718) & (!g719) & (g720) & (g721) & (!g722)) + ((g717) & (g718) & (!g719) & (g720) & (g721) & (g722)) + ((g717) & (g718) & (g719) & (!g720) & (!g721) & (g722)) + ((g717) & (g718) & (g719) & (!g720) & (g721) & (!g722)) + ((g717) & (g718) & (g719) & (g720) & (!g721) & (g722)) + ((g717) & (g718) & (g719) & (g720) & (g721) & (!g722)) + ((g717) & (g718) & (g719) & (g720) & (g721) & (g722)));
	assign g725 = (((!sk[54]) & (g723) & (!g724)) + ((!sk[54]) & (g723) & (g724)) + ((sk[54]) & (!g723) & (g724)) + ((sk[54]) & (g723) & (!g724)));
	assign g726 = (((!g711) & (!g712) & (!g713) & (!g714) & (!g721) & (g715)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g721) & (!g715)) + ((!g711) & (!g712) & (!g713) & (g714) & (g721) & (!g715)) + ((!g711) & (!g712) & (g713) & (!g714) & (g721) & (g715)) + ((!g711) & (!g712) & (g713) & (g714) & (!g721) & (g715)) + ((!g711) & (!g712) & (g713) & (g714) & (g721) & (!g715)) + ((!g711) & (g712) & (!g713) & (!g714) & (!g721) & (g715)) + ((!g711) & (g712) & (!g713) & (!g714) & (g721) & (!g715)) + ((!g711) & (g712) & (!g713) & (!g714) & (g721) & (g715)) + ((!g711) & (g712) & (g713) & (!g714) & (g721) & (g715)) + ((!g711) & (g712) & (g713) & (g714) & (g721) & (g715)) + ((g711) & (!g712) & (!g713) & (!g714) & (!g721) & (!g715)) + ((g711) & (!g712) & (!g713) & (!g714) & (g721) & (g715)) + ((g711) & (!g712) & (!g713) & (g714) & (!g721) & (!g715)) + ((g711) & (!g712) & (!g713) & (g714) & (g721) & (!g715)) + ((g711) & (!g712) & (g713) & (!g714) & (g721) & (!g715)) + ((g711) & (!g712) & (g713) & (!g714) & (g721) & (g715)) + ((g711) & (!g712) & (g713) & (g714) & (g721) & (!g715)) + ((g711) & (!g712) & (g713) & (g714) & (g721) & (g715)) + ((g711) & (g712) & (!g713) & (!g714) & (g721) & (!g715)) + ((g711) & (g712) & (!g713) & (!g714) & (g721) & (g715)) + ((g711) & (g712) & (!g713) & (g714) & (g721) & (g715)) + ((g711) & (g712) & (g713) & (!g714) & (!g721) & (!g715)) + ((g711) & (g712) & (g713) & (!g714) & (!g721) & (g715)) + ((g711) & (g712) & (g713) & (!g714) & (g721) & (!g715)) + ((g711) & (g712) & (g713) & (g714) & (!g721) & (g715)) + ((g711) & (g712) & (g713) & (g714) & (g721) & (!g715)));
	assign g727 = (((!g711) & (!g712) & (!g713) & (!g714) & (!g721) & (g715)) + ((!g711) & (!g712) & (!g713) & (!g714) & (g721) & (!g715)) + ((!g711) & (!g712) & (!g713) & (!g714) & (g721) & (g715)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g721) & (!g715)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g721) & (g715)) + ((!g711) & (!g712) & (!g713) & (g714) & (g721) & (g715)) + ((!g711) & (!g712) & (g713) & (!g714) & (g721) & (!g715)) + ((!g711) & (!g712) & (g713) & (g714) & (!g721) & (!g715)) + ((!g711) & (!g712) & (g713) & (g714) & (!g721) & (g715)) + ((!g711) & (!g712) & (g713) & (g714) & (g721) & (g715)) + ((!g711) & (g712) & (!g713) & (!g714) & (g721) & (g715)) + ((!g711) & (g712) & (!g713) & (g714) & (!g721) & (!g715)) + ((!g711) & (g712) & (!g713) & (g714) & (g721) & (!g715)) + ((!g711) & (g712) & (g713) & (!g714) & (g721) & (!g715)) + ((!g711) & (g712) & (g713) & (!g714) & (g721) & (g715)) + ((!g711) & (g712) & (g713) & (g714) & (!g721) & (!g715)) + ((g711) & (!g712) & (!g713) & (!g714) & (!g721) & (!g715)) + ((g711) & (!g712) & (!g713) & (g714) & (!g721) & (!g715)) + ((g711) & (!g712) & (!g713) & (g714) & (!g721) & (g715)) + ((g711) & (!g712) & (g713) & (!g714) & (!g721) & (g715)) + ((g711) & (!g712) & (g713) & (!g714) & (g721) & (g715)) + ((g711) & (!g712) & (g713) & (g714) & (!g721) & (!g715)) + ((g711) & (!g712) & (g713) & (g714) & (!g721) & (g715)) + ((g711) & (g712) & (!g713) & (g714) & (!g721) & (!g715)) + ((g711) & (g712) & (!g713) & (g714) & (g721) & (g715)) + ((g711) & (g712) & (g713) & (!g714) & (!g721) & (!g715)) + ((g711) & (g712) & (g713) & (!g714) & (!g721) & (g715)) + ((g711) & (g712) & (g713) & (!g714) & (g721) & (g715)) + ((g711) & (g712) & (g713) & (g714) & (!g721) & (!g715)) + ((g711) & (g712) & (g713) & (g714) & (!g721) & (g715)) + ((g711) & (g712) & (g713) & (g714) & (g721) & (!g715)));
	assign g728 = (((!g711) & (!g712) & (!g713) & (!g714) & (!g721) & (g715)) + ((!g711) & (!g712) & (!g713) & (g714) & (g721) & (!g715)) + ((!g711) & (!g712) & (g713) & (!g714) & (!g721) & (!g715)) + ((!g711) & (!g712) & (g713) & (!g714) & (g721) & (!g715)) + ((!g711) & (!g712) & (g713) & (g714) & (!g721) & (g715)) + ((!g711) & (!g712) & (g713) & (g714) & (g721) & (!g715)) + ((!g711) & (!g712) & (g713) & (g714) & (g721) & (g715)) + ((!g711) & (g712) & (!g713) & (!g714) & (!g721) & (!g715)) + ((!g711) & (g712) & (!g713) & (!g714) & (g721) & (!g715)) + ((!g711) & (g712) & (!g713) & (g714) & (!g721) & (!g715)) + ((!g711) & (g712) & (!g713) & (g714) & (g721) & (g715)) + ((!g711) & (g712) & (g713) & (!g714) & (g721) & (g715)) + ((!g711) & (g712) & (g713) & (g714) & (!g721) & (g715)) + ((!g711) & (g712) & (g713) & (g714) & (g721) & (!g715)) + ((g711) & (!g712) & (!g713) & (!g714) & (g721) & (g715)) + ((g711) & (!g712) & (!g713) & (g714) & (!g721) & (!g715)) + ((g711) & (!g712) & (!g713) & (g714) & (g721) & (!g715)) + ((g711) & (!g712) & (g713) & (!g714) & (!g721) & (!g715)) + ((g711) & (!g712) & (g713) & (!g714) & (!g721) & (g715)) + ((g711) & (!g712) & (g713) & (!g714) & (g721) & (!g715)) + ((g711) & (!g712) & (g713) & (!g714) & (g721) & (g715)) + ((g711) & (!g712) & (g713) & (g714) & (g721) & (!g715)) + ((g711) & (g712) & (!g713) & (!g714) & (!g721) & (g715)) + ((g711) & (g712) & (!g713) & (!g714) & (g721) & (g715)) + ((g711) & (g712) & (!g713) & (g714) & (!g721) & (g715)) + ((g711) & (g712) & (g713) & (!g714) & (!g721) & (!g715)) + ((g711) & (g712) & (g713) & (!g714) & (!g721) & (g715)) + ((g711) & (g712) & (g713) & (!g714) & (g721) & (g715)) + ((g711) & (g712) & (g713) & (g714) & (!g721) & (!g715)) + ((g711) & (g712) & (g713) & (g714) & (!g721) & (g715)) + ((g711) & (g712) & (g713) & (g714) & (g721) & (!g715)) + ((g711) & (g712) & (g713) & (g714) & (g721) & (g715)));
	assign g729 = (((!g711) & (!g712) & (!g713) & (!g714) & (g721) & (!g715)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g721) & (!g715)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g721) & (g715)) + ((!g711) & (!g712) & (g713) & (!g714) & (g721) & (g715)) + ((!g711) & (!g712) & (g713) & (g714) & (!g721) & (g715)) + ((!g711) & (g712) & (!g713) & (!g714) & (!g721) & (!g715)) + ((!g711) & (g712) & (!g713) & (!g714) & (g721) & (!g715)) + ((!g711) & (g712) & (!g713) & (g714) & (!g721) & (g715)) + ((!g711) & (g712) & (g713) & (!g714) & (!g721) & (g715)) + ((!g711) & (g712) & (g713) & (!g714) & (g721) & (!g715)) + ((!g711) & (g712) & (g713) & (!g714) & (g721) & (g715)) + ((!g711) & (g712) & (g713) & (g714) & (g721) & (!g715)) + ((!g711) & (g712) & (g713) & (g714) & (g721) & (g715)) + ((g711) & (!g712) & (!g713) & (!g714) & (!g721) & (!g715)) + ((g711) & (!g712) & (!g713) & (g714) & (!g721) & (!g715)) + ((g711) & (!g712) & (!g713) & (g714) & (!g721) & (g715)) + ((g711) & (!g712) & (!g713) & (g714) & (g721) & (!g715)) + ((g711) & (!g712) & (g713) & (!g714) & (!g721) & (!g715)) + ((g711) & (!g712) & (g713) & (!g714) & (g721) & (g715)) + ((g711) & (!g712) & (g713) & (g714) & (g721) & (!g715)) + ((g711) & (g712) & (!g713) & (!g714) & (!g721) & (!g715)) + ((g711) & (g712) & (!g713) & (g714) & (!g721) & (!g715)) + ((g711) & (g712) & (!g713) & (g714) & (g721) & (!g715)) + ((g711) & (g712) & (!g713) & (g714) & (g721) & (g715)) + ((g711) & (g712) & (g713) & (g714) & (!g721) & (g715)) + ((g711) & (g712) & (g713) & (g714) & (g721) & (g715)));
	assign g730 = (((!g726) & (!g727) & (!g728) & (!g729) & (!g716) & (!g722)) + ((!g726) & (!g727) & (!g728) & (!g729) & (g716) & (!g722)) + ((!g726) & (!g727) & (!g728) & (g729) & (!g716) & (!g722)) + ((!g726) & (!g727) & (!g728) & (g729) & (g716) & (!g722)) + ((!g726) & (!g727) & (!g728) & (g729) & (g716) & (g722)) + ((!g726) & (!g727) & (g728) & (!g729) & (!g716) & (!g722)) + ((!g726) & (!g727) & (g728) & (!g729) & (!g716) & (g722)) + ((!g726) & (!g727) & (g728) & (!g729) & (g716) & (!g722)) + ((!g726) & (!g727) & (g728) & (g729) & (!g716) & (!g722)) + ((!g726) & (!g727) & (g728) & (g729) & (!g716) & (g722)) + ((!g726) & (!g727) & (g728) & (g729) & (g716) & (!g722)) + ((!g726) & (!g727) & (g728) & (g729) & (g716) & (g722)) + ((!g726) & (g727) & (!g728) & (!g729) & (!g716) & (!g722)) + ((!g726) & (g727) & (!g728) & (g729) & (!g716) & (!g722)) + ((!g726) & (g727) & (!g728) & (g729) & (g716) & (g722)) + ((!g726) & (g727) & (g728) & (!g729) & (!g716) & (!g722)) + ((!g726) & (g727) & (g728) & (!g729) & (!g716) & (g722)) + ((!g726) & (g727) & (g728) & (g729) & (!g716) & (!g722)) + ((!g726) & (g727) & (g728) & (g729) & (!g716) & (g722)) + ((!g726) & (g727) & (g728) & (g729) & (g716) & (g722)) + ((g726) & (!g727) & (!g728) & (!g729) & (g716) & (!g722)) + ((g726) & (!g727) & (!g728) & (g729) & (g716) & (!g722)) + ((g726) & (!g727) & (!g728) & (g729) & (g716) & (g722)) + ((g726) & (!g727) & (g728) & (!g729) & (!g716) & (g722)) + ((g726) & (!g727) & (g728) & (!g729) & (g716) & (!g722)) + ((g726) & (!g727) & (g728) & (g729) & (!g716) & (g722)) + ((g726) & (!g727) & (g728) & (g729) & (g716) & (!g722)) + ((g726) & (!g727) & (g728) & (g729) & (g716) & (g722)) + ((g726) & (g727) & (!g728) & (g729) & (g716) & (g722)) + ((g726) & (g727) & (g728) & (!g729) & (!g716) & (g722)) + ((g726) & (g727) & (g728) & (g729) & (!g716) & (g722)) + ((g726) & (g727) & (g728) & (g729) & (g716) & (g722)));
	assign g732 = (((!g730) & (sk[60]) & (g731)) + ((g730) & (!sk[60]) & (!g731)) + ((g730) & (!sk[60]) & (g731)) + ((g730) & (sk[60]) & (!g731)));
	assign g733 = (((!g715) & (!g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((!g715) & (!g712) & (!g713) & (!g714) & (g721) & (g716)) + ((!g715) & (!g712) & (!g713) & (g714) & (!g721) & (g716)) + ((!g715) & (!g712) & (!g713) & (g714) & (g721) & (!g716)) + ((!g715) & (!g712) & (!g713) & (g714) & (g721) & (g716)) + ((!g715) & (!g712) & (g713) & (!g714) & (!g721) & (g716)) + ((!g715) & (!g712) & (g713) & (g714) & (!g721) & (!g716)) + ((!g715) & (!g712) & (g713) & (g714) & (g721) & (!g716)) + ((!g715) & (g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((!g715) & (g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((!g715) & (g712) & (!g713) & (g714) & (!g721) & (g716)) + ((!g715) & (g712) & (g713) & (!g714) & (!g721) & (!g716)) + ((!g715) & (g712) & (g713) & (!g714) & (!g721) & (g716)) + ((!g715) & (g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g715) & (g712) & (g713) & (!g714) & (g721) & (g716)) + ((g715) & (!g712) & (!g713) & (g714) & (!g721) & (g716)) + ((g715) & (!g712) & (!g713) & (g714) & (g721) & (g716)) + ((g715) & (g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((g715) & (g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((g715) & (g712) & (!g713) & (g714) & (g721) & (!g716)) + ((g715) & (g712) & (g713) & (g714) & (!g721) & (!g716)) + ((g715) & (g712) & (g713) & (g714) & (!g721) & (g716)));
	assign g734 = (((!g715) & (!g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((!g715) & (!g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((!g715) & (!g712) & (!g713) & (g714) & (g721) & (g716)) + ((!g715) & (!g712) & (g713) & (!g714) & (!g721) & (!g716)) + ((!g715) & (!g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g715) & (!g712) & (g713) & (g714) & (!g721) & (g716)) + ((!g715) & (g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((!g715) & (g712) & (!g713) & (!g714) & (g721) & (g716)) + ((!g715) & (g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((!g715) & (g712) & (!g713) & (g714) & (!g721) & (g716)) + ((!g715) & (g712) & (!g713) & (g714) & (g721) & (g716)) + ((!g715) & (g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g715) & (g712) & (g713) & (!g714) & (g721) & (g716)) + ((!g715) & (g712) & (g713) & (g714) & (g721) & (!g716)) + ((g715) & (!g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((g715) & (!g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((g715) & (!g712) & (!g713) & (!g714) & (g721) & (g716)) + ((g715) & (!g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((g715) & (!g712) & (!g713) & (g714) & (!g721) & (g716)) + ((g715) & (!g712) & (!g713) & (g714) & (g721) & (!g716)) + ((g715) & (!g712) & (g713) & (g714) & (!g721) & (!g716)) + ((g715) & (g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((g715) & (g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((g715) & (g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((g715) & (g712) & (!g713) & (g714) & (g721) & (!g716)) + ((g715) & (g712) & (!g713) & (g714) & (g721) & (g716)) + ((g715) & (g712) & (g713) & (!g714) & (!g721) & (!g716)) + ((g715) & (g712) & (g713) & (!g714) & (g721) & (!g716)) + ((g715) & (g712) & (g713) & (g714) & (!g721) & (g716)) + ((g715) & (g712) & (g713) & (g714) & (g721) & (g716)));
	assign g735 = (((!g715) & (!g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((!g715) & (!g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((!g715) & (!g712) & (!g713) & (g714) & (!g721) & (g716)) + ((!g715) & (!g712) & (g713) & (!g714) & (!g721) & (g716)) + ((!g715) & (!g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g715) & (!g712) & (g713) & (g714) & (!g721) & (g716)) + ((!g715) & (g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((!g715) & (g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((!g715) & (g712) & (!g713) & (g714) & (g721) & (!g716)) + ((!g715) & (g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g715) & (g712) & (g713) & (g714) & (!g721) & (!g716)) + ((!g715) & (g712) & (g713) & (g714) & (g721) & (!g716)) + ((g715) & (!g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((g715) & (!g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((g715) & (!g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((g715) & (!g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((g715) & (!g712) & (!g713) & (g714) & (!g721) & (g716)) + ((g715) & (!g712) & (!g713) & (g714) & (g721) & (!g716)) + ((g715) & (!g712) & (!g713) & (g714) & (g721) & (g716)) + ((g715) & (!g712) & (g713) & (!g714) & (!g721) & (g716)) + ((g715) & (!g712) & (g713) & (!g714) & (g721) & (!g716)) + ((g715) & (!g712) & (g713) & (g714) & (!g721) & (!g716)) + ((g715) & (!g712) & (g713) & (g714) & (g721) & (g716)) + ((g715) & (g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((g715) & (g712) & (!g713) & (!g714) & (g721) & (g716)) + ((g715) & (g712) & (g713) & (!g714) & (g721) & (g716)) + ((g715) & (g712) & (g713) & (g714) & (!g721) & (!g716)) + ((g715) & (g712) & (g713) & (g714) & (!g721) & (g716)) + ((g715) & (g712) & (g713) & (g714) & (g721) & (g716)));
	assign g736 = (((!g715) & (!g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((!g715) & (!g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((!g715) & (!g712) & (!g713) & (!g714) & (g721) & (g716)) + ((!g715) & (!g712) & (!g713) & (g714) & (!g721) & (g716)) + ((!g715) & (!g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g715) & (!g712) & (g713) & (g714) & (g721) & (g716)) + ((!g715) & (g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((!g715) & (g712) & (!g713) & (g714) & (!g721) & (g716)) + ((!g715) & (g712) & (!g713) & (g714) & (g721) & (g716)) + ((!g715) & (g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g715) & (g712) & (g713) & (!g714) & (g721) & (g716)) + ((!g715) & (g712) & (g713) & (g714) & (!g721) & (!g716)) + ((!g715) & (g712) & (g713) & (g714) & (!g721) & (g716)) + ((!g715) & (g712) & (g713) & (g714) & (g721) & (!g716)) + ((!g715) & (g712) & (g713) & (g714) & (g721) & (g716)) + ((g715) & (!g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((g715) & (!g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((g715) & (!g712) & (!g713) & (!g714) & (g721) & (g716)) + ((g715) & (!g712) & (!g713) & (g714) & (g721) & (g716)) + ((g715) & (!g712) & (g713) & (!g714) & (!g721) & (g716)) + ((g715) & (!g712) & (g713) & (!g714) & (g721) & (!g716)) + ((g715) & (!g712) & (g713) & (g714) & (g721) & (!g716)) + ((g715) & (g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((g715) & (g712) & (!g713) & (g714) & (!g721) & (g716)) + ((g715) & (g712) & (!g713) & (g714) & (g721) & (!g716)) + ((g715) & (g712) & (g713) & (!g714) & (g721) & (g716)) + ((g715) & (g712) & (g713) & (g714) & (!g721) & (!g716)));
	assign g737 = (((!g733) & (!g734) & (!g735) & (!g736) & (!g711) & (g722)) + ((!g733) & (!g734) & (!g735) & (!g736) & (g711) & (!g722)) + ((!g733) & (!g734) & (!g735) & (!g736) & (g711) & (g722)) + ((!g733) & (!g734) & (!g735) & (g736) & (!g711) & (g722)) + ((!g733) & (!g734) & (!g735) & (g736) & (g711) & (!g722)) + ((!g733) & (!g734) & (g735) & (!g736) & (g711) & (!g722)) + ((!g733) & (!g734) & (g735) & (!g736) & (g711) & (g722)) + ((!g733) & (!g734) & (g735) & (g736) & (g711) & (!g722)) + ((!g733) & (g734) & (!g735) & (!g736) & (!g711) & (g722)) + ((!g733) & (g734) & (!g735) & (!g736) & (g711) & (g722)) + ((!g733) & (g734) & (!g735) & (g736) & (!g711) & (g722)) + ((!g733) & (g734) & (g735) & (!g736) & (g711) & (g722)) + ((g733) & (!g734) & (!g735) & (!g736) & (!g711) & (!g722)) + ((g733) & (!g734) & (!g735) & (!g736) & (!g711) & (g722)) + ((g733) & (!g734) & (!g735) & (!g736) & (g711) & (!g722)) + ((g733) & (!g734) & (!g735) & (!g736) & (g711) & (g722)) + ((g733) & (!g734) & (!g735) & (g736) & (!g711) & (!g722)) + ((g733) & (!g734) & (!g735) & (g736) & (!g711) & (g722)) + ((g733) & (!g734) & (!g735) & (g736) & (g711) & (!g722)) + ((g733) & (!g734) & (g735) & (!g736) & (!g711) & (!g722)) + ((g733) & (!g734) & (g735) & (!g736) & (g711) & (!g722)) + ((g733) & (!g734) & (g735) & (!g736) & (g711) & (g722)) + ((g733) & (!g734) & (g735) & (g736) & (!g711) & (!g722)) + ((g733) & (!g734) & (g735) & (g736) & (g711) & (!g722)) + ((g733) & (g734) & (!g735) & (!g736) & (!g711) & (!g722)) + ((g733) & (g734) & (!g735) & (!g736) & (!g711) & (g722)) + ((g733) & (g734) & (!g735) & (!g736) & (g711) & (g722)) + ((g733) & (g734) & (!g735) & (g736) & (!g711) & (!g722)) + ((g733) & (g734) & (!g735) & (g736) & (!g711) & (g722)) + ((g733) & (g734) & (g735) & (!g736) & (!g711) & (!g722)) + ((g733) & (g734) & (g735) & (!g736) & (g711) & (g722)) + ((g733) & (g734) & (g735) & (g736) & (!g711) & (!g722)));
	assign g739 = (((!g737) & (sk[66]) & (g738)) + ((g737) & (!sk[66]) & (!g738)) + ((g737) & (!sk[66]) & (g738)) + ((g737) & (sk[66]) & (!g738)));
	assign g740 = (((!g711) & (!g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (g721) & (g716)) + ((!g711) & (!g712) & (g713) & (g714) & (!g721) & (!g716)) + ((!g711) & (!g712) & (g713) & (g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (g713) & (g714) & (g721) & (g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (g712) & (g713) & (!g714) & (!g721) & (!g716)) + ((!g711) & (g712) & (g713) & (g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((g711) & (!g712) & (g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (g713) & (!g714) & (!g721) & (g716)) + ((g711) & (!g712) & (g713) & (!g714) & (g721) & (!g716)) + ((g711) & (!g712) & (g713) & (g714) & (!g721) & (g716)) + ((g711) & (g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((g711) & (g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((g711) & (g712) & (!g713) & (g714) & (g721) & (!g716)) + ((g711) & (g712) & (g713) & (!g714) & (!g721) & (g716)) + ((g711) & (g712) & (g713) & (!g714) & (g721) & (g716)));
	assign g741 = (((!g711) & (!g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (!g713) & (!g714) & (g721) & (g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (g713) & (g714) & (!g721) & (!g716)) + ((!g711) & (!g712) & (g713) & (g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (g713) & (g714) & (g721) & (g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (g721) & (g716)) + ((!g711) & (g712) & (!g713) & (g714) & (g721) & (g716)) + ((!g711) & (g712) & (g713) & (!g714) & (!g721) & (!g716)) + ((!g711) & (g712) & (g713) & (!g714) & (!g721) & (g716)) + ((!g711) & (g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (g712) & (g713) & (g714) & (!g721) & (g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((g711) & (!g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (!g713) & (g714) & (!g721) & (g716)) + ((g711) & (!g712) & (!g713) & (g714) & (g721) & (g716)) + ((g711) & (!g712) & (g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (g713) & (!g714) & (!g721) & (g716)) + ((g711) & (!g712) & (g713) & (!g714) & (g721) & (g716)) + ((g711) & (!g712) & (g713) & (g714) & (!g721) & (g716)) + ((g711) & (g712) & (!g713) & (g714) & (!g721) & (g716)) + ((g711) & (g712) & (!g713) & (g714) & (g721) & (!g716)) + ((g711) & (g712) & (g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (g712) & (g713) & (g714) & (!g721) & (!g716)));
	assign g742 = (((!g711) & (!g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (!g713) & (!g714) & (g721) & (g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (g713) & (!g714) & (g721) & (g716)) + ((!g711) & (!g712) & (g713) & (g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (g713) & (g714) & (g721) & (g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (g721) & (g716)) + ((!g711) & (g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((!g711) & (g712) & (!g713) & (g714) & (!g721) & (g716)) + ((!g711) & (g712) & (g713) & (!g714) & (!g721) & (g716)) + ((!g711) & (g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (g712) & (g713) & (g714) & (g721) & (g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (g721) & (g716)) + ((g711) & (!g712) & (!g713) & (g714) & (g721) & (g716)) + ((g711) & (!g712) & (g713) & (g714) & (!g721) & (!g716)) + ((g711) & (g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((g711) & (g712) & (!g713) & (g714) & (g721) & (g716)) + ((g711) & (g712) & (g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (g712) & (g713) & (!g714) & (!g721) & (g716)) + ((g711) & (g712) & (g713) & (!g714) & (g721) & (g716)) + ((g711) & (g712) & (g713) & (g714) & (!g721) & (!g716)) + ((g711) & (g712) & (g713) & (g714) & (g721) & (g716)));
	assign g743 = (((!g711) & (!g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (!g713) & (g714) & (g721) & (g716)) + ((!g711) & (!g712) & (g713) & (g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (g713) & (g714) & (g721) & (g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (!g721) & (!g716)) + ((!g711) & (g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (g712) & (!g713) & (g714) & (!g721) & (!g716)) + ((!g711) & (g712) & (!g713) & (g714) & (!g721) & (g716)) + ((!g711) & (g712) & (!g713) & (g714) & (g721) & (!g716)) + ((!g711) & (g712) & (g713) & (!g714) & (!g721) & (!g716)) + ((!g711) & (g712) & (g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (g712) & (g713) & (!g714) & (g721) & (g716)) + ((g711) & (!g712) & (!g713) & (!g714) & (g721) & (g716)) + ((g711) & (!g712) & (!g713) & (g714) & (g721) & (!g716)) + ((g711) & (!g712) & (g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (g713) & (!g714) & (g721) & (!g716)) + ((g711) & (!g712) & (g713) & (!g714) & (g721) & (g716)) + ((g711) & (!g712) & (g713) & (g714) & (!g721) & (g716)) + ((g711) & (!g712) & (g713) & (g714) & (g721) & (!g716)) + ((g711) & (!g712) & (g713) & (g714) & (g721) & (g716)) + ((g711) & (g712) & (!g713) & (!g714) & (!g721) & (g716)) + ((g711) & (g712) & (!g713) & (!g714) & (g721) & (!g716)) + ((g711) & (g712) & (g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (g712) & (g713) & (!g714) & (!g721) & (g716)) + ((g711) & (g712) & (g713) & (g714) & (g721) & (g716)));
	assign g744 = (((!g740) & (!g741) & (!g742) & (!g743) & (!g722) & (g715)) + ((!g740) & (!g741) & (!g742) & (!g743) & (g722) & (!g715)) + ((!g740) & (!g741) & (!g742) & (!g743) & (g722) & (g715)) + ((!g740) & (!g741) & (!g742) & (g743) & (!g722) & (g715)) + ((!g740) & (!g741) & (!g742) & (g743) & (g722) & (!g715)) + ((!g740) & (!g741) & (g742) & (!g743) & (g722) & (!g715)) + ((!g740) & (!g741) & (g742) & (!g743) & (g722) & (g715)) + ((!g740) & (!g741) & (g742) & (g743) & (g722) & (!g715)) + ((!g740) & (g741) & (!g742) & (!g743) & (!g722) & (g715)) + ((!g740) & (g741) & (!g742) & (!g743) & (g722) & (g715)) + ((!g740) & (g741) & (!g742) & (g743) & (!g722) & (g715)) + ((!g740) & (g741) & (g742) & (!g743) & (g722) & (g715)) + ((g740) & (!g741) & (!g742) & (!g743) & (!g722) & (!g715)) + ((g740) & (!g741) & (!g742) & (!g743) & (!g722) & (g715)) + ((g740) & (!g741) & (!g742) & (!g743) & (g722) & (!g715)) + ((g740) & (!g741) & (!g742) & (!g743) & (g722) & (g715)) + ((g740) & (!g741) & (!g742) & (g743) & (!g722) & (!g715)) + ((g740) & (!g741) & (!g742) & (g743) & (!g722) & (g715)) + ((g740) & (!g741) & (!g742) & (g743) & (g722) & (!g715)) + ((g740) & (!g741) & (g742) & (!g743) & (!g722) & (!g715)) + ((g740) & (!g741) & (g742) & (!g743) & (g722) & (!g715)) + ((g740) & (!g741) & (g742) & (!g743) & (g722) & (g715)) + ((g740) & (!g741) & (g742) & (g743) & (!g722) & (!g715)) + ((g740) & (!g741) & (g742) & (g743) & (g722) & (!g715)) + ((g740) & (g741) & (!g742) & (!g743) & (!g722) & (!g715)) + ((g740) & (g741) & (!g742) & (!g743) & (!g722) & (g715)) + ((g740) & (g741) & (!g742) & (!g743) & (g722) & (g715)) + ((g740) & (g741) & (!g742) & (g743) & (!g722) & (!g715)) + ((g740) & (g741) & (!g742) & (g743) & (!g722) & (g715)) + ((g740) & (g741) & (g742) & (!g743) & (!g722) & (!g715)) + ((g740) & (g741) & (g742) & (!g743) & (g722) & (g715)) + ((g740) & (g741) & (g742) & (g743) & (!g722) & (!g715)));
	assign g746 = (((!sk[72]) & (g744) & (!g745)) + ((!sk[72]) & (g744) & (g745)) + ((sk[72]) & (!g744) & (g745)) + ((sk[72]) & (g744) & (!g745)));
	assign g747 = (((!g711) & (!g712) & (!g715) & (!g722) & (!g721) & (g716)) + ((!g711) & (!g712) & (g715) & (!g722) & (!g721) & (g716)) + ((!g711) & (!g712) & (g715) & (!g722) & (g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (!g722) & (g721) & (g716)) + ((!g711) & (!g712) & (g715) & (g722) & (!g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (g722) & (g721) & (!g716)) + ((!g711) & (g712) & (!g715) & (!g722) & (!g721) & (!g716)) + ((!g711) & (g712) & (!g715) & (!g722) & (!g721) & (g716)) + ((!g711) & (g712) & (!g715) & (g722) & (!g721) & (!g716)) + ((!g711) & (g712) & (!g715) & (g722) & (!g721) & (g716)) + ((!g711) & (g712) & (!g715) & (g722) & (g721) & (g716)) + ((!g711) & (g712) & (g715) & (g722) & (!g721) & (g716)) + ((!g711) & (g712) & (g715) & (g722) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g722) & (!g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g722) & (!g721) & (g716)) + ((g711) & (!g712) & (!g715) & (g722) & (!g721) & (g716)) + ((g711) & (!g712) & (g715) & (!g722) & (g721) & (!g716)) + ((g711) & (!g712) & (g715) & (g722) & (!g721) & (!g716)) + ((g711) & (!g712) & (g715) & (g722) & (!g721) & (g716)) + ((g711) & (!g712) & (g715) & (g722) & (g721) & (!g716)) + ((g711) & (g712) & (!g715) & (!g722) & (!g721) & (!g716)) + ((g711) & (g712) & (!g715) & (!g722) & (g721) & (!g716)) + ((g711) & (g712) & (!g715) & (g722) & (g721) & (!g716)) + ((g711) & (g712) & (g715) & (!g722) & (!g721) & (!g716)) + ((g711) & (g712) & (g715) & (!g722) & (!g721) & (g716)) + ((g711) & (g712) & (g715) & (g722) & (!g721) & (g716)));
	assign g748 = (((!g711) & (!g712) & (!g715) & (!g722) & (!g721) & (!g716)) + ((!g711) & (!g712) & (!g715) & (!g722) & (!g721) & (g716)) + ((!g711) & (!g712) & (!g715) & (!g722) & (g721) & (!g716)) + ((!g711) & (!g712) & (!g715) & (!g722) & (g721) & (g716)) + ((!g711) & (!g712) & (!g715) & (g722) & (!g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (!g722) & (!g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (!g722) & (g721) & (g716)) + ((!g711) & (!g712) & (g715) & (g722) & (!g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (g722) & (g721) & (g716)) + ((!g711) & (g712) & (!g715) & (!g722) & (!g721) & (g716)) + ((!g711) & (g712) & (!g715) & (g722) & (g721) & (!g716)) + ((!g711) & (g712) & (g715) & (!g722) & (!g721) & (!g716)) + ((!g711) & (g712) & (g715) & (!g722) & (!g721) & (g716)) + ((!g711) & (g712) & (g715) & (!g722) & (g721) & (!g716)) + ((!g711) & (g712) & (g715) & (!g722) & (g721) & (g716)) + ((!g711) & (g712) & (g715) & (g722) & (!g721) & (!g716)) + ((!g711) & (g712) & (g715) & (g722) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g722) & (!g721) & (g716)) + ((g711) & (!g712) & (!g715) & (!g722) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g722) & (g721) & (g716)) + ((g711) & (!g712) & (!g715) & (g722) & (!g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (g722) & (g721) & (g716)) + ((g711) & (!g712) & (g715) & (!g722) & (g721) & (!g716)) + ((g711) & (!g712) & (g715) & (!g722) & (g721) & (g716)) + ((g711) & (!g712) & (g715) & (g722) & (!g721) & (g716)) + ((g711) & (g712) & (!g715) & (!g722) & (g721) & (!g716)) + ((g711) & (g712) & (!g715) & (!g722) & (g721) & (g716)) + ((g711) & (g712) & (!g715) & (g722) & (!g721) & (!g716)) + ((g711) & (g712) & (!g715) & (g722) & (!g721) & (g716)) + ((g711) & (g712) & (g715) & (!g722) & (g721) & (!g716)) + ((g711) & (g712) & (g715) & (!g722) & (g721) & (g716)) + ((g711) & (g712) & (g715) & (g722) & (!g721) & (g716)));
	assign g749 = (((!g711) & (!g712) & (!g715) & (!g722) & (!g721) & (!g716)) + ((!g711) & (!g712) & (!g715) & (!g722) & (!g721) & (g716)) + ((!g711) & (!g712) & (g715) & (!g722) & (!g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (!g722) & (g721) & (g716)) + ((!g711) & (!g712) & (g715) & (g722) & (!g721) & (g716)) + ((!g711) & (g712) & (!g715) & (g722) & (!g721) & (!g716)) + ((!g711) & (g712) & (!g715) & (g722) & (g721) & (!g716)) + ((!g711) & (g712) & (!g715) & (g722) & (g721) & (g716)) + ((!g711) & (g712) & (g715) & (!g722) & (!g721) & (!g716)) + ((!g711) & (g712) & (g715) & (!g722) & (g721) & (!g716)) + ((!g711) & (g712) & (g715) & (!g722) & (g721) & (g716)) + ((!g711) & (g712) & (g715) & (g722) & (!g721) & (!g716)) + ((!g711) & (g712) & (g715) & (g722) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g722) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g722) & (g721) & (g716)) + ((g711) & (!g712) & (!g715) & (g722) & (!g721) & (g716)) + ((g711) & (!g712) & (!g715) & (g722) & (g721) & (g716)) + ((g711) & (!g712) & (g715) & (!g722) & (!g721) & (!g716)) + ((g711) & (!g712) & (g715) & (!g722) & (!g721) & (g716)) + ((g711) & (!g712) & (g715) & (!g722) & (g721) & (g716)) + ((g711) & (!g712) & (g715) & (g722) & (!g721) & (!g716)) + ((g711) & (!g712) & (g715) & (g722) & (!g721) & (g716)) + ((g711) & (!g712) & (g715) & (g722) & (g721) & (!g716)) + ((g711) & (!g712) & (g715) & (g722) & (g721) & (g716)) + ((g711) & (g712) & (!g715) & (!g722) & (!g721) & (g716)) + ((g711) & (g712) & (!g715) & (g722) & (!g721) & (!g716)) + ((g711) & (g712) & (!g715) & (g722) & (g721) & (!g716)) + ((g711) & (g712) & (g715) & (!g722) & (!g721) & (!g716)) + ((g711) & (g712) & (g715) & (!g722) & (!g721) & (g716)) + ((g711) & (g712) & (g715) & (!g722) & (g721) & (!g716)) + ((g711) & (g712) & (g715) & (g722) & (!g721) & (!g716)) + ((g711) & (g712) & (g715) & (g722) & (g721) & (!g716)));
	assign g750 = (((!g711) & (!g712) & (!g715) & (!g722) & (g721) & (g716)) + ((!g711) & (!g712) & (!g715) & (g722) & (!g721) & (!g716)) + ((!g711) & (!g712) & (!g715) & (g722) & (g721) & (g716)) + ((!g711) & (!g712) & (g715) & (!g722) & (!g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (!g722) & (g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (g722) & (!g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (g722) & (!g721) & (g716)) + ((!g711) & (!g712) & (g715) & (g722) & (g721) & (!g716)) + ((!g711) & (g712) & (!g715) & (!g722) & (!g721) & (!g716)) + ((!g711) & (g712) & (!g715) & (g722) & (!g721) & (g716)) + ((!g711) & (g712) & (!g715) & (g722) & (g721) & (!g716)) + ((!g711) & (g712) & (!g715) & (g722) & (g721) & (g716)) + ((!g711) & (g712) & (g715) & (!g722) & (!g721) & (!g716)) + ((!g711) & (g712) & (g715) & (g722) & (!g721) & (!g716)) + ((!g711) & (g712) & (g715) & (g722) & (!g721) & (g716)) + ((g711) & (!g712) & (!g715) & (!g722) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g722) & (g721) & (g716)) + ((g711) & (!g712) & (g715) & (!g722) & (!g721) & (!g716)) + ((g711) & (!g712) & (g715) & (!g722) & (g721) & (!g716)) + ((g711) & (!g712) & (g715) & (g722) & (g721) & (!g716)) + ((g711) & (g712) & (!g715) & (!g722) & (g721) & (!g716)) + ((g711) & (g712) & (!g715) & (g722) & (g721) & (g716)) + ((g711) & (g712) & (g715) & (!g722) & (!g721) & (!g716)) + ((g711) & (g712) & (g715) & (!g722) & (!g721) & (g716)) + ((g711) & (g712) & (g715) & (!g722) & (g721) & (!g716)) + ((g711) & (g712) & (g715) & (g722) & (!g721) & (!g716)));
	assign g751 = (((!g747) & (!g748) & (!g749) & (!g750) & (g713) & (g714)) + ((!g747) & (!g748) & (g749) & (!g750) & (!g713) & (g714)) + ((!g747) & (!g748) & (g749) & (!g750) & (g713) & (g714)) + ((!g747) & (!g748) & (g749) & (g750) & (!g713) & (g714)) + ((!g747) & (g748) & (!g749) & (!g750) & (g713) & (!g714)) + ((!g747) & (g748) & (!g749) & (!g750) & (g713) & (g714)) + ((!g747) & (g748) & (!g749) & (g750) & (g713) & (!g714)) + ((!g747) & (g748) & (g749) & (!g750) & (!g713) & (g714)) + ((!g747) & (g748) & (g749) & (!g750) & (g713) & (!g714)) + ((!g747) & (g748) & (g749) & (!g750) & (g713) & (g714)) + ((!g747) & (g748) & (g749) & (g750) & (!g713) & (g714)) + ((!g747) & (g748) & (g749) & (g750) & (g713) & (!g714)) + ((g747) & (!g748) & (!g749) & (!g750) & (!g713) & (!g714)) + ((g747) & (!g748) & (!g749) & (!g750) & (g713) & (g714)) + ((g747) & (!g748) & (!g749) & (g750) & (!g713) & (!g714)) + ((g747) & (!g748) & (g749) & (!g750) & (!g713) & (!g714)) + ((g747) & (!g748) & (g749) & (!g750) & (!g713) & (g714)) + ((g747) & (!g748) & (g749) & (!g750) & (g713) & (g714)) + ((g747) & (!g748) & (g749) & (g750) & (!g713) & (!g714)) + ((g747) & (!g748) & (g749) & (g750) & (!g713) & (g714)) + ((g747) & (g748) & (!g749) & (!g750) & (!g713) & (!g714)) + ((g747) & (g748) & (!g749) & (!g750) & (g713) & (!g714)) + ((g747) & (g748) & (!g749) & (!g750) & (g713) & (g714)) + ((g747) & (g748) & (!g749) & (g750) & (!g713) & (!g714)) + ((g747) & (g748) & (!g749) & (g750) & (g713) & (!g714)) + ((g747) & (g748) & (g749) & (!g750) & (!g713) & (!g714)) + ((g747) & (g748) & (g749) & (!g750) & (!g713) & (g714)) + ((g747) & (g748) & (g749) & (!g750) & (g713) & (!g714)) + ((g747) & (g748) & (g749) & (!g750) & (g713) & (g714)) + ((g747) & (g748) & (g749) & (g750) & (!g713) & (!g714)) + ((g747) & (g748) & (g749) & (g750) & (!g713) & (g714)) + ((g747) & (g748) & (g749) & (g750) & (g713) & (!g714)));
	assign g753 = (((!sk[78]) & (g751) & (!g752)) + ((!sk[78]) & (g751) & (g752)) + ((sk[78]) & (!g751) & (g752)) + ((sk[78]) & (g751) & (!g752)));
	assign g754 = (((!g711) & (!g712) & (!g715) & (!g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (!g715) & (!g714) & (g721) & (g716)) + ((!g711) & (!g712) & (!g715) & (g714) & (g721) & (g716)) + ((!g711) & (!g712) & (g715) & (!g714) & (!g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (!g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (g715) & (!g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (!g714) & (g721) & (g716)) + ((!g711) & (!g712) & (g715) & (g714) & (!g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (g714) & (!g721) & (g716)) + ((!g711) & (g712) & (!g715) & (!g714) & (!g721) & (g716)) + ((!g711) & (g712) & (!g715) & (!g714) & (g721) & (!g716)) + ((!g711) & (g712) & (!g715) & (g714) & (g721) & (g716)) + ((!g711) & (g712) & (g715) & (!g714) & (g721) & (!g716)) + ((!g711) & (g712) & (g715) & (!g714) & (g721) & (g716)) + ((!g711) & (g712) & (g715) & (g714) & (!g721) & (!g716)) + ((!g711) & (g712) & (g715) & (g714) & (!g721) & (g716)) + ((!g711) & (g712) & (g715) & (g714) & (g721) & (g716)) + ((g711) & (!g712) & (!g715) & (!g714) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g714) & (g721) & (g716)) + ((g711) & (!g712) & (!g715) & (g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (g714) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (g714) & (g721) & (g716)) + ((g711) & (!g712) & (g715) & (!g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (g715) & (!g714) & (g721) & (!g716)) + ((g711) & (!g712) & (g715) & (g714) & (g721) & (!g716)) + ((g711) & (g712) & (!g715) & (!g714) & (g721) & (g716)) + ((g711) & (g712) & (g715) & (!g714) & (!g721) & (!g716)) + ((g711) & (g712) & (g715) & (!g714) & (g721) & (g716)));
	assign g755 = (((!g711) & (!g712) & (!g715) & (!g714) & (!g721) & (!g716)) + ((!g711) & (!g712) & (!g715) & (g714) & (!g721) & (!g716)) + ((!g711) & (!g712) & (!g715) & (g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (!g715) & (g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (!g714) & (g721) & (g716)) + ((!g711) & (!g712) & (g715) & (g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (g715) & (g714) & (g721) & (g716)) + ((!g711) & (g712) & (!g715) & (!g714) & (!g721) & (!g716)) + ((!g711) & (g712) & (!g715) & (!g714) & (g721) & (!g716)) + ((!g711) & (g712) & (g715) & (!g714) & (!g721) & (g716)) + ((!g711) & (g712) & (g715) & (!g714) & (g721) & (g716)) + ((!g711) & (g712) & (g715) & (g714) & (!g721) & (g716)) + ((!g711) & (g712) & (g715) & (g714) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g714) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g714) & (g721) & (g716)) + ((g711) & (!g712) & (!g715) & (g714) & (!g721) & (g716)) + ((g711) & (!g712) & (!g715) & (g714) & (g721) & (g716)) + ((g711) & (!g712) & (g715) & (g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (g715) & (g714) & (!g721) & (g716)) + ((g711) & (!g712) & (g715) & (g714) & (g721) & (g716)) + ((g711) & (g712) & (!g715) & (!g714) & (!g721) & (g716)) + ((g711) & (g712) & (!g715) & (!g714) & (g721) & (!g716)) + ((g711) & (g712) & (!g715) & (g714) & (g721) & (!g716)) + ((g711) & (g712) & (g715) & (!g714) & (!g721) & (g716)) + ((g711) & (g712) & (g715) & (!g714) & (g721) & (g716)) + ((g711) & (g712) & (g715) & (g714) & (!g721) & (!g716)) + ((g711) & (g712) & (g715) & (g714) & (g721) & (g716)));
	assign g756 = (((!g711) & (!g712) & (!g715) & (!g714) & (g721) & (g716)) + ((!g711) & (!g712) & (!g715) & (g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (!g714) & (!g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (!g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (g715) & (!g714) & (g721) & (g716)) + ((!g711) & (!g712) & (g715) & (g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (g715) & (g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (g715) & (g714) & (g721) & (g716)) + ((!g711) & (g712) & (!g715) & (!g714) & (g721) & (!g716)) + ((!g711) & (g712) & (!g715) & (!g714) & (g721) & (g716)) + ((!g711) & (g712) & (g715) & (!g714) & (!g721) & (!g716)) + ((!g711) & (g712) & (g715) & (g714) & (!g721) & (g716)) + ((!g711) & (g712) & (g715) & (g714) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g714) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (!g714) & (g721) & (g716)) + ((g711) & (!g712) & (!g715) & (g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (g714) & (!g721) & (g716)) + ((g711) & (!g712) & (g715) & (!g714) & (!g721) & (g716)) + ((g711) & (!g712) & (g715) & (!g714) & (g721) & (g716)) + ((g711) & (!g712) & (g715) & (g714) & (g721) & (!g716)) + ((g711) & (g712) & (!g715) & (!g714) & (!g721) & (!g716)) + ((g711) & (g712) & (!g715) & (!g714) & (!g721) & (g716)) + ((g711) & (g712) & (!g715) & (!g714) & (g721) & (g716)) + ((g711) & (g712) & (!g715) & (g714) & (!g721) & (g716)) + ((g711) & (g712) & (!g715) & (g714) & (g721) & (!g716)) + ((g711) & (g712) & (g715) & (!g714) & (!g721) & (g716)) + ((g711) & (g712) & (g715) & (!g714) & (g721) & (!g716)) + ((g711) & (g712) & (g715) & (g714) & (!g721) & (!g716)) + ((g711) & (g712) & (g715) & (g714) & (g721) & (!g716)) + ((g711) & (g712) & (g715) & (g714) & (g721) & (g716)));
	assign g757 = (((!g711) & (!g712) & (!g715) & (!g714) & (g721) & (!g716)) + ((!g711) & (!g712) & (!g715) & (g714) & (!g721) & (!g716)) + ((!g711) & (!g712) & (!g715) & (g714) & (g721) & (g716)) + ((!g711) & (!g712) & (g715) & (!g714) & (!g721) & (g716)) + ((!g711) & (!g712) & (g715) & (!g714) & (g721) & (g716)) + ((!g711) & (!g712) & (g715) & (g714) & (g721) & (g716)) + ((!g711) & (g712) & (!g715) & (!g714) & (!g721) & (g716)) + ((!g711) & (g712) & (!g715) & (g714) & (!g721) & (g716)) + ((!g711) & (g712) & (!g715) & (g714) & (g721) & (g716)) + ((!g711) & (g712) & (g715) & (!g714) & (!g721) & (!g716)) + ((!g711) & (g712) & (g715) & (!g714) & (g721) & (!g716)) + ((!g711) & (g712) & (g715) & (g714) & (!g721) & (g716)) + ((!g711) & (g712) & (g715) & (g714) & (g721) & (g716)) + ((g711) & (!g712) & (!g715) & (!g714) & (g721) & (!g716)) + ((g711) & (!g712) & (!g715) & (g714) & (g721) & (g716)) + ((g711) & (!g712) & (g715) & (!g714) & (!g721) & (!g716)) + ((g711) & (!g712) & (g715) & (!g714) & (g721) & (g716)) + ((g711) & (!g712) & (g715) & (g714) & (!g721) & (!g716)) + ((g711) & (g712) & (!g715) & (!g714) & (g721) & (g716)) + ((g711) & (g712) & (!g715) & (g714) & (!g721) & (!g716)) + ((g711) & (g712) & (!g715) & (g714) & (!g721) & (g716)) + ((g711) & (g712) & (g715) & (!g714) & (g721) & (g716)));
	assign g758 = (((!g754) & (!g755) & (!g756) & (!g757) & (!g722) & (!g713)) + ((!g754) & (!g755) & (!g756) & (!g757) & (!g722) & (g713)) + ((!g754) & (!g755) & (!g756) & (!g757) & (g722) & (!g713)) + ((!g754) & (!g755) & (!g756) & (g757) & (!g722) & (!g713)) + ((!g754) & (!g755) & (!g756) & (g757) & (!g722) & (g713)) + ((!g754) & (!g755) & (!g756) & (g757) & (g722) & (!g713)) + ((!g754) & (!g755) & (!g756) & (g757) & (g722) & (g713)) + ((!g754) & (!g755) & (g756) & (!g757) & (!g722) & (!g713)) + ((!g754) & (!g755) & (g756) & (!g757) & (g722) & (!g713)) + ((!g754) & (!g755) & (g756) & (g757) & (!g722) & (!g713)) + ((!g754) & (!g755) & (g756) & (g757) & (g722) & (!g713)) + ((!g754) & (!g755) & (g756) & (g757) & (g722) & (g713)) + ((!g754) & (g755) & (!g756) & (!g757) & (!g722) & (!g713)) + ((!g754) & (g755) & (!g756) & (!g757) & (!g722) & (g713)) + ((!g754) & (g755) & (!g756) & (g757) & (!g722) & (!g713)) + ((!g754) & (g755) & (!g756) & (g757) & (!g722) & (g713)) + ((!g754) & (g755) & (!g756) & (g757) & (g722) & (g713)) + ((!g754) & (g755) & (g756) & (!g757) & (!g722) & (!g713)) + ((!g754) & (g755) & (g756) & (g757) & (!g722) & (!g713)) + ((!g754) & (g755) & (g756) & (g757) & (g722) & (g713)) + ((g754) & (!g755) & (!g756) & (!g757) & (!g722) & (g713)) + ((g754) & (!g755) & (!g756) & (!g757) & (g722) & (!g713)) + ((g754) & (!g755) & (!g756) & (g757) & (!g722) & (g713)) + ((g754) & (!g755) & (!g756) & (g757) & (g722) & (!g713)) + ((g754) & (!g755) & (!g756) & (g757) & (g722) & (g713)) + ((g754) & (!g755) & (g756) & (!g757) & (g722) & (!g713)) + ((g754) & (!g755) & (g756) & (g757) & (g722) & (!g713)) + ((g754) & (!g755) & (g756) & (g757) & (g722) & (g713)) + ((g754) & (g755) & (!g756) & (!g757) & (!g722) & (g713)) + ((g754) & (g755) & (!g756) & (g757) & (!g722) & (g713)) + ((g754) & (g755) & (!g756) & (g757) & (g722) & (g713)) + ((g754) & (g755) & (g756) & (g757) & (g722) & (g713)));
	assign g760 = (((!g758) & (sk[84]) & (g759)) + ((g758) & (!sk[84]) & (!g759)) + ((g758) & (!sk[84]) & (g759)) + ((g758) & (sk[84]) & (!g759)));
	assign g761 = (((!g711) & (!g722) & (!g713) & (!g714) & (!g721) & (g716)) + ((!g711) & (!g722) & (!g713) & (!g714) & (g721) & (g716)) + ((!g711) & (!g722) & (!g713) & (g714) & (!g721) & (!g716)) + ((!g711) & (!g722) & (!g713) & (g714) & (!g721) & (g716)) + ((!g711) & (!g722) & (!g713) & (g714) & (g721) & (!g716)) + ((!g711) & (!g722) & (!g713) & (g714) & (g721) & (g716)) + ((!g711) & (!g722) & (g713) & (!g714) & (!g721) & (g716)) + ((!g711) & (!g722) & (g713) & (!g714) & (g721) & (g716)) + ((!g711) & (!g722) & (g713) & (g714) & (g721) & (!g716)) + ((!g711) & (g722) & (g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (g722) & (g713) & (!g714) & (g721) & (g716)) + ((!g711) & (g722) & (g713) & (g714) & (!g721) & (g716)) + ((g711) & (!g722) & (!g713) & (!g714) & (g721) & (!g716)) + ((g711) & (!g722) & (!g713) & (g714) & (!g721) & (!g716)) + ((g711) & (!g722) & (!g713) & (g714) & (!g721) & (g716)) + ((g711) & (!g722) & (!g713) & (g714) & (g721) & (g716)) + ((g711) & (!g722) & (g713) & (!g714) & (!g721) & (g716)) + ((g711) & (!g722) & (g713) & (!g714) & (g721) & (g716)) + ((g711) & (!g722) & (g713) & (g714) & (g721) & (!g716)) + ((g711) & (!g722) & (g713) & (g714) & (g721) & (g716)) + ((g711) & (g722) & (!g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (g722) & (!g713) & (!g714) & (!g721) & (g716)) + ((g711) & (g722) & (!g713) & (!g714) & (g721) & (!g716)) + ((g711) & (g722) & (!g713) & (g714) & (!g721) & (!g716)) + ((g711) & (g722) & (g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (g722) & (g713) & (!g714) & (!g721) & (g716)) + ((g711) & (g722) & (g713) & (!g714) & (g721) & (!g716)) + ((g711) & (g722) & (g713) & (g714) & (!g721) & (g716)));
	assign g762 = (((!g711) & (!g722) & (!g713) & (!g714) & (!g721) & (!g716)) + ((!g711) & (!g722) & (!g713) & (g714) & (g721) & (g716)) + ((!g711) & (!g722) & (g713) & (!g714) & (!g721) & (!g716)) + ((!g711) & (!g722) & (g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (!g722) & (g713) & (!g714) & (g721) & (g716)) + ((!g711) & (!g722) & (g713) & (g714) & (!g721) & (!g716)) + ((!g711) & (!g722) & (g713) & (g714) & (g721) & (g716)) + ((!g711) & (g722) & (!g713) & (!g714) & (!g721) & (!g716)) + ((!g711) & (g722) & (!g713) & (!g714) & (g721) & (g716)) + ((!g711) & (g722) & (!g713) & (g714) & (!g721) & (g716)) + ((!g711) & (g722) & (g713) & (!g714) & (!g721) & (!g716)) + ((!g711) & (g722) & (g713) & (!g714) & (g721) & (g716)) + ((!g711) & (g722) & (g713) & (g714) & (g721) & (!g716)) + ((!g711) & (g722) & (g713) & (g714) & (g721) & (g716)) + ((g711) & (!g722) & (!g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (!g722) & (!g713) & (!g714) & (g721) & (g716)) + ((g711) & (!g722) & (!g713) & (g714) & (!g721) & (!g716)) + ((g711) & (!g722) & (!g713) & (g714) & (g721) & (g716)) + ((g711) & (!g722) & (g713) & (!g714) & (g721) & (g716)) + ((g711) & (!g722) & (g713) & (g714) & (!g721) & (g716)) + ((g711) & (g722) & (!g713) & (!g714) & (g721) & (!g716)) + ((g711) & (g722) & (!g713) & (!g714) & (g721) & (g716)) + ((g711) & (g722) & (!g713) & (g714) & (!g721) & (g716)) + ((g711) & (g722) & (!g713) & (g714) & (g721) & (!g716)) + ((g711) & (g722) & (!g713) & (g714) & (g721) & (g716)) + ((g711) & (g722) & (g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (g722) & (g713) & (!g714) & (g721) & (!g716)) + ((g711) & (g722) & (g713) & (g714) & (!g721) & (!g716)));
	assign g763 = (((!g711) & (!g722) & (!g713) & (!g714) & (!g721) & (g716)) + ((!g711) & (!g722) & (!g713) & (!g714) & (g721) & (g716)) + ((!g711) & (!g722) & (!g713) & (g714) & (g721) & (!g716)) + ((!g711) & (!g722) & (!g713) & (g714) & (g721) & (g716)) + ((!g711) & (!g722) & (g713) & (!g714) & (g721) & (g716)) + ((!g711) & (!g722) & (g713) & (g714) & (!g721) & (!g716)) + ((!g711) & (!g722) & (g713) & (g714) & (!g721) & (g716)) + ((!g711) & (!g722) & (g713) & (g714) & (g721) & (g716)) + ((!g711) & (g722) & (!g713) & (!g714) & (!g721) & (!g716)) + ((!g711) & (g722) & (!g713) & (!g714) & (!g721) & (g716)) + ((!g711) & (g722) & (!g713) & (!g714) & (g721) & (g716)) + ((!g711) & (g722) & (!g713) & (g714) & (!g721) & (g716)) + ((!g711) & (g722) & (!g713) & (g714) & (g721) & (!g716)) + ((!g711) & (g722) & (g713) & (!g714) & (!g721) & (g716)) + ((!g711) & (g722) & (g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (g722) & (g713) & (g714) & (!g721) & (!g716)) + ((!g711) & (g722) & (g713) & (g714) & (g721) & (!g716)) + ((!g711) & (g722) & (g713) & (g714) & (g721) & (g716)) + ((g711) & (!g722) & (!g713) & (!g714) & (!g721) & (g716)) + ((g711) & (!g722) & (!g713) & (g714) & (!g721) & (!g716)) + ((g711) & (!g722) & (!g713) & (g714) & (g721) & (!g716)) + ((g711) & (!g722) & (g713) & (!g714) & (g721) & (g716)) + ((g711) & (!g722) & (g713) & (g714) & (!g721) & (g716)) + ((g711) & (g722) & (!g713) & (!g714) & (!g721) & (g716)) + ((g711) & (g722) & (!g713) & (g714) & (!g721) & (!g716)) + ((g711) & (g722) & (!g713) & (g714) & (g721) & (!g716)) + ((g711) & (g722) & (g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (g722) & (g713) & (!g714) & (g721) & (!g716)) + ((g711) & (g722) & (g713) & (!g714) & (g721) & (g716)) + ((g711) & (g722) & (g713) & (g714) & (g721) & (g716)));
	assign g764 = (((!g711) & (!g722) & (!g713) & (!g714) & (g721) & (g716)) + ((!g711) & (!g722) & (!g713) & (g714) & (!g721) & (!g716)) + ((!g711) & (!g722) & (!g713) & (g714) & (g721) & (g716)) + ((!g711) & (!g722) & (g713) & (!g714) & (!g721) & (!g716)) + ((!g711) & (!g722) & (g713) & (g714) & (g721) & (!g716)) + ((!g711) & (!g722) & (g713) & (g714) & (g721) & (g716)) + ((!g711) & (g722) & (!g713) & (g714) & (!g721) & (!g716)) + ((!g711) & (g722) & (!g713) & (g714) & (g721) & (!g716)) + ((!g711) & (g722) & (g713) & (!g714) & (g721) & (!g716)) + ((!g711) & (g722) & (g713) & (!g714) & (g721) & (g716)) + ((g711) & (!g722) & (!g713) & (!g714) & (!g721) & (g716)) + ((g711) & (!g722) & (!g713) & (!g714) & (g721) & (!g716)) + ((g711) & (!g722) & (!g713) & (g714) & (!g721) & (g716)) + ((g711) & (!g722) & (g713) & (!g714) & (g721) & (!g716)) + ((g711) & (!g722) & (g713) & (!g714) & (g721) & (g716)) + ((g711) & (!g722) & (g713) & (g714) & (g721) & (!g716)) + ((g711) & (!g722) & (g713) & (g714) & (g721) & (g716)) + ((g711) & (g722) & (!g713) & (!g714) & (g721) & (!g716)) + ((g711) & (g722) & (!g713) & (g714) & (!g721) & (g716)) + ((g711) & (g722) & (g713) & (!g714) & (!g721) & (!g716)) + ((g711) & (g722) & (g713) & (!g714) & (g721) & (g716)) + ((g711) & (g722) & (g713) & (g714) & (!g721) & (g716)));
	assign g765 = (((!g761) & (!g762) & (!g763) & (!g764) & (!g715) & (!g712)) + ((!g761) & (!g762) & (!g763) & (!g764) & (!g715) & (g712)) + ((!g761) & (!g762) & (!g763) & (!g764) & (g715) & (!g712)) + ((!g761) & (!g762) & (!g763) & (g764) & (!g715) & (!g712)) + ((!g761) & (!g762) & (!g763) & (g764) & (!g715) & (g712)) + ((!g761) & (!g762) & (!g763) & (g764) & (g715) & (!g712)) + ((!g761) & (!g762) & (!g763) & (g764) & (g715) & (g712)) + ((!g761) & (!g762) & (g763) & (!g764) & (!g715) & (!g712)) + ((!g761) & (!g762) & (g763) & (!g764) & (g715) & (!g712)) + ((!g761) & (!g762) & (g763) & (g764) & (!g715) & (!g712)) + ((!g761) & (!g762) & (g763) & (g764) & (g715) & (!g712)) + ((!g761) & (!g762) & (g763) & (g764) & (g715) & (g712)) + ((!g761) & (g762) & (!g763) & (!g764) & (!g715) & (!g712)) + ((!g761) & (g762) & (!g763) & (!g764) & (!g715) & (g712)) + ((!g761) & (g762) & (!g763) & (g764) & (!g715) & (!g712)) + ((!g761) & (g762) & (!g763) & (g764) & (!g715) & (g712)) + ((!g761) & (g762) & (!g763) & (g764) & (g715) & (g712)) + ((!g761) & (g762) & (g763) & (!g764) & (!g715) & (!g712)) + ((!g761) & (g762) & (g763) & (g764) & (!g715) & (!g712)) + ((!g761) & (g762) & (g763) & (g764) & (g715) & (g712)) + ((g761) & (!g762) & (!g763) & (!g764) & (!g715) & (g712)) + ((g761) & (!g762) & (!g763) & (!g764) & (g715) & (!g712)) + ((g761) & (!g762) & (!g763) & (g764) & (!g715) & (g712)) + ((g761) & (!g762) & (!g763) & (g764) & (g715) & (!g712)) + ((g761) & (!g762) & (!g763) & (g764) & (g715) & (g712)) + ((g761) & (!g762) & (g763) & (!g764) & (g715) & (!g712)) + ((g761) & (!g762) & (g763) & (g764) & (g715) & (!g712)) + ((g761) & (!g762) & (g763) & (g764) & (g715) & (g712)) + ((g761) & (g762) & (!g763) & (!g764) & (!g715) & (g712)) + ((g761) & (g762) & (!g763) & (g764) & (!g715) & (g712)) + ((g761) & (g762) & (!g763) & (g764) & (g715) & (g712)) + ((g761) & (g762) & (g763) & (g764) & (g715) & (g712)));
	assign g767 = (((!g765) & (sk[90]) & (g766)) + ((g765) & (!sk[90]) & (!g766)) + ((g765) & (!sk[90]) & (g766)) + ((g765) & (sk[90]) & (!g766)));
	assign g768 = (((!g715) & (!g712) & (!g713) & (!g714) & (!g721) & (g722)) + ((!g715) & (!g712) & (!g713) & (!g714) & (g721) & (!g722)) + ((!g715) & (!g712) & (!g713) & (g714) & (!g721) & (g722)) + ((!g715) & (!g712) & (!g713) & (g714) & (g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (!g714) & (!g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (!g714) & (g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (g714) & (!g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (g714) & (g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (g714) & (g721) & (g722)) + ((!g715) & (g712) & (!g713) & (!g714) & (g721) & (!g722)) + ((!g715) & (g712) & (!g713) & (g714) & (g721) & (!g722)) + ((!g715) & (g712) & (!g713) & (g714) & (g721) & (g722)) + ((!g715) & (g712) & (g713) & (!g714) & (g721) & (g722)) + ((!g715) & (g712) & (g713) & (g714) & (!g721) & (!g722)) + ((g715) & (!g712) & (!g713) & (!g714) & (!g721) & (g722)) + ((g715) & (!g712) & (!g713) & (g714) & (!g721) & (g722)) + ((g715) & (!g712) & (g713) & (g714) & (g721) & (g722)) + ((g715) & (g712) & (!g713) & (!g714) & (g721) & (g722)) + ((g715) & (g712) & (!g713) & (g714) & (!g721) & (!g722)) + ((g715) & (g712) & (!g713) & (g714) & (g721) & (!g722)) + ((g715) & (g712) & (g713) & (!g714) & (!g721) & (g722)) + ((g715) & (g712) & (g713) & (!g714) & (g721) & (!g722)) + ((g715) & (g712) & (g713) & (!g714) & (g721) & (g722)) + ((g715) & (g712) & (g713) & (g714) & (!g721) & (g722)));
	assign g769 = (((!g715) & (!g712) & (!g713) & (!g714) & (!g721) & (!g722)) + ((!g715) & (!g712) & (!g713) & (!g714) & (!g721) & (g722)) + ((!g715) & (!g712) & (!g713) & (g714) & (!g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (!g714) & (!g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (!g714) & (g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (!g714) & (g721) & (g722)) + ((!g715) & (!g712) & (g713) & (g714) & (!g721) & (g722)) + ((!g715) & (!g712) & (g713) & (g714) & (g721) & (g722)) + ((!g715) & (g712) & (!g713) & (!g714) & (!g721) & (!g722)) + ((!g715) & (g712) & (!g713) & (!g714) & (g721) & (!g722)) + ((!g715) & (g712) & (!g713) & (g714) & (!g721) & (!g722)) + ((!g715) & (g712) & (!g713) & (g714) & (!g721) & (g722)) + ((!g715) & (g712) & (!g713) & (g714) & (g721) & (g722)) + ((!g715) & (g712) & (g713) & (!g714) & (!g721) & (g722)) + ((!g715) & (g712) & (g713) & (g714) & (!g721) & (!g722)) + ((!g715) & (g712) & (g713) & (g714) & (!g721) & (g722)) + ((g715) & (!g712) & (!g713) & (!g714) & (!g721) & (g722)) + ((g715) & (!g712) & (!g713) & (!g714) & (g721) & (g722)) + ((g715) & (!g712) & (!g713) & (g714) & (!g721) & (!g722)) + ((g715) & (!g712) & (!g713) & (g714) & (g721) & (g722)) + ((g715) & (!g712) & (g713) & (!g714) & (!g721) & (!g722)) + ((g715) & (!g712) & (g713) & (!g714) & (g721) & (g722)) + ((g715) & (!g712) & (g713) & (g714) & (g721) & (!g722)) + ((g715) & (g712) & (!g713) & (!g714) & (!g721) & (!g722)) + ((g715) & (g712) & (!g713) & (!g714) & (!g721) & (g722)) + ((g715) & (g712) & (!g713) & (!g714) & (g721) & (g722)) + ((g715) & (g712) & (!g713) & (g714) & (!g721) & (g722)) + ((g715) & (g712) & (!g713) & (g714) & (g721) & (!g722)) + ((g715) & (g712) & (g713) & (!g714) & (g721) & (!g722)) + ((g715) & (g712) & (g713) & (!g714) & (g721) & (g722)));
	assign g770 = (((!g715) & (!g712) & (!g713) & (!g714) & (g721) & (!g722)) + ((!g715) & (!g712) & (!g713) & (g714) & (!g721) & (!g722)) + ((!g715) & (!g712) & (!g713) & (g714) & (g721) & (!g722)) + ((!g715) & (!g712) & (!g713) & (g714) & (g721) & (g722)) + ((!g715) & (!g712) & (g713) & (!g714) & (!g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (!g714) & (!g721) & (g722)) + ((!g715) & (!g712) & (g713) & (!g714) & (g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (g714) & (!g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (g714) & (g721) & (g722)) + ((!g715) & (g712) & (!g713) & (!g714) & (!g721) & (g722)) + ((!g715) & (g712) & (!g713) & (!g714) & (g721) & (!g722)) + ((!g715) & (g712) & (!g713) & (!g714) & (g721) & (g722)) + ((!g715) & (g712) & (g713) & (!g714) & (!g721) & (g722)) + ((!g715) & (g712) & (g713) & (!g714) & (g721) & (!g722)) + ((!g715) & (g712) & (g713) & (!g714) & (g721) & (g722)) + ((!g715) & (g712) & (g713) & (g714) & (!g721) & (!g722)) + ((g715) & (!g712) & (!g713) & (!g714) & (g721) & (!g722)) + ((g715) & (!g712) & (!g713) & (g714) & (!g721) & (!g722)) + ((g715) & (!g712) & (!g713) & (g714) & (g721) & (g722)) + ((g715) & (!g712) & (g713) & (!g714) & (!g721) & (!g722)) + ((g715) & (!g712) & (g713) & (!g714) & (!g721) & (g722)) + ((g715) & (!g712) & (g713) & (g714) & (!g721) & (!g722)) + ((g715) & (!g712) & (g713) & (g714) & (g721) & (!g722)) + ((g715) & (g712) & (!g713) & (!g714) & (g721) & (!g722)) + ((g715) & (g712) & (!g713) & (g714) & (!g721) & (!g722)) + ((g715) & (g712) & (!g713) & (g714) & (g721) & (g722)) + ((g715) & (g712) & (g713) & (!g714) & (!g721) & (!g722)) + ((g715) & (g712) & (g713) & (!g714) & (g721) & (!g722)) + ((g715) & (g712) & (g713) & (!g714) & (g721) & (g722)) + ((g715) & (g712) & (g713) & (g714) & (!g721) & (g722)));
	assign g771 = (((!g715) & (!g712) & (!g713) & (!g714) & (!g721) & (g722)) + ((!g715) & (!g712) & (!g713) & (g714) & (g721) & (!g722)) + ((!g715) & (!g712) & (!g713) & (g714) & (g721) & (g722)) + ((!g715) & (!g712) & (g713) & (!g714) & (!g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (!g714) & (!g721) & (g722)) + ((!g715) & (!g712) & (g713) & (g714) & (g721) & (!g722)) + ((!g715) & (!g712) & (g713) & (g714) & (g721) & (g722)) + ((!g715) & (g712) & (!g713) & (!g714) & (!g721) & (!g722)) + ((!g715) & (g712) & (!g713) & (!g714) & (!g721) & (g722)) + ((!g715) & (g712) & (!g713) & (!g714) & (g721) & (g722)) + ((!g715) & (g712) & (!g713) & (g714) & (!g721) & (g722)) + ((!g715) & (g712) & (g713) & (!g714) & (!g721) & (g722)) + ((!g715) & (g712) & (g713) & (g714) & (!g721) & (!g722)) + ((!g715) & (g712) & (g713) & (g714) & (!g721) & (g722)) + ((!g715) & (g712) & (g713) & (g714) & (g721) & (!g722)) + ((!g715) & (g712) & (g713) & (g714) & (g721) & (g722)) + ((g715) & (!g712) & (!g713) & (g714) & (!g721) & (g722)) + ((g715) & (!g712) & (g713) & (!g714) & (!g721) & (!g722)) + ((g715) & (!g712) & (g713) & (g714) & (!g721) & (!g722)) + ((g715) & (!g712) & (g713) & (g714) & (!g721) & (g722)) + ((g715) & (!g712) & (g713) & (g714) & (g721) & (g722)) + ((g715) & (g712) & (!g713) & (!g714) & (!g721) & (g722)) + ((g715) & (g712) & (!g713) & (!g714) & (g721) & (g722)) + ((g715) & (g712) & (!g713) & (g714) & (!g721) & (!g722)) + ((g715) & (g712) & (!g713) & (g714) & (g721) & (!g722)) + ((g715) & (g712) & (!g713) & (g714) & (g721) & (g722)) + ((g715) & (g712) & (g713) & (!g714) & (g721) & (g722)) + ((g715) & (g712) & (g713) & (g714) & (g721) & (g722)));
	assign g772 = (((!g768) & (!g769) & (!g770) & (!g771) & (!g711) & (g716)) + ((!g768) & (!g769) & (!g770) & (!g771) & (g711) & (!g716)) + ((!g768) & (!g769) & (!g770) & (!g771) & (g711) & (g716)) + ((!g768) & (!g769) & (!g770) & (g771) & (!g711) & (g716)) + ((!g768) & (!g769) & (!g770) & (g771) & (g711) & (!g716)) + ((!g768) & (!g769) & (g770) & (!g771) & (g711) & (!g716)) + ((!g768) & (!g769) & (g770) & (!g771) & (g711) & (g716)) + ((!g768) & (!g769) & (g770) & (g771) & (g711) & (!g716)) + ((!g768) & (g769) & (!g770) & (!g771) & (!g711) & (g716)) + ((!g768) & (g769) & (!g770) & (!g771) & (g711) & (g716)) + ((!g768) & (g769) & (!g770) & (g771) & (!g711) & (g716)) + ((!g768) & (g769) & (g770) & (!g771) & (g711) & (g716)) + ((g768) & (!g769) & (!g770) & (!g771) & (!g711) & (!g716)) + ((g768) & (!g769) & (!g770) & (!g771) & (!g711) & (g716)) + ((g768) & (!g769) & (!g770) & (!g771) & (g711) & (!g716)) + ((g768) & (!g769) & (!g770) & (!g771) & (g711) & (g716)) + ((g768) & (!g769) & (!g770) & (g771) & (!g711) & (!g716)) + ((g768) & (!g769) & (!g770) & (g771) & (!g711) & (g716)) + ((g768) & (!g769) & (!g770) & (g771) & (g711) & (!g716)) + ((g768) & (!g769) & (g770) & (!g771) & (!g711) & (!g716)) + ((g768) & (!g769) & (g770) & (!g771) & (g711) & (!g716)) + ((g768) & (!g769) & (g770) & (!g771) & (g711) & (g716)) + ((g768) & (!g769) & (g770) & (g771) & (!g711) & (!g716)) + ((g768) & (!g769) & (g770) & (g771) & (g711) & (!g716)) + ((g768) & (g769) & (!g770) & (!g771) & (!g711) & (!g716)) + ((g768) & (g769) & (!g770) & (!g771) & (!g711) & (g716)) + ((g768) & (g769) & (!g770) & (!g771) & (g711) & (g716)) + ((g768) & (g769) & (!g770) & (g771) & (!g711) & (!g716)) + ((g768) & (g769) & (!g770) & (g771) & (!g711) & (g716)) + ((g768) & (g769) & (g770) & (!g771) & (!g711) & (!g716)) + ((g768) & (g769) & (g770) & (!g771) & (g711) & (g716)) + ((g768) & (g769) & (g770) & (g771) & (!g711) & (!g716)));
	assign g774 = (((!sk[96]) & (g772) & (!g773)) + ((!sk[96]) & (g772) & (g773)) + ((sk[96]) & (!g772) & (g773)) + ((sk[96]) & (g772) & (!g773)));
	assign g781 = (((!g775) & (!g776) & (!g777) & (!g778) & (g779) & (g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g779) & (!g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g779) & (g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (g779) & (!g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (!g779) & (!g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (!g779) & (g780)) + ((!g775) & (!g776) & (g777) & (g778) & (!g779) & (!g780)) + ((!g775) & (!g776) & (g777) & (g778) & (g779) & (g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (g779) & (!g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (g779) & (g780)) + ((!g775) & (g776) & (!g777) & (g778) & (g779) & (!g780)) + ((!g775) & (g776) & (!g777) & (g778) & (g779) & (g780)) + ((!g775) & (g776) & (g777) & (!g778) & (g779) & (!g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (!g779) & (!g780)) + ((g775) & (!g776) & (g777) & (!g778) & (g779) & (!g780)) + ((g775) & (!g776) & (g777) & (g778) & (!g779) & (g780)) + ((g775) & (!g776) & (g777) & (g778) & (g779) & (g780)) + ((g775) & (g776) & (!g777) & (!g778) & (!g779) & (g780)) + ((g775) & (g776) & (!g777) & (!g778) & (g779) & (!g780)) + ((g775) & (g776) & (g777) & (!g778) & (!g779) & (g780)) + ((g775) & (g776) & (g777) & (!g778) & (g779) & (!g780)) + ((g775) & (g776) & (g777) & (g778) & (!g779) & (!g780)) + ((g775) & (g776) & (g777) & (g778) & (g779) & (!g780)) + ((g775) & (g776) & (g777) & (g778) & (g779) & (g780)));
	assign g782 = (((!g775) & (!g776) & (!g777) & (!g778) & (g779) & (!g780)) + ((!g775) & (!g776) & (!g777) & (!g778) & (g779) & (g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g779) & (!g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g779) & (g780)) + ((!g775) & (!g776) & (g777) & (g778) & (!g779) & (g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (!g779) & (!g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (!g779) & (g780)) + ((!g775) & (g776) & (g777) & (!g778) & (!g779) & (!g780)) + ((!g775) & (g776) & (g777) & (!g778) & (!g779) & (g780)) + ((!g775) & (g776) & (g777) & (!g778) & (g779) & (!g780)) + ((!g775) & (g776) & (g777) & (g778) & (g779) & (g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (!g779) & (g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (g779) & (!g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (g779) & (g780)) + ((g775) & (!g776) & (!g777) & (g778) & (g779) & (!g780)) + ((g775) & (!g776) & (g777) & (!g778) & (!g779) & (!g780)) + ((g775) & (!g776) & (g777) & (!g778) & (g779) & (g780)) + ((g775) & (!g776) & (g777) & (g778) & (!g779) & (g780)) + ((g775) & (!g776) & (g777) & (g778) & (g779) & (g780)) + ((g775) & (g776) & (!g777) & (!g778) & (!g779) & (!g780)) + ((g775) & (g776) & (!g777) & (!g778) & (!g779) & (g780)) + ((g775) & (g776) & (!g777) & (!g778) & (g779) & (!g780)) + ((g775) & (g776) & (!g777) & (!g778) & (g779) & (g780)) + ((g775) & (g776) & (!g777) & (g778) & (!g779) & (!g780)) + ((g775) & (g776) & (!g777) & (g778) & (g779) & (!g780)) + ((g775) & (g776) & (!g777) & (g778) & (g779) & (g780)) + ((g775) & (g776) & (g777) & (!g778) & (g779) & (!g780)) + ((g775) & (g776) & (g777) & (!g778) & (g779) & (g780)) + ((g775) & (g776) & (g777) & (g778) & (!g779) & (g780)) + ((g775) & (g776) & (g777) & (g778) & (g779) & (!g780)));
	assign g783 = (((!g775) & (!g776) & (!g777) & (!g778) & (!g779) & (!g780)) + ((!g775) & (!g776) & (!g777) & (!g778) & (g779) & (g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (g779) & (g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (!g779) & (!g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (!g779) & (g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (g779) & (g780)) + ((!g775) & (!g776) & (g777) & (g778) & (!g779) & (g780)) + ((!g775) & (!g776) & (g777) & (g778) & (g779) & (!g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (!g779) & (!g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (g779) & (!g780)) + ((!g775) & (g776) & (!g777) & (g778) & (g779) & (g780)) + ((!g775) & (g776) & (g777) & (g778) & (!g779) & (!g780)) + ((!g775) & (g776) & (g777) & (g778) & (g779) & (!g780)) + ((g775) & (!g776) & (!g777) & (g778) & (!g779) & (!g780)) + ((g775) & (!g776) & (!g777) & (g778) & (!g779) & (g780)) + ((g775) & (!g776) & (!g777) & (g778) & (g779) & (!g780)) + ((g775) & (!g776) & (g777) & (!g778) & (!g779) & (!g780)) + ((g775) & (!g776) & (g777) & (!g778) & (g779) & (g780)) + ((g775) & (!g776) & (g777) & (g778) & (!g779) & (!g780)) + ((g775) & (!g776) & (g777) & (g778) & (!g779) & (g780)) + ((g775) & (!g776) & (g777) & (g778) & (g779) & (!g780)) + ((g775) & (!g776) & (g777) & (g778) & (g779) & (g780)) + ((g775) & (g776) & (!g777) & (!g778) & (g779) & (g780)) + ((g775) & (g776) & (!g777) & (g778) & (!g779) & (!g780)) + ((g775) & (g776) & (!g777) & (g778) & (g779) & (!g780)) + ((g775) & (g776) & (!g777) & (g778) & (g779) & (g780)) + ((g775) & (g776) & (g777) & (!g778) & (!g779) & (!g780)) + ((g775) & (g776) & (g777) & (g778) & (!g779) & (!g780)) + ((g775) & (g776) & (g777) & (g778) & (!g779) & (g780)) + ((g775) & (g776) & (g777) & (g778) & (g779) & (g780)));
	assign g784 = (((!g775) & (!g776) & (!g777) & (!g778) & (!g779) & (g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (g779) & (!g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (g779) & (g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (!g779) & (g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (g779) & (g780)) + ((!g775) & (!g776) & (g777) & (g778) & (!g779) & (g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (!g779) & (!g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (!g779) & (g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (g779) & (!g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (g779) & (g780)) + ((!g775) & (g776) & (!g777) & (g778) & (g779) & (!g780)) + ((!g775) & (g776) & (!g777) & (g778) & (g779) & (g780)) + ((!g775) & (g776) & (g777) & (g778) & (!g779) & (!g780)) + ((!g775) & (g776) & (g777) & (g778) & (g779) & (!g780)) + ((!g775) & (g776) & (g777) & (g778) & (g779) & (g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (!g779) & (!g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (g779) & (g780)) + ((g775) & (!g776) & (!g777) & (g778) & (g779) & (!g780)) + ((g775) & (!g776) & (!g777) & (g778) & (g779) & (g780)) + ((g775) & (!g776) & (g777) & (!g778) & (!g779) & (g780)) + ((g775) & (!g776) & (g777) & (!g778) & (g779) & (!g780)) + ((g775) & (!g776) & (g777) & (g778) & (g779) & (!g780)) + ((g775) & (g776) & (!g777) & (!g778) & (!g779) & (g780)) + ((g775) & (g776) & (!g777) & (!g778) & (g779) & (g780)) + ((g775) & (g776) & (!g777) & (g778) & (g779) & (!g780)) + ((g775) & (g776) & (!g777) & (g778) & (g779) & (g780)) + ((g775) & (g776) & (g777) & (!g778) & (!g779) & (g780)) + ((g775) & (g776) & (g777) & (g778) & (!g779) & (!g780)));
	assign g787 = (((!g781) & (!g782) & (!g783) & (!g784) & (!g785) & (!g786)) + ((!g781) & (!g782) & (!g783) & (g784) & (!g785) & (!g786)) + ((!g781) & (!g782) & (!g783) & (g784) & (g785) & (g786)) + ((!g781) & (!g782) & (g783) & (!g784) & (!g785) & (!g786)) + ((!g781) & (!g782) & (g783) & (!g784) & (!g785) & (g786)) + ((!g781) & (!g782) & (g783) & (g784) & (!g785) & (!g786)) + ((!g781) & (!g782) & (g783) & (g784) & (!g785) & (g786)) + ((!g781) & (!g782) & (g783) & (g784) & (g785) & (g786)) + ((!g781) & (g782) & (!g783) & (!g784) & (!g785) & (!g786)) + ((!g781) & (g782) & (!g783) & (!g784) & (g785) & (!g786)) + ((!g781) & (g782) & (!g783) & (g784) & (!g785) & (!g786)) + ((!g781) & (g782) & (!g783) & (g784) & (g785) & (!g786)) + ((!g781) & (g782) & (!g783) & (g784) & (g785) & (g786)) + ((!g781) & (g782) & (g783) & (!g784) & (!g785) & (!g786)) + ((!g781) & (g782) & (g783) & (!g784) & (!g785) & (g786)) + ((!g781) & (g782) & (g783) & (!g784) & (g785) & (!g786)) + ((!g781) & (g782) & (g783) & (g784) & (!g785) & (!g786)) + ((!g781) & (g782) & (g783) & (g784) & (!g785) & (g786)) + ((!g781) & (g782) & (g783) & (g784) & (g785) & (!g786)) + ((!g781) & (g782) & (g783) & (g784) & (g785) & (g786)) + ((g781) & (!g782) & (!g783) & (g784) & (g785) & (g786)) + ((g781) & (!g782) & (g783) & (!g784) & (!g785) & (g786)) + ((g781) & (!g782) & (g783) & (g784) & (!g785) & (g786)) + ((g781) & (!g782) & (g783) & (g784) & (g785) & (g786)) + ((g781) & (g782) & (!g783) & (!g784) & (g785) & (!g786)) + ((g781) & (g782) & (!g783) & (g784) & (g785) & (!g786)) + ((g781) & (g782) & (!g783) & (g784) & (g785) & (g786)) + ((g781) & (g782) & (g783) & (!g784) & (!g785) & (g786)) + ((g781) & (g782) & (g783) & (!g784) & (g785) & (!g786)) + ((g781) & (g782) & (g783) & (g784) & (!g785) & (g786)) + ((g781) & (g782) & (g783) & (g784) & (g785) & (!g786)) + ((g781) & (g782) & (g783) & (g784) & (g785) & (g786)));
	assign g789 = (((!sk[102]) & (g787) & (!g788)) + ((!sk[102]) & (g787) & (g788)) + ((sk[102]) & (!g787) & (g788)) + ((sk[102]) & (g787) & (!g788)));
	assign g790 = (((!g775) & (!g776) & (!g777) & (!g778) & (!g785) & (g779)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g785) & (!g779)) + ((!g775) & (!g776) & (!g777) & (g778) & (g785) & (!g779)) + ((!g775) & (!g776) & (g777) & (!g778) & (g785) & (g779)) + ((!g775) & (!g776) & (g777) & (g778) & (!g785) & (g779)) + ((!g775) & (!g776) & (g777) & (g778) & (g785) & (!g779)) + ((!g775) & (g776) & (!g777) & (!g778) & (!g785) & (g779)) + ((!g775) & (g776) & (!g777) & (!g778) & (g785) & (!g779)) + ((!g775) & (g776) & (!g777) & (!g778) & (g785) & (g779)) + ((!g775) & (g776) & (g777) & (!g778) & (g785) & (g779)) + ((!g775) & (g776) & (g777) & (g778) & (g785) & (g779)) + ((g775) & (!g776) & (!g777) & (!g778) & (!g785) & (!g779)) + ((g775) & (!g776) & (!g777) & (!g778) & (g785) & (g779)) + ((g775) & (!g776) & (!g777) & (g778) & (!g785) & (!g779)) + ((g775) & (!g776) & (!g777) & (g778) & (g785) & (!g779)) + ((g775) & (!g776) & (g777) & (!g778) & (g785) & (!g779)) + ((g775) & (!g776) & (g777) & (!g778) & (g785) & (g779)) + ((g775) & (!g776) & (g777) & (g778) & (g785) & (!g779)) + ((g775) & (!g776) & (g777) & (g778) & (g785) & (g779)) + ((g775) & (g776) & (!g777) & (!g778) & (g785) & (!g779)) + ((g775) & (g776) & (!g777) & (!g778) & (g785) & (g779)) + ((g775) & (g776) & (!g777) & (g778) & (g785) & (g779)) + ((g775) & (g776) & (g777) & (!g778) & (!g785) & (!g779)) + ((g775) & (g776) & (g777) & (!g778) & (!g785) & (g779)) + ((g775) & (g776) & (g777) & (!g778) & (g785) & (!g779)) + ((g775) & (g776) & (g777) & (g778) & (!g785) & (g779)) + ((g775) & (g776) & (g777) & (g778) & (g785) & (!g779)));
	assign g791 = (((!g775) & (!g776) & (!g777) & (!g778) & (!g785) & (g779)) + ((!g775) & (!g776) & (!g777) & (!g778) & (g785) & (!g779)) + ((!g775) & (!g776) & (!g777) & (!g778) & (g785) & (g779)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g785) & (!g779)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g785) & (g779)) + ((!g775) & (!g776) & (!g777) & (g778) & (g785) & (g779)) + ((!g775) & (!g776) & (g777) & (!g778) & (g785) & (!g779)) + ((!g775) & (!g776) & (g777) & (g778) & (!g785) & (!g779)) + ((!g775) & (!g776) & (g777) & (g778) & (!g785) & (g779)) + ((!g775) & (!g776) & (g777) & (g778) & (g785) & (g779)) + ((!g775) & (g776) & (!g777) & (!g778) & (g785) & (g779)) + ((!g775) & (g776) & (!g777) & (g778) & (!g785) & (!g779)) + ((!g775) & (g776) & (!g777) & (g778) & (g785) & (!g779)) + ((!g775) & (g776) & (g777) & (!g778) & (g785) & (!g779)) + ((!g775) & (g776) & (g777) & (!g778) & (g785) & (g779)) + ((!g775) & (g776) & (g777) & (g778) & (!g785) & (!g779)) + ((g775) & (!g776) & (!g777) & (!g778) & (!g785) & (!g779)) + ((g775) & (!g776) & (!g777) & (g778) & (!g785) & (!g779)) + ((g775) & (!g776) & (!g777) & (g778) & (!g785) & (g779)) + ((g775) & (!g776) & (g777) & (!g778) & (!g785) & (g779)) + ((g775) & (!g776) & (g777) & (!g778) & (g785) & (g779)) + ((g775) & (!g776) & (g777) & (g778) & (!g785) & (!g779)) + ((g775) & (!g776) & (g777) & (g778) & (!g785) & (g779)) + ((g775) & (g776) & (!g777) & (g778) & (!g785) & (!g779)) + ((g775) & (g776) & (!g777) & (g778) & (g785) & (g779)) + ((g775) & (g776) & (g777) & (!g778) & (!g785) & (!g779)) + ((g775) & (g776) & (g777) & (!g778) & (!g785) & (g779)) + ((g775) & (g776) & (g777) & (!g778) & (g785) & (g779)) + ((g775) & (g776) & (g777) & (g778) & (!g785) & (!g779)) + ((g775) & (g776) & (g777) & (g778) & (!g785) & (g779)) + ((g775) & (g776) & (g777) & (g778) & (g785) & (!g779)));
	assign g792 = (((!g775) & (!g776) & (!g777) & (!g778) & (!g785) & (g779)) + ((!g775) & (!g776) & (!g777) & (g778) & (g785) & (!g779)) + ((!g775) & (!g776) & (g777) & (!g778) & (!g785) & (!g779)) + ((!g775) & (!g776) & (g777) & (!g778) & (g785) & (!g779)) + ((!g775) & (!g776) & (g777) & (g778) & (!g785) & (g779)) + ((!g775) & (!g776) & (g777) & (g778) & (g785) & (!g779)) + ((!g775) & (!g776) & (g777) & (g778) & (g785) & (g779)) + ((!g775) & (g776) & (!g777) & (!g778) & (!g785) & (!g779)) + ((!g775) & (g776) & (!g777) & (!g778) & (g785) & (!g779)) + ((!g775) & (g776) & (!g777) & (g778) & (!g785) & (!g779)) + ((!g775) & (g776) & (!g777) & (g778) & (g785) & (g779)) + ((!g775) & (g776) & (g777) & (!g778) & (g785) & (g779)) + ((!g775) & (g776) & (g777) & (g778) & (!g785) & (g779)) + ((!g775) & (g776) & (g777) & (g778) & (g785) & (!g779)) + ((g775) & (!g776) & (!g777) & (!g778) & (g785) & (g779)) + ((g775) & (!g776) & (!g777) & (g778) & (!g785) & (!g779)) + ((g775) & (!g776) & (!g777) & (g778) & (g785) & (!g779)) + ((g775) & (!g776) & (g777) & (!g778) & (!g785) & (!g779)) + ((g775) & (!g776) & (g777) & (!g778) & (!g785) & (g779)) + ((g775) & (!g776) & (g777) & (!g778) & (g785) & (!g779)) + ((g775) & (!g776) & (g777) & (!g778) & (g785) & (g779)) + ((g775) & (!g776) & (g777) & (g778) & (g785) & (!g779)) + ((g775) & (g776) & (!g777) & (!g778) & (!g785) & (g779)) + ((g775) & (g776) & (!g777) & (!g778) & (g785) & (g779)) + ((g775) & (g776) & (!g777) & (g778) & (!g785) & (g779)) + ((g775) & (g776) & (g777) & (!g778) & (!g785) & (!g779)) + ((g775) & (g776) & (g777) & (!g778) & (!g785) & (g779)) + ((g775) & (g776) & (g777) & (!g778) & (g785) & (g779)) + ((g775) & (g776) & (g777) & (g778) & (!g785) & (!g779)) + ((g775) & (g776) & (g777) & (g778) & (!g785) & (g779)) + ((g775) & (g776) & (g777) & (g778) & (g785) & (!g779)) + ((g775) & (g776) & (g777) & (g778) & (g785) & (g779)));
	assign g793 = (((!g775) & (!g776) & (!g777) & (!g778) & (g785) & (!g779)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g785) & (!g779)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g785) & (g779)) + ((!g775) & (!g776) & (g777) & (!g778) & (g785) & (g779)) + ((!g775) & (!g776) & (g777) & (g778) & (!g785) & (g779)) + ((!g775) & (g776) & (!g777) & (!g778) & (!g785) & (!g779)) + ((!g775) & (g776) & (!g777) & (!g778) & (g785) & (!g779)) + ((!g775) & (g776) & (!g777) & (g778) & (!g785) & (g779)) + ((!g775) & (g776) & (g777) & (!g778) & (!g785) & (g779)) + ((!g775) & (g776) & (g777) & (!g778) & (g785) & (!g779)) + ((!g775) & (g776) & (g777) & (!g778) & (g785) & (g779)) + ((!g775) & (g776) & (g777) & (g778) & (g785) & (!g779)) + ((!g775) & (g776) & (g777) & (g778) & (g785) & (g779)) + ((g775) & (!g776) & (!g777) & (!g778) & (!g785) & (!g779)) + ((g775) & (!g776) & (!g777) & (g778) & (!g785) & (!g779)) + ((g775) & (!g776) & (!g777) & (g778) & (!g785) & (g779)) + ((g775) & (!g776) & (!g777) & (g778) & (g785) & (!g779)) + ((g775) & (!g776) & (g777) & (!g778) & (!g785) & (!g779)) + ((g775) & (!g776) & (g777) & (!g778) & (g785) & (g779)) + ((g775) & (!g776) & (g777) & (g778) & (g785) & (!g779)) + ((g775) & (g776) & (!g777) & (!g778) & (!g785) & (!g779)) + ((g775) & (g776) & (!g777) & (g778) & (!g785) & (!g779)) + ((g775) & (g776) & (!g777) & (g778) & (g785) & (!g779)) + ((g775) & (g776) & (!g777) & (g778) & (g785) & (g779)) + ((g775) & (g776) & (g777) & (g778) & (!g785) & (g779)) + ((g775) & (g776) & (g777) & (g778) & (g785) & (g779)));
	assign g794 = (((!g790) & (!g791) & (!g792) & (!g793) & (!g780) & (!g786)) + ((!g790) & (!g791) & (!g792) & (!g793) & (g780) & (!g786)) + ((!g790) & (!g791) & (!g792) & (g793) & (!g780) & (!g786)) + ((!g790) & (!g791) & (!g792) & (g793) & (g780) & (!g786)) + ((!g790) & (!g791) & (!g792) & (g793) & (g780) & (g786)) + ((!g790) & (!g791) & (g792) & (!g793) & (!g780) & (!g786)) + ((!g790) & (!g791) & (g792) & (!g793) & (!g780) & (g786)) + ((!g790) & (!g791) & (g792) & (!g793) & (g780) & (!g786)) + ((!g790) & (!g791) & (g792) & (g793) & (!g780) & (!g786)) + ((!g790) & (!g791) & (g792) & (g793) & (!g780) & (g786)) + ((!g790) & (!g791) & (g792) & (g793) & (g780) & (!g786)) + ((!g790) & (!g791) & (g792) & (g793) & (g780) & (g786)) + ((!g790) & (g791) & (!g792) & (!g793) & (!g780) & (!g786)) + ((!g790) & (g791) & (!g792) & (g793) & (!g780) & (!g786)) + ((!g790) & (g791) & (!g792) & (g793) & (g780) & (g786)) + ((!g790) & (g791) & (g792) & (!g793) & (!g780) & (!g786)) + ((!g790) & (g791) & (g792) & (!g793) & (!g780) & (g786)) + ((!g790) & (g791) & (g792) & (g793) & (!g780) & (!g786)) + ((!g790) & (g791) & (g792) & (g793) & (!g780) & (g786)) + ((!g790) & (g791) & (g792) & (g793) & (g780) & (g786)) + ((g790) & (!g791) & (!g792) & (!g793) & (g780) & (!g786)) + ((g790) & (!g791) & (!g792) & (g793) & (g780) & (!g786)) + ((g790) & (!g791) & (!g792) & (g793) & (g780) & (g786)) + ((g790) & (!g791) & (g792) & (!g793) & (!g780) & (g786)) + ((g790) & (!g791) & (g792) & (!g793) & (g780) & (!g786)) + ((g790) & (!g791) & (g792) & (g793) & (!g780) & (g786)) + ((g790) & (!g791) & (g792) & (g793) & (g780) & (!g786)) + ((g790) & (!g791) & (g792) & (g793) & (g780) & (g786)) + ((g790) & (g791) & (!g792) & (g793) & (g780) & (g786)) + ((g790) & (g791) & (g792) & (!g793) & (!g780) & (g786)) + ((g790) & (g791) & (g792) & (g793) & (!g780) & (g786)) + ((g790) & (g791) & (g792) & (g793) & (g780) & (g786)));
	assign g796 = (((!sk[108]) & (g794) & (!g795)) + ((!sk[108]) & (g794) & (g795)) + ((sk[108]) & (!g794) & (g795)) + ((sk[108]) & (g794) & (!g795)));
	assign g797 = (((!g779) & (!g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((!g779) & (!g776) & (!g777) & (!g778) & (g785) & (g780)) + ((!g779) & (!g776) & (!g777) & (g778) & (!g785) & (g780)) + ((!g779) & (!g776) & (!g777) & (g778) & (g785) & (!g780)) + ((!g779) & (!g776) & (!g777) & (g778) & (g785) & (g780)) + ((!g779) & (!g776) & (g777) & (!g778) & (!g785) & (g780)) + ((!g779) & (!g776) & (g777) & (g778) & (!g785) & (!g780)) + ((!g779) & (!g776) & (g777) & (g778) & (g785) & (!g780)) + ((!g779) & (g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((!g779) & (g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((!g779) & (g776) & (!g777) & (g778) & (!g785) & (g780)) + ((!g779) & (g776) & (g777) & (!g778) & (!g785) & (!g780)) + ((!g779) & (g776) & (g777) & (!g778) & (!g785) & (g780)) + ((!g779) & (g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g779) & (g776) & (g777) & (!g778) & (g785) & (g780)) + ((g779) & (!g776) & (!g777) & (g778) & (!g785) & (g780)) + ((g779) & (!g776) & (!g777) & (g778) & (g785) & (g780)) + ((g779) & (g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((g779) & (g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((g779) & (g776) & (!g777) & (g778) & (g785) & (!g780)) + ((g779) & (g776) & (g777) & (g778) & (!g785) & (!g780)) + ((g779) & (g776) & (g777) & (g778) & (!g785) & (g780)));
	assign g798 = (((!g779) & (!g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((!g779) & (!g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((!g779) & (!g776) & (!g777) & (g778) & (g785) & (g780)) + ((!g779) & (!g776) & (g777) & (!g778) & (!g785) & (!g780)) + ((!g779) & (!g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g779) & (!g776) & (g777) & (g778) & (!g785) & (g780)) + ((!g779) & (g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((!g779) & (g776) & (!g777) & (!g778) & (g785) & (g780)) + ((!g779) & (g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((!g779) & (g776) & (!g777) & (g778) & (!g785) & (g780)) + ((!g779) & (g776) & (!g777) & (g778) & (g785) & (g780)) + ((!g779) & (g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g779) & (g776) & (g777) & (!g778) & (g785) & (g780)) + ((!g779) & (g776) & (g777) & (g778) & (g785) & (!g780)) + ((g779) & (!g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((g779) & (!g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((g779) & (!g776) & (!g777) & (!g778) & (g785) & (g780)) + ((g779) & (!g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((g779) & (!g776) & (!g777) & (g778) & (!g785) & (g780)) + ((g779) & (!g776) & (!g777) & (g778) & (g785) & (!g780)) + ((g779) & (!g776) & (g777) & (g778) & (!g785) & (!g780)) + ((g779) & (g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((g779) & (g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((g779) & (g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((g779) & (g776) & (!g777) & (g778) & (g785) & (!g780)) + ((g779) & (g776) & (!g777) & (g778) & (g785) & (g780)) + ((g779) & (g776) & (g777) & (!g778) & (!g785) & (!g780)) + ((g779) & (g776) & (g777) & (!g778) & (g785) & (!g780)) + ((g779) & (g776) & (g777) & (g778) & (!g785) & (g780)) + ((g779) & (g776) & (g777) & (g778) & (g785) & (g780)));
	assign g799 = (((!g779) & (!g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((!g779) & (!g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((!g779) & (!g776) & (!g777) & (g778) & (!g785) & (g780)) + ((!g779) & (!g776) & (g777) & (!g778) & (!g785) & (g780)) + ((!g779) & (!g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g779) & (!g776) & (g777) & (g778) & (!g785) & (g780)) + ((!g779) & (g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((!g779) & (g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((!g779) & (g776) & (!g777) & (g778) & (g785) & (!g780)) + ((!g779) & (g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g779) & (g776) & (g777) & (g778) & (!g785) & (!g780)) + ((!g779) & (g776) & (g777) & (g778) & (g785) & (!g780)) + ((g779) & (!g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((g779) & (!g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((g779) & (!g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((g779) & (!g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((g779) & (!g776) & (!g777) & (g778) & (!g785) & (g780)) + ((g779) & (!g776) & (!g777) & (g778) & (g785) & (!g780)) + ((g779) & (!g776) & (!g777) & (g778) & (g785) & (g780)) + ((g779) & (!g776) & (g777) & (!g778) & (!g785) & (g780)) + ((g779) & (!g776) & (g777) & (!g778) & (g785) & (!g780)) + ((g779) & (!g776) & (g777) & (g778) & (!g785) & (!g780)) + ((g779) & (!g776) & (g777) & (g778) & (g785) & (g780)) + ((g779) & (g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((g779) & (g776) & (!g777) & (!g778) & (g785) & (g780)) + ((g779) & (g776) & (g777) & (!g778) & (g785) & (g780)) + ((g779) & (g776) & (g777) & (g778) & (!g785) & (!g780)) + ((g779) & (g776) & (g777) & (g778) & (!g785) & (g780)) + ((g779) & (g776) & (g777) & (g778) & (g785) & (g780)));
	assign g800 = (((!g779) & (!g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((!g779) & (!g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((!g779) & (!g776) & (!g777) & (!g778) & (g785) & (g780)) + ((!g779) & (!g776) & (!g777) & (g778) & (!g785) & (g780)) + ((!g779) & (!g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g779) & (!g776) & (g777) & (g778) & (g785) & (g780)) + ((!g779) & (g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((!g779) & (g776) & (!g777) & (g778) & (!g785) & (g780)) + ((!g779) & (g776) & (!g777) & (g778) & (g785) & (g780)) + ((!g779) & (g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g779) & (g776) & (g777) & (!g778) & (g785) & (g780)) + ((!g779) & (g776) & (g777) & (g778) & (!g785) & (!g780)) + ((!g779) & (g776) & (g777) & (g778) & (!g785) & (g780)) + ((!g779) & (g776) & (g777) & (g778) & (g785) & (!g780)) + ((!g779) & (g776) & (g777) & (g778) & (g785) & (g780)) + ((g779) & (!g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((g779) & (!g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((g779) & (!g776) & (!g777) & (!g778) & (g785) & (g780)) + ((g779) & (!g776) & (!g777) & (g778) & (g785) & (g780)) + ((g779) & (!g776) & (g777) & (!g778) & (!g785) & (g780)) + ((g779) & (!g776) & (g777) & (!g778) & (g785) & (!g780)) + ((g779) & (!g776) & (g777) & (g778) & (g785) & (!g780)) + ((g779) & (g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((g779) & (g776) & (!g777) & (g778) & (!g785) & (g780)) + ((g779) & (g776) & (!g777) & (g778) & (g785) & (!g780)) + ((g779) & (g776) & (g777) & (!g778) & (g785) & (g780)) + ((g779) & (g776) & (g777) & (g778) & (!g785) & (!g780)));
	assign g801 = (((!g797) & (!g798) & (!g799) & (!g800) & (!g775) & (g786)) + ((!g797) & (!g798) & (!g799) & (!g800) & (g775) & (!g786)) + ((!g797) & (!g798) & (!g799) & (!g800) & (g775) & (g786)) + ((!g797) & (!g798) & (!g799) & (g800) & (!g775) & (g786)) + ((!g797) & (!g798) & (!g799) & (g800) & (g775) & (!g786)) + ((!g797) & (!g798) & (g799) & (!g800) & (g775) & (!g786)) + ((!g797) & (!g798) & (g799) & (!g800) & (g775) & (g786)) + ((!g797) & (!g798) & (g799) & (g800) & (g775) & (!g786)) + ((!g797) & (g798) & (!g799) & (!g800) & (!g775) & (g786)) + ((!g797) & (g798) & (!g799) & (!g800) & (g775) & (g786)) + ((!g797) & (g798) & (!g799) & (g800) & (!g775) & (g786)) + ((!g797) & (g798) & (g799) & (!g800) & (g775) & (g786)) + ((g797) & (!g798) & (!g799) & (!g800) & (!g775) & (!g786)) + ((g797) & (!g798) & (!g799) & (!g800) & (!g775) & (g786)) + ((g797) & (!g798) & (!g799) & (!g800) & (g775) & (!g786)) + ((g797) & (!g798) & (!g799) & (!g800) & (g775) & (g786)) + ((g797) & (!g798) & (!g799) & (g800) & (!g775) & (!g786)) + ((g797) & (!g798) & (!g799) & (g800) & (!g775) & (g786)) + ((g797) & (!g798) & (!g799) & (g800) & (g775) & (!g786)) + ((g797) & (!g798) & (g799) & (!g800) & (!g775) & (!g786)) + ((g797) & (!g798) & (g799) & (!g800) & (g775) & (!g786)) + ((g797) & (!g798) & (g799) & (!g800) & (g775) & (g786)) + ((g797) & (!g798) & (g799) & (g800) & (!g775) & (!g786)) + ((g797) & (!g798) & (g799) & (g800) & (g775) & (!g786)) + ((g797) & (g798) & (!g799) & (!g800) & (!g775) & (!g786)) + ((g797) & (g798) & (!g799) & (!g800) & (!g775) & (g786)) + ((g797) & (g798) & (!g799) & (!g800) & (g775) & (g786)) + ((g797) & (g798) & (!g799) & (g800) & (!g775) & (!g786)) + ((g797) & (g798) & (!g799) & (g800) & (!g775) & (g786)) + ((g797) & (g798) & (g799) & (!g800) & (!g775) & (!g786)) + ((g797) & (g798) & (g799) & (!g800) & (g775) & (g786)) + ((g797) & (g798) & (g799) & (g800) & (!g775) & (!g786)));
	assign g803 = (((!g801) & (sk[114]) & (g802)) + ((g801) & (!sk[114]) & (!g802)) + ((g801) & (!sk[114]) & (g802)) + ((g801) & (sk[114]) & (!g802)));
	assign g804 = (((!g775) & (!g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (g785) & (g780)) + ((!g775) & (!g776) & (g777) & (g778) & (!g785) & (!g780)) + ((!g775) & (!g776) & (g777) & (g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (g777) & (g778) & (g785) & (g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (g776) & (g777) & (!g778) & (!g785) & (!g780)) + ((!g775) & (g776) & (g777) & (g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((g775) & (!g776) & (g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (g777) & (!g778) & (!g785) & (g780)) + ((g775) & (!g776) & (g777) & (!g778) & (g785) & (!g780)) + ((g775) & (!g776) & (g777) & (g778) & (!g785) & (g780)) + ((g775) & (g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((g775) & (g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((g775) & (g776) & (!g777) & (g778) & (g785) & (!g780)) + ((g775) & (g776) & (g777) & (!g778) & (!g785) & (g780)) + ((g775) & (g776) & (g777) & (!g778) & (g785) & (g780)));
	assign g805 = (((!g775) & (!g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (!g777) & (!g778) & (g785) & (g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (g777) & (g778) & (!g785) & (!g780)) + ((!g775) & (!g776) & (g777) & (g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (g777) & (g778) & (g785) & (g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (g785) & (g780)) + ((!g775) & (g776) & (!g777) & (g778) & (g785) & (g780)) + ((!g775) & (g776) & (g777) & (!g778) & (!g785) & (!g780)) + ((!g775) & (g776) & (g777) & (!g778) & (!g785) & (g780)) + ((!g775) & (g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (g776) & (g777) & (g778) & (!g785) & (g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((g775) & (!g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (!g777) & (g778) & (!g785) & (g780)) + ((g775) & (!g776) & (!g777) & (g778) & (g785) & (g780)) + ((g775) & (!g776) & (g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (g777) & (!g778) & (!g785) & (g780)) + ((g775) & (!g776) & (g777) & (!g778) & (g785) & (g780)) + ((g775) & (!g776) & (g777) & (g778) & (!g785) & (g780)) + ((g775) & (g776) & (!g777) & (g778) & (!g785) & (g780)) + ((g775) & (g776) & (!g777) & (g778) & (g785) & (!g780)) + ((g775) & (g776) & (g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (g776) & (g777) & (g778) & (!g785) & (!g780)));
	assign g806 = (((!g775) & (!g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (!g777) & (!g778) & (g785) & (g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (g777) & (!g778) & (g785) & (g780)) + ((!g775) & (!g776) & (g777) & (g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (g777) & (g778) & (g785) & (g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (g785) & (g780)) + ((!g775) & (g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((!g775) & (g776) & (!g777) & (g778) & (!g785) & (g780)) + ((!g775) & (g776) & (g777) & (!g778) & (!g785) & (g780)) + ((!g775) & (g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (g776) & (g777) & (g778) & (g785) & (g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (g785) & (g780)) + ((g775) & (!g776) & (!g777) & (g778) & (g785) & (g780)) + ((g775) & (!g776) & (g777) & (g778) & (!g785) & (!g780)) + ((g775) & (g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((g775) & (g776) & (!g777) & (g778) & (g785) & (g780)) + ((g775) & (g776) & (g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (g776) & (g777) & (!g778) & (!g785) & (g780)) + ((g775) & (g776) & (g777) & (!g778) & (g785) & (g780)) + ((g775) & (g776) & (g777) & (g778) & (!g785) & (!g780)) + ((g775) & (g776) & (g777) & (g778) & (g785) & (g780)));
	assign g807 = (((!g775) & (!g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (!g777) & (g778) & (g785) & (g780)) + ((!g775) & (!g776) & (g777) & (g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (g777) & (g778) & (g785) & (g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (!g785) & (!g780)) + ((!g775) & (g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (g776) & (!g777) & (g778) & (!g785) & (!g780)) + ((!g775) & (g776) & (!g777) & (g778) & (!g785) & (g780)) + ((!g775) & (g776) & (!g777) & (g778) & (g785) & (!g780)) + ((!g775) & (g776) & (g777) & (!g778) & (!g785) & (!g780)) + ((!g775) & (g776) & (g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (g776) & (g777) & (!g778) & (g785) & (g780)) + ((g775) & (!g776) & (!g777) & (!g778) & (g785) & (g780)) + ((g775) & (!g776) & (!g777) & (g778) & (g785) & (!g780)) + ((g775) & (!g776) & (g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (g777) & (!g778) & (g785) & (!g780)) + ((g775) & (!g776) & (g777) & (!g778) & (g785) & (g780)) + ((g775) & (!g776) & (g777) & (g778) & (!g785) & (g780)) + ((g775) & (!g776) & (g777) & (g778) & (g785) & (!g780)) + ((g775) & (!g776) & (g777) & (g778) & (g785) & (g780)) + ((g775) & (g776) & (!g777) & (!g778) & (!g785) & (g780)) + ((g775) & (g776) & (!g777) & (!g778) & (g785) & (!g780)) + ((g775) & (g776) & (g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (g776) & (g777) & (!g778) & (!g785) & (g780)) + ((g775) & (g776) & (g777) & (g778) & (g785) & (g780)));
	assign g808 = (((!g804) & (!g805) & (!g806) & (!g807) & (!g786) & (g779)) + ((!g804) & (!g805) & (!g806) & (!g807) & (g786) & (!g779)) + ((!g804) & (!g805) & (!g806) & (!g807) & (g786) & (g779)) + ((!g804) & (!g805) & (!g806) & (g807) & (!g786) & (g779)) + ((!g804) & (!g805) & (!g806) & (g807) & (g786) & (!g779)) + ((!g804) & (!g805) & (g806) & (!g807) & (g786) & (!g779)) + ((!g804) & (!g805) & (g806) & (!g807) & (g786) & (g779)) + ((!g804) & (!g805) & (g806) & (g807) & (g786) & (!g779)) + ((!g804) & (g805) & (!g806) & (!g807) & (!g786) & (g779)) + ((!g804) & (g805) & (!g806) & (!g807) & (g786) & (g779)) + ((!g804) & (g805) & (!g806) & (g807) & (!g786) & (g779)) + ((!g804) & (g805) & (g806) & (!g807) & (g786) & (g779)) + ((g804) & (!g805) & (!g806) & (!g807) & (!g786) & (!g779)) + ((g804) & (!g805) & (!g806) & (!g807) & (!g786) & (g779)) + ((g804) & (!g805) & (!g806) & (!g807) & (g786) & (!g779)) + ((g804) & (!g805) & (!g806) & (!g807) & (g786) & (g779)) + ((g804) & (!g805) & (!g806) & (g807) & (!g786) & (!g779)) + ((g804) & (!g805) & (!g806) & (g807) & (!g786) & (g779)) + ((g804) & (!g805) & (!g806) & (g807) & (g786) & (!g779)) + ((g804) & (!g805) & (g806) & (!g807) & (!g786) & (!g779)) + ((g804) & (!g805) & (g806) & (!g807) & (g786) & (!g779)) + ((g804) & (!g805) & (g806) & (!g807) & (g786) & (g779)) + ((g804) & (!g805) & (g806) & (g807) & (!g786) & (!g779)) + ((g804) & (!g805) & (g806) & (g807) & (g786) & (!g779)) + ((g804) & (g805) & (!g806) & (!g807) & (!g786) & (!g779)) + ((g804) & (g805) & (!g806) & (!g807) & (!g786) & (g779)) + ((g804) & (g805) & (!g806) & (!g807) & (g786) & (g779)) + ((g804) & (g805) & (!g806) & (g807) & (!g786) & (!g779)) + ((g804) & (g805) & (!g806) & (g807) & (!g786) & (g779)) + ((g804) & (g805) & (g806) & (!g807) & (!g786) & (!g779)) + ((g804) & (g805) & (g806) & (!g807) & (g786) & (g779)) + ((g804) & (g805) & (g806) & (g807) & (!g786) & (!g779)));
	assign g810 = (((!sk[120]) & (g808) & (!g809)) + ((!sk[120]) & (g808) & (g809)) + ((sk[120]) & (!g808) & (g809)) + ((sk[120]) & (g808) & (!g809)));
	assign g811 = (((!g775) & (!g776) & (!g779) & (!g786) & (!g785) & (g780)) + ((!g775) & (!g776) & (g779) & (!g786) & (!g785) & (g780)) + ((!g775) & (!g776) & (g779) & (!g786) & (g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (!g786) & (g785) & (g780)) + ((!g775) & (!g776) & (g779) & (g786) & (!g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (g786) & (g785) & (!g780)) + ((!g775) & (g776) & (!g779) & (!g786) & (!g785) & (!g780)) + ((!g775) & (g776) & (!g779) & (!g786) & (!g785) & (g780)) + ((!g775) & (g776) & (!g779) & (g786) & (!g785) & (!g780)) + ((!g775) & (g776) & (!g779) & (g786) & (!g785) & (g780)) + ((!g775) & (g776) & (!g779) & (g786) & (g785) & (g780)) + ((!g775) & (g776) & (g779) & (g786) & (!g785) & (g780)) + ((!g775) & (g776) & (g779) & (g786) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g786) & (!g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g786) & (!g785) & (g780)) + ((g775) & (!g776) & (!g779) & (g786) & (!g785) & (g780)) + ((g775) & (!g776) & (g779) & (!g786) & (g785) & (!g780)) + ((g775) & (!g776) & (g779) & (g786) & (!g785) & (!g780)) + ((g775) & (!g776) & (g779) & (g786) & (!g785) & (g780)) + ((g775) & (!g776) & (g779) & (g786) & (g785) & (!g780)) + ((g775) & (g776) & (!g779) & (!g786) & (!g785) & (!g780)) + ((g775) & (g776) & (!g779) & (!g786) & (g785) & (!g780)) + ((g775) & (g776) & (!g779) & (g786) & (g785) & (!g780)) + ((g775) & (g776) & (g779) & (!g786) & (!g785) & (!g780)) + ((g775) & (g776) & (g779) & (!g786) & (!g785) & (g780)) + ((g775) & (g776) & (g779) & (g786) & (!g785) & (g780)));
	assign g812 = (((!g775) & (!g776) & (!g779) & (!g786) & (!g785) & (!g780)) + ((!g775) & (!g776) & (!g779) & (!g786) & (!g785) & (g780)) + ((!g775) & (!g776) & (!g779) & (!g786) & (g785) & (!g780)) + ((!g775) & (!g776) & (!g779) & (!g786) & (g785) & (g780)) + ((!g775) & (!g776) & (!g779) & (g786) & (!g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (!g786) & (!g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (!g786) & (g785) & (g780)) + ((!g775) & (!g776) & (g779) & (g786) & (!g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (g786) & (g785) & (g780)) + ((!g775) & (g776) & (!g779) & (!g786) & (!g785) & (g780)) + ((!g775) & (g776) & (!g779) & (g786) & (g785) & (!g780)) + ((!g775) & (g776) & (g779) & (!g786) & (!g785) & (!g780)) + ((!g775) & (g776) & (g779) & (!g786) & (!g785) & (g780)) + ((!g775) & (g776) & (g779) & (!g786) & (g785) & (!g780)) + ((!g775) & (g776) & (g779) & (!g786) & (g785) & (g780)) + ((!g775) & (g776) & (g779) & (g786) & (!g785) & (!g780)) + ((!g775) & (g776) & (g779) & (g786) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g786) & (!g785) & (g780)) + ((g775) & (!g776) & (!g779) & (!g786) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g786) & (g785) & (g780)) + ((g775) & (!g776) & (!g779) & (g786) & (!g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (g786) & (g785) & (g780)) + ((g775) & (!g776) & (g779) & (!g786) & (g785) & (!g780)) + ((g775) & (!g776) & (g779) & (!g786) & (g785) & (g780)) + ((g775) & (!g776) & (g779) & (g786) & (!g785) & (g780)) + ((g775) & (g776) & (!g779) & (!g786) & (g785) & (!g780)) + ((g775) & (g776) & (!g779) & (!g786) & (g785) & (g780)) + ((g775) & (g776) & (!g779) & (g786) & (!g785) & (!g780)) + ((g775) & (g776) & (!g779) & (g786) & (!g785) & (g780)) + ((g775) & (g776) & (g779) & (!g786) & (g785) & (!g780)) + ((g775) & (g776) & (g779) & (!g786) & (g785) & (g780)) + ((g775) & (g776) & (g779) & (g786) & (!g785) & (g780)));
	assign g813 = (((!g775) & (!g776) & (!g779) & (!g786) & (!g785) & (!g780)) + ((!g775) & (!g776) & (!g779) & (!g786) & (!g785) & (g780)) + ((!g775) & (!g776) & (g779) & (!g786) & (!g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (!g786) & (g785) & (g780)) + ((!g775) & (!g776) & (g779) & (g786) & (!g785) & (g780)) + ((!g775) & (g776) & (!g779) & (g786) & (!g785) & (!g780)) + ((!g775) & (g776) & (!g779) & (g786) & (g785) & (!g780)) + ((!g775) & (g776) & (!g779) & (g786) & (g785) & (g780)) + ((!g775) & (g776) & (g779) & (!g786) & (!g785) & (!g780)) + ((!g775) & (g776) & (g779) & (!g786) & (g785) & (!g780)) + ((!g775) & (g776) & (g779) & (!g786) & (g785) & (g780)) + ((!g775) & (g776) & (g779) & (g786) & (!g785) & (!g780)) + ((!g775) & (g776) & (g779) & (g786) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g786) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g786) & (g785) & (g780)) + ((g775) & (!g776) & (!g779) & (g786) & (!g785) & (g780)) + ((g775) & (!g776) & (!g779) & (g786) & (g785) & (g780)) + ((g775) & (!g776) & (g779) & (!g786) & (!g785) & (!g780)) + ((g775) & (!g776) & (g779) & (!g786) & (!g785) & (g780)) + ((g775) & (!g776) & (g779) & (!g786) & (g785) & (g780)) + ((g775) & (!g776) & (g779) & (g786) & (!g785) & (!g780)) + ((g775) & (!g776) & (g779) & (g786) & (!g785) & (g780)) + ((g775) & (!g776) & (g779) & (g786) & (g785) & (!g780)) + ((g775) & (!g776) & (g779) & (g786) & (g785) & (g780)) + ((g775) & (g776) & (!g779) & (!g786) & (!g785) & (g780)) + ((g775) & (g776) & (!g779) & (g786) & (!g785) & (!g780)) + ((g775) & (g776) & (!g779) & (g786) & (g785) & (!g780)) + ((g775) & (g776) & (g779) & (!g786) & (!g785) & (!g780)) + ((g775) & (g776) & (g779) & (!g786) & (!g785) & (g780)) + ((g775) & (g776) & (g779) & (!g786) & (g785) & (!g780)) + ((g775) & (g776) & (g779) & (g786) & (!g785) & (!g780)) + ((g775) & (g776) & (g779) & (g786) & (g785) & (!g780)));
	assign g814 = (((!g775) & (!g776) & (!g779) & (!g786) & (g785) & (g780)) + ((!g775) & (!g776) & (!g779) & (g786) & (!g785) & (!g780)) + ((!g775) & (!g776) & (!g779) & (g786) & (g785) & (g780)) + ((!g775) & (!g776) & (g779) & (!g786) & (!g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (!g786) & (g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (g786) & (!g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (g786) & (!g785) & (g780)) + ((!g775) & (!g776) & (g779) & (g786) & (g785) & (!g780)) + ((!g775) & (g776) & (!g779) & (!g786) & (!g785) & (!g780)) + ((!g775) & (g776) & (!g779) & (g786) & (!g785) & (g780)) + ((!g775) & (g776) & (!g779) & (g786) & (g785) & (!g780)) + ((!g775) & (g776) & (!g779) & (g786) & (g785) & (g780)) + ((!g775) & (g776) & (g779) & (!g786) & (!g785) & (!g780)) + ((!g775) & (g776) & (g779) & (g786) & (!g785) & (!g780)) + ((!g775) & (g776) & (g779) & (g786) & (!g785) & (g780)) + ((g775) & (!g776) & (!g779) & (!g786) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g786) & (g785) & (g780)) + ((g775) & (!g776) & (g779) & (!g786) & (!g785) & (!g780)) + ((g775) & (!g776) & (g779) & (!g786) & (g785) & (!g780)) + ((g775) & (!g776) & (g779) & (g786) & (g785) & (!g780)) + ((g775) & (g776) & (!g779) & (!g786) & (g785) & (!g780)) + ((g775) & (g776) & (!g779) & (g786) & (g785) & (g780)) + ((g775) & (g776) & (g779) & (!g786) & (!g785) & (!g780)) + ((g775) & (g776) & (g779) & (!g786) & (!g785) & (g780)) + ((g775) & (g776) & (g779) & (!g786) & (g785) & (!g780)) + ((g775) & (g776) & (g779) & (g786) & (!g785) & (!g780)));
	assign g815 = (((!g811) & (!g812) & (!g813) & (!g814) & (g777) & (g778)) + ((!g811) & (!g812) & (g813) & (!g814) & (!g777) & (g778)) + ((!g811) & (!g812) & (g813) & (!g814) & (g777) & (g778)) + ((!g811) & (!g812) & (g813) & (g814) & (!g777) & (g778)) + ((!g811) & (g812) & (!g813) & (!g814) & (g777) & (!g778)) + ((!g811) & (g812) & (!g813) & (!g814) & (g777) & (g778)) + ((!g811) & (g812) & (!g813) & (g814) & (g777) & (!g778)) + ((!g811) & (g812) & (g813) & (!g814) & (!g777) & (g778)) + ((!g811) & (g812) & (g813) & (!g814) & (g777) & (!g778)) + ((!g811) & (g812) & (g813) & (!g814) & (g777) & (g778)) + ((!g811) & (g812) & (g813) & (g814) & (!g777) & (g778)) + ((!g811) & (g812) & (g813) & (g814) & (g777) & (!g778)) + ((g811) & (!g812) & (!g813) & (!g814) & (!g777) & (!g778)) + ((g811) & (!g812) & (!g813) & (!g814) & (g777) & (g778)) + ((g811) & (!g812) & (!g813) & (g814) & (!g777) & (!g778)) + ((g811) & (!g812) & (g813) & (!g814) & (!g777) & (!g778)) + ((g811) & (!g812) & (g813) & (!g814) & (!g777) & (g778)) + ((g811) & (!g812) & (g813) & (!g814) & (g777) & (g778)) + ((g811) & (!g812) & (g813) & (g814) & (!g777) & (!g778)) + ((g811) & (!g812) & (g813) & (g814) & (!g777) & (g778)) + ((g811) & (g812) & (!g813) & (!g814) & (!g777) & (!g778)) + ((g811) & (g812) & (!g813) & (!g814) & (g777) & (!g778)) + ((g811) & (g812) & (!g813) & (!g814) & (g777) & (g778)) + ((g811) & (g812) & (!g813) & (g814) & (!g777) & (!g778)) + ((g811) & (g812) & (!g813) & (g814) & (g777) & (!g778)) + ((g811) & (g812) & (g813) & (!g814) & (!g777) & (!g778)) + ((g811) & (g812) & (g813) & (!g814) & (!g777) & (g778)) + ((g811) & (g812) & (g813) & (!g814) & (g777) & (!g778)) + ((g811) & (g812) & (g813) & (!g814) & (g777) & (g778)) + ((g811) & (g812) & (g813) & (g814) & (!g777) & (!g778)) + ((g811) & (g812) & (g813) & (g814) & (!g777) & (g778)) + ((g811) & (g812) & (g813) & (g814) & (g777) & (!g778)));
	assign g817 = (((!g815) & (sk[126]) & (g816)) + ((g815) & (!sk[126]) & (!g816)) + ((g815) & (!sk[126]) & (g816)) + ((g815) & (sk[126]) & (!g816)));
	assign g818 = (((!g775) & (!g776) & (!g779) & (!g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (!g779) & (!g778) & (g785) & (g780)) + ((!g775) & (!g776) & (!g779) & (g778) & (g785) & (g780)) + ((!g775) & (!g776) & (g779) & (!g778) & (!g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (!g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (g779) & (!g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (!g778) & (g785) & (g780)) + ((!g775) & (!g776) & (g779) & (g778) & (!g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (g778) & (!g785) & (g780)) + ((!g775) & (g776) & (!g779) & (!g778) & (!g785) & (g780)) + ((!g775) & (g776) & (!g779) & (!g778) & (g785) & (!g780)) + ((!g775) & (g776) & (!g779) & (g778) & (g785) & (g780)) + ((!g775) & (g776) & (g779) & (!g778) & (g785) & (!g780)) + ((!g775) & (g776) & (g779) & (!g778) & (g785) & (g780)) + ((!g775) & (g776) & (g779) & (g778) & (!g785) & (!g780)) + ((!g775) & (g776) & (g779) & (g778) & (!g785) & (g780)) + ((!g775) & (g776) & (g779) & (g778) & (g785) & (g780)) + ((g775) & (!g776) & (!g779) & (!g778) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g778) & (g785) & (g780)) + ((g775) & (!g776) & (!g779) & (g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (g778) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (g778) & (g785) & (g780)) + ((g775) & (!g776) & (g779) & (!g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (g779) & (!g778) & (g785) & (!g780)) + ((g775) & (!g776) & (g779) & (g778) & (g785) & (!g780)) + ((g775) & (g776) & (!g779) & (!g778) & (g785) & (g780)) + ((g775) & (g776) & (g779) & (!g778) & (!g785) & (!g780)) + ((g775) & (g776) & (g779) & (!g778) & (g785) & (g780)));
	assign g819 = (((!g775) & (!g776) & (!g779) & (!g778) & (!g785) & (!g780)) + ((!g775) & (!g776) & (!g779) & (g778) & (!g785) & (!g780)) + ((!g775) & (!g776) & (!g779) & (g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (!g779) & (g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (!g778) & (g785) & (g780)) + ((!g775) & (!g776) & (g779) & (g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (g779) & (g778) & (g785) & (g780)) + ((!g775) & (g776) & (!g779) & (!g778) & (!g785) & (!g780)) + ((!g775) & (g776) & (!g779) & (!g778) & (g785) & (!g780)) + ((!g775) & (g776) & (g779) & (!g778) & (!g785) & (g780)) + ((!g775) & (g776) & (g779) & (!g778) & (g785) & (g780)) + ((!g775) & (g776) & (g779) & (g778) & (!g785) & (g780)) + ((!g775) & (g776) & (g779) & (g778) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g778) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g778) & (g785) & (g780)) + ((g775) & (!g776) & (!g779) & (g778) & (!g785) & (g780)) + ((g775) & (!g776) & (!g779) & (g778) & (g785) & (g780)) + ((g775) & (!g776) & (g779) & (g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (g779) & (g778) & (!g785) & (g780)) + ((g775) & (!g776) & (g779) & (g778) & (g785) & (g780)) + ((g775) & (g776) & (!g779) & (!g778) & (!g785) & (g780)) + ((g775) & (g776) & (!g779) & (!g778) & (g785) & (!g780)) + ((g775) & (g776) & (!g779) & (g778) & (g785) & (!g780)) + ((g775) & (g776) & (g779) & (!g778) & (!g785) & (g780)) + ((g775) & (g776) & (g779) & (!g778) & (g785) & (g780)) + ((g775) & (g776) & (g779) & (g778) & (!g785) & (!g780)) + ((g775) & (g776) & (g779) & (g778) & (g785) & (g780)));
	assign g820 = (((!g775) & (!g776) & (!g779) & (!g778) & (g785) & (g780)) + ((!g775) & (!g776) & (!g779) & (g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (!g778) & (!g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (!g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (g779) & (!g778) & (g785) & (g780)) + ((!g775) & (!g776) & (g779) & (g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (g779) & (g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (g779) & (g778) & (g785) & (g780)) + ((!g775) & (g776) & (!g779) & (!g778) & (g785) & (!g780)) + ((!g775) & (g776) & (!g779) & (!g778) & (g785) & (g780)) + ((!g775) & (g776) & (g779) & (!g778) & (!g785) & (!g780)) + ((!g775) & (g776) & (g779) & (g778) & (!g785) & (g780)) + ((!g775) & (g776) & (g779) & (g778) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g778) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (!g778) & (g785) & (g780)) + ((g775) & (!g776) & (!g779) & (g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (g778) & (!g785) & (g780)) + ((g775) & (!g776) & (g779) & (!g778) & (!g785) & (g780)) + ((g775) & (!g776) & (g779) & (!g778) & (g785) & (g780)) + ((g775) & (!g776) & (g779) & (g778) & (g785) & (!g780)) + ((g775) & (g776) & (!g779) & (!g778) & (!g785) & (!g780)) + ((g775) & (g776) & (!g779) & (!g778) & (!g785) & (g780)) + ((g775) & (g776) & (!g779) & (!g778) & (g785) & (g780)) + ((g775) & (g776) & (!g779) & (g778) & (!g785) & (g780)) + ((g775) & (g776) & (!g779) & (g778) & (g785) & (!g780)) + ((g775) & (g776) & (g779) & (!g778) & (!g785) & (g780)) + ((g775) & (g776) & (g779) & (!g778) & (g785) & (!g780)) + ((g775) & (g776) & (g779) & (g778) & (!g785) & (!g780)) + ((g775) & (g776) & (g779) & (g778) & (g785) & (!g780)) + ((g775) & (g776) & (g779) & (g778) & (g785) & (g780)));
	assign g821 = (((!g775) & (!g776) & (!g779) & (!g778) & (g785) & (!g780)) + ((!g775) & (!g776) & (!g779) & (g778) & (!g785) & (!g780)) + ((!g775) & (!g776) & (!g779) & (g778) & (g785) & (g780)) + ((!g775) & (!g776) & (g779) & (!g778) & (!g785) & (g780)) + ((!g775) & (!g776) & (g779) & (!g778) & (g785) & (g780)) + ((!g775) & (!g776) & (g779) & (g778) & (g785) & (g780)) + ((!g775) & (g776) & (!g779) & (!g778) & (!g785) & (g780)) + ((!g775) & (g776) & (!g779) & (g778) & (!g785) & (g780)) + ((!g775) & (g776) & (!g779) & (g778) & (g785) & (g780)) + ((!g775) & (g776) & (g779) & (!g778) & (!g785) & (!g780)) + ((!g775) & (g776) & (g779) & (!g778) & (g785) & (!g780)) + ((!g775) & (g776) & (g779) & (g778) & (!g785) & (g780)) + ((!g775) & (g776) & (g779) & (g778) & (g785) & (g780)) + ((g775) & (!g776) & (!g779) & (!g778) & (g785) & (!g780)) + ((g775) & (!g776) & (!g779) & (g778) & (g785) & (g780)) + ((g775) & (!g776) & (g779) & (!g778) & (!g785) & (!g780)) + ((g775) & (!g776) & (g779) & (!g778) & (g785) & (g780)) + ((g775) & (!g776) & (g779) & (g778) & (!g785) & (!g780)) + ((g775) & (g776) & (!g779) & (!g778) & (g785) & (g780)) + ((g775) & (g776) & (!g779) & (g778) & (!g785) & (!g780)) + ((g775) & (g776) & (!g779) & (g778) & (!g785) & (g780)) + ((g775) & (g776) & (g779) & (!g778) & (g785) & (g780)));
	assign g822 = (((!g818) & (!g819) & (!g820) & (!g821) & (!g786) & (!g777)) + ((!g818) & (!g819) & (!g820) & (!g821) & (!g786) & (g777)) + ((!g818) & (!g819) & (!g820) & (!g821) & (g786) & (!g777)) + ((!g818) & (!g819) & (!g820) & (g821) & (!g786) & (!g777)) + ((!g818) & (!g819) & (!g820) & (g821) & (!g786) & (g777)) + ((!g818) & (!g819) & (!g820) & (g821) & (g786) & (!g777)) + ((!g818) & (!g819) & (!g820) & (g821) & (g786) & (g777)) + ((!g818) & (!g819) & (g820) & (!g821) & (!g786) & (!g777)) + ((!g818) & (!g819) & (g820) & (!g821) & (g786) & (!g777)) + ((!g818) & (!g819) & (g820) & (g821) & (!g786) & (!g777)) + ((!g818) & (!g819) & (g820) & (g821) & (g786) & (!g777)) + ((!g818) & (!g819) & (g820) & (g821) & (g786) & (g777)) + ((!g818) & (g819) & (!g820) & (!g821) & (!g786) & (!g777)) + ((!g818) & (g819) & (!g820) & (!g821) & (!g786) & (g777)) + ((!g818) & (g819) & (!g820) & (g821) & (!g786) & (!g777)) + ((!g818) & (g819) & (!g820) & (g821) & (!g786) & (g777)) + ((!g818) & (g819) & (!g820) & (g821) & (g786) & (g777)) + ((!g818) & (g819) & (g820) & (!g821) & (!g786) & (!g777)) + ((!g818) & (g819) & (g820) & (g821) & (!g786) & (!g777)) + ((!g818) & (g819) & (g820) & (g821) & (g786) & (g777)) + ((g818) & (!g819) & (!g820) & (!g821) & (!g786) & (g777)) + ((g818) & (!g819) & (!g820) & (!g821) & (g786) & (!g777)) + ((g818) & (!g819) & (!g820) & (g821) & (!g786) & (g777)) + ((g818) & (!g819) & (!g820) & (g821) & (g786) & (!g777)) + ((g818) & (!g819) & (!g820) & (g821) & (g786) & (g777)) + ((g818) & (!g819) & (g820) & (!g821) & (g786) & (!g777)) + ((g818) & (!g819) & (g820) & (g821) & (g786) & (!g777)) + ((g818) & (!g819) & (g820) & (g821) & (g786) & (g777)) + ((g818) & (g819) & (!g820) & (!g821) & (!g786) & (g777)) + ((g818) & (g819) & (!g820) & (g821) & (!g786) & (g777)) + ((g818) & (g819) & (!g820) & (g821) & (g786) & (g777)) + ((g818) & (g819) & (g820) & (g821) & (g786) & (g777)));
	assign g824 = (((!sk[4]) & (g822) & (!g823)) + ((!sk[4]) & (g822) & (g823)) + ((sk[4]) & (!g822) & (g823)) + ((sk[4]) & (g822) & (!g823)));
	assign g825 = (((!g775) & (!g786) & (!g777) & (!g778) & (!g785) & (g780)) + ((!g775) & (!g786) & (!g777) & (!g778) & (g785) & (g780)) + ((!g775) & (!g786) & (!g777) & (g778) & (!g785) & (!g780)) + ((!g775) & (!g786) & (!g777) & (g778) & (!g785) & (g780)) + ((!g775) & (!g786) & (!g777) & (g778) & (g785) & (!g780)) + ((!g775) & (!g786) & (!g777) & (g778) & (g785) & (g780)) + ((!g775) & (!g786) & (g777) & (!g778) & (!g785) & (g780)) + ((!g775) & (!g786) & (g777) & (!g778) & (g785) & (g780)) + ((!g775) & (!g786) & (g777) & (g778) & (g785) & (!g780)) + ((!g775) & (g786) & (g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (g786) & (g777) & (!g778) & (g785) & (g780)) + ((!g775) & (g786) & (g777) & (g778) & (!g785) & (g780)) + ((g775) & (!g786) & (!g777) & (!g778) & (g785) & (!g780)) + ((g775) & (!g786) & (!g777) & (g778) & (!g785) & (!g780)) + ((g775) & (!g786) & (!g777) & (g778) & (!g785) & (g780)) + ((g775) & (!g786) & (!g777) & (g778) & (g785) & (g780)) + ((g775) & (!g786) & (g777) & (!g778) & (!g785) & (g780)) + ((g775) & (!g786) & (g777) & (!g778) & (g785) & (g780)) + ((g775) & (!g786) & (g777) & (g778) & (g785) & (!g780)) + ((g775) & (!g786) & (g777) & (g778) & (g785) & (g780)) + ((g775) & (g786) & (!g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (g786) & (!g777) & (!g778) & (!g785) & (g780)) + ((g775) & (g786) & (!g777) & (!g778) & (g785) & (!g780)) + ((g775) & (g786) & (!g777) & (g778) & (!g785) & (!g780)) + ((g775) & (g786) & (g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (g786) & (g777) & (!g778) & (!g785) & (g780)) + ((g775) & (g786) & (g777) & (!g778) & (g785) & (!g780)) + ((g775) & (g786) & (g777) & (g778) & (!g785) & (g780)));
	assign g826 = (((!g775) & (!g786) & (!g777) & (!g778) & (!g785) & (!g780)) + ((!g775) & (!g786) & (!g777) & (g778) & (g785) & (g780)) + ((!g775) & (!g786) & (g777) & (!g778) & (!g785) & (!g780)) + ((!g775) & (!g786) & (g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (!g786) & (g777) & (!g778) & (g785) & (g780)) + ((!g775) & (!g786) & (g777) & (g778) & (!g785) & (!g780)) + ((!g775) & (!g786) & (g777) & (g778) & (g785) & (g780)) + ((!g775) & (g786) & (!g777) & (!g778) & (!g785) & (!g780)) + ((!g775) & (g786) & (!g777) & (!g778) & (g785) & (g780)) + ((!g775) & (g786) & (!g777) & (g778) & (!g785) & (g780)) + ((!g775) & (g786) & (g777) & (!g778) & (!g785) & (!g780)) + ((!g775) & (g786) & (g777) & (!g778) & (g785) & (g780)) + ((!g775) & (g786) & (g777) & (g778) & (g785) & (!g780)) + ((!g775) & (g786) & (g777) & (g778) & (g785) & (g780)) + ((g775) & (!g786) & (!g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (!g786) & (!g777) & (!g778) & (g785) & (g780)) + ((g775) & (!g786) & (!g777) & (g778) & (!g785) & (!g780)) + ((g775) & (!g786) & (!g777) & (g778) & (g785) & (g780)) + ((g775) & (!g786) & (g777) & (!g778) & (g785) & (g780)) + ((g775) & (!g786) & (g777) & (g778) & (!g785) & (g780)) + ((g775) & (g786) & (!g777) & (!g778) & (g785) & (!g780)) + ((g775) & (g786) & (!g777) & (!g778) & (g785) & (g780)) + ((g775) & (g786) & (!g777) & (g778) & (!g785) & (g780)) + ((g775) & (g786) & (!g777) & (g778) & (g785) & (!g780)) + ((g775) & (g786) & (!g777) & (g778) & (g785) & (g780)) + ((g775) & (g786) & (g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (g786) & (g777) & (!g778) & (g785) & (!g780)) + ((g775) & (g786) & (g777) & (g778) & (!g785) & (!g780)));
	assign g827 = (((!g775) & (!g786) & (!g777) & (!g778) & (!g785) & (g780)) + ((!g775) & (!g786) & (!g777) & (!g778) & (g785) & (g780)) + ((!g775) & (!g786) & (!g777) & (g778) & (g785) & (!g780)) + ((!g775) & (!g786) & (!g777) & (g778) & (g785) & (g780)) + ((!g775) & (!g786) & (g777) & (!g778) & (g785) & (g780)) + ((!g775) & (!g786) & (g777) & (g778) & (!g785) & (!g780)) + ((!g775) & (!g786) & (g777) & (g778) & (!g785) & (g780)) + ((!g775) & (!g786) & (g777) & (g778) & (g785) & (g780)) + ((!g775) & (g786) & (!g777) & (!g778) & (!g785) & (!g780)) + ((!g775) & (g786) & (!g777) & (!g778) & (!g785) & (g780)) + ((!g775) & (g786) & (!g777) & (!g778) & (g785) & (g780)) + ((!g775) & (g786) & (!g777) & (g778) & (!g785) & (g780)) + ((!g775) & (g786) & (!g777) & (g778) & (g785) & (!g780)) + ((!g775) & (g786) & (g777) & (!g778) & (!g785) & (g780)) + ((!g775) & (g786) & (g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (g786) & (g777) & (g778) & (!g785) & (!g780)) + ((!g775) & (g786) & (g777) & (g778) & (g785) & (!g780)) + ((!g775) & (g786) & (g777) & (g778) & (g785) & (g780)) + ((g775) & (!g786) & (!g777) & (!g778) & (!g785) & (g780)) + ((g775) & (!g786) & (!g777) & (g778) & (!g785) & (!g780)) + ((g775) & (!g786) & (!g777) & (g778) & (g785) & (!g780)) + ((g775) & (!g786) & (g777) & (!g778) & (g785) & (g780)) + ((g775) & (!g786) & (g777) & (g778) & (!g785) & (g780)) + ((g775) & (g786) & (!g777) & (!g778) & (!g785) & (g780)) + ((g775) & (g786) & (!g777) & (g778) & (!g785) & (!g780)) + ((g775) & (g786) & (!g777) & (g778) & (g785) & (!g780)) + ((g775) & (g786) & (g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (g786) & (g777) & (!g778) & (g785) & (!g780)) + ((g775) & (g786) & (g777) & (!g778) & (g785) & (g780)) + ((g775) & (g786) & (g777) & (g778) & (g785) & (g780)));
	assign g828 = (((!g775) & (!g786) & (!g777) & (!g778) & (g785) & (g780)) + ((!g775) & (!g786) & (!g777) & (g778) & (!g785) & (!g780)) + ((!g775) & (!g786) & (!g777) & (g778) & (g785) & (g780)) + ((!g775) & (!g786) & (g777) & (!g778) & (!g785) & (!g780)) + ((!g775) & (!g786) & (g777) & (g778) & (g785) & (!g780)) + ((!g775) & (!g786) & (g777) & (g778) & (g785) & (g780)) + ((!g775) & (g786) & (!g777) & (g778) & (!g785) & (!g780)) + ((!g775) & (g786) & (!g777) & (g778) & (g785) & (!g780)) + ((!g775) & (g786) & (g777) & (!g778) & (g785) & (!g780)) + ((!g775) & (g786) & (g777) & (!g778) & (g785) & (g780)) + ((g775) & (!g786) & (!g777) & (!g778) & (!g785) & (g780)) + ((g775) & (!g786) & (!g777) & (!g778) & (g785) & (!g780)) + ((g775) & (!g786) & (!g777) & (g778) & (!g785) & (g780)) + ((g775) & (!g786) & (g777) & (!g778) & (g785) & (!g780)) + ((g775) & (!g786) & (g777) & (!g778) & (g785) & (g780)) + ((g775) & (!g786) & (g777) & (g778) & (g785) & (!g780)) + ((g775) & (!g786) & (g777) & (g778) & (g785) & (g780)) + ((g775) & (g786) & (!g777) & (!g778) & (g785) & (!g780)) + ((g775) & (g786) & (!g777) & (g778) & (!g785) & (g780)) + ((g775) & (g786) & (g777) & (!g778) & (!g785) & (!g780)) + ((g775) & (g786) & (g777) & (!g778) & (g785) & (g780)) + ((g775) & (g786) & (g777) & (g778) & (!g785) & (g780)));
	assign g829 = (((!g825) & (!g826) & (!g827) & (!g828) & (!g779) & (!g776)) + ((!g825) & (!g826) & (!g827) & (!g828) & (!g779) & (g776)) + ((!g825) & (!g826) & (!g827) & (!g828) & (g779) & (!g776)) + ((!g825) & (!g826) & (!g827) & (g828) & (!g779) & (!g776)) + ((!g825) & (!g826) & (!g827) & (g828) & (!g779) & (g776)) + ((!g825) & (!g826) & (!g827) & (g828) & (g779) & (!g776)) + ((!g825) & (!g826) & (!g827) & (g828) & (g779) & (g776)) + ((!g825) & (!g826) & (g827) & (!g828) & (!g779) & (!g776)) + ((!g825) & (!g826) & (g827) & (!g828) & (g779) & (!g776)) + ((!g825) & (!g826) & (g827) & (g828) & (!g779) & (!g776)) + ((!g825) & (!g826) & (g827) & (g828) & (g779) & (!g776)) + ((!g825) & (!g826) & (g827) & (g828) & (g779) & (g776)) + ((!g825) & (g826) & (!g827) & (!g828) & (!g779) & (!g776)) + ((!g825) & (g826) & (!g827) & (!g828) & (!g779) & (g776)) + ((!g825) & (g826) & (!g827) & (g828) & (!g779) & (!g776)) + ((!g825) & (g826) & (!g827) & (g828) & (!g779) & (g776)) + ((!g825) & (g826) & (!g827) & (g828) & (g779) & (g776)) + ((!g825) & (g826) & (g827) & (!g828) & (!g779) & (!g776)) + ((!g825) & (g826) & (g827) & (g828) & (!g779) & (!g776)) + ((!g825) & (g826) & (g827) & (g828) & (g779) & (g776)) + ((g825) & (!g826) & (!g827) & (!g828) & (!g779) & (g776)) + ((g825) & (!g826) & (!g827) & (!g828) & (g779) & (!g776)) + ((g825) & (!g826) & (!g827) & (g828) & (!g779) & (g776)) + ((g825) & (!g826) & (!g827) & (g828) & (g779) & (!g776)) + ((g825) & (!g826) & (!g827) & (g828) & (g779) & (g776)) + ((g825) & (!g826) & (g827) & (!g828) & (g779) & (!g776)) + ((g825) & (!g826) & (g827) & (g828) & (g779) & (!g776)) + ((g825) & (!g826) & (g827) & (g828) & (g779) & (g776)) + ((g825) & (g826) & (!g827) & (!g828) & (!g779) & (g776)) + ((g825) & (g826) & (!g827) & (g828) & (!g779) & (g776)) + ((g825) & (g826) & (!g827) & (g828) & (g779) & (g776)) + ((g825) & (g826) & (g827) & (g828) & (g779) & (g776)));
	assign g831 = (((!g829) & (sk[10]) & (g830)) + ((g829) & (!sk[10]) & (!g830)) + ((g829) & (!sk[10]) & (g830)) + ((g829) & (sk[10]) & (!g830)));
	assign g832 = (((!g779) & (!g776) & (!g777) & (!g778) & (!g785) & (g786)) + ((!g779) & (!g776) & (!g777) & (!g778) & (g785) & (!g786)) + ((!g779) & (!g776) & (!g777) & (g778) & (!g785) & (g786)) + ((!g779) & (!g776) & (!g777) & (g778) & (g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (!g778) & (!g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (!g778) & (g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (g778) & (!g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (g778) & (g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (g778) & (g785) & (g786)) + ((!g779) & (g776) & (!g777) & (!g778) & (g785) & (!g786)) + ((!g779) & (g776) & (!g777) & (g778) & (g785) & (!g786)) + ((!g779) & (g776) & (!g777) & (g778) & (g785) & (g786)) + ((!g779) & (g776) & (g777) & (!g778) & (g785) & (g786)) + ((!g779) & (g776) & (g777) & (g778) & (!g785) & (!g786)) + ((g779) & (!g776) & (!g777) & (!g778) & (!g785) & (g786)) + ((g779) & (!g776) & (!g777) & (g778) & (!g785) & (g786)) + ((g779) & (!g776) & (g777) & (g778) & (g785) & (g786)) + ((g779) & (g776) & (!g777) & (!g778) & (g785) & (g786)) + ((g779) & (g776) & (!g777) & (g778) & (!g785) & (!g786)) + ((g779) & (g776) & (!g777) & (g778) & (g785) & (!g786)) + ((g779) & (g776) & (g777) & (!g778) & (!g785) & (g786)) + ((g779) & (g776) & (g777) & (!g778) & (g785) & (!g786)) + ((g779) & (g776) & (g777) & (!g778) & (g785) & (g786)) + ((g779) & (g776) & (g777) & (g778) & (!g785) & (g786)));
	assign g833 = (((!g779) & (!g776) & (!g777) & (!g778) & (!g785) & (!g786)) + ((!g779) & (!g776) & (!g777) & (!g778) & (!g785) & (g786)) + ((!g779) & (!g776) & (!g777) & (g778) & (!g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (!g778) & (!g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (!g778) & (g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (!g778) & (g785) & (g786)) + ((!g779) & (!g776) & (g777) & (g778) & (!g785) & (g786)) + ((!g779) & (!g776) & (g777) & (g778) & (g785) & (g786)) + ((!g779) & (g776) & (!g777) & (!g778) & (!g785) & (!g786)) + ((!g779) & (g776) & (!g777) & (!g778) & (g785) & (!g786)) + ((!g779) & (g776) & (!g777) & (g778) & (!g785) & (!g786)) + ((!g779) & (g776) & (!g777) & (g778) & (!g785) & (g786)) + ((!g779) & (g776) & (!g777) & (g778) & (g785) & (g786)) + ((!g779) & (g776) & (g777) & (!g778) & (!g785) & (g786)) + ((!g779) & (g776) & (g777) & (g778) & (!g785) & (!g786)) + ((!g779) & (g776) & (g777) & (g778) & (!g785) & (g786)) + ((g779) & (!g776) & (!g777) & (!g778) & (!g785) & (g786)) + ((g779) & (!g776) & (!g777) & (!g778) & (g785) & (g786)) + ((g779) & (!g776) & (!g777) & (g778) & (!g785) & (!g786)) + ((g779) & (!g776) & (!g777) & (g778) & (g785) & (g786)) + ((g779) & (!g776) & (g777) & (!g778) & (!g785) & (!g786)) + ((g779) & (!g776) & (g777) & (!g778) & (g785) & (g786)) + ((g779) & (!g776) & (g777) & (g778) & (g785) & (!g786)) + ((g779) & (g776) & (!g777) & (!g778) & (!g785) & (!g786)) + ((g779) & (g776) & (!g777) & (!g778) & (!g785) & (g786)) + ((g779) & (g776) & (!g777) & (!g778) & (g785) & (g786)) + ((g779) & (g776) & (!g777) & (g778) & (!g785) & (g786)) + ((g779) & (g776) & (!g777) & (g778) & (g785) & (!g786)) + ((g779) & (g776) & (g777) & (!g778) & (g785) & (!g786)) + ((g779) & (g776) & (g777) & (!g778) & (g785) & (g786)));
	assign g834 = (((!g779) & (!g776) & (!g777) & (!g778) & (g785) & (!g786)) + ((!g779) & (!g776) & (!g777) & (g778) & (!g785) & (!g786)) + ((!g779) & (!g776) & (!g777) & (g778) & (g785) & (!g786)) + ((!g779) & (!g776) & (!g777) & (g778) & (g785) & (g786)) + ((!g779) & (!g776) & (g777) & (!g778) & (!g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (!g778) & (!g785) & (g786)) + ((!g779) & (!g776) & (g777) & (!g778) & (g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (g778) & (!g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (g778) & (g785) & (g786)) + ((!g779) & (g776) & (!g777) & (!g778) & (!g785) & (g786)) + ((!g779) & (g776) & (!g777) & (!g778) & (g785) & (!g786)) + ((!g779) & (g776) & (!g777) & (!g778) & (g785) & (g786)) + ((!g779) & (g776) & (g777) & (!g778) & (!g785) & (g786)) + ((!g779) & (g776) & (g777) & (!g778) & (g785) & (!g786)) + ((!g779) & (g776) & (g777) & (!g778) & (g785) & (g786)) + ((!g779) & (g776) & (g777) & (g778) & (!g785) & (!g786)) + ((g779) & (!g776) & (!g777) & (!g778) & (g785) & (!g786)) + ((g779) & (!g776) & (!g777) & (g778) & (!g785) & (!g786)) + ((g779) & (!g776) & (!g777) & (g778) & (g785) & (g786)) + ((g779) & (!g776) & (g777) & (!g778) & (!g785) & (!g786)) + ((g779) & (!g776) & (g777) & (!g778) & (!g785) & (g786)) + ((g779) & (!g776) & (g777) & (g778) & (!g785) & (!g786)) + ((g779) & (!g776) & (g777) & (g778) & (g785) & (!g786)) + ((g779) & (g776) & (!g777) & (!g778) & (g785) & (!g786)) + ((g779) & (g776) & (!g777) & (g778) & (!g785) & (!g786)) + ((g779) & (g776) & (!g777) & (g778) & (g785) & (g786)) + ((g779) & (g776) & (g777) & (!g778) & (!g785) & (!g786)) + ((g779) & (g776) & (g777) & (!g778) & (g785) & (!g786)) + ((g779) & (g776) & (g777) & (!g778) & (g785) & (g786)) + ((g779) & (g776) & (g777) & (g778) & (!g785) & (g786)));
	assign g835 = (((!g779) & (!g776) & (!g777) & (!g778) & (!g785) & (g786)) + ((!g779) & (!g776) & (!g777) & (g778) & (g785) & (!g786)) + ((!g779) & (!g776) & (!g777) & (g778) & (g785) & (g786)) + ((!g779) & (!g776) & (g777) & (!g778) & (!g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (!g778) & (!g785) & (g786)) + ((!g779) & (!g776) & (g777) & (g778) & (g785) & (!g786)) + ((!g779) & (!g776) & (g777) & (g778) & (g785) & (g786)) + ((!g779) & (g776) & (!g777) & (!g778) & (!g785) & (!g786)) + ((!g779) & (g776) & (!g777) & (!g778) & (!g785) & (g786)) + ((!g779) & (g776) & (!g777) & (!g778) & (g785) & (g786)) + ((!g779) & (g776) & (!g777) & (g778) & (!g785) & (g786)) + ((!g779) & (g776) & (g777) & (!g778) & (!g785) & (g786)) + ((!g779) & (g776) & (g777) & (g778) & (!g785) & (!g786)) + ((!g779) & (g776) & (g777) & (g778) & (!g785) & (g786)) + ((!g779) & (g776) & (g777) & (g778) & (g785) & (!g786)) + ((!g779) & (g776) & (g777) & (g778) & (g785) & (g786)) + ((g779) & (!g776) & (!g777) & (g778) & (!g785) & (g786)) + ((g779) & (!g776) & (g777) & (!g778) & (!g785) & (!g786)) + ((g779) & (!g776) & (g777) & (g778) & (!g785) & (!g786)) + ((g779) & (!g776) & (g777) & (g778) & (!g785) & (g786)) + ((g779) & (!g776) & (g777) & (g778) & (g785) & (g786)) + ((g779) & (g776) & (!g777) & (!g778) & (!g785) & (g786)) + ((g779) & (g776) & (!g777) & (!g778) & (g785) & (g786)) + ((g779) & (g776) & (!g777) & (g778) & (!g785) & (!g786)) + ((g779) & (g776) & (!g777) & (g778) & (g785) & (!g786)) + ((g779) & (g776) & (!g777) & (g778) & (g785) & (g786)) + ((g779) & (g776) & (g777) & (!g778) & (g785) & (g786)) + ((g779) & (g776) & (g777) & (g778) & (g785) & (g786)));
	assign g836 = (((!g832) & (!g833) & (!g834) & (!g835) & (!g775) & (g780)) + ((!g832) & (!g833) & (!g834) & (!g835) & (g775) & (!g780)) + ((!g832) & (!g833) & (!g834) & (!g835) & (g775) & (g780)) + ((!g832) & (!g833) & (!g834) & (g835) & (!g775) & (g780)) + ((!g832) & (!g833) & (!g834) & (g835) & (g775) & (!g780)) + ((!g832) & (!g833) & (g834) & (!g835) & (g775) & (!g780)) + ((!g832) & (!g833) & (g834) & (!g835) & (g775) & (g780)) + ((!g832) & (!g833) & (g834) & (g835) & (g775) & (!g780)) + ((!g832) & (g833) & (!g834) & (!g835) & (!g775) & (g780)) + ((!g832) & (g833) & (!g834) & (!g835) & (g775) & (g780)) + ((!g832) & (g833) & (!g834) & (g835) & (!g775) & (g780)) + ((!g832) & (g833) & (g834) & (!g835) & (g775) & (g780)) + ((g832) & (!g833) & (!g834) & (!g835) & (!g775) & (!g780)) + ((g832) & (!g833) & (!g834) & (!g835) & (!g775) & (g780)) + ((g832) & (!g833) & (!g834) & (!g835) & (g775) & (!g780)) + ((g832) & (!g833) & (!g834) & (!g835) & (g775) & (g780)) + ((g832) & (!g833) & (!g834) & (g835) & (!g775) & (!g780)) + ((g832) & (!g833) & (!g834) & (g835) & (!g775) & (g780)) + ((g832) & (!g833) & (!g834) & (g835) & (g775) & (!g780)) + ((g832) & (!g833) & (g834) & (!g835) & (!g775) & (!g780)) + ((g832) & (!g833) & (g834) & (!g835) & (g775) & (!g780)) + ((g832) & (!g833) & (g834) & (!g835) & (g775) & (g780)) + ((g832) & (!g833) & (g834) & (g835) & (!g775) & (!g780)) + ((g832) & (!g833) & (g834) & (g835) & (g775) & (!g780)) + ((g832) & (g833) & (!g834) & (!g835) & (!g775) & (!g780)) + ((g832) & (g833) & (!g834) & (!g835) & (!g775) & (g780)) + ((g832) & (g833) & (!g834) & (!g835) & (g775) & (g780)) + ((g832) & (g833) & (!g834) & (g835) & (!g775) & (!g780)) + ((g832) & (g833) & (!g834) & (g835) & (!g775) & (g780)) + ((g832) & (g833) & (g834) & (!g835) & (!g775) & (!g780)) + ((g832) & (g833) & (g834) & (!g835) & (g775) & (g780)) + ((g832) & (g833) & (g834) & (g835) & (!g775) & (!g780)));
	assign g838 = (((!g836) & (sk[16]) & (g837)) + ((g836) & (!sk[16]) & (!g837)) + ((g836) & (!sk[16]) & (g837)) + ((g836) & (sk[16]) & (!g837)));
	assign g845 = (((!g839) & (!g840) & (!g841) & (!g842) & (g843) & (g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g843) & (!g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g843) & (g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (g843) & (!g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (!g843) & (!g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (!g843) & (g844)) + ((!g839) & (!g840) & (g841) & (g842) & (!g843) & (!g844)) + ((!g839) & (!g840) & (g841) & (g842) & (g843) & (g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (g843) & (!g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (g843) & (g844)) + ((!g839) & (g840) & (!g841) & (g842) & (g843) & (!g844)) + ((!g839) & (g840) & (!g841) & (g842) & (g843) & (g844)) + ((!g839) & (g840) & (g841) & (!g842) & (g843) & (!g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (!g843) & (!g844)) + ((g839) & (!g840) & (g841) & (!g842) & (g843) & (!g844)) + ((g839) & (!g840) & (g841) & (g842) & (!g843) & (g844)) + ((g839) & (!g840) & (g841) & (g842) & (g843) & (g844)) + ((g839) & (g840) & (!g841) & (!g842) & (!g843) & (g844)) + ((g839) & (g840) & (!g841) & (!g842) & (g843) & (!g844)) + ((g839) & (g840) & (g841) & (!g842) & (!g843) & (g844)) + ((g839) & (g840) & (g841) & (!g842) & (g843) & (!g844)) + ((g839) & (g840) & (g841) & (g842) & (!g843) & (!g844)) + ((g839) & (g840) & (g841) & (g842) & (g843) & (!g844)) + ((g839) & (g840) & (g841) & (g842) & (g843) & (g844)));
	assign g846 = (((!g839) & (!g840) & (!g841) & (!g842) & (g843) & (!g844)) + ((!g839) & (!g840) & (!g841) & (!g842) & (g843) & (g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g843) & (!g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g843) & (g844)) + ((!g839) & (!g840) & (g841) & (g842) & (!g843) & (g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (!g843) & (!g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (!g843) & (g844)) + ((!g839) & (g840) & (g841) & (!g842) & (!g843) & (!g844)) + ((!g839) & (g840) & (g841) & (!g842) & (!g843) & (g844)) + ((!g839) & (g840) & (g841) & (!g842) & (g843) & (!g844)) + ((!g839) & (g840) & (g841) & (g842) & (g843) & (g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (!g843) & (g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (g843) & (!g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (g843) & (g844)) + ((g839) & (!g840) & (!g841) & (g842) & (g843) & (!g844)) + ((g839) & (!g840) & (g841) & (!g842) & (!g843) & (!g844)) + ((g839) & (!g840) & (g841) & (!g842) & (g843) & (g844)) + ((g839) & (!g840) & (g841) & (g842) & (!g843) & (g844)) + ((g839) & (!g840) & (g841) & (g842) & (g843) & (g844)) + ((g839) & (g840) & (!g841) & (!g842) & (!g843) & (!g844)) + ((g839) & (g840) & (!g841) & (!g842) & (!g843) & (g844)) + ((g839) & (g840) & (!g841) & (!g842) & (g843) & (!g844)) + ((g839) & (g840) & (!g841) & (!g842) & (g843) & (g844)) + ((g839) & (g840) & (!g841) & (g842) & (!g843) & (!g844)) + ((g839) & (g840) & (!g841) & (g842) & (g843) & (!g844)) + ((g839) & (g840) & (!g841) & (g842) & (g843) & (g844)) + ((g839) & (g840) & (g841) & (!g842) & (g843) & (!g844)) + ((g839) & (g840) & (g841) & (!g842) & (g843) & (g844)) + ((g839) & (g840) & (g841) & (g842) & (!g843) & (g844)) + ((g839) & (g840) & (g841) & (g842) & (g843) & (!g844)));
	assign g847 = (((!g839) & (!g840) & (!g841) & (!g842) & (!g843) & (!g844)) + ((!g839) & (!g840) & (!g841) & (!g842) & (g843) & (g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (g843) & (g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (!g843) & (!g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (!g843) & (g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (g843) & (g844)) + ((!g839) & (!g840) & (g841) & (g842) & (!g843) & (g844)) + ((!g839) & (!g840) & (g841) & (g842) & (g843) & (!g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (!g843) & (!g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (g843) & (!g844)) + ((!g839) & (g840) & (!g841) & (g842) & (g843) & (g844)) + ((!g839) & (g840) & (g841) & (g842) & (!g843) & (!g844)) + ((!g839) & (g840) & (g841) & (g842) & (g843) & (!g844)) + ((g839) & (!g840) & (!g841) & (g842) & (!g843) & (!g844)) + ((g839) & (!g840) & (!g841) & (g842) & (!g843) & (g844)) + ((g839) & (!g840) & (!g841) & (g842) & (g843) & (!g844)) + ((g839) & (!g840) & (g841) & (!g842) & (!g843) & (!g844)) + ((g839) & (!g840) & (g841) & (!g842) & (g843) & (g844)) + ((g839) & (!g840) & (g841) & (g842) & (!g843) & (!g844)) + ((g839) & (!g840) & (g841) & (g842) & (!g843) & (g844)) + ((g839) & (!g840) & (g841) & (g842) & (g843) & (!g844)) + ((g839) & (!g840) & (g841) & (g842) & (g843) & (g844)) + ((g839) & (g840) & (!g841) & (!g842) & (g843) & (g844)) + ((g839) & (g840) & (!g841) & (g842) & (!g843) & (!g844)) + ((g839) & (g840) & (!g841) & (g842) & (g843) & (!g844)) + ((g839) & (g840) & (!g841) & (g842) & (g843) & (g844)) + ((g839) & (g840) & (g841) & (!g842) & (!g843) & (!g844)) + ((g839) & (g840) & (g841) & (g842) & (!g843) & (!g844)) + ((g839) & (g840) & (g841) & (g842) & (!g843) & (g844)) + ((g839) & (g840) & (g841) & (g842) & (g843) & (g844)));
	assign g848 = (((!g839) & (!g840) & (!g841) & (!g842) & (!g843) & (g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (g843) & (!g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (g843) & (g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (!g843) & (g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (g843) & (g844)) + ((!g839) & (!g840) & (g841) & (g842) & (!g843) & (g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (!g843) & (!g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (!g843) & (g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (g843) & (!g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (g843) & (g844)) + ((!g839) & (g840) & (!g841) & (g842) & (g843) & (!g844)) + ((!g839) & (g840) & (!g841) & (g842) & (g843) & (g844)) + ((!g839) & (g840) & (g841) & (g842) & (!g843) & (!g844)) + ((!g839) & (g840) & (g841) & (g842) & (g843) & (!g844)) + ((!g839) & (g840) & (g841) & (g842) & (g843) & (g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (!g843) & (!g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (g843) & (g844)) + ((g839) & (!g840) & (!g841) & (g842) & (g843) & (!g844)) + ((g839) & (!g840) & (!g841) & (g842) & (g843) & (g844)) + ((g839) & (!g840) & (g841) & (!g842) & (!g843) & (g844)) + ((g839) & (!g840) & (g841) & (!g842) & (g843) & (!g844)) + ((g839) & (!g840) & (g841) & (g842) & (g843) & (!g844)) + ((g839) & (g840) & (!g841) & (!g842) & (!g843) & (g844)) + ((g839) & (g840) & (!g841) & (!g842) & (g843) & (g844)) + ((g839) & (g840) & (!g841) & (g842) & (g843) & (!g844)) + ((g839) & (g840) & (!g841) & (g842) & (g843) & (g844)) + ((g839) & (g840) & (g841) & (!g842) & (!g843) & (g844)) + ((g839) & (g840) & (g841) & (g842) & (!g843) & (!g844)));
	assign g851 = (((!g845) & (!g846) & (!g847) & (!g848) & (!g849) & (!g850)) + ((!g845) & (!g846) & (!g847) & (g848) & (!g849) & (!g850)) + ((!g845) & (!g846) & (!g847) & (g848) & (g849) & (g850)) + ((!g845) & (!g846) & (g847) & (!g848) & (!g849) & (!g850)) + ((!g845) & (!g846) & (g847) & (!g848) & (!g849) & (g850)) + ((!g845) & (!g846) & (g847) & (g848) & (!g849) & (!g850)) + ((!g845) & (!g846) & (g847) & (g848) & (!g849) & (g850)) + ((!g845) & (!g846) & (g847) & (g848) & (g849) & (g850)) + ((!g845) & (g846) & (!g847) & (!g848) & (!g849) & (!g850)) + ((!g845) & (g846) & (!g847) & (!g848) & (g849) & (!g850)) + ((!g845) & (g846) & (!g847) & (g848) & (!g849) & (!g850)) + ((!g845) & (g846) & (!g847) & (g848) & (g849) & (!g850)) + ((!g845) & (g846) & (!g847) & (g848) & (g849) & (g850)) + ((!g845) & (g846) & (g847) & (!g848) & (!g849) & (!g850)) + ((!g845) & (g846) & (g847) & (!g848) & (!g849) & (g850)) + ((!g845) & (g846) & (g847) & (!g848) & (g849) & (!g850)) + ((!g845) & (g846) & (g847) & (g848) & (!g849) & (!g850)) + ((!g845) & (g846) & (g847) & (g848) & (!g849) & (g850)) + ((!g845) & (g846) & (g847) & (g848) & (g849) & (!g850)) + ((!g845) & (g846) & (g847) & (g848) & (g849) & (g850)) + ((g845) & (!g846) & (!g847) & (g848) & (g849) & (g850)) + ((g845) & (!g846) & (g847) & (!g848) & (!g849) & (g850)) + ((g845) & (!g846) & (g847) & (g848) & (!g849) & (g850)) + ((g845) & (!g846) & (g847) & (g848) & (g849) & (g850)) + ((g845) & (g846) & (!g847) & (!g848) & (g849) & (!g850)) + ((g845) & (g846) & (!g847) & (g848) & (g849) & (!g850)) + ((g845) & (g846) & (!g847) & (g848) & (g849) & (g850)) + ((g845) & (g846) & (g847) & (!g848) & (!g849) & (g850)) + ((g845) & (g846) & (g847) & (!g848) & (g849) & (!g850)) + ((g845) & (g846) & (g847) & (g848) & (!g849) & (g850)) + ((g845) & (g846) & (g847) & (g848) & (g849) & (!g850)) + ((g845) & (g846) & (g847) & (g848) & (g849) & (g850)));
	assign g853 = (((!sk[22]) & (g851) & (!g852)) + ((!sk[22]) & (g851) & (g852)) + ((sk[22]) & (!g851) & (g852)) + ((sk[22]) & (g851) & (!g852)));
	assign g854 = (((!g839) & (!g840) & (!g841) & (!g842) & (!g849) & (g843)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g849) & (!g843)) + ((!g839) & (!g840) & (!g841) & (g842) & (g849) & (!g843)) + ((!g839) & (!g840) & (g841) & (!g842) & (g849) & (g843)) + ((!g839) & (!g840) & (g841) & (g842) & (!g849) & (g843)) + ((!g839) & (!g840) & (g841) & (g842) & (g849) & (!g843)) + ((!g839) & (g840) & (!g841) & (!g842) & (!g849) & (g843)) + ((!g839) & (g840) & (!g841) & (!g842) & (g849) & (!g843)) + ((!g839) & (g840) & (!g841) & (!g842) & (g849) & (g843)) + ((!g839) & (g840) & (g841) & (!g842) & (g849) & (g843)) + ((!g839) & (g840) & (g841) & (g842) & (g849) & (g843)) + ((g839) & (!g840) & (!g841) & (!g842) & (!g849) & (!g843)) + ((g839) & (!g840) & (!g841) & (!g842) & (g849) & (g843)) + ((g839) & (!g840) & (!g841) & (g842) & (!g849) & (!g843)) + ((g839) & (!g840) & (!g841) & (g842) & (g849) & (!g843)) + ((g839) & (!g840) & (g841) & (!g842) & (g849) & (!g843)) + ((g839) & (!g840) & (g841) & (!g842) & (g849) & (g843)) + ((g839) & (!g840) & (g841) & (g842) & (g849) & (!g843)) + ((g839) & (!g840) & (g841) & (g842) & (g849) & (g843)) + ((g839) & (g840) & (!g841) & (!g842) & (g849) & (!g843)) + ((g839) & (g840) & (!g841) & (!g842) & (g849) & (g843)) + ((g839) & (g840) & (!g841) & (g842) & (g849) & (g843)) + ((g839) & (g840) & (g841) & (!g842) & (!g849) & (!g843)) + ((g839) & (g840) & (g841) & (!g842) & (!g849) & (g843)) + ((g839) & (g840) & (g841) & (!g842) & (g849) & (!g843)) + ((g839) & (g840) & (g841) & (g842) & (!g849) & (g843)) + ((g839) & (g840) & (g841) & (g842) & (g849) & (!g843)));
	assign g855 = (((!g839) & (!g840) & (!g841) & (!g842) & (!g849) & (g843)) + ((!g839) & (!g840) & (!g841) & (!g842) & (g849) & (!g843)) + ((!g839) & (!g840) & (!g841) & (!g842) & (g849) & (g843)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g849) & (!g843)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g849) & (g843)) + ((!g839) & (!g840) & (!g841) & (g842) & (g849) & (g843)) + ((!g839) & (!g840) & (g841) & (!g842) & (g849) & (!g843)) + ((!g839) & (!g840) & (g841) & (g842) & (!g849) & (!g843)) + ((!g839) & (!g840) & (g841) & (g842) & (!g849) & (g843)) + ((!g839) & (!g840) & (g841) & (g842) & (g849) & (g843)) + ((!g839) & (g840) & (!g841) & (!g842) & (g849) & (g843)) + ((!g839) & (g840) & (!g841) & (g842) & (!g849) & (!g843)) + ((!g839) & (g840) & (!g841) & (g842) & (g849) & (!g843)) + ((!g839) & (g840) & (g841) & (!g842) & (g849) & (!g843)) + ((!g839) & (g840) & (g841) & (!g842) & (g849) & (g843)) + ((!g839) & (g840) & (g841) & (g842) & (!g849) & (!g843)) + ((g839) & (!g840) & (!g841) & (!g842) & (!g849) & (!g843)) + ((g839) & (!g840) & (!g841) & (g842) & (!g849) & (!g843)) + ((g839) & (!g840) & (!g841) & (g842) & (!g849) & (g843)) + ((g839) & (!g840) & (g841) & (!g842) & (!g849) & (g843)) + ((g839) & (!g840) & (g841) & (!g842) & (g849) & (g843)) + ((g839) & (!g840) & (g841) & (g842) & (!g849) & (!g843)) + ((g839) & (!g840) & (g841) & (g842) & (!g849) & (g843)) + ((g839) & (g840) & (!g841) & (g842) & (!g849) & (!g843)) + ((g839) & (g840) & (!g841) & (g842) & (g849) & (g843)) + ((g839) & (g840) & (g841) & (!g842) & (!g849) & (!g843)) + ((g839) & (g840) & (g841) & (!g842) & (!g849) & (g843)) + ((g839) & (g840) & (g841) & (!g842) & (g849) & (g843)) + ((g839) & (g840) & (g841) & (g842) & (!g849) & (!g843)) + ((g839) & (g840) & (g841) & (g842) & (!g849) & (g843)) + ((g839) & (g840) & (g841) & (g842) & (g849) & (!g843)));
	assign g856 = (((!g839) & (!g840) & (!g841) & (!g842) & (!g849) & (g843)) + ((!g839) & (!g840) & (!g841) & (g842) & (g849) & (!g843)) + ((!g839) & (!g840) & (g841) & (!g842) & (!g849) & (!g843)) + ((!g839) & (!g840) & (g841) & (!g842) & (g849) & (!g843)) + ((!g839) & (!g840) & (g841) & (g842) & (!g849) & (g843)) + ((!g839) & (!g840) & (g841) & (g842) & (g849) & (!g843)) + ((!g839) & (!g840) & (g841) & (g842) & (g849) & (g843)) + ((!g839) & (g840) & (!g841) & (!g842) & (!g849) & (!g843)) + ((!g839) & (g840) & (!g841) & (!g842) & (g849) & (!g843)) + ((!g839) & (g840) & (!g841) & (g842) & (!g849) & (!g843)) + ((!g839) & (g840) & (!g841) & (g842) & (g849) & (g843)) + ((!g839) & (g840) & (g841) & (!g842) & (g849) & (g843)) + ((!g839) & (g840) & (g841) & (g842) & (!g849) & (g843)) + ((!g839) & (g840) & (g841) & (g842) & (g849) & (!g843)) + ((g839) & (!g840) & (!g841) & (!g842) & (g849) & (g843)) + ((g839) & (!g840) & (!g841) & (g842) & (!g849) & (!g843)) + ((g839) & (!g840) & (!g841) & (g842) & (g849) & (!g843)) + ((g839) & (!g840) & (g841) & (!g842) & (!g849) & (!g843)) + ((g839) & (!g840) & (g841) & (!g842) & (!g849) & (g843)) + ((g839) & (!g840) & (g841) & (!g842) & (g849) & (!g843)) + ((g839) & (!g840) & (g841) & (!g842) & (g849) & (g843)) + ((g839) & (!g840) & (g841) & (g842) & (g849) & (!g843)) + ((g839) & (g840) & (!g841) & (!g842) & (!g849) & (g843)) + ((g839) & (g840) & (!g841) & (!g842) & (g849) & (g843)) + ((g839) & (g840) & (!g841) & (g842) & (!g849) & (g843)) + ((g839) & (g840) & (g841) & (!g842) & (!g849) & (!g843)) + ((g839) & (g840) & (g841) & (!g842) & (!g849) & (g843)) + ((g839) & (g840) & (g841) & (!g842) & (g849) & (g843)) + ((g839) & (g840) & (g841) & (g842) & (!g849) & (!g843)) + ((g839) & (g840) & (g841) & (g842) & (!g849) & (g843)) + ((g839) & (g840) & (g841) & (g842) & (g849) & (!g843)) + ((g839) & (g840) & (g841) & (g842) & (g849) & (g843)));
	assign g857 = (((!g839) & (!g840) & (!g841) & (!g842) & (g849) & (!g843)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g849) & (!g843)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g849) & (g843)) + ((!g839) & (!g840) & (g841) & (!g842) & (g849) & (g843)) + ((!g839) & (!g840) & (g841) & (g842) & (!g849) & (g843)) + ((!g839) & (g840) & (!g841) & (!g842) & (!g849) & (!g843)) + ((!g839) & (g840) & (!g841) & (!g842) & (g849) & (!g843)) + ((!g839) & (g840) & (!g841) & (g842) & (!g849) & (g843)) + ((!g839) & (g840) & (g841) & (!g842) & (!g849) & (g843)) + ((!g839) & (g840) & (g841) & (!g842) & (g849) & (!g843)) + ((!g839) & (g840) & (g841) & (!g842) & (g849) & (g843)) + ((!g839) & (g840) & (g841) & (g842) & (g849) & (!g843)) + ((!g839) & (g840) & (g841) & (g842) & (g849) & (g843)) + ((g839) & (!g840) & (!g841) & (!g842) & (!g849) & (!g843)) + ((g839) & (!g840) & (!g841) & (g842) & (!g849) & (!g843)) + ((g839) & (!g840) & (!g841) & (g842) & (!g849) & (g843)) + ((g839) & (!g840) & (!g841) & (g842) & (g849) & (!g843)) + ((g839) & (!g840) & (g841) & (!g842) & (!g849) & (!g843)) + ((g839) & (!g840) & (g841) & (!g842) & (g849) & (g843)) + ((g839) & (!g840) & (g841) & (g842) & (g849) & (!g843)) + ((g839) & (g840) & (!g841) & (!g842) & (!g849) & (!g843)) + ((g839) & (g840) & (!g841) & (g842) & (!g849) & (!g843)) + ((g839) & (g840) & (!g841) & (g842) & (g849) & (!g843)) + ((g839) & (g840) & (!g841) & (g842) & (g849) & (g843)) + ((g839) & (g840) & (g841) & (g842) & (!g849) & (g843)) + ((g839) & (g840) & (g841) & (g842) & (g849) & (g843)));
	assign g858 = (((!g854) & (!g855) & (!g856) & (!g857) & (!g844) & (!g850)) + ((!g854) & (!g855) & (!g856) & (!g857) & (g844) & (!g850)) + ((!g854) & (!g855) & (!g856) & (g857) & (!g844) & (!g850)) + ((!g854) & (!g855) & (!g856) & (g857) & (g844) & (!g850)) + ((!g854) & (!g855) & (!g856) & (g857) & (g844) & (g850)) + ((!g854) & (!g855) & (g856) & (!g857) & (!g844) & (!g850)) + ((!g854) & (!g855) & (g856) & (!g857) & (!g844) & (g850)) + ((!g854) & (!g855) & (g856) & (!g857) & (g844) & (!g850)) + ((!g854) & (!g855) & (g856) & (g857) & (!g844) & (!g850)) + ((!g854) & (!g855) & (g856) & (g857) & (!g844) & (g850)) + ((!g854) & (!g855) & (g856) & (g857) & (g844) & (!g850)) + ((!g854) & (!g855) & (g856) & (g857) & (g844) & (g850)) + ((!g854) & (g855) & (!g856) & (!g857) & (!g844) & (!g850)) + ((!g854) & (g855) & (!g856) & (g857) & (!g844) & (!g850)) + ((!g854) & (g855) & (!g856) & (g857) & (g844) & (g850)) + ((!g854) & (g855) & (g856) & (!g857) & (!g844) & (!g850)) + ((!g854) & (g855) & (g856) & (!g857) & (!g844) & (g850)) + ((!g854) & (g855) & (g856) & (g857) & (!g844) & (!g850)) + ((!g854) & (g855) & (g856) & (g857) & (!g844) & (g850)) + ((!g854) & (g855) & (g856) & (g857) & (g844) & (g850)) + ((g854) & (!g855) & (!g856) & (!g857) & (g844) & (!g850)) + ((g854) & (!g855) & (!g856) & (g857) & (g844) & (!g850)) + ((g854) & (!g855) & (!g856) & (g857) & (g844) & (g850)) + ((g854) & (!g855) & (g856) & (!g857) & (!g844) & (g850)) + ((g854) & (!g855) & (g856) & (!g857) & (g844) & (!g850)) + ((g854) & (!g855) & (g856) & (g857) & (!g844) & (g850)) + ((g854) & (!g855) & (g856) & (g857) & (g844) & (!g850)) + ((g854) & (!g855) & (g856) & (g857) & (g844) & (g850)) + ((g854) & (g855) & (!g856) & (g857) & (g844) & (g850)) + ((g854) & (g855) & (g856) & (!g857) & (!g844) & (g850)) + ((g854) & (g855) & (g856) & (g857) & (!g844) & (g850)) + ((g854) & (g855) & (g856) & (g857) & (g844) & (g850)));
	assign g860 = (((!sk[28]) & (g858) & (!g859)) + ((!sk[28]) & (g858) & (g859)) + ((sk[28]) & (!g858) & (g859)) + ((sk[28]) & (g858) & (!g859)));
	assign g861 = (((!g843) & (!g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((!g843) & (!g840) & (!g841) & (!g842) & (g849) & (g844)) + ((!g843) & (!g840) & (!g841) & (g842) & (!g849) & (g844)) + ((!g843) & (!g840) & (!g841) & (g842) & (g849) & (!g844)) + ((!g843) & (!g840) & (!g841) & (g842) & (g849) & (g844)) + ((!g843) & (!g840) & (g841) & (!g842) & (!g849) & (g844)) + ((!g843) & (!g840) & (g841) & (g842) & (!g849) & (!g844)) + ((!g843) & (!g840) & (g841) & (g842) & (g849) & (!g844)) + ((!g843) & (g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((!g843) & (g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((!g843) & (g840) & (!g841) & (g842) & (!g849) & (g844)) + ((!g843) & (g840) & (g841) & (!g842) & (!g849) & (!g844)) + ((!g843) & (g840) & (g841) & (!g842) & (!g849) & (g844)) + ((!g843) & (g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g843) & (g840) & (g841) & (!g842) & (g849) & (g844)) + ((g843) & (!g840) & (!g841) & (g842) & (!g849) & (g844)) + ((g843) & (!g840) & (!g841) & (g842) & (g849) & (g844)) + ((g843) & (g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((g843) & (g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((g843) & (g840) & (!g841) & (g842) & (g849) & (!g844)) + ((g843) & (g840) & (g841) & (g842) & (!g849) & (!g844)) + ((g843) & (g840) & (g841) & (g842) & (!g849) & (g844)));
	assign g862 = (((!g843) & (!g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((!g843) & (!g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((!g843) & (!g840) & (!g841) & (g842) & (g849) & (g844)) + ((!g843) & (!g840) & (g841) & (!g842) & (!g849) & (!g844)) + ((!g843) & (!g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g843) & (!g840) & (g841) & (g842) & (!g849) & (g844)) + ((!g843) & (g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((!g843) & (g840) & (!g841) & (!g842) & (g849) & (g844)) + ((!g843) & (g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((!g843) & (g840) & (!g841) & (g842) & (!g849) & (g844)) + ((!g843) & (g840) & (!g841) & (g842) & (g849) & (g844)) + ((!g843) & (g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g843) & (g840) & (g841) & (!g842) & (g849) & (g844)) + ((!g843) & (g840) & (g841) & (g842) & (g849) & (!g844)) + ((g843) & (!g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((g843) & (!g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((g843) & (!g840) & (!g841) & (!g842) & (g849) & (g844)) + ((g843) & (!g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((g843) & (!g840) & (!g841) & (g842) & (!g849) & (g844)) + ((g843) & (!g840) & (!g841) & (g842) & (g849) & (!g844)) + ((g843) & (!g840) & (g841) & (g842) & (!g849) & (!g844)) + ((g843) & (g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((g843) & (g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((g843) & (g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((g843) & (g840) & (!g841) & (g842) & (g849) & (!g844)) + ((g843) & (g840) & (!g841) & (g842) & (g849) & (g844)) + ((g843) & (g840) & (g841) & (!g842) & (!g849) & (!g844)) + ((g843) & (g840) & (g841) & (!g842) & (g849) & (!g844)) + ((g843) & (g840) & (g841) & (g842) & (!g849) & (g844)) + ((g843) & (g840) & (g841) & (g842) & (g849) & (g844)));
	assign g863 = (((!g843) & (!g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((!g843) & (!g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((!g843) & (!g840) & (!g841) & (g842) & (!g849) & (g844)) + ((!g843) & (!g840) & (g841) & (!g842) & (!g849) & (g844)) + ((!g843) & (!g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g843) & (!g840) & (g841) & (g842) & (!g849) & (g844)) + ((!g843) & (g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((!g843) & (g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((!g843) & (g840) & (!g841) & (g842) & (g849) & (!g844)) + ((!g843) & (g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g843) & (g840) & (g841) & (g842) & (!g849) & (!g844)) + ((!g843) & (g840) & (g841) & (g842) & (g849) & (!g844)) + ((g843) & (!g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((g843) & (!g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((g843) & (!g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((g843) & (!g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((g843) & (!g840) & (!g841) & (g842) & (!g849) & (g844)) + ((g843) & (!g840) & (!g841) & (g842) & (g849) & (!g844)) + ((g843) & (!g840) & (!g841) & (g842) & (g849) & (g844)) + ((g843) & (!g840) & (g841) & (!g842) & (!g849) & (g844)) + ((g843) & (!g840) & (g841) & (!g842) & (g849) & (!g844)) + ((g843) & (!g840) & (g841) & (g842) & (!g849) & (!g844)) + ((g843) & (!g840) & (g841) & (g842) & (g849) & (g844)) + ((g843) & (g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((g843) & (g840) & (!g841) & (!g842) & (g849) & (g844)) + ((g843) & (g840) & (g841) & (!g842) & (g849) & (g844)) + ((g843) & (g840) & (g841) & (g842) & (!g849) & (!g844)) + ((g843) & (g840) & (g841) & (g842) & (!g849) & (g844)) + ((g843) & (g840) & (g841) & (g842) & (g849) & (g844)));
	assign g864 = (((!g843) & (!g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((!g843) & (!g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((!g843) & (!g840) & (!g841) & (!g842) & (g849) & (g844)) + ((!g843) & (!g840) & (!g841) & (g842) & (!g849) & (g844)) + ((!g843) & (!g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g843) & (!g840) & (g841) & (g842) & (g849) & (g844)) + ((!g843) & (g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((!g843) & (g840) & (!g841) & (g842) & (!g849) & (g844)) + ((!g843) & (g840) & (!g841) & (g842) & (g849) & (g844)) + ((!g843) & (g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g843) & (g840) & (g841) & (!g842) & (g849) & (g844)) + ((!g843) & (g840) & (g841) & (g842) & (!g849) & (!g844)) + ((!g843) & (g840) & (g841) & (g842) & (!g849) & (g844)) + ((!g843) & (g840) & (g841) & (g842) & (g849) & (!g844)) + ((!g843) & (g840) & (g841) & (g842) & (g849) & (g844)) + ((g843) & (!g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((g843) & (!g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((g843) & (!g840) & (!g841) & (!g842) & (g849) & (g844)) + ((g843) & (!g840) & (!g841) & (g842) & (g849) & (g844)) + ((g843) & (!g840) & (g841) & (!g842) & (!g849) & (g844)) + ((g843) & (!g840) & (g841) & (!g842) & (g849) & (!g844)) + ((g843) & (!g840) & (g841) & (g842) & (g849) & (!g844)) + ((g843) & (g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((g843) & (g840) & (!g841) & (g842) & (!g849) & (g844)) + ((g843) & (g840) & (!g841) & (g842) & (g849) & (!g844)) + ((g843) & (g840) & (g841) & (!g842) & (g849) & (g844)) + ((g843) & (g840) & (g841) & (g842) & (!g849) & (!g844)));
	assign g865 = (((!g861) & (!g862) & (!g863) & (!g864) & (!g839) & (g850)) + ((!g861) & (!g862) & (!g863) & (!g864) & (g839) & (!g850)) + ((!g861) & (!g862) & (!g863) & (!g864) & (g839) & (g850)) + ((!g861) & (!g862) & (!g863) & (g864) & (!g839) & (g850)) + ((!g861) & (!g862) & (!g863) & (g864) & (g839) & (!g850)) + ((!g861) & (!g862) & (g863) & (!g864) & (g839) & (!g850)) + ((!g861) & (!g862) & (g863) & (!g864) & (g839) & (g850)) + ((!g861) & (!g862) & (g863) & (g864) & (g839) & (!g850)) + ((!g861) & (g862) & (!g863) & (!g864) & (!g839) & (g850)) + ((!g861) & (g862) & (!g863) & (!g864) & (g839) & (g850)) + ((!g861) & (g862) & (!g863) & (g864) & (!g839) & (g850)) + ((!g861) & (g862) & (g863) & (!g864) & (g839) & (g850)) + ((g861) & (!g862) & (!g863) & (!g864) & (!g839) & (!g850)) + ((g861) & (!g862) & (!g863) & (!g864) & (!g839) & (g850)) + ((g861) & (!g862) & (!g863) & (!g864) & (g839) & (!g850)) + ((g861) & (!g862) & (!g863) & (!g864) & (g839) & (g850)) + ((g861) & (!g862) & (!g863) & (g864) & (!g839) & (!g850)) + ((g861) & (!g862) & (!g863) & (g864) & (!g839) & (g850)) + ((g861) & (!g862) & (!g863) & (g864) & (g839) & (!g850)) + ((g861) & (!g862) & (g863) & (!g864) & (!g839) & (!g850)) + ((g861) & (!g862) & (g863) & (!g864) & (g839) & (!g850)) + ((g861) & (!g862) & (g863) & (!g864) & (g839) & (g850)) + ((g861) & (!g862) & (g863) & (g864) & (!g839) & (!g850)) + ((g861) & (!g862) & (g863) & (g864) & (g839) & (!g850)) + ((g861) & (g862) & (!g863) & (!g864) & (!g839) & (!g850)) + ((g861) & (g862) & (!g863) & (!g864) & (!g839) & (g850)) + ((g861) & (g862) & (!g863) & (!g864) & (g839) & (g850)) + ((g861) & (g862) & (!g863) & (g864) & (!g839) & (!g850)) + ((g861) & (g862) & (!g863) & (g864) & (!g839) & (g850)) + ((g861) & (g862) & (g863) & (!g864) & (!g839) & (!g850)) + ((g861) & (g862) & (g863) & (!g864) & (g839) & (g850)) + ((g861) & (g862) & (g863) & (g864) & (!g839) & (!g850)));
	assign g867 = (((!g865) & (sk[34]) & (g866)) + ((g865) & (!sk[34]) & (!g866)) + ((g865) & (!sk[34]) & (g866)) + ((g865) & (sk[34]) & (!g866)));
	assign g868 = (((!g839) & (!g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (g849) & (g844)) + ((!g839) & (!g840) & (g841) & (g842) & (!g849) & (!g844)) + ((!g839) & (!g840) & (g841) & (g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (g841) & (g842) & (g849) & (g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (g840) & (g841) & (!g842) & (!g849) & (!g844)) + ((!g839) & (g840) & (g841) & (g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((g839) & (!g840) & (g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (g841) & (!g842) & (!g849) & (g844)) + ((g839) & (!g840) & (g841) & (!g842) & (g849) & (!g844)) + ((g839) & (!g840) & (g841) & (g842) & (!g849) & (g844)) + ((g839) & (g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((g839) & (g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((g839) & (g840) & (!g841) & (g842) & (g849) & (!g844)) + ((g839) & (g840) & (g841) & (!g842) & (!g849) & (g844)) + ((g839) & (g840) & (g841) & (!g842) & (g849) & (g844)));
	assign g869 = (((!g839) & (!g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (!g841) & (!g842) & (g849) & (g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (g841) & (g842) & (!g849) & (!g844)) + ((!g839) & (!g840) & (g841) & (g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (g841) & (g842) & (g849) & (g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (g849) & (g844)) + ((!g839) & (g840) & (!g841) & (g842) & (g849) & (g844)) + ((!g839) & (g840) & (g841) & (!g842) & (!g849) & (!g844)) + ((!g839) & (g840) & (g841) & (!g842) & (!g849) & (g844)) + ((!g839) & (g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (g840) & (g841) & (g842) & (!g849) & (g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((g839) & (!g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (!g841) & (g842) & (!g849) & (g844)) + ((g839) & (!g840) & (!g841) & (g842) & (g849) & (g844)) + ((g839) & (!g840) & (g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (g841) & (!g842) & (!g849) & (g844)) + ((g839) & (!g840) & (g841) & (!g842) & (g849) & (g844)) + ((g839) & (!g840) & (g841) & (g842) & (!g849) & (g844)) + ((g839) & (g840) & (!g841) & (g842) & (!g849) & (g844)) + ((g839) & (g840) & (!g841) & (g842) & (g849) & (!g844)) + ((g839) & (g840) & (g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (g840) & (g841) & (g842) & (!g849) & (!g844)));
	assign g870 = (((!g839) & (!g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (!g841) & (!g842) & (g849) & (g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (g841) & (!g842) & (g849) & (g844)) + ((!g839) & (!g840) & (g841) & (g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (g841) & (g842) & (g849) & (g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (g849) & (g844)) + ((!g839) & (g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((!g839) & (g840) & (!g841) & (g842) & (!g849) & (g844)) + ((!g839) & (g840) & (g841) & (!g842) & (!g849) & (g844)) + ((!g839) & (g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (g840) & (g841) & (g842) & (g849) & (g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (g849) & (g844)) + ((g839) & (!g840) & (!g841) & (g842) & (g849) & (g844)) + ((g839) & (!g840) & (g841) & (g842) & (!g849) & (!g844)) + ((g839) & (g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((g839) & (g840) & (!g841) & (g842) & (g849) & (g844)) + ((g839) & (g840) & (g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (g840) & (g841) & (!g842) & (!g849) & (g844)) + ((g839) & (g840) & (g841) & (!g842) & (g849) & (g844)) + ((g839) & (g840) & (g841) & (g842) & (!g849) & (!g844)) + ((g839) & (g840) & (g841) & (g842) & (g849) & (g844)));
	assign g871 = (((!g839) & (!g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (!g841) & (g842) & (g849) & (g844)) + ((!g839) & (!g840) & (g841) & (g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (g841) & (g842) & (g849) & (g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (!g849) & (!g844)) + ((!g839) & (g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (g840) & (!g841) & (g842) & (!g849) & (!g844)) + ((!g839) & (g840) & (!g841) & (g842) & (!g849) & (g844)) + ((!g839) & (g840) & (!g841) & (g842) & (g849) & (!g844)) + ((!g839) & (g840) & (g841) & (!g842) & (!g849) & (!g844)) + ((!g839) & (g840) & (g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (g840) & (g841) & (!g842) & (g849) & (g844)) + ((g839) & (!g840) & (!g841) & (!g842) & (g849) & (g844)) + ((g839) & (!g840) & (!g841) & (g842) & (g849) & (!g844)) + ((g839) & (!g840) & (g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (g841) & (!g842) & (g849) & (!g844)) + ((g839) & (!g840) & (g841) & (!g842) & (g849) & (g844)) + ((g839) & (!g840) & (g841) & (g842) & (!g849) & (g844)) + ((g839) & (!g840) & (g841) & (g842) & (g849) & (!g844)) + ((g839) & (!g840) & (g841) & (g842) & (g849) & (g844)) + ((g839) & (g840) & (!g841) & (!g842) & (!g849) & (g844)) + ((g839) & (g840) & (!g841) & (!g842) & (g849) & (!g844)) + ((g839) & (g840) & (g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (g840) & (g841) & (!g842) & (!g849) & (g844)) + ((g839) & (g840) & (g841) & (g842) & (g849) & (g844)));
	assign g872 = (((!g868) & (!g869) & (!g870) & (!g871) & (!g850) & (g843)) + ((!g868) & (!g869) & (!g870) & (!g871) & (g850) & (!g843)) + ((!g868) & (!g869) & (!g870) & (!g871) & (g850) & (g843)) + ((!g868) & (!g869) & (!g870) & (g871) & (!g850) & (g843)) + ((!g868) & (!g869) & (!g870) & (g871) & (g850) & (!g843)) + ((!g868) & (!g869) & (g870) & (!g871) & (g850) & (!g843)) + ((!g868) & (!g869) & (g870) & (!g871) & (g850) & (g843)) + ((!g868) & (!g869) & (g870) & (g871) & (g850) & (!g843)) + ((!g868) & (g869) & (!g870) & (!g871) & (!g850) & (g843)) + ((!g868) & (g869) & (!g870) & (!g871) & (g850) & (g843)) + ((!g868) & (g869) & (!g870) & (g871) & (!g850) & (g843)) + ((!g868) & (g869) & (g870) & (!g871) & (g850) & (g843)) + ((g868) & (!g869) & (!g870) & (!g871) & (!g850) & (!g843)) + ((g868) & (!g869) & (!g870) & (!g871) & (!g850) & (g843)) + ((g868) & (!g869) & (!g870) & (!g871) & (g850) & (!g843)) + ((g868) & (!g869) & (!g870) & (!g871) & (g850) & (g843)) + ((g868) & (!g869) & (!g870) & (g871) & (!g850) & (!g843)) + ((g868) & (!g869) & (!g870) & (g871) & (!g850) & (g843)) + ((g868) & (!g869) & (!g870) & (g871) & (g850) & (!g843)) + ((g868) & (!g869) & (g870) & (!g871) & (!g850) & (!g843)) + ((g868) & (!g869) & (g870) & (!g871) & (g850) & (!g843)) + ((g868) & (!g869) & (g870) & (!g871) & (g850) & (g843)) + ((g868) & (!g869) & (g870) & (g871) & (!g850) & (!g843)) + ((g868) & (!g869) & (g870) & (g871) & (g850) & (!g843)) + ((g868) & (g869) & (!g870) & (!g871) & (!g850) & (!g843)) + ((g868) & (g869) & (!g870) & (!g871) & (!g850) & (g843)) + ((g868) & (g869) & (!g870) & (!g871) & (g850) & (g843)) + ((g868) & (g869) & (!g870) & (g871) & (!g850) & (!g843)) + ((g868) & (g869) & (!g870) & (g871) & (!g850) & (g843)) + ((g868) & (g869) & (g870) & (!g871) & (!g850) & (!g843)) + ((g868) & (g869) & (g870) & (!g871) & (g850) & (g843)) + ((g868) & (g869) & (g870) & (g871) & (!g850) & (!g843)));
	assign g874 = (((!g872) & (sk[40]) & (g873)) + ((g872) & (!sk[40]) & (!g873)) + ((g872) & (!sk[40]) & (g873)) + ((g872) & (sk[40]) & (!g873)));
	assign g875 = (((!g839) & (!g840) & (!g843) & (!g850) & (!g849) & (g844)) + ((!g839) & (!g840) & (g843) & (!g850) & (!g849) & (g844)) + ((!g839) & (!g840) & (g843) & (!g850) & (g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (!g850) & (g849) & (g844)) + ((!g839) & (!g840) & (g843) & (g850) & (!g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (g850) & (g849) & (!g844)) + ((!g839) & (g840) & (!g843) & (!g850) & (!g849) & (!g844)) + ((!g839) & (g840) & (!g843) & (!g850) & (!g849) & (g844)) + ((!g839) & (g840) & (!g843) & (g850) & (!g849) & (!g844)) + ((!g839) & (g840) & (!g843) & (g850) & (!g849) & (g844)) + ((!g839) & (g840) & (!g843) & (g850) & (g849) & (g844)) + ((!g839) & (g840) & (g843) & (g850) & (!g849) & (g844)) + ((!g839) & (g840) & (g843) & (g850) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g850) & (!g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g850) & (!g849) & (g844)) + ((g839) & (!g840) & (!g843) & (g850) & (!g849) & (g844)) + ((g839) & (!g840) & (g843) & (!g850) & (g849) & (!g844)) + ((g839) & (!g840) & (g843) & (g850) & (!g849) & (!g844)) + ((g839) & (!g840) & (g843) & (g850) & (!g849) & (g844)) + ((g839) & (!g840) & (g843) & (g850) & (g849) & (!g844)) + ((g839) & (g840) & (!g843) & (!g850) & (!g849) & (!g844)) + ((g839) & (g840) & (!g843) & (!g850) & (g849) & (!g844)) + ((g839) & (g840) & (!g843) & (g850) & (g849) & (!g844)) + ((g839) & (g840) & (g843) & (!g850) & (!g849) & (!g844)) + ((g839) & (g840) & (g843) & (!g850) & (!g849) & (g844)) + ((g839) & (g840) & (g843) & (g850) & (!g849) & (g844)));
	assign g876 = (((!g839) & (!g840) & (!g843) & (!g850) & (!g849) & (!g844)) + ((!g839) & (!g840) & (!g843) & (!g850) & (!g849) & (g844)) + ((!g839) & (!g840) & (!g843) & (!g850) & (g849) & (!g844)) + ((!g839) & (!g840) & (!g843) & (!g850) & (g849) & (g844)) + ((!g839) & (!g840) & (!g843) & (g850) & (!g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (!g850) & (!g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (!g850) & (g849) & (g844)) + ((!g839) & (!g840) & (g843) & (g850) & (!g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (g850) & (g849) & (g844)) + ((!g839) & (g840) & (!g843) & (!g850) & (!g849) & (g844)) + ((!g839) & (g840) & (!g843) & (g850) & (g849) & (!g844)) + ((!g839) & (g840) & (g843) & (!g850) & (!g849) & (!g844)) + ((!g839) & (g840) & (g843) & (!g850) & (!g849) & (g844)) + ((!g839) & (g840) & (g843) & (!g850) & (g849) & (!g844)) + ((!g839) & (g840) & (g843) & (!g850) & (g849) & (g844)) + ((!g839) & (g840) & (g843) & (g850) & (!g849) & (!g844)) + ((!g839) & (g840) & (g843) & (g850) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g850) & (!g849) & (g844)) + ((g839) & (!g840) & (!g843) & (!g850) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g850) & (g849) & (g844)) + ((g839) & (!g840) & (!g843) & (g850) & (!g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (g850) & (g849) & (g844)) + ((g839) & (!g840) & (g843) & (!g850) & (g849) & (!g844)) + ((g839) & (!g840) & (g843) & (!g850) & (g849) & (g844)) + ((g839) & (!g840) & (g843) & (g850) & (!g849) & (g844)) + ((g839) & (g840) & (!g843) & (!g850) & (g849) & (!g844)) + ((g839) & (g840) & (!g843) & (!g850) & (g849) & (g844)) + ((g839) & (g840) & (!g843) & (g850) & (!g849) & (!g844)) + ((g839) & (g840) & (!g843) & (g850) & (!g849) & (g844)) + ((g839) & (g840) & (g843) & (!g850) & (g849) & (!g844)) + ((g839) & (g840) & (g843) & (!g850) & (g849) & (g844)) + ((g839) & (g840) & (g843) & (g850) & (!g849) & (g844)));
	assign g877 = (((!g839) & (!g840) & (!g843) & (!g850) & (!g849) & (!g844)) + ((!g839) & (!g840) & (!g843) & (!g850) & (!g849) & (g844)) + ((!g839) & (!g840) & (g843) & (!g850) & (!g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (!g850) & (g849) & (g844)) + ((!g839) & (!g840) & (g843) & (g850) & (!g849) & (g844)) + ((!g839) & (g840) & (!g843) & (g850) & (!g849) & (!g844)) + ((!g839) & (g840) & (!g843) & (g850) & (g849) & (!g844)) + ((!g839) & (g840) & (!g843) & (g850) & (g849) & (g844)) + ((!g839) & (g840) & (g843) & (!g850) & (!g849) & (!g844)) + ((!g839) & (g840) & (g843) & (!g850) & (g849) & (!g844)) + ((!g839) & (g840) & (g843) & (!g850) & (g849) & (g844)) + ((!g839) & (g840) & (g843) & (g850) & (!g849) & (!g844)) + ((!g839) & (g840) & (g843) & (g850) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g850) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g850) & (g849) & (g844)) + ((g839) & (!g840) & (!g843) & (g850) & (!g849) & (g844)) + ((g839) & (!g840) & (!g843) & (g850) & (g849) & (g844)) + ((g839) & (!g840) & (g843) & (!g850) & (!g849) & (!g844)) + ((g839) & (!g840) & (g843) & (!g850) & (!g849) & (g844)) + ((g839) & (!g840) & (g843) & (!g850) & (g849) & (g844)) + ((g839) & (!g840) & (g843) & (g850) & (!g849) & (!g844)) + ((g839) & (!g840) & (g843) & (g850) & (!g849) & (g844)) + ((g839) & (!g840) & (g843) & (g850) & (g849) & (!g844)) + ((g839) & (!g840) & (g843) & (g850) & (g849) & (g844)) + ((g839) & (g840) & (!g843) & (!g850) & (!g849) & (g844)) + ((g839) & (g840) & (!g843) & (g850) & (!g849) & (!g844)) + ((g839) & (g840) & (!g843) & (g850) & (g849) & (!g844)) + ((g839) & (g840) & (g843) & (!g850) & (!g849) & (!g844)) + ((g839) & (g840) & (g843) & (!g850) & (!g849) & (g844)) + ((g839) & (g840) & (g843) & (!g850) & (g849) & (!g844)) + ((g839) & (g840) & (g843) & (g850) & (!g849) & (!g844)) + ((g839) & (g840) & (g843) & (g850) & (g849) & (!g844)));
	assign g878 = (((!g839) & (!g840) & (!g843) & (!g850) & (g849) & (g844)) + ((!g839) & (!g840) & (!g843) & (g850) & (!g849) & (!g844)) + ((!g839) & (!g840) & (!g843) & (g850) & (g849) & (g844)) + ((!g839) & (!g840) & (g843) & (!g850) & (!g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (!g850) & (g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (g850) & (!g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (g850) & (!g849) & (g844)) + ((!g839) & (!g840) & (g843) & (g850) & (g849) & (!g844)) + ((!g839) & (g840) & (!g843) & (!g850) & (!g849) & (!g844)) + ((!g839) & (g840) & (!g843) & (g850) & (!g849) & (g844)) + ((!g839) & (g840) & (!g843) & (g850) & (g849) & (!g844)) + ((!g839) & (g840) & (!g843) & (g850) & (g849) & (g844)) + ((!g839) & (g840) & (g843) & (!g850) & (!g849) & (!g844)) + ((!g839) & (g840) & (g843) & (g850) & (!g849) & (!g844)) + ((!g839) & (g840) & (g843) & (g850) & (!g849) & (g844)) + ((g839) & (!g840) & (!g843) & (!g850) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g850) & (g849) & (g844)) + ((g839) & (!g840) & (g843) & (!g850) & (!g849) & (!g844)) + ((g839) & (!g840) & (g843) & (!g850) & (g849) & (!g844)) + ((g839) & (!g840) & (g843) & (g850) & (g849) & (!g844)) + ((g839) & (g840) & (!g843) & (!g850) & (g849) & (!g844)) + ((g839) & (g840) & (!g843) & (g850) & (g849) & (g844)) + ((g839) & (g840) & (g843) & (!g850) & (!g849) & (!g844)) + ((g839) & (g840) & (g843) & (!g850) & (!g849) & (g844)) + ((g839) & (g840) & (g843) & (!g850) & (g849) & (!g844)) + ((g839) & (g840) & (g843) & (g850) & (!g849) & (!g844)));
	assign g879 = (((!g875) & (!g876) & (!g877) & (!g878) & (g841) & (g842)) + ((!g875) & (!g876) & (g877) & (!g878) & (!g841) & (g842)) + ((!g875) & (!g876) & (g877) & (!g878) & (g841) & (g842)) + ((!g875) & (!g876) & (g877) & (g878) & (!g841) & (g842)) + ((!g875) & (g876) & (!g877) & (!g878) & (g841) & (!g842)) + ((!g875) & (g876) & (!g877) & (!g878) & (g841) & (g842)) + ((!g875) & (g876) & (!g877) & (g878) & (g841) & (!g842)) + ((!g875) & (g876) & (g877) & (!g878) & (!g841) & (g842)) + ((!g875) & (g876) & (g877) & (!g878) & (g841) & (!g842)) + ((!g875) & (g876) & (g877) & (!g878) & (g841) & (g842)) + ((!g875) & (g876) & (g877) & (g878) & (!g841) & (g842)) + ((!g875) & (g876) & (g877) & (g878) & (g841) & (!g842)) + ((g875) & (!g876) & (!g877) & (!g878) & (!g841) & (!g842)) + ((g875) & (!g876) & (!g877) & (!g878) & (g841) & (g842)) + ((g875) & (!g876) & (!g877) & (g878) & (!g841) & (!g842)) + ((g875) & (!g876) & (g877) & (!g878) & (!g841) & (!g842)) + ((g875) & (!g876) & (g877) & (!g878) & (!g841) & (g842)) + ((g875) & (!g876) & (g877) & (!g878) & (g841) & (g842)) + ((g875) & (!g876) & (g877) & (g878) & (!g841) & (!g842)) + ((g875) & (!g876) & (g877) & (g878) & (!g841) & (g842)) + ((g875) & (g876) & (!g877) & (!g878) & (!g841) & (!g842)) + ((g875) & (g876) & (!g877) & (!g878) & (g841) & (!g842)) + ((g875) & (g876) & (!g877) & (!g878) & (g841) & (g842)) + ((g875) & (g876) & (!g877) & (g878) & (!g841) & (!g842)) + ((g875) & (g876) & (!g877) & (g878) & (g841) & (!g842)) + ((g875) & (g876) & (g877) & (!g878) & (!g841) & (!g842)) + ((g875) & (g876) & (g877) & (!g878) & (!g841) & (g842)) + ((g875) & (g876) & (g877) & (!g878) & (g841) & (!g842)) + ((g875) & (g876) & (g877) & (!g878) & (g841) & (g842)) + ((g875) & (g876) & (g877) & (g878) & (!g841) & (!g842)) + ((g875) & (g876) & (g877) & (g878) & (!g841) & (g842)) + ((g875) & (g876) & (g877) & (g878) & (g841) & (!g842)));
	assign g881 = (((!g879) & (sk[46]) & (g880)) + ((g879) & (!sk[46]) & (!g880)) + ((g879) & (!sk[46]) & (g880)) + ((g879) & (sk[46]) & (!g880)));
	assign g882 = (((!g839) & (!g840) & (!g843) & (!g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (!g843) & (!g842) & (g849) & (g844)) + ((!g839) & (!g840) & (!g843) & (g842) & (g849) & (g844)) + ((!g839) & (!g840) & (g843) & (!g842) & (!g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (!g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (g843) & (!g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (!g842) & (g849) & (g844)) + ((!g839) & (!g840) & (g843) & (g842) & (!g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (g842) & (!g849) & (g844)) + ((!g839) & (g840) & (!g843) & (!g842) & (!g849) & (g844)) + ((!g839) & (g840) & (!g843) & (!g842) & (g849) & (!g844)) + ((!g839) & (g840) & (!g843) & (g842) & (g849) & (g844)) + ((!g839) & (g840) & (g843) & (!g842) & (g849) & (!g844)) + ((!g839) & (g840) & (g843) & (!g842) & (g849) & (g844)) + ((!g839) & (g840) & (g843) & (g842) & (!g849) & (!g844)) + ((!g839) & (g840) & (g843) & (g842) & (!g849) & (g844)) + ((!g839) & (g840) & (g843) & (g842) & (g849) & (g844)) + ((g839) & (!g840) & (!g843) & (!g842) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g842) & (g849) & (g844)) + ((g839) & (!g840) & (!g843) & (g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (g842) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (g842) & (g849) & (g844)) + ((g839) & (!g840) & (g843) & (!g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (g843) & (!g842) & (g849) & (!g844)) + ((g839) & (!g840) & (g843) & (g842) & (g849) & (!g844)) + ((g839) & (g840) & (!g843) & (!g842) & (g849) & (g844)) + ((g839) & (g840) & (g843) & (!g842) & (!g849) & (!g844)) + ((g839) & (g840) & (g843) & (!g842) & (g849) & (g844)));
	assign g883 = (((!g839) & (!g840) & (!g843) & (!g842) & (!g849) & (!g844)) + ((!g839) & (!g840) & (!g843) & (g842) & (!g849) & (!g844)) + ((!g839) & (!g840) & (!g843) & (g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (!g843) & (g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (!g842) & (g849) & (g844)) + ((!g839) & (!g840) & (g843) & (g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (g843) & (g842) & (g849) & (g844)) + ((!g839) & (g840) & (!g843) & (!g842) & (!g849) & (!g844)) + ((!g839) & (g840) & (!g843) & (!g842) & (g849) & (!g844)) + ((!g839) & (g840) & (g843) & (!g842) & (!g849) & (g844)) + ((!g839) & (g840) & (g843) & (!g842) & (g849) & (g844)) + ((!g839) & (g840) & (g843) & (g842) & (!g849) & (g844)) + ((!g839) & (g840) & (g843) & (g842) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g842) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g842) & (g849) & (g844)) + ((g839) & (!g840) & (!g843) & (g842) & (!g849) & (g844)) + ((g839) & (!g840) & (!g843) & (g842) & (g849) & (g844)) + ((g839) & (!g840) & (g843) & (g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (g843) & (g842) & (!g849) & (g844)) + ((g839) & (!g840) & (g843) & (g842) & (g849) & (g844)) + ((g839) & (g840) & (!g843) & (!g842) & (!g849) & (g844)) + ((g839) & (g840) & (!g843) & (!g842) & (g849) & (!g844)) + ((g839) & (g840) & (!g843) & (g842) & (g849) & (!g844)) + ((g839) & (g840) & (g843) & (!g842) & (!g849) & (g844)) + ((g839) & (g840) & (g843) & (!g842) & (g849) & (g844)) + ((g839) & (g840) & (g843) & (g842) & (!g849) & (!g844)) + ((g839) & (g840) & (g843) & (g842) & (g849) & (g844)));
	assign g884 = (((!g839) & (!g840) & (!g843) & (!g842) & (g849) & (g844)) + ((!g839) & (!g840) & (!g843) & (g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (!g842) & (!g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (!g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (g843) & (!g842) & (g849) & (g844)) + ((!g839) & (!g840) & (g843) & (g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (g843) & (g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (g843) & (g842) & (g849) & (g844)) + ((!g839) & (g840) & (!g843) & (!g842) & (g849) & (!g844)) + ((!g839) & (g840) & (!g843) & (!g842) & (g849) & (g844)) + ((!g839) & (g840) & (g843) & (!g842) & (!g849) & (!g844)) + ((!g839) & (g840) & (g843) & (g842) & (!g849) & (g844)) + ((!g839) & (g840) & (g843) & (g842) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g842) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (!g842) & (g849) & (g844)) + ((g839) & (!g840) & (!g843) & (g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (g842) & (!g849) & (g844)) + ((g839) & (!g840) & (g843) & (!g842) & (!g849) & (g844)) + ((g839) & (!g840) & (g843) & (!g842) & (g849) & (g844)) + ((g839) & (!g840) & (g843) & (g842) & (g849) & (!g844)) + ((g839) & (g840) & (!g843) & (!g842) & (!g849) & (!g844)) + ((g839) & (g840) & (!g843) & (!g842) & (!g849) & (g844)) + ((g839) & (g840) & (!g843) & (!g842) & (g849) & (g844)) + ((g839) & (g840) & (!g843) & (g842) & (!g849) & (g844)) + ((g839) & (g840) & (!g843) & (g842) & (g849) & (!g844)) + ((g839) & (g840) & (g843) & (!g842) & (!g849) & (g844)) + ((g839) & (g840) & (g843) & (!g842) & (g849) & (!g844)) + ((g839) & (g840) & (g843) & (g842) & (!g849) & (!g844)) + ((g839) & (g840) & (g843) & (g842) & (g849) & (!g844)) + ((g839) & (g840) & (g843) & (g842) & (g849) & (g844)));
	assign g885 = (((!g839) & (!g840) & (!g843) & (!g842) & (g849) & (!g844)) + ((!g839) & (!g840) & (!g843) & (g842) & (!g849) & (!g844)) + ((!g839) & (!g840) & (!g843) & (g842) & (g849) & (g844)) + ((!g839) & (!g840) & (g843) & (!g842) & (!g849) & (g844)) + ((!g839) & (!g840) & (g843) & (!g842) & (g849) & (g844)) + ((!g839) & (!g840) & (g843) & (g842) & (g849) & (g844)) + ((!g839) & (g840) & (!g843) & (!g842) & (!g849) & (g844)) + ((!g839) & (g840) & (!g843) & (g842) & (!g849) & (g844)) + ((!g839) & (g840) & (!g843) & (g842) & (g849) & (g844)) + ((!g839) & (g840) & (g843) & (!g842) & (!g849) & (!g844)) + ((!g839) & (g840) & (g843) & (!g842) & (g849) & (!g844)) + ((!g839) & (g840) & (g843) & (g842) & (!g849) & (g844)) + ((!g839) & (g840) & (g843) & (g842) & (g849) & (g844)) + ((g839) & (!g840) & (!g843) & (!g842) & (g849) & (!g844)) + ((g839) & (!g840) & (!g843) & (g842) & (g849) & (g844)) + ((g839) & (!g840) & (g843) & (!g842) & (!g849) & (!g844)) + ((g839) & (!g840) & (g843) & (!g842) & (g849) & (g844)) + ((g839) & (!g840) & (g843) & (g842) & (!g849) & (!g844)) + ((g839) & (g840) & (!g843) & (!g842) & (g849) & (g844)) + ((g839) & (g840) & (!g843) & (g842) & (!g849) & (!g844)) + ((g839) & (g840) & (!g843) & (g842) & (!g849) & (g844)) + ((g839) & (g840) & (g843) & (!g842) & (g849) & (g844)));
	assign g886 = (((!g882) & (!g883) & (!g884) & (!g885) & (!g850) & (!g841)) + ((!g882) & (!g883) & (!g884) & (!g885) & (!g850) & (g841)) + ((!g882) & (!g883) & (!g884) & (!g885) & (g850) & (!g841)) + ((!g882) & (!g883) & (!g884) & (g885) & (!g850) & (!g841)) + ((!g882) & (!g883) & (!g884) & (g885) & (!g850) & (g841)) + ((!g882) & (!g883) & (!g884) & (g885) & (g850) & (!g841)) + ((!g882) & (!g883) & (!g884) & (g885) & (g850) & (g841)) + ((!g882) & (!g883) & (g884) & (!g885) & (!g850) & (!g841)) + ((!g882) & (!g883) & (g884) & (!g885) & (g850) & (!g841)) + ((!g882) & (!g883) & (g884) & (g885) & (!g850) & (!g841)) + ((!g882) & (!g883) & (g884) & (g885) & (g850) & (!g841)) + ((!g882) & (!g883) & (g884) & (g885) & (g850) & (g841)) + ((!g882) & (g883) & (!g884) & (!g885) & (!g850) & (!g841)) + ((!g882) & (g883) & (!g884) & (!g885) & (!g850) & (g841)) + ((!g882) & (g883) & (!g884) & (g885) & (!g850) & (!g841)) + ((!g882) & (g883) & (!g884) & (g885) & (!g850) & (g841)) + ((!g882) & (g883) & (!g884) & (g885) & (g850) & (g841)) + ((!g882) & (g883) & (g884) & (!g885) & (!g850) & (!g841)) + ((!g882) & (g883) & (g884) & (g885) & (!g850) & (!g841)) + ((!g882) & (g883) & (g884) & (g885) & (g850) & (g841)) + ((g882) & (!g883) & (!g884) & (!g885) & (!g850) & (g841)) + ((g882) & (!g883) & (!g884) & (!g885) & (g850) & (!g841)) + ((g882) & (!g883) & (!g884) & (g885) & (!g850) & (g841)) + ((g882) & (!g883) & (!g884) & (g885) & (g850) & (!g841)) + ((g882) & (!g883) & (!g884) & (g885) & (g850) & (g841)) + ((g882) & (!g883) & (g884) & (!g885) & (g850) & (!g841)) + ((g882) & (!g883) & (g884) & (g885) & (g850) & (!g841)) + ((g882) & (!g883) & (g884) & (g885) & (g850) & (g841)) + ((g882) & (g883) & (!g884) & (!g885) & (!g850) & (g841)) + ((g882) & (g883) & (!g884) & (g885) & (!g850) & (g841)) + ((g882) & (g883) & (!g884) & (g885) & (g850) & (g841)) + ((g882) & (g883) & (g884) & (g885) & (g850) & (g841)));
	assign g888 = (((!sk[52]) & (g886) & (!g887)) + ((!sk[52]) & (g886) & (g887)) + ((sk[52]) & (!g886) & (g887)) + ((sk[52]) & (g886) & (!g887)));
	assign g889 = (((!g839) & (!g850) & (!g841) & (!g842) & (!g849) & (g844)) + ((!g839) & (!g850) & (!g841) & (!g842) & (g849) & (g844)) + ((!g839) & (!g850) & (!g841) & (g842) & (!g849) & (!g844)) + ((!g839) & (!g850) & (!g841) & (g842) & (!g849) & (g844)) + ((!g839) & (!g850) & (!g841) & (g842) & (g849) & (!g844)) + ((!g839) & (!g850) & (!g841) & (g842) & (g849) & (g844)) + ((!g839) & (!g850) & (g841) & (!g842) & (!g849) & (g844)) + ((!g839) & (!g850) & (g841) & (!g842) & (g849) & (g844)) + ((!g839) & (!g850) & (g841) & (g842) & (g849) & (!g844)) + ((!g839) & (g850) & (g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (g850) & (g841) & (!g842) & (g849) & (g844)) + ((!g839) & (g850) & (g841) & (g842) & (!g849) & (g844)) + ((g839) & (!g850) & (!g841) & (!g842) & (g849) & (!g844)) + ((g839) & (!g850) & (!g841) & (g842) & (!g849) & (!g844)) + ((g839) & (!g850) & (!g841) & (g842) & (!g849) & (g844)) + ((g839) & (!g850) & (!g841) & (g842) & (g849) & (g844)) + ((g839) & (!g850) & (g841) & (!g842) & (!g849) & (g844)) + ((g839) & (!g850) & (g841) & (!g842) & (g849) & (g844)) + ((g839) & (!g850) & (g841) & (g842) & (g849) & (!g844)) + ((g839) & (!g850) & (g841) & (g842) & (g849) & (g844)) + ((g839) & (g850) & (!g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (g850) & (!g841) & (!g842) & (!g849) & (g844)) + ((g839) & (g850) & (!g841) & (!g842) & (g849) & (!g844)) + ((g839) & (g850) & (!g841) & (g842) & (!g849) & (!g844)) + ((g839) & (g850) & (g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (g850) & (g841) & (!g842) & (!g849) & (g844)) + ((g839) & (g850) & (g841) & (!g842) & (g849) & (!g844)) + ((g839) & (g850) & (g841) & (g842) & (!g849) & (g844)));
	assign g890 = (((!g839) & (!g850) & (!g841) & (!g842) & (!g849) & (!g844)) + ((!g839) & (!g850) & (!g841) & (g842) & (g849) & (g844)) + ((!g839) & (!g850) & (g841) & (!g842) & (!g849) & (!g844)) + ((!g839) & (!g850) & (g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (!g850) & (g841) & (!g842) & (g849) & (g844)) + ((!g839) & (!g850) & (g841) & (g842) & (!g849) & (!g844)) + ((!g839) & (!g850) & (g841) & (g842) & (g849) & (g844)) + ((!g839) & (g850) & (!g841) & (!g842) & (!g849) & (!g844)) + ((!g839) & (g850) & (!g841) & (!g842) & (g849) & (g844)) + ((!g839) & (g850) & (!g841) & (g842) & (!g849) & (g844)) + ((!g839) & (g850) & (g841) & (!g842) & (!g849) & (!g844)) + ((!g839) & (g850) & (g841) & (!g842) & (g849) & (g844)) + ((!g839) & (g850) & (g841) & (g842) & (g849) & (!g844)) + ((!g839) & (g850) & (g841) & (g842) & (g849) & (g844)) + ((g839) & (!g850) & (!g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (!g850) & (!g841) & (!g842) & (g849) & (g844)) + ((g839) & (!g850) & (!g841) & (g842) & (!g849) & (!g844)) + ((g839) & (!g850) & (!g841) & (g842) & (g849) & (g844)) + ((g839) & (!g850) & (g841) & (!g842) & (g849) & (g844)) + ((g839) & (!g850) & (g841) & (g842) & (!g849) & (g844)) + ((g839) & (g850) & (!g841) & (!g842) & (g849) & (!g844)) + ((g839) & (g850) & (!g841) & (!g842) & (g849) & (g844)) + ((g839) & (g850) & (!g841) & (g842) & (!g849) & (g844)) + ((g839) & (g850) & (!g841) & (g842) & (g849) & (!g844)) + ((g839) & (g850) & (!g841) & (g842) & (g849) & (g844)) + ((g839) & (g850) & (g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (g850) & (g841) & (!g842) & (g849) & (!g844)) + ((g839) & (g850) & (g841) & (g842) & (!g849) & (!g844)));
	assign g891 = (((!g839) & (!g850) & (!g841) & (!g842) & (!g849) & (g844)) + ((!g839) & (!g850) & (!g841) & (!g842) & (g849) & (g844)) + ((!g839) & (!g850) & (!g841) & (g842) & (g849) & (!g844)) + ((!g839) & (!g850) & (!g841) & (g842) & (g849) & (g844)) + ((!g839) & (!g850) & (g841) & (!g842) & (g849) & (g844)) + ((!g839) & (!g850) & (g841) & (g842) & (!g849) & (!g844)) + ((!g839) & (!g850) & (g841) & (g842) & (!g849) & (g844)) + ((!g839) & (!g850) & (g841) & (g842) & (g849) & (g844)) + ((!g839) & (g850) & (!g841) & (!g842) & (!g849) & (!g844)) + ((!g839) & (g850) & (!g841) & (!g842) & (!g849) & (g844)) + ((!g839) & (g850) & (!g841) & (!g842) & (g849) & (g844)) + ((!g839) & (g850) & (!g841) & (g842) & (!g849) & (g844)) + ((!g839) & (g850) & (!g841) & (g842) & (g849) & (!g844)) + ((!g839) & (g850) & (g841) & (!g842) & (!g849) & (g844)) + ((!g839) & (g850) & (g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (g850) & (g841) & (g842) & (!g849) & (!g844)) + ((!g839) & (g850) & (g841) & (g842) & (g849) & (!g844)) + ((!g839) & (g850) & (g841) & (g842) & (g849) & (g844)) + ((g839) & (!g850) & (!g841) & (!g842) & (!g849) & (g844)) + ((g839) & (!g850) & (!g841) & (g842) & (!g849) & (!g844)) + ((g839) & (!g850) & (!g841) & (g842) & (g849) & (!g844)) + ((g839) & (!g850) & (g841) & (!g842) & (g849) & (g844)) + ((g839) & (!g850) & (g841) & (g842) & (!g849) & (g844)) + ((g839) & (g850) & (!g841) & (!g842) & (!g849) & (g844)) + ((g839) & (g850) & (!g841) & (g842) & (!g849) & (!g844)) + ((g839) & (g850) & (!g841) & (g842) & (g849) & (!g844)) + ((g839) & (g850) & (g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (g850) & (g841) & (!g842) & (g849) & (!g844)) + ((g839) & (g850) & (g841) & (!g842) & (g849) & (g844)) + ((g839) & (g850) & (g841) & (g842) & (g849) & (g844)));
	assign g892 = (((!g839) & (!g850) & (!g841) & (!g842) & (g849) & (g844)) + ((!g839) & (!g850) & (!g841) & (g842) & (!g849) & (!g844)) + ((!g839) & (!g850) & (!g841) & (g842) & (g849) & (g844)) + ((!g839) & (!g850) & (g841) & (!g842) & (!g849) & (!g844)) + ((!g839) & (!g850) & (g841) & (g842) & (g849) & (!g844)) + ((!g839) & (!g850) & (g841) & (g842) & (g849) & (g844)) + ((!g839) & (g850) & (!g841) & (g842) & (!g849) & (!g844)) + ((!g839) & (g850) & (!g841) & (g842) & (g849) & (!g844)) + ((!g839) & (g850) & (g841) & (!g842) & (g849) & (!g844)) + ((!g839) & (g850) & (g841) & (!g842) & (g849) & (g844)) + ((g839) & (!g850) & (!g841) & (!g842) & (!g849) & (g844)) + ((g839) & (!g850) & (!g841) & (!g842) & (g849) & (!g844)) + ((g839) & (!g850) & (!g841) & (g842) & (!g849) & (g844)) + ((g839) & (!g850) & (g841) & (!g842) & (g849) & (!g844)) + ((g839) & (!g850) & (g841) & (!g842) & (g849) & (g844)) + ((g839) & (!g850) & (g841) & (g842) & (g849) & (!g844)) + ((g839) & (!g850) & (g841) & (g842) & (g849) & (g844)) + ((g839) & (g850) & (!g841) & (!g842) & (g849) & (!g844)) + ((g839) & (g850) & (!g841) & (g842) & (!g849) & (g844)) + ((g839) & (g850) & (g841) & (!g842) & (!g849) & (!g844)) + ((g839) & (g850) & (g841) & (!g842) & (g849) & (g844)) + ((g839) & (g850) & (g841) & (g842) & (!g849) & (g844)));
	assign g893 = (((!g889) & (!g890) & (!g891) & (!g892) & (!g843) & (!g840)) + ((!g889) & (!g890) & (!g891) & (!g892) & (!g843) & (g840)) + ((!g889) & (!g890) & (!g891) & (!g892) & (g843) & (!g840)) + ((!g889) & (!g890) & (!g891) & (g892) & (!g843) & (!g840)) + ((!g889) & (!g890) & (!g891) & (g892) & (!g843) & (g840)) + ((!g889) & (!g890) & (!g891) & (g892) & (g843) & (!g840)) + ((!g889) & (!g890) & (!g891) & (g892) & (g843) & (g840)) + ((!g889) & (!g890) & (g891) & (!g892) & (!g843) & (!g840)) + ((!g889) & (!g890) & (g891) & (!g892) & (g843) & (!g840)) + ((!g889) & (!g890) & (g891) & (g892) & (!g843) & (!g840)) + ((!g889) & (!g890) & (g891) & (g892) & (g843) & (!g840)) + ((!g889) & (!g890) & (g891) & (g892) & (g843) & (g840)) + ((!g889) & (g890) & (!g891) & (!g892) & (!g843) & (!g840)) + ((!g889) & (g890) & (!g891) & (!g892) & (!g843) & (g840)) + ((!g889) & (g890) & (!g891) & (g892) & (!g843) & (!g840)) + ((!g889) & (g890) & (!g891) & (g892) & (!g843) & (g840)) + ((!g889) & (g890) & (!g891) & (g892) & (g843) & (g840)) + ((!g889) & (g890) & (g891) & (!g892) & (!g843) & (!g840)) + ((!g889) & (g890) & (g891) & (g892) & (!g843) & (!g840)) + ((!g889) & (g890) & (g891) & (g892) & (g843) & (g840)) + ((g889) & (!g890) & (!g891) & (!g892) & (!g843) & (g840)) + ((g889) & (!g890) & (!g891) & (!g892) & (g843) & (!g840)) + ((g889) & (!g890) & (!g891) & (g892) & (!g843) & (g840)) + ((g889) & (!g890) & (!g891) & (g892) & (g843) & (!g840)) + ((g889) & (!g890) & (!g891) & (g892) & (g843) & (g840)) + ((g889) & (!g890) & (g891) & (!g892) & (g843) & (!g840)) + ((g889) & (!g890) & (g891) & (g892) & (g843) & (!g840)) + ((g889) & (!g890) & (g891) & (g892) & (g843) & (g840)) + ((g889) & (g890) & (!g891) & (!g892) & (!g843) & (g840)) + ((g889) & (g890) & (!g891) & (g892) & (!g843) & (g840)) + ((g889) & (g890) & (!g891) & (g892) & (g843) & (g840)) + ((g889) & (g890) & (g891) & (g892) & (g843) & (g840)));
	assign g895 = (((!sk[58]) & (g893) & (!g894)) + ((!sk[58]) & (g893) & (g894)) + ((sk[58]) & (!g893) & (g894)) + ((sk[58]) & (g893) & (!g894)));
	assign g896 = (((!g843) & (!g840) & (!g841) & (!g842) & (!g849) & (g850)) + ((!g843) & (!g840) & (!g841) & (!g842) & (g849) & (!g850)) + ((!g843) & (!g840) & (!g841) & (g842) & (!g849) & (g850)) + ((!g843) & (!g840) & (!g841) & (g842) & (g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (!g842) & (!g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (!g842) & (g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (g842) & (!g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (g842) & (g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (g842) & (g849) & (g850)) + ((!g843) & (g840) & (!g841) & (!g842) & (g849) & (!g850)) + ((!g843) & (g840) & (!g841) & (g842) & (g849) & (!g850)) + ((!g843) & (g840) & (!g841) & (g842) & (g849) & (g850)) + ((!g843) & (g840) & (g841) & (!g842) & (g849) & (g850)) + ((!g843) & (g840) & (g841) & (g842) & (!g849) & (!g850)) + ((g843) & (!g840) & (!g841) & (!g842) & (!g849) & (g850)) + ((g843) & (!g840) & (!g841) & (g842) & (!g849) & (g850)) + ((g843) & (!g840) & (g841) & (g842) & (g849) & (g850)) + ((g843) & (g840) & (!g841) & (!g842) & (g849) & (g850)) + ((g843) & (g840) & (!g841) & (g842) & (!g849) & (!g850)) + ((g843) & (g840) & (!g841) & (g842) & (g849) & (!g850)) + ((g843) & (g840) & (g841) & (!g842) & (!g849) & (g850)) + ((g843) & (g840) & (g841) & (!g842) & (g849) & (!g850)) + ((g843) & (g840) & (g841) & (!g842) & (g849) & (g850)) + ((g843) & (g840) & (g841) & (g842) & (!g849) & (g850)));
	assign g897 = (((!g843) & (!g840) & (!g841) & (!g842) & (!g849) & (!g850)) + ((!g843) & (!g840) & (!g841) & (!g842) & (!g849) & (g850)) + ((!g843) & (!g840) & (!g841) & (g842) & (!g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (!g842) & (!g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (!g842) & (g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (!g842) & (g849) & (g850)) + ((!g843) & (!g840) & (g841) & (g842) & (!g849) & (g850)) + ((!g843) & (!g840) & (g841) & (g842) & (g849) & (g850)) + ((!g843) & (g840) & (!g841) & (!g842) & (!g849) & (!g850)) + ((!g843) & (g840) & (!g841) & (!g842) & (g849) & (!g850)) + ((!g843) & (g840) & (!g841) & (g842) & (!g849) & (!g850)) + ((!g843) & (g840) & (!g841) & (g842) & (!g849) & (g850)) + ((!g843) & (g840) & (!g841) & (g842) & (g849) & (g850)) + ((!g843) & (g840) & (g841) & (!g842) & (!g849) & (g850)) + ((!g843) & (g840) & (g841) & (g842) & (!g849) & (!g850)) + ((!g843) & (g840) & (g841) & (g842) & (!g849) & (g850)) + ((g843) & (!g840) & (!g841) & (!g842) & (!g849) & (g850)) + ((g843) & (!g840) & (!g841) & (!g842) & (g849) & (g850)) + ((g843) & (!g840) & (!g841) & (g842) & (!g849) & (!g850)) + ((g843) & (!g840) & (!g841) & (g842) & (g849) & (g850)) + ((g843) & (!g840) & (g841) & (!g842) & (!g849) & (!g850)) + ((g843) & (!g840) & (g841) & (!g842) & (g849) & (g850)) + ((g843) & (!g840) & (g841) & (g842) & (g849) & (!g850)) + ((g843) & (g840) & (!g841) & (!g842) & (!g849) & (!g850)) + ((g843) & (g840) & (!g841) & (!g842) & (!g849) & (g850)) + ((g843) & (g840) & (!g841) & (!g842) & (g849) & (g850)) + ((g843) & (g840) & (!g841) & (g842) & (!g849) & (g850)) + ((g843) & (g840) & (!g841) & (g842) & (g849) & (!g850)) + ((g843) & (g840) & (g841) & (!g842) & (g849) & (!g850)) + ((g843) & (g840) & (g841) & (!g842) & (g849) & (g850)));
	assign g898 = (((!g843) & (!g840) & (!g841) & (!g842) & (g849) & (!g850)) + ((!g843) & (!g840) & (!g841) & (g842) & (!g849) & (!g850)) + ((!g843) & (!g840) & (!g841) & (g842) & (g849) & (!g850)) + ((!g843) & (!g840) & (!g841) & (g842) & (g849) & (g850)) + ((!g843) & (!g840) & (g841) & (!g842) & (!g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (!g842) & (!g849) & (g850)) + ((!g843) & (!g840) & (g841) & (!g842) & (g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (g842) & (!g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (g842) & (g849) & (g850)) + ((!g843) & (g840) & (!g841) & (!g842) & (!g849) & (g850)) + ((!g843) & (g840) & (!g841) & (!g842) & (g849) & (!g850)) + ((!g843) & (g840) & (!g841) & (!g842) & (g849) & (g850)) + ((!g843) & (g840) & (g841) & (!g842) & (!g849) & (g850)) + ((!g843) & (g840) & (g841) & (!g842) & (g849) & (!g850)) + ((!g843) & (g840) & (g841) & (!g842) & (g849) & (g850)) + ((!g843) & (g840) & (g841) & (g842) & (!g849) & (!g850)) + ((g843) & (!g840) & (!g841) & (!g842) & (g849) & (!g850)) + ((g843) & (!g840) & (!g841) & (g842) & (!g849) & (!g850)) + ((g843) & (!g840) & (!g841) & (g842) & (g849) & (g850)) + ((g843) & (!g840) & (g841) & (!g842) & (!g849) & (!g850)) + ((g843) & (!g840) & (g841) & (!g842) & (!g849) & (g850)) + ((g843) & (!g840) & (g841) & (g842) & (!g849) & (!g850)) + ((g843) & (!g840) & (g841) & (g842) & (g849) & (!g850)) + ((g843) & (g840) & (!g841) & (!g842) & (g849) & (!g850)) + ((g843) & (g840) & (!g841) & (g842) & (!g849) & (!g850)) + ((g843) & (g840) & (!g841) & (g842) & (g849) & (g850)) + ((g843) & (g840) & (g841) & (!g842) & (!g849) & (!g850)) + ((g843) & (g840) & (g841) & (!g842) & (g849) & (!g850)) + ((g843) & (g840) & (g841) & (!g842) & (g849) & (g850)) + ((g843) & (g840) & (g841) & (g842) & (!g849) & (g850)));
	assign g899 = (((!g843) & (!g840) & (!g841) & (!g842) & (!g849) & (g850)) + ((!g843) & (!g840) & (!g841) & (g842) & (g849) & (!g850)) + ((!g843) & (!g840) & (!g841) & (g842) & (g849) & (g850)) + ((!g843) & (!g840) & (g841) & (!g842) & (!g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (!g842) & (!g849) & (g850)) + ((!g843) & (!g840) & (g841) & (g842) & (g849) & (!g850)) + ((!g843) & (!g840) & (g841) & (g842) & (g849) & (g850)) + ((!g843) & (g840) & (!g841) & (!g842) & (!g849) & (!g850)) + ((!g843) & (g840) & (!g841) & (!g842) & (!g849) & (g850)) + ((!g843) & (g840) & (!g841) & (!g842) & (g849) & (g850)) + ((!g843) & (g840) & (!g841) & (g842) & (!g849) & (g850)) + ((!g843) & (g840) & (g841) & (!g842) & (!g849) & (g850)) + ((!g843) & (g840) & (g841) & (g842) & (!g849) & (!g850)) + ((!g843) & (g840) & (g841) & (g842) & (!g849) & (g850)) + ((!g843) & (g840) & (g841) & (g842) & (g849) & (!g850)) + ((!g843) & (g840) & (g841) & (g842) & (g849) & (g850)) + ((g843) & (!g840) & (!g841) & (g842) & (!g849) & (g850)) + ((g843) & (!g840) & (g841) & (!g842) & (!g849) & (!g850)) + ((g843) & (!g840) & (g841) & (g842) & (!g849) & (!g850)) + ((g843) & (!g840) & (g841) & (g842) & (!g849) & (g850)) + ((g843) & (!g840) & (g841) & (g842) & (g849) & (g850)) + ((g843) & (g840) & (!g841) & (!g842) & (!g849) & (g850)) + ((g843) & (g840) & (!g841) & (!g842) & (g849) & (g850)) + ((g843) & (g840) & (!g841) & (g842) & (!g849) & (!g850)) + ((g843) & (g840) & (!g841) & (g842) & (g849) & (!g850)) + ((g843) & (g840) & (!g841) & (g842) & (g849) & (g850)) + ((g843) & (g840) & (g841) & (!g842) & (g849) & (g850)) + ((g843) & (g840) & (g841) & (g842) & (g849) & (g850)));
	assign g900 = (((!g896) & (!g897) & (!g898) & (!g899) & (!g839) & (g844)) + ((!g896) & (!g897) & (!g898) & (!g899) & (g839) & (!g844)) + ((!g896) & (!g897) & (!g898) & (!g899) & (g839) & (g844)) + ((!g896) & (!g897) & (!g898) & (g899) & (!g839) & (g844)) + ((!g896) & (!g897) & (!g898) & (g899) & (g839) & (!g844)) + ((!g896) & (!g897) & (g898) & (!g899) & (g839) & (!g844)) + ((!g896) & (!g897) & (g898) & (!g899) & (g839) & (g844)) + ((!g896) & (!g897) & (g898) & (g899) & (g839) & (!g844)) + ((!g896) & (g897) & (!g898) & (!g899) & (!g839) & (g844)) + ((!g896) & (g897) & (!g898) & (!g899) & (g839) & (g844)) + ((!g896) & (g897) & (!g898) & (g899) & (!g839) & (g844)) + ((!g896) & (g897) & (g898) & (!g899) & (g839) & (g844)) + ((g896) & (!g897) & (!g898) & (!g899) & (!g839) & (!g844)) + ((g896) & (!g897) & (!g898) & (!g899) & (!g839) & (g844)) + ((g896) & (!g897) & (!g898) & (!g899) & (g839) & (!g844)) + ((g896) & (!g897) & (!g898) & (!g899) & (g839) & (g844)) + ((g896) & (!g897) & (!g898) & (g899) & (!g839) & (!g844)) + ((g896) & (!g897) & (!g898) & (g899) & (!g839) & (g844)) + ((g896) & (!g897) & (!g898) & (g899) & (g839) & (!g844)) + ((g896) & (!g897) & (g898) & (!g899) & (!g839) & (!g844)) + ((g896) & (!g897) & (g898) & (!g899) & (g839) & (!g844)) + ((g896) & (!g897) & (g898) & (!g899) & (g839) & (g844)) + ((g896) & (!g897) & (g898) & (g899) & (!g839) & (!g844)) + ((g896) & (!g897) & (g898) & (g899) & (g839) & (!g844)) + ((g896) & (g897) & (!g898) & (!g899) & (!g839) & (!g844)) + ((g896) & (g897) & (!g898) & (!g899) & (!g839) & (g844)) + ((g896) & (g897) & (!g898) & (!g899) & (g839) & (g844)) + ((g896) & (g897) & (!g898) & (g899) & (!g839) & (!g844)) + ((g896) & (g897) & (!g898) & (g899) & (!g839) & (g844)) + ((g896) & (g897) & (g898) & (!g899) & (!g839) & (!g844)) + ((g896) & (g897) & (g898) & (!g899) & (g839) & (g844)) + ((g896) & (g897) & (g898) & (g899) & (!g839) & (!g844)));
	assign g902 = (((!sk[64]) & (g900) & (!g901)) + ((!sk[64]) & (g900) & (g901)) + ((sk[64]) & (!g900) & (g901)) + ((sk[64]) & (g900) & (!g901)));
	assign g909 = (((!g903) & (!g904) & (!g905) & (!g906) & (g907) & (g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g907) & (!g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g907) & (g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (g907) & (!g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (!g907) & (!g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (!g907) & (g908)) + ((!g903) & (!g904) & (g905) & (g906) & (!g907) & (!g908)) + ((!g903) & (!g904) & (g905) & (g906) & (g907) & (g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (g907) & (!g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (g907) & (g908)) + ((!g903) & (g904) & (!g905) & (g906) & (g907) & (!g908)) + ((!g903) & (g904) & (!g905) & (g906) & (g907) & (g908)) + ((!g903) & (g904) & (g905) & (!g906) & (g907) & (!g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (!g907) & (!g908)) + ((g903) & (!g904) & (g905) & (!g906) & (g907) & (!g908)) + ((g903) & (!g904) & (g905) & (g906) & (!g907) & (g908)) + ((g903) & (!g904) & (g905) & (g906) & (g907) & (g908)) + ((g903) & (g904) & (!g905) & (!g906) & (!g907) & (g908)) + ((g903) & (g904) & (!g905) & (!g906) & (g907) & (!g908)) + ((g903) & (g904) & (g905) & (!g906) & (!g907) & (g908)) + ((g903) & (g904) & (g905) & (!g906) & (g907) & (!g908)) + ((g903) & (g904) & (g905) & (g906) & (!g907) & (!g908)) + ((g903) & (g904) & (g905) & (g906) & (g907) & (!g908)) + ((g903) & (g904) & (g905) & (g906) & (g907) & (g908)));
	assign g910 = (((!g903) & (!g904) & (!g905) & (!g906) & (g907) & (!g908)) + ((!g903) & (!g904) & (!g905) & (!g906) & (g907) & (g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g907) & (!g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g907) & (g908)) + ((!g903) & (!g904) & (g905) & (g906) & (!g907) & (g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (!g907) & (!g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (!g907) & (g908)) + ((!g903) & (g904) & (g905) & (!g906) & (!g907) & (!g908)) + ((!g903) & (g904) & (g905) & (!g906) & (!g907) & (g908)) + ((!g903) & (g904) & (g905) & (!g906) & (g907) & (!g908)) + ((!g903) & (g904) & (g905) & (g906) & (g907) & (g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (!g907) & (g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (g907) & (!g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (g907) & (g908)) + ((g903) & (!g904) & (!g905) & (g906) & (g907) & (!g908)) + ((g903) & (!g904) & (g905) & (!g906) & (!g907) & (!g908)) + ((g903) & (!g904) & (g905) & (!g906) & (g907) & (g908)) + ((g903) & (!g904) & (g905) & (g906) & (!g907) & (g908)) + ((g903) & (!g904) & (g905) & (g906) & (g907) & (g908)) + ((g903) & (g904) & (!g905) & (!g906) & (!g907) & (!g908)) + ((g903) & (g904) & (!g905) & (!g906) & (!g907) & (g908)) + ((g903) & (g904) & (!g905) & (!g906) & (g907) & (!g908)) + ((g903) & (g904) & (!g905) & (!g906) & (g907) & (g908)) + ((g903) & (g904) & (!g905) & (g906) & (!g907) & (!g908)) + ((g903) & (g904) & (!g905) & (g906) & (g907) & (!g908)) + ((g903) & (g904) & (!g905) & (g906) & (g907) & (g908)) + ((g903) & (g904) & (g905) & (!g906) & (g907) & (!g908)) + ((g903) & (g904) & (g905) & (!g906) & (g907) & (g908)) + ((g903) & (g904) & (g905) & (g906) & (!g907) & (g908)) + ((g903) & (g904) & (g905) & (g906) & (g907) & (!g908)));
	assign g911 = (((!g903) & (!g904) & (!g905) & (!g906) & (!g907) & (!g908)) + ((!g903) & (!g904) & (!g905) & (!g906) & (g907) & (g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (g907) & (g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (!g907) & (!g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (!g907) & (g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (g907) & (g908)) + ((!g903) & (!g904) & (g905) & (g906) & (!g907) & (g908)) + ((!g903) & (!g904) & (g905) & (g906) & (g907) & (!g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (!g907) & (!g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (g907) & (!g908)) + ((!g903) & (g904) & (!g905) & (g906) & (g907) & (g908)) + ((!g903) & (g904) & (g905) & (g906) & (!g907) & (!g908)) + ((!g903) & (g904) & (g905) & (g906) & (g907) & (!g908)) + ((g903) & (!g904) & (!g905) & (g906) & (!g907) & (!g908)) + ((g903) & (!g904) & (!g905) & (g906) & (!g907) & (g908)) + ((g903) & (!g904) & (!g905) & (g906) & (g907) & (!g908)) + ((g903) & (!g904) & (g905) & (!g906) & (!g907) & (!g908)) + ((g903) & (!g904) & (g905) & (!g906) & (g907) & (g908)) + ((g903) & (!g904) & (g905) & (g906) & (!g907) & (!g908)) + ((g903) & (!g904) & (g905) & (g906) & (!g907) & (g908)) + ((g903) & (!g904) & (g905) & (g906) & (g907) & (!g908)) + ((g903) & (!g904) & (g905) & (g906) & (g907) & (g908)) + ((g903) & (g904) & (!g905) & (!g906) & (g907) & (g908)) + ((g903) & (g904) & (!g905) & (g906) & (!g907) & (!g908)) + ((g903) & (g904) & (!g905) & (g906) & (g907) & (!g908)) + ((g903) & (g904) & (!g905) & (g906) & (g907) & (g908)) + ((g903) & (g904) & (g905) & (!g906) & (!g907) & (!g908)) + ((g903) & (g904) & (g905) & (g906) & (!g907) & (!g908)) + ((g903) & (g904) & (g905) & (g906) & (!g907) & (g908)) + ((g903) & (g904) & (g905) & (g906) & (g907) & (g908)));
	assign g912 = (((!g903) & (!g904) & (!g905) & (!g906) & (!g907) & (g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (g907) & (!g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (g907) & (g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (!g907) & (g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (g907) & (g908)) + ((!g903) & (!g904) & (g905) & (g906) & (!g907) & (g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (!g907) & (!g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (!g907) & (g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (g907) & (!g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (g907) & (g908)) + ((!g903) & (g904) & (!g905) & (g906) & (g907) & (!g908)) + ((!g903) & (g904) & (!g905) & (g906) & (g907) & (g908)) + ((!g903) & (g904) & (g905) & (g906) & (!g907) & (!g908)) + ((!g903) & (g904) & (g905) & (g906) & (g907) & (!g908)) + ((!g903) & (g904) & (g905) & (g906) & (g907) & (g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (!g907) & (!g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (g907) & (g908)) + ((g903) & (!g904) & (!g905) & (g906) & (g907) & (!g908)) + ((g903) & (!g904) & (!g905) & (g906) & (g907) & (g908)) + ((g903) & (!g904) & (g905) & (!g906) & (!g907) & (g908)) + ((g903) & (!g904) & (g905) & (!g906) & (g907) & (!g908)) + ((g903) & (!g904) & (g905) & (g906) & (g907) & (!g908)) + ((g903) & (g904) & (!g905) & (!g906) & (!g907) & (g908)) + ((g903) & (g904) & (!g905) & (!g906) & (g907) & (g908)) + ((g903) & (g904) & (!g905) & (g906) & (g907) & (!g908)) + ((g903) & (g904) & (!g905) & (g906) & (g907) & (g908)) + ((g903) & (g904) & (g905) & (!g906) & (!g907) & (g908)) + ((g903) & (g904) & (g905) & (g906) & (!g907) & (!g908)));
	assign g915 = (((!g909) & (!g910) & (!g911) & (!g912) & (!g913) & (!g914)) + ((!g909) & (!g910) & (!g911) & (g912) & (!g913) & (!g914)) + ((!g909) & (!g910) & (!g911) & (g912) & (g913) & (g914)) + ((!g909) & (!g910) & (g911) & (!g912) & (!g913) & (!g914)) + ((!g909) & (!g910) & (g911) & (!g912) & (!g913) & (g914)) + ((!g909) & (!g910) & (g911) & (g912) & (!g913) & (!g914)) + ((!g909) & (!g910) & (g911) & (g912) & (!g913) & (g914)) + ((!g909) & (!g910) & (g911) & (g912) & (g913) & (g914)) + ((!g909) & (g910) & (!g911) & (!g912) & (!g913) & (!g914)) + ((!g909) & (g910) & (!g911) & (!g912) & (g913) & (!g914)) + ((!g909) & (g910) & (!g911) & (g912) & (!g913) & (!g914)) + ((!g909) & (g910) & (!g911) & (g912) & (g913) & (!g914)) + ((!g909) & (g910) & (!g911) & (g912) & (g913) & (g914)) + ((!g909) & (g910) & (g911) & (!g912) & (!g913) & (!g914)) + ((!g909) & (g910) & (g911) & (!g912) & (!g913) & (g914)) + ((!g909) & (g910) & (g911) & (!g912) & (g913) & (!g914)) + ((!g909) & (g910) & (g911) & (g912) & (!g913) & (!g914)) + ((!g909) & (g910) & (g911) & (g912) & (!g913) & (g914)) + ((!g909) & (g910) & (g911) & (g912) & (g913) & (!g914)) + ((!g909) & (g910) & (g911) & (g912) & (g913) & (g914)) + ((g909) & (!g910) & (!g911) & (g912) & (g913) & (g914)) + ((g909) & (!g910) & (g911) & (!g912) & (!g913) & (g914)) + ((g909) & (!g910) & (g911) & (g912) & (!g913) & (g914)) + ((g909) & (!g910) & (g911) & (g912) & (g913) & (g914)) + ((g909) & (g910) & (!g911) & (!g912) & (g913) & (!g914)) + ((g909) & (g910) & (!g911) & (g912) & (g913) & (!g914)) + ((g909) & (g910) & (!g911) & (g912) & (g913) & (g914)) + ((g909) & (g910) & (g911) & (!g912) & (!g913) & (g914)) + ((g909) & (g910) & (g911) & (!g912) & (g913) & (!g914)) + ((g909) & (g910) & (g911) & (g912) & (!g913) & (g914)) + ((g909) & (g910) & (g911) & (g912) & (g913) & (!g914)) + ((g909) & (g910) & (g911) & (g912) & (g913) & (g914)));
	assign g917 = (((!g915) & (sk[70]) & (g916)) + ((g915) & (!sk[70]) & (!g916)) + ((g915) & (!sk[70]) & (g916)) + ((g915) & (sk[70]) & (!g916)));
	assign g918 = (((!g903) & (!g904) & (!g905) & (!g906) & (!g913) & (g907)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g913) & (!g907)) + ((!g903) & (!g904) & (!g905) & (g906) & (g913) & (!g907)) + ((!g903) & (!g904) & (g905) & (!g906) & (g913) & (g907)) + ((!g903) & (!g904) & (g905) & (g906) & (!g913) & (g907)) + ((!g903) & (!g904) & (g905) & (g906) & (g913) & (!g907)) + ((!g903) & (g904) & (!g905) & (!g906) & (!g913) & (g907)) + ((!g903) & (g904) & (!g905) & (!g906) & (g913) & (!g907)) + ((!g903) & (g904) & (!g905) & (!g906) & (g913) & (g907)) + ((!g903) & (g904) & (g905) & (!g906) & (g913) & (g907)) + ((!g903) & (g904) & (g905) & (g906) & (g913) & (g907)) + ((g903) & (!g904) & (!g905) & (!g906) & (!g913) & (!g907)) + ((g903) & (!g904) & (!g905) & (!g906) & (g913) & (g907)) + ((g903) & (!g904) & (!g905) & (g906) & (!g913) & (!g907)) + ((g903) & (!g904) & (!g905) & (g906) & (g913) & (!g907)) + ((g903) & (!g904) & (g905) & (!g906) & (g913) & (!g907)) + ((g903) & (!g904) & (g905) & (!g906) & (g913) & (g907)) + ((g903) & (!g904) & (g905) & (g906) & (g913) & (!g907)) + ((g903) & (!g904) & (g905) & (g906) & (g913) & (g907)) + ((g903) & (g904) & (!g905) & (!g906) & (g913) & (!g907)) + ((g903) & (g904) & (!g905) & (!g906) & (g913) & (g907)) + ((g903) & (g904) & (!g905) & (g906) & (g913) & (g907)) + ((g903) & (g904) & (g905) & (!g906) & (!g913) & (!g907)) + ((g903) & (g904) & (g905) & (!g906) & (!g913) & (g907)) + ((g903) & (g904) & (g905) & (!g906) & (g913) & (!g907)) + ((g903) & (g904) & (g905) & (g906) & (!g913) & (g907)) + ((g903) & (g904) & (g905) & (g906) & (g913) & (!g907)));
	assign g919 = (((!g903) & (!g904) & (!g905) & (!g906) & (!g913) & (g907)) + ((!g903) & (!g904) & (!g905) & (!g906) & (g913) & (!g907)) + ((!g903) & (!g904) & (!g905) & (!g906) & (g913) & (g907)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g913) & (!g907)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g913) & (g907)) + ((!g903) & (!g904) & (!g905) & (g906) & (g913) & (g907)) + ((!g903) & (!g904) & (g905) & (!g906) & (g913) & (!g907)) + ((!g903) & (!g904) & (g905) & (g906) & (!g913) & (!g907)) + ((!g903) & (!g904) & (g905) & (g906) & (!g913) & (g907)) + ((!g903) & (!g904) & (g905) & (g906) & (g913) & (g907)) + ((!g903) & (g904) & (!g905) & (!g906) & (g913) & (g907)) + ((!g903) & (g904) & (!g905) & (g906) & (!g913) & (!g907)) + ((!g903) & (g904) & (!g905) & (g906) & (g913) & (!g907)) + ((!g903) & (g904) & (g905) & (!g906) & (g913) & (!g907)) + ((!g903) & (g904) & (g905) & (!g906) & (g913) & (g907)) + ((!g903) & (g904) & (g905) & (g906) & (!g913) & (!g907)) + ((g903) & (!g904) & (!g905) & (!g906) & (!g913) & (!g907)) + ((g903) & (!g904) & (!g905) & (g906) & (!g913) & (!g907)) + ((g903) & (!g904) & (!g905) & (g906) & (!g913) & (g907)) + ((g903) & (!g904) & (g905) & (!g906) & (!g913) & (g907)) + ((g903) & (!g904) & (g905) & (!g906) & (g913) & (g907)) + ((g903) & (!g904) & (g905) & (g906) & (!g913) & (!g907)) + ((g903) & (!g904) & (g905) & (g906) & (!g913) & (g907)) + ((g903) & (g904) & (!g905) & (g906) & (!g913) & (!g907)) + ((g903) & (g904) & (!g905) & (g906) & (g913) & (g907)) + ((g903) & (g904) & (g905) & (!g906) & (!g913) & (!g907)) + ((g903) & (g904) & (g905) & (!g906) & (!g913) & (g907)) + ((g903) & (g904) & (g905) & (!g906) & (g913) & (g907)) + ((g903) & (g904) & (g905) & (g906) & (!g913) & (!g907)) + ((g903) & (g904) & (g905) & (g906) & (!g913) & (g907)) + ((g903) & (g904) & (g905) & (g906) & (g913) & (!g907)));
	assign g920 = (((!g903) & (!g904) & (!g905) & (!g906) & (!g913) & (g907)) + ((!g903) & (!g904) & (!g905) & (g906) & (g913) & (!g907)) + ((!g903) & (!g904) & (g905) & (!g906) & (!g913) & (!g907)) + ((!g903) & (!g904) & (g905) & (!g906) & (g913) & (!g907)) + ((!g903) & (!g904) & (g905) & (g906) & (!g913) & (g907)) + ((!g903) & (!g904) & (g905) & (g906) & (g913) & (!g907)) + ((!g903) & (!g904) & (g905) & (g906) & (g913) & (g907)) + ((!g903) & (g904) & (!g905) & (!g906) & (!g913) & (!g907)) + ((!g903) & (g904) & (!g905) & (!g906) & (g913) & (!g907)) + ((!g903) & (g904) & (!g905) & (g906) & (!g913) & (!g907)) + ((!g903) & (g904) & (!g905) & (g906) & (g913) & (g907)) + ((!g903) & (g904) & (g905) & (!g906) & (g913) & (g907)) + ((!g903) & (g904) & (g905) & (g906) & (!g913) & (g907)) + ((!g903) & (g904) & (g905) & (g906) & (g913) & (!g907)) + ((g903) & (!g904) & (!g905) & (!g906) & (g913) & (g907)) + ((g903) & (!g904) & (!g905) & (g906) & (!g913) & (!g907)) + ((g903) & (!g904) & (!g905) & (g906) & (g913) & (!g907)) + ((g903) & (!g904) & (g905) & (!g906) & (!g913) & (!g907)) + ((g903) & (!g904) & (g905) & (!g906) & (!g913) & (g907)) + ((g903) & (!g904) & (g905) & (!g906) & (g913) & (!g907)) + ((g903) & (!g904) & (g905) & (!g906) & (g913) & (g907)) + ((g903) & (!g904) & (g905) & (g906) & (g913) & (!g907)) + ((g903) & (g904) & (!g905) & (!g906) & (!g913) & (g907)) + ((g903) & (g904) & (!g905) & (!g906) & (g913) & (g907)) + ((g903) & (g904) & (!g905) & (g906) & (!g913) & (g907)) + ((g903) & (g904) & (g905) & (!g906) & (!g913) & (!g907)) + ((g903) & (g904) & (g905) & (!g906) & (!g913) & (g907)) + ((g903) & (g904) & (g905) & (!g906) & (g913) & (g907)) + ((g903) & (g904) & (g905) & (g906) & (!g913) & (!g907)) + ((g903) & (g904) & (g905) & (g906) & (!g913) & (g907)) + ((g903) & (g904) & (g905) & (g906) & (g913) & (!g907)) + ((g903) & (g904) & (g905) & (g906) & (g913) & (g907)));
	assign g921 = (((!g903) & (!g904) & (!g905) & (!g906) & (g913) & (!g907)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g913) & (!g907)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g913) & (g907)) + ((!g903) & (!g904) & (g905) & (!g906) & (g913) & (g907)) + ((!g903) & (!g904) & (g905) & (g906) & (!g913) & (g907)) + ((!g903) & (g904) & (!g905) & (!g906) & (!g913) & (!g907)) + ((!g903) & (g904) & (!g905) & (!g906) & (g913) & (!g907)) + ((!g903) & (g904) & (!g905) & (g906) & (!g913) & (g907)) + ((!g903) & (g904) & (g905) & (!g906) & (!g913) & (g907)) + ((!g903) & (g904) & (g905) & (!g906) & (g913) & (!g907)) + ((!g903) & (g904) & (g905) & (!g906) & (g913) & (g907)) + ((!g903) & (g904) & (g905) & (g906) & (g913) & (!g907)) + ((!g903) & (g904) & (g905) & (g906) & (g913) & (g907)) + ((g903) & (!g904) & (!g905) & (!g906) & (!g913) & (!g907)) + ((g903) & (!g904) & (!g905) & (g906) & (!g913) & (!g907)) + ((g903) & (!g904) & (!g905) & (g906) & (!g913) & (g907)) + ((g903) & (!g904) & (!g905) & (g906) & (g913) & (!g907)) + ((g903) & (!g904) & (g905) & (!g906) & (!g913) & (!g907)) + ((g903) & (!g904) & (g905) & (!g906) & (g913) & (g907)) + ((g903) & (!g904) & (g905) & (g906) & (g913) & (!g907)) + ((g903) & (g904) & (!g905) & (!g906) & (!g913) & (!g907)) + ((g903) & (g904) & (!g905) & (g906) & (!g913) & (!g907)) + ((g903) & (g904) & (!g905) & (g906) & (g913) & (!g907)) + ((g903) & (g904) & (!g905) & (g906) & (g913) & (g907)) + ((g903) & (g904) & (g905) & (g906) & (!g913) & (g907)) + ((g903) & (g904) & (g905) & (g906) & (g913) & (g907)));
	assign g922 = (((!g918) & (!g919) & (!g920) & (!g921) & (!g908) & (!g914)) + ((!g918) & (!g919) & (!g920) & (!g921) & (g908) & (!g914)) + ((!g918) & (!g919) & (!g920) & (g921) & (!g908) & (!g914)) + ((!g918) & (!g919) & (!g920) & (g921) & (g908) & (!g914)) + ((!g918) & (!g919) & (!g920) & (g921) & (g908) & (g914)) + ((!g918) & (!g919) & (g920) & (!g921) & (!g908) & (!g914)) + ((!g918) & (!g919) & (g920) & (!g921) & (!g908) & (g914)) + ((!g918) & (!g919) & (g920) & (!g921) & (g908) & (!g914)) + ((!g918) & (!g919) & (g920) & (g921) & (!g908) & (!g914)) + ((!g918) & (!g919) & (g920) & (g921) & (!g908) & (g914)) + ((!g918) & (!g919) & (g920) & (g921) & (g908) & (!g914)) + ((!g918) & (!g919) & (g920) & (g921) & (g908) & (g914)) + ((!g918) & (g919) & (!g920) & (!g921) & (!g908) & (!g914)) + ((!g918) & (g919) & (!g920) & (g921) & (!g908) & (!g914)) + ((!g918) & (g919) & (!g920) & (g921) & (g908) & (g914)) + ((!g918) & (g919) & (g920) & (!g921) & (!g908) & (!g914)) + ((!g918) & (g919) & (g920) & (!g921) & (!g908) & (g914)) + ((!g918) & (g919) & (g920) & (g921) & (!g908) & (!g914)) + ((!g918) & (g919) & (g920) & (g921) & (!g908) & (g914)) + ((!g918) & (g919) & (g920) & (g921) & (g908) & (g914)) + ((g918) & (!g919) & (!g920) & (!g921) & (g908) & (!g914)) + ((g918) & (!g919) & (!g920) & (g921) & (g908) & (!g914)) + ((g918) & (!g919) & (!g920) & (g921) & (g908) & (g914)) + ((g918) & (!g919) & (g920) & (!g921) & (!g908) & (g914)) + ((g918) & (!g919) & (g920) & (!g921) & (g908) & (!g914)) + ((g918) & (!g919) & (g920) & (g921) & (!g908) & (g914)) + ((g918) & (!g919) & (g920) & (g921) & (g908) & (!g914)) + ((g918) & (!g919) & (g920) & (g921) & (g908) & (g914)) + ((g918) & (g919) & (!g920) & (g921) & (g908) & (g914)) + ((g918) & (g919) & (g920) & (!g921) & (!g908) & (g914)) + ((g918) & (g919) & (g920) & (g921) & (!g908) & (g914)) + ((g918) & (g919) & (g920) & (g921) & (g908) & (g914)));
	assign g924 = (((!g922) & (sk[76]) & (g923)) + ((g922) & (!sk[76]) & (!g923)) + ((g922) & (!sk[76]) & (g923)) + ((g922) & (sk[76]) & (!g923)));
	assign g925 = (((!g907) & (!g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((!g907) & (!g904) & (!g905) & (!g906) & (g913) & (g908)) + ((!g907) & (!g904) & (!g905) & (g906) & (!g913) & (g908)) + ((!g907) & (!g904) & (!g905) & (g906) & (g913) & (!g908)) + ((!g907) & (!g904) & (!g905) & (g906) & (g913) & (g908)) + ((!g907) & (!g904) & (g905) & (!g906) & (!g913) & (g908)) + ((!g907) & (!g904) & (g905) & (g906) & (!g913) & (!g908)) + ((!g907) & (!g904) & (g905) & (g906) & (g913) & (!g908)) + ((!g907) & (g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((!g907) & (g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((!g907) & (g904) & (!g905) & (g906) & (!g913) & (g908)) + ((!g907) & (g904) & (g905) & (!g906) & (!g913) & (!g908)) + ((!g907) & (g904) & (g905) & (!g906) & (!g913) & (g908)) + ((!g907) & (g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g907) & (g904) & (g905) & (!g906) & (g913) & (g908)) + ((g907) & (!g904) & (!g905) & (g906) & (!g913) & (g908)) + ((g907) & (!g904) & (!g905) & (g906) & (g913) & (g908)) + ((g907) & (g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((g907) & (g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((g907) & (g904) & (!g905) & (g906) & (g913) & (!g908)) + ((g907) & (g904) & (g905) & (g906) & (!g913) & (!g908)) + ((g907) & (g904) & (g905) & (g906) & (!g913) & (g908)));
	assign g926 = (((!g907) & (!g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((!g907) & (!g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((!g907) & (!g904) & (!g905) & (g906) & (g913) & (g908)) + ((!g907) & (!g904) & (g905) & (!g906) & (!g913) & (!g908)) + ((!g907) & (!g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g907) & (!g904) & (g905) & (g906) & (!g913) & (g908)) + ((!g907) & (g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((!g907) & (g904) & (!g905) & (!g906) & (g913) & (g908)) + ((!g907) & (g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((!g907) & (g904) & (!g905) & (g906) & (!g913) & (g908)) + ((!g907) & (g904) & (!g905) & (g906) & (g913) & (g908)) + ((!g907) & (g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g907) & (g904) & (g905) & (!g906) & (g913) & (g908)) + ((!g907) & (g904) & (g905) & (g906) & (g913) & (!g908)) + ((g907) & (!g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((g907) & (!g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((g907) & (!g904) & (!g905) & (!g906) & (g913) & (g908)) + ((g907) & (!g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((g907) & (!g904) & (!g905) & (g906) & (!g913) & (g908)) + ((g907) & (!g904) & (!g905) & (g906) & (g913) & (!g908)) + ((g907) & (!g904) & (g905) & (g906) & (!g913) & (!g908)) + ((g907) & (g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((g907) & (g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((g907) & (g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((g907) & (g904) & (!g905) & (g906) & (g913) & (!g908)) + ((g907) & (g904) & (!g905) & (g906) & (g913) & (g908)) + ((g907) & (g904) & (g905) & (!g906) & (!g913) & (!g908)) + ((g907) & (g904) & (g905) & (!g906) & (g913) & (!g908)) + ((g907) & (g904) & (g905) & (g906) & (!g913) & (g908)) + ((g907) & (g904) & (g905) & (g906) & (g913) & (g908)));
	assign g927 = (((!g907) & (!g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((!g907) & (!g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((!g907) & (!g904) & (!g905) & (g906) & (!g913) & (g908)) + ((!g907) & (!g904) & (g905) & (!g906) & (!g913) & (g908)) + ((!g907) & (!g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g907) & (!g904) & (g905) & (g906) & (!g913) & (g908)) + ((!g907) & (g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((!g907) & (g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((!g907) & (g904) & (!g905) & (g906) & (g913) & (!g908)) + ((!g907) & (g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g907) & (g904) & (g905) & (g906) & (!g913) & (!g908)) + ((!g907) & (g904) & (g905) & (g906) & (g913) & (!g908)) + ((g907) & (!g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((g907) & (!g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((g907) & (!g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((g907) & (!g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((g907) & (!g904) & (!g905) & (g906) & (!g913) & (g908)) + ((g907) & (!g904) & (!g905) & (g906) & (g913) & (!g908)) + ((g907) & (!g904) & (!g905) & (g906) & (g913) & (g908)) + ((g907) & (!g904) & (g905) & (!g906) & (!g913) & (g908)) + ((g907) & (!g904) & (g905) & (!g906) & (g913) & (!g908)) + ((g907) & (!g904) & (g905) & (g906) & (!g913) & (!g908)) + ((g907) & (!g904) & (g905) & (g906) & (g913) & (g908)) + ((g907) & (g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((g907) & (g904) & (!g905) & (!g906) & (g913) & (g908)) + ((g907) & (g904) & (g905) & (!g906) & (g913) & (g908)) + ((g907) & (g904) & (g905) & (g906) & (!g913) & (!g908)) + ((g907) & (g904) & (g905) & (g906) & (!g913) & (g908)) + ((g907) & (g904) & (g905) & (g906) & (g913) & (g908)));
	assign g928 = (((!g907) & (!g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((!g907) & (!g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((!g907) & (!g904) & (!g905) & (!g906) & (g913) & (g908)) + ((!g907) & (!g904) & (!g905) & (g906) & (!g913) & (g908)) + ((!g907) & (!g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g907) & (!g904) & (g905) & (g906) & (g913) & (g908)) + ((!g907) & (g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((!g907) & (g904) & (!g905) & (g906) & (!g913) & (g908)) + ((!g907) & (g904) & (!g905) & (g906) & (g913) & (g908)) + ((!g907) & (g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g907) & (g904) & (g905) & (!g906) & (g913) & (g908)) + ((!g907) & (g904) & (g905) & (g906) & (!g913) & (!g908)) + ((!g907) & (g904) & (g905) & (g906) & (!g913) & (g908)) + ((!g907) & (g904) & (g905) & (g906) & (g913) & (!g908)) + ((!g907) & (g904) & (g905) & (g906) & (g913) & (g908)) + ((g907) & (!g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((g907) & (!g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((g907) & (!g904) & (!g905) & (!g906) & (g913) & (g908)) + ((g907) & (!g904) & (!g905) & (g906) & (g913) & (g908)) + ((g907) & (!g904) & (g905) & (!g906) & (!g913) & (g908)) + ((g907) & (!g904) & (g905) & (!g906) & (g913) & (!g908)) + ((g907) & (!g904) & (g905) & (g906) & (g913) & (!g908)) + ((g907) & (g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((g907) & (g904) & (!g905) & (g906) & (!g913) & (g908)) + ((g907) & (g904) & (!g905) & (g906) & (g913) & (!g908)) + ((g907) & (g904) & (g905) & (!g906) & (g913) & (g908)) + ((g907) & (g904) & (g905) & (g906) & (!g913) & (!g908)));
	assign g929 = (((!g925) & (!g926) & (!g927) & (!g928) & (!g903) & (g914)) + ((!g925) & (!g926) & (!g927) & (!g928) & (g903) & (!g914)) + ((!g925) & (!g926) & (!g927) & (!g928) & (g903) & (g914)) + ((!g925) & (!g926) & (!g927) & (g928) & (!g903) & (g914)) + ((!g925) & (!g926) & (!g927) & (g928) & (g903) & (!g914)) + ((!g925) & (!g926) & (g927) & (!g928) & (g903) & (!g914)) + ((!g925) & (!g926) & (g927) & (!g928) & (g903) & (g914)) + ((!g925) & (!g926) & (g927) & (g928) & (g903) & (!g914)) + ((!g925) & (g926) & (!g927) & (!g928) & (!g903) & (g914)) + ((!g925) & (g926) & (!g927) & (!g928) & (g903) & (g914)) + ((!g925) & (g926) & (!g927) & (g928) & (!g903) & (g914)) + ((!g925) & (g926) & (g927) & (!g928) & (g903) & (g914)) + ((g925) & (!g926) & (!g927) & (!g928) & (!g903) & (!g914)) + ((g925) & (!g926) & (!g927) & (!g928) & (!g903) & (g914)) + ((g925) & (!g926) & (!g927) & (!g928) & (g903) & (!g914)) + ((g925) & (!g926) & (!g927) & (!g928) & (g903) & (g914)) + ((g925) & (!g926) & (!g927) & (g928) & (!g903) & (!g914)) + ((g925) & (!g926) & (!g927) & (g928) & (!g903) & (g914)) + ((g925) & (!g926) & (!g927) & (g928) & (g903) & (!g914)) + ((g925) & (!g926) & (g927) & (!g928) & (!g903) & (!g914)) + ((g925) & (!g926) & (g927) & (!g928) & (g903) & (!g914)) + ((g925) & (!g926) & (g927) & (!g928) & (g903) & (g914)) + ((g925) & (!g926) & (g927) & (g928) & (!g903) & (!g914)) + ((g925) & (!g926) & (g927) & (g928) & (g903) & (!g914)) + ((g925) & (g926) & (!g927) & (!g928) & (!g903) & (!g914)) + ((g925) & (g926) & (!g927) & (!g928) & (!g903) & (g914)) + ((g925) & (g926) & (!g927) & (!g928) & (g903) & (g914)) + ((g925) & (g926) & (!g927) & (g928) & (!g903) & (!g914)) + ((g925) & (g926) & (!g927) & (g928) & (!g903) & (g914)) + ((g925) & (g926) & (g927) & (!g928) & (!g903) & (!g914)) + ((g925) & (g926) & (g927) & (!g928) & (g903) & (g914)) + ((g925) & (g926) & (g927) & (g928) & (!g903) & (!g914)));
	assign g931 = (((!sk[82]) & (g929) & (!g930)) + ((!sk[82]) & (g929) & (g930)) + ((sk[82]) & (!g929) & (g930)) + ((sk[82]) & (g929) & (!g930)));
	assign g932 = (((!g903) & (!g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (g913) & (g908)) + ((!g903) & (!g904) & (g905) & (g906) & (!g913) & (!g908)) + ((!g903) & (!g904) & (g905) & (g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (g905) & (g906) & (g913) & (g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (g904) & (g905) & (!g906) & (!g913) & (!g908)) + ((!g903) & (g904) & (g905) & (g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((g903) & (!g904) & (g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (g905) & (!g906) & (!g913) & (g908)) + ((g903) & (!g904) & (g905) & (!g906) & (g913) & (!g908)) + ((g903) & (!g904) & (g905) & (g906) & (!g913) & (g908)) + ((g903) & (g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((g903) & (g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((g903) & (g904) & (!g905) & (g906) & (g913) & (!g908)) + ((g903) & (g904) & (g905) & (!g906) & (!g913) & (g908)) + ((g903) & (g904) & (g905) & (!g906) & (g913) & (g908)));
	assign g933 = (((!g903) & (!g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (!g905) & (!g906) & (g913) & (g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (g905) & (g906) & (!g913) & (!g908)) + ((!g903) & (!g904) & (g905) & (g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (g905) & (g906) & (g913) & (g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (g913) & (g908)) + ((!g903) & (g904) & (!g905) & (g906) & (g913) & (g908)) + ((!g903) & (g904) & (g905) & (!g906) & (!g913) & (!g908)) + ((!g903) & (g904) & (g905) & (!g906) & (!g913) & (g908)) + ((!g903) & (g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (g904) & (g905) & (g906) & (!g913) & (g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((g903) & (!g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (!g905) & (g906) & (!g913) & (g908)) + ((g903) & (!g904) & (!g905) & (g906) & (g913) & (g908)) + ((g903) & (!g904) & (g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (g905) & (!g906) & (!g913) & (g908)) + ((g903) & (!g904) & (g905) & (!g906) & (g913) & (g908)) + ((g903) & (!g904) & (g905) & (g906) & (!g913) & (g908)) + ((g903) & (g904) & (!g905) & (g906) & (!g913) & (g908)) + ((g903) & (g904) & (!g905) & (g906) & (g913) & (!g908)) + ((g903) & (g904) & (g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (g904) & (g905) & (g906) & (!g913) & (!g908)));
	assign g934 = (((!g903) & (!g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (!g905) & (!g906) & (g913) & (g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (g905) & (!g906) & (g913) & (g908)) + ((!g903) & (!g904) & (g905) & (g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (g905) & (g906) & (g913) & (g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (g913) & (g908)) + ((!g903) & (g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((!g903) & (g904) & (!g905) & (g906) & (!g913) & (g908)) + ((!g903) & (g904) & (g905) & (!g906) & (!g913) & (g908)) + ((!g903) & (g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (g904) & (g905) & (g906) & (g913) & (g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (g913) & (g908)) + ((g903) & (!g904) & (!g905) & (g906) & (g913) & (g908)) + ((g903) & (!g904) & (g905) & (g906) & (!g913) & (!g908)) + ((g903) & (g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((g903) & (g904) & (!g905) & (g906) & (g913) & (g908)) + ((g903) & (g904) & (g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (g904) & (g905) & (!g906) & (!g913) & (g908)) + ((g903) & (g904) & (g905) & (!g906) & (g913) & (g908)) + ((g903) & (g904) & (g905) & (g906) & (!g913) & (!g908)) + ((g903) & (g904) & (g905) & (g906) & (g913) & (g908)));
	assign g935 = (((!g903) & (!g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (!g905) & (g906) & (g913) & (g908)) + ((!g903) & (!g904) & (g905) & (g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (g905) & (g906) & (g913) & (g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (!g913) & (!g908)) + ((!g903) & (g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (g904) & (!g905) & (g906) & (!g913) & (!g908)) + ((!g903) & (g904) & (!g905) & (g906) & (!g913) & (g908)) + ((!g903) & (g904) & (!g905) & (g906) & (g913) & (!g908)) + ((!g903) & (g904) & (g905) & (!g906) & (!g913) & (!g908)) + ((!g903) & (g904) & (g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (g904) & (g905) & (!g906) & (g913) & (g908)) + ((g903) & (!g904) & (!g905) & (!g906) & (g913) & (g908)) + ((g903) & (!g904) & (!g905) & (g906) & (g913) & (!g908)) + ((g903) & (!g904) & (g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (g905) & (!g906) & (g913) & (!g908)) + ((g903) & (!g904) & (g905) & (!g906) & (g913) & (g908)) + ((g903) & (!g904) & (g905) & (g906) & (!g913) & (g908)) + ((g903) & (!g904) & (g905) & (g906) & (g913) & (!g908)) + ((g903) & (!g904) & (g905) & (g906) & (g913) & (g908)) + ((g903) & (g904) & (!g905) & (!g906) & (!g913) & (g908)) + ((g903) & (g904) & (!g905) & (!g906) & (g913) & (!g908)) + ((g903) & (g904) & (g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (g904) & (g905) & (!g906) & (!g913) & (g908)) + ((g903) & (g904) & (g905) & (g906) & (g913) & (g908)));
	assign g936 = (((!g932) & (!g933) & (!g934) & (!g935) & (!g914) & (g907)) + ((!g932) & (!g933) & (!g934) & (!g935) & (g914) & (!g907)) + ((!g932) & (!g933) & (!g934) & (!g935) & (g914) & (g907)) + ((!g932) & (!g933) & (!g934) & (g935) & (!g914) & (g907)) + ((!g932) & (!g933) & (!g934) & (g935) & (g914) & (!g907)) + ((!g932) & (!g933) & (g934) & (!g935) & (g914) & (!g907)) + ((!g932) & (!g933) & (g934) & (!g935) & (g914) & (g907)) + ((!g932) & (!g933) & (g934) & (g935) & (g914) & (!g907)) + ((!g932) & (g933) & (!g934) & (!g935) & (!g914) & (g907)) + ((!g932) & (g933) & (!g934) & (!g935) & (g914) & (g907)) + ((!g932) & (g933) & (!g934) & (g935) & (!g914) & (g907)) + ((!g932) & (g933) & (g934) & (!g935) & (g914) & (g907)) + ((g932) & (!g933) & (!g934) & (!g935) & (!g914) & (!g907)) + ((g932) & (!g933) & (!g934) & (!g935) & (!g914) & (g907)) + ((g932) & (!g933) & (!g934) & (!g935) & (g914) & (!g907)) + ((g932) & (!g933) & (!g934) & (!g935) & (g914) & (g907)) + ((g932) & (!g933) & (!g934) & (g935) & (!g914) & (!g907)) + ((g932) & (!g933) & (!g934) & (g935) & (!g914) & (g907)) + ((g932) & (!g933) & (!g934) & (g935) & (g914) & (!g907)) + ((g932) & (!g933) & (g934) & (!g935) & (!g914) & (!g907)) + ((g932) & (!g933) & (g934) & (!g935) & (g914) & (!g907)) + ((g932) & (!g933) & (g934) & (!g935) & (g914) & (g907)) + ((g932) & (!g933) & (g934) & (g935) & (!g914) & (!g907)) + ((g932) & (!g933) & (g934) & (g935) & (g914) & (!g907)) + ((g932) & (g933) & (!g934) & (!g935) & (!g914) & (!g907)) + ((g932) & (g933) & (!g934) & (!g935) & (!g914) & (g907)) + ((g932) & (g933) & (!g934) & (!g935) & (g914) & (g907)) + ((g932) & (g933) & (!g934) & (g935) & (!g914) & (!g907)) + ((g932) & (g933) & (!g934) & (g935) & (!g914) & (g907)) + ((g932) & (g933) & (g934) & (!g935) & (!g914) & (!g907)) + ((g932) & (g933) & (g934) & (!g935) & (g914) & (g907)) + ((g932) & (g933) & (g934) & (g935) & (!g914) & (!g907)));
	assign g938 = (((!sk[88]) & (g936) & (!g937)) + ((!sk[88]) & (g936) & (g937)) + ((sk[88]) & (!g936) & (g937)) + ((sk[88]) & (g936) & (!g937)));
	assign g939 = (((!g903) & (!g904) & (!g907) & (!g914) & (!g913) & (g908)) + ((!g903) & (!g904) & (g907) & (!g914) & (!g913) & (g908)) + ((!g903) & (!g904) & (g907) & (!g914) & (g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (!g914) & (g913) & (g908)) + ((!g903) & (!g904) & (g907) & (g914) & (!g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (g914) & (g913) & (!g908)) + ((!g903) & (g904) & (!g907) & (!g914) & (!g913) & (!g908)) + ((!g903) & (g904) & (!g907) & (!g914) & (!g913) & (g908)) + ((!g903) & (g904) & (!g907) & (g914) & (!g913) & (!g908)) + ((!g903) & (g904) & (!g907) & (g914) & (!g913) & (g908)) + ((!g903) & (g904) & (!g907) & (g914) & (g913) & (g908)) + ((!g903) & (g904) & (g907) & (g914) & (!g913) & (g908)) + ((!g903) & (g904) & (g907) & (g914) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g914) & (!g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g914) & (!g913) & (g908)) + ((g903) & (!g904) & (!g907) & (g914) & (!g913) & (g908)) + ((g903) & (!g904) & (g907) & (!g914) & (g913) & (!g908)) + ((g903) & (!g904) & (g907) & (g914) & (!g913) & (!g908)) + ((g903) & (!g904) & (g907) & (g914) & (!g913) & (g908)) + ((g903) & (!g904) & (g907) & (g914) & (g913) & (!g908)) + ((g903) & (g904) & (!g907) & (!g914) & (!g913) & (!g908)) + ((g903) & (g904) & (!g907) & (!g914) & (g913) & (!g908)) + ((g903) & (g904) & (!g907) & (g914) & (g913) & (!g908)) + ((g903) & (g904) & (g907) & (!g914) & (!g913) & (!g908)) + ((g903) & (g904) & (g907) & (!g914) & (!g913) & (g908)) + ((g903) & (g904) & (g907) & (g914) & (!g913) & (g908)));
	assign g940 = (((!g903) & (!g904) & (!g907) & (!g914) & (!g913) & (!g908)) + ((!g903) & (!g904) & (!g907) & (!g914) & (!g913) & (g908)) + ((!g903) & (!g904) & (!g907) & (!g914) & (g913) & (!g908)) + ((!g903) & (!g904) & (!g907) & (!g914) & (g913) & (g908)) + ((!g903) & (!g904) & (!g907) & (g914) & (!g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (!g914) & (!g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (!g914) & (g913) & (g908)) + ((!g903) & (!g904) & (g907) & (g914) & (!g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (g914) & (g913) & (g908)) + ((!g903) & (g904) & (!g907) & (!g914) & (!g913) & (g908)) + ((!g903) & (g904) & (!g907) & (g914) & (g913) & (!g908)) + ((!g903) & (g904) & (g907) & (!g914) & (!g913) & (!g908)) + ((!g903) & (g904) & (g907) & (!g914) & (!g913) & (g908)) + ((!g903) & (g904) & (g907) & (!g914) & (g913) & (!g908)) + ((!g903) & (g904) & (g907) & (!g914) & (g913) & (g908)) + ((!g903) & (g904) & (g907) & (g914) & (!g913) & (!g908)) + ((!g903) & (g904) & (g907) & (g914) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g914) & (!g913) & (g908)) + ((g903) & (!g904) & (!g907) & (!g914) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g914) & (g913) & (g908)) + ((g903) & (!g904) & (!g907) & (g914) & (!g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (g914) & (g913) & (g908)) + ((g903) & (!g904) & (g907) & (!g914) & (g913) & (!g908)) + ((g903) & (!g904) & (g907) & (!g914) & (g913) & (g908)) + ((g903) & (!g904) & (g907) & (g914) & (!g913) & (g908)) + ((g903) & (g904) & (!g907) & (!g914) & (g913) & (!g908)) + ((g903) & (g904) & (!g907) & (!g914) & (g913) & (g908)) + ((g903) & (g904) & (!g907) & (g914) & (!g913) & (!g908)) + ((g903) & (g904) & (!g907) & (g914) & (!g913) & (g908)) + ((g903) & (g904) & (g907) & (!g914) & (g913) & (!g908)) + ((g903) & (g904) & (g907) & (!g914) & (g913) & (g908)) + ((g903) & (g904) & (g907) & (g914) & (!g913) & (g908)));
	assign g941 = (((!g903) & (!g904) & (!g907) & (!g914) & (!g913) & (!g908)) + ((!g903) & (!g904) & (!g907) & (!g914) & (!g913) & (g908)) + ((!g903) & (!g904) & (g907) & (!g914) & (!g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (!g914) & (g913) & (g908)) + ((!g903) & (!g904) & (g907) & (g914) & (!g913) & (g908)) + ((!g903) & (g904) & (!g907) & (g914) & (!g913) & (!g908)) + ((!g903) & (g904) & (!g907) & (g914) & (g913) & (!g908)) + ((!g903) & (g904) & (!g907) & (g914) & (g913) & (g908)) + ((!g903) & (g904) & (g907) & (!g914) & (!g913) & (!g908)) + ((!g903) & (g904) & (g907) & (!g914) & (g913) & (!g908)) + ((!g903) & (g904) & (g907) & (!g914) & (g913) & (g908)) + ((!g903) & (g904) & (g907) & (g914) & (!g913) & (!g908)) + ((!g903) & (g904) & (g907) & (g914) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g914) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g914) & (g913) & (g908)) + ((g903) & (!g904) & (!g907) & (g914) & (!g913) & (g908)) + ((g903) & (!g904) & (!g907) & (g914) & (g913) & (g908)) + ((g903) & (!g904) & (g907) & (!g914) & (!g913) & (!g908)) + ((g903) & (!g904) & (g907) & (!g914) & (!g913) & (g908)) + ((g903) & (!g904) & (g907) & (!g914) & (g913) & (g908)) + ((g903) & (!g904) & (g907) & (g914) & (!g913) & (!g908)) + ((g903) & (!g904) & (g907) & (g914) & (!g913) & (g908)) + ((g903) & (!g904) & (g907) & (g914) & (g913) & (!g908)) + ((g903) & (!g904) & (g907) & (g914) & (g913) & (g908)) + ((g903) & (g904) & (!g907) & (!g914) & (!g913) & (g908)) + ((g903) & (g904) & (!g907) & (g914) & (!g913) & (!g908)) + ((g903) & (g904) & (!g907) & (g914) & (g913) & (!g908)) + ((g903) & (g904) & (g907) & (!g914) & (!g913) & (!g908)) + ((g903) & (g904) & (g907) & (!g914) & (!g913) & (g908)) + ((g903) & (g904) & (g907) & (!g914) & (g913) & (!g908)) + ((g903) & (g904) & (g907) & (g914) & (!g913) & (!g908)) + ((g903) & (g904) & (g907) & (g914) & (g913) & (!g908)));
	assign g942 = (((!g903) & (!g904) & (!g907) & (!g914) & (g913) & (g908)) + ((!g903) & (!g904) & (!g907) & (g914) & (!g913) & (!g908)) + ((!g903) & (!g904) & (!g907) & (g914) & (g913) & (g908)) + ((!g903) & (!g904) & (g907) & (!g914) & (!g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (!g914) & (g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (g914) & (!g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (g914) & (!g913) & (g908)) + ((!g903) & (!g904) & (g907) & (g914) & (g913) & (!g908)) + ((!g903) & (g904) & (!g907) & (!g914) & (!g913) & (!g908)) + ((!g903) & (g904) & (!g907) & (g914) & (!g913) & (g908)) + ((!g903) & (g904) & (!g907) & (g914) & (g913) & (!g908)) + ((!g903) & (g904) & (!g907) & (g914) & (g913) & (g908)) + ((!g903) & (g904) & (g907) & (!g914) & (!g913) & (!g908)) + ((!g903) & (g904) & (g907) & (g914) & (!g913) & (!g908)) + ((!g903) & (g904) & (g907) & (g914) & (!g913) & (g908)) + ((g903) & (!g904) & (!g907) & (!g914) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g914) & (g913) & (g908)) + ((g903) & (!g904) & (g907) & (!g914) & (!g913) & (!g908)) + ((g903) & (!g904) & (g907) & (!g914) & (g913) & (!g908)) + ((g903) & (!g904) & (g907) & (g914) & (g913) & (!g908)) + ((g903) & (g904) & (!g907) & (!g914) & (g913) & (!g908)) + ((g903) & (g904) & (!g907) & (g914) & (g913) & (g908)) + ((g903) & (g904) & (g907) & (!g914) & (!g913) & (!g908)) + ((g903) & (g904) & (g907) & (!g914) & (!g913) & (g908)) + ((g903) & (g904) & (g907) & (!g914) & (g913) & (!g908)) + ((g903) & (g904) & (g907) & (g914) & (!g913) & (!g908)));
	assign g943 = (((!g939) & (!g940) & (!g941) & (!g942) & (g905) & (g906)) + ((!g939) & (!g940) & (g941) & (!g942) & (!g905) & (g906)) + ((!g939) & (!g940) & (g941) & (!g942) & (g905) & (g906)) + ((!g939) & (!g940) & (g941) & (g942) & (!g905) & (g906)) + ((!g939) & (g940) & (!g941) & (!g942) & (g905) & (!g906)) + ((!g939) & (g940) & (!g941) & (!g942) & (g905) & (g906)) + ((!g939) & (g940) & (!g941) & (g942) & (g905) & (!g906)) + ((!g939) & (g940) & (g941) & (!g942) & (!g905) & (g906)) + ((!g939) & (g940) & (g941) & (!g942) & (g905) & (!g906)) + ((!g939) & (g940) & (g941) & (!g942) & (g905) & (g906)) + ((!g939) & (g940) & (g941) & (g942) & (!g905) & (g906)) + ((!g939) & (g940) & (g941) & (g942) & (g905) & (!g906)) + ((g939) & (!g940) & (!g941) & (!g942) & (!g905) & (!g906)) + ((g939) & (!g940) & (!g941) & (!g942) & (g905) & (g906)) + ((g939) & (!g940) & (!g941) & (g942) & (!g905) & (!g906)) + ((g939) & (!g940) & (g941) & (!g942) & (!g905) & (!g906)) + ((g939) & (!g940) & (g941) & (!g942) & (!g905) & (g906)) + ((g939) & (!g940) & (g941) & (!g942) & (g905) & (g906)) + ((g939) & (!g940) & (g941) & (g942) & (!g905) & (!g906)) + ((g939) & (!g940) & (g941) & (g942) & (!g905) & (g906)) + ((g939) & (g940) & (!g941) & (!g942) & (!g905) & (!g906)) + ((g939) & (g940) & (!g941) & (!g942) & (g905) & (!g906)) + ((g939) & (g940) & (!g941) & (!g942) & (g905) & (g906)) + ((g939) & (g940) & (!g941) & (g942) & (!g905) & (!g906)) + ((g939) & (g940) & (!g941) & (g942) & (g905) & (!g906)) + ((g939) & (g940) & (g941) & (!g942) & (!g905) & (!g906)) + ((g939) & (g940) & (g941) & (!g942) & (!g905) & (g906)) + ((g939) & (g940) & (g941) & (!g942) & (g905) & (!g906)) + ((g939) & (g940) & (g941) & (!g942) & (g905) & (g906)) + ((g939) & (g940) & (g941) & (g942) & (!g905) & (!g906)) + ((g939) & (g940) & (g941) & (g942) & (!g905) & (g906)) + ((g939) & (g940) & (g941) & (g942) & (g905) & (!g906)));
	assign g945 = (((!g943) & (sk[94]) & (g944)) + ((g943) & (!sk[94]) & (!g944)) + ((g943) & (!sk[94]) & (g944)) + ((g943) & (sk[94]) & (!g944)));
	assign g946 = (((!g903) & (!g904) & (!g907) & (!g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (!g907) & (!g906) & (g913) & (g908)) + ((!g903) & (!g904) & (!g907) & (g906) & (g913) & (g908)) + ((!g903) & (!g904) & (g907) & (!g906) & (!g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (!g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (g907) & (!g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (!g906) & (g913) & (g908)) + ((!g903) & (!g904) & (g907) & (g906) & (!g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (g906) & (!g913) & (g908)) + ((!g903) & (g904) & (!g907) & (!g906) & (!g913) & (g908)) + ((!g903) & (g904) & (!g907) & (!g906) & (g913) & (!g908)) + ((!g903) & (g904) & (!g907) & (g906) & (g913) & (g908)) + ((!g903) & (g904) & (g907) & (!g906) & (g913) & (!g908)) + ((!g903) & (g904) & (g907) & (!g906) & (g913) & (g908)) + ((!g903) & (g904) & (g907) & (g906) & (!g913) & (!g908)) + ((!g903) & (g904) & (g907) & (g906) & (!g913) & (g908)) + ((!g903) & (g904) & (g907) & (g906) & (g913) & (g908)) + ((g903) & (!g904) & (!g907) & (!g906) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g906) & (g913) & (g908)) + ((g903) & (!g904) & (!g907) & (g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (g906) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (g906) & (g913) & (g908)) + ((g903) & (!g904) & (g907) & (!g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (g907) & (!g906) & (g913) & (!g908)) + ((g903) & (!g904) & (g907) & (g906) & (g913) & (!g908)) + ((g903) & (g904) & (!g907) & (!g906) & (g913) & (g908)) + ((g903) & (g904) & (g907) & (!g906) & (!g913) & (!g908)) + ((g903) & (g904) & (g907) & (!g906) & (g913) & (g908)));
	assign g947 = (((!g903) & (!g904) & (!g907) & (!g906) & (!g913) & (!g908)) + ((!g903) & (!g904) & (!g907) & (g906) & (!g913) & (!g908)) + ((!g903) & (!g904) & (!g907) & (g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (!g907) & (g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (!g906) & (g913) & (g908)) + ((!g903) & (!g904) & (g907) & (g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (g907) & (g906) & (g913) & (g908)) + ((!g903) & (g904) & (!g907) & (!g906) & (!g913) & (!g908)) + ((!g903) & (g904) & (!g907) & (!g906) & (g913) & (!g908)) + ((!g903) & (g904) & (g907) & (!g906) & (!g913) & (g908)) + ((!g903) & (g904) & (g907) & (!g906) & (g913) & (g908)) + ((!g903) & (g904) & (g907) & (g906) & (!g913) & (g908)) + ((!g903) & (g904) & (g907) & (g906) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g906) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g906) & (g913) & (g908)) + ((g903) & (!g904) & (!g907) & (g906) & (!g913) & (g908)) + ((g903) & (!g904) & (!g907) & (g906) & (g913) & (g908)) + ((g903) & (!g904) & (g907) & (g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (g907) & (g906) & (!g913) & (g908)) + ((g903) & (!g904) & (g907) & (g906) & (g913) & (g908)) + ((g903) & (g904) & (!g907) & (!g906) & (!g913) & (g908)) + ((g903) & (g904) & (!g907) & (!g906) & (g913) & (!g908)) + ((g903) & (g904) & (!g907) & (g906) & (g913) & (!g908)) + ((g903) & (g904) & (g907) & (!g906) & (!g913) & (g908)) + ((g903) & (g904) & (g907) & (!g906) & (g913) & (g908)) + ((g903) & (g904) & (g907) & (g906) & (!g913) & (!g908)) + ((g903) & (g904) & (g907) & (g906) & (g913) & (g908)));
	assign g948 = (((!g903) & (!g904) & (!g907) & (!g906) & (g913) & (g908)) + ((!g903) & (!g904) & (!g907) & (g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (!g906) & (!g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (!g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (g907) & (!g906) & (g913) & (g908)) + ((!g903) & (!g904) & (g907) & (g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (g907) & (g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (g907) & (g906) & (g913) & (g908)) + ((!g903) & (g904) & (!g907) & (!g906) & (g913) & (!g908)) + ((!g903) & (g904) & (!g907) & (!g906) & (g913) & (g908)) + ((!g903) & (g904) & (g907) & (!g906) & (!g913) & (!g908)) + ((!g903) & (g904) & (g907) & (g906) & (!g913) & (g908)) + ((!g903) & (g904) & (g907) & (g906) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g906) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (!g906) & (g913) & (g908)) + ((g903) & (!g904) & (!g907) & (g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (g906) & (!g913) & (g908)) + ((g903) & (!g904) & (g907) & (!g906) & (!g913) & (g908)) + ((g903) & (!g904) & (g907) & (!g906) & (g913) & (g908)) + ((g903) & (!g904) & (g907) & (g906) & (g913) & (!g908)) + ((g903) & (g904) & (!g907) & (!g906) & (!g913) & (!g908)) + ((g903) & (g904) & (!g907) & (!g906) & (!g913) & (g908)) + ((g903) & (g904) & (!g907) & (!g906) & (g913) & (g908)) + ((g903) & (g904) & (!g907) & (g906) & (!g913) & (g908)) + ((g903) & (g904) & (!g907) & (g906) & (g913) & (!g908)) + ((g903) & (g904) & (g907) & (!g906) & (!g913) & (g908)) + ((g903) & (g904) & (g907) & (!g906) & (g913) & (!g908)) + ((g903) & (g904) & (g907) & (g906) & (!g913) & (!g908)) + ((g903) & (g904) & (g907) & (g906) & (g913) & (!g908)) + ((g903) & (g904) & (g907) & (g906) & (g913) & (g908)));
	assign g949 = (((!g903) & (!g904) & (!g907) & (!g906) & (g913) & (!g908)) + ((!g903) & (!g904) & (!g907) & (g906) & (!g913) & (!g908)) + ((!g903) & (!g904) & (!g907) & (g906) & (g913) & (g908)) + ((!g903) & (!g904) & (g907) & (!g906) & (!g913) & (g908)) + ((!g903) & (!g904) & (g907) & (!g906) & (g913) & (g908)) + ((!g903) & (!g904) & (g907) & (g906) & (g913) & (g908)) + ((!g903) & (g904) & (!g907) & (!g906) & (!g913) & (g908)) + ((!g903) & (g904) & (!g907) & (g906) & (!g913) & (g908)) + ((!g903) & (g904) & (!g907) & (g906) & (g913) & (g908)) + ((!g903) & (g904) & (g907) & (!g906) & (!g913) & (!g908)) + ((!g903) & (g904) & (g907) & (!g906) & (g913) & (!g908)) + ((!g903) & (g904) & (g907) & (g906) & (!g913) & (g908)) + ((!g903) & (g904) & (g907) & (g906) & (g913) & (g908)) + ((g903) & (!g904) & (!g907) & (!g906) & (g913) & (!g908)) + ((g903) & (!g904) & (!g907) & (g906) & (g913) & (g908)) + ((g903) & (!g904) & (g907) & (!g906) & (!g913) & (!g908)) + ((g903) & (!g904) & (g907) & (!g906) & (g913) & (g908)) + ((g903) & (!g904) & (g907) & (g906) & (!g913) & (!g908)) + ((g903) & (g904) & (!g907) & (!g906) & (g913) & (g908)) + ((g903) & (g904) & (!g907) & (g906) & (!g913) & (!g908)) + ((g903) & (g904) & (!g907) & (g906) & (!g913) & (g908)) + ((g903) & (g904) & (g907) & (!g906) & (g913) & (g908)));
	assign g950 = (((!g946) & (!g947) & (!g948) & (!g949) & (!g914) & (!g905)) + ((!g946) & (!g947) & (!g948) & (!g949) & (!g914) & (g905)) + ((!g946) & (!g947) & (!g948) & (!g949) & (g914) & (!g905)) + ((!g946) & (!g947) & (!g948) & (g949) & (!g914) & (!g905)) + ((!g946) & (!g947) & (!g948) & (g949) & (!g914) & (g905)) + ((!g946) & (!g947) & (!g948) & (g949) & (g914) & (!g905)) + ((!g946) & (!g947) & (!g948) & (g949) & (g914) & (g905)) + ((!g946) & (!g947) & (g948) & (!g949) & (!g914) & (!g905)) + ((!g946) & (!g947) & (g948) & (!g949) & (g914) & (!g905)) + ((!g946) & (!g947) & (g948) & (g949) & (!g914) & (!g905)) + ((!g946) & (!g947) & (g948) & (g949) & (g914) & (!g905)) + ((!g946) & (!g947) & (g948) & (g949) & (g914) & (g905)) + ((!g946) & (g947) & (!g948) & (!g949) & (!g914) & (!g905)) + ((!g946) & (g947) & (!g948) & (!g949) & (!g914) & (g905)) + ((!g946) & (g947) & (!g948) & (g949) & (!g914) & (!g905)) + ((!g946) & (g947) & (!g948) & (g949) & (!g914) & (g905)) + ((!g946) & (g947) & (!g948) & (g949) & (g914) & (g905)) + ((!g946) & (g947) & (g948) & (!g949) & (!g914) & (!g905)) + ((!g946) & (g947) & (g948) & (g949) & (!g914) & (!g905)) + ((!g946) & (g947) & (g948) & (g949) & (g914) & (g905)) + ((g946) & (!g947) & (!g948) & (!g949) & (!g914) & (g905)) + ((g946) & (!g947) & (!g948) & (!g949) & (g914) & (!g905)) + ((g946) & (!g947) & (!g948) & (g949) & (!g914) & (g905)) + ((g946) & (!g947) & (!g948) & (g949) & (g914) & (!g905)) + ((g946) & (!g947) & (!g948) & (g949) & (g914) & (g905)) + ((g946) & (!g947) & (g948) & (!g949) & (g914) & (!g905)) + ((g946) & (!g947) & (g948) & (g949) & (g914) & (!g905)) + ((g946) & (!g947) & (g948) & (g949) & (g914) & (g905)) + ((g946) & (g947) & (!g948) & (!g949) & (!g914) & (g905)) + ((g946) & (g947) & (!g948) & (g949) & (!g914) & (g905)) + ((g946) & (g947) & (!g948) & (g949) & (g914) & (g905)) + ((g946) & (g947) & (g948) & (g949) & (g914) & (g905)));
	assign g952 = (((!g950) & (sk[100]) & (g951)) + ((g950) & (!sk[100]) & (!g951)) + ((g950) & (!sk[100]) & (g951)) + ((g950) & (sk[100]) & (!g951)));
	assign g953 = (((!g903) & (!g914) & (!g905) & (!g906) & (!g913) & (g908)) + ((!g903) & (!g914) & (!g905) & (!g906) & (g913) & (g908)) + ((!g903) & (!g914) & (!g905) & (g906) & (!g913) & (!g908)) + ((!g903) & (!g914) & (!g905) & (g906) & (!g913) & (g908)) + ((!g903) & (!g914) & (!g905) & (g906) & (g913) & (!g908)) + ((!g903) & (!g914) & (!g905) & (g906) & (g913) & (g908)) + ((!g903) & (!g914) & (g905) & (!g906) & (!g913) & (g908)) + ((!g903) & (!g914) & (g905) & (!g906) & (g913) & (g908)) + ((!g903) & (!g914) & (g905) & (g906) & (g913) & (!g908)) + ((!g903) & (g914) & (g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (g914) & (g905) & (!g906) & (g913) & (g908)) + ((!g903) & (g914) & (g905) & (g906) & (!g913) & (g908)) + ((g903) & (!g914) & (!g905) & (!g906) & (g913) & (!g908)) + ((g903) & (!g914) & (!g905) & (g906) & (!g913) & (!g908)) + ((g903) & (!g914) & (!g905) & (g906) & (!g913) & (g908)) + ((g903) & (!g914) & (!g905) & (g906) & (g913) & (g908)) + ((g903) & (!g914) & (g905) & (!g906) & (!g913) & (g908)) + ((g903) & (!g914) & (g905) & (!g906) & (g913) & (g908)) + ((g903) & (!g914) & (g905) & (g906) & (g913) & (!g908)) + ((g903) & (!g914) & (g905) & (g906) & (g913) & (g908)) + ((g903) & (g914) & (!g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (g914) & (!g905) & (!g906) & (!g913) & (g908)) + ((g903) & (g914) & (!g905) & (!g906) & (g913) & (!g908)) + ((g903) & (g914) & (!g905) & (g906) & (!g913) & (!g908)) + ((g903) & (g914) & (g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (g914) & (g905) & (!g906) & (!g913) & (g908)) + ((g903) & (g914) & (g905) & (!g906) & (g913) & (!g908)) + ((g903) & (g914) & (g905) & (g906) & (!g913) & (g908)));
	assign g954 = (((!g903) & (!g914) & (!g905) & (!g906) & (!g913) & (!g908)) + ((!g903) & (!g914) & (!g905) & (g906) & (g913) & (g908)) + ((!g903) & (!g914) & (g905) & (!g906) & (!g913) & (!g908)) + ((!g903) & (!g914) & (g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (!g914) & (g905) & (!g906) & (g913) & (g908)) + ((!g903) & (!g914) & (g905) & (g906) & (!g913) & (!g908)) + ((!g903) & (!g914) & (g905) & (g906) & (g913) & (g908)) + ((!g903) & (g914) & (!g905) & (!g906) & (!g913) & (!g908)) + ((!g903) & (g914) & (!g905) & (!g906) & (g913) & (g908)) + ((!g903) & (g914) & (!g905) & (g906) & (!g913) & (g908)) + ((!g903) & (g914) & (g905) & (!g906) & (!g913) & (!g908)) + ((!g903) & (g914) & (g905) & (!g906) & (g913) & (g908)) + ((!g903) & (g914) & (g905) & (g906) & (g913) & (!g908)) + ((!g903) & (g914) & (g905) & (g906) & (g913) & (g908)) + ((g903) & (!g914) & (!g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (!g914) & (!g905) & (!g906) & (g913) & (g908)) + ((g903) & (!g914) & (!g905) & (g906) & (!g913) & (!g908)) + ((g903) & (!g914) & (!g905) & (g906) & (g913) & (g908)) + ((g903) & (!g914) & (g905) & (!g906) & (g913) & (g908)) + ((g903) & (!g914) & (g905) & (g906) & (!g913) & (g908)) + ((g903) & (g914) & (!g905) & (!g906) & (g913) & (!g908)) + ((g903) & (g914) & (!g905) & (!g906) & (g913) & (g908)) + ((g903) & (g914) & (!g905) & (g906) & (!g913) & (g908)) + ((g903) & (g914) & (!g905) & (g906) & (g913) & (!g908)) + ((g903) & (g914) & (!g905) & (g906) & (g913) & (g908)) + ((g903) & (g914) & (g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (g914) & (g905) & (!g906) & (g913) & (!g908)) + ((g903) & (g914) & (g905) & (g906) & (!g913) & (!g908)));
	assign g955 = (((!g903) & (!g914) & (!g905) & (!g906) & (!g913) & (g908)) + ((!g903) & (!g914) & (!g905) & (!g906) & (g913) & (g908)) + ((!g903) & (!g914) & (!g905) & (g906) & (g913) & (!g908)) + ((!g903) & (!g914) & (!g905) & (g906) & (g913) & (g908)) + ((!g903) & (!g914) & (g905) & (!g906) & (g913) & (g908)) + ((!g903) & (!g914) & (g905) & (g906) & (!g913) & (!g908)) + ((!g903) & (!g914) & (g905) & (g906) & (!g913) & (g908)) + ((!g903) & (!g914) & (g905) & (g906) & (g913) & (g908)) + ((!g903) & (g914) & (!g905) & (!g906) & (!g913) & (!g908)) + ((!g903) & (g914) & (!g905) & (!g906) & (!g913) & (g908)) + ((!g903) & (g914) & (!g905) & (!g906) & (g913) & (g908)) + ((!g903) & (g914) & (!g905) & (g906) & (!g913) & (g908)) + ((!g903) & (g914) & (!g905) & (g906) & (g913) & (!g908)) + ((!g903) & (g914) & (g905) & (!g906) & (!g913) & (g908)) + ((!g903) & (g914) & (g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (g914) & (g905) & (g906) & (!g913) & (!g908)) + ((!g903) & (g914) & (g905) & (g906) & (g913) & (!g908)) + ((!g903) & (g914) & (g905) & (g906) & (g913) & (g908)) + ((g903) & (!g914) & (!g905) & (!g906) & (!g913) & (g908)) + ((g903) & (!g914) & (!g905) & (g906) & (!g913) & (!g908)) + ((g903) & (!g914) & (!g905) & (g906) & (g913) & (!g908)) + ((g903) & (!g914) & (g905) & (!g906) & (g913) & (g908)) + ((g903) & (!g914) & (g905) & (g906) & (!g913) & (g908)) + ((g903) & (g914) & (!g905) & (!g906) & (!g913) & (g908)) + ((g903) & (g914) & (!g905) & (g906) & (!g913) & (!g908)) + ((g903) & (g914) & (!g905) & (g906) & (g913) & (!g908)) + ((g903) & (g914) & (g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (g914) & (g905) & (!g906) & (g913) & (!g908)) + ((g903) & (g914) & (g905) & (!g906) & (g913) & (g908)) + ((g903) & (g914) & (g905) & (g906) & (g913) & (g908)));
	assign g956 = (((!g903) & (!g914) & (!g905) & (!g906) & (g913) & (g908)) + ((!g903) & (!g914) & (!g905) & (g906) & (!g913) & (!g908)) + ((!g903) & (!g914) & (!g905) & (g906) & (g913) & (g908)) + ((!g903) & (!g914) & (g905) & (!g906) & (!g913) & (!g908)) + ((!g903) & (!g914) & (g905) & (g906) & (g913) & (!g908)) + ((!g903) & (!g914) & (g905) & (g906) & (g913) & (g908)) + ((!g903) & (g914) & (!g905) & (g906) & (!g913) & (!g908)) + ((!g903) & (g914) & (!g905) & (g906) & (g913) & (!g908)) + ((!g903) & (g914) & (g905) & (!g906) & (g913) & (!g908)) + ((!g903) & (g914) & (g905) & (!g906) & (g913) & (g908)) + ((g903) & (!g914) & (!g905) & (!g906) & (!g913) & (g908)) + ((g903) & (!g914) & (!g905) & (!g906) & (g913) & (!g908)) + ((g903) & (!g914) & (!g905) & (g906) & (!g913) & (g908)) + ((g903) & (!g914) & (g905) & (!g906) & (g913) & (!g908)) + ((g903) & (!g914) & (g905) & (!g906) & (g913) & (g908)) + ((g903) & (!g914) & (g905) & (g906) & (g913) & (!g908)) + ((g903) & (!g914) & (g905) & (g906) & (g913) & (g908)) + ((g903) & (g914) & (!g905) & (!g906) & (g913) & (!g908)) + ((g903) & (g914) & (!g905) & (g906) & (!g913) & (g908)) + ((g903) & (g914) & (g905) & (!g906) & (!g913) & (!g908)) + ((g903) & (g914) & (g905) & (!g906) & (g913) & (g908)) + ((g903) & (g914) & (g905) & (g906) & (!g913) & (g908)));
	assign g957 = (((!g953) & (!g954) & (!g955) & (!g956) & (!g907) & (!g904)) + ((!g953) & (!g954) & (!g955) & (!g956) & (!g907) & (g904)) + ((!g953) & (!g954) & (!g955) & (!g956) & (g907) & (!g904)) + ((!g953) & (!g954) & (!g955) & (g956) & (!g907) & (!g904)) + ((!g953) & (!g954) & (!g955) & (g956) & (!g907) & (g904)) + ((!g953) & (!g954) & (!g955) & (g956) & (g907) & (!g904)) + ((!g953) & (!g954) & (!g955) & (g956) & (g907) & (g904)) + ((!g953) & (!g954) & (g955) & (!g956) & (!g907) & (!g904)) + ((!g953) & (!g954) & (g955) & (!g956) & (g907) & (!g904)) + ((!g953) & (!g954) & (g955) & (g956) & (!g907) & (!g904)) + ((!g953) & (!g954) & (g955) & (g956) & (g907) & (!g904)) + ((!g953) & (!g954) & (g955) & (g956) & (g907) & (g904)) + ((!g953) & (g954) & (!g955) & (!g956) & (!g907) & (!g904)) + ((!g953) & (g954) & (!g955) & (!g956) & (!g907) & (g904)) + ((!g953) & (g954) & (!g955) & (g956) & (!g907) & (!g904)) + ((!g953) & (g954) & (!g955) & (g956) & (!g907) & (g904)) + ((!g953) & (g954) & (!g955) & (g956) & (g907) & (g904)) + ((!g953) & (g954) & (g955) & (!g956) & (!g907) & (!g904)) + ((!g953) & (g954) & (g955) & (g956) & (!g907) & (!g904)) + ((!g953) & (g954) & (g955) & (g956) & (g907) & (g904)) + ((g953) & (!g954) & (!g955) & (!g956) & (!g907) & (g904)) + ((g953) & (!g954) & (!g955) & (!g956) & (g907) & (!g904)) + ((g953) & (!g954) & (!g955) & (g956) & (!g907) & (g904)) + ((g953) & (!g954) & (!g955) & (g956) & (g907) & (!g904)) + ((g953) & (!g954) & (!g955) & (g956) & (g907) & (g904)) + ((g953) & (!g954) & (g955) & (!g956) & (g907) & (!g904)) + ((g953) & (!g954) & (g955) & (g956) & (g907) & (!g904)) + ((g953) & (!g954) & (g955) & (g956) & (g907) & (g904)) + ((g953) & (g954) & (!g955) & (!g956) & (!g907) & (g904)) + ((g953) & (g954) & (!g955) & (g956) & (!g907) & (g904)) + ((g953) & (g954) & (!g955) & (g956) & (g907) & (g904)) + ((g953) & (g954) & (g955) & (g956) & (g907) & (g904)));
	assign g959 = (((!g957) & (sk[106]) & (g958)) + ((g957) & (!sk[106]) & (!g958)) + ((g957) & (!sk[106]) & (g958)) + ((g957) & (sk[106]) & (!g958)));
	assign g960 = (((!g907) & (!g904) & (!g905) & (!g906) & (!g913) & (g914)) + ((!g907) & (!g904) & (!g905) & (!g906) & (g913) & (!g914)) + ((!g907) & (!g904) & (!g905) & (g906) & (!g913) & (g914)) + ((!g907) & (!g904) & (!g905) & (g906) & (g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (!g906) & (!g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (!g906) & (g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (g906) & (!g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (g906) & (g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (g906) & (g913) & (g914)) + ((!g907) & (g904) & (!g905) & (!g906) & (g913) & (!g914)) + ((!g907) & (g904) & (!g905) & (g906) & (g913) & (!g914)) + ((!g907) & (g904) & (!g905) & (g906) & (g913) & (g914)) + ((!g907) & (g904) & (g905) & (!g906) & (g913) & (g914)) + ((!g907) & (g904) & (g905) & (g906) & (!g913) & (!g914)) + ((g907) & (!g904) & (!g905) & (!g906) & (!g913) & (g914)) + ((g907) & (!g904) & (!g905) & (g906) & (!g913) & (g914)) + ((g907) & (!g904) & (g905) & (g906) & (g913) & (g914)) + ((g907) & (g904) & (!g905) & (!g906) & (g913) & (g914)) + ((g907) & (g904) & (!g905) & (g906) & (!g913) & (!g914)) + ((g907) & (g904) & (!g905) & (g906) & (g913) & (!g914)) + ((g907) & (g904) & (g905) & (!g906) & (!g913) & (g914)) + ((g907) & (g904) & (g905) & (!g906) & (g913) & (!g914)) + ((g907) & (g904) & (g905) & (!g906) & (g913) & (g914)) + ((g907) & (g904) & (g905) & (g906) & (!g913) & (g914)));
	assign g961 = (((!g907) & (!g904) & (!g905) & (!g906) & (!g913) & (!g914)) + ((!g907) & (!g904) & (!g905) & (!g906) & (!g913) & (g914)) + ((!g907) & (!g904) & (!g905) & (g906) & (!g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (!g906) & (!g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (!g906) & (g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (!g906) & (g913) & (g914)) + ((!g907) & (!g904) & (g905) & (g906) & (!g913) & (g914)) + ((!g907) & (!g904) & (g905) & (g906) & (g913) & (g914)) + ((!g907) & (g904) & (!g905) & (!g906) & (!g913) & (!g914)) + ((!g907) & (g904) & (!g905) & (!g906) & (g913) & (!g914)) + ((!g907) & (g904) & (!g905) & (g906) & (!g913) & (!g914)) + ((!g907) & (g904) & (!g905) & (g906) & (!g913) & (g914)) + ((!g907) & (g904) & (!g905) & (g906) & (g913) & (g914)) + ((!g907) & (g904) & (g905) & (!g906) & (!g913) & (g914)) + ((!g907) & (g904) & (g905) & (g906) & (!g913) & (!g914)) + ((!g907) & (g904) & (g905) & (g906) & (!g913) & (g914)) + ((g907) & (!g904) & (!g905) & (!g906) & (!g913) & (g914)) + ((g907) & (!g904) & (!g905) & (!g906) & (g913) & (g914)) + ((g907) & (!g904) & (!g905) & (g906) & (!g913) & (!g914)) + ((g907) & (!g904) & (!g905) & (g906) & (g913) & (g914)) + ((g907) & (!g904) & (g905) & (!g906) & (!g913) & (!g914)) + ((g907) & (!g904) & (g905) & (!g906) & (g913) & (g914)) + ((g907) & (!g904) & (g905) & (g906) & (g913) & (!g914)) + ((g907) & (g904) & (!g905) & (!g906) & (!g913) & (!g914)) + ((g907) & (g904) & (!g905) & (!g906) & (!g913) & (g914)) + ((g907) & (g904) & (!g905) & (!g906) & (g913) & (g914)) + ((g907) & (g904) & (!g905) & (g906) & (!g913) & (g914)) + ((g907) & (g904) & (!g905) & (g906) & (g913) & (!g914)) + ((g907) & (g904) & (g905) & (!g906) & (g913) & (!g914)) + ((g907) & (g904) & (g905) & (!g906) & (g913) & (g914)));
	assign g962 = (((!g907) & (!g904) & (!g905) & (!g906) & (g913) & (!g914)) + ((!g907) & (!g904) & (!g905) & (g906) & (!g913) & (!g914)) + ((!g907) & (!g904) & (!g905) & (g906) & (g913) & (!g914)) + ((!g907) & (!g904) & (!g905) & (g906) & (g913) & (g914)) + ((!g907) & (!g904) & (g905) & (!g906) & (!g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (!g906) & (!g913) & (g914)) + ((!g907) & (!g904) & (g905) & (!g906) & (g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (g906) & (!g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (g906) & (g913) & (g914)) + ((!g907) & (g904) & (!g905) & (!g906) & (!g913) & (g914)) + ((!g907) & (g904) & (!g905) & (!g906) & (g913) & (!g914)) + ((!g907) & (g904) & (!g905) & (!g906) & (g913) & (g914)) + ((!g907) & (g904) & (g905) & (!g906) & (!g913) & (g914)) + ((!g907) & (g904) & (g905) & (!g906) & (g913) & (!g914)) + ((!g907) & (g904) & (g905) & (!g906) & (g913) & (g914)) + ((!g907) & (g904) & (g905) & (g906) & (!g913) & (!g914)) + ((g907) & (!g904) & (!g905) & (!g906) & (g913) & (!g914)) + ((g907) & (!g904) & (!g905) & (g906) & (!g913) & (!g914)) + ((g907) & (!g904) & (!g905) & (g906) & (g913) & (g914)) + ((g907) & (!g904) & (g905) & (!g906) & (!g913) & (!g914)) + ((g907) & (!g904) & (g905) & (!g906) & (!g913) & (g914)) + ((g907) & (!g904) & (g905) & (g906) & (!g913) & (!g914)) + ((g907) & (!g904) & (g905) & (g906) & (g913) & (!g914)) + ((g907) & (g904) & (!g905) & (!g906) & (g913) & (!g914)) + ((g907) & (g904) & (!g905) & (g906) & (!g913) & (!g914)) + ((g907) & (g904) & (!g905) & (g906) & (g913) & (g914)) + ((g907) & (g904) & (g905) & (!g906) & (!g913) & (!g914)) + ((g907) & (g904) & (g905) & (!g906) & (g913) & (!g914)) + ((g907) & (g904) & (g905) & (!g906) & (g913) & (g914)) + ((g907) & (g904) & (g905) & (g906) & (!g913) & (g914)));
	assign g963 = (((!g907) & (!g904) & (!g905) & (!g906) & (!g913) & (g914)) + ((!g907) & (!g904) & (!g905) & (g906) & (g913) & (!g914)) + ((!g907) & (!g904) & (!g905) & (g906) & (g913) & (g914)) + ((!g907) & (!g904) & (g905) & (!g906) & (!g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (!g906) & (!g913) & (g914)) + ((!g907) & (!g904) & (g905) & (g906) & (g913) & (!g914)) + ((!g907) & (!g904) & (g905) & (g906) & (g913) & (g914)) + ((!g907) & (g904) & (!g905) & (!g906) & (!g913) & (!g914)) + ((!g907) & (g904) & (!g905) & (!g906) & (!g913) & (g914)) + ((!g907) & (g904) & (!g905) & (!g906) & (g913) & (g914)) + ((!g907) & (g904) & (!g905) & (g906) & (!g913) & (g914)) + ((!g907) & (g904) & (g905) & (!g906) & (!g913) & (g914)) + ((!g907) & (g904) & (g905) & (g906) & (!g913) & (!g914)) + ((!g907) & (g904) & (g905) & (g906) & (!g913) & (g914)) + ((!g907) & (g904) & (g905) & (g906) & (g913) & (!g914)) + ((!g907) & (g904) & (g905) & (g906) & (g913) & (g914)) + ((g907) & (!g904) & (!g905) & (g906) & (!g913) & (g914)) + ((g907) & (!g904) & (g905) & (!g906) & (!g913) & (!g914)) + ((g907) & (!g904) & (g905) & (g906) & (!g913) & (!g914)) + ((g907) & (!g904) & (g905) & (g906) & (!g913) & (g914)) + ((g907) & (!g904) & (g905) & (g906) & (g913) & (g914)) + ((g907) & (g904) & (!g905) & (!g906) & (!g913) & (g914)) + ((g907) & (g904) & (!g905) & (!g906) & (g913) & (g914)) + ((g907) & (g904) & (!g905) & (g906) & (!g913) & (!g914)) + ((g907) & (g904) & (!g905) & (g906) & (g913) & (!g914)) + ((g907) & (g904) & (!g905) & (g906) & (g913) & (g914)) + ((g907) & (g904) & (g905) & (!g906) & (g913) & (g914)) + ((g907) & (g904) & (g905) & (g906) & (g913) & (g914)));
	assign g964 = (((!g960) & (!g961) & (!g962) & (!g963) & (!g903) & (g908)) + ((!g960) & (!g961) & (!g962) & (!g963) & (g903) & (!g908)) + ((!g960) & (!g961) & (!g962) & (!g963) & (g903) & (g908)) + ((!g960) & (!g961) & (!g962) & (g963) & (!g903) & (g908)) + ((!g960) & (!g961) & (!g962) & (g963) & (g903) & (!g908)) + ((!g960) & (!g961) & (g962) & (!g963) & (g903) & (!g908)) + ((!g960) & (!g961) & (g962) & (!g963) & (g903) & (g908)) + ((!g960) & (!g961) & (g962) & (g963) & (g903) & (!g908)) + ((!g960) & (g961) & (!g962) & (!g963) & (!g903) & (g908)) + ((!g960) & (g961) & (!g962) & (!g963) & (g903) & (g908)) + ((!g960) & (g961) & (!g962) & (g963) & (!g903) & (g908)) + ((!g960) & (g961) & (g962) & (!g963) & (g903) & (g908)) + ((g960) & (!g961) & (!g962) & (!g963) & (!g903) & (!g908)) + ((g960) & (!g961) & (!g962) & (!g963) & (!g903) & (g908)) + ((g960) & (!g961) & (!g962) & (!g963) & (g903) & (!g908)) + ((g960) & (!g961) & (!g962) & (!g963) & (g903) & (g908)) + ((g960) & (!g961) & (!g962) & (g963) & (!g903) & (!g908)) + ((g960) & (!g961) & (!g962) & (g963) & (!g903) & (g908)) + ((g960) & (!g961) & (!g962) & (g963) & (g903) & (!g908)) + ((g960) & (!g961) & (g962) & (!g963) & (!g903) & (!g908)) + ((g960) & (!g961) & (g962) & (!g963) & (g903) & (!g908)) + ((g960) & (!g961) & (g962) & (!g963) & (g903) & (g908)) + ((g960) & (!g961) & (g962) & (g963) & (!g903) & (!g908)) + ((g960) & (!g961) & (g962) & (g963) & (g903) & (!g908)) + ((g960) & (g961) & (!g962) & (!g963) & (!g903) & (!g908)) + ((g960) & (g961) & (!g962) & (!g963) & (!g903) & (g908)) + ((g960) & (g961) & (!g962) & (!g963) & (g903) & (g908)) + ((g960) & (g961) & (!g962) & (g963) & (!g903) & (!g908)) + ((g960) & (g961) & (!g962) & (g963) & (!g903) & (g908)) + ((g960) & (g961) & (g962) & (!g963) & (!g903) & (!g908)) + ((g960) & (g961) & (g962) & (!g963) & (g903) & (g908)) + ((g960) & (g961) & (g962) & (g963) & (!g903) & (!g908)));
	assign g966 = (((!sk[112]) & (g964) & (!g965)) + ((!sk[112]) & (g964) & (g965)) + ((sk[112]) & (!g964) & (g965)) + ((sk[112]) & (g964) & (!g965)));
	assign g973 = (((!g967) & (!g968) & (!g969) & (!g970) & (g971) & (g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g971) & (!g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g971) & (g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (g971) & (!g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (!g971) & (!g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (!g971) & (g972)) + ((!g967) & (!g968) & (g969) & (g970) & (!g971) & (!g972)) + ((!g967) & (!g968) & (g969) & (g970) & (g971) & (g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (g971) & (!g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (g971) & (g972)) + ((!g967) & (g968) & (!g969) & (g970) & (g971) & (!g972)) + ((!g967) & (g968) & (!g969) & (g970) & (g971) & (g972)) + ((!g967) & (g968) & (g969) & (!g970) & (g971) & (!g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (!g971) & (!g972)) + ((g967) & (!g968) & (g969) & (!g970) & (g971) & (!g972)) + ((g967) & (!g968) & (g969) & (g970) & (!g971) & (g972)) + ((g967) & (!g968) & (g969) & (g970) & (g971) & (g972)) + ((g967) & (g968) & (!g969) & (!g970) & (!g971) & (g972)) + ((g967) & (g968) & (!g969) & (!g970) & (g971) & (!g972)) + ((g967) & (g968) & (g969) & (!g970) & (!g971) & (g972)) + ((g967) & (g968) & (g969) & (!g970) & (g971) & (!g972)) + ((g967) & (g968) & (g969) & (g970) & (!g971) & (!g972)) + ((g967) & (g968) & (g969) & (g970) & (g971) & (!g972)) + ((g967) & (g968) & (g969) & (g970) & (g971) & (g972)));
	assign g974 = (((!g967) & (!g968) & (!g969) & (!g970) & (g971) & (!g972)) + ((!g967) & (!g968) & (!g969) & (!g970) & (g971) & (g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g971) & (!g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g971) & (g972)) + ((!g967) & (!g968) & (g969) & (g970) & (!g971) & (g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (!g971) & (!g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (!g971) & (g972)) + ((!g967) & (g968) & (g969) & (!g970) & (!g971) & (!g972)) + ((!g967) & (g968) & (g969) & (!g970) & (!g971) & (g972)) + ((!g967) & (g968) & (g969) & (!g970) & (g971) & (!g972)) + ((!g967) & (g968) & (g969) & (g970) & (g971) & (g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (!g971) & (g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (g971) & (!g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (g971) & (g972)) + ((g967) & (!g968) & (!g969) & (g970) & (g971) & (!g972)) + ((g967) & (!g968) & (g969) & (!g970) & (!g971) & (!g972)) + ((g967) & (!g968) & (g969) & (!g970) & (g971) & (g972)) + ((g967) & (!g968) & (g969) & (g970) & (!g971) & (g972)) + ((g967) & (!g968) & (g969) & (g970) & (g971) & (g972)) + ((g967) & (g968) & (!g969) & (!g970) & (!g971) & (!g972)) + ((g967) & (g968) & (!g969) & (!g970) & (!g971) & (g972)) + ((g967) & (g968) & (!g969) & (!g970) & (g971) & (!g972)) + ((g967) & (g968) & (!g969) & (!g970) & (g971) & (g972)) + ((g967) & (g968) & (!g969) & (g970) & (!g971) & (!g972)) + ((g967) & (g968) & (!g969) & (g970) & (g971) & (!g972)) + ((g967) & (g968) & (!g969) & (g970) & (g971) & (g972)) + ((g967) & (g968) & (g969) & (!g970) & (g971) & (!g972)) + ((g967) & (g968) & (g969) & (!g970) & (g971) & (g972)) + ((g967) & (g968) & (g969) & (g970) & (!g971) & (g972)) + ((g967) & (g968) & (g969) & (g970) & (g971) & (!g972)));
	assign g975 = (((!g967) & (!g968) & (!g969) & (!g970) & (!g971) & (!g972)) + ((!g967) & (!g968) & (!g969) & (!g970) & (g971) & (g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (g971) & (g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (!g971) & (!g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (!g971) & (g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (g971) & (g972)) + ((!g967) & (!g968) & (g969) & (g970) & (!g971) & (g972)) + ((!g967) & (!g968) & (g969) & (g970) & (g971) & (!g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (!g971) & (!g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (g971) & (!g972)) + ((!g967) & (g968) & (!g969) & (g970) & (g971) & (g972)) + ((!g967) & (g968) & (g969) & (g970) & (!g971) & (!g972)) + ((!g967) & (g968) & (g969) & (g970) & (g971) & (!g972)) + ((g967) & (!g968) & (!g969) & (g970) & (!g971) & (!g972)) + ((g967) & (!g968) & (!g969) & (g970) & (!g971) & (g972)) + ((g967) & (!g968) & (!g969) & (g970) & (g971) & (!g972)) + ((g967) & (!g968) & (g969) & (!g970) & (!g971) & (!g972)) + ((g967) & (!g968) & (g969) & (!g970) & (g971) & (g972)) + ((g967) & (!g968) & (g969) & (g970) & (!g971) & (!g972)) + ((g967) & (!g968) & (g969) & (g970) & (!g971) & (g972)) + ((g967) & (!g968) & (g969) & (g970) & (g971) & (!g972)) + ((g967) & (!g968) & (g969) & (g970) & (g971) & (g972)) + ((g967) & (g968) & (!g969) & (!g970) & (g971) & (g972)) + ((g967) & (g968) & (!g969) & (g970) & (!g971) & (!g972)) + ((g967) & (g968) & (!g969) & (g970) & (g971) & (!g972)) + ((g967) & (g968) & (!g969) & (g970) & (g971) & (g972)) + ((g967) & (g968) & (g969) & (!g970) & (!g971) & (!g972)) + ((g967) & (g968) & (g969) & (g970) & (!g971) & (!g972)) + ((g967) & (g968) & (g969) & (g970) & (!g971) & (g972)) + ((g967) & (g968) & (g969) & (g970) & (g971) & (g972)));
	assign g976 = (((!g967) & (!g968) & (!g969) & (!g970) & (!g971) & (g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (g971) & (!g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (g971) & (g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (!g971) & (g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (g971) & (g972)) + ((!g967) & (!g968) & (g969) & (g970) & (!g971) & (g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (!g971) & (!g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (!g971) & (g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (g971) & (!g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (g971) & (g972)) + ((!g967) & (g968) & (!g969) & (g970) & (g971) & (!g972)) + ((!g967) & (g968) & (!g969) & (g970) & (g971) & (g972)) + ((!g967) & (g968) & (g969) & (g970) & (!g971) & (!g972)) + ((!g967) & (g968) & (g969) & (g970) & (g971) & (!g972)) + ((!g967) & (g968) & (g969) & (g970) & (g971) & (g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (!g971) & (!g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (g971) & (g972)) + ((g967) & (!g968) & (!g969) & (g970) & (g971) & (!g972)) + ((g967) & (!g968) & (!g969) & (g970) & (g971) & (g972)) + ((g967) & (!g968) & (g969) & (!g970) & (!g971) & (g972)) + ((g967) & (!g968) & (g969) & (!g970) & (g971) & (!g972)) + ((g967) & (!g968) & (g969) & (g970) & (g971) & (!g972)) + ((g967) & (g968) & (!g969) & (!g970) & (!g971) & (g972)) + ((g967) & (g968) & (!g969) & (!g970) & (g971) & (g972)) + ((g967) & (g968) & (!g969) & (g970) & (g971) & (!g972)) + ((g967) & (g968) & (!g969) & (g970) & (g971) & (g972)) + ((g967) & (g968) & (g969) & (!g970) & (!g971) & (g972)) + ((g967) & (g968) & (g969) & (g970) & (!g971) & (!g972)));
	assign g979 = (((!g973) & (!g974) & (!g975) & (!g976) & (!g977) & (!g978)) + ((!g973) & (!g974) & (!g975) & (g976) & (!g977) & (!g978)) + ((!g973) & (!g974) & (!g975) & (g976) & (g977) & (g978)) + ((!g973) & (!g974) & (g975) & (!g976) & (!g977) & (!g978)) + ((!g973) & (!g974) & (g975) & (!g976) & (!g977) & (g978)) + ((!g973) & (!g974) & (g975) & (g976) & (!g977) & (!g978)) + ((!g973) & (!g974) & (g975) & (g976) & (!g977) & (g978)) + ((!g973) & (!g974) & (g975) & (g976) & (g977) & (g978)) + ((!g973) & (g974) & (!g975) & (!g976) & (!g977) & (!g978)) + ((!g973) & (g974) & (!g975) & (!g976) & (g977) & (!g978)) + ((!g973) & (g974) & (!g975) & (g976) & (!g977) & (!g978)) + ((!g973) & (g974) & (!g975) & (g976) & (g977) & (!g978)) + ((!g973) & (g974) & (!g975) & (g976) & (g977) & (g978)) + ((!g973) & (g974) & (g975) & (!g976) & (!g977) & (!g978)) + ((!g973) & (g974) & (g975) & (!g976) & (!g977) & (g978)) + ((!g973) & (g974) & (g975) & (!g976) & (g977) & (!g978)) + ((!g973) & (g974) & (g975) & (g976) & (!g977) & (!g978)) + ((!g973) & (g974) & (g975) & (g976) & (!g977) & (g978)) + ((!g973) & (g974) & (g975) & (g976) & (g977) & (!g978)) + ((!g973) & (g974) & (g975) & (g976) & (g977) & (g978)) + ((g973) & (!g974) & (!g975) & (g976) & (g977) & (g978)) + ((g973) & (!g974) & (g975) & (!g976) & (!g977) & (g978)) + ((g973) & (!g974) & (g975) & (g976) & (!g977) & (g978)) + ((g973) & (!g974) & (g975) & (g976) & (g977) & (g978)) + ((g973) & (g974) & (!g975) & (!g976) & (g977) & (!g978)) + ((g973) & (g974) & (!g975) & (g976) & (g977) & (!g978)) + ((g973) & (g974) & (!g975) & (g976) & (g977) & (g978)) + ((g973) & (g974) & (g975) & (!g976) & (!g977) & (g978)) + ((g973) & (g974) & (g975) & (!g976) & (g977) & (!g978)) + ((g973) & (g974) & (g975) & (g976) & (!g977) & (g978)) + ((g973) & (g974) & (g975) & (g976) & (g977) & (!g978)) + ((g973) & (g974) & (g975) & (g976) & (g977) & (g978)));
	assign g981 = (((!sk[118]) & (g979) & (!g980)) + ((!sk[118]) & (g979) & (g980)) + ((sk[118]) & (!g979) & (g980)) + ((sk[118]) & (g979) & (!g980)));
	assign g982 = (((!g967) & (!g968) & (!g969) & (!g970) & (!g977) & (g971)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g977) & (!g971)) + ((!g967) & (!g968) & (!g969) & (g970) & (g977) & (!g971)) + ((!g967) & (!g968) & (g969) & (!g970) & (g977) & (g971)) + ((!g967) & (!g968) & (g969) & (g970) & (!g977) & (g971)) + ((!g967) & (!g968) & (g969) & (g970) & (g977) & (!g971)) + ((!g967) & (g968) & (!g969) & (!g970) & (!g977) & (g971)) + ((!g967) & (g968) & (!g969) & (!g970) & (g977) & (!g971)) + ((!g967) & (g968) & (!g969) & (!g970) & (g977) & (g971)) + ((!g967) & (g968) & (g969) & (!g970) & (g977) & (g971)) + ((!g967) & (g968) & (g969) & (g970) & (g977) & (g971)) + ((g967) & (!g968) & (!g969) & (!g970) & (!g977) & (!g971)) + ((g967) & (!g968) & (!g969) & (!g970) & (g977) & (g971)) + ((g967) & (!g968) & (!g969) & (g970) & (!g977) & (!g971)) + ((g967) & (!g968) & (!g969) & (g970) & (g977) & (!g971)) + ((g967) & (!g968) & (g969) & (!g970) & (g977) & (!g971)) + ((g967) & (!g968) & (g969) & (!g970) & (g977) & (g971)) + ((g967) & (!g968) & (g969) & (g970) & (g977) & (!g971)) + ((g967) & (!g968) & (g969) & (g970) & (g977) & (g971)) + ((g967) & (g968) & (!g969) & (!g970) & (g977) & (!g971)) + ((g967) & (g968) & (!g969) & (!g970) & (g977) & (g971)) + ((g967) & (g968) & (!g969) & (g970) & (g977) & (g971)) + ((g967) & (g968) & (g969) & (!g970) & (!g977) & (!g971)) + ((g967) & (g968) & (g969) & (!g970) & (!g977) & (g971)) + ((g967) & (g968) & (g969) & (!g970) & (g977) & (!g971)) + ((g967) & (g968) & (g969) & (g970) & (!g977) & (g971)) + ((g967) & (g968) & (g969) & (g970) & (g977) & (!g971)));
	assign g983 = (((!g967) & (!g968) & (!g969) & (!g970) & (!g977) & (g971)) + ((!g967) & (!g968) & (!g969) & (!g970) & (g977) & (!g971)) + ((!g967) & (!g968) & (!g969) & (!g970) & (g977) & (g971)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g977) & (!g971)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g977) & (g971)) + ((!g967) & (!g968) & (!g969) & (g970) & (g977) & (g971)) + ((!g967) & (!g968) & (g969) & (!g970) & (g977) & (!g971)) + ((!g967) & (!g968) & (g969) & (g970) & (!g977) & (!g971)) + ((!g967) & (!g968) & (g969) & (g970) & (!g977) & (g971)) + ((!g967) & (!g968) & (g969) & (g970) & (g977) & (g971)) + ((!g967) & (g968) & (!g969) & (!g970) & (g977) & (g971)) + ((!g967) & (g968) & (!g969) & (g970) & (!g977) & (!g971)) + ((!g967) & (g968) & (!g969) & (g970) & (g977) & (!g971)) + ((!g967) & (g968) & (g969) & (!g970) & (g977) & (!g971)) + ((!g967) & (g968) & (g969) & (!g970) & (g977) & (g971)) + ((!g967) & (g968) & (g969) & (g970) & (!g977) & (!g971)) + ((g967) & (!g968) & (!g969) & (!g970) & (!g977) & (!g971)) + ((g967) & (!g968) & (!g969) & (g970) & (!g977) & (!g971)) + ((g967) & (!g968) & (!g969) & (g970) & (!g977) & (g971)) + ((g967) & (!g968) & (g969) & (!g970) & (!g977) & (g971)) + ((g967) & (!g968) & (g969) & (!g970) & (g977) & (g971)) + ((g967) & (!g968) & (g969) & (g970) & (!g977) & (!g971)) + ((g967) & (!g968) & (g969) & (g970) & (!g977) & (g971)) + ((g967) & (g968) & (!g969) & (g970) & (!g977) & (!g971)) + ((g967) & (g968) & (!g969) & (g970) & (g977) & (g971)) + ((g967) & (g968) & (g969) & (!g970) & (!g977) & (!g971)) + ((g967) & (g968) & (g969) & (!g970) & (!g977) & (g971)) + ((g967) & (g968) & (g969) & (!g970) & (g977) & (g971)) + ((g967) & (g968) & (g969) & (g970) & (!g977) & (!g971)) + ((g967) & (g968) & (g969) & (g970) & (!g977) & (g971)) + ((g967) & (g968) & (g969) & (g970) & (g977) & (!g971)));
	assign g984 = (((!g967) & (!g968) & (!g969) & (!g970) & (!g977) & (g971)) + ((!g967) & (!g968) & (!g969) & (g970) & (g977) & (!g971)) + ((!g967) & (!g968) & (g969) & (!g970) & (!g977) & (!g971)) + ((!g967) & (!g968) & (g969) & (!g970) & (g977) & (!g971)) + ((!g967) & (!g968) & (g969) & (g970) & (!g977) & (g971)) + ((!g967) & (!g968) & (g969) & (g970) & (g977) & (!g971)) + ((!g967) & (!g968) & (g969) & (g970) & (g977) & (g971)) + ((!g967) & (g968) & (!g969) & (!g970) & (!g977) & (!g971)) + ((!g967) & (g968) & (!g969) & (!g970) & (g977) & (!g971)) + ((!g967) & (g968) & (!g969) & (g970) & (!g977) & (!g971)) + ((!g967) & (g968) & (!g969) & (g970) & (g977) & (g971)) + ((!g967) & (g968) & (g969) & (!g970) & (g977) & (g971)) + ((!g967) & (g968) & (g969) & (g970) & (!g977) & (g971)) + ((!g967) & (g968) & (g969) & (g970) & (g977) & (!g971)) + ((g967) & (!g968) & (!g969) & (!g970) & (g977) & (g971)) + ((g967) & (!g968) & (!g969) & (g970) & (!g977) & (!g971)) + ((g967) & (!g968) & (!g969) & (g970) & (g977) & (!g971)) + ((g967) & (!g968) & (g969) & (!g970) & (!g977) & (!g971)) + ((g967) & (!g968) & (g969) & (!g970) & (!g977) & (g971)) + ((g967) & (!g968) & (g969) & (!g970) & (g977) & (!g971)) + ((g967) & (!g968) & (g969) & (!g970) & (g977) & (g971)) + ((g967) & (!g968) & (g969) & (g970) & (g977) & (!g971)) + ((g967) & (g968) & (!g969) & (!g970) & (!g977) & (g971)) + ((g967) & (g968) & (!g969) & (!g970) & (g977) & (g971)) + ((g967) & (g968) & (!g969) & (g970) & (!g977) & (g971)) + ((g967) & (g968) & (g969) & (!g970) & (!g977) & (!g971)) + ((g967) & (g968) & (g969) & (!g970) & (!g977) & (g971)) + ((g967) & (g968) & (g969) & (!g970) & (g977) & (g971)) + ((g967) & (g968) & (g969) & (g970) & (!g977) & (!g971)) + ((g967) & (g968) & (g969) & (g970) & (!g977) & (g971)) + ((g967) & (g968) & (g969) & (g970) & (g977) & (!g971)) + ((g967) & (g968) & (g969) & (g970) & (g977) & (g971)));
	assign g985 = (((!g967) & (!g968) & (!g969) & (!g970) & (g977) & (!g971)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g977) & (!g971)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g977) & (g971)) + ((!g967) & (!g968) & (g969) & (!g970) & (g977) & (g971)) + ((!g967) & (!g968) & (g969) & (g970) & (!g977) & (g971)) + ((!g967) & (g968) & (!g969) & (!g970) & (!g977) & (!g971)) + ((!g967) & (g968) & (!g969) & (!g970) & (g977) & (!g971)) + ((!g967) & (g968) & (!g969) & (g970) & (!g977) & (g971)) + ((!g967) & (g968) & (g969) & (!g970) & (!g977) & (g971)) + ((!g967) & (g968) & (g969) & (!g970) & (g977) & (!g971)) + ((!g967) & (g968) & (g969) & (!g970) & (g977) & (g971)) + ((!g967) & (g968) & (g969) & (g970) & (g977) & (!g971)) + ((!g967) & (g968) & (g969) & (g970) & (g977) & (g971)) + ((g967) & (!g968) & (!g969) & (!g970) & (!g977) & (!g971)) + ((g967) & (!g968) & (!g969) & (g970) & (!g977) & (!g971)) + ((g967) & (!g968) & (!g969) & (g970) & (!g977) & (g971)) + ((g967) & (!g968) & (!g969) & (g970) & (g977) & (!g971)) + ((g967) & (!g968) & (g969) & (!g970) & (!g977) & (!g971)) + ((g967) & (!g968) & (g969) & (!g970) & (g977) & (g971)) + ((g967) & (!g968) & (g969) & (g970) & (g977) & (!g971)) + ((g967) & (g968) & (!g969) & (!g970) & (!g977) & (!g971)) + ((g967) & (g968) & (!g969) & (g970) & (!g977) & (!g971)) + ((g967) & (g968) & (!g969) & (g970) & (g977) & (!g971)) + ((g967) & (g968) & (!g969) & (g970) & (g977) & (g971)) + ((g967) & (g968) & (g969) & (g970) & (!g977) & (g971)) + ((g967) & (g968) & (g969) & (g970) & (g977) & (g971)));
	assign g986 = (((!g982) & (!g983) & (!g984) & (!g985) & (!g972) & (!g978)) + ((!g982) & (!g983) & (!g984) & (!g985) & (g972) & (!g978)) + ((!g982) & (!g983) & (!g984) & (g985) & (!g972) & (!g978)) + ((!g982) & (!g983) & (!g984) & (g985) & (g972) & (!g978)) + ((!g982) & (!g983) & (!g984) & (g985) & (g972) & (g978)) + ((!g982) & (!g983) & (g984) & (!g985) & (!g972) & (!g978)) + ((!g982) & (!g983) & (g984) & (!g985) & (!g972) & (g978)) + ((!g982) & (!g983) & (g984) & (!g985) & (g972) & (!g978)) + ((!g982) & (!g983) & (g984) & (g985) & (!g972) & (!g978)) + ((!g982) & (!g983) & (g984) & (g985) & (!g972) & (g978)) + ((!g982) & (!g983) & (g984) & (g985) & (g972) & (!g978)) + ((!g982) & (!g983) & (g984) & (g985) & (g972) & (g978)) + ((!g982) & (g983) & (!g984) & (!g985) & (!g972) & (!g978)) + ((!g982) & (g983) & (!g984) & (g985) & (!g972) & (!g978)) + ((!g982) & (g983) & (!g984) & (g985) & (g972) & (g978)) + ((!g982) & (g983) & (g984) & (!g985) & (!g972) & (!g978)) + ((!g982) & (g983) & (g984) & (!g985) & (!g972) & (g978)) + ((!g982) & (g983) & (g984) & (g985) & (!g972) & (!g978)) + ((!g982) & (g983) & (g984) & (g985) & (!g972) & (g978)) + ((!g982) & (g983) & (g984) & (g985) & (g972) & (g978)) + ((g982) & (!g983) & (!g984) & (!g985) & (g972) & (!g978)) + ((g982) & (!g983) & (!g984) & (g985) & (g972) & (!g978)) + ((g982) & (!g983) & (!g984) & (g985) & (g972) & (g978)) + ((g982) & (!g983) & (g984) & (!g985) & (!g972) & (g978)) + ((g982) & (!g983) & (g984) & (!g985) & (g972) & (!g978)) + ((g982) & (!g983) & (g984) & (g985) & (!g972) & (g978)) + ((g982) & (!g983) & (g984) & (g985) & (g972) & (!g978)) + ((g982) & (!g983) & (g984) & (g985) & (g972) & (g978)) + ((g982) & (g983) & (!g984) & (g985) & (g972) & (g978)) + ((g982) & (g983) & (g984) & (!g985) & (!g972) & (g978)) + ((g982) & (g983) & (g984) & (g985) & (!g972) & (g978)) + ((g982) & (g983) & (g984) & (g985) & (g972) & (g978)));
	assign g988 = (((!g986) & (sk[124]) & (g987)) + ((g986) & (!sk[124]) & (!g987)) + ((g986) & (!sk[124]) & (g987)) + ((g986) & (sk[124]) & (!g987)));
	assign g989 = (((!g971) & (!g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((!g971) & (!g968) & (!g969) & (!g970) & (g977) & (g972)) + ((!g971) & (!g968) & (!g969) & (g970) & (!g977) & (g972)) + ((!g971) & (!g968) & (!g969) & (g970) & (g977) & (!g972)) + ((!g971) & (!g968) & (!g969) & (g970) & (g977) & (g972)) + ((!g971) & (!g968) & (g969) & (!g970) & (!g977) & (g972)) + ((!g971) & (!g968) & (g969) & (g970) & (!g977) & (!g972)) + ((!g971) & (!g968) & (g969) & (g970) & (g977) & (!g972)) + ((!g971) & (g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((!g971) & (g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((!g971) & (g968) & (!g969) & (g970) & (!g977) & (g972)) + ((!g971) & (g968) & (g969) & (!g970) & (!g977) & (!g972)) + ((!g971) & (g968) & (g969) & (!g970) & (!g977) & (g972)) + ((!g971) & (g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g971) & (g968) & (g969) & (!g970) & (g977) & (g972)) + ((g971) & (!g968) & (!g969) & (g970) & (!g977) & (g972)) + ((g971) & (!g968) & (!g969) & (g970) & (g977) & (g972)) + ((g971) & (g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((g971) & (g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((g971) & (g968) & (!g969) & (g970) & (g977) & (!g972)) + ((g971) & (g968) & (g969) & (g970) & (!g977) & (!g972)) + ((g971) & (g968) & (g969) & (g970) & (!g977) & (g972)));
	assign g990 = (((!g971) & (!g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((!g971) & (!g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((!g971) & (!g968) & (!g969) & (g970) & (g977) & (g972)) + ((!g971) & (!g968) & (g969) & (!g970) & (!g977) & (!g972)) + ((!g971) & (!g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g971) & (!g968) & (g969) & (g970) & (!g977) & (g972)) + ((!g971) & (g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((!g971) & (g968) & (!g969) & (!g970) & (g977) & (g972)) + ((!g971) & (g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((!g971) & (g968) & (!g969) & (g970) & (!g977) & (g972)) + ((!g971) & (g968) & (!g969) & (g970) & (g977) & (g972)) + ((!g971) & (g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g971) & (g968) & (g969) & (!g970) & (g977) & (g972)) + ((!g971) & (g968) & (g969) & (g970) & (g977) & (!g972)) + ((g971) & (!g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((g971) & (!g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((g971) & (!g968) & (!g969) & (!g970) & (g977) & (g972)) + ((g971) & (!g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((g971) & (!g968) & (!g969) & (g970) & (!g977) & (g972)) + ((g971) & (!g968) & (!g969) & (g970) & (g977) & (!g972)) + ((g971) & (!g968) & (g969) & (g970) & (!g977) & (!g972)) + ((g971) & (g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((g971) & (g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((g971) & (g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((g971) & (g968) & (!g969) & (g970) & (g977) & (!g972)) + ((g971) & (g968) & (!g969) & (g970) & (g977) & (g972)) + ((g971) & (g968) & (g969) & (!g970) & (!g977) & (!g972)) + ((g971) & (g968) & (g969) & (!g970) & (g977) & (!g972)) + ((g971) & (g968) & (g969) & (g970) & (!g977) & (g972)) + ((g971) & (g968) & (g969) & (g970) & (g977) & (g972)));
	assign g991 = (((!g971) & (!g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((!g971) & (!g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((!g971) & (!g968) & (!g969) & (g970) & (!g977) & (g972)) + ((!g971) & (!g968) & (g969) & (!g970) & (!g977) & (g972)) + ((!g971) & (!g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g971) & (!g968) & (g969) & (g970) & (!g977) & (g972)) + ((!g971) & (g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((!g971) & (g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((!g971) & (g968) & (!g969) & (g970) & (g977) & (!g972)) + ((!g971) & (g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g971) & (g968) & (g969) & (g970) & (!g977) & (!g972)) + ((!g971) & (g968) & (g969) & (g970) & (g977) & (!g972)) + ((g971) & (!g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((g971) & (!g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((g971) & (!g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((g971) & (!g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((g971) & (!g968) & (!g969) & (g970) & (!g977) & (g972)) + ((g971) & (!g968) & (!g969) & (g970) & (g977) & (!g972)) + ((g971) & (!g968) & (!g969) & (g970) & (g977) & (g972)) + ((g971) & (!g968) & (g969) & (!g970) & (!g977) & (g972)) + ((g971) & (!g968) & (g969) & (!g970) & (g977) & (!g972)) + ((g971) & (!g968) & (g969) & (g970) & (!g977) & (!g972)) + ((g971) & (!g968) & (g969) & (g970) & (g977) & (g972)) + ((g971) & (g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((g971) & (g968) & (!g969) & (!g970) & (g977) & (g972)) + ((g971) & (g968) & (g969) & (!g970) & (g977) & (g972)) + ((g971) & (g968) & (g969) & (g970) & (!g977) & (!g972)) + ((g971) & (g968) & (g969) & (g970) & (!g977) & (g972)) + ((g971) & (g968) & (g969) & (g970) & (g977) & (g972)));
	assign g992 = (((!g971) & (!g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((!g971) & (!g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((!g971) & (!g968) & (!g969) & (!g970) & (g977) & (g972)) + ((!g971) & (!g968) & (!g969) & (g970) & (!g977) & (g972)) + ((!g971) & (!g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g971) & (!g968) & (g969) & (g970) & (g977) & (g972)) + ((!g971) & (g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((!g971) & (g968) & (!g969) & (g970) & (!g977) & (g972)) + ((!g971) & (g968) & (!g969) & (g970) & (g977) & (g972)) + ((!g971) & (g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g971) & (g968) & (g969) & (!g970) & (g977) & (g972)) + ((!g971) & (g968) & (g969) & (g970) & (!g977) & (!g972)) + ((!g971) & (g968) & (g969) & (g970) & (!g977) & (g972)) + ((!g971) & (g968) & (g969) & (g970) & (g977) & (!g972)) + ((!g971) & (g968) & (g969) & (g970) & (g977) & (g972)) + ((g971) & (!g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((g971) & (!g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((g971) & (!g968) & (!g969) & (!g970) & (g977) & (g972)) + ((g971) & (!g968) & (!g969) & (g970) & (g977) & (g972)) + ((g971) & (!g968) & (g969) & (!g970) & (!g977) & (g972)) + ((g971) & (!g968) & (g969) & (!g970) & (g977) & (!g972)) + ((g971) & (!g968) & (g969) & (g970) & (g977) & (!g972)) + ((g971) & (g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((g971) & (g968) & (!g969) & (g970) & (!g977) & (g972)) + ((g971) & (g968) & (!g969) & (g970) & (g977) & (!g972)) + ((g971) & (g968) & (g969) & (!g970) & (g977) & (g972)) + ((g971) & (g968) & (g969) & (g970) & (!g977) & (!g972)));
	assign g993 = (((!g989) & (!g990) & (!g991) & (!g992) & (!g967) & (g978)) + ((!g989) & (!g990) & (!g991) & (!g992) & (g967) & (!g978)) + ((!g989) & (!g990) & (!g991) & (!g992) & (g967) & (g978)) + ((!g989) & (!g990) & (!g991) & (g992) & (!g967) & (g978)) + ((!g989) & (!g990) & (!g991) & (g992) & (g967) & (!g978)) + ((!g989) & (!g990) & (g991) & (!g992) & (g967) & (!g978)) + ((!g989) & (!g990) & (g991) & (!g992) & (g967) & (g978)) + ((!g989) & (!g990) & (g991) & (g992) & (g967) & (!g978)) + ((!g989) & (g990) & (!g991) & (!g992) & (!g967) & (g978)) + ((!g989) & (g990) & (!g991) & (!g992) & (g967) & (g978)) + ((!g989) & (g990) & (!g991) & (g992) & (!g967) & (g978)) + ((!g989) & (g990) & (g991) & (!g992) & (g967) & (g978)) + ((g989) & (!g990) & (!g991) & (!g992) & (!g967) & (!g978)) + ((g989) & (!g990) & (!g991) & (!g992) & (!g967) & (g978)) + ((g989) & (!g990) & (!g991) & (!g992) & (g967) & (!g978)) + ((g989) & (!g990) & (!g991) & (!g992) & (g967) & (g978)) + ((g989) & (!g990) & (!g991) & (g992) & (!g967) & (!g978)) + ((g989) & (!g990) & (!g991) & (g992) & (!g967) & (g978)) + ((g989) & (!g990) & (!g991) & (g992) & (g967) & (!g978)) + ((g989) & (!g990) & (g991) & (!g992) & (!g967) & (!g978)) + ((g989) & (!g990) & (g991) & (!g992) & (g967) & (!g978)) + ((g989) & (!g990) & (g991) & (!g992) & (g967) & (g978)) + ((g989) & (!g990) & (g991) & (g992) & (!g967) & (!g978)) + ((g989) & (!g990) & (g991) & (g992) & (g967) & (!g978)) + ((g989) & (g990) & (!g991) & (!g992) & (!g967) & (!g978)) + ((g989) & (g990) & (!g991) & (!g992) & (!g967) & (g978)) + ((g989) & (g990) & (!g991) & (!g992) & (g967) & (g978)) + ((g989) & (g990) & (!g991) & (g992) & (!g967) & (!g978)) + ((g989) & (g990) & (!g991) & (g992) & (!g967) & (g978)) + ((g989) & (g990) & (g991) & (!g992) & (!g967) & (!g978)) + ((g989) & (g990) & (g991) & (!g992) & (g967) & (g978)) + ((g989) & (g990) & (g991) & (g992) & (!g967) & (!g978)));
	assign g995 = (((!g993) & (sk[2]) & (g994)) + ((g993) & (!sk[2]) & (!g994)) + ((g993) & (!sk[2]) & (g994)) + ((g993) & (sk[2]) & (!g994)));
	assign g996 = (((!g967) & (!g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (g977) & (g972)) + ((!g967) & (!g968) & (g969) & (g970) & (!g977) & (!g972)) + ((!g967) & (!g968) & (g969) & (g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (g969) & (g970) & (g977) & (g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (g968) & (g969) & (!g970) & (!g977) & (!g972)) + ((!g967) & (g968) & (g969) & (g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((g967) & (!g968) & (g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (g969) & (!g970) & (!g977) & (g972)) + ((g967) & (!g968) & (g969) & (!g970) & (g977) & (!g972)) + ((g967) & (!g968) & (g969) & (g970) & (!g977) & (g972)) + ((g967) & (g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((g967) & (g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((g967) & (g968) & (!g969) & (g970) & (g977) & (!g972)) + ((g967) & (g968) & (g969) & (!g970) & (!g977) & (g972)) + ((g967) & (g968) & (g969) & (!g970) & (g977) & (g972)));
	assign g997 = (((!g967) & (!g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (!g969) & (!g970) & (g977) & (g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (g969) & (g970) & (!g977) & (!g972)) + ((!g967) & (!g968) & (g969) & (g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (g969) & (g970) & (g977) & (g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (g977) & (g972)) + ((!g967) & (g968) & (!g969) & (g970) & (g977) & (g972)) + ((!g967) & (g968) & (g969) & (!g970) & (!g977) & (!g972)) + ((!g967) & (g968) & (g969) & (!g970) & (!g977) & (g972)) + ((!g967) & (g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (g968) & (g969) & (g970) & (!g977) & (g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((g967) & (!g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (!g969) & (g970) & (!g977) & (g972)) + ((g967) & (!g968) & (!g969) & (g970) & (g977) & (g972)) + ((g967) & (!g968) & (g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (g969) & (!g970) & (!g977) & (g972)) + ((g967) & (!g968) & (g969) & (!g970) & (g977) & (g972)) + ((g967) & (!g968) & (g969) & (g970) & (!g977) & (g972)) + ((g967) & (g968) & (!g969) & (g970) & (!g977) & (g972)) + ((g967) & (g968) & (!g969) & (g970) & (g977) & (!g972)) + ((g967) & (g968) & (g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (g968) & (g969) & (g970) & (!g977) & (!g972)));
	assign g998 = (((!g967) & (!g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (!g969) & (!g970) & (g977) & (g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (g969) & (!g970) & (g977) & (g972)) + ((!g967) & (!g968) & (g969) & (g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (g969) & (g970) & (g977) & (g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (g977) & (g972)) + ((!g967) & (g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((!g967) & (g968) & (!g969) & (g970) & (!g977) & (g972)) + ((!g967) & (g968) & (g969) & (!g970) & (!g977) & (g972)) + ((!g967) & (g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (g968) & (g969) & (g970) & (g977) & (g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (g977) & (g972)) + ((g967) & (!g968) & (!g969) & (g970) & (g977) & (g972)) + ((g967) & (!g968) & (g969) & (g970) & (!g977) & (!g972)) + ((g967) & (g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((g967) & (g968) & (!g969) & (g970) & (g977) & (g972)) + ((g967) & (g968) & (g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (g968) & (g969) & (!g970) & (!g977) & (g972)) + ((g967) & (g968) & (g969) & (!g970) & (g977) & (g972)) + ((g967) & (g968) & (g969) & (g970) & (!g977) & (!g972)) + ((g967) & (g968) & (g969) & (g970) & (g977) & (g972)));
	assign g999 = (((!g967) & (!g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (!g969) & (g970) & (g977) & (g972)) + ((!g967) & (!g968) & (g969) & (g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (g969) & (g970) & (g977) & (g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (!g977) & (!g972)) + ((!g967) & (g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (g968) & (!g969) & (g970) & (!g977) & (!g972)) + ((!g967) & (g968) & (!g969) & (g970) & (!g977) & (g972)) + ((!g967) & (g968) & (!g969) & (g970) & (g977) & (!g972)) + ((!g967) & (g968) & (g969) & (!g970) & (!g977) & (!g972)) + ((!g967) & (g968) & (g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (g968) & (g969) & (!g970) & (g977) & (g972)) + ((g967) & (!g968) & (!g969) & (!g970) & (g977) & (g972)) + ((g967) & (!g968) & (!g969) & (g970) & (g977) & (!g972)) + ((g967) & (!g968) & (g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (g969) & (!g970) & (g977) & (!g972)) + ((g967) & (!g968) & (g969) & (!g970) & (g977) & (g972)) + ((g967) & (!g968) & (g969) & (g970) & (!g977) & (g972)) + ((g967) & (!g968) & (g969) & (g970) & (g977) & (!g972)) + ((g967) & (!g968) & (g969) & (g970) & (g977) & (g972)) + ((g967) & (g968) & (!g969) & (!g970) & (!g977) & (g972)) + ((g967) & (g968) & (!g969) & (!g970) & (g977) & (!g972)) + ((g967) & (g968) & (g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (g968) & (g969) & (!g970) & (!g977) & (g972)) + ((g967) & (g968) & (g969) & (g970) & (g977) & (g972)));
	assign g1000 = (((!g996) & (!g997) & (!g998) & (!g999) & (!g978) & (g971)) + ((!g996) & (!g997) & (!g998) & (!g999) & (g978) & (!g971)) + ((!g996) & (!g997) & (!g998) & (!g999) & (g978) & (g971)) + ((!g996) & (!g997) & (!g998) & (g999) & (!g978) & (g971)) + ((!g996) & (!g997) & (!g998) & (g999) & (g978) & (!g971)) + ((!g996) & (!g997) & (g998) & (!g999) & (g978) & (!g971)) + ((!g996) & (!g997) & (g998) & (!g999) & (g978) & (g971)) + ((!g996) & (!g997) & (g998) & (g999) & (g978) & (!g971)) + ((!g996) & (g997) & (!g998) & (!g999) & (!g978) & (g971)) + ((!g996) & (g997) & (!g998) & (!g999) & (g978) & (g971)) + ((!g996) & (g997) & (!g998) & (g999) & (!g978) & (g971)) + ((!g996) & (g997) & (g998) & (!g999) & (g978) & (g971)) + ((g996) & (!g997) & (!g998) & (!g999) & (!g978) & (!g971)) + ((g996) & (!g997) & (!g998) & (!g999) & (!g978) & (g971)) + ((g996) & (!g997) & (!g998) & (!g999) & (g978) & (!g971)) + ((g996) & (!g997) & (!g998) & (!g999) & (g978) & (g971)) + ((g996) & (!g997) & (!g998) & (g999) & (!g978) & (!g971)) + ((g996) & (!g997) & (!g998) & (g999) & (!g978) & (g971)) + ((g996) & (!g997) & (!g998) & (g999) & (g978) & (!g971)) + ((g996) & (!g997) & (g998) & (!g999) & (!g978) & (!g971)) + ((g996) & (!g997) & (g998) & (!g999) & (g978) & (!g971)) + ((g996) & (!g997) & (g998) & (!g999) & (g978) & (g971)) + ((g996) & (!g997) & (g998) & (g999) & (!g978) & (!g971)) + ((g996) & (!g997) & (g998) & (g999) & (g978) & (!g971)) + ((g996) & (g997) & (!g998) & (!g999) & (!g978) & (!g971)) + ((g996) & (g997) & (!g998) & (!g999) & (!g978) & (g971)) + ((g996) & (g997) & (!g998) & (!g999) & (g978) & (g971)) + ((g996) & (g997) & (!g998) & (g999) & (!g978) & (!g971)) + ((g996) & (g997) & (!g998) & (g999) & (!g978) & (g971)) + ((g996) & (g997) & (g998) & (!g999) & (!g978) & (!g971)) + ((g996) & (g997) & (g998) & (!g999) & (g978) & (g971)) + ((g996) & (g997) & (g998) & (g999) & (!g978) & (!g971)));
	assign g1002 = (((!sk[8]) & (g1000) & (!g1001)) + ((!sk[8]) & (g1000) & (g1001)) + ((sk[8]) & (!g1000) & (g1001)) + ((sk[8]) & (g1000) & (!g1001)));
	assign g1003 = (((!g967) & (!g968) & (!g971) & (!g978) & (!g977) & (g972)) + ((!g967) & (!g968) & (g971) & (!g978) & (!g977) & (g972)) + ((!g967) & (!g968) & (g971) & (!g978) & (g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (!g978) & (g977) & (g972)) + ((!g967) & (!g968) & (g971) & (g978) & (!g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (g978) & (g977) & (!g972)) + ((!g967) & (g968) & (!g971) & (!g978) & (!g977) & (!g972)) + ((!g967) & (g968) & (!g971) & (!g978) & (!g977) & (g972)) + ((!g967) & (g968) & (!g971) & (g978) & (!g977) & (!g972)) + ((!g967) & (g968) & (!g971) & (g978) & (!g977) & (g972)) + ((!g967) & (g968) & (!g971) & (g978) & (g977) & (g972)) + ((!g967) & (g968) & (g971) & (g978) & (!g977) & (g972)) + ((!g967) & (g968) & (g971) & (g978) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g978) & (!g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g978) & (!g977) & (g972)) + ((g967) & (!g968) & (!g971) & (g978) & (!g977) & (g972)) + ((g967) & (!g968) & (g971) & (!g978) & (g977) & (!g972)) + ((g967) & (!g968) & (g971) & (g978) & (!g977) & (!g972)) + ((g967) & (!g968) & (g971) & (g978) & (!g977) & (g972)) + ((g967) & (!g968) & (g971) & (g978) & (g977) & (!g972)) + ((g967) & (g968) & (!g971) & (!g978) & (!g977) & (!g972)) + ((g967) & (g968) & (!g971) & (!g978) & (g977) & (!g972)) + ((g967) & (g968) & (!g971) & (g978) & (g977) & (!g972)) + ((g967) & (g968) & (g971) & (!g978) & (!g977) & (!g972)) + ((g967) & (g968) & (g971) & (!g978) & (!g977) & (g972)) + ((g967) & (g968) & (g971) & (g978) & (!g977) & (g972)));
	assign g1004 = (((!g967) & (!g968) & (!g971) & (!g978) & (!g977) & (!g972)) + ((!g967) & (!g968) & (!g971) & (!g978) & (!g977) & (g972)) + ((!g967) & (!g968) & (!g971) & (!g978) & (g977) & (!g972)) + ((!g967) & (!g968) & (!g971) & (!g978) & (g977) & (g972)) + ((!g967) & (!g968) & (!g971) & (g978) & (!g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (!g978) & (!g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (!g978) & (g977) & (g972)) + ((!g967) & (!g968) & (g971) & (g978) & (!g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (g978) & (g977) & (g972)) + ((!g967) & (g968) & (!g971) & (!g978) & (!g977) & (g972)) + ((!g967) & (g968) & (!g971) & (g978) & (g977) & (!g972)) + ((!g967) & (g968) & (g971) & (!g978) & (!g977) & (!g972)) + ((!g967) & (g968) & (g971) & (!g978) & (!g977) & (g972)) + ((!g967) & (g968) & (g971) & (!g978) & (g977) & (!g972)) + ((!g967) & (g968) & (g971) & (!g978) & (g977) & (g972)) + ((!g967) & (g968) & (g971) & (g978) & (!g977) & (!g972)) + ((!g967) & (g968) & (g971) & (g978) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g978) & (!g977) & (g972)) + ((g967) & (!g968) & (!g971) & (!g978) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g978) & (g977) & (g972)) + ((g967) & (!g968) & (!g971) & (g978) & (!g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (g978) & (g977) & (g972)) + ((g967) & (!g968) & (g971) & (!g978) & (g977) & (!g972)) + ((g967) & (!g968) & (g971) & (!g978) & (g977) & (g972)) + ((g967) & (!g968) & (g971) & (g978) & (!g977) & (g972)) + ((g967) & (g968) & (!g971) & (!g978) & (g977) & (!g972)) + ((g967) & (g968) & (!g971) & (!g978) & (g977) & (g972)) + ((g967) & (g968) & (!g971) & (g978) & (!g977) & (!g972)) + ((g967) & (g968) & (!g971) & (g978) & (!g977) & (g972)) + ((g967) & (g968) & (g971) & (!g978) & (g977) & (!g972)) + ((g967) & (g968) & (g971) & (!g978) & (g977) & (g972)) + ((g967) & (g968) & (g971) & (g978) & (!g977) & (g972)));
	assign g1005 = (((!g967) & (!g968) & (!g971) & (!g978) & (!g977) & (!g972)) + ((!g967) & (!g968) & (!g971) & (!g978) & (!g977) & (g972)) + ((!g967) & (!g968) & (g971) & (!g978) & (!g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (!g978) & (g977) & (g972)) + ((!g967) & (!g968) & (g971) & (g978) & (!g977) & (g972)) + ((!g967) & (g968) & (!g971) & (g978) & (!g977) & (!g972)) + ((!g967) & (g968) & (!g971) & (g978) & (g977) & (!g972)) + ((!g967) & (g968) & (!g971) & (g978) & (g977) & (g972)) + ((!g967) & (g968) & (g971) & (!g978) & (!g977) & (!g972)) + ((!g967) & (g968) & (g971) & (!g978) & (g977) & (!g972)) + ((!g967) & (g968) & (g971) & (!g978) & (g977) & (g972)) + ((!g967) & (g968) & (g971) & (g978) & (!g977) & (!g972)) + ((!g967) & (g968) & (g971) & (g978) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g978) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g978) & (g977) & (g972)) + ((g967) & (!g968) & (!g971) & (g978) & (!g977) & (g972)) + ((g967) & (!g968) & (!g971) & (g978) & (g977) & (g972)) + ((g967) & (!g968) & (g971) & (!g978) & (!g977) & (!g972)) + ((g967) & (!g968) & (g971) & (!g978) & (!g977) & (g972)) + ((g967) & (!g968) & (g971) & (!g978) & (g977) & (g972)) + ((g967) & (!g968) & (g971) & (g978) & (!g977) & (!g972)) + ((g967) & (!g968) & (g971) & (g978) & (!g977) & (g972)) + ((g967) & (!g968) & (g971) & (g978) & (g977) & (!g972)) + ((g967) & (!g968) & (g971) & (g978) & (g977) & (g972)) + ((g967) & (g968) & (!g971) & (!g978) & (!g977) & (g972)) + ((g967) & (g968) & (!g971) & (g978) & (!g977) & (!g972)) + ((g967) & (g968) & (!g971) & (g978) & (g977) & (!g972)) + ((g967) & (g968) & (g971) & (!g978) & (!g977) & (!g972)) + ((g967) & (g968) & (g971) & (!g978) & (!g977) & (g972)) + ((g967) & (g968) & (g971) & (!g978) & (g977) & (!g972)) + ((g967) & (g968) & (g971) & (g978) & (!g977) & (!g972)) + ((g967) & (g968) & (g971) & (g978) & (g977) & (!g972)));
	assign g1006 = (((!g967) & (!g968) & (!g971) & (!g978) & (g977) & (g972)) + ((!g967) & (!g968) & (!g971) & (g978) & (!g977) & (!g972)) + ((!g967) & (!g968) & (!g971) & (g978) & (g977) & (g972)) + ((!g967) & (!g968) & (g971) & (!g978) & (!g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (!g978) & (g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (g978) & (!g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (g978) & (!g977) & (g972)) + ((!g967) & (!g968) & (g971) & (g978) & (g977) & (!g972)) + ((!g967) & (g968) & (!g971) & (!g978) & (!g977) & (!g972)) + ((!g967) & (g968) & (!g971) & (g978) & (!g977) & (g972)) + ((!g967) & (g968) & (!g971) & (g978) & (g977) & (!g972)) + ((!g967) & (g968) & (!g971) & (g978) & (g977) & (g972)) + ((!g967) & (g968) & (g971) & (!g978) & (!g977) & (!g972)) + ((!g967) & (g968) & (g971) & (g978) & (!g977) & (!g972)) + ((!g967) & (g968) & (g971) & (g978) & (!g977) & (g972)) + ((g967) & (!g968) & (!g971) & (!g978) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g978) & (g977) & (g972)) + ((g967) & (!g968) & (g971) & (!g978) & (!g977) & (!g972)) + ((g967) & (!g968) & (g971) & (!g978) & (g977) & (!g972)) + ((g967) & (!g968) & (g971) & (g978) & (g977) & (!g972)) + ((g967) & (g968) & (!g971) & (!g978) & (g977) & (!g972)) + ((g967) & (g968) & (!g971) & (g978) & (g977) & (g972)) + ((g967) & (g968) & (g971) & (!g978) & (!g977) & (!g972)) + ((g967) & (g968) & (g971) & (!g978) & (!g977) & (g972)) + ((g967) & (g968) & (g971) & (!g978) & (g977) & (!g972)) + ((g967) & (g968) & (g971) & (g978) & (!g977) & (!g972)));
	assign g1007 = (((!g1003) & (!g1004) & (!g1005) & (!g1006) & (g969) & (g970)) + ((!g1003) & (!g1004) & (g1005) & (!g1006) & (!g969) & (g970)) + ((!g1003) & (!g1004) & (g1005) & (!g1006) & (g969) & (g970)) + ((!g1003) & (!g1004) & (g1005) & (g1006) & (!g969) & (g970)) + ((!g1003) & (g1004) & (!g1005) & (!g1006) & (g969) & (!g970)) + ((!g1003) & (g1004) & (!g1005) & (!g1006) & (g969) & (g970)) + ((!g1003) & (g1004) & (!g1005) & (g1006) & (g969) & (!g970)) + ((!g1003) & (g1004) & (g1005) & (!g1006) & (!g969) & (g970)) + ((!g1003) & (g1004) & (g1005) & (!g1006) & (g969) & (!g970)) + ((!g1003) & (g1004) & (g1005) & (!g1006) & (g969) & (g970)) + ((!g1003) & (g1004) & (g1005) & (g1006) & (!g969) & (g970)) + ((!g1003) & (g1004) & (g1005) & (g1006) & (g969) & (!g970)) + ((g1003) & (!g1004) & (!g1005) & (!g1006) & (!g969) & (!g970)) + ((g1003) & (!g1004) & (!g1005) & (!g1006) & (g969) & (g970)) + ((g1003) & (!g1004) & (!g1005) & (g1006) & (!g969) & (!g970)) + ((g1003) & (!g1004) & (g1005) & (!g1006) & (!g969) & (!g970)) + ((g1003) & (!g1004) & (g1005) & (!g1006) & (!g969) & (g970)) + ((g1003) & (!g1004) & (g1005) & (!g1006) & (g969) & (g970)) + ((g1003) & (!g1004) & (g1005) & (g1006) & (!g969) & (!g970)) + ((g1003) & (!g1004) & (g1005) & (g1006) & (!g969) & (g970)) + ((g1003) & (g1004) & (!g1005) & (!g1006) & (!g969) & (!g970)) + ((g1003) & (g1004) & (!g1005) & (!g1006) & (g969) & (!g970)) + ((g1003) & (g1004) & (!g1005) & (!g1006) & (g969) & (g970)) + ((g1003) & (g1004) & (!g1005) & (g1006) & (!g969) & (!g970)) + ((g1003) & (g1004) & (!g1005) & (g1006) & (g969) & (!g970)) + ((g1003) & (g1004) & (g1005) & (!g1006) & (!g969) & (!g970)) + ((g1003) & (g1004) & (g1005) & (!g1006) & (!g969) & (g970)) + ((g1003) & (g1004) & (g1005) & (!g1006) & (g969) & (!g970)) + ((g1003) & (g1004) & (g1005) & (!g1006) & (g969) & (g970)) + ((g1003) & (g1004) & (g1005) & (g1006) & (!g969) & (!g970)) + ((g1003) & (g1004) & (g1005) & (g1006) & (!g969) & (g970)) + ((g1003) & (g1004) & (g1005) & (g1006) & (g969) & (!g970)));
	assign g1009 = (((!g1007) & (sk[14]) & (g1008)) + ((g1007) & (!sk[14]) & (!g1008)) + ((g1007) & (!sk[14]) & (g1008)) + ((g1007) & (sk[14]) & (!g1008)));
	assign g1010 = (((!g967) & (!g968) & (!g971) & (!g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (!g971) & (!g970) & (g977) & (g972)) + ((!g967) & (!g968) & (!g971) & (g970) & (g977) & (g972)) + ((!g967) & (!g968) & (g971) & (!g970) & (!g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (!g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (g971) & (!g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (!g970) & (g977) & (g972)) + ((!g967) & (!g968) & (g971) & (g970) & (!g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (g970) & (!g977) & (g972)) + ((!g967) & (g968) & (!g971) & (!g970) & (!g977) & (g972)) + ((!g967) & (g968) & (!g971) & (!g970) & (g977) & (!g972)) + ((!g967) & (g968) & (!g971) & (g970) & (g977) & (g972)) + ((!g967) & (g968) & (g971) & (!g970) & (g977) & (!g972)) + ((!g967) & (g968) & (g971) & (!g970) & (g977) & (g972)) + ((!g967) & (g968) & (g971) & (g970) & (!g977) & (!g972)) + ((!g967) & (g968) & (g971) & (g970) & (!g977) & (g972)) + ((!g967) & (g968) & (g971) & (g970) & (g977) & (g972)) + ((g967) & (!g968) & (!g971) & (!g970) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g970) & (g977) & (g972)) + ((g967) & (!g968) & (!g971) & (g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (g970) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (g970) & (g977) & (g972)) + ((g967) & (!g968) & (g971) & (!g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (g971) & (!g970) & (g977) & (!g972)) + ((g967) & (!g968) & (g971) & (g970) & (g977) & (!g972)) + ((g967) & (g968) & (!g971) & (!g970) & (g977) & (g972)) + ((g967) & (g968) & (g971) & (!g970) & (!g977) & (!g972)) + ((g967) & (g968) & (g971) & (!g970) & (g977) & (g972)));
	assign g1011 = (((!g967) & (!g968) & (!g971) & (!g970) & (!g977) & (!g972)) + ((!g967) & (!g968) & (!g971) & (g970) & (!g977) & (!g972)) + ((!g967) & (!g968) & (!g971) & (g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (!g971) & (g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (!g970) & (g977) & (g972)) + ((!g967) & (!g968) & (g971) & (g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (g971) & (g970) & (g977) & (g972)) + ((!g967) & (g968) & (!g971) & (!g970) & (!g977) & (!g972)) + ((!g967) & (g968) & (!g971) & (!g970) & (g977) & (!g972)) + ((!g967) & (g968) & (g971) & (!g970) & (!g977) & (g972)) + ((!g967) & (g968) & (g971) & (!g970) & (g977) & (g972)) + ((!g967) & (g968) & (g971) & (g970) & (!g977) & (g972)) + ((!g967) & (g968) & (g971) & (g970) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g970) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g970) & (g977) & (g972)) + ((g967) & (!g968) & (!g971) & (g970) & (!g977) & (g972)) + ((g967) & (!g968) & (!g971) & (g970) & (g977) & (g972)) + ((g967) & (!g968) & (g971) & (g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (g971) & (g970) & (!g977) & (g972)) + ((g967) & (!g968) & (g971) & (g970) & (g977) & (g972)) + ((g967) & (g968) & (!g971) & (!g970) & (!g977) & (g972)) + ((g967) & (g968) & (!g971) & (!g970) & (g977) & (!g972)) + ((g967) & (g968) & (!g971) & (g970) & (g977) & (!g972)) + ((g967) & (g968) & (g971) & (!g970) & (!g977) & (g972)) + ((g967) & (g968) & (g971) & (!g970) & (g977) & (g972)) + ((g967) & (g968) & (g971) & (g970) & (!g977) & (!g972)) + ((g967) & (g968) & (g971) & (g970) & (g977) & (g972)));
	assign g1012 = (((!g967) & (!g968) & (!g971) & (!g970) & (g977) & (g972)) + ((!g967) & (!g968) & (!g971) & (g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (!g970) & (!g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (!g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (g971) & (!g970) & (g977) & (g972)) + ((!g967) & (!g968) & (g971) & (g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (g971) & (g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (g971) & (g970) & (g977) & (g972)) + ((!g967) & (g968) & (!g971) & (!g970) & (g977) & (!g972)) + ((!g967) & (g968) & (!g971) & (!g970) & (g977) & (g972)) + ((!g967) & (g968) & (g971) & (!g970) & (!g977) & (!g972)) + ((!g967) & (g968) & (g971) & (g970) & (!g977) & (g972)) + ((!g967) & (g968) & (g971) & (g970) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g970) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (!g970) & (g977) & (g972)) + ((g967) & (!g968) & (!g971) & (g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (g970) & (!g977) & (g972)) + ((g967) & (!g968) & (g971) & (!g970) & (!g977) & (g972)) + ((g967) & (!g968) & (g971) & (!g970) & (g977) & (g972)) + ((g967) & (!g968) & (g971) & (g970) & (g977) & (!g972)) + ((g967) & (g968) & (!g971) & (!g970) & (!g977) & (!g972)) + ((g967) & (g968) & (!g971) & (!g970) & (!g977) & (g972)) + ((g967) & (g968) & (!g971) & (!g970) & (g977) & (g972)) + ((g967) & (g968) & (!g971) & (g970) & (!g977) & (g972)) + ((g967) & (g968) & (!g971) & (g970) & (g977) & (!g972)) + ((g967) & (g968) & (g971) & (!g970) & (!g977) & (g972)) + ((g967) & (g968) & (g971) & (!g970) & (g977) & (!g972)) + ((g967) & (g968) & (g971) & (g970) & (!g977) & (!g972)) + ((g967) & (g968) & (g971) & (g970) & (g977) & (!g972)) + ((g967) & (g968) & (g971) & (g970) & (g977) & (g972)));
	assign g1013 = (((!g967) & (!g968) & (!g971) & (!g970) & (g977) & (!g972)) + ((!g967) & (!g968) & (!g971) & (g970) & (!g977) & (!g972)) + ((!g967) & (!g968) & (!g971) & (g970) & (g977) & (g972)) + ((!g967) & (!g968) & (g971) & (!g970) & (!g977) & (g972)) + ((!g967) & (!g968) & (g971) & (!g970) & (g977) & (g972)) + ((!g967) & (!g968) & (g971) & (g970) & (g977) & (g972)) + ((!g967) & (g968) & (!g971) & (!g970) & (!g977) & (g972)) + ((!g967) & (g968) & (!g971) & (g970) & (!g977) & (g972)) + ((!g967) & (g968) & (!g971) & (g970) & (g977) & (g972)) + ((!g967) & (g968) & (g971) & (!g970) & (!g977) & (!g972)) + ((!g967) & (g968) & (g971) & (!g970) & (g977) & (!g972)) + ((!g967) & (g968) & (g971) & (g970) & (!g977) & (g972)) + ((!g967) & (g968) & (g971) & (g970) & (g977) & (g972)) + ((g967) & (!g968) & (!g971) & (!g970) & (g977) & (!g972)) + ((g967) & (!g968) & (!g971) & (g970) & (g977) & (g972)) + ((g967) & (!g968) & (g971) & (!g970) & (!g977) & (!g972)) + ((g967) & (!g968) & (g971) & (!g970) & (g977) & (g972)) + ((g967) & (!g968) & (g971) & (g970) & (!g977) & (!g972)) + ((g967) & (g968) & (!g971) & (!g970) & (g977) & (g972)) + ((g967) & (g968) & (!g971) & (g970) & (!g977) & (!g972)) + ((g967) & (g968) & (!g971) & (g970) & (!g977) & (g972)) + ((g967) & (g968) & (g971) & (!g970) & (g977) & (g972)));
	assign g1014 = (((!g1010) & (!g1011) & (!g1012) & (!g1013) & (!g978) & (!g969)) + ((!g1010) & (!g1011) & (!g1012) & (!g1013) & (!g978) & (g969)) + ((!g1010) & (!g1011) & (!g1012) & (!g1013) & (g978) & (!g969)) + ((!g1010) & (!g1011) & (!g1012) & (g1013) & (!g978) & (!g969)) + ((!g1010) & (!g1011) & (!g1012) & (g1013) & (!g978) & (g969)) + ((!g1010) & (!g1011) & (!g1012) & (g1013) & (g978) & (!g969)) + ((!g1010) & (!g1011) & (!g1012) & (g1013) & (g978) & (g969)) + ((!g1010) & (!g1011) & (g1012) & (!g1013) & (!g978) & (!g969)) + ((!g1010) & (!g1011) & (g1012) & (!g1013) & (g978) & (!g969)) + ((!g1010) & (!g1011) & (g1012) & (g1013) & (!g978) & (!g969)) + ((!g1010) & (!g1011) & (g1012) & (g1013) & (g978) & (!g969)) + ((!g1010) & (!g1011) & (g1012) & (g1013) & (g978) & (g969)) + ((!g1010) & (g1011) & (!g1012) & (!g1013) & (!g978) & (!g969)) + ((!g1010) & (g1011) & (!g1012) & (!g1013) & (!g978) & (g969)) + ((!g1010) & (g1011) & (!g1012) & (g1013) & (!g978) & (!g969)) + ((!g1010) & (g1011) & (!g1012) & (g1013) & (!g978) & (g969)) + ((!g1010) & (g1011) & (!g1012) & (g1013) & (g978) & (g969)) + ((!g1010) & (g1011) & (g1012) & (!g1013) & (!g978) & (!g969)) + ((!g1010) & (g1011) & (g1012) & (g1013) & (!g978) & (!g969)) + ((!g1010) & (g1011) & (g1012) & (g1013) & (g978) & (g969)) + ((g1010) & (!g1011) & (!g1012) & (!g1013) & (!g978) & (g969)) + ((g1010) & (!g1011) & (!g1012) & (!g1013) & (g978) & (!g969)) + ((g1010) & (!g1011) & (!g1012) & (g1013) & (!g978) & (g969)) + ((g1010) & (!g1011) & (!g1012) & (g1013) & (g978) & (!g969)) + ((g1010) & (!g1011) & (!g1012) & (g1013) & (g978) & (g969)) + ((g1010) & (!g1011) & (g1012) & (!g1013) & (g978) & (!g969)) + ((g1010) & (!g1011) & (g1012) & (g1013) & (g978) & (!g969)) + ((g1010) & (!g1011) & (g1012) & (g1013) & (g978) & (g969)) + ((g1010) & (g1011) & (!g1012) & (!g1013) & (!g978) & (g969)) + ((g1010) & (g1011) & (!g1012) & (g1013) & (!g978) & (g969)) + ((g1010) & (g1011) & (!g1012) & (g1013) & (g978) & (g969)) + ((g1010) & (g1011) & (g1012) & (g1013) & (g978) & (g969)));
	assign g1016 = (((!sk[20]) & (g1014) & (!g1015)) + ((!sk[20]) & (g1014) & (g1015)) + ((sk[20]) & (!g1014) & (g1015)) + ((sk[20]) & (g1014) & (!g1015)));
	assign g1017 = (((!g967) & (!g978) & (!g969) & (!g970) & (!g977) & (g972)) + ((!g967) & (!g978) & (!g969) & (!g970) & (g977) & (g972)) + ((!g967) & (!g978) & (!g969) & (g970) & (!g977) & (!g972)) + ((!g967) & (!g978) & (!g969) & (g970) & (!g977) & (g972)) + ((!g967) & (!g978) & (!g969) & (g970) & (g977) & (!g972)) + ((!g967) & (!g978) & (!g969) & (g970) & (g977) & (g972)) + ((!g967) & (!g978) & (g969) & (!g970) & (!g977) & (g972)) + ((!g967) & (!g978) & (g969) & (!g970) & (g977) & (g972)) + ((!g967) & (!g978) & (g969) & (g970) & (g977) & (!g972)) + ((!g967) & (g978) & (g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (g978) & (g969) & (!g970) & (g977) & (g972)) + ((!g967) & (g978) & (g969) & (g970) & (!g977) & (g972)) + ((g967) & (!g978) & (!g969) & (!g970) & (g977) & (!g972)) + ((g967) & (!g978) & (!g969) & (g970) & (!g977) & (!g972)) + ((g967) & (!g978) & (!g969) & (g970) & (!g977) & (g972)) + ((g967) & (!g978) & (!g969) & (g970) & (g977) & (g972)) + ((g967) & (!g978) & (g969) & (!g970) & (!g977) & (g972)) + ((g967) & (!g978) & (g969) & (!g970) & (g977) & (g972)) + ((g967) & (!g978) & (g969) & (g970) & (g977) & (!g972)) + ((g967) & (!g978) & (g969) & (g970) & (g977) & (g972)) + ((g967) & (g978) & (!g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (g978) & (!g969) & (!g970) & (!g977) & (g972)) + ((g967) & (g978) & (!g969) & (!g970) & (g977) & (!g972)) + ((g967) & (g978) & (!g969) & (g970) & (!g977) & (!g972)) + ((g967) & (g978) & (g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (g978) & (g969) & (!g970) & (!g977) & (g972)) + ((g967) & (g978) & (g969) & (!g970) & (g977) & (!g972)) + ((g967) & (g978) & (g969) & (g970) & (!g977) & (g972)));
	assign g1018 = (((!g967) & (!g978) & (!g969) & (!g970) & (!g977) & (!g972)) + ((!g967) & (!g978) & (!g969) & (g970) & (g977) & (g972)) + ((!g967) & (!g978) & (g969) & (!g970) & (!g977) & (!g972)) + ((!g967) & (!g978) & (g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (!g978) & (g969) & (!g970) & (g977) & (g972)) + ((!g967) & (!g978) & (g969) & (g970) & (!g977) & (!g972)) + ((!g967) & (!g978) & (g969) & (g970) & (g977) & (g972)) + ((!g967) & (g978) & (!g969) & (!g970) & (!g977) & (!g972)) + ((!g967) & (g978) & (!g969) & (!g970) & (g977) & (g972)) + ((!g967) & (g978) & (!g969) & (g970) & (!g977) & (g972)) + ((!g967) & (g978) & (g969) & (!g970) & (!g977) & (!g972)) + ((!g967) & (g978) & (g969) & (!g970) & (g977) & (g972)) + ((!g967) & (g978) & (g969) & (g970) & (g977) & (!g972)) + ((!g967) & (g978) & (g969) & (g970) & (g977) & (g972)) + ((g967) & (!g978) & (!g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (!g978) & (!g969) & (!g970) & (g977) & (g972)) + ((g967) & (!g978) & (!g969) & (g970) & (!g977) & (!g972)) + ((g967) & (!g978) & (!g969) & (g970) & (g977) & (g972)) + ((g967) & (!g978) & (g969) & (!g970) & (g977) & (g972)) + ((g967) & (!g978) & (g969) & (g970) & (!g977) & (g972)) + ((g967) & (g978) & (!g969) & (!g970) & (g977) & (!g972)) + ((g967) & (g978) & (!g969) & (!g970) & (g977) & (g972)) + ((g967) & (g978) & (!g969) & (g970) & (!g977) & (g972)) + ((g967) & (g978) & (!g969) & (g970) & (g977) & (!g972)) + ((g967) & (g978) & (!g969) & (g970) & (g977) & (g972)) + ((g967) & (g978) & (g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (g978) & (g969) & (!g970) & (g977) & (!g972)) + ((g967) & (g978) & (g969) & (g970) & (!g977) & (!g972)));
	assign g1019 = (((!g967) & (!g978) & (!g969) & (!g970) & (!g977) & (g972)) + ((!g967) & (!g978) & (!g969) & (!g970) & (g977) & (g972)) + ((!g967) & (!g978) & (!g969) & (g970) & (g977) & (!g972)) + ((!g967) & (!g978) & (!g969) & (g970) & (g977) & (g972)) + ((!g967) & (!g978) & (g969) & (!g970) & (g977) & (g972)) + ((!g967) & (!g978) & (g969) & (g970) & (!g977) & (!g972)) + ((!g967) & (!g978) & (g969) & (g970) & (!g977) & (g972)) + ((!g967) & (!g978) & (g969) & (g970) & (g977) & (g972)) + ((!g967) & (g978) & (!g969) & (!g970) & (!g977) & (!g972)) + ((!g967) & (g978) & (!g969) & (!g970) & (!g977) & (g972)) + ((!g967) & (g978) & (!g969) & (!g970) & (g977) & (g972)) + ((!g967) & (g978) & (!g969) & (g970) & (!g977) & (g972)) + ((!g967) & (g978) & (!g969) & (g970) & (g977) & (!g972)) + ((!g967) & (g978) & (g969) & (!g970) & (!g977) & (g972)) + ((!g967) & (g978) & (g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (g978) & (g969) & (g970) & (!g977) & (!g972)) + ((!g967) & (g978) & (g969) & (g970) & (g977) & (!g972)) + ((!g967) & (g978) & (g969) & (g970) & (g977) & (g972)) + ((g967) & (!g978) & (!g969) & (!g970) & (!g977) & (g972)) + ((g967) & (!g978) & (!g969) & (g970) & (!g977) & (!g972)) + ((g967) & (!g978) & (!g969) & (g970) & (g977) & (!g972)) + ((g967) & (!g978) & (g969) & (!g970) & (g977) & (g972)) + ((g967) & (!g978) & (g969) & (g970) & (!g977) & (g972)) + ((g967) & (g978) & (!g969) & (!g970) & (!g977) & (g972)) + ((g967) & (g978) & (!g969) & (g970) & (!g977) & (!g972)) + ((g967) & (g978) & (!g969) & (g970) & (g977) & (!g972)) + ((g967) & (g978) & (g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (g978) & (g969) & (!g970) & (g977) & (!g972)) + ((g967) & (g978) & (g969) & (!g970) & (g977) & (g972)) + ((g967) & (g978) & (g969) & (g970) & (g977) & (g972)));
	assign g1020 = (((!g967) & (!g978) & (!g969) & (!g970) & (g977) & (g972)) + ((!g967) & (!g978) & (!g969) & (g970) & (!g977) & (!g972)) + ((!g967) & (!g978) & (!g969) & (g970) & (g977) & (g972)) + ((!g967) & (!g978) & (g969) & (!g970) & (!g977) & (!g972)) + ((!g967) & (!g978) & (g969) & (g970) & (g977) & (!g972)) + ((!g967) & (!g978) & (g969) & (g970) & (g977) & (g972)) + ((!g967) & (g978) & (!g969) & (g970) & (!g977) & (!g972)) + ((!g967) & (g978) & (!g969) & (g970) & (g977) & (!g972)) + ((!g967) & (g978) & (g969) & (!g970) & (g977) & (!g972)) + ((!g967) & (g978) & (g969) & (!g970) & (g977) & (g972)) + ((g967) & (!g978) & (!g969) & (!g970) & (!g977) & (g972)) + ((g967) & (!g978) & (!g969) & (!g970) & (g977) & (!g972)) + ((g967) & (!g978) & (!g969) & (g970) & (!g977) & (g972)) + ((g967) & (!g978) & (g969) & (!g970) & (g977) & (!g972)) + ((g967) & (!g978) & (g969) & (!g970) & (g977) & (g972)) + ((g967) & (!g978) & (g969) & (g970) & (g977) & (!g972)) + ((g967) & (!g978) & (g969) & (g970) & (g977) & (g972)) + ((g967) & (g978) & (!g969) & (!g970) & (g977) & (!g972)) + ((g967) & (g978) & (!g969) & (g970) & (!g977) & (g972)) + ((g967) & (g978) & (g969) & (!g970) & (!g977) & (!g972)) + ((g967) & (g978) & (g969) & (!g970) & (g977) & (g972)) + ((g967) & (g978) & (g969) & (g970) & (!g977) & (g972)));
	assign g1021 = (((!g1017) & (!g1018) & (!g1019) & (!g1020) & (!g971) & (!g968)) + ((!g1017) & (!g1018) & (!g1019) & (!g1020) & (!g971) & (g968)) + ((!g1017) & (!g1018) & (!g1019) & (!g1020) & (g971) & (!g968)) + ((!g1017) & (!g1018) & (!g1019) & (g1020) & (!g971) & (!g968)) + ((!g1017) & (!g1018) & (!g1019) & (g1020) & (!g971) & (g968)) + ((!g1017) & (!g1018) & (!g1019) & (g1020) & (g971) & (!g968)) + ((!g1017) & (!g1018) & (!g1019) & (g1020) & (g971) & (g968)) + ((!g1017) & (!g1018) & (g1019) & (!g1020) & (!g971) & (!g968)) + ((!g1017) & (!g1018) & (g1019) & (!g1020) & (g971) & (!g968)) + ((!g1017) & (!g1018) & (g1019) & (g1020) & (!g971) & (!g968)) + ((!g1017) & (!g1018) & (g1019) & (g1020) & (g971) & (!g968)) + ((!g1017) & (!g1018) & (g1019) & (g1020) & (g971) & (g968)) + ((!g1017) & (g1018) & (!g1019) & (!g1020) & (!g971) & (!g968)) + ((!g1017) & (g1018) & (!g1019) & (!g1020) & (!g971) & (g968)) + ((!g1017) & (g1018) & (!g1019) & (g1020) & (!g971) & (!g968)) + ((!g1017) & (g1018) & (!g1019) & (g1020) & (!g971) & (g968)) + ((!g1017) & (g1018) & (!g1019) & (g1020) & (g971) & (g968)) + ((!g1017) & (g1018) & (g1019) & (!g1020) & (!g971) & (!g968)) + ((!g1017) & (g1018) & (g1019) & (g1020) & (!g971) & (!g968)) + ((!g1017) & (g1018) & (g1019) & (g1020) & (g971) & (g968)) + ((g1017) & (!g1018) & (!g1019) & (!g1020) & (!g971) & (g968)) + ((g1017) & (!g1018) & (!g1019) & (!g1020) & (g971) & (!g968)) + ((g1017) & (!g1018) & (!g1019) & (g1020) & (!g971) & (g968)) + ((g1017) & (!g1018) & (!g1019) & (g1020) & (g971) & (!g968)) + ((g1017) & (!g1018) & (!g1019) & (g1020) & (g971) & (g968)) + ((g1017) & (!g1018) & (g1019) & (!g1020) & (g971) & (!g968)) + ((g1017) & (!g1018) & (g1019) & (g1020) & (g971) & (!g968)) + ((g1017) & (!g1018) & (g1019) & (g1020) & (g971) & (g968)) + ((g1017) & (g1018) & (!g1019) & (!g1020) & (!g971) & (g968)) + ((g1017) & (g1018) & (!g1019) & (g1020) & (!g971) & (g968)) + ((g1017) & (g1018) & (!g1019) & (g1020) & (g971) & (g968)) + ((g1017) & (g1018) & (g1019) & (g1020) & (g971) & (g968)));
	assign g1023 = (((!g1021) & (sk[26]) & (g1022)) + ((g1021) & (!sk[26]) & (!g1022)) + ((g1021) & (!sk[26]) & (g1022)) + ((g1021) & (sk[26]) & (!g1022)));
	assign g1024 = (((!g971) & (!g968) & (!g969) & (!g970) & (!g977) & (g978)) + ((!g971) & (!g968) & (!g969) & (!g970) & (g977) & (!g978)) + ((!g971) & (!g968) & (!g969) & (g970) & (!g977) & (g978)) + ((!g971) & (!g968) & (!g969) & (g970) & (g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (!g970) & (!g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (!g970) & (g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (g970) & (!g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (g970) & (g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (g970) & (g977) & (g978)) + ((!g971) & (g968) & (!g969) & (!g970) & (g977) & (!g978)) + ((!g971) & (g968) & (!g969) & (g970) & (g977) & (!g978)) + ((!g971) & (g968) & (!g969) & (g970) & (g977) & (g978)) + ((!g971) & (g968) & (g969) & (!g970) & (g977) & (g978)) + ((!g971) & (g968) & (g969) & (g970) & (!g977) & (!g978)) + ((g971) & (!g968) & (!g969) & (!g970) & (!g977) & (g978)) + ((g971) & (!g968) & (!g969) & (g970) & (!g977) & (g978)) + ((g971) & (!g968) & (g969) & (g970) & (g977) & (g978)) + ((g971) & (g968) & (!g969) & (!g970) & (g977) & (g978)) + ((g971) & (g968) & (!g969) & (g970) & (!g977) & (!g978)) + ((g971) & (g968) & (!g969) & (g970) & (g977) & (!g978)) + ((g971) & (g968) & (g969) & (!g970) & (!g977) & (g978)) + ((g971) & (g968) & (g969) & (!g970) & (g977) & (!g978)) + ((g971) & (g968) & (g969) & (!g970) & (g977) & (g978)) + ((g971) & (g968) & (g969) & (g970) & (!g977) & (g978)));
	assign g1025 = (((!g971) & (!g968) & (!g969) & (!g970) & (!g977) & (!g978)) + ((!g971) & (!g968) & (!g969) & (!g970) & (!g977) & (g978)) + ((!g971) & (!g968) & (!g969) & (g970) & (!g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (!g970) & (!g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (!g970) & (g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (!g970) & (g977) & (g978)) + ((!g971) & (!g968) & (g969) & (g970) & (!g977) & (g978)) + ((!g971) & (!g968) & (g969) & (g970) & (g977) & (g978)) + ((!g971) & (g968) & (!g969) & (!g970) & (!g977) & (!g978)) + ((!g971) & (g968) & (!g969) & (!g970) & (g977) & (!g978)) + ((!g971) & (g968) & (!g969) & (g970) & (!g977) & (!g978)) + ((!g971) & (g968) & (!g969) & (g970) & (!g977) & (g978)) + ((!g971) & (g968) & (!g969) & (g970) & (g977) & (g978)) + ((!g971) & (g968) & (g969) & (!g970) & (!g977) & (g978)) + ((!g971) & (g968) & (g969) & (g970) & (!g977) & (!g978)) + ((!g971) & (g968) & (g969) & (g970) & (!g977) & (g978)) + ((g971) & (!g968) & (!g969) & (!g970) & (!g977) & (g978)) + ((g971) & (!g968) & (!g969) & (!g970) & (g977) & (g978)) + ((g971) & (!g968) & (!g969) & (g970) & (!g977) & (!g978)) + ((g971) & (!g968) & (!g969) & (g970) & (g977) & (g978)) + ((g971) & (!g968) & (g969) & (!g970) & (!g977) & (!g978)) + ((g971) & (!g968) & (g969) & (!g970) & (g977) & (g978)) + ((g971) & (!g968) & (g969) & (g970) & (g977) & (!g978)) + ((g971) & (g968) & (!g969) & (!g970) & (!g977) & (!g978)) + ((g971) & (g968) & (!g969) & (!g970) & (!g977) & (g978)) + ((g971) & (g968) & (!g969) & (!g970) & (g977) & (g978)) + ((g971) & (g968) & (!g969) & (g970) & (!g977) & (g978)) + ((g971) & (g968) & (!g969) & (g970) & (g977) & (!g978)) + ((g971) & (g968) & (g969) & (!g970) & (g977) & (!g978)) + ((g971) & (g968) & (g969) & (!g970) & (g977) & (g978)));
	assign g1026 = (((!g971) & (!g968) & (!g969) & (!g970) & (g977) & (!g978)) + ((!g971) & (!g968) & (!g969) & (g970) & (!g977) & (!g978)) + ((!g971) & (!g968) & (!g969) & (g970) & (g977) & (!g978)) + ((!g971) & (!g968) & (!g969) & (g970) & (g977) & (g978)) + ((!g971) & (!g968) & (g969) & (!g970) & (!g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (!g970) & (!g977) & (g978)) + ((!g971) & (!g968) & (g969) & (!g970) & (g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (g970) & (!g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (g970) & (g977) & (g978)) + ((!g971) & (g968) & (!g969) & (!g970) & (!g977) & (g978)) + ((!g971) & (g968) & (!g969) & (!g970) & (g977) & (!g978)) + ((!g971) & (g968) & (!g969) & (!g970) & (g977) & (g978)) + ((!g971) & (g968) & (g969) & (!g970) & (!g977) & (g978)) + ((!g971) & (g968) & (g969) & (!g970) & (g977) & (!g978)) + ((!g971) & (g968) & (g969) & (!g970) & (g977) & (g978)) + ((!g971) & (g968) & (g969) & (g970) & (!g977) & (!g978)) + ((g971) & (!g968) & (!g969) & (!g970) & (g977) & (!g978)) + ((g971) & (!g968) & (!g969) & (g970) & (!g977) & (!g978)) + ((g971) & (!g968) & (!g969) & (g970) & (g977) & (g978)) + ((g971) & (!g968) & (g969) & (!g970) & (!g977) & (!g978)) + ((g971) & (!g968) & (g969) & (!g970) & (!g977) & (g978)) + ((g971) & (!g968) & (g969) & (g970) & (!g977) & (!g978)) + ((g971) & (!g968) & (g969) & (g970) & (g977) & (!g978)) + ((g971) & (g968) & (!g969) & (!g970) & (g977) & (!g978)) + ((g971) & (g968) & (!g969) & (g970) & (!g977) & (!g978)) + ((g971) & (g968) & (!g969) & (g970) & (g977) & (g978)) + ((g971) & (g968) & (g969) & (!g970) & (!g977) & (!g978)) + ((g971) & (g968) & (g969) & (!g970) & (g977) & (!g978)) + ((g971) & (g968) & (g969) & (!g970) & (g977) & (g978)) + ((g971) & (g968) & (g969) & (g970) & (!g977) & (g978)));
	assign g1027 = (((!g971) & (!g968) & (!g969) & (!g970) & (!g977) & (g978)) + ((!g971) & (!g968) & (!g969) & (g970) & (g977) & (!g978)) + ((!g971) & (!g968) & (!g969) & (g970) & (g977) & (g978)) + ((!g971) & (!g968) & (g969) & (!g970) & (!g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (!g970) & (!g977) & (g978)) + ((!g971) & (!g968) & (g969) & (g970) & (g977) & (!g978)) + ((!g971) & (!g968) & (g969) & (g970) & (g977) & (g978)) + ((!g971) & (g968) & (!g969) & (!g970) & (!g977) & (!g978)) + ((!g971) & (g968) & (!g969) & (!g970) & (!g977) & (g978)) + ((!g971) & (g968) & (!g969) & (!g970) & (g977) & (g978)) + ((!g971) & (g968) & (!g969) & (g970) & (!g977) & (g978)) + ((!g971) & (g968) & (g969) & (!g970) & (!g977) & (g978)) + ((!g971) & (g968) & (g969) & (g970) & (!g977) & (!g978)) + ((!g971) & (g968) & (g969) & (g970) & (!g977) & (g978)) + ((!g971) & (g968) & (g969) & (g970) & (g977) & (!g978)) + ((!g971) & (g968) & (g969) & (g970) & (g977) & (g978)) + ((g971) & (!g968) & (!g969) & (g970) & (!g977) & (g978)) + ((g971) & (!g968) & (g969) & (!g970) & (!g977) & (!g978)) + ((g971) & (!g968) & (g969) & (g970) & (!g977) & (!g978)) + ((g971) & (!g968) & (g969) & (g970) & (!g977) & (g978)) + ((g971) & (!g968) & (g969) & (g970) & (g977) & (g978)) + ((g971) & (g968) & (!g969) & (!g970) & (!g977) & (g978)) + ((g971) & (g968) & (!g969) & (!g970) & (g977) & (g978)) + ((g971) & (g968) & (!g969) & (g970) & (!g977) & (!g978)) + ((g971) & (g968) & (!g969) & (g970) & (g977) & (!g978)) + ((g971) & (g968) & (!g969) & (g970) & (g977) & (g978)) + ((g971) & (g968) & (g969) & (!g970) & (g977) & (g978)) + ((g971) & (g968) & (g969) & (g970) & (g977) & (g978)));
	assign g1028 = (((!g1024) & (!g1025) & (!g1026) & (!g1027) & (!g967) & (g972)) + ((!g1024) & (!g1025) & (!g1026) & (!g1027) & (g967) & (!g972)) + ((!g1024) & (!g1025) & (!g1026) & (!g1027) & (g967) & (g972)) + ((!g1024) & (!g1025) & (!g1026) & (g1027) & (!g967) & (g972)) + ((!g1024) & (!g1025) & (!g1026) & (g1027) & (g967) & (!g972)) + ((!g1024) & (!g1025) & (g1026) & (!g1027) & (g967) & (!g972)) + ((!g1024) & (!g1025) & (g1026) & (!g1027) & (g967) & (g972)) + ((!g1024) & (!g1025) & (g1026) & (g1027) & (g967) & (!g972)) + ((!g1024) & (g1025) & (!g1026) & (!g1027) & (!g967) & (g972)) + ((!g1024) & (g1025) & (!g1026) & (!g1027) & (g967) & (g972)) + ((!g1024) & (g1025) & (!g1026) & (g1027) & (!g967) & (g972)) + ((!g1024) & (g1025) & (g1026) & (!g1027) & (g967) & (g972)) + ((g1024) & (!g1025) & (!g1026) & (!g1027) & (!g967) & (!g972)) + ((g1024) & (!g1025) & (!g1026) & (!g1027) & (!g967) & (g972)) + ((g1024) & (!g1025) & (!g1026) & (!g1027) & (g967) & (!g972)) + ((g1024) & (!g1025) & (!g1026) & (!g1027) & (g967) & (g972)) + ((g1024) & (!g1025) & (!g1026) & (g1027) & (!g967) & (!g972)) + ((g1024) & (!g1025) & (!g1026) & (g1027) & (!g967) & (g972)) + ((g1024) & (!g1025) & (!g1026) & (g1027) & (g967) & (!g972)) + ((g1024) & (!g1025) & (g1026) & (!g1027) & (!g967) & (!g972)) + ((g1024) & (!g1025) & (g1026) & (!g1027) & (g967) & (!g972)) + ((g1024) & (!g1025) & (g1026) & (!g1027) & (g967) & (g972)) + ((g1024) & (!g1025) & (g1026) & (g1027) & (!g967) & (!g972)) + ((g1024) & (!g1025) & (g1026) & (g1027) & (g967) & (!g972)) + ((g1024) & (g1025) & (!g1026) & (!g1027) & (!g967) & (!g972)) + ((g1024) & (g1025) & (!g1026) & (!g1027) & (!g967) & (g972)) + ((g1024) & (g1025) & (!g1026) & (!g1027) & (g967) & (g972)) + ((g1024) & (g1025) & (!g1026) & (g1027) & (!g967) & (!g972)) + ((g1024) & (g1025) & (!g1026) & (g1027) & (!g967) & (g972)) + ((g1024) & (g1025) & (g1026) & (!g1027) & (!g967) & (!g972)) + ((g1024) & (g1025) & (g1026) & (!g1027) & (g967) & (g972)) + ((g1024) & (g1025) & (g1026) & (g1027) & (!g967) & (!g972)));
	assign g1030 = (((!sk[32]) & (g1028) & (!g1029)) + ((!sk[32]) & (g1028) & (g1029)) + ((sk[32]) & (!g1028) & (g1029)) + ((sk[32]) & (g1028) & (!g1029)));
	assign g1037 = (((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1035) & (g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1035) & (!g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1035) & (g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (g1035) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (!g1035) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (!g1035) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1035) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (g1035) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1035) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1035) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (g1035) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (g1035) & (g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (g1035) & (!g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1035) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1035) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (!g1035) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (g1035) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (!g1035) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (g1035) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1035) & (g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (g1035) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1035) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (g1035) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (g1035) & (g1036)));
	assign g1038 = (((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1035) & (!g1036)) + ((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1035) & (g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1035) & (!g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1035) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1035) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (!g1035) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (!g1035) & (g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (!g1035) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (!g1035) & (g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (g1035) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (g1035) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1035) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (g1035) & (!g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (g1035) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (g1035) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (!g1035) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1035) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (!g1035) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (g1035) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (!g1035) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (!g1035) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (g1035) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (g1035) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (!g1035) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1035) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1035) & (g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (g1035) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (g1035) & (g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1035) & (g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (g1035) & (!g1036)));
	assign g1039 = (((!g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1035) & (!g1036)) + ((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1035) & (g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (g1035) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (!g1035) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (!g1035) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (g1035) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1035) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (g1035) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (!g1035) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1035) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (g1035) & (g1036)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (!g1035) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (g1035) & (!g1036)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (!g1035) & (!g1036)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (!g1035) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (g1035) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (!g1035) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1035) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (!g1035) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (!g1035) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (g1035) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (g1035) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (g1035) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (!g1035) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1035) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1035) & (g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1035) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1035) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1035) & (g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (g1035) & (g1036)));
	assign g1040 = (((!g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1035) & (g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (g1035) & (!g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (g1035) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (!g1035) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (g1035) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1035) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (!g1035) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (!g1035) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1035) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1035) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (g1035) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (g1035) & (g1036)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (!g1035) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (g1035) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (g1035) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1035) & (!g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (g1035) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (g1035) & (!g1036)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (g1035) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (!g1035) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1035) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (g1035) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (!g1035) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (g1035) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1035) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1035) & (g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1035) & (g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1035) & (!g1036)));
	assign g1043 = (((!g1037) & (!g1038) & (!g1039) & (!g1040) & (!g1041) & (!g1042)) + ((!g1037) & (!g1038) & (!g1039) & (g1040) & (!g1041) & (!g1042)) + ((!g1037) & (!g1038) & (!g1039) & (g1040) & (g1041) & (g1042)) + ((!g1037) & (!g1038) & (g1039) & (!g1040) & (!g1041) & (!g1042)) + ((!g1037) & (!g1038) & (g1039) & (!g1040) & (!g1041) & (g1042)) + ((!g1037) & (!g1038) & (g1039) & (g1040) & (!g1041) & (!g1042)) + ((!g1037) & (!g1038) & (g1039) & (g1040) & (!g1041) & (g1042)) + ((!g1037) & (!g1038) & (g1039) & (g1040) & (g1041) & (g1042)) + ((!g1037) & (g1038) & (!g1039) & (!g1040) & (!g1041) & (!g1042)) + ((!g1037) & (g1038) & (!g1039) & (!g1040) & (g1041) & (!g1042)) + ((!g1037) & (g1038) & (!g1039) & (g1040) & (!g1041) & (!g1042)) + ((!g1037) & (g1038) & (!g1039) & (g1040) & (g1041) & (!g1042)) + ((!g1037) & (g1038) & (!g1039) & (g1040) & (g1041) & (g1042)) + ((!g1037) & (g1038) & (g1039) & (!g1040) & (!g1041) & (!g1042)) + ((!g1037) & (g1038) & (g1039) & (!g1040) & (!g1041) & (g1042)) + ((!g1037) & (g1038) & (g1039) & (!g1040) & (g1041) & (!g1042)) + ((!g1037) & (g1038) & (g1039) & (g1040) & (!g1041) & (!g1042)) + ((!g1037) & (g1038) & (g1039) & (g1040) & (!g1041) & (g1042)) + ((!g1037) & (g1038) & (g1039) & (g1040) & (g1041) & (!g1042)) + ((!g1037) & (g1038) & (g1039) & (g1040) & (g1041) & (g1042)) + ((g1037) & (!g1038) & (!g1039) & (g1040) & (g1041) & (g1042)) + ((g1037) & (!g1038) & (g1039) & (!g1040) & (!g1041) & (g1042)) + ((g1037) & (!g1038) & (g1039) & (g1040) & (!g1041) & (g1042)) + ((g1037) & (!g1038) & (g1039) & (g1040) & (g1041) & (g1042)) + ((g1037) & (g1038) & (!g1039) & (!g1040) & (g1041) & (!g1042)) + ((g1037) & (g1038) & (!g1039) & (g1040) & (g1041) & (!g1042)) + ((g1037) & (g1038) & (!g1039) & (g1040) & (g1041) & (g1042)) + ((g1037) & (g1038) & (g1039) & (!g1040) & (!g1041) & (g1042)) + ((g1037) & (g1038) & (g1039) & (!g1040) & (g1041) & (!g1042)) + ((g1037) & (g1038) & (g1039) & (g1040) & (!g1041) & (g1042)) + ((g1037) & (g1038) & (g1039) & (g1040) & (g1041) & (!g1042)) + ((g1037) & (g1038) & (g1039) & (g1040) & (g1041) & (g1042)));
	assign g1045 = (((!g1043) & (sk[38]) & (g1044)) + ((g1043) & (!sk[38]) & (!g1044)) + ((g1043) & (!sk[38]) & (g1044)) + ((g1043) & (sk[38]) & (!g1044)));
	assign g1046 = (((!g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1035)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1035)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1035)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (g1035)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1035)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1035)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (g1035)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1035)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1035)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1035)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (g1041) & (g1035)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1035)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (g1035)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1035)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1035)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1035)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (g1035)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1035)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1035)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1035)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1035)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (!g1035)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1035)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (g1034) & (g1041) & (!g1035)));
	assign g1047 = (((!g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1035)) + ((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1035)) + ((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (g1035)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1035)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1035)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1035)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1035)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (!g1035)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1035)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1035)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1035)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1035)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1035)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1035)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1035)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1035)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1035)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1035)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1035)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (g1035)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (g1035)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (!g1035)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1035)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1035)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (!g1035)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1035)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (g1034) & (g1041) & (!g1035)));
	assign g1048 = (((!g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1035)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1035)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1035)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1035)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1035)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1035)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1035)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1035)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1035)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1035)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1035)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1035)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1035)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (g1041) & (!g1035)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (g1035)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1035)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1035)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1035)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (g1035)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1035)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (g1035)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1035)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (g1035)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1035)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (!g1035)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1035)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (g1034) & (g1041) & (!g1035)) + ((g1031) & (g1032) & (g1033) & (g1034) & (g1041) & (g1035)));
	assign g1049 = (((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1035)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1035)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1035)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (g1035)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1035)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1035)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1035)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (g1035)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1035)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1035)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1035)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (g1041) & (!g1035)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (g1041) & (g1035)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1035)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1035)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1035)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1035)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1035)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (g1035)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1035)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1035)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1035)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1035)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1035)) + ((g1031) & (g1032) & (g1033) & (g1034) & (g1041) & (g1035)));
	assign g1050 = (((!g1046) & (!g1047) & (!g1048) & (!g1049) & (!g1036) & (!g1042)) + ((!g1046) & (!g1047) & (!g1048) & (!g1049) & (g1036) & (!g1042)) + ((!g1046) & (!g1047) & (!g1048) & (g1049) & (!g1036) & (!g1042)) + ((!g1046) & (!g1047) & (!g1048) & (g1049) & (g1036) & (!g1042)) + ((!g1046) & (!g1047) & (!g1048) & (g1049) & (g1036) & (g1042)) + ((!g1046) & (!g1047) & (g1048) & (!g1049) & (!g1036) & (!g1042)) + ((!g1046) & (!g1047) & (g1048) & (!g1049) & (!g1036) & (g1042)) + ((!g1046) & (!g1047) & (g1048) & (!g1049) & (g1036) & (!g1042)) + ((!g1046) & (!g1047) & (g1048) & (g1049) & (!g1036) & (!g1042)) + ((!g1046) & (!g1047) & (g1048) & (g1049) & (!g1036) & (g1042)) + ((!g1046) & (!g1047) & (g1048) & (g1049) & (g1036) & (!g1042)) + ((!g1046) & (!g1047) & (g1048) & (g1049) & (g1036) & (g1042)) + ((!g1046) & (g1047) & (!g1048) & (!g1049) & (!g1036) & (!g1042)) + ((!g1046) & (g1047) & (!g1048) & (g1049) & (!g1036) & (!g1042)) + ((!g1046) & (g1047) & (!g1048) & (g1049) & (g1036) & (g1042)) + ((!g1046) & (g1047) & (g1048) & (!g1049) & (!g1036) & (!g1042)) + ((!g1046) & (g1047) & (g1048) & (!g1049) & (!g1036) & (g1042)) + ((!g1046) & (g1047) & (g1048) & (g1049) & (!g1036) & (!g1042)) + ((!g1046) & (g1047) & (g1048) & (g1049) & (!g1036) & (g1042)) + ((!g1046) & (g1047) & (g1048) & (g1049) & (g1036) & (g1042)) + ((g1046) & (!g1047) & (!g1048) & (!g1049) & (g1036) & (!g1042)) + ((g1046) & (!g1047) & (!g1048) & (g1049) & (g1036) & (!g1042)) + ((g1046) & (!g1047) & (!g1048) & (g1049) & (g1036) & (g1042)) + ((g1046) & (!g1047) & (g1048) & (!g1049) & (!g1036) & (g1042)) + ((g1046) & (!g1047) & (g1048) & (!g1049) & (g1036) & (!g1042)) + ((g1046) & (!g1047) & (g1048) & (g1049) & (!g1036) & (g1042)) + ((g1046) & (!g1047) & (g1048) & (g1049) & (g1036) & (!g1042)) + ((g1046) & (!g1047) & (g1048) & (g1049) & (g1036) & (g1042)) + ((g1046) & (g1047) & (!g1048) & (g1049) & (g1036) & (g1042)) + ((g1046) & (g1047) & (g1048) & (!g1049) & (!g1036) & (g1042)) + ((g1046) & (g1047) & (g1048) & (g1049) & (!g1036) & (g1042)) + ((g1046) & (g1047) & (g1048) & (g1049) & (g1036) & (g1042)));
	assign g1052 = (((!g1050) & (sk[44]) & (g1051)) + ((g1050) & (!sk[44]) & (!g1051)) + ((g1050) & (!sk[44]) & (g1051)) + ((g1050) & (sk[44]) & (!g1051)));
	assign g1053 = (((!g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1036)));
	assign g1054 = (((!g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((g1035) & (!g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((g1035) & (g1032) & (g1033) & (g1034) & (g1041) & (g1036)));
	assign g1055 = (((!g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1035) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1035) & (!g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1036)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((g1035) & (g1032) & (g1033) & (g1034) & (g1041) & (g1036)));
	assign g1056 = (((!g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1036)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (g1041) & (g1036)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1035) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)));
	assign g1057 = (((!g1053) & (!g1054) & (!g1055) & (!g1056) & (!g1031) & (g1042)) + ((!g1053) & (!g1054) & (!g1055) & (!g1056) & (g1031) & (!g1042)) + ((!g1053) & (!g1054) & (!g1055) & (!g1056) & (g1031) & (g1042)) + ((!g1053) & (!g1054) & (!g1055) & (g1056) & (!g1031) & (g1042)) + ((!g1053) & (!g1054) & (!g1055) & (g1056) & (g1031) & (!g1042)) + ((!g1053) & (!g1054) & (g1055) & (!g1056) & (g1031) & (!g1042)) + ((!g1053) & (!g1054) & (g1055) & (!g1056) & (g1031) & (g1042)) + ((!g1053) & (!g1054) & (g1055) & (g1056) & (g1031) & (!g1042)) + ((!g1053) & (g1054) & (!g1055) & (!g1056) & (!g1031) & (g1042)) + ((!g1053) & (g1054) & (!g1055) & (!g1056) & (g1031) & (g1042)) + ((!g1053) & (g1054) & (!g1055) & (g1056) & (!g1031) & (g1042)) + ((!g1053) & (g1054) & (g1055) & (!g1056) & (g1031) & (g1042)) + ((g1053) & (!g1054) & (!g1055) & (!g1056) & (!g1031) & (!g1042)) + ((g1053) & (!g1054) & (!g1055) & (!g1056) & (!g1031) & (g1042)) + ((g1053) & (!g1054) & (!g1055) & (!g1056) & (g1031) & (!g1042)) + ((g1053) & (!g1054) & (!g1055) & (!g1056) & (g1031) & (g1042)) + ((g1053) & (!g1054) & (!g1055) & (g1056) & (!g1031) & (!g1042)) + ((g1053) & (!g1054) & (!g1055) & (g1056) & (!g1031) & (g1042)) + ((g1053) & (!g1054) & (!g1055) & (g1056) & (g1031) & (!g1042)) + ((g1053) & (!g1054) & (g1055) & (!g1056) & (!g1031) & (!g1042)) + ((g1053) & (!g1054) & (g1055) & (!g1056) & (g1031) & (!g1042)) + ((g1053) & (!g1054) & (g1055) & (!g1056) & (g1031) & (g1042)) + ((g1053) & (!g1054) & (g1055) & (g1056) & (!g1031) & (!g1042)) + ((g1053) & (!g1054) & (g1055) & (g1056) & (g1031) & (!g1042)) + ((g1053) & (g1054) & (!g1055) & (!g1056) & (!g1031) & (!g1042)) + ((g1053) & (g1054) & (!g1055) & (!g1056) & (!g1031) & (g1042)) + ((g1053) & (g1054) & (!g1055) & (!g1056) & (g1031) & (g1042)) + ((g1053) & (g1054) & (!g1055) & (g1056) & (!g1031) & (!g1042)) + ((g1053) & (g1054) & (!g1055) & (g1056) & (!g1031) & (g1042)) + ((g1053) & (g1054) & (g1055) & (!g1056) & (!g1031) & (!g1042)) + ((g1053) & (g1054) & (g1055) & (!g1056) & (g1031) & (g1042)) + ((g1053) & (g1054) & (g1055) & (g1056) & (!g1031) & (!g1042)));
	assign g1059 = (((!g1057) & (sk[50]) & (g1058)) + ((g1057) & (!sk[50]) & (!g1058)) + ((g1057) & (!sk[50]) & (g1058)) + ((g1057) & (sk[50]) & (!g1058)));
	assign g1060 = (((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1036)));
	assign g1061 = (((!g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)));
	assign g1062 = (((!g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (g1041) & (g1036)));
	assign g1063 = (((!g1031) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (g1033) & (g1034) & (g1041) & (g1036)));
	assign g1064 = (((!g1060) & (!g1061) & (!g1062) & (!g1063) & (!g1042) & (g1035)) + ((!g1060) & (!g1061) & (!g1062) & (!g1063) & (g1042) & (!g1035)) + ((!g1060) & (!g1061) & (!g1062) & (!g1063) & (g1042) & (g1035)) + ((!g1060) & (!g1061) & (!g1062) & (g1063) & (!g1042) & (g1035)) + ((!g1060) & (!g1061) & (!g1062) & (g1063) & (g1042) & (!g1035)) + ((!g1060) & (!g1061) & (g1062) & (!g1063) & (g1042) & (!g1035)) + ((!g1060) & (!g1061) & (g1062) & (!g1063) & (g1042) & (g1035)) + ((!g1060) & (!g1061) & (g1062) & (g1063) & (g1042) & (!g1035)) + ((!g1060) & (g1061) & (!g1062) & (!g1063) & (!g1042) & (g1035)) + ((!g1060) & (g1061) & (!g1062) & (!g1063) & (g1042) & (g1035)) + ((!g1060) & (g1061) & (!g1062) & (g1063) & (!g1042) & (g1035)) + ((!g1060) & (g1061) & (g1062) & (!g1063) & (g1042) & (g1035)) + ((g1060) & (!g1061) & (!g1062) & (!g1063) & (!g1042) & (!g1035)) + ((g1060) & (!g1061) & (!g1062) & (!g1063) & (!g1042) & (g1035)) + ((g1060) & (!g1061) & (!g1062) & (!g1063) & (g1042) & (!g1035)) + ((g1060) & (!g1061) & (!g1062) & (!g1063) & (g1042) & (g1035)) + ((g1060) & (!g1061) & (!g1062) & (g1063) & (!g1042) & (!g1035)) + ((g1060) & (!g1061) & (!g1062) & (g1063) & (!g1042) & (g1035)) + ((g1060) & (!g1061) & (!g1062) & (g1063) & (g1042) & (!g1035)) + ((g1060) & (!g1061) & (g1062) & (!g1063) & (!g1042) & (!g1035)) + ((g1060) & (!g1061) & (g1062) & (!g1063) & (g1042) & (!g1035)) + ((g1060) & (!g1061) & (g1062) & (!g1063) & (g1042) & (g1035)) + ((g1060) & (!g1061) & (g1062) & (g1063) & (!g1042) & (!g1035)) + ((g1060) & (!g1061) & (g1062) & (g1063) & (g1042) & (!g1035)) + ((g1060) & (g1061) & (!g1062) & (!g1063) & (!g1042) & (!g1035)) + ((g1060) & (g1061) & (!g1062) & (!g1063) & (!g1042) & (g1035)) + ((g1060) & (g1061) & (!g1062) & (!g1063) & (g1042) & (g1035)) + ((g1060) & (g1061) & (!g1062) & (g1063) & (!g1042) & (!g1035)) + ((g1060) & (g1061) & (!g1062) & (g1063) & (!g1042) & (g1035)) + ((g1060) & (g1061) & (g1062) & (!g1063) & (!g1042) & (!g1035)) + ((g1060) & (g1061) & (g1062) & (!g1063) & (g1042) & (g1035)) + ((g1060) & (g1061) & (g1062) & (g1063) & (!g1042) & (!g1035)));
	assign g1066 = (((!g1064) & (sk[56]) & (g1065)) + ((g1064) & (!sk[56]) & (!g1065)) + ((g1064) & (!sk[56]) & (g1065)) + ((g1064) & (sk[56]) & (!g1065)));
	assign g1067 = (((!g1031) & (!g1032) & (!g1035) & (!g1042) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1042) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1042) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1042) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1042) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1042) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1035) & (!g1042) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1035) & (!g1042) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1042) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1042) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1042) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (g1042) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (g1042) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1042) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1042) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1042) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1042) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1035) & (g1042) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1035) & (g1042) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (g1042) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1042) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1042) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (g1042) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (!g1042) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (!g1042) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (g1035) & (g1042) & (!g1041) & (g1036)));
	assign g1068 = (((!g1031) & (!g1032) & (!g1035) & (!g1042) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1035) & (!g1042) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (!g1035) & (!g1042) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1035) & (!g1042) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (!g1035) & (g1042) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1042) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1042) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1042) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1042) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (!g1042) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1042) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1042) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1042) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1042) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1042) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (g1042) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (g1042) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1042) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1042) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1042) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1042) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1042) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1042) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1042) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (g1042) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1042) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1042) & (g1041) & (g1036)) + ((g1031) & (g1032) & (!g1035) & (g1042) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (g1042) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (g1035) & (!g1042) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (!g1042) & (g1041) & (g1036)) + ((g1031) & (g1032) & (g1035) & (g1042) & (!g1041) & (g1036)));
	assign g1069 = (((!g1031) & (!g1032) & (!g1035) & (!g1042) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1035) & (!g1042) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1042) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1042) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1042) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1042) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1042) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1042) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1042) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1042) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1042) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (g1042) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (g1042) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1042) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1042) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1042) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1042) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1042) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1042) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1042) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (g1042) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1035) & (g1042) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (g1042) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1035) & (g1042) & (g1041) & (g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1042) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (!g1035) & (g1042) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (g1042) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (!g1042) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (!g1042) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (g1035) & (!g1042) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (g1042) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (g1042) & (g1041) & (!g1036)));
	assign g1070 = (((!g1031) & (!g1032) & (!g1035) & (!g1042) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (!g1035) & (g1042) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1035) & (g1042) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1042) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1042) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1042) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1042) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1042) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1035) & (!g1042) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1042) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1042) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1042) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1042) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (g1042) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (g1042) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1042) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1042) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1042) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1042) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1035) & (g1042) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1042) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (g1042) & (g1041) & (g1036)) + ((g1031) & (g1032) & (g1035) & (!g1042) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (!g1042) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (g1035) & (!g1042) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (g1042) & (!g1041) & (!g1036)));
	assign g1071 = (((!g1067) & (!g1068) & (!g1069) & (!g1070) & (g1033) & (g1034)) + ((!g1067) & (!g1068) & (g1069) & (!g1070) & (!g1033) & (g1034)) + ((!g1067) & (!g1068) & (g1069) & (!g1070) & (g1033) & (g1034)) + ((!g1067) & (!g1068) & (g1069) & (g1070) & (!g1033) & (g1034)) + ((!g1067) & (g1068) & (!g1069) & (!g1070) & (g1033) & (!g1034)) + ((!g1067) & (g1068) & (!g1069) & (!g1070) & (g1033) & (g1034)) + ((!g1067) & (g1068) & (!g1069) & (g1070) & (g1033) & (!g1034)) + ((!g1067) & (g1068) & (g1069) & (!g1070) & (!g1033) & (g1034)) + ((!g1067) & (g1068) & (g1069) & (!g1070) & (g1033) & (!g1034)) + ((!g1067) & (g1068) & (g1069) & (!g1070) & (g1033) & (g1034)) + ((!g1067) & (g1068) & (g1069) & (g1070) & (!g1033) & (g1034)) + ((!g1067) & (g1068) & (g1069) & (g1070) & (g1033) & (!g1034)) + ((g1067) & (!g1068) & (!g1069) & (!g1070) & (!g1033) & (!g1034)) + ((g1067) & (!g1068) & (!g1069) & (!g1070) & (g1033) & (g1034)) + ((g1067) & (!g1068) & (!g1069) & (g1070) & (!g1033) & (!g1034)) + ((g1067) & (!g1068) & (g1069) & (!g1070) & (!g1033) & (!g1034)) + ((g1067) & (!g1068) & (g1069) & (!g1070) & (!g1033) & (g1034)) + ((g1067) & (!g1068) & (g1069) & (!g1070) & (g1033) & (g1034)) + ((g1067) & (!g1068) & (g1069) & (g1070) & (!g1033) & (!g1034)) + ((g1067) & (!g1068) & (g1069) & (g1070) & (!g1033) & (g1034)) + ((g1067) & (g1068) & (!g1069) & (!g1070) & (!g1033) & (!g1034)) + ((g1067) & (g1068) & (!g1069) & (!g1070) & (g1033) & (!g1034)) + ((g1067) & (g1068) & (!g1069) & (!g1070) & (g1033) & (g1034)) + ((g1067) & (g1068) & (!g1069) & (g1070) & (!g1033) & (!g1034)) + ((g1067) & (g1068) & (!g1069) & (g1070) & (g1033) & (!g1034)) + ((g1067) & (g1068) & (g1069) & (!g1070) & (!g1033) & (!g1034)) + ((g1067) & (g1068) & (g1069) & (!g1070) & (!g1033) & (g1034)) + ((g1067) & (g1068) & (g1069) & (!g1070) & (g1033) & (!g1034)) + ((g1067) & (g1068) & (g1069) & (!g1070) & (g1033) & (g1034)) + ((g1067) & (g1068) & (g1069) & (g1070) & (!g1033) & (!g1034)) + ((g1067) & (g1068) & (g1069) & (g1070) & (!g1033) & (g1034)) + ((g1067) & (g1068) & (g1069) & (g1070) & (g1033) & (!g1034)));
	assign g1073 = (((!g1071) & (sk[62]) & (g1072)) + ((g1071) & (!sk[62]) & (!g1072)) + ((g1071) & (!sk[62]) & (g1072)) + ((g1071) & (sk[62]) & (!g1072)));
	assign g1074 = (((!g1031) & (!g1032) & (!g1035) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1035) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (!g1035) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1035) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (g1032) & (g1035) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (!g1034) & (g1041) & (g1036)));
	assign g1075 = (((!g1031) & (!g1032) & (!g1035) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1035) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1035) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (!g1035) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1035) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1035) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (g1034) & (g1041) & (g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (g1035) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (g1032) & (g1035) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (g1034) & (g1041) & (g1036)));
	assign g1076 = (((!g1031) & (!g1032) & (!g1035) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (!g1035) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (!g1035) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (g1032) & (!g1035) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (!g1035) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (g1035) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (g1032) & (g1035) & (g1034) & (g1041) & (g1036)));
	assign g1077 = (((!g1031) & (!g1032) & (!g1035) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1035) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1032) & (!g1035) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1032) & (g1035) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (!g1035) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1032) & (g1035) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1032) & (g1035) & (g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (!g1035) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1032) & (!g1035) & (g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1032) & (g1035) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1032) & (g1035) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (g1032) & (!g1035) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1032) & (!g1035) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (g1032) & (g1035) & (!g1034) & (g1041) & (g1036)));
	assign g1078 = (((!g1074) & (!g1075) & (!g1076) & (!g1077) & (!g1042) & (!g1033)) + ((!g1074) & (!g1075) & (!g1076) & (!g1077) & (!g1042) & (g1033)) + ((!g1074) & (!g1075) & (!g1076) & (!g1077) & (g1042) & (!g1033)) + ((!g1074) & (!g1075) & (!g1076) & (g1077) & (!g1042) & (!g1033)) + ((!g1074) & (!g1075) & (!g1076) & (g1077) & (!g1042) & (g1033)) + ((!g1074) & (!g1075) & (!g1076) & (g1077) & (g1042) & (!g1033)) + ((!g1074) & (!g1075) & (!g1076) & (g1077) & (g1042) & (g1033)) + ((!g1074) & (!g1075) & (g1076) & (!g1077) & (!g1042) & (!g1033)) + ((!g1074) & (!g1075) & (g1076) & (!g1077) & (g1042) & (!g1033)) + ((!g1074) & (!g1075) & (g1076) & (g1077) & (!g1042) & (!g1033)) + ((!g1074) & (!g1075) & (g1076) & (g1077) & (g1042) & (!g1033)) + ((!g1074) & (!g1075) & (g1076) & (g1077) & (g1042) & (g1033)) + ((!g1074) & (g1075) & (!g1076) & (!g1077) & (!g1042) & (!g1033)) + ((!g1074) & (g1075) & (!g1076) & (!g1077) & (!g1042) & (g1033)) + ((!g1074) & (g1075) & (!g1076) & (g1077) & (!g1042) & (!g1033)) + ((!g1074) & (g1075) & (!g1076) & (g1077) & (!g1042) & (g1033)) + ((!g1074) & (g1075) & (!g1076) & (g1077) & (g1042) & (g1033)) + ((!g1074) & (g1075) & (g1076) & (!g1077) & (!g1042) & (!g1033)) + ((!g1074) & (g1075) & (g1076) & (g1077) & (!g1042) & (!g1033)) + ((!g1074) & (g1075) & (g1076) & (g1077) & (g1042) & (g1033)) + ((g1074) & (!g1075) & (!g1076) & (!g1077) & (!g1042) & (g1033)) + ((g1074) & (!g1075) & (!g1076) & (!g1077) & (g1042) & (!g1033)) + ((g1074) & (!g1075) & (!g1076) & (g1077) & (!g1042) & (g1033)) + ((g1074) & (!g1075) & (!g1076) & (g1077) & (g1042) & (!g1033)) + ((g1074) & (!g1075) & (!g1076) & (g1077) & (g1042) & (g1033)) + ((g1074) & (!g1075) & (g1076) & (!g1077) & (g1042) & (!g1033)) + ((g1074) & (!g1075) & (g1076) & (g1077) & (g1042) & (!g1033)) + ((g1074) & (!g1075) & (g1076) & (g1077) & (g1042) & (g1033)) + ((g1074) & (g1075) & (!g1076) & (!g1077) & (!g1042) & (g1033)) + ((g1074) & (g1075) & (!g1076) & (g1077) & (!g1042) & (g1033)) + ((g1074) & (g1075) & (!g1076) & (g1077) & (g1042) & (g1033)) + ((g1074) & (g1075) & (g1076) & (g1077) & (g1042) & (g1033)));
	assign g1080 = (((!g1078) & (sk[68]) & (g1079)) + ((g1078) & (!sk[68]) & (!g1079)) + ((g1078) & (!sk[68]) & (g1079)) + ((g1078) & (sk[68]) & (!g1079)));
	assign g1081 = (((!g1031) & (!g1042) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1042) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1042) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1042) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1042) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1042) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1042) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1042) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1042) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1042) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1042) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (g1042) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1042) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1042) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1042) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1042) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((g1031) & (!g1042) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1042) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1042) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1042) & (g1033) & (g1034) & (g1041) & (g1036)) + ((g1031) & (g1042) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1042) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (g1042) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (g1042) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1042) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1042) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (g1042) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (g1042) & (g1033) & (g1034) & (!g1041) & (g1036)));
	assign g1082 = (((!g1031) & (!g1042) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1042) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1042) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1042) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1042) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1042) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1042) & (g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1042) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1042) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (g1042) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1042) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1042) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (g1042) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1042) & (g1033) & (g1034) & (g1041) & (g1036)) + ((g1031) & (!g1042) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1042) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1042) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1042) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((g1031) & (!g1042) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1042) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (g1042) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (g1042) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (g1042) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (g1042) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (g1042) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((g1031) & (g1042) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1042) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (g1042) & (g1033) & (g1034) & (!g1041) & (!g1036)));
	assign g1083 = (((!g1031) & (!g1042) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1042) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1042) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1042) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1042) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1042) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1042) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (!g1042) & (g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1042) & (!g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1042) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1042) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (g1042) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1042) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1042) & (g1033) & (!g1034) & (!g1041) & (g1036)) + ((!g1031) & (g1042) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1042) & (g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1042) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1042) & (g1033) & (g1034) & (g1041) & (g1036)) + ((g1031) & (!g1042) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1042) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (!g1042) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1042) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1042) & (g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (g1042) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (g1042) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1042) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (g1042) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1042) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (g1042) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (g1042) & (g1033) & (g1034) & (g1041) & (g1036)));
	assign g1084 = (((!g1031) & (!g1042) & (!g1033) & (!g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1042) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1042) & (!g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (!g1042) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((!g1031) & (!g1042) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (!g1042) & (g1033) & (g1034) & (g1041) & (g1036)) + ((!g1031) & (g1042) & (!g1033) & (g1034) & (!g1041) & (!g1036)) + ((!g1031) & (g1042) & (!g1033) & (g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1042) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((!g1031) & (g1042) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1042) & (!g1033) & (!g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1042) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1042) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (!g1042) & (g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1042) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (!g1042) & (g1033) & (g1034) & (g1041) & (!g1036)) + ((g1031) & (!g1042) & (g1033) & (g1034) & (g1041) & (g1036)) + ((g1031) & (g1042) & (!g1033) & (!g1034) & (g1041) & (!g1036)) + ((g1031) & (g1042) & (!g1033) & (g1034) & (!g1041) & (g1036)) + ((g1031) & (g1042) & (g1033) & (!g1034) & (!g1041) & (!g1036)) + ((g1031) & (g1042) & (g1033) & (!g1034) & (g1041) & (g1036)) + ((g1031) & (g1042) & (g1033) & (g1034) & (!g1041) & (g1036)));
	assign g1085 = (((!g1081) & (!g1082) & (!g1083) & (!g1084) & (!g1035) & (!g1032)) + ((!g1081) & (!g1082) & (!g1083) & (!g1084) & (!g1035) & (g1032)) + ((!g1081) & (!g1082) & (!g1083) & (!g1084) & (g1035) & (!g1032)) + ((!g1081) & (!g1082) & (!g1083) & (g1084) & (!g1035) & (!g1032)) + ((!g1081) & (!g1082) & (!g1083) & (g1084) & (!g1035) & (g1032)) + ((!g1081) & (!g1082) & (!g1083) & (g1084) & (g1035) & (!g1032)) + ((!g1081) & (!g1082) & (!g1083) & (g1084) & (g1035) & (g1032)) + ((!g1081) & (!g1082) & (g1083) & (!g1084) & (!g1035) & (!g1032)) + ((!g1081) & (!g1082) & (g1083) & (!g1084) & (g1035) & (!g1032)) + ((!g1081) & (!g1082) & (g1083) & (g1084) & (!g1035) & (!g1032)) + ((!g1081) & (!g1082) & (g1083) & (g1084) & (g1035) & (!g1032)) + ((!g1081) & (!g1082) & (g1083) & (g1084) & (g1035) & (g1032)) + ((!g1081) & (g1082) & (!g1083) & (!g1084) & (!g1035) & (!g1032)) + ((!g1081) & (g1082) & (!g1083) & (!g1084) & (!g1035) & (g1032)) + ((!g1081) & (g1082) & (!g1083) & (g1084) & (!g1035) & (!g1032)) + ((!g1081) & (g1082) & (!g1083) & (g1084) & (!g1035) & (g1032)) + ((!g1081) & (g1082) & (!g1083) & (g1084) & (g1035) & (g1032)) + ((!g1081) & (g1082) & (g1083) & (!g1084) & (!g1035) & (!g1032)) + ((!g1081) & (g1082) & (g1083) & (g1084) & (!g1035) & (!g1032)) + ((!g1081) & (g1082) & (g1083) & (g1084) & (g1035) & (g1032)) + ((g1081) & (!g1082) & (!g1083) & (!g1084) & (!g1035) & (g1032)) + ((g1081) & (!g1082) & (!g1083) & (!g1084) & (g1035) & (!g1032)) + ((g1081) & (!g1082) & (!g1083) & (g1084) & (!g1035) & (g1032)) + ((g1081) & (!g1082) & (!g1083) & (g1084) & (g1035) & (!g1032)) + ((g1081) & (!g1082) & (!g1083) & (g1084) & (g1035) & (g1032)) + ((g1081) & (!g1082) & (g1083) & (!g1084) & (g1035) & (!g1032)) + ((g1081) & (!g1082) & (g1083) & (g1084) & (g1035) & (!g1032)) + ((g1081) & (!g1082) & (g1083) & (g1084) & (g1035) & (g1032)) + ((g1081) & (g1082) & (!g1083) & (!g1084) & (!g1035) & (g1032)) + ((g1081) & (g1082) & (!g1083) & (g1084) & (!g1035) & (g1032)) + ((g1081) & (g1082) & (!g1083) & (g1084) & (g1035) & (g1032)) + ((g1081) & (g1082) & (g1083) & (g1084) & (g1035) & (g1032)));
	assign g1087 = (((!g1085) & (sk[74]) & (g1086)) + ((g1085) & (!sk[74]) & (!g1086)) + ((g1085) & (!sk[74]) & (g1086)) + ((g1085) & (sk[74]) & (!g1086)));
	assign g1088 = (((!g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1042)) + ((!g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1042)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1042)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (!g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1042)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1042)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1042)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1042)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1042)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1042)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1042)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1042)) + ((g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1042)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1042)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1042)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1042)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1042)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1042)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1042)) + ((g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1042)));
	assign g1089 = (((!g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1042)) + ((!g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1042)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (g1041) & (g1042)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1042)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1042)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1042)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1042)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1042)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (g1042)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1042)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1042)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1042)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1042)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1042)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (g1042)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1042)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1042)) + ((g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1042)) + ((g1035) & (!g1032) & (g1033) & (!g1034) & (g1041) & (g1042)) + ((g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1042)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1042)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (g1042)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1042)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (g1042)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1042)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1042)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1042)));
	assign g1090 = (((!g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1042)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1042)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1042)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1042)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (g1042)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (!g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1042)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (g1042)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1042)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1042)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1042)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1042)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1042)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1042)) + ((g1035) & (!g1032) & (!g1033) & (!g1034) & (g1041) & (!g1042)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (!g1042)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1042)) + ((g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1042)) + ((g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (g1042)) + ((g1035) & (!g1032) & (g1033) & (g1034) & (!g1041) & (!g1042)) + ((g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1042)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (g1041) & (!g1042)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1042)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1042)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (!g1041) & (!g1042)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (!g1042)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1042)) + ((g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1042)));
	assign g1091 = (((!g1035) & (!g1032) & (!g1033) & (!g1034) & (!g1041) & (g1042)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (!g1042)) + ((!g1035) & (!g1032) & (!g1033) & (g1034) & (g1041) & (g1042)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (g1042)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (!g1042)) + ((!g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1042)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (!g1042)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (g1042)) + ((!g1035) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1042)) + ((!g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (g1042)) + ((!g1035) & (g1032) & (g1033) & (!g1034) & (!g1041) & (g1042)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (!g1042)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (!g1041) & (g1042)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (g1041) & (!g1042)) + ((!g1035) & (g1032) & (g1033) & (g1034) & (g1041) & (g1042)) + ((g1035) & (!g1032) & (!g1033) & (g1034) & (!g1041) & (g1042)) + ((g1035) & (!g1032) & (g1033) & (!g1034) & (!g1041) & (!g1042)) + ((g1035) & (!g1032) & (g1033) & (g1034) & (!g1041) & (!g1042)) + ((g1035) & (!g1032) & (g1033) & (g1034) & (!g1041) & (g1042)) + ((g1035) & (!g1032) & (g1033) & (g1034) & (g1041) & (g1042)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (!g1041) & (g1042)) + ((g1035) & (g1032) & (!g1033) & (!g1034) & (g1041) & (g1042)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (!g1041) & (!g1042)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (!g1042)) + ((g1035) & (g1032) & (!g1033) & (g1034) & (g1041) & (g1042)) + ((g1035) & (g1032) & (g1033) & (!g1034) & (g1041) & (g1042)) + ((g1035) & (g1032) & (g1033) & (g1034) & (g1041) & (g1042)));
	assign g1092 = (((!g1088) & (!g1089) & (!g1090) & (!g1091) & (!g1031) & (g1036)) + ((!g1088) & (!g1089) & (!g1090) & (!g1091) & (g1031) & (!g1036)) + ((!g1088) & (!g1089) & (!g1090) & (!g1091) & (g1031) & (g1036)) + ((!g1088) & (!g1089) & (!g1090) & (g1091) & (!g1031) & (g1036)) + ((!g1088) & (!g1089) & (!g1090) & (g1091) & (g1031) & (!g1036)) + ((!g1088) & (!g1089) & (g1090) & (!g1091) & (g1031) & (!g1036)) + ((!g1088) & (!g1089) & (g1090) & (!g1091) & (g1031) & (g1036)) + ((!g1088) & (!g1089) & (g1090) & (g1091) & (g1031) & (!g1036)) + ((!g1088) & (g1089) & (!g1090) & (!g1091) & (!g1031) & (g1036)) + ((!g1088) & (g1089) & (!g1090) & (!g1091) & (g1031) & (g1036)) + ((!g1088) & (g1089) & (!g1090) & (g1091) & (!g1031) & (g1036)) + ((!g1088) & (g1089) & (g1090) & (!g1091) & (g1031) & (g1036)) + ((g1088) & (!g1089) & (!g1090) & (!g1091) & (!g1031) & (!g1036)) + ((g1088) & (!g1089) & (!g1090) & (!g1091) & (!g1031) & (g1036)) + ((g1088) & (!g1089) & (!g1090) & (!g1091) & (g1031) & (!g1036)) + ((g1088) & (!g1089) & (!g1090) & (!g1091) & (g1031) & (g1036)) + ((g1088) & (!g1089) & (!g1090) & (g1091) & (!g1031) & (!g1036)) + ((g1088) & (!g1089) & (!g1090) & (g1091) & (!g1031) & (g1036)) + ((g1088) & (!g1089) & (!g1090) & (g1091) & (g1031) & (!g1036)) + ((g1088) & (!g1089) & (g1090) & (!g1091) & (!g1031) & (!g1036)) + ((g1088) & (!g1089) & (g1090) & (!g1091) & (g1031) & (!g1036)) + ((g1088) & (!g1089) & (g1090) & (!g1091) & (g1031) & (g1036)) + ((g1088) & (!g1089) & (g1090) & (g1091) & (!g1031) & (!g1036)) + ((g1088) & (!g1089) & (g1090) & (g1091) & (g1031) & (!g1036)) + ((g1088) & (g1089) & (!g1090) & (!g1091) & (!g1031) & (!g1036)) + ((g1088) & (g1089) & (!g1090) & (!g1091) & (!g1031) & (g1036)) + ((g1088) & (g1089) & (!g1090) & (!g1091) & (g1031) & (g1036)) + ((g1088) & (g1089) & (!g1090) & (g1091) & (!g1031) & (!g1036)) + ((g1088) & (g1089) & (!g1090) & (g1091) & (!g1031) & (g1036)) + ((g1088) & (g1089) & (g1090) & (!g1091) & (!g1031) & (!g1036)) + ((g1088) & (g1089) & (g1090) & (!g1091) & (g1031) & (g1036)) + ((g1088) & (g1089) & (g1090) & (g1091) & (!g1031) & (!g1036)));
	assign g1094 = (((!g1092) & (sk[80]) & (g1093)) + ((g1092) & (!sk[80]) & (!g1093)) + ((g1092) & (!sk[80]) & (g1093)) + ((g1092) & (sk[80]) & (!g1093)));
	assign g1101 = (((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1099) & (g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1099) & (!g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1099) & (g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (g1099) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (!g1099) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (!g1099) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1099) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (g1099) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1099) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1099) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (g1099) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (g1099) & (g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (g1099) & (!g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1099) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1099) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (!g1099) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (g1099) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (!g1099) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (g1099) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1099) & (g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (g1099) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1099) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (g1099) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (g1099) & (g1100)));
	assign g1102 = (((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1099) & (!g1100)) + ((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1099) & (g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1099) & (!g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1099) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1099) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (!g1099) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (!g1099) & (g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (!g1099) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (!g1099) & (g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (g1099) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (g1099) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1099) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (g1099) & (!g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (g1099) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (g1099) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (!g1099) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1099) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (!g1099) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (g1099) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (!g1099) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (!g1099) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (g1099) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (g1099) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (!g1099) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1099) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1099) & (g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (g1099) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (g1099) & (g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1099) & (g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (g1099) & (!g1100)));
	assign g1103 = (((!g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1099) & (!g1100)) + ((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1099) & (g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (g1099) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (!g1099) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (!g1099) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (g1099) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1099) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (g1099) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (!g1099) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1099) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (g1099) & (g1100)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (!g1099) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (g1099) & (!g1100)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (!g1099) & (!g1100)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (!g1099) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (g1099) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (!g1099) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1099) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (!g1099) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (!g1099) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (g1099) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (g1099) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (g1099) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (!g1099) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1099) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1099) & (g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1099) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1099) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1099) & (g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (g1099) & (g1100)));
	assign g1104 = (((!g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1099) & (g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (g1099) & (!g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (g1099) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (!g1099) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (g1099) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1099) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (!g1099) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (!g1099) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1099) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1099) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (g1099) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (g1099) & (g1100)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (!g1099) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (g1099) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (g1099) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1099) & (!g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (g1099) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (g1099) & (!g1100)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (g1099) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (!g1099) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1099) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (g1099) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (!g1099) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (g1099) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1099) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1099) & (g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1099) & (g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1099) & (!g1100)));
	assign g1107 = (((!g1101) & (!g1102) & (!g1103) & (!g1104) & (!g1105) & (!g1106)) + ((!g1101) & (!g1102) & (!g1103) & (g1104) & (!g1105) & (!g1106)) + ((!g1101) & (!g1102) & (!g1103) & (g1104) & (g1105) & (g1106)) + ((!g1101) & (!g1102) & (g1103) & (!g1104) & (!g1105) & (!g1106)) + ((!g1101) & (!g1102) & (g1103) & (!g1104) & (!g1105) & (g1106)) + ((!g1101) & (!g1102) & (g1103) & (g1104) & (!g1105) & (!g1106)) + ((!g1101) & (!g1102) & (g1103) & (g1104) & (!g1105) & (g1106)) + ((!g1101) & (!g1102) & (g1103) & (g1104) & (g1105) & (g1106)) + ((!g1101) & (g1102) & (!g1103) & (!g1104) & (!g1105) & (!g1106)) + ((!g1101) & (g1102) & (!g1103) & (!g1104) & (g1105) & (!g1106)) + ((!g1101) & (g1102) & (!g1103) & (g1104) & (!g1105) & (!g1106)) + ((!g1101) & (g1102) & (!g1103) & (g1104) & (g1105) & (!g1106)) + ((!g1101) & (g1102) & (!g1103) & (g1104) & (g1105) & (g1106)) + ((!g1101) & (g1102) & (g1103) & (!g1104) & (!g1105) & (!g1106)) + ((!g1101) & (g1102) & (g1103) & (!g1104) & (!g1105) & (g1106)) + ((!g1101) & (g1102) & (g1103) & (!g1104) & (g1105) & (!g1106)) + ((!g1101) & (g1102) & (g1103) & (g1104) & (!g1105) & (!g1106)) + ((!g1101) & (g1102) & (g1103) & (g1104) & (!g1105) & (g1106)) + ((!g1101) & (g1102) & (g1103) & (g1104) & (g1105) & (!g1106)) + ((!g1101) & (g1102) & (g1103) & (g1104) & (g1105) & (g1106)) + ((g1101) & (!g1102) & (!g1103) & (g1104) & (g1105) & (g1106)) + ((g1101) & (!g1102) & (g1103) & (!g1104) & (!g1105) & (g1106)) + ((g1101) & (!g1102) & (g1103) & (g1104) & (!g1105) & (g1106)) + ((g1101) & (!g1102) & (g1103) & (g1104) & (g1105) & (g1106)) + ((g1101) & (g1102) & (!g1103) & (!g1104) & (g1105) & (!g1106)) + ((g1101) & (g1102) & (!g1103) & (g1104) & (g1105) & (!g1106)) + ((g1101) & (g1102) & (!g1103) & (g1104) & (g1105) & (g1106)) + ((g1101) & (g1102) & (g1103) & (!g1104) & (!g1105) & (g1106)) + ((g1101) & (g1102) & (g1103) & (!g1104) & (g1105) & (!g1106)) + ((g1101) & (g1102) & (g1103) & (g1104) & (!g1105) & (g1106)) + ((g1101) & (g1102) & (g1103) & (g1104) & (g1105) & (!g1106)) + ((g1101) & (g1102) & (g1103) & (g1104) & (g1105) & (g1106)));
	assign g1109 = (((!g1107) & (sk[86]) & (g1108)) + ((g1107) & (!sk[86]) & (!g1108)) + ((g1107) & (!sk[86]) & (g1108)) + ((g1107) & (sk[86]) & (!g1108)));
	assign g1110 = (((!g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1099)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1099)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1099)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (g1099)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1099)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1099)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (g1099)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1099)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1099)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1099)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (g1105) & (g1099)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1099)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (g1099)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1099)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1099)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1099)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (g1099)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1099)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1099)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1099)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1099)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (!g1099)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1099)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (g1098) & (g1105) & (!g1099)));
	assign g1111 = (((!g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1099)) + ((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1099)) + ((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (g1099)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1099)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1099)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1099)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1099)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (!g1099)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1099)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1099)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1099)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1099)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1099)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1099)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1099)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1099)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1099)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1099)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1099)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (g1099)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (g1099)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (!g1099)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1099)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1099)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (!g1099)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1099)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (g1098) & (g1105) & (!g1099)));
	assign g1112 = (((!g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1099)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1099)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1099)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1099)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1099)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1099)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1099)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1099)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1099)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1099)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1099)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1099)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1099)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (g1105) & (!g1099)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (g1099)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1099)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1099)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1099)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (g1099)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1099)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (g1099)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1099)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (g1099)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1099)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (!g1099)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1099)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (g1098) & (g1105) & (!g1099)) + ((g1095) & (g1096) & (g1097) & (g1098) & (g1105) & (g1099)));
	assign g1113 = (((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1099)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1099)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1099)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (g1099)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1099)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1099)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1099)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (g1099)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1099)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1099)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1099)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (g1105) & (!g1099)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (g1105) & (g1099)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1099)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1099)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1099)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1099)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1099)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (g1099)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1099)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1099)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1099)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1099)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1099)) + ((g1095) & (g1096) & (g1097) & (g1098) & (g1105) & (g1099)));
	assign g1114 = (((!g1110) & (!g1111) & (!g1112) & (!g1113) & (!g1100) & (!g1106)) + ((!g1110) & (!g1111) & (!g1112) & (!g1113) & (g1100) & (!g1106)) + ((!g1110) & (!g1111) & (!g1112) & (g1113) & (!g1100) & (!g1106)) + ((!g1110) & (!g1111) & (!g1112) & (g1113) & (g1100) & (!g1106)) + ((!g1110) & (!g1111) & (!g1112) & (g1113) & (g1100) & (g1106)) + ((!g1110) & (!g1111) & (g1112) & (!g1113) & (!g1100) & (!g1106)) + ((!g1110) & (!g1111) & (g1112) & (!g1113) & (!g1100) & (g1106)) + ((!g1110) & (!g1111) & (g1112) & (!g1113) & (g1100) & (!g1106)) + ((!g1110) & (!g1111) & (g1112) & (g1113) & (!g1100) & (!g1106)) + ((!g1110) & (!g1111) & (g1112) & (g1113) & (!g1100) & (g1106)) + ((!g1110) & (!g1111) & (g1112) & (g1113) & (g1100) & (!g1106)) + ((!g1110) & (!g1111) & (g1112) & (g1113) & (g1100) & (g1106)) + ((!g1110) & (g1111) & (!g1112) & (!g1113) & (!g1100) & (!g1106)) + ((!g1110) & (g1111) & (!g1112) & (g1113) & (!g1100) & (!g1106)) + ((!g1110) & (g1111) & (!g1112) & (g1113) & (g1100) & (g1106)) + ((!g1110) & (g1111) & (g1112) & (!g1113) & (!g1100) & (!g1106)) + ((!g1110) & (g1111) & (g1112) & (!g1113) & (!g1100) & (g1106)) + ((!g1110) & (g1111) & (g1112) & (g1113) & (!g1100) & (!g1106)) + ((!g1110) & (g1111) & (g1112) & (g1113) & (!g1100) & (g1106)) + ((!g1110) & (g1111) & (g1112) & (g1113) & (g1100) & (g1106)) + ((g1110) & (!g1111) & (!g1112) & (!g1113) & (g1100) & (!g1106)) + ((g1110) & (!g1111) & (!g1112) & (g1113) & (g1100) & (!g1106)) + ((g1110) & (!g1111) & (!g1112) & (g1113) & (g1100) & (g1106)) + ((g1110) & (!g1111) & (g1112) & (!g1113) & (!g1100) & (g1106)) + ((g1110) & (!g1111) & (g1112) & (!g1113) & (g1100) & (!g1106)) + ((g1110) & (!g1111) & (g1112) & (g1113) & (!g1100) & (g1106)) + ((g1110) & (!g1111) & (g1112) & (g1113) & (g1100) & (!g1106)) + ((g1110) & (!g1111) & (g1112) & (g1113) & (g1100) & (g1106)) + ((g1110) & (g1111) & (!g1112) & (g1113) & (g1100) & (g1106)) + ((g1110) & (g1111) & (g1112) & (!g1113) & (!g1100) & (g1106)) + ((g1110) & (g1111) & (g1112) & (g1113) & (!g1100) & (g1106)) + ((g1110) & (g1111) & (g1112) & (g1113) & (g1100) & (g1106)));
	assign g1116 = (((!sk[92]) & (g1114) & (!g1115)) + ((!sk[92]) & (g1114) & (g1115)) + ((sk[92]) & (!g1114) & (g1115)) + ((sk[92]) & (g1114) & (!g1115)));
	assign g1117 = (((!g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1100)));
	assign g1118 = (((!g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((g1099) & (!g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((g1099) & (g1096) & (g1097) & (g1098) & (g1105) & (g1100)));
	assign g1119 = (((!g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1099) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1099) & (!g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1100)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((g1099) & (g1096) & (g1097) & (g1098) & (g1105) & (g1100)));
	assign g1120 = (((!g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1100)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (g1105) & (g1100)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1099) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)));
	assign g1121 = (((!g1117) & (!g1118) & (!g1119) & (!g1120) & (!g1095) & (g1106)) + ((!g1117) & (!g1118) & (!g1119) & (!g1120) & (g1095) & (!g1106)) + ((!g1117) & (!g1118) & (!g1119) & (!g1120) & (g1095) & (g1106)) + ((!g1117) & (!g1118) & (!g1119) & (g1120) & (!g1095) & (g1106)) + ((!g1117) & (!g1118) & (!g1119) & (g1120) & (g1095) & (!g1106)) + ((!g1117) & (!g1118) & (g1119) & (!g1120) & (g1095) & (!g1106)) + ((!g1117) & (!g1118) & (g1119) & (!g1120) & (g1095) & (g1106)) + ((!g1117) & (!g1118) & (g1119) & (g1120) & (g1095) & (!g1106)) + ((!g1117) & (g1118) & (!g1119) & (!g1120) & (!g1095) & (g1106)) + ((!g1117) & (g1118) & (!g1119) & (!g1120) & (g1095) & (g1106)) + ((!g1117) & (g1118) & (!g1119) & (g1120) & (!g1095) & (g1106)) + ((!g1117) & (g1118) & (g1119) & (!g1120) & (g1095) & (g1106)) + ((g1117) & (!g1118) & (!g1119) & (!g1120) & (!g1095) & (!g1106)) + ((g1117) & (!g1118) & (!g1119) & (!g1120) & (!g1095) & (g1106)) + ((g1117) & (!g1118) & (!g1119) & (!g1120) & (g1095) & (!g1106)) + ((g1117) & (!g1118) & (!g1119) & (!g1120) & (g1095) & (g1106)) + ((g1117) & (!g1118) & (!g1119) & (g1120) & (!g1095) & (!g1106)) + ((g1117) & (!g1118) & (!g1119) & (g1120) & (!g1095) & (g1106)) + ((g1117) & (!g1118) & (!g1119) & (g1120) & (g1095) & (!g1106)) + ((g1117) & (!g1118) & (g1119) & (!g1120) & (!g1095) & (!g1106)) + ((g1117) & (!g1118) & (g1119) & (!g1120) & (g1095) & (!g1106)) + ((g1117) & (!g1118) & (g1119) & (!g1120) & (g1095) & (g1106)) + ((g1117) & (!g1118) & (g1119) & (g1120) & (!g1095) & (!g1106)) + ((g1117) & (!g1118) & (g1119) & (g1120) & (g1095) & (!g1106)) + ((g1117) & (g1118) & (!g1119) & (!g1120) & (!g1095) & (!g1106)) + ((g1117) & (g1118) & (!g1119) & (!g1120) & (!g1095) & (g1106)) + ((g1117) & (g1118) & (!g1119) & (!g1120) & (g1095) & (g1106)) + ((g1117) & (g1118) & (!g1119) & (g1120) & (!g1095) & (!g1106)) + ((g1117) & (g1118) & (!g1119) & (g1120) & (!g1095) & (g1106)) + ((g1117) & (g1118) & (g1119) & (!g1120) & (!g1095) & (!g1106)) + ((g1117) & (g1118) & (g1119) & (!g1120) & (g1095) & (g1106)) + ((g1117) & (g1118) & (g1119) & (g1120) & (!g1095) & (!g1106)));
	assign g1123 = (((!g1121) & (sk[98]) & (g1122)) + ((g1121) & (!sk[98]) & (!g1122)) + ((g1121) & (!sk[98]) & (g1122)) + ((g1121) & (sk[98]) & (!g1122)));
	assign g1124 = (((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1100)));
	assign g1125 = (((!g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)));
	assign g1126 = (((!g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (g1105) & (g1100)));
	assign g1127 = (((!g1095) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (g1097) & (g1098) & (g1105) & (g1100)));
	assign g1128 = (((!g1124) & (!g1125) & (!g1126) & (!g1127) & (!g1106) & (g1099)) + ((!g1124) & (!g1125) & (!g1126) & (!g1127) & (g1106) & (!g1099)) + ((!g1124) & (!g1125) & (!g1126) & (!g1127) & (g1106) & (g1099)) + ((!g1124) & (!g1125) & (!g1126) & (g1127) & (!g1106) & (g1099)) + ((!g1124) & (!g1125) & (!g1126) & (g1127) & (g1106) & (!g1099)) + ((!g1124) & (!g1125) & (g1126) & (!g1127) & (g1106) & (!g1099)) + ((!g1124) & (!g1125) & (g1126) & (!g1127) & (g1106) & (g1099)) + ((!g1124) & (!g1125) & (g1126) & (g1127) & (g1106) & (!g1099)) + ((!g1124) & (g1125) & (!g1126) & (!g1127) & (!g1106) & (g1099)) + ((!g1124) & (g1125) & (!g1126) & (!g1127) & (g1106) & (g1099)) + ((!g1124) & (g1125) & (!g1126) & (g1127) & (!g1106) & (g1099)) + ((!g1124) & (g1125) & (g1126) & (!g1127) & (g1106) & (g1099)) + ((g1124) & (!g1125) & (!g1126) & (!g1127) & (!g1106) & (!g1099)) + ((g1124) & (!g1125) & (!g1126) & (!g1127) & (!g1106) & (g1099)) + ((g1124) & (!g1125) & (!g1126) & (!g1127) & (g1106) & (!g1099)) + ((g1124) & (!g1125) & (!g1126) & (!g1127) & (g1106) & (g1099)) + ((g1124) & (!g1125) & (!g1126) & (g1127) & (!g1106) & (!g1099)) + ((g1124) & (!g1125) & (!g1126) & (g1127) & (!g1106) & (g1099)) + ((g1124) & (!g1125) & (!g1126) & (g1127) & (g1106) & (!g1099)) + ((g1124) & (!g1125) & (g1126) & (!g1127) & (!g1106) & (!g1099)) + ((g1124) & (!g1125) & (g1126) & (!g1127) & (g1106) & (!g1099)) + ((g1124) & (!g1125) & (g1126) & (!g1127) & (g1106) & (g1099)) + ((g1124) & (!g1125) & (g1126) & (g1127) & (!g1106) & (!g1099)) + ((g1124) & (!g1125) & (g1126) & (g1127) & (g1106) & (!g1099)) + ((g1124) & (g1125) & (!g1126) & (!g1127) & (!g1106) & (!g1099)) + ((g1124) & (g1125) & (!g1126) & (!g1127) & (!g1106) & (g1099)) + ((g1124) & (g1125) & (!g1126) & (!g1127) & (g1106) & (g1099)) + ((g1124) & (g1125) & (!g1126) & (g1127) & (!g1106) & (!g1099)) + ((g1124) & (g1125) & (!g1126) & (g1127) & (!g1106) & (g1099)) + ((g1124) & (g1125) & (g1126) & (!g1127) & (!g1106) & (!g1099)) + ((g1124) & (g1125) & (g1126) & (!g1127) & (g1106) & (g1099)) + ((g1124) & (g1125) & (g1126) & (g1127) & (!g1106) & (!g1099)));
	assign g1130 = (((!sk[104]) & (g1128) & (!g1129)) + ((!sk[104]) & (g1128) & (g1129)) + ((sk[104]) & (!g1128) & (g1129)) + ((sk[104]) & (g1128) & (!g1129)));
	assign g1131 = (((!g1095) & (!g1096) & (!g1099) & (!g1106) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1106) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1106) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1106) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1106) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1106) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1099) & (!g1106) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1099) & (!g1106) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1106) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1106) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1106) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (g1106) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (g1106) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1106) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1106) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1106) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1106) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1099) & (g1106) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1099) & (g1106) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (g1106) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1106) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1106) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (g1106) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (!g1106) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (!g1106) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (g1099) & (g1106) & (!g1105) & (g1100)));
	assign g1132 = (((!g1095) & (!g1096) & (!g1099) & (!g1106) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1099) & (!g1106) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (!g1099) & (!g1106) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1099) & (!g1106) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (!g1099) & (g1106) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1106) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1106) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1106) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1106) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (!g1106) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1106) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1106) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1106) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1106) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1106) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (g1106) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (g1106) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1106) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1106) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1106) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1106) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1106) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1106) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1106) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (g1106) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1106) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1106) & (g1105) & (g1100)) + ((g1095) & (g1096) & (!g1099) & (g1106) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (g1106) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (g1099) & (!g1106) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (!g1106) & (g1105) & (g1100)) + ((g1095) & (g1096) & (g1099) & (g1106) & (!g1105) & (g1100)));
	assign g1133 = (((!g1095) & (!g1096) & (!g1099) & (!g1106) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1099) & (!g1106) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1106) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1106) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1106) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1106) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1106) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1106) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1106) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1106) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1106) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (g1106) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (g1106) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1106) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1106) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1106) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1106) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1106) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1106) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1106) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (g1106) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1099) & (g1106) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (g1106) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1099) & (g1106) & (g1105) & (g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1106) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (!g1099) & (g1106) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (g1106) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (!g1106) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (!g1106) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (g1099) & (!g1106) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (g1106) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (g1106) & (g1105) & (!g1100)));
	assign g1134 = (((!g1095) & (!g1096) & (!g1099) & (!g1106) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (!g1099) & (g1106) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1099) & (g1106) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1106) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1106) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1106) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1106) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1106) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1099) & (!g1106) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1106) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1106) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1106) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1106) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (g1106) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (g1106) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1106) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1106) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1106) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1106) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1099) & (g1106) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1106) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (g1106) & (g1105) & (g1100)) + ((g1095) & (g1096) & (g1099) & (!g1106) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (!g1106) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (g1099) & (!g1106) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (g1106) & (!g1105) & (!g1100)));
	assign g1135 = (((!g1131) & (!g1132) & (!g1133) & (!g1134) & (g1097) & (g1098)) + ((!g1131) & (!g1132) & (g1133) & (!g1134) & (!g1097) & (g1098)) + ((!g1131) & (!g1132) & (g1133) & (!g1134) & (g1097) & (g1098)) + ((!g1131) & (!g1132) & (g1133) & (g1134) & (!g1097) & (g1098)) + ((!g1131) & (g1132) & (!g1133) & (!g1134) & (g1097) & (!g1098)) + ((!g1131) & (g1132) & (!g1133) & (!g1134) & (g1097) & (g1098)) + ((!g1131) & (g1132) & (!g1133) & (g1134) & (g1097) & (!g1098)) + ((!g1131) & (g1132) & (g1133) & (!g1134) & (!g1097) & (g1098)) + ((!g1131) & (g1132) & (g1133) & (!g1134) & (g1097) & (!g1098)) + ((!g1131) & (g1132) & (g1133) & (!g1134) & (g1097) & (g1098)) + ((!g1131) & (g1132) & (g1133) & (g1134) & (!g1097) & (g1098)) + ((!g1131) & (g1132) & (g1133) & (g1134) & (g1097) & (!g1098)) + ((g1131) & (!g1132) & (!g1133) & (!g1134) & (!g1097) & (!g1098)) + ((g1131) & (!g1132) & (!g1133) & (!g1134) & (g1097) & (g1098)) + ((g1131) & (!g1132) & (!g1133) & (g1134) & (!g1097) & (!g1098)) + ((g1131) & (!g1132) & (g1133) & (!g1134) & (!g1097) & (!g1098)) + ((g1131) & (!g1132) & (g1133) & (!g1134) & (!g1097) & (g1098)) + ((g1131) & (!g1132) & (g1133) & (!g1134) & (g1097) & (g1098)) + ((g1131) & (!g1132) & (g1133) & (g1134) & (!g1097) & (!g1098)) + ((g1131) & (!g1132) & (g1133) & (g1134) & (!g1097) & (g1098)) + ((g1131) & (g1132) & (!g1133) & (!g1134) & (!g1097) & (!g1098)) + ((g1131) & (g1132) & (!g1133) & (!g1134) & (g1097) & (!g1098)) + ((g1131) & (g1132) & (!g1133) & (!g1134) & (g1097) & (g1098)) + ((g1131) & (g1132) & (!g1133) & (g1134) & (!g1097) & (!g1098)) + ((g1131) & (g1132) & (!g1133) & (g1134) & (g1097) & (!g1098)) + ((g1131) & (g1132) & (g1133) & (!g1134) & (!g1097) & (!g1098)) + ((g1131) & (g1132) & (g1133) & (!g1134) & (!g1097) & (g1098)) + ((g1131) & (g1132) & (g1133) & (!g1134) & (g1097) & (!g1098)) + ((g1131) & (g1132) & (g1133) & (!g1134) & (g1097) & (g1098)) + ((g1131) & (g1132) & (g1133) & (g1134) & (!g1097) & (!g1098)) + ((g1131) & (g1132) & (g1133) & (g1134) & (!g1097) & (g1098)) + ((g1131) & (g1132) & (g1133) & (g1134) & (g1097) & (!g1098)));
	assign g1137 = (((!g1135) & (sk[110]) & (g1136)) + ((g1135) & (!sk[110]) & (!g1136)) + ((g1135) & (!sk[110]) & (g1136)) + ((g1135) & (sk[110]) & (!g1136)));
	assign g1138 = (((!g1095) & (!g1096) & (!g1099) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1099) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (!g1099) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1099) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (g1096) & (g1099) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (!g1098) & (g1105) & (g1100)));
	assign g1139 = (((!g1095) & (!g1096) & (!g1099) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1099) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1099) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (!g1099) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1099) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1099) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (g1098) & (g1105) & (g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (g1099) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (g1096) & (g1099) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (g1098) & (g1105) & (g1100)));
	assign g1140 = (((!g1095) & (!g1096) & (!g1099) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (!g1099) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (!g1099) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (g1096) & (!g1099) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (!g1099) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (g1099) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (g1096) & (g1099) & (g1098) & (g1105) & (g1100)));
	assign g1141 = (((!g1095) & (!g1096) & (!g1099) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1099) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1096) & (!g1099) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1096) & (g1099) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (!g1099) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1096) & (g1099) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1096) & (g1099) & (g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (!g1099) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1096) & (!g1099) & (g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1096) & (g1099) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1096) & (g1099) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (g1096) & (!g1099) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1096) & (!g1099) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (g1096) & (g1099) & (!g1098) & (g1105) & (g1100)));
	assign g1142 = (((!g1138) & (!g1139) & (!g1140) & (!g1141) & (!g1106) & (!g1097)) + ((!g1138) & (!g1139) & (!g1140) & (!g1141) & (!g1106) & (g1097)) + ((!g1138) & (!g1139) & (!g1140) & (!g1141) & (g1106) & (!g1097)) + ((!g1138) & (!g1139) & (!g1140) & (g1141) & (!g1106) & (!g1097)) + ((!g1138) & (!g1139) & (!g1140) & (g1141) & (!g1106) & (g1097)) + ((!g1138) & (!g1139) & (!g1140) & (g1141) & (g1106) & (!g1097)) + ((!g1138) & (!g1139) & (!g1140) & (g1141) & (g1106) & (g1097)) + ((!g1138) & (!g1139) & (g1140) & (!g1141) & (!g1106) & (!g1097)) + ((!g1138) & (!g1139) & (g1140) & (!g1141) & (g1106) & (!g1097)) + ((!g1138) & (!g1139) & (g1140) & (g1141) & (!g1106) & (!g1097)) + ((!g1138) & (!g1139) & (g1140) & (g1141) & (g1106) & (!g1097)) + ((!g1138) & (!g1139) & (g1140) & (g1141) & (g1106) & (g1097)) + ((!g1138) & (g1139) & (!g1140) & (!g1141) & (!g1106) & (!g1097)) + ((!g1138) & (g1139) & (!g1140) & (!g1141) & (!g1106) & (g1097)) + ((!g1138) & (g1139) & (!g1140) & (g1141) & (!g1106) & (!g1097)) + ((!g1138) & (g1139) & (!g1140) & (g1141) & (!g1106) & (g1097)) + ((!g1138) & (g1139) & (!g1140) & (g1141) & (g1106) & (g1097)) + ((!g1138) & (g1139) & (g1140) & (!g1141) & (!g1106) & (!g1097)) + ((!g1138) & (g1139) & (g1140) & (g1141) & (!g1106) & (!g1097)) + ((!g1138) & (g1139) & (g1140) & (g1141) & (g1106) & (g1097)) + ((g1138) & (!g1139) & (!g1140) & (!g1141) & (!g1106) & (g1097)) + ((g1138) & (!g1139) & (!g1140) & (!g1141) & (g1106) & (!g1097)) + ((g1138) & (!g1139) & (!g1140) & (g1141) & (!g1106) & (g1097)) + ((g1138) & (!g1139) & (!g1140) & (g1141) & (g1106) & (!g1097)) + ((g1138) & (!g1139) & (!g1140) & (g1141) & (g1106) & (g1097)) + ((g1138) & (!g1139) & (g1140) & (!g1141) & (g1106) & (!g1097)) + ((g1138) & (!g1139) & (g1140) & (g1141) & (g1106) & (!g1097)) + ((g1138) & (!g1139) & (g1140) & (g1141) & (g1106) & (g1097)) + ((g1138) & (g1139) & (!g1140) & (!g1141) & (!g1106) & (g1097)) + ((g1138) & (g1139) & (!g1140) & (g1141) & (!g1106) & (g1097)) + ((g1138) & (g1139) & (!g1140) & (g1141) & (g1106) & (g1097)) + ((g1138) & (g1139) & (g1140) & (g1141) & (g1106) & (g1097)));
	assign g1144 = (((!sk[116]) & (g1142) & (!g1143)) + ((!sk[116]) & (g1142) & (g1143)) + ((sk[116]) & (!g1142) & (g1143)) + ((sk[116]) & (g1142) & (!g1143)));
	assign g1145 = (((!g1095) & (!g1106) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1106) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1106) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1106) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1106) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1106) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1106) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1106) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1106) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1106) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1106) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (g1106) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1106) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1106) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1106) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1106) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((g1095) & (!g1106) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1106) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1106) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1106) & (g1097) & (g1098) & (g1105) & (g1100)) + ((g1095) & (g1106) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1106) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (g1106) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (g1106) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1106) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1106) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (g1106) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (g1106) & (g1097) & (g1098) & (!g1105) & (g1100)));
	assign g1146 = (((!g1095) & (!g1106) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1106) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1106) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1106) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1106) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1106) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1106) & (g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1106) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1106) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (g1106) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1106) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1106) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (g1106) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1106) & (g1097) & (g1098) & (g1105) & (g1100)) + ((g1095) & (!g1106) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1106) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1106) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1106) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((g1095) & (!g1106) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1106) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (g1106) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (g1106) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (g1106) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (g1106) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (g1106) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((g1095) & (g1106) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1106) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (g1106) & (g1097) & (g1098) & (!g1105) & (!g1100)));
	assign g1147 = (((!g1095) & (!g1106) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1106) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1106) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1106) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1106) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1106) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1106) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (!g1106) & (g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1106) & (!g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1106) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1106) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (g1106) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1106) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1106) & (g1097) & (!g1098) & (!g1105) & (g1100)) + ((!g1095) & (g1106) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1106) & (g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1106) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1106) & (g1097) & (g1098) & (g1105) & (g1100)) + ((g1095) & (!g1106) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1106) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (!g1106) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1106) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1106) & (g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (g1106) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (g1106) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1106) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (g1106) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1106) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (g1106) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (g1106) & (g1097) & (g1098) & (g1105) & (g1100)));
	assign g1148 = (((!g1095) & (!g1106) & (!g1097) & (!g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1106) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1106) & (!g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (!g1106) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((!g1095) & (!g1106) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (!g1106) & (g1097) & (g1098) & (g1105) & (g1100)) + ((!g1095) & (g1106) & (!g1097) & (g1098) & (!g1105) & (!g1100)) + ((!g1095) & (g1106) & (!g1097) & (g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1106) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((!g1095) & (g1106) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1106) & (!g1097) & (!g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1106) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1106) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (!g1106) & (g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1106) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (!g1106) & (g1097) & (g1098) & (g1105) & (!g1100)) + ((g1095) & (!g1106) & (g1097) & (g1098) & (g1105) & (g1100)) + ((g1095) & (g1106) & (!g1097) & (!g1098) & (g1105) & (!g1100)) + ((g1095) & (g1106) & (!g1097) & (g1098) & (!g1105) & (g1100)) + ((g1095) & (g1106) & (g1097) & (!g1098) & (!g1105) & (!g1100)) + ((g1095) & (g1106) & (g1097) & (!g1098) & (g1105) & (g1100)) + ((g1095) & (g1106) & (g1097) & (g1098) & (!g1105) & (g1100)));
	assign g1149 = (((!g1145) & (!g1146) & (!g1147) & (!g1148) & (!g1099) & (!g1096)) + ((!g1145) & (!g1146) & (!g1147) & (!g1148) & (!g1099) & (g1096)) + ((!g1145) & (!g1146) & (!g1147) & (!g1148) & (g1099) & (!g1096)) + ((!g1145) & (!g1146) & (!g1147) & (g1148) & (!g1099) & (!g1096)) + ((!g1145) & (!g1146) & (!g1147) & (g1148) & (!g1099) & (g1096)) + ((!g1145) & (!g1146) & (!g1147) & (g1148) & (g1099) & (!g1096)) + ((!g1145) & (!g1146) & (!g1147) & (g1148) & (g1099) & (g1096)) + ((!g1145) & (!g1146) & (g1147) & (!g1148) & (!g1099) & (!g1096)) + ((!g1145) & (!g1146) & (g1147) & (!g1148) & (g1099) & (!g1096)) + ((!g1145) & (!g1146) & (g1147) & (g1148) & (!g1099) & (!g1096)) + ((!g1145) & (!g1146) & (g1147) & (g1148) & (g1099) & (!g1096)) + ((!g1145) & (!g1146) & (g1147) & (g1148) & (g1099) & (g1096)) + ((!g1145) & (g1146) & (!g1147) & (!g1148) & (!g1099) & (!g1096)) + ((!g1145) & (g1146) & (!g1147) & (!g1148) & (!g1099) & (g1096)) + ((!g1145) & (g1146) & (!g1147) & (g1148) & (!g1099) & (!g1096)) + ((!g1145) & (g1146) & (!g1147) & (g1148) & (!g1099) & (g1096)) + ((!g1145) & (g1146) & (!g1147) & (g1148) & (g1099) & (g1096)) + ((!g1145) & (g1146) & (g1147) & (!g1148) & (!g1099) & (!g1096)) + ((!g1145) & (g1146) & (g1147) & (g1148) & (!g1099) & (!g1096)) + ((!g1145) & (g1146) & (g1147) & (g1148) & (g1099) & (g1096)) + ((g1145) & (!g1146) & (!g1147) & (!g1148) & (!g1099) & (g1096)) + ((g1145) & (!g1146) & (!g1147) & (!g1148) & (g1099) & (!g1096)) + ((g1145) & (!g1146) & (!g1147) & (g1148) & (!g1099) & (g1096)) + ((g1145) & (!g1146) & (!g1147) & (g1148) & (g1099) & (!g1096)) + ((g1145) & (!g1146) & (!g1147) & (g1148) & (g1099) & (g1096)) + ((g1145) & (!g1146) & (g1147) & (!g1148) & (g1099) & (!g1096)) + ((g1145) & (!g1146) & (g1147) & (g1148) & (g1099) & (!g1096)) + ((g1145) & (!g1146) & (g1147) & (g1148) & (g1099) & (g1096)) + ((g1145) & (g1146) & (!g1147) & (!g1148) & (!g1099) & (g1096)) + ((g1145) & (g1146) & (!g1147) & (g1148) & (!g1099) & (g1096)) + ((g1145) & (g1146) & (!g1147) & (g1148) & (g1099) & (g1096)) + ((g1145) & (g1146) & (g1147) & (g1148) & (g1099) & (g1096)));
	assign g1151 = (((!sk[122]) & (g1149) & (!g1150)) + ((!sk[122]) & (g1149) & (g1150)) + ((sk[122]) & (!g1149) & (g1150)) + ((sk[122]) & (g1149) & (!g1150)));
	assign g1152 = (((!g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1106)) + ((!g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1106)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1106)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (!g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1106)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1106)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1106)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1106)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1106)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1106)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1106)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1106)) + ((g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1106)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1106)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1106)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1106)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1106)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1106)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1106)) + ((g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1106)));
	assign g1153 = (((!g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1106)) + ((!g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1106)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (g1105) & (g1106)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1106)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1106)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1106)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1106)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1106)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (g1106)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1106)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1106)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1106)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1106)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1106)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (g1106)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1106)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1106)) + ((g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1106)) + ((g1099) & (!g1096) & (g1097) & (!g1098) & (g1105) & (g1106)) + ((g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1106)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1106)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (g1106)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1106)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (g1106)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1106)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1106)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1106)));
	assign g1154 = (((!g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1106)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1106)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1106)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1106)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (g1106)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (!g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1106)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (g1106)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1106)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1106)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1106)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1106)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1106)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1106)) + ((g1099) & (!g1096) & (!g1097) & (!g1098) & (g1105) & (!g1106)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (!g1106)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1106)) + ((g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1106)) + ((g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (g1106)) + ((g1099) & (!g1096) & (g1097) & (g1098) & (!g1105) & (!g1106)) + ((g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1106)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (g1105) & (!g1106)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1106)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1106)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (!g1105) & (!g1106)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (!g1106)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1106)) + ((g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1106)));
	assign g1155 = (((!g1099) & (!g1096) & (!g1097) & (!g1098) & (!g1105) & (g1106)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (!g1106)) + ((!g1099) & (!g1096) & (!g1097) & (g1098) & (g1105) & (g1106)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (g1106)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (!g1106)) + ((!g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1106)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (!g1106)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (g1106)) + ((!g1099) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1106)) + ((!g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (g1106)) + ((!g1099) & (g1096) & (g1097) & (!g1098) & (!g1105) & (g1106)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (!g1106)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (!g1105) & (g1106)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (g1105) & (!g1106)) + ((!g1099) & (g1096) & (g1097) & (g1098) & (g1105) & (g1106)) + ((g1099) & (!g1096) & (!g1097) & (g1098) & (!g1105) & (g1106)) + ((g1099) & (!g1096) & (g1097) & (!g1098) & (!g1105) & (!g1106)) + ((g1099) & (!g1096) & (g1097) & (g1098) & (!g1105) & (!g1106)) + ((g1099) & (!g1096) & (g1097) & (g1098) & (!g1105) & (g1106)) + ((g1099) & (!g1096) & (g1097) & (g1098) & (g1105) & (g1106)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (!g1105) & (g1106)) + ((g1099) & (g1096) & (!g1097) & (!g1098) & (g1105) & (g1106)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (!g1105) & (!g1106)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (!g1106)) + ((g1099) & (g1096) & (!g1097) & (g1098) & (g1105) & (g1106)) + ((g1099) & (g1096) & (g1097) & (!g1098) & (g1105) & (g1106)) + ((g1099) & (g1096) & (g1097) & (g1098) & (g1105) & (g1106)));
	assign g1156 = (((!g1152) & (!g1153) & (!g1154) & (!g1155) & (!g1095) & (g1100)) + ((!g1152) & (!g1153) & (!g1154) & (!g1155) & (g1095) & (!g1100)) + ((!g1152) & (!g1153) & (!g1154) & (!g1155) & (g1095) & (g1100)) + ((!g1152) & (!g1153) & (!g1154) & (g1155) & (!g1095) & (g1100)) + ((!g1152) & (!g1153) & (!g1154) & (g1155) & (g1095) & (!g1100)) + ((!g1152) & (!g1153) & (g1154) & (!g1155) & (g1095) & (!g1100)) + ((!g1152) & (!g1153) & (g1154) & (!g1155) & (g1095) & (g1100)) + ((!g1152) & (!g1153) & (g1154) & (g1155) & (g1095) & (!g1100)) + ((!g1152) & (g1153) & (!g1154) & (!g1155) & (!g1095) & (g1100)) + ((!g1152) & (g1153) & (!g1154) & (!g1155) & (g1095) & (g1100)) + ((!g1152) & (g1153) & (!g1154) & (g1155) & (!g1095) & (g1100)) + ((!g1152) & (g1153) & (g1154) & (!g1155) & (g1095) & (g1100)) + ((g1152) & (!g1153) & (!g1154) & (!g1155) & (!g1095) & (!g1100)) + ((g1152) & (!g1153) & (!g1154) & (!g1155) & (!g1095) & (g1100)) + ((g1152) & (!g1153) & (!g1154) & (!g1155) & (g1095) & (!g1100)) + ((g1152) & (!g1153) & (!g1154) & (!g1155) & (g1095) & (g1100)) + ((g1152) & (!g1153) & (!g1154) & (g1155) & (!g1095) & (!g1100)) + ((g1152) & (!g1153) & (!g1154) & (g1155) & (!g1095) & (g1100)) + ((g1152) & (!g1153) & (!g1154) & (g1155) & (g1095) & (!g1100)) + ((g1152) & (!g1153) & (g1154) & (!g1155) & (!g1095) & (!g1100)) + ((g1152) & (!g1153) & (g1154) & (!g1155) & (g1095) & (!g1100)) + ((g1152) & (!g1153) & (g1154) & (!g1155) & (g1095) & (g1100)) + ((g1152) & (!g1153) & (g1154) & (g1155) & (!g1095) & (!g1100)) + ((g1152) & (!g1153) & (g1154) & (g1155) & (g1095) & (!g1100)) + ((g1152) & (g1153) & (!g1154) & (!g1155) & (!g1095) & (!g1100)) + ((g1152) & (g1153) & (!g1154) & (!g1155) & (!g1095) & (g1100)) + ((g1152) & (g1153) & (!g1154) & (!g1155) & (g1095) & (g1100)) + ((g1152) & (g1153) & (!g1154) & (g1155) & (!g1095) & (!g1100)) + ((g1152) & (g1153) & (!g1154) & (g1155) & (!g1095) & (g1100)) + ((g1152) & (g1153) & (g1154) & (!g1155) & (!g1095) & (!g1100)) + ((g1152) & (g1153) & (g1154) & (!g1155) & (g1095) & (g1100)) + ((g1152) & (g1153) & (g1154) & (g1155) & (!g1095) & (!g1100)));
	assign g1158 = (((!g1156) & (sk[0]) & (g1157)) + ((g1156) & (!sk[0]) & (!g1157)) + ((g1156) & (!sk[0]) & (g1157)) + ((g1156) & (sk[0]) & (!g1157)));
	assign g1159 = (((!g130) & (!g131) & (!g132) & (!g133) & (ld) & (rst)) + ((!g130) & (!g131) & (!g132) & (g133) & (!ld) & (rst)) + ((!g130) & (!g131) & (!g132) & (g133) & (ld) & (rst)) + ((!g130) & (!g131) & (g132) & (!g133) & (!ld) & (rst)) + ((!g130) & (!g131) & (g132) & (!g133) & (ld) & (rst)) + ((!g130) & (!g131) & (g132) & (g133) & (!ld) & (rst)) + ((!g130) & (!g131) & (g132) & (g133) & (ld) & (rst)) + ((!g130) & (g131) & (!g132) & (!g133) & (!ld) & (rst)) + ((!g130) & (g131) & (!g132) & (!g133) & (ld) & (rst)) + ((!g130) & (g131) & (!g132) & (g133) & (!ld) & (rst)) + ((!g130) & (g131) & (!g132) & (g133) & (ld) & (rst)) + ((!g130) & (g131) & (g132) & (!g133) & (!ld) & (rst)) + ((!g130) & (g131) & (g132) & (!g133) & (ld) & (rst)) + ((!g130) & (g131) & (g132) & (g133) & (!ld) & (rst)) + ((!g130) & (g131) & (g132) & (g133) & (ld) & (rst)) + ((g130) & (!g131) & (!g132) & (!g133) & (ld) & (rst)) + ((g130) & (!g131) & (!g132) & (g133) & (ld) & (rst)) + ((g130) & (!g131) & (g132) & (!g133) & (ld) & (rst)) + ((g130) & (!g131) & (g132) & (g133) & (ld) & (rst)) + ((g130) & (g131) & (!g132) & (!g133) & (ld) & (rst)) + ((g130) & (g131) & (!g132) & (g133) & (ld) & (rst)) + ((g130) & (g131) & (g132) & (!g133) & (ld) & (rst)) + ((g130) & (g131) & (g132) & (g133) & (ld) & (rst)));
	assign g1160 = (((!g130) & (!g131) & (!g132) & (!g133) & (ld) & (rst)) + ((!g130) & (!g131) & (!g132) & (g133) & (!ld) & (rst)) + ((!g130) & (!g131) & (!g132) & (g133) & (ld) & (rst)) + ((!g130) & (!g131) & (g132) & (!g133) & (!ld) & (rst)) + ((!g130) & (!g131) & (g132) & (!g133) & (ld) & (rst)) + ((!g130) & (!g131) & (g132) & (g133) & (!ld) & (rst)) + ((!g130) & (!g131) & (g132) & (g133) & (ld) & (rst)) + ((!g130) & (g131) & (!g132) & (!g133) & (ld) & (rst)) + ((!g130) & (g131) & (!g132) & (g133) & (ld) & (rst)) + ((!g130) & (g131) & (g132) & (!g133) & (ld) & (rst)) + ((!g130) & (g131) & (g132) & (g133) & (ld) & (rst)) + ((g130) & (!g131) & (!g132) & (!g133) & (ld) & (rst)) + ((g130) & (!g131) & (!g132) & (g133) & (ld) & (rst)) + ((g130) & (!g131) & (g132) & (!g133) & (ld) & (rst)) + ((g130) & (!g131) & (g132) & (g133) & (ld) & (rst)) + ((g130) & (g131) & (!g132) & (!g133) & (!ld) & (rst)) + ((g130) & (g131) & (!g132) & (!g133) & (ld) & (rst)) + ((g130) & (g131) & (!g132) & (g133) & (!ld) & (rst)) + ((g130) & (g131) & (!g132) & (g133) & (ld) & (rst)) + ((g130) & (g131) & (g132) & (!g133) & (!ld) & (rst)) + ((g130) & (g131) & (g132) & (!g133) & (ld) & (rst)) + ((g130) & (g131) & (g132) & (g133) & (!ld) & (rst)) + ((g130) & (g131) & (g132) & (g133) & (ld) & (rst)));
	assign g1161 = (((!g130) & (!g131) & (!g132) & (g133) & (!ld) & (rst)) + ((!g130) & (g131) & (g132) & (!g133) & (!ld) & (rst)) + ((!g130) & (g131) & (g132) & (g133) & (!ld) & (rst)) + ((g130) & (!g131) & (g132) & (!g133) & (!ld) & (rst)) + ((g130) & (!g131) & (g132) & (g133) & (!ld) & (rst)) + ((g130) & (g131) & (g132) & (!g133) & (!ld) & (rst)) + ((g130) & (g131) & (g132) & (g133) & (!ld) & (rst)));
	assign g1162 = (((!g130) & (!g131) & (!g132) & (!g133) & (ld) & (rst)) + ((!g130) & (!g131) & (!g132) & (g133) & (ld) & (rst)) + ((!g130) & (!g131) & (g132) & (!g133) & (ld) & (rst)) + ((!g130) & (!g131) & (g132) & (g133) & (!ld) & (rst)) + ((!g130) & (!g131) & (g132) & (g133) & (ld) & (rst)) + ((!g130) & (g131) & (!g132) & (!g133) & (ld) & (rst)) + ((!g130) & (g131) & (!g132) & (g133) & (!ld) & (rst)) + ((!g130) & (g131) & (!g132) & (g133) & (ld) & (rst)) + ((!g130) & (g131) & (g132) & (!g133) & (ld) & (rst)) + ((!g130) & (g131) & (g132) & (g133) & (!ld) & (rst)) + ((!g130) & (g131) & (g132) & (g133) & (ld) & (rst)) + ((g130) & (!g131) & (!g132) & (!g133) & (ld) & (rst)) + ((g130) & (!g131) & (!g132) & (g133) & (!ld) & (rst)) + ((g130) & (!g131) & (!g132) & (g133) & (ld) & (rst)) + ((g130) & (!g131) & (g132) & (!g133) & (ld) & (rst)) + ((g130) & (!g131) & (g132) & (g133) & (!ld) & (rst)) + ((g130) & (!g131) & (g132) & (g133) & (ld) & (rst)) + ((g130) & (g131) & (!g132) & (!g133) & (ld) & (rst)) + ((g130) & (g131) & (!g132) & (g133) & (!ld) & (rst)) + ((g130) & (g131) & (!g132) & (g133) & (ld) & (rst)) + ((g130) & (g131) & (g132) & (!g133) & (ld) & (rst)) + ((g130) & (g131) & (g132) & (g133) & (!ld) & (rst)) + ((g130) & (g131) & (g132) & (g133) & (ld) & (rst)));
	assign g2082 = (((!ld) & (!sk[5]) & (text_inx32x) & (!g1164)) + ((!ld) & (!sk[5]) & (text_inx32x) & (g1164)) + ((!ld) & (sk[5]) & (!text_inx32x) & (g1164)) + ((!ld) & (sk[5]) & (text_inx32x) & (g1164)) + ((ld) & (!sk[5]) & (!text_inx32x) & (!g1164)) + ((ld) & (!sk[5]) & (!text_inx32x) & (g1164)) + ((ld) & (!sk[5]) & (text_inx32x) & (!g1164)) + ((ld) & (!sk[5]) & (text_inx32x) & (g1164)) + ((ld) & (sk[5]) & (text_inx32x) & (!g1164)) + ((ld) & (sk[5]) & (text_inx32x) & (g1164)));
	assign g1165 = (((!sk[6]) & (!g404) & (!g452) & (g467) & (!g644)) + ((!sk[6]) & (!g404) & (!g452) & (g467) & (g644)) + ((!sk[6]) & (!g404) & (g452) & (!g467) & (!g644)) + ((!sk[6]) & (!g404) & (g452) & (!g467) & (g644)) + ((!sk[6]) & (!g404) & (g452) & (g467) & (!g644)) + ((!sk[6]) & (!g404) & (g452) & (g467) & (g644)) + ((!sk[6]) & (g404) & (!g452) & (g467) & (!g644)) + ((!sk[6]) & (g404) & (!g452) & (g467) & (g644)) + ((!sk[6]) & (g404) & (g452) & (!g467) & (!g644)) + ((!sk[6]) & (g404) & (g452) & (!g467) & (g644)) + ((!sk[6]) & (g404) & (g452) & (g467) & (!g644)) + ((!sk[6]) & (g404) & (g452) & (g467) & (g644)) + ((sk[6]) & (!g404) & (!g452) & (!g467) & (g644)) + ((sk[6]) & (!g404) & (!g452) & (g467) & (!g644)) + ((sk[6]) & (!g404) & (g452) & (!g467) & (!g644)) + ((sk[6]) & (!g404) & (g452) & (g467) & (g644)) + ((sk[6]) & (g404) & (!g452) & (!g467) & (!g644)) + ((sk[6]) & (g404) & (!g452) & (g467) & (g644)) + ((sk[6]) & (g404) & (g452) & (!g467) & (g644)) + ((sk[6]) & (g404) & (g452) & (g467) & (!g644)));
	assign g1166 = (((!g404) & (!g531) & (!g595) & (!g1163) & (!g1164) & (g1165)) + ((!g404) & (!g531) & (!g595) & (!g1163) & (g1164) & (g1165)) + ((!g404) & (!g531) & (!g595) & (g1163) & (g1164) & (!g1165)) + ((!g404) & (!g531) & (!g595) & (g1163) & (g1164) & (g1165)) + ((!g404) & (!g531) & (g595) & (!g1163) & (!g1164) & (!g1165)) + ((!g404) & (!g531) & (g595) & (!g1163) & (g1164) & (!g1165)) + ((!g404) & (!g531) & (g595) & (g1163) & (g1164) & (!g1165)) + ((!g404) & (!g531) & (g595) & (g1163) & (g1164) & (g1165)) + ((!g404) & (g531) & (!g595) & (!g1163) & (!g1164) & (!g1165)) + ((!g404) & (g531) & (!g595) & (!g1163) & (g1164) & (!g1165)) + ((!g404) & (g531) & (!g595) & (g1163) & (g1164) & (!g1165)) + ((!g404) & (g531) & (!g595) & (g1163) & (g1164) & (g1165)) + ((!g404) & (g531) & (g595) & (!g1163) & (!g1164) & (g1165)) + ((!g404) & (g531) & (g595) & (!g1163) & (g1164) & (g1165)) + ((!g404) & (g531) & (g595) & (g1163) & (g1164) & (!g1165)) + ((!g404) & (g531) & (g595) & (g1163) & (g1164) & (g1165)) + ((g404) & (!g531) & (!g595) & (!g1163) & (!g1164) & (g1165)) + ((g404) & (!g531) & (!g595) & (!g1163) & (g1164) & (g1165)) + ((g404) & (!g531) & (!g595) & (g1163) & (!g1164) & (!g1165)) + ((g404) & (!g531) & (!g595) & (g1163) & (!g1164) & (g1165)) + ((g404) & (!g531) & (g595) & (!g1163) & (!g1164) & (!g1165)) + ((g404) & (!g531) & (g595) & (!g1163) & (g1164) & (!g1165)) + ((g404) & (!g531) & (g595) & (g1163) & (!g1164) & (!g1165)) + ((g404) & (!g531) & (g595) & (g1163) & (!g1164) & (g1165)) + ((g404) & (g531) & (!g595) & (!g1163) & (!g1164) & (!g1165)) + ((g404) & (g531) & (!g595) & (!g1163) & (g1164) & (!g1165)) + ((g404) & (g531) & (!g595) & (g1163) & (!g1164) & (!g1165)) + ((g404) & (g531) & (!g595) & (g1163) & (!g1164) & (g1165)) + ((g404) & (g531) & (g595) & (!g1163) & (!g1164) & (g1165)) + ((g404) & (g531) & (g595) & (!g1163) & (g1164) & (g1165)) + ((g404) & (g531) & (g595) & (g1163) & (!g1164) & (!g1165)) + ((g404) & (g531) & (g595) & (g1163) & (!g1164) & (g1165)));
	assign g2083 = (((!ld) & (!sk[8]) & (text_inx33x) & (!g1167)) + ((!ld) & (!sk[8]) & (text_inx33x) & (g1167)) + ((!ld) & (sk[8]) & (!text_inx33x) & (g1167)) + ((!ld) & (sk[8]) & (text_inx33x) & (g1167)) + ((ld) & (!sk[8]) & (!text_inx33x) & (!g1167)) + ((ld) & (!sk[8]) & (!text_inx33x) & (g1167)) + ((ld) & (!sk[8]) & (text_inx33x) & (!g1167)) + ((ld) & (!sk[8]) & (text_inx33x) & (g1167)) + ((ld) & (sk[8]) & (text_inx33x) & (!g1167)) + ((ld) & (sk[8]) & (text_inx33x) & (g1167)));
	assign g1168 = (((!g474) & (!sk[9]) & (g538) & (!g595)) + ((!g474) & (!sk[9]) & (g538) & (g595)) + ((!g474) & (sk[9]) & (!g538) & (g595)) + ((!g474) & (sk[9]) & (g538) & (!g595)) + ((g474) & (!sk[9]) & (!g538) & (!g595)) + ((g474) & (!sk[9]) & (!g538) & (g595)) + ((g474) & (!sk[9]) & (g538) & (!g595)) + ((g474) & (!sk[9]) & (g538) & (g595)) + ((g474) & (sk[9]) & (!g538) & (!g595)) + ((g474) & (sk[9]) & (g538) & (g595)));
	assign g1169 = (((!g403) & (!g411) & (!g452) & (!sk[10]) & (!g602) & (g644)) + ((!g403) & (!g411) & (!g452) & (!sk[10]) & (g602) & (g644)) + ((!g403) & (!g411) & (!g452) & (sk[10]) & (!g602) & (g644)) + ((!g403) & (!g411) & (!g452) & (sk[10]) & (g602) & (!g644)) + ((!g403) & (!g411) & (g452) & (!sk[10]) & (!g602) & (g644)) + ((!g403) & (!g411) & (g452) & (!sk[10]) & (g602) & (g644)) + ((!g403) & (!g411) & (g452) & (sk[10]) & (!g602) & (!g644)) + ((!g403) & (!g411) & (g452) & (sk[10]) & (g602) & (g644)) + ((!g403) & (g411) & (!g452) & (!sk[10]) & (!g602) & (!g644)) + ((!g403) & (g411) & (!g452) & (!sk[10]) & (!g602) & (g644)) + ((!g403) & (g411) & (!g452) & (!sk[10]) & (g602) & (!g644)) + ((!g403) & (g411) & (!g452) & (!sk[10]) & (g602) & (g644)) + ((!g403) & (g411) & (!g452) & (sk[10]) & (!g602) & (!g644)) + ((!g403) & (g411) & (!g452) & (sk[10]) & (g602) & (g644)) + ((!g403) & (g411) & (g452) & (!sk[10]) & (!g602) & (!g644)) + ((!g403) & (g411) & (g452) & (!sk[10]) & (!g602) & (g644)) + ((!g403) & (g411) & (g452) & (!sk[10]) & (g602) & (!g644)) + ((!g403) & (g411) & (g452) & (!sk[10]) & (g602) & (g644)) + ((!g403) & (g411) & (g452) & (sk[10]) & (!g602) & (g644)) + ((!g403) & (g411) & (g452) & (sk[10]) & (g602) & (!g644)) + ((g403) & (!g411) & (!g452) & (!sk[10]) & (!g602) & (g644)) + ((g403) & (!g411) & (!g452) & (!sk[10]) & (g602) & (!g644)) + ((g403) & (!g411) & (!g452) & (!sk[10]) & (g602) & (g644)) + ((g403) & (!g411) & (!g452) & (sk[10]) & (!g602) & (!g644)) + ((g403) & (!g411) & (!g452) & (sk[10]) & (g602) & (g644)) + ((g403) & (!g411) & (g452) & (!sk[10]) & (!g602) & (g644)) + ((g403) & (!g411) & (g452) & (!sk[10]) & (g602) & (!g644)) + ((g403) & (!g411) & (g452) & (!sk[10]) & (g602) & (g644)) + ((g403) & (!g411) & (g452) & (sk[10]) & (!g602) & (g644)) + ((g403) & (!g411) & (g452) & (sk[10]) & (g602) & (!g644)) + ((g403) & (g411) & (!g452) & (!sk[10]) & (!g602) & (!g644)) + ((g403) & (g411) & (!g452) & (!sk[10]) & (!g602) & (g644)) + ((g403) & (g411) & (!g452) & (!sk[10]) & (g602) & (!g644)) + ((g403) & (g411) & (!g452) & (!sk[10]) & (g602) & (g644)) + ((g403) & (g411) & (!g452) & (sk[10]) & (!g602) & (g644)) + ((g403) & (g411) & (!g452) & (sk[10]) & (g602) & (!g644)) + ((g403) & (g411) & (g452) & (!sk[10]) & (!g602) & (!g644)) + ((g403) & (g411) & (g452) & (!sk[10]) & (!g602) & (g644)) + ((g403) & (g411) & (g452) & (!sk[10]) & (g602) & (!g644)) + ((g403) & (g411) & (g452) & (!sk[10]) & (g602) & (g644)) + ((g403) & (g411) & (g452) & (sk[10]) & (!g602) & (!g644)) + ((g403) & (g411) & (g452) & (sk[10]) & (g602) & (g644)));
	assign g1170 = (((!g411) & (!g1163) & (!sk[11]) & (!g1167) & (!g1168) & (g1169)) + ((!g411) & (!g1163) & (!sk[11]) & (!g1167) & (g1168) & (g1169)) + ((!g411) & (!g1163) & (!sk[11]) & (g1167) & (!g1168) & (g1169)) + ((!g411) & (!g1163) & (!sk[11]) & (g1167) & (g1168) & (g1169)) + ((!g411) & (!g1163) & (sk[11]) & (!g1167) & (!g1168) & (g1169)) + ((!g411) & (!g1163) & (sk[11]) & (!g1167) & (g1168) & (!g1169)) + ((!g411) & (!g1163) & (sk[11]) & (g1167) & (!g1168) & (g1169)) + ((!g411) & (!g1163) & (sk[11]) & (g1167) & (g1168) & (!g1169)) + ((!g411) & (g1163) & (!sk[11]) & (!g1167) & (!g1168) & (!g1169)) + ((!g411) & (g1163) & (!sk[11]) & (!g1167) & (!g1168) & (g1169)) + ((!g411) & (g1163) & (!sk[11]) & (!g1167) & (g1168) & (!g1169)) + ((!g411) & (g1163) & (!sk[11]) & (!g1167) & (g1168) & (g1169)) + ((!g411) & (g1163) & (!sk[11]) & (g1167) & (!g1168) & (!g1169)) + ((!g411) & (g1163) & (!sk[11]) & (g1167) & (!g1168) & (g1169)) + ((!g411) & (g1163) & (!sk[11]) & (g1167) & (g1168) & (!g1169)) + ((!g411) & (g1163) & (!sk[11]) & (g1167) & (g1168) & (g1169)) + ((!g411) & (g1163) & (sk[11]) & (g1167) & (!g1168) & (!g1169)) + ((!g411) & (g1163) & (sk[11]) & (g1167) & (!g1168) & (g1169)) + ((!g411) & (g1163) & (sk[11]) & (g1167) & (g1168) & (!g1169)) + ((!g411) & (g1163) & (sk[11]) & (g1167) & (g1168) & (g1169)) + ((g411) & (!g1163) & (!sk[11]) & (!g1167) & (!g1168) & (g1169)) + ((g411) & (!g1163) & (!sk[11]) & (!g1167) & (g1168) & (!g1169)) + ((g411) & (!g1163) & (!sk[11]) & (!g1167) & (g1168) & (g1169)) + ((g411) & (!g1163) & (!sk[11]) & (g1167) & (!g1168) & (g1169)) + ((g411) & (!g1163) & (!sk[11]) & (g1167) & (g1168) & (!g1169)) + ((g411) & (!g1163) & (!sk[11]) & (g1167) & (g1168) & (g1169)) + ((g411) & (!g1163) & (sk[11]) & (!g1167) & (!g1168) & (g1169)) + ((g411) & (!g1163) & (sk[11]) & (!g1167) & (g1168) & (!g1169)) + ((g411) & (!g1163) & (sk[11]) & (g1167) & (!g1168) & (g1169)) + ((g411) & (!g1163) & (sk[11]) & (g1167) & (g1168) & (!g1169)) + ((g411) & (g1163) & (!sk[11]) & (!g1167) & (!g1168) & (!g1169)) + ((g411) & (g1163) & (!sk[11]) & (!g1167) & (!g1168) & (g1169)) + ((g411) & (g1163) & (!sk[11]) & (!g1167) & (g1168) & (!g1169)) + ((g411) & (g1163) & (!sk[11]) & (!g1167) & (g1168) & (g1169)) + ((g411) & (g1163) & (!sk[11]) & (g1167) & (!g1168) & (!g1169)) + ((g411) & (g1163) & (!sk[11]) & (g1167) & (!g1168) & (g1169)) + ((g411) & (g1163) & (!sk[11]) & (g1167) & (g1168) & (!g1169)) + ((g411) & (g1163) & (!sk[11]) & (g1167) & (g1168) & (g1169)) + ((g411) & (g1163) & (sk[11]) & (!g1167) & (!g1168) & (!g1169)) + ((g411) & (g1163) & (sk[11]) & (!g1167) & (!g1168) & (g1169)) + ((g411) & (g1163) & (sk[11]) & (!g1167) & (g1168) & (!g1169)) + ((g411) & (g1163) & (sk[11]) & (!g1167) & (g1168) & (g1169)));
	assign g2084 = (((!ld) & (!text_inx34x) & (sk[12]) & (g1171)) + ((!ld) & (text_inx34x) & (!sk[12]) & (!g1171)) + ((!ld) & (text_inx34x) & (!sk[12]) & (g1171)) + ((!ld) & (text_inx34x) & (sk[12]) & (g1171)) + ((ld) & (!text_inx34x) & (!sk[12]) & (!g1171)) + ((ld) & (!text_inx34x) & (!sk[12]) & (g1171)) + ((ld) & (text_inx34x) & (!sk[12]) & (!g1171)) + ((ld) & (text_inx34x) & (!sk[12]) & (g1171)) + ((ld) & (text_inx34x) & (sk[12]) & (!g1171)) + ((ld) & (text_inx34x) & (sk[12]) & (g1171)));
	assign g1172 = (((!g410) & (!sk[13]) & (g545) & (!g609)) + ((!g410) & (!sk[13]) & (g545) & (g609)) + ((!g410) & (sk[13]) & (!g545) & (g609)) + ((!g410) & (sk[13]) & (g545) & (!g609)) + ((g410) & (!sk[13]) & (!g545) & (!g609)) + ((g410) & (!sk[13]) & (!g545) & (g609)) + ((g410) & (!sk[13]) & (g545) & (!g609)) + ((g410) & (!sk[13]) & (g545) & (g609)) + ((g410) & (sk[13]) & (!g545) & (!g609)) + ((g410) & (sk[13]) & (g545) & (g609)));
	assign g1173 = (((!g418) & (!g481) & (!g602) & (!g1163) & (!g1171) & (g1172)) + ((!g418) & (!g481) & (!g602) & (!g1163) & (g1171) & (g1172)) + ((!g418) & (!g481) & (!g602) & (g1163) & (g1171) & (!g1172)) + ((!g418) & (!g481) & (!g602) & (g1163) & (g1171) & (g1172)) + ((!g418) & (!g481) & (g602) & (!g1163) & (!g1171) & (!g1172)) + ((!g418) & (!g481) & (g602) & (!g1163) & (g1171) & (!g1172)) + ((!g418) & (!g481) & (g602) & (g1163) & (g1171) & (!g1172)) + ((!g418) & (!g481) & (g602) & (g1163) & (g1171) & (g1172)) + ((!g418) & (g481) & (!g602) & (!g1163) & (!g1171) & (!g1172)) + ((!g418) & (g481) & (!g602) & (!g1163) & (g1171) & (!g1172)) + ((!g418) & (g481) & (!g602) & (g1163) & (g1171) & (!g1172)) + ((!g418) & (g481) & (!g602) & (g1163) & (g1171) & (g1172)) + ((!g418) & (g481) & (g602) & (!g1163) & (!g1171) & (g1172)) + ((!g418) & (g481) & (g602) & (!g1163) & (g1171) & (g1172)) + ((!g418) & (g481) & (g602) & (g1163) & (g1171) & (!g1172)) + ((!g418) & (g481) & (g602) & (g1163) & (g1171) & (g1172)) + ((g418) & (!g481) & (!g602) & (!g1163) & (!g1171) & (!g1172)) + ((g418) & (!g481) & (!g602) & (!g1163) & (g1171) & (!g1172)) + ((g418) & (!g481) & (!g602) & (g1163) & (!g1171) & (!g1172)) + ((g418) & (!g481) & (!g602) & (g1163) & (!g1171) & (g1172)) + ((g418) & (!g481) & (g602) & (!g1163) & (!g1171) & (g1172)) + ((g418) & (!g481) & (g602) & (!g1163) & (g1171) & (g1172)) + ((g418) & (!g481) & (g602) & (g1163) & (!g1171) & (!g1172)) + ((g418) & (!g481) & (g602) & (g1163) & (!g1171) & (g1172)) + ((g418) & (g481) & (!g602) & (!g1163) & (!g1171) & (g1172)) + ((g418) & (g481) & (!g602) & (!g1163) & (g1171) & (g1172)) + ((g418) & (g481) & (!g602) & (g1163) & (!g1171) & (!g1172)) + ((g418) & (g481) & (!g602) & (g1163) & (!g1171) & (g1172)) + ((g418) & (g481) & (g602) & (!g1163) & (!g1171) & (!g1172)) + ((g418) & (g481) & (g602) & (!g1163) & (g1171) & (!g1172)) + ((g418) & (g481) & (g602) & (g1163) & (!g1171) & (!g1172)) + ((g418) & (g481) & (g602) & (g1163) & (!g1171) & (g1172)));
	assign g2085 = (((!ld) & (!sk[15]) & (text_inx35x) & (!g1174)) + ((!ld) & (!sk[15]) & (text_inx35x) & (g1174)) + ((!ld) & (sk[15]) & (!text_inx35x) & (g1174)) + ((!ld) & (sk[15]) & (text_inx35x) & (g1174)) + ((ld) & (!sk[15]) & (!text_inx35x) & (!g1174)) + ((ld) & (!sk[15]) & (!text_inx35x) & (g1174)) + ((ld) & (!sk[15]) & (text_inx35x) & (!g1174)) + ((ld) & (!sk[15]) & (text_inx35x) & (g1174)) + ((ld) & (sk[15]) & (text_inx35x) & (!g1174)) + ((ld) & (sk[15]) & (text_inx35x) & (g1174)));
	assign g1175 = (((!g488) & (!g552) & (!sk[16]) & (g609) & (!g644)) + ((!g488) & (!g552) & (!sk[16]) & (g609) & (g644)) + ((!g488) & (!g552) & (sk[16]) & (!g609) & (g644)) + ((!g488) & (!g552) & (sk[16]) & (g609) & (!g644)) + ((!g488) & (g552) & (!sk[16]) & (!g609) & (!g644)) + ((!g488) & (g552) & (!sk[16]) & (!g609) & (g644)) + ((!g488) & (g552) & (!sk[16]) & (g609) & (!g644)) + ((!g488) & (g552) & (!sk[16]) & (g609) & (g644)) + ((!g488) & (g552) & (sk[16]) & (!g609) & (!g644)) + ((!g488) & (g552) & (sk[16]) & (g609) & (g644)) + ((g488) & (!g552) & (!sk[16]) & (g609) & (!g644)) + ((g488) & (!g552) & (!sk[16]) & (g609) & (g644)) + ((g488) & (!g552) & (sk[16]) & (!g609) & (!g644)) + ((g488) & (!g552) & (sk[16]) & (g609) & (g644)) + ((g488) & (g552) & (!sk[16]) & (!g609) & (!g644)) + ((g488) & (g552) & (!sk[16]) & (!g609) & (g644)) + ((g488) & (g552) & (!sk[16]) & (g609) & (!g644)) + ((g488) & (g552) & (!sk[16]) & (g609) & (g644)) + ((g488) & (g552) & (sk[16]) & (!g609) & (g644)) + ((g488) & (g552) & (sk[16]) & (g609) & (!g644)));
	assign g2086 = (((!sk[17]) & (!ld) & (text_inx38x) & (!g1176)) + ((!sk[17]) & (!ld) & (text_inx38x) & (g1176)) + ((!sk[17]) & (ld) & (!text_inx38x) & (!g1176)) + ((!sk[17]) & (ld) & (!text_inx38x) & (g1176)) + ((!sk[17]) & (ld) & (text_inx38x) & (!g1176)) + ((!sk[17]) & (ld) & (text_inx38x) & (g1176)) + ((sk[17]) & (!ld) & (!text_inx38x) & (g1176)) + ((sk[17]) & (!ld) & (text_inx38x) & (g1176)) + ((sk[17]) & (ld) & (text_inx38x) & (!g1176)) + ((sk[17]) & (ld) & (text_inx38x) & (g1176)));
	assign g1177 = (((!sk[18]) & (!g438) & (g573) & (!g637)) + ((!sk[18]) & (!g438) & (g573) & (g637)) + ((!sk[18]) & (g438) & (!g573) & (!g637)) + ((!sk[18]) & (g438) & (!g573) & (g637)) + ((!sk[18]) & (g438) & (g573) & (!g637)) + ((!sk[18]) & (g438) & (g573) & (g637)) + ((sk[18]) & (!g438) & (!g573) & (g637)) + ((sk[18]) & (!g438) & (g573) & (!g637)) + ((sk[18]) & (g438) & (!g573) & (!g637)) + ((sk[18]) & (g438) & (g573) & (g637)));
	assign g1178 = (((!g446) & (!g509) & (!g630) & (!g1163) & (!g1176) & (g1177)) + ((!g446) & (!g509) & (!g630) & (!g1163) & (g1176) & (g1177)) + ((!g446) & (!g509) & (!g630) & (g1163) & (g1176) & (!g1177)) + ((!g446) & (!g509) & (!g630) & (g1163) & (g1176) & (g1177)) + ((!g446) & (!g509) & (g630) & (!g1163) & (!g1176) & (!g1177)) + ((!g446) & (!g509) & (g630) & (!g1163) & (g1176) & (!g1177)) + ((!g446) & (!g509) & (g630) & (g1163) & (g1176) & (!g1177)) + ((!g446) & (!g509) & (g630) & (g1163) & (g1176) & (g1177)) + ((!g446) & (g509) & (!g630) & (!g1163) & (!g1176) & (!g1177)) + ((!g446) & (g509) & (!g630) & (!g1163) & (g1176) & (!g1177)) + ((!g446) & (g509) & (!g630) & (g1163) & (g1176) & (!g1177)) + ((!g446) & (g509) & (!g630) & (g1163) & (g1176) & (g1177)) + ((!g446) & (g509) & (g630) & (!g1163) & (!g1176) & (g1177)) + ((!g446) & (g509) & (g630) & (!g1163) & (g1176) & (g1177)) + ((!g446) & (g509) & (g630) & (g1163) & (g1176) & (!g1177)) + ((!g446) & (g509) & (g630) & (g1163) & (g1176) & (g1177)) + ((g446) & (!g509) & (!g630) & (!g1163) & (!g1176) & (!g1177)) + ((g446) & (!g509) & (!g630) & (!g1163) & (g1176) & (!g1177)) + ((g446) & (!g509) & (!g630) & (g1163) & (!g1176) & (!g1177)) + ((g446) & (!g509) & (!g630) & (g1163) & (!g1176) & (g1177)) + ((g446) & (!g509) & (g630) & (!g1163) & (!g1176) & (g1177)) + ((g446) & (!g509) & (g630) & (!g1163) & (g1176) & (g1177)) + ((g446) & (!g509) & (g630) & (g1163) & (!g1176) & (!g1177)) + ((g446) & (!g509) & (g630) & (g1163) & (!g1176) & (g1177)) + ((g446) & (g509) & (!g630) & (!g1163) & (!g1176) & (g1177)) + ((g446) & (g509) & (!g630) & (!g1163) & (g1176) & (g1177)) + ((g446) & (g509) & (!g630) & (g1163) & (!g1176) & (!g1177)) + ((g446) & (g509) & (!g630) & (g1163) & (!g1176) & (g1177)) + ((g446) & (g509) & (g630) & (!g1163) & (!g1176) & (!g1177)) + ((g446) & (g509) & (g630) & (!g1163) & (g1176) & (!g1177)) + ((g446) & (g509) & (g630) & (g1163) & (!g1176) & (!g1177)) + ((g446) & (g509) & (g630) & (g1163) & (!g1176) & (g1177)));
	assign g2087 = (((!ld) & (!text_inx37x) & (sk[20]) & (g1179)) + ((!ld) & (text_inx37x) & (!sk[20]) & (!g1179)) + ((!ld) & (text_inx37x) & (!sk[20]) & (g1179)) + ((!ld) & (text_inx37x) & (sk[20]) & (g1179)) + ((ld) & (!text_inx37x) & (!sk[20]) & (!g1179)) + ((ld) & (!text_inx37x) & (!sk[20]) & (g1179)) + ((ld) & (text_inx37x) & (!sk[20]) & (!g1179)) + ((ld) & (text_inx37x) & (!sk[20]) & (g1179)) + ((ld) & (text_inx37x) & (sk[20]) & (!g1179)) + ((ld) & (text_inx37x) & (sk[20]) & (g1179)));
	assign g1180 = (((!g431) & (!sk[21]) & (g566) & (!g630)) + ((!g431) & (!sk[21]) & (g566) & (g630)) + ((!g431) & (sk[21]) & (!g566) & (g630)) + ((!g431) & (sk[21]) & (g566) & (!g630)) + ((g431) & (!sk[21]) & (!g566) & (!g630)) + ((g431) & (!sk[21]) & (!g566) & (g630)) + ((g431) & (!sk[21]) & (g566) & (!g630)) + ((g431) & (!sk[21]) & (g566) & (g630)) + ((g431) & (sk[21]) & (!g566) & (!g630)) + ((g431) & (sk[21]) & (g566) & (g630)));
	assign g1181 = (((!g439) & (!g502) & (!g623) & (!g1163) & (!g1179) & (g1180)) + ((!g439) & (!g502) & (!g623) & (!g1163) & (g1179) & (g1180)) + ((!g439) & (!g502) & (!g623) & (g1163) & (g1179) & (!g1180)) + ((!g439) & (!g502) & (!g623) & (g1163) & (g1179) & (g1180)) + ((!g439) & (!g502) & (g623) & (!g1163) & (!g1179) & (!g1180)) + ((!g439) & (!g502) & (g623) & (!g1163) & (g1179) & (!g1180)) + ((!g439) & (!g502) & (g623) & (g1163) & (g1179) & (!g1180)) + ((!g439) & (!g502) & (g623) & (g1163) & (g1179) & (g1180)) + ((!g439) & (g502) & (!g623) & (!g1163) & (!g1179) & (!g1180)) + ((!g439) & (g502) & (!g623) & (!g1163) & (g1179) & (!g1180)) + ((!g439) & (g502) & (!g623) & (g1163) & (g1179) & (!g1180)) + ((!g439) & (g502) & (!g623) & (g1163) & (g1179) & (g1180)) + ((!g439) & (g502) & (g623) & (!g1163) & (!g1179) & (g1180)) + ((!g439) & (g502) & (g623) & (!g1163) & (g1179) & (g1180)) + ((!g439) & (g502) & (g623) & (g1163) & (g1179) & (!g1180)) + ((!g439) & (g502) & (g623) & (g1163) & (g1179) & (g1180)) + ((g439) & (!g502) & (!g623) & (!g1163) & (!g1179) & (!g1180)) + ((g439) & (!g502) & (!g623) & (!g1163) & (g1179) & (!g1180)) + ((g439) & (!g502) & (!g623) & (g1163) & (!g1179) & (!g1180)) + ((g439) & (!g502) & (!g623) & (g1163) & (!g1179) & (g1180)) + ((g439) & (!g502) & (g623) & (!g1163) & (!g1179) & (g1180)) + ((g439) & (!g502) & (g623) & (!g1163) & (g1179) & (g1180)) + ((g439) & (!g502) & (g623) & (g1163) & (!g1179) & (!g1180)) + ((g439) & (!g502) & (g623) & (g1163) & (!g1179) & (g1180)) + ((g439) & (g502) & (!g623) & (!g1163) & (!g1179) & (g1180)) + ((g439) & (g502) & (!g623) & (!g1163) & (g1179) & (g1180)) + ((g439) & (g502) & (!g623) & (g1163) & (!g1179) & (!g1180)) + ((g439) & (g502) & (!g623) & (g1163) & (!g1179) & (g1180)) + ((g439) & (g502) & (g623) & (!g1163) & (!g1179) & (!g1180)) + ((g439) & (g502) & (g623) & (!g1163) & (g1179) & (!g1180)) + ((g439) & (g502) & (g623) & (g1163) & (!g1179) & (!g1180)) + ((g439) & (g502) & (g623) & (g1163) & (!g1179) & (g1180)));
	assign g2088 = (((!sk[23]) & (!ld) & (text_inx36x) & (!g1182)) + ((!sk[23]) & (!ld) & (text_inx36x) & (g1182)) + ((!sk[23]) & (ld) & (!text_inx36x) & (!g1182)) + ((!sk[23]) & (ld) & (!text_inx36x) & (g1182)) + ((!sk[23]) & (ld) & (text_inx36x) & (!g1182)) + ((!sk[23]) & (ld) & (text_inx36x) & (g1182)) + ((sk[23]) & (!ld) & (!text_inx36x) & (g1182)) + ((sk[23]) & (!ld) & (text_inx36x) & (g1182)) + ((sk[23]) & (ld) & (text_inx36x) & (!g1182)) + ((sk[23]) & (ld) & (text_inx36x) & (g1182)));
	assign g1183 = (((!g424) & (!sk[24]) & (g559) & (!g623)) + ((!g424) & (!sk[24]) & (g559) & (g623)) + ((!g424) & (sk[24]) & (!g559) & (g623)) + ((!g424) & (sk[24]) & (g559) & (!g623)) + ((g424) & (!sk[24]) & (!g559) & (!g623)) + ((g424) & (!sk[24]) & (!g559) & (g623)) + ((g424) & (!sk[24]) & (g559) & (!g623)) + ((g424) & (!sk[24]) & (g559) & (g623)) + ((g424) & (sk[24]) & (!g559) & (!g623)) + ((g424) & (sk[24]) & (g559) & (g623)));
	assign g1184 = (((!g432) & (!g452) & (!g495) & (!sk[25]) & (!g616) & (g644)) + ((!g432) & (!g452) & (!g495) & (!sk[25]) & (g616) & (g644)) + ((!g432) & (!g452) & (!g495) & (sk[25]) & (!g616) & (g644)) + ((!g432) & (!g452) & (!g495) & (sk[25]) & (g616) & (!g644)) + ((!g432) & (!g452) & (g495) & (!sk[25]) & (!g616) & (g644)) + ((!g432) & (!g452) & (g495) & (!sk[25]) & (g616) & (g644)) + ((!g432) & (!g452) & (g495) & (sk[25]) & (!g616) & (!g644)) + ((!g432) & (!g452) & (g495) & (sk[25]) & (g616) & (g644)) + ((!g432) & (g452) & (!g495) & (!sk[25]) & (!g616) & (!g644)) + ((!g432) & (g452) & (!g495) & (!sk[25]) & (!g616) & (g644)) + ((!g432) & (g452) & (!g495) & (!sk[25]) & (g616) & (!g644)) + ((!g432) & (g452) & (!g495) & (!sk[25]) & (g616) & (g644)) + ((!g432) & (g452) & (!g495) & (sk[25]) & (!g616) & (!g644)) + ((!g432) & (g452) & (!g495) & (sk[25]) & (g616) & (g644)) + ((!g432) & (g452) & (g495) & (!sk[25]) & (!g616) & (!g644)) + ((!g432) & (g452) & (g495) & (!sk[25]) & (!g616) & (g644)) + ((!g432) & (g452) & (g495) & (!sk[25]) & (g616) & (!g644)) + ((!g432) & (g452) & (g495) & (!sk[25]) & (g616) & (g644)) + ((!g432) & (g452) & (g495) & (sk[25]) & (!g616) & (g644)) + ((!g432) & (g452) & (g495) & (sk[25]) & (g616) & (!g644)) + ((g432) & (!g452) & (!g495) & (!sk[25]) & (!g616) & (g644)) + ((g432) & (!g452) & (!g495) & (!sk[25]) & (g616) & (!g644)) + ((g432) & (!g452) & (!g495) & (!sk[25]) & (g616) & (g644)) + ((g432) & (!g452) & (!g495) & (sk[25]) & (!g616) & (!g644)) + ((g432) & (!g452) & (!g495) & (sk[25]) & (g616) & (g644)) + ((g432) & (!g452) & (g495) & (!sk[25]) & (!g616) & (g644)) + ((g432) & (!g452) & (g495) & (!sk[25]) & (g616) & (!g644)) + ((g432) & (!g452) & (g495) & (!sk[25]) & (g616) & (g644)) + ((g432) & (!g452) & (g495) & (sk[25]) & (!g616) & (g644)) + ((g432) & (!g452) & (g495) & (sk[25]) & (g616) & (!g644)) + ((g432) & (g452) & (!g495) & (!sk[25]) & (!g616) & (!g644)) + ((g432) & (g452) & (!g495) & (!sk[25]) & (!g616) & (g644)) + ((g432) & (g452) & (!g495) & (!sk[25]) & (g616) & (!g644)) + ((g432) & (g452) & (!g495) & (!sk[25]) & (g616) & (g644)) + ((g432) & (g452) & (!g495) & (sk[25]) & (!g616) & (g644)) + ((g432) & (g452) & (!g495) & (sk[25]) & (g616) & (!g644)) + ((g432) & (g452) & (g495) & (!sk[25]) & (!g616) & (!g644)) + ((g432) & (g452) & (g495) & (!sk[25]) & (!g616) & (g644)) + ((g432) & (g452) & (g495) & (!sk[25]) & (g616) & (!g644)) + ((g432) & (g452) & (g495) & (!sk[25]) & (g616) & (g644)) + ((g432) & (g452) & (g495) & (sk[25]) & (!g616) & (!g644)) + ((g432) & (g452) & (g495) & (sk[25]) & (g616) & (g644)));
	assign g1185 = (((!g432) & (!g1163) & (!sk[26]) & (!g1182) & (!g1183) & (g1184)) + ((!g432) & (!g1163) & (!sk[26]) & (!g1182) & (g1183) & (g1184)) + ((!g432) & (!g1163) & (!sk[26]) & (g1182) & (!g1183) & (g1184)) + ((!g432) & (!g1163) & (!sk[26]) & (g1182) & (g1183) & (g1184)) + ((!g432) & (!g1163) & (sk[26]) & (!g1182) & (!g1183) & (g1184)) + ((!g432) & (!g1163) & (sk[26]) & (!g1182) & (g1183) & (!g1184)) + ((!g432) & (!g1163) & (sk[26]) & (g1182) & (!g1183) & (g1184)) + ((!g432) & (!g1163) & (sk[26]) & (g1182) & (g1183) & (!g1184)) + ((!g432) & (g1163) & (!sk[26]) & (!g1182) & (!g1183) & (!g1184)) + ((!g432) & (g1163) & (!sk[26]) & (!g1182) & (!g1183) & (g1184)) + ((!g432) & (g1163) & (!sk[26]) & (!g1182) & (g1183) & (!g1184)) + ((!g432) & (g1163) & (!sk[26]) & (!g1182) & (g1183) & (g1184)) + ((!g432) & (g1163) & (!sk[26]) & (g1182) & (!g1183) & (!g1184)) + ((!g432) & (g1163) & (!sk[26]) & (g1182) & (!g1183) & (g1184)) + ((!g432) & (g1163) & (!sk[26]) & (g1182) & (g1183) & (!g1184)) + ((!g432) & (g1163) & (!sk[26]) & (g1182) & (g1183) & (g1184)) + ((!g432) & (g1163) & (sk[26]) & (g1182) & (!g1183) & (!g1184)) + ((!g432) & (g1163) & (sk[26]) & (g1182) & (!g1183) & (g1184)) + ((!g432) & (g1163) & (sk[26]) & (g1182) & (g1183) & (!g1184)) + ((!g432) & (g1163) & (sk[26]) & (g1182) & (g1183) & (g1184)) + ((g432) & (!g1163) & (!sk[26]) & (!g1182) & (!g1183) & (g1184)) + ((g432) & (!g1163) & (!sk[26]) & (!g1182) & (g1183) & (!g1184)) + ((g432) & (!g1163) & (!sk[26]) & (!g1182) & (g1183) & (g1184)) + ((g432) & (!g1163) & (!sk[26]) & (g1182) & (!g1183) & (g1184)) + ((g432) & (!g1163) & (!sk[26]) & (g1182) & (g1183) & (!g1184)) + ((g432) & (!g1163) & (!sk[26]) & (g1182) & (g1183) & (g1184)) + ((g432) & (!g1163) & (sk[26]) & (!g1182) & (!g1183) & (g1184)) + ((g432) & (!g1163) & (sk[26]) & (!g1182) & (g1183) & (!g1184)) + ((g432) & (!g1163) & (sk[26]) & (g1182) & (!g1183) & (g1184)) + ((g432) & (!g1163) & (sk[26]) & (g1182) & (g1183) & (!g1184)) + ((g432) & (g1163) & (!sk[26]) & (!g1182) & (!g1183) & (!g1184)) + ((g432) & (g1163) & (!sk[26]) & (!g1182) & (!g1183) & (g1184)) + ((g432) & (g1163) & (!sk[26]) & (!g1182) & (g1183) & (!g1184)) + ((g432) & (g1163) & (!sk[26]) & (!g1182) & (g1183) & (g1184)) + ((g432) & (g1163) & (!sk[26]) & (g1182) & (!g1183) & (!g1184)) + ((g432) & (g1163) & (!sk[26]) & (g1182) & (!g1183) & (g1184)) + ((g432) & (g1163) & (!sk[26]) & (g1182) & (g1183) & (!g1184)) + ((g432) & (g1163) & (!sk[26]) & (g1182) & (g1183) & (g1184)) + ((g432) & (g1163) & (sk[26]) & (!g1182) & (!g1183) & (!g1184)) + ((g432) & (g1163) & (sk[26]) & (!g1182) & (!g1183) & (g1184)) + ((g432) & (g1163) & (sk[26]) & (!g1182) & (g1183) & (!g1184)) + ((g432) & (g1163) & (sk[26]) & (!g1182) & (g1183) & (g1184)));
	assign g2089 = (((!ld) & (!text_inx39x) & (sk[27]) & (g1186)) + ((!ld) & (text_inx39x) & (!sk[27]) & (!g1186)) + ((!ld) & (text_inx39x) & (!sk[27]) & (g1186)) + ((!ld) & (text_inx39x) & (sk[27]) & (g1186)) + ((ld) & (!text_inx39x) & (!sk[27]) & (g1186)) + ((ld) & (text_inx39x) & (!sk[27]) & (!g1186)) + ((ld) & (text_inx39x) & (!sk[27]) & (g1186)) + ((ld) & (text_inx39x) & (sk[27]) & (!g1186)) + ((ld) & (text_inx39x) & (sk[27]) & (g1186)));
	assign g1187 = (((!sk[28]) & (!g445) & (g580) & (!g644)) + ((!sk[28]) & (!g445) & (g580) & (g644)) + ((!sk[28]) & (g445) & (!g580) & (g644)) + ((!sk[28]) & (g445) & (g580) & (!g644)) + ((!sk[28]) & (g445) & (g580) & (g644)) + ((sk[28]) & (!g445) & (!g580) & (g644)) + ((sk[28]) & (!g445) & (g580) & (!g644)) + ((sk[28]) & (g445) & (!g580) & (!g644)) + ((sk[28]) & (g445) & (g580) & (g644)));
	assign g1188 = (((!g453) & (!g516) & (!g637) & (!g1163) & (!g1186) & (g1187)) + ((!g453) & (!g516) & (!g637) & (!g1163) & (g1186) & (g1187)) + ((!g453) & (!g516) & (!g637) & (g1163) & (g1186) & (!g1187)) + ((!g453) & (!g516) & (!g637) & (g1163) & (g1186) & (g1187)) + ((!g453) & (!g516) & (g637) & (!g1163) & (!g1186) & (!g1187)) + ((!g453) & (!g516) & (g637) & (!g1163) & (g1186) & (!g1187)) + ((!g453) & (!g516) & (g637) & (g1163) & (g1186) & (!g1187)) + ((!g453) & (!g516) & (g637) & (g1163) & (g1186) & (g1187)) + ((!g453) & (g516) & (!g637) & (!g1163) & (!g1186) & (!g1187)) + ((!g453) & (g516) & (!g637) & (!g1163) & (g1186) & (!g1187)) + ((!g453) & (g516) & (!g637) & (g1163) & (g1186) & (!g1187)) + ((!g453) & (g516) & (!g637) & (g1163) & (g1186) & (g1187)) + ((!g453) & (g516) & (g637) & (!g1163) & (!g1186) & (g1187)) + ((!g453) & (g516) & (g637) & (!g1163) & (g1186) & (g1187)) + ((!g453) & (g516) & (g637) & (g1163) & (g1186) & (!g1187)) + ((!g453) & (g516) & (g637) & (g1163) & (g1186) & (g1187)) + ((g453) & (!g516) & (!g637) & (!g1163) & (!g1186) & (!g1187)) + ((g453) & (!g516) & (!g637) & (!g1163) & (g1186) & (!g1187)) + ((g453) & (!g516) & (!g637) & (g1163) & (!g1186) & (!g1187)) + ((g453) & (!g516) & (!g637) & (g1163) & (!g1186) & (g1187)) + ((g453) & (!g516) & (g637) & (!g1163) & (!g1186) & (g1187)) + ((g453) & (!g516) & (g637) & (!g1163) & (g1186) & (g1187)) + ((g453) & (!g516) & (g637) & (g1163) & (!g1186) & (!g1187)) + ((g453) & (!g516) & (g637) & (g1163) & (!g1186) & (g1187)) + ((g453) & (g516) & (!g637) & (!g1163) & (!g1186) & (g1187)) + ((g453) & (g516) & (!g637) & (!g1163) & (g1186) & (g1187)) + ((g453) & (g516) & (!g637) & (g1163) & (!g1186) & (!g1187)) + ((g453) & (g516) & (!g637) & (g1163) & (!g1186) & (g1187)) + ((g453) & (g516) & (g637) & (!g1163) & (!g1186) & (!g1187)) + ((g453) & (g516) & (g637) & (!g1163) & (g1186) & (!g1187)) + ((g453) & (g516) & (g637) & (g1163) & (!g1186) & (!g1187)) + ((g453) & (g516) & (g637) & (g1163) & (!g1186) & (g1187)));
	assign g1189 = (((!g340) & (!g347) & (!g354) & (!g361) & (g382) & (g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g382) & (!g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g382) & (g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (g382) & (!g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (!g382) & (!g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (!g382) & (g375)) + ((!g340) & (!g347) & (g354) & (g361) & (!g382) & (!g375)) + ((!g340) & (!g347) & (g354) & (g361) & (g382) & (g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (g382) & (!g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (g382) & (g375)) + ((!g340) & (g347) & (!g354) & (g361) & (g382) & (!g375)) + ((!g340) & (g347) & (!g354) & (g361) & (g382) & (g375)) + ((!g340) & (g347) & (g354) & (!g361) & (g382) & (!g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (!g382) & (!g375)) + ((g340) & (!g347) & (g354) & (!g361) & (g382) & (!g375)) + ((g340) & (!g347) & (g354) & (g361) & (!g382) & (g375)) + ((g340) & (!g347) & (g354) & (g361) & (g382) & (g375)) + ((g340) & (g347) & (!g354) & (!g361) & (!g382) & (g375)) + ((g340) & (g347) & (!g354) & (!g361) & (g382) & (!g375)) + ((g340) & (g347) & (g354) & (!g361) & (!g382) & (g375)) + ((g340) & (g347) & (g354) & (!g361) & (g382) & (!g375)) + ((g340) & (g347) & (g354) & (g361) & (!g382) & (!g375)) + ((g340) & (g347) & (g354) & (g361) & (g382) & (!g375)) + ((g340) & (g347) & (g354) & (g361) & (g382) & (g375)));
	assign g1190 = (((!g340) & (!g347) & (!g354) & (!g361) & (g382) & (!g375)) + ((!g340) & (!g347) & (!g354) & (!g361) & (g382) & (g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g382) & (!g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g382) & (g375)) + ((!g340) & (!g347) & (g354) & (g361) & (!g382) & (g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (!g382) & (!g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (!g382) & (g375)) + ((!g340) & (g347) & (g354) & (!g361) & (!g382) & (!g375)) + ((!g340) & (g347) & (g354) & (!g361) & (!g382) & (g375)) + ((!g340) & (g347) & (g354) & (!g361) & (g382) & (!g375)) + ((!g340) & (g347) & (g354) & (g361) & (g382) & (g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (!g382) & (g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (g382) & (!g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (g382) & (g375)) + ((g340) & (!g347) & (!g354) & (g361) & (g382) & (!g375)) + ((g340) & (!g347) & (g354) & (!g361) & (!g382) & (!g375)) + ((g340) & (!g347) & (g354) & (!g361) & (g382) & (g375)) + ((g340) & (!g347) & (g354) & (g361) & (!g382) & (g375)) + ((g340) & (!g347) & (g354) & (g361) & (g382) & (g375)) + ((g340) & (g347) & (!g354) & (!g361) & (!g382) & (!g375)) + ((g340) & (g347) & (!g354) & (!g361) & (!g382) & (g375)) + ((g340) & (g347) & (!g354) & (!g361) & (g382) & (!g375)) + ((g340) & (g347) & (!g354) & (!g361) & (g382) & (g375)) + ((g340) & (g347) & (!g354) & (g361) & (!g382) & (!g375)) + ((g340) & (g347) & (!g354) & (g361) & (g382) & (!g375)) + ((g340) & (g347) & (!g354) & (g361) & (g382) & (g375)) + ((g340) & (g347) & (g354) & (!g361) & (g382) & (!g375)) + ((g340) & (g347) & (g354) & (!g361) & (g382) & (g375)) + ((g340) & (g347) & (g354) & (g361) & (!g382) & (g375)) + ((g340) & (g347) & (g354) & (g361) & (g382) & (!g375)));
	assign g1191 = (((!g340) & (!g347) & (!g354) & (!g361) & (!g382) & (!g375)) + ((!g340) & (!g347) & (!g354) & (!g361) & (g382) & (g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (g382) & (g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (!g382) & (!g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (!g382) & (g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (g382) & (g375)) + ((!g340) & (!g347) & (g354) & (g361) & (!g382) & (g375)) + ((!g340) & (!g347) & (g354) & (g361) & (g382) & (!g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (!g382) & (!g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (g382) & (!g375)) + ((!g340) & (g347) & (!g354) & (g361) & (g382) & (g375)) + ((!g340) & (g347) & (g354) & (g361) & (!g382) & (!g375)) + ((!g340) & (g347) & (g354) & (g361) & (g382) & (!g375)) + ((g340) & (!g347) & (!g354) & (g361) & (!g382) & (!g375)) + ((g340) & (!g347) & (!g354) & (g361) & (!g382) & (g375)) + ((g340) & (!g347) & (!g354) & (g361) & (g382) & (!g375)) + ((g340) & (!g347) & (g354) & (!g361) & (!g382) & (!g375)) + ((g340) & (!g347) & (g354) & (!g361) & (g382) & (g375)) + ((g340) & (!g347) & (g354) & (g361) & (!g382) & (!g375)) + ((g340) & (!g347) & (g354) & (g361) & (!g382) & (g375)) + ((g340) & (!g347) & (g354) & (g361) & (g382) & (!g375)) + ((g340) & (!g347) & (g354) & (g361) & (g382) & (g375)) + ((g340) & (g347) & (!g354) & (!g361) & (g382) & (g375)) + ((g340) & (g347) & (!g354) & (g361) & (!g382) & (!g375)) + ((g340) & (g347) & (!g354) & (g361) & (g382) & (!g375)) + ((g340) & (g347) & (!g354) & (g361) & (g382) & (g375)) + ((g340) & (g347) & (g354) & (!g361) & (!g382) & (!g375)) + ((g340) & (g347) & (g354) & (g361) & (!g382) & (!g375)) + ((g340) & (g347) & (g354) & (g361) & (!g382) & (g375)) + ((g340) & (g347) & (g354) & (g361) & (g382) & (g375)));
	assign g1192 = (((!g340) & (!g347) & (!g354) & (!g361) & (!g382) & (g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (g382) & (!g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (g382) & (g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (!g382) & (g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (g382) & (g375)) + ((!g340) & (!g347) & (g354) & (g361) & (!g382) & (g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (!g382) & (!g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (!g382) & (g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (g382) & (!g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (g382) & (g375)) + ((!g340) & (g347) & (!g354) & (g361) & (g382) & (!g375)) + ((!g340) & (g347) & (!g354) & (g361) & (g382) & (g375)) + ((!g340) & (g347) & (g354) & (g361) & (!g382) & (!g375)) + ((!g340) & (g347) & (g354) & (g361) & (g382) & (!g375)) + ((!g340) & (g347) & (g354) & (g361) & (g382) & (g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (!g382) & (!g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (g382) & (g375)) + ((g340) & (!g347) & (!g354) & (g361) & (g382) & (!g375)) + ((g340) & (!g347) & (!g354) & (g361) & (g382) & (g375)) + ((g340) & (!g347) & (g354) & (!g361) & (!g382) & (g375)) + ((g340) & (!g347) & (g354) & (!g361) & (g382) & (!g375)) + ((g340) & (!g347) & (g354) & (g361) & (g382) & (!g375)) + ((g340) & (g347) & (!g354) & (!g361) & (!g382) & (g375)) + ((g340) & (g347) & (!g354) & (!g361) & (g382) & (g375)) + ((g340) & (g347) & (!g354) & (g361) & (g382) & (!g375)) + ((g340) & (g347) & (!g354) & (g361) & (g382) & (g375)) + ((g340) & (g347) & (g354) & (!g361) & (!g382) & (g375)) + ((g340) & (g347) & (g354) & (g361) & (!g382) & (!g375)));
	assign g1193 = (((!g1189) & (!g1190) & (!g1191) & (!g1192) & (!g368) & (!g389)) + ((!g1189) & (!g1190) & (!g1191) & (g1192) & (!g368) & (!g389)) + ((!g1189) & (!g1190) & (!g1191) & (g1192) & (g368) & (g389)) + ((!g1189) & (!g1190) & (g1191) & (!g1192) & (!g368) & (!g389)) + ((!g1189) & (!g1190) & (g1191) & (!g1192) & (!g368) & (g389)) + ((!g1189) & (!g1190) & (g1191) & (g1192) & (!g368) & (!g389)) + ((!g1189) & (!g1190) & (g1191) & (g1192) & (!g368) & (g389)) + ((!g1189) & (!g1190) & (g1191) & (g1192) & (g368) & (g389)) + ((!g1189) & (g1190) & (!g1191) & (!g1192) & (!g368) & (!g389)) + ((!g1189) & (g1190) & (!g1191) & (!g1192) & (g368) & (!g389)) + ((!g1189) & (g1190) & (!g1191) & (g1192) & (!g368) & (!g389)) + ((!g1189) & (g1190) & (!g1191) & (g1192) & (g368) & (!g389)) + ((!g1189) & (g1190) & (!g1191) & (g1192) & (g368) & (g389)) + ((!g1189) & (g1190) & (g1191) & (!g1192) & (!g368) & (!g389)) + ((!g1189) & (g1190) & (g1191) & (!g1192) & (!g368) & (g389)) + ((!g1189) & (g1190) & (g1191) & (!g1192) & (g368) & (!g389)) + ((!g1189) & (g1190) & (g1191) & (g1192) & (!g368) & (!g389)) + ((!g1189) & (g1190) & (g1191) & (g1192) & (!g368) & (g389)) + ((!g1189) & (g1190) & (g1191) & (g1192) & (g368) & (!g389)) + ((!g1189) & (g1190) & (g1191) & (g1192) & (g368) & (g389)) + ((g1189) & (!g1190) & (!g1191) & (g1192) & (g368) & (g389)) + ((g1189) & (!g1190) & (g1191) & (!g1192) & (!g368) & (g389)) + ((g1189) & (!g1190) & (g1191) & (g1192) & (!g368) & (g389)) + ((g1189) & (!g1190) & (g1191) & (g1192) & (g368) & (g389)) + ((g1189) & (g1190) & (!g1191) & (!g1192) & (g368) & (!g389)) + ((g1189) & (g1190) & (!g1191) & (g1192) & (g368) & (!g389)) + ((g1189) & (g1190) & (!g1191) & (g1192) & (g368) & (g389)) + ((g1189) & (g1190) & (g1191) & (!g1192) & (!g368) & (g389)) + ((g1189) & (g1190) & (g1191) & (!g1192) & (g368) & (!g389)) + ((g1189) & (g1190) & (g1191) & (g1192) & (!g368) & (g389)) + ((g1189) & (g1190) & (g1191) & (g1192) & (g368) & (!g389)) + ((g1189) & (g1190) & (g1191) & (g1192) & (g368) & (g389)));
	assign g1194 = (((!g404) & (!g660) & (!g916) & (sk[35]) & (g1193)) + ((!g404) & (!g660) & (g916) & (!sk[35]) & (!g1193)) + ((!g404) & (!g660) & (g916) & (!sk[35]) & (g1193)) + ((!g404) & (!g660) & (g916) & (sk[35]) & (!g1193)) + ((!g404) & (g660) & (!g916) & (!sk[35]) & (!g1193)) + ((!g404) & (g660) & (!g916) & (!sk[35]) & (g1193)) + ((!g404) & (g660) & (!g916) & (sk[35]) & (!g1193)) + ((!g404) & (g660) & (g916) & (!sk[35]) & (!g1193)) + ((!g404) & (g660) & (g916) & (!sk[35]) & (g1193)) + ((!g404) & (g660) & (g916) & (sk[35]) & (g1193)) + ((g404) & (!g660) & (!g916) & (sk[35]) & (!g1193)) + ((g404) & (!g660) & (g916) & (!sk[35]) & (!g1193)) + ((g404) & (!g660) & (g916) & (!sk[35]) & (g1193)) + ((g404) & (!g660) & (g916) & (sk[35]) & (g1193)) + ((g404) & (g660) & (!g916) & (!sk[35]) & (!g1193)) + ((g404) & (g660) & (!g916) & (!sk[35]) & (g1193)) + ((g404) & (g660) & (!g916) & (sk[35]) & (g1193)) + ((g404) & (g660) & (g916) & (!sk[35]) & (!g1193)) + ((g404) & (g660) & (g916) & (!sk[35]) & (g1193)) + ((g404) & (g660) & (g916) & (sk[35]) & (!g1193)));
	assign g1195 = (((!ld) & (!g148) & (g1194) & (!sk[36]) & (!keyx0x)) + ((!ld) & (!g148) & (g1194) & (!sk[36]) & (keyx0x)) + ((!ld) & (!g148) & (g1194) & (sk[36]) & (!keyx0x)) + ((!ld) & (!g148) & (g1194) & (sk[36]) & (keyx0x)) + ((!ld) & (g148) & (!g1194) & (!sk[36]) & (!keyx0x)) + ((!ld) & (g148) & (!g1194) & (!sk[36]) & (keyx0x)) + ((!ld) & (g148) & (!g1194) & (sk[36]) & (!keyx0x)) + ((!ld) & (g148) & (!g1194) & (sk[36]) & (keyx0x)) + ((!ld) & (g148) & (g1194) & (!sk[36]) & (!keyx0x)) + ((!ld) & (g148) & (g1194) & (!sk[36]) & (keyx0x)) + ((ld) & (!g148) & (!g1194) & (sk[36]) & (keyx0x)) + ((ld) & (!g148) & (g1194) & (!sk[36]) & (!keyx0x)) + ((ld) & (!g148) & (g1194) & (!sk[36]) & (keyx0x)) + ((ld) & (!g148) & (g1194) & (sk[36]) & (keyx0x)) + ((ld) & (g148) & (!g1194) & (!sk[36]) & (!keyx0x)) + ((ld) & (g148) & (!g1194) & (!sk[36]) & (keyx0x)) + ((ld) & (g148) & (!g1194) & (sk[36]) & (keyx0x)) + ((ld) & (g148) & (g1194) & (!sk[36]) & (!keyx0x)) + ((ld) & (g148) & (g1194) & (!sk[36]) & (keyx0x)) + ((ld) & (g148) & (g1194) & (sk[36]) & (keyx0x)));
	assign g1196 = (((!g340) & (!g347) & (!g354) & (!g361) & (!g368) & (g382)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g368) & (!g382)) + ((!g340) & (!g347) & (!g354) & (g361) & (g368) & (!g382)) + ((!g340) & (!g347) & (g354) & (!g361) & (g368) & (g382)) + ((!g340) & (!g347) & (g354) & (g361) & (!g368) & (g382)) + ((!g340) & (!g347) & (g354) & (g361) & (g368) & (!g382)) + ((!g340) & (g347) & (!g354) & (!g361) & (!g368) & (g382)) + ((!g340) & (g347) & (!g354) & (!g361) & (g368) & (!g382)) + ((!g340) & (g347) & (!g354) & (!g361) & (g368) & (g382)) + ((!g340) & (g347) & (g354) & (!g361) & (g368) & (g382)) + ((!g340) & (g347) & (g354) & (g361) & (g368) & (g382)) + ((g340) & (!g347) & (!g354) & (!g361) & (!g368) & (!g382)) + ((g340) & (!g347) & (!g354) & (!g361) & (g368) & (g382)) + ((g340) & (!g347) & (!g354) & (g361) & (!g368) & (!g382)) + ((g340) & (!g347) & (!g354) & (g361) & (g368) & (!g382)) + ((g340) & (!g347) & (g354) & (!g361) & (g368) & (!g382)) + ((g340) & (!g347) & (g354) & (!g361) & (g368) & (g382)) + ((g340) & (!g347) & (g354) & (g361) & (g368) & (!g382)) + ((g340) & (!g347) & (g354) & (g361) & (g368) & (g382)) + ((g340) & (g347) & (!g354) & (!g361) & (g368) & (!g382)) + ((g340) & (g347) & (!g354) & (!g361) & (g368) & (g382)) + ((g340) & (g347) & (!g354) & (g361) & (g368) & (g382)) + ((g340) & (g347) & (g354) & (!g361) & (!g368) & (!g382)) + ((g340) & (g347) & (g354) & (!g361) & (!g368) & (g382)) + ((g340) & (g347) & (g354) & (!g361) & (g368) & (!g382)) + ((g340) & (g347) & (g354) & (g361) & (!g368) & (g382)) + ((g340) & (g347) & (g354) & (g361) & (g368) & (!g382)));
	assign g1197 = (((!g340) & (!g347) & (!g354) & (!g361) & (!g368) & (g382)) + ((!g340) & (!g347) & (!g354) & (!g361) & (g368) & (!g382)) + ((!g340) & (!g347) & (!g354) & (!g361) & (g368) & (g382)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g368) & (!g382)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g368) & (g382)) + ((!g340) & (!g347) & (!g354) & (g361) & (g368) & (g382)) + ((!g340) & (!g347) & (g354) & (!g361) & (g368) & (!g382)) + ((!g340) & (!g347) & (g354) & (g361) & (!g368) & (!g382)) + ((!g340) & (!g347) & (g354) & (g361) & (!g368) & (g382)) + ((!g340) & (!g347) & (g354) & (g361) & (g368) & (g382)) + ((!g340) & (g347) & (!g354) & (!g361) & (g368) & (g382)) + ((!g340) & (g347) & (!g354) & (g361) & (!g368) & (!g382)) + ((!g340) & (g347) & (!g354) & (g361) & (g368) & (!g382)) + ((!g340) & (g347) & (g354) & (!g361) & (g368) & (!g382)) + ((!g340) & (g347) & (g354) & (!g361) & (g368) & (g382)) + ((!g340) & (g347) & (g354) & (g361) & (!g368) & (!g382)) + ((g340) & (!g347) & (!g354) & (!g361) & (!g368) & (!g382)) + ((g340) & (!g347) & (!g354) & (g361) & (!g368) & (!g382)) + ((g340) & (!g347) & (!g354) & (g361) & (!g368) & (g382)) + ((g340) & (!g347) & (g354) & (!g361) & (!g368) & (g382)) + ((g340) & (!g347) & (g354) & (!g361) & (g368) & (g382)) + ((g340) & (!g347) & (g354) & (g361) & (!g368) & (!g382)) + ((g340) & (!g347) & (g354) & (g361) & (!g368) & (g382)) + ((g340) & (g347) & (!g354) & (g361) & (!g368) & (!g382)) + ((g340) & (g347) & (!g354) & (g361) & (g368) & (g382)) + ((g340) & (g347) & (g354) & (!g361) & (!g368) & (!g382)) + ((g340) & (g347) & (g354) & (!g361) & (!g368) & (g382)) + ((g340) & (g347) & (g354) & (!g361) & (g368) & (g382)) + ((g340) & (g347) & (g354) & (g361) & (!g368) & (!g382)) + ((g340) & (g347) & (g354) & (g361) & (!g368) & (g382)) + ((g340) & (g347) & (g354) & (g361) & (g368) & (!g382)));
	assign g1198 = (((!g340) & (!g347) & (!g354) & (!g361) & (!g368) & (g382)) + ((!g340) & (!g347) & (!g354) & (g361) & (g368) & (!g382)) + ((!g340) & (!g347) & (g354) & (!g361) & (!g368) & (!g382)) + ((!g340) & (!g347) & (g354) & (!g361) & (g368) & (!g382)) + ((!g340) & (!g347) & (g354) & (g361) & (!g368) & (g382)) + ((!g340) & (!g347) & (g354) & (g361) & (g368) & (!g382)) + ((!g340) & (!g347) & (g354) & (g361) & (g368) & (g382)) + ((!g340) & (g347) & (!g354) & (!g361) & (!g368) & (!g382)) + ((!g340) & (g347) & (!g354) & (!g361) & (g368) & (!g382)) + ((!g340) & (g347) & (!g354) & (g361) & (!g368) & (!g382)) + ((!g340) & (g347) & (!g354) & (g361) & (g368) & (g382)) + ((!g340) & (g347) & (g354) & (!g361) & (g368) & (g382)) + ((!g340) & (g347) & (g354) & (g361) & (!g368) & (g382)) + ((!g340) & (g347) & (g354) & (g361) & (g368) & (!g382)) + ((g340) & (!g347) & (!g354) & (!g361) & (g368) & (g382)) + ((g340) & (!g347) & (!g354) & (g361) & (!g368) & (!g382)) + ((g340) & (!g347) & (!g354) & (g361) & (g368) & (!g382)) + ((g340) & (!g347) & (g354) & (!g361) & (!g368) & (!g382)) + ((g340) & (!g347) & (g354) & (!g361) & (!g368) & (g382)) + ((g340) & (!g347) & (g354) & (!g361) & (g368) & (!g382)) + ((g340) & (!g347) & (g354) & (!g361) & (g368) & (g382)) + ((g340) & (!g347) & (g354) & (g361) & (g368) & (!g382)) + ((g340) & (g347) & (!g354) & (!g361) & (!g368) & (g382)) + ((g340) & (g347) & (!g354) & (!g361) & (g368) & (g382)) + ((g340) & (g347) & (!g354) & (g361) & (!g368) & (g382)) + ((g340) & (g347) & (g354) & (!g361) & (!g368) & (!g382)) + ((g340) & (g347) & (g354) & (!g361) & (!g368) & (g382)) + ((g340) & (g347) & (g354) & (!g361) & (g368) & (g382)) + ((g340) & (g347) & (g354) & (g361) & (!g368) & (!g382)) + ((g340) & (g347) & (g354) & (g361) & (!g368) & (g382)) + ((g340) & (g347) & (g354) & (g361) & (g368) & (!g382)) + ((g340) & (g347) & (g354) & (g361) & (g368) & (g382)));
	assign g1199 = (((!g340) & (!g347) & (!g354) & (!g361) & (g368) & (!g382)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g368) & (!g382)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g368) & (g382)) + ((!g340) & (!g347) & (g354) & (!g361) & (g368) & (g382)) + ((!g340) & (!g347) & (g354) & (g361) & (!g368) & (g382)) + ((!g340) & (g347) & (!g354) & (!g361) & (!g368) & (!g382)) + ((!g340) & (g347) & (!g354) & (!g361) & (g368) & (!g382)) + ((!g340) & (g347) & (!g354) & (g361) & (!g368) & (g382)) + ((!g340) & (g347) & (g354) & (!g361) & (!g368) & (g382)) + ((!g340) & (g347) & (g354) & (!g361) & (g368) & (!g382)) + ((!g340) & (g347) & (g354) & (!g361) & (g368) & (g382)) + ((!g340) & (g347) & (g354) & (g361) & (g368) & (!g382)) + ((!g340) & (g347) & (g354) & (g361) & (g368) & (g382)) + ((g340) & (!g347) & (!g354) & (!g361) & (!g368) & (!g382)) + ((g340) & (!g347) & (!g354) & (g361) & (!g368) & (!g382)) + ((g340) & (!g347) & (!g354) & (g361) & (!g368) & (g382)) + ((g340) & (!g347) & (!g354) & (g361) & (g368) & (!g382)) + ((g340) & (!g347) & (g354) & (!g361) & (!g368) & (!g382)) + ((g340) & (!g347) & (g354) & (!g361) & (g368) & (g382)) + ((g340) & (!g347) & (g354) & (g361) & (g368) & (!g382)) + ((g340) & (g347) & (!g354) & (!g361) & (!g368) & (!g382)) + ((g340) & (g347) & (!g354) & (g361) & (!g368) & (!g382)) + ((g340) & (g347) & (!g354) & (g361) & (g368) & (!g382)) + ((g340) & (g347) & (!g354) & (g361) & (g368) & (g382)) + ((g340) & (g347) & (g354) & (g361) & (!g368) & (g382)) + ((g340) & (g347) & (g354) & (g361) & (g368) & (g382)));
	assign g1200 = (((!g1196) & (!g1197) & (!g1198) & (!g1199) & (!g375) & (!g389)) + ((!g1196) & (!g1197) & (!g1198) & (!g1199) & (g375) & (!g389)) + ((!g1196) & (!g1197) & (!g1198) & (g1199) & (!g375) & (!g389)) + ((!g1196) & (!g1197) & (!g1198) & (g1199) & (g375) & (!g389)) + ((!g1196) & (!g1197) & (!g1198) & (g1199) & (g375) & (g389)) + ((!g1196) & (!g1197) & (g1198) & (!g1199) & (!g375) & (!g389)) + ((!g1196) & (!g1197) & (g1198) & (!g1199) & (!g375) & (g389)) + ((!g1196) & (!g1197) & (g1198) & (!g1199) & (g375) & (!g389)) + ((!g1196) & (!g1197) & (g1198) & (g1199) & (!g375) & (!g389)) + ((!g1196) & (!g1197) & (g1198) & (g1199) & (!g375) & (g389)) + ((!g1196) & (!g1197) & (g1198) & (g1199) & (g375) & (!g389)) + ((!g1196) & (!g1197) & (g1198) & (g1199) & (g375) & (g389)) + ((!g1196) & (g1197) & (!g1198) & (!g1199) & (!g375) & (!g389)) + ((!g1196) & (g1197) & (!g1198) & (g1199) & (!g375) & (!g389)) + ((!g1196) & (g1197) & (!g1198) & (g1199) & (g375) & (g389)) + ((!g1196) & (g1197) & (g1198) & (!g1199) & (!g375) & (!g389)) + ((!g1196) & (g1197) & (g1198) & (!g1199) & (!g375) & (g389)) + ((!g1196) & (g1197) & (g1198) & (g1199) & (!g375) & (!g389)) + ((!g1196) & (g1197) & (g1198) & (g1199) & (!g375) & (g389)) + ((!g1196) & (g1197) & (g1198) & (g1199) & (g375) & (g389)) + ((g1196) & (!g1197) & (!g1198) & (!g1199) & (g375) & (!g389)) + ((g1196) & (!g1197) & (!g1198) & (g1199) & (g375) & (!g389)) + ((g1196) & (!g1197) & (!g1198) & (g1199) & (g375) & (g389)) + ((g1196) & (!g1197) & (g1198) & (!g1199) & (!g375) & (g389)) + ((g1196) & (!g1197) & (g1198) & (!g1199) & (g375) & (!g389)) + ((g1196) & (!g1197) & (g1198) & (g1199) & (!g375) & (g389)) + ((g1196) & (!g1197) & (g1198) & (g1199) & (g375) & (!g389)) + ((g1196) & (!g1197) & (g1198) & (g1199) & (g375) & (g389)) + ((g1196) & (g1197) & (!g1198) & (g1199) & (g375) & (g389)) + ((g1196) & (g1197) & (g1198) & (!g1199) & (!g375) & (g389)) + ((g1196) & (g1197) & (g1198) & (g1199) & (!g375) & (g389)) + ((g1196) & (g1197) & (g1198) & (g1199) & (g375) & (g389)));
	assign g1201 = (((!g411) & (!g667) & (!sk[42]) & (g923) & (!g1200)) + ((!g411) & (!g667) & (!sk[42]) & (g923) & (g1200)) + ((!g411) & (!g667) & (sk[42]) & (!g923) & (g1200)) + ((!g411) & (!g667) & (sk[42]) & (g923) & (!g1200)) + ((!g411) & (g667) & (!sk[42]) & (!g923) & (!g1200)) + ((!g411) & (g667) & (!sk[42]) & (!g923) & (g1200)) + ((!g411) & (g667) & (!sk[42]) & (g923) & (!g1200)) + ((!g411) & (g667) & (!sk[42]) & (g923) & (g1200)) + ((!g411) & (g667) & (sk[42]) & (!g923) & (!g1200)) + ((!g411) & (g667) & (sk[42]) & (g923) & (g1200)) + ((g411) & (!g667) & (!sk[42]) & (g923) & (!g1200)) + ((g411) & (!g667) & (!sk[42]) & (g923) & (g1200)) + ((g411) & (!g667) & (sk[42]) & (!g923) & (!g1200)) + ((g411) & (!g667) & (sk[42]) & (g923) & (g1200)) + ((g411) & (g667) & (!sk[42]) & (!g923) & (!g1200)) + ((g411) & (g667) & (!sk[42]) & (!g923) & (g1200)) + ((g411) & (g667) & (!sk[42]) & (g923) & (!g1200)) + ((g411) & (g667) & (!sk[42]) & (g923) & (g1200)) + ((g411) & (g667) & (sk[42]) & (!g923) & (g1200)) + ((g411) & (g667) & (sk[42]) & (g923) & (!g1200)));
	assign g1202 = (((!sk[43]) & (!ld) & (!g155) & (g1201) & (!keyx1x)) + ((!sk[43]) & (!ld) & (!g155) & (g1201) & (keyx1x)) + ((!sk[43]) & (!ld) & (g155) & (!g1201) & (!keyx1x)) + ((!sk[43]) & (!ld) & (g155) & (!g1201) & (keyx1x)) + ((!sk[43]) & (!ld) & (g155) & (g1201) & (!keyx1x)) + ((!sk[43]) & (!ld) & (g155) & (g1201) & (keyx1x)) + ((!sk[43]) & (ld) & (!g155) & (g1201) & (!keyx1x)) + ((!sk[43]) & (ld) & (!g155) & (g1201) & (keyx1x)) + ((!sk[43]) & (ld) & (g155) & (!g1201) & (!keyx1x)) + ((!sk[43]) & (ld) & (g155) & (!g1201) & (keyx1x)) + ((!sk[43]) & (ld) & (g155) & (g1201) & (!keyx1x)) + ((!sk[43]) & (ld) & (g155) & (g1201) & (keyx1x)) + ((sk[43]) & (!ld) & (!g155) & (g1201) & (!keyx1x)) + ((sk[43]) & (!ld) & (!g155) & (g1201) & (keyx1x)) + ((sk[43]) & (!ld) & (g155) & (!g1201) & (!keyx1x)) + ((sk[43]) & (!ld) & (g155) & (!g1201) & (keyx1x)) + ((sk[43]) & (ld) & (!g155) & (!g1201) & (keyx1x)) + ((sk[43]) & (ld) & (!g155) & (g1201) & (keyx1x)) + ((sk[43]) & (ld) & (g155) & (!g1201) & (keyx1x)) + ((sk[43]) & (ld) & (g155) & (g1201) & (keyx1x)));
	assign g1203 = (((!g382) & (!g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((!g382) & (!g347) & (!g354) & (!g361) & (g368) & (g375)) + ((!g382) & (!g347) & (!g354) & (g361) & (!g368) & (g375)) + ((!g382) & (!g347) & (!g354) & (g361) & (g368) & (!g375)) + ((!g382) & (!g347) & (!g354) & (g361) & (g368) & (g375)) + ((!g382) & (!g347) & (g354) & (!g361) & (!g368) & (g375)) + ((!g382) & (!g347) & (g354) & (g361) & (!g368) & (!g375)) + ((!g382) & (!g347) & (g354) & (g361) & (g368) & (!g375)) + ((!g382) & (g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((!g382) & (g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((!g382) & (g347) & (!g354) & (g361) & (!g368) & (g375)) + ((!g382) & (g347) & (g354) & (!g361) & (!g368) & (!g375)) + ((!g382) & (g347) & (g354) & (!g361) & (!g368) & (g375)) + ((!g382) & (g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g382) & (g347) & (g354) & (!g361) & (g368) & (g375)) + ((g382) & (!g347) & (!g354) & (g361) & (!g368) & (g375)) + ((g382) & (!g347) & (!g354) & (g361) & (g368) & (g375)) + ((g382) & (g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((g382) & (g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((g382) & (g347) & (!g354) & (g361) & (g368) & (!g375)) + ((g382) & (g347) & (g354) & (g361) & (!g368) & (!g375)) + ((g382) & (g347) & (g354) & (g361) & (!g368) & (g375)));
	assign g1204 = (((!g382) & (!g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((!g382) & (!g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((!g382) & (!g347) & (!g354) & (g361) & (g368) & (g375)) + ((!g382) & (!g347) & (g354) & (!g361) & (!g368) & (!g375)) + ((!g382) & (!g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g382) & (!g347) & (g354) & (g361) & (!g368) & (g375)) + ((!g382) & (g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((!g382) & (g347) & (!g354) & (!g361) & (g368) & (g375)) + ((!g382) & (g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((!g382) & (g347) & (!g354) & (g361) & (!g368) & (g375)) + ((!g382) & (g347) & (!g354) & (g361) & (g368) & (g375)) + ((!g382) & (g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g382) & (g347) & (g354) & (!g361) & (g368) & (g375)) + ((!g382) & (g347) & (g354) & (g361) & (g368) & (!g375)) + ((g382) & (!g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((g382) & (!g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((g382) & (!g347) & (!g354) & (!g361) & (g368) & (g375)) + ((g382) & (!g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((g382) & (!g347) & (!g354) & (g361) & (!g368) & (g375)) + ((g382) & (!g347) & (!g354) & (g361) & (g368) & (!g375)) + ((g382) & (!g347) & (g354) & (g361) & (!g368) & (!g375)) + ((g382) & (g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((g382) & (g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((g382) & (g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((g382) & (g347) & (!g354) & (g361) & (g368) & (!g375)) + ((g382) & (g347) & (!g354) & (g361) & (g368) & (g375)) + ((g382) & (g347) & (g354) & (!g361) & (!g368) & (!g375)) + ((g382) & (g347) & (g354) & (!g361) & (g368) & (!g375)) + ((g382) & (g347) & (g354) & (g361) & (!g368) & (g375)) + ((g382) & (g347) & (g354) & (g361) & (g368) & (g375)));
	assign g1205 = (((!g382) & (!g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((!g382) & (!g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((!g382) & (!g347) & (!g354) & (g361) & (!g368) & (g375)) + ((!g382) & (!g347) & (g354) & (!g361) & (!g368) & (g375)) + ((!g382) & (!g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g382) & (!g347) & (g354) & (g361) & (!g368) & (g375)) + ((!g382) & (g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((!g382) & (g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((!g382) & (g347) & (!g354) & (g361) & (g368) & (!g375)) + ((!g382) & (g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g382) & (g347) & (g354) & (g361) & (!g368) & (!g375)) + ((!g382) & (g347) & (g354) & (g361) & (g368) & (!g375)) + ((g382) & (!g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((g382) & (!g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((g382) & (!g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((g382) & (!g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((g382) & (!g347) & (!g354) & (g361) & (!g368) & (g375)) + ((g382) & (!g347) & (!g354) & (g361) & (g368) & (!g375)) + ((g382) & (!g347) & (!g354) & (g361) & (g368) & (g375)) + ((g382) & (!g347) & (g354) & (!g361) & (!g368) & (g375)) + ((g382) & (!g347) & (g354) & (!g361) & (g368) & (!g375)) + ((g382) & (!g347) & (g354) & (g361) & (!g368) & (!g375)) + ((g382) & (!g347) & (g354) & (g361) & (g368) & (g375)) + ((g382) & (g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((g382) & (g347) & (!g354) & (!g361) & (g368) & (g375)) + ((g382) & (g347) & (g354) & (!g361) & (g368) & (g375)) + ((g382) & (g347) & (g354) & (g361) & (!g368) & (!g375)) + ((g382) & (g347) & (g354) & (g361) & (!g368) & (g375)) + ((g382) & (g347) & (g354) & (g361) & (g368) & (g375)));
	assign g1206 = (((!g382) & (!g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((!g382) & (!g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((!g382) & (!g347) & (!g354) & (!g361) & (g368) & (g375)) + ((!g382) & (!g347) & (!g354) & (g361) & (!g368) & (g375)) + ((!g382) & (!g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g382) & (!g347) & (g354) & (g361) & (g368) & (g375)) + ((!g382) & (g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((!g382) & (g347) & (!g354) & (g361) & (!g368) & (g375)) + ((!g382) & (g347) & (!g354) & (g361) & (g368) & (g375)) + ((!g382) & (g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g382) & (g347) & (g354) & (!g361) & (g368) & (g375)) + ((!g382) & (g347) & (g354) & (g361) & (!g368) & (!g375)) + ((!g382) & (g347) & (g354) & (g361) & (!g368) & (g375)) + ((!g382) & (g347) & (g354) & (g361) & (g368) & (!g375)) + ((!g382) & (g347) & (g354) & (g361) & (g368) & (g375)) + ((g382) & (!g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((g382) & (!g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((g382) & (!g347) & (!g354) & (!g361) & (g368) & (g375)) + ((g382) & (!g347) & (!g354) & (g361) & (g368) & (g375)) + ((g382) & (!g347) & (g354) & (!g361) & (!g368) & (g375)) + ((g382) & (!g347) & (g354) & (!g361) & (g368) & (!g375)) + ((g382) & (!g347) & (g354) & (g361) & (g368) & (!g375)) + ((g382) & (g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((g382) & (g347) & (!g354) & (g361) & (!g368) & (g375)) + ((g382) & (g347) & (!g354) & (g361) & (g368) & (!g375)) + ((g382) & (g347) & (g354) & (!g361) & (g368) & (g375)) + ((g382) & (g347) & (g354) & (g361) & (!g368) & (!g375)));
	assign g1207 = (((!g1203) & (!g1204) & (!g1205) & (!g1206) & (!g340) & (g389)) + ((!g1203) & (!g1204) & (!g1205) & (!g1206) & (g340) & (!g389)) + ((!g1203) & (!g1204) & (!g1205) & (!g1206) & (g340) & (g389)) + ((!g1203) & (!g1204) & (!g1205) & (g1206) & (!g340) & (g389)) + ((!g1203) & (!g1204) & (!g1205) & (g1206) & (g340) & (!g389)) + ((!g1203) & (!g1204) & (g1205) & (!g1206) & (g340) & (!g389)) + ((!g1203) & (!g1204) & (g1205) & (!g1206) & (g340) & (g389)) + ((!g1203) & (!g1204) & (g1205) & (g1206) & (g340) & (!g389)) + ((!g1203) & (g1204) & (!g1205) & (!g1206) & (!g340) & (g389)) + ((!g1203) & (g1204) & (!g1205) & (!g1206) & (g340) & (g389)) + ((!g1203) & (g1204) & (!g1205) & (g1206) & (!g340) & (g389)) + ((!g1203) & (g1204) & (g1205) & (!g1206) & (g340) & (g389)) + ((g1203) & (!g1204) & (!g1205) & (!g1206) & (!g340) & (!g389)) + ((g1203) & (!g1204) & (!g1205) & (!g1206) & (!g340) & (g389)) + ((g1203) & (!g1204) & (!g1205) & (!g1206) & (g340) & (!g389)) + ((g1203) & (!g1204) & (!g1205) & (!g1206) & (g340) & (g389)) + ((g1203) & (!g1204) & (!g1205) & (g1206) & (!g340) & (!g389)) + ((g1203) & (!g1204) & (!g1205) & (g1206) & (!g340) & (g389)) + ((g1203) & (!g1204) & (!g1205) & (g1206) & (g340) & (!g389)) + ((g1203) & (!g1204) & (g1205) & (!g1206) & (!g340) & (!g389)) + ((g1203) & (!g1204) & (g1205) & (!g1206) & (g340) & (!g389)) + ((g1203) & (!g1204) & (g1205) & (!g1206) & (g340) & (g389)) + ((g1203) & (!g1204) & (g1205) & (g1206) & (!g340) & (!g389)) + ((g1203) & (!g1204) & (g1205) & (g1206) & (g340) & (!g389)) + ((g1203) & (g1204) & (!g1205) & (!g1206) & (!g340) & (!g389)) + ((g1203) & (g1204) & (!g1205) & (!g1206) & (!g340) & (g389)) + ((g1203) & (g1204) & (!g1205) & (!g1206) & (g340) & (g389)) + ((g1203) & (g1204) & (!g1205) & (g1206) & (!g340) & (!g389)) + ((g1203) & (g1204) & (!g1205) & (g1206) & (!g340) & (g389)) + ((g1203) & (g1204) & (g1205) & (!g1206) & (!g340) & (!g389)) + ((g1203) & (g1204) & (g1205) & (!g1206) & (g340) & (g389)) + ((g1203) & (g1204) & (g1205) & (g1206) & (!g340) & (!g389)));
	assign g1208 = (((!sk[49]) & (!g418) & (!g674) & (g930) & (!g1207)) + ((!sk[49]) & (!g418) & (!g674) & (g930) & (g1207)) + ((!sk[49]) & (!g418) & (g674) & (!g930) & (!g1207)) + ((!sk[49]) & (!g418) & (g674) & (!g930) & (g1207)) + ((!sk[49]) & (!g418) & (g674) & (g930) & (!g1207)) + ((!sk[49]) & (!g418) & (g674) & (g930) & (g1207)) + ((!sk[49]) & (g418) & (!g674) & (g930) & (!g1207)) + ((!sk[49]) & (g418) & (!g674) & (g930) & (g1207)) + ((!sk[49]) & (g418) & (g674) & (!g930) & (!g1207)) + ((!sk[49]) & (g418) & (g674) & (!g930) & (g1207)) + ((!sk[49]) & (g418) & (g674) & (g930) & (!g1207)) + ((!sk[49]) & (g418) & (g674) & (g930) & (g1207)) + ((sk[49]) & (!g418) & (!g674) & (!g930) & (g1207)) + ((sk[49]) & (!g418) & (!g674) & (g930) & (!g1207)) + ((sk[49]) & (!g418) & (g674) & (!g930) & (!g1207)) + ((sk[49]) & (!g418) & (g674) & (g930) & (g1207)) + ((sk[49]) & (g418) & (!g674) & (!g930) & (!g1207)) + ((sk[49]) & (g418) & (!g674) & (g930) & (g1207)) + ((sk[49]) & (g418) & (g674) & (!g930) & (g1207)) + ((sk[49]) & (g418) & (g674) & (g930) & (!g1207)));
	assign g1209 = (((!sk[50]) & (!ld) & (!g162) & (g1208) & (!keyx2x)) + ((!sk[50]) & (!ld) & (!g162) & (g1208) & (keyx2x)) + ((!sk[50]) & (!ld) & (g162) & (!g1208) & (!keyx2x)) + ((!sk[50]) & (!ld) & (g162) & (!g1208) & (keyx2x)) + ((!sk[50]) & (!ld) & (g162) & (g1208) & (!keyx2x)) + ((!sk[50]) & (!ld) & (g162) & (g1208) & (keyx2x)) + ((!sk[50]) & (ld) & (!g162) & (g1208) & (!keyx2x)) + ((!sk[50]) & (ld) & (!g162) & (g1208) & (keyx2x)) + ((!sk[50]) & (ld) & (g162) & (!g1208) & (!keyx2x)) + ((!sk[50]) & (ld) & (g162) & (!g1208) & (keyx2x)) + ((!sk[50]) & (ld) & (g162) & (g1208) & (!keyx2x)) + ((!sk[50]) & (ld) & (g162) & (g1208) & (keyx2x)) + ((sk[50]) & (!ld) & (!g162) & (g1208) & (!keyx2x)) + ((sk[50]) & (!ld) & (!g162) & (g1208) & (keyx2x)) + ((sk[50]) & (!ld) & (g162) & (!g1208) & (!keyx2x)) + ((sk[50]) & (!ld) & (g162) & (!g1208) & (keyx2x)) + ((sk[50]) & (ld) & (!g162) & (!g1208) & (keyx2x)) + ((sk[50]) & (ld) & (!g162) & (g1208) & (keyx2x)) + ((sk[50]) & (ld) & (g162) & (!g1208) & (keyx2x)) + ((sk[50]) & (ld) & (g162) & (g1208) & (keyx2x)));
	assign g1210 = (((!g340) & (!g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (g368) & (g375)) + ((!g340) & (!g347) & (g354) & (g361) & (!g368) & (!g375)) + ((!g340) & (!g347) & (g354) & (g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (g354) & (g361) & (g368) & (g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (g347) & (g354) & (!g361) & (!g368) & (!g375)) + ((!g340) & (g347) & (g354) & (g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((g340) & (!g347) & (g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (g354) & (!g361) & (!g368) & (g375)) + ((g340) & (!g347) & (g354) & (!g361) & (g368) & (!g375)) + ((g340) & (!g347) & (g354) & (g361) & (!g368) & (g375)) + ((g340) & (g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((g340) & (g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((g340) & (g347) & (!g354) & (g361) & (g368) & (!g375)) + ((g340) & (g347) & (g354) & (!g361) & (!g368) & (g375)) + ((g340) & (g347) & (g354) & (!g361) & (g368) & (g375)));
	assign g1211 = (((!g340) & (!g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (!g354) & (!g361) & (g368) & (g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (g354) & (g361) & (!g368) & (!g375)) + ((!g340) & (!g347) & (g354) & (g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (g354) & (g361) & (g368) & (g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (g368) & (g375)) + ((!g340) & (g347) & (!g354) & (g361) & (g368) & (g375)) + ((!g340) & (g347) & (g354) & (!g361) & (!g368) & (!g375)) + ((!g340) & (g347) & (g354) & (!g361) & (!g368) & (g375)) + ((!g340) & (g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (g347) & (g354) & (g361) & (!g368) & (g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((g340) & (!g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (!g354) & (g361) & (!g368) & (g375)) + ((g340) & (!g347) & (!g354) & (g361) & (g368) & (g375)) + ((g340) & (!g347) & (g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (g354) & (!g361) & (!g368) & (g375)) + ((g340) & (!g347) & (g354) & (!g361) & (g368) & (g375)) + ((g340) & (!g347) & (g354) & (g361) & (!g368) & (g375)) + ((g340) & (g347) & (!g354) & (g361) & (!g368) & (g375)) + ((g340) & (g347) & (!g354) & (g361) & (g368) & (!g375)) + ((g340) & (g347) & (g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (g347) & (g354) & (g361) & (!g368) & (!g375)));
	assign g1212 = (((!g340) & (!g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (!g354) & (!g361) & (g368) & (g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (g354) & (!g361) & (g368) & (g375)) + ((!g340) & (!g347) & (g354) & (g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (g354) & (g361) & (g368) & (g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (g368) & (g375)) + ((!g340) & (g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((!g340) & (g347) & (!g354) & (g361) & (!g368) & (g375)) + ((!g340) & (g347) & (g354) & (!g361) & (!g368) & (g375)) + ((!g340) & (g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (g347) & (g354) & (g361) & (g368) & (g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (g368) & (g375)) + ((g340) & (!g347) & (!g354) & (g361) & (g368) & (g375)) + ((g340) & (!g347) & (g354) & (g361) & (!g368) & (!g375)) + ((g340) & (g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((g340) & (g347) & (!g354) & (g361) & (g368) & (g375)) + ((g340) & (g347) & (g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (g347) & (g354) & (!g361) & (!g368) & (g375)) + ((g340) & (g347) & (g354) & (!g361) & (g368) & (g375)) + ((g340) & (g347) & (g354) & (g361) & (!g368) & (!g375)) + ((g340) & (g347) & (g354) & (g361) & (g368) & (g375)));
	assign g1213 = (((!g340) & (!g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (!g354) & (g361) & (g368) & (g375)) + ((!g340) & (!g347) & (g354) & (g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (g354) & (g361) & (g368) & (g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (!g368) & (!g375)) + ((!g340) & (g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (g347) & (!g354) & (g361) & (!g368) & (!g375)) + ((!g340) & (g347) & (!g354) & (g361) & (!g368) & (g375)) + ((!g340) & (g347) & (!g354) & (g361) & (g368) & (!g375)) + ((!g340) & (g347) & (g354) & (!g361) & (!g368) & (!g375)) + ((!g340) & (g347) & (g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (g347) & (g354) & (!g361) & (g368) & (g375)) + ((g340) & (!g347) & (!g354) & (!g361) & (g368) & (g375)) + ((g340) & (!g347) & (!g354) & (g361) & (g368) & (!g375)) + ((g340) & (!g347) & (g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (g354) & (!g361) & (g368) & (!g375)) + ((g340) & (!g347) & (g354) & (!g361) & (g368) & (g375)) + ((g340) & (!g347) & (g354) & (g361) & (!g368) & (g375)) + ((g340) & (!g347) & (g354) & (g361) & (g368) & (!g375)) + ((g340) & (!g347) & (g354) & (g361) & (g368) & (g375)) + ((g340) & (g347) & (!g354) & (!g361) & (!g368) & (g375)) + ((g340) & (g347) & (!g354) & (!g361) & (g368) & (!g375)) + ((g340) & (g347) & (g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (g347) & (g354) & (!g361) & (!g368) & (g375)) + ((g340) & (g347) & (g354) & (g361) & (g368) & (g375)));
	assign g1214 = (((!g1210) & (!g1211) & (!g1212) & (!g1213) & (!g389) & (g382)) + ((!g1210) & (!g1211) & (!g1212) & (!g1213) & (g389) & (!g382)) + ((!g1210) & (!g1211) & (!g1212) & (!g1213) & (g389) & (g382)) + ((!g1210) & (!g1211) & (!g1212) & (g1213) & (!g389) & (g382)) + ((!g1210) & (!g1211) & (!g1212) & (g1213) & (g389) & (!g382)) + ((!g1210) & (!g1211) & (g1212) & (!g1213) & (g389) & (!g382)) + ((!g1210) & (!g1211) & (g1212) & (!g1213) & (g389) & (g382)) + ((!g1210) & (!g1211) & (g1212) & (g1213) & (g389) & (!g382)) + ((!g1210) & (g1211) & (!g1212) & (!g1213) & (!g389) & (g382)) + ((!g1210) & (g1211) & (!g1212) & (!g1213) & (g389) & (g382)) + ((!g1210) & (g1211) & (!g1212) & (g1213) & (!g389) & (g382)) + ((!g1210) & (g1211) & (g1212) & (!g1213) & (g389) & (g382)) + ((g1210) & (!g1211) & (!g1212) & (!g1213) & (!g389) & (!g382)) + ((g1210) & (!g1211) & (!g1212) & (!g1213) & (!g389) & (g382)) + ((g1210) & (!g1211) & (!g1212) & (!g1213) & (g389) & (!g382)) + ((g1210) & (!g1211) & (!g1212) & (!g1213) & (g389) & (g382)) + ((g1210) & (!g1211) & (!g1212) & (g1213) & (!g389) & (!g382)) + ((g1210) & (!g1211) & (!g1212) & (g1213) & (!g389) & (g382)) + ((g1210) & (!g1211) & (!g1212) & (g1213) & (g389) & (!g382)) + ((g1210) & (!g1211) & (g1212) & (!g1213) & (!g389) & (!g382)) + ((g1210) & (!g1211) & (g1212) & (!g1213) & (g389) & (!g382)) + ((g1210) & (!g1211) & (g1212) & (!g1213) & (g389) & (g382)) + ((g1210) & (!g1211) & (g1212) & (g1213) & (!g389) & (!g382)) + ((g1210) & (!g1211) & (g1212) & (g1213) & (g389) & (!g382)) + ((g1210) & (g1211) & (!g1212) & (!g1213) & (!g389) & (!g382)) + ((g1210) & (g1211) & (!g1212) & (!g1213) & (!g389) & (g382)) + ((g1210) & (g1211) & (!g1212) & (!g1213) & (g389) & (g382)) + ((g1210) & (g1211) & (!g1212) & (g1213) & (!g389) & (!g382)) + ((g1210) & (g1211) & (!g1212) & (g1213) & (!g389) & (g382)) + ((g1210) & (g1211) & (g1212) & (!g1213) & (!g389) & (!g382)) + ((g1210) & (g1211) & (g1212) & (!g1213) & (g389) & (g382)) + ((g1210) & (g1211) & (g1212) & (g1213) & (!g389) & (!g382)));
	assign g1215 = (((!g425) & (!sk[56]) & (!g681) & (g937) & (!g1214)) + ((!g425) & (!sk[56]) & (!g681) & (g937) & (g1214)) + ((!g425) & (!sk[56]) & (g681) & (!g937) & (!g1214)) + ((!g425) & (!sk[56]) & (g681) & (!g937) & (g1214)) + ((!g425) & (!sk[56]) & (g681) & (g937) & (!g1214)) + ((!g425) & (!sk[56]) & (g681) & (g937) & (g1214)) + ((!g425) & (sk[56]) & (!g681) & (!g937) & (g1214)) + ((!g425) & (sk[56]) & (!g681) & (g937) & (!g1214)) + ((!g425) & (sk[56]) & (g681) & (!g937) & (!g1214)) + ((!g425) & (sk[56]) & (g681) & (g937) & (g1214)) + ((g425) & (!sk[56]) & (!g681) & (g937) & (!g1214)) + ((g425) & (!sk[56]) & (!g681) & (g937) & (g1214)) + ((g425) & (!sk[56]) & (g681) & (!g937) & (!g1214)) + ((g425) & (!sk[56]) & (g681) & (!g937) & (g1214)) + ((g425) & (!sk[56]) & (g681) & (g937) & (!g1214)) + ((g425) & (!sk[56]) & (g681) & (g937) & (g1214)) + ((g425) & (sk[56]) & (!g681) & (!g937) & (!g1214)) + ((g425) & (sk[56]) & (!g681) & (g937) & (g1214)) + ((g425) & (sk[56]) & (g681) & (!g937) & (g1214)) + ((g425) & (sk[56]) & (g681) & (g937) & (!g1214)));
	assign g1216 = (((!ld) & (!sk[57]) & (!g169) & (g1215) & (!keyx3x)) + ((!ld) & (!sk[57]) & (!g169) & (g1215) & (keyx3x)) + ((!ld) & (!sk[57]) & (g169) & (!g1215) & (!keyx3x)) + ((!ld) & (!sk[57]) & (g169) & (!g1215) & (keyx3x)) + ((!ld) & (!sk[57]) & (g169) & (g1215) & (!keyx3x)) + ((!ld) & (!sk[57]) & (g169) & (g1215) & (keyx3x)) + ((!ld) & (sk[57]) & (!g169) & (g1215) & (!keyx3x)) + ((!ld) & (sk[57]) & (!g169) & (g1215) & (keyx3x)) + ((!ld) & (sk[57]) & (g169) & (!g1215) & (!keyx3x)) + ((!ld) & (sk[57]) & (g169) & (!g1215) & (keyx3x)) + ((ld) & (!sk[57]) & (!g169) & (g1215) & (!keyx3x)) + ((ld) & (!sk[57]) & (!g169) & (g1215) & (keyx3x)) + ((ld) & (!sk[57]) & (g169) & (!g1215) & (!keyx3x)) + ((ld) & (!sk[57]) & (g169) & (!g1215) & (keyx3x)) + ((ld) & (!sk[57]) & (g169) & (g1215) & (!keyx3x)) + ((ld) & (!sk[57]) & (g169) & (g1215) & (keyx3x)) + ((ld) & (sk[57]) & (!g169) & (!g1215) & (keyx3x)) + ((ld) & (sk[57]) & (!g169) & (g1215) & (keyx3x)) + ((ld) & (sk[57]) & (g169) & (!g1215) & (keyx3x)) + ((ld) & (sk[57]) & (g169) & (g1215) & (keyx3x)));
	assign g1217 = (((!g340) & (!g347) & (!g382) & (!g389) & (!g368) & (g375)) + ((!g340) & (!g347) & (g382) & (!g389) & (!g368) & (g375)) + ((!g340) & (!g347) & (g382) & (!g389) & (g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (!g389) & (g368) & (g375)) + ((!g340) & (!g347) & (g382) & (g389) & (!g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (g389) & (g368) & (!g375)) + ((!g340) & (g347) & (!g382) & (!g389) & (!g368) & (!g375)) + ((!g340) & (g347) & (!g382) & (!g389) & (!g368) & (g375)) + ((!g340) & (g347) & (!g382) & (g389) & (!g368) & (!g375)) + ((!g340) & (g347) & (!g382) & (g389) & (!g368) & (g375)) + ((!g340) & (g347) & (!g382) & (g389) & (g368) & (g375)) + ((!g340) & (g347) & (g382) & (g389) & (!g368) & (g375)) + ((!g340) & (g347) & (g382) & (g389) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g389) & (!g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g389) & (!g368) & (g375)) + ((g340) & (!g347) & (!g382) & (g389) & (!g368) & (g375)) + ((g340) & (!g347) & (g382) & (!g389) & (g368) & (!g375)) + ((g340) & (!g347) & (g382) & (g389) & (!g368) & (!g375)) + ((g340) & (!g347) & (g382) & (g389) & (!g368) & (g375)) + ((g340) & (!g347) & (g382) & (g389) & (g368) & (!g375)) + ((g340) & (g347) & (!g382) & (!g389) & (!g368) & (!g375)) + ((g340) & (g347) & (!g382) & (!g389) & (g368) & (!g375)) + ((g340) & (g347) & (!g382) & (g389) & (g368) & (!g375)) + ((g340) & (g347) & (g382) & (!g389) & (!g368) & (!g375)) + ((g340) & (g347) & (g382) & (!g389) & (!g368) & (g375)) + ((g340) & (g347) & (g382) & (g389) & (!g368) & (g375)));
	assign g1218 = (((!g340) & (!g347) & (!g382) & (!g389) & (!g368) & (!g375)) + ((!g340) & (!g347) & (!g382) & (!g389) & (!g368) & (g375)) + ((!g340) & (!g347) & (!g382) & (!g389) & (g368) & (!g375)) + ((!g340) & (!g347) & (!g382) & (!g389) & (g368) & (g375)) + ((!g340) & (!g347) & (!g382) & (g389) & (!g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (!g389) & (!g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (!g389) & (g368) & (g375)) + ((!g340) & (!g347) & (g382) & (g389) & (!g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (g389) & (g368) & (g375)) + ((!g340) & (g347) & (!g382) & (!g389) & (!g368) & (g375)) + ((!g340) & (g347) & (!g382) & (g389) & (g368) & (!g375)) + ((!g340) & (g347) & (g382) & (!g389) & (!g368) & (!g375)) + ((!g340) & (g347) & (g382) & (!g389) & (!g368) & (g375)) + ((!g340) & (g347) & (g382) & (!g389) & (g368) & (!g375)) + ((!g340) & (g347) & (g382) & (!g389) & (g368) & (g375)) + ((!g340) & (g347) & (g382) & (g389) & (!g368) & (!g375)) + ((!g340) & (g347) & (g382) & (g389) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g389) & (!g368) & (g375)) + ((g340) & (!g347) & (!g382) & (!g389) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g389) & (g368) & (g375)) + ((g340) & (!g347) & (!g382) & (g389) & (!g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (g389) & (g368) & (g375)) + ((g340) & (!g347) & (g382) & (!g389) & (g368) & (!g375)) + ((g340) & (!g347) & (g382) & (!g389) & (g368) & (g375)) + ((g340) & (!g347) & (g382) & (g389) & (!g368) & (g375)) + ((g340) & (g347) & (!g382) & (!g389) & (g368) & (!g375)) + ((g340) & (g347) & (!g382) & (!g389) & (g368) & (g375)) + ((g340) & (g347) & (!g382) & (g389) & (!g368) & (!g375)) + ((g340) & (g347) & (!g382) & (g389) & (!g368) & (g375)) + ((g340) & (g347) & (g382) & (!g389) & (g368) & (!g375)) + ((g340) & (g347) & (g382) & (!g389) & (g368) & (g375)) + ((g340) & (g347) & (g382) & (g389) & (!g368) & (g375)));
	assign g1219 = (((!g340) & (!g347) & (!g382) & (!g389) & (!g368) & (!g375)) + ((!g340) & (!g347) & (!g382) & (!g389) & (!g368) & (g375)) + ((!g340) & (!g347) & (g382) & (!g389) & (!g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (!g389) & (g368) & (g375)) + ((!g340) & (!g347) & (g382) & (g389) & (!g368) & (g375)) + ((!g340) & (g347) & (!g382) & (g389) & (!g368) & (!g375)) + ((!g340) & (g347) & (!g382) & (g389) & (g368) & (!g375)) + ((!g340) & (g347) & (!g382) & (g389) & (g368) & (g375)) + ((!g340) & (g347) & (g382) & (!g389) & (!g368) & (!g375)) + ((!g340) & (g347) & (g382) & (!g389) & (g368) & (!g375)) + ((!g340) & (g347) & (g382) & (!g389) & (g368) & (g375)) + ((!g340) & (g347) & (g382) & (g389) & (!g368) & (!g375)) + ((!g340) & (g347) & (g382) & (g389) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g389) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g389) & (g368) & (g375)) + ((g340) & (!g347) & (!g382) & (g389) & (!g368) & (g375)) + ((g340) & (!g347) & (!g382) & (g389) & (g368) & (g375)) + ((g340) & (!g347) & (g382) & (!g389) & (!g368) & (!g375)) + ((g340) & (!g347) & (g382) & (!g389) & (!g368) & (g375)) + ((g340) & (!g347) & (g382) & (!g389) & (g368) & (g375)) + ((g340) & (!g347) & (g382) & (g389) & (!g368) & (!g375)) + ((g340) & (!g347) & (g382) & (g389) & (!g368) & (g375)) + ((g340) & (!g347) & (g382) & (g389) & (g368) & (!g375)) + ((g340) & (!g347) & (g382) & (g389) & (g368) & (g375)) + ((g340) & (g347) & (!g382) & (!g389) & (!g368) & (g375)) + ((g340) & (g347) & (!g382) & (g389) & (!g368) & (!g375)) + ((g340) & (g347) & (!g382) & (g389) & (g368) & (!g375)) + ((g340) & (g347) & (g382) & (!g389) & (!g368) & (!g375)) + ((g340) & (g347) & (g382) & (!g389) & (!g368) & (g375)) + ((g340) & (g347) & (g382) & (!g389) & (g368) & (!g375)) + ((g340) & (g347) & (g382) & (g389) & (!g368) & (!g375)) + ((g340) & (g347) & (g382) & (g389) & (g368) & (!g375)));
	assign g1220 = (((!g340) & (!g347) & (!g382) & (!g389) & (g368) & (g375)) + ((!g340) & (!g347) & (!g382) & (g389) & (!g368) & (!g375)) + ((!g340) & (!g347) & (!g382) & (g389) & (g368) & (g375)) + ((!g340) & (!g347) & (g382) & (!g389) & (!g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (!g389) & (g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (g389) & (!g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (g389) & (!g368) & (g375)) + ((!g340) & (!g347) & (g382) & (g389) & (g368) & (!g375)) + ((!g340) & (g347) & (!g382) & (!g389) & (!g368) & (!g375)) + ((!g340) & (g347) & (!g382) & (g389) & (!g368) & (g375)) + ((!g340) & (g347) & (!g382) & (g389) & (g368) & (!g375)) + ((!g340) & (g347) & (!g382) & (g389) & (g368) & (g375)) + ((!g340) & (g347) & (g382) & (!g389) & (!g368) & (!g375)) + ((!g340) & (g347) & (g382) & (g389) & (!g368) & (!g375)) + ((!g340) & (g347) & (g382) & (g389) & (!g368) & (g375)) + ((g340) & (!g347) & (!g382) & (!g389) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g389) & (g368) & (g375)) + ((g340) & (!g347) & (g382) & (!g389) & (!g368) & (!g375)) + ((g340) & (!g347) & (g382) & (!g389) & (g368) & (!g375)) + ((g340) & (!g347) & (g382) & (g389) & (g368) & (!g375)) + ((g340) & (g347) & (!g382) & (!g389) & (g368) & (!g375)) + ((g340) & (g347) & (!g382) & (g389) & (g368) & (g375)) + ((g340) & (g347) & (g382) & (!g389) & (!g368) & (!g375)) + ((g340) & (g347) & (g382) & (!g389) & (!g368) & (g375)) + ((g340) & (g347) & (g382) & (!g389) & (g368) & (!g375)) + ((g340) & (g347) & (g382) & (g389) & (!g368) & (!g375)));
	assign g1221 = (((!g1217) & (!g1218) & (!g1219) & (!g1220) & (g354) & (g361)) + ((!g1217) & (!g1218) & (g1219) & (!g1220) & (!g354) & (g361)) + ((!g1217) & (!g1218) & (g1219) & (!g1220) & (g354) & (g361)) + ((!g1217) & (!g1218) & (g1219) & (g1220) & (!g354) & (g361)) + ((!g1217) & (g1218) & (!g1219) & (!g1220) & (g354) & (!g361)) + ((!g1217) & (g1218) & (!g1219) & (!g1220) & (g354) & (g361)) + ((!g1217) & (g1218) & (!g1219) & (g1220) & (g354) & (!g361)) + ((!g1217) & (g1218) & (g1219) & (!g1220) & (!g354) & (g361)) + ((!g1217) & (g1218) & (g1219) & (!g1220) & (g354) & (!g361)) + ((!g1217) & (g1218) & (g1219) & (!g1220) & (g354) & (g361)) + ((!g1217) & (g1218) & (g1219) & (g1220) & (!g354) & (g361)) + ((!g1217) & (g1218) & (g1219) & (g1220) & (g354) & (!g361)) + ((g1217) & (!g1218) & (!g1219) & (!g1220) & (!g354) & (!g361)) + ((g1217) & (!g1218) & (!g1219) & (!g1220) & (g354) & (g361)) + ((g1217) & (!g1218) & (!g1219) & (g1220) & (!g354) & (!g361)) + ((g1217) & (!g1218) & (g1219) & (!g1220) & (!g354) & (!g361)) + ((g1217) & (!g1218) & (g1219) & (!g1220) & (!g354) & (g361)) + ((g1217) & (!g1218) & (g1219) & (!g1220) & (g354) & (g361)) + ((g1217) & (!g1218) & (g1219) & (g1220) & (!g354) & (!g361)) + ((g1217) & (!g1218) & (g1219) & (g1220) & (!g354) & (g361)) + ((g1217) & (g1218) & (!g1219) & (!g1220) & (!g354) & (!g361)) + ((g1217) & (g1218) & (!g1219) & (!g1220) & (g354) & (!g361)) + ((g1217) & (g1218) & (!g1219) & (!g1220) & (g354) & (g361)) + ((g1217) & (g1218) & (!g1219) & (g1220) & (!g354) & (!g361)) + ((g1217) & (g1218) & (!g1219) & (g1220) & (g354) & (!g361)) + ((g1217) & (g1218) & (g1219) & (!g1220) & (!g354) & (!g361)) + ((g1217) & (g1218) & (g1219) & (!g1220) & (!g354) & (g361)) + ((g1217) & (g1218) & (g1219) & (!g1220) & (g354) & (!g361)) + ((g1217) & (g1218) & (g1219) & (!g1220) & (g354) & (g361)) + ((g1217) & (g1218) & (g1219) & (g1220) & (!g354) & (!g361)) + ((g1217) & (g1218) & (g1219) & (g1220) & (!g354) & (g361)) + ((g1217) & (g1218) & (g1219) & (g1220) & (g354) & (!g361)));
	assign g1222 = (((!g432) & (!g688) & (!g944) & (sk[63]) & (g1221)) + ((!g432) & (!g688) & (g944) & (!sk[63]) & (!g1221)) + ((!g432) & (!g688) & (g944) & (!sk[63]) & (g1221)) + ((!g432) & (!g688) & (g944) & (sk[63]) & (!g1221)) + ((!g432) & (g688) & (!g944) & (!sk[63]) & (!g1221)) + ((!g432) & (g688) & (!g944) & (!sk[63]) & (g1221)) + ((!g432) & (g688) & (!g944) & (sk[63]) & (!g1221)) + ((!g432) & (g688) & (g944) & (!sk[63]) & (!g1221)) + ((!g432) & (g688) & (g944) & (!sk[63]) & (g1221)) + ((!g432) & (g688) & (g944) & (sk[63]) & (g1221)) + ((g432) & (!g688) & (!g944) & (sk[63]) & (!g1221)) + ((g432) & (!g688) & (g944) & (!sk[63]) & (!g1221)) + ((g432) & (!g688) & (g944) & (!sk[63]) & (g1221)) + ((g432) & (!g688) & (g944) & (sk[63]) & (g1221)) + ((g432) & (g688) & (!g944) & (!sk[63]) & (!g1221)) + ((g432) & (g688) & (!g944) & (!sk[63]) & (g1221)) + ((g432) & (g688) & (!g944) & (sk[63]) & (g1221)) + ((g432) & (g688) & (g944) & (!sk[63]) & (!g1221)) + ((g432) & (g688) & (g944) & (!sk[63]) & (g1221)) + ((g432) & (g688) & (g944) & (sk[63]) & (!g1221)));
	assign g1223 = (((!ld) & (!g176) & (!sk[64]) & (g1222) & (!keyx4x)) + ((!ld) & (!g176) & (!sk[64]) & (g1222) & (keyx4x)) + ((!ld) & (!g176) & (sk[64]) & (g1222) & (!keyx4x)) + ((!ld) & (!g176) & (sk[64]) & (g1222) & (keyx4x)) + ((!ld) & (g176) & (!sk[64]) & (!g1222) & (!keyx4x)) + ((!ld) & (g176) & (!sk[64]) & (!g1222) & (keyx4x)) + ((!ld) & (g176) & (!sk[64]) & (g1222) & (!keyx4x)) + ((!ld) & (g176) & (!sk[64]) & (g1222) & (keyx4x)) + ((!ld) & (g176) & (sk[64]) & (!g1222) & (!keyx4x)) + ((!ld) & (g176) & (sk[64]) & (!g1222) & (keyx4x)) + ((ld) & (!g176) & (!sk[64]) & (g1222) & (!keyx4x)) + ((ld) & (!g176) & (!sk[64]) & (g1222) & (keyx4x)) + ((ld) & (!g176) & (sk[64]) & (!g1222) & (keyx4x)) + ((ld) & (!g176) & (sk[64]) & (g1222) & (keyx4x)) + ((ld) & (g176) & (!sk[64]) & (!g1222) & (!keyx4x)) + ((ld) & (g176) & (!sk[64]) & (!g1222) & (keyx4x)) + ((ld) & (g176) & (!sk[64]) & (g1222) & (!keyx4x)) + ((ld) & (g176) & (!sk[64]) & (g1222) & (keyx4x)) + ((ld) & (g176) & (sk[64]) & (!g1222) & (keyx4x)) + ((ld) & (g176) & (sk[64]) & (g1222) & (keyx4x)));
	assign g1224 = (((!g340) & (!g347) & (!g382) & (!g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (!g382) & (!g361) & (g368) & (g375)) + ((!g340) & (!g347) & (!g382) & (g361) & (g368) & (g375)) + ((!g340) & (!g347) & (g382) & (!g361) & (!g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (!g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (g382) & (!g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (!g361) & (g368) & (g375)) + ((!g340) & (!g347) & (g382) & (g361) & (!g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (g361) & (!g368) & (g375)) + ((!g340) & (g347) & (!g382) & (!g361) & (!g368) & (g375)) + ((!g340) & (g347) & (!g382) & (!g361) & (g368) & (!g375)) + ((!g340) & (g347) & (!g382) & (g361) & (g368) & (g375)) + ((!g340) & (g347) & (g382) & (!g361) & (g368) & (!g375)) + ((!g340) & (g347) & (g382) & (!g361) & (g368) & (g375)) + ((!g340) & (g347) & (g382) & (g361) & (!g368) & (!g375)) + ((!g340) & (g347) & (g382) & (g361) & (!g368) & (g375)) + ((!g340) & (g347) & (g382) & (g361) & (g368) & (g375)) + ((g340) & (!g347) & (!g382) & (!g361) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g361) & (g368) & (g375)) + ((g340) & (!g347) & (!g382) & (g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (g361) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (g361) & (g368) & (g375)) + ((g340) & (!g347) & (g382) & (!g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (g382) & (!g361) & (g368) & (!g375)) + ((g340) & (!g347) & (g382) & (g361) & (g368) & (!g375)) + ((g340) & (g347) & (!g382) & (!g361) & (g368) & (g375)) + ((g340) & (g347) & (g382) & (!g361) & (!g368) & (!g375)) + ((g340) & (g347) & (g382) & (!g361) & (g368) & (g375)));
	assign g1225 = (((!g340) & (!g347) & (!g382) & (!g361) & (!g368) & (!g375)) + ((!g340) & (!g347) & (!g382) & (g361) & (!g368) & (!g375)) + ((!g340) & (!g347) & (!g382) & (g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (!g382) & (g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (!g361) & (g368) & (g375)) + ((!g340) & (!g347) & (g382) & (g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (g382) & (g361) & (g368) & (g375)) + ((!g340) & (g347) & (!g382) & (!g361) & (!g368) & (!g375)) + ((!g340) & (g347) & (!g382) & (!g361) & (g368) & (!g375)) + ((!g340) & (g347) & (g382) & (!g361) & (!g368) & (g375)) + ((!g340) & (g347) & (g382) & (!g361) & (g368) & (g375)) + ((!g340) & (g347) & (g382) & (g361) & (!g368) & (g375)) + ((!g340) & (g347) & (g382) & (g361) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g361) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g361) & (g368) & (g375)) + ((g340) & (!g347) & (!g382) & (g361) & (!g368) & (g375)) + ((g340) & (!g347) & (!g382) & (g361) & (g368) & (g375)) + ((g340) & (!g347) & (g382) & (g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (g382) & (g361) & (!g368) & (g375)) + ((g340) & (!g347) & (g382) & (g361) & (g368) & (g375)) + ((g340) & (g347) & (!g382) & (!g361) & (!g368) & (g375)) + ((g340) & (g347) & (!g382) & (!g361) & (g368) & (!g375)) + ((g340) & (g347) & (!g382) & (g361) & (g368) & (!g375)) + ((g340) & (g347) & (g382) & (!g361) & (!g368) & (g375)) + ((g340) & (g347) & (g382) & (!g361) & (g368) & (g375)) + ((g340) & (g347) & (g382) & (g361) & (!g368) & (!g375)) + ((g340) & (g347) & (g382) & (g361) & (g368) & (g375)));
	assign g1226 = (((!g340) & (!g347) & (!g382) & (!g361) & (g368) & (g375)) + ((!g340) & (!g347) & (!g382) & (g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (!g361) & (!g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (!g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (g382) & (!g361) & (g368) & (g375)) + ((!g340) & (!g347) & (g382) & (g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (g382) & (g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (g382) & (g361) & (g368) & (g375)) + ((!g340) & (g347) & (!g382) & (!g361) & (g368) & (!g375)) + ((!g340) & (g347) & (!g382) & (!g361) & (g368) & (g375)) + ((!g340) & (g347) & (g382) & (!g361) & (!g368) & (!g375)) + ((!g340) & (g347) & (g382) & (g361) & (!g368) & (g375)) + ((!g340) & (g347) & (g382) & (g361) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g361) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (!g361) & (g368) & (g375)) + ((g340) & (!g347) & (!g382) & (g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (g361) & (!g368) & (g375)) + ((g340) & (!g347) & (g382) & (!g361) & (!g368) & (g375)) + ((g340) & (!g347) & (g382) & (!g361) & (g368) & (g375)) + ((g340) & (!g347) & (g382) & (g361) & (g368) & (!g375)) + ((g340) & (g347) & (!g382) & (!g361) & (!g368) & (!g375)) + ((g340) & (g347) & (!g382) & (!g361) & (!g368) & (g375)) + ((g340) & (g347) & (!g382) & (!g361) & (g368) & (g375)) + ((g340) & (g347) & (!g382) & (g361) & (!g368) & (g375)) + ((g340) & (g347) & (!g382) & (g361) & (g368) & (!g375)) + ((g340) & (g347) & (g382) & (!g361) & (!g368) & (g375)) + ((g340) & (g347) & (g382) & (!g361) & (g368) & (!g375)) + ((g340) & (g347) & (g382) & (g361) & (!g368) & (!g375)) + ((g340) & (g347) & (g382) & (g361) & (g368) & (!g375)) + ((g340) & (g347) & (g382) & (g361) & (g368) & (g375)));
	assign g1227 = (((!g340) & (!g347) & (!g382) & (!g361) & (g368) & (!g375)) + ((!g340) & (!g347) & (!g382) & (g361) & (!g368) & (!g375)) + ((!g340) & (!g347) & (!g382) & (g361) & (g368) & (g375)) + ((!g340) & (!g347) & (g382) & (!g361) & (!g368) & (g375)) + ((!g340) & (!g347) & (g382) & (!g361) & (g368) & (g375)) + ((!g340) & (!g347) & (g382) & (g361) & (g368) & (g375)) + ((!g340) & (g347) & (!g382) & (!g361) & (!g368) & (g375)) + ((!g340) & (g347) & (!g382) & (g361) & (!g368) & (g375)) + ((!g340) & (g347) & (!g382) & (g361) & (g368) & (g375)) + ((!g340) & (g347) & (g382) & (!g361) & (!g368) & (!g375)) + ((!g340) & (g347) & (g382) & (!g361) & (g368) & (!g375)) + ((!g340) & (g347) & (g382) & (g361) & (!g368) & (g375)) + ((!g340) & (g347) & (g382) & (g361) & (g368) & (g375)) + ((g340) & (!g347) & (!g382) & (!g361) & (g368) & (!g375)) + ((g340) & (!g347) & (!g382) & (g361) & (g368) & (g375)) + ((g340) & (!g347) & (g382) & (!g361) & (!g368) & (!g375)) + ((g340) & (!g347) & (g382) & (!g361) & (g368) & (g375)) + ((g340) & (!g347) & (g382) & (g361) & (!g368) & (!g375)) + ((g340) & (g347) & (!g382) & (!g361) & (g368) & (g375)) + ((g340) & (g347) & (!g382) & (g361) & (!g368) & (!g375)) + ((g340) & (g347) & (!g382) & (g361) & (!g368) & (g375)) + ((g340) & (g347) & (g382) & (!g361) & (g368) & (g375)));
	assign g1228 = (((!g1224) & (!g1225) & (!g1226) & (!g1227) & (!g389) & (!g354)) + ((!g1224) & (!g1225) & (!g1226) & (!g1227) & (!g389) & (g354)) + ((!g1224) & (!g1225) & (!g1226) & (!g1227) & (g389) & (!g354)) + ((!g1224) & (!g1225) & (!g1226) & (g1227) & (!g389) & (!g354)) + ((!g1224) & (!g1225) & (!g1226) & (g1227) & (!g389) & (g354)) + ((!g1224) & (!g1225) & (!g1226) & (g1227) & (g389) & (!g354)) + ((!g1224) & (!g1225) & (!g1226) & (g1227) & (g389) & (g354)) + ((!g1224) & (!g1225) & (g1226) & (!g1227) & (!g389) & (!g354)) + ((!g1224) & (!g1225) & (g1226) & (!g1227) & (g389) & (!g354)) + ((!g1224) & (!g1225) & (g1226) & (g1227) & (!g389) & (!g354)) + ((!g1224) & (!g1225) & (g1226) & (g1227) & (g389) & (!g354)) + ((!g1224) & (!g1225) & (g1226) & (g1227) & (g389) & (g354)) + ((!g1224) & (g1225) & (!g1226) & (!g1227) & (!g389) & (!g354)) + ((!g1224) & (g1225) & (!g1226) & (!g1227) & (!g389) & (g354)) + ((!g1224) & (g1225) & (!g1226) & (g1227) & (!g389) & (!g354)) + ((!g1224) & (g1225) & (!g1226) & (g1227) & (!g389) & (g354)) + ((!g1224) & (g1225) & (!g1226) & (g1227) & (g389) & (g354)) + ((!g1224) & (g1225) & (g1226) & (!g1227) & (!g389) & (!g354)) + ((!g1224) & (g1225) & (g1226) & (g1227) & (!g389) & (!g354)) + ((!g1224) & (g1225) & (g1226) & (g1227) & (g389) & (g354)) + ((g1224) & (!g1225) & (!g1226) & (!g1227) & (!g389) & (g354)) + ((g1224) & (!g1225) & (!g1226) & (!g1227) & (g389) & (!g354)) + ((g1224) & (!g1225) & (!g1226) & (g1227) & (!g389) & (g354)) + ((g1224) & (!g1225) & (!g1226) & (g1227) & (g389) & (!g354)) + ((g1224) & (!g1225) & (!g1226) & (g1227) & (g389) & (g354)) + ((g1224) & (!g1225) & (g1226) & (!g1227) & (g389) & (!g354)) + ((g1224) & (!g1225) & (g1226) & (g1227) & (g389) & (!g354)) + ((g1224) & (!g1225) & (g1226) & (g1227) & (g389) & (g354)) + ((g1224) & (g1225) & (!g1226) & (!g1227) & (!g389) & (g354)) + ((g1224) & (g1225) & (!g1226) & (g1227) & (!g389) & (g354)) + ((g1224) & (g1225) & (!g1226) & (g1227) & (g389) & (g354)) + ((g1224) & (g1225) & (g1226) & (g1227) & (g389) & (g354)));
	assign g1229 = (((!g439) & (!sk[70]) & (!g695) & (g951) & (!g1228)) + ((!g439) & (!sk[70]) & (!g695) & (g951) & (g1228)) + ((!g439) & (!sk[70]) & (g695) & (!g951) & (!g1228)) + ((!g439) & (!sk[70]) & (g695) & (!g951) & (g1228)) + ((!g439) & (!sk[70]) & (g695) & (g951) & (!g1228)) + ((!g439) & (!sk[70]) & (g695) & (g951) & (g1228)) + ((!g439) & (sk[70]) & (!g695) & (!g951) & (g1228)) + ((!g439) & (sk[70]) & (!g695) & (g951) & (!g1228)) + ((!g439) & (sk[70]) & (g695) & (!g951) & (!g1228)) + ((!g439) & (sk[70]) & (g695) & (g951) & (g1228)) + ((g439) & (!sk[70]) & (!g695) & (g951) & (!g1228)) + ((g439) & (!sk[70]) & (!g695) & (g951) & (g1228)) + ((g439) & (!sk[70]) & (g695) & (!g951) & (!g1228)) + ((g439) & (!sk[70]) & (g695) & (!g951) & (g1228)) + ((g439) & (!sk[70]) & (g695) & (g951) & (!g1228)) + ((g439) & (!sk[70]) & (g695) & (g951) & (g1228)) + ((g439) & (sk[70]) & (!g695) & (!g951) & (!g1228)) + ((g439) & (sk[70]) & (!g695) & (g951) & (g1228)) + ((g439) & (sk[70]) & (g695) & (!g951) & (g1228)) + ((g439) & (sk[70]) & (g695) & (g951) & (!g1228)));
	assign g1230 = (((!ld) & (!g183) & (!sk[71]) & (g1229) & (!keyx5x)) + ((!ld) & (!g183) & (!sk[71]) & (g1229) & (keyx5x)) + ((!ld) & (!g183) & (sk[71]) & (g1229) & (!keyx5x)) + ((!ld) & (!g183) & (sk[71]) & (g1229) & (keyx5x)) + ((!ld) & (g183) & (!sk[71]) & (!g1229) & (!keyx5x)) + ((!ld) & (g183) & (!sk[71]) & (!g1229) & (keyx5x)) + ((!ld) & (g183) & (!sk[71]) & (g1229) & (!keyx5x)) + ((!ld) & (g183) & (!sk[71]) & (g1229) & (keyx5x)) + ((!ld) & (g183) & (sk[71]) & (!g1229) & (!keyx5x)) + ((!ld) & (g183) & (sk[71]) & (!g1229) & (keyx5x)) + ((ld) & (!g183) & (!sk[71]) & (g1229) & (!keyx5x)) + ((ld) & (!g183) & (!sk[71]) & (g1229) & (keyx5x)) + ((ld) & (!g183) & (sk[71]) & (!g1229) & (keyx5x)) + ((ld) & (!g183) & (sk[71]) & (g1229) & (keyx5x)) + ((ld) & (g183) & (!sk[71]) & (!g1229) & (!keyx5x)) + ((ld) & (g183) & (!sk[71]) & (!g1229) & (keyx5x)) + ((ld) & (g183) & (!sk[71]) & (g1229) & (!keyx5x)) + ((ld) & (g183) & (!sk[71]) & (g1229) & (keyx5x)) + ((ld) & (g183) & (sk[71]) & (!g1229) & (keyx5x)) + ((ld) & (g183) & (sk[71]) & (g1229) & (keyx5x)));
	assign g1231 = (((!g340) & (!g389) & (!g354) & (!g361) & (!g368) & (g375)) + ((!g340) & (!g389) & (!g354) & (!g361) & (g368) & (g375)) + ((!g340) & (!g389) & (!g354) & (g361) & (!g368) & (!g375)) + ((!g340) & (!g389) & (!g354) & (g361) & (!g368) & (g375)) + ((!g340) & (!g389) & (!g354) & (g361) & (g368) & (!g375)) + ((!g340) & (!g389) & (!g354) & (g361) & (g368) & (g375)) + ((!g340) & (!g389) & (g354) & (!g361) & (!g368) & (g375)) + ((!g340) & (!g389) & (g354) & (!g361) & (g368) & (g375)) + ((!g340) & (!g389) & (g354) & (g361) & (g368) & (!g375)) + ((!g340) & (g389) & (g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (g389) & (g354) & (!g361) & (g368) & (g375)) + ((!g340) & (g389) & (g354) & (g361) & (!g368) & (g375)) + ((g340) & (!g389) & (!g354) & (!g361) & (g368) & (!g375)) + ((g340) & (!g389) & (!g354) & (g361) & (!g368) & (!g375)) + ((g340) & (!g389) & (!g354) & (g361) & (!g368) & (g375)) + ((g340) & (!g389) & (!g354) & (g361) & (g368) & (g375)) + ((g340) & (!g389) & (g354) & (!g361) & (!g368) & (g375)) + ((g340) & (!g389) & (g354) & (!g361) & (g368) & (g375)) + ((g340) & (!g389) & (g354) & (g361) & (g368) & (!g375)) + ((g340) & (!g389) & (g354) & (g361) & (g368) & (g375)) + ((g340) & (g389) & (!g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (g389) & (!g354) & (!g361) & (!g368) & (g375)) + ((g340) & (g389) & (!g354) & (!g361) & (g368) & (!g375)) + ((g340) & (g389) & (!g354) & (g361) & (!g368) & (!g375)) + ((g340) & (g389) & (g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (g389) & (g354) & (!g361) & (!g368) & (g375)) + ((g340) & (g389) & (g354) & (!g361) & (g368) & (!g375)) + ((g340) & (g389) & (g354) & (g361) & (!g368) & (g375)));
	assign g1232 = (((!g340) & (!g389) & (!g354) & (!g361) & (!g368) & (!g375)) + ((!g340) & (!g389) & (!g354) & (g361) & (g368) & (g375)) + ((!g340) & (!g389) & (g354) & (!g361) & (!g368) & (!g375)) + ((!g340) & (!g389) & (g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (!g389) & (g354) & (!g361) & (g368) & (g375)) + ((!g340) & (!g389) & (g354) & (g361) & (!g368) & (!g375)) + ((!g340) & (!g389) & (g354) & (g361) & (g368) & (g375)) + ((!g340) & (g389) & (!g354) & (!g361) & (!g368) & (!g375)) + ((!g340) & (g389) & (!g354) & (!g361) & (g368) & (g375)) + ((!g340) & (g389) & (!g354) & (g361) & (!g368) & (g375)) + ((!g340) & (g389) & (g354) & (!g361) & (!g368) & (!g375)) + ((!g340) & (g389) & (g354) & (!g361) & (g368) & (g375)) + ((!g340) & (g389) & (g354) & (g361) & (g368) & (!g375)) + ((!g340) & (g389) & (g354) & (g361) & (g368) & (g375)) + ((g340) & (!g389) & (!g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (!g389) & (!g354) & (!g361) & (g368) & (g375)) + ((g340) & (!g389) & (!g354) & (g361) & (!g368) & (!g375)) + ((g340) & (!g389) & (!g354) & (g361) & (g368) & (g375)) + ((g340) & (!g389) & (g354) & (!g361) & (g368) & (g375)) + ((g340) & (!g389) & (g354) & (g361) & (!g368) & (g375)) + ((g340) & (g389) & (!g354) & (!g361) & (g368) & (!g375)) + ((g340) & (g389) & (!g354) & (!g361) & (g368) & (g375)) + ((g340) & (g389) & (!g354) & (g361) & (!g368) & (g375)) + ((g340) & (g389) & (!g354) & (g361) & (g368) & (!g375)) + ((g340) & (g389) & (!g354) & (g361) & (g368) & (g375)) + ((g340) & (g389) & (g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (g389) & (g354) & (!g361) & (g368) & (!g375)) + ((g340) & (g389) & (g354) & (g361) & (!g368) & (!g375)));
	assign g1233 = (((!g340) & (!g389) & (!g354) & (!g361) & (!g368) & (g375)) + ((!g340) & (!g389) & (!g354) & (!g361) & (g368) & (g375)) + ((!g340) & (!g389) & (!g354) & (g361) & (g368) & (!g375)) + ((!g340) & (!g389) & (!g354) & (g361) & (g368) & (g375)) + ((!g340) & (!g389) & (g354) & (!g361) & (g368) & (g375)) + ((!g340) & (!g389) & (g354) & (g361) & (!g368) & (!g375)) + ((!g340) & (!g389) & (g354) & (g361) & (!g368) & (g375)) + ((!g340) & (!g389) & (g354) & (g361) & (g368) & (g375)) + ((!g340) & (g389) & (!g354) & (!g361) & (!g368) & (!g375)) + ((!g340) & (g389) & (!g354) & (!g361) & (!g368) & (g375)) + ((!g340) & (g389) & (!g354) & (!g361) & (g368) & (g375)) + ((!g340) & (g389) & (!g354) & (g361) & (!g368) & (g375)) + ((!g340) & (g389) & (!g354) & (g361) & (g368) & (!g375)) + ((!g340) & (g389) & (g354) & (!g361) & (!g368) & (g375)) + ((!g340) & (g389) & (g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (g389) & (g354) & (g361) & (!g368) & (!g375)) + ((!g340) & (g389) & (g354) & (g361) & (g368) & (!g375)) + ((!g340) & (g389) & (g354) & (g361) & (g368) & (g375)) + ((g340) & (!g389) & (!g354) & (!g361) & (!g368) & (g375)) + ((g340) & (!g389) & (!g354) & (g361) & (!g368) & (!g375)) + ((g340) & (!g389) & (!g354) & (g361) & (g368) & (!g375)) + ((g340) & (!g389) & (g354) & (!g361) & (g368) & (g375)) + ((g340) & (!g389) & (g354) & (g361) & (!g368) & (g375)) + ((g340) & (g389) & (!g354) & (!g361) & (!g368) & (g375)) + ((g340) & (g389) & (!g354) & (g361) & (!g368) & (!g375)) + ((g340) & (g389) & (!g354) & (g361) & (g368) & (!g375)) + ((g340) & (g389) & (g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (g389) & (g354) & (!g361) & (g368) & (!g375)) + ((g340) & (g389) & (g354) & (!g361) & (g368) & (g375)) + ((g340) & (g389) & (g354) & (g361) & (g368) & (g375)));
	assign g1234 = (((!g340) & (!g389) & (!g354) & (!g361) & (g368) & (g375)) + ((!g340) & (!g389) & (!g354) & (g361) & (!g368) & (!g375)) + ((!g340) & (!g389) & (!g354) & (g361) & (g368) & (g375)) + ((!g340) & (!g389) & (g354) & (!g361) & (!g368) & (!g375)) + ((!g340) & (!g389) & (g354) & (g361) & (g368) & (!g375)) + ((!g340) & (!g389) & (g354) & (g361) & (g368) & (g375)) + ((!g340) & (g389) & (!g354) & (g361) & (!g368) & (!g375)) + ((!g340) & (g389) & (!g354) & (g361) & (g368) & (!g375)) + ((!g340) & (g389) & (g354) & (!g361) & (g368) & (!g375)) + ((!g340) & (g389) & (g354) & (!g361) & (g368) & (g375)) + ((g340) & (!g389) & (!g354) & (!g361) & (!g368) & (g375)) + ((g340) & (!g389) & (!g354) & (!g361) & (g368) & (!g375)) + ((g340) & (!g389) & (!g354) & (g361) & (!g368) & (g375)) + ((g340) & (!g389) & (g354) & (!g361) & (g368) & (!g375)) + ((g340) & (!g389) & (g354) & (!g361) & (g368) & (g375)) + ((g340) & (!g389) & (g354) & (g361) & (g368) & (!g375)) + ((g340) & (!g389) & (g354) & (g361) & (g368) & (g375)) + ((g340) & (g389) & (!g354) & (!g361) & (g368) & (!g375)) + ((g340) & (g389) & (!g354) & (g361) & (!g368) & (g375)) + ((g340) & (g389) & (g354) & (!g361) & (!g368) & (!g375)) + ((g340) & (g389) & (g354) & (!g361) & (g368) & (g375)) + ((g340) & (g389) & (g354) & (g361) & (!g368) & (g375)));
	assign g1235 = (((!g1231) & (!g1232) & (!g1233) & (!g1234) & (!g382) & (!g347)) + ((!g1231) & (!g1232) & (!g1233) & (!g1234) & (!g382) & (g347)) + ((!g1231) & (!g1232) & (!g1233) & (!g1234) & (g382) & (!g347)) + ((!g1231) & (!g1232) & (!g1233) & (g1234) & (!g382) & (!g347)) + ((!g1231) & (!g1232) & (!g1233) & (g1234) & (!g382) & (g347)) + ((!g1231) & (!g1232) & (!g1233) & (g1234) & (g382) & (!g347)) + ((!g1231) & (!g1232) & (!g1233) & (g1234) & (g382) & (g347)) + ((!g1231) & (!g1232) & (g1233) & (!g1234) & (!g382) & (!g347)) + ((!g1231) & (!g1232) & (g1233) & (!g1234) & (g382) & (!g347)) + ((!g1231) & (!g1232) & (g1233) & (g1234) & (!g382) & (!g347)) + ((!g1231) & (!g1232) & (g1233) & (g1234) & (g382) & (!g347)) + ((!g1231) & (!g1232) & (g1233) & (g1234) & (g382) & (g347)) + ((!g1231) & (g1232) & (!g1233) & (!g1234) & (!g382) & (!g347)) + ((!g1231) & (g1232) & (!g1233) & (!g1234) & (!g382) & (g347)) + ((!g1231) & (g1232) & (!g1233) & (g1234) & (!g382) & (!g347)) + ((!g1231) & (g1232) & (!g1233) & (g1234) & (!g382) & (g347)) + ((!g1231) & (g1232) & (!g1233) & (g1234) & (g382) & (g347)) + ((!g1231) & (g1232) & (g1233) & (!g1234) & (!g382) & (!g347)) + ((!g1231) & (g1232) & (g1233) & (g1234) & (!g382) & (!g347)) + ((!g1231) & (g1232) & (g1233) & (g1234) & (g382) & (g347)) + ((g1231) & (!g1232) & (!g1233) & (!g1234) & (!g382) & (g347)) + ((g1231) & (!g1232) & (!g1233) & (!g1234) & (g382) & (!g347)) + ((g1231) & (!g1232) & (!g1233) & (g1234) & (!g382) & (g347)) + ((g1231) & (!g1232) & (!g1233) & (g1234) & (g382) & (!g347)) + ((g1231) & (!g1232) & (!g1233) & (g1234) & (g382) & (g347)) + ((g1231) & (!g1232) & (g1233) & (!g1234) & (g382) & (!g347)) + ((g1231) & (!g1232) & (g1233) & (g1234) & (g382) & (!g347)) + ((g1231) & (!g1232) & (g1233) & (g1234) & (g382) & (g347)) + ((g1231) & (g1232) & (!g1233) & (!g1234) & (!g382) & (g347)) + ((g1231) & (g1232) & (!g1233) & (g1234) & (!g382) & (g347)) + ((g1231) & (g1232) & (!g1233) & (g1234) & (g382) & (g347)) + ((g1231) & (g1232) & (g1233) & (g1234) & (g382) & (g347)));
	assign g1236 = (((!g446) & (!sk[77]) & (!g702) & (g958) & (!g1235)) + ((!g446) & (!sk[77]) & (!g702) & (g958) & (g1235)) + ((!g446) & (!sk[77]) & (g702) & (!g958) & (!g1235)) + ((!g446) & (!sk[77]) & (g702) & (!g958) & (g1235)) + ((!g446) & (!sk[77]) & (g702) & (g958) & (!g1235)) + ((!g446) & (!sk[77]) & (g702) & (g958) & (g1235)) + ((!g446) & (sk[77]) & (!g702) & (!g958) & (g1235)) + ((!g446) & (sk[77]) & (!g702) & (g958) & (!g1235)) + ((!g446) & (sk[77]) & (g702) & (!g958) & (!g1235)) + ((!g446) & (sk[77]) & (g702) & (g958) & (g1235)) + ((g446) & (!sk[77]) & (!g702) & (g958) & (!g1235)) + ((g446) & (!sk[77]) & (!g702) & (g958) & (g1235)) + ((g446) & (!sk[77]) & (g702) & (!g958) & (!g1235)) + ((g446) & (!sk[77]) & (g702) & (!g958) & (g1235)) + ((g446) & (!sk[77]) & (g702) & (g958) & (!g1235)) + ((g446) & (!sk[77]) & (g702) & (g958) & (g1235)) + ((g446) & (sk[77]) & (!g702) & (!g958) & (!g1235)) + ((g446) & (sk[77]) & (!g702) & (g958) & (g1235)) + ((g446) & (sk[77]) & (g702) & (!g958) & (g1235)) + ((g446) & (sk[77]) & (g702) & (g958) & (!g1235)));
	assign g1237 = (((!ld) & (!g190) & (g1236) & (!sk[78]) & (!keyx6x)) + ((!ld) & (!g190) & (g1236) & (!sk[78]) & (keyx6x)) + ((!ld) & (!g190) & (g1236) & (sk[78]) & (!keyx6x)) + ((!ld) & (!g190) & (g1236) & (sk[78]) & (keyx6x)) + ((!ld) & (g190) & (!g1236) & (!sk[78]) & (!keyx6x)) + ((!ld) & (g190) & (!g1236) & (!sk[78]) & (keyx6x)) + ((!ld) & (g190) & (!g1236) & (sk[78]) & (!keyx6x)) + ((!ld) & (g190) & (!g1236) & (sk[78]) & (keyx6x)) + ((!ld) & (g190) & (g1236) & (!sk[78]) & (!keyx6x)) + ((!ld) & (g190) & (g1236) & (!sk[78]) & (keyx6x)) + ((ld) & (!g190) & (!g1236) & (sk[78]) & (keyx6x)) + ((ld) & (!g190) & (g1236) & (!sk[78]) & (!keyx6x)) + ((ld) & (!g190) & (g1236) & (!sk[78]) & (keyx6x)) + ((ld) & (!g190) & (g1236) & (sk[78]) & (keyx6x)) + ((ld) & (g190) & (!g1236) & (!sk[78]) & (!keyx6x)) + ((ld) & (g190) & (!g1236) & (!sk[78]) & (keyx6x)) + ((ld) & (g190) & (!g1236) & (sk[78]) & (keyx6x)) + ((ld) & (g190) & (g1236) & (!sk[78]) & (!keyx6x)) + ((ld) & (g190) & (g1236) & (!sk[78]) & (keyx6x)) + ((ld) & (g190) & (g1236) & (sk[78]) & (keyx6x)));
	assign g1238 = (((!g382) & (!g347) & (!g354) & (!g361) & (!g368) & (g389)) + ((!g382) & (!g347) & (!g354) & (!g361) & (g368) & (!g389)) + ((!g382) & (!g347) & (!g354) & (g361) & (!g368) & (g389)) + ((!g382) & (!g347) & (!g354) & (g361) & (g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (!g361) & (!g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (!g361) & (g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (g361) & (!g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (g361) & (g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (g361) & (g368) & (g389)) + ((!g382) & (g347) & (!g354) & (!g361) & (g368) & (!g389)) + ((!g382) & (g347) & (!g354) & (g361) & (g368) & (!g389)) + ((!g382) & (g347) & (!g354) & (g361) & (g368) & (g389)) + ((!g382) & (g347) & (g354) & (!g361) & (g368) & (g389)) + ((!g382) & (g347) & (g354) & (g361) & (!g368) & (!g389)) + ((g382) & (!g347) & (!g354) & (!g361) & (!g368) & (g389)) + ((g382) & (!g347) & (!g354) & (g361) & (!g368) & (g389)) + ((g382) & (!g347) & (g354) & (g361) & (g368) & (g389)) + ((g382) & (g347) & (!g354) & (!g361) & (g368) & (g389)) + ((g382) & (g347) & (!g354) & (g361) & (!g368) & (!g389)) + ((g382) & (g347) & (!g354) & (g361) & (g368) & (!g389)) + ((g382) & (g347) & (g354) & (!g361) & (!g368) & (g389)) + ((g382) & (g347) & (g354) & (!g361) & (g368) & (!g389)) + ((g382) & (g347) & (g354) & (!g361) & (g368) & (g389)) + ((g382) & (g347) & (g354) & (g361) & (!g368) & (g389)));
	assign g1239 = (((!g382) & (!g347) & (!g354) & (!g361) & (!g368) & (!g389)) + ((!g382) & (!g347) & (!g354) & (!g361) & (!g368) & (g389)) + ((!g382) & (!g347) & (!g354) & (g361) & (!g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (!g361) & (!g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (!g361) & (g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (!g361) & (g368) & (g389)) + ((!g382) & (!g347) & (g354) & (g361) & (!g368) & (g389)) + ((!g382) & (!g347) & (g354) & (g361) & (g368) & (g389)) + ((!g382) & (g347) & (!g354) & (!g361) & (!g368) & (!g389)) + ((!g382) & (g347) & (!g354) & (!g361) & (g368) & (!g389)) + ((!g382) & (g347) & (!g354) & (g361) & (!g368) & (!g389)) + ((!g382) & (g347) & (!g354) & (g361) & (!g368) & (g389)) + ((!g382) & (g347) & (!g354) & (g361) & (g368) & (g389)) + ((!g382) & (g347) & (g354) & (!g361) & (!g368) & (g389)) + ((!g382) & (g347) & (g354) & (g361) & (!g368) & (!g389)) + ((!g382) & (g347) & (g354) & (g361) & (!g368) & (g389)) + ((g382) & (!g347) & (!g354) & (!g361) & (!g368) & (g389)) + ((g382) & (!g347) & (!g354) & (!g361) & (g368) & (g389)) + ((g382) & (!g347) & (!g354) & (g361) & (!g368) & (!g389)) + ((g382) & (!g347) & (!g354) & (g361) & (g368) & (g389)) + ((g382) & (!g347) & (g354) & (!g361) & (!g368) & (!g389)) + ((g382) & (!g347) & (g354) & (!g361) & (g368) & (g389)) + ((g382) & (!g347) & (g354) & (g361) & (g368) & (!g389)) + ((g382) & (g347) & (!g354) & (!g361) & (!g368) & (!g389)) + ((g382) & (g347) & (!g354) & (!g361) & (!g368) & (g389)) + ((g382) & (g347) & (!g354) & (!g361) & (g368) & (g389)) + ((g382) & (g347) & (!g354) & (g361) & (!g368) & (g389)) + ((g382) & (g347) & (!g354) & (g361) & (g368) & (!g389)) + ((g382) & (g347) & (g354) & (!g361) & (g368) & (!g389)) + ((g382) & (g347) & (g354) & (!g361) & (g368) & (g389)));
	assign g1240 = (((!g382) & (!g347) & (!g354) & (!g361) & (g368) & (!g389)) + ((!g382) & (!g347) & (!g354) & (g361) & (!g368) & (!g389)) + ((!g382) & (!g347) & (!g354) & (g361) & (g368) & (!g389)) + ((!g382) & (!g347) & (!g354) & (g361) & (g368) & (g389)) + ((!g382) & (!g347) & (g354) & (!g361) & (!g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (!g361) & (!g368) & (g389)) + ((!g382) & (!g347) & (g354) & (!g361) & (g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (g361) & (!g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (g361) & (g368) & (g389)) + ((!g382) & (g347) & (!g354) & (!g361) & (!g368) & (g389)) + ((!g382) & (g347) & (!g354) & (!g361) & (g368) & (!g389)) + ((!g382) & (g347) & (!g354) & (!g361) & (g368) & (g389)) + ((!g382) & (g347) & (g354) & (!g361) & (!g368) & (g389)) + ((!g382) & (g347) & (g354) & (!g361) & (g368) & (!g389)) + ((!g382) & (g347) & (g354) & (!g361) & (g368) & (g389)) + ((!g382) & (g347) & (g354) & (g361) & (!g368) & (!g389)) + ((g382) & (!g347) & (!g354) & (!g361) & (g368) & (!g389)) + ((g382) & (!g347) & (!g354) & (g361) & (!g368) & (!g389)) + ((g382) & (!g347) & (!g354) & (g361) & (g368) & (g389)) + ((g382) & (!g347) & (g354) & (!g361) & (!g368) & (!g389)) + ((g382) & (!g347) & (g354) & (!g361) & (!g368) & (g389)) + ((g382) & (!g347) & (g354) & (g361) & (!g368) & (!g389)) + ((g382) & (!g347) & (g354) & (g361) & (g368) & (!g389)) + ((g382) & (g347) & (!g354) & (!g361) & (g368) & (!g389)) + ((g382) & (g347) & (!g354) & (g361) & (!g368) & (!g389)) + ((g382) & (g347) & (!g354) & (g361) & (g368) & (g389)) + ((g382) & (g347) & (g354) & (!g361) & (!g368) & (!g389)) + ((g382) & (g347) & (g354) & (!g361) & (g368) & (!g389)) + ((g382) & (g347) & (g354) & (!g361) & (g368) & (g389)) + ((g382) & (g347) & (g354) & (g361) & (!g368) & (g389)));
	assign g1241 = (((!g382) & (!g347) & (!g354) & (!g361) & (!g368) & (g389)) + ((!g382) & (!g347) & (!g354) & (g361) & (g368) & (!g389)) + ((!g382) & (!g347) & (!g354) & (g361) & (g368) & (g389)) + ((!g382) & (!g347) & (g354) & (!g361) & (!g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (!g361) & (!g368) & (g389)) + ((!g382) & (!g347) & (g354) & (g361) & (g368) & (!g389)) + ((!g382) & (!g347) & (g354) & (g361) & (g368) & (g389)) + ((!g382) & (g347) & (!g354) & (!g361) & (!g368) & (!g389)) + ((!g382) & (g347) & (!g354) & (!g361) & (!g368) & (g389)) + ((!g382) & (g347) & (!g354) & (!g361) & (g368) & (g389)) + ((!g382) & (g347) & (!g354) & (g361) & (!g368) & (g389)) + ((!g382) & (g347) & (g354) & (!g361) & (!g368) & (g389)) + ((!g382) & (g347) & (g354) & (g361) & (!g368) & (!g389)) + ((!g382) & (g347) & (g354) & (g361) & (!g368) & (g389)) + ((!g382) & (g347) & (g354) & (g361) & (g368) & (!g389)) + ((!g382) & (g347) & (g354) & (g361) & (g368) & (g389)) + ((g382) & (!g347) & (!g354) & (g361) & (!g368) & (g389)) + ((g382) & (!g347) & (g354) & (!g361) & (!g368) & (!g389)) + ((g382) & (!g347) & (g354) & (g361) & (!g368) & (!g389)) + ((g382) & (!g347) & (g354) & (g361) & (!g368) & (g389)) + ((g382) & (!g347) & (g354) & (g361) & (g368) & (g389)) + ((g382) & (g347) & (!g354) & (!g361) & (!g368) & (g389)) + ((g382) & (g347) & (!g354) & (!g361) & (g368) & (g389)) + ((g382) & (g347) & (!g354) & (g361) & (!g368) & (!g389)) + ((g382) & (g347) & (!g354) & (g361) & (g368) & (!g389)) + ((g382) & (g347) & (!g354) & (g361) & (g368) & (g389)) + ((g382) & (g347) & (g354) & (!g361) & (g368) & (g389)) + ((g382) & (g347) & (g354) & (g361) & (g368) & (g389)));
	assign g1242 = (((!g1238) & (!g1239) & (!g1240) & (!g1241) & (!g340) & (g375)) + ((!g1238) & (!g1239) & (!g1240) & (!g1241) & (g340) & (!g375)) + ((!g1238) & (!g1239) & (!g1240) & (!g1241) & (g340) & (g375)) + ((!g1238) & (!g1239) & (!g1240) & (g1241) & (!g340) & (g375)) + ((!g1238) & (!g1239) & (!g1240) & (g1241) & (g340) & (!g375)) + ((!g1238) & (!g1239) & (g1240) & (!g1241) & (g340) & (!g375)) + ((!g1238) & (!g1239) & (g1240) & (!g1241) & (g340) & (g375)) + ((!g1238) & (!g1239) & (g1240) & (g1241) & (g340) & (!g375)) + ((!g1238) & (g1239) & (!g1240) & (!g1241) & (!g340) & (g375)) + ((!g1238) & (g1239) & (!g1240) & (!g1241) & (g340) & (g375)) + ((!g1238) & (g1239) & (!g1240) & (g1241) & (!g340) & (g375)) + ((!g1238) & (g1239) & (g1240) & (!g1241) & (g340) & (g375)) + ((g1238) & (!g1239) & (!g1240) & (!g1241) & (!g340) & (!g375)) + ((g1238) & (!g1239) & (!g1240) & (!g1241) & (!g340) & (g375)) + ((g1238) & (!g1239) & (!g1240) & (!g1241) & (g340) & (!g375)) + ((g1238) & (!g1239) & (!g1240) & (!g1241) & (g340) & (g375)) + ((g1238) & (!g1239) & (!g1240) & (g1241) & (!g340) & (!g375)) + ((g1238) & (!g1239) & (!g1240) & (g1241) & (!g340) & (g375)) + ((g1238) & (!g1239) & (!g1240) & (g1241) & (g340) & (!g375)) + ((g1238) & (!g1239) & (g1240) & (!g1241) & (!g340) & (!g375)) + ((g1238) & (!g1239) & (g1240) & (!g1241) & (g340) & (!g375)) + ((g1238) & (!g1239) & (g1240) & (!g1241) & (g340) & (g375)) + ((g1238) & (!g1239) & (g1240) & (g1241) & (!g340) & (!g375)) + ((g1238) & (!g1239) & (g1240) & (g1241) & (g340) & (!g375)) + ((g1238) & (g1239) & (!g1240) & (!g1241) & (!g340) & (!g375)) + ((g1238) & (g1239) & (!g1240) & (!g1241) & (!g340) & (g375)) + ((g1238) & (g1239) & (!g1240) & (!g1241) & (g340) & (g375)) + ((g1238) & (g1239) & (!g1240) & (g1241) & (!g340) & (!g375)) + ((g1238) & (g1239) & (!g1240) & (g1241) & (!g340) & (g375)) + ((g1238) & (g1239) & (g1240) & (!g1241) & (!g340) & (!g375)) + ((g1238) & (g1239) & (g1240) & (!g1241) & (g340) & (g375)) + ((g1238) & (g1239) & (g1240) & (g1241) & (!g340) & (!g375)));
	assign g1243 = (((!g453) & (!g709) & (!g965) & (sk[84]) & (g1242)) + ((!g453) & (!g709) & (g965) & (!sk[84]) & (!g1242)) + ((!g453) & (!g709) & (g965) & (!sk[84]) & (g1242)) + ((!g453) & (!g709) & (g965) & (sk[84]) & (!g1242)) + ((!g453) & (g709) & (!g965) & (!sk[84]) & (!g1242)) + ((!g453) & (g709) & (!g965) & (!sk[84]) & (g1242)) + ((!g453) & (g709) & (!g965) & (sk[84]) & (!g1242)) + ((!g453) & (g709) & (g965) & (!sk[84]) & (!g1242)) + ((!g453) & (g709) & (g965) & (!sk[84]) & (g1242)) + ((!g453) & (g709) & (g965) & (sk[84]) & (g1242)) + ((g453) & (!g709) & (!g965) & (sk[84]) & (!g1242)) + ((g453) & (!g709) & (g965) & (!sk[84]) & (!g1242)) + ((g453) & (!g709) & (g965) & (!sk[84]) & (g1242)) + ((g453) & (!g709) & (g965) & (sk[84]) & (g1242)) + ((g453) & (g709) & (!g965) & (!sk[84]) & (!g1242)) + ((g453) & (g709) & (!g965) & (!sk[84]) & (g1242)) + ((g453) & (g709) & (!g965) & (sk[84]) & (g1242)) + ((g453) & (g709) & (g965) & (!sk[84]) & (!g1242)) + ((g453) & (g709) & (g965) & (!sk[84]) & (g1242)) + ((g453) & (g709) & (g965) & (sk[84]) & (!g1242)));
	assign g1244 = (((!ld) & (!g197) & (!sk[85]) & (g1243) & (!keyx7x)) + ((!ld) & (!g197) & (!sk[85]) & (g1243) & (keyx7x)) + ((!ld) & (!g197) & (sk[85]) & (g1243) & (!keyx7x)) + ((!ld) & (!g197) & (sk[85]) & (g1243) & (keyx7x)) + ((!ld) & (g197) & (!sk[85]) & (!g1243) & (!keyx7x)) + ((!ld) & (g197) & (!sk[85]) & (!g1243) & (keyx7x)) + ((!ld) & (g197) & (!sk[85]) & (g1243) & (!keyx7x)) + ((!ld) & (g197) & (!sk[85]) & (g1243) & (keyx7x)) + ((!ld) & (g197) & (sk[85]) & (!g1243) & (!keyx7x)) + ((!ld) & (g197) & (sk[85]) & (!g1243) & (keyx7x)) + ((ld) & (!g197) & (!sk[85]) & (g1243) & (!keyx7x)) + ((ld) & (!g197) & (!sk[85]) & (g1243) & (keyx7x)) + ((ld) & (!g197) & (sk[85]) & (!g1243) & (keyx7x)) + ((ld) & (!g197) & (sk[85]) & (g1243) & (keyx7x)) + ((ld) & (g197) & (!sk[85]) & (!g1243) & (!keyx7x)) + ((ld) & (g197) & (!sk[85]) & (!g1243) & (keyx7x)) + ((ld) & (g197) & (!sk[85]) & (g1243) & (!keyx7x)) + ((ld) & (g197) & (!sk[85]) & (g1243) & (keyx7x)) + ((ld) & (g197) & (sk[85]) & (!g1243) & (keyx7x)) + ((ld) & (g197) & (sk[85]) & (g1243) & (keyx7x)));
	assign g2090 = (((!ld) & (!sk[86]) & (text_inx72x) & (!g1245)) + ((!ld) & (!sk[86]) & (text_inx72x) & (g1245)) + ((!ld) & (sk[86]) & (!text_inx72x) & (g1245)) + ((!ld) & (sk[86]) & (text_inx72x) & (g1245)) + ((ld) & (!sk[86]) & (!text_inx72x) & (g1245)) + ((ld) & (!sk[86]) & (text_inx72x) & (!g1245)) + ((ld) & (!sk[86]) & (text_inx72x) & (g1245)) + ((ld) & (sk[86]) & (text_inx72x) & (!g1245)) + ((ld) & (sk[86]) & (text_inx72x) & (g1245)));
	assign g1246 = (((!g708) & (!sk[87]) & (g772)) + ((!g708) & (sk[87]) & (g772)) + ((g708) & (!sk[87]) & (g772)) + ((g708) & (sk[87]) & (!g772)));
	assign g1247 = (((!sk[88]) & (!g787) & (g851)) + ((!sk[88]) & (g787) & (g851)) + ((sk[88]) & (!g787) & (g851)) + ((sk[88]) & (g787) & (!g851)));
	assign g1248 = (((!g659) & (!g724) & (!g1163) & (!g1245) & (!g1246) & (g1247)) + ((!g659) & (!g724) & (!g1163) & (!g1245) & (g1246) & (!g1247)) + ((!g659) & (!g724) & (!g1163) & (g1245) & (!g1246) & (g1247)) + ((!g659) & (!g724) & (!g1163) & (g1245) & (g1246) & (!g1247)) + ((!g659) & (!g724) & (g1163) & (g1245) & (!g1246) & (!g1247)) + ((!g659) & (!g724) & (g1163) & (g1245) & (!g1246) & (g1247)) + ((!g659) & (!g724) & (g1163) & (g1245) & (g1246) & (!g1247)) + ((!g659) & (!g724) & (g1163) & (g1245) & (g1246) & (g1247)) + ((!g659) & (g724) & (!g1163) & (!g1245) & (!g1246) & (!g1247)) + ((!g659) & (g724) & (!g1163) & (!g1245) & (g1246) & (g1247)) + ((!g659) & (g724) & (!g1163) & (g1245) & (!g1246) & (!g1247)) + ((!g659) & (g724) & (!g1163) & (g1245) & (g1246) & (g1247)) + ((!g659) & (g724) & (g1163) & (!g1245) & (!g1246) & (!g1247)) + ((!g659) & (g724) & (g1163) & (!g1245) & (!g1246) & (g1247)) + ((!g659) & (g724) & (g1163) & (!g1245) & (g1246) & (!g1247)) + ((!g659) & (g724) & (g1163) & (!g1245) & (g1246) & (g1247)) + ((g659) & (!g724) & (!g1163) & (!g1245) & (!g1246) & (!g1247)) + ((g659) & (!g724) & (!g1163) & (!g1245) & (g1246) & (g1247)) + ((g659) & (!g724) & (!g1163) & (g1245) & (!g1246) & (!g1247)) + ((g659) & (!g724) & (!g1163) & (g1245) & (g1246) & (g1247)) + ((g659) & (!g724) & (g1163) & (g1245) & (!g1246) & (!g1247)) + ((g659) & (!g724) & (g1163) & (g1245) & (!g1246) & (g1247)) + ((g659) & (!g724) & (g1163) & (g1245) & (g1246) & (!g1247)) + ((g659) & (!g724) & (g1163) & (g1245) & (g1246) & (g1247)) + ((g659) & (g724) & (!g1163) & (!g1245) & (!g1246) & (g1247)) + ((g659) & (g724) & (!g1163) & (!g1245) & (g1246) & (!g1247)) + ((g659) & (g724) & (!g1163) & (g1245) & (!g1246) & (g1247)) + ((g659) & (g724) & (!g1163) & (g1245) & (g1246) & (!g1247)) + ((g659) & (g724) & (g1163) & (!g1245) & (!g1246) & (!g1247)) + ((g659) & (g724) & (g1163) & (!g1245) & (!g1246) & (g1247)) + ((g659) & (g724) & (g1163) & (!g1245) & (g1246) & (!g1247)) + ((g659) & (g724) & (g1163) & (!g1245) & (g1246) & (g1247)));
	assign g2091 = (((!ld) & (!sk[90]) & (text_inx73x) & (!g1249)) + ((!ld) & (!sk[90]) & (text_inx73x) & (g1249)) + ((!ld) & (sk[90]) & (!text_inx73x) & (g1249)) + ((!ld) & (sk[90]) & (text_inx73x) & (g1249)) + ((ld) & (!sk[90]) & (!text_inx73x) & (g1249)) + ((ld) & (!sk[90]) & (text_inx73x) & (!g1249)) + ((ld) & (!sk[90]) & (text_inx73x) & (g1249)) + ((ld) & (sk[90]) & (text_inx73x) & (!g1249)) + ((ld) & (sk[90]) & (text_inx73x) & (g1249)));
	assign g1250 = (((!sk[91]) & (!g666) & (g858)) + ((!sk[91]) & (g666) & (g858)) + ((sk[91]) & (!g666) & (g858)) + ((sk[91]) & (g666) & (!g858)));
	assign g1251 = (((!g659) & (!g708) & (!g723) & (!g731) & (!g772) & (g794)) + ((!g659) & (!g708) & (!g723) & (!g731) & (g772) & (!g794)) + ((!g659) & (!g708) & (!g723) & (g731) & (!g772) & (!g794)) + ((!g659) & (!g708) & (!g723) & (g731) & (g772) & (g794)) + ((!g659) & (!g708) & (g723) & (!g731) & (!g772) & (!g794)) + ((!g659) & (!g708) & (g723) & (!g731) & (g772) & (g794)) + ((!g659) & (!g708) & (g723) & (g731) & (!g772) & (g794)) + ((!g659) & (!g708) & (g723) & (g731) & (g772) & (!g794)) + ((!g659) & (g708) & (!g723) & (!g731) & (!g772) & (!g794)) + ((!g659) & (g708) & (!g723) & (!g731) & (g772) & (g794)) + ((!g659) & (g708) & (!g723) & (g731) & (!g772) & (g794)) + ((!g659) & (g708) & (!g723) & (g731) & (g772) & (!g794)) + ((!g659) & (g708) & (g723) & (!g731) & (!g772) & (g794)) + ((!g659) & (g708) & (g723) & (!g731) & (g772) & (!g794)) + ((!g659) & (g708) & (g723) & (g731) & (!g772) & (!g794)) + ((!g659) & (g708) & (g723) & (g731) & (g772) & (g794)) + ((g659) & (!g708) & (!g723) & (!g731) & (!g772) & (!g794)) + ((g659) & (!g708) & (!g723) & (!g731) & (g772) & (g794)) + ((g659) & (!g708) & (!g723) & (g731) & (!g772) & (g794)) + ((g659) & (!g708) & (!g723) & (g731) & (g772) & (!g794)) + ((g659) & (!g708) & (g723) & (!g731) & (!g772) & (g794)) + ((g659) & (!g708) & (g723) & (!g731) & (g772) & (!g794)) + ((g659) & (!g708) & (g723) & (g731) & (!g772) & (!g794)) + ((g659) & (!g708) & (g723) & (g731) & (g772) & (g794)) + ((g659) & (g708) & (!g723) & (!g731) & (!g772) & (g794)) + ((g659) & (g708) & (!g723) & (!g731) & (g772) & (!g794)) + ((g659) & (g708) & (!g723) & (g731) & (!g772) & (!g794)) + ((g659) & (g708) & (!g723) & (g731) & (g772) & (g794)) + ((g659) & (g708) & (g723) & (!g731) & (!g772) & (!g794)) + ((g659) & (g708) & (g723) & (!g731) & (g772) & (g794)) + ((g659) & (g708) & (g723) & (g731) & (!g772) & (g794)) + ((g659) & (g708) & (g723) & (g731) & (g772) & (!g794)));
	assign g1252 = (((!sk[93]) & (!g731) & (g1163) & (!g1249) & (!g1250) & (!g1251)) + ((!sk[93]) & (!g731) & (g1163) & (!g1249) & (!g1250) & (g1251)) + ((!sk[93]) & (!g731) & (g1163) & (!g1249) & (g1250) & (!g1251)) + ((!sk[93]) & (!g731) & (g1163) & (!g1249) & (g1250) & (g1251)) + ((!sk[93]) & (!g731) & (g1163) & (g1249) & (!g1250) & (!g1251)) + ((!sk[93]) & (!g731) & (g1163) & (g1249) & (!g1250) & (g1251)) + ((!sk[93]) & (!g731) & (g1163) & (g1249) & (g1250) & (!g1251)) + ((!sk[93]) & (!g731) & (g1163) & (g1249) & (g1250) & (g1251)) + ((!sk[93]) & (g731) & (!g1163) & (!g1249) & (!g1250) & (!g1251)) + ((!sk[93]) & (g731) & (!g1163) & (!g1249) & (!g1250) & (g1251)) + ((!sk[93]) & (g731) & (!g1163) & (!g1249) & (g1250) & (!g1251)) + ((!sk[93]) & (g731) & (!g1163) & (!g1249) & (g1250) & (g1251)) + ((!sk[93]) & (g731) & (!g1163) & (g1249) & (!g1250) & (!g1251)) + ((!sk[93]) & (g731) & (!g1163) & (g1249) & (!g1250) & (g1251)) + ((!sk[93]) & (g731) & (!g1163) & (g1249) & (g1250) & (!g1251)) + ((!sk[93]) & (g731) & (!g1163) & (g1249) & (g1250) & (g1251)) + ((!sk[93]) & (g731) & (g1163) & (!g1249) & (!g1250) & (!g1251)) + ((!sk[93]) & (g731) & (g1163) & (!g1249) & (!g1250) & (g1251)) + ((!sk[93]) & (g731) & (g1163) & (!g1249) & (g1250) & (!g1251)) + ((!sk[93]) & (g731) & (g1163) & (!g1249) & (g1250) & (g1251)) + ((!sk[93]) & (g731) & (g1163) & (g1249) & (!g1250) & (!g1251)) + ((!sk[93]) & (g731) & (g1163) & (g1249) & (!g1250) & (g1251)) + ((!sk[93]) & (g731) & (g1163) & (g1249) & (g1250) & (!g1251)) + ((!sk[93]) & (g731) & (g1163) & (g1249) & (g1250) & (g1251)) + ((sk[93]) & (!g731) & (!g1163) & (!g1249) & (!g1250) & (g1251)) + ((sk[93]) & (!g731) & (!g1163) & (!g1249) & (g1250) & (!g1251)) + ((sk[93]) & (!g731) & (!g1163) & (g1249) & (!g1250) & (g1251)) + ((sk[93]) & (!g731) & (!g1163) & (g1249) & (g1250) & (!g1251)) + ((sk[93]) & (!g731) & (g1163) & (g1249) & (!g1250) & (!g1251)) + ((sk[93]) & (!g731) & (g1163) & (g1249) & (!g1250) & (g1251)) + ((sk[93]) & (!g731) & (g1163) & (g1249) & (g1250) & (!g1251)) + ((sk[93]) & (!g731) & (g1163) & (g1249) & (g1250) & (g1251)) + ((sk[93]) & (g731) & (!g1163) & (!g1249) & (!g1250) & (g1251)) + ((sk[93]) & (g731) & (!g1163) & (!g1249) & (g1250) & (!g1251)) + ((sk[93]) & (g731) & (!g1163) & (g1249) & (!g1250) & (g1251)) + ((sk[93]) & (g731) & (!g1163) & (g1249) & (g1250) & (!g1251)) + ((sk[93]) & (g731) & (g1163) & (!g1249) & (!g1250) & (!g1251)) + ((sk[93]) & (g731) & (g1163) & (!g1249) & (!g1250) & (g1251)) + ((sk[93]) & (g731) & (g1163) & (!g1249) & (g1250) & (!g1251)) + ((sk[93]) & (g731) & (g1163) & (!g1249) & (g1250) & (g1251)));
	assign g2092 = (((!sk[94]) & (!ld) & (text_inx74x) & (!g1253)) + ((!sk[94]) & (!ld) & (text_inx74x) & (g1253)) + ((!sk[94]) & (ld) & (!text_inx74x) & (g1253)) + ((!sk[94]) & (ld) & (text_inx74x) & (!g1253)) + ((!sk[94]) & (ld) & (text_inx74x) & (g1253)) + ((sk[94]) & (!ld) & (!text_inx74x) & (g1253)) + ((sk[94]) & (!ld) & (text_inx74x) & (g1253)) + ((sk[94]) & (ld) & (text_inx74x) & (!g1253)) + ((sk[94]) & (ld) & (text_inx74x) & (g1253)));
	assign g1254 = (((!sk[95]) & (!g666) & (g801) & (!g865)) + ((!sk[95]) & (!g666) & (g801) & (g865)) + ((!sk[95]) & (g666) & (!g801) & (g865)) + ((!sk[95]) & (g666) & (g801) & (!g865)) + ((!sk[95]) & (g666) & (g801) & (g865)) + ((sk[95]) & (!g666) & (!g801) & (g865)) + ((sk[95]) & (!g666) & (g801) & (!g865)) + ((sk[95]) & (g666) & (!g801) & (!g865)) + ((sk[95]) & (g666) & (g801) & (g865)));
	assign g1255 = (((!g673) & (!g730) & (!g738) & (!g1163) & (!g1253) & (g1254)) + ((!g673) & (!g730) & (!g738) & (!g1163) & (g1253) & (g1254)) + ((!g673) & (!g730) & (!g738) & (g1163) & (g1253) & (!g1254)) + ((!g673) & (!g730) & (!g738) & (g1163) & (g1253) & (g1254)) + ((!g673) & (!g730) & (g738) & (!g1163) & (!g1253) & (!g1254)) + ((!g673) & (!g730) & (g738) & (!g1163) & (g1253) & (!g1254)) + ((!g673) & (!g730) & (g738) & (g1163) & (!g1253) & (!g1254)) + ((!g673) & (!g730) & (g738) & (g1163) & (!g1253) & (g1254)) + ((!g673) & (g730) & (!g738) & (!g1163) & (!g1253) & (!g1254)) + ((!g673) & (g730) & (!g738) & (!g1163) & (g1253) & (!g1254)) + ((!g673) & (g730) & (!g738) & (g1163) & (g1253) & (!g1254)) + ((!g673) & (g730) & (!g738) & (g1163) & (g1253) & (g1254)) + ((!g673) & (g730) & (g738) & (!g1163) & (!g1253) & (g1254)) + ((!g673) & (g730) & (g738) & (!g1163) & (g1253) & (g1254)) + ((!g673) & (g730) & (g738) & (g1163) & (!g1253) & (!g1254)) + ((!g673) & (g730) & (g738) & (g1163) & (!g1253) & (g1254)) + ((g673) & (!g730) & (!g738) & (!g1163) & (!g1253) & (!g1254)) + ((g673) & (!g730) & (!g738) & (!g1163) & (g1253) & (!g1254)) + ((g673) & (!g730) & (!g738) & (g1163) & (g1253) & (!g1254)) + ((g673) & (!g730) & (!g738) & (g1163) & (g1253) & (g1254)) + ((g673) & (!g730) & (g738) & (!g1163) & (!g1253) & (g1254)) + ((g673) & (!g730) & (g738) & (!g1163) & (g1253) & (g1254)) + ((g673) & (!g730) & (g738) & (g1163) & (!g1253) & (!g1254)) + ((g673) & (!g730) & (g738) & (g1163) & (!g1253) & (g1254)) + ((g673) & (g730) & (!g738) & (!g1163) & (!g1253) & (g1254)) + ((g673) & (g730) & (!g738) & (!g1163) & (g1253) & (g1254)) + ((g673) & (g730) & (!g738) & (g1163) & (g1253) & (!g1254)) + ((g673) & (g730) & (!g738) & (g1163) & (g1253) & (g1254)) + ((g673) & (g730) & (g738) & (!g1163) & (!g1253) & (!g1254)) + ((g673) & (g730) & (g738) & (!g1163) & (g1253) & (!g1254)) + ((g673) & (g730) & (g738) & (g1163) & (!g1253) & (!g1254)) + ((g673) & (g730) & (g738) & (g1163) & (!g1253) & (g1254)));
	assign g2093 = (((!ld) & (!text_inx75x) & (sk[97]) & (g1256)) + ((!ld) & (text_inx75x) & (!sk[97]) & (!g1256)) + ((!ld) & (text_inx75x) & (!sk[97]) & (g1256)) + ((!ld) & (text_inx75x) & (sk[97]) & (g1256)) + ((ld) & (!text_inx75x) & (!sk[97]) & (g1256)) + ((ld) & (text_inx75x) & (!sk[97]) & (!g1256)) + ((ld) & (text_inx75x) & (!sk[97]) & (g1256)) + ((ld) & (text_inx75x) & (sk[97]) & (!g1256)) + ((ld) & (text_inx75x) & (sk[97]) & (g1256)));
	assign g1257 = (((!g673) & (!g708) & (!g737) & (!g745) & (!g772) & (g808)) + ((!g673) & (!g708) & (!g737) & (!g745) & (g772) & (!g808)) + ((!g673) & (!g708) & (!g737) & (g745) & (!g772) & (!g808)) + ((!g673) & (!g708) & (!g737) & (g745) & (g772) & (g808)) + ((!g673) & (!g708) & (g737) & (!g745) & (!g772) & (!g808)) + ((!g673) & (!g708) & (g737) & (!g745) & (g772) & (g808)) + ((!g673) & (!g708) & (g737) & (g745) & (!g772) & (g808)) + ((!g673) & (!g708) & (g737) & (g745) & (g772) & (!g808)) + ((!g673) & (g708) & (!g737) & (!g745) & (!g772) & (!g808)) + ((!g673) & (g708) & (!g737) & (!g745) & (g772) & (g808)) + ((!g673) & (g708) & (!g737) & (g745) & (!g772) & (g808)) + ((!g673) & (g708) & (!g737) & (g745) & (g772) & (!g808)) + ((!g673) & (g708) & (g737) & (!g745) & (!g772) & (g808)) + ((!g673) & (g708) & (g737) & (!g745) & (g772) & (!g808)) + ((!g673) & (g708) & (g737) & (g745) & (!g772) & (!g808)) + ((!g673) & (g708) & (g737) & (g745) & (g772) & (g808)) + ((g673) & (!g708) & (!g737) & (!g745) & (!g772) & (!g808)) + ((g673) & (!g708) & (!g737) & (!g745) & (g772) & (g808)) + ((g673) & (!g708) & (!g737) & (g745) & (!g772) & (g808)) + ((g673) & (!g708) & (!g737) & (g745) & (g772) & (!g808)) + ((g673) & (!g708) & (g737) & (!g745) & (!g772) & (g808)) + ((g673) & (!g708) & (g737) & (!g745) & (g772) & (!g808)) + ((g673) & (!g708) & (g737) & (g745) & (!g772) & (!g808)) + ((g673) & (!g708) & (g737) & (g745) & (g772) & (g808)) + ((g673) & (g708) & (!g737) & (!g745) & (!g772) & (g808)) + ((g673) & (g708) & (!g737) & (!g745) & (g772) & (!g808)) + ((g673) & (g708) & (!g737) & (g745) & (!g772) & (!g808)) + ((g673) & (g708) & (!g737) & (g745) & (g772) & (g808)) + ((g673) & (g708) & (g737) & (!g745) & (!g772) & (!g808)) + ((g673) & (g708) & (g737) & (!g745) & (g772) & (g808)) + ((g673) & (g708) & (g737) & (g745) & (!g772) & (g808)) + ((g673) & (g708) & (g737) & (g745) & (g772) & (!g808)));
	assign g1258 = (((!g680) & (!g745) & (!g872) & (!g1163) & (!g1256) & (g1257)) + ((!g680) & (!g745) & (!g872) & (!g1163) & (g1256) & (g1257)) + ((!g680) & (!g745) & (!g872) & (g1163) & (g1256) & (!g1257)) + ((!g680) & (!g745) & (!g872) & (g1163) & (g1256) & (g1257)) + ((!g680) & (!g745) & (g872) & (!g1163) & (!g1256) & (!g1257)) + ((!g680) & (!g745) & (g872) & (!g1163) & (g1256) & (!g1257)) + ((!g680) & (!g745) & (g872) & (g1163) & (g1256) & (!g1257)) + ((!g680) & (!g745) & (g872) & (g1163) & (g1256) & (g1257)) + ((!g680) & (g745) & (!g872) & (!g1163) & (!g1256) & (g1257)) + ((!g680) & (g745) & (!g872) & (!g1163) & (g1256) & (g1257)) + ((!g680) & (g745) & (!g872) & (g1163) & (!g1256) & (!g1257)) + ((!g680) & (g745) & (!g872) & (g1163) & (!g1256) & (g1257)) + ((!g680) & (g745) & (g872) & (!g1163) & (!g1256) & (!g1257)) + ((!g680) & (g745) & (g872) & (!g1163) & (g1256) & (!g1257)) + ((!g680) & (g745) & (g872) & (g1163) & (!g1256) & (!g1257)) + ((!g680) & (g745) & (g872) & (g1163) & (!g1256) & (g1257)) + ((g680) & (!g745) & (!g872) & (!g1163) & (!g1256) & (!g1257)) + ((g680) & (!g745) & (!g872) & (!g1163) & (g1256) & (!g1257)) + ((g680) & (!g745) & (!g872) & (g1163) & (g1256) & (!g1257)) + ((g680) & (!g745) & (!g872) & (g1163) & (g1256) & (g1257)) + ((g680) & (!g745) & (g872) & (!g1163) & (!g1256) & (g1257)) + ((g680) & (!g745) & (g872) & (!g1163) & (g1256) & (g1257)) + ((g680) & (!g745) & (g872) & (g1163) & (g1256) & (!g1257)) + ((g680) & (!g745) & (g872) & (g1163) & (g1256) & (g1257)) + ((g680) & (g745) & (!g872) & (!g1163) & (!g1256) & (!g1257)) + ((g680) & (g745) & (!g872) & (!g1163) & (g1256) & (!g1257)) + ((g680) & (g745) & (!g872) & (g1163) & (!g1256) & (!g1257)) + ((g680) & (g745) & (!g872) & (g1163) & (!g1256) & (g1257)) + ((g680) & (g745) & (g872) & (!g1163) & (!g1256) & (g1257)) + ((g680) & (g745) & (g872) & (!g1163) & (g1256) & (g1257)) + ((g680) & (g745) & (g872) & (g1163) & (!g1256) & (!g1257)) + ((g680) & (g745) & (g872) & (g1163) & (!g1256) & (g1257)));
	assign g2094 = (((!ld) & (!sk[100]) & (text_inx78x) & (!g1259)) + ((!ld) & (!sk[100]) & (text_inx78x) & (g1259)) + ((!ld) & (sk[100]) & (!text_inx78x) & (g1259)) + ((!ld) & (sk[100]) & (text_inx78x) & (g1259)) + ((ld) & (!sk[100]) & (!text_inx78x) & (g1259)) + ((ld) & (!sk[100]) & (text_inx78x) & (!g1259)) + ((ld) & (!sk[100]) & (text_inx78x) & (g1259)) + ((ld) & (sk[100]) & (text_inx78x) & (!g1259)) + ((ld) & (sk[100]) & (text_inx78x) & (g1259)));
	assign g1260 = (((!sk[101]) & (!g694) & (g829) & (!g893)) + ((!sk[101]) & (!g694) & (g829) & (g893)) + ((!sk[101]) & (g694) & (!g829) & (g893)) + ((!sk[101]) & (g694) & (g829) & (!g893)) + ((!sk[101]) & (g694) & (g829) & (g893)) + ((sk[101]) & (!g694) & (!g829) & (g893)) + ((sk[101]) & (!g694) & (g829) & (!g893)) + ((sk[101]) & (g694) & (!g829) & (!g893)) + ((sk[101]) & (g694) & (g829) & (g893)));
	assign g1261 = (((!g701) & (!g758) & (!g766) & (!g1163) & (!g1259) & (g1260)) + ((!g701) & (!g758) & (!g766) & (!g1163) & (g1259) & (g1260)) + ((!g701) & (!g758) & (!g766) & (g1163) & (g1259) & (!g1260)) + ((!g701) & (!g758) & (!g766) & (g1163) & (g1259) & (g1260)) + ((!g701) & (!g758) & (g766) & (!g1163) & (!g1259) & (!g1260)) + ((!g701) & (!g758) & (g766) & (!g1163) & (g1259) & (!g1260)) + ((!g701) & (!g758) & (g766) & (g1163) & (!g1259) & (!g1260)) + ((!g701) & (!g758) & (g766) & (g1163) & (!g1259) & (g1260)) + ((!g701) & (g758) & (!g766) & (!g1163) & (!g1259) & (!g1260)) + ((!g701) & (g758) & (!g766) & (!g1163) & (g1259) & (!g1260)) + ((!g701) & (g758) & (!g766) & (g1163) & (g1259) & (!g1260)) + ((!g701) & (g758) & (!g766) & (g1163) & (g1259) & (g1260)) + ((!g701) & (g758) & (g766) & (!g1163) & (!g1259) & (g1260)) + ((!g701) & (g758) & (g766) & (!g1163) & (g1259) & (g1260)) + ((!g701) & (g758) & (g766) & (g1163) & (!g1259) & (!g1260)) + ((!g701) & (g758) & (g766) & (g1163) & (!g1259) & (g1260)) + ((g701) & (!g758) & (!g766) & (!g1163) & (!g1259) & (!g1260)) + ((g701) & (!g758) & (!g766) & (!g1163) & (g1259) & (!g1260)) + ((g701) & (!g758) & (!g766) & (g1163) & (g1259) & (!g1260)) + ((g701) & (!g758) & (!g766) & (g1163) & (g1259) & (g1260)) + ((g701) & (!g758) & (g766) & (!g1163) & (!g1259) & (g1260)) + ((g701) & (!g758) & (g766) & (!g1163) & (g1259) & (g1260)) + ((g701) & (!g758) & (g766) & (g1163) & (!g1259) & (!g1260)) + ((g701) & (!g758) & (g766) & (g1163) & (!g1259) & (g1260)) + ((g701) & (g758) & (!g766) & (!g1163) & (!g1259) & (g1260)) + ((g701) & (g758) & (!g766) & (!g1163) & (g1259) & (g1260)) + ((g701) & (g758) & (!g766) & (g1163) & (g1259) & (!g1260)) + ((g701) & (g758) & (!g766) & (g1163) & (g1259) & (g1260)) + ((g701) & (g758) & (g766) & (!g1163) & (!g1259) & (!g1260)) + ((g701) & (g758) & (g766) & (!g1163) & (g1259) & (!g1260)) + ((g701) & (g758) & (g766) & (g1163) & (!g1259) & (!g1260)) + ((g701) & (g758) & (g766) & (g1163) & (!g1259) & (g1260)));
	assign g2095 = (((!sk[103]) & (!ld) & (text_inx77x) & (!g1262)) + ((!sk[103]) & (!ld) & (text_inx77x) & (g1262)) + ((!sk[103]) & (ld) & (!text_inx77x) & (g1262)) + ((!sk[103]) & (ld) & (text_inx77x) & (!g1262)) + ((!sk[103]) & (ld) & (text_inx77x) & (g1262)) + ((sk[103]) & (!ld) & (!text_inx77x) & (g1262)) + ((sk[103]) & (!ld) & (text_inx77x) & (g1262)) + ((sk[103]) & (ld) & (text_inx77x) & (!g1262)) + ((sk[103]) & (ld) & (text_inx77x) & (g1262)));
	assign g1263 = (((!sk[104]) & (!g687) & (g822) & (!g886)) + ((!sk[104]) & (!g687) & (g822) & (g886)) + ((!sk[104]) & (g687) & (!g822) & (g886)) + ((!sk[104]) & (g687) & (g822) & (!g886)) + ((!sk[104]) & (g687) & (g822) & (g886)) + ((sk[104]) & (!g687) & (!g822) & (g886)) + ((sk[104]) & (!g687) & (g822) & (!g886)) + ((sk[104]) & (g687) & (!g822) & (!g886)) + ((sk[104]) & (g687) & (g822) & (g886)));
	assign g1264 = (((!g694) & (!g751) & (!g759) & (!g1163) & (!g1262) & (g1263)) + ((!g694) & (!g751) & (!g759) & (!g1163) & (g1262) & (g1263)) + ((!g694) & (!g751) & (!g759) & (g1163) & (g1262) & (!g1263)) + ((!g694) & (!g751) & (!g759) & (g1163) & (g1262) & (g1263)) + ((!g694) & (!g751) & (g759) & (!g1163) & (!g1262) & (!g1263)) + ((!g694) & (!g751) & (g759) & (!g1163) & (g1262) & (!g1263)) + ((!g694) & (!g751) & (g759) & (g1163) & (!g1262) & (!g1263)) + ((!g694) & (!g751) & (g759) & (g1163) & (!g1262) & (g1263)) + ((!g694) & (g751) & (!g759) & (!g1163) & (!g1262) & (!g1263)) + ((!g694) & (g751) & (!g759) & (!g1163) & (g1262) & (!g1263)) + ((!g694) & (g751) & (!g759) & (g1163) & (g1262) & (!g1263)) + ((!g694) & (g751) & (!g759) & (g1163) & (g1262) & (g1263)) + ((!g694) & (g751) & (g759) & (!g1163) & (!g1262) & (g1263)) + ((!g694) & (g751) & (g759) & (!g1163) & (g1262) & (g1263)) + ((!g694) & (g751) & (g759) & (g1163) & (!g1262) & (!g1263)) + ((!g694) & (g751) & (g759) & (g1163) & (!g1262) & (g1263)) + ((g694) & (!g751) & (!g759) & (!g1163) & (!g1262) & (!g1263)) + ((g694) & (!g751) & (!g759) & (!g1163) & (g1262) & (!g1263)) + ((g694) & (!g751) & (!g759) & (g1163) & (g1262) & (!g1263)) + ((g694) & (!g751) & (!g759) & (g1163) & (g1262) & (g1263)) + ((g694) & (!g751) & (g759) & (!g1163) & (!g1262) & (g1263)) + ((g694) & (!g751) & (g759) & (!g1163) & (g1262) & (g1263)) + ((g694) & (!g751) & (g759) & (g1163) & (!g1262) & (!g1263)) + ((g694) & (!g751) & (g759) & (g1163) & (!g1262) & (g1263)) + ((g694) & (g751) & (!g759) & (!g1163) & (!g1262) & (g1263)) + ((g694) & (g751) & (!g759) & (!g1163) & (g1262) & (g1263)) + ((g694) & (g751) & (!g759) & (g1163) & (g1262) & (!g1263)) + ((g694) & (g751) & (!g759) & (g1163) & (g1262) & (g1263)) + ((g694) & (g751) & (g759) & (!g1163) & (!g1262) & (!g1263)) + ((g694) & (g751) & (g759) & (!g1163) & (g1262) & (!g1263)) + ((g694) & (g751) & (g759) & (g1163) & (!g1262) & (!g1263)) + ((g694) & (g751) & (g759) & (g1163) & (!g1262) & (g1263)));
	assign g2096 = (((!ld) & (!sk[106]) & (text_inx76x) & (!g1265)) + ((!ld) & (!sk[106]) & (text_inx76x) & (g1265)) + ((!ld) & (sk[106]) & (!text_inx76x) & (g1265)) + ((!ld) & (sk[106]) & (text_inx76x) & (g1265)) + ((ld) & (!sk[106]) & (!text_inx76x) & (g1265)) + ((ld) & (!sk[106]) & (text_inx76x) & (!g1265)) + ((ld) & (!sk[106]) & (text_inx76x) & (g1265)) + ((ld) & (sk[106]) & (text_inx76x) & (!g1265)) + ((ld) & (sk[106]) & (text_inx76x) & (g1265)));
	assign g1266 = (((!g680) & (!g687) & (!g708) & (!g744) & (!g752) & (g772)) + ((!g680) & (!g687) & (!g708) & (!g744) & (g752) & (!g772)) + ((!g680) & (!g687) & (!g708) & (g744) & (!g752) & (!g772)) + ((!g680) & (!g687) & (!g708) & (g744) & (g752) & (g772)) + ((!g680) & (!g687) & (g708) & (!g744) & (!g752) & (!g772)) + ((!g680) & (!g687) & (g708) & (!g744) & (g752) & (g772)) + ((!g680) & (!g687) & (g708) & (g744) & (!g752) & (g772)) + ((!g680) & (!g687) & (g708) & (g744) & (g752) & (!g772)) + ((!g680) & (g687) & (!g708) & (!g744) & (!g752) & (!g772)) + ((!g680) & (g687) & (!g708) & (!g744) & (g752) & (g772)) + ((!g680) & (g687) & (!g708) & (g744) & (!g752) & (g772)) + ((!g680) & (g687) & (!g708) & (g744) & (g752) & (!g772)) + ((!g680) & (g687) & (g708) & (!g744) & (!g752) & (g772)) + ((!g680) & (g687) & (g708) & (!g744) & (g752) & (!g772)) + ((!g680) & (g687) & (g708) & (g744) & (!g752) & (!g772)) + ((!g680) & (g687) & (g708) & (g744) & (g752) & (g772)) + ((g680) & (!g687) & (!g708) & (!g744) & (!g752) & (!g772)) + ((g680) & (!g687) & (!g708) & (!g744) & (g752) & (g772)) + ((g680) & (!g687) & (!g708) & (g744) & (!g752) & (g772)) + ((g680) & (!g687) & (!g708) & (g744) & (g752) & (!g772)) + ((g680) & (!g687) & (g708) & (!g744) & (!g752) & (g772)) + ((g680) & (!g687) & (g708) & (!g744) & (g752) & (!g772)) + ((g680) & (!g687) & (g708) & (g744) & (!g752) & (!g772)) + ((g680) & (!g687) & (g708) & (g744) & (g752) & (g772)) + ((g680) & (g687) & (!g708) & (!g744) & (!g752) & (g772)) + ((g680) & (g687) & (!g708) & (!g744) & (g752) & (!g772)) + ((g680) & (g687) & (!g708) & (g744) & (!g752) & (!g772)) + ((g680) & (g687) & (!g708) & (g744) & (g752) & (g772)) + ((g680) & (g687) & (g708) & (!g744) & (!g752) & (!g772)) + ((g680) & (g687) & (g708) & (!g744) & (g752) & (g772)) + ((g680) & (g687) & (g708) & (g744) & (!g752) & (g772)) + ((g680) & (g687) & (g708) & (g744) & (g752) & (!g772)));
	assign g1267 = (((!g752) & (!g815) & (!g879) & (!g1163) & (!g1265) & (g1266)) + ((!g752) & (!g815) & (!g879) & (!g1163) & (g1265) & (g1266)) + ((!g752) & (!g815) & (!g879) & (g1163) & (g1265) & (!g1266)) + ((!g752) & (!g815) & (!g879) & (g1163) & (g1265) & (g1266)) + ((!g752) & (!g815) & (g879) & (!g1163) & (!g1265) & (!g1266)) + ((!g752) & (!g815) & (g879) & (!g1163) & (g1265) & (!g1266)) + ((!g752) & (!g815) & (g879) & (g1163) & (g1265) & (!g1266)) + ((!g752) & (!g815) & (g879) & (g1163) & (g1265) & (g1266)) + ((!g752) & (g815) & (!g879) & (!g1163) & (!g1265) & (!g1266)) + ((!g752) & (g815) & (!g879) & (!g1163) & (g1265) & (!g1266)) + ((!g752) & (g815) & (!g879) & (g1163) & (g1265) & (!g1266)) + ((!g752) & (g815) & (!g879) & (g1163) & (g1265) & (g1266)) + ((!g752) & (g815) & (g879) & (!g1163) & (!g1265) & (g1266)) + ((!g752) & (g815) & (g879) & (!g1163) & (g1265) & (g1266)) + ((!g752) & (g815) & (g879) & (g1163) & (g1265) & (!g1266)) + ((!g752) & (g815) & (g879) & (g1163) & (g1265) & (g1266)) + ((g752) & (!g815) & (!g879) & (!g1163) & (!g1265) & (g1266)) + ((g752) & (!g815) & (!g879) & (!g1163) & (g1265) & (g1266)) + ((g752) & (!g815) & (!g879) & (g1163) & (!g1265) & (!g1266)) + ((g752) & (!g815) & (!g879) & (g1163) & (!g1265) & (g1266)) + ((g752) & (!g815) & (g879) & (!g1163) & (!g1265) & (!g1266)) + ((g752) & (!g815) & (g879) & (!g1163) & (g1265) & (!g1266)) + ((g752) & (!g815) & (g879) & (g1163) & (!g1265) & (!g1266)) + ((g752) & (!g815) & (g879) & (g1163) & (!g1265) & (g1266)) + ((g752) & (g815) & (!g879) & (!g1163) & (!g1265) & (!g1266)) + ((g752) & (g815) & (!g879) & (!g1163) & (g1265) & (!g1266)) + ((g752) & (g815) & (!g879) & (g1163) & (!g1265) & (!g1266)) + ((g752) & (g815) & (!g879) & (g1163) & (!g1265) & (g1266)) + ((g752) & (g815) & (g879) & (!g1163) & (!g1265) & (g1266)) + ((g752) & (g815) & (g879) & (!g1163) & (g1265) & (g1266)) + ((g752) & (g815) & (g879) & (g1163) & (!g1265) & (!g1266)) + ((g752) & (g815) & (g879) & (g1163) & (!g1265) & (g1266)));
	assign g2097 = (((!ld) & (!sk[109]) & (text_inx79x) & (!g1268)) + ((!ld) & (!sk[109]) & (text_inx79x) & (g1268)) + ((!ld) & (sk[109]) & (!text_inx79x) & (g1268)) + ((!ld) & (sk[109]) & (text_inx79x) & (g1268)) + ((ld) & (!sk[109]) & (!text_inx79x) & (g1268)) + ((ld) & (!sk[109]) & (text_inx79x) & (!g1268)) + ((ld) & (!sk[109]) & (text_inx79x) & (g1268)) + ((ld) & (sk[109]) & (text_inx79x) & (!g1268)) + ((ld) & (sk[109]) & (text_inx79x) & (g1268)));
	assign g1269 = (((!sk[110]) & (!g708) & (g900)) + ((!sk[110]) & (g708) & (g900)) + ((sk[110]) & (!g708) & (g900)) + ((sk[110]) & (g708) & (!g900)));
	assign g1270 = (((!g701) & (!sk[111]) & (g765)) + ((!g701) & (sk[111]) & (g765)) + ((g701) & (!sk[111]) & (g765)) + ((g701) & (sk[111]) & (!g765)));
	assign g1271 = (((!g773) & (!g836) & (!g1163) & (!g1268) & (!g1269) & (g1270)) + ((!g773) & (!g836) & (!g1163) & (!g1268) & (g1269) & (!g1270)) + ((!g773) & (!g836) & (!g1163) & (g1268) & (!g1269) & (g1270)) + ((!g773) & (!g836) & (!g1163) & (g1268) & (g1269) & (!g1270)) + ((!g773) & (!g836) & (g1163) & (g1268) & (!g1269) & (!g1270)) + ((!g773) & (!g836) & (g1163) & (g1268) & (!g1269) & (g1270)) + ((!g773) & (!g836) & (g1163) & (g1268) & (g1269) & (!g1270)) + ((!g773) & (!g836) & (g1163) & (g1268) & (g1269) & (g1270)) + ((!g773) & (g836) & (!g1163) & (!g1268) & (!g1269) & (!g1270)) + ((!g773) & (g836) & (!g1163) & (!g1268) & (g1269) & (g1270)) + ((!g773) & (g836) & (!g1163) & (g1268) & (!g1269) & (!g1270)) + ((!g773) & (g836) & (!g1163) & (g1268) & (g1269) & (g1270)) + ((!g773) & (g836) & (g1163) & (g1268) & (!g1269) & (!g1270)) + ((!g773) & (g836) & (g1163) & (g1268) & (!g1269) & (g1270)) + ((!g773) & (g836) & (g1163) & (g1268) & (g1269) & (!g1270)) + ((!g773) & (g836) & (g1163) & (g1268) & (g1269) & (g1270)) + ((g773) & (!g836) & (!g1163) & (!g1268) & (!g1269) & (!g1270)) + ((g773) & (!g836) & (!g1163) & (!g1268) & (g1269) & (g1270)) + ((g773) & (!g836) & (!g1163) & (g1268) & (!g1269) & (!g1270)) + ((g773) & (!g836) & (!g1163) & (g1268) & (g1269) & (g1270)) + ((g773) & (!g836) & (g1163) & (!g1268) & (!g1269) & (!g1270)) + ((g773) & (!g836) & (g1163) & (!g1268) & (!g1269) & (g1270)) + ((g773) & (!g836) & (g1163) & (!g1268) & (g1269) & (!g1270)) + ((g773) & (!g836) & (g1163) & (!g1268) & (g1269) & (g1270)) + ((g773) & (g836) & (!g1163) & (!g1268) & (!g1269) & (g1270)) + ((g773) & (g836) & (!g1163) & (!g1268) & (g1269) & (!g1270)) + ((g773) & (g836) & (!g1163) & (g1268) & (!g1269) & (g1270)) + ((g773) & (g836) & (!g1163) & (g1268) & (g1269) & (!g1270)) + ((g773) & (g836) & (g1163) & (!g1268) & (!g1269) & (!g1270)) + ((g773) & (g836) & (g1163) & (!g1268) & (!g1269) & (g1270)) + ((g773) & (g836) & (g1163) & (!g1268) & (g1269) & (!g1270)) + ((g773) & (g836) & (g1163) & (!g1268) & (g1269) & (g1270)));
	assign g1272 = (((!g148) & (!g155) & (!g162) & (!g169) & (g190) & (g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g190) & (!g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g190) & (g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (g190) & (!g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (!g190) & (!g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (!g190) & (g183)) + ((!g148) & (!g155) & (g162) & (g169) & (!g190) & (!g183)) + ((!g148) & (!g155) & (g162) & (g169) & (g190) & (g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (g190) & (!g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (g190) & (g183)) + ((!g148) & (g155) & (!g162) & (g169) & (g190) & (!g183)) + ((!g148) & (g155) & (!g162) & (g169) & (g190) & (g183)) + ((!g148) & (g155) & (g162) & (!g169) & (g190) & (!g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (!g190) & (!g183)) + ((g148) & (!g155) & (g162) & (!g169) & (g190) & (!g183)) + ((g148) & (!g155) & (g162) & (g169) & (!g190) & (g183)) + ((g148) & (!g155) & (g162) & (g169) & (g190) & (g183)) + ((g148) & (g155) & (!g162) & (!g169) & (!g190) & (g183)) + ((g148) & (g155) & (!g162) & (!g169) & (g190) & (!g183)) + ((g148) & (g155) & (g162) & (!g169) & (!g190) & (g183)) + ((g148) & (g155) & (g162) & (!g169) & (g190) & (!g183)) + ((g148) & (g155) & (g162) & (g169) & (!g190) & (!g183)) + ((g148) & (g155) & (g162) & (g169) & (g190) & (!g183)) + ((g148) & (g155) & (g162) & (g169) & (g190) & (g183)));
	assign g1273 = (((!g148) & (!g155) & (!g162) & (!g169) & (g190) & (!g183)) + ((!g148) & (!g155) & (!g162) & (!g169) & (g190) & (g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g190) & (!g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g190) & (g183)) + ((!g148) & (!g155) & (g162) & (g169) & (!g190) & (g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (!g190) & (!g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (!g190) & (g183)) + ((!g148) & (g155) & (g162) & (!g169) & (!g190) & (!g183)) + ((!g148) & (g155) & (g162) & (!g169) & (!g190) & (g183)) + ((!g148) & (g155) & (g162) & (!g169) & (g190) & (!g183)) + ((!g148) & (g155) & (g162) & (g169) & (g190) & (g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (!g190) & (g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (g190) & (!g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (g190) & (g183)) + ((g148) & (!g155) & (!g162) & (g169) & (g190) & (!g183)) + ((g148) & (!g155) & (g162) & (!g169) & (!g190) & (!g183)) + ((g148) & (!g155) & (g162) & (!g169) & (g190) & (g183)) + ((g148) & (!g155) & (g162) & (g169) & (!g190) & (g183)) + ((g148) & (!g155) & (g162) & (g169) & (g190) & (g183)) + ((g148) & (g155) & (!g162) & (!g169) & (!g190) & (!g183)) + ((g148) & (g155) & (!g162) & (!g169) & (!g190) & (g183)) + ((g148) & (g155) & (!g162) & (!g169) & (g190) & (!g183)) + ((g148) & (g155) & (!g162) & (!g169) & (g190) & (g183)) + ((g148) & (g155) & (!g162) & (g169) & (!g190) & (!g183)) + ((g148) & (g155) & (!g162) & (g169) & (g190) & (!g183)) + ((g148) & (g155) & (!g162) & (g169) & (g190) & (g183)) + ((g148) & (g155) & (g162) & (!g169) & (g190) & (!g183)) + ((g148) & (g155) & (g162) & (!g169) & (g190) & (g183)) + ((g148) & (g155) & (g162) & (g169) & (!g190) & (g183)) + ((g148) & (g155) & (g162) & (g169) & (g190) & (!g183)));
	assign g1274 = (((!g148) & (!g155) & (!g162) & (!g169) & (!g190) & (!g183)) + ((!g148) & (!g155) & (!g162) & (!g169) & (g190) & (g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (g190) & (g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (!g190) & (!g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (!g190) & (g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (g190) & (g183)) + ((!g148) & (!g155) & (g162) & (g169) & (!g190) & (g183)) + ((!g148) & (!g155) & (g162) & (g169) & (g190) & (!g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (!g190) & (!g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (g190) & (!g183)) + ((!g148) & (g155) & (!g162) & (g169) & (g190) & (g183)) + ((!g148) & (g155) & (g162) & (g169) & (!g190) & (!g183)) + ((!g148) & (g155) & (g162) & (g169) & (g190) & (!g183)) + ((g148) & (!g155) & (!g162) & (g169) & (!g190) & (!g183)) + ((g148) & (!g155) & (!g162) & (g169) & (!g190) & (g183)) + ((g148) & (!g155) & (!g162) & (g169) & (g190) & (!g183)) + ((g148) & (!g155) & (g162) & (!g169) & (!g190) & (!g183)) + ((g148) & (!g155) & (g162) & (!g169) & (g190) & (g183)) + ((g148) & (!g155) & (g162) & (g169) & (!g190) & (!g183)) + ((g148) & (!g155) & (g162) & (g169) & (!g190) & (g183)) + ((g148) & (!g155) & (g162) & (g169) & (g190) & (!g183)) + ((g148) & (!g155) & (g162) & (g169) & (g190) & (g183)) + ((g148) & (g155) & (!g162) & (!g169) & (g190) & (g183)) + ((g148) & (g155) & (!g162) & (g169) & (!g190) & (!g183)) + ((g148) & (g155) & (!g162) & (g169) & (g190) & (!g183)) + ((g148) & (g155) & (!g162) & (g169) & (g190) & (g183)) + ((g148) & (g155) & (g162) & (!g169) & (!g190) & (!g183)) + ((g148) & (g155) & (g162) & (g169) & (!g190) & (!g183)) + ((g148) & (g155) & (g162) & (g169) & (!g190) & (g183)) + ((g148) & (g155) & (g162) & (g169) & (g190) & (g183)));
	assign g1275 = (((!g148) & (!g155) & (!g162) & (!g169) & (!g190) & (g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (g190) & (!g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (g190) & (g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (!g190) & (g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (g190) & (g183)) + ((!g148) & (!g155) & (g162) & (g169) & (!g190) & (g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (!g190) & (!g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (!g190) & (g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (g190) & (!g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (g190) & (g183)) + ((!g148) & (g155) & (!g162) & (g169) & (g190) & (!g183)) + ((!g148) & (g155) & (!g162) & (g169) & (g190) & (g183)) + ((!g148) & (g155) & (g162) & (g169) & (!g190) & (!g183)) + ((!g148) & (g155) & (g162) & (g169) & (g190) & (!g183)) + ((!g148) & (g155) & (g162) & (g169) & (g190) & (g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (!g190) & (!g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (g190) & (g183)) + ((g148) & (!g155) & (!g162) & (g169) & (g190) & (!g183)) + ((g148) & (!g155) & (!g162) & (g169) & (g190) & (g183)) + ((g148) & (!g155) & (g162) & (!g169) & (!g190) & (g183)) + ((g148) & (!g155) & (g162) & (!g169) & (g190) & (!g183)) + ((g148) & (!g155) & (g162) & (g169) & (g190) & (!g183)) + ((g148) & (g155) & (!g162) & (!g169) & (!g190) & (g183)) + ((g148) & (g155) & (!g162) & (!g169) & (g190) & (g183)) + ((g148) & (g155) & (!g162) & (g169) & (g190) & (!g183)) + ((g148) & (g155) & (!g162) & (g169) & (g190) & (g183)) + ((g148) & (g155) & (g162) & (!g169) & (!g190) & (g183)) + ((g148) & (g155) & (g162) & (g169) & (!g190) & (!g183)));
	assign g1276 = (((!g1272) & (!g1273) & (!g1274) & (!g1275) & (!g176) & (!g197)) + ((!g1272) & (!g1273) & (!g1274) & (g1275) & (!g176) & (!g197)) + ((!g1272) & (!g1273) & (!g1274) & (g1275) & (g176) & (g197)) + ((!g1272) & (!g1273) & (g1274) & (!g1275) & (!g176) & (!g197)) + ((!g1272) & (!g1273) & (g1274) & (!g1275) & (!g176) & (g197)) + ((!g1272) & (!g1273) & (g1274) & (g1275) & (!g176) & (!g197)) + ((!g1272) & (!g1273) & (g1274) & (g1275) & (!g176) & (g197)) + ((!g1272) & (!g1273) & (g1274) & (g1275) & (g176) & (g197)) + ((!g1272) & (g1273) & (!g1274) & (!g1275) & (!g176) & (!g197)) + ((!g1272) & (g1273) & (!g1274) & (!g1275) & (g176) & (!g197)) + ((!g1272) & (g1273) & (!g1274) & (g1275) & (!g176) & (!g197)) + ((!g1272) & (g1273) & (!g1274) & (g1275) & (g176) & (!g197)) + ((!g1272) & (g1273) & (!g1274) & (g1275) & (g176) & (g197)) + ((!g1272) & (g1273) & (g1274) & (!g1275) & (!g176) & (!g197)) + ((!g1272) & (g1273) & (g1274) & (!g1275) & (!g176) & (g197)) + ((!g1272) & (g1273) & (g1274) & (!g1275) & (g176) & (!g197)) + ((!g1272) & (g1273) & (g1274) & (g1275) & (!g176) & (!g197)) + ((!g1272) & (g1273) & (g1274) & (g1275) & (!g176) & (g197)) + ((!g1272) & (g1273) & (g1274) & (g1275) & (g176) & (!g197)) + ((!g1272) & (g1273) & (g1274) & (g1275) & (g176) & (g197)) + ((g1272) & (!g1273) & (!g1274) & (g1275) & (g176) & (g197)) + ((g1272) & (!g1273) & (g1274) & (!g1275) & (!g176) & (g197)) + ((g1272) & (!g1273) & (g1274) & (g1275) & (!g176) & (g197)) + ((g1272) & (!g1273) & (g1274) & (g1275) & (g176) & (g197)) + ((g1272) & (g1273) & (!g1274) & (!g1275) & (g176) & (!g197)) + ((g1272) & (g1273) & (!g1274) & (g1275) & (g176) & (!g197)) + ((g1272) & (g1273) & (!g1274) & (g1275) & (g176) & (g197)) + ((g1272) & (g1273) & (g1274) & (!g1275) & (!g176) & (g197)) + ((g1272) & (g1273) & (g1274) & (!g1275) & (g176) & (!g197)) + ((g1272) & (g1273) & (g1274) & (g1275) & (!g176) & (g197)) + ((g1272) & (g1273) & (g1274) & (g1275) & (g176) & (!g197)) + ((g1272) & (g1273) & (g1274) & (g1275) & (g176) & (g197)));
	assign g1277 = (((!sk[118]) & (!g468) & (!g724) & (g980) & (!g1276)) + ((!sk[118]) & (!g468) & (!g724) & (g980) & (g1276)) + ((!sk[118]) & (!g468) & (g724) & (!g980) & (!g1276)) + ((!sk[118]) & (!g468) & (g724) & (!g980) & (g1276)) + ((!sk[118]) & (!g468) & (g724) & (g980) & (!g1276)) + ((!sk[118]) & (!g468) & (g724) & (g980) & (g1276)) + ((!sk[118]) & (g468) & (!g724) & (g980) & (!g1276)) + ((!sk[118]) & (g468) & (!g724) & (g980) & (g1276)) + ((!sk[118]) & (g468) & (g724) & (!g980) & (!g1276)) + ((!sk[118]) & (g468) & (g724) & (!g980) & (g1276)) + ((!sk[118]) & (g468) & (g724) & (g980) & (!g1276)) + ((!sk[118]) & (g468) & (g724) & (g980) & (g1276)) + ((sk[118]) & (!g468) & (!g724) & (!g980) & (g1276)) + ((sk[118]) & (!g468) & (!g724) & (g980) & (!g1276)) + ((sk[118]) & (!g468) & (g724) & (!g980) & (!g1276)) + ((sk[118]) & (!g468) & (g724) & (g980) & (g1276)) + ((sk[118]) & (g468) & (!g724) & (!g980) & (!g1276)) + ((sk[118]) & (g468) & (!g724) & (g980) & (g1276)) + ((sk[118]) & (g468) & (g724) & (!g980) & (g1276)) + ((sk[118]) & (g468) & (g724) & (g980) & (!g1276)));
	assign g1278 = (((!sk[119]) & (!ld) & (!g212) & (g1277) & (!keyx8x)) + ((!sk[119]) & (!ld) & (!g212) & (g1277) & (keyx8x)) + ((!sk[119]) & (!ld) & (g212) & (!g1277) & (!keyx8x)) + ((!sk[119]) & (!ld) & (g212) & (!g1277) & (keyx8x)) + ((!sk[119]) & (!ld) & (g212) & (g1277) & (!keyx8x)) + ((!sk[119]) & (!ld) & (g212) & (g1277) & (keyx8x)) + ((!sk[119]) & (ld) & (!g212) & (g1277) & (!keyx8x)) + ((!sk[119]) & (ld) & (!g212) & (g1277) & (keyx8x)) + ((!sk[119]) & (ld) & (g212) & (!g1277) & (!keyx8x)) + ((!sk[119]) & (ld) & (g212) & (!g1277) & (keyx8x)) + ((!sk[119]) & (ld) & (g212) & (g1277) & (!keyx8x)) + ((!sk[119]) & (ld) & (g212) & (g1277) & (keyx8x)) + ((sk[119]) & (!ld) & (!g212) & (g1277) & (!keyx8x)) + ((sk[119]) & (!ld) & (!g212) & (g1277) & (keyx8x)) + ((sk[119]) & (!ld) & (g212) & (!g1277) & (!keyx8x)) + ((sk[119]) & (!ld) & (g212) & (!g1277) & (keyx8x)) + ((sk[119]) & (ld) & (!g212) & (!g1277) & (keyx8x)) + ((sk[119]) & (ld) & (!g212) & (g1277) & (keyx8x)) + ((sk[119]) & (ld) & (g212) & (!g1277) & (keyx8x)) + ((sk[119]) & (ld) & (g212) & (g1277) & (keyx8x)));
	assign g1279 = (((!g148) & (!g155) & (!g162) & (!g169) & (!g176) & (g190)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g176) & (!g190)) + ((!g148) & (!g155) & (!g162) & (g169) & (g176) & (!g190)) + ((!g148) & (!g155) & (g162) & (!g169) & (g176) & (g190)) + ((!g148) & (!g155) & (g162) & (g169) & (!g176) & (g190)) + ((!g148) & (!g155) & (g162) & (g169) & (g176) & (!g190)) + ((!g148) & (g155) & (!g162) & (!g169) & (!g176) & (g190)) + ((!g148) & (g155) & (!g162) & (!g169) & (g176) & (!g190)) + ((!g148) & (g155) & (!g162) & (!g169) & (g176) & (g190)) + ((!g148) & (g155) & (g162) & (!g169) & (g176) & (g190)) + ((!g148) & (g155) & (g162) & (g169) & (g176) & (g190)) + ((g148) & (!g155) & (!g162) & (!g169) & (!g176) & (!g190)) + ((g148) & (!g155) & (!g162) & (!g169) & (g176) & (g190)) + ((g148) & (!g155) & (!g162) & (g169) & (!g176) & (!g190)) + ((g148) & (!g155) & (!g162) & (g169) & (g176) & (!g190)) + ((g148) & (!g155) & (g162) & (!g169) & (g176) & (!g190)) + ((g148) & (!g155) & (g162) & (!g169) & (g176) & (g190)) + ((g148) & (!g155) & (g162) & (g169) & (g176) & (!g190)) + ((g148) & (!g155) & (g162) & (g169) & (g176) & (g190)) + ((g148) & (g155) & (!g162) & (!g169) & (g176) & (!g190)) + ((g148) & (g155) & (!g162) & (!g169) & (g176) & (g190)) + ((g148) & (g155) & (!g162) & (g169) & (g176) & (g190)) + ((g148) & (g155) & (g162) & (!g169) & (!g176) & (!g190)) + ((g148) & (g155) & (g162) & (!g169) & (!g176) & (g190)) + ((g148) & (g155) & (g162) & (!g169) & (g176) & (!g190)) + ((g148) & (g155) & (g162) & (g169) & (!g176) & (g190)) + ((g148) & (g155) & (g162) & (g169) & (g176) & (!g190)));
	assign g1280 = (((!g148) & (!g155) & (!g162) & (!g169) & (!g176) & (g190)) + ((!g148) & (!g155) & (!g162) & (!g169) & (g176) & (!g190)) + ((!g148) & (!g155) & (!g162) & (!g169) & (g176) & (g190)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g176) & (!g190)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g176) & (g190)) + ((!g148) & (!g155) & (!g162) & (g169) & (g176) & (g190)) + ((!g148) & (!g155) & (g162) & (!g169) & (g176) & (!g190)) + ((!g148) & (!g155) & (g162) & (g169) & (!g176) & (!g190)) + ((!g148) & (!g155) & (g162) & (g169) & (!g176) & (g190)) + ((!g148) & (!g155) & (g162) & (g169) & (g176) & (g190)) + ((!g148) & (g155) & (!g162) & (!g169) & (g176) & (g190)) + ((!g148) & (g155) & (!g162) & (g169) & (!g176) & (!g190)) + ((!g148) & (g155) & (!g162) & (g169) & (g176) & (!g190)) + ((!g148) & (g155) & (g162) & (!g169) & (g176) & (!g190)) + ((!g148) & (g155) & (g162) & (!g169) & (g176) & (g190)) + ((!g148) & (g155) & (g162) & (g169) & (!g176) & (!g190)) + ((g148) & (!g155) & (!g162) & (!g169) & (!g176) & (!g190)) + ((g148) & (!g155) & (!g162) & (g169) & (!g176) & (!g190)) + ((g148) & (!g155) & (!g162) & (g169) & (!g176) & (g190)) + ((g148) & (!g155) & (g162) & (!g169) & (!g176) & (g190)) + ((g148) & (!g155) & (g162) & (!g169) & (g176) & (g190)) + ((g148) & (!g155) & (g162) & (g169) & (!g176) & (!g190)) + ((g148) & (!g155) & (g162) & (g169) & (!g176) & (g190)) + ((g148) & (g155) & (!g162) & (g169) & (!g176) & (!g190)) + ((g148) & (g155) & (!g162) & (g169) & (g176) & (g190)) + ((g148) & (g155) & (g162) & (!g169) & (!g176) & (!g190)) + ((g148) & (g155) & (g162) & (!g169) & (!g176) & (g190)) + ((g148) & (g155) & (g162) & (!g169) & (g176) & (g190)) + ((g148) & (g155) & (g162) & (g169) & (!g176) & (!g190)) + ((g148) & (g155) & (g162) & (g169) & (!g176) & (g190)) + ((g148) & (g155) & (g162) & (g169) & (g176) & (!g190)));
	assign g1281 = (((!g148) & (!g155) & (!g162) & (!g169) & (!g176) & (g190)) + ((!g148) & (!g155) & (!g162) & (g169) & (g176) & (!g190)) + ((!g148) & (!g155) & (g162) & (!g169) & (!g176) & (!g190)) + ((!g148) & (!g155) & (g162) & (!g169) & (g176) & (!g190)) + ((!g148) & (!g155) & (g162) & (g169) & (!g176) & (g190)) + ((!g148) & (!g155) & (g162) & (g169) & (g176) & (!g190)) + ((!g148) & (!g155) & (g162) & (g169) & (g176) & (g190)) + ((!g148) & (g155) & (!g162) & (!g169) & (!g176) & (!g190)) + ((!g148) & (g155) & (!g162) & (!g169) & (g176) & (!g190)) + ((!g148) & (g155) & (!g162) & (g169) & (!g176) & (!g190)) + ((!g148) & (g155) & (!g162) & (g169) & (g176) & (g190)) + ((!g148) & (g155) & (g162) & (!g169) & (g176) & (g190)) + ((!g148) & (g155) & (g162) & (g169) & (!g176) & (g190)) + ((!g148) & (g155) & (g162) & (g169) & (g176) & (!g190)) + ((g148) & (!g155) & (!g162) & (!g169) & (g176) & (g190)) + ((g148) & (!g155) & (!g162) & (g169) & (!g176) & (!g190)) + ((g148) & (!g155) & (!g162) & (g169) & (g176) & (!g190)) + ((g148) & (!g155) & (g162) & (!g169) & (!g176) & (!g190)) + ((g148) & (!g155) & (g162) & (!g169) & (!g176) & (g190)) + ((g148) & (!g155) & (g162) & (!g169) & (g176) & (!g190)) + ((g148) & (!g155) & (g162) & (!g169) & (g176) & (g190)) + ((g148) & (!g155) & (g162) & (g169) & (g176) & (!g190)) + ((g148) & (g155) & (!g162) & (!g169) & (!g176) & (g190)) + ((g148) & (g155) & (!g162) & (!g169) & (g176) & (g190)) + ((g148) & (g155) & (!g162) & (g169) & (!g176) & (g190)) + ((g148) & (g155) & (g162) & (!g169) & (!g176) & (!g190)) + ((g148) & (g155) & (g162) & (!g169) & (!g176) & (g190)) + ((g148) & (g155) & (g162) & (!g169) & (g176) & (g190)) + ((g148) & (g155) & (g162) & (g169) & (!g176) & (!g190)) + ((g148) & (g155) & (g162) & (g169) & (!g176) & (g190)) + ((g148) & (g155) & (g162) & (g169) & (g176) & (!g190)) + ((g148) & (g155) & (g162) & (g169) & (g176) & (g190)));
	assign g1282 = (((!g148) & (!g155) & (!g162) & (!g169) & (g176) & (!g190)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g176) & (!g190)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g176) & (g190)) + ((!g148) & (!g155) & (g162) & (!g169) & (g176) & (g190)) + ((!g148) & (!g155) & (g162) & (g169) & (!g176) & (g190)) + ((!g148) & (g155) & (!g162) & (!g169) & (!g176) & (!g190)) + ((!g148) & (g155) & (!g162) & (!g169) & (g176) & (!g190)) + ((!g148) & (g155) & (!g162) & (g169) & (!g176) & (g190)) + ((!g148) & (g155) & (g162) & (!g169) & (!g176) & (g190)) + ((!g148) & (g155) & (g162) & (!g169) & (g176) & (!g190)) + ((!g148) & (g155) & (g162) & (!g169) & (g176) & (g190)) + ((!g148) & (g155) & (g162) & (g169) & (g176) & (!g190)) + ((!g148) & (g155) & (g162) & (g169) & (g176) & (g190)) + ((g148) & (!g155) & (!g162) & (!g169) & (!g176) & (!g190)) + ((g148) & (!g155) & (!g162) & (g169) & (!g176) & (!g190)) + ((g148) & (!g155) & (!g162) & (g169) & (!g176) & (g190)) + ((g148) & (!g155) & (!g162) & (g169) & (g176) & (!g190)) + ((g148) & (!g155) & (g162) & (!g169) & (!g176) & (!g190)) + ((g148) & (!g155) & (g162) & (!g169) & (g176) & (g190)) + ((g148) & (!g155) & (g162) & (g169) & (g176) & (!g190)) + ((g148) & (g155) & (!g162) & (!g169) & (!g176) & (!g190)) + ((g148) & (g155) & (!g162) & (g169) & (!g176) & (!g190)) + ((g148) & (g155) & (!g162) & (g169) & (g176) & (!g190)) + ((g148) & (g155) & (!g162) & (g169) & (g176) & (g190)) + ((g148) & (g155) & (g162) & (g169) & (!g176) & (g190)) + ((g148) & (g155) & (g162) & (g169) & (g176) & (g190)));
	assign g1283 = (((!g1279) & (!g1280) & (!g1281) & (!g1282) & (!g183) & (!g197)) + ((!g1279) & (!g1280) & (!g1281) & (!g1282) & (g183) & (!g197)) + ((!g1279) & (!g1280) & (!g1281) & (g1282) & (!g183) & (!g197)) + ((!g1279) & (!g1280) & (!g1281) & (g1282) & (g183) & (!g197)) + ((!g1279) & (!g1280) & (!g1281) & (g1282) & (g183) & (g197)) + ((!g1279) & (!g1280) & (g1281) & (!g1282) & (!g183) & (!g197)) + ((!g1279) & (!g1280) & (g1281) & (!g1282) & (!g183) & (g197)) + ((!g1279) & (!g1280) & (g1281) & (!g1282) & (g183) & (!g197)) + ((!g1279) & (!g1280) & (g1281) & (g1282) & (!g183) & (!g197)) + ((!g1279) & (!g1280) & (g1281) & (g1282) & (!g183) & (g197)) + ((!g1279) & (!g1280) & (g1281) & (g1282) & (g183) & (!g197)) + ((!g1279) & (!g1280) & (g1281) & (g1282) & (g183) & (g197)) + ((!g1279) & (g1280) & (!g1281) & (!g1282) & (!g183) & (!g197)) + ((!g1279) & (g1280) & (!g1281) & (g1282) & (!g183) & (!g197)) + ((!g1279) & (g1280) & (!g1281) & (g1282) & (g183) & (g197)) + ((!g1279) & (g1280) & (g1281) & (!g1282) & (!g183) & (!g197)) + ((!g1279) & (g1280) & (g1281) & (!g1282) & (!g183) & (g197)) + ((!g1279) & (g1280) & (g1281) & (g1282) & (!g183) & (!g197)) + ((!g1279) & (g1280) & (g1281) & (g1282) & (!g183) & (g197)) + ((!g1279) & (g1280) & (g1281) & (g1282) & (g183) & (g197)) + ((g1279) & (!g1280) & (!g1281) & (!g1282) & (g183) & (!g197)) + ((g1279) & (!g1280) & (!g1281) & (g1282) & (g183) & (!g197)) + ((g1279) & (!g1280) & (!g1281) & (g1282) & (g183) & (g197)) + ((g1279) & (!g1280) & (g1281) & (!g1282) & (!g183) & (g197)) + ((g1279) & (!g1280) & (g1281) & (!g1282) & (g183) & (!g197)) + ((g1279) & (!g1280) & (g1281) & (g1282) & (!g183) & (g197)) + ((g1279) & (!g1280) & (g1281) & (g1282) & (g183) & (!g197)) + ((g1279) & (!g1280) & (g1281) & (g1282) & (g183) & (g197)) + ((g1279) & (g1280) & (!g1281) & (g1282) & (g183) & (g197)) + ((g1279) & (g1280) & (g1281) & (!g1282) & (!g183) & (g197)) + ((g1279) & (g1280) & (g1281) & (g1282) & (!g183) & (g197)) + ((g1279) & (g1280) & (g1281) & (g1282) & (g183) & (g197)));
	assign g1284 = (((!g475) & (!g731) & (!sk[125]) & (g987) & (!g1283)) + ((!g475) & (!g731) & (!sk[125]) & (g987) & (g1283)) + ((!g475) & (!g731) & (sk[125]) & (!g987) & (g1283)) + ((!g475) & (!g731) & (sk[125]) & (g987) & (!g1283)) + ((!g475) & (g731) & (!sk[125]) & (!g987) & (!g1283)) + ((!g475) & (g731) & (!sk[125]) & (!g987) & (g1283)) + ((!g475) & (g731) & (!sk[125]) & (g987) & (!g1283)) + ((!g475) & (g731) & (!sk[125]) & (g987) & (g1283)) + ((!g475) & (g731) & (sk[125]) & (!g987) & (!g1283)) + ((!g475) & (g731) & (sk[125]) & (g987) & (g1283)) + ((g475) & (!g731) & (!sk[125]) & (g987) & (!g1283)) + ((g475) & (!g731) & (!sk[125]) & (g987) & (g1283)) + ((g475) & (!g731) & (sk[125]) & (!g987) & (!g1283)) + ((g475) & (!g731) & (sk[125]) & (g987) & (g1283)) + ((g475) & (g731) & (!sk[125]) & (!g987) & (!g1283)) + ((g475) & (g731) & (!sk[125]) & (!g987) & (g1283)) + ((g475) & (g731) & (!sk[125]) & (g987) & (!g1283)) + ((g475) & (g731) & (!sk[125]) & (g987) & (g1283)) + ((g475) & (g731) & (sk[125]) & (!g987) & (g1283)) + ((g475) & (g731) & (sk[125]) & (g987) & (!g1283)));
	assign g1285 = (((!ld) & (!sk[126]) & (!g219) & (g1284) & (!keyx9x)) + ((!ld) & (!sk[126]) & (!g219) & (g1284) & (keyx9x)) + ((!ld) & (!sk[126]) & (g219) & (!g1284) & (!keyx9x)) + ((!ld) & (!sk[126]) & (g219) & (!g1284) & (keyx9x)) + ((!ld) & (!sk[126]) & (g219) & (g1284) & (!keyx9x)) + ((!ld) & (!sk[126]) & (g219) & (g1284) & (keyx9x)) + ((!ld) & (sk[126]) & (!g219) & (g1284) & (!keyx9x)) + ((!ld) & (sk[126]) & (!g219) & (g1284) & (keyx9x)) + ((!ld) & (sk[126]) & (g219) & (!g1284) & (!keyx9x)) + ((!ld) & (sk[126]) & (g219) & (!g1284) & (keyx9x)) + ((ld) & (!sk[126]) & (!g219) & (g1284) & (!keyx9x)) + ((ld) & (!sk[126]) & (!g219) & (g1284) & (keyx9x)) + ((ld) & (!sk[126]) & (g219) & (!g1284) & (!keyx9x)) + ((ld) & (!sk[126]) & (g219) & (!g1284) & (keyx9x)) + ((ld) & (!sk[126]) & (g219) & (g1284) & (!keyx9x)) + ((ld) & (!sk[126]) & (g219) & (g1284) & (keyx9x)) + ((ld) & (sk[126]) & (!g219) & (!g1284) & (keyx9x)) + ((ld) & (sk[126]) & (!g219) & (g1284) & (keyx9x)) + ((ld) & (sk[126]) & (g219) & (!g1284) & (keyx9x)) + ((ld) & (sk[126]) & (g219) & (g1284) & (keyx9x)));
	assign g1286 = (((!g190) & (!g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((!g190) & (!g155) & (!g162) & (!g169) & (g176) & (g183)) + ((!g190) & (!g155) & (!g162) & (g169) & (!g176) & (g183)) + ((!g190) & (!g155) & (!g162) & (g169) & (g176) & (!g183)) + ((!g190) & (!g155) & (!g162) & (g169) & (g176) & (g183)) + ((!g190) & (!g155) & (g162) & (!g169) & (!g176) & (g183)) + ((!g190) & (!g155) & (g162) & (g169) & (!g176) & (!g183)) + ((!g190) & (!g155) & (g162) & (g169) & (g176) & (!g183)) + ((!g190) & (g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((!g190) & (g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((!g190) & (g155) & (!g162) & (g169) & (!g176) & (g183)) + ((!g190) & (g155) & (g162) & (!g169) & (!g176) & (!g183)) + ((!g190) & (g155) & (g162) & (!g169) & (!g176) & (g183)) + ((!g190) & (g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g190) & (g155) & (g162) & (!g169) & (g176) & (g183)) + ((g190) & (!g155) & (!g162) & (g169) & (!g176) & (g183)) + ((g190) & (!g155) & (!g162) & (g169) & (g176) & (g183)) + ((g190) & (g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((g190) & (g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((g190) & (g155) & (!g162) & (g169) & (g176) & (!g183)) + ((g190) & (g155) & (g162) & (g169) & (!g176) & (!g183)) + ((g190) & (g155) & (g162) & (g169) & (!g176) & (g183)));
	assign g1287 = (((!g190) & (!g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((!g190) & (!g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((!g190) & (!g155) & (!g162) & (g169) & (g176) & (g183)) + ((!g190) & (!g155) & (g162) & (!g169) & (!g176) & (!g183)) + ((!g190) & (!g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g190) & (!g155) & (g162) & (g169) & (!g176) & (g183)) + ((!g190) & (g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((!g190) & (g155) & (!g162) & (!g169) & (g176) & (g183)) + ((!g190) & (g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((!g190) & (g155) & (!g162) & (g169) & (!g176) & (g183)) + ((!g190) & (g155) & (!g162) & (g169) & (g176) & (g183)) + ((!g190) & (g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g190) & (g155) & (g162) & (!g169) & (g176) & (g183)) + ((!g190) & (g155) & (g162) & (g169) & (g176) & (!g183)) + ((g190) & (!g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((g190) & (!g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((g190) & (!g155) & (!g162) & (!g169) & (g176) & (g183)) + ((g190) & (!g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((g190) & (!g155) & (!g162) & (g169) & (!g176) & (g183)) + ((g190) & (!g155) & (!g162) & (g169) & (g176) & (!g183)) + ((g190) & (!g155) & (g162) & (g169) & (!g176) & (!g183)) + ((g190) & (g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((g190) & (g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((g190) & (g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((g190) & (g155) & (!g162) & (g169) & (g176) & (!g183)) + ((g190) & (g155) & (!g162) & (g169) & (g176) & (g183)) + ((g190) & (g155) & (g162) & (!g169) & (!g176) & (!g183)) + ((g190) & (g155) & (g162) & (!g169) & (g176) & (!g183)) + ((g190) & (g155) & (g162) & (g169) & (!g176) & (g183)) + ((g190) & (g155) & (g162) & (g169) & (g176) & (g183)));
	assign g1288 = (((!g190) & (!g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((!g190) & (!g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((!g190) & (!g155) & (!g162) & (g169) & (!g176) & (g183)) + ((!g190) & (!g155) & (g162) & (!g169) & (!g176) & (g183)) + ((!g190) & (!g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g190) & (!g155) & (g162) & (g169) & (!g176) & (g183)) + ((!g190) & (g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((!g190) & (g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((!g190) & (g155) & (!g162) & (g169) & (g176) & (!g183)) + ((!g190) & (g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g190) & (g155) & (g162) & (g169) & (!g176) & (!g183)) + ((!g190) & (g155) & (g162) & (g169) & (g176) & (!g183)) + ((g190) & (!g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((g190) & (!g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((g190) & (!g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((g190) & (!g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((g190) & (!g155) & (!g162) & (g169) & (!g176) & (g183)) + ((g190) & (!g155) & (!g162) & (g169) & (g176) & (!g183)) + ((g190) & (!g155) & (!g162) & (g169) & (g176) & (g183)) + ((g190) & (!g155) & (g162) & (!g169) & (!g176) & (g183)) + ((g190) & (!g155) & (g162) & (!g169) & (g176) & (!g183)) + ((g190) & (!g155) & (g162) & (g169) & (!g176) & (!g183)) + ((g190) & (!g155) & (g162) & (g169) & (g176) & (g183)) + ((g190) & (g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((g190) & (g155) & (!g162) & (!g169) & (g176) & (g183)) + ((g190) & (g155) & (g162) & (!g169) & (g176) & (g183)) + ((g190) & (g155) & (g162) & (g169) & (!g176) & (!g183)) + ((g190) & (g155) & (g162) & (g169) & (!g176) & (g183)) + ((g190) & (g155) & (g162) & (g169) & (g176) & (g183)));
	assign g1289 = (((!g190) & (!g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((!g190) & (!g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((!g190) & (!g155) & (!g162) & (!g169) & (g176) & (g183)) + ((!g190) & (!g155) & (!g162) & (g169) & (!g176) & (g183)) + ((!g190) & (!g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g190) & (!g155) & (g162) & (g169) & (g176) & (g183)) + ((!g190) & (g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((!g190) & (g155) & (!g162) & (g169) & (!g176) & (g183)) + ((!g190) & (g155) & (!g162) & (g169) & (g176) & (g183)) + ((!g190) & (g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g190) & (g155) & (g162) & (!g169) & (g176) & (g183)) + ((!g190) & (g155) & (g162) & (g169) & (!g176) & (!g183)) + ((!g190) & (g155) & (g162) & (g169) & (!g176) & (g183)) + ((!g190) & (g155) & (g162) & (g169) & (g176) & (!g183)) + ((!g190) & (g155) & (g162) & (g169) & (g176) & (g183)) + ((g190) & (!g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((g190) & (!g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((g190) & (!g155) & (!g162) & (!g169) & (g176) & (g183)) + ((g190) & (!g155) & (!g162) & (g169) & (g176) & (g183)) + ((g190) & (!g155) & (g162) & (!g169) & (!g176) & (g183)) + ((g190) & (!g155) & (g162) & (!g169) & (g176) & (!g183)) + ((g190) & (!g155) & (g162) & (g169) & (g176) & (!g183)) + ((g190) & (g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((g190) & (g155) & (!g162) & (g169) & (!g176) & (g183)) + ((g190) & (g155) & (!g162) & (g169) & (g176) & (!g183)) + ((g190) & (g155) & (g162) & (!g169) & (g176) & (g183)) + ((g190) & (g155) & (g162) & (g169) & (!g176) & (!g183)));
	assign g1290 = (((!g1286) & (!g1287) & (!g1288) & (!g1289) & (!g148) & (g197)) + ((!g1286) & (!g1287) & (!g1288) & (!g1289) & (g148) & (!g197)) + ((!g1286) & (!g1287) & (!g1288) & (!g1289) & (g148) & (g197)) + ((!g1286) & (!g1287) & (!g1288) & (g1289) & (!g148) & (g197)) + ((!g1286) & (!g1287) & (!g1288) & (g1289) & (g148) & (!g197)) + ((!g1286) & (!g1287) & (g1288) & (!g1289) & (g148) & (!g197)) + ((!g1286) & (!g1287) & (g1288) & (!g1289) & (g148) & (g197)) + ((!g1286) & (!g1287) & (g1288) & (g1289) & (g148) & (!g197)) + ((!g1286) & (g1287) & (!g1288) & (!g1289) & (!g148) & (g197)) + ((!g1286) & (g1287) & (!g1288) & (!g1289) & (g148) & (g197)) + ((!g1286) & (g1287) & (!g1288) & (g1289) & (!g148) & (g197)) + ((!g1286) & (g1287) & (g1288) & (!g1289) & (g148) & (g197)) + ((g1286) & (!g1287) & (!g1288) & (!g1289) & (!g148) & (!g197)) + ((g1286) & (!g1287) & (!g1288) & (!g1289) & (!g148) & (g197)) + ((g1286) & (!g1287) & (!g1288) & (!g1289) & (g148) & (!g197)) + ((g1286) & (!g1287) & (!g1288) & (!g1289) & (g148) & (g197)) + ((g1286) & (!g1287) & (!g1288) & (g1289) & (!g148) & (!g197)) + ((g1286) & (!g1287) & (!g1288) & (g1289) & (!g148) & (g197)) + ((g1286) & (!g1287) & (!g1288) & (g1289) & (g148) & (!g197)) + ((g1286) & (!g1287) & (g1288) & (!g1289) & (!g148) & (!g197)) + ((g1286) & (!g1287) & (g1288) & (!g1289) & (g148) & (!g197)) + ((g1286) & (!g1287) & (g1288) & (!g1289) & (g148) & (g197)) + ((g1286) & (!g1287) & (g1288) & (g1289) & (!g148) & (!g197)) + ((g1286) & (!g1287) & (g1288) & (g1289) & (g148) & (!g197)) + ((g1286) & (g1287) & (!g1288) & (!g1289) & (!g148) & (!g197)) + ((g1286) & (g1287) & (!g1288) & (!g1289) & (!g148) & (g197)) + ((g1286) & (g1287) & (!g1288) & (!g1289) & (g148) & (g197)) + ((g1286) & (g1287) & (!g1288) & (g1289) & (!g148) & (!g197)) + ((g1286) & (g1287) & (!g1288) & (g1289) & (!g148) & (g197)) + ((g1286) & (g1287) & (g1288) & (!g1289) & (!g148) & (!g197)) + ((g1286) & (g1287) & (g1288) & (!g1289) & (g148) & (g197)) + ((g1286) & (g1287) & (g1288) & (g1289) & (!g148) & (!g197)));
	assign g1291 = (((!g482) & (!sk[4]) & (!g738) & (g994) & (!g1290)) + ((!g482) & (!sk[4]) & (!g738) & (g994) & (g1290)) + ((!g482) & (!sk[4]) & (g738) & (!g994) & (!g1290)) + ((!g482) & (!sk[4]) & (g738) & (!g994) & (g1290)) + ((!g482) & (!sk[4]) & (g738) & (g994) & (!g1290)) + ((!g482) & (!sk[4]) & (g738) & (g994) & (g1290)) + ((!g482) & (sk[4]) & (!g738) & (!g994) & (g1290)) + ((!g482) & (sk[4]) & (!g738) & (g994) & (!g1290)) + ((!g482) & (sk[4]) & (g738) & (!g994) & (!g1290)) + ((!g482) & (sk[4]) & (g738) & (g994) & (g1290)) + ((g482) & (!sk[4]) & (!g738) & (g994) & (!g1290)) + ((g482) & (!sk[4]) & (!g738) & (g994) & (g1290)) + ((g482) & (!sk[4]) & (g738) & (!g994) & (!g1290)) + ((g482) & (!sk[4]) & (g738) & (!g994) & (g1290)) + ((g482) & (!sk[4]) & (g738) & (g994) & (!g1290)) + ((g482) & (!sk[4]) & (g738) & (g994) & (g1290)) + ((g482) & (sk[4]) & (!g738) & (!g994) & (!g1290)) + ((g482) & (sk[4]) & (!g738) & (g994) & (g1290)) + ((g482) & (sk[4]) & (g738) & (!g994) & (g1290)) + ((g482) & (sk[4]) & (g738) & (g994) & (!g1290)));
	assign g1292 = (((!ld) & (!sk[5]) & (!g226) & (g1291) & (!keyx10x)) + ((!ld) & (!sk[5]) & (!g226) & (g1291) & (keyx10x)) + ((!ld) & (!sk[5]) & (g226) & (!g1291) & (!keyx10x)) + ((!ld) & (!sk[5]) & (g226) & (!g1291) & (keyx10x)) + ((!ld) & (!sk[5]) & (g226) & (g1291) & (!keyx10x)) + ((!ld) & (!sk[5]) & (g226) & (g1291) & (keyx10x)) + ((!ld) & (sk[5]) & (!g226) & (g1291) & (!keyx10x)) + ((!ld) & (sk[5]) & (!g226) & (g1291) & (keyx10x)) + ((!ld) & (sk[5]) & (g226) & (!g1291) & (!keyx10x)) + ((!ld) & (sk[5]) & (g226) & (!g1291) & (keyx10x)) + ((ld) & (!sk[5]) & (!g226) & (g1291) & (!keyx10x)) + ((ld) & (!sk[5]) & (!g226) & (g1291) & (keyx10x)) + ((ld) & (!sk[5]) & (g226) & (!g1291) & (!keyx10x)) + ((ld) & (!sk[5]) & (g226) & (!g1291) & (keyx10x)) + ((ld) & (!sk[5]) & (g226) & (g1291) & (!keyx10x)) + ((ld) & (!sk[5]) & (g226) & (g1291) & (keyx10x)) + ((ld) & (sk[5]) & (!g226) & (!g1291) & (keyx10x)) + ((ld) & (sk[5]) & (!g226) & (g1291) & (keyx10x)) + ((ld) & (sk[5]) & (g226) & (!g1291) & (keyx10x)) + ((ld) & (sk[5]) & (g226) & (g1291) & (keyx10x)));
	assign g1293 = (((!g148) & (!g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (g176) & (g183)) + ((!g148) & (!g155) & (g162) & (g169) & (!g176) & (!g183)) + ((!g148) & (!g155) & (g162) & (g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (g162) & (g169) & (g176) & (g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (g155) & (g162) & (!g169) & (!g176) & (!g183)) + ((!g148) & (g155) & (g162) & (g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((g148) & (!g155) & (g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (g162) & (!g169) & (!g176) & (g183)) + ((g148) & (!g155) & (g162) & (!g169) & (g176) & (!g183)) + ((g148) & (!g155) & (g162) & (g169) & (!g176) & (g183)) + ((g148) & (g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((g148) & (g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((g148) & (g155) & (!g162) & (g169) & (g176) & (!g183)) + ((g148) & (g155) & (g162) & (!g169) & (!g176) & (g183)) + ((g148) & (g155) & (g162) & (!g169) & (g176) & (g183)));
	assign g1294 = (((!g148) & (!g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (!g162) & (!g169) & (g176) & (g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (g162) & (g169) & (!g176) & (!g183)) + ((!g148) & (!g155) & (g162) & (g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (g162) & (g169) & (g176) & (g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (g176) & (g183)) + ((!g148) & (g155) & (!g162) & (g169) & (g176) & (g183)) + ((!g148) & (g155) & (g162) & (!g169) & (!g176) & (!g183)) + ((!g148) & (g155) & (g162) & (!g169) & (!g176) & (g183)) + ((!g148) & (g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (g155) & (g162) & (g169) & (!g176) & (g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((g148) & (!g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (!g162) & (g169) & (!g176) & (g183)) + ((g148) & (!g155) & (!g162) & (g169) & (g176) & (g183)) + ((g148) & (!g155) & (g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (g162) & (!g169) & (!g176) & (g183)) + ((g148) & (!g155) & (g162) & (!g169) & (g176) & (g183)) + ((g148) & (!g155) & (g162) & (g169) & (!g176) & (g183)) + ((g148) & (g155) & (!g162) & (g169) & (!g176) & (g183)) + ((g148) & (g155) & (!g162) & (g169) & (g176) & (!g183)) + ((g148) & (g155) & (g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (g155) & (g162) & (g169) & (!g176) & (!g183)));
	assign g1295 = (((!g148) & (!g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (!g162) & (!g169) & (g176) & (g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (g162) & (!g169) & (g176) & (g183)) + ((!g148) & (!g155) & (g162) & (g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (g162) & (g169) & (g176) & (g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (g176) & (g183)) + ((!g148) & (g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((!g148) & (g155) & (!g162) & (g169) & (!g176) & (g183)) + ((!g148) & (g155) & (g162) & (!g169) & (!g176) & (g183)) + ((!g148) & (g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (g155) & (g162) & (g169) & (g176) & (g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (g176) & (g183)) + ((g148) & (!g155) & (!g162) & (g169) & (g176) & (g183)) + ((g148) & (!g155) & (g162) & (g169) & (!g176) & (!g183)) + ((g148) & (g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((g148) & (g155) & (!g162) & (g169) & (g176) & (g183)) + ((g148) & (g155) & (g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (g155) & (g162) & (!g169) & (!g176) & (g183)) + ((g148) & (g155) & (g162) & (!g169) & (g176) & (g183)) + ((g148) & (g155) & (g162) & (g169) & (!g176) & (!g183)) + ((g148) & (g155) & (g162) & (g169) & (g176) & (g183)));
	assign g1296 = (((!g148) & (!g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (!g162) & (g169) & (g176) & (g183)) + ((!g148) & (!g155) & (g162) & (g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (g162) & (g169) & (g176) & (g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (!g176) & (!g183)) + ((!g148) & (g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (g155) & (!g162) & (g169) & (!g176) & (!g183)) + ((!g148) & (g155) & (!g162) & (g169) & (!g176) & (g183)) + ((!g148) & (g155) & (!g162) & (g169) & (g176) & (!g183)) + ((!g148) & (g155) & (g162) & (!g169) & (!g176) & (!g183)) + ((!g148) & (g155) & (g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (g155) & (g162) & (!g169) & (g176) & (g183)) + ((g148) & (!g155) & (!g162) & (!g169) & (g176) & (g183)) + ((g148) & (!g155) & (!g162) & (g169) & (g176) & (!g183)) + ((g148) & (!g155) & (g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (g162) & (!g169) & (g176) & (!g183)) + ((g148) & (!g155) & (g162) & (!g169) & (g176) & (g183)) + ((g148) & (!g155) & (g162) & (g169) & (!g176) & (g183)) + ((g148) & (!g155) & (g162) & (g169) & (g176) & (!g183)) + ((g148) & (!g155) & (g162) & (g169) & (g176) & (g183)) + ((g148) & (g155) & (!g162) & (!g169) & (!g176) & (g183)) + ((g148) & (g155) & (!g162) & (!g169) & (g176) & (!g183)) + ((g148) & (g155) & (g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (g155) & (g162) & (!g169) & (!g176) & (g183)) + ((g148) & (g155) & (g162) & (g169) & (g176) & (g183)));
	assign g1297 = (((!g1293) & (!g1294) & (!g1295) & (!g1296) & (!g197) & (g190)) + ((!g1293) & (!g1294) & (!g1295) & (!g1296) & (g197) & (!g190)) + ((!g1293) & (!g1294) & (!g1295) & (!g1296) & (g197) & (g190)) + ((!g1293) & (!g1294) & (!g1295) & (g1296) & (!g197) & (g190)) + ((!g1293) & (!g1294) & (!g1295) & (g1296) & (g197) & (!g190)) + ((!g1293) & (!g1294) & (g1295) & (!g1296) & (g197) & (!g190)) + ((!g1293) & (!g1294) & (g1295) & (!g1296) & (g197) & (g190)) + ((!g1293) & (!g1294) & (g1295) & (g1296) & (g197) & (!g190)) + ((!g1293) & (g1294) & (!g1295) & (!g1296) & (!g197) & (g190)) + ((!g1293) & (g1294) & (!g1295) & (!g1296) & (g197) & (g190)) + ((!g1293) & (g1294) & (!g1295) & (g1296) & (!g197) & (g190)) + ((!g1293) & (g1294) & (g1295) & (!g1296) & (g197) & (g190)) + ((g1293) & (!g1294) & (!g1295) & (!g1296) & (!g197) & (!g190)) + ((g1293) & (!g1294) & (!g1295) & (!g1296) & (!g197) & (g190)) + ((g1293) & (!g1294) & (!g1295) & (!g1296) & (g197) & (!g190)) + ((g1293) & (!g1294) & (!g1295) & (!g1296) & (g197) & (g190)) + ((g1293) & (!g1294) & (!g1295) & (g1296) & (!g197) & (!g190)) + ((g1293) & (!g1294) & (!g1295) & (g1296) & (!g197) & (g190)) + ((g1293) & (!g1294) & (!g1295) & (g1296) & (g197) & (!g190)) + ((g1293) & (!g1294) & (g1295) & (!g1296) & (!g197) & (!g190)) + ((g1293) & (!g1294) & (g1295) & (!g1296) & (g197) & (!g190)) + ((g1293) & (!g1294) & (g1295) & (!g1296) & (g197) & (g190)) + ((g1293) & (!g1294) & (g1295) & (g1296) & (!g197) & (!g190)) + ((g1293) & (!g1294) & (g1295) & (g1296) & (g197) & (!g190)) + ((g1293) & (g1294) & (!g1295) & (!g1296) & (!g197) & (!g190)) + ((g1293) & (g1294) & (!g1295) & (!g1296) & (!g197) & (g190)) + ((g1293) & (g1294) & (!g1295) & (!g1296) & (g197) & (g190)) + ((g1293) & (g1294) & (!g1295) & (g1296) & (!g197) & (!g190)) + ((g1293) & (g1294) & (!g1295) & (g1296) & (!g197) & (g190)) + ((g1293) & (g1294) & (g1295) & (!g1296) & (!g197) & (!g190)) + ((g1293) & (g1294) & (g1295) & (!g1296) & (g197) & (g190)) + ((g1293) & (g1294) & (g1295) & (g1296) & (!g197) & (!g190)));
	assign g1298 = (((!g489) & (!g745) & (!sk[11]) & (g1001) & (!g1297)) + ((!g489) & (!g745) & (!sk[11]) & (g1001) & (g1297)) + ((!g489) & (!g745) & (sk[11]) & (!g1001) & (g1297)) + ((!g489) & (!g745) & (sk[11]) & (g1001) & (!g1297)) + ((!g489) & (g745) & (!sk[11]) & (!g1001) & (!g1297)) + ((!g489) & (g745) & (!sk[11]) & (!g1001) & (g1297)) + ((!g489) & (g745) & (!sk[11]) & (g1001) & (!g1297)) + ((!g489) & (g745) & (!sk[11]) & (g1001) & (g1297)) + ((!g489) & (g745) & (sk[11]) & (!g1001) & (!g1297)) + ((!g489) & (g745) & (sk[11]) & (g1001) & (g1297)) + ((g489) & (!g745) & (!sk[11]) & (g1001) & (!g1297)) + ((g489) & (!g745) & (!sk[11]) & (g1001) & (g1297)) + ((g489) & (!g745) & (sk[11]) & (!g1001) & (!g1297)) + ((g489) & (!g745) & (sk[11]) & (g1001) & (g1297)) + ((g489) & (g745) & (!sk[11]) & (!g1001) & (!g1297)) + ((g489) & (g745) & (!sk[11]) & (!g1001) & (g1297)) + ((g489) & (g745) & (!sk[11]) & (g1001) & (!g1297)) + ((g489) & (g745) & (!sk[11]) & (g1001) & (g1297)) + ((g489) & (g745) & (sk[11]) & (!g1001) & (g1297)) + ((g489) & (g745) & (sk[11]) & (g1001) & (!g1297)));
	assign g1299 = (((!ld) & (!sk[12]) & (!g233) & (g1298) & (!keyx11x)) + ((!ld) & (!sk[12]) & (!g233) & (g1298) & (keyx11x)) + ((!ld) & (!sk[12]) & (g233) & (!g1298) & (!keyx11x)) + ((!ld) & (!sk[12]) & (g233) & (!g1298) & (keyx11x)) + ((!ld) & (!sk[12]) & (g233) & (g1298) & (!keyx11x)) + ((!ld) & (!sk[12]) & (g233) & (g1298) & (keyx11x)) + ((!ld) & (sk[12]) & (!g233) & (g1298) & (!keyx11x)) + ((!ld) & (sk[12]) & (!g233) & (g1298) & (keyx11x)) + ((!ld) & (sk[12]) & (g233) & (!g1298) & (!keyx11x)) + ((!ld) & (sk[12]) & (g233) & (!g1298) & (keyx11x)) + ((ld) & (!sk[12]) & (!g233) & (g1298) & (!keyx11x)) + ((ld) & (!sk[12]) & (!g233) & (g1298) & (keyx11x)) + ((ld) & (!sk[12]) & (g233) & (!g1298) & (!keyx11x)) + ((ld) & (!sk[12]) & (g233) & (!g1298) & (keyx11x)) + ((ld) & (!sk[12]) & (g233) & (g1298) & (!keyx11x)) + ((ld) & (!sk[12]) & (g233) & (g1298) & (keyx11x)) + ((ld) & (sk[12]) & (!g233) & (!g1298) & (keyx11x)) + ((ld) & (sk[12]) & (!g233) & (g1298) & (keyx11x)) + ((ld) & (sk[12]) & (g233) & (!g1298) & (keyx11x)) + ((ld) & (sk[12]) & (g233) & (g1298) & (keyx11x)));
	assign g1300 = (((!g148) & (!g155) & (!g190) & (!g197) & (!g176) & (g183)) + ((!g148) & (!g155) & (g190) & (!g197) & (!g176) & (g183)) + ((!g148) & (!g155) & (g190) & (!g197) & (g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (!g197) & (g176) & (g183)) + ((!g148) & (!g155) & (g190) & (g197) & (!g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (g197) & (g176) & (!g183)) + ((!g148) & (g155) & (!g190) & (!g197) & (!g176) & (!g183)) + ((!g148) & (g155) & (!g190) & (!g197) & (!g176) & (g183)) + ((!g148) & (g155) & (!g190) & (g197) & (!g176) & (!g183)) + ((!g148) & (g155) & (!g190) & (g197) & (!g176) & (g183)) + ((!g148) & (g155) & (!g190) & (g197) & (g176) & (g183)) + ((!g148) & (g155) & (g190) & (g197) & (!g176) & (g183)) + ((!g148) & (g155) & (g190) & (g197) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g197) & (!g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g197) & (!g176) & (g183)) + ((g148) & (!g155) & (!g190) & (g197) & (!g176) & (g183)) + ((g148) & (!g155) & (g190) & (!g197) & (g176) & (!g183)) + ((g148) & (!g155) & (g190) & (g197) & (!g176) & (!g183)) + ((g148) & (!g155) & (g190) & (g197) & (!g176) & (g183)) + ((g148) & (!g155) & (g190) & (g197) & (g176) & (!g183)) + ((g148) & (g155) & (!g190) & (!g197) & (!g176) & (!g183)) + ((g148) & (g155) & (!g190) & (!g197) & (g176) & (!g183)) + ((g148) & (g155) & (!g190) & (g197) & (g176) & (!g183)) + ((g148) & (g155) & (g190) & (!g197) & (!g176) & (!g183)) + ((g148) & (g155) & (g190) & (!g197) & (!g176) & (g183)) + ((g148) & (g155) & (g190) & (g197) & (!g176) & (g183)));
	assign g1301 = (((!g148) & (!g155) & (!g190) & (!g197) & (!g176) & (!g183)) + ((!g148) & (!g155) & (!g190) & (!g197) & (!g176) & (g183)) + ((!g148) & (!g155) & (!g190) & (!g197) & (g176) & (!g183)) + ((!g148) & (!g155) & (!g190) & (!g197) & (g176) & (g183)) + ((!g148) & (!g155) & (!g190) & (g197) & (!g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (!g197) & (!g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (!g197) & (g176) & (g183)) + ((!g148) & (!g155) & (g190) & (g197) & (!g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (g197) & (g176) & (g183)) + ((!g148) & (g155) & (!g190) & (!g197) & (!g176) & (g183)) + ((!g148) & (g155) & (!g190) & (g197) & (g176) & (!g183)) + ((!g148) & (g155) & (g190) & (!g197) & (!g176) & (!g183)) + ((!g148) & (g155) & (g190) & (!g197) & (!g176) & (g183)) + ((!g148) & (g155) & (g190) & (!g197) & (g176) & (!g183)) + ((!g148) & (g155) & (g190) & (!g197) & (g176) & (g183)) + ((!g148) & (g155) & (g190) & (g197) & (!g176) & (!g183)) + ((!g148) & (g155) & (g190) & (g197) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g197) & (!g176) & (g183)) + ((g148) & (!g155) & (!g190) & (!g197) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g197) & (g176) & (g183)) + ((g148) & (!g155) & (!g190) & (g197) & (!g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (g197) & (g176) & (g183)) + ((g148) & (!g155) & (g190) & (!g197) & (g176) & (!g183)) + ((g148) & (!g155) & (g190) & (!g197) & (g176) & (g183)) + ((g148) & (!g155) & (g190) & (g197) & (!g176) & (g183)) + ((g148) & (g155) & (!g190) & (!g197) & (g176) & (!g183)) + ((g148) & (g155) & (!g190) & (!g197) & (g176) & (g183)) + ((g148) & (g155) & (!g190) & (g197) & (!g176) & (!g183)) + ((g148) & (g155) & (!g190) & (g197) & (!g176) & (g183)) + ((g148) & (g155) & (g190) & (!g197) & (g176) & (!g183)) + ((g148) & (g155) & (g190) & (!g197) & (g176) & (g183)) + ((g148) & (g155) & (g190) & (g197) & (!g176) & (g183)));
	assign g1302 = (((!g148) & (!g155) & (!g190) & (!g197) & (!g176) & (!g183)) + ((!g148) & (!g155) & (!g190) & (!g197) & (!g176) & (g183)) + ((!g148) & (!g155) & (g190) & (!g197) & (!g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (!g197) & (g176) & (g183)) + ((!g148) & (!g155) & (g190) & (g197) & (!g176) & (g183)) + ((!g148) & (g155) & (!g190) & (g197) & (!g176) & (!g183)) + ((!g148) & (g155) & (!g190) & (g197) & (g176) & (!g183)) + ((!g148) & (g155) & (!g190) & (g197) & (g176) & (g183)) + ((!g148) & (g155) & (g190) & (!g197) & (!g176) & (!g183)) + ((!g148) & (g155) & (g190) & (!g197) & (g176) & (!g183)) + ((!g148) & (g155) & (g190) & (!g197) & (g176) & (g183)) + ((!g148) & (g155) & (g190) & (g197) & (!g176) & (!g183)) + ((!g148) & (g155) & (g190) & (g197) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g197) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g197) & (g176) & (g183)) + ((g148) & (!g155) & (!g190) & (g197) & (!g176) & (g183)) + ((g148) & (!g155) & (!g190) & (g197) & (g176) & (g183)) + ((g148) & (!g155) & (g190) & (!g197) & (!g176) & (!g183)) + ((g148) & (!g155) & (g190) & (!g197) & (!g176) & (g183)) + ((g148) & (!g155) & (g190) & (!g197) & (g176) & (g183)) + ((g148) & (!g155) & (g190) & (g197) & (!g176) & (!g183)) + ((g148) & (!g155) & (g190) & (g197) & (!g176) & (g183)) + ((g148) & (!g155) & (g190) & (g197) & (g176) & (!g183)) + ((g148) & (!g155) & (g190) & (g197) & (g176) & (g183)) + ((g148) & (g155) & (!g190) & (!g197) & (!g176) & (g183)) + ((g148) & (g155) & (!g190) & (g197) & (!g176) & (!g183)) + ((g148) & (g155) & (!g190) & (g197) & (g176) & (!g183)) + ((g148) & (g155) & (g190) & (!g197) & (!g176) & (!g183)) + ((g148) & (g155) & (g190) & (!g197) & (!g176) & (g183)) + ((g148) & (g155) & (g190) & (!g197) & (g176) & (!g183)) + ((g148) & (g155) & (g190) & (g197) & (!g176) & (!g183)) + ((g148) & (g155) & (g190) & (g197) & (g176) & (!g183)));
	assign g1303 = (((!g148) & (!g155) & (!g190) & (!g197) & (g176) & (g183)) + ((!g148) & (!g155) & (!g190) & (g197) & (!g176) & (!g183)) + ((!g148) & (!g155) & (!g190) & (g197) & (g176) & (g183)) + ((!g148) & (!g155) & (g190) & (!g197) & (!g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (!g197) & (g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (g197) & (!g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (g197) & (!g176) & (g183)) + ((!g148) & (!g155) & (g190) & (g197) & (g176) & (!g183)) + ((!g148) & (g155) & (!g190) & (!g197) & (!g176) & (!g183)) + ((!g148) & (g155) & (!g190) & (g197) & (!g176) & (g183)) + ((!g148) & (g155) & (!g190) & (g197) & (g176) & (!g183)) + ((!g148) & (g155) & (!g190) & (g197) & (g176) & (g183)) + ((!g148) & (g155) & (g190) & (!g197) & (!g176) & (!g183)) + ((!g148) & (g155) & (g190) & (g197) & (!g176) & (!g183)) + ((!g148) & (g155) & (g190) & (g197) & (!g176) & (g183)) + ((g148) & (!g155) & (!g190) & (!g197) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g197) & (g176) & (g183)) + ((g148) & (!g155) & (g190) & (!g197) & (!g176) & (!g183)) + ((g148) & (!g155) & (g190) & (!g197) & (g176) & (!g183)) + ((g148) & (!g155) & (g190) & (g197) & (g176) & (!g183)) + ((g148) & (g155) & (!g190) & (!g197) & (g176) & (!g183)) + ((g148) & (g155) & (!g190) & (g197) & (g176) & (g183)) + ((g148) & (g155) & (g190) & (!g197) & (!g176) & (!g183)) + ((g148) & (g155) & (g190) & (!g197) & (!g176) & (g183)) + ((g148) & (g155) & (g190) & (!g197) & (g176) & (!g183)) + ((g148) & (g155) & (g190) & (g197) & (!g176) & (!g183)));
	assign g1304 = (((!g1300) & (!g1301) & (!g1302) & (!g1303) & (g162) & (g169)) + ((!g1300) & (!g1301) & (g1302) & (!g1303) & (!g162) & (g169)) + ((!g1300) & (!g1301) & (g1302) & (!g1303) & (g162) & (g169)) + ((!g1300) & (!g1301) & (g1302) & (g1303) & (!g162) & (g169)) + ((!g1300) & (g1301) & (!g1302) & (!g1303) & (g162) & (!g169)) + ((!g1300) & (g1301) & (!g1302) & (!g1303) & (g162) & (g169)) + ((!g1300) & (g1301) & (!g1302) & (g1303) & (g162) & (!g169)) + ((!g1300) & (g1301) & (g1302) & (!g1303) & (!g162) & (g169)) + ((!g1300) & (g1301) & (g1302) & (!g1303) & (g162) & (!g169)) + ((!g1300) & (g1301) & (g1302) & (!g1303) & (g162) & (g169)) + ((!g1300) & (g1301) & (g1302) & (g1303) & (!g162) & (g169)) + ((!g1300) & (g1301) & (g1302) & (g1303) & (g162) & (!g169)) + ((g1300) & (!g1301) & (!g1302) & (!g1303) & (!g162) & (!g169)) + ((g1300) & (!g1301) & (!g1302) & (!g1303) & (g162) & (g169)) + ((g1300) & (!g1301) & (!g1302) & (g1303) & (!g162) & (!g169)) + ((g1300) & (!g1301) & (g1302) & (!g1303) & (!g162) & (!g169)) + ((g1300) & (!g1301) & (g1302) & (!g1303) & (!g162) & (g169)) + ((g1300) & (!g1301) & (g1302) & (!g1303) & (g162) & (g169)) + ((g1300) & (!g1301) & (g1302) & (g1303) & (!g162) & (!g169)) + ((g1300) & (!g1301) & (g1302) & (g1303) & (!g162) & (g169)) + ((g1300) & (g1301) & (!g1302) & (!g1303) & (!g162) & (!g169)) + ((g1300) & (g1301) & (!g1302) & (!g1303) & (g162) & (!g169)) + ((g1300) & (g1301) & (!g1302) & (!g1303) & (g162) & (g169)) + ((g1300) & (g1301) & (!g1302) & (g1303) & (!g162) & (!g169)) + ((g1300) & (g1301) & (!g1302) & (g1303) & (g162) & (!g169)) + ((g1300) & (g1301) & (g1302) & (!g1303) & (!g162) & (!g169)) + ((g1300) & (g1301) & (g1302) & (!g1303) & (!g162) & (g169)) + ((g1300) & (g1301) & (g1302) & (!g1303) & (g162) & (!g169)) + ((g1300) & (g1301) & (g1302) & (!g1303) & (g162) & (g169)) + ((g1300) & (g1301) & (g1302) & (g1303) & (!g162) & (!g169)) + ((g1300) & (g1301) & (g1302) & (g1303) & (!g162) & (g169)) + ((g1300) & (g1301) & (g1302) & (g1303) & (g162) & (!g169)));
	assign g1305 = (((!g496) & (!sk[18]) & (!g752) & (g1008) & (!g1304)) + ((!g496) & (!sk[18]) & (!g752) & (g1008) & (g1304)) + ((!g496) & (!sk[18]) & (g752) & (!g1008) & (!g1304)) + ((!g496) & (!sk[18]) & (g752) & (!g1008) & (g1304)) + ((!g496) & (!sk[18]) & (g752) & (g1008) & (!g1304)) + ((!g496) & (!sk[18]) & (g752) & (g1008) & (g1304)) + ((!g496) & (sk[18]) & (!g752) & (!g1008) & (g1304)) + ((!g496) & (sk[18]) & (!g752) & (g1008) & (!g1304)) + ((!g496) & (sk[18]) & (g752) & (!g1008) & (!g1304)) + ((!g496) & (sk[18]) & (g752) & (g1008) & (g1304)) + ((g496) & (!sk[18]) & (!g752) & (g1008) & (!g1304)) + ((g496) & (!sk[18]) & (!g752) & (g1008) & (g1304)) + ((g496) & (!sk[18]) & (g752) & (!g1008) & (!g1304)) + ((g496) & (!sk[18]) & (g752) & (!g1008) & (g1304)) + ((g496) & (!sk[18]) & (g752) & (g1008) & (!g1304)) + ((g496) & (!sk[18]) & (g752) & (g1008) & (g1304)) + ((g496) & (sk[18]) & (!g752) & (!g1008) & (!g1304)) + ((g496) & (sk[18]) & (!g752) & (g1008) & (g1304)) + ((g496) & (sk[18]) & (g752) & (!g1008) & (g1304)) + ((g496) & (sk[18]) & (g752) & (g1008) & (!g1304)));
	assign g1306 = (((!ld) & (!g240) & (!sk[19]) & (g1305) & (!keyx12x)) + ((!ld) & (!g240) & (!sk[19]) & (g1305) & (keyx12x)) + ((!ld) & (!g240) & (sk[19]) & (g1305) & (!keyx12x)) + ((!ld) & (!g240) & (sk[19]) & (g1305) & (keyx12x)) + ((!ld) & (g240) & (!sk[19]) & (!g1305) & (!keyx12x)) + ((!ld) & (g240) & (!sk[19]) & (!g1305) & (keyx12x)) + ((!ld) & (g240) & (!sk[19]) & (g1305) & (!keyx12x)) + ((!ld) & (g240) & (!sk[19]) & (g1305) & (keyx12x)) + ((!ld) & (g240) & (sk[19]) & (!g1305) & (!keyx12x)) + ((!ld) & (g240) & (sk[19]) & (!g1305) & (keyx12x)) + ((ld) & (!g240) & (!sk[19]) & (g1305) & (!keyx12x)) + ((ld) & (!g240) & (!sk[19]) & (g1305) & (keyx12x)) + ((ld) & (!g240) & (sk[19]) & (!g1305) & (keyx12x)) + ((ld) & (!g240) & (sk[19]) & (g1305) & (keyx12x)) + ((ld) & (g240) & (!sk[19]) & (!g1305) & (!keyx12x)) + ((ld) & (g240) & (!sk[19]) & (!g1305) & (keyx12x)) + ((ld) & (g240) & (!sk[19]) & (g1305) & (!keyx12x)) + ((ld) & (g240) & (!sk[19]) & (g1305) & (keyx12x)) + ((ld) & (g240) & (sk[19]) & (!g1305) & (keyx12x)) + ((ld) & (g240) & (sk[19]) & (g1305) & (keyx12x)));
	assign g1307 = (((!g148) & (!g155) & (!g190) & (!g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (!g190) & (!g169) & (g176) & (g183)) + ((!g148) & (!g155) & (!g190) & (g169) & (g176) & (g183)) + ((!g148) & (!g155) & (g190) & (!g169) & (!g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (!g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (g190) & (!g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (!g169) & (g176) & (g183)) + ((!g148) & (!g155) & (g190) & (g169) & (!g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (g169) & (!g176) & (g183)) + ((!g148) & (g155) & (!g190) & (!g169) & (!g176) & (g183)) + ((!g148) & (g155) & (!g190) & (!g169) & (g176) & (!g183)) + ((!g148) & (g155) & (!g190) & (g169) & (g176) & (g183)) + ((!g148) & (g155) & (g190) & (!g169) & (g176) & (!g183)) + ((!g148) & (g155) & (g190) & (!g169) & (g176) & (g183)) + ((!g148) & (g155) & (g190) & (g169) & (!g176) & (!g183)) + ((!g148) & (g155) & (g190) & (g169) & (!g176) & (g183)) + ((!g148) & (g155) & (g190) & (g169) & (g176) & (g183)) + ((g148) & (!g155) & (!g190) & (!g169) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g169) & (g176) & (g183)) + ((g148) & (!g155) & (!g190) & (g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (g169) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (g169) & (g176) & (g183)) + ((g148) & (!g155) & (g190) & (!g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (g190) & (!g169) & (g176) & (!g183)) + ((g148) & (!g155) & (g190) & (g169) & (g176) & (!g183)) + ((g148) & (g155) & (!g190) & (!g169) & (g176) & (g183)) + ((g148) & (g155) & (g190) & (!g169) & (!g176) & (!g183)) + ((g148) & (g155) & (g190) & (!g169) & (g176) & (g183)));
	assign g1308 = (((!g148) & (!g155) & (!g190) & (!g169) & (!g176) & (!g183)) + ((!g148) & (!g155) & (!g190) & (g169) & (!g176) & (!g183)) + ((!g148) & (!g155) & (!g190) & (g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (!g190) & (g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (!g169) & (g176) & (g183)) + ((!g148) & (!g155) & (g190) & (g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (g190) & (g169) & (g176) & (g183)) + ((!g148) & (g155) & (!g190) & (!g169) & (!g176) & (!g183)) + ((!g148) & (g155) & (!g190) & (!g169) & (g176) & (!g183)) + ((!g148) & (g155) & (g190) & (!g169) & (!g176) & (g183)) + ((!g148) & (g155) & (g190) & (!g169) & (g176) & (g183)) + ((!g148) & (g155) & (g190) & (g169) & (!g176) & (g183)) + ((!g148) & (g155) & (g190) & (g169) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g169) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g169) & (g176) & (g183)) + ((g148) & (!g155) & (!g190) & (g169) & (!g176) & (g183)) + ((g148) & (!g155) & (!g190) & (g169) & (g176) & (g183)) + ((g148) & (!g155) & (g190) & (g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (g190) & (g169) & (!g176) & (g183)) + ((g148) & (!g155) & (g190) & (g169) & (g176) & (g183)) + ((g148) & (g155) & (!g190) & (!g169) & (!g176) & (g183)) + ((g148) & (g155) & (!g190) & (!g169) & (g176) & (!g183)) + ((g148) & (g155) & (!g190) & (g169) & (g176) & (!g183)) + ((g148) & (g155) & (g190) & (!g169) & (!g176) & (g183)) + ((g148) & (g155) & (g190) & (!g169) & (g176) & (g183)) + ((g148) & (g155) & (g190) & (g169) & (!g176) & (!g183)) + ((g148) & (g155) & (g190) & (g169) & (g176) & (g183)));
	assign g1309 = (((!g148) & (!g155) & (!g190) & (!g169) & (g176) & (g183)) + ((!g148) & (!g155) & (!g190) & (g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (!g169) & (!g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (!g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (g190) & (!g169) & (g176) & (g183)) + ((!g148) & (!g155) & (g190) & (g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (g190) & (g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (g190) & (g169) & (g176) & (g183)) + ((!g148) & (g155) & (!g190) & (!g169) & (g176) & (!g183)) + ((!g148) & (g155) & (!g190) & (!g169) & (g176) & (g183)) + ((!g148) & (g155) & (g190) & (!g169) & (!g176) & (!g183)) + ((!g148) & (g155) & (g190) & (g169) & (!g176) & (g183)) + ((!g148) & (g155) & (g190) & (g169) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g169) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (!g169) & (g176) & (g183)) + ((g148) & (!g155) & (!g190) & (g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (g169) & (!g176) & (g183)) + ((g148) & (!g155) & (g190) & (!g169) & (!g176) & (g183)) + ((g148) & (!g155) & (g190) & (!g169) & (g176) & (g183)) + ((g148) & (!g155) & (g190) & (g169) & (g176) & (!g183)) + ((g148) & (g155) & (!g190) & (!g169) & (!g176) & (!g183)) + ((g148) & (g155) & (!g190) & (!g169) & (!g176) & (g183)) + ((g148) & (g155) & (!g190) & (!g169) & (g176) & (g183)) + ((g148) & (g155) & (!g190) & (g169) & (!g176) & (g183)) + ((g148) & (g155) & (!g190) & (g169) & (g176) & (!g183)) + ((g148) & (g155) & (g190) & (!g169) & (!g176) & (g183)) + ((g148) & (g155) & (g190) & (!g169) & (g176) & (!g183)) + ((g148) & (g155) & (g190) & (g169) & (!g176) & (!g183)) + ((g148) & (g155) & (g190) & (g169) & (g176) & (!g183)) + ((g148) & (g155) & (g190) & (g169) & (g176) & (g183)));
	assign g1310 = (((!g148) & (!g155) & (!g190) & (!g169) & (g176) & (!g183)) + ((!g148) & (!g155) & (!g190) & (g169) & (!g176) & (!g183)) + ((!g148) & (!g155) & (!g190) & (g169) & (g176) & (g183)) + ((!g148) & (!g155) & (g190) & (!g169) & (!g176) & (g183)) + ((!g148) & (!g155) & (g190) & (!g169) & (g176) & (g183)) + ((!g148) & (!g155) & (g190) & (g169) & (g176) & (g183)) + ((!g148) & (g155) & (!g190) & (!g169) & (!g176) & (g183)) + ((!g148) & (g155) & (!g190) & (g169) & (!g176) & (g183)) + ((!g148) & (g155) & (!g190) & (g169) & (g176) & (g183)) + ((!g148) & (g155) & (g190) & (!g169) & (!g176) & (!g183)) + ((!g148) & (g155) & (g190) & (!g169) & (g176) & (!g183)) + ((!g148) & (g155) & (g190) & (g169) & (!g176) & (g183)) + ((!g148) & (g155) & (g190) & (g169) & (g176) & (g183)) + ((g148) & (!g155) & (!g190) & (!g169) & (g176) & (!g183)) + ((g148) & (!g155) & (!g190) & (g169) & (g176) & (g183)) + ((g148) & (!g155) & (g190) & (!g169) & (!g176) & (!g183)) + ((g148) & (!g155) & (g190) & (!g169) & (g176) & (g183)) + ((g148) & (!g155) & (g190) & (g169) & (!g176) & (!g183)) + ((g148) & (g155) & (!g190) & (!g169) & (g176) & (g183)) + ((g148) & (g155) & (!g190) & (g169) & (!g176) & (!g183)) + ((g148) & (g155) & (!g190) & (g169) & (!g176) & (g183)) + ((g148) & (g155) & (g190) & (!g169) & (g176) & (g183)));
	assign g1311 = (((!g1307) & (!g1308) & (!g1309) & (!g1310) & (!g197) & (!g162)) + ((!g1307) & (!g1308) & (!g1309) & (!g1310) & (!g197) & (g162)) + ((!g1307) & (!g1308) & (!g1309) & (!g1310) & (g197) & (!g162)) + ((!g1307) & (!g1308) & (!g1309) & (g1310) & (!g197) & (!g162)) + ((!g1307) & (!g1308) & (!g1309) & (g1310) & (!g197) & (g162)) + ((!g1307) & (!g1308) & (!g1309) & (g1310) & (g197) & (!g162)) + ((!g1307) & (!g1308) & (!g1309) & (g1310) & (g197) & (g162)) + ((!g1307) & (!g1308) & (g1309) & (!g1310) & (!g197) & (!g162)) + ((!g1307) & (!g1308) & (g1309) & (!g1310) & (g197) & (!g162)) + ((!g1307) & (!g1308) & (g1309) & (g1310) & (!g197) & (!g162)) + ((!g1307) & (!g1308) & (g1309) & (g1310) & (g197) & (!g162)) + ((!g1307) & (!g1308) & (g1309) & (g1310) & (g197) & (g162)) + ((!g1307) & (g1308) & (!g1309) & (!g1310) & (!g197) & (!g162)) + ((!g1307) & (g1308) & (!g1309) & (!g1310) & (!g197) & (g162)) + ((!g1307) & (g1308) & (!g1309) & (g1310) & (!g197) & (!g162)) + ((!g1307) & (g1308) & (!g1309) & (g1310) & (!g197) & (g162)) + ((!g1307) & (g1308) & (!g1309) & (g1310) & (g197) & (g162)) + ((!g1307) & (g1308) & (g1309) & (!g1310) & (!g197) & (!g162)) + ((!g1307) & (g1308) & (g1309) & (g1310) & (!g197) & (!g162)) + ((!g1307) & (g1308) & (g1309) & (g1310) & (g197) & (g162)) + ((g1307) & (!g1308) & (!g1309) & (!g1310) & (!g197) & (g162)) + ((g1307) & (!g1308) & (!g1309) & (!g1310) & (g197) & (!g162)) + ((g1307) & (!g1308) & (!g1309) & (g1310) & (!g197) & (g162)) + ((g1307) & (!g1308) & (!g1309) & (g1310) & (g197) & (!g162)) + ((g1307) & (!g1308) & (!g1309) & (g1310) & (g197) & (g162)) + ((g1307) & (!g1308) & (g1309) & (!g1310) & (g197) & (!g162)) + ((g1307) & (!g1308) & (g1309) & (g1310) & (g197) & (!g162)) + ((g1307) & (!g1308) & (g1309) & (g1310) & (g197) & (g162)) + ((g1307) & (g1308) & (!g1309) & (!g1310) & (!g197) & (g162)) + ((g1307) & (g1308) & (!g1309) & (g1310) & (!g197) & (g162)) + ((g1307) & (g1308) & (!g1309) & (g1310) & (g197) & (g162)) + ((g1307) & (g1308) & (g1309) & (g1310) & (g197) & (g162)));
	assign g1312 = (((!g503) & (!g759) & (!g1015) & (sk[25]) & (g1311)) + ((!g503) & (!g759) & (g1015) & (!sk[25]) & (!g1311)) + ((!g503) & (!g759) & (g1015) & (!sk[25]) & (g1311)) + ((!g503) & (!g759) & (g1015) & (sk[25]) & (!g1311)) + ((!g503) & (g759) & (!g1015) & (!sk[25]) & (!g1311)) + ((!g503) & (g759) & (!g1015) & (!sk[25]) & (g1311)) + ((!g503) & (g759) & (!g1015) & (sk[25]) & (!g1311)) + ((!g503) & (g759) & (g1015) & (!sk[25]) & (!g1311)) + ((!g503) & (g759) & (g1015) & (!sk[25]) & (g1311)) + ((!g503) & (g759) & (g1015) & (sk[25]) & (g1311)) + ((g503) & (!g759) & (!g1015) & (sk[25]) & (!g1311)) + ((g503) & (!g759) & (g1015) & (!sk[25]) & (!g1311)) + ((g503) & (!g759) & (g1015) & (!sk[25]) & (g1311)) + ((g503) & (!g759) & (g1015) & (sk[25]) & (g1311)) + ((g503) & (g759) & (!g1015) & (!sk[25]) & (!g1311)) + ((g503) & (g759) & (!g1015) & (!sk[25]) & (g1311)) + ((g503) & (g759) & (!g1015) & (sk[25]) & (g1311)) + ((g503) & (g759) & (g1015) & (!sk[25]) & (!g1311)) + ((g503) & (g759) & (g1015) & (!sk[25]) & (g1311)) + ((g503) & (g759) & (g1015) & (sk[25]) & (!g1311)));
	assign g1313 = (((!ld) & (!sk[26]) & (!g247) & (g1312) & (!keyx13x)) + ((!ld) & (!sk[26]) & (!g247) & (g1312) & (keyx13x)) + ((!ld) & (!sk[26]) & (g247) & (!g1312) & (!keyx13x)) + ((!ld) & (!sk[26]) & (g247) & (!g1312) & (keyx13x)) + ((!ld) & (!sk[26]) & (g247) & (g1312) & (!keyx13x)) + ((!ld) & (!sk[26]) & (g247) & (g1312) & (keyx13x)) + ((!ld) & (sk[26]) & (!g247) & (g1312) & (!keyx13x)) + ((!ld) & (sk[26]) & (!g247) & (g1312) & (keyx13x)) + ((!ld) & (sk[26]) & (g247) & (!g1312) & (!keyx13x)) + ((!ld) & (sk[26]) & (g247) & (!g1312) & (keyx13x)) + ((ld) & (!sk[26]) & (!g247) & (g1312) & (!keyx13x)) + ((ld) & (!sk[26]) & (!g247) & (g1312) & (keyx13x)) + ((ld) & (!sk[26]) & (g247) & (!g1312) & (!keyx13x)) + ((ld) & (!sk[26]) & (g247) & (!g1312) & (keyx13x)) + ((ld) & (!sk[26]) & (g247) & (g1312) & (!keyx13x)) + ((ld) & (!sk[26]) & (g247) & (g1312) & (keyx13x)) + ((ld) & (sk[26]) & (!g247) & (!g1312) & (keyx13x)) + ((ld) & (sk[26]) & (!g247) & (g1312) & (keyx13x)) + ((ld) & (sk[26]) & (g247) & (!g1312) & (keyx13x)) + ((ld) & (sk[26]) & (g247) & (g1312) & (keyx13x)));
	assign g1314 = (((!g148) & (!g197) & (!g162) & (!g169) & (!g176) & (g183)) + ((!g148) & (!g197) & (!g162) & (!g169) & (g176) & (g183)) + ((!g148) & (!g197) & (!g162) & (g169) & (!g176) & (!g183)) + ((!g148) & (!g197) & (!g162) & (g169) & (!g176) & (g183)) + ((!g148) & (!g197) & (!g162) & (g169) & (g176) & (!g183)) + ((!g148) & (!g197) & (!g162) & (g169) & (g176) & (g183)) + ((!g148) & (!g197) & (g162) & (!g169) & (!g176) & (g183)) + ((!g148) & (!g197) & (g162) & (!g169) & (g176) & (g183)) + ((!g148) & (!g197) & (g162) & (g169) & (g176) & (!g183)) + ((!g148) & (g197) & (g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (g197) & (g162) & (!g169) & (g176) & (g183)) + ((!g148) & (g197) & (g162) & (g169) & (!g176) & (g183)) + ((g148) & (!g197) & (!g162) & (!g169) & (g176) & (!g183)) + ((g148) & (!g197) & (!g162) & (g169) & (!g176) & (!g183)) + ((g148) & (!g197) & (!g162) & (g169) & (!g176) & (g183)) + ((g148) & (!g197) & (!g162) & (g169) & (g176) & (g183)) + ((g148) & (!g197) & (g162) & (!g169) & (!g176) & (g183)) + ((g148) & (!g197) & (g162) & (!g169) & (g176) & (g183)) + ((g148) & (!g197) & (g162) & (g169) & (g176) & (!g183)) + ((g148) & (!g197) & (g162) & (g169) & (g176) & (g183)) + ((g148) & (g197) & (!g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (g197) & (!g162) & (!g169) & (!g176) & (g183)) + ((g148) & (g197) & (!g162) & (!g169) & (g176) & (!g183)) + ((g148) & (g197) & (!g162) & (g169) & (!g176) & (!g183)) + ((g148) & (g197) & (g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (g197) & (g162) & (!g169) & (!g176) & (g183)) + ((g148) & (g197) & (g162) & (!g169) & (g176) & (!g183)) + ((g148) & (g197) & (g162) & (g169) & (!g176) & (g183)));
	assign g1315 = (((!g148) & (!g197) & (!g162) & (!g169) & (!g176) & (!g183)) + ((!g148) & (!g197) & (!g162) & (g169) & (g176) & (g183)) + ((!g148) & (!g197) & (g162) & (!g169) & (!g176) & (!g183)) + ((!g148) & (!g197) & (g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (!g197) & (g162) & (!g169) & (g176) & (g183)) + ((!g148) & (!g197) & (g162) & (g169) & (!g176) & (!g183)) + ((!g148) & (!g197) & (g162) & (g169) & (g176) & (g183)) + ((!g148) & (g197) & (!g162) & (!g169) & (!g176) & (!g183)) + ((!g148) & (g197) & (!g162) & (!g169) & (g176) & (g183)) + ((!g148) & (g197) & (!g162) & (g169) & (!g176) & (g183)) + ((!g148) & (g197) & (g162) & (!g169) & (!g176) & (!g183)) + ((!g148) & (g197) & (g162) & (!g169) & (g176) & (g183)) + ((!g148) & (g197) & (g162) & (g169) & (g176) & (!g183)) + ((!g148) & (g197) & (g162) & (g169) & (g176) & (g183)) + ((g148) & (!g197) & (!g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (!g197) & (!g162) & (!g169) & (g176) & (g183)) + ((g148) & (!g197) & (!g162) & (g169) & (!g176) & (!g183)) + ((g148) & (!g197) & (!g162) & (g169) & (g176) & (g183)) + ((g148) & (!g197) & (g162) & (!g169) & (g176) & (g183)) + ((g148) & (!g197) & (g162) & (g169) & (!g176) & (g183)) + ((g148) & (g197) & (!g162) & (!g169) & (g176) & (!g183)) + ((g148) & (g197) & (!g162) & (!g169) & (g176) & (g183)) + ((g148) & (g197) & (!g162) & (g169) & (!g176) & (g183)) + ((g148) & (g197) & (!g162) & (g169) & (g176) & (!g183)) + ((g148) & (g197) & (!g162) & (g169) & (g176) & (g183)) + ((g148) & (g197) & (g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (g197) & (g162) & (!g169) & (g176) & (!g183)) + ((g148) & (g197) & (g162) & (g169) & (!g176) & (!g183)));
	assign g1316 = (((!g148) & (!g197) & (!g162) & (!g169) & (!g176) & (g183)) + ((!g148) & (!g197) & (!g162) & (!g169) & (g176) & (g183)) + ((!g148) & (!g197) & (!g162) & (g169) & (g176) & (!g183)) + ((!g148) & (!g197) & (!g162) & (g169) & (g176) & (g183)) + ((!g148) & (!g197) & (g162) & (!g169) & (g176) & (g183)) + ((!g148) & (!g197) & (g162) & (g169) & (!g176) & (!g183)) + ((!g148) & (!g197) & (g162) & (g169) & (!g176) & (g183)) + ((!g148) & (!g197) & (g162) & (g169) & (g176) & (g183)) + ((!g148) & (g197) & (!g162) & (!g169) & (!g176) & (!g183)) + ((!g148) & (g197) & (!g162) & (!g169) & (!g176) & (g183)) + ((!g148) & (g197) & (!g162) & (!g169) & (g176) & (g183)) + ((!g148) & (g197) & (!g162) & (g169) & (!g176) & (g183)) + ((!g148) & (g197) & (!g162) & (g169) & (g176) & (!g183)) + ((!g148) & (g197) & (g162) & (!g169) & (!g176) & (g183)) + ((!g148) & (g197) & (g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (g197) & (g162) & (g169) & (!g176) & (!g183)) + ((!g148) & (g197) & (g162) & (g169) & (g176) & (!g183)) + ((!g148) & (g197) & (g162) & (g169) & (g176) & (g183)) + ((g148) & (!g197) & (!g162) & (!g169) & (!g176) & (g183)) + ((g148) & (!g197) & (!g162) & (g169) & (!g176) & (!g183)) + ((g148) & (!g197) & (!g162) & (g169) & (g176) & (!g183)) + ((g148) & (!g197) & (g162) & (!g169) & (g176) & (g183)) + ((g148) & (!g197) & (g162) & (g169) & (!g176) & (g183)) + ((g148) & (g197) & (!g162) & (!g169) & (!g176) & (g183)) + ((g148) & (g197) & (!g162) & (g169) & (!g176) & (!g183)) + ((g148) & (g197) & (!g162) & (g169) & (g176) & (!g183)) + ((g148) & (g197) & (g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (g197) & (g162) & (!g169) & (g176) & (!g183)) + ((g148) & (g197) & (g162) & (!g169) & (g176) & (g183)) + ((g148) & (g197) & (g162) & (g169) & (g176) & (g183)));
	assign g1317 = (((!g148) & (!g197) & (!g162) & (!g169) & (g176) & (g183)) + ((!g148) & (!g197) & (!g162) & (g169) & (!g176) & (!g183)) + ((!g148) & (!g197) & (!g162) & (g169) & (g176) & (g183)) + ((!g148) & (!g197) & (g162) & (!g169) & (!g176) & (!g183)) + ((!g148) & (!g197) & (g162) & (g169) & (g176) & (!g183)) + ((!g148) & (!g197) & (g162) & (g169) & (g176) & (g183)) + ((!g148) & (g197) & (!g162) & (g169) & (!g176) & (!g183)) + ((!g148) & (g197) & (!g162) & (g169) & (g176) & (!g183)) + ((!g148) & (g197) & (g162) & (!g169) & (g176) & (!g183)) + ((!g148) & (g197) & (g162) & (!g169) & (g176) & (g183)) + ((g148) & (!g197) & (!g162) & (!g169) & (!g176) & (g183)) + ((g148) & (!g197) & (!g162) & (!g169) & (g176) & (!g183)) + ((g148) & (!g197) & (!g162) & (g169) & (!g176) & (g183)) + ((g148) & (!g197) & (g162) & (!g169) & (g176) & (!g183)) + ((g148) & (!g197) & (g162) & (!g169) & (g176) & (g183)) + ((g148) & (!g197) & (g162) & (g169) & (g176) & (!g183)) + ((g148) & (!g197) & (g162) & (g169) & (g176) & (g183)) + ((g148) & (g197) & (!g162) & (!g169) & (g176) & (!g183)) + ((g148) & (g197) & (!g162) & (g169) & (!g176) & (g183)) + ((g148) & (g197) & (g162) & (!g169) & (!g176) & (!g183)) + ((g148) & (g197) & (g162) & (!g169) & (g176) & (g183)) + ((g148) & (g197) & (g162) & (g169) & (!g176) & (g183)));
	assign g1318 = (((!g1314) & (!g1315) & (!g1316) & (!g1317) & (!g190) & (!g155)) + ((!g1314) & (!g1315) & (!g1316) & (!g1317) & (!g190) & (g155)) + ((!g1314) & (!g1315) & (!g1316) & (!g1317) & (g190) & (!g155)) + ((!g1314) & (!g1315) & (!g1316) & (g1317) & (!g190) & (!g155)) + ((!g1314) & (!g1315) & (!g1316) & (g1317) & (!g190) & (g155)) + ((!g1314) & (!g1315) & (!g1316) & (g1317) & (g190) & (!g155)) + ((!g1314) & (!g1315) & (!g1316) & (g1317) & (g190) & (g155)) + ((!g1314) & (!g1315) & (g1316) & (!g1317) & (!g190) & (!g155)) + ((!g1314) & (!g1315) & (g1316) & (!g1317) & (g190) & (!g155)) + ((!g1314) & (!g1315) & (g1316) & (g1317) & (!g190) & (!g155)) + ((!g1314) & (!g1315) & (g1316) & (g1317) & (g190) & (!g155)) + ((!g1314) & (!g1315) & (g1316) & (g1317) & (g190) & (g155)) + ((!g1314) & (g1315) & (!g1316) & (!g1317) & (!g190) & (!g155)) + ((!g1314) & (g1315) & (!g1316) & (!g1317) & (!g190) & (g155)) + ((!g1314) & (g1315) & (!g1316) & (g1317) & (!g190) & (!g155)) + ((!g1314) & (g1315) & (!g1316) & (g1317) & (!g190) & (g155)) + ((!g1314) & (g1315) & (!g1316) & (g1317) & (g190) & (g155)) + ((!g1314) & (g1315) & (g1316) & (!g1317) & (!g190) & (!g155)) + ((!g1314) & (g1315) & (g1316) & (g1317) & (!g190) & (!g155)) + ((!g1314) & (g1315) & (g1316) & (g1317) & (g190) & (g155)) + ((g1314) & (!g1315) & (!g1316) & (!g1317) & (!g190) & (g155)) + ((g1314) & (!g1315) & (!g1316) & (!g1317) & (g190) & (!g155)) + ((g1314) & (!g1315) & (!g1316) & (g1317) & (!g190) & (g155)) + ((g1314) & (!g1315) & (!g1316) & (g1317) & (g190) & (!g155)) + ((g1314) & (!g1315) & (!g1316) & (g1317) & (g190) & (g155)) + ((g1314) & (!g1315) & (g1316) & (!g1317) & (g190) & (!g155)) + ((g1314) & (!g1315) & (g1316) & (g1317) & (g190) & (!g155)) + ((g1314) & (!g1315) & (g1316) & (g1317) & (g190) & (g155)) + ((g1314) & (g1315) & (!g1316) & (!g1317) & (!g190) & (g155)) + ((g1314) & (g1315) & (!g1316) & (g1317) & (!g190) & (g155)) + ((g1314) & (g1315) & (!g1316) & (g1317) & (g190) & (g155)) + ((g1314) & (g1315) & (g1316) & (g1317) & (g190) & (g155)));
	assign g1319 = (((!g510) & (!sk[32]) & (!g766) & (g1022) & (!g1318)) + ((!g510) & (!sk[32]) & (!g766) & (g1022) & (g1318)) + ((!g510) & (!sk[32]) & (g766) & (!g1022) & (!g1318)) + ((!g510) & (!sk[32]) & (g766) & (!g1022) & (g1318)) + ((!g510) & (!sk[32]) & (g766) & (g1022) & (!g1318)) + ((!g510) & (!sk[32]) & (g766) & (g1022) & (g1318)) + ((!g510) & (sk[32]) & (!g766) & (!g1022) & (g1318)) + ((!g510) & (sk[32]) & (!g766) & (g1022) & (!g1318)) + ((!g510) & (sk[32]) & (g766) & (!g1022) & (!g1318)) + ((!g510) & (sk[32]) & (g766) & (g1022) & (g1318)) + ((g510) & (!sk[32]) & (!g766) & (g1022) & (!g1318)) + ((g510) & (!sk[32]) & (!g766) & (g1022) & (g1318)) + ((g510) & (!sk[32]) & (g766) & (!g1022) & (!g1318)) + ((g510) & (!sk[32]) & (g766) & (!g1022) & (g1318)) + ((g510) & (!sk[32]) & (g766) & (g1022) & (!g1318)) + ((g510) & (!sk[32]) & (g766) & (g1022) & (g1318)) + ((g510) & (sk[32]) & (!g766) & (!g1022) & (!g1318)) + ((g510) & (sk[32]) & (!g766) & (g1022) & (g1318)) + ((g510) & (sk[32]) & (g766) & (!g1022) & (g1318)) + ((g510) & (sk[32]) & (g766) & (g1022) & (!g1318)));
	assign g1320 = (((!ld) & (!g254) & (!sk[33]) & (g1319) & (!keyx14x)) + ((!ld) & (!g254) & (!sk[33]) & (g1319) & (keyx14x)) + ((!ld) & (!g254) & (sk[33]) & (g1319) & (!keyx14x)) + ((!ld) & (!g254) & (sk[33]) & (g1319) & (keyx14x)) + ((!ld) & (g254) & (!sk[33]) & (!g1319) & (!keyx14x)) + ((!ld) & (g254) & (!sk[33]) & (!g1319) & (keyx14x)) + ((!ld) & (g254) & (!sk[33]) & (g1319) & (!keyx14x)) + ((!ld) & (g254) & (!sk[33]) & (g1319) & (keyx14x)) + ((!ld) & (g254) & (sk[33]) & (!g1319) & (!keyx14x)) + ((!ld) & (g254) & (sk[33]) & (!g1319) & (keyx14x)) + ((ld) & (!g254) & (!sk[33]) & (g1319) & (!keyx14x)) + ((ld) & (!g254) & (!sk[33]) & (g1319) & (keyx14x)) + ((ld) & (!g254) & (sk[33]) & (!g1319) & (keyx14x)) + ((ld) & (!g254) & (sk[33]) & (g1319) & (keyx14x)) + ((ld) & (g254) & (!sk[33]) & (!g1319) & (!keyx14x)) + ((ld) & (g254) & (!sk[33]) & (!g1319) & (keyx14x)) + ((ld) & (g254) & (!sk[33]) & (g1319) & (!keyx14x)) + ((ld) & (g254) & (!sk[33]) & (g1319) & (keyx14x)) + ((ld) & (g254) & (sk[33]) & (!g1319) & (keyx14x)) + ((ld) & (g254) & (sk[33]) & (g1319) & (keyx14x)));
	assign g1321 = (((!g190) & (!g155) & (!g162) & (!g169) & (!g176) & (g197)) + ((!g190) & (!g155) & (!g162) & (!g169) & (g176) & (!g197)) + ((!g190) & (!g155) & (!g162) & (g169) & (!g176) & (g197)) + ((!g190) & (!g155) & (!g162) & (g169) & (g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (!g169) & (!g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (!g169) & (g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (g169) & (!g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (g169) & (g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (g169) & (g176) & (g197)) + ((!g190) & (g155) & (!g162) & (!g169) & (g176) & (!g197)) + ((!g190) & (g155) & (!g162) & (g169) & (g176) & (!g197)) + ((!g190) & (g155) & (!g162) & (g169) & (g176) & (g197)) + ((!g190) & (g155) & (g162) & (!g169) & (g176) & (g197)) + ((!g190) & (g155) & (g162) & (g169) & (!g176) & (!g197)) + ((g190) & (!g155) & (!g162) & (!g169) & (!g176) & (g197)) + ((g190) & (!g155) & (!g162) & (g169) & (!g176) & (g197)) + ((g190) & (!g155) & (g162) & (g169) & (g176) & (g197)) + ((g190) & (g155) & (!g162) & (!g169) & (g176) & (g197)) + ((g190) & (g155) & (!g162) & (g169) & (!g176) & (!g197)) + ((g190) & (g155) & (!g162) & (g169) & (g176) & (!g197)) + ((g190) & (g155) & (g162) & (!g169) & (!g176) & (g197)) + ((g190) & (g155) & (g162) & (!g169) & (g176) & (!g197)) + ((g190) & (g155) & (g162) & (!g169) & (g176) & (g197)) + ((g190) & (g155) & (g162) & (g169) & (!g176) & (g197)));
	assign g1322 = (((!g190) & (!g155) & (!g162) & (!g169) & (!g176) & (!g197)) + ((!g190) & (!g155) & (!g162) & (!g169) & (!g176) & (g197)) + ((!g190) & (!g155) & (!g162) & (g169) & (!g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (!g169) & (!g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (!g169) & (g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (!g169) & (g176) & (g197)) + ((!g190) & (!g155) & (g162) & (g169) & (!g176) & (g197)) + ((!g190) & (!g155) & (g162) & (g169) & (g176) & (g197)) + ((!g190) & (g155) & (!g162) & (!g169) & (!g176) & (!g197)) + ((!g190) & (g155) & (!g162) & (!g169) & (g176) & (!g197)) + ((!g190) & (g155) & (!g162) & (g169) & (!g176) & (!g197)) + ((!g190) & (g155) & (!g162) & (g169) & (!g176) & (g197)) + ((!g190) & (g155) & (!g162) & (g169) & (g176) & (g197)) + ((!g190) & (g155) & (g162) & (!g169) & (!g176) & (g197)) + ((!g190) & (g155) & (g162) & (g169) & (!g176) & (!g197)) + ((!g190) & (g155) & (g162) & (g169) & (!g176) & (g197)) + ((g190) & (!g155) & (!g162) & (!g169) & (!g176) & (g197)) + ((g190) & (!g155) & (!g162) & (!g169) & (g176) & (g197)) + ((g190) & (!g155) & (!g162) & (g169) & (!g176) & (!g197)) + ((g190) & (!g155) & (!g162) & (g169) & (g176) & (g197)) + ((g190) & (!g155) & (g162) & (!g169) & (!g176) & (!g197)) + ((g190) & (!g155) & (g162) & (!g169) & (g176) & (g197)) + ((g190) & (!g155) & (g162) & (g169) & (g176) & (!g197)) + ((g190) & (g155) & (!g162) & (!g169) & (!g176) & (!g197)) + ((g190) & (g155) & (!g162) & (!g169) & (!g176) & (g197)) + ((g190) & (g155) & (!g162) & (!g169) & (g176) & (g197)) + ((g190) & (g155) & (!g162) & (g169) & (!g176) & (g197)) + ((g190) & (g155) & (!g162) & (g169) & (g176) & (!g197)) + ((g190) & (g155) & (g162) & (!g169) & (g176) & (!g197)) + ((g190) & (g155) & (g162) & (!g169) & (g176) & (g197)));
	assign g1323 = (((!g190) & (!g155) & (!g162) & (!g169) & (g176) & (!g197)) + ((!g190) & (!g155) & (!g162) & (g169) & (!g176) & (!g197)) + ((!g190) & (!g155) & (!g162) & (g169) & (g176) & (!g197)) + ((!g190) & (!g155) & (!g162) & (g169) & (g176) & (g197)) + ((!g190) & (!g155) & (g162) & (!g169) & (!g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (!g169) & (!g176) & (g197)) + ((!g190) & (!g155) & (g162) & (!g169) & (g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (g169) & (!g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (g169) & (g176) & (g197)) + ((!g190) & (g155) & (!g162) & (!g169) & (!g176) & (g197)) + ((!g190) & (g155) & (!g162) & (!g169) & (g176) & (!g197)) + ((!g190) & (g155) & (!g162) & (!g169) & (g176) & (g197)) + ((!g190) & (g155) & (g162) & (!g169) & (!g176) & (g197)) + ((!g190) & (g155) & (g162) & (!g169) & (g176) & (!g197)) + ((!g190) & (g155) & (g162) & (!g169) & (g176) & (g197)) + ((!g190) & (g155) & (g162) & (g169) & (!g176) & (!g197)) + ((g190) & (!g155) & (!g162) & (!g169) & (g176) & (!g197)) + ((g190) & (!g155) & (!g162) & (g169) & (!g176) & (!g197)) + ((g190) & (!g155) & (!g162) & (g169) & (g176) & (g197)) + ((g190) & (!g155) & (g162) & (!g169) & (!g176) & (!g197)) + ((g190) & (!g155) & (g162) & (!g169) & (!g176) & (g197)) + ((g190) & (!g155) & (g162) & (g169) & (!g176) & (!g197)) + ((g190) & (!g155) & (g162) & (g169) & (g176) & (!g197)) + ((g190) & (g155) & (!g162) & (!g169) & (g176) & (!g197)) + ((g190) & (g155) & (!g162) & (g169) & (!g176) & (!g197)) + ((g190) & (g155) & (!g162) & (g169) & (g176) & (g197)) + ((g190) & (g155) & (g162) & (!g169) & (!g176) & (!g197)) + ((g190) & (g155) & (g162) & (!g169) & (g176) & (!g197)) + ((g190) & (g155) & (g162) & (!g169) & (g176) & (g197)) + ((g190) & (g155) & (g162) & (g169) & (!g176) & (g197)));
	assign g1324 = (((!g190) & (!g155) & (!g162) & (!g169) & (!g176) & (g197)) + ((!g190) & (!g155) & (!g162) & (g169) & (g176) & (!g197)) + ((!g190) & (!g155) & (!g162) & (g169) & (g176) & (g197)) + ((!g190) & (!g155) & (g162) & (!g169) & (!g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (!g169) & (!g176) & (g197)) + ((!g190) & (!g155) & (g162) & (g169) & (g176) & (!g197)) + ((!g190) & (!g155) & (g162) & (g169) & (g176) & (g197)) + ((!g190) & (g155) & (!g162) & (!g169) & (!g176) & (!g197)) + ((!g190) & (g155) & (!g162) & (!g169) & (!g176) & (g197)) + ((!g190) & (g155) & (!g162) & (!g169) & (g176) & (g197)) + ((!g190) & (g155) & (!g162) & (g169) & (!g176) & (g197)) + ((!g190) & (g155) & (g162) & (!g169) & (!g176) & (g197)) + ((!g190) & (g155) & (g162) & (g169) & (!g176) & (!g197)) + ((!g190) & (g155) & (g162) & (g169) & (!g176) & (g197)) + ((!g190) & (g155) & (g162) & (g169) & (g176) & (!g197)) + ((!g190) & (g155) & (g162) & (g169) & (g176) & (g197)) + ((g190) & (!g155) & (!g162) & (g169) & (!g176) & (g197)) + ((g190) & (!g155) & (g162) & (!g169) & (!g176) & (!g197)) + ((g190) & (!g155) & (g162) & (g169) & (!g176) & (!g197)) + ((g190) & (!g155) & (g162) & (g169) & (!g176) & (g197)) + ((g190) & (!g155) & (g162) & (g169) & (g176) & (g197)) + ((g190) & (g155) & (!g162) & (!g169) & (!g176) & (g197)) + ((g190) & (g155) & (!g162) & (!g169) & (g176) & (g197)) + ((g190) & (g155) & (!g162) & (g169) & (!g176) & (!g197)) + ((g190) & (g155) & (!g162) & (g169) & (g176) & (!g197)) + ((g190) & (g155) & (!g162) & (g169) & (g176) & (g197)) + ((g190) & (g155) & (g162) & (!g169) & (g176) & (g197)) + ((g190) & (g155) & (g162) & (g169) & (g176) & (g197)));
	assign g1325 = (((!g1321) & (!g1322) & (!g1323) & (!g1324) & (!g148) & (g183)) + ((!g1321) & (!g1322) & (!g1323) & (!g1324) & (g148) & (!g183)) + ((!g1321) & (!g1322) & (!g1323) & (!g1324) & (g148) & (g183)) + ((!g1321) & (!g1322) & (!g1323) & (g1324) & (!g148) & (g183)) + ((!g1321) & (!g1322) & (!g1323) & (g1324) & (g148) & (!g183)) + ((!g1321) & (!g1322) & (g1323) & (!g1324) & (g148) & (!g183)) + ((!g1321) & (!g1322) & (g1323) & (!g1324) & (g148) & (g183)) + ((!g1321) & (!g1322) & (g1323) & (g1324) & (g148) & (!g183)) + ((!g1321) & (g1322) & (!g1323) & (!g1324) & (!g148) & (g183)) + ((!g1321) & (g1322) & (!g1323) & (!g1324) & (g148) & (g183)) + ((!g1321) & (g1322) & (!g1323) & (g1324) & (!g148) & (g183)) + ((!g1321) & (g1322) & (g1323) & (!g1324) & (g148) & (g183)) + ((g1321) & (!g1322) & (!g1323) & (!g1324) & (!g148) & (!g183)) + ((g1321) & (!g1322) & (!g1323) & (!g1324) & (!g148) & (g183)) + ((g1321) & (!g1322) & (!g1323) & (!g1324) & (g148) & (!g183)) + ((g1321) & (!g1322) & (!g1323) & (!g1324) & (g148) & (g183)) + ((g1321) & (!g1322) & (!g1323) & (g1324) & (!g148) & (!g183)) + ((g1321) & (!g1322) & (!g1323) & (g1324) & (!g148) & (g183)) + ((g1321) & (!g1322) & (!g1323) & (g1324) & (g148) & (!g183)) + ((g1321) & (!g1322) & (g1323) & (!g1324) & (!g148) & (!g183)) + ((g1321) & (!g1322) & (g1323) & (!g1324) & (g148) & (!g183)) + ((g1321) & (!g1322) & (g1323) & (!g1324) & (g148) & (g183)) + ((g1321) & (!g1322) & (g1323) & (g1324) & (!g148) & (!g183)) + ((g1321) & (!g1322) & (g1323) & (g1324) & (g148) & (!g183)) + ((g1321) & (g1322) & (!g1323) & (!g1324) & (!g148) & (!g183)) + ((g1321) & (g1322) & (!g1323) & (!g1324) & (!g148) & (g183)) + ((g1321) & (g1322) & (!g1323) & (!g1324) & (g148) & (g183)) + ((g1321) & (g1322) & (!g1323) & (g1324) & (!g148) & (!g183)) + ((g1321) & (g1322) & (!g1323) & (g1324) & (!g148) & (g183)) + ((g1321) & (g1322) & (g1323) & (!g1324) & (!g148) & (!g183)) + ((g1321) & (g1322) & (g1323) & (!g1324) & (g148) & (g183)) + ((g1321) & (g1322) & (g1323) & (g1324) & (!g148) & (!g183)));
	assign g1326 = (((!g517) & (!g773) & (!g1029) & (sk[39]) & (g1325)) + ((!g517) & (!g773) & (g1029) & (!sk[39]) & (!g1325)) + ((!g517) & (!g773) & (g1029) & (!sk[39]) & (g1325)) + ((!g517) & (!g773) & (g1029) & (sk[39]) & (!g1325)) + ((!g517) & (g773) & (!g1029) & (!sk[39]) & (!g1325)) + ((!g517) & (g773) & (!g1029) & (!sk[39]) & (g1325)) + ((!g517) & (g773) & (!g1029) & (sk[39]) & (!g1325)) + ((!g517) & (g773) & (g1029) & (!sk[39]) & (!g1325)) + ((!g517) & (g773) & (g1029) & (!sk[39]) & (g1325)) + ((!g517) & (g773) & (g1029) & (sk[39]) & (g1325)) + ((g517) & (!g773) & (!g1029) & (sk[39]) & (!g1325)) + ((g517) & (!g773) & (g1029) & (!sk[39]) & (!g1325)) + ((g517) & (!g773) & (g1029) & (!sk[39]) & (g1325)) + ((g517) & (!g773) & (g1029) & (sk[39]) & (g1325)) + ((g517) & (g773) & (!g1029) & (!sk[39]) & (!g1325)) + ((g517) & (g773) & (!g1029) & (!sk[39]) & (g1325)) + ((g517) & (g773) & (!g1029) & (sk[39]) & (g1325)) + ((g517) & (g773) & (g1029) & (!sk[39]) & (!g1325)) + ((g517) & (g773) & (g1029) & (!sk[39]) & (g1325)) + ((g517) & (g773) & (g1029) & (sk[39]) & (!g1325)));
	assign g1327 = (((!ld) & (!g261) & (g1326) & (!sk[40]) & (!keyx15x)) + ((!ld) & (!g261) & (g1326) & (!sk[40]) & (keyx15x)) + ((!ld) & (!g261) & (g1326) & (sk[40]) & (!keyx15x)) + ((!ld) & (!g261) & (g1326) & (sk[40]) & (keyx15x)) + ((!ld) & (g261) & (!g1326) & (!sk[40]) & (!keyx15x)) + ((!ld) & (g261) & (!g1326) & (!sk[40]) & (keyx15x)) + ((!ld) & (g261) & (!g1326) & (sk[40]) & (!keyx15x)) + ((!ld) & (g261) & (!g1326) & (sk[40]) & (keyx15x)) + ((!ld) & (g261) & (g1326) & (!sk[40]) & (!keyx15x)) + ((!ld) & (g261) & (g1326) & (!sk[40]) & (keyx15x)) + ((ld) & (!g261) & (!g1326) & (sk[40]) & (keyx15x)) + ((ld) & (!g261) & (g1326) & (!sk[40]) & (!keyx15x)) + ((ld) & (!g261) & (g1326) & (!sk[40]) & (keyx15x)) + ((ld) & (!g261) & (g1326) & (sk[40]) & (keyx15x)) + ((ld) & (g261) & (!g1326) & (!sk[40]) & (!keyx15x)) + ((ld) & (g261) & (!g1326) & (!sk[40]) & (keyx15x)) + ((ld) & (g261) & (!g1326) & (sk[40]) & (keyx15x)) + ((ld) & (g261) & (g1326) & (!sk[40]) & (!keyx15x)) + ((ld) & (g261) & (g1326) & (!sk[40]) & (keyx15x)) + ((ld) & (g261) & (g1326) & (sk[40]) & (keyx15x)));
	assign g2098 = (((!ld) & (!sk[41]) & (text_inx112x) & (!g1328)) + ((!ld) & (!sk[41]) & (text_inx112x) & (g1328)) + ((!ld) & (sk[41]) & (!text_inx112x) & (g1328)) + ((!ld) & (sk[41]) & (text_inx112x) & (g1328)) + ((ld) & (!sk[41]) & (!text_inx112x) & (g1328)) + ((ld) & (!sk[41]) & (text_inx112x) & (!g1328)) + ((ld) & (!sk[41]) & (text_inx112x) & (g1328)) + ((ld) & (sk[41]) & (text_inx112x) & (!g1328)) + ((ld) & (sk[41]) & (text_inx112x) & (g1328)));
	assign g1329 = (((!g1028) & (!sk[42]) & (g1092)) + ((!g1028) & (sk[42]) & (g1092)) + ((g1028) & (!sk[42]) & (g1092)) + ((g1028) & (sk[42]) & (!g1092)));
	assign g1330 = (((!g915) & (!sk[43]) & (g979)) + ((!g915) & (sk[43]) & (g979)) + ((g915) & (!sk[43]) & (g979)) + ((g915) & (sk[43]) & (!g979)));
	assign g1331 = (((!g1044) & (!g1107) & (!g1163) & (!g1328) & (!g1329) & (g1330)) + ((!g1044) & (!g1107) & (!g1163) & (!g1328) & (g1329) & (!g1330)) + ((!g1044) & (!g1107) & (!g1163) & (g1328) & (!g1329) & (g1330)) + ((!g1044) & (!g1107) & (!g1163) & (g1328) & (g1329) & (!g1330)) + ((!g1044) & (!g1107) & (g1163) & (g1328) & (!g1329) & (!g1330)) + ((!g1044) & (!g1107) & (g1163) & (g1328) & (!g1329) & (g1330)) + ((!g1044) & (!g1107) & (g1163) & (g1328) & (g1329) & (!g1330)) + ((!g1044) & (!g1107) & (g1163) & (g1328) & (g1329) & (g1330)) + ((!g1044) & (g1107) & (!g1163) & (!g1328) & (!g1329) & (!g1330)) + ((!g1044) & (g1107) & (!g1163) & (!g1328) & (g1329) & (g1330)) + ((!g1044) & (g1107) & (!g1163) & (g1328) & (!g1329) & (!g1330)) + ((!g1044) & (g1107) & (!g1163) & (g1328) & (g1329) & (g1330)) + ((!g1044) & (g1107) & (g1163) & (g1328) & (!g1329) & (!g1330)) + ((!g1044) & (g1107) & (g1163) & (g1328) & (!g1329) & (g1330)) + ((!g1044) & (g1107) & (g1163) & (g1328) & (g1329) & (!g1330)) + ((!g1044) & (g1107) & (g1163) & (g1328) & (g1329) & (g1330)) + ((g1044) & (!g1107) & (!g1163) & (!g1328) & (!g1329) & (!g1330)) + ((g1044) & (!g1107) & (!g1163) & (!g1328) & (g1329) & (g1330)) + ((g1044) & (!g1107) & (!g1163) & (g1328) & (!g1329) & (!g1330)) + ((g1044) & (!g1107) & (!g1163) & (g1328) & (g1329) & (g1330)) + ((g1044) & (!g1107) & (g1163) & (!g1328) & (!g1329) & (!g1330)) + ((g1044) & (!g1107) & (g1163) & (!g1328) & (!g1329) & (g1330)) + ((g1044) & (!g1107) & (g1163) & (!g1328) & (g1329) & (!g1330)) + ((g1044) & (!g1107) & (g1163) & (!g1328) & (g1329) & (g1330)) + ((g1044) & (g1107) & (!g1163) & (!g1328) & (!g1329) & (g1330)) + ((g1044) & (g1107) & (!g1163) & (!g1328) & (g1329) & (!g1330)) + ((g1044) & (g1107) & (!g1163) & (g1328) & (!g1329) & (g1330)) + ((g1044) & (g1107) & (!g1163) & (g1328) & (g1329) & (!g1330)) + ((g1044) & (g1107) & (g1163) & (!g1328) & (!g1329) & (!g1330)) + ((g1044) & (g1107) & (g1163) & (!g1328) & (!g1329) & (g1330)) + ((g1044) & (g1107) & (g1163) & (!g1328) & (g1329) & (!g1330)) + ((g1044) & (g1107) & (g1163) & (!g1328) & (g1329) & (g1330)));
	assign g2099 = (((!sk[45]) & (!ld) & (text_inx113x) & (!g1332)) + ((!sk[45]) & (!ld) & (text_inx113x) & (g1332)) + ((!sk[45]) & (ld) & (!text_inx113x) & (g1332)) + ((!sk[45]) & (ld) & (text_inx113x) & (!g1332)) + ((!sk[45]) & (ld) & (text_inx113x) & (g1332)) + ((sk[45]) & (!ld) & (!text_inx113x) & (g1332)) + ((sk[45]) & (!ld) & (text_inx113x) & (g1332)) + ((sk[45]) & (ld) & (text_inx113x) & (!g1332)) + ((sk[45]) & (ld) & (text_inx113x) & (g1332)));
	assign g1333 = (((!sk[46]) & (!g979) & (g1043)) + ((!sk[46]) & (g979) & (g1043)) + ((sk[46]) & (!g979) & (g1043)) + ((sk[46]) & (g979) & (!g1043)));
	assign g1334 = (((!sk[47]) & (!g922) & (!g986) & (g1051) & (!g1114)) + ((!sk[47]) & (!g922) & (!g986) & (g1051) & (g1114)) + ((!sk[47]) & (!g922) & (g986) & (!g1051) & (!g1114)) + ((!sk[47]) & (!g922) & (g986) & (!g1051) & (g1114)) + ((!sk[47]) & (!g922) & (g986) & (g1051) & (!g1114)) + ((!sk[47]) & (!g922) & (g986) & (g1051) & (g1114)) + ((!sk[47]) & (g922) & (!g986) & (g1051) & (!g1114)) + ((!sk[47]) & (g922) & (!g986) & (g1051) & (g1114)) + ((!sk[47]) & (g922) & (g986) & (!g1051) & (!g1114)) + ((!sk[47]) & (g922) & (g986) & (!g1051) & (g1114)) + ((!sk[47]) & (g922) & (g986) & (g1051) & (!g1114)) + ((!sk[47]) & (g922) & (g986) & (g1051) & (g1114)) + ((sk[47]) & (!g922) & (!g986) & (!g1051) & (g1114)) + ((sk[47]) & (!g922) & (!g986) & (g1051) & (!g1114)) + ((sk[47]) & (!g922) & (g986) & (!g1051) & (!g1114)) + ((sk[47]) & (!g922) & (g986) & (g1051) & (g1114)) + ((sk[47]) & (g922) & (!g986) & (!g1051) & (!g1114)) + ((sk[47]) & (g922) & (!g986) & (g1051) & (g1114)) + ((sk[47]) & (g922) & (g986) & (!g1051) & (g1114)) + ((sk[47]) & (g922) & (g986) & (g1051) & (!g1114)));
	assign g1335 = (((!g1051) & (!g1163) & (!g1329) & (!g1332) & (!g1333) & (g1334)) + ((!g1051) & (!g1163) & (!g1329) & (!g1332) & (g1333) & (!g1334)) + ((!g1051) & (!g1163) & (!g1329) & (g1332) & (!g1333) & (g1334)) + ((!g1051) & (!g1163) & (!g1329) & (g1332) & (g1333) & (!g1334)) + ((!g1051) & (!g1163) & (g1329) & (!g1332) & (!g1333) & (!g1334)) + ((!g1051) & (!g1163) & (g1329) & (!g1332) & (g1333) & (g1334)) + ((!g1051) & (!g1163) & (g1329) & (g1332) & (!g1333) & (!g1334)) + ((!g1051) & (!g1163) & (g1329) & (g1332) & (g1333) & (g1334)) + ((!g1051) & (g1163) & (!g1329) & (g1332) & (!g1333) & (!g1334)) + ((!g1051) & (g1163) & (!g1329) & (g1332) & (!g1333) & (g1334)) + ((!g1051) & (g1163) & (!g1329) & (g1332) & (g1333) & (!g1334)) + ((!g1051) & (g1163) & (!g1329) & (g1332) & (g1333) & (g1334)) + ((!g1051) & (g1163) & (g1329) & (g1332) & (!g1333) & (!g1334)) + ((!g1051) & (g1163) & (g1329) & (g1332) & (!g1333) & (g1334)) + ((!g1051) & (g1163) & (g1329) & (g1332) & (g1333) & (!g1334)) + ((!g1051) & (g1163) & (g1329) & (g1332) & (g1333) & (g1334)) + ((g1051) & (!g1163) & (!g1329) & (!g1332) & (!g1333) & (g1334)) + ((g1051) & (!g1163) & (!g1329) & (!g1332) & (g1333) & (!g1334)) + ((g1051) & (!g1163) & (!g1329) & (g1332) & (!g1333) & (g1334)) + ((g1051) & (!g1163) & (!g1329) & (g1332) & (g1333) & (!g1334)) + ((g1051) & (!g1163) & (g1329) & (!g1332) & (!g1333) & (!g1334)) + ((g1051) & (!g1163) & (g1329) & (!g1332) & (g1333) & (g1334)) + ((g1051) & (!g1163) & (g1329) & (g1332) & (!g1333) & (!g1334)) + ((g1051) & (!g1163) & (g1329) & (g1332) & (g1333) & (g1334)) + ((g1051) & (g1163) & (!g1329) & (!g1332) & (!g1333) & (!g1334)) + ((g1051) & (g1163) & (!g1329) & (!g1332) & (!g1333) & (g1334)) + ((g1051) & (g1163) & (!g1329) & (!g1332) & (g1333) & (!g1334)) + ((g1051) & (g1163) & (!g1329) & (!g1332) & (g1333) & (g1334)) + ((g1051) & (g1163) & (g1329) & (!g1332) & (!g1333) & (!g1334)) + ((g1051) & (g1163) & (g1329) & (!g1332) & (!g1333) & (g1334)) + ((g1051) & (g1163) & (g1329) & (!g1332) & (g1333) & (!g1334)) + ((g1051) & (g1163) & (g1329) & (!g1332) & (g1333) & (g1334)));
	assign g2100 = (((!ld) & (!sk[49]) & (text_inx114x) & (!g1336)) + ((!ld) & (!sk[49]) & (text_inx114x) & (g1336)) + ((!ld) & (sk[49]) & (!text_inx114x) & (g1336)) + ((!ld) & (sk[49]) & (text_inx114x) & (g1336)) + ((ld) & (!sk[49]) & (!text_inx114x) & (g1336)) + ((ld) & (!sk[49]) & (text_inx114x) & (!g1336)) + ((ld) & (!sk[49]) & (text_inx114x) & (g1336)) + ((ld) & (sk[49]) & (text_inx114x) & (!g1336)) + ((ld) & (sk[49]) & (text_inx114x) & (g1336)));
	assign g1337 = (((!g929) & (!sk[50]) & (g993) & (!g1050)) + ((!g929) & (!sk[50]) & (g993) & (g1050)) + ((!g929) & (sk[50]) & (!g993) & (g1050)) + ((!g929) & (sk[50]) & (g993) & (!g1050)) + ((g929) & (!sk[50]) & (!g993) & (g1050)) + ((g929) & (!sk[50]) & (g993) & (!g1050)) + ((g929) & (!sk[50]) & (g993) & (g1050)) + ((g929) & (sk[50]) & (!g993) & (!g1050)) + ((g929) & (sk[50]) & (g993) & (g1050)));
	assign g1338 = (((!g986) & (!g1058) & (!g1121) & (!g1163) & (!g1336) & (g1337)) + ((!g986) & (!g1058) & (!g1121) & (!g1163) & (g1336) & (g1337)) + ((!g986) & (!g1058) & (!g1121) & (g1163) & (g1336) & (!g1337)) + ((!g986) & (!g1058) & (!g1121) & (g1163) & (g1336) & (g1337)) + ((!g986) & (!g1058) & (g1121) & (!g1163) & (!g1336) & (!g1337)) + ((!g986) & (!g1058) & (g1121) & (!g1163) & (g1336) & (!g1337)) + ((!g986) & (!g1058) & (g1121) & (g1163) & (g1336) & (!g1337)) + ((!g986) & (!g1058) & (g1121) & (g1163) & (g1336) & (g1337)) + ((!g986) & (g1058) & (!g1121) & (!g1163) & (!g1336) & (!g1337)) + ((!g986) & (g1058) & (!g1121) & (!g1163) & (g1336) & (!g1337)) + ((!g986) & (g1058) & (!g1121) & (g1163) & (!g1336) & (!g1337)) + ((!g986) & (g1058) & (!g1121) & (g1163) & (!g1336) & (g1337)) + ((!g986) & (g1058) & (g1121) & (!g1163) & (!g1336) & (g1337)) + ((!g986) & (g1058) & (g1121) & (!g1163) & (g1336) & (g1337)) + ((!g986) & (g1058) & (g1121) & (g1163) & (!g1336) & (!g1337)) + ((!g986) & (g1058) & (g1121) & (g1163) & (!g1336) & (g1337)) + ((g986) & (!g1058) & (!g1121) & (!g1163) & (!g1336) & (!g1337)) + ((g986) & (!g1058) & (!g1121) & (!g1163) & (g1336) & (!g1337)) + ((g986) & (!g1058) & (!g1121) & (g1163) & (g1336) & (!g1337)) + ((g986) & (!g1058) & (!g1121) & (g1163) & (g1336) & (g1337)) + ((g986) & (!g1058) & (g1121) & (!g1163) & (!g1336) & (g1337)) + ((g986) & (!g1058) & (g1121) & (!g1163) & (g1336) & (g1337)) + ((g986) & (!g1058) & (g1121) & (g1163) & (g1336) & (!g1337)) + ((g986) & (!g1058) & (g1121) & (g1163) & (g1336) & (g1337)) + ((g986) & (g1058) & (!g1121) & (!g1163) & (!g1336) & (g1337)) + ((g986) & (g1058) & (!g1121) & (!g1163) & (g1336) & (g1337)) + ((g986) & (g1058) & (!g1121) & (g1163) & (!g1336) & (!g1337)) + ((g986) & (g1058) & (!g1121) & (g1163) & (!g1336) & (g1337)) + ((g986) & (g1058) & (g1121) & (!g1163) & (!g1336) & (!g1337)) + ((g986) & (g1058) & (g1121) & (!g1163) & (g1336) & (!g1337)) + ((g986) & (g1058) & (g1121) & (g1163) & (!g1336) & (!g1337)) + ((g986) & (g1058) & (g1121) & (g1163) & (!g1336) & (g1337)));
	assign g2101 = (((!ld) & (!sk[52]) & (text_inx115x) & (!g1339)) + ((!ld) & (!sk[52]) & (text_inx115x) & (g1339)) + ((!ld) & (sk[52]) & (!text_inx115x) & (g1339)) + ((!ld) & (sk[52]) & (text_inx115x) & (g1339)) + ((ld) & (!sk[52]) & (!text_inx115x) & (g1339)) + ((ld) & (!sk[52]) & (text_inx115x) & (!g1339)) + ((ld) & (!sk[52]) & (text_inx115x) & (g1339)) + ((ld) & (sk[52]) & (text_inx115x) & (!g1339)) + ((ld) & (sk[52]) & (text_inx115x) & (g1339)));
	assign g1340 = (((!g936) & (!sk[53]) & (!g1000) & (g1057) & (!g1092)) + ((!g936) & (!sk[53]) & (!g1000) & (g1057) & (g1092)) + ((!g936) & (!sk[53]) & (g1000) & (!g1057) & (!g1092)) + ((!g936) & (!sk[53]) & (g1000) & (!g1057) & (g1092)) + ((!g936) & (!sk[53]) & (g1000) & (g1057) & (!g1092)) + ((!g936) & (!sk[53]) & (g1000) & (g1057) & (g1092)) + ((!g936) & (sk[53]) & (!g1000) & (!g1057) & (g1092)) + ((!g936) & (sk[53]) & (!g1000) & (g1057) & (!g1092)) + ((!g936) & (sk[53]) & (g1000) & (!g1057) & (!g1092)) + ((!g936) & (sk[53]) & (g1000) & (g1057) & (g1092)) + ((g936) & (!sk[53]) & (!g1000) & (g1057) & (!g1092)) + ((g936) & (!sk[53]) & (!g1000) & (g1057) & (g1092)) + ((g936) & (!sk[53]) & (g1000) & (!g1057) & (!g1092)) + ((g936) & (!sk[53]) & (g1000) & (!g1057) & (g1092)) + ((g936) & (!sk[53]) & (g1000) & (g1057) & (!g1092)) + ((g936) & (!sk[53]) & (g1000) & (g1057) & (g1092)) + ((g936) & (sk[53]) & (!g1000) & (!g1057) & (!g1092)) + ((g936) & (sk[53]) & (!g1000) & (g1057) & (g1092)) + ((g936) & (sk[53]) & (g1000) & (!g1057) & (g1092)) + ((g936) & (sk[53]) & (g1000) & (g1057) & (!g1092)));
	assign g2102 = (((!ld) & (!sk[54]) & (text_inx118x) & (!g1341)) + ((!ld) & (!sk[54]) & (text_inx118x) & (g1341)) + ((!ld) & (sk[54]) & (!text_inx118x) & (g1341)) + ((!ld) & (sk[54]) & (text_inx118x) & (g1341)) + ((ld) & (!sk[54]) & (!text_inx118x) & (g1341)) + ((ld) & (!sk[54]) & (text_inx118x) & (!g1341)) + ((ld) & (!sk[54]) & (text_inx118x) & (g1341)) + ((ld) & (sk[54]) & (text_inx118x) & (!g1341)) + ((ld) & (sk[54]) & (text_inx118x) & (g1341)));
	assign g1342 = (((!g957) & (!g1021) & (sk[55]) & (g1078)) + ((!g957) & (g1021) & (!sk[55]) & (!g1078)) + ((!g957) & (g1021) & (!sk[55]) & (g1078)) + ((!g957) & (g1021) & (sk[55]) & (!g1078)) + ((g957) & (!g1021) & (!sk[55]) & (g1078)) + ((g957) & (!g1021) & (sk[55]) & (!g1078)) + ((g957) & (g1021) & (!sk[55]) & (!g1078)) + ((g957) & (g1021) & (!sk[55]) & (g1078)) + ((g957) & (g1021) & (sk[55]) & (g1078)));
	assign g1343 = (((!g1014) & (!g1086) & (!g1149) & (!g1163) & (!g1341) & (g1342)) + ((!g1014) & (!g1086) & (!g1149) & (!g1163) & (g1341) & (g1342)) + ((!g1014) & (!g1086) & (!g1149) & (g1163) & (g1341) & (!g1342)) + ((!g1014) & (!g1086) & (!g1149) & (g1163) & (g1341) & (g1342)) + ((!g1014) & (!g1086) & (g1149) & (!g1163) & (!g1341) & (!g1342)) + ((!g1014) & (!g1086) & (g1149) & (!g1163) & (g1341) & (!g1342)) + ((!g1014) & (!g1086) & (g1149) & (g1163) & (g1341) & (!g1342)) + ((!g1014) & (!g1086) & (g1149) & (g1163) & (g1341) & (g1342)) + ((!g1014) & (g1086) & (!g1149) & (!g1163) & (!g1341) & (!g1342)) + ((!g1014) & (g1086) & (!g1149) & (!g1163) & (g1341) & (!g1342)) + ((!g1014) & (g1086) & (!g1149) & (g1163) & (!g1341) & (!g1342)) + ((!g1014) & (g1086) & (!g1149) & (g1163) & (!g1341) & (g1342)) + ((!g1014) & (g1086) & (g1149) & (!g1163) & (!g1341) & (g1342)) + ((!g1014) & (g1086) & (g1149) & (!g1163) & (g1341) & (g1342)) + ((!g1014) & (g1086) & (g1149) & (g1163) & (!g1341) & (!g1342)) + ((!g1014) & (g1086) & (g1149) & (g1163) & (!g1341) & (g1342)) + ((g1014) & (!g1086) & (!g1149) & (!g1163) & (!g1341) & (!g1342)) + ((g1014) & (!g1086) & (!g1149) & (!g1163) & (g1341) & (!g1342)) + ((g1014) & (!g1086) & (!g1149) & (g1163) & (g1341) & (!g1342)) + ((g1014) & (!g1086) & (!g1149) & (g1163) & (g1341) & (g1342)) + ((g1014) & (!g1086) & (g1149) & (!g1163) & (!g1341) & (g1342)) + ((g1014) & (!g1086) & (g1149) & (!g1163) & (g1341) & (g1342)) + ((g1014) & (!g1086) & (g1149) & (g1163) & (g1341) & (!g1342)) + ((g1014) & (!g1086) & (g1149) & (g1163) & (g1341) & (g1342)) + ((g1014) & (g1086) & (!g1149) & (!g1163) & (!g1341) & (g1342)) + ((g1014) & (g1086) & (!g1149) & (!g1163) & (g1341) & (g1342)) + ((g1014) & (g1086) & (!g1149) & (g1163) & (!g1341) & (!g1342)) + ((g1014) & (g1086) & (!g1149) & (g1163) & (!g1341) & (g1342)) + ((g1014) & (g1086) & (g1149) & (!g1163) & (!g1341) & (!g1342)) + ((g1014) & (g1086) & (g1149) & (!g1163) & (g1341) & (!g1342)) + ((g1014) & (g1086) & (g1149) & (g1163) & (!g1341) & (!g1342)) + ((g1014) & (g1086) & (g1149) & (g1163) & (!g1341) & (g1342)));
	assign g2103 = (((!sk[57]) & (!ld) & (text_inx117x) & (!g1344)) + ((!sk[57]) & (!ld) & (text_inx117x) & (g1344)) + ((!sk[57]) & (ld) & (!text_inx117x) & (g1344)) + ((!sk[57]) & (ld) & (text_inx117x) & (!g1344)) + ((!sk[57]) & (ld) & (text_inx117x) & (g1344)) + ((sk[57]) & (!ld) & (!text_inx117x) & (g1344)) + ((sk[57]) & (!ld) & (text_inx117x) & (g1344)) + ((sk[57]) & (ld) & (text_inx117x) & (!g1344)) + ((sk[57]) & (ld) & (text_inx117x) & (g1344)));
	assign g1345 = (((!g950) & (!g1014) & (sk[58]) & (g1071)) + ((!g950) & (g1014) & (!sk[58]) & (!g1071)) + ((!g950) & (g1014) & (!sk[58]) & (g1071)) + ((!g950) & (g1014) & (sk[58]) & (!g1071)) + ((g950) & (!g1014) & (!sk[58]) & (g1071)) + ((g950) & (!g1014) & (sk[58]) & (!g1071)) + ((g950) & (g1014) & (!sk[58]) & (!g1071)) + ((g950) & (g1014) & (!sk[58]) & (g1071)) + ((g950) & (g1014) & (sk[58]) & (g1071)));
	assign g1346 = (((!g1007) & (!g1079) & (!g1142) & (!g1163) & (!g1344) & (g1345)) + ((!g1007) & (!g1079) & (!g1142) & (!g1163) & (g1344) & (g1345)) + ((!g1007) & (!g1079) & (!g1142) & (g1163) & (g1344) & (!g1345)) + ((!g1007) & (!g1079) & (!g1142) & (g1163) & (g1344) & (g1345)) + ((!g1007) & (!g1079) & (g1142) & (!g1163) & (!g1344) & (!g1345)) + ((!g1007) & (!g1079) & (g1142) & (!g1163) & (g1344) & (!g1345)) + ((!g1007) & (!g1079) & (g1142) & (g1163) & (g1344) & (!g1345)) + ((!g1007) & (!g1079) & (g1142) & (g1163) & (g1344) & (g1345)) + ((!g1007) & (g1079) & (!g1142) & (!g1163) & (!g1344) & (!g1345)) + ((!g1007) & (g1079) & (!g1142) & (!g1163) & (g1344) & (!g1345)) + ((!g1007) & (g1079) & (!g1142) & (g1163) & (!g1344) & (!g1345)) + ((!g1007) & (g1079) & (!g1142) & (g1163) & (!g1344) & (g1345)) + ((!g1007) & (g1079) & (g1142) & (!g1163) & (!g1344) & (g1345)) + ((!g1007) & (g1079) & (g1142) & (!g1163) & (g1344) & (g1345)) + ((!g1007) & (g1079) & (g1142) & (g1163) & (!g1344) & (!g1345)) + ((!g1007) & (g1079) & (g1142) & (g1163) & (!g1344) & (g1345)) + ((g1007) & (!g1079) & (!g1142) & (!g1163) & (!g1344) & (!g1345)) + ((g1007) & (!g1079) & (!g1142) & (!g1163) & (g1344) & (!g1345)) + ((g1007) & (!g1079) & (!g1142) & (g1163) & (g1344) & (!g1345)) + ((g1007) & (!g1079) & (!g1142) & (g1163) & (g1344) & (g1345)) + ((g1007) & (!g1079) & (g1142) & (!g1163) & (!g1344) & (g1345)) + ((g1007) & (!g1079) & (g1142) & (!g1163) & (g1344) & (g1345)) + ((g1007) & (!g1079) & (g1142) & (g1163) & (g1344) & (!g1345)) + ((g1007) & (!g1079) & (g1142) & (g1163) & (g1344) & (g1345)) + ((g1007) & (g1079) & (!g1142) & (!g1163) & (!g1344) & (g1345)) + ((g1007) & (g1079) & (!g1142) & (!g1163) & (g1344) & (g1345)) + ((g1007) & (g1079) & (!g1142) & (g1163) & (!g1344) & (!g1345)) + ((g1007) & (g1079) & (!g1142) & (g1163) & (!g1344) & (g1345)) + ((g1007) & (g1079) & (g1142) & (!g1163) & (!g1344) & (!g1345)) + ((g1007) & (g1079) & (g1142) & (!g1163) & (g1344) & (!g1345)) + ((g1007) & (g1079) & (g1142) & (g1163) & (!g1344) & (!g1345)) + ((g1007) & (g1079) & (g1142) & (g1163) & (!g1344) & (g1345)));
	assign g2104 = (((!ld) & (!sk[60]) & (text_inx116x) & (!g1347)) + ((!ld) & (!sk[60]) & (text_inx116x) & (g1347)) + ((!ld) & (sk[60]) & (!text_inx116x) & (g1347)) + ((!ld) & (sk[60]) & (text_inx116x) & (g1347)) + ((ld) & (!sk[60]) & (!text_inx116x) & (g1347)) + ((ld) & (!sk[60]) & (text_inx116x) & (!g1347)) + ((ld) & (!sk[60]) & (text_inx116x) & (g1347)) + ((ld) & (sk[60]) & (text_inx116x) & (!g1347)) + ((ld) & (sk[60]) & (text_inx116x) & (g1347)));
	assign g1348 = (((!g943) & (!g1000) & (sk[61]) & (g1135)) + ((!g943) & (g1000) & (!sk[61]) & (!g1135)) + ((!g943) & (g1000) & (!sk[61]) & (g1135)) + ((!g943) & (g1000) & (sk[61]) & (!g1135)) + ((g943) & (!g1000) & (!sk[61]) & (g1135)) + ((g943) & (!g1000) & (sk[61]) & (!g1135)) + ((g943) & (g1000) & (!sk[61]) & (!g1135)) + ((g943) & (g1000) & (!sk[61]) & (g1135)) + ((g943) & (g1000) & (sk[61]) & (g1135)));
	assign g1349 = (((!g1007) & (!g1028) & (!g1064) & (!g1072) & (sk[62]) & (g1092)) + ((!g1007) & (!g1028) & (!g1064) & (g1072) & (sk[62]) & (!g1092)) + ((!g1007) & (!g1028) & (g1064) & (!g1072) & (sk[62]) & (!g1092)) + ((!g1007) & (!g1028) & (g1064) & (g1072) & (sk[62]) & (g1092)) + ((!g1007) & (g1028) & (!g1064) & (!g1072) & (!sk[62]) & (!g1092)) + ((!g1007) & (g1028) & (!g1064) & (!g1072) & (!sk[62]) & (g1092)) + ((!g1007) & (g1028) & (!g1064) & (!g1072) & (sk[62]) & (!g1092)) + ((!g1007) & (g1028) & (!g1064) & (g1072) & (!sk[62]) & (!g1092)) + ((!g1007) & (g1028) & (!g1064) & (g1072) & (!sk[62]) & (g1092)) + ((!g1007) & (g1028) & (!g1064) & (g1072) & (sk[62]) & (g1092)) + ((!g1007) & (g1028) & (g1064) & (!g1072) & (!sk[62]) & (!g1092)) + ((!g1007) & (g1028) & (g1064) & (!g1072) & (!sk[62]) & (g1092)) + ((!g1007) & (g1028) & (g1064) & (!g1072) & (sk[62]) & (g1092)) + ((!g1007) & (g1028) & (g1064) & (g1072) & (!sk[62]) & (!g1092)) + ((!g1007) & (g1028) & (g1064) & (g1072) & (!sk[62]) & (g1092)) + ((!g1007) & (g1028) & (g1064) & (g1072) & (sk[62]) & (!g1092)) + ((g1007) & (!g1028) & (!g1064) & (!g1072) & (!sk[62]) & (!g1092)) + ((g1007) & (!g1028) & (!g1064) & (!g1072) & (!sk[62]) & (g1092)) + ((g1007) & (!g1028) & (!g1064) & (!g1072) & (sk[62]) & (!g1092)) + ((g1007) & (!g1028) & (!g1064) & (g1072) & (!sk[62]) & (!g1092)) + ((g1007) & (!g1028) & (!g1064) & (g1072) & (!sk[62]) & (g1092)) + ((g1007) & (!g1028) & (!g1064) & (g1072) & (sk[62]) & (g1092)) + ((g1007) & (!g1028) & (g1064) & (!g1072) & (!sk[62]) & (!g1092)) + ((g1007) & (!g1028) & (g1064) & (!g1072) & (!sk[62]) & (g1092)) + ((g1007) & (!g1028) & (g1064) & (!g1072) & (sk[62]) & (g1092)) + ((g1007) & (!g1028) & (g1064) & (g1072) & (!sk[62]) & (!g1092)) + ((g1007) & (!g1028) & (g1064) & (g1072) & (!sk[62]) & (g1092)) + ((g1007) & (!g1028) & (g1064) & (g1072) & (sk[62]) & (!g1092)) + ((g1007) & (g1028) & (!g1064) & (!g1072) & (!sk[62]) & (!g1092)) + ((g1007) & (g1028) & (!g1064) & (!g1072) & (!sk[62]) & (g1092)) + ((g1007) & (g1028) & (!g1064) & (!g1072) & (sk[62]) & (g1092)) + ((g1007) & (g1028) & (!g1064) & (g1072) & (!sk[62]) & (!g1092)) + ((g1007) & (g1028) & (!g1064) & (g1072) & (!sk[62]) & (g1092)) + ((g1007) & (g1028) & (!g1064) & (g1072) & (sk[62]) & (!g1092)) + ((g1007) & (g1028) & (g1064) & (!g1072) & (!sk[62]) & (!g1092)) + ((g1007) & (g1028) & (g1064) & (!g1072) & (!sk[62]) & (g1092)) + ((g1007) & (g1028) & (g1064) & (!g1072) & (sk[62]) & (!g1092)) + ((g1007) & (g1028) & (g1064) & (g1072) & (!sk[62]) & (!g1092)) + ((g1007) & (g1028) & (g1064) & (g1072) & (!sk[62]) & (g1092)) + ((g1007) & (g1028) & (g1064) & (g1072) & (sk[62]) & (g1092)));
	assign g1350 = (((!sk[63]) & (!g1072) & (g1163) & (!g1347) & (!g1348) & (!g1349)) + ((!sk[63]) & (!g1072) & (g1163) & (!g1347) & (!g1348) & (g1349)) + ((!sk[63]) & (!g1072) & (g1163) & (!g1347) & (g1348) & (!g1349)) + ((!sk[63]) & (!g1072) & (g1163) & (!g1347) & (g1348) & (g1349)) + ((!sk[63]) & (!g1072) & (g1163) & (g1347) & (!g1348) & (!g1349)) + ((!sk[63]) & (!g1072) & (g1163) & (g1347) & (!g1348) & (g1349)) + ((!sk[63]) & (!g1072) & (g1163) & (g1347) & (g1348) & (!g1349)) + ((!sk[63]) & (!g1072) & (g1163) & (g1347) & (g1348) & (g1349)) + ((!sk[63]) & (g1072) & (!g1163) & (!g1347) & (!g1348) & (!g1349)) + ((!sk[63]) & (g1072) & (!g1163) & (!g1347) & (!g1348) & (g1349)) + ((!sk[63]) & (g1072) & (!g1163) & (!g1347) & (g1348) & (!g1349)) + ((!sk[63]) & (g1072) & (!g1163) & (!g1347) & (g1348) & (g1349)) + ((!sk[63]) & (g1072) & (!g1163) & (g1347) & (!g1348) & (!g1349)) + ((!sk[63]) & (g1072) & (!g1163) & (g1347) & (!g1348) & (g1349)) + ((!sk[63]) & (g1072) & (!g1163) & (g1347) & (g1348) & (!g1349)) + ((!sk[63]) & (g1072) & (!g1163) & (g1347) & (g1348) & (g1349)) + ((!sk[63]) & (g1072) & (g1163) & (!g1347) & (!g1348) & (!g1349)) + ((!sk[63]) & (g1072) & (g1163) & (!g1347) & (!g1348) & (g1349)) + ((!sk[63]) & (g1072) & (g1163) & (!g1347) & (g1348) & (!g1349)) + ((!sk[63]) & (g1072) & (g1163) & (!g1347) & (g1348) & (g1349)) + ((!sk[63]) & (g1072) & (g1163) & (g1347) & (!g1348) & (!g1349)) + ((!sk[63]) & (g1072) & (g1163) & (g1347) & (!g1348) & (g1349)) + ((!sk[63]) & (g1072) & (g1163) & (g1347) & (g1348) & (!g1349)) + ((!sk[63]) & (g1072) & (g1163) & (g1347) & (g1348) & (g1349)) + ((sk[63]) & (!g1072) & (!g1163) & (!g1347) & (!g1348) & (g1349)) + ((sk[63]) & (!g1072) & (!g1163) & (!g1347) & (g1348) & (!g1349)) + ((sk[63]) & (!g1072) & (!g1163) & (g1347) & (!g1348) & (g1349)) + ((sk[63]) & (!g1072) & (!g1163) & (g1347) & (g1348) & (!g1349)) + ((sk[63]) & (!g1072) & (g1163) & (g1347) & (!g1348) & (!g1349)) + ((sk[63]) & (!g1072) & (g1163) & (g1347) & (!g1348) & (g1349)) + ((sk[63]) & (!g1072) & (g1163) & (g1347) & (g1348) & (!g1349)) + ((sk[63]) & (!g1072) & (g1163) & (g1347) & (g1348) & (g1349)) + ((sk[63]) & (g1072) & (!g1163) & (!g1347) & (!g1348) & (g1349)) + ((sk[63]) & (g1072) & (!g1163) & (!g1347) & (g1348) & (!g1349)) + ((sk[63]) & (g1072) & (!g1163) & (g1347) & (!g1348) & (g1349)) + ((sk[63]) & (g1072) & (!g1163) & (g1347) & (g1348) & (!g1349)) + ((sk[63]) & (g1072) & (g1163) & (!g1347) & (!g1348) & (!g1349)) + ((sk[63]) & (g1072) & (g1163) & (!g1347) & (!g1348) & (g1349)) + ((sk[63]) & (g1072) & (g1163) & (!g1347) & (g1348) & (!g1349)) + ((sk[63]) & (g1072) & (g1163) & (!g1347) & (g1348) & (g1349)));
	assign g2105 = (((!ld) & (!sk[64]) & (text_inx119x) & (!g1351)) + ((!ld) & (!sk[64]) & (text_inx119x) & (g1351)) + ((!ld) & (sk[64]) & (!text_inx119x) & (g1351)) + ((!ld) & (sk[64]) & (text_inx119x) & (g1351)) + ((ld) & (!sk[64]) & (!text_inx119x) & (g1351)) + ((ld) & (!sk[64]) & (text_inx119x) & (!g1351)) + ((ld) & (!sk[64]) & (text_inx119x) & (g1351)) + ((ld) & (sk[64]) & (text_inx119x) & (!g1351)) + ((ld) & (sk[64]) & (text_inx119x) & (g1351)));
	assign g1352 = (((!g964) & (!sk[65]) & (g1021) & (!g1156)) + ((!g964) & (!sk[65]) & (g1021) & (g1156)) + ((!g964) & (sk[65]) & (!g1021) & (g1156)) + ((!g964) & (sk[65]) & (g1021) & (!g1156)) + ((g964) & (!sk[65]) & (!g1021) & (g1156)) + ((g964) & (!sk[65]) & (g1021) & (!g1156)) + ((g964) & (!sk[65]) & (g1021) & (g1156)) + ((g964) & (sk[65]) & (!g1021) & (!g1156)) + ((g964) & (sk[65]) & (g1021) & (g1156)));
	assign g1353 = (((!g1028) & (!g1085) & (!g1093) & (!g1163) & (!g1351) & (g1352)) + ((!g1028) & (!g1085) & (!g1093) & (!g1163) & (g1351) & (g1352)) + ((!g1028) & (!g1085) & (!g1093) & (g1163) & (g1351) & (!g1352)) + ((!g1028) & (!g1085) & (!g1093) & (g1163) & (g1351) & (g1352)) + ((!g1028) & (!g1085) & (g1093) & (!g1163) & (!g1351) & (!g1352)) + ((!g1028) & (!g1085) & (g1093) & (!g1163) & (g1351) & (!g1352)) + ((!g1028) & (!g1085) & (g1093) & (g1163) & (!g1351) & (!g1352)) + ((!g1028) & (!g1085) & (g1093) & (g1163) & (!g1351) & (g1352)) + ((!g1028) & (g1085) & (!g1093) & (!g1163) & (!g1351) & (!g1352)) + ((!g1028) & (g1085) & (!g1093) & (!g1163) & (g1351) & (!g1352)) + ((!g1028) & (g1085) & (!g1093) & (g1163) & (g1351) & (!g1352)) + ((!g1028) & (g1085) & (!g1093) & (g1163) & (g1351) & (g1352)) + ((!g1028) & (g1085) & (g1093) & (!g1163) & (!g1351) & (g1352)) + ((!g1028) & (g1085) & (g1093) & (!g1163) & (g1351) & (g1352)) + ((!g1028) & (g1085) & (g1093) & (g1163) & (!g1351) & (!g1352)) + ((!g1028) & (g1085) & (g1093) & (g1163) & (!g1351) & (g1352)) + ((g1028) & (!g1085) & (!g1093) & (!g1163) & (!g1351) & (!g1352)) + ((g1028) & (!g1085) & (!g1093) & (!g1163) & (g1351) & (!g1352)) + ((g1028) & (!g1085) & (!g1093) & (g1163) & (g1351) & (!g1352)) + ((g1028) & (!g1085) & (!g1093) & (g1163) & (g1351) & (g1352)) + ((g1028) & (!g1085) & (g1093) & (!g1163) & (!g1351) & (g1352)) + ((g1028) & (!g1085) & (g1093) & (!g1163) & (g1351) & (g1352)) + ((g1028) & (!g1085) & (g1093) & (g1163) & (!g1351) & (!g1352)) + ((g1028) & (!g1085) & (g1093) & (g1163) & (!g1351) & (g1352)) + ((g1028) & (g1085) & (!g1093) & (!g1163) & (!g1351) & (g1352)) + ((g1028) & (g1085) & (!g1093) & (!g1163) & (g1351) & (g1352)) + ((g1028) & (g1085) & (!g1093) & (g1163) & (g1351) & (!g1352)) + ((g1028) & (g1085) & (!g1093) & (g1163) & (g1351) & (g1352)) + ((g1028) & (g1085) & (g1093) & (!g1163) & (!g1351) & (!g1352)) + ((g1028) & (g1085) & (g1093) & (!g1163) & (g1351) & (!g1352)) + ((g1028) & (g1085) & (g1093) & (g1163) & (!g1351) & (!g1352)) + ((g1028) & (g1085) & (g1093) & (g1163) & (!g1351) & (g1352)));
	assign g1354 = (((!g212) & (!g219) & (!g226) & (!g233) & (g254) & (g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g254) & (!g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g254) & (g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (g254) & (!g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (!g254) & (!g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (!g254) & (g247)) + ((!g212) & (!g219) & (g226) & (g233) & (!g254) & (!g247)) + ((!g212) & (!g219) & (g226) & (g233) & (g254) & (g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (g254) & (!g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (g254) & (g247)) + ((!g212) & (g219) & (!g226) & (g233) & (g254) & (!g247)) + ((!g212) & (g219) & (!g226) & (g233) & (g254) & (g247)) + ((!g212) & (g219) & (g226) & (!g233) & (g254) & (!g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (!g254) & (!g247)) + ((g212) & (!g219) & (g226) & (!g233) & (g254) & (!g247)) + ((g212) & (!g219) & (g226) & (g233) & (!g254) & (g247)) + ((g212) & (!g219) & (g226) & (g233) & (g254) & (g247)) + ((g212) & (g219) & (!g226) & (!g233) & (!g254) & (g247)) + ((g212) & (g219) & (!g226) & (!g233) & (g254) & (!g247)) + ((g212) & (g219) & (g226) & (!g233) & (!g254) & (g247)) + ((g212) & (g219) & (g226) & (!g233) & (g254) & (!g247)) + ((g212) & (g219) & (g226) & (g233) & (!g254) & (!g247)) + ((g212) & (g219) & (g226) & (g233) & (g254) & (!g247)) + ((g212) & (g219) & (g226) & (g233) & (g254) & (g247)));
	assign g1355 = (((!g212) & (!g219) & (!g226) & (!g233) & (g254) & (!g247)) + ((!g212) & (!g219) & (!g226) & (!g233) & (g254) & (g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g254) & (!g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g254) & (g247)) + ((!g212) & (!g219) & (g226) & (g233) & (!g254) & (g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (!g254) & (!g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (!g254) & (g247)) + ((!g212) & (g219) & (g226) & (!g233) & (!g254) & (!g247)) + ((!g212) & (g219) & (g226) & (!g233) & (!g254) & (g247)) + ((!g212) & (g219) & (g226) & (!g233) & (g254) & (!g247)) + ((!g212) & (g219) & (g226) & (g233) & (g254) & (g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (!g254) & (g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (g254) & (!g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (g254) & (g247)) + ((g212) & (!g219) & (!g226) & (g233) & (g254) & (!g247)) + ((g212) & (!g219) & (g226) & (!g233) & (!g254) & (!g247)) + ((g212) & (!g219) & (g226) & (!g233) & (g254) & (g247)) + ((g212) & (!g219) & (g226) & (g233) & (!g254) & (g247)) + ((g212) & (!g219) & (g226) & (g233) & (g254) & (g247)) + ((g212) & (g219) & (!g226) & (!g233) & (!g254) & (!g247)) + ((g212) & (g219) & (!g226) & (!g233) & (!g254) & (g247)) + ((g212) & (g219) & (!g226) & (!g233) & (g254) & (!g247)) + ((g212) & (g219) & (!g226) & (!g233) & (g254) & (g247)) + ((g212) & (g219) & (!g226) & (g233) & (!g254) & (!g247)) + ((g212) & (g219) & (!g226) & (g233) & (g254) & (!g247)) + ((g212) & (g219) & (!g226) & (g233) & (g254) & (g247)) + ((g212) & (g219) & (g226) & (!g233) & (g254) & (!g247)) + ((g212) & (g219) & (g226) & (!g233) & (g254) & (g247)) + ((g212) & (g219) & (g226) & (g233) & (!g254) & (g247)) + ((g212) & (g219) & (g226) & (g233) & (g254) & (!g247)));
	assign g1356 = (((!g212) & (!g219) & (!g226) & (!g233) & (!g254) & (!g247)) + ((!g212) & (!g219) & (!g226) & (!g233) & (g254) & (g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (g254) & (g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (!g254) & (!g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (!g254) & (g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (g254) & (g247)) + ((!g212) & (!g219) & (g226) & (g233) & (!g254) & (g247)) + ((!g212) & (!g219) & (g226) & (g233) & (g254) & (!g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (!g254) & (!g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (g254) & (!g247)) + ((!g212) & (g219) & (!g226) & (g233) & (g254) & (g247)) + ((!g212) & (g219) & (g226) & (g233) & (!g254) & (!g247)) + ((!g212) & (g219) & (g226) & (g233) & (g254) & (!g247)) + ((g212) & (!g219) & (!g226) & (g233) & (!g254) & (!g247)) + ((g212) & (!g219) & (!g226) & (g233) & (!g254) & (g247)) + ((g212) & (!g219) & (!g226) & (g233) & (g254) & (!g247)) + ((g212) & (!g219) & (g226) & (!g233) & (!g254) & (!g247)) + ((g212) & (!g219) & (g226) & (!g233) & (g254) & (g247)) + ((g212) & (!g219) & (g226) & (g233) & (!g254) & (!g247)) + ((g212) & (!g219) & (g226) & (g233) & (!g254) & (g247)) + ((g212) & (!g219) & (g226) & (g233) & (g254) & (!g247)) + ((g212) & (!g219) & (g226) & (g233) & (g254) & (g247)) + ((g212) & (g219) & (!g226) & (!g233) & (g254) & (g247)) + ((g212) & (g219) & (!g226) & (g233) & (!g254) & (!g247)) + ((g212) & (g219) & (!g226) & (g233) & (g254) & (!g247)) + ((g212) & (g219) & (!g226) & (g233) & (g254) & (g247)) + ((g212) & (g219) & (g226) & (!g233) & (!g254) & (!g247)) + ((g212) & (g219) & (g226) & (g233) & (!g254) & (!g247)) + ((g212) & (g219) & (g226) & (g233) & (!g254) & (g247)) + ((g212) & (g219) & (g226) & (g233) & (g254) & (g247)));
	assign g1357 = (((!g212) & (!g219) & (!g226) & (!g233) & (!g254) & (g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (g254) & (!g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (g254) & (g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (!g254) & (g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (g254) & (g247)) + ((!g212) & (!g219) & (g226) & (g233) & (!g254) & (g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (!g254) & (!g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (!g254) & (g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (g254) & (!g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (g254) & (g247)) + ((!g212) & (g219) & (!g226) & (g233) & (g254) & (!g247)) + ((!g212) & (g219) & (!g226) & (g233) & (g254) & (g247)) + ((!g212) & (g219) & (g226) & (g233) & (!g254) & (!g247)) + ((!g212) & (g219) & (g226) & (g233) & (g254) & (!g247)) + ((!g212) & (g219) & (g226) & (g233) & (g254) & (g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (!g254) & (!g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (g254) & (g247)) + ((g212) & (!g219) & (!g226) & (g233) & (g254) & (!g247)) + ((g212) & (!g219) & (!g226) & (g233) & (g254) & (g247)) + ((g212) & (!g219) & (g226) & (!g233) & (!g254) & (g247)) + ((g212) & (!g219) & (g226) & (!g233) & (g254) & (!g247)) + ((g212) & (!g219) & (g226) & (g233) & (g254) & (!g247)) + ((g212) & (g219) & (!g226) & (!g233) & (!g254) & (g247)) + ((g212) & (g219) & (!g226) & (!g233) & (g254) & (g247)) + ((g212) & (g219) & (!g226) & (g233) & (g254) & (!g247)) + ((g212) & (g219) & (!g226) & (g233) & (g254) & (g247)) + ((g212) & (g219) & (g226) & (!g233) & (!g254) & (g247)) + ((g212) & (g219) & (g226) & (g233) & (!g254) & (!g247)));
	assign g1358 = (((!g1354) & (!g1355) & (!g1356) & (!g1357) & (!g240) & (!g261)) + ((!g1354) & (!g1355) & (!g1356) & (g1357) & (!g240) & (!g261)) + ((!g1354) & (!g1355) & (!g1356) & (g1357) & (g240) & (g261)) + ((!g1354) & (!g1355) & (g1356) & (!g1357) & (!g240) & (!g261)) + ((!g1354) & (!g1355) & (g1356) & (!g1357) & (!g240) & (g261)) + ((!g1354) & (!g1355) & (g1356) & (g1357) & (!g240) & (!g261)) + ((!g1354) & (!g1355) & (g1356) & (g1357) & (!g240) & (g261)) + ((!g1354) & (!g1355) & (g1356) & (g1357) & (g240) & (g261)) + ((!g1354) & (g1355) & (!g1356) & (!g1357) & (!g240) & (!g261)) + ((!g1354) & (g1355) & (!g1356) & (!g1357) & (g240) & (!g261)) + ((!g1354) & (g1355) & (!g1356) & (g1357) & (!g240) & (!g261)) + ((!g1354) & (g1355) & (!g1356) & (g1357) & (g240) & (!g261)) + ((!g1354) & (g1355) & (!g1356) & (g1357) & (g240) & (g261)) + ((!g1354) & (g1355) & (g1356) & (!g1357) & (!g240) & (!g261)) + ((!g1354) & (g1355) & (g1356) & (!g1357) & (!g240) & (g261)) + ((!g1354) & (g1355) & (g1356) & (!g1357) & (g240) & (!g261)) + ((!g1354) & (g1355) & (g1356) & (g1357) & (!g240) & (!g261)) + ((!g1354) & (g1355) & (g1356) & (g1357) & (!g240) & (g261)) + ((!g1354) & (g1355) & (g1356) & (g1357) & (g240) & (!g261)) + ((!g1354) & (g1355) & (g1356) & (g1357) & (g240) & (g261)) + ((g1354) & (!g1355) & (!g1356) & (g1357) & (g240) & (g261)) + ((g1354) & (!g1355) & (g1356) & (!g1357) & (!g240) & (g261)) + ((g1354) & (!g1355) & (g1356) & (g1357) & (!g240) & (g261)) + ((g1354) & (!g1355) & (g1356) & (g1357) & (g240) & (g261)) + ((g1354) & (g1355) & (!g1356) & (!g1357) & (g240) & (!g261)) + ((g1354) & (g1355) & (!g1356) & (g1357) & (g240) & (!g261)) + ((g1354) & (g1355) & (!g1356) & (g1357) & (g240) & (g261)) + ((g1354) & (g1355) & (g1356) & (!g1357) & (!g240) & (g261)) + ((g1354) & (g1355) & (g1356) & (!g1357) & (g240) & (!g261)) + ((g1354) & (g1355) & (g1356) & (g1357) & (!g240) & (g261)) + ((g1354) & (g1355) & (g1356) & (g1357) & (g240) & (!g261)) + ((g1354) & (g1355) & (g1356) & (g1357) & (g240) & (g261)));
	assign g1359 = (((!g532) & (!sk[72]) & (!g788) & (g1044) & (!g1358)) + ((!g532) & (!sk[72]) & (!g788) & (g1044) & (g1358)) + ((!g532) & (!sk[72]) & (g788) & (!g1044) & (!g1358)) + ((!g532) & (!sk[72]) & (g788) & (!g1044) & (g1358)) + ((!g532) & (!sk[72]) & (g788) & (g1044) & (!g1358)) + ((!g532) & (!sk[72]) & (g788) & (g1044) & (g1358)) + ((!g532) & (sk[72]) & (!g788) & (!g1044) & (g1358)) + ((!g532) & (sk[72]) & (!g788) & (g1044) & (!g1358)) + ((!g532) & (sk[72]) & (g788) & (!g1044) & (!g1358)) + ((!g532) & (sk[72]) & (g788) & (g1044) & (g1358)) + ((g532) & (!sk[72]) & (!g788) & (g1044) & (!g1358)) + ((g532) & (!sk[72]) & (!g788) & (g1044) & (g1358)) + ((g532) & (!sk[72]) & (g788) & (!g1044) & (!g1358)) + ((g532) & (!sk[72]) & (g788) & (!g1044) & (g1358)) + ((g532) & (!sk[72]) & (g788) & (g1044) & (!g1358)) + ((g532) & (!sk[72]) & (g788) & (g1044) & (g1358)) + ((g532) & (sk[72]) & (!g788) & (!g1044) & (!g1358)) + ((g532) & (sk[72]) & (!g788) & (g1044) & (g1358)) + ((g532) & (sk[72]) & (g788) & (!g1044) & (g1358)) + ((g532) & (sk[72]) & (g788) & (g1044) & (!g1358)));
	assign g1360 = (((!sk[73]) & (!ld) & (!g276) & (g1359) & (!keyx16x)) + ((!sk[73]) & (!ld) & (!g276) & (g1359) & (keyx16x)) + ((!sk[73]) & (!ld) & (g276) & (!g1359) & (!keyx16x)) + ((!sk[73]) & (!ld) & (g276) & (!g1359) & (keyx16x)) + ((!sk[73]) & (!ld) & (g276) & (g1359) & (!keyx16x)) + ((!sk[73]) & (!ld) & (g276) & (g1359) & (keyx16x)) + ((!sk[73]) & (ld) & (!g276) & (g1359) & (!keyx16x)) + ((!sk[73]) & (ld) & (!g276) & (g1359) & (keyx16x)) + ((!sk[73]) & (ld) & (g276) & (!g1359) & (!keyx16x)) + ((!sk[73]) & (ld) & (g276) & (!g1359) & (keyx16x)) + ((!sk[73]) & (ld) & (g276) & (g1359) & (!keyx16x)) + ((!sk[73]) & (ld) & (g276) & (g1359) & (keyx16x)) + ((sk[73]) & (!ld) & (!g276) & (g1359) & (!keyx16x)) + ((sk[73]) & (!ld) & (!g276) & (g1359) & (keyx16x)) + ((sk[73]) & (!ld) & (g276) & (!g1359) & (!keyx16x)) + ((sk[73]) & (!ld) & (g276) & (!g1359) & (keyx16x)) + ((sk[73]) & (ld) & (!g276) & (!g1359) & (keyx16x)) + ((sk[73]) & (ld) & (!g276) & (g1359) & (keyx16x)) + ((sk[73]) & (ld) & (g276) & (!g1359) & (keyx16x)) + ((sk[73]) & (ld) & (g276) & (g1359) & (keyx16x)));
	assign g1361 = (((!g212) & (!g219) & (!g226) & (!g233) & (!g240) & (g254)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g240) & (!g254)) + ((!g212) & (!g219) & (!g226) & (g233) & (g240) & (!g254)) + ((!g212) & (!g219) & (g226) & (!g233) & (g240) & (g254)) + ((!g212) & (!g219) & (g226) & (g233) & (!g240) & (g254)) + ((!g212) & (!g219) & (g226) & (g233) & (g240) & (!g254)) + ((!g212) & (g219) & (!g226) & (!g233) & (!g240) & (g254)) + ((!g212) & (g219) & (!g226) & (!g233) & (g240) & (!g254)) + ((!g212) & (g219) & (!g226) & (!g233) & (g240) & (g254)) + ((!g212) & (g219) & (g226) & (!g233) & (g240) & (g254)) + ((!g212) & (g219) & (g226) & (g233) & (g240) & (g254)) + ((g212) & (!g219) & (!g226) & (!g233) & (!g240) & (!g254)) + ((g212) & (!g219) & (!g226) & (!g233) & (g240) & (g254)) + ((g212) & (!g219) & (!g226) & (g233) & (!g240) & (!g254)) + ((g212) & (!g219) & (!g226) & (g233) & (g240) & (!g254)) + ((g212) & (!g219) & (g226) & (!g233) & (g240) & (!g254)) + ((g212) & (!g219) & (g226) & (!g233) & (g240) & (g254)) + ((g212) & (!g219) & (g226) & (g233) & (g240) & (!g254)) + ((g212) & (!g219) & (g226) & (g233) & (g240) & (g254)) + ((g212) & (g219) & (!g226) & (!g233) & (g240) & (!g254)) + ((g212) & (g219) & (!g226) & (!g233) & (g240) & (g254)) + ((g212) & (g219) & (!g226) & (g233) & (g240) & (g254)) + ((g212) & (g219) & (g226) & (!g233) & (!g240) & (!g254)) + ((g212) & (g219) & (g226) & (!g233) & (!g240) & (g254)) + ((g212) & (g219) & (g226) & (!g233) & (g240) & (!g254)) + ((g212) & (g219) & (g226) & (g233) & (!g240) & (g254)) + ((g212) & (g219) & (g226) & (g233) & (g240) & (!g254)));
	assign g1362 = (((!g212) & (!g219) & (!g226) & (!g233) & (!g240) & (g254)) + ((!g212) & (!g219) & (!g226) & (!g233) & (g240) & (!g254)) + ((!g212) & (!g219) & (!g226) & (!g233) & (g240) & (g254)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g240) & (!g254)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g240) & (g254)) + ((!g212) & (!g219) & (!g226) & (g233) & (g240) & (g254)) + ((!g212) & (!g219) & (g226) & (!g233) & (g240) & (!g254)) + ((!g212) & (!g219) & (g226) & (g233) & (!g240) & (!g254)) + ((!g212) & (!g219) & (g226) & (g233) & (!g240) & (g254)) + ((!g212) & (!g219) & (g226) & (g233) & (g240) & (g254)) + ((!g212) & (g219) & (!g226) & (!g233) & (g240) & (g254)) + ((!g212) & (g219) & (!g226) & (g233) & (!g240) & (!g254)) + ((!g212) & (g219) & (!g226) & (g233) & (g240) & (!g254)) + ((!g212) & (g219) & (g226) & (!g233) & (g240) & (!g254)) + ((!g212) & (g219) & (g226) & (!g233) & (g240) & (g254)) + ((!g212) & (g219) & (g226) & (g233) & (!g240) & (!g254)) + ((g212) & (!g219) & (!g226) & (!g233) & (!g240) & (!g254)) + ((g212) & (!g219) & (!g226) & (g233) & (!g240) & (!g254)) + ((g212) & (!g219) & (!g226) & (g233) & (!g240) & (g254)) + ((g212) & (!g219) & (g226) & (!g233) & (!g240) & (g254)) + ((g212) & (!g219) & (g226) & (!g233) & (g240) & (g254)) + ((g212) & (!g219) & (g226) & (g233) & (!g240) & (!g254)) + ((g212) & (!g219) & (g226) & (g233) & (!g240) & (g254)) + ((g212) & (g219) & (!g226) & (g233) & (!g240) & (!g254)) + ((g212) & (g219) & (!g226) & (g233) & (g240) & (g254)) + ((g212) & (g219) & (g226) & (!g233) & (!g240) & (!g254)) + ((g212) & (g219) & (g226) & (!g233) & (!g240) & (g254)) + ((g212) & (g219) & (g226) & (!g233) & (g240) & (g254)) + ((g212) & (g219) & (g226) & (g233) & (!g240) & (!g254)) + ((g212) & (g219) & (g226) & (g233) & (!g240) & (g254)) + ((g212) & (g219) & (g226) & (g233) & (g240) & (!g254)));
	assign g1363 = (((!g212) & (!g219) & (!g226) & (!g233) & (!g240) & (g254)) + ((!g212) & (!g219) & (!g226) & (g233) & (g240) & (!g254)) + ((!g212) & (!g219) & (g226) & (!g233) & (!g240) & (!g254)) + ((!g212) & (!g219) & (g226) & (!g233) & (g240) & (!g254)) + ((!g212) & (!g219) & (g226) & (g233) & (!g240) & (g254)) + ((!g212) & (!g219) & (g226) & (g233) & (g240) & (!g254)) + ((!g212) & (!g219) & (g226) & (g233) & (g240) & (g254)) + ((!g212) & (g219) & (!g226) & (!g233) & (!g240) & (!g254)) + ((!g212) & (g219) & (!g226) & (!g233) & (g240) & (!g254)) + ((!g212) & (g219) & (!g226) & (g233) & (!g240) & (!g254)) + ((!g212) & (g219) & (!g226) & (g233) & (g240) & (g254)) + ((!g212) & (g219) & (g226) & (!g233) & (g240) & (g254)) + ((!g212) & (g219) & (g226) & (g233) & (!g240) & (g254)) + ((!g212) & (g219) & (g226) & (g233) & (g240) & (!g254)) + ((g212) & (!g219) & (!g226) & (!g233) & (g240) & (g254)) + ((g212) & (!g219) & (!g226) & (g233) & (!g240) & (!g254)) + ((g212) & (!g219) & (!g226) & (g233) & (g240) & (!g254)) + ((g212) & (!g219) & (g226) & (!g233) & (!g240) & (!g254)) + ((g212) & (!g219) & (g226) & (!g233) & (!g240) & (g254)) + ((g212) & (!g219) & (g226) & (!g233) & (g240) & (!g254)) + ((g212) & (!g219) & (g226) & (!g233) & (g240) & (g254)) + ((g212) & (!g219) & (g226) & (g233) & (g240) & (!g254)) + ((g212) & (g219) & (!g226) & (!g233) & (!g240) & (g254)) + ((g212) & (g219) & (!g226) & (!g233) & (g240) & (g254)) + ((g212) & (g219) & (!g226) & (g233) & (!g240) & (g254)) + ((g212) & (g219) & (g226) & (!g233) & (!g240) & (!g254)) + ((g212) & (g219) & (g226) & (!g233) & (!g240) & (g254)) + ((g212) & (g219) & (g226) & (!g233) & (g240) & (g254)) + ((g212) & (g219) & (g226) & (g233) & (!g240) & (!g254)) + ((g212) & (g219) & (g226) & (g233) & (!g240) & (g254)) + ((g212) & (g219) & (g226) & (g233) & (g240) & (!g254)) + ((g212) & (g219) & (g226) & (g233) & (g240) & (g254)));
	assign g1364 = (((!g212) & (!g219) & (!g226) & (!g233) & (g240) & (!g254)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g240) & (!g254)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g240) & (g254)) + ((!g212) & (!g219) & (g226) & (!g233) & (g240) & (g254)) + ((!g212) & (!g219) & (g226) & (g233) & (!g240) & (g254)) + ((!g212) & (g219) & (!g226) & (!g233) & (!g240) & (!g254)) + ((!g212) & (g219) & (!g226) & (!g233) & (g240) & (!g254)) + ((!g212) & (g219) & (!g226) & (g233) & (!g240) & (g254)) + ((!g212) & (g219) & (g226) & (!g233) & (!g240) & (g254)) + ((!g212) & (g219) & (g226) & (!g233) & (g240) & (!g254)) + ((!g212) & (g219) & (g226) & (!g233) & (g240) & (g254)) + ((!g212) & (g219) & (g226) & (g233) & (g240) & (!g254)) + ((!g212) & (g219) & (g226) & (g233) & (g240) & (g254)) + ((g212) & (!g219) & (!g226) & (!g233) & (!g240) & (!g254)) + ((g212) & (!g219) & (!g226) & (g233) & (!g240) & (!g254)) + ((g212) & (!g219) & (!g226) & (g233) & (!g240) & (g254)) + ((g212) & (!g219) & (!g226) & (g233) & (g240) & (!g254)) + ((g212) & (!g219) & (g226) & (!g233) & (!g240) & (!g254)) + ((g212) & (!g219) & (g226) & (!g233) & (g240) & (g254)) + ((g212) & (!g219) & (g226) & (g233) & (g240) & (!g254)) + ((g212) & (g219) & (!g226) & (!g233) & (!g240) & (!g254)) + ((g212) & (g219) & (!g226) & (g233) & (!g240) & (!g254)) + ((g212) & (g219) & (!g226) & (g233) & (g240) & (!g254)) + ((g212) & (g219) & (!g226) & (g233) & (g240) & (g254)) + ((g212) & (g219) & (g226) & (g233) & (!g240) & (g254)) + ((g212) & (g219) & (g226) & (g233) & (g240) & (g254)));
	assign g1365 = (((!g1361) & (!g1362) & (!g1363) & (!g1364) & (!g247) & (!g261)) + ((!g1361) & (!g1362) & (!g1363) & (!g1364) & (g247) & (!g261)) + ((!g1361) & (!g1362) & (!g1363) & (g1364) & (!g247) & (!g261)) + ((!g1361) & (!g1362) & (!g1363) & (g1364) & (g247) & (!g261)) + ((!g1361) & (!g1362) & (!g1363) & (g1364) & (g247) & (g261)) + ((!g1361) & (!g1362) & (g1363) & (!g1364) & (!g247) & (!g261)) + ((!g1361) & (!g1362) & (g1363) & (!g1364) & (!g247) & (g261)) + ((!g1361) & (!g1362) & (g1363) & (!g1364) & (g247) & (!g261)) + ((!g1361) & (!g1362) & (g1363) & (g1364) & (!g247) & (!g261)) + ((!g1361) & (!g1362) & (g1363) & (g1364) & (!g247) & (g261)) + ((!g1361) & (!g1362) & (g1363) & (g1364) & (g247) & (!g261)) + ((!g1361) & (!g1362) & (g1363) & (g1364) & (g247) & (g261)) + ((!g1361) & (g1362) & (!g1363) & (!g1364) & (!g247) & (!g261)) + ((!g1361) & (g1362) & (!g1363) & (g1364) & (!g247) & (!g261)) + ((!g1361) & (g1362) & (!g1363) & (g1364) & (g247) & (g261)) + ((!g1361) & (g1362) & (g1363) & (!g1364) & (!g247) & (!g261)) + ((!g1361) & (g1362) & (g1363) & (!g1364) & (!g247) & (g261)) + ((!g1361) & (g1362) & (g1363) & (g1364) & (!g247) & (!g261)) + ((!g1361) & (g1362) & (g1363) & (g1364) & (!g247) & (g261)) + ((!g1361) & (g1362) & (g1363) & (g1364) & (g247) & (g261)) + ((g1361) & (!g1362) & (!g1363) & (!g1364) & (g247) & (!g261)) + ((g1361) & (!g1362) & (!g1363) & (g1364) & (g247) & (!g261)) + ((g1361) & (!g1362) & (!g1363) & (g1364) & (g247) & (g261)) + ((g1361) & (!g1362) & (g1363) & (!g1364) & (!g247) & (g261)) + ((g1361) & (!g1362) & (g1363) & (!g1364) & (g247) & (!g261)) + ((g1361) & (!g1362) & (g1363) & (g1364) & (!g247) & (g261)) + ((g1361) & (!g1362) & (g1363) & (g1364) & (g247) & (!g261)) + ((g1361) & (!g1362) & (g1363) & (g1364) & (g247) & (g261)) + ((g1361) & (g1362) & (!g1363) & (g1364) & (g247) & (g261)) + ((g1361) & (g1362) & (g1363) & (!g1364) & (!g247) & (g261)) + ((g1361) & (g1362) & (g1363) & (g1364) & (!g247) & (g261)) + ((g1361) & (g1362) & (g1363) & (g1364) & (g247) & (g261)));
	assign g1366 = (((!g539) & (!sk[79]) & (!g795) & (g1051) & (!g1365)) + ((!g539) & (!sk[79]) & (!g795) & (g1051) & (g1365)) + ((!g539) & (!sk[79]) & (g795) & (!g1051) & (!g1365)) + ((!g539) & (!sk[79]) & (g795) & (!g1051) & (g1365)) + ((!g539) & (!sk[79]) & (g795) & (g1051) & (!g1365)) + ((!g539) & (!sk[79]) & (g795) & (g1051) & (g1365)) + ((!g539) & (sk[79]) & (!g795) & (!g1051) & (g1365)) + ((!g539) & (sk[79]) & (!g795) & (g1051) & (!g1365)) + ((!g539) & (sk[79]) & (g795) & (!g1051) & (!g1365)) + ((!g539) & (sk[79]) & (g795) & (g1051) & (g1365)) + ((g539) & (!sk[79]) & (!g795) & (g1051) & (!g1365)) + ((g539) & (!sk[79]) & (!g795) & (g1051) & (g1365)) + ((g539) & (!sk[79]) & (g795) & (!g1051) & (!g1365)) + ((g539) & (!sk[79]) & (g795) & (!g1051) & (g1365)) + ((g539) & (!sk[79]) & (g795) & (g1051) & (!g1365)) + ((g539) & (!sk[79]) & (g795) & (g1051) & (g1365)) + ((g539) & (sk[79]) & (!g795) & (!g1051) & (!g1365)) + ((g539) & (sk[79]) & (!g795) & (g1051) & (g1365)) + ((g539) & (sk[79]) & (g795) & (!g1051) & (g1365)) + ((g539) & (sk[79]) & (g795) & (g1051) & (!g1365)));
	assign g1367 = (((!ld) & (!g283) & (!sk[80]) & (g1366) & (!keyx17x)) + ((!ld) & (!g283) & (!sk[80]) & (g1366) & (keyx17x)) + ((!ld) & (!g283) & (sk[80]) & (g1366) & (!keyx17x)) + ((!ld) & (!g283) & (sk[80]) & (g1366) & (keyx17x)) + ((!ld) & (g283) & (!sk[80]) & (!g1366) & (!keyx17x)) + ((!ld) & (g283) & (!sk[80]) & (!g1366) & (keyx17x)) + ((!ld) & (g283) & (!sk[80]) & (g1366) & (!keyx17x)) + ((!ld) & (g283) & (!sk[80]) & (g1366) & (keyx17x)) + ((!ld) & (g283) & (sk[80]) & (!g1366) & (!keyx17x)) + ((!ld) & (g283) & (sk[80]) & (!g1366) & (keyx17x)) + ((ld) & (!g283) & (!sk[80]) & (g1366) & (!keyx17x)) + ((ld) & (!g283) & (!sk[80]) & (g1366) & (keyx17x)) + ((ld) & (!g283) & (sk[80]) & (!g1366) & (keyx17x)) + ((ld) & (!g283) & (sk[80]) & (g1366) & (keyx17x)) + ((ld) & (g283) & (!sk[80]) & (!g1366) & (!keyx17x)) + ((ld) & (g283) & (!sk[80]) & (!g1366) & (keyx17x)) + ((ld) & (g283) & (!sk[80]) & (g1366) & (!keyx17x)) + ((ld) & (g283) & (!sk[80]) & (g1366) & (keyx17x)) + ((ld) & (g283) & (sk[80]) & (!g1366) & (keyx17x)) + ((ld) & (g283) & (sk[80]) & (g1366) & (keyx17x)));
	assign g1368 = (((!g254) & (!g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((!g254) & (!g219) & (!g226) & (!g233) & (g240) & (g247)) + ((!g254) & (!g219) & (!g226) & (g233) & (!g240) & (g247)) + ((!g254) & (!g219) & (!g226) & (g233) & (g240) & (!g247)) + ((!g254) & (!g219) & (!g226) & (g233) & (g240) & (g247)) + ((!g254) & (!g219) & (g226) & (!g233) & (!g240) & (g247)) + ((!g254) & (!g219) & (g226) & (g233) & (!g240) & (!g247)) + ((!g254) & (!g219) & (g226) & (g233) & (g240) & (!g247)) + ((!g254) & (g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((!g254) & (g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((!g254) & (g219) & (!g226) & (g233) & (!g240) & (g247)) + ((!g254) & (g219) & (g226) & (!g233) & (!g240) & (!g247)) + ((!g254) & (g219) & (g226) & (!g233) & (!g240) & (g247)) + ((!g254) & (g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g254) & (g219) & (g226) & (!g233) & (g240) & (g247)) + ((g254) & (!g219) & (!g226) & (g233) & (!g240) & (g247)) + ((g254) & (!g219) & (!g226) & (g233) & (g240) & (g247)) + ((g254) & (g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((g254) & (g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((g254) & (g219) & (!g226) & (g233) & (g240) & (!g247)) + ((g254) & (g219) & (g226) & (g233) & (!g240) & (!g247)) + ((g254) & (g219) & (g226) & (g233) & (!g240) & (g247)));
	assign g1369 = (((!g254) & (!g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((!g254) & (!g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((!g254) & (!g219) & (!g226) & (g233) & (g240) & (g247)) + ((!g254) & (!g219) & (g226) & (!g233) & (!g240) & (!g247)) + ((!g254) & (!g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g254) & (!g219) & (g226) & (g233) & (!g240) & (g247)) + ((!g254) & (g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((!g254) & (g219) & (!g226) & (!g233) & (g240) & (g247)) + ((!g254) & (g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((!g254) & (g219) & (!g226) & (g233) & (!g240) & (g247)) + ((!g254) & (g219) & (!g226) & (g233) & (g240) & (g247)) + ((!g254) & (g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g254) & (g219) & (g226) & (!g233) & (g240) & (g247)) + ((!g254) & (g219) & (g226) & (g233) & (g240) & (!g247)) + ((g254) & (!g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((g254) & (!g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((g254) & (!g219) & (!g226) & (!g233) & (g240) & (g247)) + ((g254) & (!g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((g254) & (!g219) & (!g226) & (g233) & (!g240) & (g247)) + ((g254) & (!g219) & (!g226) & (g233) & (g240) & (!g247)) + ((g254) & (!g219) & (g226) & (g233) & (!g240) & (!g247)) + ((g254) & (g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((g254) & (g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((g254) & (g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((g254) & (g219) & (!g226) & (g233) & (g240) & (!g247)) + ((g254) & (g219) & (!g226) & (g233) & (g240) & (g247)) + ((g254) & (g219) & (g226) & (!g233) & (!g240) & (!g247)) + ((g254) & (g219) & (g226) & (!g233) & (g240) & (!g247)) + ((g254) & (g219) & (g226) & (g233) & (!g240) & (g247)) + ((g254) & (g219) & (g226) & (g233) & (g240) & (g247)));
	assign g1370 = (((!g254) & (!g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((!g254) & (!g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((!g254) & (!g219) & (!g226) & (g233) & (!g240) & (g247)) + ((!g254) & (!g219) & (g226) & (!g233) & (!g240) & (g247)) + ((!g254) & (!g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g254) & (!g219) & (g226) & (g233) & (!g240) & (g247)) + ((!g254) & (g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((!g254) & (g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((!g254) & (g219) & (!g226) & (g233) & (g240) & (!g247)) + ((!g254) & (g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g254) & (g219) & (g226) & (g233) & (!g240) & (!g247)) + ((!g254) & (g219) & (g226) & (g233) & (g240) & (!g247)) + ((g254) & (!g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((g254) & (!g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((g254) & (!g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((g254) & (!g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((g254) & (!g219) & (!g226) & (g233) & (!g240) & (g247)) + ((g254) & (!g219) & (!g226) & (g233) & (g240) & (!g247)) + ((g254) & (!g219) & (!g226) & (g233) & (g240) & (g247)) + ((g254) & (!g219) & (g226) & (!g233) & (!g240) & (g247)) + ((g254) & (!g219) & (g226) & (!g233) & (g240) & (!g247)) + ((g254) & (!g219) & (g226) & (g233) & (!g240) & (!g247)) + ((g254) & (!g219) & (g226) & (g233) & (g240) & (g247)) + ((g254) & (g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((g254) & (g219) & (!g226) & (!g233) & (g240) & (g247)) + ((g254) & (g219) & (g226) & (!g233) & (g240) & (g247)) + ((g254) & (g219) & (g226) & (g233) & (!g240) & (!g247)) + ((g254) & (g219) & (g226) & (g233) & (!g240) & (g247)) + ((g254) & (g219) & (g226) & (g233) & (g240) & (g247)));
	assign g1371 = (((!g254) & (!g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((!g254) & (!g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((!g254) & (!g219) & (!g226) & (!g233) & (g240) & (g247)) + ((!g254) & (!g219) & (!g226) & (g233) & (!g240) & (g247)) + ((!g254) & (!g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g254) & (!g219) & (g226) & (g233) & (g240) & (g247)) + ((!g254) & (g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((!g254) & (g219) & (!g226) & (g233) & (!g240) & (g247)) + ((!g254) & (g219) & (!g226) & (g233) & (g240) & (g247)) + ((!g254) & (g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g254) & (g219) & (g226) & (!g233) & (g240) & (g247)) + ((!g254) & (g219) & (g226) & (g233) & (!g240) & (!g247)) + ((!g254) & (g219) & (g226) & (g233) & (!g240) & (g247)) + ((!g254) & (g219) & (g226) & (g233) & (g240) & (!g247)) + ((!g254) & (g219) & (g226) & (g233) & (g240) & (g247)) + ((g254) & (!g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((g254) & (!g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((g254) & (!g219) & (!g226) & (!g233) & (g240) & (g247)) + ((g254) & (!g219) & (!g226) & (g233) & (g240) & (g247)) + ((g254) & (!g219) & (g226) & (!g233) & (!g240) & (g247)) + ((g254) & (!g219) & (g226) & (!g233) & (g240) & (!g247)) + ((g254) & (!g219) & (g226) & (g233) & (g240) & (!g247)) + ((g254) & (g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((g254) & (g219) & (!g226) & (g233) & (!g240) & (g247)) + ((g254) & (g219) & (!g226) & (g233) & (g240) & (!g247)) + ((g254) & (g219) & (g226) & (!g233) & (g240) & (g247)) + ((g254) & (g219) & (g226) & (g233) & (!g240) & (!g247)));
	assign g1372 = (((!g1368) & (!g1369) & (!g1370) & (!g1371) & (!g212) & (g261)) + ((!g1368) & (!g1369) & (!g1370) & (!g1371) & (g212) & (!g261)) + ((!g1368) & (!g1369) & (!g1370) & (!g1371) & (g212) & (g261)) + ((!g1368) & (!g1369) & (!g1370) & (g1371) & (!g212) & (g261)) + ((!g1368) & (!g1369) & (!g1370) & (g1371) & (g212) & (!g261)) + ((!g1368) & (!g1369) & (g1370) & (!g1371) & (g212) & (!g261)) + ((!g1368) & (!g1369) & (g1370) & (!g1371) & (g212) & (g261)) + ((!g1368) & (!g1369) & (g1370) & (g1371) & (g212) & (!g261)) + ((!g1368) & (g1369) & (!g1370) & (!g1371) & (!g212) & (g261)) + ((!g1368) & (g1369) & (!g1370) & (!g1371) & (g212) & (g261)) + ((!g1368) & (g1369) & (!g1370) & (g1371) & (!g212) & (g261)) + ((!g1368) & (g1369) & (g1370) & (!g1371) & (g212) & (g261)) + ((g1368) & (!g1369) & (!g1370) & (!g1371) & (!g212) & (!g261)) + ((g1368) & (!g1369) & (!g1370) & (!g1371) & (!g212) & (g261)) + ((g1368) & (!g1369) & (!g1370) & (!g1371) & (g212) & (!g261)) + ((g1368) & (!g1369) & (!g1370) & (!g1371) & (g212) & (g261)) + ((g1368) & (!g1369) & (!g1370) & (g1371) & (!g212) & (!g261)) + ((g1368) & (!g1369) & (!g1370) & (g1371) & (!g212) & (g261)) + ((g1368) & (!g1369) & (!g1370) & (g1371) & (g212) & (!g261)) + ((g1368) & (!g1369) & (g1370) & (!g1371) & (!g212) & (!g261)) + ((g1368) & (!g1369) & (g1370) & (!g1371) & (g212) & (!g261)) + ((g1368) & (!g1369) & (g1370) & (!g1371) & (g212) & (g261)) + ((g1368) & (!g1369) & (g1370) & (g1371) & (!g212) & (!g261)) + ((g1368) & (!g1369) & (g1370) & (g1371) & (g212) & (!g261)) + ((g1368) & (g1369) & (!g1370) & (!g1371) & (!g212) & (!g261)) + ((g1368) & (g1369) & (!g1370) & (!g1371) & (!g212) & (g261)) + ((g1368) & (g1369) & (!g1370) & (!g1371) & (g212) & (g261)) + ((g1368) & (g1369) & (!g1370) & (g1371) & (!g212) & (!g261)) + ((g1368) & (g1369) & (!g1370) & (g1371) & (!g212) & (g261)) + ((g1368) & (g1369) & (g1370) & (!g1371) & (!g212) & (!g261)) + ((g1368) & (g1369) & (g1370) & (!g1371) & (g212) & (g261)) + ((g1368) & (g1369) & (g1370) & (g1371) & (!g212) & (!g261)));
	assign g1373 = (((!g546) & (!g802) & (!sk[86]) & (g1058) & (!g1372)) + ((!g546) & (!g802) & (!sk[86]) & (g1058) & (g1372)) + ((!g546) & (!g802) & (sk[86]) & (!g1058) & (g1372)) + ((!g546) & (!g802) & (sk[86]) & (g1058) & (!g1372)) + ((!g546) & (g802) & (!sk[86]) & (!g1058) & (!g1372)) + ((!g546) & (g802) & (!sk[86]) & (!g1058) & (g1372)) + ((!g546) & (g802) & (!sk[86]) & (g1058) & (!g1372)) + ((!g546) & (g802) & (!sk[86]) & (g1058) & (g1372)) + ((!g546) & (g802) & (sk[86]) & (!g1058) & (!g1372)) + ((!g546) & (g802) & (sk[86]) & (g1058) & (g1372)) + ((g546) & (!g802) & (!sk[86]) & (g1058) & (!g1372)) + ((g546) & (!g802) & (!sk[86]) & (g1058) & (g1372)) + ((g546) & (!g802) & (sk[86]) & (!g1058) & (!g1372)) + ((g546) & (!g802) & (sk[86]) & (g1058) & (g1372)) + ((g546) & (g802) & (!sk[86]) & (!g1058) & (!g1372)) + ((g546) & (g802) & (!sk[86]) & (!g1058) & (g1372)) + ((g546) & (g802) & (!sk[86]) & (g1058) & (!g1372)) + ((g546) & (g802) & (!sk[86]) & (g1058) & (g1372)) + ((g546) & (g802) & (sk[86]) & (!g1058) & (g1372)) + ((g546) & (g802) & (sk[86]) & (g1058) & (!g1372)));
	assign g1374 = (((!sk[87]) & (!ld) & (!g290) & (g1373) & (!keyx18x)) + ((!sk[87]) & (!ld) & (!g290) & (g1373) & (keyx18x)) + ((!sk[87]) & (!ld) & (g290) & (!g1373) & (!keyx18x)) + ((!sk[87]) & (!ld) & (g290) & (!g1373) & (keyx18x)) + ((!sk[87]) & (!ld) & (g290) & (g1373) & (!keyx18x)) + ((!sk[87]) & (!ld) & (g290) & (g1373) & (keyx18x)) + ((!sk[87]) & (ld) & (!g290) & (g1373) & (!keyx18x)) + ((!sk[87]) & (ld) & (!g290) & (g1373) & (keyx18x)) + ((!sk[87]) & (ld) & (g290) & (!g1373) & (!keyx18x)) + ((!sk[87]) & (ld) & (g290) & (!g1373) & (keyx18x)) + ((!sk[87]) & (ld) & (g290) & (g1373) & (!keyx18x)) + ((!sk[87]) & (ld) & (g290) & (g1373) & (keyx18x)) + ((sk[87]) & (!ld) & (!g290) & (g1373) & (!keyx18x)) + ((sk[87]) & (!ld) & (!g290) & (g1373) & (keyx18x)) + ((sk[87]) & (!ld) & (g290) & (!g1373) & (!keyx18x)) + ((sk[87]) & (!ld) & (g290) & (!g1373) & (keyx18x)) + ((sk[87]) & (ld) & (!g290) & (!g1373) & (keyx18x)) + ((sk[87]) & (ld) & (!g290) & (g1373) & (keyx18x)) + ((sk[87]) & (ld) & (g290) & (!g1373) & (keyx18x)) + ((sk[87]) & (ld) & (g290) & (g1373) & (keyx18x)));
	assign g1375 = (((!g212) & (!g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (g240) & (g247)) + ((!g212) & (!g219) & (g226) & (g233) & (!g240) & (!g247)) + ((!g212) & (!g219) & (g226) & (g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (g226) & (g233) & (g240) & (g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (g219) & (g226) & (!g233) & (!g240) & (!g247)) + ((!g212) & (g219) & (g226) & (g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((g212) & (!g219) & (g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (g226) & (!g233) & (!g240) & (g247)) + ((g212) & (!g219) & (g226) & (!g233) & (g240) & (!g247)) + ((g212) & (!g219) & (g226) & (g233) & (!g240) & (g247)) + ((g212) & (g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((g212) & (g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((g212) & (g219) & (!g226) & (g233) & (g240) & (!g247)) + ((g212) & (g219) & (g226) & (!g233) & (!g240) & (g247)) + ((g212) & (g219) & (g226) & (!g233) & (g240) & (g247)));
	assign g1376 = (((!g212) & (!g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (!g226) & (!g233) & (g240) & (g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (g226) & (g233) & (!g240) & (!g247)) + ((!g212) & (!g219) & (g226) & (g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (g226) & (g233) & (g240) & (g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (g240) & (g247)) + ((!g212) & (g219) & (!g226) & (g233) & (g240) & (g247)) + ((!g212) & (g219) & (g226) & (!g233) & (!g240) & (!g247)) + ((!g212) & (g219) & (g226) & (!g233) & (!g240) & (g247)) + ((!g212) & (g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (g219) & (g226) & (g233) & (!g240) & (g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((g212) & (!g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (!g226) & (g233) & (!g240) & (g247)) + ((g212) & (!g219) & (!g226) & (g233) & (g240) & (g247)) + ((g212) & (!g219) & (g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (g226) & (!g233) & (!g240) & (g247)) + ((g212) & (!g219) & (g226) & (!g233) & (g240) & (g247)) + ((g212) & (!g219) & (g226) & (g233) & (!g240) & (g247)) + ((g212) & (g219) & (!g226) & (g233) & (!g240) & (g247)) + ((g212) & (g219) & (!g226) & (g233) & (g240) & (!g247)) + ((g212) & (g219) & (g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (g219) & (g226) & (g233) & (!g240) & (!g247)));
	assign g1377 = (((!g212) & (!g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (!g226) & (!g233) & (g240) & (g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (g226) & (!g233) & (g240) & (g247)) + ((!g212) & (!g219) & (g226) & (g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (g226) & (g233) & (g240) & (g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (g240) & (g247)) + ((!g212) & (g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((!g212) & (g219) & (!g226) & (g233) & (!g240) & (g247)) + ((!g212) & (g219) & (g226) & (!g233) & (!g240) & (g247)) + ((!g212) & (g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (g219) & (g226) & (g233) & (g240) & (g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (g240) & (g247)) + ((g212) & (!g219) & (!g226) & (g233) & (g240) & (g247)) + ((g212) & (!g219) & (g226) & (g233) & (!g240) & (!g247)) + ((g212) & (g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((g212) & (g219) & (!g226) & (g233) & (g240) & (g247)) + ((g212) & (g219) & (g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (g219) & (g226) & (!g233) & (!g240) & (g247)) + ((g212) & (g219) & (g226) & (!g233) & (g240) & (g247)) + ((g212) & (g219) & (g226) & (g233) & (!g240) & (!g247)) + ((g212) & (g219) & (g226) & (g233) & (g240) & (g247)));
	assign g1378 = (((!g212) & (!g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (!g226) & (g233) & (g240) & (g247)) + ((!g212) & (!g219) & (g226) & (g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (g226) & (g233) & (g240) & (g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (!g240) & (!g247)) + ((!g212) & (g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (g219) & (!g226) & (g233) & (!g240) & (!g247)) + ((!g212) & (g219) & (!g226) & (g233) & (!g240) & (g247)) + ((!g212) & (g219) & (!g226) & (g233) & (g240) & (!g247)) + ((!g212) & (g219) & (g226) & (!g233) & (!g240) & (!g247)) + ((!g212) & (g219) & (g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (g219) & (g226) & (!g233) & (g240) & (g247)) + ((g212) & (!g219) & (!g226) & (!g233) & (g240) & (g247)) + ((g212) & (!g219) & (!g226) & (g233) & (g240) & (!g247)) + ((g212) & (!g219) & (g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (g226) & (!g233) & (g240) & (!g247)) + ((g212) & (!g219) & (g226) & (!g233) & (g240) & (g247)) + ((g212) & (!g219) & (g226) & (g233) & (!g240) & (g247)) + ((g212) & (!g219) & (g226) & (g233) & (g240) & (!g247)) + ((g212) & (!g219) & (g226) & (g233) & (g240) & (g247)) + ((g212) & (g219) & (!g226) & (!g233) & (!g240) & (g247)) + ((g212) & (g219) & (!g226) & (!g233) & (g240) & (!g247)) + ((g212) & (g219) & (g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (g219) & (g226) & (!g233) & (!g240) & (g247)) + ((g212) & (g219) & (g226) & (g233) & (g240) & (g247)));
	assign g1379 = (((!g1375) & (!g1376) & (!g1377) & (!g1378) & (!g261) & (g254)) + ((!g1375) & (!g1376) & (!g1377) & (!g1378) & (g261) & (!g254)) + ((!g1375) & (!g1376) & (!g1377) & (!g1378) & (g261) & (g254)) + ((!g1375) & (!g1376) & (!g1377) & (g1378) & (!g261) & (g254)) + ((!g1375) & (!g1376) & (!g1377) & (g1378) & (g261) & (!g254)) + ((!g1375) & (!g1376) & (g1377) & (!g1378) & (g261) & (!g254)) + ((!g1375) & (!g1376) & (g1377) & (!g1378) & (g261) & (g254)) + ((!g1375) & (!g1376) & (g1377) & (g1378) & (g261) & (!g254)) + ((!g1375) & (g1376) & (!g1377) & (!g1378) & (!g261) & (g254)) + ((!g1375) & (g1376) & (!g1377) & (!g1378) & (g261) & (g254)) + ((!g1375) & (g1376) & (!g1377) & (g1378) & (!g261) & (g254)) + ((!g1375) & (g1376) & (g1377) & (!g1378) & (g261) & (g254)) + ((g1375) & (!g1376) & (!g1377) & (!g1378) & (!g261) & (!g254)) + ((g1375) & (!g1376) & (!g1377) & (!g1378) & (!g261) & (g254)) + ((g1375) & (!g1376) & (!g1377) & (!g1378) & (g261) & (!g254)) + ((g1375) & (!g1376) & (!g1377) & (!g1378) & (g261) & (g254)) + ((g1375) & (!g1376) & (!g1377) & (g1378) & (!g261) & (!g254)) + ((g1375) & (!g1376) & (!g1377) & (g1378) & (!g261) & (g254)) + ((g1375) & (!g1376) & (!g1377) & (g1378) & (g261) & (!g254)) + ((g1375) & (!g1376) & (g1377) & (!g1378) & (!g261) & (!g254)) + ((g1375) & (!g1376) & (g1377) & (!g1378) & (g261) & (!g254)) + ((g1375) & (!g1376) & (g1377) & (!g1378) & (g261) & (g254)) + ((g1375) & (!g1376) & (g1377) & (g1378) & (!g261) & (!g254)) + ((g1375) & (!g1376) & (g1377) & (g1378) & (g261) & (!g254)) + ((g1375) & (g1376) & (!g1377) & (!g1378) & (!g261) & (!g254)) + ((g1375) & (g1376) & (!g1377) & (!g1378) & (!g261) & (g254)) + ((g1375) & (g1376) & (!g1377) & (!g1378) & (g261) & (g254)) + ((g1375) & (g1376) & (!g1377) & (g1378) & (!g261) & (!g254)) + ((g1375) & (g1376) & (!g1377) & (g1378) & (!g261) & (g254)) + ((g1375) & (g1376) & (g1377) & (!g1378) & (!g261) & (!g254)) + ((g1375) & (g1376) & (g1377) & (!g1378) & (g261) & (g254)) + ((g1375) & (g1376) & (g1377) & (g1378) & (!g261) & (!g254)));
	assign g1380 = (((!g553) & (!g809) & (!sk[93]) & (g1065) & (!g1379)) + ((!g553) & (!g809) & (!sk[93]) & (g1065) & (g1379)) + ((!g553) & (!g809) & (sk[93]) & (!g1065) & (g1379)) + ((!g553) & (!g809) & (sk[93]) & (g1065) & (!g1379)) + ((!g553) & (g809) & (!sk[93]) & (!g1065) & (!g1379)) + ((!g553) & (g809) & (!sk[93]) & (!g1065) & (g1379)) + ((!g553) & (g809) & (!sk[93]) & (g1065) & (!g1379)) + ((!g553) & (g809) & (!sk[93]) & (g1065) & (g1379)) + ((!g553) & (g809) & (sk[93]) & (!g1065) & (!g1379)) + ((!g553) & (g809) & (sk[93]) & (g1065) & (g1379)) + ((g553) & (!g809) & (!sk[93]) & (g1065) & (!g1379)) + ((g553) & (!g809) & (!sk[93]) & (g1065) & (g1379)) + ((g553) & (!g809) & (sk[93]) & (!g1065) & (!g1379)) + ((g553) & (!g809) & (sk[93]) & (g1065) & (g1379)) + ((g553) & (g809) & (!sk[93]) & (!g1065) & (!g1379)) + ((g553) & (g809) & (!sk[93]) & (!g1065) & (g1379)) + ((g553) & (g809) & (!sk[93]) & (g1065) & (!g1379)) + ((g553) & (g809) & (!sk[93]) & (g1065) & (g1379)) + ((g553) & (g809) & (sk[93]) & (!g1065) & (g1379)) + ((g553) & (g809) & (sk[93]) & (g1065) & (!g1379)));
	assign g1381 = (((!ld) & (!g297) & (!sk[94]) & (g1380) & (!keyx19x)) + ((!ld) & (!g297) & (!sk[94]) & (g1380) & (keyx19x)) + ((!ld) & (!g297) & (sk[94]) & (g1380) & (!keyx19x)) + ((!ld) & (!g297) & (sk[94]) & (g1380) & (keyx19x)) + ((!ld) & (g297) & (!sk[94]) & (!g1380) & (!keyx19x)) + ((!ld) & (g297) & (!sk[94]) & (!g1380) & (keyx19x)) + ((!ld) & (g297) & (!sk[94]) & (g1380) & (!keyx19x)) + ((!ld) & (g297) & (!sk[94]) & (g1380) & (keyx19x)) + ((!ld) & (g297) & (sk[94]) & (!g1380) & (!keyx19x)) + ((!ld) & (g297) & (sk[94]) & (!g1380) & (keyx19x)) + ((ld) & (!g297) & (!sk[94]) & (g1380) & (!keyx19x)) + ((ld) & (!g297) & (!sk[94]) & (g1380) & (keyx19x)) + ((ld) & (!g297) & (sk[94]) & (!g1380) & (keyx19x)) + ((ld) & (!g297) & (sk[94]) & (g1380) & (keyx19x)) + ((ld) & (g297) & (!sk[94]) & (!g1380) & (!keyx19x)) + ((ld) & (g297) & (!sk[94]) & (!g1380) & (keyx19x)) + ((ld) & (g297) & (!sk[94]) & (g1380) & (!keyx19x)) + ((ld) & (g297) & (!sk[94]) & (g1380) & (keyx19x)) + ((ld) & (g297) & (sk[94]) & (!g1380) & (keyx19x)) + ((ld) & (g297) & (sk[94]) & (g1380) & (keyx19x)));
	assign g1382 = (((!g212) & (!g219) & (!g254) & (!g261) & (!g240) & (g247)) + ((!g212) & (!g219) & (g254) & (!g261) & (!g240) & (g247)) + ((!g212) & (!g219) & (g254) & (!g261) & (g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (!g261) & (g240) & (g247)) + ((!g212) & (!g219) & (g254) & (g261) & (!g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (g261) & (g240) & (!g247)) + ((!g212) & (g219) & (!g254) & (!g261) & (!g240) & (!g247)) + ((!g212) & (g219) & (!g254) & (!g261) & (!g240) & (g247)) + ((!g212) & (g219) & (!g254) & (g261) & (!g240) & (!g247)) + ((!g212) & (g219) & (!g254) & (g261) & (!g240) & (g247)) + ((!g212) & (g219) & (!g254) & (g261) & (g240) & (g247)) + ((!g212) & (g219) & (g254) & (g261) & (!g240) & (g247)) + ((!g212) & (g219) & (g254) & (g261) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g261) & (!g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g261) & (!g240) & (g247)) + ((g212) & (!g219) & (!g254) & (g261) & (!g240) & (g247)) + ((g212) & (!g219) & (g254) & (!g261) & (g240) & (!g247)) + ((g212) & (!g219) & (g254) & (g261) & (!g240) & (!g247)) + ((g212) & (!g219) & (g254) & (g261) & (!g240) & (g247)) + ((g212) & (!g219) & (g254) & (g261) & (g240) & (!g247)) + ((g212) & (g219) & (!g254) & (!g261) & (!g240) & (!g247)) + ((g212) & (g219) & (!g254) & (!g261) & (g240) & (!g247)) + ((g212) & (g219) & (!g254) & (g261) & (g240) & (!g247)) + ((g212) & (g219) & (g254) & (!g261) & (!g240) & (!g247)) + ((g212) & (g219) & (g254) & (!g261) & (!g240) & (g247)) + ((g212) & (g219) & (g254) & (g261) & (!g240) & (g247)));
	assign g1383 = (((!g212) & (!g219) & (!g254) & (!g261) & (!g240) & (!g247)) + ((!g212) & (!g219) & (!g254) & (!g261) & (!g240) & (g247)) + ((!g212) & (!g219) & (!g254) & (!g261) & (g240) & (!g247)) + ((!g212) & (!g219) & (!g254) & (!g261) & (g240) & (g247)) + ((!g212) & (!g219) & (!g254) & (g261) & (!g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (!g261) & (!g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (!g261) & (g240) & (g247)) + ((!g212) & (!g219) & (g254) & (g261) & (!g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (g261) & (g240) & (g247)) + ((!g212) & (g219) & (!g254) & (!g261) & (!g240) & (g247)) + ((!g212) & (g219) & (!g254) & (g261) & (g240) & (!g247)) + ((!g212) & (g219) & (g254) & (!g261) & (!g240) & (!g247)) + ((!g212) & (g219) & (g254) & (!g261) & (!g240) & (g247)) + ((!g212) & (g219) & (g254) & (!g261) & (g240) & (!g247)) + ((!g212) & (g219) & (g254) & (!g261) & (g240) & (g247)) + ((!g212) & (g219) & (g254) & (g261) & (!g240) & (!g247)) + ((!g212) & (g219) & (g254) & (g261) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g261) & (!g240) & (g247)) + ((g212) & (!g219) & (!g254) & (!g261) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g261) & (g240) & (g247)) + ((g212) & (!g219) & (!g254) & (g261) & (!g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (g261) & (g240) & (g247)) + ((g212) & (!g219) & (g254) & (!g261) & (g240) & (!g247)) + ((g212) & (!g219) & (g254) & (!g261) & (g240) & (g247)) + ((g212) & (!g219) & (g254) & (g261) & (!g240) & (g247)) + ((g212) & (g219) & (!g254) & (!g261) & (g240) & (!g247)) + ((g212) & (g219) & (!g254) & (!g261) & (g240) & (g247)) + ((g212) & (g219) & (!g254) & (g261) & (!g240) & (!g247)) + ((g212) & (g219) & (!g254) & (g261) & (!g240) & (g247)) + ((g212) & (g219) & (g254) & (!g261) & (g240) & (!g247)) + ((g212) & (g219) & (g254) & (!g261) & (g240) & (g247)) + ((g212) & (g219) & (g254) & (g261) & (!g240) & (g247)));
	assign g1384 = (((!g212) & (!g219) & (!g254) & (!g261) & (!g240) & (!g247)) + ((!g212) & (!g219) & (!g254) & (!g261) & (!g240) & (g247)) + ((!g212) & (!g219) & (g254) & (!g261) & (!g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (!g261) & (g240) & (g247)) + ((!g212) & (!g219) & (g254) & (g261) & (!g240) & (g247)) + ((!g212) & (g219) & (!g254) & (g261) & (!g240) & (!g247)) + ((!g212) & (g219) & (!g254) & (g261) & (g240) & (!g247)) + ((!g212) & (g219) & (!g254) & (g261) & (g240) & (g247)) + ((!g212) & (g219) & (g254) & (!g261) & (!g240) & (!g247)) + ((!g212) & (g219) & (g254) & (!g261) & (g240) & (!g247)) + ((!g212) & (g219) & (g254) & (!g261) & (g240) & (g247)) + ((!g212) & (g219) & (g254) & (g261) & (!g240) & (!g247)) + ((!g212) & (g219) & (g254) & (g261) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g261) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g261) & (g240) & (g247)) + ((g212) & (!g219) & (!g254) & (g261) & (!g240) & (g247)) + ((g212) & (!g219) & (!g254) & (g261) & (g240) & (g247)) + ((g212) & (!g219) & (g254) & (!g261) & (!g240) & (!g247)) + ((g212) & (!g219) & (g254) & (!g261) & (!g240) & (g247)) + ((g212) & (!g219) & (g254) & (!g261) & (g240) & (g247)) + ((g212) & (!g219) & (g254) & (g261) & (!g240) & (!g247)) + ((g212) & (!g219) & (g254) & (g261) & (!g240) & (g247)) + ((g212) & (!g219) & (g254) & (g261) & (g240) & (!g247)) + ((g212) & (!g219) & (g254) & (g261) & (g240) & (g247)) + ((g212) & (g219) & (!g254) & (!g261) & (!g240) & (g247)) + ((g212) & (g219) & (!g254) & (g261) & (!g240) & (!g247)) + ((g212) & (g219) & (!g254) & (g261) & (g240) & (!g247)) + ((g212) & (g219) & (g254) & (!g261) & (!g240) & (!g247)) + ((g212) & (g219) & (g254) & (!g261) & (!g240) & (g247)) + ((g212) & (g219) & (g254) & (!g261) & (g240) & (!g247)) + ((g212) & (g219) & (g254) & (g261) & (!g240) & (!g247)) + ((g212) & (g219) & (g254) & (g261) & (g240) & (!g247)));
	assign g1385 = (((!g212) & (!g219) & (!g254) & (!g261) & (g240) & (g247)) + ((!g212) & (!g219) & (!g254) & (g261) & (!g240) & (!g247)) + ((!g212) & (!g219) & (!g254) & (g261) & (g240) & (g247)) + ((!g212) & (!g219) & (g254) & (!g261) & (!g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (!g261) & (g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (g261) & (!g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (g261) & (!g240) & (g247)) + ((!g212) & (!g219) & (g254) & (g261) & (g240) & (!g247)) + ((!g212) & (g219) & (!g254) & (!g261) & (!g240) & (!g247)) + ((!g212) & (g219) & (!g254) & (g261) & (!g240) & (g247)) + ((!g212) & (g219) & (!g254) & (g261) & (g240) & (!g247)) + ((!g212) & (g219) & (!g254) & (g261) & (g240) & (g247)) + ((!g212) & (g219) & (g254) & (!g261) & (!g240) & (!g247)) + ((!g212) & (g219) & (g254) & (g261) & (!g240) & (!g247)) + ((!g212) & (g219) & (g254) & (g261) & (!g240) & (g247)) + ((g212) & (!g219) & (!g254) & (!g261) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g261) & (g240) & (g247)) + ((g212) & (!g219) & (g254) & (!g261) & (!g240) & (!g247)) + ((g212) & (!g219) & (g254) & (!g261) & (g240) & (!g247)) + ((g212) & (!g219) & (g254) & (g261) & (g240) & (!g247)) + ((g212) & (g219) & (!g254) & (!g261) & (g240) & (!g247)) + ((g212) & (g219) & (!g254) & (g261) & (g240) & (g247)) + ((g212) & (g219) & (g254) & (!g261) & (!g240) & (!g247)) + ((g212) & (g219) & (g254) & (!g261) & (!g240) & (g247)) + ((g212) & (g219) & (g254) & (!g261) & (g240) & (!g247)) + ((g212) & (g219) & (g254) & (g261) & (!g240) & (!g247)));
	assign g1386 = (((!g1382) & (!g1383) & (!g1384) & (!g1385) & (g226) & (g233)) + ((!g1382) & (!g1383) & (g1384) & (!g1385) & (!g226) & (g233)) + ((!g1382) & (!g1383) & (g1384) & (!g1385) & (g226) & (g233)) + ((!g1382) & (!g1383) & (g1384) & (g1385) & (!g226) & (g233)) + ((!g1382) & (g1383) & (!g1384) & (!g1385) & (g226) & (!g233)) + ((!g1382) & (g1383) & (!g1384) & (!g1385) & (g226) & (g233)) + ((!g1382) & (g1383) & (!g1384) & (g1385) & (g226) & (!g233)) + ((!g1382) & (g1383) & (g1384) & (!g1385) & (!g226) & (g233)) + ((!g1382) & (g1383) & (g1384) & (!g1385) & (g226) & (!g233)) + ((!g1382) & (g1383) & (g1384) & (!g1385) & (g226) & (g233)) + ((!g1382) & (g1383) & (g1384) & (g1385) & (!g226) & (g233)) + ((!g1382) & (g1383) & (g1384) & (g1385) & (g226) & (!g233)) + ((g1382) & (!g1383) & (!g1384) & (!g1385) & (!g226) & (!g233)) + ((g1382) & (!g1383) & (!g1384) & (!g1385) & (g226) & (g233)) + ((g1382) & (!g1383) & (!g1384) & (g1385) & (!g226) & (!g233)) + ((g1382) & (!g1383) & (g1384) & (!g1385) & (!g226) & (!g233)) + ((g1382) & (!g1383) & (g1384) & (!g1385) & (!g226) & (g233)) + ((g1382) & (!g1383) & (g1384) & (!g1385) & (g226) & (g233)) + ((g1382) & (!g1383) & (g1384) & (g1385) & (!g226) & (!g233)) + ((g1382) & (!g1383) & (g1384) & (g1385) & (!g226) & (g233)) + ((g1382) & (g1383) & (!g1384) & (!g1385) & (!g226) & (!g233)) + ((g1382) & (g1383) & (!g1384) & (!g1385) & (g226) & (!g233)) + ((g1382) & (g1383) & (!g1384) & (!g1385) & (g226) & (g233)) + ((g1382) & (g1383) & (!g1384) & (g1385) & (!g226) & (!g233)) + ((g1382) & (g1383) & (!g1384) & (g1385) & (g226) & (!g233)) + ((g1382) & (g1383) & (g1384) & (!g1385) & (!g226) & (!g233)) + ((g1382) & (g1383) & (g1384) & (!g1385) & (!g226) & (g233)) + ((g1382) & (g1383) & (g1384) & (!g1385) & (g226) & (!g233)) + ((g1382) & (g1383) & (g1384) & (!g1385) & (g226) & (g233)) + ((g1382) & (g1383) & (g1384) & (g1385) & (!g226) & (!g233)) + ((g1382) & (g1383) & (g1384) & (g1385) & (!g226) & (g233)) + ((g1382) & (g1383) & (g1384) & (g1385) & (g226) & (!g233)));
	assign g1387 = (((!sk[100]) & (!g560) & (!g816) & (g1072) & (!g1386)) + ((!sk[100]) & (!g560) & (!g816) & (g1072) & (g1386)) + ((!sk[100]) & (!g560) & (g816) & (!g1072) & (!g1386)) + ((!sk[100]) & (!g560) & (g816) & (!g1072) & (g1386)) + ((!sk[100]) & (!g560) & (g816) & (g1072) & (!g1386)) + ((!sk[100]) & (!g560) & (g816) & (g1072) & (g1386)) + ((!sk[100]) & (g560) & (!g816) & (g1072) & (!g1386)) + ((!sk[100]) & (g560) & (!g816) & (g1072) & (g1386)) + ((!sk[100]) & (g560) & (g816) & (!g1072) & (!g1386)) + ((!sk[100]) & (g560) & (g816) & (!g1072) & (g1386)) + ((!sk[100]) & (g560) & (g816) & (g1072) & (!g1386)) + ((!sk[100]) & (g560) & (g816) & (g1072) & (g1386)) + ((sk[100]) & (!g560) & (!g816) & (!g1072) & (g1386)) + ((sk[100]) & (!g560) & (!g816) & (g1072) & (!g1386)) + ((sk[100]) & (!g560) & (g816) & (!g1072) & (!g1386)) + ((sk[100]) & (!g560) & (g816) & (g1072) & (g1386)) + ((sk[100]) & (g560) & (!g816) & (!g1072) & (!g1386)) + ((sk[100]) & (g560) & (!g816) & (g1072) & (g1386)) + ((sk[100]) & (g560) & (g816) & (!g1072) & (g1386)) + ((sk[100]) & (g560) & (g816) & (g1072) & (!g1386)));
	assign g1388 = (((!ld) & (!g304) & (g1387) & (!sk[101]) & (!keyx20x)) + ((!ld) & (!g304) & (g1387) & (!sk[101]) & (keyx20x)) + ((!ld) & (!g304) & (g1387) & (sk[101]) & (!keyx20x)) + ((!ld) & (!g304) & (g1387) & (sk[101]) & (keyx20x)) + ((!ld) & (g304) & (!g1387) & (!sk[101]) & (!keyx20x)) + ((!ld) & (g304) & (!g1387) & (!sk[101]) & (keyx20x)) + ((!ld) & (g304) & (!g1387) & (sk[101]) & (!keyx20x)) + ((!ld) & (g304) & (!g1387) & (sk[101]) & (keyx20x)) + ((!ld) & (g304) & (g1387) & (!sk[101]) & (!keyx20x)) + ((!ld) & (g304) & (g1387) & (!sk[101]) & (keyx20x)) + ((ld) & (!g304) & (!g1387) & (sk[101]) & (keyx20x)) + ((ld) & (!g304) & (g1387) & (!sk[101]) & (!keyx20x)) + ((ld) & (!g304) & (g1387) & (!sk[101]) & (keyx20x)) + ((ld) & (!g304) & (g1387) & (sk[101]) & (keyx20x)) + ((ld) & (g304) & (!g1387) & (!sk[101]) & (!keyx20x)) + ((ld) & (g304) & (!g1387) & (!sk[101]) & (keyx20x)) + ((ld) & (g304) & (!g1387) & (sk[101]) & (keyx20x)) + ((ld) & (g304) & (g1387) & (!sk[101]) & (!keyx20x)) + ((ld) & (g304) & (g1387) & (!sk[101]) & (keyx20x)) + ((ld) & (g304) & (g1387) & (sk[101]) & (keyx20x)));
	assign g1389 = (((!g212) & (!g219) & (!g254) & (!g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (!g254) & (!g233) & (g240) & (g247)) + ((!g212) & (!g219) & (!g254) & (g233) & (g240) & (g247)) + ((!g212) & (!g219) & (g254) & (!g233) & (!g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (!g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (g254) & (!g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (!g233) & (g240) & (g247)) + ((!g212) & (!g219) & (g254) & (g233) & (!g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (g233) & (!g240) & (g247)) + ((!g212) & (g219) & (!g254) & (!g233) & (!g240) & (g247)) + ((!g212) & (g219) & (!g254) & (!g233) & (g240) & (!g247)) + ((!g212) & (g219) & (!g254) & (g233) & (g240) & (g247)) + ((!g212) & (g219) & (g254) & (!g233) & (g240) & (!g247)) + ((!g212) & (g219) & (g254) & (!g233) & (g240) & (g247)) + ((!g212) & (g219) & (g254) & (g233) & (!g240) & (!g247)) + ((!g212) & (g219) & (g254) & (g233) & (!g240) & (g247)) + ((!g212) & (g219) & (g254) & (g233) & (g240) & (g247)) + ((g212) & (!g219) & (!g254) & (!g233) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g233) & (g240) & (g247)) + ((g212) & (!g219) & (!g254) & (g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (g233) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (g233) & (g240) & (g247)) + ((g212) & (!g219) & (g254) & (!g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (g254) & (!g233) & (g240) & (!g247)) + ((g212) & (!g219) & (g254) & (g233) & (g240) & (!g247)) + ((g212) & (g219) & (!g254) & (!g233) & (g240) & (g247)) + ((g212) & (g219) & (g254) & (!g233) & (!g240) & (!g247)) + ((g212) & (g219) & (g254) & (!g233) & (g240) & (g247)));
	assign g1390 = (((!g212) & (!g219) & (!g254) & (!g233) & (!g240) & (!g247)) + ((!g212) & (!g219) & (!g254) & (g233) & (!g240) & (!g247)) + ((!g212) & (!g219) & (!g254) & (g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (!g254) & (g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (!g233) & (g240) & (g247)) + ((!g212) & (!g219) & (g254) & (g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (g254) & (g233) & (g240) & (g247)) + ((!g212) & (g219) & (!g254) & (!g233) & (!g240) & (!g247)) + ((!g212) & (g219) & (!g254) & (!g233) & (g240) & (!g247)) + ((!g212) & (g219) & (g254) & (!g233) & (!g240) & (g247)) + ((!g212) & (g219) & (g254) & (!g233) & (g240) & (g247)) + ((!g212) & (g219) & (g254) & (g233) & (!g240) & (g247)) + ((!g212) & (g219) & (g254) & (g233) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g233) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g233) & (g240) & (g247)) + ((g212) & (!g219) & (!g254) & (g233) & (!g240) & (g247)) + ((g212) & (!g219) & (!g254) & (g233) & (g240) & (g247)) + ((g212) & (!g219) & (g254) & (g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (g254) & (g233) & (!g240) & (g247)) + ((g212) & (!g219) & (g254) & (g233) & (g240) & (g247)) + ((g212) & (g219) & (!g254) & (!g233) & (!g240) & (g247)) + ((g212) & (g219) & (!g254) & (!g233) & (g240) & (!g247)) + ((g212) & (g219) & (!g254) & (g233) & (g240) & (!g247)) + ((g212) & (g219) & (g254) & (!g233) & (!g240) & (g247)) + ((g212) & (g219) & (g254) & (!g233) & (g240) & (g247)) + ((g212) & (g219) & (g254) & (g233) & (!g240) & (!g247)) + ((g212) & (g219) & (g254) & (g233) & (g240) & (g247)));
	assign g1391 = (((!g212) & (!g219) & (!g254) & (!g233) & (g240) & (g247)) + ((!g212) & (!g219) & (!g254) & (g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (!g233) & (!g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (!g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (g254) & (!g233) & (g240) & (g247)) + ((!g212) & (!g219) & (g254) & (g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (g254) & (g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (g254) & (g233) & (g240) & (g247)) + ((!g212) & (g219) & (!g254) & (!g233) & (g240) & (!g247)) + ((!g212) & (g219) & (!g254) & (!g233) & (g240) & (g247)) + ((!g212) & (g219) & (g254) & (!g233) & (!g240) & (!g247)) + ((!g212) & (g219) & (g254) & (g233) & (!g240) & (g247)) + ((!g212) & (g219) & (g254) & (g233) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g233) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (!g233) & (g240) & (g247)) + ((g212) & (!g219) & (!g254) & (g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (g233) & (!g240) & (g247)) + ((g212) & (!g219) & (g254) & (!g233) & (!g240) & (g247)) + ((g212) & (!g219) & (g254) & (!g233) & (g240) & (g247)) + ((g212) & (!g219) & (g254) & (g233) & (g240) & (!g247)) + ((g212) & (g219) & (!g254) & (!g233) & (!g240) & (!g247)) + ((g212) & (g219) & (!g254) & (!g233) & (!g240) & (g247)) + ((g212) & (g219) & (!g254) & (!g233) & (g240) & (g247)) + ((g212) & (g219) & (!g254) & (g233) & (!g240) & (g247)) + ((g212) & (g219) & (!g254) & (g233) & (g240) & (!g247)) + ((g212) & (g219) & (g254) & (!g233) & (!g240) & (g247)) + ((g212) & (g219) & (g254) & (!g233) & (g240) & (!g247)) + ((g212) & (g219) & (g254) & (g233) & (!g240) & (!g247)) + ((g212) & (g219) & (g254) & (g233) & (g240) & (!g247)) + ((g212) & (g219) & (g254) & (g233) & (g240) & (g247)));
	assign g1392 = (((!g212) & (!g219) & (!g254) & (!g233) & (g240) & (!g247)) + ((!g212) & (!g219) & (!g254) & (g233) & (!g240) & (!g247)) + ((!g212) & (!g219) & (!g254) & (g233) & (g240) & (g247)) + ((!g212) & (!g219) & (g254) & (!g233) & (!g240) & (g247)) + ((!g212) & (!g219) & (g254) & (!g233) & (g240) & (g247)) + ((!g212) & (!g219) & (g254) & (g233) & (g240) & (g247)) + ((!g212) & (g219) & (!g254) & (!g233) & (!g240) & (g247)) + ((!g212) & (g219) & (!g254) & (g233) & (!g240) & (g247)) + ((!g212) & (g219) & (!g254) & (g233) & (g240) & (g247)) + ((!g212) & (g219) & (g254) & (!g233) & (!g240) & (!g247)) + ((!g212) & (g219) & (g254) & (!g233) & (g240) & (!g247)) + ((!g212) & (g219) & (g254) & (g233) & (!g240) & (g247)) + ((!g212) & (g219) & (g254) & (g233) & (g240) & (g247)) + ((g212) & (!g219) & (!g254) & (!g233) & (g240) & (!g247)) + ((g212) & (!g219) & (!g254) & (g233) & (g240) & (g247)) + ((g212) & (!g219) & (g254) & (!g233) & (!g240) & (!g247)) + ((g212) & (!g219) & (g254) & (!g233) & (g240) & (g247)) + ((g212) & (!g219) & (g254) & (g233) & (!g240) & (!g247)) + ((g212) & (g219) & (!g254) & (!g233) & (g240) & (g247)) + ((g212) & (g219) & (!g254) & (g233) & (!g240) & (!g247)) + ((g212) & (g219) & (!g254) & (g233) & (!g240) & (g247)) + ((g212) & (g219) & (g254) & (!g233) & (g240) & (g247)));
	assign g1393 = (((!g1389) & (!g1390) & (!g1391) & (!g1392) & (!g261) & (!g226)) + ((!g1389) & (!g1390) & (!g1391) & (!g1392) & (!g261) & (g226)) + ((!g1389) & (!g1390) & (!g1391) & (!g1392) & (g261) & (!g226)) + ((!g1389) & (!g1390) & (!g1391) & (g1392) & (!g261) & (!g226)) + ((!g1389) & (!g1390) & (!g1391) & (g1392) & (!g261) & (g226)) + ((!g1389) & (!g1390) & (!g1391) & (g1392) & (g261) & (!g226)) + ((!g1389) & (!g1390) & (!g1391) & (g1392) & (g261) & (g226)) + ((!g1389) & (!g1390) & (g1391) & (!g1392) & (!g261) & (!g226)) + ((!g1389) & (!g1390) & (g1391) & (!g1392) & (g261) & (!g226)) + ((!g1389) & (!g1390) & (g1391) & (g1392) & (!g261) & (!g226)) + ((!g1389) & (!g1390) & (g1391) & (g1392) & (g261) & (!g226)) + ((!g1389) & (!g1390) & (g1391) & (g1392) & (g261) & (g226)) + ((!g1389) & (g1390) & (!g1391) & (!g1392) & (!g261) & (!g226)) + ((!g1389) & (g1390) & (!g1391) & (!g1392) & (!g261) & (g226)) + ((!g1389) & (g1390) & (!g1391) & (g1392) & (!g261) & (!g226)) + ((!g1389) & (g1390) & (!g1391) & (g1392) & (!g261) & (g226)) + ((!g1389) & (g1390) & (!g1391) & (g1392) & (g261) & (g226)) + ((!g1389) & (g1390) & (g1391) & (!g1392) & (!g261) & (!g226)) + ((!g1389) & (g1390) & (g1391) & (g1392) & (!g261) & (!g226)) + ((!g1389) & (g1390) & (g1391) & (g1392) & (g261) & (g226)) + ((g1389) & (!g1390) & (!g1391) & (!g1392) & (!g261) & (g226)) + ((g1389) & (!g1390) & (!g1391) & (!g1392) & (g261) & (!g226)) + ((g1389) & (!g1390) & (!g1391) & (g1392) & (!g261) & (g226)) + ((g1389) & (!g1390) & (!g1391) & (g1392) & (g261) & (!g226)) + ((g1389) & (!g1390) & (!g1391) & (g1392) & (g261) & (g226)) + ((g1389) & (!g1390) & (g1391) & (!g1392) & (g261) & (!g226)) + ((g1389) & (!g1390) & (g1391) & (g1392) & (g261) & (!g226)) + ((g1389) & (!g1390) & (g1391) & (g1392) & (g261) & (g226)) + ((g1389) & (g1390) & (!g1391) & (!g1392) & (!g261) & (g226)) + ((g1389) & (g1390) & (!g1391) & (g1392) & (!g261) & (g226)) + ((g1389) & (g1390) & (!g1391) & (g1392) & (g261) & (g226)) + ((g1389) & (g1390) & (g1391) & (g1392) & (g261) & (g226)));
	assign g1394 = (((!g567) & (!sk[107]) & (!g823) & (g1079) & (!g1393)) + ((!g567) & (!sk[107]) & (!g823) & (g1079) & (g1393)) + ((!g567) & (!sk[107]) & (g823) & (!g1079) & (!g1393)) + ((!g567) & (!sk[107]) & (g823) & (!g1079) & (g1393)) + ((!g567) & (!sk[107]) & (g823) & (g1079) & (!g1393)) + ((!g567) & (!sk[107]) & (g823) & (g1079) & (g1393)) + ((!g567) & (sk[107]) & (!g823) & (!g1079) & (g1393)) + ((!g567) & (sk[107]) & (!g823) & (g1079) & (!g1393)) + ((!g567) & (sk[107]) & (g823) & (!g1079) & (!g1393)) + ((!g567) & (sk[107]) & (g823) & (g1079) & (g1393)) + ((g567) & (!sk[107]) & (!g823) & (g1079) & (!g1393)) + ((g567) & (!sk[107]) & (!g823) & (g1079) & (g1393)) + ((g567) & (!sk[107]) & (g823) & (!g1079) & (!g1393)) + ((g567) & (!sk[107]) & (g823) & (!g1079) & (g1393)) + ((g567) & (!sk[107]) & (g823) & (g1079) & (!g1393)) + ((g567) & (!sk[107]) & (g823) & (g1079) & (g1393)) + ((g567) & (sk[107]) & (!g823) & (!g1079) & (!g1393)) + ((g567) & (sk[107]) & (!g823) & (g1079) & (g1393)) + ((g567) & (sk[107]) & (g823) & (!g1079) & (g1393)) + ((g567) & (sk[107]) & (g823) & (g1079) & (!g1393)));
	assign g1395 = (((!sk[108]) & (!ld) & (!g311) & (g1394) & (!keyx21x)) + ((!sk[108]) & (!ld) & (!g311) & (g1394) & (keyx21x)) + ((!sk[108]) & (!ld) & (g311) & (!g1394) & (!keyx21x)) + ((!sk[108]) & (!ld) & (g311) & (!g1394) & (keyx21x)) + ((!sk[108]) & (!ld) & (g311) & (g1394) & (!keyx21x)) + ((!sk[108]) & (!ld) & (g311) & (g1394) & (keyx21x)) + ((!sk[108]) & (ld) & (!g311) & (g1394) & (!keyx21x)) + ((!sk[108]) & (ld) & (!g311) & (g1394) & (keyx21x)) + ((!sk[108]) & (ld) & (g311) & (!g1394) & (!keyx21x)) + ((!sk[108]) & (ld) & (g311) & (!g1394) & (keyx21x)) + ((!sk[108]) & (ld) & (g311) & (g1394) & (!keyx21x)) + ((!sk[108]) & (ld) & (g311) & (g1394) & (keyx21x)) + ((sk[108]) & (!ld) & (!g311) & (g1394) & (!keyx21x)) + ((sk[108]) & (!ld) & (!g311) & (g1394) & (keyx21x)) + ((sk[108]) & (!ld) & (g311) & (!g1394) & (!keyx21x)) + ((sk[108]) & (!ld) & (g311) & (!g1394) & (keyx21x)) + ((sk[108]) & (ld) & (!g311) & (!g1394) & (keyx21x)) + ((sk[108]) & (ld) & (!g311) & (g1394) & (keyx21x)) + ((sk[108]) & (ld) & (g311) & (!g1394) & (keyx21x)) + ((sk[108]) & (ld) & (g311) & (g1394) & (keyx21x)));
	assign g1396 = (((!g212) & (!g261) & (!g226) & (!g233) & (!g240) & (g247)) + ((!g212) & (!g261) & (!g226) & (!g233) & (g240) & (g247)) + ((!g212) & (!g261) & (!g226) & (g233) & (!g240) & (!g247)) + ((!g212) & (!g261) & (!g226) & (g233) & (!g240) & (g247)) + ((!g212) & (!g261) & (!g226) & (g233) & (g240) & (!g247)) + ((!g212) & (!g261) & (!g226) & (g233) & (g240) & (g247)) + ((!g212) & (!g261) & (g226) & (!g233) & (!g240) & (g247)) + ((!g212) & (!g261) & (g226) & (!g233) & (g240) & (g247)) + ((!g212) & (!g261) & (g226) & (g233) & (g240) & (!g247)) + ((!g212) & (g261) & (g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (g261) & (g226) & (!g233) & (g240) & (g247)) + ((!g212) & (g261) & (g226) & (g233) & (!g240) & (g247)) + ((g212) & (!g261) & (!g226) & (!g233) & (g240) & (!g247)) + ((g212) & (!g261) & (!g226) & (g233) & (!g240) & (!g247)) + ((g212) & (!g261) & (!g226) & (g233) & (!g240) & (g247)) + ((g212) & (!g261) & (!g226) & (g233) & (g240) & (g247)) + ((g212) & (!g261) & (g226) & (!g233) & (!g240) & (g247)) + ((g212) & (!g261) & (g226) & (!g233) & (g240) & (g247)) + ((g212) & (!g261) & (g226) & (g233) & (g240) & (!g247)) + ((g212) & (!g261) & (g226) & (g233) & (g240) & (g247)) + ((g212) & (g261) & (!g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (g261) & (!g226) & (!g233) & (!g240) & (g247)) + ((g212) & (g261) & (!g226) & (!g233) & (g240) & (!g247)) + ((g212) & (g261) & (!g226) & (g233) & (!g240) & (!g247)) + ((g212) & (g261) & (g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (g261) & (g226) & (!g233) & (!g240) & (g247)) + ((g212) & (g261) & (g226) & (!g233) & (g240) & (!g247)) + ((g212) & (g261) & (g226) & (g233) & (!g240) & (g247)));
	assign g1397 = (((!g212) & (!g261) & (!g226) & (!g233) & (!g240) & (!g247)) + ((!g212) & (!g261) & (!g226) & (g233) & (g240) & (g247)) + ((!g212) & (!g261) & (g226) & (!g233) & (!g240) & (!g247)) + ((!g212) & (!g261) & (g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (!g261) & (g226) & (!g233) & (g240) & (g247)) + ((!g212) & (!g261) & (g226) & (g233) & (!g240) & (!g247)) + ((!g212) & (!g261) & (g226) & (g233) & (g240) & (g247)) + ((!g212) & (g261) & (!g226) & (!g233) & (!g240) & (!g247)) + ((!g212) & (g261) & (!g226) & (!g233) & (g240) & (g247)) + ((!g212) & (g261) & (!g226) & (g233) & (!g240) & (g247)) + ((!g212) & (g261) & (g226) & (!g233) & (!g240) & (!g247)) + ((!g212) & (g261) & (g226) & (!g233) & (g240) & (g247)) + ((!g212) & (g261) & (g226) & (g233) & (g240) & (!g247)) + ((!g212) & (g261) & (g226) & (g233) & (g240) & (g247)) + ((g212) & (!g261) & (!g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (!g261) & (!g226) & (!g233) & (g240) & (g247)) + ((g212) & (!g261) & (!g226) & (g233) & (!g240) & (!g247)) + ((g212) & (!g261) & (!g226) & (g233) & (g240) & (g247)) + ((g212) & (!g261) & (g226) & (!g233) & (g240) & (g247)) + ((g212) & (!g261) & (g226) & (g233) & (!g240) & (g247)) + ((g212) & (g261) & (!g226) & (!g233) & (g240) & (!g247)) + ((g212) & (g261) & (!g226) & (!g233) & (g240) & (g247)) + ((g212) & (g261) & (!g226) & (g233) & (!g240) & (g247)) + ((g212) & (g261) & (!g226) & (g233) & (g240) & (!g247)) + ((g212) & (g261) & (!g226) & (g233) & (g240) & (g247)) + ((g212) & (g261) & (g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (g261) & (g226) & (!g233) & (g240) & (!g247)) + ((g212) & (g261) & (g226) & (g233) & (!g240) & (!g247)));
	assign g1398 = (((!g212) & (!g261) & (!g226) & (!g233) & (!g240) & (g247)) + ((!g212) & (!g261) & (!g226) & (!g233) & (g240) & (g247)) + ((!g212) & (!g261) & (!g226) & (g233) & (g240) & (!g247)) + ((!g212) & (!g261) & (!g226) & (g233) & (g240) & (g247)) + ((!g212) & (!g261) & (g226) & (!g233) & (g240) & (g247)) + ((!g212) & (!g261) & (g226) & (g233) & (!g240) & (!g247)) + ((!g212) & (!g261) & (g226) & (g233) & (!g240) & (g247)) + ((!g212) & (!g261) & (g226) & (g233) & (g240) & (g247)) + ((!g212) & (g261) & (!g226) & (!g233) & (!g240) & (!g247)) + ((!g212) & (g261) & (!g226) & (!g233) & (!g240) & (g247)) + ((!g212) & (g261) & (!g226) & (!g233) & (g240) & (g247)) + ((!g212) & (g261) & (!g226) & (g233) & (!g240) & (g247)) + ((!g212) & (g261) & (!g226) & (g233) & (g240) & (!g247)) + ((!g212) & (g261) & (g226) & (!g233) & (!g240) & (g247)) + ((!g212) & (g261) & (g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (g261) & (g226) & (g233) & (!g240) & (!g247)) + ((!g212) & (g261) & (g226) & (g233) & (g240) & (!g247)) + ((!g212) & (g261) & (g226) & (g233) & (g240) & (g247)) + ((g212) & (!g261) & (!g226) & (!g233) & (!g240) & (g247)) + ((g212) & (!g261) & (!g226) & (g233) & (!g240) & (!g247)) + ((g212) & (!g261) & (!g226) & (g233) & (g240) & (!g247)) + ((g212) & (!g261) & (g226) & (!g233) & (g240) & (g247)) + ((g212) & (!g261) & (g226) & (g233) & (!g240) & (g247)) + ((g212) & (g261) & (!g226) & (!g233) & (!g240) & (g247)) + ((g212) & (g261) & (!g226) & (g233) & (!g240) & (!g247)) + ((g212) & (g261) & (!g226) & (g233) & (g240) & (!g247)) + ((g212) & (g261) & (g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (g261) & (g226) & (!g233) & (g240) & (!g247)) + ((g212) & (g261) & (g226) & (!g233) & (g240) & (g247)) + ((g212) & (g261) & (g226) & (g233) & (g240) & (g247)));
	assign g1399 = (((!g212) & (!g261) & (!g226) & (!g233) & (g240) & (g247)) + ((!g212) & (!g261) & (!g226) & (g233) & (!g240) & (!g247)) + ((!g212) & (!g261) & (!g226) & (g233) & (g240) & (g247)) + ((!g212) & (!g261) & (g226) & (!g233) & (!g240) & (!g247)) + ((!g212) & (!g261) & (g226) & (g233) & (g240) & (!g247)) + ((!g212) & (!g261) & (g226) & (g233) & (g240) & (g247)) + ((!g212) & (g261) & (!g226) & (g233) & (!g240) & (!g247)) + ((!g212) & (g261) & (!g226) & (g233) & (g240) & (!g247)) + ((!g212) & (g261) & (g226) & (!g233) & (g240) & (!g247)) + ((!g212) & (g261) & (g226) & (!g233) & (g240) & (g247)) + ((g212) & (!g261) & (!g226) & (!g233) & (!g240) & (g247)) + ((g212) & (!g261) & (!g226) & (!g233) & (g240) & (!g247)) + ((g212) & (!g261) & (!g226) & (g233) & (!g240) & (g247)) + ((g212) & (!g261) & (g226) & (!g233) & (g240) & (!g247)) + ((g212) & (!g261) & (g226) & (!g233) & (g240) & (g247)) + ((g212) & (!g261) & (g226) & (g233) & (g240) & (!g247)) + ((g212) & (!g261) & (g226) & (g233) & (g240) & (g247)) + ((g212) & (g261) & (!g226) & (!g233) & (g240) & (!g247)) + ((g212) & (g261) & (!g226) & (g233) & (!g240) & (g247)) + ((g212) & (g261) & (g226) & (!g233) & (!g240) & (!g247)) + ((g212) & (g261) & (g226) & (!g233) & (g240) & (g247)) + ((g212) & (g261) & (g226) & (g233) & (!g240) & (g247)));
	assign g1400 = (((!g1396) & (!g1397) & (!g1398) & (!g1399) & (!g254) & (!g219)) + ((!g1396) & (!g1397) & (!g1398) & (!g1399) & (!g254) & (g219)) + ((!g1396) & (!g1397) & (!g1398) & (!g1399) & (g254) & (!g219)) + ((!g1396) & (!g1397) & (!g1398) & (g1399) & (!g254) & (!g219)) + ((!g1396) & (!g1397) & (!g1398) & (g1399) & (!g254) & (g219)) + ((!g1396) & (!g1397) & (!g1398) & (g1399) & (g254) & (!g219)) + ((!g1396) & (!g1397) & (!g1398) & (g1399) & (g254) & (g219)) + ((!g1396) & (!g1397) & (g1398) & (!g1399) & (!g254) & (!g219)) + ((!g1396) & (!g1397) & (g1398) & (!g1399) & (g254) & (!g219)) + ((!g1396) & (!g1397) & (g1398) & (g1399) & (!g254) & (!g219)) + ((!g1396) & (!g1397) & (g1398) & (g1399) & (g254) & (!g219)) + ((!g1396) & (!g1397) & (g1398) & (g1399) & (g254) & (g219)) + ((!g1396) & (g1397) & (!g1398) & (!g1399) & (!g254) & (!g219)) + ((!g1396) & (g1397) & (!g1398) & (!g1399) & (!g254) & (g219)) + ((!g1396) & (g1397) & (!g1398) & (g1399) & (!g254) & (!g219)) + ((!g1396) & (g1397) & (!g1398) & (g1399) & (!g254) & (g219)) + ((!g1396) & (g1397) & (!g1398) & (g1399) & (g254) & (g219)) + ((!g1396) & (g1397) & (g1398) & (!g1399) & (!g254) & (!g219)) + ((!g1396) & (g1397) & (g1398) & (g1399) & (!g254) & (!g219)) + ((!g1396) & (g1397) & (g1398) & (g1399) & (g254) & (g219)) + ((g1396) & (!g1397) & (!g1398) & (!g1399) & (!g254) & (g219)) + ((g1396) & (!g1397) & (!g1398) & (!g1399) & (g254) & (!g219)) + ((g1396) & (!g1397) & (!g1398) & (g1399) & (!g254) & (g219)) + ((g1396) & (!g1397) & (!g1398) & (g1399) & (g254) & (!g219)) + ((g1396) & (!g1397) & (!g1398) & (g1399) & (g254) & (g219)) + ((g1396) & (!g1397) & (g1398) & (!g1399) & (g254) & (!g219)) + ((g1396) & (!g1397) & (g1398) & (g1399) & (g254) & (!g219)) + ((g1396) & (!g1397) & (g1398) & (g1399) & (g254) & (g219)) + ((g1396) & (g1397) & (!g1398) & (!g1399) & (!g254) & (g219)) + ((g1396) & (g1397) & (!g1398) & (g1399) & (!g254) & (g219)) + ((g1396) & (g1397) & (!g1398) & (g1399) & (g254) & (g219)) + ((g1396) & (g1397) & (g1398) & (g1399) & (g254) & (g219)));
	assign g1401 = (((!g574) & (!sk[114]) & (!g830) & (g1086) & (!g1400)) + ((!g574) & (!sk[114]) & (!g830) & (g1086) & (g1400)) + ((!g574) & (!sk[114]) & (g830) & (!g1086) & (!g1400)) + ((!g574) & (!sk[114]) & (g830) & (!g1086) & (g1400)) + ((!g574) & (!sk[114]) & (g830) & (g1086) & (!g1400)) + ((!g574) & (!sk[114]) & (g830) & (g1086) & (g1400)) + ((!g574) & (sk[114]) & (!g830) & (!g1086) & (g1400)) + ((!g574) & (sk[114]) & (!g830) & (g1086) & (!g1400)) + ((!g574) & (sk[114]) & (g830) & (!g1086) & (!g1400)) + ((!g574) & (sk[114]) & (g830) & (g1086) & (g1400)) + ((g574) & (!sk[114]) & (!g830) & (g1086) & (!g1400)) + ((g574) & (!sk[114]) & (!g830) & (g1086) & (g1400)) + ((g574) & (!sk[114]) & (g830) & (!g1086) & (!g1400)) + ((g574) & (!sk[114]) & (g830) & (!g1086) & (g1400)) + ((g574) & (!sk[114]) & (g830) & (g1086) & (!g1400)) + ((g574) & (!sk[114]) & (g830) & (g1086) & (g1400)) + ((g574) & (sk[114]) & (!g830) & (!g1086) & (!g1400)) + ((g574) & (sk[114]) & (!g830) & (g1086) & (g1400)) + ((g574) & (sk[114]) & (g830) & (!g1086) & (g1400)) + ((g574) & (sk[114]) & (g830) & (g1086) & (!g1400)));
	assign g1402 = (((!ld) & (!sk[115]) & (!g318) & (g1401) & (!keyx22x)) + ((!ld) & (!sk[115]) & (!g318) & (g1401) & (keyx22x)) + ((!ld) & (!sk[115]) & (g318) & (!g1401) & (!keyx22x)) + ((!ld) & (!sk[115]) & (g318) & (!g1401) & (keyx22x)) + ((!ld) & (!sk[115]) & (g318) & (g1401) & (!keyx22x)) + ((!ld) & (!sk[115]) & (g318) & (g1401) & (keyx22x)) + ((!ld) & (sk[115]) & (!g318) & (g1401) & (!keyx22x)) + ((!ld) & (sk[115]) & (!g318) & (g1401) & (keyx22x)) + ((!ld) & (sk[115]) & (g318) & (!g1401) & (!keyx22x)) + ((!ld) & (sk[115]) & (g318) & (!g1401) & (keyx22x)) + ((ld) & (!sk[115]) & (!g318) & (g1401) & (!keyx22x)) + ((ld) & (!sk[115]) & (!g318) & (g1401) & (keyx22x)) + ((ld) & (!sk[115]) & (g318) & (!g1401) & (!keyx22x)) + ((ld) & (!sk[115]) & (g318) & (!g1401) & (keyx22x)) + ((ld) & (!sk[115]) & (g318) & (g1401) & (!keyx22x)) + ((ld) & (!sk[115]) & (g318) & (g1401) & (keyx22x)) + ((ld) & (sk[115]) & (!g318) & (!g1401) & (keyx22x)) + ((ld) & (sk[115]) & (!g318) & (g1401) & (keyx22x)) + ((ld) & (sk[115]) & (g318) & (!g1401) & (keyx22x)) + ((ld) & (sk[115]) & (g318) & (g1401) & (keyx22x)));
	assign g1403 = (((!g254) & (!g219) & (!g226) & (!g233) & (!g240) & (g261)) + ((!g254) & (!g219) & (!g226) & (!g233) & (g240) & (!g261)) + ((!g254) & (!g219) & (!g226) & (g233) & (!g240) & (g261)) + ((!g254) & (!g219) & (!g226) & (g233) & (g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (!g233) & (!g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (!g233) & (g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (g233) & (!g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (g233) & (g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (g233) & (g240) & (g261)) + ((!g254) & (g219) & (!g226) & (!g233) & (g240) & (!g261)) + ((!g254) & (g219) & (!g226) & (g233) & (g240) & (!g261)) + ((!g254) & (g219) & (!g226) & (g233) & (g240) & (g261)) + ((!g254) & (g219) & (g226) & (!g233) & (g240) & (g261)) + ((!g254) & (g219) & (g226) & (g233) & (!g240) & (!g261)) + ((g254) & (!g219) & (!g226) & (!g233) & (!g240) & (g261)) + ((g254) & (!g219) & (!g226) & (g233) & (!g240) & (g261)) + ((g254) & (!g219) & (g226) & (g233) & (g240) & (g261)) + ((g254) & (g219) & (!g226) & (!g233) & (g240) & (g261)) + ((g254) & (g219) & (!g226) & (g233) & (!g240) & (!g261)) + ((g254) & (g219) & (!g226) & (g233) & (g240) & (!g261)) + ((g254) & (g219) & (g226) & (!g233) & (!g240) & (g261)) + ((g254) & (g219) & (g226) & (!g233) & (g240) & (!g261)) + ((g254) & (g219) & (g226) & (!g233) & (g240) & (g261)) + ((g254) & (g219) & (g226) & (g233) & (!g240) & (g261)));
	assign g1404 = (((!g254) & (!g219) & (!g226) & (!g233) & (!g240) & (!g261)) + ((!g254) & (!g219) & (!g226) & (!g233) & (!g240) & (g261)) + ((!g254) & (!g219) & (!g226) & (g233) & (!g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (!g233) & (!g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (!g233) & (g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (!g233) & (g240) & (g261)) + ((!g254) & (!g219) & (g226) & (g233) & (!g240) & (g261)) + ((!g254) & (!g219) & (g226) & (g233) & (g240) & (g261)) + ((!g254) & (g219) & (!g226) & (!g233) & (!g240) & (!g261)) + ((!g254) & (g219) & (!g226) & (!g233) & (g240) & (!g261)) + ((!g254) & (g219) & (!g226) & (g233) & (!g240) & (!g261)) + ((!g254) & (g219) & (!g226) & (g233) & (!g240) & (g261)) + ((!g254) & (g219) & (!g226) & (g233) & (g240) & (g261)) + ((!g254) & (g219) & (g226) & (!g233) & (!g240) & (g261)) + ((!g254) & (g219) & (g226) & (g233) & (!g240) & (!g261)) + ((!g254) & (g219) & (g226) & (g233) & (!g240) & (g261)) + ((g254) & (!g219) & (!g226) & (!g233) & (!g240) & (g261)) + ((g254) & (!g219) & (!g226) & (!g233) & (g240) & (g261)) + ((g254) & (!g219) & (!g226) & (g233) & (!g240) & (!g261)) + ((g254) & (!g219) & (!g226) & (g233) & (g240) & (g261)) + ((g254) & (!g219) & (g226) & (!g233) & (!g240) & (!g261)) + ((g254) & (!g219) & (g226) & (!g233) & (g240) & (g261)) + ((g254) & (!g219) & (g226) & (g233) & (g240) & (!g261)) + ((g254) & (g219) & (!g226) & (!g233) & (!g240) & (!g261)) + ((g254) & (g219) & (!g226) & (!g233) & (!g240) & (g261)) + ((g254) & (g219) & (!g226) & (!g233) & (g240) & (g261)) + ((g254) & (g219) & (!g226) & (g233) & (!g240) & (g261)) + ((g254) & (g219) & (!g226) & (g233) & (g240) & (!g261)) + ((g254) & (g219) & (g226) & (!g233) & (g240) & (!g261)) + ((g254) & (g219) & (g226) & (!g233) & (g240) & (g261)));
	assign g1405 = (((!g254) & (!g219) & (!g226) & (!g233) & (g240) & (!g261)) + ((!g254) & (!g219) & (!g226) & (g233) & (!g240) & (!g261)) + ((!g254) & (!g219) & (!g226) & (g233) & (g240) & (!g261)) + ((!g254) & (!g219) & (!g226) & (g233) & (g240) & (g261)) + ((!g254) & (!g219) & (g226) & (!g233) & (!g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (!g233) & (!g240) & (g261)) + ((!g254) & (!g219) & (g226) & (!g233) & (g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (g233) & (!g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (g233) & (g240) & (g261)) + ((!g254) & (g219) & (!g226) & (!g233) & (!g240) & (g261)) + ((!g254) & (g219) & (!g226) & (!g233) & (g240) & (!g261)) + ((!g254) & (g219) & (!g226) & (!g233) & (g240) & (g261)) + ((!g254) & (g219) & (g226) & (!g233) & (!g240) & (g261)) + ((!g254) & (g219) & (g226) & (!g233) & (g240) & (!g261)) + ((!g254) & (g219) & (g226) & (!g233) & (g240) & (g261)) + ((!g254) & (g219) & (g226) & (g233) & (!g240) & (!g261)) + ((g254) & (!g219) & (!g226) & (!g233) & (g240) & (!g261)) + ((g254) & (!g219) & (!g226) & (g233) & (!g240) & (!g261)) + ((g254) & (!g219) & (!g226) & (g233) & (g240) & (g261)) + ((g254) & (!g219) & (g226) & (!g233) & (!g240) & (!g261)) + ((g254) & (!g219) & (g226) & (!g233) & (!g240) & (g261)) + ((g254) & (!g219) & (g226) & (g233) & (!g240) & (!g261)) + ((g254) & (!g219) & (g226) & (g233) & (g240) & (!g261)) + ((g254) & (g219) & (!g226) & (!g233) & (g240) & (!g261)) + ((g254) & (g219) & (!g226) & (g233) & (!g240) & (!g261)) + ((g254) & (g219) & (!g226) & (g233) & (g240) & (g261)) + ((g254) & (g219) & (g226) & (!g233) & (!g240) & (!g261)) + ((g254) & (g219) & (g226) & (!g233) & (g240) & (!g261)) + ((g254) & (g219) & (g226) & (!g233) & (g240) & (g261)) + ((g254) & (g219) & (g226) & (g233) & (!g240) & (g261)));
	assign g1406 = (((!g254) & (!g219) & (!g226) & (!g233) & (!g240) & (g261)) + ((!g254) & (!g219) & (!g226) & (g233) & (g240) & (!g261)) + ((!g254) & (!g219) & (!g226) & (g233) & (g240) & (g261)) + ((!g254) & (!g219) & (g226) & (!g233) & (!g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (!g233) & (!g240) & (g261)) + ((!g254) & (!g219) & (g226) & (g233) & (g240) & (!g261)) + ((!g254) & (!g219) & (g226) & (g233) & (g240) & (g261)) + ((!g254) & (g219) & (!g226) & (!g233) & (!g240) & (!g261)) + ((!g254) & (g219) & (!g226) & (!g233) & (!g240) & (g261)) + ((!g254) & (g219) & (!g226) & (!g233) & (g240) & (g261)) + ((!g254) & (g219) & (!g226) & (g233) & (!g240) & (g261)) + ((!g254) & (g219) & (g226) & (!g233) & (!g240) & (g261)) + ((!g254) & (g219) & (g226) & (g233) & (!g240) & (!g261)) + ((!g254) & (g219) & (g226) & (g233) & (!g240) & (g261)) + ((!g254) & (g219) & (g226) & (g233) & (g240) & (!g261)) + ((!g254) & (g219) & (g226) & (g233) & (g240) & (g261)) + ((g254) & (!g219) & (!g226) & (g233) & (!g240) & (g261)) + ((g254) & (!g219) & (g226) & (!g233) & (!g240) & (!g261)) + ((g254) & (!g219) & (g226) & (g233) & (!g240) & (!g261)) + ((g254) & (!g219) & (g226) & (g233) & (!g240) & (g261)) + ((g254) & (!g219) & (g226) & (g233) & (g240) & (g261)) + ((g254) & (g219) & (!g226) & (!g233) & (!g240) & (g261)) + ((g254) & (g219) & (!g226) & (!g233) & (g240) & (g261)) + ((g254) & (g219) & (!g226) & (g233) & (!g240) & (!g261)) + ((g254) & (g219) & (!g226) & (g233) & (g240) & (!g261)) + ((g254) & (g219) & (!g226) & (g233) & (g240) & (g261)) + ((g254) & (g219) & (g226) & (!g233) & (g240) & (g261)) + ((g254) & (g219) & (g226) & (g233) & (g240) & (g261)));
	assign g1407 = (((!g1403) & (!g1404) & (!g1405) & (!g1406) & (!g212) & (g247)) + ((!g1403) & (!g1404) & (!g1405) & (!g1406) & (g212) & (!g247)) + ((!g1403) & (!g1404) & (!g1405) & (!g1406) & (g212) & (g247)) + ((!g1403) & (!g1404) & (!g1405) & (g1406) & (!g212) & (g247)) + ((!g1403) & (!g1404) & (!g1405) & (g1406) & (g212) & (!g247)) + ((!g1403) & (!g1404) & (g1405) & (!g1406) & (g212) & (!g247)) + ((!g1403) & (!g1404) & (g1405) & (!g1406) & (g212) & (g247)) + ((!g1403) & (!g1404) & (g1405) & (g1406) & (g212) & (!g247)) + ((!g1403) & (g1404) & (!g1405) & (!g1406) & (!g212) & (g247)) + ((!g1403) & (g1404) & (!g1405) & (!g1406) & (g212) & (g247)) + ((!g1403) & (g1404) & (!g1405) & (g1406) & (!g212) & (g247)) + ((!g1403) & (g1404) & (g1405) & (!g1406) & (g212) & (g247)) + ((g1403) & (!g1404) & (!g1405) & (!g1406) & (!g212) & (!g247)) + ((g1403) & (!g1404) & (!g1405) & (!g1406) & (!g212) & (g247)) + ((g1403) & (!g1404) & (!g1405) & (!g1406) & (g212) & (!g247)) + ((g1403) & (!g1404) & (!g1405) & (!g1406) & (g212) & (g247)) + ((g1403) & (!g1404) & (!g1405) & (g1406) & (!g212) & (!g247)) + ((g1403) & (!g1404) & (!g1405) & (g1406) & (!g212) & (g247)) + ((g1403) & (!g1404) & (!g1405) & (g1406) & (g212) & (!g247)) + ((g1403) & (!g1404) & (g1405) & (!g1406) & (!g212) & (!g247)) + ((g1403) & (!g1404) & (g1405) & (!g1406) & (g212) & (!g247)) + ((g1403) & (!g1404) & (g1405) & (!g1406) & (g212) & (g247)) + ((g1403) & (!g1404) & (g1405) & (g1406) & (!g212) & (!g247)) + ((g1403) & (!g1404) & (g1405) & (g1406) & (g212) & (!g247)) + ((g1403) & (g1404) & (!g1405) & (!g1406) & (!g212) & (!g247)) + ((g1403) & (g1404) & (!g1405) & (!g1406) & (!g212) & (g247)) + ((g1403) & (g1404) & (!g1405) & (!g1406) & (g212) & (g247)) + ((g1403) & (g1404) & (!g1405) & (g1406) & (!g212) & (!g247)) + ((g1403) & (g1404) & (!g1405) & (g1406) & (!g212) & (g247)) + ((g1403) & (g1404) & (g1405) & (!g1406) & (!g212) & (!g247)) + ((g1403) & (g1404) & (g1405) & (!g1406) & (g212) & (g247)) + ((g1403) & (g1404) & (g1405) & (g1406) & (!g212) & (!g247)));
	assign g1408 = (((!g581) & (!g837) & (!g1093) & (sk[121]) & (g1407)) + ((!g581) & (!g837) & (g1093) & (!sk[121]) & (!g1407)) + ((!g581) & (!g837) & (g1093) & (!sk[121]) & (g1407)) + ((!g581) & (!g837) & (g1093) & (sk[121]) & (!g1407)) + ((!g581) & (g837) & (!g1093) & (!sk[121]) & (!g1407)) + ((!g581) & (g837) & (!g1093) & (!sk[121]) & (g1407)) + ((!g581) & (g837) & (!g1093) & (sk[121]) & (!g1407)) + ((!g581) & (g837) & (g1093) & (!sk[121]) & (!g1407)) + ((!g581) & (g837) & (g1093) & (!sk[121]) & (g1407)) + ((!g581) & (g837) & (g1093) & (sk[121]) & (g1407)) + ((g581) & (!g837) & (!g1093) & (sk[121]) & (!g1407)) + ((g581) & (!g837) & (g1093) & (!sk[121]) & (!g1407)) + ((g581) & (!g837) & (g1093) & (!sk[121]) & (g1407)) + ((g581) & (!g837) & (g1093) & (sk[121]) & (g1407)) + ((g581) & (g837) & (!g1093) & (!sk[121]) & (!g1407)) + ((g581) & (g837) & (!g1093) & (!sk[121]) & (g1407)) + ((g581) & (g837) & (!g1093) & (sk[121]) & (g1407)) + ((g581) & (g837) & (g1093) & (!sk[121]) & (!g1407)) + ((g581) & (g837) & (g1093) & (!sk[121]) & (g1407)) + ((g581) & (g837) & (g1093) & (sk[121]) & (!g1407)));
	assign g1409 = (((!ld) & (!g325) & (!sk[122]) & (g1408) & (!keyx23x)) + ((!ld) & (!g325) & (!sk[122]) & (g1408) & (keyx23x)) + ((!ld) & (!g325) & (sk[122]) & (g1408) & (!keyx23x)) + ((!ld) & (!g325) & (sk[122]) & (g1408) & (keyx23x)) + ((!ld) & (g325) & (!sk[122]) & (!g1408) & (!keyx23x)) + ((!ld) & (g325) & (!sk[122]) & (!g1408) & (keyx23x)) + ((!ld) & (g325) & (!sk[122]) & (g1408) & (!keyx23x)) + ((!ld) & (g325) & (!sk[122]) & (g1408) & (keyx23x)) + ((!ld) & (g325) & (sk[122]) & (!g1408) & (!keyx23x)) + ((!ld) & (g325) & (sk[122]) & (!g1408) & (keyx23x)) + ((ld) & (!g325) & (!sk[122]) & (g1408) & (!keyx23x)) + ((ld) & (!g325) & (!sk[122]) & (g1408) & (keyx23x)) + ((ld) & (!g325) & (sk[122]) & (!g1408) & (keyx23x)) + ((ld) & (!g325) & (sk[122]) & (g1408) & (keyx23x)) + ((ld) & (g325) & (!sk[122]) & (!g1408) & (!keyx23x)) + ((ld) & (g325) & (!sk[122]) & (!g1408) & (keyx23x)) + ((ld) & (g325) & (!sk[122]) & (g1408) & (!keyx23x)) + ((ld) & (g325) & (!sk[122]) & (g1408) & (keyx23x)) + ((ld) & (g325) & (sk[122]) & (!g1408) & (keyx23x)) + ((ld) & (g325) & (sk[122]) & (g1408) & (keyx23x)));
	assign g2106 = (((!ld) & (!text_inx24x) & (sk[123]) & (g1410)) + ((!ld) & (text_inx24x) & (!sk[123]) & (!g1410)) + ((!ld) & (text_inx24x) & (!sk[123]) & (g1410)) + ((!ld) & (text_inx24x) & (sk[123]) & (g1410)) + ((ld) & (!text_inx24x) & (!sk[123]) & (g1410)) + ((ld) & (text_inx24x) & (!sk[123]) & (!g1410)) + ((ld) & (text_inx24x) & (!sk[123]) & (g1410)) + ((ld) & (text_inx24x) & (sk[123]) & (!g1410)) + ((ld) & (text_inx24x) & (sk[123]) & (g1410)));
	assign g1411 = (((!sk[124]) & (!g147) & (g211)) + ((!sk[124]) & (g147) & (g211)) + ((sk[124]) & (!g147) & (g211)) + ((sk[124]) & (g147) & (!g211)));
	assign g1412 = (((!sk[125]) & (!g275) & (g324)) + ((!sk[125]) & (g275) & (g324)) + ((sk[125]) & (!g275) & (g324)) + ((sk[125]) & (g275) & (!g324)));
	assign g1413 = (((!g340) & (!g388) & (!g1163) & (!g1410) & (!g1411) & (g1412)) + ((!g340) & (!g388) & (!g1163) & (!g1410) & (g1411) & (!g1412)) + ((!g340) & (!g388) & (!g1163) & (g1410) & (!g1411) & (g1412)) + ((!g340) & (!g388) & (!g1163) & (g1410) & (g1411) & (!g1412)) + ((!g340) & (!g388) & (g1163) & (g1410) & (!g1411) & (!g1412)) + ((!g340) & (!g388) & (g1163) & (g1410) & (!g1411) & (g1412)) + ((!g340) & (!g388) & (g1163) & (g1410) & (g1411) & (!g1412)) + ((!g340) & (!g388) & (g1163) & (g1410) & (g1411) & (g1412)) + ((!g340) & (g388) & (!g1163) & (!g1410) & (!g1411) & (!g1412)) + ((!g340) & (g388) & (!g1163) & (!g1410) & (g1411) & (g1412)) + ((!g340) & (g388) & (!g1163) & (g1410) & (!g1411) & (!g1412)) + ((!g340) & (g388) & (!g1163) & (g1410) & (g1411) & (g1412)) + ((!g340) & (g388) & (g1163) & (g1410) & (!g1411) & (!g1412)) + ((!g340) & (g388) & (g1163) & (g1410) & (!g1411) & (g1412)) + ((!g340) & (g388) & (g1163) & (g1410) & (g1411) & (!g1412)) + ((!g340) & (g388) & (g1163) & (g1410) & (g1411) & (g1412)) + ((g340) & (!g388) & (!g1163) & (!g1410) & (!g1411) & (!g1412)) + ((g340) & (!g388) & (!g1163) & (!g1410) & (g1411) & (g1412)) + ((g340) & (!g388) & (!g1163) & (g1410) & (!g1411) & (!g1412)) + ((g340) & (!g388) & (!g1163) & (g1410) & (g1411) & (g1412)) + ((g340) & (!g388) & (g1163) & (!g1410) & (!g1411) & (!g1412)) + ((g340) & (!g388) & (g1163) & (!g1410) & (!g1411) & (g1412)) + ((g340) & (!g388) & (g1163) & (!g1410) & (g1411) & (!g1412)) + ((g340) & (!g388) & (g1163) & (!g1410) & (g1411) & (g1412)) + ((g340) & (g388) & (!g1163) & (!g1410) & (!g1411) & (g1412)) + ((g340) & (g388) & (!g1163) & (!g1410) & (g1411) & (!g1412)) + ((g340) & (g388) & (!g1163) & (g1410) & (!g1411) & (g1412)) + ((g340) & (g388) & (!g1163) & (g1410) & (g1411) & (!g1412)) + ((g340) & (g388) & (g1163) & (!g1410) & (!g1411) & (!g1412)) + ((g340) & (g388) & (g1163) & (!g1410) & (!g1411) & (g1412)) + ((g340) & (g388) & (g1163) & (!g1410) & (g1411) & (!g1412)) + ((g340) & (g388) & (g1163) & (!g1410) & (g1411) & (g1412)));
	assign g2107 = (((!sk[127]) & (!ld) & (text_inx25x) & (!g1414)) + ((!sk[127]) & (!ld) & (text_inx25x) & (g1414)) + ((!sk[127]) & (ld) & (!text_inx25x) & (g1414)) + ((!sk[127]) & (ld) & (text_inx25x) & (!g1414)) + ((!sk[127]) & (ld) & (text_inx25x) & (g1414)) + ((sk[127]) & (!ld) & (!text_inx25x) & (g1414)) + ((sk[127]) & (!ld) & (text_inx25x) & (g1414)) + ((sk[127]) & (ld) & (text_inx25x) & (!g1414)) + ((sk[127]) & (ld) & (text_inx25x) & (g1414)));
	assign g1415 = (((!g154) & (!g218) & (!sk[0]) & (g275) & (!g324)) + ((!g154) & (!g218) & (!sk[0]) & (g275) & (g324)) + ((!g154) & (!g218) & (sk[0]) & (!g275) & (g324)) + ((!g154) & (!g218) & (sk[0]) & (g275) & (!g324)) + ((!g154) & (g218) & (!sk[0]) & (!g275) & (!g324)) + ((!g154) & (g218) & (!sk[0]) & (!g275) & (g324)) + ((!g154) & (g218) & (!sk[0]) & (g275) & (!g324)) + ((!g154) & (g218) & (!sk[0]) & (g275) & (g324)) + ((!g154) & (g218) & (sk[0]) & (!g275) & (!g324)) + ((!g154) & (g218) & (sk[0]) & (g275) & (g324)) + ((g154) & (!g218) & (!sk[0]) & (g275) & (!g324)) + ((g154) & (!g218) & (!sk[0]) & (g275) & (g324)) + ((g154) & (!g218) & (sk[0]) & (!g275) & (!g324)) + ((g154) & (!g218) & (sk[0]) & (g275) & (g324)) + ((g154) & (g218) & (!sk[0]) & (!g275) & (!g324)) + ((g154) & (g218) & (!sk[0]) & (!g275) & (g324)) + ((g154) & (g218) & (!sk[0]) & (g275) & (!g324)) + ((g154) & (g218) & (!sk[0]) & (g275) & (g324)) + ((g154) & (g218) & (sk[0]) & (!g275) & (g324)) + ((g154) & (g218) & (sk[0]) & (g275) & (!g324)));
	assign g2108 = (((!ld) & (!text_inx26x) & (sk[1]) & (g1416)) + ((!ld) & (text_inx26x) & (!sk[1]) & (!g1416)) + ((!ld) & (text_inx26x) & (!sk[1]) & (g1416)) + ((!ld) & (text_inx26x) & (sk[1]) & (g1416)) + ((ld) & (!text_inx26x) & (!sk[1]) & (g1416)) + ((ld) & (text_inx26x) & (!sk[1]) & (!g1416)) + ((ld) & (text_inx26x) & (!sk[1]) & (g1416)) + ((ld) & (text_inx26x) & (sk[1]) & (!g1416)) + ((ld) & (text_inx26x) & (sk[1]) & (g1416)));
	assign g1417 = (((!g161) & (!g225) & (sk[2]) & (g282)) + ((!g161) & (g225) & (!sk[2]) & (!g282)) + ((!g161) & (g225) & (!sk[2]) & (g282)) + ((!g161) & (g225) & (sk[2]) & (!g282)) + ((g161) & (!g225) & (!sk[2]) & (g282)) + ((g161) & (!g225) & (sk[2]) & (!g282)) + ((g161) & (g225) & (!sk[2]) & (!g282)) + ((g161) & (g225) & (!sk[2]) & (g282)) + ((g161) & (g225) & (sk[2]) & (g282)));
	assign g1418 = (((!g289) & (!g346) & (!g354) & (!g1163) & (!g1416) & (g1417)) + ((!g289) & (!g346) & (!g354) & (!g1163) & (g1416) & (g1417)) + ((!g289) & (!g346) & (!g354) & (g1163) & (g1416) & (!g1417)) + ((!g289) & (!g346) & (!g354) & (g1163) & (g1416) & (g1417)) + ((!g289) & (!g346) & (g354) & (!g1163) & (!g1416) & (!g1417)) + ((!g289) & (!g346) & (g354) & (!g1163) & (g1416) & (!g1417)) + ((!g289) & (!g346) & (g354) & (g1163) & (!g1416) & (!g1417)) + ((!g289) & (!g346) & (g354) & (g1163) & (!g1416) & (g1417)) + ((!g289) & (g346) & (!g354) & (!g1163) & (!g1416) & (!g1417)) + ((!g289) & (g346) & (!g354) & (!g1163) & (g1416) & (!g1417)) + ((!g289) & (g346) & (!g354) & (g1163) & (g1416) & (!g1417)) + ((!g289) & (g346) & (!g354) & (g1163) & (g1416) & (g1417)) + ((!g289) & (g346) & (g354) & (!g1163) & (!g1416) & (g1417)) + ((!g289) & (g346) & (g354) & (!g1163) & (g1416) & (g1417)) + ((!g289) & (g346) & (g354) & (g1163) & (!g1416) & (!g1417)) + ((!g289) & (g346) & (g354) & (g1163) & (!g1416) & (g1417)) + ((g289) & (!g346) & (!g354) & (!g1163) & (!g1416) & (!g1417)) + ((g289) & (!g346) & (!g354) & (!g1163) & (g1416) & (!g1417)) + ((g289) & (!g346) & (!g354) & (g1163) & (g1416) & (!g1417)) + ((g289) & (!g346) & (!g354) & (g1163) & (g1416) & (g1417)) + ((g289) & (!g346) & (g354) & (!g1163) & (!g1416) & (g1417)) + ((g289) & (!g346) & (g354) & (!g1163) & (g1416) & (g1417)) + ((g289) & (!g346) & (g354) & (g1163) & (!g1416) & (!g1417)) + ((g289) & (!g346) & (g354) & (g1163) & (!g1416) & (g1417)) + ((g289) & (g346) & (!g354) & (!g1163) & (!g1416) & (g1417)) + ((g289) & (g346) & (!g354) & (!g1163) & (g1416) & (g1417)) + ((g289) & (g346) & (!g354) & (g1163) & (g1416) & (!g1417)) + ((g289) & (g346) & (!g354) & (g1163) & (g1416) & (g1417)) + ((g289) & (g346) & (g354) & (!g1163) & (!g1416) & (!g1417)) + ((g289) & (g346) & (g354) & (!g1163) & (g1416) & (!g1417)) + ((g289) & (g346) & (g354) & (g1163) & (!g1416) & (!g1417)) + ((g289) & (g346) & (g354) & (g1163) & (!g1416) & (g1417)));
	assign g2109 = (((!sk[4]) & (!ld) & (text_inx27x) & (!g1419)) + ((!sk[4]) & (!ld) & (text_inx27x) & (g1419)) + ((!sk[4]) & (ld) & (!text_inx27x) & (g1419)) + ((!sk[4]) & (ld) & (text_inx27x) & (!g1419)) + ((!sk[4]) & (ld) & (text_inx27x) & (g1419)) + ((sk[4]) & (!ld) & (!text_inx27x) & (g1419)) + ((sk[4]) & (!ld) & (text_inx27x) & (g1419)) + ((sk[4]) & (ld) & (text_inx27x) & (!g1419)) + ((sk[4]) & (ld) & (text_inx27x) & (g1419)));
	assign g1420 = (((!g168) & (!g232) & (!g289) & (!g353) & (!g361) & (g388)) + ((!g168) & (!g232) & (!g289) & (!g353) & (g361) & (!g388)) + ((!g168) & (!g232) & (!g289) & (g353) & (!g361) & (!g388)) + ((!g168) & (!g232) & (!g289) & (g353) & (g361) & (g388)) + ((!g168) & (!g232) & (g289) & (!g353) & (!g361) & (!g388)) + ((!g168) & (!g232) & (g289) & (!g353) & (g361) & (g388)) + ((!g168) & (!g232) & (g289) & (g353) & (!g361) & (g388)) + ((!g168) & (!g232) & (g289) & (g353) & (g361) & (!g388)) + ((!g168) & (g232) & (!g289) & (!g353) & (!g361) & (!g388)) + ((!g168) & (g232) & (!g289) & (!g353) & (g361) & (g388)) + ((!g168) & (g232) & (!g289) & (g353) & (!g361) & (g388)) + ((!g168) & (g232) & (!g289) & (g353) & (g361) & (!g388)) + ((!g168) & (g232) & (g289) & (!g353) & (!g361) & (g388)) + ((!g168) & (g232) & (g289) & (!g353) & (g361) & (!g388)) + ((!g168) & (g232) & (g289) & (g353) & (!g361) & (!g388)) + ((!g168) & (g232) & (g289) & (g353) & (g361) & (g388)) + ((g168) & (!g232) & (!g289) & (!g353) & (!g361) & (!g388)) + ((g168) & (!g232) & (!g289) & (!g353) & (g361) & (g388)) + ((g168) & (!g232) & (!g289) & (g353) & (!g361) & (g388)) + ((g168) & (!g232) & (!g289) & (g353) & (g361) & (!g388)) + ((g168) & (!g232) & (g289) & (!g353) & (!g361) & (g388)) + ((g168) & (!g232) & (g289) & (!g353) & (g361) & (!g388)) + ((g168) & (!g232) & (g289) & (g353) & (!g361) & (!g388)) + ((g168) & (!g232) & (g289) & (g353) & (g361) & (g388)) + ((g168) & (g232) & (!g289) & (!g353) & (!g361) & (g388)) + ((g168) & (g232) & (!g289) & (!g353) & (g361) & (!g388)) + ((g168) & (g232) & (!g289) & (g353) & (!g361) & (!g388)) + ((g168) & (g232) & (!g289) & (g353) & (g361) & (g388)) + ((g168) & (g232) & (g289) & (!g353) & (!g361) & (!g388)) + ((g168) & (g232) & (g289) & (!g353) & (g361) & (g388)) + ((g168) & (g232) & (g289) & (g353) & (!g361) & (g388)) + ((g168) & (g232) & (g289) & (g353) & (g361) & (!g388)));
	assign g1421 = (((!g296) & (!g324) & (!g361) & (!g1163) & (!g1419) & (g1420)) + ((!g296) & (!g324) & (!g361) & (!g1163) & (g1419) & (g1420)) + ((!g296) & (!g324) & (!g361) & (g1163) & (g1419) & (!g1420)) + ((!g296) & (!g324) & (!g361) & (g1163) & (g1419) & (g1420)) + ((!g296) & (!g324) & (g361) & (!g1163) & (!g1419) & (g1420)) + ((!g296) & (!g324) & (g361) & (!g1163) & (g1419) & (g1420)) + ((!g296) & (!g324) & (g361) & (g1163) & (!g1419) & (!g1420)) + ((!g296) & (!g324) & (g361) & (g1163) & (!g1419) & (g1420)) + ((!g296) & (g324) & (!g361) & (!g1163) & (!g1419) & (!g1420)) + ((!g296) & (g324) & (!g361) & (!g1163) & (g1419) & (!g1420)) + ((!g296) & (g324) & (!g361) & (g1163) & (g1419) & (!g1420)) + ((!g296) & (g324) & (!g361) & (g1163) & (g1419) & (g1420)) + ((!g296) & (g324) & (g361) & (!g1163) & (!g1419) & (!g1420)) + ((!g296) & (g324) & (g361) & (!g1163) & (g1419) & (!g1420)) + ((!g296) & (g324) & (g361) & (g1163) & (!g1419) & (!g1420)) + ((!g296) & (g324) & (g361) & (g1163) & (!g1419) & (g1420)) + ((g296) & (!g324) & (!g361) & (!g1163) & (!g1419) & (!g1420)) + ((g296) & (!g324) & (!g361) & (!g1163) & (g1419) & (!g1420)) + ((g296) & (!g324) & (!g361) & (g1163) & (g1419) & (!g1420)) + ((g296) & (!g324) & (!g361) & (g1163) & (g1419) & (g1420)) + ((g296) & (!g324) & (g361) & (!g1163) & (!g1419) & (!g1420)) + ((g296) & (!g324) & (g361) & (!g1163) & (g1419) & (!g1420)) + ((g296) & (!g324) & (g361) & (g1163) & (!g1419) & (!g1420)) + ((g296) & (!g324) & (g361) & (g1163) & (!g1419) & (g1420)) + ((g296) & (g324) & (!g361) & (!g1163) & (!g1419) & (g1420)) + ((g296) & (g324) & (!g361) & (!g1163) & (g1419) & (g1420)) + ((g296) & (g324) & (!g361) & (g1163) & (g1419) & (!g1420)) + ((g296) & (g324) & (!g361) & (g1163) & (g1419) & (g1420)) + ((g296) & (g324) & (g361) & (!g1163) & (!g1419) & (g1420)) + ((g296) & (g324) & (g361) & (!g1163) & (g1419) & (g1420)) + ((g296) & (g324) & (g361) & (g1163) & (!g1419) & (!g1420)) + ((g296) & (g324) & (g361) & (g1163) & (!g1419) & (g1420)));
	assign g2110 = (((!sk[7]) & (!ld) & (text_inx30x) & (!g1422)) + ((!sk[7]) & (!ld) & (text_inx30x) & (g1422)) + ((!sk[7]) & (ld) & (!text_inx30x) & (g1422)) + ((!sk[7]) & (ld) & (text_inx30x) & (!g1422)) + ((!sk[7]) & (ld) & (text_inx30x) & (g1422)) + ((sk[7]) & (!ld) & (!text_inx30x) & (g1422)) + ((sk[7]) & (!ld) & (text_inx30x) & (g1422)) + ((sk[7]) & (ld) & (text_inx30x) & (!g1422)) + ((sk[7]) & (ld) & (text_inx30x) & (g1422)));
	assign g1423 = (((!g189) & (!g253) & (sk[8]) & (g310)) + ((!g189) & (g253) & (!sk[8]) & (!g310)) + ((!g189) & (g253) & (!sk[8]) & (g310)) + ((!g189) & (g253) & (sk[8]) & (!g310)) + ((g189) & (!g253) & (!sk[8]) & (g310)) + ((g189) & (!g253) & (sk[8]) & (!g310)) + ((g189) & (g253) & (!sk[8]) & (!g310)) + ((g189) & (g253) & (!sk[8]) & (g310)) + ((g189) & (g253) & (sk[8]) & (g310)));
	assign g1424 = (((!g317) & (!g374) & (!g382) & (!g1163) & (!g1422) & (g1423)) + ((!g317) & (!g374) & (!g382) & (!g1163) & (g1422) & (g1423)) + ((!g317) & (!g374) & (!g382) & (g1163) & (g1422) & (!g1423)) + ((!g317) & (!g374) & (!g382) & (g1163) & (g1422) & (g1423)) + ((!g317) & (!g374) & (g382) & (!g1163) & (!g1422) & (!g1423)) + ((!g317) & (!g374) & (g382) & (!g1163) & (g1422) & (!g1423)) + ((!g317) & (!g374) & (g382) & (g1163) & (!g1422) & (!g1423)) + ((!g317) & (!g374) & (g382) & (g1163) & (!g1422) & (g1423)) + ((!g317) & (g374) & (!g382) & (!g1163) & (!g1422) & (!g1423)) + ((!g317) & (g374) & (!g382) & (!g1163) & (g1422) & (!g1423)) + ((!g317) & (g374) & (!g382) & (g1163) & (g1422) & (!g1423)) + ((!g317) & (g374) & (!g382) & (g1163) & (g1422) & (g1423)) + ((!g317) & (g374) & (g382) & (!g1163) & (!g1422) & (g1423)) + ((!g317) & (g374) & (g382) & (!g1163) & (g1422) & (g1423)) + ((!g317) & (g374) & (g382) & (g1163) & (!g1422) & (!g1423)) + ((!g317) & (g374) & (g382) & (g1163) & (!g1422) & (g1423)) + ((g317) & (!g374) & (!g382) & (!g1163) & (!g1422) & (!g1423)) + ((g317) & (!g374) & (!g382) & (!g1163) & (g1422) & (!g1423)) + ((g317) & (!g374) & (!g382) & (g1163) & (g1422) & (!g1423)) + ((g317) & (!g374) & (!g382) & (g1163) & (g1422) & (g1423)) + ((g317) & (!g374) & (g382) & (!g1163) & (!g1422) & (g1423)) + ((g317) & (!g374) & (g382) & (!g1163) & (g1422) & (g1423)) + ((g317) & (!g374) & (g382) & (g1163) & (!g1422) & (!g1423)) + ((g317) & (!g374) & (g382) & (g1163) & (!g1422) & (g1423)) + ((g317) & (g374) & (!g382) & (!g1163) & (!g1422) & (g1423)) + ((g317) & (g374) & (!g382) & (!g1163) & (g1422) & (g1423)) + ((g317) & (g374) & (!g382) & (g1163) & (g1422) & (!g1423)) + ((g317) & (g374) & (!g382) & (g1163) & (g1422) & (g1423)) + ((g317) & (g374) & (g382) & (!g1163) & (!g1422) & (!g1423)) + ((g317) & (g374) & (g382) & (!g1163) & (g1422) & (!g1423)) + ((g317) & (g374) & (g382) & (g1163) & (!g1422) & (!g1423)) + ((g317) & (g374) & (g382) & (g1163) & (!g1422) & (g1423)));
	assign g2111 = (((!sk[10]) & (!ld) & (text_inx29x) & (!g1425)) + ((!sk[10]) & (!ld) & (text_inx29x) & (g1425)) + ((!sk[10]) & (ld) & (!text_inx29x) & (g1425)) + ((!sk[10]) & (ld) & (text_inx29x) & (!g1425)) + ((!sk[10]) & (ld) & (text_inx29x) & (g1425)) + ((sk[10]) & (!ld) & (!text_inx29x) & (g1425)) + ((sk[10]) & (!ld) & (text_inx29x) & (g1425)) + ((sk[10]) & (ld) & (text_inx29x) & (!g1425)) + ((sk[10]) & (ld) & (text_inx29x) & (g1425)));
	assign g1426 = (((!g182) & (!sk[11]) & (g246) & (!g303)) + ((!g182) & (!sk[11]) & (g246) & (g303)) + ((!g182) & (sk[11]) & (!g246) & (g303)) + ((!g182) & (sk[11]) & (g246) & (!g303)) + ((g182) & (!sk[11]) & (!g246) & (g303)) + ((g182) & (!sk[11]) & (g246) & (!g303)) + ((g182) & (!sk[11]) & (g246) & (g303)) + ((g182) & (sk[11]) & (!g246) & (!g303)) + ((g182) & (sk[11]) & (g246) & (g303)));
	assign g1427 = (((!g310) & (!g367) & (!g375) & (!g1163) & (!g1425) & (g1426)) + ((!g310) & (!g367) & (!g375) & (!g1163) & (g1425) & (g1426)) + ((!g310) & (!g367) & (!g375) & (g1163) & (g1425) & (!g1426)) + ((!g310) & (!g367) & (!g375) & (g1163) & (g1425) & (g1426)) + ((!g310) & (!g367) & (g375) & (!g1163) & (!g1425) & (!g1426)) + ((!g310) & (!g367) & (g375) & (!g1163) & (g1425) & (!g1426)) + ((!g310) & (!g367) & (g375) & (g1163) & (!g1425) & (!g1426)) + ((!g310) & (!g367) & (g375) & (g1163) & (!g1425) & (g1426)) + ((!g310) & (g367) & (!g375) & (!g1163) & (!g1425) & (!g1426)) + ((!g310) & (g367) & (!g375) & (!g1163) & (g1425) & (!g1426)) + ((!g310) & (g367) & (!g375) & (g1163) & (g1425) & (!g1426)) + ((!g310) & (g367) & (!g375) & (g1163) & (g1425) & (g1426)) + ((!g310) & (g367) & (g375) & (!g1163) & (!g1425) & (g1426)) + ((!g310) & (g367) & (g375) & (!g1163) & (g1425) & (g1426)) + ((!g310) & (g367) & (g375) & (g1163) & (!g1425) & (!g1426)) + ((!g310) & (g367) & (g375) & (g1163) & (!g1425) & (g1426)) + ((g310) & (!g367) & (!g375) & (!g1163) & (!g1425) & (!g1426)) + ((g310) & (!g367) & (!g375) & (!g1163) & (g1425) & (!g1426)) + ((g310) & (!g367) & (!g375) & (g1163) & (g1425) & (!g1426)) + ((g310) & (!g367) & (!g375) & (g1163) & (g1425) & (g1426)) + ((g310) & (!g367) & (g375) & (!g1163) & (!g1425) & (g1426)) + ((g310) & (!g367) & (g375) & (!g1163) & (g1425) & (g1426)) + ((g310) & (!g367) & (g375) & (g1163) & (!g1425) & (!g1426)) + ((g310) & (!g367) & (g375) & (g1163) & (!g1425) & (g1426)) + ((g310) & (g367) & (!g375) & (!g1163) & (!g1425) & (g1426)) + ((g310) & (g367) & (!g375) & (!g1163) & (g1425) & (g1426)) + ((g310) & (g367) & (!g375) & (g1163) & (g1425) & (!g1426)) + ((g310) & (g367) & (!g375) & (g1163) & (g1425) & (g1426)) + ((g310) & (g367) & (g375) & (!g1163) & (!g1425) & (!g1426)) + ((g310) & (g367) & (g375) & (!g1163) & (g1425) & (!g1426)) + ((g310) & (g367) & (g375) & (g1163) & (!g1425) & (!g1426)) + ((g310) & (g367) & (g375) & (g1163) & (!g1425) & (g1426)));
	assign g2112 = (((!sk[13]) & (!ld) & (text_inx28x) & (!g1428)) + ((!sk[13]) & (!ld) & (text_inx28x) & (g1428)) + ((!sk[13]) & (ld) & (!text_inx28x) & (g1428)) + ((!sk[13]) & (ld) & (text_inx28x) & (!g1428)) + ((!sk[13]) & (ld) & (text_inx28x) & (g1428)) + ((sk[13]) & (!ld) & (!text_inx28x) & (g1428)) + ((sk[13]) & (!ld) & (text_inx28x) & (g1428)) + ((sk[13]) & (ld) & (text_inx28x) & (!g1428)) + ((sk[13]) & (ld) & (text_inx28x) & (g1428)));
	assign g1429 = (((!sk[14]) & (!g175) & (!g239) & (g296) & (!g324)) + ((!sk[14]) & (!g175) & (!g239) & (g296) & (g324)) + ((!sk[14]) & (!g175) & (g239) & (!g296) & (!g324)) + ((!sk[14]) & (!g175) & (g239) & (!g296) & (g324)) + ((!sk[14]) & (!g175) & (g239) & (g296) & (!g324)) + ((!sk[14]) & (!g175) & (g239) & (g296) & (g324)) + ((!sk[14]) & (g175) & (!g239) & (g296) & (!g324)) + ((!sk[14]) & (g175) & (!g239) & (g296) & (g324)) + ((!sk[14]) & (g175) & (g239) & (!g296) & (!g324)) + ((!sk[14]) & (g175) & (g239) & (!g296) & (g324)) + ((!sk[14]) & (g175) & (g239) & (g296) & (!g324)) + ((!sk[14]) & (g175) & (g239) & (g296) & (g324)) + ((sk[14]) & (!g175) & (!g239) & (!g296) & (g324)) + ((sk[14]) & (!g175) & (!g239) & (g296) & (!g324)) + ((sk[14]) & (!g175) & (g239) & (!g296) & (!g324)) + ((sk[14]) & (!g175) & (g239) & (g296) & (g324)) + ((sk[14]) & (g175) & (!g239) & (!g296) & (!g324)) + ((sk[14]) & (g175) & (!g239) & (g296) & (g324)) + ((sk[14]) & (g175) & (g239) & (!g296) & (g324)) + ((sk[14]) & (g175) & (g239) & (g296) & (!g324)));
	assign g2113 = (((!ld) & (!sk[15]) & (text_inx31x) & (!g1430)) + ((!ld) & (!sk[15]) & (text_inx31x) & (g1430)) + ((!ld) & (sk[15]) & (!text_inx31x) & (g1430)) + ((!ld) & (sk[15]) & (text_inx31x) & (g1430)) + ((ld) & (!sk[15]) & (!text_inx31x) & (g1430)) + ((ld) & (!sk[15]) & (text_inx31x) & (!g1430)) + ((ld) & (!sk[15]) & (text_inx31x) & (g1430)) + ((ld) & (sk[15]) & (text_inx31x) & (!g1430)) + ((ld) & (sk[15]) & (text_inx31x) & (g1430)));
	assign g1431 = (((!sk[16]) & (!g196) & (g260)) + ((!sk[16]) & (g196) & (g260)) + ((sk[16]) & (!g196) & (g260)) + ((sk[16]) & (g196) & (!g260)));
	assign g1432 = (((!sk[17]) & (!g317) & (g381)) + ((!sk[17]) & (g317) & (g381)) + ((sk[17]) & (!g317) & (g381)) + ((sk[17]) & (g317) & (!g381)));
	assign g1433 = (((!g324) & (!g389) & (!g1163) & (!g1430) & (!g1431) & (g1432)) + ((!g324) & (!g389) & (!g1163) & (!g1430) & (g1431) & (!g1432)) + ((!g324) & (!g389) & (!g1163) & (g1430) & (!g1431) & (g1432)) + ((!g324) & (!g389) & (!g1163) & (g1430) & (g1431) & (!g1432)) + ((!g324) & (!g389) & (g1163) & (g1430) & (!g1431) & (!g1432)) + ((!g324) & (!g389) & (g1163) & (g1430) & (!g1431) & (g1432)) + ((!g324) & (!g389) & (g1163) & (g1430) & (g1431) & (!g1432)) + ((!g324) & (!g389) & (g1163) & (g1430) & (g1431) & (g1432)) + ((!g324) & (g389) & (!g1163) & (!g1430) & (!g1431) & (!g1432)) + ((!g324) & (g389) & (!g1163) & (!g1430) & (g1431) & (g1432)) + ((!g324) & (g389) & (!g1163) & (g1430) & (!g1431) & (!g1432)) + ((!g324) & (g389) & (!g1163) & (g1430) & (g1431) & (g1432)) + ((!g324) & (g389) & (g1163) & (!g1430) & (!g1431) & (!g1432)) + ((!g324) & (g389) & (g1163) & (!g1430) & (!g1431) & (g1432)) + ((!g324) & (g389) & (g1163) & (!g1430) & (g1431) & (!g1432)) + ((!g324) & (g389) & (g1163) & (!g1430) & (g1431) & (g1432)) + ((g324) & (!g389) & (!g1163) & (!g1430) & (!g1431) & (!g1432)) + ((g324) & (!g389) & (!g1163) & (!g1430) & (g1431) & (g1432)) + ((g324) & (!g389) & (!g1163) & (g1430) & (!g1431) & (!g1432)) + ((g324) & (!g389) & (!g1163) & (g1430) & (g1431) & (g1432)) + ((g324) & (!g389) & (g1163) & (g1430) & (!g1431) & (!g1432)) + ((g324) & (!g389) & (g1163) & (g1430) & (!g1431) & (g1432)) + ((g324) & (!g389) & (g1163) & (g1430) & (g1431) & (!g1432)) + ((g324) & (!g389) & (g1163) & (g1430) & (g1431) & (g1432)) + ((g324) & (g389) & (!g1163) & (!g1430) & (!g1431) & (g1432)) + ((g324) & (g389) & (!g1163) & (!g1430) & (g1431) & (!g1432)) + ((g324) & (g389) & (!g1163) & (g1430) & (!g1431) & (g1432)) + ((g324) & (g389) & (!g1163) & (g1430) & (g1431) & (!g1432)) + ((g324) & (g389) & (g1163) & (!g1430) & (!g1431) & (!g1432)) + ((g324) & (g389) & (g1163) & (!g1430) & (!g1431) & (g1432)) + ((g324) & (g389) & (g1163) & (!g1430) & (g1431) & (!g1432)) + ((g324) & (g389) & (g1163) & (!g1430) & (g1431) & (g1432)));
	assign g1434 = (((!g276) & (!g283) & (!g290) & (!g297) & (g318) & (g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g318) & (!g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g318) & (g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (g318) & (!g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (!g318) & (!g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (!g318) & (g311)) + ((!g276) & (!g283) & (g290) & (g297) & (!g318) & (!g311)) + ((!g276) & (!g283) & (g290) & (g297) & (g318) & (g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (g318) & (!g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (g318) & (g311)) + ((!g276) & (g283) & (!g290) & (g297) & (g318) & (!g311)) + ((!g276) & (g283) & (!g290) & (g297) & (g318) & (g311)) + ((!g276) & (g283) & (g290) & (!g297) & (g318) & (!g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (!g318) & (!g311)) + ((g276) & (!g283) & (g290) & (!g297) & (g318) & (!g311)) + ((g276) & (!g283) & (g290) & (g297) & (!g318) & (g311)) + ((g276) & (!g283) & (g290) & (g297) & (g318) & (g311)) + ((g276) & (g283) & (!g290) & (!g297) & (!g318) & (g311)) + ((g276) & (g283) & (!g290) & (!g297) & (g318) & (!g311)) + ((g276) & (g283) & (g290) & (!g297) & (!g318) & (g311)) + ((g276) & (g283) & (g290) & (!g297) & (g318) & (!g311)) + ((g276) & (g283) & (g290) & (g297) & (!g318) & (!g311)) + ((g276) & (g283) & (g290) & (g297) & (g318) & (!g311)) + ((g276) & (g283) & (g290) & (g297) & (g318) & (g311)));
	assign g1435 = (((!g276) & (!g283) & (!g290) & (!g297) & (g318) & (!g311)) + ((!g276) & (!g283) & (!g290) & (!g297) & (g318) & (g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g318) & (!g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g318) & (g311)) + ((!g276) & (!g283) & (g290) & (g297) & (!g318) & (g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (!g318) & (!g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (!g318) & (g311)) + ((!g276) & (g283) & (g290) & (!g297) & (!g318) & (!g311)) + ((!g276) & (g283) & (g290) & (!g297) & (!g318) & (g311)) + ((!g276) & (g283) & (g290) & (!g297) & (g318) & (!g311)) + ((!g276) & (g283) & (g290) & (g297) & (g318) & (g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (!g318) & (g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (g318) & (!g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (g318) & (g311)) + ((g276) & (!g283) & (!g290) & (g297) & (g318) & (!g311)) + ((g276) & (!g283) & (g290) & (!g297) & (!g318) & (!g311)) + ((g276) & (!g283) & (g290) & (!g297) & (g318) & (g311)) + ((g276) & (!g283) & (g290) & (g297) & (!g318) & (g311)) + ((g276) & (!g283) & (g290) & (g297) & (g318) & (g311)) + ((g276) & (g283) & (!g290) & (!g297) & (!g318) & (!g311)) + ((g276) & (g283) & (!g290) & (!g297) & (!g318) & (g311)) + ((g276) & (g283) & (!g290) & (!g297) & (g318) & (!g311)) + ((g276) & (g283) & (!g290) & (!g297) & (g318) & (g311)) + ((g276) & (g283) & (!g290) & (g297) & (!g318) & (!g311)) + ((g276) & (g283) & (!g290) & (g297) & (g318) & (!g311)) + ((g276) & (g283) & (!g290) & (g297) & (g318) & (g311)) + ((g276) & (g283) & (g290) & (!g297) & (g318) & (!g311)) + ((g276) & (g283) & (g290) & (!g297) & (g318) & (g311)) + ((g276) & (g283) & (g290) & (g297) & (!g318) & (g311)) + ((g276) & (g283) & (g290) & (g297) & (g318) & (!g311)));
	assign g1436 = (((!g276) & (!g283) & (!g290) & (!g297) & (!g318) & (!g311)) + ((!g276) & (!g283) & (!g290) & (!g297) & (g318) & (g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (g318) & (g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (!g318) & (!g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (!g318) & (g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (g318) & (g311)) + ((!g276) & (!g283) & (g290) & (g297) & (!g318) & (g311)) + ((!g276) & (!g283) & (g290) & (g297) & (g318) & (!g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (!g318) & (!g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (g318) & (!g311)) + ((!g276) & (g283) & (!g290) & (g297) & (g318) & (g311)) + ((!g276) & (g283) & (g290) & (g297) & (!g318) & (!g311)) + ((!g276) & (g283) & (g290) & (g297) & (g318) & (!g311)) + ((g276) & (!g283) & (!g290) & (g297) & (!g318) & (!g311)) + ((g276) & (!g283) & (!g290) & (g297) & (!g318) & (g311)) + ((g276) & (!g283) & (!g290) & (g297) & (g318) & (!g311)) + ((g276) & (!g283) & (g290) & (!g297) & (!g318) & (!g311)) + ((g276) & (!g283) & (g290) & (!g297) & (g318) & (g311)) + ((g276) & (!g283) & (g290) & (g297) & (!g318) & (!g311)) + ((g276) & (!g283) & (g290) & (g297) & (!g318) & (g311)) + ((g276) & (!g283) & (g290) & (g297) & (g318) & (!g311)) + ((g276) & (!g283) & (g290) & (g297) & (g318) & (g311)) + ((g276) & (g283) & (!g290) & (!g297) & (g318) & (g311)) + ((g276) & (g283) & (!g290) & (g297) & (!g318) & (!g311)) + ((g276) & (g283) & (!g290) & (g297) & (g318) & (!g311)) + ((g276) & (g283) & (!g290) & (g297) & (g318) & (g311)) + ((g276) & (g283) & (g290) & (!g297) & (!g318) & (!g311)) + ((g276) & (g283) & (g290) & (g297) & (!g318) & (!g311)) + ((g276) & (g283) & (g290) & (g297) & (!g318) & (g311)) + ((g276) & (g283) & (g290) & (g297) & (g318) & (g311)));
	assign g1437 = (((!g276) & (!g283) & (!g290) & (!g297) & (!g318) & (g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (g318) & (!g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (g318) & (g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (!g318) & (g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (g318) & (g311)) + ((!g276) & (!g283) & (g290) & (g297) & (!g318) & (g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (!g318) & (!g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (!g318) & (g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (g318) & (!g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (g318) & (g311)) + ((!g276) & (g283) & (!g290) & (g297) & (g318) & (!g311)) + ((!g276) & (g283) & (!g290) & (g297) & (g318) & (g311)) + ((!g276) & (g283) & (g290) & (g297) & (!g318) & (!g311)) + ((!g276) & (g283) & (g290) & (g297) & (g318) & (!g311)) + ((!g276) & (g283) & (g290) & (g297) & (g318) & (g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (!g318) & (!g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (g318) & (g311)) + ((g276) & (!g283) & (!g290) & (g297) & (g318) & (!g311)) + ((g276) & (!g283) & (!g290) & (g297) & (g318) & (g311)) + ((g276) & (!g283) & (g290) & (!g297) & (!g318) & (g311)) + ((g276) & (!g283) & (g290) & (!g297) & (g318) & (!g311)) + ((g276) & (!g283) & (g290) & (g297) & (g318) & (!g311)) + ((g276) & (g283) & (!g290) & (!g297) & (!g318) & (g311)) + ((g276) & (g283) & (!g290) & (!g297) & (g318) & (g311)) + ((g276) & (g283) & (!g290) & (g297) & (g318) & (!g311)) + ((g276) & (g283) & (!g290) & (g297) & (g318) & (g311)) + ((g276) & (g283) & (g290) & (!g297) & (!g318) & (g311)) + ((g276) & (g283) & (g290) & (g297) & (!g318) & (!g311)));
	assign g1438 = (((!g1434) & (!g1435) & (!g1436) & (!g1437) & (!g304) & (!g325)) + ((!g1434) & (!g1435) & (!g1436) & (g1437) & (!g304) & (!g325)) + ((!g1434) & (!g1435) & (!g1436) & (g1437) & (g304) & (g325)) + ((!g1434) & (!g1435) & (g1436) & (!g1437) & (!g304) & (!g325)) + ((!g1434) & (!g1435) & (g1436) & (!g1437) & (!g304) & (g325)) + ((!g1434) & (!g1435) & (g1436) & (g1437) & (!g304) & (!g325)) + ((!g1434) & (!g1435) & (g1436) & (g1437) & (!g304) & (g325)) + ((!g1434) & (!g1435) & (g1436) & (g1437) & (g304) & (g325)) + ((!g1434) & (g1435) & (!g1436) & (!g1437) & (!g304) & (!g325)) + ((!g1434) & (g1435) & (!g1436) & (!g1437) & (g304) & (!g325)) + ((!g1434) & (g1435) & (!g1436) & (g1437) & (!g304) & (!g325)) + ((!g1434) & (g1435) & (!g1436) & (g1437) & (g304) & (!g325)) + ((!g1434) & (g1435) & (!g1436) & (g1437) & (g304) & (g325)) + ((!g1434) & (g1435) & (g1436) & (!g1437) & (!g304) & (!g325)) + ((!g1434) & (g1435) & (g1436) & (!g1437) & (!g304) & (g325)) + ((!g1434) & (g1435) & (g1436) & (!g1437) & (g304) & (!g325)) + ((!g1434) & (g1435) & (g1436) & (g1437) & (!g304) & (!g325)) + ((!g1434) & (g1435) & (g1436) & (g1437) & (!g304) & (g325)) + ((!g1434) & (g1435) & (g1436) & (g1437) & (g304) & (!g325)) + ((!g1434) & (g1435) & (g1436) & (g1437) & (g304) & (g325)) + ((g1434) & (!g1435) & (!g1436) & (g1437) & (g304) & (g325)) + ((g1434) & (!g1435) & (g1436) & (!g1437) & (!g304) & (g325)) + ((g1434) & (!g1435) & (g1436) & (g1437) & (!g304) & (g325)) + ((g1434) & (!g1435) & (g1436) & (g1437) & (g304) & (g325)) + ((g1434) & (g1435) & (!g1436) & (!g1437) & (g304) & (!g325)) + ((g1434) & (g1435) & (!g1436) & (g1437) & (g304) & (!g325)) + ((g1434) & (g1435) & (!g1436) & (g1437) & (g304) & (g325)) + ((g1434) & (g1435) & (g1436) & (!g1437) & (!g304) & (g325)) + ((g1434) & (g1435) & (g1436) & (!g1437) & (g304) & (!g325)) + ((g1434) & (g1435) & (g1436) & (g1437) & (!g304) & (g325)) + ((g1434) & (g1435) & (g1436) & (g1437) & (g304) & (!g325)) + ((g1434) & (g1435) & (g1436) & (g1437) & (g304) & (g325)));
	assign g1440 = (((!sk[24]) & (!g1108) & (g1439)) + ((!sk[24]) & (g1108) & (g1439)) + ((sk[24]) & (!g1108) & (g1439)) + ((sk[24]) & (g1108) & (!g1439)));
	assign g1441 = (((!g596) & (!sk[25]) & (!g852) & (g1438) & (!g1440)) + ((!g596) & (!sk[25]) & (!g852) & (g1438) & (g1440)) + ((!g596) & (!sk[25]) & (g852) & (!g1438) & (!g1440)) + ((!g596) & (!sk[25]) & (g852) & (!g1438) & (g1440)) + ((!g596) & (!sk[25]) & (g852) & (g1438) & (!g1440)) + ((!g596) & (!sk[25]) & (g852) & (g1438) & (g1440)) + ((!g596) & (sk[25]) & (!g852) & (!g1438) & (g1440)) + ((!g596) & (sk[25]) & (!g852) & (g1438) & (!g1440)) + ((!g596) & (sk[25]) & (g852) & (!g1438) & (!g1440)) + ((!g596) & (sk[25]) & (g852) & (g1438) & (g1440)) + ((g596) & (!sk[25]) & (!g852) & (g1438) & (!g1440)) + ((g596) & (!sk[25]) & (!g852) & (g1438) & (g1440)) + ((g596) & (!sk[25]) & (g852) & (!g1438) & (!g1440)) + ((g596) & (!sk[25]) & (g852) & (!g1438) & (g1440)) + ((g596) & (!sk[25]) & (g852) & (g1438) & (!g1440)) + ((g596) & (!sk[25]) & (g852) & (g1438) & (g1440)) + ((g596) & (sk[25]) & (!g852) & (!g1438) & (!g1440)) + ((g596) & (sk[25]) & (!g852) & (g1438) & (g1440)) + ((g596) & (sk[25]) & (g852) & (!g1438) & (g1440)) + ((g596) & (sk[25]) & (g852) & (g1438) & (!g1440)));
	assign g1442 = (((!ld) & (!sk[26]) & (!g340) & (g1441) & (!keyx24x)) + ((!ld) & (!sk[26]) & (!g340) & (g1441) & (keyx24x)) + ((!ld) & (!sk[26]) & (g340) & (!g1441) & (!keyx24x)) + ((!ld) & (!sk[26]) & (g340) & (!g1441) & (keyx24x)) + ((!ld) & (!sk[26]) & (g340) & (g1441) & (!keyx24x)) + ((!ld) & (!sk[26]) & (g340) & (g1441) & (keyx24x)) + ((!ld) & (sk[26]) & (!g340) & (g1441) & (!keyx24x)) + ((!ld) & (sk[26]) & (!g340) & (g1441) & (keyx24x)) + ((!ld) & (sk[26]) & (g340) & (!g1441) & (!keyx24x)) + ((!ld) & (sk[26]) & (g340) & (!g1441) & (keyx24x)) + ((ld) & (!sk[26]) & (!g340) & (g1441) & (!keyx24x)) + ((ld) & (!sk[26]) & (!g340) & (g1441) & (keyx24x)) + ((ld) & (!sk[26]) & (g340) & (!g1441) & (!keyx24x)) + ((ld) & (!sk[26]) & (g340) & (!g1441) & (keyx24x)) + ((ld) & (!sk[26]) & (g340) & (g1441) & (!keyx24x)) + ((ld) & (!sk[26]) & (g340) & (g1441) & (keyx24x)) + ((ld) & (sk[26]) & (!g340) & (!g1441) & (keyx24x)) + ((ld) & (sk[26]) & (!g340) & (g1441) & (keyx24x)) + ((ld) & (sk[26]) & (g340) & (!g1441) & (keyx24x)) + ((ld) & (sk[26]) & (g340) & (g1441) & (keyx24x)));
	assign g1443 = (((!g276) & (!g283) & (!g290) & (!g297) & (!g304) & (g318)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g304) & (!g318)) + ((!g276) & (!g283) & (!g290) & (g297) & (g304) & (!g318)) + ((!g276) & (!g283) & (g290) & (!g297) & (g304) & (g318)) + ((!g276) & (!g283) & (g290) & (g297) & (!g304) & (g318)) + ((!g276) & (!g283) & (g290) & (g297) & (g304) & (!g318)) + ((!g276) & (g283) & (!g290) & (!g297) & (!g304) & (g318)) + ((!g276) & (g283) & (!g290) & (!g297) & (g304) & (!g318)) + ((!g276) & (g283) & (!g290) & (!g297) & (g304) & (g318)) + ((!g276) & (g283) & (g290) & (!g297) & (g304) & (g318)) + ((!g276) & (g283) & (g290) & (g297) & (g304) & (g318)) + ((g276) & (!g283) & (!g290) & (!g297) & (!g304) & (!g318)) + ((g276) & (!g283) & (!g290) & (!g297) & (g304) & (g318)) + ((g276) & (!g283) & (!g290) & (g297) & (!g304) & (!g318)) + ((g276) & (!g283) & (!g290) & (g297) & (g304) & (!g318)) + ((g276) & (!g283) & (g290) & (!g297) & (g304) & (!g318)) + ((g276) & (!g283) & (g290) & (!g297) & (g304) & (g318)) + ((g276) & (!g283) & (g290) & (g297) & (g304) & (!g318)) + ((g276) & (!g283) & (g290) & (g297) & (g304) & (g318)) + ((g276) & (g283) & (!g290) & (!g297) & (g304) & (!g318)) + ((g276) & (g283) & (!g290) & (!g297) & (g304) & (g318)) + ((g276) & (g283) & (!g290) & (g297) & (g304) & (g318)) + ((g276) & (g283) & (g290) & (!g297) & (!g304) & (!g318)) + ((g276) & (g283) & (g290) & (!g297) & (!g304) & (g318)) + ((g276) & (g283) & (g290) & (!g297) & (g304) & (!g318)) + ((g276) & (g283) & (g290) & (g297) & (!g304) & (g318)) + ((g276) & (g283) & (g290) & (g297) & (g304) & (!g318)));
	assign g1444 = (((!g276) & (!g283) & (!g290) & (!g297) & (!g304) & (g318)) + ((!g276) & (!g283) & (!g290) & (!g297) & (g304) & (!g318)) + ((!g276) & (!g283) & (!g290) & (!g297) & (g304) & (g318)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g304) & (!g318)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g304) & (g318)) + ((!g276) & (!g283) & (!g290) & (g297) & (g304) & (g318)) + ((!g276) & (!g283) & (g290) & (!g297) & (g304) & (!g318)) + ((!g276) & (!g283) & (g290) & (g297) & (!g304) & (!g318)) + ((!g276) & (!g283) & (g290) & (g297) & (!g304) & (g318)) + ((!g276) & (!g283) & (g290) & (g297) & (g304) & (g318)) + ((!g276) & (g283) & (!g290) & (!g297) & (g304) & (g318)) + ((!g276) & (g283) & (!g290) & (g297) & (!g304) & (!g318)) + ((!g276) & (g283) & (!g290) & (g297) & (g304) & (!g318)) + ((!g276) & (g283) & (g290) & (!g297) & (g304) & (!g318)) + ((!g276) & (g283) & (g290) & (!g297) & (g304) & (g318)) + ((!g276) & (g283) & (g290) & (g297) & (!g304) & (!g318)) + ((g276) & (!g283) & (!g290) & (!g297) & (!g304) & (!g318)) + ((g276) & (!g283) & (!g290) & (g297) & (!g304) & (!g318)) + ((g276) & (!g283) & (!g290) & (g297) & (!g304) & (g318)) + ((g276) & (!g283) & (g290) & (!g297) & (!g304) & (g318)) + ((g276) & (!g283) & (g290) & (!g297) & (g304) & (g318)) + ((g276) & (!g283) & (g290) & (g297) & (!g304) & (!g318)) + ((g276) & (!g283) & (g290) & (g297) & (!g304) & (g318)) + ((g276) & (g283) & (!g290) & (g297) & (!g304) & (!g318)) + ((g276) & (g283) & (!g290) & (g297) & (g304) & (g318)) + ((g276) & (g283) & (g290) & (!g297) & (!g304) & (!g318)) + ((g276) & (g283) & (g290) & (!g297) & (!g304) & (g318)) + ((g276) & (g283) & (g290) & (!g297) & (g304) & (g318)) + ((g276) & (g283) & (g290) & (g297) & (!g304) & (!g318)) + ((g276) & (g283) & (g290) & (g297) & (!g304) & (g318)) + ((g276) & (g283) & (g290) & (g297) & (g304) & (!g318)));
	assign g1445 = (((!g276) & (!g283) & (!g290) & (!g297) & (!g304) & (g318)) + ((!g276) & (!g283) & (!g290) & (g297) & (g304) & (!g318)) + ((!g276) & (!g283) & (g290) & (!g297) & (!g304) & (!g318)) + ((!g276) & (!g283) & (g290) & (!g297) & (g304) & (!g318)) + ((!g276) & (!g283) & (g290) & (g297) & (!g304) & (g318)) + ((!g276) & (!g283) & (g290) & (g297) & (g304) & (!g318)) + ((!g276) & (!g283) & (g290) & (g297) & (g304) & (g318)) + ((!g276) & (g283) & (!g290) & (!g297) & (!g304) & (!g318)) + ((!g276) & (g283) & (!g290) & (!g297) & (g304) & (!g318)) + ((!g276) & (g283) & (!g290) & (g297) & (!g304) & (!g318)) + ((!g276) & (g283) & (!g290) & (g297) & (g304) & (g318)) + ((!g276) & (g283) & (g290) & (!g297) & (g304) & (g318)) + ((!g276) & (g283) & (g290) & (g297) & (!g304) & (g318)) + ((!g276) & (g283) & (g290) & (g297) & (g304) & (!g318)) + ((g276) & (!g283) & (!g290) & (!g297) & (g304) & (g318)) + ((g276) & (!g283) & (!g290) & (g297) & (!g304) & (!g318)) + ((g276) & (!g283) & (!g290) & (g297) & (g304) & (!g318)) + ((g276) & (!g283) & (g290) & (!g297) & (!g304) & (!g318)) + ((g276) & (!g283) & (g290) & (!g297) & (!g304) & (g318)) + ((g276) & (!g283) & (g290) & (!g297) & (g304) & (!g318)) + ((g276) & (!g283) & (g290) & (!g297) & (g304) & (g318)) + ((g276) & (!g283) & (g290) & (g297) & (g304) & (!g318)) + ((g276) & (g283) & (!g290) & (!g297) & (!g304) & (g318)) + ((g276) & (g283) & (!g290) & (!g297) & (g304) & (g318)) + ((g276) & (g283) & (!g290) & (g297) & (!g304) & (g318)) + ((g276) & (g283) & (g290) & (!g297) & (!g304) & (!g318)) + ((g276) & (g283) & (g290) & (!g297) & (!g304) & (g318)) + ((g276) & (g283) & (g290) & (!g297) & (g304) & (g318)) + ((g276) & (g283) & (g290) & (g297) & (!g304) & (!g318)) + ((g276) & (g283) & (g290) & (g297) & (!g304) & (g318)) + ((g276) & (g283) & (g290) & (g297) & (g304) & (!g318)) + ((g276) & (g283) & (g290) & (g297) & (g304) & (g318)));
	assign g1446 = (((!g276) & (!g283) & (!g290) & (!g297) & (g304) & (!g318)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g304) & (!g318)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g304) & (g318)) + ((!g276) & (!g283) & (g290) & (!g297) & (g304) & (g318)) + ((!g276) & (!g283) & (g290) & (g297) & (!g304) & (g318)) + ((!g276) & (g283) & (!g290) & (!g297) & (!g304) & (!g318)) + ((!g276) & (g283) & (!g290) & (!g297) & (g304) & (!g318)) + ((!g276) & (g283) & (!g290) & (g297) & (!g304) & (g318)) + ((!g276) & (g283) & (g290) & (!g297) & (!g304) & (g318)) + ((!g276) & (g283) & (g290) & (!g297) & (g304) & (!g318)) + ((!g276) & (g283) & (g290) & (!g297) & (g304) & (g318)) + ((!g276) & (g283) & (g290) & (g297) & (g304) & (!g318)) + ((!g276) & (g283) & (g290) & (g297) & (g304) & (g318)) + ((g276) & (!g283) & (!g290) & (!g297) & (!g304) & (!g318)) + ((g276) & (!g283) & (!g290) & (g297) & (!g304) & (!g318)) + ((g276) & (!g283) & (!g290) & (g297) & (!g304) & (g318)) + ((g276) & (!g283) & (!g290) & (g297) & (g304) & (!g318)) + ((g276) & (!g283) & (g290) & (!g297) & (!g304) & (!g318)) + ((g276) & (!g283) & (g290) & (!g297) & (g304) & (g318)) + ((g276) & (!g283) & (g290) & (g297) & (g304) & (!g318)) + ((g276) & (g283) & (!g290) & (!g297) & (!g304) & (!g318)) + ((g276) & (g283) & (!g290) & (g297) & (!g304) & (!g318)) + ((g276) & (g283) & (!g290) & (g297) & (g304) & (!g318)) + ((g276) & (g283) & (!g290) & (g297) & (g304) & (g318)) + ((g276) & (g283) & (g290) & (g297) & (!g304) & (g318)) + ((g276) & (g283) & (g290) & (g297) & (g304) & (g318)));
	assign g1447 = (((!g1443) & (!g1444) & (!g1445) & (!g1446) & (!g311) & (!g325)) + ((!g1443) & (!g1444) & (!g1445) & (!g1446) & (g311) & (!g325)) + ((!g1443) & (!g1444) & (!g1445) & (g1446) & (!g311) & (!g325)) + ((!g1443) & (!g1444) & (!g1445) & (g1446) & (g311) & (!g325)) + ((!g1443) & (!g1444) & (!g1445) & (g1446) & (g311) & (g325)) + ((!g1443) & (!g1444) & (g1445) & (!g1446) & (!g311) & (!g325)) + ((!g1443) & (!g1444) & (g1445) & (!g1446) & (!g311) & (g325)) + ((!g1443) & (!g1444) & (g1445) & (!g1446) & (g311) & (!g325)) + ((!g1443) & (!g1444) & (g1445) & (g1446) & (!g311) & (!g325)) + ((!g1443) & (!g1444) & (g1445) & (g1446) & (!g311) & (g325)) + ((!g1443) & (!g1444) & (g1445) & (g1446) & (g311) & (!g325)) + ((!g1443) & (!g1444) & (g1445) & (g1446) & (g311) & (g325)) + ((!g1443) & (g1444) & (!g1445) & (!g1446) & (!g311) & (!g325)) + ((!g1443) & (g1444) & (!g1445) & (g1446) & (!g311) & (!g325)) + ((!g1443) & (g1444) & (!g1445) & (g1446) & (g311) & (g325)) + ((!g1443) & (g1444) & (g1445) & (!g1446) & (!g311) & (!g325)) + ((!g1443) & (g1444) & (g1445) & (!g1446) & (!g311) & (g325)) + ((!g1443) & (g1444) & (g1445) & (g1446) & (!g311) & (!g325)) + ((!g1443) & (g1444) & (g1445) & (g1446) & (!g311) & (g325)) + ((!g1443) & (g1444) & (g1445) & (g1446) & (g311) & (g325)) + ((g1443) & (!g1444) & (!g1445) & (!g1446) & (g311) & (!g325)) + ((g1443) & (!g1444) & (!g1445) & (g1446) & (g311) & (!g325)) + ((g1443) & (!g1444) & (!g1445) & (g1446) & (g311) & (g325)) + ((g1443) & (!g1444) & (g1445) & (!g1446) & (!g311) & (g325)) + ((g1443) & (!g1444) & (g1445) & (!g1446) & (g311) & (!g325)) + ((g1443) & (!g1444) & (g1445) & (g1446) & (!g311) & (g325)) + ((g1443) & (!g1444) & (g1445) & (g1446) & (g311) & (!g325)) + ((g1443) & (!g1444) & (g1445) & (g1446) & (g311) & (g325)) + ((g1443) & (g1444) & (!g1445) & (g1446) & (g311) & (g325)) + ((g1443) & (g1444) & (g1445) & (!g1446) & (!g311) & (g325)) + ((g1443) & (g1444) & (g1445) & (g1446) & (!g311) & (g325)) + ((g1443) & (g1444) & (g1445) & (g1446) & (g311) & (g325)));
	assign g1449 = (((!g1115) & (!sk[32]) & (g1448)) + ((!g1115) & (sk[32]) & (g1448)) + ((g1115) & (!sk[32]) & (g1448)) + ((g1115) & (sk[32]) & (!g1448)));
	assign g1450 = (((!sk[33]) & (!g603) & (!g859) & (g1447) & (!g1449)) + ((!sk[33]) & (!g603) & (!g859) & (g1447) & (g1449)) + ((!sk[33]) & (!g603) & (g859) & (!g1447) & (!g1449)) + ((!sk[33]) & (!g603) & (g859) & (!g1447) & (g1449)) + ((!sk[33]) & (!g603) & (g859) & (g1447) & (!g1449)) + ((!sk[33]) & (!g603) & (g859) & (g1447) & (g1449)) + ((!sk[33]) & (g603) & (!g859) & (g1447) & (!g1449)) + ((!sk[33]) & (g603) & (!g859) & (g1447) & (g1449)) + ((!sk[33]) & (g603) & (g859) & (!g1447) & (!g1449)) + ((!sk[33]) & (g603) & (g859) & (!g1447) & (g1449)) + ((!sk[33]) & (g603) & (g859) & (g1447) & (!g1449)) + ((!sk[33]) & (g603) & (g859) & (g1447) & (g1449)) + ((sk[33]) & (!g603) & (!g859) & (!g1447) & (g1449)) + ((sk[33]) & (!g603) & (!g859) & (g1447) & (!g1449)) + ((sk[33]) & (!g603) & (g859) & (!g1447) & (!g1449)) + ((sk[33]) & (!g603) & (g859) & (g1447) & (g1449)) + ((sk[33]) & (g603) & (!g859) & (!g1447) & (!g1449)) + ((sk[33]) & (g603) & (!g859) & (g1447) & (g1449)) + ((sk[33]) & (g603) & (g859) & (!g1447) & (g1449)) + ((sk[33]) & (g603) & (g859) & (g1447) & (!g1449)));
	assign g1451 = (((!ld) & (!sk[34]) & (!g347) & (g1450) & (!keyx25x)) + ((!ld) & (!sk[34]) & (!g347) & (g1450) & (keyx25x)) + ((!ld) & (!sk[34]) & (g347) & (!g1450) & (!keyx25x)) + ((!ld) & (!sk[34]) & (g347) & (!g1450) & (keyx25x)) + ((!ld) & (!sk[34]) & (g347) & (g1450) & (!keyx25x)) + ((!ld) & (!sk[34]) & (g347) & (g1450) & (keyx25x)) + ((!ld) & (sk[34]) & (!g347) & (g1450) & (!keyx25x)) + ((!ld) & (sk[34]) & (!g347) & (g1450) & (keyx25x)) + ((!ld) & (sk[34]) & (g347) & (!g1450) & (!keyx25x)) + ((!ld) & (sk[34]) & (g347) & (!g1450) & (keyx25x)) + ((ld) & (!sk[34]) & (!g347) & (g1450) & (!keyx25x)) + ((ld) & (!sk[34]) & (!g347) & (g1450) & (keyx25x)) + ((ld) & (!sk[34]) & (g347) & (!g1450) & (!keyx25x)) + ((ld) & (!sk[34]) & (g347) & (!g1450) & (keyx25x)) + ((ld) & (!sk[34]) & (g347) & (g1450) & (!keyx25x)) + ((ld) & (!sk[34]) & (g347) & (g1450) & (keyx25x)) + ((ld) & (sk[34]) & (!g347) & (!g1450) & (keyx25x)) + ((ld) & (sk[34]) & (!g347) & (g1450) & (keyx25x)) + ((ld) & (sk[34]) & (g347) & (!g1450) & (keyx25x)) + ((ld) & (sk[34]) & (g347) & (g1450) & (keyx25x)));
	assign g1452 = (((!g318) & (!g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((!g318) & (!g283) & (!g290) & (!g297) & (g304) & (g311)) + ((!g318) & (!g283) & (!g290) & (g297) & (!g304) & (g311)) + ((!g318) & (!g283) & (!g290) & (g297) & (g304) & (!g311)) + ((!g318) & (!g283) & (!g290) & (g297) & (g304) & (g311)) + ((!g318) & (!g283) & (g290) & (!g297) & (!g304) & (g311)) + ((!g318) & (!g283) & (g290) & (g297) & (!g304) & (!g311)) + ((!g318) & (!g283) & (g290) & (g297) & (g304) & (!g311)) + ((!g318) & (g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((!g318) & (g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((!g318) & (g283) & (!g290) & (g297) & (!g304) & (g311)) + ((!g318) & (g283) & (g290) & (!g297) & (!g304) & (!g311)) + ((!g318) & (g283) & (g290) & (!g297) & (!g304) & (g311)) + ((!g318) & (g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g318) & (g283) & (g290) & (!g297) & (g304) & (g311)) + ((g318) & (!g283) & (!g290) & (g297) & (!g304) & (g311)) + ((g318) & (!g283) & (!g290) & (g297) & (g304) & (g311)) + ((g318) & (g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((g318) & (g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((g318) & (g283) & (!g290) & (g297) & (g304) & (!g311)) + ((g318) & (g283) & (g290) & (g297) & (!g304) & (!g311)) + ((g318) & (g283) & (g290) & (g297) & (!g304) & (g311)));
	assign g1453 = (((!g318) & (!g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((!g318) & (!g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((!g318) & (!g283) & (!g290) & (g297) & (g304) & (g311)) + ((!g318) & (!g283) & (g290) & (!g297) & (!g304) & (!g311)) + ((!g318) & (!g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g318) & (!g283) & (g290) & (g297) & (!g304) & (g311)) + ((!g318) & (g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((!g318) & (g283) & (!g290) & (!g297) & (g304) & (g311)) + ((!g318) & (g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((!g318) & (g283) & (!g290) & (g297) & (!g304) & (g311)) + ((!g318) & (g283) & (!g290) & (g297) & (g304) & (g311)) + ((!g318) & (g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g318) & (g283) & (g290) & (!g297) & (g304) & (g311)) + ((!g318) & (g283) & (g290) & (g297) & (g304) & (!g311)) + ((g318) & (!g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((g318) & (!g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((g318) & (!g283) & (!g290) & (!g297) & (g304) & (g311)) + ((g318) & (!g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((g318) & (!g283) & (!g290) & (g297) & (!g304) & (g311)) + ((g318) & (!g283) & (!g290) & (g297) & (g304) & (!g311)) + ((g318) & (!g283) & (g290) & (g297) & (!g304) & (!g311)) + ((g318) & (g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((g318) & (g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((g318) & (g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((g318) & (g283) & (!g290) & (g297) & (g304) & (!g311)) + ((g318) & (g283) & (!g290) & (g297) & (g304) & (g311)) + ((g318) & (g283) & (g290) & (!g297) & (!g304) & (!g311)) + ((g318) & (g283) & (g290) & (!g297) & (g304) & (!g311)) + ((g318) & (g283) & (g290) & (g297) & (!g304) & (g311)) + ((g318) & (g283) & (g290) & (g297) & (g304) & (g311)));
	assign g1454 = (((!g318) & (!g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((!g318) & (!g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((!g318) & (!g283) & (!g290) & (g297) & (!g304) & (g311)) + ((!g318) & (!g283) & (g290) & (!g297) & (!g304) & (g311)) + ((!g318) & (!g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g318) & (!g283) & (g290) & (g297) & (!g304) & (g311)) + ((!g318) & (g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((!g318) & (g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((!g318) & (g283) & (!g290) & (g297) & (g304) & (!g311)) + ((!g318) & (g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g318) & (g283) & (g290) & (g297) & (!g304) & (!g311)) + ((!g318) & (g283) & (g290) & (g297) & (g304) & (!g311)) + ((g318) & (!g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((g318) & (!g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((g318) & (!g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((g318) & (!g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((g318) & (!g283) & (!g290) & (g297) & (!g304) & (g311)) + ((g318) & (!g283) & (!g290) & (g297) & (g304) & (!g311)) + ((g318) & (!g283) & (!g290) & (g297) & (g304) & (g311)) + ((g318) & (!g283) & (g290) & (!g297) & (!g304) & (g311)) + ((g318) & (!g283) & (g290) & (!g297) & (g304) & (!g311)) + ((g318) & (!g283) & (g290) & (g297) & (!g304) & (!g311)) + ((g318) & (!g283) & (g290) & (g297) & (g304) & (g311)) + ((g318) & (g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((g318) & (g283) & (!g290) & (!g297) & (g304) & (g311)) + ((g318) & (g283) & (g290) & (!g297) & (g304) & (g311)) + ((g318) & (g283) & (g290) & (g297) & (!g304) & (!g311)) + ((g318) & (g283) & (g290) & (g297) & (!g304) & (g311)) + ((g318) & (g283) & (g290) & (g297) & (g304) & (g311)));
	assign g1455 = (((!g318) & (!g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((!g318) & (!g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((!g318) & (!g283) & (!g290) & (!g297) & (g304) & (g311)) + ((!g318) & (!g283) & (!g290) & (g297) & (!g304) & (g311)) + ((!g318) & (!g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g318) & (!g283) & (g290) & (g297) & (g304) & (g311)) + ((!g318) & (g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((!g318) & (g283) & (!g290) & (g297) & (!g304) & (g311)) + ((!g318) & (g283) & (!g290) & (g297) & (g304) & (g311)) + ((!g318) & (g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g318) & (g283) & (g290) & (!g297) & (g304) & (g311)) + ((!g318) & (g283) & (g290) & (g297) & (!g304) & (!g311)) + ((!g318) & (g283) & (g290) & (g297) & (!g304) & (g311)) + ((!g318) & (g283) & (g290) & (g297) & (g304) & (!g311)) + ((!g318) & (g283) & (g290) & (g297) & (g304) & (g311)) + ((g318) & (!g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((g318) & (!g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((g318) & (!g283) & (!g290) & (!g297) & (g304) & (g311)) + ((g318) & (!g283) & (!g290) & (g297) & (g304) & (g311)) + ((g318) & (!g283) & (g290) & (!g297) & (!g304) & (g311)) + ((g318) & (!g283) & (g290) & (!g297) & (g304) & (!g311)) + ((g318) & (!g283) & (g290) & (g297) & (g304) & (!g311)) + ((g318) & (g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((g318) & (g283) & (!g290) & (g297) & (!g304) & (g311)) + ((g318) & (g283) & (!g290) & (g297) & (g304) & (!g311)) + ((g318) & (g283) & (g290) & (!g297) & (g304) & (g311)) + ((g318) & (g283) & (g290) & (g297) & (!g304) & (!g311)));
	assign g1456 = (((!g1452) & (!g1453) & (!g1454) & (!g1455) & (!g276) & (g325)) + ((!g1452) & (!g1453) & (!g1454) & (!g1455) & (g276) & (!g325)) + ((!g1452) & (!g1453) & (!g1454) & (!g1455) & (g276) & (g325)) + ((!g1452) & (!g1453) & (!g1454) & (g1455) & (!g276) & (g325)) + ((!g1452) & (!g1453) & (!g1454) & (g1455) & (g276) & (!g325)) + ((!g1452) & (!g1453) & (g1454) & (!g1455) & (g276) & (!g325)) + ((!g1452) & (!g1453) & (g1454) & (!g1455) & (g276) & (g325)) + ((!g1452) & (!g1453) & (g1454) & (g1455) & (g276) & (!g325)) + ((!g1452) & (g1453) & (!g1454) & (!g1455) & (!g276) & (g325)) + ((!g1452) & (g1453) & (!g1454) & (!g1455) & (g276) & (g325)) + ((!g1452) & (g1453) & (!g1454) & (g1455) & (!g276) & (g325)) + ((!g1452) & (g1453) & (g1454) & (!g1455) & (g276) & (g325)) + ((g1452) & (!g1453) & (!g1454) & (!g1455) & (!g276) & (!g325)) + ((g1452) & (!g1453) & (!g1454) & (!g1455) & (!g276) & (g325)) + ((g1452) & (!g1453) & (!g1454) & (!g1455) & (g276) & (!g325)) + ((g1452) & (!g1453) & (!g1454) & (!g1455) & (g276) & (g325)) + ((g1452) & (!g1453) & (!g1454) & (g1455) & (!g276) & (!g325)) + ((g1452) & (!g1453) & (!g1454) & (g1455) & (!g276) & (g325)) + ((g1452) & (!g1453) & (!g1454) & (g1455) & (g276) & (!g325)) + ((g1452) & (!g1453) & (g1454) & (!g1455) & (!g276) & (!g325)) + ((g1452) & (!g1453) & (g1454) & (!g1455) & (g276) & (!g325)) + ((g1452) & (!g1453) & (g1454) & (!g1455) & (g276) & (g325)) + ((g1452) & (!g1453) & (g1454) & (g1455) & (!g276) & (!g325)) + ((g1452) & (!g1453) & (g1454) & (g1455) & (g276) & (!g325)) + ((g1452) & (g1453) & (!g1454) & (!g1455) & (!g276) & (!g325)) + ((g1452) & (g1453) & (!g1454) & (!g1455) & (!g276) & (g325)) + ((g1452) & (g1453) & (!g1454) & (!g1455) & (g276) & (g325)) + ((g1452) & (g1453) & (!g1454) & (g1455) & (!g276) & (!g325)) + ((g1452) & (g1453) & (!g1454) & (g1455) & (!g276) & (g325)) + ((g1452) & (g1453) & (g1454) & (!g1455) & (!g276) & (!g325)) + ((g1452) & (g1453) & (g1454) & (!g1455) & (g276) & (g325)) + ((g1452) & (g1453) & (g1454) & (g1455) & (!g276) & (!g325)));
	assign g1458 = (((!sk[40]) & (!g1122) & (g1457)) + ((!sk[40]) & (g1122) & (g1457)) + ((sk[40]) & (!g1122) & (g1457)) + ((sk[40]) & (g1122) & (!g1457)));
	assign g1459 = (((!g610) & (!g866) & (!sk[41]) & (g1456) & (!g1458)) + ((!g610) & (!g866) & (!sk[41]) & (g1456) & (g1458)) + ((!g610) & (!g866) & (sk[41]) & (!g1456) & (g1458)) + ((!g610) & (!g866) & (sk[41]) & (g1456) & (!g1458)) + ((!g610) & (g866) & (!sk[41]) & (!g1456) & (!g1458)) + ((!g610) & (g866) & (!sk[41]) & (!g1456) & (g1458)) + ((!g610) & (g866) & (!sk[41]) & (g1456) & (!g1458)) + ((!g610) & (g866) & (!sk[41]) & (g1456) & (g1458)) + ((!g610) & (g866) & (sk[41]) & (!g1456) & (!g1458)) + ((!g610) & (g866) & (sk[41]) & (g1456) & (g1458)) + ((g610) & (!g866) & (!sk[41]) & (g1456) & (!g1458)) + ((g610) & (!g866) & (!sk[41]) & (g1456) & (g1458)) + ((g610) & (!g866) & (sk[41]) & (!g1456) & (!g1458)) + ((g610) & (!g866) & (sk[41]) & (g1456) & (g1458)) + ((g610) & (g866) & (!sk[41]) & (!g1456) & (!g1458)) + ((g610) & (g866) & (!sk[41]) & (!g1456) & (g1458)) + ((g610) & (g866) & (!sk[41]) & (g1456) & (!g1458)) + ((g610) & (g866) & (!sk[41]) & (g1456) & (g1458)) + ((g610) & (g866) & (sk[41]) & (!g1456) & (g1458)) + ((g610) & (g866) & (sk[41]) & (g1456) & (!g1458)));
	assign g1460 = (((!ld) & (!g354) & (g1459) & (!sk[42]) & (!keyx26x)) + ((!ld) & (!g354) & (g1459) & (!sk[42]) & (keyx26x)) + ((!ld) & (!g354) & (g1459) & (sk[42]) & (!keyx26x)) + ((!ld) & (!g354) & (g1459) & (sk[42]) & (keyx26x)) + ((!ld) & (g354) & (!g1459) & (!sk[42]) & (!keyx26x)) + ((!ld) & (g354) & (!g1459) & (!sk[42]) & (keyx26x)) + ((!ld) & (g354) & (!g1459) & (sk[42]) & (!keyx26x)) + ((!ld) & (g354) & (!g1459) & (sk[42]) & (keyx26x)) + ((!ld) & (g354) & (g1459) & (!sk[42]) & (!keyx26x)) + ((!ld) & (g354) & (g1459) & (!sk[42]) & (keyx26x)) + ((ld) & (!g354) & (!g1459) & (sk[42]) & (keyx26x)) + ((ld) & (!g354) & (g1459) & (!sk[42]) & (!keyx26x)) + ((ld) & (!g354) & (g1459) & (!sk[42]) & (keyx26x)) + ((ld) & (!g354) & (g1459) & (sk[42]) & (keyx26x)) + ((ld) & (g354) & (!g1459) & (!sk[42]) & (!keyx26x)) + ((ld) & (g354) & (!g1459) & (!sk[42]) & (keyx26x)) + ((ld) & (g354) & (!g1459) & (sk[42]) & (keyx26x)) + ((ld) & (g354) & (g1459) & (!sk[42]) & (!keyx26x)) + ((ld) & (g354) & (g1459) & (!sk[42]) & (keyx26x)) + ((ld) & (g354) & (g1459) & (sk[42]) & (keyx26x)));
	assign g1461 = (((!g276) & (!g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (g304) & (g311)) + ((!g276) & (!g283) & (g290) & (g297) & (!g304) & (!g311)) + ((!g276) & (!g283) & (g290) & (g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (g290) & (g297) & (g304) & (g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (g283) & (g290) & (!g297) & (!g304) & (!g311)) + ((!g276) & (g283) & (g290) & (g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((g276) & (!g283) & (g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (g290) & (!g297) & (!g304) & (g311)) + ((g276) & (!g283) & (g290) & (!g297) & (g304) & (!g311)) + ((g276) & (!g283) & (g290) & (g297) & (!g304) & (g311)) + ((g276) & (g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((g276) & (g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((g276) & (g283) & (!g290) & (g297) & (g304) & (!g311)) + ((g276) & (g283) & (g290) & (!g297) & (!g304) & (g311)) + ((g276) & (g283) & (g290) & (!g297) & (g304) & (g311)));
	assign g1462 = (((!g276) & (!g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (!g290) & (!g297) & (g304) & (g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (g290) & (g297) & (!g304) & (!g311)) + ((!g276) & (!g283) & (g290) & (g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (g290) & (g297) & (g304) & (g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (g304) & (g311)) + ((!g276) & (g283) & (!g290) & (g297) & (g304) & (g311)) + ((!g276) & (g283) & (g290) & (!g297) & (!g304) & (!g311)) + ((!g276) & (g283) & (g290) & (!g297) & (!g304) & (g311)) + ((!g276) & (g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (g283) & (g290) & (g297) & (!g304) & (g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((g276) & (!g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (!g290) & (g297) & (!g304) & (g311)) + ((g276) & (!g283) & (!g290) & (g297) & (g304) & (g311)) + ((g276) & (!g283) & (g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (g290) & (!g297) & (!g304) & (g311)) + ((g276) & (!g283) & (g290) & (!g297) & (g304) & (g311)) + ((g276) & (!g283) & (g290) & (g297) & (!g304) & (g311)) + ((g276) & (g283) & (!g290) & (g297) & (!g304) & (g311)) + ((g276) & (g283) & (!g290) & (g297) & (g304) & (!g311)) + ((g276) & (g283) & (g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (g283) & (g290) & (g297) & (!g304) & (!g311)));
	assign g1463 = (((!g276) & (!g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (!g290) & (!g297) & (g304) & (g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (g290) & (!g297) & (g304) & (g311)) + ((!g276) & (!g283) & (g290) & (g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (g290) & (g297) & (g304) & (g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (g304) & (g311)) + ((!g276) & (g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((!g276) & (g283) & (!g290) & (g297) & (!g304) & (g311)) + ((!g276) & (g283) & (g290) & (!g297) & (!g304) & (g311)) + ((!g276) & (g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (g283) & (g290) & (g297) & (g304) & (g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (g304) & (g311)) + ((g276) & (!g283) & (!g290) & (g297) & (g304) & (g311)) + ((g276) & (!g283) & (g290) & (g297) & (!g304) & (!g311)) + ((g276) & (g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((g276) & (g283) & (!g290) & (g297) & (g304) & (g311)) + ((g276) & (g283) & (g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (g283) & (g290) & (!g297) & (!g304) & (g311)) + ((g276) & (g283) & (g290) & (!g297) & (g304) & (g311)) + ((g276) & (g283) & (g290) & (g297) & (!g304) & (!g311)) + ((g276) & (g283) & (g290) & (g297) & (g304) & (g311)));
	assign g1464 = (((!g276) & (!g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (!g290) & (g297) & (g304) & (g311)) + ((!g276) & (!g283) & (g290) & (g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (g290) & (g297) & (g304) & (g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (!g304) & (!g311)) + ((!g276) & (g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (g283) & (!g290) & (g297) & (!g304) & (!g311)) + ((!g276) & (g283) & (!g290) & (g297) & (!g304) & (g311)) + ((!g276) & (g283) & (!g290) & (g297) & (g304) & (!g311)) + ((!g276) & (g283) & (g290) & (!g297) & (!g304) & (!g311)) + ((!g276) & (g283) & (g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (g283) & (g290) & (!g297) & (g304) & (g311)) + ((g276) & (!g283) & (!g290) & (!g297) & (g304) & (g311)) + ((g276) & (!g283) & (!g290) & (g297) & (g304) & (!g311)) + ((g276) & (!g283) & (g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (g290) & (!g297) & (g304) & (!g311)) + ((g276) & (!g283) & (g290) & (!g297) & (g304) & (g311)) + ((g276) & (!g283) & (g290) & (g297) & (!g304) & (g311)) + ((g276) & (!g283) & (g290) & (g297) & (g304) & (!g311)) + ((g276) & (!g283) & (g290) & (g297) & (g304) & (g311)) + ((g276) & (g283) & (!g290) & (!g297) & (!g304) & (g311)) + ((g276) & (g283) & (!g290) & (!g297) & (g304) & (!g311)) + ((g276) & (g283) & (g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (g283) & (g290) & (!g297) & (!g304) & (g311)) + ((g276) & (g283) & (g290) & (g297) & (g304) & (g311)));
	assign g1465 = (((!g1461) & (!g1462) & (!g1463) & (!g1464) & (!g325) & (g318)) + ((!g1461) & (!g1462) & (!g1463) & (!g1464) & (g325) & (!g318)) + ((!g1461) & (!g1462) & (!g1463) & (!g1464) & (g325) & (g318)) + ((!g1461) & (!g1462) & (!g1463) & (g1464) & (!g325) & (g318)) + ((!g1461) & (!g1462) & (!g1463) & (g1464) & (g325) & (!g318)) + ((!g1461) & (!g1462) & (g1463) & (!g1464) & (g325) & (!g318)) + ((!g1461) & (!g1462) & (g1463) & (!g1464) & (g325) & (g318)) + ((!g1461) & (!g1462) & (g1463) & (g1464) & (g325) & (!g318)) + ((!g1461) & (g1462) & (!g1463) & (!g1464) & (!g325) & (g318)) + ((!g1461) & (g1462) & (!g1463) & (!g1464) & (g325) & (g318)) + ((!g1461) & (g1462) & (!g1463) & (g1464) & (!g325) & (g318)) + ((!g1461) & (g1462) & (g1463) & (!g1464) & (g325) & (g318)) + ((g1461) & (!g1462) & (!g1463) & (!g1464) & (!g325) & (!g318)) + ((g1461) & (!g1462) & (!g1463) & (!g1464) & (!g325) & (g318)) + ((g1461) & (!g1462) & (!g1463) & (!g1464) & (g325) & (!g318)) + ((g1461) & (!g1462) & (!g1463) & (!g1464) & (g325) & (g318)) + ((g1461) & (!g1462) & (!g1463) & (g1464) & (!g325) & (!g318)) + ((g1461) & (!g1462) & (!g1463) & (g1464) & (!g325) & (g318)) + ((g1461) & (!g1462) & (!g1463) & (g1464) & (g325) & (!g318)) + ((g1461) & (!g1462) & (g1463) & (!g1464) & (!g325) & (!g318)) + ((g1461) & (!g1462) & (g1463) & (!g1464) & (g325) & (!g318)) + ((g1461) & (!g1462) & (g1463) & (!g1464) & (g325) & (g318)) + ((g1461) & (!g1462) & (g1463) & (g1464) & (!g325) & (!g318)) + ((g1461) & (!g1462) & (g1463) & (g1464) & (g325) & (!g318)) + ((g1461) & (g1462) & (!g1463) & (!g1464) & (!g325) & (!g318)) + ((g1461) & (g1462) & (!g1463) & (!g1464) & (!g325) & (g318)) + ((g1461) & (g1462) & (!g1463) & (!g1464) & (g325) & (g318)) + ((g1461) & (g1462) & (!g1463) & (g1464) & (!g325) & (!g318)) + ((g1461) & (g1462) & (!g1463) & (g1464) & (!g325) & (g318)) + ((g1461) & (g1462) & (g1463) & (!g1464) & (!g325) & (!g318)) + ((g1461) & (g1462) & (g1463) & (!g1464) & (g325) & (g318)) + ((g1461) & (g1462) & (g1463) & (g1464) & (!g325) & (!g318)));
	assign g1467 = (((!sk[48]) & (!g1129) & (g1466)) + ((!sk[48]) & (g1129) & (g1466)) + ((sk[48]) & (!g1129) & (g1466)) + ((sk[48]) & (g1129) & (!g1466)));
	assign g1468 = (((!g617) & (!g873) & (!g1465) & (sk[49]) & (g1467)) + ((!g617) & (!g873) & (g1465) & (!sk[49]) & (!g1467)) + ((!g617) & (!g873) & (g1465) & (!sk[49]) & (g1467)) + ((!g617) & (!g873) & (g1465) & (sk[49]) & (!g1467)) + ((!g617) & (g873) & (!g1465) & (!sk[49]) & (!g1467)) + ((!g617) & (g873) & (!g1465) & (!sk[49]) & (g1467)) + ((!g617) & (g873) & (!g1465) & (sk[49]) & (!g1467)) + ((!g617) & (g873) & (g1465) & (!sk[49]) & (!g1467)) + ((!g617) & (g873) & (g1465) & (!sk[49]) & (g1467)) + ((!g617) & (g873) & (g1465) & (sk[49]) & (g1467)) + ((g617) & (!g873) & (!g1465) & (sk[49]) & (!g1467)) + ((g617) & (!g873) & (g1465) & (!sk[49]) & (!g1467)) + ((g617) & (!g873) & (g1465) & (!sk[49]) & (g1467)) + ((g617) & (!g873) & (g1465) & (sk[49]) & (g1467)) + ((g617) & (g873) & (!g1465) & (!sk[49]) & (!g1467)) + ((g617) & (g873) & (!g1465) & (!sk[49]) & (g1467)) + ((g617) & (g873) & (!g1465) & (sk[49]) & (g1467)) + ((g617) & (g873) & (g1465) & (!sk[49]) & (!g1467)) + ((g617) & (g873) & (g1465) & (!sk[49]) & (g1467)) + ((g617) & (g873) & (g1465) & (sk[49]) & (!g1467)));
	assign g1469 = (((!sk[50]) & (!ld) & (!g361) & (g1468) & (!keyx27x)) + ((!sk[50]) & (!ld) & (!g361) & (g1468) & (keyx27x)) + ((!sk[50]) & (!ld) & (g361) & (!g1468) & (!keyx27x)) + ((!sk[50]) & (!ld) & (g361) & (!g1468) & (keyx27x)) + ((!sk[50]) & (!ld) & (g361) & (g1468) & (!keyx27x)) + ((!sk[50]) & (!ld) & (g361) & (g1468) & (keyx27x)) + ((!sk[50]) & (ld) & (!g361) & (g1468) & (!keyx27x)) + ((!sk[50]) & (ld) & (!g361) & (g1468) & (keyx27x)) + ((!sk[50]) & (ld) & (g361) & (!g1468) & (!keyx27x)) + ((!sk[50]) & (ld) & (g361) & (!g1468) & (keyx27x)) + ((!sk[50]) & (ld) & (g361) & (g1468) & (!keyx27x)) + ((!sk[50]) & (ld) & (g361) & (g1468) & (keyx27x)) + ((sk[50]) & (!ld) & (!g361) & (g1468) & (!keyx27x)) + ((sk[50]) & (!ld) & (!g361) & (g1468) & (keyx27x)) + ((sk[50]) & (!ld) & (g361) & (!g1468) & (!keyx27x)) + ((sk[50]) & (!ld) & (g361) & (!g1468) & (keyx27x)) + ((sk[50]) & (ld) & (!g361) & (!g1468) & (keyx27x)) + ((sk[50]) & (ld) & (!g361) & (g1468) & (keyx27x)) + ((sk[50]) & (ld) & (g361) & (!g1468) & (keyx27x)) + ((sk[50]) & (ld) & (g361) & (g1468) & (keyx27x)));
	assign g1470 = (((!g276) & (!g283) & (!g318) & (!g325) & (!g304) & (g311)) + ((!g276) & (!g283) & (g318) & (!g325) & (!g304) & (g311)) + ((!g276) & (!g283) & (g318) & (!g325) & (g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (!g325) & (g304) & (g311)) + ((!g276) & (!g283) & (g318) & (g325) & (!g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (g325) & (g304) & (!g311)) + ((!g276) & (g283) & (!g318) & (!g325) & (!g304) & (!g311)) + ((!g276) & (g283) & (!g318) & (!g325) & (!g304) & (g311)) + ((!g276) & (g283) & (!g318) & (g325) & (!g304) & (!g311)) + ((!g276) & (g283) & (!g318) & (g325) & (!g304) & (g311)) + ((!g276) & (g283) & (!g318) & (g325) & (g304) & (g311)) + ((!g276) & (g283) & (g318) & (g325) & (!g304) & (g311)) + ((!g276) & (g283) & (g318) & (g325) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g325) & (!g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g325) & (!g304) & (g311)) + ((g276) & (!g283) & (!g318) & (g325) & (!g304) & (g311)) + ((g276) & (!g283) & (g318) & (!g325) & (g304) & (!g311)) + ((g276) & (!g283) & (g318) & (g325) & (!g304) & (!g311)) + ((g276) & (!g283) & (g318) & (g325) & (!g304) & (g311)) + ((g276) & (!g283) & (g318) & (g325) & (g304) & (!g311)) + ((g276) & (g283) & (!g318) & (!g325) & (!g304) & (!g311)) + ((g276) & (g283) & (!g318) & (!g325) & (g304) & (!g311)) + ((g276) & (g283) & (!g318) & (g325) & (g304) & (!g311)) + ((g276) & (g283) & (g318) & (!g325) & (!g304) & (!g311)) + ((g276) & (g283) & (g318) & (!g325) & (!g304) & (g311)) + ((g276) & (g283) & (g318) & (g325) & (!g304) & (g311)));
	assign g1471 = (((!g276) & (!g283) & (!g318) & (!g325) & (!g304) & (!g311)) + ((!g276) & (!g283) & (!g318) & (!g325) & (!g304) & (g311)) + ((!g276) & (!g283) & (!g318) & (!g325) & (g304) & (!g311)) + ((!g276) & (!g283) & (!g318) & (!g325) & (g304) & (g311)) + ((!g276) & (!g283) & (!g318) & (g325) & (!g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (!g325) & (!g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (!g325) & (g304) & (g311)) + ((!g276) & (!g283) & (g318) & (g325) & (!g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (g325) & (g304) & (g311)) + ((!g276) & (g283) & (!g318) & (!g325) & (!g304) & (g311)) + ((!g276) & (g283) & (!g318) & (g325) & (g304) & (!g311)) + ((!g276) & (g283) & (g318) & (!g325) & (!g304) & (!g311)) + ((!g276) & (g283) & (g318) & (!g325) & (!g304) & (g311)) + ((!g276) & (g283) & (g318) & (!g325) & (g304) & (!g311)) + ((!g276) & (g283) & (g318) & (!g325) & (g304) & (g311)) + ((!g276) & (g283) & (g318) & (g325) & (!g304) & (!g311)) + ((!g276) & (g283) & (g318) & (g325) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g325) & (!g304) & (g311)) + ((g276) & (!g283) & (!g318) & (!g325) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g325) & (g304) & (g311)) + ((g276) & (!g283) & (!g318) & (g325) & (!g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (g325) & (g304) & (g311)) + ((g276) & (!g283) & (g318) & (!g325) & (g304) & (!g311)) + ((g276) & (!g283) & (g318) & (!g325) & (g304) & (g311)) + ((g276) & (!g283) & (g318) & (g325) & (!g304) & (g311)) + ((g276) & (g283) & (!g318) & (!g325) & (g304) & (!g311)) + ((g276) & (g283) & (!g318) & (!g325) & (g304) & (g311)) + ((g276) & (g283) & (!g318) & (g325) & (!g304) & (!g311)) + ((g276) & (g283) & (!g318) & (g325) & (!g304) & (g311)) + ((g276) & (g283) & (g318) & (!g325) & (g304) & (!g311)) + ((g276) & (g283) & (g318) & (!g325) & (g304) & (g311)) + ((g276) & (g283) & (g318) & (g325) & (!g304) & (g311)));
	assign g1472 = (((!g276) & (!g283) & (!g318) & (!g325) & (!g304) & (!g311)) + ((!g276) & (!g283) & (!g318) & (!g325) & (!g304) & (g311)) + ((!g276) & (!g283) & (g318) & (!g325) & (!g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (!g325) & (g304) & (g311)) + ((!g276) & (!g283) & (g318) & (g325) & (!g304) & (g311)) + ((!g276) & (g283) & (!g318) & (g325) & (!g304) & (!g311)) + ((!g276) & (g283) & (!g318) & (g325) & (g304) & (!g311)) + ((!g276) & (g283) & (!g318) & (g325) & (g304) & (g311)) + ((!g276) & (g283) & (g318) & (!g325) & (!g304) & (!g311)) + ((!g276) & (g283) & (g318) & (!g325) & (g304) & (!g311)) + ((!g276) & (g283) & (g318) & (!g325) & (g304) & (g311)) + ((!g276) & (g283) & (g318) & (g325) & (!g304) & (!g311)) + ((!g276) & (g283) & (g318) & (g325) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g325) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g325) & (g304) & (g311)) + ((g276) & (!g283) & (!g318) & (g325) & (!g304) & (g311)) + ((g276) & (!g283) & (!g318) & (g325) & (g304) & (g311)) + ((g276) & (!g283) & (g318) & (!g325) & (!g304) & (!g311)) + ((g276) & (!g283) & (g318) & (!g325) & (!g304) & (g311)) + ((g276) & (!g283) & (g318) & (!g325) & (g304) & (g311)) + ((g276) & (!g283) & (g318) & (g325) & (!g304) & (!g311)) + ((g276) & (!g283) & (g318) & (g325) & (!g304) & (g311)) + ((g276) & (!g283) & (g318) & (g325) & (g304) & (!g311)) + ((g276) & (!g283) & (g318) & (g325) & (g304) & (g311)) + ((g276) & (g283) & (!g318) & (!g325) & (!g304) & (g311)) + ((g276) & (g283) & (!g318) & (g325) & (!g304) & (!g311)) + ((g276) & (g283) & (!g318) & (g325) & (g304) & (!g311)) + ((g276) & (g283) & (g318) & (!g325) & (!g304) & (!g311)) + ((g276) & (g283) & (g318) & (!g325) & (!g304) & (g311)) + ((g276) & (g283) & (g318) & (!g325) & (g304) & (!g311)) + ((g276) & (g283) & (g318) & (g325) & (!g304) & (!g311)) + ((g276) & (g283) & (g318) & (g325) & (g304) & (!g311)));
	assign g1473 = (((!g276) & (!g283) & (!g318) & (!g325) & (g304) & (g311)) + ((!g276) & (!g283) & (!g318) & (g325) & (!g304) & (!g311)) + ((!g276) & (!g283) & (!g318) & (g325) & (g304) & (g311)) + ((!g276) & (!g283) & (g318) & (!g325) & (!g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (!g325) & (g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (g325) & (!g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (g325) & (!g304) & (g311)) + ((!g276) & (!g283) & (g318) & (g325) & (g304) & (!g311)) + ((!g276) & (g283) & (!g318) & (!g325) & (!g304) & (!g311)) + ((!g276) & (g283) & (!g318) & (g325) & (!g304) & (g311)) + ((!g276) & (g283) & (!g318) & (g325) & (g304) & (!g311)) + ((!g276) & (g283) & (!g318) & (g325) & (g304) & (g311)) + ((!g276) & (g283) & (g318) & (!g325) & (!g304) & (!g311)) + ((!g276) & (g283) & (g318) & (g325) & (!g304) & (!g311)) + ((!g276) & (g283) & (g318) & (g325) & (!g304) & (g311)) + ((g276) & (!g283) & (!g318) & (!g325) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g325) & (g304) & (g311)) + ((g276) & (!g283) & (g318) & (!g325) & (!g304) & (!g311)) + ((g276) & (!g283) & (g318) & (!g325) & (g304) & (!g311)) + ((g276) & (!g283) & (g318) & (g325) & (g304) & (!g311)) + ((g276) & (g283) & (!g318) & (!g325) & (g304) & (!g311)) + ((g276) & (g283) & (!g318) & (g325) & (g304) & (g311)) + ((g276) & (g283) & (g318) & (!g325) & (!g304) & (!g311)) + ((g276) & (g283) & (g318) & (!g325) & (!g304) & (g311)) + ((g276) & (g283) & (g318) & (!g325) & (g304) & (!g311)) + ((g276) & (g283) & (g318) & (g325) & (!g304) & (!g311)));
	assign g1474 = (((!g1470) & (!g1471) & (!g1472) & (!g1473) & (g290) & (g297)) + ((!g1470) & (!g1471) & (g1472) & (!g1473) & (!g290) & (g297)) + ((!g1470) & (!g1471) & (g1472) & (!g1473) & (g290) & (g297)) + ((!g1470) & (!g1471) & (g1472) & (g1473) & (!g290) & (g297)) + ((!g1470) & (g1471) & (!g1472) & (!g1473) & (g290) & (!g297)) + ((!g1470) & (g1471) & (!g1472) & (!g1473) & (g290) & (g297)) + ((!g1470) & (g1471) & (!g1472) & (g1473) & (g290) & (!g297)) + ((!g1470) & (g1471) & (g1472) & (!g1473) & (!g290) & (g297)) + ((!g1470) & (g1471) & (g1472) & (!g1473) & (g290) & (!g297)) + ((!g1470) & (g1471) & (g1472) & (!g1473) & (g290) & (g297)) + ((!g1470) & (g1471) & (g1472) & (g1473) & (!g290) & (g297)) + ((!g1470) & (g1471) & (g1472) & (g1473) & (g290) & (!g297)) + ((g1470) & (!g1471) & (!g1472) & (!g1473) & (!g290) & (!g297)) + ((g1470) & (!g1471) & (!g1472) & (!g1473) & (g290) & (g297)) + ((g1470) & (!g1471) & (!g1472) & (g1473) & (!g290) & (!g297)) + ((g1470) & (!g1471) & (g1472) & (!g1473) & (!g290) & (!g297)) + ((g1470) & (!g1471) & (g1472) & (!g1473) & (!g290) & (g297)) + ((g1470) & (!g1471) & (g1472) & (!g1473) & (g290) & (g297)) + ((g1470) & (!g1471) & (g1472) & (g1473) & (!g290) & (!g297)) + ((g1470) & (!g1471) & (g1472) & (g1473) & (!g290) & (g297)) + ((g1470) & (g1471) & (!g1472) & (!g1473) & (!g290) & (!g297)) + ((g1470) & (g1471) & (!g1472) & (!g1473) & (g290) & (!g297)) + ((g1470) & (g1471) & (!g1472) & (!g1473) & (g290) & (g297)) + ((g1470) & (g1471) & (!g1472) & (g1473) & (!g290) & (!g297)) + ((g1470) & (g1471) & (!g1472) & (g1473) & (g290) & (!g297)) + ((g1470) & (g1471) & (g1472) & (!g1473) & (!g290) & (!g297)) + ((g1470) & (g1471) & (g1472) & (!g1473) & (!g290) & (g297)) + ((g1470) & (g1471) & (g1472) & (!g1473) & (g290) & (!g297)) + ((g1470) & (g1471) & (g1472) & (!g1473) & (g290) & (g297)) + ((g1470) & (g1471) & (g1472) & (g1473) & (!g290) & (!g297)) + ((g1470) & (g1471) & (g1472) & (g1473) & (!g290) & (g297)) + ((g1470) & (g1471) & (g1472) & (g1473) & (g290) & (!g297)));
	assign g1476 = (((!sk[56]) & (!g1136) & (g1475)) + ((!sk[56]) & (g1136) & (g1475)) + ((sk[56]) & (!g1136) & (g1475)) + ((sk[56]) & (g1136) & (!g1475)));
	assign g1477 = (((!g624) & (!g880) & (!sk[57]) & (g1474) & (!g1476)) + ((!g624) & (!g880) & (!sk[57]) & (g1474) & (g1476)) + ((!g624) & (!g880) & (sk[57]) & (!g1474) & (g1476)) + ((!g624) & (!g880) & (sk[57]) & (g1474) & (!g1476)) + ((!g624) & (g880) & (!sk[57]) & (!g1474) & (!g1476)) + ((!g624) & (g880) & (!sk[57]) & (!g1474) & (g1476)) + ((!g624) & (g880) & (!sk[57]) & (g1474) & (!g1476)) + ((!g624) & (g880) & (!sk[57]) & (g1474) & (g1476)) + ((!g624) & (g880) & (sk[57]) & (!g1474) & (!g1476)) + ((!g624) & (g880) & (sk[57]) & (g1474) & (g1476)) + ((g624) & (!g880) & (!sk[57]) & (g1474) & (!g1476)) + ((g624) & (!g880) & (!sk[57]) & (g1474) & (g1476)) + ((g624) & (!g880) & (sk[57]) & (!g1474) & (!g1476)) + ((g624) & (!g880) & (sk[57]) & (g1474) & (g1476)) + ((g624) & (g880) & (!sk[57]) & (!g1474) & (!g1476)) + ((g624) & (g880) & (!sk[57]) & (!g1474) & (g1476)) + ((g624) & (g880) & (!sk[57]) & (g1474) & (!g1476)) + ((g624) & (g880) & (!sk[57]) & (g1474) & (g1476)) + ((g624) & (g880) & (sk[57]) & (!g1474) & (g1476)) + ((g624) & (g880) & (sk[57]) & (g1474) & (!g1476)));
	assign g1478 = (((!ld) & (!g368) & (!sk[58]) & (g1477) & (!keyx28x)) + ((!ld) & (!g368) & (!sk[58]) & (g1477) & (keyx28x)) + ((!ld) & (!g368) & (sk[58]) & (g1477) & (!keyx28x)) + ((!ld) & (!g368) & (sk[58]) & (g1477) & (keyx28x)) + ((!ld) & (g368) & (!sk[58]) & (!g1477) & (!keyx28x)) + ((!ld) & (g368) & (!sk[58]) & (!g1477) & (keyx28x)) + ((!ld) & (g368) & (!sk[58]) & (g1477) & (!keyx28x)) + ((!ld) & (g368) & (!sk[58]) & (g1477) & (keyx28x)) + ((!ld) & (g368) & (sk[58]) & (!g1477) & (!keyx28x)) + ((!ld) & (g368) & (sk[58]) & (!g1477) & (keyx28x)) + ((ld) & (!g368) & (!sk[58]) & (g1477) & (!keyx28x)) + ((ld) & (!g368) & (!sk[58]) & (g1477) & (keyx28x)) + ((ld) & (!g368) & (sk[58]) & (!g1477) & (keyx28x)) + ((ld) & (!g368) & (sk[58]) & (g1477) & (keyx28x)) + ((ld) & (g368) & (!sk[58]) & (!g1477) & (!keyx28x)) + ((ld) & (g368) & (!sk[58]) & (!g1477) & (keyx28x)) + ((ld) & (g368) & (!sk[58]) & (g1477) & (!keyx28x)) + ((ld) & (g368) & (!sk[58]) & (g1477) & (keyx28x)) + ((ld) & (g368) & (sk[58]) & (!g1477) & (keyx28x)) + ((ld) & (g368) & (sk[58]) & (g1477) & (keyx28x)));
	assign g1479 = (((!g276) & (!g283) & (!g318) & (!g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (!g318) & (!g297) & (g304) & (g311)) + ((!g276) & (!g283) & (!g318) & (g297) & (g304) & (g311)) + ((!g276) & (!g283) & (g318) & (!g297) & (!g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (!g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (g318) & (!g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (!g297) & (g304) & (g311)) + ((!g276) & (!g283) & (g318) & (g297) & (!g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (g297) & (!g304) & (g311)) + ((!g276) & (g283) & (!g318) & (!g297) & (!g304) & (g311)) + ((!g276) & (g283) & (!g318) & (!g297) & (g304) & (!g311)) + ((!g276) & (g283) & (!g318) & (g297) & (g304) & (g311)) + ((!g276) & (g283) & (g318) & (!g297) & (g304) & (!g311)) + ((!g276) & (g283) & (g318) & (!g297) & (g304) & (g311)) + ((!g276) & (g283) & (g318) & (g297) & (!g304) & (!g311)) + ((!g276) & (g283) & (g318) & (g297) & (!g304) & (g311)) + ((!g276) & (g283) & (g318) & (g297) & (g304) & (g311)) + ((g276) & (!g283) & (!g318) & (!g297) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g297) & (g304) & (g311)) + ((g276) & (!g283) & (!g318) & (g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (g297) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (g297) & (g304) & (g311)) + ((g276) & (!g283) & (g318) & (!g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (g318) & (!g297) & (g304) & (!g311)) + ((g276) & (!g283) & (g318) & (g297) & (g304) & (!g311)) + ((g276) & (g283) & (!g318) & (!g297) & (g304) & (g311)) + ((g276) & (g283) & (g318) & (!g297) & (!g304) & (!g311)) + ((g276) & (g283) & (g318) & (!g297) & (g304) & (g311)));
	assign g1480 = (((!g276) & (!g283) & (!g318) & (!g297) & (!g304) & (!g311)) + ((!g276) & (!g283) & (!g318) & (g297) & (!g304) & (!g311)) + ((!g276) & (!g283) & (!g318) & (g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (!g318) & (g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (!g297) & (g304) & (g311)) + ((!g276) & (!g283) & (g318) & (g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (g318) & (g297) & (g304) & (g311)) + ((!g276) & (g283) & (!g318) & (!g297) & (!g304) & (!g311)) + ((!g276) & (g283) & (!g318) & (!g297) & (g304) & (!g311)) + ((!g276) & (g283) & (g318) & (!g297) & (!g304) & (g311)) + ((!g276) & (g283) & (g318) & (!g297) & (g304) & (g311)) + ((!g276) & (g283) & (g318) & (g297) & (!g304) & (g311)) + ((!g276) & (g283) & (g318) & (g297) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g297) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g297) & (g304) & (g311)) + ((g276) & (!g283) & (!g318) & (g297) & (!g304) & (g311)) + ((g276) & (!g283) & (!g318) & (g297) & (g304) & (g311)) + ((g276) & (!g283) & (g318) & (g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (g318) & (g297) & (!g304) & (g311)) + ((g276) & (!g283) & (g318) & (g297) & (g304) & (g311)) + ((g276) & (g283) & (!g318) & (!g297) & (!g304) & (g311)) + ((g276) & (g283) & (!g318) & (!g297) & (g304) & (!g311)) + ((g276) & (g283) & (!g318) & (g297) & (g304) & (!g311)) + ((g276) & (g283) & (g318) & (!g297) & (!g304) & (g311)) + ((g276) & (g283) & (g318) & (!g297) & (g304) & (g311)) + ((g276) & (g283) & (g318) & (g297) & (!g304) & (!g311)) + ((g276) & (g283) & (g318) & (g297) & (g304) & (g311)));
	assign g1481 = (((!g276) & (!g283) & (!g318) & (!g297) & (g304) & (g311)) + ((!g276) & (!g283) & (!g318) & (g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (!g297) & (!g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (!g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (g318) & (!g297) & (g304) & (g311)) + ((!g276) & (!g283) & (g318) & (g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (g318) & (g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (g318) & (g297) & (g304) & (g311)) + ((!g276) & (g283) & (!g318) & (!g297) & (g304) & (!g311)) + ((!g276) & (g283) & (!g318) & (!g297) & (g304) & (g311)) + ((!g276) & (g283) & (g318) & (!g297) & (!g304) & (!g311)) + ((!g276) & (g283) & (g318) & (g297) & (!g304) & (g311)) + ((!g276) & (g283) & (g318) & (g297) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g297) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (!g297) & (g304) & (g311)) + ((g276) & (!g283) & (!g318) & (g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (g297) & (!g304) & (g311)) + ((g276) & (!g283) & (g318) & (!g297) & (!g304) & (g311)) + ((g276) & (!g283) & (g318) & (!g297) & (g304) & (g311)) + ((g276) & (!g283) & (g318) & (g297) & (g304) & (!g311)) + ((g276) & (g283) & (!g318) & (!g297) & (!g304) & (!g311)) + ((g276) & (g283) & (!g318) & (!g297) & (!g304) & (g311)) + ((g276) & (g283) & (!g318) & (!g297) & (g304) & (g311)) + ((g276) & (g283) & (!g318) & (g297) & (!g304) & (g311)) + ((g276) & (g283) & (!g318) & (g297) & (g304) & (!g311)) + ((g276) & (g283) & (g318) & (!g297) & (!g304) & (g311)) + ((g276) & (g283) & (g318) & (!g297) & (g304) & (!g311)) + ((g276) & (g283) & (g318) & (g297) & (!g304) & (!g311)) + ((g276) & (g283) & (g318) & (g297) & (g304) & (!g311)) + ((g276) & (g283) & (g318) & (g297) & (g304) & (g311)));
	assign g1482 = (((!g276) & (!g283) & (!g318) & (!g297) & (g304) & (!g311)) + ((!g276) & (!g283) & (!g318) & (g297) & (!g304) & (!g311)) + ((!g276) & (!g283) & (!g318) & (g297) & (g304) & (g311)) + ((!g276) & (!g283) & (g318) & (!g297) & (!g304) & (g311)) + ((!g276) & (!g283) & (g318) & (!g297) & (g304) & (g311)) + ((!g276) & (!g283) & (g318) & (g297) & (g304) & (g311)) + ((!g276) & (g283) & (!g318) & (!g297) & (!g304) & (g311)) + ((!g276) & (g283) & (!g318) & (g297) & (!g304) & (g311)) + ((!g276) & (g283) & (!g318) & (g297) & (g304) & (g311)) + ((!g276) & (g283) & (g318) & (!g297) & (!g304) & (!g311)) + ((!g276) & (g283) & (g318) & (!g297) & (g304) & (!g311)) + ((!g276) & (g283) & (g318) & (g297) & (!g304) & (g311)) + ((!g276) & (g283) & (g318) & (g297) & (g304) & (g311)) + ((g276) & (!g283) & (!g318) & (!g297) & (g304) & (!g311)) + ((g276) & (!g283) & (!g318) & (g297) & (g304) & (g311)) + ((g276) & (!g283) & (g318) & (!g297) & (!g304) & (!g311)) + ((g276) & (!g283) & (g318) & (!g297) & (g304) & (g311)) + ((g276) & (!g283) & (g318) & (g297) & (!g304) & (!g311)) + ((g276) & (g283) & (!g318) & (!g297) & (g304) & (g311)) + ((g276) & (g283) & (!g318) & (g297) & (!g304) & (!g311)) + ((g276) & (g283) & (!g318) & (g297) & (!g304) & (g311)) + ((g276) & (g283) & (g318) & (!g297) & (g304) & (g311)));
	assign g1483 = (((!g1479) & (!g1480) & (!g1481) & (!g1482) & (!g325) & (!g290)) + ((!g1479) & (!g1480) & (!g1481) & (!g1482) & (!g325) & (g290)) + ((!g1479) & (!g1480) & (!g1481) & (!g1482) & (g325) & (!g290)) + ((!g1479) & (!g1480) & (!g1481) & (g1482) & (!g325) & (!g290)) + ((!g1479) & (!g1480) & (!g1481) & (g1482) & (!g325) & (g290)) + ((!g1479) & (!g1480) & (!g1481) & (g1482) & (g325) & (!g290)) + ((!g1479) & (!g1480) & (!g1481) & (g1482) & (g325) & (g290)) + ((!g1479) & (!g1480) & (g1481) & (!g1482) & (!g325) & (!g290)) + ((!g1479) & (!g1480) & (g1481) & (!g1482) & (g325) & (!g290)) + ((!g1479) & (!g1480) & (g1481) & (g1482) & (!g325) & (!g290)) + ((!g1479) & (!g1480) & (g1481) & (g1482) & (g325) & (!g290)) + ((!g1479) & (!g1480) & (g1481) & (g1482) & (g325) & (g290)) + ((!g1479) & (g1480) & (!g1481) & (!g1482) & (!g325) & (!g290)) + ((!g1479) & (g1480) & (!g1481) & (!g1482) & (!g325) & (g290)) + ((!g1479) & (g1480) & (!g1481) & (g1482) & (!g325) & (!g290)) + ((!g1479) & (g1480) & (!g1481) & (g1482) & (!g325) & (g290)) + ((!g1479) & (g1480) & (!g1481) & (g1482) & (g325) & (g290)) + ((!g1479) & (g1480) & (g1481) & (!g1482) & (!g325) & (!g290)) + ((!g1479) & (g1480) & (g1481) & (g1482) & (!g325) & (!g290)) + ((!g1479) & (g1480) & (g1481) & (g1482) & (g325) & (g290)) + ((g1479) & (!g1480) & (!g1481) & (!g1482) & (!g325) & (g290)) + ((g1479) & (!g1480) & (!g1481) & (!g1482) & (g325) & (!g290)) + ((g1479) & (!g1480) & (!g1481) & (g1482) & (!g325) & (g290)) + ((g1479) & (!g1480) & (!g1481) & (g1482) & (g325) & (!g290)) + ((g1479) & (!g1480) & (!g1481) & (g1482) & (g325) & (g290)) + ((g1479) & (!g1480) & (g1481) & (!g1482) & (g325) & (!g290)) + ((g1479) & (!g1480) & (g1481) & (g1482) & (g325) & (!g290)) + ((g1479) & (!g1480) & (g1481) & (g1482) & (g325) & (g290)) + ((g1479) & (g1480) & (!g1481) & (!g1482) & (!g325) & (g290)) + ((g1479) & (g1480) & (!g1481) & (g1482) & (!g325) & (g290)) + ((g1479) & (g1480) & (!g1481) & (g1482) & (g325) & (g290)) + ((g1479) & (g1480) & (g1481) & (g1482) & (g325) & (g290)));
	assign g1485 = (((!sk[64]) & (!g1143) & (g1484)) + ((!sk[64]) & (g1143) & (g1484)) + ((sk[64]) & (!g1143) & (g1484)) + ((sk[64]) & (g1143) & (!g1484)));
	assign g1486 = (((!g631) & (!g887) & (!g1483) & (sk[65]) & (g1485)) + ((!g631) & (!g887) & (g1483) & (!sk[65]) & (!g1485)) + ((!g631) & (!g887) & (g1483) & (!sk[65]) & (g1485)) + ((!g631) & (!g887) & (g1483) & (sk[65]) & (!g1485)) + ((!g631) & (g887) & (!g1483) & (!sk[65]) & (!g1485)) + ((!g631) & (g887) & (!g1483) & (!sk[65]) & (g1485)) + ((!g631) & (g887) & (!g1483) & (sk[65]) & (!g1485)) + ((!g631) & (g887) & (g1483) & (!sk[65]) & (!g1485)) + ((!g631) & (g887) & (g1483) & (!sk[65]) & (g1485)) + ((!g631) & (g887) & (g1483) & (sk[65]) & (g1485)) + ((g631) & (!g887) & (!g1483) & (sk[65]) & (!g1485)) + ((g631) & (!g887) & (g1483) & (!sk[65]) & (!g1485)) + ((g631) & (!g887) & (g1483) & (!sk[65]) & (g1485)) + ((g631) & (!g887) & (g1483) & (sk[65]) & (g1485)) + ((g631) & (g887) & (!g1483) & (!sk[65]) & (!g1485)) + ((g631) & (g887) & (!g1483) & (!sk[65]) & (g1485)) + ((g631) & (g887) & (!g1483) & (sk[65]) & (g1485)) + ((g631) & (g887) & (g1483) & (!sk[65]) & (!g1485)) + ((g631) & (g887) & (g1483) & (!sk[65]) & (g1485)) + ((g631) & (g887) & (g1483) & (sk[65]) & (!g1485)));
	assign g1487 = (((!ld) & (!g375) & (g1486) & (!sk[66]) & (!keyx29x)) + ((!ld) & (!g375) & (g1486) & (!sk[66]) & (keyx29x)) + ((!ld) & (!g375) & (g1486) & (sk[66]) & (!keyx29x)) + ((!ld) & (!g375) & (g1486) & (sk[66]) & (keyx29x)) + ((!ld) & (g375) & (!g1486) & (!sk[66]) & (!keyx29x)) + ((!ld) & (g375) & (!g1486) & (!sk[66]) & (keyx29x)) + ((!ld) & (g375) & (!g1486) & (sk[66]) & (!keyx29x)) + ((!ld) & (g375) & (!g1486) & (sk[66]) & (keyx29x)) + ((!ld) & (g375) & (g1486) & (!sk[66]) & (!keyx29x)) + ((!ld) & (g375) & (g1486) & (!sk[66]) & (keyx29x)) + ((ld) & (!g375) & (!g1486) & (sk[66]) & (keyx29x)) + ((ld) & (!g375) & (g1486) & (!sk[66]) & (!keyx29x)) + ((ld) & (!g375) & (g1486) & (!sk[66]) & (keyx29x)) + ((ld) & (!g375) & (g1486) & (sk[66]) & (keyx29x)) + ((ld) & (g375) & (!g1486) & (!sk[66]) & (!keyx29x)) + ((ld) & (g375) & (!g1486) & (!sk[66]) & (keyx29x)) + ((ld) & (g375) & (!g1486) & (sk[66]) & (keyx29x)) + ((ld) & (g375) & (g1486) & (!sk[66]) & (!keyx29x)) + ((ld) & (g375) & (g1486) & (!sk[66]) & (keyx29x)) + ((ld) & (g375) & (g1486) & (sk[66]) & (keyx29x)));
	assign g1488 = (((!g276) & (!g325) & (!g290) & (!g297) & (!g304) & (g311)) + ((!g276) & (!g325) & (!g290) & (!g297) & (g304) & (g311)) + ((!g276) & (!g325) & (!g290) & (g297) & (!g304) & (!g311)) + ((!g276) & (!g325) & (!g290) & (g297) & (!g304) & (g311)) + ((!g276) & (!g325) & (!g290) & (g297) & (g304) & (!g311)) + ((!g276) & (!g325) & (!g290) & (g297) & (g304) & (g311)) + ((!g276) & (!g325) & (g290) & (!g297) & (!g304) & (g311)) + ((!g276) & (!g325) & (g290) & (!g297) & (g304) & (g311)) + ((!g276) & (!g325) & (g290) & (g297) & (g304) & (!g311)) + ((!g276) & (g325) & (g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (g325) & (g290) & (!g297) & (g304) & (g311)) + ((!g276) & (g325) & (g290) & (g297) & (!g304) & (g311)) + ((g276) & (!g325) & (!g290) & (!g297) & (g304) & (!g311)) + ((g276) & (!g325) & (!g290) & (g297) & (!g304) & (!g311)) + ((g276) & (!g325) & (!g290) & (g297) & (!g304) & (g311)) + ((g276) & (!g325) & (!g290) & (g297) & (g304) & (g311)) + ((g276) & (!g325) & (g290) & (!g297) & (!g304) & (g311)) + ((g276) & (!g325) & (g290) & (!g297) & (g304) & (g311)) + ((g276) & (!g325) & (g290) & (g297) & (g304) & (!g311)) + ((g276) & (!g325) & (g290) & (g297) & (g304) & (g311)) + ((g276) & (g325) & (!g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (g325) & (!g290) & (!g297) & (!g304) & (g311)) + ((g276) & (g325) & (!g290) & (!g297) & (g304) & (!g311)) + ((g276) & (g325) & (!g290) & (g297) & (!g304) & (!g311)) + ((g276) & (g325) & (g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (g325) & (g290) & (!g297) & (!g304) & (g311)) + ((g276) & (g325) & (g290) & (!g297) & (g304) & (!g311)) + ((g276) & (g325) & (g290) & (g297) & (!g304) & (g311)));
	assign g1489 = (((!g276) & (!g325) & (!g290) & (!g297) & (!g304) & (!g311)) + ((!g276) & (!g325) & (!g290) & (g297) & (g304) & (g311)) + ((!g276) & (!g325) & (g290) & (!g297) & (!g304) & (!g311)) + ((!g276) & (!g325) & (g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (!g325) & (g290) & (!g297) & (g304) & (g311)) + ((!g276) & (!g325) & (g290) & (g297) & (!g304) & (!g311)) + ((!g276) & (!g325) & (g290) & (g297) & (g304) & (g311)) + ((!g276) & (g325) & (!g290) & (!g297) & (!g304) & (!g311)) + ((!g276) & (g325) & (!g290) & (!g297) & (g304) & (g311)) + ((!g276) & (g325) & (!g290) & (g297) & (!g304) & (g311)) + ((!g276) & (g325) & (g290) & (!g297) & (!g304) & (!g311)) + ((!g276) & (g325) & (g290) & (!g297) & (g304) & (g311)) + ((!g276) & (g325) & (g290) & (g297) & (g304) & (!g311)) + ((!g276) & (g325) & (g290) & (g297) & (g304) & (g311)) + ((g276) & (!g325) & (!g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (!g325) & (!g290) & (!g297) & (g304) & (g311)) + ((g276) & (!g325) & (!g290) & (g297) & (!g304) & (!g311)) + ((g276) & (!g325) & (!g290) & (g297) & (g304) & (g311)) + ((g276) & (!g325) & (g290) & (!g297) & (g304) & (g311)) + ((g276) & (!g325) & (g290) & (g297) & (!g304) & (g311)) + ((g276) & (g325) & (!g290) & (!g297) & (g304) & (!g311)) + ((g276) & (g325) & (!g290) & (!g297) & (g304) & (g311)) + ((g276) & (g325) & (!g290) & (g297) & (!g304) & (g311)) + ((g276) & (g325) & (!g290) & (g297) & (g304) & (!g311)) + ((g276) & (g325) & (!g290) & (g297) & (g304) & (g311)) + ((g276) & (g325) & (g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (g325) & (g290) & (!g297) & (g304) & (!g311)) + ((g276) & (g325) & (g290) & (g297) & (!g304) & (!g311)));
	assign g1490 = (((!g276) & (!g325) & (!g290) & (!g297) & (!g304) & (g311)) + ((!g276) & (!g325) & (!g290) & (!g297) & (g304) & (g311)) + ((!g276) & (!g325) & (!g290) & (g297) & (g304) & (!g311)) + ((!g276) & (!g325) & (!g290) & (g297) & (g304) & (g311)) + ((!g276) & (!g325) & (g290) & (!g297) & (g304) & (g311)) + ((!g276) & (!g325) & (g290) & (g297) & (!g304) & (!g311)) + ((!g276) & (!g325) & (g290) & (g297) & (!g304) & (g311)) + ((!g276) & (!g325) & (g290) & (g297) & (g304) & (g311)) + ((!g276) & (g325) & (!g290) & (!g297) & (!g304) & (!g311)) + ((!g276) & (g325) & (!g290) & (!g297) & (!g304) & (g311)) + ((!g276) & (g325) & (!g290) & (!g297) & (g304) & (g311)) + ((!g276) & (g325) & (!g290) & (g297) & (!g304) & (g311)) + ((!g276) & (g325) & (!g290) & (g297) & (g304) & (!g311)) + ((!g276) & (g325) & (g290) & (!g297) & (!g304) & (g311)) + ((!g276) & (g325) & (g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (g325) & (g290) & (g297) & (!g304) & (!g311)) + ((!g276) & (g325) & (g290) & (g297) & (g304) & (!g311)) + ((!g276) & (g325) & (g290) & (g297) & (g304) & (g311)) + ((g276) & (!g325) & (!g290) & (!g297) & (!g304) & (g311)) + ((g276) & (!g325) & (!g290) & (g297) & (!g304) & (!g311)) + ((g276) & (!g325) & (!g290) & (g297) & (g304) & (!g311)) + ((g276) & (!g325) & (g290) & (!g297) & (g304) & (g311)) + ((g276) & (!g325) & (g290) & (g297) & (!g304) & (g311)) + ((g276) & (g325) & (!g290) & (!g297) & (!g304) & (g311)) + ((g276) & (g325) & (!g290) & (g297) & (!g304) & (!g311)) + ((g276) & (g325) & (!g290) & (g297) & (g304) & (!g311)) + ((g276) & (g325) & (g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (g325) & (g290) & (!g297) & (g304) & (!g311)) + ((g276) & (g325) & (g290) & (!g297) & (g304) & (g311)) + ((g276) & (g325) & (g290) & (g297) & (g304) & (g311)));
	assign g1491 = (((!g276) & (!g325) & (!g290) & (!g297) & (g304) & (g311)) + ((!g276) & (!g325) & (!g290) & (g297) & (!g304) & (!g311)) + ((!g276) & (!g325) & (!g290) & (g297) & (g304) & (g311)) + ((!g276) & (!g325) & (g290) & (!g297) & (!g304) & (!g311)) + ((!g276) & (!g325) & (g290) & (g297) & (g304) & (!g311)) + ((!g276) & (!g325) & (g290) & (g297) & (g304) & (g311)) + ((!g276) & (g325) & (!g290) & (g297) & (!g304) & (!g311)) + ((!g276) & (g325) & (!g290) & (g297) & (g304) & (!g311)) + ((!g276) & (g325) & (g290) & (!g297) & (g304) & (!g311)) + ((!g276) & (g325) & (g290) & (!g297) & (g304) & (g311)) + ((g276) & (!g325) & (!g290) & (!g297) & (!g304) & (g311)) + ((g276) & (!g325) & (!g290) & (!g297) & (g304) & (!g311)) + ((g276) & (!g325) & (!g290) & (g297) & (!g304) & (g311)) + ((g276) & (!g325) & (g290) & (!g297) & (g304) & (!g311)) + ((g276) & (!g325) & (g290) & (!g297) & (g304) & (g311)) + ((g276) & (!g325) & (g290) & (g297) & (g304) & (!g311)) + ((g276) & (!g325) & (g290) & (g297) & (g304) & (g311)) + ((g276) & (g325) & (!g290) & (!g297) & (g304) & (!g311)) + ((g276) & (g325) & (!g290) & (g297) & (!g304) & (g311)) + ((g276) & (g325) & (g290) & (!g297) & (!g304) & (!g311)) + ((g276) & (g325) & (g290) & (!g297) & (g304) & (g311)) + ((g276) & (g325) & (g290) & (g297) & (!g304) & (g311)));
	assign g1492 = (((!g1488) & (!g1489) & (!g1490) & (!g1491) & (!g318) & (!g283)) + ((!g1488) & (!g1489) & (!g1490) & (!g1491) & (!g318) & (g283)) + ((!g1488) & (!g1489) & (!g1490) & (!g1491) & (g318) & (!g283)) + ((!g1488) & (!g1489) & (!g1490) & (g1491) & (!g318) & (!g283)) + ((!g1488) & (!g1489) & (!g1490) & (g1491) & (!g318) & (g283)) + ((!g1488) & (!g1489) & (!g1490) & (g1491) & (g318) & (!g283)) + ((!g1488) & (!g1489) & (!g1490) & (g1491) & (g318) & (g283)) + ((!g1488) & (!g1489) & (g1490) & (!g1491) & (!g318) & (!g283)) + ((!g1488) & (!g1489) & (g1490) & (!g1491) & (g318) & (!g283)) + ((!g1488) & (!g1489) & (g1490) & (g1491) & (!g318) & (!g283)) + ((!g1488) & (!g1489) & (g1490) & (g1491) & (g318) & (!g283)) + ((!g1488) & (!g1489) & (g1490) & (g1491) & (g318) & (g283)) + ((!g1488) & (g1489) & (!g1490) & (!g1491) & (!g318) & (!g283)) + ((!g1488) & (g1489) & (!g1490) & (!g1491) & (!g318) & (g283)) + ((!g1488) & (g1489) & (!g1490) & (g1491) & (!g318) & (!g283)) + ((!g1488) & (g1489) & (!g1490) & (g1491) & (!g318) & (g283)) + ((!g1488) & (g1489) & (!g1490) & (g1491) & (g318) & (g283)) + ((!g1488) & (g1489) & (g1490) & (!g1491) & (!g318) & (!g283)) + ((!g1488) & (g1489) & (g1490) & (g1491) & (!g318) & (!g283)) + ((!g1488) & (g1489) & (g1490) & (g1491) & (g318) & (g283)) + ((g1488) & (!g1489) & (!g1490) & (!g1491) & (!g318) & (g283)) + ((g1488) & (!g1489) & (!g1490) & (!g1491) & (g318) & (!g283)) + ((g1488) & (!g1489) & (!g1490) & (g1491) & (!g318) & (g283)) + ((g1488) & (!g1489) & (!g1490) & (g1491) & (g318) & (!g283)) + ((g1488) & (!g1489) & (!g1490) & (g1491) & (g318) & (g283)) + ((g1488) & (!g1489) & (g1490) & (!g1491) & (g318) & (!g283)) + ((g1488) & (!g1489) & (g1490) & (g1491) & (g318) & (!g283)) + ((g1488) & (!g1489) & (g1490) & (g1491) & (g318) & (g283)) + ((g1488) & (g1489) & (!g1490) & (!g1491) & (!g318) & (g283)) + ((g1488) & (g1489) & (!g1490) & (g1491) & (!g318) & (g283)) + ((g1488) & (g1489) & (!g1490) & (g1491) & (g318) & (g283)) + ((g1488) & (g1489) & (g1490) & (g1491) & (g318) & (g283)));
	assign g1494 = (((!g1150) & (!sk[72]) & (g1493)) + ((!g1150) & (sk[72]) & (g1493)) + ((g1150) & (!sk[72]) & (g1493)) + ((g1150) & (sk[72]) & (!g1493)));
	assign g1495 = (((!g638) & (!g894) & (!g1492) & (sk[73]) & (g1494)) + ((!g638) & (!g894) & (g1492) & (!sk[73]) & (!g1494)) + ((!g638) & (!g894) & (g1492) & (!sk[73]) & (g1494)) + ((!g638) & (!g894) & (g1492) & (sk[73]) & (!g1494)) + ((!g638) & (g894) & (!g1492) & (!sk[73]) & (!g1494)) + ((!g638) & (g894) & (!g1492) & (!sk[73]) & (g1494)) + ((!g638) & (g894) & (!g1492) & (sk[73]) & (!g1494)) + ((!g638) & (g894) & (g1492) & (!sk[73]) & (!g1494)) + ((!g638) & (g894) & (g1492) & (!sk[73]) & (g1494)) + ((!g638) & (g894) & (g1492) & (sk[73]) & (g1494)) + ((g638) & (!g894) & (!g1492) & (sk[73]) & (!g1494)) + ((g638) & (!g894) & (g1492) & (!sk[73]) & (!g1494)) + ((g638) & (!g894) & (g1492) & (!sk[73]) & (g1494)) + ((g638) & (!g894) & (g1492) & (sk[73]) & (g1494)) + ((g638) & (g894) & (!g1492) & (!sk[73]) & (!g1494)) + ((g638) & (g894) & (!g1492) & (!sk[73]) & (g1494)) + ((g638) & (g894) & (!g1492) & (sk[73]) & (g1494)) + ((g638) & (g894) & (g1492) & (!sk[73]) & (!g1494)) + ((g638) & (g894) & (g1492) & (!sk[73]) & (g1494)) + ((g638) & (g894) & (g1492) & (sk[73]) & (!g1494)));
	assign g1496 = (((!ld) & (!sk[74]) & (!g382) & (g1495) & (!keyx30x)) + ((!ld) & (!sk[74]) & (!g382) & (g1495) & (keyx30x)) + ((!ld) & (!sk[74]) & (g382) & (!g1495) & (!keyx30x)) + ((!ld) & (!sk[74]) & (g382) & (!g1495) & (keyx30x)) + ((!ld) & (!sk[74]) & (g382) & (g1495) & (!keyx30x)) + ((!ld) & (!sk[74]) & (g382) & (g1495) & (keyx30x)) + ((!ld) & (sk[74]) & (!g382) & (g1495) & (!keyx30x)) + ((!ld) & (sk[74]) & (!g382) & (g1495) & (keyx30x)) + ((!ld) & (sk[74]) & (g382) & (!g1495) & (!keyx30x)) + ((!ld) & (sk[74]) & (g382) & (!g1495) & (keyx30x)) + ((ld) & (!sk[74]) & (!g382) & (g1495) & (!keyx30x)) + ((ld) & (!sk[74]) & (!g382) & (g1495) & (keyx30x)) + ((ld) & (!sk[74]) & (g382) & (!g1495) & (!keyx30x)) + ((ld) & (!sk[74]) & (g382) & (!g1495) & (keyx30x)) + ((ld) & (!sk[74]) & (g382) & (g1495) & (!keyx30x)) + ((ld) & (!sk[74]) & (g382) & (g1495) & (keyx30x)) + ((ld) & (sk[74]) & (!g382) & (!g1495) & (keyx30x)) + ((ld) & (sk[74]) & (!g382) & (g1495) & (keyx30x)) + ((ld) & (sk[74]) & (g382) & (!g1495) & (keyx30x)) + ((ld) & (sk[74]) & (g382) & (g1495) & (keyx30x)));
	assign g1497 = (((!g318) & (!g283) & (!g290) & (!g297) & (!g304) & (g325)) + ((!g318) & (!g283) & (!g290) & (!g297) & (g304) & (!g325)) + ((!g318) & (!g283) & (!g290) & (g297) & (!g304) & (g325)) + ((!g318) & (!g283) & (!g290) & (g297) & (g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (!g297) & (!g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (!g297) & (g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (g297) & (!g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (g297) & (g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (g297) & (g304) & (g325)) + ((!g318) & (g283) & (!g290) & (!g297) & (g304) & (!g325)) + ((!g318) & (g283) & (!g290) & (g297) & (g304) & (!g325)) + ((!g318) & (g283) & (!g290) & (g297) & (g304) & (g325)) + ((!g318) & (g283) & (g290) & (!g297) & (g304) & (g325)) + ((!g318) & (g283) & (g290) & (g297) & (!g304) & (!g325)) + ((g318) & (!g283) & (!g290) & (!g297) & (!g304) & (g325)) + ((g318) & (!g283) & (!g290) & (g297) & (!g304) & (g325)) + ((g318) & (!g283) & (g290) & (g297) & (g304) & (g325)) + ((g318) & (g283) & (!g290) & (!g297) & (g304) & (g325)) + ((g318) & (g283) & (!g290) & (g297) & (!g304) & (!g325)) + ((g318) & (g283) & (!g290) & (g297) & (g304) & (!g325)) + ((g318) & (g283) & (g290) & (!g297) & (!g304) & (g325)) + ((g318) & (g283) & (g290) & (!g297) & (g304) & (!g325)) + ((g318) & (g283) & (g290) & (!g297) & (g304) & (g325)) + ((g318) & (g283) & (g290) & (g297) & (!g304) & (g325)));
	assign g1498 = (((!g318) & (!g283) & (!g290) & (!g297) & (!g304) & (!g325)) + ((!g318) & (!g283) & (!g290) & (!g297) & (!g304) & (g325)) + ((!g318) & (!g283) & (!g290) & (g297) & (!g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (!g297) & (!g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (!g297) & (g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (!g297) & (g304) & (g325)) + ((!g318) & (!g283) & (g290) & (g297) & (!g304) & (g325)) + ((!g318) & (!g283) & (g290) & (g297) & (g304) & (g325)) + ((!g318) & (g283) & (!g290) & (!g297) & (!g304) & (!g325)) + ((!g318) & (g283) & (!g290) & (!g297) & (g304) & (!g325)) + ((!g318) & (g283) & (!g290) & (g297) & (!g304) & (!g325)) + ((!g318) & (g283) & (!g290) & (g297) & (!g304) & (g325)) + ((!g318) & (g283) & (!g290) & (g297) & (g304) & (g325)) + ((!g318) & (g283) & (g290) & (!g297) & (!g304) & (g325)) + ((!g318) & (g283) & (g290) & (g297) & (!g304) & (!g325)) + ((!g318) & (g283) & (g290) & (g297) & (!g304) & (g325)) + ((g318) & (!g283) & (!g290) & (!g297) & (!g304) & (g325)) + ((g318) & (!g283) & (!g290) & (!g297) & (g304) & (g325)) + ((g318) & (!g283) & (!g290) & (g297) & (!g304) & (!g325)) + ((g318) & (!g283) & (!g290) & (g297) & (g304) & (g325)) + ((g318) & (!g283) & (g290) & (!g297) & (!g304) & (!g325)) + ((g318) & (!g283) & (g290) & (!g297) & (g304) & (g325)) + ((g318) & (!g283) & (g290) & (g297) & (g304) & (!g325)) + ((g318) & (g283) & (!g290) & (!g297) & (!g304) & (!g325)) + ((g318) & (g283) & (!g290) & (!g297) & (!g304) & (g325)) + ((g318) & (g283) & (!g290) & (!g297) & (g304) & (g325)) + ((g318) & (g283) & (!g290) & (g297) & (!g304) & (g325)) + ((g318) & (g283) & (!g290) & (g297) & (g304) & (!g325)) + ((g318) & (g283) & (g290) & (!g297) & (g304) & (!g325)) + ((g318) & (g283) & (g290) & (!g297) & (g304) & (g325)));
	assign g1499 = (((!g318) & (!g283) & (!g290) & (!g297) & (g304) & (!g325)) + ((!g318) & (!g283) & (!g290) & (g297) & (!g304) & (!g325)) + ((!g318) & (!g283) & (!g290) & (g297) & (g304) & (!g325)) + ((!g318) & (!g283) & (!g290) & (g297) & (g304) & (g325)) + ((!g318) & (!g283) & (g290) & (!g297) & (!g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (!g297) & (!g304) & (g325)) + ((!g318) & (!g283) & (g290) & (!g297) & (g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (g297) & (!g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (g297) & (g304) & (g325)) + ((!g318) & (g283) & (!g290) & (!g297) & (!g304) & (g325)) + ((!g318) & (g283) & (!g290) & (!g297) & (g304) & (!g325)) + ((!g318) & (g283) & (!g290) & (!g297) & (g304) & (g325)) + ((!g318) & (g283) & (g290) & (!g297) & (!g304) & (g325)) + ((!g318) & (g283) & (g290) & (!g297) & (g304) & (!g325)) + ((!g318) & (g283) & (g290) & (!g297) & (g304) & (g325)) + ((!g318) & (g283) & (g290) & (g297) & (!g304) & (!g325)) + ((g318) & (!g283) & (!g290) & (!g297) & (g304) & (!g325)) + ((g318) & (!g283) & (!g290) & (g297) & (!g304) & (!g325)) + ((g318) & (!g283) & (!g290) & (g297) & (g304) & (g325)) + ((g318) & (!g283) & (g290) & (!g297) & (!g304) & (!g325)) + ((g318) & (!g283) & (g290) & (!g297) & (!g304) & (g325)) + ((g318) & (!g283) & (g290) & (g297) & (!g304) & (!g325)) + ((g318) & (!g283) & (g290) & (g297) & (g304) & (!g325)) + ((g318) & (g283) & (!g290) & (!g297) & (g304) & (!g325)) + ((g318) & (g283) & (!g290) & (g297) & (!g304) & (!g325)) + ((g318) & (g283) & (!g290) & (g297) & (g304) & (g325)) + ((g318) & (g283) & (g290) & (!g297) & (!g304) & (!g325)) + ((g318) & (g283) & (g290) & (!g297) & (g304) & (!g325)) + ((g318) & (g283) & (g290) & (!g297) & (g304) & (g325)) + ((g318) & (g283) & (g290) & (g297) & (!g304) & (g325)));
	assign g1500 = (((!g318) & (!g283) & (!g290) & (!g297) & (!g304) & (g325)) + ((!g318) & (!g283) & (!g290) & (g297) & (g304) & (!g325)) + ((!g318) & (!g283) & (!g290) & (g297) & (g304) & (g325)) + ((!g318) & (!g283) & (g290) & (!g297) & (!g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (!g297) & (!g304) & (g325)) + ((!g318) & (!g283) & (g290) & (g297) & (g304) & (!g325)) + ((!g318) & (!g283) & (g290) & (g297) & (g304) & (g325)) + ((!g318) & (g283) & (!g290) & (!g297) & (!g304) & (!g325)) + ((!g318) & (g283) & (!g290) & (!g297) & (!g304) & (g325)) + ((!g318) & (g283) & (!g290) & (!g297) & (g304) & (g325)) + ((!g318) & (g283) & (!g290) & (g297) & (!g304) & (g325)) + ((!g318) & (g283) & (g290) & (!g297) & (!g304) & (g325)) + ((!g318) & (g283) & (g290) & (g297) & (!g304) & (!g325)) + ((!g318) & (g283) & (g290) & (g297) & (!g304) & (g325)) + ((!g318) & (g283) & (g290) & (g297) & (g304) & (!g325)) + ((!g318) & (g283) & (g290) & (g297) & (g304) & (g325)) + ((g318) & (!g283) & (!g290) & (g297) & (!g304) & (g325)) + ((g318) & (!g283) & (g290) & (!g297) & (!g304) & (!g325)) + ((g318) & (!g283) & (g290) & (g297) & (!g304) & (!g325)) + ((g318) & (!g283) & (g290) & (g297) & (!g304) & (g325)) + ((g318) & (!g283) & (g290) & (g297) & (g304) & (g325)) + ((g318) & (g283) & (!g290) & (!g297) & (!g304) & (g325)) + ((g318) & (g283) & (!g290) & (!g297) & (g304) & (g325)) + ((g318) & (g283) & (!g290) & (g297) & (!g304) & (!g325)) + ((g318) & (g283) & (!g290) & (g297) & (g304) & (!g325)) + ((g318) & (g283) & (!g290) & (g297) & (g304) & (g325)) + ((g318) & (g283) & (g290) & (!g297) & (g304) & (g325)) + ((g318) & (g283) & (g290) & (g297) & (g304) & (g325)));
	assign g1501 = (((!g1497) & (!g1498) & (!g1499) & (!g1500) & (!g276) & (g311)) + ((!g1497) & (!g1498) & (!g1499) & (!g1500) & (g276) & (!g311)) + ((!g1497) & (!g1498) & (!g1499) & (!g1500) & (g276) & (g311)) + ((!g1497) & (!g1498) & (!g1499) & (g1500) & (!g276) & (g311)) + ((!g1497) & (!g1498) & (!g1499) & (g1500) & (g276) & (!g311)) + ((!g1497) & (!g1498) & (g1499) & (!g1500) & (g276) & (!g311)) + ((!g1497) & (!g1498) & (g1499) & (!g1500) & (g276) & (g311)) + ((!g1497) & (!g1498) & (g1499) & (g1500) & (g276) & (!g311)) + ((!g1497) & (g1498) & (!g1499) & (!g1500) & (!g276) & (g311)) + ((!g1497) & (g1498) & (!g1499) & (!g1500) & (g276) & (g311)) + ((!g1497) & (g1498) & (!g1499) & (g1500) & (!g276) & (g311)) + ((!g1497) & (g1498) & (g1499) & (!g1500) & (g276) & (g311)) + ((g1497) & (!g1498) & (!g1499) & (!g1500) & (!g276) & (!g311)) + ((g1497) & (!g1498) & (!g1499) & (!g1500) & (!g276) & (g311)) + ((g1497) & (!g1498) & (!g1499) & (!g1500) & (g276) & (!g311)) + ((g1497) & (!g1498) & (!g1499) & (!g1500) & (g276) & (g311)) + ((g1497) & (!g1498) & (!g1499) & (g1500) & (!g276) & (!g311)) + ((g1497) & (!g1498) & (!g1499) & (g1500) & (!g276) & (g311)) + ((g1497) & (!g1498) & (!g1499) & (g1500) & (g276) & (!g311)) + ((g1497) & (!g1498) & (g1499) & (!g1500) & (!g276) & (!g311)) + ((g1497) & (!g1498) & (g1499) & (!g1500) & (g276) & (!g311)) + ((g1497) & (!g1498) & (g1499) & (!g1500) & (g276) & (g311)) + ((g1497) & (!g1498) & (g1499) & (g1500) & (!g276) & (!g311)) + ((g1497) & (!g1498) & (g1499) & (g1500) & (g276) & (!g311)) + ((g1497) & (g1498) & (!g1499) & (!g1500) & (!g276) & (!g311)) + ((g1497) & (g1498) & (!g1499) & (!g1500) & (!g276) & (g311)) + ((g1497) & (g1498) & (!g1499) & (!g1500) & (g276) & (g311)) + ((g1497) & (g1498) & (!g1499) & (g1500) & (!g276) & (!g311)) + ((g1497) & (g1498) & (!g1499) & (g1500) & (!g276) & (g311)) + ((g1497) & (g1498) & (g1499) & (!g1500) & (!g276) & (!g311)) + ((g1497) & (g1498) & (g1499) & (!g1500) & (g276) & (g311)) + ((g1497) & (g1498) & (g1499) & (g1500) & (!g276) & (!g311)));
	assign g1503 = (((!sk[80]) & (!g1157) & (g1502)) + ((!sk[80]) & (g1157) & (g1502)) + ((sk[80]) & (!g1157) & (g1502)) + ((sk[80]) & (g1157) & (!g1502)));
	assign g1504 = (((!g645) & (!sk[81]) & (!g901) & (g1501) & (!g1503)) + ((!g645) & (!sk[81]) & (!g901) & (g1501) & (g1503)) + ((!g645) & (!sk[81]) & (g901) & (!g1501) & (!g1503)) + ((!g645) & (!sk[81]) & (g901) & (!g1501) & (g1503)) + ((!g645) & (!sk[81]) & (g901) & (g1501) & (!g1503)) + ((!g645) & (!sk[81]) & (g901) & (g1501) & (g1503)) + ((!g645) & (sk[81]) & (!g901) & (!g1501) & (g1503)) + ((!g645) & (sk[81]) & (!g901) & (g1501) & (!g1503)) + ((!g645) & (sk[81]) & (g901) & (!g1501) & (!g1503)) + ((!g645) & (sk[81]) & (g901) & (g1501) & (g1503)) + ((g645) & (!sk[81]) & (!g901) & (g1501) & (!g1503)) + ((g645) & (!sk[81]) & (!g901) & (g1501) & (g1503)) + ((g645) & (!sk[81]) & (g901) & (!g1501) & (!g1503)) + ((g645) & (!sk[81]) & (g901) & (!g1501) & (g1503)) + ((g645) & (!sk[81]) & (g901) & (g1501) & (!g1503)) + ((g645) & (!sk[81]) & (g901) & (g1501) & (g1503)) + ((g645) & (sk[81]) & (!g901) & (!g1501) & (!g1503)) + ((g645) & (sk[81]) & (!g901) & (g1501) & (g1503)) + ((g645) & (sk[81]) & (g901) & (!g1501) & (g1503)) + ((g645) & (sk[81]) & (g901) & (g1501) & (!g1503)));
	assign g1505 = (((!ld) & (!sk[82]) & (!g389) & (g1504) & (!keyx31x)) + ((!ld) & (!sk[82]) & (!g389) & (g1504) & (keyx31x)) + ((!ld) & (!sk[82]) & (g389) & (!g1504) & (!keyx31x)) + ((!ld) & (!sk[82]) & (g389) & (!g1504) & (keyx31x)) + ((!ld) & (!sk[82]) & (g389) & (g1504) & (!keyx31x)) + ((!ld) & (!sk[82]) & (g389) & (g1504) & (keyx31x)) + ((!ld) & (sk[82]) & (!g389) & (g1504) & (!keyx31x)) + ((!ld) & (sk[82]) & (!g389) & (g1504) & (keyx31x)) + ((!ld) & (sk[82]) & (g389) & (!g1504) & (!keyx31x)) + ((!ld) & (sk[82]) & (g389) & (!g1504) & (keyx31x)) + ((ld) & (!sk[82]) & (!g389) & (g1504) & (!keyx31x)) + ((ld) & (!sk[82]) & (!g389) & (g1504) & (keyx31x)) + ((ld) & (!sk[82]) & (g389) & (!g1504) & (!keyx31x)) + ((ld) & (!sk[82]) & (g389) & (!g1504) & (keyx31x)) + ((ld) & (!sk[82]) & (g389) & (g1504) & (!keyx31x)) + ((ld) & (!sk[82]) & (g389) & (g1504) & (keyx31x)) + ((ld) & (sk[82]) & (!g389) & (!g1504) & (keyx31x)) + ((ld) & (sk[82]) & (!g389) & (g1504) & (keyx31x)) + ((ld) & (sk[82]) & (g389) & (!g1504) & (keyx31x)) + ((ld) & (sk[82]) & (g389) & (g1504) & (keyx31x)));
	assign g2114 = (((!sk[83]) & (!ld) & (text_inx64x) & (!g1506)) + ((!sk[83]) & (!ld) & (text_inx64x) & (g1506)) + ((!sk[83]) & (ld) & (!text_inx64x) & (g1506)) + ((!sk[83]) & (ld) & (text_inx64x) & (!g1506)) + ((!sk[83]) & (ld) & (text_inx64x) & (g1506)) + ((sk[83]) & (!ld) & (!text_inx64x) & (g1506)) + ((sk[83]) & (!ld) & (text_inx64x) & (g1506)) + ((sk[83]) & (ld) & (text_inx64x) & (!g1506)) + ((sk[83]) & (ld) & (text_inx64x) & (g1506)));
	assign g1507 = (((!g660) & (!g723) & (!g1163) & (!g1247) & (g1269) & (!g1506)) + ((!g660) & (!g723) & (!g1163) & (!g1247) & (g1269) & (g1506)) + ((!g660) & (!g723) & (!g1163) & (g1247) & (!g1269) & (!g1506)) + ((!g660) & (!g723) & (!g1163) & (g1247) & (!g1269) & (g1506)) + ((!g660) & (!g723) & (g1163) & (!g1247) & (!g1269) & (g1506)) + ((!g660) & (!g723) & (g1163) & (!g1247) & (g1269) & (g1506)) + ((!g660) & (!g723) & (g1163) & (g1247) & (!g1269) & (g1506)) + ((!g660) & (!g723) & (g1163) & (g1247) & (g1269) & (g1506)) + ((!g660) & (g723) & (!g1163) & (!g1247) & (!g1269) & (!g1506)) + ((!g660) & (g723) & (!g1163) & (!g1247) & (!g1269) & (g1506)) + ((!g660) & (g723) & (!g1163) & (g1247) & (g1269) & (!g1506)) + ((!g660) & (g723) & (!g1163) & (g1247) & (g1269) & (g1506)) + ((!g660) & (g723) & (g1163) & (!g1247) & (!g1269) & (g1506)) + ((!g660) & (g723) & (g1163) & (!g1247) & (g1269) & (g1506)) + ((!g660) & (g723) & (g1163) & (g1247) & (!g1269) & (g1506)) + ((!g660) & (g723) & (g1163) & (g1247) & (g1269) & (g1506)) + ((g660) & (!g723) & (!g1163) & (!g1247) & (!g1269) & (!g1506)) + ((g660) & (!g723) & (!g1163) & (!g1247) & (!g1269) & (g1506)) + ((g660) & (!g723) & (!g1163) & (g1247) & (g1269) & (!g1506)) + ((g660) & (!g723) & (!g1163) & (g1247) & (g1269) & (g1506)) + ((g660) & (!g723) & (g1163) & (!g1247) & (!g1269) & (!g1506)) + ((g660) & (!g723) & (g1163) & (!g1247) & (g1269) & (!g1506)) + ((g660) & (!g723) & (g1163) & (g1247) & (!g1269) & (!g1506)) + ((g660) & (!g723) & (g1163) & (g1247) & (g1269) & (!g1506)) + ((g660) & (g723) & (!g1163) & (!g1247) & (g1269) & (!g1506)) + ((g660) & (g723) & (!g1163) & (!g1247) & (g1269) & (g1506)) + ((g660) & (g723) & (!g1163) & (g1247) & (!g1269) & (!g1506)) + ((g660) & (g723) & (!g1163) & (g1247) & (!g1269) & (g1506)) + ((g660) & (g723) & (g1163) & (!g1247) & (!g1269) & (!g1506)) + ((g660) & (g723) & (g1163) & (!g1247) & (g1269) & (!g1506)) + ((g660) & (g723) & (g1163) & (g1247) & (!g1269) & (!g1506)) + ((g660) & (g723) & (g1163) & (g1247) & (g1269) & (!g1506)));
	assign g2115 = (((!ld) & (!sk[85]) & (text_inx65x) & (!g1508)) + ((!ld) & (!sk[85]) & (text_inx65x) & (g1508)) + ((!ld) & (sk[85]) & (!text_inx65x) & (g1508)) + ((!ld) & (sk[85]) & (text_inx65x) & (g1508)) + ((ld) & (!sk[85]) & (!text_inx65x) & (g1508)) + ((ld) & (!sk[85]) & (text_inx65x) & (!g1508)) + ((ld) & (!sk[85]) & (text_inx65x) & (g1508)) + ((ld) & (sk[85]) & (text_inx65x) & (!g1508)) + ((ld) & (sk[85]) & (text_inx65x) & (g1508)));
	assign g1509 = (((!sk[86]) & (!g659) & (g667) & (!g730) & (!g794) & (!g851)) + ((!sk[86]) & (!g659) & (g667) & (!g730) & (!g794) & (g851)) + ((!sk[86]) & (!g659) & (g667) & (!g730) & (g794) & (!g851)) + ((!sk[86]) & (!g659) & (g667) & (!g730) & (g794) & (g851)) + ((!sk[86]) & (!g659) & (g667) & (g730) & (!g794) & (!g851)) + ((!sk[86]) & (!g659) & (g667) & (g730) & (!g794) & (g851)) + ((!sk[86]) & (!g659) & (g667) & (g730) & (g794) & (!g851)) + ((!sk[86]) & (!g659) & (g667) & (g730) & (g794) & (g851)) + ((!sk[86]) & (g659) & (!g667) & (!g730) & (!g794) & (!g851)) + ((!sk[86]) & (g659) & (!g667) & (!g730) & (!g794) & (g851)) + ((!sk[86]) & (g659) & (!g667) & (!g730) & (g794) & (!g851)) + ((!sk[86]) & (g659) & (!g667) & (!g730) & (g794) & (g851)) + ((!sk[86]) & (g659) & (!g667) & (g730) & (!g794) & (!g851)) + ((!sk[86]) & (g659) & (!g667) & (g730) & (!g794) & (g851)) + ((!sk[86]) & (g659) & (!g667) & (g730) & (g794) & (!g851)) + ((!sk[86]) & (g659) & (!g667) & (g730) & (g794) & (g851)) + ((!sk[86]) & (g659) & (g667) & (!g730) & (!g794) & (!g851)) + ((!sk[86]) & (g659) & (g667) & (!g730) & (!g794) & (g851)) + ((!sk[86]) & (g659) & (g667) & (!g730) & (g794) & (!g851)) + ((!sk[86]) & (g659) & (g667) & (!g730) & (g794) & (g851)) + ((!sk[86]) & (g659) & (g667) & (g730) & (!g794) & (!g851)) + ((!sk[86]) & (g659) & (g667) & (g730) & (!g794) & (g851)) + ((!sk[86]) & (g659) & (g667) & (g730) & (g794) & (!g851)) + ((!sk[86]) & (g659) & (g667) & (g730) & (g794) & (g851)) + ((sk[86]) & (!g659) & (!g667) & (!g730) & (!g794) & (g851)) + ((sk[86]) & (!g659) & (!g667) & (!g730) & (g794) & (!g851)) + ((sk[86]) & (!g659) & (!g667) & (g730) & (!g794) & (!g851)) + ((sk[86]) & (!g659) & (!g667) & (g730) & (g794) & (g851)) + ((sk[86]) & (!g659) & (g667) & (!g730) & (!g794) & (!g851)) + ((sk[86]) & (!g659) & (g667) & (!g730) & (g794) & (g851)) + ((sk[86]) & (!g659) & (g667) & (g730) & (!g794) & (g851)) + ((sk[86]) & (!g659) & (g667) & (g730) & (g794) & (!g851)) + ((sk[86]) & (g659) & (!g667) & (!g730) & (!g794) & (!g851)) + ((sk[86]) & (g659) & (!g667) & (!g730) & (g794) & (g851)) + ((sk[86]) & (g659) & (!g667) & (g730) & (!g794) & (g851)) + ((sk[86]) & (g659) & (!g667) & (g730) & (g794) & (!g851)) + ((sk[86]) & (g659) & (g667) & (!g730) & (!g794) & (g851)) + ((sk[86]) & (g659) & (g667) & (!g730) & (g794) & (!g851)) + ((sk[86]) & (g659) & (g667) & (g730) & (!g794) & (!g851)) + ((sk[86]) & (g659) & (g667) & (g730) & (g794) & (g851)));
	assign g1510 = (((!g667) & (!g858) & (!g1163) & (!g1269) & (!g1508) & (g1509)) + ((!g667) & (!g858) & (!g1163) & (!g1269) & (g1508) & (g1509)) + ((!g667) & (!g858) & (!g1163) & (g1269) & (!g1508) & (!g1509)) + ((!g667) & (!g858) & (!g1163) & (g1269) & (g1508) & (!g1509)) + ((!g667) & (!g858) & (g1163) & (!g1269) & (g1508) & (!g1509)) + ((!g667) & (!g858) & (g1163) & (!g1269) & (g1508) & (g1509)) + ((!g667) & (!g858) & (g1163) & (g1269) & (g1508) & (!g1509)) + ((!g667) & (!g858) & (g1163) & (g1269) & (g1508) & (g1509)) + ((!g667) & (g858) & (!g1163) & (!g1269) & (!g1508) & (!g1509)) + ((!g667) & (g858) & (!g1163) & (!g1269) & (g1508) & (!g1509)) + ((!g667) & (g858) & (!g1163) & (g1269) & (!g1508) & (g1509)) + ((!g667) & (g858) & (!g1163) & (g1269) & (g1508) & (g1509)) + ((!g667) & (g858) & (g1163) & (!g1269) & (g1508) & (!g1509)) + ((!g667) & (g858) & (g1163) & (!g1269) & (g1508) & (g1509)) + ((!g667) & (g858) & (g1163) & (g1269) & (g1508) & (!g1509)) + ((!g667) & (g858) & (g1163) & (g1269) & (g1508) & (g1509)) + ((g667) & (!g858) & (!g1163) & (!g1269) & (!g1508) & (g1509)) + ((g667) & (!g858) & (!g1163) & (!g1269) & (g1508) & (g1509)) + ((g667) & (!g858) & (!g1163) & (g1269) & (!g1508) & (!g1509)) + ((g667) & (!g858) & (!g1163) & (g1269) & (g1508) & (!g1509)) + ((g667) & (!g858) & (g1163) & (!g1269) & (!g1508) & (!g1509)) + ((g667) & (!g858) & (g1163) & (!g1269) & (!g1508) & (g1509)) + ((g667) & (!g858) & (g1163) & (g1269) & (!g1508) & (!g1509)) + ((g667) & (!g858) & (g1163) & (g1269) & (!g1508) & (g1509)) + ((g667) & (g858) & (!g1163) & (!g1269) & (!g1508) & (!g1509)) + ((g667) & (g858) & (!g1163) & (!g1269) & (g1508) & (!g1509)) + ((g667) & (g858) & (!g1163) & (g1269) & (!g1508) & (g1509)) + ((g667) & (g858) & (!g1163) & (g1269) & (g1508) & (g1509)) + ((g667) & (g858) & (g1163) & (!g1269) & (!g1508) & (!g1509)) + ((g667) & (g858) & (g1163) & (!g1269) & (!g1508) & (g1509)) + ((g667) & (g858) & (g1163) & (g1269) & (!g1508) & (!g1509)) + ((g667) & (g858) & (g1163) & (g1269) & (!g1508) & (g1509)));
	assign g2116 = (((!sk[88]) & (!ld) & (text_inx66x) & (!g1511)) + ((!sk[88]) & (!ld) & (text_inx66x) & (g1511)) + ((!sk[88]) & (ld) & (!text_inx66x) & (g1511)) + ((!sk[88]) & (ld) & (text_inx66x) & (!g1511)) + ((!sk[88]) & (ld) & (text_inx66x) & (g1511)) + ((sk[88]) & (!ld) & (!text_inx66x) & (g1511)) + ((sk[88]) & (!ld) & (text_inx66x) & (g1511)) + ((sk[88]) & (ld) & (text_inx66x) & (!g1511)) + ((sk[88]) & (ld) & (text_inx66x) & (g1511)));
	assign g1512 = (((!g674) & (!g737) & (!g858) & (!g1163) & (g1254) & (!g1511)) + ((!g674) & (!g737) & (!g858) & (!g1163) & (g1254) & (g1511)) + ((!g674) & (!g737) & (!g858) & (g1163) & (!g1254) & (g1511)) + ((!g674) & (!g737) & (!g858) & (g1163) & (g1254) & (g1511)) + ((!g674) & (!g737) & (g858) & (!g1163) & (!g1254) & (!g1511)) + ((!g674) & (!g737) & (g858) & (!g1163) & (!g1254) & (g1511)) + ((!g674) & (!g737) & (g858) & (g1163) & (!g1254) & (g1511)) + ((!g674) & (!g737) & (g858) & (g1163) & (g1254) & (g1511)) + ((!g674) & (g737) & (!g858) & (!g1163) & (!g1254) & (!g1511)) + ((!g674) & (g737) & (!g858) & (!g1163) & (!g1254) & (g1511)) + ((!g674) & (g737) & (!g858) & (g1163) & (!g1254) & (g1511)) + ((!g674) & (g737) & (!g858) & (g1163) & (g1254) & (g1511)) + ((!g674) & (g737) & (g858) & (!g1163) & (g1254) & (!g1511)) + ((!g674) & (g737) & (g858) & (!g1163) & (g1254) & (g1511)) + ((!g674) & (g737) & (g858) & (g1163) & (!g1254) & (g1511)) + ((!g674) & (g737) & (g858) & (g1163) & (g1254) & (g1511)) + ((g674) & (!g737) & (!g858) & (!g1163) & (!g1254) & (!g1511)) + ((g674) & (!g737) & (!g858) & (!g1163) & (!g1254) & (g1511)) + ((g674) & (!g737) & (!g858) & (g1163) & (!g1254) & (!g1511)) + ((g674) & (!g737) & (!g858) & (g1163) & (g1254) & (!g1511)) + ((g674) & (!g737) & (g858) & (!g1163) & (g1254) & (!g1511)) + ((g674) & (!g737) & (g858) & (!g1163) & (g1254) & (g1511)) + ((g674) & (!g737) & (g858) & (g1163) & (!g1254) & (!g1511)) + ((g674) & (!g737) & (g858) & (g1163) & (g1254) & (!g1511)) + ((g674) & (g737) & (!g858) & (!g1163) & (g1254) & (!g1511)) + ((g674) & (g737) & (!g858) & (!g1163) & (g1254) & (g1511)) + ((g674) & (g737) & (!g858) & (g1163) & (!g1254) & (!g1511)) + ((g674) & (g737) & (!g858) & (g1163) & (g1254) & (!g1511)) + ((g674) & (g737) & (g858) & (!g1163) & (!g1254) & (!g1511)) + ((g674) & (g737) & (g858) & (!g1163) & (!g1254) & (g1511)) + ((g674) & (g737) & (g858) & (g1163) & (!g1254) & (!g1511)) + ((g674) & (g737) & (g858) & (g1163) & (g1254) & (!g1511)));
	assign g2117 = (((!sk[90]) & (!ld) & (text_inx67x) & (!g1513)) + ((!sk[90]) & (!ld) & (text_inx67x) & (g1513)) + ((!sk[90]) & (ld) & (!text_inx67x) & (g1513)) + ((!sk[90]) & (ld) & (text_inx67x) & (!g1513)) + ((!sk[90]) & (ld) & (text_inx67x) & (g1513)) + ((sk[90]) & (!ld) & (!text_inx67x) & (g1513)) + ((sk[90]) & (!ld) & (text_inx67x) & (g1513)) + ((sk[90]) & (ld) & (text_inx67x) & (!g1513)) + ((sk[90]) & (ld) & (text_inx67x) & (g1513)));
	assign g1514 = (((!g744) & (!g808) & (!sk[91]) & (g865) & (!g900)) + ((!g744) & (!g808) & (!sk[91]) & (g865) & (g900)) + ((!g744) & (!g808) & (sk[91]) & (!g865) & (g900)) + ((!g744) & (!g808) & (sk[91]) & (g865) & (!g900)) + ((!g744) & (g808) & (!sk[91]) & (!g865) & (!g900)) + ((!g744) & (g808) & (!sk[91]) & (!g865) & (g900)) + ((!g744) & (g808) & (!sk[91]) & (g865) & (!g900)) + ((!g744) & (g808) & (!sk[91]) & (g865) & (g900)) + ((!g744) & (g808) & (sk[91]) & (!g865) & (!g900)) + ((!g744) & (g808) & (sk[91]) & (g865) & (g900)) + ((g744) & (!g808) & (!sk[91]) & (g865) & (!g900)) + ((g744) & (!g808) & (!sk[91]) & (g865) & (g900)) + ((g744) & (!g808) & (sk[91]) & (!g865) & (!g900)) + ((g744) & (!g808) & (sk[91]) & (g865) & (g900)) + ((g744) & (g808) & (!sk[91]) & (!g865) & (!g900)) + ((g744) & (g808) & (!sk[91]) & (!g865) & (g900)) + ((g744) & (g808) & (!sk[91]) & (g865) & (!g900)) + ((g744) & (g808) & (!sk[91]) & (g865) & (g900)) + ((g744) & (g808) & (sk[91]) & (!g865) & (g900)) + ((g744) & (g808) & (sk[91]) & (g865) & (!g900)));
	assign g2118 = (((!sk[92]) & (!ld) & (text_inx70x) & (!g1515)) + ((!sk[92]) & (!ld) & (text_inx70x) & (g1515)) + ((!sk[92]) & (ld) & (!text_inx70x) & (g1515)) + ((!sk[92]) & (ld) & (text_inx70x) & (!g1515)) + ((!sk[92]) & (ld) & (text_inx70x) & (g1515)) + ((sk[92]) & (!ld) & (!text_inx70x) & (g1515)) + ((sk[92]) & (!ld) & (text_inx70x) & (g1515)) + ((sk[92]) & (ld) & (text_inx70x) & (!g1515)) + ((sk[92]) & (ld) & (text_inx70x) & (g1515)));
	assign g1516 = (((!g702) & (!g765) & (!g886) & (!g1163) & (g1260) & (!g1515)) + ((!g702) & (!g765) & (!g886) & (!g1163) & (g1260) & (g1515)) + ((!g702) & (!g765) & (!g886) & (g1163) & (!g1260) & (g1515)) + ((!g702) & (!g765) & (!g886) & (g1163) & (g1260) & (g1515)) + ((!g702) & (!g765) & (g886) & (!g1163) & (!g1260) & (!g1515)) + ((!g702) & (!g765) & (g886) & (!g1163) & (!g1260) & (g1515)) + ((!g702) & (!g765) & (g886) & (g1163) & (!g1260) & (g1515)) + ((!g702) & (!g765) & (g886) & (g1163) & (g1260) & (g1515)) + ((!g702) & (g765) & (!g886) & (!g1163) & (!g1260) & (!g1515)) + ((!g702) & (g765) & (!g886) & (!g1163) & (!g1260) & (g1515)) + ((!g702) & (g765) & (!g886) & (g1163) & (!g1260) & (g1515)) + ((!g702) & (g765) & (!g886) & (g1163) & (g1260) & (g1515)) + ((!g702) & (g765) & (g886) & (!g1163) & (g1260) & (!g1515)) + ((!g702) & (g765) & (g886) & (!g1163) & (g1260) & (g1515)) + ((!g702) & (g765) & (g886) & (g1163) & (!g1260) & (g1515)) + ((!g702) & (g765) & (g886) & (g1163) & (g1260) & (g1515)) + ((g702) & (!g765) & (!g886) & (!g1163) & (!g1260) & (!g1515)) + ((g702) & (!g765) & (!g886) & (!g1163) & (!g1260) & (g1515)) + ((g702) & (!g765) & (!g886) & (g1163) & (!g1260) & (!g1515)) + ((g702) & (!g765) & (!g886) & (g1163) & (g1260) & (!g1515)) + ((g702) & (!g765) & (g886) & (!g1163) & (g1260) & (!g1515)) + ((g702) & (!g765) & (g886) & (!g1163) & (g1260) & (g1515)) + ((g702) & (!g765) & (g886) & (g1163) & (!g1260) & (!g1515)) + ((g702) & (!g765) & (g886) & (g1163) & (g1260) & (!g1515)) + ((g702) & (g765) & (!g886) & (!g1163) & (g1260) & (!g1515)) + ((g702) & (g765) & (!g886) & (!g1163) & (g1260) & (g1515)) + ((g702) & (g765) & (!g886) & (g1163) & (!g1260) & (!g1515)) + ((g702) & (g765) & (!g886) & (g1163) & (g1260) & (!g1515)) + ((g702) & (g765) & (g886) & (!g1163) & (!g1260) & (!g1515)) + ((g702) & (g765) & (g886) & (!g1163) & (!g1260) & (g1515)) + ((g702) & (g765) & (g886) & (g1163) & (!g1260) & (!g1515)) + ((g702) & (g765) & (g886) & (g1163) & (g1260) & (!g1515)));
	assign g2119 = (((!ld) & (!sk[94]) & (text_inx69x) & (!g1517)) + ((!ld) & (!sk[94]) & (text_inx69x) & (g1517)) + ((!ld) & (sk[94]) & (!text_inx69x) & (g1517)) + ((!ld) & (sk[94]) & (text_inx69x) & (g1517)) + ((ld) & (!sk[94]) & (!text_inx69x) & (g1517)) + ((ld) & (!sk[94]) & (text_inx69x) & (!g1517)) + ((ld) & (!sk[94]) & (text_inx69x) & (g1517)) + ((ld) & (sk[94]) & (text_inx69x) & (!g1517)) + ((ld) & (sk[94]) & (text_inx69x) & (g1517)));
	assign g1518 = (((!g695) & (!g758) & (!g879) & (!g1163) & (g1263) & (!g1517)) + ((!g695) & (!g758) & (!g879) & (!g1163) & (g1263) & (g1517)) + ((!g695) & (!g758) & (!g879) & (g1163) & (!g1263) & (g1517)) + ((!g695) & (!g758) & (!g879) & (g1163) & (g1263) & (g1517)) + ((!g695) & (!g758) & (g879) & (!g1163) & (!g1263) & (!g1517)) + ((!g695) & (!g758) & (g879) & (!g1163) & (!g1263) & (g1517)) + ((!g695) & (!g758) & (g879) & (g1163) & (!g1263) & (g1517)) + ((!g695) & (!g758) & (g879) & (g1163) & (g1263) & (g1517)) + ((!g695) & (g758) & (!g879) & (!g1163) & (!g1263) & (!g1517)) + ((!g695) & (g758) & (!g879) & (!g1163) & (!g1263) & (g1517)) + ((!g695) & (g758) & (!g879) & (g1163) & (!g1263) & (g1517)) + ((!g695) & (g758) & (!g879) & (g1163) & (g1263) & (g1517)) + ((!g695) & (g758) & (g879) & (!g1163) & (g1263) & (!g1517)) + ((!g695) & (g758) & (g879) & (!g1163) & (g1263) & (g1517)) + ((!g695) & (g758) & (g879) & (g1163) & (!g1263) & (g1517)) + ((!g695) & (g758) & (g879) & (g1163) & (g1263) & (g1517)) + ((g695) & (!g758) & (!g879) & (!g1163) & (!g1263) & (!g1517)) + ((g695) & (!g758) & (!g879) & (!g1163) & (!g1263) & (g1517)) + ((g695) & (!g758) & (!g879) & (g1163) & (!g1263) & (!g1517)) + ((g695) & (!g758) & (!g879) & (g1163) & (g1263) & (!g1517)) + ((g695) & (!g758) & (g879) & (!g1163) & (g1263) & (!g1517)) + ((g695) & (!g758) & (g879) & (!g1163) & (g1263) & (g1517)) + ((g695) & (!g758) & (g879) & (g1163) & (!g1263) & (!g1517)) + ((g695) & (!g758) & (g879) & (g1163) & (g1263) & (!g1517)) + ((g695) & (g758) & (!g879) & (!g1163) & (g1263) & (!g1517)) + ((g695) & (g758) & (!g879) & (!g1163) & (g1263) & (g1517)) + ((g695) & (g758) & (!g879) & (g1163) & (!g1263) & (!g1517)) + ((g695) & (g758) & (!g879) & (g1163) & (g1263) & (!g1517)) + ((g695) & (g758) & (g879) & (!g1163) & (!g1263) & (!g1517)) + ((g695) & (g758) & (g879) & (!g1163) & (!g1263) & (g1517)) + ((g695) & (g758) & (g879) & (g1163) & (!g1263) & (!g1517)) + ((g695) & (g758) & (g879) & (g1163) & (g1263) & (!g1517)));
	assign g2120 = (((!ld) & (!text_inx68x) & (sk[96]) & (g1519)) + ((!ld) & (text_inx68x) & (!sk[96]) & (!g1519)) + ((!ld) & (text_inx68x) & (!sk[96]) & (g1519)) + ((!ld) & (text_inx68x) & (sk[96]) & (g1519)) + ((ld) & (!text_inx68x) & (!sk[96]) & (g1519)) + ((ld) & (text_inx68x) & (!sk[96]) & (!g1519)) + ((ld) & (text_inx68x) & (!sk[96]) & (g1519)) + ((ld) & (text_inx68x) & (sk[96]) & (!g1519)) + ((ld) & (text_inx68x) & (sk[96]) & (g1519)));
	assign g1520 = (((!g680) & (!g688) & (!g708) & (!g751) & (!g872) & (g900)) + ((!g680) & (!g688) & (!g708) & (!g751) & (g872) & (!g900)) + ((!g680) & (!g688) & (!g708) & (g751) & (!g872) & (!g900)) + ((!g680) & (!g688) & (!g708) & (g751) & (g872) & (g900)) + ((!g680) & (!g688) & (g708) & (!g751) & (!g872) & (!g900)) + ((!g680) & (!g688) & (g708) & (!g751) & (g872) & (g900)) + ((!g680) & (!g688) & (g708) & (g751) & (!g872) & (g900)) + ((!g680) & (!g688) & (g708) & (g751) & (g872) & (!g900)) + ((!g680) & (g688) & (!g708) & (!g751) & (!g872) & (!g900)) + ((!g680) & (g688) & (!g708) & (!g751) & (g872) & (g900)) + ((!g680) & (g688) & (!g708) & (g751) & (!g872) & (g900)) + ((!g680) & (g688) & (!g708) & (g751) & (g872) & (!g900)) + ((!g680) & (g688) & (g708) & (!g751) & (!g872) & (g900)) + ((!g680) & (g688) & (g708) & (!g751) & (g872) & (!g900)) + ((!g680) & (g688) & (g708) & (g751) & (!g872) & (!g900)) + ((!g680) & (g688) & (g708) & (g751) & (g872) & (g900)) + ((g680) & (!g688) & (!g708) & (!g751) & (!g872) & (!g900)) + ((g680) & (!g688) & (!g708) & (!g751) & (g872) & (g900)) + ((g680) & (!g688) & (!g708) & (g751) & (!g872) & (g900)) + ((g680) & (!g688) & (!g708) & (g751) & (g872) & (!g900)) + ((g680) & (!g688) & (g708) & (!g751) & (!g872) & (g900)) + ((g680) & (!g688) & (g708) & (!g751) & (g872) & (!g900)) + ((g680) & (!g688) & (g708) & (g751) & (!g872) & (!g900)) + ((g680) & (!g688) & (g708) & (g751) & (g872) & (g900)) + ((g680) & (g688) & (!g708) & (!g751) & (!g872) & (g900)) + ((g680) & (g688) & (!g708) & (!g751) & (g872) & (!g900)) + ((g680) & (g688) & (!g708) & (g751) & (!g872) & (!g900)) + ((g680) & (g688) & (!g708) & (g751) & (g872) & (g900)) + ((g680) & (g688) & (g708) & (!g751) & (!g872) & (!g900)) + ((g680) & (g688) & (g708) & (!g751) & (g872) & (g900)) + ((g680) & (g688) & (g708) & (g751) & (!g872) & (g900)) + ((g680) & (g688) & (g708) & (g751) & (g872) & (!g900)));
	assign g1521 = (((!g688) & (!g815) & (!g879) & (!g1163) & (!g1519) & (g1520)) + ((!g688) & (!g815) & (!g879) & (!g1163) & (g1519) & (g1520)) + ((!g688) & (!g815) & (!g879) & (g1163) & (g1519) & (!g1520)) + ((!g688) & (!g815) & (!g879) & (g1163) & (g1519) & (g1520)) + ((!g688) & (!g815) & (g879) & (!g1163) & (!g1519) & (!g1520)) + ((!g688) & (!g815) & (g879) & (!g1163) & (g1519) & (!g1520)) + ((!g688) & (!g815) & (g879) & (g1163) & (g1519) & (!g1520)) + ((!g688) & (!g815) & (g879) & (g1163) & (g1519) & (g1520)) + ((!g688) & (g815) & (!g879) & (!g1163) & (!g1519) & (!g1520)) + ((!g688) & (g815) & (!g879) & (!g1163) & (g1519) & (!g1520)) + ((!g688) & (g815) & (!g879) & (g1163) & (g1519) & (!g1520)) + ((!g688) & (g815) & (!g879) & (g1163) & (g1519) & (g1520)) + ((!g688) & (g815) & (g879) & (!g1163) & (!g1519) & (g1520)) + ((!g688) & (g815) & (g879) & (!g1163) & (g1519) & (g1520)) + ((!g688) & (g815) & (g879) & (g1163) & (g1519) & (!g1520)) + ((!g688) & (g815) & (g879) & (g1163) & (g1519) & (g1520)) + ((g688) & (!g815) & (!g879) & (!g1163) & (!g1519) & (g1520)) + ((g688) & (!g815) & (!g879) & (!g1163) & (g1519) & (g1520)) + ((g688) & (!g815) & (!g879) & (g1163) & (!g1519) & (!g1520)) + ((g688) & (!g815) & (!g879) & (g1163) & (!g1519) & (g1520)) + ((g688) & (!g815) & (g879) & (!g1163) & (!g1519) & (!g1520)) + ((g688) & (!g815) & (g879) & (!g1163) & (g1519) & (!g1520)) + ((g688) & (!g815) & (g879) & (g1163) & (!g1519) & (!g1520)) + ((g688) & (!g815) & (g879) & (g1163) & (!g1519) & (g1520)) + ((g688) & (g815) & (!g879) & (!g1163) & (!g1519) & (!g1520)) + ((g688) & (g815) & (!g879) & (!g1163) & (g1519) & (!g1520)) + ((g688) & (g815) & (!g879) & (g1163) & (!g1519) & (!g1520)) + ((g688) & (g815) & (!g879) & (g1163) & (!g1519) & (g1520)) + ((g688) & (g815) & (g879) & (!g1163) & (!g1519) & (g1520)) + ((g688) & (g815) & (g879) & (!g1163) & (g1519) & (g1520)) + ((g688) & (g815) & (g879) & (g1163) & (!g1519) & (!g1520)) + ((g688) & (g815) & (g879) & (g1163) & (!g1519) & (g1520)));
	assign g2121 = (((!ld) & (!text_inx71x) & (sk[99]) & (g1522)) + ((!ld) & (text_inx71x) & (!sk[99]) & (!g1522)) + ((!ld) & (text_inx71x) & (!sk[99]) & (g1522)) + ((!ld) & (text_inx71x) & (sk[99]) & (g1522)) + ((ld) & (!text_inx71x) & (!sk[99]) & (g1522)) + ((ld) & (text_inx71x) & (!sk[99]) & (!g1522)) + ((ld) & (text_inx71x) & (!sk[99]) & (g1522)) + ((ld) & (text_inx71x) & (sk[99]) & (!g1522)) + ((ld) & (text_inx71x) & (sk[99]) & (g1522)));
	assign g1523 = (((!sk[100]) & (!g701) & (!g709) & (g893) & (!g900)) + ((!sk[100]) & (!g701) & (!g709) & (g893) & (g900)) + ((!sk[100]) & (!g701) & (g709) & (!g893) & (!g900)) + ((!sk[100]) & (!g701) & (g709) & (!g893) & (g900)) + ((!sk[100]) & (!g701) & (g709) & (g893) & (!g900)) + ((!sk[100]) & (!g701) & (g709) & (g893) & (g900)) + ((!sk[100]) & (g701) & (!g709) & (g893) & (!g900)) + ((!sk[100]) & (g701) & (!g709) & (g893) & (g900)) + ((!sk[100]) & (g701) & (g709) & (!g893) & (!g900)) + ((!sk[100]) & (g701) & (g709) & (!g893) & (g900)) + ((!sk[100]) & (g701) & (g709) & (g893) & (!g900)) + ((!sk[100]) & (g701) & (g709) & (g893) & (g900)) + ((sk[100]) & (!g701) & (!g709) & (!g893) & (g900)) + ((sk[100]) & (!g701) & (!g709) & (g893) & (!g900)) + ((sk[100]) & (!g701) & (g709) & (!g893) & (!g900)) + ((sk[100]) & (!g701) & (g709) & (g893) & (g900)) + ((sk[100]) & (g701) & (!g709) & (!g893) & (!g900)) + ((sk[100]) & (g701) & (!g709) & (g893) & (g900)) + ((sk[100]) & (g701) & (g709) & (!g893) & (g900)) + ((sk[100]) & (g701) & (g709) & (g893) & (!g900)));
	assign g1524 = (((!g709) & (!g772) & (!g836) & (!g1163) & (!g1522) & (g1523)) + ((!g709) & (!g772) & (!g836) & (!g1163) & (g1522) & (g1523)) + ((!g709) & (!g772) & (!g836) & (g1163) & (g1522) & (!g1523)) + ((!g709) & (!g772) & (!g836) & (g1163) & (g1522) & (g1523)) + ((!g709) & (!g772) & (g836) & (!g1163) & (!g1522) & (!g1523)) + ((!g709) & (!g772) & (g836) & (!g1163) & (g1522) & (!g1523)) + ((!g709) & (!g772) & (g836) & (g1163) & (g1522) & (!g1523)) + ((!g709) & (!g772) & (g836) & (g1163) & (g1522) & (g1523)) + ((!g709) & (g772) & (!g836) & (!g1163) & (!g1522) & (!g1523)) + ((!g709) & (g772) & (!g836) & (!g1163) & (g1522) & (!g1523)) + ((!g709) & (g772) & (!g836) & (g1163) & (g1522) & (!g1523)) + ((!g709) & (g772) & (!g836) & (g1163) & (g1522) & (g1523)) + ((!g709) & (g772) & (g836) & (!g1163) & (!g1522) & (g1523)) + ((!g709) & (g772) & (g836) & (!g1163) & (g1522) & (g1523)) + ((!g709) & (g772) & (g836) & (g1163) & (g1522) & (!g1523)) + ((!g709) & (g772) & (g836) & (g1163) & (g1522) & (g1523)) + ((g709) & (!g772) & (!g836) & (!g1163) & (!g1522) & (g1523)) + ((g709) & (!g772) & (!g836) & (!g1163) & (g1522) & (g1523)) + ((g709) & (!g772) & (!g836) & (g1163) & (!g1522) & (!g1523)) + ((g709) & (!g772) & (!g836) & (g1163) & (!g1522) & (g1523)) + ((g709) & (!g772) & (g836) & (!g1163) & (!g1522) & (!g1523)) + ((g709) & (!g772) & (g836) & (!g1163) & (g1522) & (!g1523)) + ((g709) & (!g772) & (g836) & (g1163) & (!g1522) & (!g1523)) + ((g709) & (!g772) & (g836) & (g1163) & (!g1522) & (g1523)) + ((g709) & (g772) & (!g836) & (!g1163) & (!g1522) & (!g1523)) + ((g709) & (g772) & (!g836) & (!g1163) & (g1522) & (!g1523)) + ((g709) & (g772) & (!g836) & (g1163) & (!g1522) & (!g1523)) + ((g709) & (g772) & (!g836) & (g1163) & (!g1522) & (g1523)) + ((g709) & (g772) & (g836) & (!g1163) & (!g1522) & (g1523)) + ((g709) & (g772) & (g836) & (!g1163) & (g1522) & (g1523)) + ((g709) & (g772) & (g836) & (g1163) & (!g1522) & (!g1523)) + ((g709) & (g772) & (g836) & (g1163) & (!g1522) & (g1523)));
	assign g1525 = (((!ld) & (!g404) & (!g660) & (!g916) & (g1193) & (!keyx32x)) + ((!ld) & (!g404) & (!g660) & (!g916) & (g1193) & (keyx32x)) + ((!ld) & (!g404) & (!g660) & (g916) & (!g1193) & (!keyx32x)) + ((!ld) & (!g404) & (!g660) & (g916) & (!g1193) & (keyx32x)) + ((!ld) & (!g404) & (g660) & (!g916) & (!g1193) & (!keyx32x)) + ((!ld) & (!g404) & (g660) & (!g916) & (!g1193) & (keyx32x)) + ((!ld) & (!g404) & (g660) & (g916) & (g1193) & (!keyx32x)) + ((!ld) & (!g404) & (g660) & (g916) & (g1193) & (keyx32x)) + ((!ld) & (g404) & (!g660) & (!g916) & (!g1193) & (!keyx32x)) + ((!ld) & (g404) & (!g660) & (!g916) & (!g1193) & (keyx32x)) + ((!ld) & (g404) & (!g660) & (g916) & (g1193) & (!keyx32x)) + ((!ld) & (g404) & (!g660) & (g916) & (g1193) & (keyx32x)) + ((!ld) & (g404) & (g660) & (!g916) & (g1193) & (!keyx32x)) + ((!ld) & (g404) & (g660) & (!g916) & (g1193) & (keyx32x)) + ((!ld) & (g404) & (g660) & (g916) & (!g1193) & (!keyx32x)) + ((!ld) & (g404) & (g660) & (g916) & (!g1193) & (keyx32x)) + ((ld) & (!g404) & (!g660) & (!g916) & (!g1193) & (keyx32x)) + ((ld) & (!g404) & (!g660) & (!g916) & (g1193) & (keyx32x)) + ((ld) & (!g404) & (!g660) & (g916) & (!g1193) & (keyx32x)) + ((ld) & (!g404) & (!g660) & (g916) & (g1193) & (keyx32x)) + ((ld) & (!g404) & (g660) & (!g916) & (!g1193) & (keyx32x)) + ((ld) & (!g404) & (g660) & (!g916) & (g1193) & (keyx32x)) + ((ld) & (!g404) & (g660) & (g916) & (!g1193) & (keyx32x)) + ((ld) & (!g404) & (g660) & (g916) & (g1193) & (keyx32x)) + ((ld) & (g404) & (!g660) & (!g916) & (!g1193) & (keyx32x)) + ((ld) & (g404) & (!g660) & (!g916) & (g1193) & (keyx32x)) + ((ld) & (g404) & (!g660) & (g916) & (!g1193) & (keyx32x)) + ((ld) & (g404) & (!g660) & (g916) & (g1193) & (keyx32x)) + ((ld) & (g404) & (g660) & (!g916) & (!g1193) & (keyx32x)) + ((ld) & (g404) & (g660) & (!g916) & (g1193) & (keyx32x)) + ((ld) & (g404) & (g660) & (g916) & (!g1193) & (keyx32x)) + ((ld) & (g404) & (g660) & (g916) & (g1193) & (keyx32x)));
	assign g1526 = (((!ld) & (!g411) & (!g667) & (!g923) & (g1200) & (!keyx33x)) + ((!ld) & (!g411) & (!g667) & (!g923) & (g1200) & (keyx33x)) + ((!ld) & (!g411) & (!g667) & (g923) & (!g1200) & (!keyx33x)) + ((!ld) & (!g411) & (!g667) & (g923) & (!g1200) & (keyx33x)) + ((!ld) & (!g411) & (g667) & (!g923) & (!g1200) & (!keyx33x)) + ((!ld) & (!g411) & (g667) & (!g923) & (!g1200) & (keyx33x)) + ((!ld) & (!g411) & (g667) & (g923) & (g1200) & (!keyx33x)) + ((!ld) & (!g411) & (g667) & (g923) & (g1200) & (keyx33x)) + ((!ld) & (g411) & (!g667) & (!g923) & (!g1200) & (!keyx33x)) + ((!ld) & (g411) & (!g667) & (!g923) & (!g1200) & (keyx33x)) + ((!ld) & (g411) & (!g667) & (g923) & (g1200) & (!keyx33x)) + ((!ld) & (g411) & (!g667) & (g923) & (g1200) & (keyx33x)) + ((!ld) & (g411) & (g667) & (!g923) & (g1200) & (!keyx33x)) + ((!ld) & (g411) & (g667) & (!g923) & (g1200) & (keyx33x)) + ((!ld) & (g411) & (g667) & (g923) & (!g1200) & (!keyx33x)) + ((!ld) & (g411) & (g667) & (g923) & (!g1200) & (keyx33x)) + ((ld) & (!g411) & (!g667) & (!g923) & (!g1200) & (keyx33x)) + ((ld) & (!g411) & (!g667) & (!g923) & (g1200) & (keyx33x)) + ((ld) & (!g411) & (!g667) & (g923) & (!g1200) & (keyx33x)) + ((ld) & (!g411) & (!g667) & (g923) & (g1200) & (keyx33x)) + ((ld) & (!g411) & (g667) & (!g923) & (!g1200) & (keyx33x)) + ((ld) & (!g411) & (g667) & (!g923) & (g1200) & (keyx33x)) + ((ld) & (!g411) & (g667) & (g923) & (!g1200) & (keyx33x)) + ((ld) & (!g411) & (g667) & (g923) & (g1200) & (keyx33x)) + ((ld) & (g411) & (!g667) & (!g923) & (!g1200) & (keyx33x)) + ((ld) & (g411) & (!g667) & (!g923) & (g1200) & (keyx33x)) + ((ld) & (g411) & (!g667) & (g923) & (!g1200) & (keyx33x)) + ((ld) & (g411) & (!g667) & (g923) & (g1200) & (keyx33x)) + ((ld) & (g411) & (g667) & (!g923) & (!g1200) & (keyx33x)) + ((ld) & (g411) & (g667) & (!g923) & (g1200) & (keyx33x)) + ((ld) & (g411) & (g667) & (g923) & (!g1200) & (keyx33x)) + ((ld) & (g411) & (g667) & (g923) & (g1200) & (keyx33x)));
	assign g1527 = (((!ld) & (!g418) & (!g674) & (!g930) & (g1207) & (!keyx34x)) + ((!ld) & (!g418) & (!g674) & (!g930) & (g1207) & (keyx34x)) + ((!ld) & (!g418) & (!g674) & (g930) & (!g1207) & (!keyx34x)) + ((!ld) & (!g418) & (!g674) & (g930) & (!g1207) & (keyx34x)) + ((!ld) & (!g418) & (g674) & (!g930) & (!g1207) & (!keyx34x)) + ((!ld) & (!g418) & (g674) & (!g930) & (!g1207) & (keyx34x)) + ((!ld) & (!g418) & (g674) & (g930) & (g1207) & (!keyx34x)) + ((!ld) & (!g418) & (g674) & (g930) & (g1207) & (keyx34x)) + ((!ld) & (g418) & (!g674) & (!g930) & (!g1207) & (!keyx34x)) + ((!ld) & (g418) & (!g674) & (!g930) & (!g1207) & (keyx34x)) + ((!ld) & (g418) & (!g674) & (g930) & (g1207) & (!keyx34x)) + ((!ld) & (g418) & (!g674) & (g930) & (g1207) & (keyx34x)) + ((!ld) & (g418) & (g674) & (!g930) & (g1207) & (!keyx34x)) + ((!ld) & (g418) & (g674) & (!g930) & (g1207) & (keyx34x)) + ((!ld) & (g418) & (g674) & (g930) & (!g1207) & (!keyx34x)) + ((!ld) & (g418) & (g674) & (g930) & (!g1207) & (keyx34x)) + ((ld) & (!g418) & (!g674) & (!g930) & (!g1207) & (keyx34x)) + ((ld) & (!g418) & (!g674) & (!g930) & (g1207) & (keyx34x)) + ((ld) & (!g418) & (!g674) & (g930) & (!g1207) & (keyx34x)) + ((ld) & (!g418) & (!g674) & (g930) & (g1207) & (keyx34x)) + ((ld) & (!g418) & (g674) & (!g930) & (!g1207) & (keyx34x)) + ((ld) & (!g418) & (g674) & (!g930) & (g1207) & (keyx34x)) + ((ld) & (!g418) & (g674) & (g930) & (!g1207) & (keyx34x)) + ((ld) & (!g418) & (g674) & (g930) & (g1207) & (keyx34x)) + ((ld) & (g418) & (!g674) & (!g930) & (!g1207) & (keyx34x)) + ((ld) & (g418) & (!g674) & (!g930) & (g1207) & (keyx34x)) + ((ld) & (g418) & (!g674) & (g930) & (!g1207) & (keyx34x)) + ((ld) & (g418) & (!g674) & (g930) & (g1207) & (keyx34x)) + ((ld) & (g418) & (g674) & (!g930) & (!g1207) & (keyx34x)) + ((ld) & (g418) & (g674) & (!g930) & (g1207) & (keyx34x)) + ((ld) & (g418) & (g674) & (g930) & (!g1207) & (keyx34x)) + ((ld) & (g418) & (g674) & (g930) & (g1207) & (keyx34x)));
	assign g1528 = (((!ld) & (!g425) & (!g681) & (!g937) & (g1214) & (!keyx35x)) + ((!ld) & (!g425) & (!g681) & (!g937) & (g1214) & (keyx35x)) + ((!ld) & (!g425) & (!g681) & (g937) & (!g1214) & (!keyx35x)) + ((!ld) & (!g425) & (!g681) & (g937) & (!g1214) & (keyx35x)) + ((!ld) & (!g425) & (g681) & (!g937) & (!g1214) & (!keyx35x)) + ((!ld) & (!g425) & (g681) & (!g937) & (!g1214) & (keyx35x)) + ((!ld) & (!g425) & (g681) & (g937) & (g1214) & (!keyx35x)) + ((!ld) & (!g425) & (g681) & (g937) & (g1214) & (keyx35x)) + ((!ld) & (g425) & (!g681) & (!g937) & (!g1214) & (!keyx35x)) + ((!ld) & (g425) & (!g681) & (!g937) & (!g1214) & (keyx35x)) + ((!ld) & (g425) & (!g681) & (g937) & (g1214) & (!keyx35x)) + ((!ld) & (g425) & (!g681) & (g937) & (g1214) & (keyx35x)) + ((!ld) & (g425) & (g681) & (!g937) & (g1214) & (!keyx35x)) + ((!ld) & (g425) & (g681) & (!g937) & (g1214) & (keyx35x)) + ((!ld) & (g425) & (g681) & (g937) & (!g1214) & (!keyx35x)) + ((!ld) & (g425) & (g681) & (g937) & (!g1214) & (keyx35x)) + ((ld) & (!g425) & (!g681) & (!g937) & (!g1214) & (keyx35x)) + ((ld) & (!g425) & (!g681) & (!g937) & (g1214) & (keyx35x)) + ((ld) & (!g425) & (!g681) & (g937) & (!g1214) & (keyx35x)) + ((ld) & (!g425) & (!g681) & (g937) & (g1214) & (keyx35x)) + ((ld) & (!g425) & (g681) & (!g937) & (!g1214) & (keyx35x)) + ((ld) & (!g425) & (g681) & (!g937) & (g1214) & (keyx35x)) + ((ld) & (!g425) & (g681) & (g937) & (!g1214) & (keyx35x)) + ((ld) & (!g425) & (g681) & (g937) & (g1214) & (keyx35x)) + ((ld) & (g425) & (!g681) & (!g937) & (!g1214) & (keyx35x)) + ((ld) & (g425) & (!g681) & (!g937) & (g1214) & (keyx35x)) + ((ld) & (g425) & (!g681) & (g937) & (!g1214) & (keyx35x)) + ((ld) & (g425) & (!g681) & (g937) & (g1214) & (keyx35x)) + ((ld) & (g425) & (g681) & (!g937) & (!g1214) & (keyx35x)) + ((ld) & (g425) & (g681) & (!g937) & (g1214) & (keyx35x)) + ((ld) & (g425) & (g681) & (g937) & (!g1214) & (keyx35x)) + ((ld) & (g425) & (g681) & (g937) & (g1214) & (keyx35x)));
	assign g1529 = (((!ld) & (!g432) & (!g688) & (!g944) & (g1221) & (!keyx36x)) + ((!ld) & (!g432) & (!g688) & (!g944) & (g1221) & (keyx36x)) + ((!ld) & (!g432) & (!g688) & (g944) & (!g1221) & (!keyx36x)) + ((!ld) & (!g432) & (!g688) & (g944) & (!g1221) & (keyx36x)) + ((!ld) & (!g432) & (g688) & (!g944) & (!g1221) & (!keyx36x)) + ((!ld) & (!g432) & (g688) & (!g944) & (!g1221) & (keyx36x)) + ((!ld) & (!g432) & (g688) & (g944) & (g1221) & (!keyx36x)) + ((!ld) & (!g432) & (g688) & (g944) & (g1221) & (keyx36x)) + ((!ld) & (g432) & (!g688) & (!g944) & (!g1221) & (!keyx36x)) + ((!ld) & (g432) & (!g688) & (!g944) & (!g1221) & (keyx36x)) + ((!ld) & (g432) & (!g688) & (g944) & (g1221) & (!keyx36x)) + ((!ld) & (g432) & (!g688) & (g944) & (g1221) & (keyx36x)) + ((!ld) & (g432) & (g688) & (!g944) & (g1221) & (!keyx36x)) + ((!ld) & (g432) & (g688) & (!g944) & (g1221) & (keyx36x)) + ((!ld) & (g432) & (g688) & (g944) & (!g1221) & (!keyx36x)) + ((!ld) & (g432) & (g688) & (g944) & (!g1221) & (keyx36x)) + ((ld) & (!g432) & (!g688) & (!g944) & (!g1221) & (keyx36x)) + ((ld) & (!g432) & (!g688) & (!g944) & (g1221) & (keyx36x)) + ((ld) & (!g432) & (!g688) & (g944) & (!g1221) & (keyx36x)) + ((ld) & (!g432) & (!g688) & (g944) & (g1221) & (keyx36x)) + ((ld) & (!g432) & (g688) & (!g944) & (!g1221) & (keyx36x)) + ((ld) & (!g432) & (g688) & (!g944) & (g1221) & (keyx36x)) + ((ld) & (!g432) & (g688) & (g944) & (!g1221) & (keyx36x)) + ((ld) & (!g432) & (g688) & (g944) & (g1221) & (keyx36x)) + ((ld) & (g432) & (!g688) & (!g944) & (!g1221) & (keyx36x)) + ((ld) & (g432) & (!g688) & (!g944) & (g1221) & (keyx36x)) + ((ld) & (g432) & (!g688) & (g944) & (!g1221) & (keyx36x)) + ((ld) & (g432) & (!g688) & (g944) & (g1221) & (keyx36x)) + ((ld) & (g432) & (g688) & (!g944) & (!g1221) & (keyx36x)) + ((ld) & (g432) & (g688) & (!g944) & (g1221) & (keyx36x)) + ((ld) & (g432) & (g688) & (g944) & (!g1221) & (keyx36x)) + ((ld) & (g432) & (g688) & (g944) & (g1221) & (keyx36x)));
	assign g1530 = (((!ld) & (!g439) & (!g695) & (!g951) & (g1228) & (!keyx37x)) + ((!ld) & (!g439) & (!g695) & (!g951) & (g1228) & (keyx37x)) + ((!ld) & (!g439) & (!g695) & (g951) & (!g1228) & (!keyx37x)) + ((!ld) & (!g439) & (!g695) & (g951) & (!g1228) & (keyx37x)) + ((!ld) & (!g439) & (g695) & (!g951) & (!g1228) & (!keyx37x)) + ((!ld) & (!g439) & (g695) & (!g951) & (!g1228) & (keyx37x)) + ((!ld) & (!g439) & (g695) & (g951) & (g1228) & (!keyx37x)) + ((!ld) & (!g439) & (g695) & (g951) & (g1228) & (keyx37x)) + ((!ld) & (g439) & (!g695) & (!g951) & (!g1228) & (!keyx37x)) + ((!ld) & (g439) & (!g695) & (!g951) & (!g1228) & (keyx37x)) + ((!ld) & (g439) & (!g695) & (g951) & (g1228) & (!keyx37x)) + ((!ld) & (g439) & (!g695) & (g951) & (g1228) & (keyx37x)) + ((!ld) & (g439) & (g695) & (!g951) & (g1228) & (!keyx37x)) + ((!ld) & (g439) & (g695) & (!g951) & (g1228) & (keyx37x)) + ((!ld) & (g439) & (g695) & (g951) & (!g1228) & (!keyx37x)) + ((!ld) & (g439) & (g695) & (g951) & (!g1228) & (keyx37x)) + ((ld) & (!g439) & (!g695) & (!g951) & (!g1228) & (keyx37x)) + ((ld) & (!g439) & (!g695) & (!g951) & (g1228) & (keyx37x)) + ((ld) & (!g439) & (!g695) & (g951) & (!g1228) & (keyx37x)) + ((ld) & (!g439) & (!g695) & (g951) & (g1228) & (keyx37x)) + ((ld) & (!g439) & (g695) & (!g951) & (!g1228) & (keyx37x)) + ((ld) & (!g439) & (g695) & (!g951) & (g1228) & (keyx37x)) + ((ld) & (!g439) & (g695) & (g951) & (!g1228) & (keyx37x)) + ((ld) & (!g439) & (g695) & (g951) & (g1228) & (keyx37x)) + ((ld) & (g439) & (!g695) & (!g951) & (!g1228) & (keyx37x)) + ((ld) & (g439) & (!g695) & (!g951) & (g1228) & (keyx37x)) + ((ld) & (g439) & (!g695) & (g951) & (!g1228) & (keyx37x)) + ((ld) & (g439) & (!g695) & (g951) & (g1228) & (keyx37x)) + ((ld) & (g439) & (g695) & (!g951) & (!g1228) & (keyx37x)) + ((ld) & (g439) & (g695) & (!g951) & (g1228) & (keyx37x)) + ((ld) & (g439) & (g695) & (g951) & (!g1228) & (keyx37x)) + ((ld) & (g439) & (g695) & (g951) & (g1228) & (keyx37x)));
	assign g1531 = (((!ld) & (!g446) & (!g702) & (!g958) & (g1235) & (!keyx38x)) + ((!ld) & (!g446) & (!g702) & (!g958) & (g1235) & (keyx38x)) + ((!ld) & (!g446) & (!g702) & (g958) & (!g1235) & (!keyx38x)) + ((!ld) & (!g446) & (!g702) & (g958) & (!g1235) & (keyx38x)) + ((!ld) & (!g446) & (g702) & (!g958) & (!g1235) & (!keyx38x)) + ((!ld) & (!g446) & (g702) & (!g958) & (!g1235) & (keyx38x)) + ((!ld) & (!g446) & (g702) & (g958) & (g1235) & (!keyx38x)) + ((!ld) & (!g446) & (g702) & (g958) & (g1235) & (keyx38x)) + ((!ld) & (g446) & (!g702) & (!g958) & (!g1235) & (!keyx38x)) + ((!ld) & (g446) & (!g702) & (!g958) & (!g1235) & (keyx38x)) + ((!ld) & (g446) & (!g702) & (g958) & (g1235) & (!keyx38x)) + ((!ld) & (g446) & (!g702) & (g958) & (g1235) & (keyx38x)) + ((!ld) & (g446) & (g702) & (!g958) & (g1235) & (!keyx38x)) + ((!ld) & (g446) & (g702) & (!g958) & (g1235) & (keyx38x)) + ((!ld) & (g446) & (g702) & (g958) & (!g1235) & (!keyx38x)) + ((!ld) & (g446) & (g702) & (g958) & (!g1235) & (keyx38x)) + ((ld) & (!g446) & (!g702) & (!g958) & (!g1235) & (keyx38x)) + ((ld) & (!g446) & (!g702) & (!g958) & (g1235) & (keyx38x)) + ((ld) & (!g446) & (!g702) & (g958) & (!g1235) & (keyx38x)) + ((ld) & (!g446) & (!g702) & (g958) & (g1235) & (keyx38x)) + ((ld) & (!g446) & (g702) & (!g958) & (!g1235) & (keyx38x)) + ((ld) & (!g446) & (g702) & (!g958) & (g1235) & (keyx38x)) + ((ld) & (!g446) & (g702) & (g958) & (!g1235) & (keyx38x)) + ((ld) & (!g446) & (g702) & (g958) & (g1235) & (keyx38x)) + ((ld) & (g446) & (!g702) & (!g958) & (!g1235) & (keyx38x)) + ((ld) & (g446) & (!g702) & (!g958) & (g1235) & (keyx38x)) + ((ld) & (g446) & (!g702) & (g958) & (!g1235) & (keyx38x)) + ((ld) & (g446) & (!g702) & (g958) & (g1235) & (keyx38x)) + ((ld) & (g446) & (g702) & (!g958) & (!g1235) & (keyx38x)) + ((ld) & (g446) & (g702) & (!g958) & (g1235) & (keyx38x)) + ((ld) & (g446) & (g702) & (g958) & (!g1235) & (keyx38x)) + ((ld) & (g446) & (g702) & (g958) & (g1235) & (keyx38x)));
	assign g1532 = (((!ld) & (!g453) & (!g709) & (!g965) & (g1242) & (!keyx39x)) + ((!ld) & (!g453) & (!g709) & (!g965) & (g1242) & (keyx39x)) + ((!ld) & (!g453) & (!g709) & (g965) & (!g1242) & (!keyx39x)) + ((!ld) & (!g453) & (!g709) & (g965) & (!g1242) & (keyx39x)) + ((!ld) & (!g453) & (g709) & (!g965) & (!g1242) & (!keyx39x)) + ((!ld) & (!g453) & (g709) & (!g965) & (!g1242) & (keyx39x)) + ((!ld) & (!g453) & (g709) & (g965) & (g1242) & (!keyx39x)) + ((!ld) & (!g453) & (g709) & (g965) & (g1242) & (keyx39x)) + ((!ld) & (g453) & (!g709) & (!g965) & (!g1242) & (!keyx39x)) + ((!ld) & (g453) & (!g709) & (!g965) & (!g1242) & (keyx39x)) + ((!ld) & (g453) & (!g709) & (g965) & (g1242) & (!keyx39x)) + ((!ld) & (g453) & (!g709) & (g965) & (g1242) & (keyx39x)) + ((!ld) & (g453) & (g709) & (!g965) & (g1242) & (!keyx39x)) + ((!ld) & (g453) & (g709) & (!g965) & (g1242) & (keyx39x)) + ((!ld) & (g453) & (g709) & (g965) & (!g1242) & (!keyx39x)) + ((!ld) & (g453) & (g709) & (g965) & (!g1242) & (keyx39x)) + ((ld) & (!g453) & (!g709) & (!g965) & (!g1242) & (keyx39x)) + ((ld) & (!g453) & (!g709) & (!g965) & (g1242) & (keyx39x)) + ((ld) & (!g453) & (!g709) & (g965) & (!g1242) & (keyx39x)) + ((ld) & (!g453) & (!g709) & (g965) & (g1242) & (keyx39x)) + ((ld) & (!g453) & (g709) & (!g965) & (!g1242) & (keyx39x)) + ((ld) & (!g453) & (g709) & (!g965) & (g1242) & (keyx39x)) + ((ld) & (!g453) & (g709) & (g965) & (!g1242) & (keyx39x)) + ((ld) & (!g453) & (g709) & (g965) & (g1242) & (keyx39x)) + ((ld) & (g453) & (!g709) & (!g965) & (!g1242) & (keyx39x)) + ((ld) & (g453) & (!g709) & (!g965) & (g1242) & (keyx39x)) + ((ld) & (g453) & (!g709) & (g965) & (!g1242) & (keyx39x)) + ((ld) & (g453) & (!g709) & (g965) & (g1242) & (keyx39x)) + ((ld) & (g453) & (g709) & (!g965) & (!g1242) & (keyx39x)) + ((ld) & (g453) & (g709) & (!g965) & (g1242) & (keyx39x)) + ((ld) & (g453) & (g709) & (g965) & (!g1242) & (keyx39x)) + ((ld) & (g453) & (g709) & (g965) & (g1242) & (keyx39x)));
	assign g2122 = (((!ld) & (!text_inx104x) & (sk[110]) & (g1533)) + ((!ld) & (text_inx104x) & (!sk[110]) & (!g1533)) + ((!ld) & (text_inx104x) & (!sk[110]) & (g1533)) + ((!ld) & (text_inx104x) & (sk[110]) & (g1533)) + ((ld) & (!text_inx104x) & (!sk[110]) & (g1533)) + ((ld) & (text_inx104x) & (!sk[110]) & (!g1533)) + ((ld) & (text_inx104x) & (!sk[110]) & (g1533)) + ((ld) & (text_inx104x) & (sk[110]) & (!g1533)) + ((ld) & (text_inx104x) & (sk[110]) & (g1533)));
	assign g1534 = (((!g915) & (!g980) & (!sk[111]) & (g1043) & (!g1107)) + ((!g915) & (!g980) & (!sk[111]) & (g1043) & (g1107)) + ((!g915) & (!g980) & (sk[111]) & (!g1043) & (g1107)) + ((!g915) & (!g980) & (sk[111]) & (g1043) & (!g1107)) + ((!g915) & (g980) & (!sk[111]) & (!g1043) & (!g1107)) + ((!g915) & (g980) & (!sk[111]) & (!g1043) & (g1107)) + ((!g915) & (g980) & (!sk[111]) & (g1043) & (!g1107)) + ((!g915) & (g980) & (!sk[111]) & (g1043) & (g1107)) + ((!g915) & (g980) & (sk[111]) & (!g1043) & (!g1107)) + ((!g915) & (g980) & (sk[111]) & (g1043) & (g1107)) + ((g915) & (!g980) & (!sk[111]) & (g1043) & (!g1107)) + ((g915) & (!g980) & (!sk[111]) & (g1043) & (g1107)) + ((g915) & (!g980) & (sk[111]) & (!g1043) & (!g1107)) + ((g915) & (!g980) & (sk[111]) & (g1043) & (g1107)) + ((g915) & (g980) & (!sk[111]) & (!g1043) & (!g1107)) + ((g915) & (g980) & (!sk[111]) & (!g1043) & (g1107)) + ((g915) & (g980) & (!sk[111]) & (g1043) & (!g1107)) + ((g915) & (g980) & (!sk[111]) & (g1043) & (g1107)) + ((g915) & (g980) & (sk[111]) & (!g1043) & (g1107)) + ((g915) & (g980) & (sk[111]) & (g1043) & (!g1107)));
	assign g1535 = (((!g964) & (!g980) & (!g1028) & (!g1163) & (!g1533) & (g1534)) + ((!g964) & (!g980) & (!g1028) & (!g1163) & (g1533) & (g1534)) + ((!g964) & (!g980) & (!g1028) & (g1163) & (g1533) & (!g1534)) + ((!g964) & (!g980) & (!g1028) & (g1163) & (g1533) & (g1534)) + ((!g964) & (!g980) & (g1028) & (!g1163) & (!g1533) & (!g1534)) + ((!g964) & (!g980) & (g1028) & (!g1163) & (g1533) & (!g1534)) + ((!g964) & (!g980) & (g1028) & (g1163) & (g1533) & (!g1534)) + ((!g964) & (!g980) & (g1028) & (g1163) & (g1533) & (g1534)) + ((!g964) & (g980) & (!g1028) & (!g1163) & (!g1533) & (g1534)) + ((!g964) & (g980) & (!g1028) & (!g1163) & (g1533) & (g1534)) + ((!g964) & (g980) & (!g1028) & (g1163) & (!g1533) & (!g1534)) + ((!g964) & (g980) & (!g1028) & (g1163) & (!g1533) & (g1534)) + ((!g964) & (g980) & (g1028) & (!g1163) & (!g1533) & (!g1534)) + ((!g964) & (g980) & (g1028) & (!g1163) & (g1533) & (!g1534)) + ((!g964) & (g980) & (g1028) & (g1163) & (!g1533) & (!g1534)) + ((!g964) & (g980) & (g1028) & (g1163) & (!g1533) & (g1534)) + ((g964) & (!g980) & (!g1028) & (!g1163) & (!g1533) & (!g1534)) + ((g964) & (!g980) & (!g1028) & (!g1163) & (g1533) & (!g1534)) + ((g964) & (!g980) & (!g1028) & (g1163) & (g1533) & (!g1534)) + ((g964) & (!g980) & (!g1028) & (g1163) & (g1533) & (g1534)) + ((g964) & (!g980) & (g1028) & (!g1163) & (!g1533) & (g1534)) + ((g964) & (!g980) & (g1028) & (!g1163) & (g1533) & (g1534)) + ((g964) & (!g980) & (g1028) & (g1163) & (g1533) & (!g1534)) + ((g964) & (!g980) & (g1028) & (g1163) & (g1533) & (g1534)) + ((g964) & (g980) & (!g1028) & (!g1163) & (!g1533) & (!g1534)) + ((g964) & (g980) & (!g1028) & (!g1163) & (g1533) & (!g1534)) + ((g964) & (g980) & (!g1028) & (g1163) & (!g1533) & (!g1534)) + ((g964) & (g980) & (!g1028) & (g1163) & (!g1533) & (g1534)) + ((g964) & (g980) & (g1028) & (!g1163) & (!g1533) & (g1534)) + ((g964) & (g980) & (g1028) & (!g1163) & (g1533) & (g1534)) + ((g964) & (g980) & (g1028) & (g1163) & (!g1533) & (!g1534)) + ((g964) & (g980) & (g1028) & (g1163) & (!g1533) & (g1534)));
	assign g2123 = (((!ld) & (!text_inx105x) & (sk[113]) & (g1536)) + ((!ld) & (text_inx105x) & (!sk[113]) & (!g1536)) + ((!ld) & (text_inx105x) & (!sk[113]) & (g1536)) + ((!ld) & (text_inx105x) & (sk[113]) & (g1536)) + ((ld) & (!text_inx105x) & (!sk[113]) & (g1536)) + ((ld) & (text_inx105x) & (!sk[113]) & (!g1536)) + ((ld) & (text_inx105x) & (!sk[113]) & (g1536)) + ((ld) & (text_inx105x) & (sk[113]) & (!g1536)) + ((ld) & (text_inx105x) & (sk[113]) & (g1536)));
	assign g1537 = (((!g987) & (!sk[114]) & (g1536)) + ((!g987) & (sk[114]) & (g1536)) + ((g987) & (!sk[114]) & (g1536)) + ((g987) & (sk[114]) & (!g1536)));
	assign g1538 = (((!g922) & (!g987) & (!g1050) & (sk[115]) & (g1114)) + ((!g922) & (!g987) & (g1050) & (!sk[115]) & (!g1114)) + ((!g922) & (!g987) & (g1050) & (!sk[115]) & (g1114)) + ((!g922) & (!g987) & (g1050) & (sk[115]) & (!g1114)) + ((!g922) & (g987) & (!g1050) & (!sk[115]) & (!g1114)) + ((!g922) & (g987) & (!g1050) & (!sk[115]) & (g1114)) + ((!g922) & (g987) & (!g1050) & (sk[115]) & (!g1114)) + ((!g922) & (g987) & (g1050) & (!sk[115]) & (!g1114)) + ((!g922) & (g987) & (g1050) & (!sk[115]) & (g1114)) + ((!g922) & (g987) & (g1050) & (sk[115]) & (g1114)) + ((g922) & (!g987) & (!g1050) & (sk[115]) & (!g1114)) + ((g922) & (!g987) & (g1050) & (!sk[115]) & (!g1114)) + ((g922) & (!g987) & (g1050) & (!sk[115]) & (g1114)) + ((g922) & (!g987) & (g1050) & (sk[115]) & (g1114)) + ((g922) & (g987) & (!g1050) & (!sk[115]) & (!g1114)) + ((g922) & (g987) & (!g1050) & (!sk[115]) & (g1114)) + ((g922) & (g987) & (!g1050) & (sk[115]) & (g1114)) + ((g922) & (g987) & (g1050) & (!sk[115]) & (!g1114)) + ((g922) & (g987) & (g1050) & (!sk[115]) & (g1114)) + ((g922) & (g987) & (g1050) & (sk[115]) & (!g1114)));
	assign g1539 = (((!g964) & (!g1028) & (!g1163) & (!g1330) & (!g1537) & (g1538)) + ((!g964) & (!g1028) & (!g1163) & (!g1330) & (g1537) & (g1538)) + ((!g964) & (!g1028) & (!g1163) & (g1330) & (!g1537) & (!g1538)) + ((!g964) & (!g1028) & (!g1163) & (g1330) & (g1537) & (!g1538)) + ((!g964) & (!g1028) & (g1163) & (!g1330) & (g1537) & (!g1538)) + ((!g964) & (!g1028) & (g1163) & (!g1330) & (g1537) & (g1538)) + ((!g964) & (!g1028) & (g1163) & (g1330) & (g1537) & (!g1538)) + ((!g964) & (!g1028) & (g1163) & (g1330) & (g1537) & (g1538)) + ((!g964) & (g1028) & (!g1163) & (!g1330) & (!g1537) & (!g1538)) + ((!g964) & (g1028) & (!g1163) & (!g1330) & (g1537) & (!g1538)) + ((!g964) & (g1028) & (!g1163) & (g1330) & (!g1537) & (g1538)) + ((!g964) & (g1028) & (!g1163) & (g1330) & (g1537) & (g1538)) + ((!g964) & (g1028) & (g1163) & (!g1330) & (g1537) & (!g1538)) + ((!g964) & (g1028) & (g1163) & (!g1330) & (g1537) & (g1538)) + ((!g964) & (g1028) & (g1163) & (g1330) & (g1537) & (!g1538)) + ((!g964) & (g1028) & (g1163) & (g1330) & (g1537) & (g1538)) + ((g964) & (!g1028) & (!g1163) & (!g1330) & (!g1537) & (!g1538)) + ((g964) & (!g1028) & (!g1163) & (!g1330) & (g1537) & (!g1538)) + ((g964) & (!g1028) & (!g1163) & (g1330) & (!g1537) & (g1538)) + ((g964) & (!g1028) & (!g1163) & (g1330) & (g1537) & (g1538)) + ((g964) & (!g1028) & (g1163) & (!g1330) & (g1537) & (!g1538)) + ((g964) & (!g1028) & (g1163) & (!g1330) & (g1537) & (g1538)) + ((g964) & (!g1028) & (g1163) & (g1330) & (g1537) & (!g1538)) + ((g964) & (!g1028) & (g1163) & (g1330) & (g1537) & (g1538)) + ((g964) & (g1028) & (!g1163) & (!g1330) & (!g1537) & (g1538)) + ((g964) & (g1028) & (!g1163) & (!g1330) & (g1537) & (g1538)) + ((g964) & (g1028) & (!g1163) & (g1330) & (!g1537) & (!g1538)) + ((g964) & (g1028) & (!g1163) & (g1330) & (g1537) & (!g1538)) + ((g964) & (g1028) & (g1163) & (!g1330) & (g1537) & (!g1538)) + ((g964) & (g1028) & (g1163) & (!g1330) & (g1537) & (g1538)) + ((g964) & (g1028) & (g1163) & (g1330) & (g1537) & (!g1538)) + ((g964) & (g1028) & (g1163) & (g1330) & (g1537) & (g1538)));
	assign g2124 = (((!ld) & (!text_inx106x) & (sk[117]) & (g1540)) + ((!ld) & (text_inx106x) & (!sk[117]) & (!g1540)) + ((!ld) & (text_inx106x) & (!sk[117]) & (g1540)) + ((!ld) & (text_inx106x) & (sk[117]) & (g1540)) + ((ld) & (!text_inx106x) & (!sk[117]) & (g1540)) + ((ld) & (text_inx106x) & (!sk[117]) & (!g1540)) + ((ld) & (text_inx106x) & (!sk[117]) & (g1540)) + ((ld) & (text_inx106x) & (sk[117]) & (!g1540)) + ((ld) & (text_inx106x) & (sk[117]) & (g1540)));
	assign g1541 = (((!g922) & (!sk[118]) & (g1057) & (!g1121)) + ((!g922) & (!sk[118]) & (g1057) & (g1121)) + ((!g922) & (sk[118]) & (!g1057) & (g1121)) + ((!g922) & (sk[118]) & (g1057) & (!g1121)) + ((g922) & (!sk[118]) & (!g1057) & (g1121)) + ((g922) & (!sk[118]) & (g1057) & (!g1121)) + ((g922) & (!sk[118]) & (g1057) & (g1121)) + ((g922) & (sk[118]) & (!g1057) & (!g1121)) + ((g922) & (sk[118]) & (g1057) & (g1121)));
	assign g1542 = (((!g929) & (!g986) & (!g994) & (!g1163) & (!g1540) & (g1541)) + ((!g929) & (!g986) & (!g994) & (!g1163) & (g1540) & (g1541)) + ((!g929) & (!g986) & (!g994) & (g1163) & (g1540) & (!g1541)) + ((!g929) & (!g986) & (!g994) & (g1163) & (g1540) & (g1541)) + ((!g929) & (!g986) & (g994) & (!g1163) & (!g1540) & (!g1541)) + ((!g929) & (!g986) & (g994) & (!g1163) & (g1540) & (!g1541)) + ((!g929) & (!g986) & (g994) & (g1163) & (!g1540) & (!g1541)) + ((!g929) & (!g986) & (g994) & (g1163) & (!g1540) & (g1541)) + ((!g929) & (g986) & (!g994) & (!g1163) & (!g1540) & (!g1541)) + ((!g929) & (g986) & (!g994) & (!g1163) & (g1540) & (!g1541)) + ((!g929) & (g986) & (!g994) & (g1163) & (g1540) & (!g1541)) + ((!g929) & (g986) & (!g994) & (g1163) & (g1540) & (g1541)) + ((!g929) & (g986) & (g994) & (!g1163) & (!g1540) & (g1541)) + ((!g929) & (g986) & (g994) & (!g1163) & (g1540) & (g1541)) + ((!g929) & (g986) & (g994) & (g1163) & (!g1540) & (!g1541)) + ((!g929) & (g986) & (g994) & (g1163) & (!g1540) & (g1541)) + ((g929) & (!g986) & (!g994) & (!g1163) & (!g1540) & (!g1541)) + ((g929) & (!g986) & (!g994) & (!g1163) & (g1540) & (!g1541)) + ((g929) & (!g986) & (!g994) & (g1163) & (g1540) & (!g1541)) + ((g929) & (!g986) & (!g994) & (g1163) & (g1540) & (g1541)) + ((g929) & (!g986) & (g994) & (!g1163) & (!g1540) & (g1541)) + ((g929) & (!g986) & (g994) & (!g1163) & (g1540) & (g1541)) + ((g929) & (!g986) & (g994) & (g1163) & (!g1540) & (!g1541)) + ((g929) & (!g986) & (g994) & (g1163) & (!g1540) & (g1541)) + ((g929) & (g986) & (!g994) & (!g1163) & (!g1540) & (g1541)) + ((g929) & (g986) & (!g994) & (!g1163) & (g1540) & (g1541)) + ((g929) & (g986) & (!g994) & (g1163) & (g1540) & (!g1541)) + ((g929) & (g986) & (!g994) & (g1163) & (g1540) & (g1541)) + ((g929) & (g986) & (g994) & (!g1163) & (!g1540) & (!g1541)) + ((g929) & (g986) & (g994) & (!g1163) & (g1540) & (!g1541)) + ((g929) & (g986) & (g994) & (g1163) & (!g1540) & (!g1541)) + ((g929) & (g986) & (g994) & (g1163) & (!g1540) & (g1541)));
	assign g2125 = (((!ld) & (!sk[120]) & (text_inx107x) & (!g1543)) + ((!ld) & (!sk[120]) & (text_inx107x) & (g1543)) + ((!ld) & (sk[120]) & (!text_inx107x) & (g1543)) + ((!ld) & (sk[120]) & (text_inx107x) & (g1543)) + ((ld) & (!sk[120]) & (!text_inx107x) & (g1543)) + ((ld) & (!sk[120]) & (text_inx107x) & (!g1543)) + ((ld) & (!sk[120]) & (text_inx107x) & (g1543)) + ((ld) & (sk[120]) & (text_inx107x) & (!g1543)) + ((ld) & (sk[120]) & (text_inx107x) & (g1543)));
	assign g1544 = (((!g936) & (!sk[121]) & (g964) & (!g1028)) + ((!g936) & (!sk[121]) & (g964) & (g1028)) + ((!g936) & (sk[121]) & (!g964) & (g1028)) + ((!g936) & (sk[121]) & (g964) & (!g1028)) + ((g936) & (!sk[121]) & (!g964) & (g1028)) + ((g936) & (!sk[121]) & (g964) & (!g1028)) + ((g936) & (!sk[121]) & (g964) & (g1028)) + ((g936) & (sk[121]) & (!g964) & (!g1028)) + ((g936) & (sk[121]) & (g964) & (g1028)));
	assign g1545 = (((!sk[122]) & (!g929) & (g993) & (!g1001) & (!g1064) & (!g1128)) + ((!sk[122]) & (!g929) & (g993) & (!g1001) & (!g1064) & (g1128)) + ((!sk[122]) & (!g929) & (g993) & (!g1001) & (g1064) & (!g1128)) + ((!sk[122]) & (!g929) & (g993) & (!g1001) & (g1064) & (g1128)) + ((!sk[122]) & (!g929) & (g993) & (g1001) & (!g1064) & (!g1128)) + ((!sk[122]) & (!g929) & (g993) & (g1001) & (!g1064) & (g1128)) + ((!sk[122]) & (!g929) & (g993) & (g1001) & (g1064) & (!g1128)) + ((!sk[122]) & (!g929) & (g993) & (g1001) & (g1064) & (g1128)) + ((!sk[122]) & (g929) & (!g993) & (!g1001) & (!g1064) & (!g1128)) + ((!sk[122]) & (g929) & (!g993) & (!g1001) & (!g1064) & (g1128)) + ((!sk[122]) & (g929) & (!g993) & (!g1001) & (g1064) & (!g1128)) + ((!sk[122]) & (g929) & (!g993) & (!g1001) & (g1064) & (g1128)) + ((!sk[122]) & (g929) & (!g993) & (g1001) & (!g1064) & (!g1128)) + ((!sk[122]) & (g929) & (!g993) & (g1001) & (!g1064) & (g1128)) + ((!sk[122]) & (g929) & (!g993) & (g1001) & (g1064) & (!g1128)) + ((!sk[122]) & (g929) & (!g993) & (g1001) & (g1064) & (g1128)) + ((!sk[122]) & (g929) & (g993) & (!g1001) & (!g1064) & (!g1128)) + ((!sk[122]) & (g929) & (g993) & (!g1001) & (!g1064) & (g1128)) + ((!sk[122]) & (g929) & (g993) & (!g1001) & (g1064) & (!g1128)) + ((!sk[122]) & (g929) & (g993) & (!g1001) & (g1064) & (g1128)) + ((!sk[122]) & (g929) & (g993) & (g1001) & (!g1064) & (!g1128)) + ((!sk[122]) & (g929) & (g993) & (g1001) & (!g1064) & (g1128)) + ((!sk[122]) & (g929) & (g993) & (g1001) & (g1064) & (!g1128)) + ((!sk[122]) & (g929) & (g993) & (g1001) & (g1064) & (g1128)) + ((sk[122]) & (!g929) & (!g993) & (!g1001) & (!g1064) & (g1128)) + ((sk[122]) & (!g929) & (!g993) & (!g1001) & (g1064) & (!g1128)) + ((sk[122]) & (!g929) & (!g993) & (g1001) & (!g1064) & (!g1128)) + ((sk[122]) & (!g929) & (!g993) & (g1001) & (g1064) & (g1128)) + ((sk[122]) & (!g929) & (g993) & (!g1001) & (!g1064) & (!g1128)) + ((sk[122]) & (!g929) & (g993) & (!g1001) & (g1064) & (g1128)) + ((sk[122]) & (!g929) & (g993) & (g1001) & (!g1064) & (g1128)) + ((sk[122]) & (!g929) & (g993) & (g1001) & (g1064) & (!g1128)) + ((sk[122]) & (g929) & (!g993) & (!g1001) & (!g1064) & (!g1128)) + ((sk[122]) & (g929) & (!g993) & (!g1001) & (g1064) & (g1128)) + ((sk[122]) & (g929) & (!g993) & (g1001) & (!g1064) & (g1128)) + ((sk[122]) & (g929) & (!g993) & (g1001) & (g1064) & (!g1128)) + ((sk[122]) & (g929) & (g993) & (!g1001) & (!g1064) & (g1128)) + ((sk[122]) & (g929) & (g993) & (!g1001) & (g1064) & (!g1128)) + ((sk[122]) & (g929) & (g993) & (g1001) & (!g1064) & (!g1128)) + ((sk[122]) & (g929) & (g993) & (g1001) & (g1064) & (g1128)));
	assign g1546 = (((!sk[123]) & (!g1001) & (g1163) & (!g1543) & (!g1544) & (!g1545)) + ((!sk[123]) & (!g1001) & (g1163) & (!g1543) & (!g1544) & (g1545)) + ((!sk[123]) & (!g1001) & (g1163) & (!g1543) & (g1544) & (!g1545)) + ((!sk[123]) & (!g1001) & (g1163) & (!g1543) & (g1544) & (g1545)) + ((!sk[123]) & (!g1001) & (g1163) & (g1543) & (!g1544) & (!g1545)) + ((!sk[123]) & (!g1001) & (g1163) & (g1543) & (!g1544) & (g1545)) + ((!sk[123]) & (!g1001) & (g1163) & (g1543) & (g1544) & (!g1545)) + ((!sk[123]) & (!g1001) & (g1163) & (g1543) & (g1544) & (g1545)) + ((!sk[123]) & (g1001) & (!g1163) & (!g1543) & (!g1544) & (!g1545)) + ((!sk[123]) & (g1001) & (!g1163) & (!g1543) & (!g1544) & (g1545)) + ((!sk[123]) & (g1001) & (!g1163) & (!g1543) & (g1544) & (!g1545)) + ((!sk[123]) & (g1001) & (!g1163) & (!g1543) & (g1544) & (g1545)) + ((!sk[123]) & (g1001) & (!g1163) & (g1543) & (!g1544) & (!g1545)) + ((!sk[123]) & (g1001) & (!g1163) & (g1543) & (!g1544) & (g1545)) + ((!sk[123]) & (g1001) & (!g1163) & (g1543) & (g1544) & (!g1545)) + ((!sk[123]) & (g1001) & (!g1163) & (g1543) & (g1544) & (g1545)) + ((!sk[123]) & (g1001) & (g1163) & (!g1543) & (!g1544) & (!g1545)) + ((!sk[123]) & (g1001) & (g1163) & (!g1543) & (!g1544) & (g1545)) + ((!sk[123]) & (g1001) & (g1163) & (!g1543) & (g1544) & (!g1545)) + ((!sk[123]) & (g1001) & (g1163) & (!g1543) & (g1544) & (g1545)) + ((!sk[123]) & (g1001) & (g1163) & (g1543) & (!g1544) & (!g1545)) + ((!sk[123]) & (g1001) & (g1163) & (g1543) & (!g1544) & (g1545)) + ((!sk[123]) & (g1001) & (g1163) & (g1543) & (g1544) & (!g1545)) + ((!sk[123]) & (g1001) & (g1163) & (g1543) & (g1544) & (g1545)) + ((sk[123]) & (!g1001) & (!g1163) & (!g1543) & (!g1544) & (g1545)) + ((sk[123]) & (!g1001) & (!g1163) & (!g1543) & (g1544) & (!g1545)) + ((sk[123]) & (!g1001) & (!g1163) & (g1543) & (!g1544) & (g1545)) + ((sk[123]) & (!g1001) & (!g1163) & (g1543) & (g1544) & (!g1545)) + ((sk[123]) & (!g1001) & (g1163) & (g1543) & (!g1544) & (!g1545)) + ((sk[123]) & (!g1001) & (g1163) & (g1543) & (!g1544) & (g1545)) + ((sk[123]) & (!g1001) & (g1163) & (g1543) & (g1544) & (!g1545)) + ((sk[123]) & (!g1001) & (g1163) & (g1543) & (g1544) & (g1545)) + ((sk[123]) & (g1001) & (!g1163) & (!g1543) & (!g1544) & (g1545)) + ((sk[123]) & (g1001) & (!g1163) & (!g1543) & (g1544) & (!g1545)) + ((sk[123]) & (g1001) & (!g1163) & (g1543) & (!g1544) & (g1545)) + ((sk[123]) & (g1001) & (!g1163) & (g1543) & (g1544) & (!g1545)) + ((sk[123]) & (g1001) & (g1163) & (!g1543) & (!g1544) & (!g1545)) + ((sk[123]) & (g1001) & (g1163) & (!g1543) & (!g1544) & (g1545)) + ((sk[123]) & (g1001) & (g1163) & (!g1543) & (g1544) & (!g1545)) + ((sk[123]) & (g1001) & (g1163) & (!g1543) & (g1544) & (g1545)));
	assign g2126 = (((!ld) & (!sk[124]) & (text_inx110x) & (!g1547)) + ((!ld) & (!sk[124]) & (text_inx110x) & (g1547)) + ((!ld) & (sk[124]) & (!text_inx110x) & (g1547)) + ((!ld) & (sk[124]) & (text_inx110x) & (g1547)) + ((ld) & (!sk[124]) & (!text_inx110x) & (g1547)) + ((ld) & (!sk[124]) & (text_inx110x) & (!g1547)) + ((ld) & (!sk[124]) & (text_inx110x) & (g1547)) + ((ld) & (sk[124]) & (text_inx110x) & (!g1547)) + ((ld) & (sk[124]) & (text_inx110x) & (g1547)));
	assign g1548 = (((!sk[125]) & (!g950) & (g1085) & (!g1149)) + ((!sk[125]) & (!g950) & (g1085) & (g1149)) + ((!sk[125]) & (g950) & (!g1085) & (g1149)) + ((!sk[125]) & (g950) & (g1085) & (!g1149)) + ((!sk[125]) & (g950) & (g1085) & (g1149)) + ((sk[125]) & (!g950) & (!g1085) & (g1149)) + ((sk[125]) & (!g950) & (g1085) & (!g1149)) + ((sk[125]) & (g950) & (!g1085) & (!g1149)) + ((sk[125]) & (g950) & (g1085) & (g1149)));
	assign g1549 = (((!g957) & (!g1014) & (!g1022) & (!g1163) & (!g1547) & (g1548)) + ((!g957) & (!g1014) & (!g1022) & (!g1163) & (g1547) & (g1548)) + ((!g957) & (!g1014) & (!g1022) & (g1163) & (g1547) & (!g1548)) + ((!g957) & (!g1014) & (!g1022) & (g1163) & (g1547) & (g1548)) + ((!g957) & (!g1014) & (g1022) & (!g1163) & (!g1547) & (!g1548)) + ((!g957) & (!g1014) & (g1022) & (!g1163) & (g1547) & (!g1548)) + ((!g957) & (!g1014) & (g1022) & (g1163) & (!g1547) & (!g1548)) + ((!g957) & (!g1014) & (g1022) & (g1163) & (!g1547) & (g1548)) + ((!g957) & (g1014) & (!g1022) & (!g1163) & (!g1547) & (!g1548)) + ((!g957) & (g1014) & (!g1022) & (!g1163) & (g1547) & (!g1548)) + ((!g957) & (g1014) & (!g1022) & (g1163) & (g1547) & (!g1548)) + ((!g957) & (g1014) & (!g1022) & (g1163) & (g1547) & (g1548)) + ((!g957) & (g1014) & (g1022) & (!g1163) & (!g1547) & (g1548)) + ((!g957) & (g1014) & (g1022) & (!g1163) & (g1547) & (g1548)) + ((!g957) & (g1014) & (g1022) & (g1163) & (!g1547) & (!g1548)) + ((!g957) & (g1014) & (g1022) & (g1163) & (!g1547) & (g1548)) + ((g957) & (!g1014) & (!g1022) & (!g1163) & (!g1547) & (!g1548)) + ((g957) & (!g1014) & (!g1022) & (!g1163) & (g1547) & (!g1548)) + ((g957) & (!g1014) & (!g1022) & (g1163) & (g1547) & (!g1548)) + ((g957) & (!g1014) & (!g1022) & (g1163) & (g1547) & (g1548)) + ((g957) & (!g1014) & (g1022) & (!g1163) & (!g1547) & (g1548)) + ((g957) & (!g1014) & (g1022) & (!g1163) & (g1547) & (g1548)) + ((g957) & (!g1014) & (g1022) & (g1163) & (!g1547) & (!g1548)) + ((g957) & (!g1014) & (g1022) & (g1163) & (!g1547) & (g1548)) + ((g957) & (g1014) & (!g1022) & (!g1163) & (!g1547) & (g1548)) + ((g957) & (g1014) & (!g1022) & (!g1163) & (g1547) & (g1548)) + ((g957) & (g1014) & (!g1022) & (g1163) & (g1547) & (!g1548)) + ((g957) & (g1014) & (!g1022) & (g1163) & (g1547) & (g1548)) + ((g957) & (g1014) & (g1022) & (!g1163) & (!g1547) & (!g1548)) + ((g957) & (g1014) & (g1022) & (!g1163) & (g1547) & (!g1548)) + ((g957) & (g1014) & (g1022) & (g1163) & (!g1547) & (!g1548)) + ((g957) & (g1014) & (g1022) & (g1163) & (!g1547) & (g1548)));
	assign g2127 = (((!ld) & (!sk[127]) & (text_inx109x) & (!g1550)) + ((!ld) & (!sk[127]) & (text_inx109x) & (g1550)) + ((!ld) & (sk[127]) & (!text_inx109x) & (g1550)) + ((!ld) & (sk[127]) & (text_inx109x) & (g1550)) + ((ld) & (!sk[127]) & (!text_inx109x) & (g1550)) + ((ld) & (!sk[127]) & (text_inx109x) & (!g1550)) + ((ld) & (!sk[127]) & (text_inx109x) & (g1550)) + ((ld) & (sk[127]) & (text_inx109x) & (!g1550)) + ((ld) & (sk[127]) & (text_inx109x) & (g1550)));
	assign g1551 = (((!g943) & (!sk[0]) & (g1078) & (!g1142)) + ((!g943) & (!sk[0]) & (g1078) & (g1142)) + ((!g943) & (sk[0]) & (!g1078) & (g1142)) + ((!g943) & (sk[0]) & (g1078) & (!g1142)) + ((g943) & (!sk[0]) & (!g1078) & (g1142)) + ((g943) & (!sk[0]) & (g1078) & (!g1142)) + ((g943) & (!sk[0]) & (g1078) & (g1142)) + ((g943) & (sk[0]) & (!g1078) & (!g1142)) + ((g943) & (sk[0]) & (g1078) & (g1142)));
	assign g1552 = (((!g950) & (!g1007) & (!g1015) & (!g1163) & (!g1550) & (g1551)) + ((!g950) & (!g1007) & (!g1015) & (!g1163) & (g1550) & (g1551)) + ((!g950) & (!g1007) & (!g1015) & (g1163) & (g1550) & (!g1551)) + ((!g950) & (!g1007) & (!g1015) & (g1163) & (g1550) & (g1551)) + ((!g950) & (!g1007) & (g1015) & (!g1163) & (!g1550) & (!g1551)) + ((!g950) & (!g1007) & (g1015) & (!g1163) & (g1550) & (!g1551)) + ((!g950) & (!g1007) & (g1015) & (g1163) & (!g1550) & (!g1551)) + ((!g950) & (!g1007) & (g1015) & (g1163) & (!g1550) & (g1551)) + ((!g950) & (g1007) & (!g1015) & (!g1163) & (!g1550) & (!g1551)) + ((!g950) & (g1007) & (!g1015) & (!g1163) & (g1550) & (!g1551)) + ((!g950) & (g1007) & (!g1015) & (g1163) & (g1550) & (!g1551)) + ((!g950) & (g1007) & (!g1015) & (g1163) & (g1550) & (g1551)) + ((!g950) & (g1007) & (g1015) & (!g1163) & (!g1550) & (g1551)) + ((!g950) & (g1007) & (g1015) & (!g1163) & (g1550) & (g1551)) + ((!g950) & (g1007) & (g1015) & (g1163) & (!g1550) & (!g1551)) + ((!g950) & (g1007) & (g1015) & (g1163) & (!g1550) & (g1551)) + ((g950) & (!g1007) & (!g1015) & (!g1163) & (!g1550) & (!g1551)) + ((g950) & (!g1007) & (!g1015) & (!g1163) & (g1550) & (!g1551)) + ((g950) & (!g1007) & (!g1015) & (g1163) & (g1550) & (!g1551)) + ((g950) & (!g1007) & (!g1015) & (g1163) & (g1550) & (g1551)) + ((g950) & (!g1007) & (g1015) & (!g1163) & (!g1550) & (g1551)) + ((g950) & (!g1007) & (g1015) & (!g1163) & (g1550) & (g1551)) + ((g950) & (!g1007) & (g1015) & (g1163) & (!g1550) & (!g1551)) + ((g950) & (!g1007) & (g1015) & (g1163) & (!g1550) & (g1551)) + ((g950) & (g1007) & (!g1015) & (!g1163) & (!g1550) & (g1551)) + ((g950) & (g1007) & (!g1015) & (!g1163) & (g1550) & (g1551)) + ((g950) & (g1007) & (!g1015) & (g1163) & (g1550) & (!g1551)) + ((g950) & (g1007) & (!g1015) & (g1163) & (g1550) & (g1551)) + ((g950) & (g1007) & (g1015) & (!g1163) & (!g1550) & (!g1551)) + ((g950) & (g1007) & (g1015) & (!g1163) & (g1550) & (!g1551)) + ((g950) & (g1007) & (g1015) & (g1163) & (!g1550) & (!g1551)) + ((g950) & (g1007) & (g1015) & (g1163) & (!g1550) & (g1551)));
	assign g2128 = (((!sk[2]) & (!ld) & (text_inx108x) & (!g1553)) + ((!sk[2]) & (!ld) & (text_inx108x) & (g1553)) + ((!sk[2]) & (ld) & (!text_inx108x) & (g1553)) + ((!sk[2]) & (ld) & (text_inx108x) & (!g1553)) + ((!sk[2]) & (ld) & (text_inx108x) & (g1553)) + ((sk[2]) & (!ld) & (!text_inx108x) & (g1553)) + ((sk[2]) & (!ld) & (text_inx108x) & (g1553)) + ((sk[2]) & (ld) & (text_inx108x) & (!g1553)) + ((sk[2]) & (ld) & (text_inx108x) & (g1553)));
	assign g1554 = (((!g1008) & (!g1071) & (!g1163) & (!g1348) & (g1544) & (!g1553)) + ((!g1008) & (!g1071) & (!g1163) & (!g1348) & (g1544) & (g1553)) + ((!g1008) & (!g1071) & (!g1163) & (g1348) & (!g1544) & (!g1553)) + ((!g1008) & (!g1071) & (!g1163) & (g1348) & (!g1544) & (g1553)) + ((!g1008) & (!g1071) & (g1163) & (!g1348) & (!g1544) & (g1553)) + ((!g1008) & (!g1071) & (g1163) & (!g1348) & (g1544) & (g1553)) + ((!g1008) & (!g1071) & (g1163) & (g1348) & (!g1544) & (g1553)) + ((!g1008) & (!g1071) & (g1163) & (g1348) & (g1544) & (g1553)) + ((!g1008) & (g1071) & (!g1163) & (!g1348) & (!g1544) & (!g1553)) + ((!g1008) & (g1071) & (!g1163) & (!g1348) & (!g1544) & (g1553)) + ((!g1008) & (g1071) & (!g1163) & (g1348) & (g1544) & (!g1553)) + ((!g1008) & (g1071) & (!g1163) & (g1348) & (g1544) & (g1553)) + ((!g1008) & (g1071) & (g1163) & (!g1348) & (!g1544) & (g1553)) + ((!g1008) & (g1071) & (g1163) & (!g1348) & (g1544) & (g1553)) + ((!g1008) & (g1071) & (g1163) & (g1348) & (!g1544) & (g1553)) + ((!g1008) & (g1071) & (g1163) & (g1348) & (g1544) & (g1553)) + ((g1008) & (!g1071) & (!g1163) & (!g1348) & (!g1544) & (!g1553)) + ((g1008) & (!g1071) & (!g1163) & (!g1348) & (!g1544) & (g1553)) + ((g1008) & (!g1071) & (!g1163) & (g1348) & (g1544) & (!g1553)) + ((g1008) & (!g1071) & (!g1163) & (g1348) & (g1544) & (g1553)) + ((g1008) & (!g1071) & (g1163) & (!g1348) & (!g1544) & (!g1553)) + ((g1008) & (!g1071) & (g1163) & (!g1348) & (g1544) & (!g1553)) + ((g1008) & (!g1071) & (g1163) & (g1348) & (!g1544) & (!g1553)) + ((g1008) & (!g1071) & (g1163) & (g1348) & (g1544) & (!g1553)) + ((g1008) & (g1071) & (!g1163) & (!g1348) & (g1544) & (!g1553)) + ((g1008) & (g1071) & (!g1163) & (!g1348) & (g1544) & (g1553)) + ((g1008) & (g1071) & (!g1163) & (g1348) & (!g1544) & (!g1553)) + ((g1008) & (g1071) & (!g1163) & (g1348) & (!g1544) & (g1553)) + ((g1008) & (g1071) & (g1163) & (!g1348) & (!g1544) & (!g1553)) + ((g1008) & (g1071) & (g1163) & (!g1348) & (g1544) & (!g1553)) + ((g1008) & (g1071) & (g1163) & (g1348) & (!g1544) & (!g1553)) + ((g1008) & (g1071) & (g1163) & (g1348) & (g1544) & (!g1553)));
	assign g2129 = (((!sk[4]) & (!ld) & (text_inx111x) & (!g1555)) + ((!sk[4]) & (!ld) & (text_inx111x) & (g1555)) + ((!sk[4]) & (ld) & (!text_inx111x) & (g1555)) + ((!sk[4]) & (ld) & (text_inx111x) & (!g1555)) + ((!sk[4]) & (ld) & (text_inx111x) & (g1555)) + ((sk[4]) & (!ld) & (!text_inx111x) & (g1555)) + ((sk[4]) & (!ld) & (text_inx111x) & (g1555)) + ((sk[4]) & (ld) & (text_inx111x) & (!g1555)) + ((sk[4]) & (ld) & (text_inx111x) & (g1555)));
	assign g1556 = (((!g957) & (!g1029) & (!g1092) & (!g1163) & (g1352) & (!g1555)) + ((!g957) & (!g1029) & (!g1092) & (!g1163) & (g1352) & (g1555)) + ((!g957) & (!g1029) & (!g1092) & (g1163) & (!g1352) & (g1555)) + ((!g957) & (!g1029) & (!g1092) & (g1163) & (g1352) & (g1555)) + ((!g957) & (!g1029) & (g1092) & (!g1163) & (!g1352) & (!g1555)) + ((!g957) & (!g1029) & (g1092) & (!g1163) & (!g1352) & (g1555)) + ((!g957) & (!g1029) & (g1092) & (g1163) & (!g1352) & (g1555)) + ((!g957) & (!g1029) & (g1092) & (g1163) & (g1352) & (g1555)) + ((!g957) & (g1029) & (!g1092) & (!g1163) & (!g1352) & (!g1555)) + ((!g957) & (g1029) & (!g1092) & (!g1163) & (!g1352) & (g1555)) + ((!g957) & (g1029) & (!g1092) & (g1163) & (!g1352) & (!g1555)) + ((!g957) & (g1029) & (!g1092) & (g1163) & (g1352) & (!g1555)) + ((!g957) & (g1029) & (g1092) & (!g1163) & (g1352) & (!g1555)) + ((!g957) & (g1029) & (g1092) & (!g1163) & (g1352) & (g1555)) + ((!g957) & (g1029) & (g1092) & (g1163) & (!g1352) & (!g1555)) + ((!g957) & (g1029) & (g1092) & (g1163) & (g1352) & (!g1555)) + ((g957) & (!g1029) & (!g1092) & (!g1163) & (!g1352) & (!g1555)) + ((g957) & (!g1029) & (!g1092) & (!g1163) & (!g1352) & (g1555)) + ((g957) & (!g1029) & (!g1092) & (g1163) & (!g1352) & (g1555)) + ((g957) & (!g1029) & (!g1092) & (g1163) & (g1352) & (g1555)) + ((g957) & (!g1029) & (g1092) & (!g1163) & (g1352) & (!g1555)) + ((g957) & (!g1029) & (g1092) & (!g1163) & (g1352) & (g1555)) + ((g957) & (!g1029) & (g1092) & (g1163) & (!g1352) & (g1555)) + ((g957) & (!g1029) & (g1092) & (g1163) & (g1352) & (g1555)) + ((g957) & (g1029) & (!g1092) & (!g1163) & (g1352) & (!g1555)) + ((g957) & (g1029) & (!g1092) & (!g1163) & (g1352) & (g1555)) + ((g957) & (g1029) & (!g1092) & (g1163) & (!g1352) & (!g1555)) + ((g957) & (g1029) & (!g1092) & (g1163) & (g1352) & (!g1555)) + ((g957) & (g1029) & (g1092) & (!g1163) & (!g1352) & (!g1555)) + ((g957) & (g1029) & (g1092) & (!g1163) & (!g1352) & (g1555)) + ((g957) & (g1029) & (g1092) & (g1163) & (!g1352) & (!g1555)) + ((g957) & (g1029) & (g1092) & (g1163) & (g1352) & (!g1555)));
	assign g1557 = (((!ld) & (!g468) & (!g724) & (!g980) & (g1276) & (!keyx40x)) + ((!ld) & (!g468) & (!g724) & (!g980) & (g1276) & (keyx40x)) + ((!ld) & (!g468) & (!g724) & (g980) & (!g1276) & (!keyx40x)) + ((!ld) & (!g468) & (!g724) & (g980) & (!g1276) & (keyx40x)) + ((!ld) & (!g468) & (g724) & (!g980) & (!g1276) & (!keyx40x)) + ((!ld) & (!g468) & (g724) & (!g980) & (!g1276) & (keyx40x)) + ((!ld) & (!g468) & (g724) & (g980) & (g1276) & (!keyx40x)) + ((!ld) & (!g468) & (g724) & (g980) & (g1276) & (keyx40x)) + ((!ld) & (g468) & (!g724) & (!g980) & (!g1276) & (!keyx40x)) + ((!ld) & (g468) & (!g724) & (!g980) & (!g1276) & (keyx40x)) + ((!ld) & (g468) & (!g724) & (g980) & (g1276) & (!keyx40x)) + ((!ld) & (g468) & (!g724) & (g980) & (g1276) & (keyx40x)) + ((!ld) & (g468) & (g724) & (!g980) & (g1276) & (!keyx40x)) + ((!ld) & (g468) & (g724) & (!g980) & (g1276) & (keyx40x)) + ((!ld) & (g468) & (g724) & (g980) & (!g1276) & (!keyx40x)) + ((!ld) & (g468) & (g724) & (g980) & (!g1276) & (keyx40x)) + ((ld) & (!g468) & (!g724) & (!g980) & (!g1276) & (keyx40x)) + ((ld) & (!g468) & (!g724) & (!g980) & (g1276) & (keyx40x)) + ((ld) & (!g468) & (!g724) & (g980) & (!g1276) & (keyx40x)) + ((ld) & (!g468) & (!g724) & (g980) & (g1276) & (keyx40x)) + ((ld) & (!g468) & (g724) & (!g980) & (!g1276) & (keyx40x)) + ((ld) & (!g468) & (g724) & (!g980) & (g1276) & (keyx40x)) + ((ld) & (!g468) & (g724) & (g980) & (!g1276) & (keyx40x)) + ((ld) & (!g468) & (g724) & (g980) & (g1276) & (keyx40x)) + ((ld) & (g468) & (!g724) & (!g980) & (!g1276) & (keyx40x)) + ((ld) & (g468) & (!g724) & (!g980) & (g1276) & (keyx40x)) + ((ld) & (g468) & (!g724) & (g980) & (!g1276) & (keyx40x)) + ((ld) & (g468) & (!g724) & (g980) & (g1276) & (keyx40x)) + ((ld) & (g468) & (g724) & (!g980) & (!g1276) & (keyx40x)) + ((ld) & (g468) & (g724) & (!g980) & (g1276) & (keyx40x)) + ((ld) & (g468) & (g724) & (g980) & (!g1276) & (keyx40x)) + ((ld) & (g468) & (g724) & (g980) & (g1276) & (keyx40x)));
	assign g1558 = (((!ld) & (!g475) & (!g731) & (!g987) & (g1283) & (!keyx41x)) + ((!ld) & (!g475) & (!g731) & (!g987) & (g1283) & (keyx41x)) + ((!ld) & (!g475) & (!g731) & (g987) & (!g1283) & (!keyx41x)) + ((!ld) & (!g475) & (!g731) & (g987) & (!g1283) & (keyx41x)) + ((!ld) & (!g475) & (g731) & (!g987) & (!g1283) & (!keyx41x)) + ((!ld) & (!g475) & (g731) & (!g987) & (!g1283) & (keyx41x)) + ((!ld) & (!g475) & (g731) & (g987) & (g1283) & (!keyx41x)) + ((!ld) & (!g475) & (g731) & (g987) & (g1283) & (keyx41x)) + ((!ld) & (g475) & (!g731) & (!g987) & (!g1283) & (!keyx41x)) + ((!ld) & (g475) & (!g731) & (!g987) & (!g1283) & (keyx41x)) + ((!ld) & (g475) & (!g731) & (g987) & (g1283) & (!keyx41x)) + ((!ld) & (g475) & (!g731) & (g987) & (g1283) & (keyx41x)) + ((!ld) & (g475) & (g731) & (!g987) & (g1283) & (!keyx41x)) + ((!ld) & (g475) & (g731) & (!g987) & (g1283) & (keyx41x)) + ((!ld) & (g475) & (g731) & (g987) & (!g1283) & (!keyx41x)) + ((!ld) & (g475) & (g731) & (g987) & (!g1283) & (keyx41x)) + ((ld) & (!g475) & (!g731) & (!g987) & (!g1283) & (keyx41x)) + ((ld) & (!g475) & (!g731) & (!g987) & (g1283) & (keyx41x)) + ((ld) & (!g475) & (!g731) & (g987) & (!g1283) & (keyx41x)) + ((ld) & (!g475) & (!g731) & (g987) & (g1283) & (keyx41x)) + ((ld) & (!g475) & (g731) & (!g987) & (!g1283) & (keyx41x)) + ((ld) & (!g475) & (g731) & (!g987) & (g1283) & (keyx41x)) + ((ld) & (!g475) & (g731) & (g987) & (!g1283) & (keyx41x)) + ((ld) & (!g475) & (g731) & (g987) & (g1283) & (keyx41x)) + ((ld) & (g475) & (!g731) & (!g987) & (!g1283) & (keyx41x)) + ((ld) & (g475) & (!g731) & (!g987) & (g1283) & (keyx41x)) + ((ld) & (g475) & (!g731) & (g987) & (!g1283) & (keyx41x)) + ((ld) & (g475) & (!g731) & (g987) & (g1283) & (keyx41x)) + ((ld) & (g475) & (g731) & (!g987) & (!g1283) & (keyx41x)) + ((ld) & (g475) & (g731) & (!g987) & (g1283) & (keyx41x)) + ((ld) & (g475) & (g731) & (g987) & (!g1283) & (keyx41x)) + ((ld) & (g475) & (g731) & (g987) & (g1283) & (keyx41x)));
	assign g1559 = (((!ld) & (!g482) & (!g738) & (!g994) & (g1290) & (!keyx42x)) + ((!ld) & (!g482) & (!g738) & (!g994) & (g1290) & (keyx42x)) + ((!ld) & (!g482) & (!g738) & (g994) & (!g1290) & (!keyx42x)) + ((!ld) & (!g482) & (!g738) & (g994) & (!g1290) & (keyx42x)) + ((!ld) & (!g482) & (g738) & (!g994) & (!g1290) & (!keyx42x)) + ((!ld) & (!g482) & (g738) & (!g994) & (!g1290) & (keyx42x)) + ((!ld) & (!g482) & (g738) & (g994) & (g1290) & (!keyx42x)) + ((!ld) & (!g482) & (g738) & (g994) & (g1290) & (keyx42x)) + ((!ld) & (g482) & (!g738) & (!g994) & (!g1290) & (!keyx42x)) + ((!ld) & (g482) & (!g738) & (!g994) & (!g1290) & (keyx42x)) + ((!ld) & (g482) & (!g738) & (g994) & (g1290) & (!keyx42x)) + ((!ld) & (g482) & (!g738) & (g994) & (g1290) & (keyx42x)) + ((!ld) & (g482) & (g738) & (!g994) & (g1290) & (!keyx42x)) + ((!ld) & (g482) & (g738) & (!g994) & (g1290) & (keyx42x)) + ((!ld) & (g482) & (g738) & (g994) & (!g1290) & (!keyx42x)) + ((!ld) & (g482) & (g738) & (g994) & (!g1290) & (keyx42x)) + ((ld) & (!g482) & (!g738) & (!g994) & (!g1290) & (keyx42x)) + ((ld) & (!g482) & (!g738) & (!g994) & (g1290) & (keyx42x)) + ((ld) & (!g482) & (!g738) & (g994) & (!g1290) & (keyx42x)) + ((ld) & (!g482) & (!g738) & (g994) & (g1290) & (keyx42x)) + ((ld) & (!g482) & (g738) & (!g994) & (!g1290) & (keyx42x)) + ((ld) & (!g482) & (g738) & (!g994) & (g1290) & (keyx42x)) + ((ld) & (!g482) & (g738) & (g994) & (!g1290) & (keyx42x)) + ((ld) & (!g482) & (g738) & (g994) & (g1290) & (keyx42x)) + ((ld) & (g482) & (!g738) & (!g994) & (!g1290) & (keyx42x)) + ((ld) & (g482) & (!g738) & (!g994) & (g1290) & (keyx42x)) + ((ld) & (g482) & (!g738) & (g994) & (!g1290) & (keyx42x)) + ((ld) & (g482) & (!g738) & (g994) & (g1290) & (keyx42x)) + ((ld) & (g482) & (g738) & (!g994) & (!g1290) & (keyx42x)) + ((ld) & (g482) & (g738) & (!g994) & (g1290) & (keyx42x)) + ((ld) & (g482) & (g738) & (g994) & (!g1290) & (keyx42x)) + ((ld) & (g482) & (g738) & (g994) & (g1290) & (keyx42x)));
	assign g1560 = (((!ld) & (!g489) & (!g745) & (!g1001) & (g1297) & (!keyx43x)) + ((!ld) & (!g489) & (!g745) & (!g1001) & (g1297) & (keyx43x)) + ((!ld) & (!g489) & (!g745) & (g1001) & (!g1297) & (!keyx43x)) + ((!ld) & (!g489) & (!g745) & (g1001) & (!g1297) & (keyx43x)) + ((!ld) & (!g489) & (g745) & (!g1001) & (!g1297) & (!keyx43x)) + ((!ld) & (!g489) & (g745) & (!g1001) & (!g1297) & (keyx43x)) + ((!ld) & (!g489) & (g745) & (g1001) & (g1297) & (!keyx43x)) + ((!ld) & (!g489) & (g745) & (g1001) & (g1297) & (keyx43x)) + ((!ld) & (g489) & (!g745) & (!g1001) & (!g1297) & (!keyx43x)) + ((!ld) & (g489) & (!g745) & (!g1001) & (!g1297) & (keyx43x)) + ((!ld) & (g489) & (!g745) & (g1001) & (g1297) & (!keyx43x)) + ((!ld) & (g489) & (!g745) & (g1001) & (g1297) & (keyx43x)) + ((!ld) & (g489) & (g745) & (!g1001) & (g1297) & (!keyx43x)) + ((!ld) & (g489) & (g745) & (!g1001) & (g1297) & (keyx43x)) + ((!ld) & (g489) & (g745) & (g1001) & (!g1297) & (!keyx43x)) + ((!ld) & (g489) & (g745) & (g1001) & (!g1297) & (keyx43x)) + ((ld) & (!g489) & (!g745) & (!g1001) & (!g1297) & (keyx43x)) + ((ld) & (!g489) & (!g745) & (!g1001) & (g1297) & (keyx43x)) + ((ld) & (!g489) & (!g745) & (g1001) & (!g1297) & (keyx43x)) + ((ld) & (!g489) & (!g745) & (g1001) & (g1297) & (keyx43x)) + ((ld) & (!g489) & (g745) & (!g1001) & (!g1297) & (keyx43x)) + ((ld) & (!g489) & (g745) & (!g1001) & (g1297) & (keyx43x)) + ((ld) & (!g489) & (g745) & (g1001) & (!g1297) & (keyx43x)) + ((ld) & (!g489) & (g745) & (g1001) & (g1297) & (keyx43x)) + ((ld) & (g489) & (!g745) & (!g1001) & (!g1297) & (keyx43x)) + ((ld) & (g489) & (!g745) & (!g1001) & (g1297) & (keyx43x)) + ((ld) & (g489) & (!g745) & (g1001) & (!g1297) & (keyx43x)) + ((ld) & (g489) & (!g745) & (g1001) & (g1297) & (keyx43x)) + ((ld) & (g489) & (g745) & (!g1001) & (!g1297) & (keyx43x)) + ((ld) & (g489) & (g745) & (!g1001) & (g1297) & (keyx43x)) + ((ld) & (g489) & (g745) & (g1001) & (!g1297) & (keyx43x)) + ((ld) & (g489) & (g745) & (g1001) & (g1297) & (keyx43x)));
	assign g1561 = (((!ld) & (!g496) & (!g752) & (!g1008) & (g1304) & (!keyx44x)) + ((!ld) & (!g496) & (!g752) & (!g1008) & (g1304) & (keyx44x)) + ((!ld) & (!g496) & (!g752) & (g1008) & (!g1304) & (!keyx44x)) + ((!ld) & (!g496) & (!g752) & (g1008) & (!g1304) & (keyx44x)) + ((!ld) & (!g496) & (g752) & (!g1008) & (!g1304) & (!keyx44x)) + ((!ld) & (!g496) & (g752) & (!g1008) & (!g1304) & (keyx44x)) + ((!ld) & (!g496) & (g752) & (g1008) & (g1304) & (!keyx44x)) + ((!ld) & (!g496) & (g752) & (g1008) & (g1304) & (keyx44x)) + ((!ld) & (g496) & (!g752) & (!g1008) & (!g1304) & (!keyx44x)) + ((!ld) & (g496) & (!g752) & (!g1008) & (!g1304) & (keyx44x)) + ((!ld) & (g496) & (!g752) & (g1008) & (g1304) & (!keyx44x)) + ((!ld) & (g496) & (!g752) & (g1008) & (g1304) & (keyx44x)) + ((!ld) & (g496) & (g752) & (!g1008) & (g1304) & (!keyx44x)) + ((!ld) & (g496) & (g752) & (!g1008) & (g1304) & (keyx44x)) + ((!ld) & (g496) & (g752) & (g1008) & (!g1304) & (!keyx44x)) + ((!ld) & (g496) & (g752) & (g1008) & (!g1304) & (keyx44x)) + ((ld) & (!g496) & (!g752) & (!g1008) & (!g1304) & (keyx44x)) + ((ld) & (!g496) & (!g752) & (!g1008) & (g1304) & (keyx44x)) + ((ld) & (!g496) & (!g752) & (g1008) & (!g1304) & (keyx44x)) + ((ld) & (!g496) & (!g752) & (g1008) & (g1304) & (keyx44x)) + ((ld) & (!g496) & (g752) & (!g1008) & (!g1304) & (keyx44x)) + ((ld) & (!g496) & (g752) & (!g1008) & (g1304) & (keyx44x)) + ((ld) & (!g496) & (g752) & (g1008) & (!g1304) & (keyx44x)) + ((ld) & (!g496) & (g752) & (g1008) & (g1304) & (keyx44x)) + ((ld) & (g496) & (!g752) & (!g1008) & (!g1304) & (keyx44x)) + ((ld) & (g496) & (!g752) & (!g1008) & (g1304) & (keyx44x)) + ((ld) & (g496) & (!g752) & (g1008) & (!g1304) & (keyx44x)) + ((ld) & (g496) & (!g752) & (g1008) & (g1304) & (keyx44x)) + ((ld) & (g496) & (g752) & (!g1008) & (!g1304) & (keyx44x)) + ((ld) & (g496) & (g752) & (!g1008) & (g1304) & (keyx44x)) + ((ld) & (g496) & (g752) & (g1008) & (!g1304) & (keyx44x)) + ((ld) & (g496) & (g752) & (g1008) & (g1304) & (keyx44x)));
	assign g1562 = (((!ld) & (!g503) & (!g759) & (!g1015) & (g1311) & (!keyx45x)) + ((!ld) & (!g503) & (!g759) & (!g1015) & (g1311) & (keyx45x)) + ((!ld) & (!g503) & (!g759) & (g1015) & (!g1311) & (!keyx45x)) + ((!ld) & (!g503) & (!g759) & (g1015) & (!g1311) & (keyx45x)) + ((!ld) & (!g503) & (g759) & (!g1015) & (!g1311) & (!keyx45x)) + ((!ld) & (!g503) & (g759) & (!g1015) & (!g1311) & (keyx45x)) + ((!ld) & (!g503) & (g759) & (g1015) & (g1311) & (!keyx45x)) + ((!ld) & (!g503) & (g759) & (g1015) & (g1311) & (keyx45x)) + ((!ld) & (g503) & (!g759) & (!g1015) & (!g1311) & (!keyx45x)) + ((!ld) & (g503) & (!g759) & (!g1015) & (!g1311) & (keyx45x)) + ((!ld) & (g503) & (!g759) & (g1015) & (g1311) & (!keyx45x)) + ((!ld) & (g503) & (!g759) & (g1015) & (g1311) & (keyx45x)) + ((!ld) & (g503) & (g759) & (!g1015) & (g1311) & (!keyx45x)) + ((!ld) & (g503) & (g759) & (!g1015) & (g1311) & (keyx45x)) + ((!ld) & (g503) & (g759) & (g1015) & (!g1311) & (!keyx45x)) + ((!ld) & (g503) & (g759) & (g1015) & (!g1311) & (keyx45x)) + ((ld) & (!g503) & (!g759) & (!g1015) & (!g1311) & (keyx45x)) + ((ld) & (!g503) & (!g759) & (!g1015) & (g1311) & (keyx45x)) + ((ld) & (!g503) & (!g759) & (g1015) & (!g1311) & (keyx45x)) + ((ld) & (!g503) & (!g759) & (g1015) & (g1311) & (keyx45x)) + ((ld) & (!g503) & (g759) & (!g1015) & (!g1311) & (keyx45x)) + ((ld) & (!g503) & (g759) & (!g1015) & (g1311) & (keyx45x)) + ((ld) & (!g503) & (g759) & (g1015) & (!g1311) & (keyx45x)) + ((ld) & (!g503) & (g759) & (g1015) & (g1311) & (keyx45x)) + ((ld) & (g503) & (!g759) & (!g1015) & (!g1311) & (keyx45x)) + ((ld) & (g503) & (!g759) & (!g1015) & (g1311) & (keyx45x)) + ((ld) & (g503) & (!g759) & (g1015) & (!g1311) & (keyx45x)) + ((ld) & (g503) & (!g759) & (g1015) & (g1311) & (keyx45x)) + ((ld) & (g503) & (g759) & (!g1015) & (!g1311) & (keyx45x)) + ((ld) & (g503) & (g759) & (!g1015) & (g1311) & (keyx45x)) + ((ld) & (g503) & (g759) & (g1015) & (!g1311) & (keyx45x)) + ((ld) & (g503) & (g759) & (g1015) & (g1311) & (keyx45x)));
	assign g1563 = (((!ld) & (!g510) & (!g766) & (!g1022) & (g1318) & (!keyx46x)) + ((!ld) & (!g510) & (!g766) & (!g1022) & (g1318) & (keyx46x)) + ((!ld) & (!g510) & (!g766) & (g1022) & (!g1318) & (!keyx46x)) + ((!ld) & (!g510) & (!g766) & (g1022) & (!g1318) & (keyx46x)) + ((!ld) & (!g510) & (g766) & (!g1022) & (!g1318) & (!keyx46x)) + ((!ld) & (!g510) & (g766) & (!g1022) & (!g1318) & (keyx46x)) + ((!ld) & (!g510) & (g766) & (g1022) & (g1318) & (!keyx46x)) + ((!ld) & (!g510) & (g766) & (g1022) & (g1318) & (keyx46x)) + ((!ld) & (g510) & (!g766) & (!g1022) & (!g1318) & (!keyx46x)) + ((!ld) & (g510) & (!g766) & (!g1022) & (!g1318) & (keyx46x)) + ((!ld) & (g510) & (!g766) & (g1022) & (g1318) & (!keyx46x)) + ((!ld) & (g510) & (!g766) & (g1022) & (g1318) & (keyx46x)) + ((!ld) & (g510) & (g766) & (!g1022) & (g1318) & (!keyx46x)) + ((!ld) & (g510) & (g766) & (!g1022) & (g1318) & (keyx46x)) + ((!ld) & (g510) & (g766) & (g1022) & (!g1318) & (!keyx46x)) + ((!ld) & (g510) & (g766) & (g1022) & (!g1318) & (keyx46x)) + ((ld) & (!g510) & (!g766) & (!g1022) & (!g1318) & (keyx46x)) + ((ld) & (!g510) & (!g766) & (!g1022) & (g1318) & (keyx46x)) + ((ld) & (!g510) & (!g766) & (g1022) & (!g1318) & (keyx46x)) + ((ld) & (!g510) & (!g766) & (g1022) & (g1318) & (keyx46x)) + ((ld) & (!g510) & (g766) & (!g1022) & (!g1318) & (keyx46x)) + ((ld) & (!g510) & (g766) & (!g1022) & (g1318) & (keyx46x)) + ((ld) & (!g510) & (g766) & (g1022) & (!g1318) & (keyx46x)) + ((ld) & (!g510) & (g766) & (g1022) & (g1318) & (keyx46x)) + ((ld) & (g510) & (!g766) & (!g1022) & (!g1318) & (keyx46x)) + ((ld) & (g510) & (!g766) & (!g1022) & (g1318) & (keyx46x)) + ((ld) & (g510) & (!g766) & (g1022) & (!g1318) & (keyx46x)) + ((ld) & (g510) & (!g766) & (g1022) & (g1318) & (keyx46x)) + ((ld) & (g510) & (g766) & (!g1022) & (!g1318) & (keyx46x)) + ((ld) & (g510) & (g766) & (!g1022) & (g1318) & (keyx46x)) + ((ld) & (g510) & (g766) & (g1022) & (!g1318) & (keyx46x)) + ((ld) & (g510) & (g766) & (g1022) & (g1318) & (keyx46x)));
	assign g1564 = (((!ld) & (!g517) & (!g773) & (!g1029) & (g1325) & (!keyx47x)) + ((!ld) & (!g517) & (!g773) & (!g1029) & (g1325) & (keyx47x)) + ((!ld) & (!g517) & (!g773) & (g1029) & (!g1325) & (!keyx47x)) + ((!ld) & (!g517) & (!g773) & (g1029) & (!g1325) & (keyx47x)) + ((!ld) & (!g517) & (g773) & (!g1029) & (!g1325) & (!keyx47x)) + ((!ld) & (!g517) & (g773) & (!g1029) & (!g1325) & (keyx47x)) + ((!ld) & (!g517) & (g773) & (g1029) & (g1325) & (!keyx47x)) + ((!ld) & (!g517) & (g773) & (g1029) & (g1325) & (keyx47x)) + ((!ld) & (g517) & (!g773) & (!g1029) & (!g1325) & (!keyx47x)) + ((!ld) & (g517) & (!g773) & (!g1029) & (!g1325) & (keyx47x)) + ((!ld) & (g517) & (!g773) & (g1029) & (g1325) & (!keyx47x)) + ((!ld) & (g517) & (!g773) & (g1029) & (g1325) & (keyx47x)) + ((!ld) & (g517) & (g773) & (!g1029) & (g1325) & (!keyx47x)) + ((!ld) & (g517) & (g773) & (!g1029) & (g1325) & (keyx47x)) + ((!ld) & (g517) & (g773) & (g1029) & (!g1325) & (!keyx47x)) + ((!ld) & (g517) & (g773) & (g1029) & (!g1325) & (keyx47x)) + ((ld) & (!g517) & (!g773) & (!g1029) & (!g1325) & (keyx47x)) + ((ld) & (!g517) & (!g773) & (!g1029) & (g1325) & (keyx47x)) + ((ld) & (!g517) & (!g773) & (g1029) & (!g1325) & (keyx47x)) + ((ld) & (!g517) & (!g773) & (g1029) & (g1325) & (keyx47x)) + ((ld) & (!g517) & (g773) & (!g1029) & (!g1325) & (keyx47x)) + ((ld) & (!g517) & (g773) & (!g1029) & (g1325) & (keyx47x)) + ((ld) & (!g517) & (g773) & (g1029) & (!g1325) & (keyx47x)) + ((ld) & (!g517) & (g773) & (g1029) & (g1325) & (keyx47x)) + ((ld) & (g517) & (!g773) & (!g1029) & (!g1325) & (keyx47x)) + ((ld) & (g517) & (!g773) & (!g1029) & (g1325) & (keyx47x)) + ((ld) & (g517) & (!g773) & (g1029) & (!g1325) & (keyx47x)) + ((ld) & (g517) & (!g773) & (g1029) & (g1325) & (keyx47x)) + ((ld) & (g517) & (g773) & (!g1029) & (!g1325) & (keyx47x)) + ((ld) & (g517) & (g773) & (!g1029) & (g1325) & (keyx47x)) + ((ld) & (g517) & (g773) & (g1029) & (!g1325) & (keyx47x)) + ((ld) & (g517) & (g773) & (g1029) & (g1325) & (keyx47x)));
	assign g2130 = (((!ld) & (!text_inx16x) & (sk[14]) & (g1565)) + ((!ld) & (text_inx16x) & (!sk[14]) & (!g1565)) + ((!ld) & (text_inx16x) & (!sk[14]) & (g1565)) + ((!ld) & (text_inx16x) & (sk[14]) & (g1565)) + ((ld) & (!text_inx16x) & (!sk[14]) & (g1565)) + ((ld) & (text_inx16x) & (!sk[14]) & (!g1565)) + ((ld) & (text_inx16x) & (!sk[14]) & (g1565)) + ((ld) & (text_inx16x) & (sk[14]) & (!g1565)) + ((ld) & (text_inx16x) & (sk[14]) & (g1565)));
	assign g1566 = (((!g260) & (!sk[15]) & (g324)) + ((!g260) & (sk[15]) & (g324)) + ((g260) & (!sk[15]) & (g324)) + ((g260) & (sk[15]) & (!g324)));
	assign g1567 = (((!g276) & (!g339) & (!g1163) & (!g1411) & (!g1565) & (g1566)) + ((!g276) & (!g339) & (!g1163) & (!g1411) & (g1565) & (g1566)) + ((!g276) & (!g339) & (!g1163) & (g1411) & (!g1565) & (!g1566)) + ((!g276) & (!g339) & (!g1163) & (g1411) & (g1565) & (!g1566)) + ((!g276) & (!g339) & (g1163) & (!g1411) & (g1565) & (!g1566)) + ((!g276) & (!g339) & (g1163) & (!g1411) & (g1565) & (g1566)) + ((!g276) & (!g339) & (g1163) & (g1411) & (g1565) & (!g1566)) + ((!g276) & (!g339) & (g1163) & (g1411) & (g1565) & (g1566)) + ((!g276) & (g339) & (!g1163) & (!g1411) & (!g1565) & (!g1566)) + ((!g276) & (g339) & (!g1163) & (!g1411) & (g1565) & (!g1566)) + ((!g276) & (g339) & (!g1163) & (g1411) & (!g1565) & (g1566)) + ((!g276) & (g339) & (!g1163) & (g1411) & (g1565) & (g1566)) + ((!g276) & (g339) & (g1163) & (!g1411) & (g1565) & (!g1566)) + ((!g276) & (g339) & (g1163) & (!g1411) & (g1565) & (g1566)) + ((!g276) & (g339) & (g1163) & (g1411) & (g1565) & (!g1566)) + ((!g276) & (g339) & (g1163) & (g1411) & (g1565) & (g1566)) + ((g276) & (!g339) & (!g1163) & (!g1411) & (!g1565) & (!g1566)) + ((g276) & (!g339) & (!g1163) & (!g1411) & (g1565) & (!g1566)) + ((g276) & (!g339) & (!g1163) & (g1411) & (!g1565) & (g1566)) + ((g276) & (!g339) & (!g1163) & (g1411) & (g1565) & (g1566)) + ((g276) & (!g339) & (g1163) & (!g1411) & (!g1565) & (!g1566)) + ((g276) & (!g339) & (g1163) & (!g1411) & (!g1565) & (g1566)) + ((g276) & (!g339) & (g1163) & (g1411) & (!g1565) & (!g1566)) + ((g276) & (!g339) & (g1163) & (g1411) & (!g1565) & (g1566)) + ((g276) & (g339) & (!g1163) & (!g1411) & (!g1565) & (g1566)) + ((g276) & (g339) & (!g1163) & (!g1411) & (g1565) & (g1566)) + ((g276) & (g339) & (!g1163) & (g1411) & (!g1565) & (!g1566)) + ((g276) & (g339) & (!g1163) & (g1411) & (g1565) & (!g1566)) + ((g276) & (g339) & (g1163) & (!g1411) & (!g1565) & (!g1566)) + ((g276) & (g339) & (g1163) & (!g1411) & (!g1565) & (g1566)) + ((g276) & (g339) & (g1163) & (g1411) & (!g1565) & (!g1566)) + ((g276) & (g339) & (g1163) & (g1411) & (!g1565) & (g1566)));
	assign g2131 = (((!ld) & (!text_inx17x) & (sk[17]) & (g1568)) + ((!ld) & (text_inx17x) & (!sk[17]) & (!g1568)) + ((!ld) & (text_inx17x) & (!sk[17]) & (g1568)) + ((!ld) & (text_inx17x) & (sk[17]) & (g1568)) + ((ld) & (!text_inx17x) & (!sk[17]) & (g1568)) + ((ld) & (text_inx17x) & (!sk[17]) & (!g1568)) + ((ld) & (text_inx17x) & (!sk[17]) & (g1568)) + ((ld) & (text_inx17x) & (sk[17]) & (!g1568)) + ((ld) & (text_inx17x) & (sk[17]) & (g1568)));
	assign g2132 = (((!sk[18]) & (!ld) & (text_inx18x) & (!g1569)) + ((!sk[18]) & (!ld) & (text_inx18x) & (g1569)) + ((!sk[18]) & (ld) & (!text_inx18x) & (g1569)) + ((!sk[18]) & (ld) & (text_inx18x) & (!g1569)) + ((!sk[18]) & (ld) & (text_inx18x) & (g1569)) + ((sk[18]) & (!ld) & (!text_inx18x) & (g1569)) + ((sk[18]) & (!ld) & (text_inx18x) & (g1569)) + ((sk[18]) & (ld) & (text_inx18x) & (!g1569)) + ((sk[18]) & (ld) & (text_inx18x) & (g1569)));
	assign g1570 = (((!g218) & (!g290) & (!g353) & (!g1163) & (g1417) & (!g1569)) + ((!g218) & (!g290) & (!g353) & (!g1163) & (g1417) & (g1569)) + ((!g218) & (!g290) & (!g353) & (g1163) & (!g1417) & (g1569)) + ((!g218) & (!g290) & (!g353) & (g1163) & (g1417) & (g1569)) + ((!g218) & (!g290) & (g353) & (!g1163) & (!g1417) & (!g1569)) + ((!g218) & (!g290) & (g353) & (!g1163) & (!g1417) & (g1569)) + ((!g218) & (!g290) & (g353) & (g1163) & (!g1417) & (g1569)) + ((!g218) & (!g290) & (g353) & (g1163) & (g1417) & (g1569)) + ((!g218) & (g290) & (!g353) & (!g1163) & (!g1417) & (!g1569)) + ((!g218) & (g290) & (!g353) & (!g1163) & (!g1417) & (g1569)) + ((!g218) & (g290) & (!g353) & (g1163) & (!g1417) & (!g1569)) + ((!g218) & (g290) & (!g353) & (g1163) & (g1417) & (!g1569)) + ((!g218) & (g290) & (g353) & (!g1163) & (g1417) & (!g1569)) + ((!g218) & (g290) & (g353) & (!g1163) & (g1417) & (g1569)) + ((!g218) & (g290) & (g353) & (g1163) & (!g1417) & (!g1569)) + ((!g218) & (g290) & (g353) & (g1163) & (g1417) & (!g1569)) + ((g218) & (!g290) & (!g353) & (!g1163) & (!g1417) & (!g1569)) + ((g218) & (!g290) & (!g353) & (!g1163) & (!g1417) & (g1569)) + ((g218) & (!g290) & (!g353) & (g1163) & (!g1417) & (g1569)) + ((g218) & (!g290) & (!g353) & (g1163) & (g1417) & (g1569)) + ((g218) & (!g290) & (g353) & (!g1163) & (g1417) & (!g1569)) + ((g218) & (!g290) & (g353) & (!g1163) & (g1417) & (g1569)) + ((g218) & (!g290) & (g353) & (g1163) & (!g1417) & (g1569)) + ((g218) & (!g290) & (g353) & (g1163) & (g1417) & (g1569)) + ((g218) & (g290) & (!g353) & (!g1163) & (g1417) & (!g1569)) + ((g218) & (g290) & (!g353) & (!g1163) & (g1417) & (g1569)) + ((g218) & (g290) & (!g353) & (g1163) & (!g1417) & (!g1569)) + ((g218) & (g290) & (!g353) & (g1163) & (g1417) & (!g1569)) + ((g218) & (g290) & (g353) & (!g1163) & (!g1417) & (!g1569)) + ((g218) & (g290) & (g353) & (!g1163) & (!g1417) & (g1569)) + ((g218) & (g290) & (g353) & (g1163) & (!g1417) & (!g1569)) + ((g218) & (g290) & (g353) & (g1163) & (g1417) & (!g1569)));
	assign g2133 = (((!sk[20]) & (!ld) & (text_inx19x) & (!g1571)) + ((!sk[20]) & (!ld) & (text_inx19x) & (g1571)) + ((!sk[20]) & (ld) & (!text_inx19x) & (g1571)) + ((!sk[20]) & (ld) & (text_inx19x) & (!g1571)) + ((!sk[20]) & (ld) & (text_inx19x) & (g1571)) + ((sk[20]) & (!ld) & (!text_inx19x) & (g1571)) + ((sk[20]) & (!ld) & (text_inx19x) & (g1571)) + ((sk[20]) & (ld) & (text_inx19x) & (!g1571)) + ((sk[20]) & (ld) & (text_inx19x) & (g1571)));
	assign g1572 = (((!g168) & (!g225) & (!g232) & (!g289) & (sk[21]) & (g297)) + ((!g168) & (!g225) & (!g232) & (g289) & (sk[21]) & (!g297)) + ((!g168) & (!g225) & (g232) & (!g289) & (sk[21]) & (!g297)) + ((!g168) & (!g225) & (g232) & (g289) & (sk[21]) & (g297)) + ((!g168) & (g225) & (!g232) & (!g289) & (!sk[21]) & (!g297)) + ((!g168) & (g225) & (!g232) & (!g289) & (!sk[21]) & (g297)) + ((!g168) & (g225) & (!g232) & (!g289) & (sk[21]) & (!g297)) + ((!g168) & (g225) & (!g232) & (g289) & (!sk[21]) & (!g297)) + ((!g168) & (g225) & (!g232) & (g289) & (!sk[21]) & (g297)) + ((!g168) & (g225) & (!g232) & (g289) & (sk[21]) & (g297)) + ((!g168) & (g225) & (g232) & (!g289) & (!sk[21]) & (!g297)) + ((!g168) & (g225) & (g232) & (!g289) & (!sk[21]) & (g297)) + ((!g168) & (g225) & (g232) & (!g289) & (sk[21]) & (g297)) + ((!g168) & (g225) & (g232) & (g289) & (!sk[21]) & (!g297)) + ((!g168) & (g225) & (g232) & (g289) & (!sk[21]) & (g297)) + ((!g168) & (g225) & (g232) & (g289) & (sk[21]) & (!g297)) + ((g168) & (!g225) & (!g232) & (!g289) & (!sk[21]) & (!g297)) + ((g168) & (!g225) & (!g232) & (!g289) & (!sk[21]) & (g297)) + ((g168) & (!g225) & (!g232) & (!g289) & (sk[21]) & (!g297)) + ((g168) & (!g225) & (!g232) & (g289) & (!sk[21]) & (!g297)) + ((g168) & (!g225) & (!g232) & (g289) & (!sk[21]) & (g297)) + ((g168) & (!g225) & (!g232) & (g289) & (sk[21]) & (g297)) + ((g168) & (!g225) & (g232) & (!g289) & (!sk[21]) & (!g297)) + ((g168) & (!g225) & (g232) & (!g289) & (!sk[21]) & (g297)) + ((g168) & (!g225) & (g232) & (!g289) & (sk[21]) & (g297)) + ((g168) & (!g225) & (g232) & (g289) & (!sk[21]) & (!g297)) + ((g168) & (!g225) & (g232) & (g289) & (!sk[21]) & (g297)) + ((g168) & (!g225) & (g232) & (g289) & (sk[21]) & (!g297)) + ((g168) & (g225) & (!g232) & (!g289) & (!sk[21]) & (!g297)) + ((g168) & (g225) & (!g232) & (!g289) & (!sk[21]) & (g297)) + ((g168) & (g225) & (!g232) & (!g289) & (sk[21]) & (g297)) + ((g168) & (g225) & (!g232) & (g289) & (!sk[21]) & (!g297)) + ((g168) & (g225) & (!g232) & (g289) & (!sk[21]) & (g297)) + ((g168) & (g225) & (!g232) & (g289) & (sk[21]) & (!g297)) + ((g168) & (g225) & (g232) & (!g289) & (!sk[21]) & (!g297)) + ((g168) & (g225) & (g232) & (!g289) & (!sk[21]) & (g297)) + ((g168) & (g225) & (g232) & (!g289) & (sk[21]) & (!g297)) + ((g168) & (g225) & (g232) & (g289) & (!sk[21]) & (!g297)) + ((g168) & (g225) & (g232) & (g289) & (!sk[21]) & (g297)) + ((g168) & (g225) & (g232) & (g289) & (sk[21]) & (g297)));
	assign g1573 = (((!g297) & (!g360) & (!g1163) & (!g1566) & (!g1571) & (g1572)) + ((!g297) & (!g360) & (!g1163) & (!g1566) & (g1571) & (g1572)) + ((!g297) & (!g360) & (!g1163) & (g1566) & (!g1571) & (!g1572)) + ((!g297) & (!g360) & (!g1163) & (g1566) & (g1571) & (!g1572)) + ((!g297) & (!g360) & (g1163) & (!g1566) & (g1571) & (!g1572)) + ((!g297) & (!g360) & (g1163) & (!g1566) & (g1571) & (g1572)) + ((!g297) & (!g360) & (g1163) & (g1566) & (g1571) & (!g1572)) + ((!g297) & (!g360) & (g1163) & (g1566) & (g1571) & (g1572)) + ((!g297) & (g360) & (!g1163) & (!g1566) & (!g1571) & (!g1572)) + ((!g297) & (g360) & (!g1163) & (!g1566) & (g1571) & (!g1572)) + ((!g297) & (g360) & (!g1163) & (g1566) & (!g1571) & (g1572)) + ((!g297) & (g360) & (!g1163) & (g1566) & (g1571) & (g1572)) + ((!g297) & (g360) & (g1163) & (!g1566) & (g1571) & (!g1572)) + ((!g297) & (g360) & (g1163) & (!g1566) & (g1571) & (g1572)) + ((!g297) & (g360) & (g1163) & (g1566) & (g1571) & (!g1572)) + ((!g297) & (g360) & (g1163) & (g1566) & (g1571) & (g1572)) + ((g297) & (!g360) & (!g1163) & (!g1566) & (!g1571) & (g1572)) + ((g297) & (!g360) & (!g1163) & (!g1566) & (g1571) & (g1572)) + ((g297) & (!g360) & (!g1163) & (g1566) & (!g1571) & (!g1572)) + ((g297) & (!g360) & (!g1163) & (g1566) & (g1571) & (!g1572)) + ((g297) & (!g360) & (g1163) & (!g1566) & (!g1571) & (!g1572)) + ((g297) & (!g360) & (g1163) & (!g1566) & (!g1571) & (g1572)) + ((g297) & (!g360) & (g1163) & (g1566) & (!g1571) & (!g1572)) + ((g297) & (!g360) & (g1163) & (g1566) & (!g1571) & (g1572)) + ((g297) & (g360) & (!g1163) & (!g1566) & (!g1571) & (!g1572)) + ((g297) & (g360) & (!g1163) & (!g1566) & (g1571) & (!g1572)) + ((g297) & (g360) & (!g1163) & (g1566) & (!g1571) & (g1572)) + ((g297) & (g360) & (!g1163) & (g1566) & (g1571) & (g1572)) + ((g297) & (g360) & (g1163) & (!g1566) & (!g1571) & (!g1572)) + ((g297) & (g360) & (g1163) & (!g1566) & (!g1571) & (g1572)) + ((g297) & (g360) & (g1163) & (g1566) & (!g1571) & (!g1572)) + ((g297) & (g360) & (g1163) & (g1566) & (!g1571) & (g1572)));
	assign g2134 = (((!ld) & (!sk[23]) & (text_inx22x) & (!g1574)) + ((!ld) & (!sk[23]) & (text_inx22x) & (g1574)) + ((!ld) & (sk[23]) & (!text_inx22x) & (g1574)) + ((!ld) & (sk[23]) & (text_inx22x) & (g1574)) + ((ld) & (!sk[23]) & (!text_inx22x) & (g1574)) + ((ld) & (!sk[23]) & (text_inx22x) & (!g1574)) + ((ld) & (!sk[23]) & (text_inx22x) & (g1574)) + ((ld) & (sk[23]) & (text_inx22x) & (!g1574)) + ((ld) & (sk[23]) & (text_inx22x) & (g1574)));
	assign g1575 = (((!g246) & (!g318) & (!g381) & (!g1163) & (g1423) & (!g1574)) + ((!g246) & (!g318) & (!g381) & (!g1163) & (g1423) & (g1574)) + ((!g246) & (!g318) & (!g381) & (g1163) & (!g1423) & (g1574)) + ((!g246) & (!g318) & (!g381) & (g1163) & (g1423) & (g1574)) + ((!g246) & (!g318) & (g381) & (!g1163) & (!g1423) & (!g1574)) + ((!g246) & (!g318) & (g381) & (!g1163) & (!g1423) & (g1574)) + ((!g246) & (!g318) & (g381) & (g1163) & (!g1423) & (g1574)) + ((!g246) & (!g318) & (g381) & (g1163) & (g1423) & (g1574)) + ((!g246) & (g318) & (!g381) & (!g1163) & (!g1423) & (!g1574)) + ((!g246) & (g318) & (!g381) & (!g1163) & (!g1423) & (g1574)) + ((!g246) & (g318) & (!g381) & (g1163) & (!g1423) & (!g1574)) + ((!g246) & (g318) & (!g381) & (g1163) & (g1423) & (!g1574)) + ((!g246) & (g318) & (g381) & (!g1163) & (g1423) & (!g1574)) + ((!g246) & (g318) & (g381) & (!g1163) & (g1423) & (g1574)) + ((!g246) & (g318) & (g381) & (g1163) & (!g1423) & (!g1574)) + ((!g246) & (g318) & (g381) & (g1163) & (g1423) & (!g1574)) + ((g246) & (!g318) & (!g381) & (!g1163) & (!g1423) & (!g1574)) + ((g246) & (!g318) & (!g381) & (!g1163) & (!g1423) & (g1574)) + ((g246) & (!g318) & (!g381) & (g1163) & (!g1423) & (g1574)) + ((g246) & (!g318) & (!g381) & (g1163) & (g1423) & (g1574)) + ((g246) & (!g318) & (g381) & (!g1163) & (g1423) & (!g1574)) + ((g246) & (!g318) & (g381) & (!g1163) & (g1423) & (g1574)) + ((g246) & (!g318) & (g381) & (g1163) & (!g1423) & (g1574)) + ((g246) & (!g318) & (g381) & (g1163) & (g1423) & (g1574)) + ((g246) & (g318) & (!g381) & (!g1163) & (g1423) & (!g1574)) + ((g246) & (g318) & (!g381) & (!g1163) & (g1423) & (g1574)) + ((g246) & (g318) & (!g381) & (g1163) & (!g1423) & (!g1574)) + ((g246) & (g318) & (!g381) & (g1163) & (g1423) & (!g1574)) + ((g246) & (g318) & (g381) & (!g1163) & (!g1423) & (!g1574)) + ((g246) & (g318) & (g381) & (!g1163) & (!g1423) & (g1574)) + ((g246) & (g318) & (g381) & (g1163) & (!g1423) & (!g1574)) + ((g246) & (g318) & (g381) & (g1163) & (g1423) & (!g1574)));
	assign g2135 = (((!ld) & (!text_inx21x) & (sk[25]) & (g1576)) + ((!ld) & (text_inx21x) & (!sk[25]) & (!g1576)) + ((!ld) & (text_inx21x) & (!sk[25]) & (g1576)) + ((!ld) & (text_inx21x) & (sk[25]) & (g1576)) + ((ld) & (!text_inx21x) & (!sk[25]) & (g1576)) + ((ld) & (text_inx21x) & (!sk[25]) & (!g1576)) + ((ld) & (text_inx21x) & (!sk[25]) & (g1576)) + ((ld) & (text_inx21x) & (sk[25]) & (!g1576)) + ((ld) & (text_inx21x) & (sk[25]) & (g1576)));
	assign g1577 = (((!g239) & (!g311) & (!g374) & (!g1163) & (g1426) & (!g1576)) + ((!g239) & (!g311) & (!g374) & (!g1163) & (g1426) & (g1576)) + ((!g239) & (!g311) & (!g374) & (g1163) & (!g1426) & (g1576)) + ((!g239) & (!g311) & (!g374) & (g1163) & (g1426) & (g1576)) + ((!g239) & (!g311) & (g374) & (!g1163) & (!g1426) & (!g1576)) + ((!g239) & (!g311) & (g374) & (!g1163) & (!g1426) & (g1576)) + ((!g239) & (!g311) & (g374) & (g1163) & (!g1426) & (g1576)) + ((!g239) & (!g311) & (g374) & (g1163) & (g1426) & (g1576)) + ((!g239) & (g311) & (!g374) & (!g1163) & (!g1426) & (!g1576)) + ((!g239) & (g311) & (!g374) & (!g1163) & (!g1426) & (g1576)) + ((!g239) & (g311) & (!g374) & (g1163) & (!g1426) & (!g1576)) + ((!g239) & (g311) & (!g374) & (g1163) & (g1426) & (!g1576)) + ((!g239) & (g311) & (g374) & (!g1163) & (g1426) & (!g1576)) + ((!g239) & (g311) & (g374) & (!g1163) & (g1426) & (g1576)) + ((!g239) & (g311) & (g374) & (g1163) & (!g1426) & (!g1576)) + ((!g239) & (g311) & (g374) & (g1163) & (g1426) & (!g1576)) + ((g239) & (!g311) & (!g374) & (!g1163) & (!g1426) & (!g1576)) + ((g239) & (!g311) & (!g374) & (!g1163) & (!g1426) & (g1576)) + ((g239) & (!g311) & (!g374) & (g1163) & (!g1426) & (g1576)) + ((g239) & (!g311) & (!g374) & (g1163) & (g1426) & (g1576)) + ((g239) & (!g311) & (g374) & (!g1163) & (g1426) & (!g1576)) + ((g239) & (!g311) & (g374) & (!g1163) & (g1426) & (g1576)) + ((g239) & (!g311) & (g374) & (g1163) & (!g1426) & (g1576)) + ((g239) & (!g311) & (g374) & (g1163) & (g1426) & (g1576)) + ((g239) & (g311) & (!g374) & (!g1163) & (g1426) & (!g1576)) + ((g239) & (g311) & (!g374) & (!g1163) & (g1426) & (g1576)) + ((g239) & (g311) & (!g374) & (g1163) & (!g1426) & (!g1576)) + ((g239) & (g311) & (!g374) & (g1163) & (g1426) & (!g1576)) + ((g239) & (g311) & (g374) & (!g1163) & (!g1426) & (!g1576)) + ((g239) & (g311) & (g374) & (!g1163) & (!g1426) & (g1576)) + ((g239) & (g311) & (g374) & (g1163) & (!g1426) & (!g1576)) + ((g239) & (g311) & (g374) & (g1163) & (g1426) & (!g1576)));
	assign g2136 = (((!ld) & (!sk[27]) & (text_inx20x) & (!g1578)) + ((!ld) & (!sk[27]) & (text_inx20x) & (g1578)) + ((!ld) & (sk[27]) & (!text_inx20x) & (g1578)) + ((!ld) & (sk[27]) & (text_inx20x) & (g1578)) + ((ld) & (!sk[27]) & (!text_inx20x) & (g1578)) + ((ld) & (!sk[27]) & (text_inx20x) & (!g1578)) + ((ld) & (!sk[27]) & (text_inx20x) & (g1578)) + ((ld) & (sk[27]) & (text_inx20x) & (!g1578)) + ((ld) & (sk[27]) & (text_inx20x) & (g1578)));
	assign g2137 = (((!sk[28]) & (!ld) & (text_inx23x) & (!g1579)) + ((!sk[28]) & (!ld) & (text_inx23x) & (g1579)) + ((!sk[28]) & (ld) & (!text_inx23x) & (g1579)) + ((!sk[28]) & (ld) & (text_inx23x) & (!g1579)) + ((!sk[28]) & (ld) & (text_inx23x) & (g1579)) + ((sk[28]) & (!ld) & (!text_inx23x) & (g1579)) + ((sk[28]) & (!ld) & (text_inx23x) & (g1579)) + ((sk[28]) & (ld) & (text_inx23x) & (!g1579)) + ((sk[28]) & (ld) & (text_inx23x) & (g1579)));
	assign g1580 = (((!ld) & (!g532) & (!g788) & (!g1044) & (g1358) & (!keyx48x)) + ((!ld) & (!g532) & (!g788) & (!g1044) & (g1358) & (keyx48x)) + ((!ld) & (!g532) & (!g788) & (g1044) & (!g1358) & (!keyx48x)) + ((!ld) & (!g532) & (!g788) & (g1044) & (!g1358) & (keyx48x)) + ((!ld) & (!g532) & (g788) & (!g1044) & (!g1358) & (!keyx48x)) + ((!ld) & (!g532) & (g788) & (!g1044) & (!g1358) & (keyx48x)) + ((!ld) & (!g532) & (g788) & (g1044) & (g1358) & (!keyx48x)) + ((!ld) & (!g532) & (g788) & (g1044) & (g1358) & (keyx48x)) + ((!ld) & (g532) & (!g788) & (!g1044) & (!g1358) & (!keyx48x)) + ((!ld) & (g532) & (!g788) & (!g1044) & (!g1358) & (keyx48x)) + ((!ld) & (g532) & (!g788) & (g1044) & (g1358) & (!keyx48x)) + ((!ld) & (g532) & (!g788) & (g1044) & (g1358) & (keyx48x)) + ((!ld) & (g532) & (g788) & (!g1044) & (g1358) & (!keyx48x)) + ((!ld) & (g532) & (g788) & (!g1044) & (g1358) & (keyx48x)) + ((!ld) & (g532) & (g788) & (g1044) & (!g1358) & (!keyx48x)) + ((!ld) & (g532) & (g788) & (g1044) & (!g1358) & (keyx48x)) + ((ld) & (!g532) & (!g788) & (!g1044) & (!g1358) & (keyx48x)) + ((ld) & (!g532) & (!g788) & (!g1044) & (g1358) & (keyx48x)) + ((ld) & (!g532) & (!g788) & (g1044) & (!g1358) & (keyx48x)) + ((ld) & (!g532) & (!g788) & (g1044) & (g1358) & (keyx48x)) + ((ld) & (!g532) & (g788) & (!g1044) & (!g1358) & (keyx48x)) + ((ld) & (!g532) & (g788) & (!g1044) & (g1358) & (keyx48x)) + ((ld) & (!g532) & (g788) & (g1044) & (!g1358) & (keyx48x)) + ((ld) & (!g532) & (g788) & (g1044) & (g1358) & (keyx48x)) + ((ld) & (g532) & (!g788) & (!g1044) & (!g1358) & (keyx48x)) + ((ld) & (g532) & (!g788) & (!g1044) & (g1358) & (keyx48x)) + ((ld) & (g532) & (!g788) & (g1044) & (!g1358) & (keyx48x)) + ((ld) & (g532) & (!g788) & (g1044) & (g1358) & (keyx48x)) + ((ld) & (g532) & (g788) & (!g1044) & (!g1358) & (keyx48x)) + ((ld) & (g532) & (g788) & (!g1044) & (g1358) & (keyx48x)) + ((ld) & (g532) & (g788) & (g1044) & (!g1358) & (keyx48x)) + ((ld) & (g532) & (g788) & (g1044) & (g1358) & (keyx48x)));
	assign g1581 = (((!ld) & (!g539) & (!g795) & (!g1051) & (g1365) & (!keyx49x)) + ((!ld) & (!g539) & (!g795) & (!g1051) & (g1365) & (keyx49x)) + ((!ld) & (!g539) & (!g795) & (g1051) & (!g1365) & (!keyx49x)) + ((!ld) & (!g539) & (!g795) & (g1051) & (!g1365) & (keyx49x)) + ((!ld) & (!g539) & (g795) & (!g1051) & (!g1365) & (!keyx49x)) + ((!ld) & (!g539) & (g795) & (!g1051) & (!g1365) & (keyx49x)) + ((!ld) & (!g539) & (g795) & (g1051) & (g1365) & (!keyx49x)) + ((!ld) & (!g539) & (g795) & (g1051) & (g1365) & (keyx49x)) + ((!ld) & (g539) & (!g795) & (!g1051) & (!g1365) & (!keyx49x)) + ((!ld) & (g539) & (!g795) & (!g1051) & (!g1365) & (keyx49x)) + ((!ld) & (g539) & (!g795) & (g1051) & (g1365) & (!keyx49x)) + ((!ld) & (g539) & (!g795) & (g1051) & (g1365) & (keyx49x)) + ((!ld) & (g539) & (g795) & (!g1051) & (g1365) & (!keyx49x)) + ((!ld) & (g539) & (g795) & (!g1051) & (g1365) & (keyx49x)) + ((!ld) & (g539) & (g795) & (g1051) & (!g1365) & (!keyx49x)) + ((!ld) & (g539) & (g795) & (g1051) & (!g1365) & (keyx49x)) + ((ld) & (!g539) & (!g795) & (!g1051) & (!g1365) & (keyx49x)) + ((ld) & (!g539) & (!g795) & (!g1051) & (g1365) & (keyx49x)) + ((ld) & (!g539) & (!g795) & (g1051) & (!g1365) & (keyx49x)) + ((ld) & (!g539) & (!g795) & (g1051) & (g1365) & (keyx49x)) + ((ld) & (!g539) & (g795) & (!g1051) & (!g1365) & (keyx49x)) + ((ld) & (!g539) & (g795) & (!g1051) & (g1365) & (keyx49x)) + ((ld) & (!g539) & (g795) & (g1051) & (!g1365) & (keyx49x)) + ((ld) & (!g539) & (g795) & (g1051) & (g1365) & (keyx49x)) + ((ld) & (g539) & (!g795) & (!g1051) & (!g1365) & (keyx49x)) + ((ld) & (g539) & (!g795) & (!g1051) & (g1365) & (keyx49x)) + ((ld) & (g539) & (!g795) & (g1051) & (!g1365) & (keyx49x)) + ((ld) & (g539) & (!g795) & (g1051) & (g1365) & (keyx49x)) + ((ld) & (g539) & (g795) & (!g1051) & (!g1365) & (keyx49x)) + ((ld) & (g539) & (g795) & (!g1051) & (g1365) & (keyx49x)) + ((ld) & (g539) & (g795) & (g1051) & (!g1365) & (keyx49x)) + ((ld) & (g539) & (g795) & (g1051) & (g1365) & (keyx49x)));
	assign g1582 = (((!ld) & (!g546) & (!g802) & (!g1058) & (g1372) & (!keyx50x)) + ((!ld) & (!g546) & (!g802) & (!g1058) & (g1372) & (keyx50x)) + ((!ld) & (!g546) & (!g802) & (g1058) & (!g1372) & (!keyx50x)) + ((!ld) & (!g546) & (!g802) & (g1058) & (!g1372) & (keyx50x)) + ((!ld) & (!g546) & (g802) & (!g1058) & (!g1372) & (!keyx50x)) + ((!ld) & (!g546) & (g802) & (!g1058) & (!g1372) & (keyx50x)) + ((!ld) & (!g546) & (g802) & (g1058) & (g1372) & (!keyx50x)) + ((!ld) & (!g546) & (g802) & (g1058) & (g1372) & (keyx50x)) + ((!ld) & (g546) & (!g802) & (!g1058) & (!g1372) & (!keyx50x)) + ((!ld) & (g546) & (!g802) & (!g1058) & (!g1372) & (keyx50x)) + ((!ld) & (g546) & (!g802) & (g1058) & (g1372) & (!keyx50x)) + ((!ld) & (g546) & (!g802) & (g1058) & (g1372) & (keyx50x)) + ((!ld) & (g546) & (g802) & (!g1058) & (g1372) & (!keyx50x)) + ((!ld) & (g546) & (g802) & (!g1058) & (g1372) & (keyx50x)) + ((!ld) & (g546) & (g802) & (g1058) & (!g1372) & (!keyx50x)) + ((!ld) & (g546) & (g802) & (g1058) & (!g1372) & (keyx50x)) + ((ld) & (!g546) & (!g802) & (!g1058) & (!g1372) & (keyx50x)) + ((ld) & (!g546) & (!g802) & (!g1058) & (g1372) & (keyx50x)) + ((ld) & (!g546) & (!g802) & (g1058) & (!g1372) & (keyx50x)) + ((ld) & (!g546) & (!g802) & (g1058) & (g1372) & (keyx50x)) + ((ld) & (!g546) & (g802) & (!g1058) & (!g1372) & (keyx50x)) + ((ld) & (!g546) & (g802) & (!g1058) & (g1372) & (keyx50x)) + ((ld) & (!g546) & (g802) & (g1058) & (!g1372) & (keyx50x)) + ((ld) & (!g546) & (g802) & (g1058) & (g1372) & (keyx50x)) + ((ld) & (g546) & (!g802) & (!g1058) & (!g1372) & (keyx50x)) + ((ld) & (g546) & (!g802) & (!g1058) & (g1372) & (keyx50x)) + ((ld) & (g546) & (!g802) & (g1058) & (!g1372) & (keyx50x)) + ((ld) & (g546) & (!g802) & (g1058) & (g1372) & (keyx50x)) + ((ld) & (g546) & (g802) & (!g1058) & (!g1372) & (keyx50x)) + ((ld) & (g546) & (g802) & (!g1058) & (g1372) & (keyx50x)) + ((ld) & (g546) & (g802) & (g1058) & (!g1372) & (keyx50x)) + ((ld) & (g546) & (g802) & (g1058) & (g1372) & (keyx50x)));
	assign g1583 = (((!ld) & (!g553) & (!g809) & (!g1065) & (g1379) & (!keyx51x)) + ((!ld) & (!g553) & (!g809) & (!g1065) & (g1379) & (keyx51x)) + ((!ld) & (!g553) & (!g809) & (g1065) & (!g1379) & (!keyx51x)) + ((!ld) & (!g553) & (!g809) & (g1065) & (!g1379) & (keyx51x)) + ((!ld) & (!g553) & (g809) & (!g1065) & (!g1379) & (!keyx51x)) + ((!ld) & (!g553) & (g809) & (!g1065) & (!g1379) & (keyx51x)) + ((!ld) & (!g553) & (g809) & (g1065) & (g1379) & (!keyx51x)) + ((!ld) & (!g553) & (g809) & (g1065) & (g1379) & (keyx51x)) + ((!ld) & (g553) & (!g809) & (!g1065) & (!g1379) & (!keyx51x)) + ((!ld) & (g553) & (!g809) & (!g1065) & (!g1379) & (keyx51x)) + ((!ld) & (g553) & (!g809) & (g1065) & (g1379) & (!keyx51x)) + ((!ld) & (g553) & (!g809) & (g1065) & (g1379) & (keyx51x)) + ((!ld) & (g553) & (g809) & (!g1065) & (g1379) & (!keyx51x)) + ((!ld) & (g553) & (g809) & (!g1065) & (g1379) & (keyx51x)) + ((!ld) & (g553) & (g809) & (g1065) & (!g1379) & (!keyx51x)) + ((!ld) & (g553) & (g809) & (g1065) & (!g1379) & (keyx51x)) + ((ld) & (!g553) & (!g809) & (!g1065) & (!g1379) & (keyx51x)) + ((ld) & (!g553) & (!g809) & (!g1065) & (g1379) & (keyx51x)) + ((ld) & (!g553) & (!g809) & (g1065) & (!g1379) & (keyx51x)) + ((ld) & (!g553) & (!g809) & (g1065) & (g1379) & (keyx51x)) + ((ld) & (!g553) & (g809) & (!g1065) & (!g1379) & (keyx51x)) + ((ld) & (!g553) & (g809) & (!g1065) & (g1379) & (keyx51x)) + ((ld) & (!g553) & (g809) & (g1065) & (!g1379) & (keyx51x)) + ((ld) & (!g553) & (g809) & (g1065) & (g1379) & (keyx51x)) + ((ld) & (g553) & (!g809) & (!g1065) & (!g1379) & (keyx51x)) + ((ld) & (g553) & (!g809) & (!g1065) & (g1379) & (keyx51x)) + ((ld) & (g553) & (!g809) & (g1065) & (!g1379) & (keyx51x)) + ((ld) & (g553) & (!g809) & (g1065) & (g1379) & (keyx51x)) + ((ld) & (g553) & (g809) & (!g1065) & (!g1379) & (keyx51x)) + ((ld) & (g553) & (g809) & (!g1065) & (g1379) & (keyx51x)) + ((ld) & (g553) & (g809) & (g1065) & (!g1379) & (keyx51x)) + ((ld) & (g553) & (g809) & (g1065) & (g1379) & (keyx51x)));
	assign g1584 = (((!ld) & (!g560) & (!g816) & (!g1072) & (g1386) & (!keyx52x)) + ((!ld) & (!g560) & (!g816) & (!g1072) & (g1386) & (keyx52x)) + ((!ld) & (!g560) & (!g816) & (g1072) & (!g1386) & (!keyx52x)) + ((!ld) & (!g560) & (!g816) & (g1072) & (!g1386) & (keyx52x)) + ((!ld) & (!g560) & (g816) & (!g1072) & (!g1386) & (!keyx52x)) + ((!ld) & (!g560) & (g816) & (!g1072) & (!g1386) & (keyx52x)) + ((!ld) & (!g560) & (g816) & (g1072) & (g1386) & (!keyx52x)) + ((!ld) & (!g560) & (g816) & (g1072) & (g1386) & (keyx52x)) + ((!ld) & (g560) & (!g816) & (!g1072) & (!g1386) & (!keyx52x)) + ((!ld) & (g560) & (!g816) & (!g1072) & (!g1386) & (keyx52x)) + ((!ld) & (g560) & (!g816) & (g1072) & (g1386) & (!keyx52x)) + ((!ld) & (g560) & (!g816) & (g1072) & (g1386) & (keyx52x)) + ((!ld) & (g560) & (g816) & (!g1072) & (g1386) & (!keyx52x)) + ((!ld) & (g560) & (g816) & (!g1072) & (g1386) & (keyx52x)) + ((!ld) & (g560) & (g816) & (g1072) & (!g1386) & (!keyx52x)) + ((!ld) & (g560) & (g816) & (g1072) & (!g1386) & (keyx52x)) + ((ld) & (!g560) & (!g816) & (!g1072) & (!g1386) & (keyx52x)) + ((ld) & (!g560) & (!g816) & (!g1072) & (g1386) & (keyx52x)) + ((ld) & (!g560) & (!g816) & (g1072) & (!g1386) & (keyx52x)) + ((ld) & (!g560) & (!g816) & (g1072) & (g1386) & (keyx52x)) + ((ld) & (!g560) & (g816) & (!g1072) & (!g1386) & (keyx52x)) + ((ld) & (!g560) & (g816) & (!g1072) & (g1386) & (keyx52x)) + ((ld) & (!g560) & (g816) & (g1072) & (!g1386) & (keyx52x)) + ((ld) & (!g560) & (g816) & (g1072) & (g1386) & (keyx52x)) + ((ld) & (g560) & (!g816) & (!g1072) & (!g1386) & (keyx52x)) + ((ld) & (g560) & (!g816) & (!g1072) & (g1386) & (keyx52x)) + ((ld) & (g560) & (!g816) & (g1072) & (!g1386) & (keyx52x)) + ((ld) & (g560) & (!g816) & (g1072) & (g1386) & (keyx52x)) + ((ld) & (g560) & (g816) & (!g1072) & (!g1386) & (keyx52x)) + ((ld) & (g560) & (g816) & (!g1072) & (g1386) & (keyx52x)) + ((ld) & (g560) & (g816) & (g1072) & (!g1386) & (keyx52x)) + ((ld) & (g560) & (g816) & (g1072) & (g1386) & (keyx52x)));
	assign g1585 = (((!ld) & (!g567) & (!g823) & (!g1079) & (g1393) & (!keyx53x)) + ((!ld) & (!g567) & (!g823) & (!g1079) & (g1393) & (keyx53x)) + ((!ld) & (!g567) & (!g823) & (g1079) & (!g1393) & (!keyx53x)) + ((!ld) & (!g567) & (!g823) & (g1079) & (!g1393) & (keyx53x)) + ((!ld) & (!g567) & (g823) & (!g1079) & (!g1393) & (!keyx53x)) + ((!ld) & (!g567) & (g823) & (!g1079) & (!g1393) & (keyx53x)) + ((!ld) & (!g567) & (g823) & (g1079) & (g1393) & (!keyx53x)) + ((!ld) & (!g567) & (g823) & (g1079) & (g1393) & (keyx53x)) + ((!ld) & (g567) & (!g823) & (!g1079) & (!g1393) & (!keyx53x)) + ((!ld) & (g567) & (!g823) & (!g1079) & (!g1393) & (keyx53x)) + ((!ld) & (g567) & (!g823) & (g1079) & (g1393) & (!keyx53x)) + ((!ld) & (g567) & (!g823) & (g1079) & (g1393) & (keyx53x)) + ((!ld) & (g567) & (g823) & (!g1079) & (g1393) & (!keyx53x)) + ((!ld) & (g567) & (g823) & (!g1079) & (g1393) & (keyx53x)) + ((!ld) & (g567) & (g823) & (g1079) & (!g1393) & (!keyx53x)) + ((!ld) & (g567) & (g823) & (g1079) & (!g1393) & (keyx53x)) + ((ld) & (!g567) & (!g823) & (!g1079) & (!g1393) & (keyx53x)) + ((ld) & (!g567) & (!g823) & (!g1079) & (g1393) & (keyx53x)) + ((ld) & (!g567) & (!g823) & (g1079) & (!g1393) & (keyx53x)) + ((ld) & (!g567) & (!g823) & (g1079) & (g1393) & (keyx53x)) + ((ld) & (!g567) & (g823) & (!g1079) & (!g1393) & (keyx53x)) + ((ld) & (!g567) & (g823) & (!g1079) & (g1393) & (keyx53x)) + ((ld) & (!g567) & (g823) & (g1079) & (!g1393) & (keyx53x)) + ((ld) & (!g567) & (g823) & (g1079) & (g1393) & (keyx53x)) + ((ld) & (g567) & (!g823) & (!g1079) & (!g1393) & (keyx53x)) + ((ld) & (g567) & (!g823) & (!g1079) & (g1393) & (keyx53x)) + ((ld) & (g567) & (!g823) & (g1079) & (!g1393) & (keyx53x)) + ((ld) & (g567) & (!g823) & (g1079) & (g1393) & (keyx53x)) + ((ld) & (g567) & (g823) & (!g1079) & (!g1393) & (keyx53x)) + ((ld) & (g567) & (g823) & (!g1079) & (g1393) & (keyx53x)) + ((ld) & (g567) & (g823) & (g1079) & (!g1393) & (keyx53x)) + ((ld) & (g567) & (g823) & (g1079) & (g1393) & (keyx53x)));
	assign g1586 = (((!ld) & (!g574) & (!g830) & (!g1086) & (g1400) & (!keyx54x)) + ((!ld) & (!g574) & (!g830) & (!g1086) & (g1400) & (keyx54x)) + ((!ld) & (!g574) & (!g830) & (g1086) & (!g1400) & (!keyx54x)) + ((!ld) & (!g574) & (!g830) & (g1086) & (!g1400) & (keyx54x)) + ((!ld) & (!g574) & (g830) & (!g1086) & (!g1400) & (!keyx54x)) + ((!ld) & (!g574) & (g830) & (!g1086) & (!g1400) & (keyx54x)) + ((!ld) & (!g574) & (g830) & (g1086) & (g1400) & (!keyx54x)) + ((!ld) & (!g574) & (g830) & (g1086) & (g1400) & (keyx54x)) + ((!ld) & (g574) & (!g830) & (!g1086) & (!g1400) & (!keyx54x)) + ((!ld) & (g574) & (!g830) & (!g1086) & (!g1400) & (keyx54x)) + ((!ld) & (g574) & (!g830) & (g1086) & (g1400) & (!keyx54x)) + ((!ld) & (g574) & (!g830) & (g1086) & (g1400) & (keyx54x)) + ((!ld) & (g574) & (g830) & (!g1086) & (g1400) & (!keyx54x)) + ((!ld) & (g574) & (g830) & (!g1086) & (g1400) & (keyx54x)) + ((!ld) & (g574) & (g830) & (g1086) & (!g1400) & (!keyx54x)) + ((!ld) & (g574) & (g830) & (g1086) & (!g1400) & (keyx54x)) + ((ld) & (!g574) & (!g830) & (!g1086) & (!g1400) & (keyx54x)) + ((ld) & (!g574) & (!g830) & (!g1086) & (g1400) & (keyx54x)) + ((ld) & (!g574) & (!g830) & (g1086) & (!g1400) & (keyx54x)) + ((ld) & (!g574) & (!g830) & (g1086) & (g1400) & (keyx54x)) + ((ld) & (!g574) & (g830) & (!g1086) & (!g1400) & (keyx54x)) + ((ld) & (!g574) & (g830) & (!g1086) & (g1400) & (keyx54x)) + ((ld) & (!g574) & (g830) & (g1086) & (!g1400) & (keyx54x)) + ((ld) & (!g574) & (g830) & (g1086) & (g1400) & (keyx54x)) + ((ld) & (g574) & (!g830) & (!g1086) & (!g1400) & (keyx54x)) + ((ld) & (g574) & (!g830) & (!g1086) & (g1400) & (keyx54x)) + ((ld) & (g574) & (!g830) & (g1086) & (!g1400) & (keyx54x)) + ((ld) & (g574) & (!g830) & (g1086) & (g1400) & (keyx54x)) + ((ld) & (g574) & (g830) & (!g1086) & (!g1400) & (keyx54x)) + ((ld) & (g574) & (g830) & (!g1086) & (g1400) & (keyx54x)) + ((ld) & (g574) & (g830) & (g1086) & (!g1400) & (keyx54x)) + ((ld) & (g574) & (g830) & (g1086) & (g1400) & (keyx54x)));
	assign g1587 = (((!ld) & (!g581) & (!g837) & (!g1093) & (g1407) & (!keyx55x)) + ((!ld) & (!g581) & (!g837) & (!g1093) & (g1407) & (keyx55x)) + ((!ld) & (!g581) & (!g837) & (g1093) & (!g1407) & (!keyx55x)) + ((!ld) & (!g581) & (!g837) & (g1093) & (!g1407) & (keyx55x)) + ((!ld) & (!g581) & (g837) & (!g1093) & (!g1407) & (!keyx55x)) + ((!ld) & (!g581) & (g837) & (!g1093) & (!g1407) & (keyx55x)) + ((!ld) & (!g581) & (g837) & (g1093) & (g1407) & (!keyx55x)) + ((!ld) & (!g581) & (g837) & (g1093) & (g1407) & (keyx55x)) + ((!ld) & (g581) & (!g837) & (!g1093) & (!g1407) & (!keyx55x)) + ((!ld) & (g581) & (!g837) & (!g1093) & (!g1407) & (keyx55x)) + ((!ld) & (g581) & (!g837) & (g1093) & (g1407) & (!keyx55x)) + ((!ld) & (g581) & (!g837) & (g1093) & (g1407) & (keyx55x)) + ((!ld) & (g581) & (g837) & (!g1093) & (g1407) & (!keyx55x)) + ((!ld) & (g581) & (g837) & (!g1093) & (g1407) & (keyx55x)) + ((!ld) & (g581) & (g837) & (g1093) & (!g1407) & (!keyx55x)) + ((!ld) & (g581) & (g837) & (g1093) & (!g1407) & (keyx55x)) + ((ld) & (!g581) & (!g837) & (!g1093) & (!g1407) & (keyx55x)) + ((ld) & (!g581) & (!g837) & (!g1093) & (g1407) & (keyx55x)) + ((ld) & (!g581) & (!g837) & (g1093) & (!g1407) & (keyx55x)) + ((ld) & (!g581) & (!g837) & (g1093) & (g1407) & (keyx55x)) + ((ld) & (!g581) & (g837) & (!g1093) & (!g1407) & (keyx55x)) + ((ld) & (!g581) & (g837) & (!g1093) & (g1407) & (keyx55x)) + ((ld) & (!g581) & (g837) & (g1093) & (!g1407) & (keyx55x)) + ((ld) & (!g581) & (g837) & (g1093) & (g1407) & (keyx55x)) + ((ld) & (g581) & (!g837) & (!g1093) & (!g1407) & (keyx55x)) + ((ld) & (g581) & (!g837) & (!g1093) & (g1407) & (keyx55x)) + ((ld) & (g581) & (!g837) & (g1093) & (!g1407) & (keyx55x)) + ((ld) & (g581) & (!g837) & (g1093) & (g1407) & (keyx55x)) + ((ld) & (g581) & (g837) & (!g1093) & (!g1407) & (keyx55x)) + ((ld) & (g581) & (g837) & (!g1093) & (g1407) & (keyx55x)) + ((ld) & (g581) & (g837) & (g1093) & (!g1407) & (keyx55x)) + ((ld) & (g581) & (g837) & (g1093) & (g1407) & (keyx55x)));
	assign g2138 = (((!ld) & (!sk[37]) & (text_inx56x) & (!g1588)) + ((!ld) & (!sk[37]) & (text_inx56x) & (g1588)) + ((!ld) & (sk[37]) & (!text_inx56x) & (g1588)) + ((!ld) & (sk[37]) & (text_inx56x) & (g1588)) + ((ld) & (!sk[37]) & (!text_inx56x) & (g1588)) + ((ld) & (!sk[37]) & (text_inx56x) & (!g1588)) + ((ld) & (!sk[37]) & (text_inx56x) & (g1588)) + ((ld) & (sk[37]) & (text_inx56x) & (!g1588)) + ((ld) & (sk[37]) & (text_inx56x) & (g1588)));
	assign g1589 = (((!g531) & (!sk[38]) & (g580) & (!g644)) + ((!g531) & (!sk[38]) & (g580) & (g644)) + ((!g531) & (sk[38]) & (!g580) & (g644)) + ((!g531) & (sk[38]) & (g580) & (!g644)) + ((g531) & (!sk[38]) & (!g580) & (g644)) + ((g531) & (!sk[38]) & (g580) & (!g644)) + ((g531) & (!sk[38]) & (g580) & (g644)) + ((g531) & (sk[38]) & (!g580) & (!g644)) + ((g531) & (sk[38]) & (g580) & (g644)));
	assign g1590 = (((!g403) & (!g467) & (!g596) & (!g1163) & (!g1588) & (g1589)) + ((!g403) & (!g467) & (!g596) & (!g1163) & (g1588) & (g1589)) + ((!g403) & (!g467) & (!g596) & (g1163) & (g1588) & (!g1589)) + ((!g403) & (!g467) & (!g596) & (g1163) & (g1588) & (g1589)) + ((!g403) & (!g467) & (g596) & (!g1163) & (!g1588) & (!g1589)) + ((!g403) & (!g467) & (g596) & (!g1163) & (g1588) & (!g1589)) + ((!g403) & (!g467) & (g596) & (g1163) & (!g1588) & (!g1589)) + ((!g403) & (!g467) & (g596) & (g1163) & (!g1588) & (g1589)) + ((!g403) & (g467) & (!g596) & (!g1163) & (!g1588) & (!g1589)) + ((!g403) & (g467) & (!g596) & (!g1163) & (g1588) & (!g1589)) + ((!g403) & (g467) & (!g596) & (g1163) & (g1588) & (!g1589)) + ((!g403) & (g467) & (!g596) & (g1163) & (g1588) & (g1589)) + ((!g403) & (g467) & (g596) & (!g1163) & (!g1588) & (g1589)) + ((!g403) & (g467) & (g596) & (!g1163) & (g1588) & (g1589)) + ((!g403) & (g467) & (g596) & (g1163) & (!g1588) & (!g1589)) + ((!g403) & (g467) & (g596) & (g1163) & (!g1588) & (g1589)) + ((g403) & (!g467) & (!g596) & (!g1163) & (!g1588) & (!g1589)) + ((g403) & (!g467) & (!g596) & (!g1163) & (g1588) & (!g1589)) + ((g403) & (!g467) & (!g596) & (g1163) & (g1588) & (!g1589)) + ((g403) & (!g467) & (!g596) & (g1163) & (g1588) & (g1589)) + ((g403) & (!g467) & (g596) & (!g1163) & (!g1588) & (g1589)) + ((g403) & (!g467) & (g596) & (!g1163) & (g1588) & (g1589)) + ((g403) & (!g467) & (g596) & (g1163) & (!g1588) & (!g1589)) + ((g403) & (!g467) & (g596) & (g1163) & (!g1588) & (g1589)) + ((g403) & (g467) & (!g596) & (!g1163) & (!g1588) & (g1589)) + ((g403) & (g467) & (!g596) & (!g1163) & (g1588) & (g1589)) + ((g403) & (g467) & (!g596) & (g1163) & (g1588) & (!g1589)) + ((g403) & (g467) & (!g596) & (g1163) & (g1588) & (g1589)) + ((g403) & (g467) & (g596) & (!g1163) & (!g1588) & (!g1589)) + ((g403) & (g467) & (g596) & (!g1163) & (g1588) & (!g1589)) + ((g403) & (g467) & (g596) & (g1163) & (!g1588) & (!g1589)) + ((g403) & (g467) & (g596) & (g1163) & (!g1588) & (g1589)));
	assign g2139 = (((!ld) & (!sk[40]) & (text_inx57x) & (!g1591)) + ((!ld) & (!sk[40]) & (text_inx57x) & (g1591)) + ((!ld) & (sk[40]) & (!text_inx57x) & (g1591)) + ((!ld) & (sk[40]) & (text_inx57x) & (g1591)) + ((ld) & (!sk[40]) & (!text_inx57x) & (g1591)) + ((ld) & (!sk[40]) & (text_inx57x) & (!g1591)) + ((ld) & (!sk[40]) & (text_inx57x) & (g1591)) + ((ld) & (sk[40]) & (text_inx57x) & (!g1591)) + ((ld) & (sk[40]) & (text_inx57x) & (g1591)));
	assign g1592 = (((!g410) & (!g603) & (!g1163) & (!g1168) & (g1589) & (!g1591)) + ((!g410) & (!g603) & (!g1163) & (!g1168) & (g1589) & (g1591)) + ((!g410) & (!g603) & (!g1163) & (g1168) & (!g1589) & (!g1591)) + ((!g410) & (!g603) & (!g1163) & (g1168) & (!g1589) & (g1591)) + ((!g410) & (!g603) & (g1163) & (!g1168) & (!g1589) & (g1591)) + ((!g410) & (!g603) & (g1163) & (!g1168) & (g1589) & (g1591)) + ((!g410) & (!g603) & (g1163) & (g1168) & (!g1589) & (g1591)) + ((!g410) & (!g603) & (g1163) & (g1168) & (g1589) & (g1591)) + ((!g410) & (g603) & (!g1163) & (!g1168) & (!g1589) & (!g1591)) + ((!g410) & (g603) & (!g1163) & (!g1168) & (!g1589) & (g1591)) + ((!g410) & (g603) & (!g1163) & (g1168) & (g1589) & (!g1591)) + ((!g410) & (g603) & (!g1163) & (g1168) & (g1589) & (g1591)) + ((!g410) & (g603) & (g1163) & (!g1168) & (!g1589) & (!g1591)) + ((!g410) & (g603) & (g1163) & (!g1168) & (g1589) & (!g1591)) + ((!g410) & (g603) & (g1163) & (g1168) & (!g1589) & (!g1591)) + ((!g410) & (g603) & (g1163) & (g1168) & (g1589) & (!g1591)) + ((g410) & (!g603) & (!g1163) & (!g1168) & (!g1589) & (!g1591)) + ((g410) & (!g603) & (!g1163) & (!g1168) & (!g1589) & (g1591)) + ((g410) & (!g603) & (!g1163) & (g1168) & (g1589) & (!g1591)) + ((g410) & (!g603) & (!g1163) & (g1168) & (g1589) & (g1591)) + ((g410) & (!g603) & (g1163) & (!g1168) & (!g1589) & (g1591)) + ((g410) & (!g603) & (g1163) & (!g1168) & (g1589) & (g1591)) + ((g410) & (!g603) & (g1163) & (g1168) & (!g1589) & (g1591)) + ((g410) & (!g603) & (g1163) & (g1168) & (g1589) & (g1591)) + ((g410) & (g603) & (!g1163) & (!g1168) & (g1589) & (!g1591)) + ((g410) & (g603) & (!g1163) & (!g1168) & (g1589) & (g1591)) + ((g410) & (g603) & (!g1163) & (g1168) & (!g1589) & (!g1591)) + ((g410) & (g603) & (!g1163) & (g1168) & (!g1589) & (g1591)) + ((g410) & (g603) & (g1163) & (!g1168) & (!g1589) & (!g1591)) + ((g410) & (g603) & (g1163) & (!g1168) & (g1589) & (!g1591)) + ((g410) & (g603) & (g1163) & (g1168) & (!g1589) & (!g1591)) + ((g410) & (g603) & (g1163) & (g1168) & (g1589) & (!g1591)));
	assign g2140 = (((!ld) & (!sk[42]) & (text_inx58x) & (!g1593)) + ((!ld) & (!sk[42]) & (text_inx58x) & (g1593)) + ((!ld) & (sk[42]) & (!text_inx58x) & (g1593)) + ((!ld) & (sk[42]) & (text_inx58x) & (g1593)) + ((ld) & (!sk[42]) & (!text_inx58x) & (g1593)) + ((ld) & (!sk[42]) & (text_inx58x) & (!g1593)) + ((ld) & (!sk[42]) & (text_inx58x) & (g1593)) + ((ld) & (sk[42]) & (text_inx58x) & (!g1593)) + ((ld) & (sk[42]) & (text_inx58x) & (g1593)));
	assign g1594 = (((!sk[43]) & (!g417) & (g481) & (!g538)) + ((!sk[43]) & (!g417) & (g481) & (g538)) + ((!sk[43]) & (g417) & (!g481) & (g538)) + ((!sk[43]) & (g417) & (g481) & (!g538)) + ((!sk[43]) & (g417) & (g481) & (g538)) + ((sk[43]) & (!g417) & (!g481) & (g538)) + ((sk[43]) & (!g417) & (g481) & (!g538)) + ((sk[43]) & (g417) & (!g481) & (!g538)) + ((sk[43]) & (g417) & (g481) & (g538)));
	assign g1595 = (((!g545) & (!g602) & (!g610) & (!g1163) & (!g1593) & (g1594)) + ((!g545) & (!g602) & (!g610) & (!g1163) & (g1593) & (g1594)) + ((!g545) & (!g602) & (!g610) & (g1163) & (g1593) & (!g1594)) + ((!g545) & (!g602) & (!g610) & (g1163) & (g1593) & (g1594)) + ((!g545) & (!g602) & (g610) & (!g1163) & (!g1593) & (!g1594)) + ((!g545) & (!g602) & (g610) & (!g1163) & (g1593) & (!g1594)) + ((!g545) & (!g602) & (g610) & (g1163) & (!g1593) & (!g1594)) + ((!g545) & (!g602) & (g610) & (g1163) & (!g1593) & (g1594)) + ((!g545) & (g602) & (!g610) & (!g1163) & (!g1593) & (!g1594)) + ((!g545) & (g602) & (!g610) & (!g1163) & (g1593) & (!g1594)) + ((!g545) & (g602) & (!g610) & (g1163) & (g1593) & (!g1594)) + ((!g545) & (g602) & (!g610) & (g1163) & (g1593) & (g1594)) + ((!g545) & (g602) & (g610) & (!g1163) & (!g1593) & (g1594)) + ((!g545) & (g602) & (g610) & (!g1163) & (g1593) & (g1594)) + ((!g545) & (g602) & (g610) & (g1163) & (!g1593) & (!g1594)) + ((!g545) & (g602) & (g610) & (g1163) & (!g1593) & (g1594)) + ((g545) & (!g602) & (!g610) & (!g1163) & (!g1593) & (!g1594)) + ((g545) & (!g602) & (!g610) & (!g1163) & (g1593) & (!g1594)) + ((g545) & (!g602) & (!g610) & (g1163) & (g1593) & (!g1594)) + ((g545) & (!g602) & (!g610) & (g1163) & (g1593) & (g1594)) + ((g545) & (!g602) & (g610) & (!g1163) & (!g1593) & (g1594)) + ((g545) & (!g602) & (g610) & (!g1163) & (g1593) & (g1594)) + ((g545) & (!g602) & (g610) & (g1163) & (!g1593) & (!g1594)) + ((g545) & (!g602) & (g610) & (g1163) & (!g1593) & (g1594)) + ((g545) & (g602) & (!g610) & (!g1163) & (!g1593) & (g1594)) + ((g545) & (g602) & (!g610) & (!g1163) & (g1593) & (g1594)) + ((g545) & (g602) & (!g610) & (g1163) & (g1593) & (!g1594)) + ((g545) & (g602) & (!g610) & (g1163) & (g1593) & (g1594)) + ((g545) & (g602) & (g610) & (!g1163) & (!g1593) & (!g1594)) + ((g545) & (g602) & (g610) & (!g1163) & (g1593) & (!g1594)) + ((g545) & (g602) & (g610) & (g1163) & (!g1593) & (!g1594)) + ((g545) & (g602) & (g610) & (g1163) & (!g1593) & (g1594)));
	assign g2141 = (((!ld) & (!text_inx59x) & (sk[45]) & (g1596)) + ((!ld) & (text_inx59x) & (!sk[45]) & (!g1596)) + ((!ld) & (text_inx59x) & (!sk[45]) & (g1596)) + ((!ld) & (text_inx59x) & (sk[45]) & (g1596)) + ((ld) & (!text_inx59x) & (!sk[45]) & (g1596)) + ((ld) & (text_inx59x) & (!sk[45]) & (!g1596)) + ((ld) & (text_inx59x) & (!sk[45]) & (g1596)) + ((ld) & (text_inx59x) & (sk[45]) & (!g1596)) + ((ld) & (text_inx59x) & (sk[45]) & (g1596)));
	assign g2142 = (((!ld) & (!sk[46]) & (text_inx62x) & (!g1597)) + ((!ld) & (!sk[46]) & (text_inx62x) & (g1597)) + ((!ld) & (sk[46]) & (!text_inx62x) & (g1597)) + ((!ld) & (sk[46]) & (text_inx62x) & (g1597)) + ((ld) & (!sk[46]) & (!text_inx62x) & (g1597)) + ((ld) & (!sk[46]) & (text_inx62x) & (!g1597)) + ((ld) & (!sk[46]) & (text_inx62x) & (g1597)) + ((ld) & (sk[46]) & (text_inx62x) & (!g1597)) + ((ld) & (sk[46]) & (text_inx62x) & (g1597)));
	assign g1598 = (((!g445) & (!g509) & (sk[47]) & (g566)) + ((!g445) & (g509) & (!sk[47]) & (!g566)) + ((!g445) & (g509) & (!sk[47]) & (g566)) + ((!g445) & (g509) & (sk[47]) & (!g566)) + ((g445) & (!g509) & (!sk[47]) & (g566)) + ((g445) & (!g509) & (sk[47]) & (!g566)) + ((g445) & (g509) & (!sk[47]) & (!g566)) + ((g445) & (g509) & (!sk[47]) & (g566)) + ((g445) & (g509) & (sk[47]) & (g566)));
	assign g1599 = (((!g573) & (!g630) & (!g638) & (!g1163) & (!g1597) & (g1598)) + ((!g573) & (!g630) & (!g638) & (!g1163) & (g1597) & (g1598)) + ((!g573) & (!g630) & (!g638) & (g1163) & (g1597) & (!g1598)) + ((!g573) & (!g630) & (!g638) & (g1163) & (g1597) & (g1598)) + ((!g573) & (!g630) & (g638) & (!g1163) & (!g1597) & (!g1598)) + ((!g573) & (!g630) & (g638) & (!g1163) & (g1597) & (!g1598)) + ((!g573) & (!g630) & (g638) & (g1163) & (!g1597) & (!g1598)) + ((!g573) & (!g630) & (g638) & (g1163) & (!g1597) & (g1598)) + ((!g573) & (g630) & (!g638) & (!g1163) & (!g1597) & (!g1598)) + ((!g573) & (g630) & (!g638) & (!g1163) & (g1597) & (!g1598)) + ((!g573) & (g630) & (!g638) & (g1163) & (g1597) & (!g1598)) + ((!g573) & (g630) & (!g638) & (g1163) & (g1597) & (g1598)) + ((!g573) & (g630) & (g638) & (!g1163) & (!g1597) & (g1598)) + ((!g573) & (g630) & (g638) & (!g1163) & (g1597) & (g1598)) + ((!g573) & (g630) & (g638) & (g1163) & (!g1597) & (!g1598)) + ((!g573) & (g630) & (g638) & (g1163) & (!g1597) & (g1598)) + ((g573) & (!g630) & (!g638) & (!g1163) & (!g1597) & (!g1598)) + ((g573) & (!g630) & (!g638) & (!g1163) & (g1597) & (!g1598)) + ((g573) & (!g630) & (!g638) & (g1163) & (g1597) & (!g1598)) + ((g573) & (!g630) & (!g638) & (g1163) & (g1597) & (g1598)) + ((g573) & (!g630) & (g638) & (!g1163) & (!g1597) & (g1598)) + ((g573) & (!g630) & (g638) & (!g1163) & (g1597) & (g1598)) + ((g573) & (!g630) & (g638) & (g1163) & (!g1597) & (!g1598)) + ((g573) & (!g630) & (g638) & (g1163) & (!g1597) & (g1598)) + ((g573) & (g630) & (!g638) & (!g1163) & (!g1597) & (g1598)) + ((g573) & (g630) & (!g638) & (!g1163) & (g1597) & (g1598)) + ((g573) & (g630) & (!g638) & (g1163) & (g1597) & (!g1598)) + ((g573) & (g630) & (!g638) & (g1163) & (g1597) & (g1598)) + ((g573) & (g630) & (g638) & (!g1163) & (!g1597) & (!g1598)) + ((g573) & (g630) & (g638) & (!g1163) & (g1597) & (!g1598)) + ((g573) & (g630) & (g638) & (g1163) & (!g1597) & (!g1598)) + ((g573) & (g630) & (g638) & (g1163) & (!g1597) & (g1598)));
	assign g2143 = (((!ld) & (!sk[49]) & (text_inx61x) & (!g1600)) + ((!ld) & (!sk[49]) & (text_inx61x) & (g1600)) + ((!ld) & (sk[49]) & (!text_inx61x) & (g1600)) + ((!ld) & (sk[49]) & (text_inx61x) & (g1600)) + ((ld) & (!sk[49]) & (!text_inx61x) & (g1600)) + ((ld) & (!sk[49]) & (text_inx61x) & (!g1600)) + ((ld) & (!sk[49]) & (text_inx61x) & (g1600)) + ((ld) & (sk[49]) & (text_inx61x) & (!g1600)) + ((ld) & (sk[49]) & (text_inx61x) & (g1600)));
	assign g1601 = (((!sk[50]) & (!g438) & (g502) & (!g559)) + ((!sk[50]) & (!g438) & (g502) & (g559)) + ((!sk[50]) & (g438) & (!g502) & (g559)) + ((!sk[50]) & (g438) & (g502) & (!g559)) + ((!sk[50]) & (g438) & (g502) & (g559)) + ((sk[50]) & (!g438) & (!g502) & (g559)) + ((sk[50]) & (!g438) & (g502) & (!g559)) + ((sk[50]) & (g438) & (!g502) & (!g559)) + ((sk[50]) & (g438) & (g502) & (g559)));
	assign g1602 = (((!g566) & (!g623) & (!g631) & (!g1163) & (!g1600) & (g1601)) + ((!g566) & (!g623) & (!g631) & (!g1163) & (g1600) & (g1601)) + ((!g566) & (!g623) & (!g631) & (g1163) & (g1600) & (!g1601)) + ((!g566) & (!g623) & (!g631) & (g1163) & (g1600) & (g1601)) + ((!g566) & (!g623) & (g631) & (!g1163) & (!g1600) & (!g1601)) + ((!g566) & (!g623) & (g631) & (!g1163) & (g1600) & (!g1601)) + ((!g566) & (!g623) & (g631) & (g1163) & (!g1600) & (!g1601)) + ((!g566) & (!g623) & (g631) & (g1163) & (!g1600) & (g1601)) + ((!g566) & (g623) & (!g631) & (!g1163) & (!g1600) & (!g1601)) + ((!g566) & (g623) & (!g631) & (!g1163) & (g1600) & (!g1601)) + ((!g566) & (g623) & (!g631) & (g1163) & (g1600) & (!g1601)) + ((!g566) & (g623) & (!g631) & (g1163) & (g1600) & (g1601)) + ((!g566) & (g623) & (g631) & (!g1163) & (!g1600) & (g1601)) + ((!g566) & (g623) & (g631) & (!g1163) & (g1600) & (g1601)) + ((!g566) & (g623) & (g631) & (g1163) & (!g1600) & (!g1601)) + ((!g566) & (g623) & (g631) & (g1163) & (!g1600) & (g1601)) + ((g566) & (!g623) & (!g631) & (!g1163) & (!g1600) & (!g1601)) + ((g566) & (!g623) & (!g631) & (!g1163) & (g1600) & (!g1601)) + ((g566) & (!g623) & (!g631) & (g1163) & (g1600) & (!g1601)) + ((g566) & (!g623) & (!g631) & (g1163) & (g1600) & (g1601)) + ((g566) & (!g623) & (g631) & (!g1163) & (!g1600) & (g1601)) + ((g566) & (!g623) & (g631) & (!g1163) & (g1600) & (g1601)) + ((g566) & (!g623) & (g631) & (g1163) & (!g1600) & (!g1601)) + ((g566) & (!g623) & (g631) & (g1163) & (!g1600) & (g1601)) + ((g566) & (g623) & (!g631) & (!g1163) & (!g1600) & (g1601)) + ((g566) & (g623) & (!g631) & (!g1163) & (g1600) & (g1601)) + ((g566) & (g623) & (!g631) & (g1163) & (g1600) & (!g1601)) + ((g566) & (g623) & (!g631) & (g1163) & (g1600) & (g1601)) + ((g566) & (g623) & (g631) & (!g1163) & (!g1600) & (!g1601)) + ((g566) & (g623) & (g631) & (!g1163) & (g1600) & (!g1601)) + ((g566) & (g623) & (g631) & (g1163) & (!g1600) & (!g1601)) + ((g566) & (g623) & (g631) & (g1163) & (!g1600) & (g1601)));
	assign g2144 = (((!ld) & (!sk[52]) & (text_inx60x) & (!g1603)) + ((!ld) & (!sk[52]) & (text_inx60x) & (g1603)) + ((!ld) & (sk[52]) & (!text_inx60x) & (g1603)) + ((!ld) & (sk[52]) & (text_inx60x) & (g1603)) + ((ld) & (!sk[52]) & (!text_inx60x) & (g1603)) + ((ld) & (!sk[52]) & (text_inx60x) & (!g1603)) + ((ld) & (!sk[52]) & (text_inx60x) & (g1603)) + ((ld) & (sk[52]) & (text_inx60x) & (!g1603)) + ((ld) & (sk[52]) & (text_inx60x) & (g1603)));
	assign g1604 = (((!g431) & (!g495) & (sk[53]) & (g552)) + ((!g431) & (g495) & (!sk[53]) & (!g552)) + ((!g431) & (g495) & (!sk[53]) & (g552)) + ((!g431) & (g495) & (sk[53]) & (!g552)) + ((g431) & (!g495) & (!sk[53]) & (g552)) + ((g431) & (!g495) & (sk[53]) & (!g552)) + ((g431) & (g495) & (!sk[53]) & (!g552)) + ((g431) & (g495) & (!sk[53]) & (g552)) + ((g431) & (g495) & (sk[53]) & (g552)));
	assign g1605 = (((!sk[54]) & (!g559) & (g580) & (!g616) & (!g624) & (!g644)) + ((!sk[54]) & (!g559) & (g580) & (!g616) & (!g624) & (g644)) + ((!sk[54]) & (!g559) & (g580) & (!g616) & (g624) & (!g644)) + ((!sk[54]) & (!g559) & (g580) & (!g616) & (g624) & (g644)) + ((!sk[54]) & (!g559) & (g580) & (g616) & (!g624) & (!g644)) + ((!sk[54]) & (!g559) & (g580) & (g616) & (!g624) & (g644)) + ((!sk[54]) & (!g559) & (g580) & (g616) & (g624) & (!g644)) + ((!sk[54]) & (!g559) & (g580) & (g616) & (g624) & (g644)) + ((!sk[54]) & (g559) & (!g580) & (!g616) & (!g624) & (!g644)) + ((!sk[54]) & (g559) & (!g580) & (!g616) & (!g624) & (g644)) + ((!sk[54]) & (g559) & (!g580) & (!g616) & (g624) & (!g644)) + ((!sk[54]) & (g559) & (!g580) & (!g616) & (g624) & (g644)) + ((!sk[54]) & (g559) & (!g580) & (g616) & (!g624) & (!g644)) + ((!sk[54]) & (g559) & (!g580) & (g616) & (!g624) & (g644)) + ((!sk[54]) & (g559) & (!g580) & (g616) & (g624) & (!g644)) + ((!sk[54]) & (g559) & (!g580) & (g616) & (g624) & (g644)) + ((!sk[54]) & (g559) & (g580) & (!g616) & (!g624) & (!g644)) + ((!sk[54]) & (g559) & (g580) & (!g616) & (!g624) & (g644)) + ((!sk[54]) & (g559) & (g580) & (!g616) & (g624) & (!g644)) + ((!sk[54]) & (g559) & (g580) & (!g616) & (g624) & (g644)) + ((!sk[54]) & (g559) & (g580) & (g616) & (!g624) & (!g644)) + ((!sk[54]) & (g559) & (g580) & (g616) & (!g624) & (g644)) + ((!sk[54]) & (g559) & (g580) & (g616) & (g624) & (!g644)) + ((!sk[54]) & (g559) & (g580) & (g616) & (g624) & (g644)) + ((sk[54]) & (!g559) & (!g580) & (!g616) & (!g624) & (g644)) + ((sk[54]) & (!g559) & (!g580) & (!g616) & (g624) & (!g644)) + ((sk[54]) & (!g559) & (!g580) & (g616) & (!g624) & (!g644)) + ((sk[54]) & (!g559) & (!g580) & (g616) & (g624) & (g644)) + ((sk[54]) & (!g559) & (g580) & (!g616) & (!g624) & (!g644)) + ((sk[54]) & (!g559) & (g580) & (!g616) & (g624) & (g644)) + ((sk[54]) & (!g559) & (g580) & (g616) & (!g624) & (g644)) + ((sk[54]) & (!g559) & (g580) & (g616) & (g624) & (!g644)) + ((sk[54]) & (g559) & (!g580) & (!g616) & (!g624) & (!g644)) + ((sk[54]) & (g559) & (!g580) & (!g616) & (g624) & (g644)) + ((sk[54]) & (g559) & (!g580) & (g616) & (!g624) & (g644)) + ((sk[54]) & (g559) & (!g580) & (g616) & (g624) & (!g644)) + ((sk[54]) & (g559) & (g580) & (!g616) & (!g624) & (g644)) + ((sk[54]) & (g559) & (g580) & (!g616) & (g624) & (!g644)) + ((sk[54]) & (g559) & (g580) & (g616) & (!g624) & (!g644)) + ((sk[54]) & (g559) & (g580) & (g616) & (g624) & (g644)));
	assign g1606 = (((!g624) & (!g1163) & (!g1603) & (!g1604) & (sk[55]) & (g1605)) + ((!g624) & (!g1163) & (!g1603) & (g1604) & (sk[55]) & (!g1605)) + ((!g624) & (!g1163) & (g1603) & (!g1604) & (sk[55]) & (g1605)) + ((!g624) & (!g1163) & (g1603) & (g1604) & (sk[55]) & (!g1605)) + ((!g624) & (g1163) & (!g1603) & (!g1604) & (!sk[55]) & (!g1605)) + ((!g624) & (g1163) & (!g1603) & (!g1604) & (!sk[55]) & (g1605)) + ((!g624) & (g1163) & (!g1603) & (g1604) & (!sk[55]) & (!g1605)) + ((!g624) & (g1163) & (!g1603) & (g1604) & (!sk[55]) & (g1605)) + ((!g624) & (g1163) & (g1603) & (!g1604) & (!sk[55]) & (!g1605)) + ((!g624) & (g1163) & (g1603) & (!g1604) & (!sk[55]) & (g1605)) + ((!g624) & (g1163) & (g1603) & (!g1604) & (sk[55]) & (!g1605)) + ((!g624) & (g1163) & (g1603) & (!g1604) & (sk[55]) & (g1605)) + ((!g624) & (g1163) & (g1603) & (g1604) & (!sk[55]) & (!g1605)) + ((!g624) & (g1163) & (g1603) & (g1604) & (!sk[55]) & (g1605)) + ((!g624) & (g1163) & (g1603) & (g1604) & (sk[55]) & (!g1605)) + ((!g624) & (g1163) & (g1603) & (g1604) & (sk[55]) & (g1605)) + ((g624) & (!g1163) & (!g1603) & (!g1604) & (!sk[55]) & (!g1605)) + ((g624) & (!g1163) & (!g1603) & (!g1604) & (!sk[55]) & (g1605)) + ((g624) & (!g1163) & (!g1603) & (!g1604) & (sk[55]) & (g1605)) + ((g624) & (!g1163) & (!g1603) & (g1604) & (!sk[55]) & (!g1605)) + ((g624) & (!g1163) & (!g1603) & (g1604) & (!sk[55]) & (g1605)) + ((g624) & (!g1163) & (!g1603) & (g1604) & (sk[55]) & (!g1605)) + ((g624) & (!g1163) & (g1603) & (!g1604) & (!sk[55]) & (!g1605)) + ((g624) & (!g1163) & (g1603) & (!g1604) & (!sk[55]) & (g1605)) + ((g624) & (!g1163) & (g1603) & (!g1604) & (sk[55]) & (g1605)) + ((g624) & (!g1163) & (g1603) & (g1604) & (!sk[55]) & (!g1605)) + ((g624) & (!g1163) & (g1603) & (g1604) & (!sk[55]) & (g1605)) + ((g624) & (!g1163) & (g1603) & (g1604) & (sk[55]) & (!g1605)) + ((g624) & (g1163) & (!g1603) & (!g1604) & (!sk[55]) & (!g1605)) + ((g624) & (g1163) & (!g1603) & (!g1604) & (!sk[55]) & (g1605)) + ((g624) & (g1163) & (!g1603) & (!g1604) & (sk[55]) & (!g1605)) + ((g624) & (g1163) & (!g1603) & (!g1604) & (sk[55]) & (g1605)) + ((g624) & (g1163) & (!g1603) & (g1604) & (!sk[55]) & (!g1605)) + ((g624) & (g1163) & (!g1603) & (g1604) & (!sk[55]) & (g1605)) + ((g624) & (g1163) & (!g1603) & (g1604) & (sk[55]) & (!g1605)) + ((g624) & (g1163) & (!g1603) & (g1604) & (sk[55]) & (g1605)) + ((g624) & (g1163) & (g1603) & (!g1604) & (!sk[55]) & (!g1605)) + ((g624) & (g1163) & (g1603) & (!g1604) & (!sk[55]) & (g1605)) + ((g624) & (g1163) & (g1603) & (g1604) & (!sk[55]) & (!g1605)) + ((g624) & (g1163) & (g1603) & (g1604) & (!sk[55]) & (g1605)));
	assign g2145 = (((!ld) & (!sk[56]) & (text_inx63x) & (!g1607)) + ((!ld) & (!sk[56]) & (text_inx63x) & (g1607)) + ((!ld) & (sk[56]) & (!text_inx63x) & (g1607)) + ((!ld) & (sk[56]) & (text_inx63x) & (g1607)) + ((ld) & (!sk[56]) & (!text_inx63x) & (g1607)) + ((ld) & (!sk[56]) & (text_inx63x) & (!g1607)) + ((ld) & (!sk[56]) & (text_inx63x) & (g1607)) + ((ld) & (sk[56]) & (text_inx63x) & (!g1607)) + ((ld) & (sk[56]) & (text_inx63x) & (g1607)));
	assign g1608 = (((!g452) & (!g516) & (sk[57]) & (g573)) + ((!g452) & (g516) & (!sk[57]) & (!g573)) + ((!g452) & (g516) & (!sk[57]) & (g573)) + ((!g452) & (g516) & (sk[57]) & (!g573)) + ((g452) & (!g516) & (!sk[57]) & (g573)) + ((g452) & (!g516) & (sk[57]) & (!g573)) + ((g452) & (g516) & (!sk[57]) & (!g573)) + ((g452) & (g516) & (!sk[57]) & (g573)) + ((g452) & (g516) & (sk[57]) & (g573)));
	assign g1609 = (((!g580) & (!g637) & (!g645) & (!g1163) & (!g1607) & (g1608)) + ((!g580) & (!g637) & (!g645) & (!g1163) & (g1607) & (g1608)) + ((!g580) & (!g637) & (!g645) & (g1163) & (g1607) & (!g1608)) + ((!g580) & (!g637) & (!g645) & (g1163) & (g1607) & (g1608)) + ((!g580) & (!g637) & (g645) & (!g1163) & (!g1607) & (!g1608)) + ((!g580) & (!g637) & (g645) & (!g1163) & (g1607) & (!g1608)) + ((!g580) & (!g637) & (g645) & (g1163) & (!g1607) & (!g1608)) + ((!g580) & (!g637) & (g645) & (g1163) & (!g1607) & (g1608)) + ((!g580) & (g637) & (!g645) & (!g1163) & (!g1607) & (!g1608)) + ((!g580) & (g637) & (!g645) & (!g1163) & (g1607) & (!g1608)) + ((!g580) & (g637) & (!g645) & (g1163) & (g1607) & (!g1608)) + ((!g580) & (g637) & (!g645) & (g1163) & (g1607) & (g1608)) + ((!g580) & (g637) & (g645) & (!g1163) & (!g1607) & (g1608)) + ((!g580) & (g637) & (g645) & (!g1163) & (g1607) & (g1608)) + ((!g580) & (g637) & (g645) & (g1163) & (!g1607) & (!g1608)) + ((!g580) & (g637) & (g645) & (g1163) & (!g1607) & (g1608)) + ((g580) & (!g637) & (!g645) & (!g1163) & (!g1607) & (!g1608)) + ((g580) & (!g637) & (!g645) & (!g1163) & (g1607) & (!g1608)) + ((g580) & (!g637) & (!g645) & (g1163) & (g1607) & (!g1608)) + ((g580) & (!g637) & (!g645) & (g1163) & (g1607) & (g1608)) + ((g580) & (!g637) & (g645) & (!g1163) & (!g1607) & (g1608)) + ((g580) & (!g637) & (g645) & (!g1163) & (g1607) & (g1608)) + ((g580) & (!g637) & (g645) & (g1163) & (!g1607) & (!g1608)) + ((g580) & (!g637) & (g645) & (g1163) & (!g1607) & (g1608)) + ((g580) & (g637) & (!g645) & (!g1163) & (!g1607) & (g1608)) + ((g580) & (g637) & (!g645) & (!g1163) & (g1607) & (g1608)) + ((g580) & (g637) & (!g645) & (g1163) & (g1607) & (!g1608)) + ((g580) & (g637) & (!g645) & (g1163) & (g1607) & (g1608)) + ((g580) & (g637) & (g645) & (!g1163) & (!g1607) & (!g1608)) + ((g580) & (g637) & (g645) & (!g1163) & (g1607) & (!g1608)) + ((g580) & (g637) & (g645) & (g1163) & (!g1607) & (!g1608)) + ((g580) & (g637) & (g645) & (g1163) & (!g1607) & (g1608)));
	assign g1610 = (((!ld) & (!g596) & (!g852) & (!g1438) & (g1440) & (!keyx56x)) + ((!ld) & (!g596) & (!g852) & (!g1438) & (g1440) & (keyx56x)) + ((!ld) & (!g596) & (!g852) & (g1438) & (!g1440) & (!keyx56x)) + ((!ld) & (!g596) & (!g852) & (g1438) & (!g1440) & (keyx56x)) + ((!ld) & (!g596) & (g852) & (!g1438) & (!g1440) & (!keyx56x)) + ((!ld) & (!g596) & (g852) & (!g1438) & (!g1440) & (keyx56x)) + ((!ld) & (!g596) & (g852) & (g1438) & (g1440) & (!keyx56x)) + ((!ld) & (!g596) & (g852) & (g1438) & (g1440) & (keyx56x)) + ((!ld) & (g596) & (!g852) & (!g1438) & (!g1440) & (!keyx56x)) + ((!ld) & (g596) & (!g852) & (!g1438) & (!g1440) & (keyx56x)) + ((!ld) & (g596) & (!g852) & (g1438) & (g1440) & (!keyx56x)) + ((!ld) & (g596) & (!g852) & (g1438) & (g1440) & (keyx56x)) + ((!ld) & (g596) & (g852) & (!g1438) & (g1440) & (!keyx56x)) + ((!ld) & (g596) & (g852) & (!g1438) & (g1440) & (keyx56x)) + ((!ld) & (g596) & (g852) & (g1438) & (!g1440) & (!keyx56x)) + ((!ld) & (g596) & (g852) & (g1438) & (!g1440) & (keyx56x)) + ((ld) & (!g596) & (!g852) & (!g1438) & (!g1440) & (keyx56x)) + ((ld) & (!g596) & (!g852) & (!g1438) & (g1440) & (keyx56x)) + ((ld) & (!g596) & (!g852) & (g1438) & (!g1440) & (keyx56x)) + ((ld) & (!g596) & (!g852) & (g1438) & (g1440) & (keyx56x)) + ((ld) & (!g596) & (g852) & (!g1438) & (!g1440) & (keyx56x)) + ((ld) & (!g596) & (g852) & (!g1438) & (g1440) & (keyx56x)) + ((ld) & (!g596) & (g852) & (g1438) & (!g1440) & (keyx56x)) + ((ld) & (!g596) & (g852) & (g1438) & (g1440) & (keyx56x)) + ((ld) & (g596) & (!g852) & (!g1438) & (!g1440) & (keyx56x)) + ((ld) & (g596) & (!g852) & (!g1438) & (g1440) & (keyx56x)) + ((ld) & (g596) & (!g852) & (g1438) & (!g1440) & (keyx56x)) + ((ld) & (g596) & (!g852) & (g1438) & (g1440) & (keyx56x)) + ((ld) & (g596) & (g852) & (!g1438) & (!g1440) & (keyx56x)) + ((ld) & (g596) & (g852) & (!g1438) & (g1440) & (keyx56x)) + ((ld) & (g596) & (g852) & (g1438) & (!g1440) & (keyx56x)) + ((ld) & (g596) & (g852) & (g1438) & (g1440) & (keyx56x)));
	assign g1611 = (((!ld) & (!g603) & (!g859) & (!g1447) & (g1449) & (!keyx57x)) + ((!ld) & (!g603) & (!g859) & (!g1447) & (g1449) & (keyx57x)) + ((!ld) & (!g603) & (!g859) & (g1447) & (!g1449) & (!keyx57x)) + ((!ld) & (!g603) & (!g859) & (g1447) & (!g1449) & (keyx57x)) + ((!ld) & (!g603) & (g859) & (!g1447) & (!g1449) & (!keyx57x)) + ((!ld) & (!g603) & (g859) & (!g1447) & (!g1449) & (keyx57x)) + ((!ld) & (!g603) & (g859) & (g1447) & (g1449) & (!keyx57x)) + ((!ld) & (!g603) & (g859) & (g1447) & (g1449) & (keyx57x)) + ((!ld) & (g603) & (!g859) & (!g1447) & (!g1449) & (!keyx57x)) + ((!ld) & (g603) & (!g859) & (!g1447) & (!g1449) & (keyx57x)) + ((!ld) & (g603) & (!g859) & (g1447) & (g1449) & (!keyx57x)) + ((!ld) & (g603) & (!g859) & (g1447) & (g1449) & (keyx57x)) + ((!ld) & (g603) & (g859) & (!g1447) & (g1449) & (!keyx57x)) + ((!ld) & (g603) & (g859) & (!g1447) & (g1449) & (keyx57x)) + ((!ld) & (g603) & (g859) & (g1447) & (!g1449) & (!keyx57x)) + ((!ld) & (g603) & (g859) & (g1447) & (!g1449) & (keyx57x)) + ((ld) & (!g603) & (!g859) & (!g1447) & (!g1449) & (keyx57x)) + ((ld) & (!g603) & (!g859) & (!g1447) & (g1449) & (keyx57x)) + ((ld) & (!g603) & (!g859) & (g1447) & (!g1449) & (keyx57x)) + ((ld) & (!g603) & (!g859) & (g1447) & (g1449) & (keyx57x)) + ((ld) & (!g603) & (g859) & (!g1447) & (!g1449) & (keyx57x)) + ((ld) & (!g603) & (g859) & (!g1447) & (g1449) & (keyx57x)) + ((ld) & (!g603) & (g859) & (g1447) & (!g1449) & (keyx57x)) + ((ld) & (!g603) & (g859) & (g1447) & (g1449) & (keyx57x)) + ((ld) & (g603) & (!g859) & (!g1447) & (!g1449) & (keyx57x)) + ((ld) & (g603) & (!g859) & (!g1447) & (g1449) & (keyx57x)) + ((ld) & (g603) & (!g859) & (g1447) & (!g1449) & (keyx57x)) + ((ld) & (g603) & (!g859) & (g1447) & (g1449) & (keyx57x)) + ((ld) & (g603) & (g859) & (!g1447) & (!g1449) & (keyx57x)) + ((ld) & (g603) & (g859) & (!g1447) & (g1449) & (keyx57x)) + ((ld) & (g603) & (g859) & (g1447) & (!g1449) & (keyx57x)) + ((ld) & (g603) & (g859) & (g1447) & (g1449) & (keyx57x)));
	assign g1612 = (((!ld) & (!g610) & (!g866) & (!g1456) & (g1458) & (!keyx58x)) + ((!ld) & (!g610) & (!g866) & (!g1456) & (g1458) & (keyx58x)) + ((!ld) & (!g610) & (!g866) & (g1456) & (!g1458) & (!keyx58x)) + ((!ld) & (!g610) & (!g866) & (g1456) & (!g1458) & (keyx58x)) + ((!ld) & (!g610) & (g866) & (!g1456) & (!g1458) & (!keyx58x)) + ((!ld) & (!g610) & (g866) & (!g1456) & (!g1458) & (keyx58x)) + ((!ld) & (!g610) & (g866) & (g1456) & (g1458) & (!keyx58x)) + ((!ld) & (!g610) & (g866) & (g1456) & (g1458) & (keyx58x)) + ((!ld) & (g610) & (!g866) & (!g1456) & (!g1458) & (!keyx58x)) + ((!ld) & (g610) & (!g866) & (!g1456) & (!g1458) & (keyx58x)) + ((!ld) & (g610) & (!g866) & (g1456) & (g1458) & (!keyx58x)) + ((!ld) & (g610) & (!g866) & (g1456) & (g1458) & (keyx58x)) + ((!ld) & (g610) & (g866) & (!g1456) & (g1458) & (!keyx58x)) + ((!ld) & (g610) & (g866) & (!g1456) & (g1458) & (keyx58x)) + ((!ld) & (g610) & (g866) & (g1456) & (!g1458) & (!keyx58x)) + ((!ld) & (g610) & (g866) & (g1456) & (!g1458) & (keyx58x)) + ((ld) & (!g610) & (!g866) & (!g1456) & (!g1458) & (keyx58x)) + ((ld) & (!g610) & (!g866) & (!g1456) & (g1458) & (keyx58x)) + ((ld) & (!g610) & (!g866) & (g1456) & (!g1458) & (keyx58x)) + ((ld) & (!g610) & (!g866) & (g1456) & (g1458) & (keyx58x)) + ((ld) & (!g610) & (g866) & (!g1456) & (!g1458) & (keyx58x)) + ((ld) & (!g610) & (g866) & (!g1456) & (g1458) & (keyx58x)) + ((ld) & (!g610) & (g866) & (g1456) & (!g1458) & (keyx58x)) + ((ld) & (!g610) & (g866) & (g1456) & (g1458) & (keyx58x)) + ((ld) & (g610) & (!g866) & (!g1456) & (!g1458) & (keyx58x)) + ((ld) & (g610) & (!g866) & (!g1456) & (g1458) & (keyx58x)) + ((ld) & (g610) & (!g866) & (g1456) & (!g1458) & (keyx58x)) + ((ld) & (g610) & (!g866) & (g1456) & (g1458) & (keyx58x)) + ((ld) & (g610) & (g866) & (!g1456) & (!g1458) & (keyx58x)) + ((ld) & (g610) & (g866) & (!g1456) & (g1458) & (keyx58x)) + ((ld) & (g610) & (g866) & (g1456) & (!g1458) & (keyx58x)) + ((ld) & (g610) & (g866) & (g1456) & (g1458) & (keyx58x)));
	assign g1613 = (((!ld) & (!g617) & (!g873) & (!g1465) & (g1467) & (!keyx59x)) + ((!ld) & (!g617) & (!g873) & (!g1465) & (g1467) & (keyx59x)) + ((!ld) & (!g617) & (!g873) & (g1465) & (!g1467) & (!keyx59x)) + ((!ld) & (!g617) & (!g873) & (g1465) & (!g1467) & (keyx59x)) + ((!ld) & (!g617) & (g873) & (!g1465) & (!g1467) & (!keyx59x)) + ((!ld) & (!g617) & (g873) & (!g1465) & (!g1467) & (keyx59x)) + ((!ld) & (!g617) & (g873) & (g1465) & (g1467) & (!keyx59x)) + ((!ld) & (!g617) & (g873) & (g1465) & (g1467) & (keyx59x)) + ((!ld) & (g617) & (!g873) & (!g1465) & (!g1467) & (!keyx59x)) + ((!ld) & (g617) & (!g873) & (!g1465) & (!g1467) & (keyx59x)) + ((!ld) & (g617) & (!g873) & (g1465) & (g1467) & (!keyx59x)) + ((!ld) & (g617) & (!g873) & (g1465) & (g1467) & (keyx59x)) + ((!ld) & (g617) & (g873) & (!g1465) & (g1467) & (!keyx59x)) + ((!ld) & (g617) & (g873) & (!g1465) & (g1467) & (keyx59x)) + ((!ld) & (g617) & (g873) & (g1465) & (!g1467) & (!keyx59x)) + ((!ld) & (g617) & (g873) & (g1465) & (!g1467) & (keyx59x)) + ((ld) & (!g617) & (!g873) & (!g1465) & (!g1467) & (keyx59x)) + ((ld) & (!g617) & (!g873) & (!g1465) & (g1467) & (keyx59x)) + ((ld) & (!g617) & (!g873) & (g1465) & (!g1467) & (keyx59x)) + ((ld) & (!g617) & (!g873) & (g1465) & (g1467) & (keyx59x)) + ((ld) & (!g617) & (g873) & (!g1465) & (!g1467) & (keyx59x)) + ((ld) & (!g617) & (g873) & (!g1465) & (g1467) & (keyx59x)) + ((ld) & (!g617) & (g873) & (g1465) & (!g1467) & (keyx59x)) + ((ld) & (!g617) & (g873) & (g1465) & (g1467) & (keyx59x)) + ((ld) & (g617) & (!g873) & (!g1465) & (!g1467) & (keyx59x)) + ((ld) & (g617) & (!g873) & (!g1465) & (g1467) & (keyx59x)) + ((ld) & (g617) & (!g873) & (g1465) & (!g1467) & (keyx59x)) + ((ld) & (g617) & (!g873) & (g1465) & (g1467) & (keyx59x)) + ((ld) & (g617) & (g873) & (!g1465) & (!g1467) & (keyx59x)) + ((ld) & (g617) & (g873) & (!g1465) & (g1467) & (keyx59x)) + ((ld) & (g617) & (g873) & (g1465) & (!g1467) & (keyx59x)) + ((ld) & (g617) & (g873) & (g1465) & (g1467) & (keyx59x)));
	assign g1614 = (((!ld) & (!g624) & (!g880) & (!g1474) & (g1476) & (!keyx60x)) + ((!ld) & (!g624) & (!g880) & (!g1474) & (g1476) & (keyx60x)) + ((!ld) & (!g624) & (!g880) & (g1474) & (!g1476) & (!keyx60x)) + ((!ld) & (!g624) & (!g880) & (g1474) & (!g1476) & (keyx60x)) + ((!ld) & (!g624) & (g880) & (!g1474) & (!g1476) & (!keyx60x)) + ((!ld) & (!g624) & (g880) & (!g1474) & (!g1476) & (keyx60x)) + ((!ld) & (!g624) & (g880) & (g1474) & (g1476) & (!keyx60x)) + ((!ld) & (!g624) & (g880) & (g1474) & (g1476) & (keyx60x)) + ((!ld) & (g624) & (!g880) & (!g1474) & (!g1476) & (!keyx60x)) + ((!ld) & (g624) & (!g880) & (!g1474) & (!g1476) & (keyx60x)) + ((!ld) & (g624) & (!g880) & (g1474) & (g1476) & (!keyx60x)) + ((!ld) & (g624) & (!g880) & (g1474) & (g1476) & (keyx60x)) + ((!ld) & (g624) & (g880) & (!g1474) & (g1476) & (!keyx60x)) + ((!ld) & (g624) & (g880) & (!g1474) & (g1476) & (keyx60x)) + ((!ld) & (g624) & (g880) & (g1474) & (!g1476) & (!keyx60x)) + ((!ld) & (g624) & (g880) & (g1474) & (!g1476) & (keyx60x)) + ((ld) & (!g624) & (!g880) & (!g1474) & (!g1476) & (keyx60x)) + ((ld) & (!g624) & (!g880) & (!g1474) & (g1476) & (keyx60x)) + ((ld) & (!g624) & (!g880) & (g1474) & (!g1476) & (keyx60x)) + ((ld) & (!g624) & (!g880) & (g1474) & (g1476) & (keyx60x)) + ((ld) & (!g624) & (g880) & (!g1474) & (!g1476) & (keyx60x)) + ((ld) & (!g624) & (g880) & (!g1474) & (g1476) & (keyx60x)) + ((ld) & (!g624) & (g880) & (g1474) & (!g1476) & (keyx60x)) + ((ld) & (!g624) & (g880) & (g1474) & (g1476) & (keyx60x)) + ((ld) & (g624) & (!g880) & (!g1474) & (!g1476) & (keyx60x)) + ((ld) & (g624) & (!g880) & (!g1474) & (g1476) & (keyx60x)) + ((ld) & (g624) & (!g880) & (g1474) & (!g1476) & (keyx60x)) + ((ld) & (g624) & (!g880) & (g1474) & (g1476) & (keyx60x)) + ((ld) & (g624) & (g880) & (!g1474) & (!g1476) & (keyx60x)) + ((ld) & (g624) & (g880) & (!g1474) & (g1476) & (keyx60x)) + ((ld) & (g624) & (g880) & (g1474) & (!g1476) & (keyx60x)) + ((ld) & (g624) & (g880) & (g1474) & (g1476) & (keyx60x)));
	assign g1615 = (((!ld) & (!g631) & (!g887) & (!g1483) & (g1485) & (!keyx61x)) + ((!ld) & (!g631) & (!g887) & (!g1483) & (g1485) & (keyx61x)) + ((!ld) & (!g631) & (!g887) & (g1483) & (!g1485) & (!keyx61x)) + ((!ld) & (!g631) & (!g887) & (g1483) & (!g1485) & (keyx61x)) + ((!ld) & (!g631) & (g887) & (!g1483) & (!g1485) & (!keyx61x)) + ((!ld) & (!g631) & (g887) & (!g1483) & (!g1485) & (keyx61x)) + ((!ld) & (!g631) & (g887) & (g1483) & (g1485) & (!keyx61x)) + ((!ld) & (!g631) & (g887) & (g1483) & (g1485) & (keyx61x)) + ((!ld) & (g631) & (!g887) & (!g1483) & (!g1485) & (!keyx61x)) + ((!ld) & (g631) & (!g887) & (!g1483) & (!g1485) & (keyx61x)) + ((!ld) & (g631) & (!g887) & (g1483) & (g1485) & (!keyx61x)) + ((!ld) & (g631) & (!g887) & (g1483) & (g1485) & (keyx61x)) + ((!ld) & (g631) & (g887) & (!g1483) & (g1485) & (!keyx61x)) + ((!ld) & (g631) & (g887) & (!g1483) & (g1485) & (keyx61x)) + ((!ld) & (g631) & (g887) & (g1483) & (!g1485) & (!keyx61x)) + ((!ld) & (g631) & (g887) & (g1483) & (!g1485) & (keyx61x)) + ((ld) & (!g631) & (!g887) & (!g1483) & (!g1485) & (keyx61x)) + ((ld) & (!g631) & (!g887) & (!g1483) & (g1485) & (keyx61x)) + ((ld) & (!g631) & (!g887) & (g1483) & (!g1485) & (keyx61x)) + ((ld) & (!g631) & (!g887) & (g1483) & (g1485) & (keyx61x)) + ((ld) & (!g631) & (g887) & (!g1483) & (!g1485) & (keyx61x)) + ((ld) & (!g631) & (g887) & (!g1483) & (g1485) & (keyx61x)) + ((ld) & (!g631) & (g887) & (g1483) & (!g1485) & (keyx61x)) + ((ld) & (!g631) & (g887) & (g1483) & (g1485) & (keyx61x)) + ((ld) & (g631) & (!g887) & (!g1483) & (!g1485) & (keyx61x)) + ((ld) & (g631) & (!g887) & (!g1483) & (g1485) & (keyx61x)) + ((ld) & (g631) & (!g887) & (g1483) & (!g1485) & (keyx61x)) + ((ld) & (g631) & (!g887) & (g1483) & (g1485) & (keyx61x)) + ((ld) & (g631) & (g887) & (!g1483) & (!g1485) & (keyx61x)) + ((ld) & (g631) & (g887) & (!g1483) & (g1485) & (keyx61x)) + ((ld) & (g631) & (g887) & (g1483) & (!g1485) & (keyx61x)) + ((ld) & (g631) & (g887) & (g1483) & (g1485) & (keyx61x)));
	assign g1616 = (((!ld) & (!g638) & (!g894) & (!g1492) & (g1494) & (!keyx62x)) + ((!ld) & (!g638) & (!g894) & (!g1492) & (g1494) & (keyx62x)) + ((!ld) & (!g638) & (!g894) & (g1492) & (!g1494) & (!keyx62x)) + ((!ld) & (!g638) & (!g894) & (g1492) & (!g1494) & (keyx62x)) + ((!ld) & (!g638) & (g894) & (!g1492) & (!g1494) & (!keyx62x)) + ((!ld) & (!g638) & (g894) & (!g1492) & (!g1494) & (keyx62x)) + ((!ld) & (!g638) & (g894) & (g1492) & (g1494) & (!keyx62x)) + ((!ld) & (!g638) & (g894) & (g1492) & (g1494) & (keyx62x)) + ((!ld) & (g638) & (!g894) & (!g1492) & (!g1494) & (!keyx62x)) + ((!ld) & (g638) & (!g894) & (!g1492) & (!g1494) & (keyx62x)) + ((!ld) & (g638) & (!g894) & (g1492) & (g1494) & (!keyx62x)) + ((!ld) & (g638) & (!g894) & (g1492) & (g1494) & (keyx62x)) + ((!ld) & (g638) & (g894) & (!g1492) & (g1494) & (!keyx62x)) + ((!ld) & (g638) & (g894) & (!g1492) & (g1494) & (keyx62x)) + ((!ld) & (g638) & (g894) & (g1492) & (!g1494) & (!keyx62x)) + ((!ld) & (g638) & (g894) & (g1492) & (!g1494) & (keyx62x)) + ((ld) & (!g638) & (!g894) & (!g1492) & (!g1494) & (keyx62x)) + ((ld) & (!g638) & (!g894) & (!g1492) & (g1494) & (keyx62x)) + ((ld) & (!g638) & (!g894) & (g1492) & (!g1494) & (keyx62x)) + ((ld) & (!g638) & (!g894) & (g1492) & (g1494) & (keyx62x)) + ((ld) & (!g638) & (g894) & (!g1492) & (!g1494) & (keyx62x)) + ((ld) & (!g638) & (g894) & (!g1492) & (g1494) & (keyx62x)) + ((ld) & (!g638) & (g894) & (g1492) & (!g1494) & (keyx62x)) + ((ld) & (!g638) & (g894) & (g1492) & (g1494) & (keyx62x)) + ((ld) & (g638) & (!g894) & (!g1492) & (!g1494) & (keyx62x)) + ((ld) & (g638) & (!g894) & (!g1492) & (g1494) & (keyx62x)) + ((ld) & (g638) & (!g894) & (g1492) & (!g1494) & (keyx62x)) + ((ld) & (g638) & (!g894) & (g1492) & (g1494) & (keyx62x)) + ((ld) & (g638) & (g894) & (!g1492) & (!g1494) & (keyx62x)) + ((ld) & (g638) & (g894) & (!g1492) & (g1494) & (keyx62x)) + ((ld) & (g638) & (g894) & (g1492) & (!g1494) & (keyx62x)) + ((ld) & (g638) & (g894) & (g1492) & (g1494) & (keyx62x)));
	assign g1617 = (((!ld) & (!g645) & (!g901) & (!g1501) & (g1503) & (!keyx63x)) + ((!ld) & (!g645) & (!g901) & (!g1501) & (g1503) & (keyx63x)) + ((!ld) & (!g645) & (!g901) & (g1501) & (!g1503) & (!keyx63x)) + ((!ld) & (!g645) & (!g901) & (g1501) & (!g1503) & (keyx63x)) + ((!ld) & (!g645) & (g901) & (!g1501) & (!g1503) & (!keyx63x)) + ((!ld) & (!g645) & (g901) & (!g1501) & (!g1503) & (keyx63x)) + ((!ld) & (!g645) & (g901) & (g1501) & (g1503) & (!keyx63x)) + ((!ld) & (!g645) & (g901) & (g1501) & (g1503) & (keyx63x)) + ((!ld) & (g645) & (!g901) & (!g1501) & (!g1503) & (!keyx63x)) + ((!ld) & (g645) & (!g901) & (!g1501) & (!g1503) & (keyx63x)) + ((!ld) & (g645) & (!g901) & (g1501) & (g1503) & (!keyx63x)) + ((!ld) & (g645) & (!g901) & (g1501) & (g1503) & (keyx63x)) + ((!ld) & (g645) & (g901) & (!g1501) & (g1503) & (!keyx63x)) + ((!ld) & (g645) & (g901) & (!g1501) & (g1503) & (keyx63x)) + ((!ld) & (g645) & (g901) & (g1501) & (!g1503) & (!keyx63x)) + ((!ld) & (g645) & (g901) & (g1501) & (!g1503) & (keyx63x)) + ((ld) & (!g645) & (!g901) & (!g1501) & (!g1503) & (keyx63x)) + ((ld) & (!g645) & (!g901) & (!g1501) & (g1503) & (keyx63x)) + ((ld) & (!g645) & (!g901) & (g1501) & (!g1503) & (keyx63x)) + ((ld) & (!g645) & (!g901) & (g1501) & (g1503) & (keyx63x)) + ((ld) & (!g645) & (g901) & (!g1501) & (!g1503) & (keyx63x)) + ((ld) & (!g645) & (g901) & (!g1501) & (g1503) & (keyx63x)) + ((ld) & (!g645) & (g901) & (g1501) & (!g1503) & (keyx63x)) + ((ld) & (!g645) & (g901) & (g1501) & (g1503) & (keyx63x)) + ((ld) & (g645) & (!g901) & (!g1501) & (!g1503) & (keyx63x)) + ((ld) & (g645) & (!g901) & (!g1501) & (g1503) & (keyx63x)) + ((ld) & (g645) & (!g901) & (g1501) & (!g1503) & (keyx63x)) + ((ld) & (g645) & (!g901) & (g1501) & (g1503) & (keyx63x)) + ((ld) & (g645) & (g901) & (!g1501) & (!g1503) & (keyx63x)) + ((ld) & (g645) & (g901) & (!g1501) & (g1503) & (keyx63x)) + ((ld) & (g645) & (g901) & (g1501) & (!g1503) & (keyx63x)) + ((ld) & (g645) & (g901) & (g1501) & (g1503) & (keyx63x)));
	assign g1618 = (((!sk[67]) & (!g964) & (g1156)) + ((!sk[67]) & (g964) & (g1156)) + ((sk[67]) & (!g964) & (g1156)) + ((sk[67]) & (g964) & (!g1156)));
	assign g2146 = (((!sk[68]) & (!ld) & (text_inx96x) & (!g1619)) + ((!sk[68]) & (!ld) & (text_inx96x) & (g1619)) + ((!sk[68]) & (ld) & (!text_inx96x) & (g1619)) + ((!sk[68]) & (ld) & (text_inx96x) & (!g1619)) + ((!sk[68]) & (ld) & (text_inx96x) & (g1619)) + ((sk[68]) & (!ld) & (!text_inx96x) & (g1619)) + ((sk[68]) & (!ld) & (text_inx96x) & (g1619)) + ((sk[68]) & (ld) & (text_inx96x) & (!g1619)) + ((sk[68]) & (ld) & (text_inx96x) & (g1619)));
	assign g1620 = (((!g916) & (!g1107) & (!g1163) & (!g1333) & (g1618) & (!g1619)) + ((!g916) & (!g1107) & (!g1163) & (!g1333) & (g1618) & (g1619)) + ((!g916) & (!g1107) & (!g1163) & (g1333) & (!g1618) & (!g1619)) + ((!g916) & (!g1107) & (!g1163) & (g1333) & (!g1618) & (g1619)) + ((!g916) & (!g1107) & (g1163) & (!g1333) & (!g1618) & (g1619)) + ((!g916) & (!g1107) & (g1163) & (!g1333) & (g1618) & (g1619)) + ((!g916) & (!g1107) & (g1163) & (g1333) & (!g1618) & (g1619)) + ((!g916) & (!g1107) & (g1163) & (g1333) & (g1618) & (g1619)) + ((!g916) & (g1107) & (!g1163) & (!g1333) & (!g1618) & (!g1619)) + ((!g916) & (g1107) & (!g1163) & (!g1333) & (!g1618) & (g1619)) + ((!g916) & (g1107) & (!g1163) & (g1333) & (g1618) & (!g1619)) + ((!g916) & (g1107) & (!g1163) & (g1333) & (g1618) & (g1619)) + ((!g916) & (g1107) & (g1163) & (!g1333) & (!g1618) & (g1619)) + ((!g916) & (g1107) & (g1163) & (!g1333) & (g1618) & (g1619)) + ((!g916) & (g1107) & (g1163) & (g1333) & (!g1618) & (g1619)) + ((!g916) & (g1107) & (g1163) & (g1333) & (g1618) & (g1619)) + ((g916) & (!g1107) & (!g1163) & (!g1333) & (!g1618) & (!g1619)) + ((g916) & (!g1107) & (!g1163) & (!g1333) & (!g1618) & (g1619)) + ((g916) & (!g1107) & (!g1163) & (g1333) & (g1618) & (!g1619)) + ((g916) & (!g1107) & (!g1163) & (g1333) & (g1618) & (g1619)) + ((g916) & (!g1107) & (g1163) & (!g1333) & (!g1618) & (!g1619)) + ((g916) & (!g1107) & (g1163) & (!g1333) & (g1618) & (!g1619)) + ((g916) & (!g1107) & (g1163) & (g1333) & (!g1618) & (!g1619)) + ((g916) & (!g1107) & (g1163) & (g1333) & (g1618) & (!g1619)) + ((g916) & (g1107) & (!g1163) & (!g1333) & (g1618) & (!g1619)) + ((g916) & (g1107) & (!g1163) & (!g1333) & (g1618) & (g1619)) + ((g916) & (g1107) & (!g1163) & (g1333) & (!g1618) & (!g1619)) + ((g916) & (g1107) & (!g1163) & (g1333) & (!g1618) & (g1619)) + ((g916) & (g1107) & (g1163) & (!g1333) & (!g1618) & (!g1619)) + ((g916) & (g1107) & (g1163) & (!g1333) & (g1618) & (!g1619)) + ((g916) & (g1107) & (g1163) & (g1333) & (!g1618) & (!g1619)) + ((g916) & (g1107) & (g1163) & (g1333) & (g1618) & (!g1619)));
	assign g2147 = (((!ld) & (!text_inx97x) & (sk[70]) & (g1621)) + ((!ld) & (text_inx97x) & (!sk[70]) & (!g1621)) + ((!ld) & (text_inx97x) & (!sk[70]) & (g1621)) + ((!ld) & (text_inx97x) & (sk[70]) & (g1621)) + ((ld) & (!text_inx97x) & (!sk[70]) & (g1621)) + ((ld) & (text_inx97x) & (!sk[70]) & (!g1621)) + ((ld) & (text_inx97x) & (!sk[70]) & (g1621)) + ((ld) & (text_inx97x) & (sk[70]) & (!g1621)) + ((ld) & (text_inx97x) & (sk[70]) & (g1621)));
	assign g1622 = (((!g986) & (!g1050) & (sk[71]) & (g1107)) + ((!g986) & (g1050) & (!sk[71]) & (!g1107)) + ((!g986) & (g1050) & (!sk[71]) & (g1107)) + ((!g986) & (g1050) & (sk[71]) & (!g1107)) + ((g986) & (!g1050) & (!sk[71]) & (g1107)) + ((g986) & (!g1050) & (sk[71]) & (!g1107)) + ((g986) & (g1050) & (!sk[71]) & (!g1107)) + ((g986) & (g1050) & (!sk[71]) & (g1107)) + ((g986) & (g1050) & (sk[71]) & (g1107)));
	assign g1623 = (((!g915) & (!g923) & (!g964) & (sk[72]) & (!g1114) & (g1156)) + ((!g915) & (!g923) & (!g964) & (sk[72]) & (g1114) & (!g1156)) + ((!g915) & (!g923) & (g964) & (sk[72]) & (!g1114) & (!g1156)) + ((!g915) & (!g923) & (g964) & (sk[72]) & (g1114) & (g1156)) + ((!g915) & (g923) & (!g964) & (!sk[72]) & (!g1114) & (!g1156)) + ((!g915) & (g923) & (!g964) & (!sk[72]) & (!g1114) & (g1156)) + ((!g915) & (g923) & (!g964) & (!sk[72]) & (g1114) & (!g1156)) + ((!g915) & (g923) & (!g964) & (!sk[72]) & (g1114) & (g1156)) + ((!g915) & (g923) & (!g964) & (sk[72]) & (!g1114) & (!g1156)) + ((!g915) & (g923) & (!g964) & (sk[72]) & (g1114) & (g1156)) + ((!g915) & (g923) & (g964) & (!sk[72]) & (!g1114) & (!g1156)) + ((!g915) & (g923) & (g964) & (!sk[72]) & (!g1114) & (g1156)) + ((!g915) & (g923) & (g964) & (!sk[72]) & (g1114) & (!g1156)) + ((!g915) & (g923) & (g964) & (!sk[72]) & (g1114) & (g1156)) + ((!g915) & (g923) & (g964) & (sk[72]) & (!g1114) & (g1156)) + ((!g915) & (g923) & (g964) & (sk[72]) & (g1114) & (!g1156)) + ((g915) & (!g923) & (!g964) & (!sk[72]) & (!g1114) & (!g1156)) + ((g915) & (!g923) & (!g964) & (!sk[72]) & (!g1114) & (g1156)) + ((g915) & (!g923) & (!g964) & (!sk[72]) & (g1114) & (!g1156)) + ((g915) & (!g923) & (!g964) & (!sk[72]) & (g1114) & (g1156)) + ((g915) & (!g923) & (!g964) & (sk[72]) & (!g1114) & (!g1156)) + ((g915) & (!g923) & (!g964) & (sk[72]) & (g1114) & (g1156)) + ((g915) & (!g923) & (g964) & (!sk[72]) & (!g1114) & (!g1156)) + ((g915) & (!g923) & (g964) & (!sk[72]) & (!g1114) & (g1156)) + ((g915) & (!g923) & (g964) & (!sk[72]) & (g1114) & (!g1156)) + ((g915) & (!g923) & (g964) & (!sk[72]) & (g1114) & (g1156)) + ((g915) & (!g923) & (g964) & (sk[72]) & (!g1114) & (g1156)) + ((g915) & (!g923) & (g964) & (sk[72]) & (g1114) & (!g1156)) + ((g915) & (g923) & (!g964) & (!sk[72]) & (!g1114) & (!g1156)) + ((g915) & (g923) & (!g964) & (!sk[72]) & (!g1114) & (g1156)) + ((g915) & (g923) & (!g964) & (!sk[72]) & (g1114) & (!g1156)) + ((g915) & (g923) & (!g964) & (!sk[72]) & (g1114) & (g1156)) + ((g915) & (g923) & (!g964) & (sk[72]) & (!g1114) & (g1156)) + ((g915) & (g923) & (!g964) & (sk[72]) & (g1114) & (!g1156)) + ((g915) & (g923) & (g964) & (!sk[72]) & (!g1114) & (!g1156)) + ((g915) & (g923) & (g964) & (!sk[72]) & (!g1114) & (g1156)) + ((g915) & (g923) & (g964) & (!sk[72]) & (g1114) & (!g1156)) + ((g915) & (g923) & (g964) & (!sk[72]) & (g1114) & (g1156)) + ((g915) & (g923) & (g964) & (sk[72]) & (!g1114) & (!g1156)) + ((g915) & (g923) & (g964) & (sk[72]) & (g1114) & (g1156)));
	assign g1624 = (((!g923) & (!g1163) & (!g1621) & (!g1622) & (sk[73]) & (g1623)) + ((!g923) & (!g1163) & (!g1621) & (g1622) & (sk[73]) & (!g1623)) + ((!g923) & (!g1163) & (g1621) & (!g1622) & (sk[73]) & (g1623)) + ((!g923) & (!g1163) & (g1621) & (g1622) & (sk[73]) & (!g1623)) + ((!g923) & (g1163) & (!g1621) & (!g1622) & (!sk[73]) & (!g1623)) + ((!g923) & (g1163) & (!g1621) & (!g1622) & (!sk[73]) & (g1623)) + ((!g923) & (g1163) & (!g1621) & (g1622) & (!sk[73]) & (!g1623)) + ((!g923) & (g1163) & (!g1621) & (g1622) & (!sk[73]) & (g1623)) + ((!g923) & (g1163) & (g1621) & (!g1622) & (!sk[73]) & (!g1623)) + ((!g923) & (g1163) & (g1621) & (!g1622) & (!sk[73]) & (g1623)) + ((!g923) & (g1163) & (g1621) & (!g1622) & (sk[73]) & (!g1623)) + ((!g923) & (g1163) & (g1621) & (!g1622) & (sk[73]) & (g1623)) + ((!g923) & (g1163) & (g1621) & (g1622) & (!sk[73]) & (!g1623)) + ((!g923) & (g1163) & (g1621) & (g1622) & (!sk[73]) & (g1623)) + ((!g923) & (g1163) & (g1621) & (g1622) & (sk[73]) & (!g1623)) + ((!g923) & (g1163) & (g1621) & (g1622) & (sk[73]) & (g1623)) + ((g923) & (!g1163) & (!g1621) & (!g1622) & (!sk[73]) & (!g1623)) + ((g923) & (!g1163) & (!g1621) & (!g1622) & (!sk[73]) & (g1623)) + ((g923) & (!g1163) & (!g1621) & (!g1622) & (sk[73]) & (g1623)) + ((g923) & (!g1163) & (!g1621) & (g1622) & (!sk[73]) & (!g1623)) + ((g923) & (!g1163) & (!g1621) & (g1622) & (!sk[73]) & (g1623)) + ((g923) & (!g1163) & (!g1621) & (g1622) & (sk[73]) & (!g1623)) + ((g923) & (!g1163) & (g1621) & (!g1622) & (!sk[73]) & (!g1623)) + ((g923) & (!g1163) & (g1621) & (!g1622) & (!sk[73]) & (g1623)) + ((g923) & (!g1163) & (g1621) & (!g1622) & (sk[73]) & (g1623)) + ((g923) & (!g1163) & (g1621) & (g1622) & (!sk[73]) & (!g1623)) + ((g923) & (!g1163) & (g1621) & (g1622) & (!sk[73]) & (g1623)) + ((g923) & (!g1163) & (g1621) & (g1622) & (sk[73]) & (!g1623)) + ((g923) & (g1163) & (!g1621) & (!g1622) & (!sk[73]) & (!g1623)) + ((g923) & (g1163) & (!g1621) & (!g1622) & (!sk[73]) & (g1623)) + ((g923) & (g1163) & (!g1621) & (!g1622) & (sk[73]) & (!g1623)) + ((g923) & (g1163) & (!g1621) & (!g1622) & (sk[73]) & (g1623)) + ((g923) & (g1163) & (!g1621) & (g1622) & (!sk[73]) & (!g1623)) + ((g923) & (g1163) & (!g1621) & (g1622) & (!sk[73]) & (g1623)) + ((g923) & (g1163) & (!g1621) & (g1622) & (sk[73]) & (!g1623)) + ((g923) & (g1163) & (!g1621) & (g1622) & (sk[73]) & (g1623)) + ((g923) & (g1163) & (g1621) & (!g1622) & (!sk[73]) & (!g1623)) + ((g923) & (g1163) & (g1621) & (!g1622) & (!sk[73]) & (g1623)) + ((g923) & (g1163) & (g1621) & (g1622) & (!sk[73]) & (!g1623)) + ((g923) & (g1163) & (g1621) & (g1622) & (!sk[73]) & (g1623)));
	assign g2148 = (((!ld) & (!sk[74]) & (text_inx98x) & (!g1625)) + ((!ld) & (!sk[74]) & (text_inx98x) & (g1625)) + ((!ld) & (sk[74]) & (!text_inx98x) & (g1625)) + ((!ld) & (sk[74]) & (text_inx98x) & (g1625)) + ((ld) & (!sk[74]) & (!text_inx98x) & (g1625)) + ((ld) & (!sk[74]) & (text_inx98x) & (!g1625)) + ((ld) & (!sk[74]) & (text_inx98x) & (g1625)) + ((ld) & (sk[74]) & (text_inx98x) & (!g1625)) + ((ld) & (sk[74]) & (text_inx98x) & (g1625)));
	assign g1626 = (((!g930) & (!g993) & (!g1114) & (!g1163) & (g1541) & (!g1625)) + ((!g930) & (!g993) & (!g1114) & (!g1163) & (g1541) & (g1625)) + ((!g930) & (!g993) & (!g1114) & (g1163) & (!g1541) & (g1625)) + ((!g930) & (!g993) & (!g1114) & (g1163) & (g1541) & (g1625)) + ((!g930) & (!g993) & (g1114) & (!g1163) & (!g1541) & (!g1625)) + ((!g930) & (!g993) & (g1114) & (!g1163) & (!g1541) & (g1625)) + ((!g930) & (!g993) & (g1114) & (g1163) & (!g1541) & (g1625)) + ((!g930) & (!g993) & (g1114) & (g1163) & (g1541) & (g1625)) + ((!g930) & (g993) & (!g1114) & (!g1163) & (!g1541) & (!g1625)) + ((!g930) & (g993) & (!g1114) & (!g1163) & (!g1541) & (g1625)) + ((!g930) & (g993) & (!g1114) & (g1163) & (!g1541) & (g1625)) + ((!g930) & (g993) & (!g1114) & (g1163) & (g1541) & (g1625)) + ((!g930) & (g993) & (g1114) & (!g1163) & (g1541) & (!g1625)) + ((!g930) & (g993) & (g1114) & (!g1163) & (g1541) & (g1625)) + ((!g930) & (g993) & (g1114) & (g1163) & (!g1541) & (g1625)) + ((!g930) & (g993) & (g1114) & (g1163) & (g1541) & (g1625)) + ((g930) & (!g993) & (!g1114) & (!g1163) & (!g1541) & (!g1625)) + ((g930) & (!g993) & (!g1114) & (!g1163) & (!g1541) & (g1625)) + ((g930) & (!g993) & (!g1114) & (g1163) & (!g1541) & (!g1625)) + ((g930) & (!g993) & (!g1114) & (g1163) & (g1541) & (!g1625)) + ((g930) & (!g993) & (g1114) & (!g1163) & (g1541) & (!g1625)) + ((g930) & (!g993) & (g1114) & (!g1163) & (g1541) & (g1625)) + ((g930) & (!g993) & (g1114) & (g1163) & (!g1541) & (!g1625)) + ((g930) & (!g993) & (g1114) & (g1163) & (g1541) & (!g1625)) + ((g930) & (g993) & (!g1114) & (!g1163) & (g1541) & (!g1625)) + ((g930) & (g993) & (!g1114) & (!g1163) & (g1541) & (g1625)) + ((g930) & (g993) & (!g1114) & (g1163) & (!g1541) & (!g1625)) + ((g930) & (g993) & (!g1114) & (g1163) & (g1541) & (!g1625)) + ((g930) & (g993) & (g1114) & (!g1163) & (!g1541) & (!g1625)) + ((g930) & (g993) & (g1114) & (!g1163) & (!g1541) & (g1625)) + ((g930) & (g993) & (g1114) & (g1163) & (!g1541) & (!g1625)) + ((g930) & (g993) & (g1114) & (g1163) & (g1541) & (!g1625)));
	assign g2149 = (((!sk[76]) & (!ld) & (text_inx99x) & (!g1627)) + ((!sk[76]) & (!ld) & (text_inx99x) & (g1627)) + ((!sk[76]) & (ld) & (!text_inx99x) & (g1627)) + ((!sk[76]) & (ld) & (text_inx99x) & (!g1627)) + ((!sk[76]) & (ld) & (text_inx99x) & (g1627)) + ((sk[76]) & (!ld) & (!text_inx99x) & (g1627)) + ((sk[76]) & (!ld) & (text_inx99x) & (g1627)) + ((sk[76]) & (ld) & (text_inx99x) & (!g1627)) + ((sk[76]) & (ld) & (text_inx99x) & (g1627)));
	assign g1628 = (((!g929) & (!g937) & (!g1000) & (sk[77]) & (!g1064) & (g1128)) + ((!g929) & (!g937) & (!g1000) & (sk[77]) & (g1064) & (!g1128)) + ((!g929) & (!g937) & (g1000) & (sk[77]) & (!g1064) & (!g1128)) + ((!g929) & (!g937) & (g1000) & (sk[77]) & (g1064) & (g1128)) + ((!g929) & (g937) & (!g1000) & (!sk[77]) & (!g1064) & (!g1128)) + ((!g929) & (g937) & (!g1000) & (!sk[77]) & (!g1064) & (g1128)) + ((!g929) & (g937) & (!g1000) & (!sk[77]) & (g1064) & (!g1128)) + ((!g929) & (g937) & (!g1000) & (!sk[77]) & (g1064) & (g1128)) + ((!g929) & (g937) & (!g1000) & (sk[77]) & (!g1064) & (!g1128)) + ((!g929) & (g937) & (!g1000) & (sk[77]) & (g1064) & (g1128)) + ((!g929) & (g937) & (g1000) & (!sk[77]) & (!g1064) & (!g1128)) + ((!g929) & (g937) & (g1000) & (!sk[77]) & (!g1064) & (g1128)) + ((!g929) & (g937) & (g1000) & (!sk[77]) & (g1064) & (!g1128)) + ((!g929) & (g937) & (g1000) & (!sk[77]) & (g1064) & (g1128)) + ((!g929) & (g937) & (g1000) & (sk[77]) & (!g1064) & (g1128)) + ((!g929) & (g937) & (g1000) & (sk[77]) & (g1064) & (!g1128)) + ((g929) & (!g937) & (!g1000) & (!sk[77]) & (!g1064) & (!g1128)) + ((g929) & (!g937) & (!g1000) & (!sk[77]) & (!g1064) & (g1128)) + ((g929) & (!g937) & (!g1000) & (!sk[77]) & (g1064) & (!g1128)) + ((g929) & (!g937) & (!g1000) & (!sk[77]) & (g1064) & (g1128)) + ((g929) & (!g937) & (!g1000) & (sk[77]) & (!g1064) & (!g1128)) + ((g929) & (!g937) & (!g1000) & (sk[77]) & (g1064) & (g1128)) + ((g929) & (!g937) & (g1000) & (!sk[77]) & (!g1064) & (!g1128)) + ((g929) & (!g937) & (g1000) & (!sk[77]) & (!g1064) & (g1128)) + ((g929) & (!g937) & (g1000) & (!sk[77]) & (g1064) & (!g1128)) + ((g929) & (!g937) & (g1000) & (!sk[77]) & (g1064) & (g1128)) + ((g929) & (!g937) & (g1000) & (sk[77]) & (!g1064) & (g1128)) + ((g929) & (!g937) & (g1000) & (sk[77]) & (g1064) & (!g1128)) + ((g929) & (g937) & (!g1000) & (!sk[77]) & (!g1064) & (!g1128)) + ((g929) & (g937) & (!g1000) & (!sk[77]) & (!g1064) & (g1128)) + ((g929) & (g937) & (!g1000) & (!sk[77]) & (g1064) & (!g1128)) + ((g929) & (g937) & (!g1000) & (!sk[77]) & (g1064) & (g1128)) + ((g929) & (g937) & (!g1000) & (sk[77]) & (!g1064) & (g1128)) + ((g929) & (g937) & (!g1000) & (sk[77]) & (g1064) & (!g1128)) + ((g929) & (g937) & (g1000) & (!sk[77]) & (!g1064) & (!g1128)) + ((g929) & (g937) & (g1000) & (!sk[77]) & (!g1064) & (g1128)) + ((g929) & (g937) & (g1000) & (!sk[77]) & (g1064) & (!g1128)) + ((g929) & (g937) & (g1000) & (!sk[77]) & (g1064) & (g1128)) + ((g929) & (g937) & (g1000) & (sk[77]) & (!g1064) & (!g1128)) + ((g929) & (g937) & (g1000) & (sk[77]) & (g1064) & (g1128)));
	assign g1629 = (((!g937) & (!g1121) & (!g1163) & (!g1618) & (!g1627) & (g1628)) + ((!g937) & (!g1121) & (!g1163) & (!g1618) & (g1627) & (g1628)) + ((!g937) & (!g1121) & (!g1163) & (g1618) & (!g1627) & (!g1628)) + ((!g937) & (!g1121) & (!g1163) & (g1618) & (g1627) & (!g1628)) + ((!g937) & (!g1121) & (g1163) & (!g1618) & (g1627) & (!g1628)) + ((!g937) & (!g1121) & (g1163) & (!g1618) & (g1627) & (g1628)) + ((!g937) & (!g1121) & (g1163) & (g1618) & (g1627) & (!g1628)) + ((!g937) & (!g1121) & (g1163) & (g1618) & (g1627) & (g1628)) + ((!g937) & (g1121) & (!g1163) & (!g1618) & (!g1627) & (!g1628)) + ((!g937) & (g1121) & (!g1163) & (!g1618) & (g1627) & (!g1628)) + ((!g937) & (g1121) & (!g1163) & (g1618) & (!g1627) & (g1628)) + ((!g937) & (g1121) & (!g1163) & (g1618) & (g1627) & (g1628)) + ((!g937) & (g1121) & (g1163) & (!g1618) & (g1627) & (!g1628)) + ((!g937) & (g1121) & (g1163) & (!g1618) & (g1627) & (g1628)) + ((!g937) & (g1121) & (g1163) & (g1618) & (g1627) & (!g1628)) + ((!g937) & (g1121) & (g1163) & (g1618) & (g1627) & (g1628)) + ((g937) & (!g1121) & (!g1163) & (!g1618) & (!g1627) & (g1628)) + ((g937) & (!g1121) & (!g1163) & (!g1618) & (g1627) & (g1628)) + ((g937) & (!g1121) & (!g1163) & (g1618) & (!g1627) & (!g1628)) + ((g937) & (!g1121) & (!g1163) & (g1618) & (g1627) & (!g1628)) + ((g937) & (!g1121) & (g1163) & (!g1618) & (!g1627) & (!g1628)) + ((g937) & (!g1121) & (g1163) & (!g1618) & (!g1627) & (g1628)) + ((g937) & (!g1121) & (g1163) & (g1618) & (!g1627) & (!g1628)) + ((g937) & (!g1121) & (g1163) & (g1618) & (!g1627) & (g1628)) + ((g937) & (g1121) & (!g1163) & (!g1618) & (!g1627) & (!g1628)) + ((g937) & (g1121) & (!g1163) & (!g1618) & (g1627) & (!g1628)) + ((g937) & (g1121) & (!g1163) & (g1618) & (!g1627) & (g1628)) + ((g937) & (g1121) & (!g1163) & (g1618) & (g1627) & (g1628)) + ((g937) & (g1121) & (g1163) & (!g1618) & (!g1627) & (!g1628)) + ((g937) & (g1121) & (g1163) & (!g1618) & (!g1627) & (g1628)) + ((g937) & (g1121) & (g1163) & (g1618) & (!g1627) & (!g1628)) + ((g937) & (g1121) & (g1163) & (g1618) & (!g1627) & (g1628)));
	assign g2150 = (((!sk[79]) & (!ld) & (text_inx102x) & (!g1630)) + ((!sk[79]) & (!ld) & (text_inx102x) & (g1630)) + ((!sk[79]) & (ld) & (!text_inx102x) & (g1630)) + ((!sk[79]) & (ld) & (text_inx102x) & (!g1630)) + ((!sk[79]) & (ld) & (text_inx102x) & (g1630)) + ((sk[79]) & (!ld) & (!text_inx102x) & (g1630)) + ((sk[79]) & (!ld) & (text_inx102x) & (g1630)) + ((sk[79]) & (ld) & (text_inx102x) & (!g1630)) + ((sk[79]) & (ld) & (text_inx102x) & (g1630)));
	assign g1631 = (((!g958) & (!g1021) & (!g1142) & (!g1163) & (g1548) & (!g1630)) + ((!g958) & (!g1021) & (!g1142) & (!g1163) & (g1548) & (g1630)) + ((!g958) & (!g1021) & (!g1142) & (g1163) & (!g1548) & (g1630)) + ((!g958) & (!g1021) & (!g1142) & (g1163) & (g1548) & (g1630)) + ((!g958) & (!g1021) & (g1142) & (!g1163) & (!g1548) & (!g1630)) + ((!g958) & (!g1021) & (g1142) & (!g1163) & (!g1548) & (g1630)) + ((!g958) & (!g1021) & (g1142) & (g1163) & (!g1548) & (g1630)) + ((!g958) & (!g1021) & (g1142) & (g1163) & (g1548) & (g1630)) + ((!g958) & (g1021) & (!g1142) & (!g1163) & (!g1548) & (!g1630)) + ((!g958) & (g1021) & (!g1142) & (!g1163) & (!g1548) & (g1630)) + ((!g958) & (g1021) & (!g1142) & (g1163) & (!g1548) & (g1630)) + ((!g958) & (g1021) & (!g1142) & (g1163) & (g1548) & (g1630)) + ((!g958) & (g1021) & (g1142) & (!g1163) & (g1548) & (!g1630)) + ((!g958) & (g1021) & (g1142) & (!g1163) & (g1548) & (g1630)) + ((!g958) & (g1021) & (g1142) & (g1163) & (!g1548) & (g1630)) + ((!g958) & (g1021) & (g1142) & (g1163) & (g1548) & (g1630)) + ((g958) & (!g1021) & (!g1142) & (!g1163) & (!g1548) & (!g1630)) + ((g958) & (!g1021) & (!g1142) & (!g1163) & (!g1548) & (g1630)) + ((g958) & (!g1021) & (!g1142) & (g1163) & (!g1548) & (!g1630)) + ((g958) & (!g1021) & (!g1142) & (g1163) & (g1548) & (!g1630)) + ((g958) & (!g1021) & (g1142) & (!g1163) & (g1548) & (!g1630)) + ((g958) & (!g1021) & (g1142) & (!g1163) & (g1548) & (g1630)) + ((g958) & (!g1021) & (g1142) & (g1163) & (!g1548) & (!g1630)) + ((g958) & (!g1021) & (g1142) & (g1163) & (g1548) & (!g1630)) + ((g958) & (g1021) & (!g1142) & (!g1163) & (g1548) & (!g1630)) + ((g958) & (g1021) & (!g1142) & (!g1163) & (g1548) & (g1630)) + ((g958) & (g1021) & (!g1142) & (g1163) & (!g1548) & (!g1630)) + ((g958) & (g1021) & (!g1142) & (g1163) & (g1548) & (!g1630)) + ((g958) & (g1021) & (g1142) & (!g1163) & (!g1548) & (!g1630)) + ((g958) & (g1021) & (g1142) & (!g1163) & (!g1548) & (g1630)) + ((g958) & (g1021) & (g1142) & (g1163) & (!g1548) & (!g1630)) + ((g958) & (g1021) & (g1142) & (g1163) & (g1548) & (!g1630)));
	assign g2151 = (((!ld) & (!text_inx101x) & (sk[81]) & (g1632)) + ((!ld) & (text_inx101x) & (!sk[81]) & (!g1632)) + ((!ld) & (text_inx101x) & (!sk[81]) & (g1632)) + ((!ld) & (text_inx101x) & (sk[81]) & (g1632)) + ((ld) & (!text_inx101x) & (!sk[81]) & (g1632)) + ((ld) & (text_inx101x) & (!sk[81]) & (!g1632)) + ((ld) & (text_inx101x) & (!sk[81]) & (g1632)) + ((ld) & (text_inx101x) & (sk[81]) & (!g1632)) + ((ld) & (text_inx101x) & (sk[81]) & (g1632)));
	assign g1633 = (((!g951) & (!g1014) & (!g1135) & (!g1163) & (g1551) & (!g1632)) + ((!g951) & (!g1014) & (!g1135) & (!g1163) & (g1551) & (g1632)) + ((!g951) & (!g1014) & (!g1135) & (g1163) & (!g1551) & (g1632)) + ((!g951) & (!g1014) & (!g1135) & (g1163) & (g1551) & (g1632)) + ((!g951) & (!g1014) & (g1135) & (!g1163) & (!g1551) & (!g1632)) + ((!g951) & (!g1014) & (g1135) & (!g1163) & (!g1551) & (g1632)) + ((!g951) & (!g1014) & (g1135) & (g1163) & (!g1551) & (g1632)) + ((!g951) & (!g1014) & (g1135) & (g1163) & (g1551) & (g1632)) + ((!g951) & (g1014) & (!g1135) & (!g1163) & (!g1551) & (!g1632)) + ((!g951) & (g1014) & (!g1135) & (!g1163) & (!g1551) & (g1632)) + ((!g951) & (g1014) & (!g1135) & (g1163) & (!g1551) & (g1632)) + ((!g951) & (g1014) & (!g1135) & (g1163) & (g1551) & (g1632)) + ((!g951) & (g1014) & (g1135) & (!g1163) & (g1551) & (!g1632)) + ((!g951) & (g1014) & (g1135) & (!g1163) & (g1551) & (g1632)) + ((!g951) & (g1014) & (g1135) & (g1163) & (!g1551) & (g1632)) + ((!g951) & (g1014) & (g1135) & (g1163) & (g1551) & (g1632)) + ((g951) & (!g1014) & (!g1135) & (!g1163) & (!g1551) & (!g1632)) + ((g951) & (!g1014) & (!g1135) & (!g1163) & (!g1551) & (g1632)) + ((g951) & (!g1014) & (!g1135) & (g1163) & (!g1551) & (!g1632)) + ((g951) & (!g1014) & (!g1135) & (g1163) & (g1551) & (!g1632)) + ((g951) & (!g1014) & (g1135) & (!g1163) & (g1551) & (!g1632)) + ((g951) & (!g1014) & (g1135) & (!g1163) & (g1551) & (g1632)) + ((g951) & (!g1014) & (g1135) & (g1163) & (!g1551) & (!g1632)) + ((g951) & (!g1014) & (g1135) & (g1163) & (g1551) & (!g1632)) + ((g951) & (g1014) & (!g1135) & (!g1163) & (g1551) & (!g1632)) + ((g951) & (g1014) & (!g1135) & (!g1163) & (g1551) & (g1632)) + ((g951) & (g1014) & (!g1135) & (g1163) & (!g1551) & (!g1632)) + ((g951) & (g1014) & (!g1135) & (g1163) & (g1551) & (!g1632)) + ((g951) & (g1014) & (g1135) & (!g1163) & (!g1551) & (!g1632)) + ((g951) & (g1014) & (g1135) & (!g1163) & (!g1551) & (g1632)) + ((g951) & (g1014) & (g1135) & (g1163) & (!g1551) & (!g1632)) + ((g951) & (g1014) & (g1135) & (g1163) & (g1551) & (!g1632)));
	assign g2152 = (((!ld) & (!text_inx100x) & (sk[83]) & (g1634)) + ((!ld) & (text_inx100x) & (!sk[83]) & (!g1634)) + ((!ld) & (text_inx100x) & (!sk[83]) & (g1634)) + ((!ld) & (text_inx100x) & (sk[83]) & (g1634)) + ((ld) & (!text_inx100x) & (!sk[83]) & (g1634)) + ((ld) & (text_inx100x) & (!sk[83]) & (!g1634)) + ((ld) & (text_inx100x) & (!sk[83]) & (g1634)) + ((ld) & (text_inx100x) & (sk[83]) & (!g1634)) + ((ld) & (text_inx100x) & (sk[83]) & (g1634)));
	assign g1635 = (((!g1007) & (!g1071) & (!sk[84]) & (g1128) & (!g1156)) + ((!g1007) & (!g1071) & (!sk[84]) & (g1128) & (g1156)) + ((!g1007) & (!g1071) & (sk[84]) & (!g1128) & (g1156)) + ((!g1007) & (!g1071) & (sk[84]) & (g1128) & (!g1156)) + ((!g1007) & (g1071) & (!sk[84]) & (!g1128) & (!g1156)) + ((!g1007) & (g1071) & (!sk[84]) & (!g1128) & (g1156)) + ((!g1007) & (g1071) & (!sk[84]) & (g1128) & (!g1156)) + ((!g1007) & (g1071) & (!sk[84]) & (g1128) & (g1156)) + ((!g1007) & (g1071) & (sk[84]) & (!g1128) & (!g1156)) + ((!g1007) & (g1071) & (sk[84]) & (g1128) & (g1156)) + ((g1007) & (!g1071) & (!sk[84]) & (g1128) & (!g1156)) + ((g1007) & (!g1071) & (!sk[84]) & (g1128) & (g1156)) + ((g1007) & (!g1071) & (sk[84]) & (!g1128) & (!g1156)) + ((g1007) & (!g1071) & (sk[84]) & (g1128) & (g1156)) + ((g1007) & (g1071) & (!sk[84]) & (!g1128) & (!g1156)) + ((g1007) & (g1071) & (!sk[84]) & (!g1128) & (g1156)) + ((g1007) & (g1071) & (!sk[84]) & (g1128) & (!g1156)) + ((g1007) & (g1071) & (!sk[84]) & (g1128) & (g1156)) + ((g1007) & (g1071) & (sk[84]) & (!g1128) & (g1156)) + ((g1007) & (g1071) & (sk[84]) & (g1128) & (!g1156)));
	assign g2153 = (((!ld) & (!sk[85]) & (text_inx103x) & (!g1636)) + ((!ld) & (!sk[85]) & (text_inx103x) & (g1636)) + ((!ld) & (sk[85]) & (!text_inx103x) & (g1636)) + ((!ld) & (sk[85]) & (text_inx103x) & (g1636)) + ((ld) & (!sk[85]) & (!text_inx103x) & (g1636)) + ((ld) & (!sk[85]) & (text_inx103x) & (!g1636)) + ((ld) & (!sk[85]) & (text_inx103x) & (g1636)) + ((ld) & (sk[85]) & (text_inx103x) & (!g1636)) + ((ld) & (sk[85]) & (text_inx103x) & (g1636)));
	assign g1637 = (((!ld) & (!g660) & (sk[86]) & (!g916) & (g1193) & (!keyx64x)) + ((!ld) & (!g660) & (sk[86]) & (!g916) & (g1193) & (keyx64x)) + ((!ld) & (!g660) & (sk[86]) & (g916) & (!g1193) & (!keyx64x)) + ((!ld) & (!g660) & (sk[86]) & (g916) & (!g1193) & (keyx64x)) + ((!ld) & (g660) & (!sk[86]) & (!g916) & (!g1193) & (!keyx64x)) + ((!ld) & (g660) & (!sk[86]) & (!g916) & (!g1193) & (keyx64x)) + ((!ld) & (g660) & (!sk[86]) & (!g916) & (g1193) & (!keyx64x)) + ((!ld) & (g660) & (!sk[86]) & (!g916) & (g1193) & (keyx64x)) + ((!ld) & (g660) & (!sk[86]) & (g916) & (!g1193) & (!keyx64x)) + ((!ld) & (g660) & (!sk[86]) & (g916) & (!g1193) & (keyx64x)) + ((!ld) & (g660) & (!sk[86]) & (g916) & (g1193) & (!keyx64x)) + ((!ld) & (g660) & (!sk[86]) & (g916) & (g1193) & (keyx64x)) + ((!ld) & (g660) & (sk[86]) & (!g916) & (!g1193) & (!keyx64x)) + ((!ld) & (g660) & (sk[86]) & (!g916) & (!g1193) & (keyx64x)) + ((!ld) & (g660) & (sk[86]) & (g916) & (g1193) & (!keyx64x)) + ((!ld) & (g660) & (sk[86]) & (g916) & (g1193) & (keyx64x)) + ((ld) & (!g660) & (!sk[86]) & (!g916) & (!g1193) & (!keyx64x)) + ((ld) & (!g660) & (!sk[86]) & (!g916) & (!g1193) & (keyx64x)) + ((ld) & (!g660) & (!sk[86]) & (!g916) & (g1193) & (!keyx64x)) + ((ld) & (!g660) & (!sk[86]) & (!g916) & (g1193) & (keyx64x)) + ((ld) & (!g660) & (!sk[86]) & (g916) & (!g1193) & (!keyx64x)) + ((ld) & (!g660) & (!sk[86]) & (g916) & (!g1193) & (keyx64x)) + ((ld) & (!g660) & (!sk[86]) & (g916) & (g1193) & (!keyx64x)) + ((ld) & (!g660) & (!sk[86]) & (g916) & (g1193) & (keyx64x)) + ((ld) & (!g660) & (sk[86]) & (!g916) & (!g1193) & (keyx64x)) + ((ld) & (!g660) & (sk[86]) & (!g916) & (g1193) & (keyx64x)) + ((ld) & (!g660) & (sk[86]) & (g916) & (!g1193) & (keyx64x)) + ((ld) & (!g660) & (sk[86]) & (g916) & (g1193) & (keyx64x)) + ((ld) & (g660) & (!sk[86]) & (!g916) & (!g1193) & (!keyx64x)) + ((ld) & (g660) & (!sk[86]) & (!g916) & (!g1193) & (keyx64x)) + ((ld) & (g660) & (!sk[86]) & (!g916) & (g1193) & (!keyx64x)) + ((ld) & (g660) & (!sk[86]) & (!g916) & (g1193) & (keyx64x)) + ((ld) & (g660) & (!sk[86]) & (g916) & (!g1193) & (!keyx64x)) + ((ld) & (g660) & (!sk[86]) & (g916) & (!g1193) & (keyx64x)) + ((ld) & (g660) & (!sk[86]) & (g916) & (g1193) & (!keyx64x)) + ((ld) & (g660) & (!sk[86]) & (g916) & (g1193) & (keyx64x)) + ((ld) & (g660) & (sk[86]) & (!g916) & (!g1193) & (keyx64x)) + ((ld) & (g660) & (sk[86]) & (!g916) & (g1193) & (keyx64x)) + ((ld) & (g660) & (sk[86]) & (g916) & (!g1193) & (keyx64x)) + ((ld) & (g660) & (sk[86]) & (g916) & (g1193) & (keyx64x)));
	assign g1638 = (((!ld) & (!g667) & (!g923) & (g1200) & (sk[87]) & (!keyx65x)) + ((!ld) & (!g667) & (!g923) & (g1200) & (sk[87]) & (keyx65x)) + ((!ld) & (!g667) & (g923) & (!g1200) & (sk[87]) & (!keyx65x)) + ((!ld) & (!g667) & (g923) & (!g1200) & (sk[87]) & (keyx65x)) + ((!ld) & (g667) & (!g923) & (!g1200) & (!sk[87]) & (!keyx65x)) + ((!ld) & (g667) & (!g923) & (!g1200) & (!sk[87]) & (keyx65x)) + ((!ld) & (g667) & (!g923) & (!g1200) & (sk[87]) & (!keyx65x)) + ((!ld) & (g667) & (!g923) & (!g1200) & (sk[87]) & (keyx65x)) + ((!ld) & (g667) & (!g923) & (g1200) & (!sk[87]) & (!keyx65x)) + ((!ld) & (g667) & (!g923) & (g1200) & (!sk[87]) & (keyx65x)) + ((!ld) & (g667) & (g923) & (!g1200) & (!sk[87]) & (!keyx65x)) + ((!ld) & (g667) & (g923) & (!g1200) & (!sk[87]) & (keyx65x)) + ((!ld) & (g667) & (g923) & (g1200) & (!sk[87]) & (!keyx65x)) + ((!ld) & (g667) & (g923) & (g1200) & (!sk[87]) & (keyx65x)) + ((!ld) & (g667) & (g923) & (g1200) & (sk[87]) & (!keyx65x)) + ((!ld) & (g667) & (g923) & (g1200) & (sk[87]) & (keyx65x)) + ((ld) & (!g667) & (!g923) & (!g1200) & (!sk[87]) & (!keyx65x)) + ((ld) & (!g667) & (!g923) & (!g1200) & (!sk[87]) & (keyx65x)) + ((ld) & (!g667) & (!g923) & (!g1200) & (sk[87]) & (keyx65x)) + ((ld) & (!g667) & (!g923) & (g1200) & (!sk[87]) & (!keyx65x)) + ((ld) & (!g667) & (!g923) & (g1200) & (!sk[87]) & (keyx65x)) + ((ld) & (!g667) & (!g923) & (g1200) & (sk[87]) & (keyx65x)) + ((ld) & (!g667) & (g923) & (!g1200) & (!sk[87]) & (!keyx65x)) + ((ld) & (!g667) & (g923) & (!g1200) & (!sk[87]) & (keyx65x)) + ((ld) & (!g667) & (g923) & (!g1200) & (sk[87]) & (keyx65x)) + ((ld) & (!g667) & (g923) & (g1200) & (!sk[87]) & (!keyx65x)) + ((ld) & (!g667) & (g923) & (g1200) & (!sk[87]) & (keyx65x)) + ((ld) & (!g667) & (g923) & (g1200) & (sk[87]) & (keyx65x)) + ((ld) & (g667) & (!g923) & (!g1200) & (!sk[87]) & (!keyx65x)) + ((ld) & (g667) & (!g923) & (!g1200) & (!sk[87]) & (keyx65x)) + ((ld) & (g667) & (!g923) & (!g1200) & (sk[87]) & (keyx65x)) + ((ld) & (g667) & (!g923) & (g1200) & (!sk[87]) & (!keyx65x)) + ((ld) & (g667) & (!g923) & (g1200) & (!sk[87]) & (keyx65x)) + ((ld) & (g667) & (!g923) & (g1200) & (sk[87]) & (keyx65x)) + ((ld) & (g667) & (g923) & (!g1200) & (!sk[87]) & (!keyx65x)) + ((ld) & (g667) & (g923) & (!g1200) & (!sk[87]) & (keyx65x)) + ((ld) & (g667) & (g923) & (!g1200) & (sk[87]) & (keyx65x)) + ((ld) & (g667) & (g923) & (g1200) & (!sk[87]) & (!keyx65x)) + ((ld) & (g667) & (g923) & (g1200) & (!sk[87]) & (keyx65x)) + ((ld) & (g667) & (g923) & (g1200) & (sk[87]) & (keyx65x)));
	assign g1639 = (((!ld) & (!g674) & (sk[88]) & (!g930) & (g1207) & (!keyx66x)) + ((!ld) & (!g674) & (sk[88]) & (!g930) & (g1207) & (keyx66x)) + ((!ld) & (!g674) & (sk[88]) & (g930) & (!g1207) & (!keyx66x)) + ((!ld) & (!g674) & (sk[88]) & (g930) & (!g1207) & (keyx66x)) + ((!ld) & (g674) & (!sk[88]) & (!g930) & (!g1207) & (!keyx66x)) + ((!ld) & (g674) & (!sk[88]) & (!g930) & (!g1207) & (keyx66x)) + ((!ld) & (g674) & (!sk[88]) & (!g930) & (g1207) & (!keyx66x)) + ((!ld) & (g674) & (!sk[88]) & (!g930) & (g1207) & (keyx66x)) + ((!ld) & (g674) & (!sk[88]) & (g930) & (!g1207) & (!keyx66x)) + ((!ld) & (g674) & (!sk[88]) & (g930) & (!g1207) & (keyx66x)) + ((!ld) & (g674) & (!sk[88]) & (g930) & (g1207) & (!keyx66x)) + ((!ld) & (g674) & (!sk[88]) & (g930) & (g1207) & (keyx66x)) + ((!ld) & (g674) & (sk[88]) & (!g930) & (!g1207) & (!keyx66x)) + ((!ld) & (g674) & (sk[88]) & (!g930) & (!g1207) & (keyx66x)) + ((!ld) & (g674) & (sk[88]) & (g930) & (g1207) & (!keyx66x)) + ((!ld) & (g674) & (sk[88]) & (g930) & (g1207) & (keyx66x)) + ((ld) & (!g674) & (!sk[88]) & (!g930) & (!g1207) & (!keyx66x)) + ((ld) & (!g674) & (!sk[88]) & (!g930) & (!g1207) & (keyx66x)) + ((ld) & (!g674) & (!sk[88]) & (!g930) & (g1207) & (!keyx66x)) + ((ld) & (!g674) & (!sk[88]) & (!g930) & (g1207) & (keyx66x)) + ((ld) & (!g674) & (!sk[88]) & (g930) & (!g1207) & (!keyx66x)) + ((ld) & (!g674) & (!sk[88]) & (g930) & (!g1207) & (keyx66x)) + ((ld) & (!g674) & (!sk[88]) & (g930) & (g1207) & (!keyx66x)) + ((ld) & (!g674) & (!sk[88]) & (g930) & (g1207) & (keyx66x)) + ((ld) & (!g674) & (sk[88]) & (!g930) & (!g1207) & (keyx66x)) + ((ld) & (!g674) & (sk[88]) & (!g930) & (g1207) & (keyx66x)) + ((ld) & (!g674) & (sk[88]) & (g930) & (!g1207) & (keyx66x)) + ((ld) & (!g674) & (sk[88]) & (g930) & (g1207) & (keyx66x)) + ((ld) & (g674) & (!sk[88]) & (!g930) & (!g1207) & (!keyx66x)) + ((ld) & (g674) & (!sk[88]) & (!g930) & (!g1207) & (keyx66x)) + ((ld) & (g674) & (!sk[88]) & (!g930) & (g1207) & (!keyx66x)) + ((ld) & (g674) & (!sk[88]) & (!g930) & (g1207) & (keyx66x)) + ((ld) & (g674) & (!sk[88]) & (g930) & (!g1207) & (!keyx66x)) + ((ld) & (g674) & (!sk[88]) & (g930) & (!g1207) & (keyx66x)) + ((ld) & (g674) & (!sk[88]) & (g930) & (g1207) & (!keyx66x)) + ((ld) & (g674) & (!sk[88]) & (g930) & (g1207) & (keyx66x)) + ((ld) & (g674) & (sk[88]) & (!g930) & (!g1207) & (keyx66x)) + ((ld) & (g674) & (sk[88]) & (!g930) & (g1207) & (keyx66x)) + ((ld) & (g674) & (sk[88]) & (g930) & (!g1207) & (keyx66x)) + ((ld) & (g674) & (sk[88]) & (g930) & (g1207) & (keyx66x)));
	assign g1640 = (((!ld) & (!g681) & (sk[89]) & (!g937) & (g1214) & (!keyx67x)) + ((!ld) & (!g681) & (sk[89]) & (!g937) & (g1214) & (keyx67x)) + ((!ld) & (!g681) & (sk[89]) & (g937) & (!g1214) & (!keyx67x)) + ((!ld) & (!g681) & (sk[89]) & (g937) & (!g1214) & (keyx67x)) + ((!ld) & (g681) & (!sk[89]) & (!g937) & (!g1214) & (!keyx67x)) + ((!ld) & (g681) & (!sk[89]) & (!g937) & (!g1214) & (keyx67x)) + ((!ld) & (g681) & (!sk[89]) & (!g937) & (g1214) & (!keyx67x)) + ((!ld) & (g681) & (!sk[89]) & (!g937) & (g1214) & (keyx67x)) + ((!ld) & (g681) & (!sk[89]) & (g937) & (!g1214) & (!keyx67x)) + ((!ld) & (g681) & (!sk[89]) & (g937) & (!g1214) & (keyx67x)) + ((!ld) & (g681) & (!sk[89]) & (g937) & (g1214) & (!keyx67x)) + ((!ld) & (g681) & (!sk[89]) & (g937) & (g1214) & (keyx67x)) + ((!ld) & (g681) & (sk[89]) & (!g937) & (!g1214) & (!keyx67x)) + ((!ld) & (g681) & (sk[89]) & (!g937) & (!g1214) & (keyx67x)) + ((!ld) & (g681) & (sk[89]) & (g937) & (g1214) & (!keyx67x)) + ((!ld) & (g681) & (sk[89]) & (g937) & (g1214) & (keyx67x)) + ((ld) & (!g681) & (!sk[89]) & (!g937) & (!g1214) & (!keyx67x)) + ((ld) & (!g681) & (!sk[89]) & (!g937) & (!g1214) & (keyx67x)) + ((ld) & (!g681) & (!sk[89]) & (!g937) & (g1214) & (!keyx67x)) + ((ld) & (!g681) & (!sk[89]) & (!g937) & (g1214) & (keyx67x)) + ((ld) & (!g681) & (!sk[89]) & (g937) & (!g1214) & (!keyx67x)) + ((ld) & (!g681) & (!sk[89]) & (g937) & (!g1214) & (keyx67x)) + ((ld) & (!g681) & (!sk[89]) & (g937) & (g1214) & (!keyx67x)) + ((ld) & (!g681) & (!sk[89]) & (g937) & (g1214) & (keyx67x)) + ((ld) & (!g681) & (sk[89]) & (!g937) & (!g1214) & (keyx67x)) + ((ld) & (!g681) & (sk[89]) & (!g937) & (g1214) & (keyx67x)) + ((ld) & (!g681) & (sk[89]) & (g937) & (!g1214) & (keyx67x)) + ((ld) & (!g681) & (sk[89]) & (g937) & (g1214) & (keyx67x)) + ((ld) & (g681) & (!sk[89]) & (!g937) & (!g1214) & (!keyx67x)) + ((ld) & (g681) & (!sk[89]) & (!g937) & (!g1214) & (keyx67x)) + ((ld) & (g681) & (!sk[89]) & (!g937) & (g1214) & (!keyx67x)) + ((ld) & (g681) & (!sk[89]) & (!g937) & (g1214) & (keyx67x)) + ((ld) & (g681) & (!sk[89]) & (g937) & (!g1214) & (!keyx67x)) + ((ld) & (g681) & (!sk[89]) & (g937) & (!g1214) & (keyx67x)) + ((ld) & (g681) & (!sk[89]) & (g937) & (g1214) & (!keyx67x)) + ((ld) & (g681) & (!sk[89]) & (g937) & (g1214) & (keyx67x)) + ((ld) & (g681) & (sk[89]) & (!g937) & (!g1214) & (keyx67x)) + ((ld) & (g681) & (sk[89]) & (!g937) & (g1214) & (keyx67x)) + ((ld) & (g681) & (sk[89]) & (g937) & (!g1214) & (keyx67x)) + ((ld) & (g681) & (sk[89]) & (g937) & (g1214) & (keyx67x)));
	assign g1641 = (((!sk[90]) & (!ld) & (g688) & (!g944) & (!g1221) & (!keyx68x)) + ((!sk[90]) & (!ld) & (g688) & (!g944) & (!g1221) & (keyx68x)) + ((!sk[90]) & (!ld) & (g688) & (!g944) & (g1221) & (!keyx68x)) + ((!sk[90]) & (!ld) & (g688) & (!g944) & (g1221) & (keyx68x)) + ((!sk[90]) & (!ld) & (g688) & (g944) & (!g1221) & (!keyx68x)) + ((!sk[90]) & (!ld) & (g688) & (g944) & (!g1221) & (keyx68x)) + ((!sk[90]) & (!ld) & (g688) & (g944) & (g1221) & (!keyx68x)) + ((!sk[90]) & (!ld) & (g688) & (g944) & (g1221) & (keyx68x)) + ((!sk[90]) & (ld) & (!g688) & (!g944) & (!g1221) & (!keyx68x)) + ((!sk[90]) & (ld) & (!g688) & (!g944) & (!g1221) & (keyx68x)) + ((!sk[90]) & (ld) & (!g688) & (!g944) & (g1221) & (!keyx68x)) + ((!sk[90]) & (ld) & (!g688) & (!g944) & (g1221) & (keyx68x)) + ((!sk[90]) & (ld) & (!g688) & (g944) & (!g1221) & (!keyx68x)) + ((!sk[90]) & (ld) & (!g688) & (g944) & (!g1221) & (keyx68x)) + ((!sk[90]) & (ld) & (!g688) & (g944) & (g1221) & (!keyx68x)) + ((!sk[90]) & (ld) & (!g688) & (g944) & (g1221) & (keyx68x)) + ((!sk[90]) & (ld) & (g688) & (!g944) & (!g1221) & (!keyx68x)) + ((!sk[90]) & (ld) & (g688) & (!g944) & (!g1221) & (keyx68x)) + ((!sk[90]) & (ld) & (g688) & (!g944) & (g1221) & (!keyx68x)) + ((!sk[90]) & (ld) & (g688) & (!g944) & (g1221) & (keyx68x)) + ((!sk[90]) & (ld) & (g688) & (g944) & (!g1221) & (!keyx68x)) + ((!sk[90]) & (ld) & (g688) & (g944) & (!g1221) & (keyx68x)) + ((!sk[90]) & (ld) & (g688) & (g944) & (g1221) & (!keyx68x)) + ((!sk[90]) & (ld) & (g688) & (g944) & (g1221) & (keyx68x)) + ((sk[90]) & (!ld) & (!g688) & (!g944) & (g1221) & (!keyx68x)) + ((sk[90]) & (!ld) & (!g688) & (!g944) & (g1221) & (keyx68x)) + ((sk[90]) & (!ld) & (!g688) & (g944) & (!g1221) & (!keyx68x)) + ((sk[90]) & (!ld) & (!g688) & (g944) & (!g1221) & (keyx68x)) + ((sk[90]) & (!ld) & (g688) & (!g944) & (!g1221) & (!keyx68x)) + ((sk[90]) & (!ld) & (g688) & (!g944) & (!g1221) & (keyx68x)) + ((sk[90]) & (!ld) & (g688) & (g944) & (g1221) & (!keyx68x)) + ((sk[90]) & (!ld) & (g688) & (g944) & (g1221) & (keyx68x)) + ((sk[90]) & (ld) & (!g688) & (!g944) & (!g1221) & (keyx68x)) + ((sk[90]) & (ld) & (!g688) & (!g944) & (g1221) & (keyx68x)) + ((sk[90]) & (ld) & (!g688) & (g944) & (!g1221) & (keyx68x)) + ((sk[90]) & (ld) & (!g688) & (g944) & (g1221) & (keyx68x)) + ((sk[90]) & (ld) & (g688) & (!g944) & (!g1221) & (keyx68x)) + ((sk[90]) & (ld) & (g688) & (!g944) & (g1221) & (keyx68x)) + ((sk[90]) & (ld) & (g688) & (g944) & (!g1221) & (keyx68x)) + ((sk[90]) & (ld) & (g688) & (g944) & (g1221) & (keyx68x)));
	assign g1642 = (((!sk[91]) & (!ld) & (g695) & (!g951) & (!g1228) & (!keyx69x)) + ((!sk[91]) & (!ld) & (g695) & (!g951) & (!g1228) & (keyx69x)) + ((!sk[91]) & (!ld) & (g695) & (!g951) & (g1228) & (!keyx69x)) + ((!sk[91]) & (!ld) & (g695) & (!g951) & (g1228) & (keyx69x)) + ((!sk[91]) & (!ld) & (g695) & (g951) & (!g1228) & (!keyx69x)) + ((!sk[91]) & (!ld) & (g695) & (g951) & (!g1228) & (keyx69x)) + ((!sk[91]) & (!ld) & (g695) & (g951) & (g1228) & (!keyx69x)) + ((!sk[91]) & (!ld) & (g695) & (g951) & (g1228) & (keyx69x)) + ((!sk[91]) & (ld) & (!g695) & (!g951) & (!g1228) & (!keyx69x)) + ((!sk[91]) & (ld) & (!g695) & (!g951) & (!g1228) & (keyx69x)) + ((!sk[91]) & (ld) & (!g695) & (!g951) & (g1228) & (!keyx69x)) + ((!sk[91]) & (ld) & (!g695) & (!g951) & (g1228) & (keyx69x)) + ((!sk[91]) & (ld) & (!g695) & (g951) & (!g1228) & (!keyx69x)) + ((!sk[91]) & (ld) & (!g695) & (g951) & (!g1228) & (keyx69x)) + ((!sk[91]) & (ld) & (!g695) & (g951) & (g1228) & (!keyx69x)) + ((!sk[91]) & (ld) & (!g695) & (g951) & (g1228) & (keyx69x)) + ((!sk[91]) & (ld) & (g695) & (!g951) & (!g1228) & (!keyx69x)) + ((!sk[91]) & (ld) & (g695) & (!g951) & (!g1228) & (keyx69x)) + ((!sk[91]) & (ld) & (g695) & (!g951) & (g1228) & (!keyx69x)) + ((!sk[91]) & (ld) & (g695) & (!g951) & (g1228) & (keyx69x)) + ((!sk[91]) & (ld) & (g695) & (g951) & (!g1228) & (!keyx69x)) + ((!sk[91]) & (ld) & (g695) & (g951) & (!g1228) & (keyx69x)) + ((!sk[91]) & (ld) & (g695) & (g951) & (g1228) & (!keyx69x)) + ((!sk[91]) & (ld) & (g695) & (g951) & (g1228) & (keyx69x)) + ((sk[91]) & (!ld) & (!g695) & (!g951) & (g1228) & (!keyx69x)) + ((sk[91]) & (!ld) & (!g695) & (!g951) & (g1228) & (keyx69x)) + ((sk[91]) & (!ld) & (!g695) & (g951) & (!g1228) & (!keyx69x)) + ((sk[91]) & (!ld) & (!g695) & (g951) & (!g1228) & (keyx69x)) + ((sk[91]) & (!ld) & (g695) & (!g951) & (!g1228) & (!keyx69x)) + ((sk[91]) & (!ld) & (g695) & (!g951) & (!g1228) & (keyx69x)) + ((sk[91]) & (!ld) & (g695) & (g951) & (g1228) & (!keyx69x)) + ((sk[91]) & (!ld) & (g695) & (g951) & (g1228) & (keyx69x)) + ((sk[91]) & (ld) & (!g695) & (!g951) & (!g1228) & (keyx69x)) + ((sk[91]) & (ld) & (!g695) & (!g951) & (g1228) & (keyx69x)) + ((sk[91]) & (ld) & (!g695) & (g951) & (!g1228) & (keyx69x)) + ((sk[91]) & (ld) & (!g695) & (g951) & (g1228) & (keyx69x)) + ((sk[91]) & (ld) & (g695) & (!g951) & (!g1228) & (keyx69x)) + ((sk[91]) & (ld) & (g695) & (!g951) & (g1228) & (keyx69x)) + ((sk[91]) & (ld) & (g695) & (g951) & (!g1228) & (keyx69x)) + ((sk[91]) & (ld) & (g695) & (g951) & (g1228) & (keyx69x)));
	assign g1643 = (((!sk[92]) & (!ld) & (g702) & (!g958) & (!g1235) & (!keyx70x)) + ((!sk[92]) & (!ld) & (g702) & (!g958) & (!g1235) & (keyx70x)) + ((!sk[92]) & (!ld) & (g702) & (!g958) & (g1235) & (!keyx70x)) + ((!sk[92]) & (!ld) & (g702) & (!g958) & (g1235) & (keyx70x)) + ((!sk[92]) & (!ld) & (g702) & (g958) & (!g1235) & (!keyx70x)) + ((!sk[92]) & (!ld) & (g702) & (g958) & (!g1235) & (keyx70x)) + ((!sk[92]) & (!ld) & (g702) & (g958) & (g1235) & (!keyx70x)) + ((!sk[92]) & (!ld) & (g702) & (g958) & (g1235) & (keyx70x)) + ((!sk[92]) & (ld) & (!g702) & (!g958) & (!g1235) & (!keyx70x)) + ((!sk[92]) & (ld) & (!g702) & (!g958) & (!g1235) & (keyx70x)) + ((!sk[92]) & (ld) & (!g702) & (!g958) & (g1235) & (!keyx70x)) + ((!sk[92]) & (ld) & (!g702) & (!g958) & (g1235) & (keyx70x)) + ((!sk[92]) & (ld) & (!g702) & (g958) & (!g1235) & (!keyx70x)) + ((!sk[92]) & (ld) & (!g702) & (g958) & (!g1235) & (keyx70x)) + ((!sk[92]) & (ld) & (!g702) & (g958) & (g1235) & (!keyx70x)) + ((!sk[92]) & (ld) & (!g702) & (g958) & (g1235) & (keyx70x)) + ((!sk[92]) & (ld) & (g702) & (!g958) & (!g1235) & (!keyx70x)) + ((!sk[92]) & (ld) & (g702) & (!g958) & (!g1235) & (keyx70x)) + ((!sk[92]) & (ld) & (g702) & (!g958) & (g1235) & (!keyx70x)) + ((!sk[92]) & (ld) & (g702) & (!g958) & (g1235) & (keyx70x)) + ((!sk[92]) & (ld) & (g702) & (g958) & (!g1235) & (!keyx70x)) + ((!sk[92]) & (ld) & (g702) & (g958) & (!g1235) & (keyx70x)) + ((!sk[92]) & (ld) & (g702) & (g958) & (g1235) & (!keyx70x)) + ((!sk[92]) & (ld) & (g702) & (g958) & (g1235) & (keyx70x)) + ((sk[92]) & (!ld) & (!g702) & (!g958) & (g1235) & (!keyx70x)) + ((sk[92]) & (!ld) & (!g702) & (!g958) & (g1235) & (keyx70x)) + ((sk[92]) & (!ld) & (!g702) & (g958) & (!g1235) & (!keyx70x)) + ((sk[92]) & (!ld) & (!g702) & (g958) & (!g1235) & (keyx70x)) + ((sk[92]) & (!ld) & (g702) & (!g958) & (!g1235) & (!keyx70x)) + ((sk[92]) & (!ld) & (g702) & (!g958) & (!g1235) & (keyx70x)) + ((sk[92]) & (!ld) & (g702) & (g958) & (g1235) & (!keyx70x)) + ((sk[92]) & (!ld) & (g702) & (g958) & (g1235) & (keyx70x)) + ((sk[92]) & (ld) & (!g702) & (!g958) & (!g1235) & (keyx70x)) + ((sk[92]) & (ld) & (!g702) & (!g958) & (g1235) & (keyx70x)) + ((sk[92]) & (ld) & (!g702) & (g958) & (!g1235) & (keyx70x)) + ((sk[92]) & (ld) & (!g702) & (g958) & (g1235) & (keyx70x)) + ((sk[92]) & (ld) & (g702) & (!g958) & (!g1235) & (keyx70x)) + ((sk[92]) & (ld) & (g702) & (!g958) & (g1235) & (keyx70x)) + ((sk[92]) & (ld) & (g702) & (g958) & (!g1235) & (keyx70x)) + ((sk[92]) & (ld) & (g702) & (g958) & (g1235) & (keyx70x)));
	assign g1644 = (((!ld) & (!g709) & (!g965) & (sk[93]) & (g1242) & (!keyx71x)) + ((!ld) & (!g709) & (!g965) & (sk[93]) & (g1242) & (keyx71x)) + ((!ld) & (!g709) & (g965) & (sk[93]) & (!g1242) & (!keyx71x)) + ((!ld) & (!g709) & (g965) & (sk[93]) & (!g1242) & (keyx71x)) + ((!ld) & (g709) & (!g965) & (!sk[93]) & (!g1242) & (!keyx71x)) + ((!ld) & (g709) & (!g965) & (!sk[93]) & (!g1242) & (keyx71x)) + ((!ld) & (g709) & (!g965) & (!sk[93]) & (g1242) & (!keyx71x)) + ((!ld) & (g709) & (!g965) & (!sk[93]) & (g1242) & (keyx71x)) + ((!ld) & (g709) & (!g965) & (sk[93]) & (!g1242) & (!keyx71x)) + ((!ld) & (g709) & (!g965) & (sk[93]) & (!g1242) & (keyx71x)) + ((!ld) & (g709) & (g965) & (!sk[93]) & (!g1242) & (!keyx71x)) + ((!ld) & (g709) & (g965) & (!sk[93]) & (!g1242) & (keyx71x)) + ((!ld) & (g709) & (g965) & (!sk[93]) & (g1242) & (!keyx71x)) + ((!ld) & (g709) & (g965) & (!sk[93]) & (g1242) & (keyx71x)) + ((!ld) & (g709) & (g965) & (sk[93]) & (g1242) & (!keyx71x)) + ((!ld) & (g709) & (g965) & (sk[93]) & (g1242) & (keyx71x)) + ((ld) & (!g709) & (!g965) & (!sk[93]) & (!g1242) & (!keyx71x)) + ((ld) & (!g709) & (!g965) & (!sk[93]) & (!g1242) & (keyx71x)) + ((ld) & (!g709) & (!g965) & (!sk[93]) & (g1242) & (!keyx71x)) + ((ld) & (!g709) & (!g965) & (!sk[93]) & (g1242) & (keyx71x)) + ((ld) & (!g709) & (!g965) & (sk[93]) & (!g1242) & (keyx71x)) + ((ld) & (!g709) & (!g965) & (sk[93]) & (g1242) & (keyx71x)) + ((ld) & (!g709) & (g965) & (!sk[93]) & (!g1242) & (!keyx71x)) + ((ld) & (!g709) & (g965) & (!sk[93]) & (!g1242) & (keyx71x)) + ((ld) & (!g709) & (g965) & (!sk[93]) & (g1242) & (!keyx71x)) + ((ld) & (!g709) & (g965) & (!sk[93]) & (g1242) & (keyx71x)) + ((ld) & (!g709) & (g965) & (sk[93]) & (!g1242) & (keyx71x)) + ((ld) & (!g709) & (g965) & (sk[93]) & (g1242) & (keyx71x)) + ((ld) & (g709) & (!g965) & (!sk[93]) & (!g1242) & (!keyx71x)) + ((ld) & (g709) & (!g965) & (!sk[93]) & (!g1242) & (keyx71x)) + ((ld) & (g709) & (!g965) & (!sk[93]) & (g1242) & (!keyx71x)) + ((ld) & (g709) & (!g965) & (!sk[93]) & (g1242) & (keyx71x)) + ((ld) & (g709) & (!g965) & (sk[93]) & (!g1242) & (keyx71x)) + ((ld) & (g709) & (!g965) & (sk[93]) & (g1242) & (keyx71x)) + ((ld) & (g709) & (g965) & (!sk[93]) & (!g1242) & (!keyx71x)) + ((ld) & (g709) & (g965) & (!sk[93]) & (!g1242) & (keyx71x)) + ((ld) & (g709) & (g965) & (!sk[93]) & (g1242) & (!keyx71x)) + ((ld) & (g709) & (g965) & (!sk[93]) & (g1242) & (keyx71x)) + ((ld) & (g709) & (g965) & (sk[93]) & (!g1242) & (keyx71x)) + ((ld) & (g709) & (g965) & (sk[93]) & (g1242) & (keyx71x)));
	assign g2154 = (((!ld) & (!text_inx8x) & (sk[94]) & (g1645)) + ((!ld) & (text_inx8x) & (!sk[94]) & (!g1645)) + ((!ld) & (text_inx8x) & (!sk[94]) & (g1645)) + ((!ld) & (text_inx8x) & (sk[94]) & (g1645)) + ((ld) & (!text_inx8x) & (!sk[94]) & (g1645)) + ((ld) & (text_inx8x) & (!sk[94]) & (!g1645)) + ((ld) & (text_inx8x) & (!sk[94]) & (g1645)) + ((ld) & (text_inx8x) & (sk[94]) & (!g1645)) + ((ld) & (text_inx8x) & (sk[94]) & (g1645)));
	assign g2155 = (((!ld) & (!text_inx9x) & (sk[95]) & (g1646)) + ((!ld) & (text_inx9x) & (!sk[95]) & (!g1646)) + ((!ld) & (text_inx9x) & (!sk[95]) & (g1646)) + ((!ld) & (text_inx9x) & (sk[95]) & (g1646)) + ((ld) & (!text_inx9x) & (!sk[95]) & (g1646)) + ((ld) & (text_inx9x) & (!sk[95]) & (!g1646)) + ((ld) & (text_inx9x) & (!sk[95]) & (g1646)) + ((ld) & (text_inx9x) & (sk[95]) & (!g1646)) + ((ld) & (text_inx9x) & (sk[95]) & (g1646)));
	assign g1647 = (((!g147) & (!sk[96]) & (g282) & (!g346)) + ((!g147) & (!sk[96]) & (g282) & (g346)) + ((!g147) & (sk[96]) & (!g282) & (g346)) + ((!g147) & (sk[96]) & (g282) & (!g346)) + ((g147) & (!sk[96]) & (!g282) & (g346)) + ((g147) & (!sk[96]) & (g282) & (!g346)) + ((g147) & (!sk[96]) & (g282) & (g346)) + ((g147) & (sk[96]) & (!g282) & (!g346)) + ((g147) & (sk[96]) & (g282) & (g346)));
	assign g1648 = (((!g154) & (!g196) & (sk[97]) & (!g211) & (!g219) & (g260)) + ((!g154) & (!g196) & (sk[97]) & (!g211) & (g219) & (!g260)) + ((!g154) & (!g196) & (sk[97]) & (g211) & (!g219) & (!g260)) + ((!g154) & (!g196) & (sk[97]) & (g211) & (g219) & (g260)) + ((!g154) & (g196) & (!sk[97]) & (!g211) & (!g219) & (!g260)) + ((!g154) & (g196) & (!sk[97]) & (!g211) & (!g219) & (g260)) + ((!g154) & (g196) & (!sk[97]) & (!g211) & (g219) & (!g260)) + ((!g154) & (g196) & (!sk[97]) & (!g211) & (g219) & (g260)) + ((!g154) & (g196) & (!sk[97]) & (g211) & (!g219) & (!g260)) + ((!g154) & (g196) & (!sk[97]) & (g211) & (!g219) & (g260)) + ((!g154) & (g196) & (!sk[97]) & (g211) & (g219) & (!g260)) + ((!g154) & (g196) & (!sk[97]) & (g211) & (g219) & (g260)) + ((!g154) & (g196) & (sk[97]) & (!g211) & (!g219) & (!g260)) + ((!g154) & (g196) & (sk[97]) & (!g211) & (g219) & (g260)) + ((!g154) & (g196) & (sk[97]) & (g211) & (!g219) & (g260)) + ((!g154) & (g196) & (sk[97]) & (g211) & (g219) & (!g260)) + ((g154) & (!g196) & (!sk[97]) & (!g211) & (!g219) & (!g260)) + ((g154) & (!g196) & (!sk[97]) & (!g211) & (!g219) & (g260)) + ((g154) & (!g196) & (!sk[97]) & (!g211) & (g219) & (!g260)) + ((g154) & (!g196) & (!sk[97]) & (!g211) & (g219) & (g260)) + ((g154) & (!g196) & (!sk[97]) & (g211) & (!g219) & (!g260)) + ((g154) & (!g196) & (!sk[97]) & (g211) & (!g219) & (g260)) + ((g154) & (!g196) & (!sk[97]) & (g211) & (g219) & (!g260)) + ((g154) & (!g196) & (!sk[97]) & (g211) & (g219) & (g260)) + ((g154) & (!g196) & (sk[97]) & (!g211) & (!g219) & (!g260)) + ((g154) & (!g196) & (sk[97]) & (!g211) & (g219) & (g260)) + ((g154) & (!g196) & (sk[97]) & (g211) & (!g219) & (g260)) + ((g154) & (!g196) & (sk[97]) & (g211) & (g219) & (!g260)) + ((g154) & (g196) & (!sk[97]) & (!g211) & (!g219) & (!g260)) + ((g154) & (g196) & (!sk[97]) & (!g211) & (!g219) & (g260)) + ((g154) & (g196) & (!sk[97]) & (!g211) & (g219) & (!g260)) + ((g154) & (g196) & (!sk[97]) & (!g211) & (g219) & (g260)) + ((g154) & (g196) & (!sk[97]) & (g211) & (!g219) & (!g260)) + ((g154) & (g196) & (!sk[97]) & (g211) & (!g219) & (g260)) + ((g154) & (g196) & (!sk[97]) & (g211) & (g219) & (!g260)) + ((g154) & (g196) & (!sk[97]) & (g211) & (g219) & (g260)) + ((g154) & (g196) & (sk[97]) & (!g211) & (!g219) & (g260)) + ((g154) & (g196) & (sk[97]) & (!g211) & (g219) & (!g260)) + ((g154) & (g196) & (sk[97]) & (g211) & (!g219) & (!g260)) + ((g154) & (g196) & (sk[97]) & (g211) & (g219) & (g260)));
	assign g1649 = (((!g219) & (!g1163) & (!g1646) & (!g1647) & (sk[98]) & (g1648)) + ((!g219) & (!g1163) & (!g1646) & (g1647) & (sk[98]) & (!g1648)) + ((!g219) & (!g1163) & (g1646) & (!g1647) & (sk[98]) & (g1648)) + ((!g219) & (!g1163) & (g1646) & (g1647) & (sk[98]) & (!g1648)) + ((!g219) & (g1163) & (!g1646) & (!g1647) & (!sk[98]) & (!g1648)) + ((!g219) & (g1163) & (!g1646) & (!g1647) & (!sk[98]) & (g1648)) + ((!g219) & (g1163) & (!g1646) & (g1647) & (!sk[98]) & (!g1648)) + ((!g219) & (g1163) & (!g1646) & (g1647) & (!sk[98]) & (g1648)) + ((!g219) & (g1163) & (g1646) & (!g1647) & (!sk[98]) & (!g1648)) + ((!g219) & (g1163) & (g1646) & (!g1647) & (!sk[98]) & (g1648)) + ((!g219) & (g1163) & (g1646) & (!g1647) & (sk[98]) & (!g1648)) + ((!g219) & (g1163) & (g1646) & (!g1647) & (sk[98]) & (g1648)) + ((!g219) & (g1163) & (g1646) & (g1647) & (!sk[98]) & (!g1648)) + ((!g219) & (g1163) & (g1646) & (g1647) & (!sk[98]) & (g1648)) + ((!g219) & (g1163) & (g1646) & (g1647) & (sk[98]) & (!g1648)) + ((!g219) & (g1163) & (g1646) & (g1647) & (sk[98]) & (g1648)) + ((g219) & (!g1163) & (!g1646) & (!g1647) & (!sk[98]) & (!g1648)) + ((g219) & (!g1163) & (!g1646) & (!g1647) & (!sk[98]) & (g1648)) + ((g219) & (!g1163) & (!g1646) & (!g1647) & (sk[98]) & (g1648)) + ((g219) & (!g1163) & (!g1646) & (g1647) & (!sk[98]) & (!g1648)) + ((g219) & (!g1163) & (!g1646) & (g1647) & (!sk[98]) & (g1648)) + ((g219) & (!g1163) & (!g1646) & (g1647) & (sk[98]) & (!g1648)) + ((g219) & (!g1163) & (g1646) & (!g1647) & (!sk[98]) & (!g1648)) + ((g219) & (!g1163) & (g1646) & (!g1647) & (!sk[98]) & (g1648)) + ((g219) & (!g1163) & (g1646) & (!g1647) & (sk[98]) & (g1648)) + ((g219) & (!g1163) & (g1646) & (g1647) & (!sk[98]) & (!g1648)) + ((g219) & (!g1163) & (g1646) & (g1647) & (!sk[98]) & (g1648)) + ((g219) & (!g1163) & (g1646) & (g1647) & (sk[98]) & (!g1648)) + ((g219) & (g1163) & (!g1646) & (!g1647) & (!sk[98]) & (!g1648)) + ((g219) & (g1163) & (!g1646) & (!g1647) & (!sk[98]) & (g1648)) + ((g219) & (g1163) & (!g1646) & (!g1647) & (sk[98]) & (!g1648)) + ((g219) & (g1163) & (!g1646) & (!g1647) & (sk[98]) & (g1648)) + ((g219) & (g1163) & (!g1646) & (g1647) & (!sk[98]) & (!g1648)) + ((g219) & (g1163) & (!g1646) & (g1647) & (!sk[98]) & (g1648)) + ((g219) & (g1163) & (!g1646) & (g1647) & (sk[98]) & (!g1648)) + ((g219) & (g1163) & (!g1646) & (g1647) & (sk[98]) & (g1648)) + ((g219) & (g1163) & (g1646) & (!g1647) & (!sk[98]) & (!g1648)) + ((g219) & (g1163) & (g1646) & (!g1647) & (!sk[98]) & (g1648)) + ((g219) & (g1163) & (g1646) & (g1647) & (!sk[98]) & (!g1648)) + ((g219) & (g1163) & (g1646) & (g1647) & (!sk[98]) & (g1648)));
	assign g2156 = (((!sk[99]) & (!ld) & (text_inx10x) & (!g1650)) + ((!sk[99]) & (!ld) & (text_inx10x) & (g1650)) + ((!sk[99]) & (ld) & (!text_inx10x) & (g1650)) + ((!sk[99]) & (ld) & (text_inx10x) & (!g1650)) + ((!sk[99]) & (ld) & (text_inx10x) & (g1650)) + ((sk[99]) & (!ld) & (!text_inx10x) & (g1650)) + ((sk[99]) & (!ld) & (text_inx10x) & (g1650)) + ((sk[99]) & (ld) & (text_inx10x) & (!g1650)) + ((sk[99]) & (ld) & (text_inx10x) & (g1650)));
	assign g1651 = (((!g154) & (!g289) & (sk[100]) & (g353)) + ((!g154) & (g289) & (!sk[100]) & (!g353)) + ((!g154) & (g289) & (!sk[100]) & (g353)) + ((!g154) & (g289) & (sk[100]) & (!g353)) + ((g154) & (!g289) & (!sk[100]) & (g353)) + ((g154) & (!g289) & (sk[100]) & (!g353)) + ((g154) & (g289) & (!sk[100]) & (!g353)) + ((g154) & (g289) & (!sk[100]) & (g353)) + ((g154) & (g289) & (sk[100]) & (g353)));
	assign g1652 = (((!g161) & (!g218) & (!g226) & (!g1163) & (!g1650) & (g1651)) + ((!g161) & (!g218) & (!g226) & (!g1163) & (g1650) & (g1651)) + ((!g161) & (!g218) & (!g226) & (g1163) & (g1650) & (!g1651)) + ((!g161) & (!g218) & (!g226) & (g1163) & (g1650) & (g1651)) + ((!g161) & (!g218) & (g226) & (!g1163) & (!g1650) & (!g1651)) + ((!g161) & (!g218) & (g226) & (!g1163) & (g1650) & (!g1651)) + ((!g161) & (!g218) & (g226) & (g1163) & (!g1650) & (!g1651)) + ((!g161) & (!g218) & (g226) & (g1163) & (!g1650) & (g1651)) + ((!g161) & (g218) & (!g226) & (!g1163) & (!g1650) & (!g1651)) + ((!g161) & (g218) & (!g226) & (!g1163) & (g1650) & (!g1651)) + ((!g161) & (g218) & (!g226) & (g1163) & (g1650) & (!g1651)) + ((!g161) & (g218) & (!g226) & (g1163) & (g1650) & (g1651)) + ((!g161) & (g218) & (g226) & (!g1163) & (!g1650) & (g1651)) + ((!g161) & (g218) & (g226) & (!g1163) & (g1650) & (g1651)) + ((!g161) & (g218) & (g226) & (g1163) & (!g1650) & (!g1651)) + ((!g161) & (g218) & (g226) & (g1163) & (!g1650) & (g1651)) + ((g161) & (!g218) & (!g226) & (!g1163) & (!g1650) & (!g1651)) + ((g161) & (!g218) & (!g226) & (!g1163) & (g1650) & (!g1651)) + ((g161) & (!g218) & (!g226) & (g1163) & (g1650) & (!g1651)) + ((g161) & (!g218) & (!g226) & (g1163) & (g1650) & (g1651)) + ((g161) & (!g218) & (g226) & (!g1163) & (!g1650) & (g1651)) + ((g161) & (!g218) & (g226) & (!g1163) & (g1650) & (g1651)) + ((g161) & (!g218) & (g226) & (g1163) & (!g1650) & (!g1651)) + ((g161) & (!g218) & (g226) & (g1163) & (!g1650) & (g1651)) + ((g161) & (g218) & (!g226) & (!g1163) & (!g1650) & (g1651)) + ((g161) & (g218) & (!g226) & (!g1163) & (g1650) & (g1651)) + ((g161) & (g218) & (!g226) & (g1163) & (g1650) & (!g1651)) + ((g161) & (g218) & (!g226) & (g1163) & (g1650) & (g1651)) + ((g161) & (g218) & (g226) & (!g1163) & (!g1650) & (!g1651)) + ((g161) & (g218) & (g226) & (!g1163) & (g1650) & (!g1651)) + ((g161) & (g218) & (g226) & (g1163) & (!g1650) & (!g1651)) + ((g161) & (g218) & (g226) & (g1163) & (!g1650) & (g1651)));
	assign g2157 = (((!sk[102]) & (!ld) & (text_inx11x) & (!g1653)) + ((!sk[102]) & (!ld) & (text_inx11x) & (g1653)) + ((!sk[102]) & (ld) & (!text_inx11x) & (g1653)) + ((!sk[102]) & (ld) & (text_inx11x) & (!g1653)) + ((!sk[102]) & (ld) & (text_inx11x) & (g1653)) + ((sk[102]) & (!ld) & (!text_inx11x) & (g1653)) + ((sk[102]) & (!ld) & (text_inx11x) & (g1653)) + ((sk[102]) & (ld) & (text_inx11x) & (!g1653)) + ((sk[102]) & (ld) & (text_inx11x) & (g1653)));
	assign g1654 = (((!sk[103]) & (!g161) & (g296) & (!g360)) + ((!sk[103]) & (!g161) & (g296) & (g360)) + ((!sk[103]) & (g161) & (!g296) & (g360)) + ((!sk[103]) & (g161) & (g296) & (!g360)) + ((!sk[103]) & (g161) & (g296) & (g360)) + ((sk[103]) & (!g161) & (!g296) & (g360)) + ((sk[103]) & (!g161) & (g296) & (!g360)) + ((sk[103]) & (g161) & (!g296) & (!g360)) + ((sk[103]) & (g161) & (g296) & (g360)));
	assign g1655 = (((!sk[104]) & (!g168) & (g196) & (!g225) & (!g233) & (!g260)) + ((!sk[104]) & (!g168) & (g196) & (!g225) & (!g233) & (g260)) + ((!sk[104]) & (!g168) & (g196) & (!g225) & (g233) & (!g260)) + ((!sk[104]) & (!g168) & (g196) & (!g225) & (g233) & (g260)) + ((!sk[104]) & (!g168) & (g196) & (g225) & (!g233) & (!g260)) + ((!sk[104]) & (!g168) & (g196) & (g225) & (!g233) & (g260)) + ((!sk[104]) & (!g168) & (g196) & (g225) & (g233) & (!g260)) + ((!sk[104]) & (!g168) & (g196) & (g225) & (g233) & (g260)) + ((!sk[104]) & (g168) & (!g196) & (!g225) & (!g233) & (!g260)) + ((!sk[104]) & (g168) & (!g196) & (!g225) & (!g233) & (g260)) + ((!sk[104]) & (g168) & (!g196) & (!g225) & (g233) & (!g260)) + ((!sk[104]) & (g168) & (!g196) & (!g225) & (g233) & (g260)) + ((!sk[104]) & (g168) & (!g196) & (g225) & (!g233) & (!g260)) + ((!sk[104]) & (g168) & (!g196) & (g225) & (!g233) & (g260)) + ((!sk[104]) & (g168) & (!g196) & (g225) & (g233) & (!g260)) + ((!sk[104]) & (g168) & (!g196) & (g225) & (g233) & (g260)) + ((!sk[104]) & (g168) & (g196) & (!g225) & (!g233) & (!g260)) + ((!sk[104]) & (g168) & (g196) & (!g225) & (!g233) & (g260)) + ((!sk[104]) & (g168) & (g196) & (!g225) & (g233) & (!g260)) + ((!sk[104]) & (g168) & (g196) & (!g225) & (g233) & (g260)) + ((!sk[104]) & (g168) & (g196) & (g225) & (!g233) & (!g260)) + ((!sk[104]) & (g168) & (g196) & (g225) & (!g233) & (g260)) + ((!sk[104]) & (g168) & (g196) & (g225) & (g233) & (!g260)) + ((!sk[104]) & (g168) & (g196) & (g225) & (g233) & (g260)) + ((sk[104]) & (!g168) & (!g196) & (!g225) & (!g233) & (g260)) + ((sk[104]) & (!g168) & (!g196) & (!g225) & (g233) & (!g260)) + ((sk[104]) & (!g168) & (!g196) & (g225) & (!g233) & (!g260)) + ((sk[104]) & (!g168) & (!g196) & (g225) & (g233) & (g260)) + ((sk[104]) & (!g168) & (g196) & (!g225) & (!g233) & (!g260)) + ((sk[104]) & (!g168) & (g196) & (!g225) & (g233) & (g260)) + ((sk[104]) & (!g168) & (g196) & (g225) & (!g233) & (g260)) + ((sk[104]) & (!g168) & (g196) & (g225) & (g233) & (!g260)) + ((sk[104]) & (g168) & (!g196) & (!g225) & (!g233) & (!g260)) + ((sk[104]) & (g168) & (!g196) & (!g225) & (g233) & (g260)) + ((sk[104]) & (g168) & (!g196) & (g225) & (!g233) & (g260)) + ((sk[104]) & (g168) & (!g196) & (g225) & (g233) & (!g260)) + ((sk[104]) & (g168) & (g196) & (!g225) & (!g233) & (g260)) + ((sk[104]) & (g168) & (g196) & (!g225) & (g233) & (!g260)) + ((sk[104]) & (g168) & (g196) & (g225) & (!g233) & (!g260)) + ((sk[104]) & (g168) & (g196) & (g225) & (g233) & (g260)));
	assign g1656 = (((!g233) & (!g1163) & (!g1653) & (sk[105]) & (!g1654) & (g1655)) + ((!g233) & (!g1163) & (!g1653) & (sk[105]) & (g1654) & (!g1655)) + ((!g233) & (!g1163) & (g1653) & (sk[105]) & (!g1654) & (g1655)) + ((!g233) & (!g1163) & (g1653) & (sk[105]) & (g1654) & (!g1655)) + ((!g233) & (g1163) & (!g1653) & (!sk[105]) & (!g1654) & (!g1655)) + ((!g233) & (g1163) & (!g1653) & (!sk[105]) & (!g1654) & (g1655)) + ((!g233) & (g1163) & (!g1653) & (!sk[105]) & (g1654) & (!g1655)) + ((!g233) & (g1163) & (!g1653) & (!sk[105]) & (g1654) & (g1655)) + ((!g233) & (g1163) & (g1653) & (!sk[105]) & (!g1654) & (!g1655)) + ((!g233) & (g1163) & (g1653) & (!sk[105]) & (!g1654) & (g1655)) + ((!g233) & (g1163) & (g1653) & (!sk[105]) & (g1654) & (!g1655)) + ((!g233) & (g1163) & (g1653) & (!sk[105]) & (g1654) & (g1655)) + ((!g233) & (g1163) & (g1653) & (sk[105]) & (!g1654) & (!g1655)) + ((!g233) & (g1163) & (g1653) & (sk[105]) & (!g1654) & (g1655)) + ((!g233) & (g1163) & (g1653) & (sk[105]) & (g1654) & (!g1655)) + ((!g233) & (g1163) & (g1653) & (sk[105]) & (g1654) & (g1655)) + ((g233) & (!g1163) & (!g1653) & (!sk[105]) & (!g1654) & (!g1655)) + ((g233) & (!g1163) & (!g1653) & (!sk[105]) & (!g1654) & (g1655)) + ((g233) & (!g1163) & (!g1653) & (!sk[105]) & (g1654) & (!g1655)) + ((g233) & (!g1163) & (!g1653) & (!sk[105]) & (g1654) & (g1655)) + ((g233) & (!g1163) & (!g1653) & (sk[105]) & (!g1654) & (g1655)) + ((g233) & (!g1163) & (!g1653) & (sk[105]) & (g1654) & (!g1655)) + ((g233) & (!g1163) & (g1653) & (!sk[105]) & (!g1654) & (!g1655)) + ((g233) & (!g1163) & (g1653) & (!sk[105]) & (!g1654) & (g1655)) + ((g233) & (!g1163) & (g1653) & (!sk[105]) & (g1654) & (!g1655)) + ((g233) & (!g1163) & (g1653) & (!sk[105]) & (g1654) & (g1655)) + ((g233) & (!g1163) & (g1653) & (sk[105]) & (!g1654) & (g1655)) + ((g233) & (!g1163) & (g1653) & (sk[105]) & (g1654) & (!g1655)) + ((g233) & (g1163) & (!g1653) & (!sk[105]) & (!g1654) & (!g1655)) + ((g233) & (g1163) & (!g1653) & (!sk[105]) & (!g1654) & (g1655)) + ((g233) & (g1163) & (!g1653) & (!sk[105]) & (g1654) & (!g1655)) + ((g233) & (g1163) & (!g1653) & (!sk[105]) & (g1654) & (g1655)) + ((g233) & (g1163) & (!g1653) & (sk[105]) & (!g1654) & (!g1655)) + ((g233) & (g1163) & (!g1653) & (sk[105]) & (!g1654) & (g1655)) + ((g233) & (g1163) & (!g1653) & (sk[105]) & (g1654) & (!g1655)) + ((g233) & (g1163) & (!g1653) & (sk[105]) & (g1654) & (g1655)) + ((g233) & (g1163) & (g1653) & (!sk[105]) & (!g1654) & (!g1655)) + ((g233) & (g1163) & (g1653) & (!sk[105]) & (!g1654) & (g1655)) + ((g233) & (g1163) & (g1653) & (!sk[105]) & (g1654) & (!g1655)) + ((g233) & (g1163) & (g1653) & (!sk[105]) & (g1654) & (g1655)));
	assign g2158 = (((!ld) & (!sk[106]) & (text_inx14x) & (!g1657)) + ((!ld) & (!sk[106]) & (text_inx14x) & (g1657)) + ((!ld) & (sk[106]) & (!text_inx14x) & (g1657)) + ((!ld) & (sk[106]) & (text_inx14x) & (g1657)) + ((ld) & (!sk[106]) & (!text_inx14x) & (g1657)) + ((ld) & (!sk[106]) & (text_inx14x) & (!g1657)) + ((ld) & (!sk[106]) & (text_inx14x) & (g1657)) + ((ld) & (sk[106]) & (text_inx14x) & (!g1657)) + ((ld) & (sk[106]) & (text_inx14x) & (g1657)));
	assign g1658 = (((!g182) & (!g317) & (sk[107]) & (g381)) + ((!g182) & (g317) & (!sk[107]) & (!g381)) + ((!g182) & (g317) & (!sk[107]) & (g381)) + ((!g182) & (g317) & (sk[107]) & (!g381)) + ((g182) & (!g317) & (!sk[107]) & (g381)) + ((g182) & (!g317) & (sk[107]) & (!g381)) + ((g182) & (g317) & (!sk[107]) & (!g381)) + ((g182) & (g317) & (!sk[107]) & (g381)) + ((g182) & (g317) & (sk[107]) & (g381)));
	assign g1659 = (((!g189) & (!g246) & (!g254) & (!g1163) & (!g1657) & (g1658)) + ((!g189) & (!g246) & (!g254) & (!g1163) & (g1657) & (g1658)) + ((!g189) & (!g246) & (!g254) & (g1163) & (g1657) & (!g1658)) + ((!g189) & (!g246) & (!g254) & (g1163) & (g1657) & (g1658)) + ((!g189) & (!g246) & (g254) & (!g1163) & (!g1657) & (!g1658)) + ((!g189) & (!g246) & (g254) & (!g1163) & (g1657) & (!g1658)) + ((!g189) & (!g246) & (g254) & (g1163) & (!g1657) & (!g1658)) + ((!g189) & (!g246) & (g254) & (g1163) & (!g1657) & (g1658)) + ((!g189) & (g246) & (!g254) & (!g1163) & (!g1657) & (!g1658)) + ((!g189) & (g246) & (!g254) & (!g1163) & (g1657) & (!g1658)) + ((!g189) & (g246) & (!g254) & (g1163) & (g1657) & (!g1658)) + ((!g189) & (g246) & (!g254) & (g1163) & (g1657) & (g1658)) + ((!g189) & (g246) & (g254) & (!g1163) & (!g1657) & (g1658)) + ((!g189) & (g246) & (g254) & (!g1163) & (g1657) & (g1658)) + ((!g189) & (g246) & (g254) & (g1163) & (!g1657) & (!g1658)) + ((!g189) & (g246) & (g254) & (g1163) & (!g1657) & (g1658)) + ((g189) & (!g246) & (!g254) & (!g1163) & (!g1657) & (!g1658)) + ((g189) & (!g246) & (!g254) & (!g1163) & (g1657) & (!g1658)) + ((g189) & (!g246) & (!g254) & (g1163) & (g1657) & (!g1658)) + ((g189) & (!g246) & (!g254) & (g1163) & (g1657) & (g1658)) + ((g189) & (!g246) & (g254) & (!g1163) & (!g1657) & (g1658)) + ((g189) & (!g246) & (g254) & (!g1163) & (g1657) & (g1658)) + ((g189) & (!g246) & (g254) & (g1163) & (!g1657) & (!g1658)) + ((g189) & (!g246) & (g254) & (g1163) & (!g1657) & (g1658)) + ((g189) & (g246) & (!g254) & (!g1163) & (!g1657) & (g1658)) + ((g189) & (g246) & (!g254) & (!g1163) & (g1657) & (g1658)) + ((g189) & (g246) & (!g254) & (g1163) & (g1657) & (!g1658)) + ((g189) & (g246) & (!g254) & (g1163) & (g1657) & (g1658)) + ((g189) & (g246) & (g254) & (!g1163) & (!g1657) & (!g1658)) + ((g189) & (g246) & (g254) & (!g1163) & (g1657) & (!g1658)) + ((g189) & (g246) & (g254) & (g1163) & (!g1657) & (!g1658)) + ((g189) & (g246) & (g254) & (g1163) & (!g1657) & (g1658)));
	assign g2159 = (((!sk[109]) & (!ld) & (text_inx13x) & (!g1660)) + ((!sk[109]) & (!ld) & (text_inx13x) & (g1660)) + ((!sk[109]) & (ld) & (!text_inx13x) & (g1660)) + ((!sk[109]) & (ld) & (text_inx13x) & (!g1660)) + ((!sk[109]) & (ld) & (text_inx13x) & (g1660)) + ((sk[109]) & (!ld) & (!text_inx13x) & (g1660)) + ((sk[109]) & (!ld) & (text_inx13x) & (g1660)) + ((sk[109]) & (ld) & (text_inx13x) & (!g1660)) + ((sk[109]) & (ld) & (text_inx13x) & (g1660)));
	assign g1661 = (((!g175) & (!g310) & (sk[110]) & (g374)) + ((!g175) & (g310) & (!sk[110]) & (!g374)) + ((!g175) & (g310) & (!sk[110]) & (g374)) + ((!g175) & (g310) & (sk[110]) & (!g374)) + ((g175) & (!g310) & (!sk[110]) & (g374)) + ((g175) & (!g310) & (sk[110]) & (!g374)) + ((g175) & (g310) & (!sk[110]) & (!g374)) + ((g175) & (g310) & (!sk[110]) & (g374)) + ((g175) & (g310) & (sk[110]) & (g374)));
	assign g1662 = (((!g182) & (!g239) & (!g247) & (!g1163) & (!g1660) & (g1661)) + ((!g182) & (!g239) & (!g247) & (!g1163) & (g1660) & (g1661)) + ((!g182) & (!g239) & (!g247) & (g1163) & (g1660) & (!g1661)) + ((!g182) & (!g239) & (!g247) & (g1163) & (g1660) & (g1661)) + ((!g182) & (!g239) & (g247) & (!g1163) & (!g1660) & (!g1661)) + ((!g182) & (!g239) & (g247) & (!g1163) & (g1660) & (!g1661)) + ((!g182) & (!g239) & (g247) & (g1163) & (!g1660) & (!g1661)) + ((!g182) & (!g239) & (g247) & (g1163) & (!g1660) & (g1661)) + ((!g182) & (g239) & (!g247) & (!g1163) & (!g1660) & (!g1661)) + ((!g182) & (g239) & (!g247) & (!g1163) & (g1660) & (!g1661)) + ((!g182) & (g239) & (!g247) & (g1163) & (g1660) & (!g1661)) + ((!g182) & (g239) & (!g247) & (g1163) & (g1660) & (g1661)) + ((!g182) & (g239) & (g247) & (!g1163) & (!g1660) & (g1661)) + ((!g182) & (g239) & (g247) & (!g1163) & (g1660) & (g1661)) + ((!g182) & (g239) & (g247) & (g1163) & (!g1660) & (!g1661)) + ((!g182) & (g239) & (g247) & (g1163) & (!g1660) & (g1661)) + ((g182) & (!g239) & (!g247) & (!g1163) & (!g1660) & (!g1661)) + ((g182) & (!g239) & (!g247) & (!g1163) & (g1660) & (!g1661)) + ((g182) & (!g239) & (!g247) & (g1163) & (g1660) & (!g1661)) + ((g182) & (!g239) & (!g247) & (g1163) & (g1660) & (g1661)) + ((g182) & (!g239) & (g247) & (!g1163) & (!g1660) & (g1661)) + ((g182) & (!g239) & (g247) & (!g1163) & (g1660) & (g1661)) + ((g182) & (!g239) & (g247) & (g1163) & (!g1660) & (!g1661)) + ((g182) & (!g239) & (g247) & (g1163) & (!g1660) & (g1661)) + ((g182) & (g239) & (!g247) & (!g1163) & (!g1660) & (g1661)) + ((g182) & (g239) & (!g247) & (!g1163) & (g1660) & (g1661)) + ((g182) & (g239) & (!g247) & (g1163) & (g1660) & (!g1661)) + ((g182) & (g239) & (!g247) & (g1163) & (g1660) & (g1661)) + ((g182) & (g239) & (g247) & (!g1163) & (!g1660) & (!g1661)) + ((g182) & (g239) & (g247) & (!g1163) & (g1660) & (!g1661)) + ((g182) & (g239) & (g247) & (g1163) & (!g1660) & (!g1661)) + ((g182) & (g239) & (g247) & (g1163) & (!g1660) & (g1661)));
	assign g2160 = (((!ld) & (!sk[112]) & (text_inx12x) & (!g1663)) + ((!ld) & (!sk[112]) & (text_inx12x) & (g1663)) + ((!ld) & (sk[112]) & (!text_inx12x) & (g1663)) + ((!ld) & (sk[112]) & (text_inx12x) & (g1663)) + ((ld) & (!sk[112]) & (!text_inx12x) & (g1663)) + ((ld) & (!sk[112]) & (text_inx12x) & (!g1663)) + ((ld) & (!sk[112]) & (text_inx12x) & (g1663)) + ((ld) & (sk[112]) & (text_inx12x) & (!g1663)) + ((ld) & (sk[112]) & (text_inx12x) & (g1663)));
	assign g1664 = (((!g303) & (!sk[113]) & (g367)) + ((!g303) & (sk[113]) & (g367)) + ((g303) & (!sk[113]) & (g367)) + ((g303) & (sk[113]) & (!g367)));
	assign g1665 = (((!g168) & (!g175) & (!sk[114]) & (g232) & (!g240)) + ((!g168) & (!g175) & (!sk[114]) & (g232) & (g240)) + ((!g168) & (!g175) & (sk[114]) & (!g232) & (g240)) + ((!g168) & (!g175) & (sk[114]) & (g232) & (!g240)) + ((!g168) & (g175) & (!sk[114]) & (!g232) & (!g240)) + ((!g168) & (g175) & (!sk[114]) & (!g232) & (g240)) + ((!g168) & (g175) & (!sk[114]) & (g232) & (!g240)) + ((!g168) & (g175) & (!sk[114]) & (g232) & (g240)) + ((!g168) & (g175) & (sk[114]) & (!g232) & (!g240)) + ((!g168) & (g175) & (sk[114]) & (g232) & (g240)) + ((g168) & (!g175) & (!sk[114]) & (g232) & (!g240)) + ((g168) & (!g175) & (!sk[114]) & (g232) & (g240)) + ((g168) & (!g175) & (sk[114]) & (!g232) & (!g240)) + ((g168) & (!g175) & (sk[114]) & (g232) & (g240)) + ((g168) & (g175) & (!sk[114]) & (!g232) & (!g240)) + ((g168) & (g175) & (!sk[114]) & (!g232) & (g240)) + ((g168) & (g175) & (!sk[114]) & (g232) & (!g240)) + ((g168) & (g175) & (!sk[114]) & (g232) & (g240)) + ((g168) & (g175) & (sk[114]) & (!g232) & (g240)) + ((g168) & (g175) & (sk[114]) & (g232) & (!g240)));
	assign g1666 = (((!g240) & (!g1163) & (!g1431) & (!g1663) & (!g1664) & (g1665)) + ((!g240) & (!g1163) & (!g1431) & (!g1663) & (g1664) & (!g1665)) + ((!g240) & (!g1163) & (!g1431) & (g1663) & (!g1664) & (g1665)) + ((!g240) & (!g1163) & (!g1431) & (g1663) & (g1664) & (!g1665)) + ((!g240) & (!g1163) & (g1431) & (!g1663) & (!g1664) & (!g1665)) + ((!g240) & (!g1163) & (g1431) & (!g1663) & (g1664) & (g1665)) + ((!g240) & (!g1163) & (g1431) & (g1663) & (!g1664) & (!g1665)) + ((!g240) & (!g1163) & (g1431) & (g1663) & (g1664) & (g1665)) + ((!g240) & (g1163) & (!g1431) & (g1663) & (!g1664) & (!g1665)) + ((!g240) & (g1163) & (!g1431) & (g1663) & (!g1664) & (g1665)) + ((!g240) & (g1163) & (!g1431) & (g1663) & (g1664) & (!g1665)) + ((!g240) & (g1163) & (!g1431) & (g1663) & (g1664) & (g1665)) + ((!g240) & (g1163) & (g1431) & (g1663) & (!g1664) & (!g1665)) + ((!g240) & (g1163) & (g1431) & (g1663) & (!g1664) & (g1665)) + ((!g240) & (g1163) & (g1431) & (g1663) & (g1664) & (!g1665)) + ((!g240) & (g1163) & (g1431) & (g1663) & (g1664) & (g1665)) + ((g240) & (!g1163) & (!g1431) & (!g1663) & (!g1664) & (g1665)) + ((g240) & (!g1163) & (!g1431) & (!g1663) & (g1664) & (!g1665)) + ((g240) & (!g1163) & (!g1431) & (g1663) & (!g1664) & (g1665)) + ((g240) & (!g1163) & (!g1431) & (g1663) & (g1664) & (!g1665)) + ((g240) & (!g1163) & (g1431) & (!g1663) & (!g1664) & (!g1665)) + ((g240) & (!g1163) & (g1431) & (!g1663) & (g1664) & (g1665)) + ((g240) & (!g1163) & (g1431) & (g1663) & (!g1664) & (!g1665)) + ((g240) & (!g1163) & (g1431) & (g1663) & (g1664) & (g1665)) + ((g240) & (g1163) & (!g1431) & (!g1663) & (!g1664) & (!g1665)) + ((g240) & (g1163) & (!g1431) & (!g1663) & (!g1664) & (g1665)) + ((g240) & (g1163) & (!g1431) & (!g1663) & (g1664) & (!g1665)) + ((g240) & (g1163) & (!g1431) & (!g1663) & (g1664) & (g1665)) + ((g240) & (g1163) & (g1431) & (!g1663) & (!g1664) & (!g1665)) + ((g240) & (g1163) & (g1431) & (!g1663) & (!g1664) & (g1665)) + ((g240) & (g1163) & (g1431) & (!g1663) & (g1664) & (!g1665)) + ((g240) & (g1163) & (g1431) & (!g1663) & (g1664) & (g1665)));
	assign g2161 = (((!sk[116]) & (!ld) & (text_inx15x) & (!g1667)) + ((!sk[116]) & (!ld) & (text_inx15x) & (g1667)) + ((!sk[116]) & (ld) & (!text_inx15x) & (g1667)) + ((!sk[116]) & (ld) & (text_inx15x) & (!g1667)) + ((!sk[116]) & (ld) & (text_inx15x) & (g1667)) + ((sk[116]) & (!ld) & (!text_inx15x) & (g1667)) + ((sk[116]) & (!ld) & (text_inx15x) & (g1667)) + ((sk[116]) & (ld) & (text_inx15x) & (!g1667)) + ((sk[116]) & (ld) & (text_inx15x) & (g1667)));
	assign g1668 = (((!g196) & (!sk[117]) & (!g261) & (g324) & (!g388)) + ((!g196) & (!sk[117]) & (!g261) & (g324) & (g388)) + ((!g196) & (!sk[117]) & (g261) & (!g324) & (!g388)) + ((!g196) & (!sk[117]) & (g261) & (!g324) & (g388)) + ((!g196) & (!sk[117]) & (g261) & (g324) & (!g388)) + ((!g196) & (!sk[117]) & (g261) & (g324) & (g388)) + ((!g196) & (sk[117]) & (!g261) & (!g324) & (g388)) + ((!g196) & (sk[117]) & (!g261) & (g324) & (!g388)) + ((!g196) & (sk[117]) & (g261) & (!g324) & (!g388)) + ((!g196) & (sk[117]) & (g261) & (g324) & (g388)) + ((g196) & (!sk[117]) & (!g261) & (g324) & (!g388)) + ((g196) & (!sk[117]) & (!g261) & (g324) & (g388)) + ((g196) & (!sk[117]) & (g261) & (!g324) & (!g388)) + ((g196) & (!sk[117]) & (g261) & (!g324) & (g388)) + ((g196) & (!sk[117]) & (g261) & (g324) & (!g388)) + ((g196) & (!sk[117]) & (g261) & (g324) & (g388)) + ((g196) & (sk[117]) & (!g261) & (!g324) & (!g388)) + ((g196) & (sk[117]) & (!g261) & (g324) & (g388)) + ((g196) & (sk[117]) & (g261) & (!g324) & (g388)) + ((g196) & (sk[117]) & (g261) & (g324) & (!g388)));
	assign g1669 = (((!g189) & (!g253) & (!g261) & (!g1163) & (!g1667) & (g1668)) + ((!g189) & (!g253) & (!g261) & (!g1163) & (g1667) & (g1668)) + ((!g189) & (!g253) & (!g261) & (g1163) & (g1667) & (!g1668)) + ((!g189) & (!g253) & (!g261) & (g1163) & (g1667) & (g1668)) + ((!g189) & (!g253) & (g261) & (!g1163) & (!g1667) & (g1668)) + ((!g189) & (!g253) & (g261) & (!g1163) & (g1667) & (g1668)) + ((!g189) & (!g253) & (g261) & (g1163) & (!g1667) & (!g1668)) + ((!g189) & (!g253) & (g261) & (g1163) & (!g1667) & (g1668)) + ((!g189) & (g253) & (!g261) & (!g1163) & (!g1667) & (!g1668)) + ((!g189) & (g253) & (!g261) & (!g1163) & (g1667) & (!g1668)) + ((!g189) & (g253) & (!g261) & (g1163) & (g1667) & (!g1668)) + ((!g189) & (g253) & (!g261) & (g1163) & (g1667) & (g1668)) + ((!g189) & (g253) & (g261) & (!g1163) & (!g1667) & (!g1668)) + ((!g189) & (g253) & (g261) & (!g1163) & (g1667) & (!g1668)) + ((!g189) & (g253) & (g261) & (g1163) & (!g1667) & (!g1668)) + ((!g189) & (g253) & (g261) & (g1163) & (!g1667) & (g1668)) + ((g189) & (!g253) & (!g261) & (!g1163) & (!g1667) & (!g1668)) + ((g189) & (!g253) & (!g261) & (!g1163) & (g1667) & (!g1668)) + ((g189) & (!g253) & (!g261) & (g1163) & (g1667) & (!g1668)) + ((g189) & (!g253) & (!g261) & (g1163) & (g1667) & (g1668)) + ((g189) & (!g253) & (g261) & (!g1163) & (!g1667) & (!g1668)) + ((g189) & (!g253) & (g261) & (!g1163) & (g1667) & (!g1668)) + ((g189) & (!g253) & (g261) & (g1163) & (!g1667) & (!g1668)) + ((g189) & (!g253) & (g261) & (g1163) & (!g1667) & (g1668)) + ((g189) & (g253) & (!g261) & (!g1163) & (!g1667) & (g1668)) + ((g189) & (g253) & (!g261) & (!g1163) & (g1667) & (g1668)) + ((g189) & (g253) & (!g261) & (g1163) & (g1667) & (!g1668)) + ((g189) & (g253) & (!g261) & (g1163) & (g1667) & (g1668)) + ((g189) & (g253) & (g261) & (!g1163) & (!g1667) & (g1668)) + ((g189) & (g253) & (g261) & (!g1163) & (g1667) & (g1668)) + ((g189) & (g253) & (g261) & (g1163) & (!g1667) & (!g1668)) + ((g189) & (g253) & (g261) & (g1163) & (!g1667) & (g1668)));
	assign g1670 = (((!ld) & (!g724) & (!g980) & (sk[119]) & (g1276) & (!keyx72x)) + ((!ld) & (!g724) & (!g980) & (sk[119]) & (g1276) & (keyx72x)) + ((!ld) & (!g724) & (g980) & (sk[119]) & (!g1276) & (!keyx72x)) + ((!ld) & (!g724) & (g980) & (sk[119]) & (!g1276) & (keyx72x)) + ((!ld) & (g724) & (!g980) & (!sk[119]) & (!g1276) & (!keyx72x)) + ((!ld) & (g724) & (!g980) & (!sk[119]) & (!g1276) & (keyx72x)) + ((!ld) & (g724) & (!g980) & (!sk[119]) & (g1276) & (!keyx72x)) + ((!ld) & (g724) & (!g980) & (!sk[119]) & (g1276) & (keyx72x)) + ((!ld) & (g724) & (!g980) & (sk[119]) & (!g1276) & (!keyx72x)) + ((!ld) & (g724) & (!g980) & (sk[119]) & (!g1276) & (keyx72x)) + ((!ld) & (g724) & (g980) & (!sk[119]) & (!g1276) & (!keyx72x)) + ((!ld) & (g724) & (g980) & (!sk[119]) & (!g1276) & (keyx72x)) + ((!ld) & (g724) & (g980) & (!sk[119]) & (g1276) & (!keyx72x)) + ((!ld) & (g724) & (g980) & (!sk[119]) & (g1276) & (keyx72x)) + ((!ld) & (g724) & (g980) & (sk[119]) & (g1276) & (!keyx72x)) + ((!ld) & (g724) & (g980) & (sk[119]) & (g1276) & (keyx72x)) + ((ld) & (!g724) & (!g980) & (!sk[119]) & (!g1276) & (!keyx72x)) + ((ld) & (!g724) & (!g980) & (!sk[119]) & (!g1276) & (keyx72x)) + ((ld) & (!g724) & (!g980) & (!sk[119]) & (g1276) & (!keyx72x)) + ((ld) & (!g724) & (!g980) & (!sk[119]) & (g1276) & (keyx72x)) + ((ld) & (!g724) & (!g980) & (sk[119]) & (!g1276) & (keyx72x)) + ((ld) & (!g724) & (!g980) & (sk[119]) & (g1276) & (keyx72x)) + ((ld) & (!g724) & (g980) & (!sk[119]) & (!g1276) & (!keyx72x)) + ((ld) & (!g724) & (g980) & (!sk[119]) & (!g1276) & (keyx72x)) + ((ld) & (!g724) & (g980) & (!sk[119]) & (g1276) & (!keyx72x)) + ((ld) & (!g724) & (g980) & (!sk[119]) & (g1276) & (keyx72x)) + ((ld) & (!g724) & (g980) & (sk[119]) & (!g1276) & (keyx72x)) + ((ld) & (!g724) & (g980) & (sk[119]) & (g1276) & (keyx72x)) + ((ld) & (g724) & (!g980) & (!sk[119]) & (!g1276) & (!keyx72x)) + ((ld) & (g724) & (!g980) & (!sk[119]) & (!g1276) & (keyx72x)) + ((ld) & (g724) & (!g980) & (!sk[119]) & (g1276) & (!keyx72x)) + ((ld) & (g724) & (!g980) & (!sk[119]) & (g1276) & (keyx72x)) + ((ld) & (g724) & (!g980) & (sk[119]) & (!g1276) & (keyx72x)) + ((ld) & (g724) & (!g980) & (sk[119]) & (g1276) & (keyx72x)) + ((ld) & (g724) & (g980) & (!sk[119]) & (!g1276) & (!keyx72x)) + ((ld) & (g724) & (g980) & (!sk[119]) & (!g1276) & (keyx72x)) + ((ld) & (g724) & (g980) & (!sk[119]) & (g1276) & (!keyx72x)) + ((ld) & (g724) & (g980) & (!sk[119]) & (g1276) & (keyx72x)) + ((ld) & (g724) & (g980) & (sk[119]) & (!g1276) & (keyx72x)) + ((ld) & (g724) & (g980) & (sk[119]) & (g1276) & (keyx72x)));
	assign g1671 = (((!ld) & (!g731) & (!g987) & (g1283) & (sk[120]) & (!keyx73x)) + ((!ld) & (!g731) & (!g987) & (g1283) & (sk[120]) & (keyx73x)) + ((!ld) & (!g731) & (g987) & (!g1283) & (sk[120]) & (!keyx73x)) + ((!ld) & (!g731) & (g987) & (!g1283) & (sk[120]) & (keyx73x)) + ((!ld) & (g731) & (!g987) & (!g1283) & (!sk[120]) & (!keyx73x)) + ((!ld) & (g731) & (!g987) & (!g1283) & (!sk[120]) & (keyx73x)) + ((!ld) & (g731) & (!g987) & (!g1283) & (sk[120]) & (!keyx73x)) + ((!ld) & (g731) & (!g987) & (!g1283) & (sk[120]) & (keyx73x)) + ((!ld) & (g731) & (!g987) & (g1283) & (!sk[120]) & (!keyx73x)) + ((!ld) & (g731) & (!g987) & (g1283) & (!sk[120]) & (keyx73x)) + ((!ld) & (g731) & (g987) & (!g1283) & (!sk[120]) & (!keyx73x)) + ((!ld) & (g731) & (g987) & (!g1283) & (!sk[120]) & (keyx73x)) + ((!ld) & (g731) & (g987) & (g1283) & (!sk[120]) & (!keyx73x)) + ((!ld) & (g731) & (g987) & (g1283) & (!sk[120]) & (keyx73x)) + ((!ld) & (g731) & (g987) & (g1283) & (sk[120]) & (!keyx73x)) + ((!ld) & (g731) & (g987) & (g1283) & (sk[120]) & (keyx73x)) + ((ld) & (!g731) & (!g987) & (!g1283) & (!sk[120]) & (!keyx73x)) + ((ld) & (!g731) & (!g987) & (!g1283) & (!sk[120]) & (keyx73x)) + ((ld) & (!g731) & (!g987) & (!g1283) & (sk[120]) & (keyx73x)) + ((ld) & (!g731) & (!g987) & (g1283) & (!sk[120]) & (!keyx73x)) + ((ld) & (!g731) & (!g987) & (g1283) & (!sk[120]) & (keyx73x)) + ((ld) & (!g731) & (!g987) & (g1283) & (sk[120]) & (keyx73x)) + ((ld) & (!g731) & (g987) & (!g1283) & (!sk[120]) & (!keyx73x)) + ((ld) & (!g731) & (g987) & (!g1283) & (!sk[120]) & (keyx73x)) + ((ld) & (!g731) & (g987) & (!g1283) & (sk[120]) & (keyx73x)) + ((ld) & (!g731) & (g987) & (g1283) & (!sk[120]) & (!keyx73x)) + ((ld) & (!g731) & (g987) & (g1283) & (!sk[120]) & (keyx73x)) + ((ld) & (!g731) & (g987) & (g1283) & (sk[120]) & (keyx73x)) + ((ld) & (g731) & (!g987) & (!g1283) & (!sk[120]) & (!keyx73x)) + ((ld) & (g731) & (!g987) & (!g1283) & (!sk[120]) & (keyx73x)) + ((ld) & (g731) & (!g987) & (!g1283) & (sk[120]) & (keyx73x)) + ((ld) & (g731) & (!g987) & (g1283) & (!sk[120]) & (!keyx73x)) + ((ld) & (g731) & (!g987) & (g1283) & (!sk[120]) & (keyx73x)) + ((ld) & (g731) & (!g987) & (g1283) & (sk[120]) & (keyx73x)) + ((ld) & (g731) & (g987) & (!g1283) & (!sk[120]) & (!keyx73x)) + ((ld) & (g731) & (g987) & (!g1283) & (!sk[120]) & (keyx73x)) + ((ld) & (g731) & (g987) & (!g1283) & (sk[120]) & (keyx73x)) + ((ld) & (g731) & (g987) & (g1283) & (!sk[120]) & (!keyx73x)) + ((ld) & (g731) & (g987) & (g1283) & (!sk[120]) & (keyx73x)) + ((ld) & (g731) & (g987) & (g1283) & (sk[120]) & (keyx73x)));
	assign g1672 = (((!ld) & (!g738) & (!g994) & (g1290) & (sk[121]) & (!keyx74x)) + ((!ld) & (!g738) & (!g994) & (g1290) & (sk[121]) & (keyx74x)) + ((!ld) & (!g738) & (g994) & (!g1290) & (sk[121]) & (!keyx74x)) + ((!ld) & (!g738) & (g994) & (!g1290) & (sk[121]) & (keyx74x)) + ((!ld) & (g738) & (!g994) & (!g1290) & (!sk[121]) & (!keyx74x)) + ((!ld) & (g738) & (!g994) & (!g1290) & (!sk[121]) & (keyx74x)) + ((!ld) & (g738) & (!g994) & (!g1290) & (sk[121]) & (!keyx74x)) + ((!ld) & (g738) & (!g994) & (!g1290) & (sk[121]) & (keyx74x)) + ((!ld) & (g738) & (!g994) & (g1290) & (!sk[121]) & (!keyx74x)) + ((!ld) & (g738) & (!g994) & (g1290) & (!sk[121]) & (keyx74x)) + ((!ld) & (g738) & (g994) & (!g1290) & (!sk[121]) & (!keyx74x)) + ((!ld) & (g738) & (g994) & (!g1290) & (!sk[121]) & (keyx74x)) + ((!ld) & (g738) & (g994) & (g1290) & (!sk[121]) & (!keyx74x)) + ((!ld) & (g738) & (g994) & (g1290) & (!sk[121]) & (keyx74x)) + ((!ld) & (g738) & (g994) & (g1290) & (sk[121]) & (!keyx74x)) + ((!ld) & (g738) & (g994) & (g1290) & (sk[121]) & (keyx74x)) + ((ld) & (!g738) & (!g994) & (!g1290) & (!sk[121]) & (!keyx74x)) + ((ld) & (!g738) & (!g994) & (!g1290) & (!sk[121]) & (keyx74x)) + ((ld) & (!g738) & (!g994) & (!g1290) & (sk[121]) & (keyx74x)) + ((ld) & (!g738) & (!g994) & (g1290) & (!sk[121]) & (!keyx74x)) + ((ld) & (!g738) & (!g994) & (g1290) & (!sk[121]) & (keyx74x)) + ((ld) & (!g738) & (!g994) & (g1290) & (sk[121]) & (keyx74x)) + ((ld) & (!g738) & (g994) & (!g1290) & (!sk[121]) & (!keyx74x)) + ((ld) & (!g738) & (g994) & (!g1290) & (!sk[121]) & (keyx74x)) + ((ld) & (!g738) & (g994) & (!g1290) & (sk[121]) & (keyx74x)) + ((ld) & (!g738) & (g994) & (g1290) & (!sk[121]) & (!keyx74x)) + ((ld) & (!g738) & (g994) & (g1290) & (!sk[121]) & (keyx74x)) + ((ld) & (!g738) & (g994) & (g1290) & (sk[121]) & (keyx74x)) + ((ld) & (g738) & (!g994) & (!g1290) & (!sk[121]) & (!keyx74x)) + ((ld) & (g738) & (!g994) & (!g1290) & (!sk[121]) & (keyx74x)) + ((ld) & (g738) & (!g994) & (!g1290) & (sk[121]) & (keyx74x)) + ((ld) & (g738) & (!g994) & (g1290) & (!sk[121]) & (!keyx74x)) + ((ld) & (g738) & (!g994) & (g1290) & (!sk[121]) & (keyx74x)) + ((ld) & (g738) & (!g994) & (g1290) & (sk[121]) & (keyx74x)) + ((ld) & (g738) & (g994) & (!g1290) & (!sk[121]) & (!keyx74x)) + ((ld) & (g738) & (g994) & (!g1290) & (!sk[121]) & (keyx74x)) + ((ld) & (g738) & (g994) & (!g1290) & (sk[121]) & (keyx74x)) + ((ld) & (g738) & (g994) & (g1290) & (!sk[121]) & (!keyx74x)) + ((ld) & (g738) & (g994) & (g1290) & (!sk[121]) & (keyx74x)) + ((ld) & (g738) & (g994) & (g1290) & (sk[121]) & (keyx74x)));
	assign g1673 = (((!ld) & (!g745) & (!g1001) & (sk[122]) & (g1297) & (!keyx75x)) + ((!ld) & (!g745) & (!g1001) & (sk[122]) & (g1297) & (keyx75x)) + ((!ld) & (!g745) & (g1001) & (sk[122]) & (!g1297) & (!keyx75x)) + ((!ld) & (!g745) & (g1001) & (sk[122]) & (!g1297) & (keyx75x)) + ((!ld) & (g745) & (!g1001) & (!sk[122]) & (!g1297) & (!keyx75x)) + ((!ld) & (g745) & (!g1001) & (!sk[122]) & (!g1297) & (keyx75x)) + ((!ld) & (g745) & (!g1001) & (!sk[122]) & (g1297) & (!keyx75x)) + ((!ld) & (g745) & (!g1001) & (!sk[122]) & (g1297) & (keyx75x)) + ((!ld) & (g745) & (!g1001) & (sk[122]) & (!g1297) & (!keyx75x)) + ((!ld) & (g745) & (!g1001) & (sk[122]) & (!g1297) & (keyx75x)) + ((!ld) & (g745) & (g1001) & (!sk[122]) & (!g1297) & (!keyx75x)) + ((!ld) & (g745) & (g1001) & (!sk[122]) & (!g1297) & (keyx75x)) + ((!ld) & (g745) & (g1001) & (!sk[122]) & (g1297) & (!keyx75x)) + ((!ld) & (g745) & (g1001) & (!sk[122]) & (g1297) & (keyx75x)) + ((!ld) & (g745) & (g1001) & (sk[122]) & (g1297) & (!keyx75x)) + ((!ld) & (g745) & (g1001) & (sk[122]) & (g1297) & (keyx75x)) + ((ld) & (!g745) & (!g1001) & (!sk[122]) & (!g1297) & (!keyx75x)) + ((ld) & (!g745) & (!g1001) & (!sk[122]) & (!g1297) & (keyx75x)) + ((ld) & (!g745) & (!g1001) & (!sk[122]) & (g1297) & (!keyx75x)) + ((ld) & (!g745) & (!g1001) & (!sk[122]) & (g1297) & (keyx75x)) + ((ld) & (!g745) & (!g1001) & (sk[122]) & (!g1297) & (keyx75x)) + ((ld) & (!g745) & (!g1001) & (sk[122]) & (g1297) & (keyx75x)) + ((ld) & (!g745) & (g1001) & (!sk[122]) & (!g1297) & (!keyx75x)) + ((ld) & (!g745) & (g1001) & (!sk[122]) & (!g1297) & (keyx75x)) + ((ld) & (!g745) & (g1001) & (!sk[122]) & (g1297) & (!keyx75x)) + ((ld) & (!g745) & (g1001) & (!sk[122]) & (g1297) & (keyx75x)) + ((ld) & (!g745) & (g1001) & (sk[122]) & (!g1297) & (keyx75x)) + ((ld) & (!g745) & (g1001) & (sk[122]) & (g1297) & (keyx75x)) + ((ld) & (g745) & (!g1001) & (!sk[122]) & (!g1297) & (!keyx75x)) + ((ld) & (g745) & (!g1001) & (!sk[122]) & (!g1297) & (keyx75x)) + ((ld) & (g745) & (!g1001) & (!sk[122]) & (g1297) & (!keyx75x)) + ((ld) & (g745) & (!g1001) & (!sk[122]) & (g1297) & (keyx75x)) + ((ld) & (g745) & (!g1001) & (sk[122]) & (!g1297) & (keyx75x)) + ((ld) & (g745) & (!g1001) & (sk[122]) & (g1297) & (keyx75x)) + ((ld) & (g745) & (g1001) & (!sk[122]) & (!g1297) & (!keyx75x)) + ((ld) & (g745) & (g1001) & (!sk[122]) & (!g1297) & (keyx75x)) + ((ld) & (g745) & (g1001) & (!sk[122]) & (g1297) & (!keyx75x)) + ((ld) & (g745) & (g1001) & (!sk[122]) & (g1297) & (keyx75x)) + ((ld) & (g745) & (g1001) & (sk[122]) & (!g1297) & (keyx75x)) + ((ld) & (g745) & (g1001) & (sk[122]) & (g1297) & (keyx75x)));
	assign g1674 = (((!sk[123]) & (!ld) & (g752) & (!g1008) & (!g1304) & (!keyx76x)) + ((!sk[123]) & (!ld) & (g752) & (!g1008) & (!g1304) & (keyx76x)) + ((!sk[123]) & (!ld) & (g752) & (!g1008) & (g1304) & (!keyx76x)) + ((!sk[123]) & (!ld) & (g752) & (!g1008) & (g1304) & (keyx76x)) + ((!sk[123]) & (!ld) & (g752) & (g1008) & (!g1304) & (!keyx76x)) + ((!sk[123]) & (!ld) & (g752) & (g1008) & (!g1304) & (keyx76x)) + ((!sk[123]) & (!ld) & (g752) & (g1008) & (g1304) & (!keyx76x)) + ((!sk[123]) & (!ld) & (g752) & (g1008) & (g1304) & (keyx76x)) + ((!sk[123]) & (ld) & (!g752) & (!g1008) & (!g1304) & (!keyx76x)) + ((!sk[123]) & (ld) & (!g752) & (!g1008) & (!g1304) & (keyx76x)) + ((!sk[123]) & (ld) & (!g752) & (!g1008) & (g1304) & (!keyx76x)) + ((!sk[123]) & (ld) & (!g752) & (!g1008) & (g1304) & (keyx76x)) + ((!sk[123]) & (ld) & (!g752) & (g1008) & (!g1304) & (!keyx76x)) + ((!sk[123]) & (ld) & (!g752) & (g1008) & (!g1304) & (keyx76x)) + ((!sk[123]) & (ld) & (!g752) & (g1008) & (g1304) & (!keyx76x)) + ((!sk[123]) & (ld) & (!g752) & (g1008) & (g1304) & (keyx76x)) + ((!sk[123]) & (ld) & (g752) & (!g1008) & (!g1304) & (!keyx76x)) + ((!sk[123]) & (ld) & (g752) & (!g1008) & (!g1304) & (keyx76x)) + ((!sk[123]) & (ld) & (g752) & (!g1008) & (g1304) & (!keyx76x)) + ((!sk[123]) & (ld) & (g752) & (!g1008) & (g1304) & (keyx76x)) + ((!sk[123]) & (ld) & (g752) & (g1008) & (!g1304) & (!keyx76x)) + ((!sk[123]) & (ld) & (g752) & (g1008) & (!g1304) & (keyx76x)) + ((!sk[123]) & (ld) & (g752) & (g1008) & (g1304) & (!keyx76x)) + ((!sk[123]) & (ld) & (g752) & (g1008) & (g1304) & (keyx76x)) + ((sk[123]) & (!ld) & (!g752) & (!g1008) & (g1304) & (!keyx76x)) + ((sk[123]) & (!ld) & (!g752) & (!g1008) & (g1304) & (keyx76x)) + ((sk[123]) & (!ld) & (!g752) & (g1008) & (!g1304) & (!keyx76x)) + ((sk[123]) & (!ld) & (!g752) & (g1008) & (!g1304) & (keyx76x)) + ((sk[123]) & (!ld) & (g752) & (!g1008) & (!g1304) & (!keyx76x)) + ((sk[123]) & (!ld) & (g752) & (!g1008) & (!g1304) & (keyx76x)) + ((sk[123]) & (!ld) & (g752) & (g1008) & (g1304) & (!keyx76x)) + ((sk[123]) & (!ld) & (g752) & (g1008) & (g1304) & (keyx76x)) + ((sk[123]) & (ld) & (!g752) & (!g1008) & (!g1304) & (keyx76x)) + ((sk[123]) & (ld) & (!g752) & (!g1008) & (g1304) & (keyx76x)) + ((sk[123]) & (ld) & (!g752) & (g1008) & (!g1304) & (keyx76x)) + ((sk[123]) & (ld) & (!g752) & (g1008) & (g1304) & (keyx76x)) + ((sk[123]) & (ld) & (g752) & (!g1008) & (!g1304) & (keyx76x)) + ((sk[123]) & (ld) & (g752) & (!g1008) & (g1304) & (keyx76x)) + ((sk[123]) & (ld) & (g752) & (g1008) & (!g1304) & (keyx76x)) + ((sk[123]) & (ld) & (g752) & (g1008) & (g1304) & (keyx76x)));
	assign g1675 = (((!ld) & (!g759) & (!g1015) & (g1311) & (sk[124]) & (!keyx77x)) + ((!ld) & (!g759) & (!g1015) & (g1311) & (sk[124]) & (keyx77x)) + ((!ld) & (!g759) & (g1015) & (!g1311) & (sk[124]) & (!keyx77x)) + ((!ld) & (!g759) & (g1015) & (!g1311) & (sk[124]) & (keyx77x)) + ((!ld) & (g759) & (!g1015) & (!g1311) & (!sk[124]) & (!keyx77x)) + ((!ld) & (g759) & (!g1015) & (!g1311) & (!sk[124]) & (keyx77x)) + ((!ld) & (g759) & (!g1015) & (!g1311) & (sk[124]) & (!keyx77x)) + ((!ld) & (g759) & (!g1015) & (!g1311) & (sk[124]) & (keyx77x)) + ((!ld) & (g759) & (!g1015) & (g1311) & (!sk[124]) & (!keyx77x)) + ((!ld) & (g759) & (!g1015) & (g1311) & (!sk[124]) & (keyx77x)) + ((!ld) & (g759) & (g1015) & (!g1311) & (!sk[124]) & (!keyx77x)) + ((!ld) & (g759) & (g1015) & (!g1311) & (!sk[124]) & (keyx77x)) + ((!ld) & (g759) & (g1015) & (g1311) & (!sk[124]) & (!keyx77x)) + ((!ld) & (g759) & (g1015) & (g1311) & (!sk[124]) & (keyx77x)) + ((!ld) & (g759) & (g1015) & (g1311) & (sk[124]) & (!keyx77x)) + ((!ld) & (g759) & (g1015) & (g1311) & (sk[124]) & (keyx77x)) + ((ld) & (!g759) & (!g1015) & (!g1311) & (!sk[124]) & (!keyx77x)) + ((ld) & (!g759) & (!g1015) & (!g1311) & (!sk[124]) & (keyx77x)) + ((ld) & (!g759) & (!g1015) & (!g1311) & (sk[124]) & (keyx77x)) + ((ld) & (!g759) & (!g1015) & (g1311) & (!sk[124]) & (!keyx77x)) + ((ld) & (!g759) & (!g1015) & (g1311) & (!sk[124]) & (keyx77x)) + ((ld) & (!g759) & (!g1015) & (g1311) & (sk[124]) & (keyx77x)) + ((ld) & (!g759) & (g1015) & (!g1311) & (!sk[124]) & (!keyx77x)) + ((ld) & (!g759) & (g1015) & (!g1311) & (!sk[124]) & (keyx77x)) + ((ld) & (!g759) & (g1015) & (!g1311) & (sk[124]) & (keyx77x)) + ((ld) & (!g759) & (g1015) & (g1311) & (!sk[124]) & (!keyx77x)) + ((ld) & (!g759) & (g1015) & (g1311) & (!sk[124]) & (keyx77x)) + ((ld) & (!g759) & (g1015) & (g1311) & (sk[124]) & (keyx77x)) + ((ld) & (g759) & (!g1015) & (!g1311) & (!sk[124]) & (!keyx77x)) + ((ld) & (g759) & (!g1015) & (!g1311) & (!sk[124]) & (keyx77x)) + ((ld) & (g759) & (!g1015) & (!g1311) & (sk[124]) & (keyx77x)) + ((ld) & (g759) & (!g1015) & (g1311) & (!sk[124]) & (!keyx77x)) + ((ld) & (g759) & (!g1015) & (g1311) & (!sk[124]) & (keyx77x)) + ((ld) & (g759) & (!g1015) & (g1311) & (sk[124]) & (keyx77x)) + ((ld) & (g759) & (g1015) & (!g1311) & (!sk[124]) & (!keyx77x)) + ((ld) & (g759) & (g1015) & (!g1311) & (!sk[124]) & (keyx77x)) + ((ld) & (g759) & (g1015) & (!g1311) & (sk[124]) & (keyx77x)) + ((ld) & (g759) & (g1015) & (g1311) & (!sk[124]) & (!keyx77x)) + ((ld) & (g759) & (g1015) & (g1311) & (!sk[124]) & (keyx77x)) + ((ld) & (g759) & (g1015) & (g1311) & (sk[124]) & (keyx77x)));
	assign g1676 = (((!ld) & (!g766) & (sk[125]) & (!g1022) & (g1318) & (!keyx78x)) + ((!ld) & (!g766) & (sk[125]) & (!g1022) & (g1318) & (keyx78x)) + ((!ld) & (!g766) & (sk[125]) & (g1022) & (!g1318) & (!keyx78x)) + ((!ld) & (!g766) & (sk[125]) & (g1022) & (!g1318) & (keyx78x)) + ((!ld) & (g766) & (!sk[125]) & (!g1022) & (!g1318) & (!keyx78x)) + ((!ld) & (g766) & (!sk[125]) & (!g1022) & (!g1318) & (keyx78x)) + ((!ld) & (g766) & (!sk[125]) & (!g1022) & (g1318) & (!keyx78x)) + ((!ld) & (g766) & (!sk[125]) & (!g1022) & (g1318) & (keyx78x)) + ((!ld) & (g766) & (!sk[125]) & (g1022) & (!g1318) & (!keyx78x)) + ((!ld) & (g766) & (!sk[125]) & (g1022) & (!g1318) & (keyx78x)) + ((!ld) & (g766) & (!sk[125]) & (g1022) & (g1318) & (!keyx78x)) + ((!ld) & (g766) & (!sk[125]) & (g1022) & (g1318) & (keyx78x)) + ((!ld) & (g766) & (sk[125]) & (!g1022) & (!g1318) & (!keyx78x)) + ((!ld) & (g766) & (sk[125]) & (!g1022) & (!g1318) & (keyx78x)) + ((!ld) & (g766) & (sk[125]) & (g1022) & (g1318) & (!keyx78x)) + ((!ld) & (g766) & (sk[125]) & (g1022) & (g1318) & (keyx78x)) + ((ld) & (!g766) & (!sk[125]) & (!g1022) & (!g1318) & (!keyx78x)) + ((ld) & (!g766) & (!sk[125]) & (!g1022) & (!g1318) & (keyx78x)) + ((ld) & (!g766) & (!sk[125]) & (!g1022) & (g1318) & (!keyx78x)) + ((ld) & (!g766) & (!sk[125]) & (!g1022) & (g1318) & (keyx78x)) + ((ld) & (!g766) & (!sk[125]) & (g1022) & (!g1318) & (!keyx78x)) + ((ld) & (!g766) & (!sk[125]) & (g1022) & (!g1318) & (keyx78x)) + ((ld) & (!g766) & (!sk[125]) & (g1022) & (g1318) & (!keyx78x)) + ((ld) & (!g766) & (!sk[125]) & (g1022) & (g1318) & (keyx78x)) + ((ld) & (!g766) & (sk[125]) & (!g1022) & (!g1318) & (keyx78x)) + ((ld) & (!g766) & (sk[125]) & (!g1022) & (g1318) & (keyx78x)) + ((ld) & (!g766) & (sk[125]) & (g1022) & (!g1318) & (keyx78x)) + ((ld) & (!g766) & (sk[125]) & (g1022) & (g1318) & (keyx78x)) + ((ld) & (g766) & (!sk[125]) & (!g1022) & (!g1318) & (!keyx78x)) + ((ld) & (g766) & (!sk[125]) & (!g1022) & (!g1318) & (keyx78x)) + ((ld) & (g766) & (!sk[125]) & (!g1022) & (g1318) & (!keyx78x)) + ((ld) & (g766) & (!sk[125]) & (!g1022) & (g1318) & (keyx78x)) + ((ld) & (g766) & (!sk[125]) & (g1022) & (!g1318) & (!keyx78x)) + ((ld) & (g766) & (!sk[125]) & (g1022) & (!g1318) & (keyx78x)) + ((ld) & (g766) & (!sk[125]) & (g1022) & (g1318) & (!keyx78x)) + ((ld) & (g766) & (!sk[125]) & (g1022) & (g1318) & (keyx78x)) + ((ld) & (g766) & (sk[125]) & (!g1022) & (!g1318) & (keyx78x)) + ((ld) & (g766) & (sk[125]) & (!g1022) & (g1318) & (keyx78x)) + ((ld) & (g766) & (sk[125]) & (g1022) & (!g1318) & (keyx78x)) + ((ld) & (g766) & (sk[125]) & (g1022) & (g1318) & (keyx78x)));
	assign g1677 = (((!ld) & (!g773) & (sk[126]) & (!g1029) & (g1325) & (!keyx79x)) + ((!ld) & (!g773) & (sk[126]) & (!g1029) & (g1325) & (keyx79x)) + ((!ld) & (!g773) & (sk[126]) & (g1029) & (!g1325) & (!keyx79x)) + ((!ld) & (!g773) & (sk[126]) & (g1029) & (!g1325) & (keyx79x)) + ((!ld) & (g773) & (!sk[126]) & (!g1029) & (!g1325) & (!keyx79x)) + ((!ld) & (g773) & (!sk[126]) & (!g1029) & (!g1325) & (keyx79x)) + ((!ld) & (g773) & (!sk[126]) & (!g1029) & (g1325) & (!keyx79x)) + ((!ld) & (g773) & (!sk[126]) & (!g1029) & (g1325) & (keyx79x)) + ((!ld) & (g773) & (!sk[126]) & (g1029) & (!g1325) & (!keyx79x)) + ((!ld) & (g773) & (!sk[126]) & (g1029) & (!g1325) & (keyx79x)) + ((!ld) & (g773) & (!sk[126]) & (g1029) & (g1325) & (!keyx79x)) + ((!ld) & (g773) & (!sk[126]) & (g1029) & (g1325) & (keyx79x)) + ((!ld) & (g773) & (sk[126]) & (!g1029) & (!g1325) & (!keyx79x)) + ((!ld) & (g773) & (sk[126]) & (!g1029) & (!g1325) & (keyx79x)) + ((!ld) & (g773) & (sk[126]) & (g1029) & (g1325) & (!keyx79x)) + ((!ld) & (g773) & (sk[126]) & (g1029) & (g1325) & (keyx79x)) + ((ld) & (!g773) & (!sk[126]) & (!g1029) & (!g1325) & (!keyx79x)) + ((ld) & (!g773) & (!sk[126]) & (!g1029) & (!g1325) & (keyx79x)) + ((ld) & (!g773) & (!sk[126]) & (!g1029) & (g1325) & (!keyx79x)) + ((ld) & (!g773) & (!sk[126]) & (!g1029) & (g1325) & (keyx79x)) + ((ld) & (!g773) & (!sk[126]) & (g1029) & (!g1325) & (!keyx79x)) + ((ld) & (!g773) & (!sk[126]) & (g1029) & (!g1325) & (keyx79x)) + ((ld) & (!g773) & (!sk[126]) & (g1029) & (g1325) & (!keyx79x)) + ((ld) & (!g773) & (!sk[126]) & (g1029) & (g1325) & (keyx79x)) + ((ld) & (!g773) & (sk[126]) & (!g1029) & (!g1325) & (keyx79x)) + ((ld) & (!g773) & (sk[126]) & (!g1029) & (g1325) & (keyx79x)) + ((ld) & (!g773) & (sk[126]) & (g1029) & (!g1325) & (keyx79x)) + ((ld) & (!g773) & (sk[126]) & (g1029) & (g1325) & (keyx79x)) + ((ld) & (g773) & (!sk[126]) & (!g1029) & (!g1325) & (!keyx79x)) + ((ld) & (g773) & (!sk[126]) & (!g1029) & (!g1325) & (keyx79x)) + ((ld) & (g773) & (!sk[126]) & (!g1029) & (g1325) & (!keyx79x)) + ((ld) & (g773) & (!sk[126]) & (!g1029) & (g1325) & (keyx79x)) + ((ld) & (g773) & (!sk[126]) & (g1029) & (!g1325) & (!keyx79x)) + ((ld) & (g773) & (!sk[126]) & (g1029) & (!g1325) & (keyx79x)) + ((ld) & (g773) & (!sk[126]) & (g1029) & (g1325) & (!keyx79x)) + ((ld) & (g773) & (!sk[126]) & (g1029) & (g1325) & (keyx79x)) + ((ld) & (g773) & (sk[126]) & (!g1029) & (!g1325) & (keyx79x)) + ((ld) & (g773) & (sk[126]) & (!g1029) & (g1325) & (keyx79x)) + ((ld) & (g773) & (sk[126]) & (g1029) & (!g1325) & (keyx79x)) + ((ld) & (g773) & (sk[126]) & (g1029) & (g1325) & (keyx79x)));
	assign g2162 = (((!ld) & (!sk[127]) & (text_inx48x) & (!g1678)) + ((!ld) & (!sk[127]) & (text_inx48x) & (g1678)) + ((!ld) & (sk[127]) & (!text_inx48x) & (g1678)) + ((!ld) & (sk[127]) & (text_inx48x) & (g1678)) + ((ld) & (!sk[127]) & (!text_inx48x) & (g1678)) + ((ld) & (!sk[127]) & (text_inx48x) & (!g1678)) + ((ld) & (!sk[127]) & (text_inx48x) & (g1678)) + ((ld) & (sk[127]) & (text_inx48x) & (!g1678)) + ((ld) & (sk[127]) & (text_inx48x) & (g1678)));
	assign g1679 = (((!g403) & (!g467) & (!sk[0]) & (g532) & (!g595)) + ((!g403) & (!g467) & (!sk[0]) & (g532) & (g595)) + ((!g403) & (!g467) & (sk[0]) & (!g532) & (g595)) + ((!g403) & (!g467) & (sk[0]) & (g532) & (!g595)) + ((!g403) & (g467) & (!sk[0]) & (!g532) & (!g595)) + ((!g403) & (g467) & (!sk[0]) & (!g532) & (g595)) + ((!g403) & (g467) & (!sk[0]) & (g532) & (!g595)) + ((!g403) & (g467) & (!sk[0]) & (g532) & (g595)) + ((!g403) & (g467) & (sk[0]) & (!g532) & (!g595)) + ((!g403) & (g467) & (sk[0]) & (g532) & (g595)) + ((g403) & (!g467) & (!sk[0]) & (g532) & (!g595)) + ((g403) & (!g467) & (!sk[0]) & (g532) & (g595)) + ((g403) & (!g467) & (sk[0]) & (!g532) & (!g595)) + ((g403) & (!g467) & (sk[0]) & (g532) & (g595)) + ((g403) & (g467) & (!sk[0]) & (!g532) & (!g595)) + ((g403) & (g467) & (!sk[0]) & (!g532) & (g595)) + ((g403) & (g467) & (!sk[0]) & (g532) & (!g595)) + ((g403) & (g467) & (!sk[0]) & (g532) & (g595)) + ((g403) & (g467) & (sk[0]) & (!g532) & (g595)) + ((g403) & (g467) & (sk[0]) & (g532) & (!g595)));
	assign g1680 = (((!g516) & (!g532) & (!g580) & (!g1163) & (!g1678) & (g1679)) + ((!g516) & (!g532) & (!g580) & (!g1163) & (g1678) & (g1679)) + ((!g516) & (!g532) & (!g580) & (g1163) & (g1678) & (!g1679)) + ((!g516) & (!g532) & (!g580) & (g1163) & (g1678) & (g1679)) + ((!g516) & (!g532) & (g580) & (!g1163) & (!g1678) & (!g1679)) + ((!g516) & (!g532) & (g580) & (!g1163) & (g1678) & (!g1679)) + ((!g516) & (!g532) & (g580) & (g1163) & (g1678) & (!g1679)) + ((!g516) & (!g532) & (g580) & (g1163) & (g1678) & (g1679)) + ((!g516) & (g532) & (!g580) & (!g1163) & (!g1678) & (g1679)) + ((!g516) & (g532) & (!g580) & (!g1163) & (g1678) & (g1679)) + ((!g516) & (g532) & (!g580) & (g1163) & (!g1678) & (!g1679)) + ((!g516) & (g532) & (!g580) & (g1163) & (!g1678) & (g1679)) + ((!g516) & (g532) & (g580) & (!g1163) & (!g1678) & (!g1679)) + ((!g516) & (g532) & (g580) & (!g1163) & (g1678) & (!g1679)) + ((!g516) & (g532) & (g580) & (g1163) & (!g1678) & (!g1679)) + ((!g516) & (g532) & (g580) & (g1163) & (!g1678) & (g1679)) + ((g516) & (!g532) & (!g580) & (!g1163) & (!g1678) & (!g1679)) + ((g516) & (!g532) & (!g580) & (!g1163) & (g1678) & (!g1679)) + ((g516) & (!g532) & (!g580) & (g1163) & (g1678) & (!g1679)) + ((g516) & (!g532) & (!g580) & (g1163) & (g1678) & (g1679)) + ((g516) & (!g532) & (g580) & (!g1163) & (!g1678) & (g1679)) + ((g516) & (!g532) & (g580) & (!g1163) & (g1678) & (g1679)) + ((g516) & (!g532) & (g580) & (g1163) & (g1678) & (!g1679)) + ((g516) & (!g532) & (g580) & (g1163) & (g1678) & (g1679)) + ((g516) & (g532) & (!g580) & (!g1163) & (!g1678) & (!g1679)) + ((g516) & (g532) & (!g580) & (!g1163) & (g1678) & (!g1679)) + ((g516) & (g532) & (!g580) & (g1163) & (!g1678) & (!g1679)) + ((g516) & (g532) & (!g580) & (g1163) & (!g1678) & (g1679)) + ((g516) & (g532) & (g580) & (!g1163) & (!g1678) & (g1679)) + ((g516) & (g532) & (g580) & (!g1163) & (g1678) & (g1679)) + ((g516) & (g532) & (g580) & (g1163) & (!g1678) & (!g1679)) + ((g516) & (g532) & (g580) & (g1163) & (!g1678) & (g1679)));
	assign g2163 = (((!ld) & (!text_inx49x) & (sk[2]) & (g1681)) + ((!ld) & (text_inx49x) & (!sk[2]) & (!g1681)) + ((!ld) & (text_inx49x) & (!sk[2]) & (g1681)) + ((!ld) & (text_inx49x) & (sk[2]) & (g1681)) + ((ld) & (!text_inx49x) & (!sk[2]) & (g1681)) + ((ld) & (text_inx49x) & (!sk[2]) & (!g1681)) + ((ld) & (text_inx49x) & (!sk[2]) & (g1681)) + ((ld) & (text_inx49x) & (sk[2]) & (!g1681)) + ((ld) & (text_inx49x) & (sk[2]) & (g1681)));
	assign g1682 = (((!g410) & (!sk[3]) & (!g467) & (g516) & (!g602)) + ((!g410) & (!sk[3]) & (!g467) & (g516) & (g602)) + ((!g410) & (!sk[3]) & (g467) & (!g516) & (!g602)) + ((!g410) & (!sk[3]) & (g467) & (!g516) & (g602)) + ((!g410) & (!sk[3]) & (g467) & (g516) & (!g602)) + ((!g410) & (!sk[3]) & (g467) & (g516) & (g602)) + ((!g410) & (sk[3]) & (!g467) & (!g516) & (g602)) + ((!g410) & (sk[3]) & (!g467) & (g516) & (!g602)) + ((!g410) & (sk[3]) & (g467) & (!g516) & (!g602)) + ((!g410) & (sk[3]) & (g467) & (g516) & (g602)) + ((g410) & (!sk[3]) & (!g467) & (g516) & (!g602)) + ((g410) & (!sk[3]) & (!g467) & (g516) & (g602)) + ((g410) & (!sk[3]) & (g467) & (!g516) & (!g602)) + ((g410) & (!sk[3]) & (g467) & (!g516) & (g602)) + ((g410) & (!sk[3]) & (g467) & (g516) & (!g602)) + ((g410) & (!sk[3]) & (g467) & (g516) & (g602)) + ((g410) & (sk[3]) & (!g467) & (!g516) & (!g602)) + ((g410) & (sk[3]) & (!g467) & (g516) & (g602)) + ((g410) & (sk[3]) & (g467) & (!g516) & (g602)) + ((g410) & (sk[3]) & (g467) & (g516) & (!g602)));
	assign g2164 = (((!ld) & (!text_inx50x) & (sk[4]) & (g1683)) + ((!ld) & (text_inx50x) & (!sk[4]) & (!g1683)) + ((!ld) & (text_inx50x) & (!sk[4]) & (g1683)) + ((!ld) & (text_inx50x) & (sk[4]) & (g1683)) + ((ld) & (!text_inx50x) & (!sk[4]) & (g1683)) + ((ld) & (text_inx50x) & (!sk[4]) & (!g1683)) + ((ld) & (text_inx50x) & (!sk[4]) & (g1683)) + ((ld) & (text_inx50x) & (sk[4]) & (!g1683)) + ((ld) & (text_inx50x) & (sk[4]) & (g1683)));
	assign g1684 = (((!g474) & (!g546) & (!g609) & (!g1163) & (g1594) & (!g1683)) + ((!g474) & (!g546) & (!g609) & (!g1163) & (g1594) & (g1683)) + ((!g474) & (!g546) & (!g609) & (g1163) & (!g1594) & (g1683)) + ((!g474) & (!g546) & (!g609) & (g1163) & (g1594) & (g1683)) + ((!g474) & (!g546) & (g609) & (!g1163) & (!g1594) & (!g1683)) + ((!g474) & (!g546) & (g609) & (!g1163) & (!g1594) & (g1683)) + ((!g474) & (!g546) & (g609) & (g1163) & (!g1594) & (g1683)) + ((!g474) & (!g546) & (g609) & (g1163) & (g1594) & (g1683)) + ((!g474) & (g546) & (!g609) & (!g1163) & (!g1594) & (!g1683)) + ((!g474) & (g546) & (!g609) & (!g1163) & (!g1594) & (g1683)) + ((!g474) & (g546) & (!g609) & (g1163) & (!g1594) & (!g1683)) + ((!g474) & (g546) & (!g609) & (g1163) & (g1594) & (!g1683)) + ((!g474) & (g546) & (g609) & (!g1163) & (g1594) & (!g1683)) + ((!g474) & (g546) & (g609) & (!g1163) & (g1594) & (g1683)) + ((!g474) & (g546) & (g609) & (g1163) & (!g1594) & (!g1683)) + ((!g474) & (g546) & (g609) & (g1163) & (g1594) & (!g1683)) + ((g474) & (!g546) & (!g609) & (!g1163) & (!g1594) & (!g1683)) + ((g474) & (!g546) & (!g609) & (!g1163) & (!g1594) & (g1683)) + ((g474) & (!g546) & (!g609) & (g1163) & (!g1594) & (g1683)) + ((g474) & (!g546) & (!g609) & (g1163) & (g1594) & (g1683)) + ((g474) & (!g546) & (g609) & (!g1163) & (g1594) & (!g1683)) + ((g474) & (!g546) & (g609) & (!g1163) & (g1594) & (g1683)) + ((g474) & (!g546) & (g609) & (g1163) & (!g1594) & (g1683)) + ((g474) & (!g546) & (g609) & (g1163) & (g1594) & (g1683)) + ((g474) & (g546) & (!g609) & (!g1163) & (g1594) & (!g1683)) + ((g474) & (g546) & (!g609) & (!g1163) & (g1594) & (g1683)) + ((g474) & (g546) & (!g609) & (g1163) & (!g1594) & (!g1683)) + ((g474) & (g546) & (!g609) & (g1163) & (g1594) & (!g1683)) + ((g474) & (g546) & (g609) & (!g1163) & (!g1594) & (!g1683)) + ((g474) & (g546) & (g609) & (!g1163) & (!g1594) & (g1683)) + ((g474) & (g546) & (g609) & (g1163) & (!g1594) & (!g1683)) + ((g474) & (g546) & (g609) & (g1163) & (g1594) & (!g1683)));
	assign g2165 = (((!ld) & (!sk[6]) & (text_inx51x) & (!g1685)) + ((!ld) & (!sk[6]) & (text_inx51x) & (g1685)) + ((!ld) & (sk[6]) & (!text_inx51x) & (g1685)) + ((!ld) & (sk[6]) & (text_inx51x) & (g1685)) + ((ld) & (!sk[6]) & (!text_inx51x) & (g1685)) + ((ld) & (!sk[6]) & (text_inx51x) & (!g1685)) + ((ld) & (!sk[6]) & (text_inx51x) & (g1685)) + ((ld) & (sk[6]) & (text_inx51x) & (!g1685)) + ((ld) & (sk[6]) & (text_inx51x) & (g1685)));
	assign g1686 = (((!sk[7]) & (!g424) & (g481) & (!g616)) + ((!sk[7]) & (!g424) & (g481) & (g616)) + ((!sk[7]) & (g424) & (!g481) & (g616)) + ((!sk[7]) & (g424) & (g481) & (!g616)) + ((!sk[7]) & (g424) & (g481) & (g616)) + ((sk[7]) & (!g424) & (!g481) & (g616)) + ((sk[7]) & (!g424) & (g481) & (!g616)) + ((sk[7]) & (g424) & (!g481) & (!g616)) + ((sk[7]) & (g424) & (g481) & (g616)));
	assign g1687 = (((!g488) & (!g516) & (!g545) & (!g553) & (sk[8]) & (g580)) + ((!g488) & (!g516) & (!g545) & (g553) & (sk[8]) & (!g580)) + ((!g488) & (!g516) & (g545) & (!g553) & (sk[8]) & (!g580)) + ((!g488) & (!g516) & (g545) & (g553) & (sk[8]) & (g580)) + ((!g488) & (g516) & (!g545) & (!g553) & (!sk[8]) & (!g580)) + ((!g488) & (g516) & (!g545) & (!g553) & (!sk[8]) & (g580)) + ((!g488) & (g516) & (!g545) & (!g553) & (sk[8]) & (!g580)) + ((!g488) & (g516) & (!g545) & (g553) & (!sk[8]) & (!g580)) + ((!g488) & (g516) & (!g545) & (g553) & (!sk[8]) & (g580)) + ((!g488) & (g516) & (!g545) & (g553) & (sk[8]) & (g580)) + ((!g488) & (g516) & (g545) & (!g553) & (!sk[8]) & (!g580)) + ((!g488) & (g516) & (g545) & (!g553) & (!sk[8]) & (g580)) + ((!g488) & (g516) & (g545) & (!g553) & (sk[8]) & (g580)) + ((!g488) & (g516) & (g545) & (g553) & (!sk[8]) & (!g580)) + ((!g488) & (g516) & (g545) & (g553) & (!sk[8]) & (g580)) + ((!g488) & (g516) & (g545) & (g553) & (sk[8]) & (!g580)) + ((g488) & (!g516) & (!g545) & (!g553) & (!sk[8]) & (!g580)) + ((g488) & (!g516) & (!g545) & (!g553) & (!sk[8]) & (g580)) + ((g488) & (!g516) & (!g545) & (!g553) & (sk[8]) & (!g580)) + ((g488) & (!g516) & (!g545) & (g553) & (!sk[8]) & (!g580)) + ((g488) & (!g516) & (!g545) & (g553) & (!sk[8]) & (g580)) + ((g488) & (!g516) & (!g545) & (g553) & (sk[8]) & (g580)) + ((g488) & (!g516) & (g545) & (!g553) & (!sk[8]) & (!g580)) + ((g488) & (!g516) & (g545) & (!g553) & (!sk[8]) & (g580)) + ((g488) & (!g516) & (g545) & (!g553) & (sk[8]) & (g580)) + ((g488) & (!g516) & (g545) & (g553) & (!sk[8]) & (!g580)) + ((g488) & (!g516) & (g545) & (g553) & (!sk[8]) & (g580)) + ((g488) & (!g516) & (g545) & (g553) & (sk[8]) & (!g580)) + ((g488) & (g516) & (!g545) & (!g553) & (!sk[8]) & (!g580)) + ((g488) & (g516) & (!g545) & (!g553) & (!sk[8]) & (g580)) + ((g488) & (g516) & (!g545) & (!g553) & (sk[8]) & (g580)) + ((g488) & (g516) & (!g545) & (g553) & (!sk[8]) & (!g580)) + ((g488) & (g516) & (!g545) & (g553) & (!sk[8]) & (g580)) + ((g488) & (g516) & (!g545) & (g553) & (sk[8]) & (!g580)) + ((g488) & (g516) & (g545) & (!g553) & (!sk[8]) & (!g580)) + ((g488) & (g516) & (g545) & (!g553) & (!sk[8]) & (g580)) + ((g488) & (g516) & (g545) & (!g553) & (sk[8]) & (!g580)) + ((g488) & (g516) & (g545) & (g553) & (!sk[8]) & (!g580)) + ((g488) & (g516) & (g545) & (g553) & (!sk[8]) & (g580)) + ((g488) & (g516) & (g545) & (g553) & (sk[8]) & (g580)));
	assign g1688 = (((!g553) & (!g1163) & (sk[9]) & (!g1685) & (!g1686) & (g1687)) + ((!g553) & (!g1163) & (sk[9]) & (!g1685) & (g1686) & (!g1687)) + ((!g553) & (!g1163) & (sk[9]) & (g1685) & (!g1686) & (g1687)) + ((!g553) & (!g1163) & (sk[9]) & (g1685) & (g1686) & (!g1687)) + ((!g553) & (g1163) & (!sk[9]) & (!g1685) & (!g1686) & (!g1687)) + ((!g553) & (g1163) & (!sk[9]) & (!g1685) & (!g1686) & (g1687)) + ((!g553) & (g1163) & (!sk[9]) & (!g1685) & (g1686) & (!g1687)) + ((!g553) & (g1163) & (!sk[9]) & (!g1685) & (g1686) & (g1687)) + ((!g553) & (g1163) & (!sk[9]) & (g1685) & (!g1686) & (!g1687)) + ((!g553) & (g1163) & (!sk[9]) & (g1685) & (!g1686) & (g1687)) + ((!g553) & (g1163) & (!sk[9]) & (g1685) & (g1686) & (!g1687)) + ((!g553) & (g1163) & (!sk[9]) & (g1685) & (g1686) & (g1687)) + ((!g553) & (g1163) & (sk[9]) & (g1685) & (!g1686) & (!g1687)) + ((!g553) & (g1163) & (sk[9]) & (g1685) & (!g1686) & (g1687)) + ((!g553) & (g1163) & (sk[9]) & (g1685) & (g1686) & (!g1687)) + ((!g553) & (g1163) & (sk[9]) & (g1685) & (g1686) & (g1687)) + ((g553) & (!g1163) & (!sk[9]) & (!g1685) & (!g1686) & (!g1687)) + ((g553) & (!g1163) & (!sk[9]) & (!g1685) & (!g1686) & (g1687)) + ((g553) & (!g1163) & (!sk[9]) & (!g1685) & (g1686) & (!g1687)) + ((g553) & (!g1163) & (!sk[9]) & (!g1685) & (g1686) & (g1687)) + ((g553) & (!g1163) & (!sk[9]) & (g1685) & (!g1686) & (!g1687)) + ((g553) & (!g1163) & (!sk[9]) & (g1685) & (!g1686) & (g1687)) + ((g553) & (!g1163) & (!sk[9]) & (g1685) & (g1686) & (!g1687)) + ((g553) & (!g1163) & (!sk[9]) & (g1685) & (g1686) & (g1687)) + ((g553) & (!g1163) & (sk[9]) & (!g1685) & (!g1686) & (g1687)) + ((g553) & (!g1163) & (sk[9]) & (!g1685) & (g1686) & (!g1687)) + ((g553) & (!g1163) & (sk[9]) & (g1685) & (!g1686) & (g1687)) + ((g553) & (!g1163) & (sk[9]) & (g1685) & (g1686) & (!g1687)) + ((g553) & (g1163) & (!sk[9]) & (!g1685) & (!g1686) & (!g1687)) + ((g553) & (g1163) & (!sk[9]) & (!g1685) & (!g1686) & (g1687)) + ((g553) & (g1163) & (!sk[9]) & (!g1685) & (g1686) & (!g1687)) + ((g553) & (g1163) & (!sk[9]) & (!g1685) & (g1686) & (g1687)) + ((g553) & (g1163) & (!sk[9]) & (g1685) & (!g1686) & (!g1687)) + ((g553) & (g1163) & (!sk[9]) & (g1685) & (!g1686) & (g1687)) + ((g553) & (g1163) & (!sk[9]) & (g1685) & (g1686) & (!g1687)) + ((g553) & (g1163) & (!sk[9]) & (g1685) & (g1686) & (g1687)) + ((g553) & (g1163) & (sk[9]) & (!g1685) & (!g1686) & (!g1687)) + ((g553) & (g1163) & (sk[9]) & (!g1685) & (!g1686) & (g1687)) + ((g553) & (g1163) & (sk[9]) & (!g1685) & (g1686) & (!g1687)) + ((g553) & (g1163) & (sk[9]) & (!g1685) & (g1686) & (g1687)));
	assign g2166 = (((!sk[10]) & (!ld) & (text_inx54x) & (!g1689)) + ((!sk[10]) & (!ld) & (text_inx54x) & (g1689)) + ((!sk[10]) & (ld) & (!text_inx54x) & (g1689)) + ((!sk[10]) & (ld) & (text_inx54x) & (!g1689)) + ((!sk[10]) & (ld) & (text_inx54x) & (g1689)) + ((sk[10]) & (!ld) & (!text_inx54x) & (g1689)) + ((sk[10]) & (!ld) & (text_inx54x) & (g1689)) + ((sk[10]) & (ld) & (text_inx54x) & (!g1689)) + ((sk[10]) & (ld) & (text_inx54x) & (g1689)));
	assign g1690 = (((!g502) & (!g574) & (!g637) & (!g1163) & (g1598) & (!g1689)) + ((!g502) & (!g574) & (!g637) & (!g1163) & (g1598) & (g1689)) + ((!g502) & (!g574) & (!g637) & (g1163) & (!g1598) & (g1689)) + ((!g502) & (!g574) & (!g637) & (g1163) & (g1598) & (g1689)) + ((!g502) & (!g574) & (g637) & (!g1163) & (!g1598) & (!g1689)) + ((!g502) & (!g574) & (g637) & (!g1163) & (!g1598) & (g1689)) + ((!g502) & (!g574) & (g637) & (g1163) & (!g1598) & (g1689)) + ((!g502) & (!g574) & (g637) & (g1163) & (g1598) & (g1689)) + ((!g502) & (g574) & (!g637) & (!g1163) & (!g1598) & (!g1689)) + ((!g502) & (g574) & (!g637) & (!g1163) & (!g1598) & (g1689)) + ((!g502) & (g574) & (!g637) & (g1163) & (!g1598) & (!g1689)) + ((!g502) & (g574) & (!g637) & (g1163) & (g1598) & (!g1689)) + ((!g502) & (g574) & (g637) & (!g1163) & (g1598) & (!g1689)) + ((!g502) & (g574) & (g637) & (!g1163) & (g1598) & (g1689)) + ((!g502) & (g574) & (g637) & (g1163) & (!g1598) & (!g1689)) + ((!g502) & (g574) & (g637) & (g1163) & (g1598) & (!g1689)) + ((g502) & (!g574) & (!g637) & (!g1163) & (!g1598) & (!g1689)) + ((g502) & (!g574) & (!g637) & (!g1163) & (!g1598) & (g1689)) + ((g502) & (!g574) & (!g637) & (g1163) & (!g1598) & (g1689)) + ((g502) & (!g574) & (!g637) & (g1163) & (g1598) & (g1689)) + ((g502) & (!g574) & (g637) & (!g1163) & (g1598) & (!g1689)) + ((g502) & (!g574) & (g637) & (!g1163) & (g1598) & (g1689)) + ((g502) & (!g574) & (g637) & (g1163) & (!g1598) & (g1689)) + ((g502) & (!g574) & (g637) & (g1163) & (g1598) & (g1689)) + ((g502) & (g574) & (!g637) & (!g1163) & (g1598) & (!g1689)) + ((g502) & (g574) & (!g637) & (!g1163) & (g1598) & (g1689)) + ((g502) & (g574) & (!g637) & (g1163) & (!g1598) & (!g1689)) + ((g502) & (g574) & (!g637) & (g1163) & (g1598) & (!g1689)) + ((g502) & (g574) & (g637) & (!g1163) & (!g1598) & (!g1689)) + ((g502) & (g574) & (g637) & (!g1163) & (!g1598) & (g1689)) + ((g502) & (g574) & (g637) & (g1163) & (!g1598) & (!g1689)) + ((g502) & (g574) & (g637) & (g1163) & (g1598) & (!g1689)));
	assign g2167 = (((!sk[12]) & (!ld) & (text_inx53x) & (!g1691)) + ((!sk[12]) & (!ld) & (text_inx53x) & (g1691)) + ((!sk[12]) & (ld) & (!text_inx53x) & (g1691)) + ((!sk[12]) & (ld) & (text_inx53x) & (!g1691)) + ((!sk[12]) & (ld) & (text_inx53x) & (g1691)) + ((sk[12]) & (!ld) & (!text_inx53x) & (g1691)) + ((sk[12]) & (!ld) & (text_inx53x) & (g1691)) + ((sk[12]) & (ld) & (text_inx53x) & (!g1691)) + ((sk[12]) & (ld) & (text_inx53x) & (g1691)));
	assign g1692 = (((!g495) & (!g567) & (!g630) & (!g1163) & (g1601) & (!g1691)) + ((!g495) & (!g567) & (!g630) & (!g1163) & (g1601) & (g1691)) + ((!g495) & (!g567) & (!g630) & (g1163) & (!g1601) & (g1691)) + ((!g495) & (!g567) & (!g630) & (g1163) & (g1601) & (g1691)) + ((!g495) & (!g567) & (g630) & (!g1163) & (!g1601) & (!g1691)) + ((!g495) & (!g567) & (g630) & (!g1163) & (!g1601) & (g1691)) + ((!g495) & (!g567) & (g630) & (g1163) & (!g1601) & (g1691)) + ((!g495) & (!g567) & (g630) & (g1163) & (g1601) & (g1691)) + ((!g495) & (g567) & (!g630) & (!g1163) & (!g1601) & (!g1691)) + ((!g495) & (g567) & (!g630) & (!g1163) & (!g1601) & (g1691)) + ((!g495) & (g567) & (!g630) & (g1163) & (!g1601) & (!g1691)) + ((!g495) & (g567) & (!g630) & (g1163) & (g1601) & (!g1691)) + ((!g495) & (g567) & (g630) & (!g1163) & (g1601) & (!g1691)) + ((!g495) & (g567) & (g630) & (!g1163) & (g1601) & (g1691)) + ((!g495) & (g567) & (g630) & (g1163) & (!g1601) & (!g1691)) + ((!g495) & (g567) & (g630) & (g1163) & (g1601) & (!g1691)) + ((g495) & (!g567) & (!g630) & (!g1163) & (!g1601) & (!g1691)) + ((g495) & (!g567) & (!g630) & (!g1163) & (!g1601) & (g1691)) + ((g495) & (!g567) & (!g630) & (g1163) & (!g1601) & (g1691)) + ((g495) & (!g567) & (!g630) & (g1163) & (g1601) & (g1691)) + ((g495) & (!g567) & (g630) & (!g1163) & (g1601) & (!g1691)) + ((g495) & (!g567) & (g630) & (!g1163) & (g1601) & (g1691)) + ((g495) & (!g567) & (g630) & (g1163) & (!g1601) & (g1691)) + ((g495) & (!g567) & (g630) & (g1163) & (g1601) & (g1691)) + ((g495) & (g567) & (!g630) & (!g1163) & (g1601) & (!g1691)) + ((g495) & (g567) & (!g630) & (!g1163) & (g1601) & (g1691)) + ((g495) & (g567) & (!g630) & (g1163) & (!g1601) & (!g1691)) + ((g495) & (g567) & (!g630) & (g1163) & (g1601) & (!g1691)) + ((g495) & (g567) & (g630) & (!g1163) & (!g1601) & (!g1691)) + ((g495) & (g567) & (g630) & (!g1163) & (!g1601) & (g1691)) + ((g495) & (g567) & (g630) & (g1163) & (!g1601) & (!g1691)) + ((g495) & (g567) & (g630) & (g1163) & (g1601) & (!g1691)));
	assign g2168 = (((!sk[14]) & (!ld) & (text_inx52x) & (!g1693)) + ((!sk[14]) & (!ld) & (text_inx52x) & (g1693)) + ((!sk[14]) & (ld) & (!text_inx52x) & (g1693)) + ((!sk[14]) & (ld) & (text_inx52x) & (!g1693)) + ((!sk[14]) & (ld) & (text_inx52x) & (g1693)) + ((sk[14]) & (!ld) & (!text_inx52x) & (g1693)) + ((sk[14]) & (!ld) & (text_inx52x) & (g1693)) + ((sk[14]) & (ld) & (text_inx52x) & (!g1693)) + ((sk[14]) & (ld) & (text_inx52x) & (g1693)));
	assign g1694 = (((!g488) & (!sk[15]) & (g516) & (!g560) & (!g580) & (!g623)) + ((!g488) & (!sk[15]) & (g516) & (!g560) & (!g580) & (g623)) + ((!g488) & (!sk[15]) & (g516) & (!g560) & (g580) & (!g623)) + ((!g488) & (!sk[15]) & (g516) & (!g560) & (g580) & (g623)) + ((!g488) & (!sk[15]) & (g516) & (g560) & (!g580) & (!g623)) + ((!g488) & (!sk[15]) & (g516) & (g560) & (!g580) & (g623)) + ((!g488) & (!sk[15]) & (g516) & (g560) & (g580) & (!g623)) + ((!g488) & (!sk[15]) & (g516) & (g560) & (g580) & (g623)) + ((!g488) & (sk[15]) & (!g516) & (!g560) & (!g580) & (g623)) + ((!g488) & (sk[15]) & (!g516) & (!g560) & (g580) & (!g623)) + ((!g488) & (sk[15]) & (!g516) & (g560) & (!g580) & (!g623)) + ((!g488) & (sk[15]) & (!g516) & (g560) & (g580) & (g623)) + ((!g488) & (sk[15]) & (g516) & (!g560) & (!g580) & (!g623)) + ((!g488) & (sk[15]) & (g516) & (!g560) & (g580) & (g623)) + ((!g488) & (sk[15]) & (g516) & (g560) & (!g580) & (g623)) + ((!g488) & (sk[15]) & (g516) & (g560) & (g580) & (!g623)) + ((g488) & (!sk[15]) & (!g516) & (!g560) & (!g580) & (!g623)) + ((g488) & (!sk[15]) & (!g516) & (!g560) & (!g580) & (g623)) + ((g488) & (!sk[15]) & (!g516) & (!g560) & (g580) & (!g623)) + ((g488) & (!sk[15]) & (!g516) & (!g560) & (g580) & (g623)) + ((g488) & (!sk[15]) & (!g516) & (g560) & (!g580) & (!g623)) + ((g488) & (!sk[15]) & (!g516) & (g560) & (!g580) & (g623)) + ((g488) & (!sk[15]) & (!g516) & (g560) & (g580) & (!g623)) + ((g488) & (!sk[15]) & (!g516) & (g560) & (g580) & (g623)) + ((g488) & (!sk[15]) & (g516) & (!g560) & (!g580) & (!g623)) + ((g488) & (!sk[15]) & (g516) & (!g560) & (!g580) & (g623)) + ((g488) & (!sk[15]) & (g516) & (!g560) & (g580) & (!g623)) + ((g488) & (!sk[15]) & (g516) & (!g560) & (g580) & (g623)) + ((g488) & (!sk[15]) & (g516) & (g560) & (!g580) & (!g623)) + ((g488) & (!sk[15]) & (g516) & (g560) & (!g580) & (g623)) + ((g488) & (!sk[15]) & (g516) & (g560) & (g580) & (!g623)) + ((g488) & (!sk[15]) & (g516) & (g560) & (g580) & (g623)) + ((g488) & (sk[15]) & (!g516) & (!g560) & (!g580) & (!g623)) + ((g488) & (sk[15]) & (!g516) & (!g560) & (g580) & (g623)) + ((g488) & (sk[15]) & (!g516) & (g560) & (!g580) & (g623)) + ((g488) & (sk[15]) & (!g516) & (g560) & (g580) & (!g623)) + ((g488) & (sk[15]) & (g516) & (!g560) & (!g580) & (g623)) + ((g488) & (sk[15]) & (g516) & (!g560) & (g580) & (!g623)) + ((g488) & (sk[15]) & (g516) & (g560) & (!g580) & (!g623)) + ((g488) & (sk[15]) & (g516) & (g560) & (g580) & (g623)));
	assign g1695 = (((!g560) & (!g1163) & (!g1604) & (sk[16]) & (!g1693) & (g1694)) + ((!g560) & (!g1163) & (!g1604) & (sk[16]) & (g1693) & (g1694)) + ((!g560) & (!g1163) & (g1604) & (sk[16]) & (!g1693) & (!g1694)) + ((!g560) & (!g1163) & (g1604) & (sk[16]) & (g1693) & (!g1694)) + ((!g560) & (g1163) & (!g1604) & (!sk[16]) & (!g1693) & (!g1694)) + ((!g560) & (g1163) & (!g1604) & (!sk[16]) & (!g1693) & (g1694)) + ((!g560) & (g1163) & (!g1604) & (!sk[16]) & (g1693) & (!g1694)) + ((!g560) & (g1163) & (!g1604) & (!sk[16]) & (g1693) & (g1694)) + ((!g560) & (g1163) & (!g1604) & (sk[16]) & (g1693) & (!g1694)) + ((!g560) & (g1163) & (!g1604) & (sk[16]) & (g1693) & (g1694)) + ((!g560) & (g1163) & (g1604) & (!sk[16]) & (!g1693) & (!g1694)) + ((!g560) & (g1163) & (g1604) & (!sk[16]) & (!g1693) & (g1694)) + ((!g560) & (g1163) & (g1604) & (!sk[16]) & (g1693) & (!g1694)) + ((!g560) & (g1163) & (g1604) & (!sk[16]) & (g1693) & (g1694)) + ((!g560) & (g1163) & (g1604) & (sk[16]) & (g1693) & (!g1694)) + ((!g560) & (g1163) & (g1604) & (sk[16]) & (g1693) & (g1694)) + ((g560) & (!g1163) & (!g1604) & (!sk[16]) & (!g1693) & (!g1694)) + ((g560) & (!g1163) & (!g1604) & (!sk[16]) & (!g1693) & (g1694)) + ((g560) & (!g1163) & (!g1604) & (!sk[16]) & (g1693) & (!g1694)) + ((g560) & (!g1163) & (!g1604) & (!sk[16]) & (g1693) & (g1694)) + ((g560) & (!g1163) & (!g1604) & (sk[16]) & (!g1693) & (g1694)) + ((g560) & (!g1163) & (!g1604) & (sk[16]) & (g1693) & (g1694)) + ((g560) & (!g1163) & (g1604) & (!sk[16]) & (!g1693) & (!g1694)) + ((g560) & (!g1163) & (g1604) & (!sk[16]) & (!g1693) & (g1694)) + ((g560) & (!g1163) & (g1604) & (!sk[16]) & (g1693) & (!g1694)) + ((g560) & (!g1163) & (g1604) & (!sk[16]) & (g1693) & (g1694)) + ((g560) & (!g1163) & (g1604) & (sk[16]) & (!g1693) & (!g1694)) + ((g560) & (!g1163) & (g1604) & (sk[16]) & (g1693) & (!g1694)) + ((g560) & (g1163) & (!g1604) & (!sk[16]) & (!g1693) & (!g1694)) + ((g560) & (g1163) & (!g1604) & (!sk[16]) & (!g1693) & (g1694)) + ((g560) & (g1163) & (!g1604) & (!sk[16]) & (g1693) & (!g1694)) + ((g560) & (g1163) & (!g1604) & (!sk[16]) & (g1693) & (g1694)) + ((g560) & (g1163) & (!g1604) & (sk[16]) & (!g1693) & (!g1694)) + ((g560) & (g1163) & (!g1604) & (sk[16]) & (!g1693) & (g1694)) + ((g560) & (g1163) & (g1604) & (!sk[16]) & (!g1693) & (!g1694)) + ((g560) & (g1163) & (g1604) & (!sk[16]) & (!g1693) & (g1694)) + ((g560) & (g1163) & (g1604) & (!sk[16]) & (g1693) & (!g1694)) + ((g560) & (g1163) & (g1604) & (!sk[16]) & (g1693) & (g1694)) + ((g560) & (g1163) & (g1604) & (sk[16]) & (!g1693) & (!g1694)) + ((g560) & (g1163) & (g1604) & (sk[16]) & (!g1693) & (g1694)));
	assign g2169 = (((!ld) & (!text_inx55x) & (sk[17]) & (g1696)) + ((!ld) & (text_inx55x) & (!sk[17]) & (!g1696)) + ((!ld) & (text_inx55x) & (!sk[17]) & (g1696)) + ((!ld) & (text_inx55x) & (sk[17]) & (g1696)) + ((ld) & (!text_inx55x) & (!sk[17]) & (g1696)) + ((ld) & (text_inx55x) & (!sk[17]) & (!g1696)) + ((ld) & (text_inx55x) & (!sk[17]) & (g1696)) + ((ld) & (text_inx55x) & (sk[17]) & (!g1696)) + ((ld) & (text_inx55x) & (sk[17]) & (g1696)));
	assign g1697 = (((!g509) & (!g581) & (!g644) & (!g1163) & (g1608) & (!g1696)) + ((!g509) & (!g581) & (!g644) & (!g1163) & (g1608) & (g1696)) + ((!g509) & (!g581) & (!g644) & (g1163) & (!g1608) & (g1696)) + ((!g509) & (!g581) & (!g644) & (g1163) & (g1608) & (g1696)) + ((!g509) & (!g581) & (g644) & (!g1163) & (!g1608) & (!g1696)) + ((!g509) & (!g581) & (g644) & (!g1163) & (!g1608) & (g1696)) + ((!g509) & (!g581) & (g644) & (g1163) & (!g1608) & (g1696)) + ((!g509) & (!g581) & (g644) & (g1163) & (g1608) & (g1696)) + ((!g509) & (g581) & (!g644) & (!g1163) & (!g1608) & (!g1696)) + ((!g509) & (g581) & (!g644) & (!g1163) & (!g1608) & (g1696)) + ((!g509) & (g581) & (!g644) & (g1163) & (!g1608) & (!g1696)) + ((!g509) & (g581) & (!g644) & (g1163) & (g1608) & (!g1696)) + ((!g509) & (g581) & (g644) & (!g1163) & (g1608) & (!g1696)) + ((!g509) & (g581) & (g644) & (!g1163) & (g1608) & (g1696)) + ((!g509) & (g581) & (g644) & (g1163) & (!g1608) & (!g1696)) + ((!g509) & (g581) & (g644) & (g1163) & (g1608) & (!g1696)) + ((g509) & (!g581) & (!g644) & (!g1163) & (!g1608) & (!g1696)) + ((g509) & (!g581) & (!g644) & (!g1163) & (!g1608) & (g1696)) + ((g509) & (!g581) & (!g644) & (g1163) & (!g1608) & (g1696)) + ((g509) & (!g581) & (!g644) & (g1163) & (g1608) & (g1696)) + ((g509) & (!g581) & (g644) & (!g1163) & (g1608) & (!g1696)) + ((g509) & (!g581) & (g644) & (!g1163) & (g1608) & (g1696)) + ((g509) & (!g581) & (g644) & (g1163) & (!g1608) & (g1696)) + ((g509) & (!g581) & (g644) & (g1163) & (g1608) & (g1696)) + ((g509) & (g581) & (!g644) & (!g1163) & (g1608) & (!g1696)) + ((g509) & (g581) & (!g644) & (!g1163) & (g1608) & (g1696)) + ((g509) & (g581) & (!g644) & (g1163) & (!g1608) & (!g1696)) + ((g509) & (g581) & (!g644) & (g1163) & (g1608) & (!g1696)) + ((g509) & (g581) & (g644) & (!g1163) & (!g1608) & (!g1696)) + ((g509) & (g581) & (g644) & (!g1163) & (!g1608) & (g1696)) + ((g509) & (g581) & (g644) & (g1163) & (!g1608) & (!g1696)) + ((g509) & (g581) & (g644) & (g1163) & (g1608) & (!g1696)));
	assign g1698 = (((!ld) & (!g788) & (!g1044) & (g1358) & (sk[19]) & (!keyx80x)) + ((!ld) & (!g788) & (!g1044) & (g1358) & (sk[19]) & (keyx80x)) + ((!ld) & (!g788) & (g1044) & (!g1358) & (sk[19]) & (!keyx80x)) + ((!ld) & (!g788) & (g1044) & (!g1358) & (sk[19]) & (keyx80x)) + ((!ld) & (g788) & (!g1044) & (!g1358) & (!sk[19]) & (!keyx80x)) + ((!ld) & (g788) & (!g1044) & (!g1358) & (!sk[19]) & (keyx80x)) + ((!ld) & (g788) & (!g1044) & (!g1358) & (sk[19]) & (!keyx80x)) + ((!ld) & (g788) & (!g1044) & (!g1358) & (sk[19]) & (keyx80x)) + ((!ld) & (g788) & (!g1044) & (g1358) & (!sk[19]) & (!keyx80x)) + ((!ld) & (g788) & (!g1044) & (g1358) & (!sk[19]) & (keyx80x)) + ((!ld) & (g788) & (g1044) & (!g1358) & (!sk[19]) & (!keyx80x)) + ((!ld) & (g788) & (g1044) & (!g1358) & (!sk[19]) & (keyx80x)) + ((!ld) & (g788) & (g1044) & (g1358) & (!sk[19]) & (!keyx80x)) + ((!ld) & (g788) & (g1044) & (g1358) & (!sk[19]) & (keyx80x)) + ((!ld) & (g788) & (g1044) & (g1358) & (sk[19]) & (!keyx80x)) + ((!ld) & (g788) & (g1044) & (g1358) & (sk[19]) & (keyx80x)) + ((ld) & (!g788) & (!g1044) & (!g1358) & (!sk[19]) & (!keyx80x)) + ((ld) & (!g788) & (!g1044) & (!g1358) & (!sk[19]) & (keyx80x)) + ((ld) & (!g788) & (!g1044) & (!g1358) & (sk[19]) & (keyx80x)) + ((ld) & (!g788) & (!g1044) & (g1358) & (!sk[19]) & (!keyx80x)) + ((ld) & (!g788) & (!g1044) & (g1358) & (!sk[19]) & (keyx80x)) + ((ld) & (!g788) & (!g1044) & (g1358) & (sk[19]) & (keyx80x)) + ((ld) & (!g788) & (g1044) & (!g1358) & (!sk[19]) & (!keyx80x)) + ((ld) & (!g788) & (g1044) & (!g1358) & (!sk[19]) & (keyx80x)) + ((ld) & (!g788) & (g1044) & (!g1358) & (sk[19]) & (keyx80x)) + ((ld) & (!g788) & (g1044) & (g1358) & (!sk[19]) & (!keyx80x)) + ((ld) & (!g788) & (g1044) & (g1358) & (!sk[19]) & (keyx80x)) + ((ld) & (!g788) & (g1044) & (g1358) & (sk[19]) & (keyx80x)) + ((ld) & (g788) & (!g1044) & (!g1358) & (!sk[19]) & (!keyx80x)) + ((ld) & (g788) & (!g1044) & (!g1358) & (!sk[19]) & (keyx80x)) + ((ld) & (g788) & (!g1044) & (!g1358) & (sk[19]) & (keyx80x)) + ((ld) & (g788) & (!g1044) & (g1358) & (!sk[19]) & (!keyx80x)) + ((ld) & (g788) & (!g1044) & (g1358) & (!sk[19]) & (keyx80x)) + ((ld) & (g788) & (!g1044) & (g1358) & (sk[19]) & (keyx80x)) + ((ld) & (g788) & (g1044) & (!g1358) & (!sk[19]) & (!keyx80x)) + ((ld) & (g788) & (g1044) & (!g1358) & (!sk[19]) & (keyx80x)) + ((ld) & (g788) & (g1044) & (!g1358) & (sk[19]) & (keyx80x)) + ((ld) & (g788) & (g1044) & (g1358) & (!sk[19]) & (!keyx80x)) + ((ld) & (g788) & (g1044) & (g1358) & (!sk[19]) & (keyx80x)) + ((ld) & (g788) & (g1044) & (g1358) & (sk[19]) & (keyx80x)));
	assign g1699 = (((!ld) & (!sk[20]) & (g795) & (!g1051) & (!g1365) & (!keyx81x)) + ((!ld) & (!sk[20]) & (g795) & (!g1051) & (!g1365) & (keyx81x)) + ((!ld) & (!sk[20]) & (g795) & (!g1051) & (g1365) & (!keyx81x)) + ((!ld) & (!sk[20]) & (g795) & (!g1051) & (g1365) & (keyx81x)) + ((!ld) & (!sk[20]) & (g795) & (g1051) & (!g1365) & (!keyx81x)) + ((!ld) & (!sk[20]) & (g795) & (g1051) & (!g1365) & (keyx81x)) + ((!ld) & (!sk[20]) & (g795) & (g1051) & (g1365) & (!keyx81x)) + ((!ld) & (!sk[20]) & (g795) & (g1051) & (g1365) & (keyx81x)) + ((!ld) & (sk[20]) & (!g795) & (!g1051) & (g1365) & (!keyx81x)) + ((!ld) & (sk[20]) & (!g795) & (!g1051) & (g1365) & (keyx81x)) + ((!ld) & (sk[20]) & (!g795) & (g1051) & (!g1365) & (!keyx81x)) + ((!ld) & (sk[20]) & (!g795) & (g1051) & (!g1365) & (keyx81x)) + ((!ld) & (sk[20]) & (g795) & (!g1051) & (!g1365) & (!keyx81x)) + ((!ld) & (sk[20]) & (g795) & (!g1051) & (!g1365) & (keyx81x)) + ((!ld) & (sk[20]) & (g795) & (g1051) & (g1365) & (!keyx81x)) + ((!ld) & (sk[20]) & (g795) & (g1051) & (g1365) & (keyx81x)) + ((ld) & (!sk[20]) & (!g795) & (!g1051) & (!g1365) & (!keyx81x)) + ((ld) & (!sk[20]) & (!g795) & (!g1051) & (!g1365) & (keyx81x)) + ((ld) & (!sk[20]) & (!g795) & (!g1051) & (g1365) & (!keyx81x)) + ((ld) & (!sk[20]) & (!g795) & (!g1051) & (g1365) & (keyx81x)) + ((ld) & (!sk[20]) & (!g795) & (g1051) & (!g1365) & (!keyx81x)) + ((ld) & (!sk[20]) & (!g795) & (g1051) & (!g1365) & (keyx81x)) + ((ld) & (!sk[20]) & (!g795) & (g1051) & (g1365) & (!keyx81x)) + ((ld) & (!sk[20]) & (!g795) & (g1051) & (g1365) & (keyx81x)) + ((ld) & (!sk[20]) & (g795) & (!g1051) & (!g1365) & (!keyx81x)) + ((ld) & (!sk[20]) & (g795) & (!g1051) & (!g1365) & (keyx81x)) + ((ld) & (!sk[20]) & (g795) & (!g1051) & (g1365) & (!keyx81x)) + ((ld) & (!sk[20]) & (g795) & (!g1051) & (g1365) & (keyx81x)) + ((ld) & (!sk[20]) & (g795) & (g1051) & (!g1365) & (!keyx81x)) + ((ld) & (!sk[20]) & (g795) & (g1051) & (!g1365) & (keyx81x)) + ((ld) & (!sk[20]) & (g795) & (g1051) & (g1365) & (!keyx81x)) + ((ld) & (!sk[20]) & (g795) & (g1051) & (g1365) & (keyx81x)) + ((ld) & (sk[20]) & (!g795) & (!g1051) & (!g1365) & (keyx81x)) + ((ld) & (sk[20]) & (!g795) & (!g1051) & (g1365) & (keyx81x)) + ((ld) & (sk[20]) & (!g795) & (g1051) & (!g1365) & (keyx81x)) + ((ld) & (sk[20]) & (!g795) & (g1051) & (g1365) & (keyx81x)) + ((ld) & (sk[20]) & (g795) & (!g1051) & (!g1365) & (keyx81x)) + ((ld) & (sk[20]) & (g795) & (!g1051) & (g1365) & (keyx81x)) + ((ld) & (sk[20]) & (g795) & (g1051) & (!g1365) & (keyx81x)) + ((ld) & (sk[20]) & (g795) & (g1051) & (g1365) & (keyx81x)));
	assign g1700 = (((!ld) & (!sk[21]) & (g802) & (!g1058) & (!g1372) & (!keyx82x)) + ((!ld) & (!sk[21]) & (g802) & (!g1058) & (!g1372) & (keyx82x)) + ((!ld) & (!sk[21]) & (g802) & (!g1058) & (g1372) & (!keyx82x)) + ((!ld) & (!sk[21]) & (g802) & (!g1058) & (g1372) & (keyx82x)) + ((!ld) & (!sk[21]) & (g802) & (g1058) & (!g1372) & (!keyx82x)) + ((!ld) & (!sk[21]) & (g802) & (g1058) & (!g1372) & (keyx82x)) + ((!ld) & (!sk[21]) & (g802) & (g1058) & (g1372) & (!keyx82x)) + ((!ld) & (!sk[21]) & (g802) & (g1058) & (g1372) & (keyx82x)) + ((!ld) & (sk[21]) & (!g802) & (!g1058) & (g1372) & (!keyx82x)) + ((!ld) & (sk[21]) & (!g802) & (!g1058) & (g1372) & (keyx82x)) + ((!ld) & (sk[21]) & (!g802) & (g1058) & (!g1372) & (!keyx82x)) + ((!ld) & (sk[21]) & (!g802) & (g1058) & (!g1372) & (keyx82x)) + ((!ld) & (sk[21]) & (g802) & (!g1058) & (!g1372) & (!keyx82x)) + ((!ld) & (sk[21]) & (g802) & (!g1058) & (!g1372) & (keyx82x)) + ((!ld) & (sk[21]) & (g802) & (g1058) & (g1372) & (!keyx82x)) + ((!ld) & (sk[21]) & (g802) & (g1058) & (g1372) & (keyx82x)) + ((ld) & (!sk[21]) & (!g802) & (!g1058) & (!g1372) & (!keyx82x)) + ((ld) & (!sk[21]) & (!g802) & (!g1058) & (!g1372) & (keyx82x)) + ((ld) & (!sk[21]) & (!g802) & (!g1058) & (g1372) & (!keyx82x)) + ((ld) & (!sk[21]) & (!g802) & (!g1058) & (g1372) & (keyx82x)) + ((ld) & (!sk[21]) & (!g802) & (g1058) & (!g1372) & (!keyx82x)) + ((ld) & (!sk[21]) & (!g802) & (g1058) & (!g1372) & (keyx82x)) + ((ld) & (!sk[21]) & (!g802) & (g1058) & (g1372) & (!keyx82x)) + ((ld) & (!sk[21]) & (!g802) & (g1058) & (g1372) & (keyx82x)) + ((ld) & (!sk[21]) & (g802) & (!g1058) & (!g1372) & (!keyx82x)) + ((ld) & (!sk[21]) & (g802) & (!g1058) & (!g1372) & (keyx82x)) + ((ld) & (!sk[21]) & (g802) & (!g1058) & (g1372) & (!keyx82x)) + ((ld) & (!sk[21]) & (g802) & (!g1058) & (g1372) & (keyx82x)) + ((ld) & (!sk[21]) & (g802) & (g1058) & (!g1372) & (!keyx82x)) + ((ld) & (!sk[21]) & (g802) & (g1058) & (!g1372) & (keyx82x)) + ((ld) & (!sk[21]) & (g802) & (g1058) & (g1372) & (!keyx82x)) + ((ld) & (!sk[21]) & (g802) & (g1058) & (g1372) & (keyx82x)) + ((ld) & (sk[21]) & (!g802) & (!g1058) & (!g1372) & (keyx82x)) + ((ld) & (sk[21]) & (!g802) & (!g1058) & (g1372) & (keyx82x)) + ((ld) & (sk[21]) & (!g802) & (g1058) & (!g1372) & (keyx82x)) + ((ld) & (sk[21]) & (!g802) & (g1058) & (g1372) & (keyx82x)) + ((ld) & (sk[21]) & (g802) & (!g1058) & (!g1372) & (keyx82x)) + ((ld) & (sk[21]) & (g802) & (!g1058) & (g1372) & (keyx82x)) + ((ld) & (sk[21]) & (g802) & (g1058) & (!g1372) & (keyx82x)) + ((ld) & (sk[21]) & (g802) & (g1058) & (g1372) & (keyx82x)));
	assign g1701 = (((!ld) & (!g809) & (!g1065) & (g1379) & (sk[22]) & (!keyx83x)) + ((!ld) & (!g809) & (!g1065) & (g1379) & (sk[22]) & (keyx83x)) + ((!ld) & (!g809) & (g1065) & (!g1379) & (sk[22]) & (!keyx83x)) + ((!ld) & (!g809) & (g1065) & (!g1379) & (sk[22]) & (keyx83x)) + ((!ld) & (g809) & (!g1065) & (!g1379) & (!sk[22]) & (!keyx83x)) + ((!ld) & (g809) & (!g1065) & (!g1379) & (!sk[22]) & (keyx83x)) + ((!ld) & (g809) & (!g1065) & (!g1379) & (sk[22]) & (!keyx83x)) + ((!ld) & (g809) & (!g1065) & (!g1379) & (sk[22]) & (keyx83x)) + ((!ld) & (g809) & (!g1065) & (g1379) & (!sk[22]) & (!keyx83x)) + ((!ld) & (g809) & (!g1065) & (g1379) & (!sk[22]) & (keyx83x)) + ((!ld) & (g809) & (g1065) & (!g1379) & (!sk[22]) & (!keyx83x)) + ((!ld) & (g809) & (g1065) & (!g1379) & (!sk[22]) & (keyx83x)) + ((!ld) & (g809) & (g1065) & (g1379) & (!sk[22]) & (!keyx83x)) + ((!ld) & (g809) & (g1065) & (g1379) & (!sk[22]) & (keyx83x)) + ((!ld) & (g809) & (g1065) & (g1379) & (sk[22]) & (!keyx83x)) + ((!ld) & (g809) & (g1065) & (g1379) & (sk[22]) & (keyx83x)) + ((ld) & (!g809) & (!g1065) & (!g1379) & (!sk[22]) & (!keyx83x)) + ((ld) & (!g809) & (!g1065) & (!g1379) & (!sk[22]) & (keyx83x)) + ((ld) & (!g809) & (!g1065) & (!g1379) & (sk[22]) & (keyx83x)) + ((ld) & (!g809) & (!g1065) & (g1379) & (!sk[22]) & (!keyx83x)) + ((ld) & (!g809) & (!g1065) & (g1379) & (!sk[22]) & (keyx83x)) + ((ld) & (!g809) & (!g1065) & (g1379) & (sk[22]) & (keyx83x)) + ((ld) & (!g809) & (g1065) & (!g1379) & (!sk[22]) & (!keyx83x)) + ((ld) & (!g809) & (g1065) & (!g1379) & (!sk[22]) & (keyx83x)) + ((ld) & (!g809) & (g1065) & (!g1379) & (sk[22]) & (keyx83x)) + ((ld) & (!g809) & (g1065) & (g1379) & (!sk[22]) & (!keyx83x)) + ((ld) & (!g809) & (g1065) & (g1379) & (!sk[22]) & (keyx83x)) + ((ld) & (!g809) & (g1065) & (g1379) & (sk[22]) & (keyx83x)) + ((ld) & (g809) & (!g1065) & (!g1379) & (!sk[22]) & (!keyx83x)) + ((ld) & (g809) & (!g1065) & (!g1379) & (!sk[22]) & (keyx83x)) + ((ld) & (g809) & (!g1065) & (!g1379) & (sk[22]) & (keyx83x)) + ((ld) & (g809) & (!g1065) & (g1379) & (!sk[22]) & (!keyx83x)) + ((ld) & (g809) & (!g1065) & (g1379) & (!sk[22]) & (keyx83x)) + ((ld) & (g809) & (!g1065) & (g1379) & (sk[22]) & (keyx83x)) + ((ld) & (g809) & (g1065) & (!g1379) & (!sk[22]) & (!keyx83x)) + ((ld) & (g809) & (g1065) & (!g1379) & (!sk[22]) & (keyx83x)) + ((ld) & (g809) & (g1065) & (!g1379) & (sk[22]) & (keyx83x)) + ((ld) & (g809) & (g1065) & (g1379) & (!sk[22]) & (!keyx83x)) + ((ld) & (g809) & (g1065) & (g1379) & (!sk[22]) & (keyx83x)) + ((ld) & (g809) & (g1065) & (g1379) & (sk[22]) & (keyx83x)));
	assign g1702 = (((!ld) & (!sk[23]) & (g816) & (!g1072) & (!g1386) & (!keyx84x)) + ((!ld) & (!sk[23]) & (g816) & (!g1072) & (!g1386) & (keyx84x)) + ((!ld) & (!sk[23]) & (g816) & (!g1072) & (g1386) & (!keyx84x)) + ((!ld) & (!sk[23]) & (g816) & (!g1072) & (g1386) & (keyx84x)) + ((!ld) & (!sk[23]) & (g816) & (g1072) & (!g1386) & (!keyx84x)) + ((!ld) & (!sk[23]) & (g816) & (g1072) & (!g1386) & (keyx84x)) + ((!ld) & (!sk[23]) & (g816) & (g1072) & (g1386) & (!keyx84x)) + ((!ld) & (!sk[23]) & (g816) & (g1072) & (g1386) & (keyx84x)) + ((!ld) & (sk[23]) & (!g816) & (!g1072) & (g1386) & (!keyx84x)) + ((!ld) & (sk[23]) & (!g816) & (!g1072) & (g1386) & (keyx84x)) + ((!ld) & (sk[23]) & (!g816) & (g1072) & (!g1386) & (!keyx84x)) + ((!ld) & (sk[23]) & (!g816) & (g1072) & (!g1386) & (keyx84x)) + ((!ld) & (sk[23]) & (g816) & (!g1072) & (!g1386) & (!keyx84x)) + ((!ld) & (sk[23]) & (g816) & (!g1072) & (!g1386) & (keyx84x)) + ((!ld) & (sk[23]) & (g816) & (g1072) & (g1386) & (!keyx84x)) + ((!ld) & (sk[23]) & (g816) & (g1072) & (g1386) & (keyx84x)) + ((ld) & (!sk[23]) & (!g816) & (!g1072) & (!g1386) & (!keyx84x)) + ((ld) & (!sk[23]) & (!g816) & (!g1072) & (!g1386) & (keyx84x)) + ((ld) & (!sk[23]) & (!g816) & (!g1072) & (g1386) & (!keyx84x)) + ((ld) & (!sk[23]) & (!g816) & (!g1072) & (g1386) & (keyx84x)) + ((ld) & (!sk[23]) & (!g816) & (g1072) & (!g1386) & (!keyx84x)) + ((ld) & (!sk[23]) & (!g816) & (g1072) & (!g1386) & (keyx84x)) + ((ld) & (!sk[23]) & (!g816) & (g1072) & (g1386) & (!keyx84x)) + ((ld) & (!sk[23]) & (!g816) & (g1072) & (g1386) & (keyx84x)) + ((ld) & (!sk[23]) & (g816) & (!g1072) & (!g1386) & (!keyx84x)) + ((ld) & (!sk[23]) & (g816) & (!g1072) & (!g1386) & (keyx84x)) + ((ld) & (!sk[23]) & (g816) & (!g1072) & (g1386) & (!keyx84x)) + ((ld) & (!sk[23]) & (g816) & (!g1072) & (g1386) & (keyx84x)) + ((ld) & (!sk[23]) & (g816) & (g1072) & (!g1386) & (!keyx84x)) + ((ld) & (!sk[23]) & (g816) & (g1072) & (!g1386) & (keyx84x)) + ((ld) & (!sk[23]) & (g816) & (g1072) & (g1386) & (!keyx84x)) + ((ld) & (!sk[23]) & (g816) & (g1072) & (g1386) & (keyx84x)) + ((ld) & (sk[23]) & (!g816) & (!g1072) & (!g1386) & (keyx84x)) + ((ld) & (sk[23]) & (!g816) & (!g1072) & (g1386) & (keyx84x)) + ((ld) & (sk[23]) & (!g816) & (g1072) & (!g1386) & (keyx84x)) + ((ld) & (sk[23]) & (!g816) & (g1072) & (g1386) & (keyx84x)) + ((ld) & (sk[23]) & (g816) & (!g1072) & (!g1386) & (keyx84x)) + ((ld) & (sk[23]) & (g816) & (!g1072) & (g1386) & (keyx84x)) + ((ld) & (sk[23]) & (g816) & (g1072) & (!g1386) & (keyx84x)) + ((ld) & (sk[23]) & (g816) & (g1072) & (g1386) & (keyx84x)));
	assign g1703 = (((!ld) & (!g823) & (!g1079) & (g1393) & (sk[24]) & (!keyx85x)) + ((!ld) & (!g823) & (!g1079) & (g1393) & (sk[24]) & (keyx85x)) + ((!ld) & (!g823) & (g1079) & (!g1393) & (sk[24]) & (!keyx85x)) + ((!ld) & (!g823) & (g1079) & (!g1393) & (sk[24]) & (keyx85x)) + ((!ld) & (g823) & (!g1079) & (!g1393) & (!sk[24]) & (!keyx85x)) + ((!ld) & (g823) & (!g1079) & (!g1393) & (!sk[24]) & (keyx85x)) + ((!ld) & (g823) & (!g1079) & (!g1393) & (sk[24]) & (!keyx85x)) + ((!ld) & (g823) & (!g1079) & (!g1393) & (sk[24]) & (keyx85x)) + ((!ld) & (g823) & (!g1079) & (g1393) & (!sk[24]) & (!keyx85x)) + ((!ld) & (g823) & (!g1079) & (g1393) & (!sk[24]) & (keyx85x)) + ((!ld) & (g823) & (g1079) & (!g1393) & (!sk[24]) & (!keyx85x)) + ((!ld) & (g823) & (g1079) & (!g1393) & (!sk[24]) & (keyx85x)) + ((!ld) & (g823) & (g1079) & (g1393) & (!sk[24]) & (!keyx85x)) + ((!ld) & (g823) & (g1079) & (g1393) & (!sk[24]) & (keyx85x)) + ((!ld) & (g823) & (g1079) & (g1393) & (sk[24]) & (!keyx85x)) + ((!ld) & (g823) & (g1079) & (g1393) & (sk[24]) & (keyx85x)) + ((ld) & (!g823) & (!g1079) & (!g1393) & (!sk[24]) & (!keyx85x)) + ((ld) & (!g823) & (!g1079) & (!g1393) & (!sk[24]) & (keyx85x)) + ((ld) & (!g823) & (!g1079) & (!g1393) & (sk[24]) & (keyx85x)) + ((ld) & (!g823) & (!g1079) & (g1393) & (!sk[24]) & (!keyx85x)) + ((ld) & (!g823) & (!g1079) & (g1393) & (!sk[24]) & (keyx85x)) + ((ld) & (!g823) & (!g1079) & (g1393) & (sk[24]) & (keyx85x)) + ((ld) & (!g823) & (g1079) & (!g1393) & (!sk[24]) & (!keyx85x)) + ((ld) & (!g823) & (g1079) & (!g1393) & (!sk[24]) & (keyx85x)) + ((ld) & (!g823) & (g1079) & (!g1393) & (sk[24]) & (keyx85x)) + ((ld) & (!g823) & (g1079) & (g1393) & (!sk[24]) & (!keyx85x)) + ((ld) & (!g823) & (g1079) & (g1393) & (!sk[24]) & (keyx85x)) + ((ld) & (!g823) & (g1079) & (g1393) & (sk[24]) & (keyx85x)) + ((ld) & (g823) & (!g1079) & (!g1393) & (!sk[24]) & (!keyx85x)) + ((ld) & (g823) & (!g1079) & (!g1393) & (!sk[24]) & (keyx85x)) + ((ld) & (g823) & (!g1079) & (!g1393) & (sk[24]) & (keyx85x)) + ((ld) & (g823) & (!g1079) & (g1393) & (!sk[24]) & (!keyx85x)) + ((ld) & (g823) & (!g1079) & (g1393) & (!sk[24]) & (keyx85x)) + ((ld) & (g823) & (!g1079) & (g1393) & (sk[24]) & (keyx85x)) + ((ld) & (g823) & (g1079) & (!g1393) & (!sk[24]) & (!keyx85x)) + ((ld) & (g823) & (g1079) & (!g1393) & (!sk[24]) & (keyx85x)) + ((ld) & (g823) & (g1079) & (!g1393) & (sk[24]) & (keyx85x)) + ((ld) & (g823) & (g1079) & (g1393) & (!sk[24]) & (!keyx85x)) + ((ld) & (g823) & (g1079) & (g1393) & (!sk[24]) & (keyx85x)) + ((ld) & (g823) & (g1079) & (g1393) & (sk[24]) & (keyx85x)));
	assign g1704 = (((!ld) & (!g830) & (!g1086) & (g1400) & (sk[25]) & (!keyx86x)) + ((!ld) & (!g830) & (!g1086) & (g1400) & (sk[25]) & (keyx86x)) + ((!ld) & (!g830) & (g1086) & (!g1400) & (sk[25]) & (!keyx86x)) + ((!ld) & (!g830) & (g1086) & (!g1400) & (sk[25]) & (keyx86x)) + ((!ld) & (g830) & (!g1086) & (!g1400) & (!sk[25]) & (!keyx86x)) + ((!ld) & (g830) & (!g1086) & (!g1400) & (!sk[25]) & (keyx86x)) + ((!ld) & (g830) & (!g1086) & (!g1400) & (sk[25]) & (!keyx86x)) + ((!ld) & (g830) & (!g1086) & (!g1400) & (sk[25]) & (keyx86x)) + ((!ld) & (g830) & (!g1086) & (g1400) & (!sk[25]) & (!keyx86x)) + ((!ld) & (g830) & (!g1086) & (g1400) & (!sk[25]) & (keyx86x)) + ((!ld) & (g830) & (g1086) & (!g1400) & (!sk[25]) & (!keyx86x)) + ((!ld) & (g830) & (g1086) & (!g1400) & (!sk[25]) & (keyx86x)) + ((!ld) & (g830) & (g1086) & (g1400) & (!sk[25]) & (!keyx86x)) + ((!ld) & (g830) & (g1086) & (g1400) & (!sk[25]) & (keyx86x)) + ((!ld) & (g830) & (g1086) & (g1400) & (sk[25]) & (!keyx86x)) + ((!ld) & (g830) & (g1086) & (g1400) & (sk[25]) & (keyx86x)) + ((ld) & (!g830) & (!g1086) & (!g1400) & (!sk[25]) & (!keyx86x)) + ((ld) & (!g830) & (!g1086) & (!g1400) & (!sk[25]) & (keyx86x)) + ((ld) & (!g830) & (!g1086) & (!g1400) & (sk[25]) & (keyx86x)) + ((ld) & (!g830) & (!g1086) & (g1400) & (!sk[25]) & (!keyx86x)) + ((ld) & (!g830) & (!g1086) & (g1400) & (!sk[25]) & (keyx86x)) + ((ld) & (!g830) & (!g1086) & (g1400) & (sk[25]) & (keyx86x)) + ((ld) & (!g830) & (g1086) & (!g1400) & (!sk[25]) & (!keyx86x)) + ((ld) & (!g830) & (g1086) & (!g1400) & (!sk[25]) & (keyx86x)) + ((ld) & (!g830) & (g1086) & (!g1400) & (sk[25]) & (keyx86x)) + ((ld) & (!g830) & (g1086) & (g1400) & (!sk[25]) & (!keyx86x)) + ((ld) & (!g830) & (g1086) & (g1400) & (!sk[25]) & (keyx86x)) + ((ld) & (!g830) & (g1086) & (g1400) & (sk[25]) & (keyx86x)) + ((ld) & (g830) & (!g1086) & (!g1400) & (!sk[25]) & (!keyx86x)) + ((ld) & (g830) & (!g1086) & (!g1400) & (!sk[25]) & (keyx86x)) + ((ld) & (g830) & (!g1086) & (!g1400) & (sk[25]) & (keyx86x)) + ((ld) & (g830) & (!g1086) & (g1400) & (!sk[25]) & (!keyx86x)) + ((ld) & (g830) & (!g1086) & (g1400) & (!sk[25]) & (keyx86x)) + ((ld) & (g830) & (!g1086) & (g1400) & (sk[25]) & (keyx86x)) + ((ld) & (g830) & (g1086) & (!g1400) & (!sk[25]) & (!keyx86x)) + ((ld) & (g830) & (g1086) & (!g1400) & (!sk[25]) & (keyx86x)) + ((ld) & (g830) & (g1086) & (!g1400) & (sk[25]) & (keyx86x)) + ((ld) & (g830) & (g1086) & (g1400) & (!sk[25]) & (!keyx86x)) + ((ld) & (g830) & (g1086) & (g1400) & (!sk[25]) & (keyx86x)) + ((ld) & (g830) & (g1086) & (g1400) & (sk[25]) & (keyx86x)));
	assign g1705 = (((!ld) & (!g837) & (!g1093) & (sk[26]) & (g1407) & (!keyx87x)) + ((!ld) & (!g837) & (!g1093) & (sk[26]) & (g1407) & (keyx87x)) + ((!ld) & (!g837) & (g1093) & (sk[26]) & (!g1407) & (!keyx87x)) + ((!ld) & (!g837) & (g1093) & (sk[26]) & (!g1407) & (keyx87x)) + ((!ld) & (g837) & (!g1093) & (!sk[26]) & (!g1407) & (!keyx87x)) + ((!ld) & (g837) & (!g1093) & (!sk[26]) & (!g1407) & (keyx87x)) + ((!ld) & (g837) & (!g1093) & (!sk[26]) & (g1407) & (!keyx87x)) + ((!ld) & (g837) & (!g1093) & (!sk[26]) & (g1407) & (keyx87x)) + ((!ld) & (g837) & (!g1093) & (sk[26]) & (!g1407) & (!keyx87x)) + ((!ld) & (g837) & (!g1093) & (sk[26]) & (!g1407) & (keyx87x)) + ((!ld) & (g837) & (g1093) & (!sk[26]) & (!g1407) & (!keyx87x)) + ((!ld) & (g837) & (g1093) & (!sk[26]) & (!g1407) & (keyx87x)) + ((!ld) & (g837) & (g1093) & (!sk[26]) & (g1407) & (!keyx87x)) + ((!ld) & (g837) & (g1093) & (!sk[26]) & (g1407) & (keyx87x)) + ((!ld) & (g837) & (g1093) & (sk[26]) & (g1407) & (!keyx87x)) + ((!ld) & (g837) & (g1093) & (sk[26]) & (g1407) & (keyx87x)) + ((ld) & (!g837) & (!g1093) & (!sk[26]) & (!g1407) & (!keyx87x)) + ((ld) & (!g837) & (!g1093) & (!sk[26]) & (!g1407) & (keyx87x)) + ((ld) & (!g837) & (!g1093) & (!sk[26]) & (g1407) & (!keyx87x)) + ((ld) & (!g837) & (!g1093) & (!sk[26]) & (g1407) & (keyx87x)) + ((ld) & (!g837) & (!g1093) & (sk[26]) & (!g1407) & (keyx87x)) + ((ld) & (!g837) & (!g1093) & (sk[26]) & (g1407) & (keyx87x)) + ((ld) & (!g837) & (g1093) & (!sk[26]) & (!g1407) & (!keyx87x)) + ((ld) & (!g837) & (g1093) & (!sk[26]) & (!g1407) & (keyx87x)) + ((ld) & (!g837) & (g1093) & (!sk[26]) & (g1407) & (!keyx87x)) + ((ld) & (!g837) & (g1093) & (!sk[26]) & (g1407) & (keyx87x)) + ((ld) & (!g837) & (g1093) & (sk[26]) & (!g1407) & (keyx87x)) + ((ld) & (!g837) & (g1093) & (sk[26]) & (g1407) & (keyx87x)) + ((ld) & (g837) & (!g1093) & (!sk[26]) & (!g1407) & (!keyx87x)) + ((ld) & (g837) & (!g1093) & (!sk[26]) & (!g1407) & (keyx87x)) + ((ld) & (g837) & (!g1093) & (!sk[26]) & (g1407) & (!keyx87x)) + ((ld) & (g837) & (!g1093) & (!sk[26]) & (g1407) & (keyx87x)) + ((ld) & (g837) & (!g1093) & (sk[26]) & (!g1407) & (keyx87x)) + ((ld) & (g837) & (!g1093) & (sk[26]) & (g1407) & (keyx87x)) + ((ld) & (g837) & (g1093) & (!sk[26]) & (!g1407) & (!keyx87x)) + ((ld) & (g837) & (g1093) & (!sk[26]) & (!g1407) & (keyx87x)) + ((ld) & (g837) & (g1093) & (!sk[26]) & (g1407) & (!keyx87x)) + ((ld) & (g837) & (g1093) & (!sk[26]) & (g1407) & (keyx87x)) + ((ld) & (g837) & (g1093) & (sk[26]) & (!g1407) & (keyx87x)) + ((ld) & (g837) & (g1093) & (sk[26]) & (g1407) & (keyx87x)));
	assign g2170 = (((!ld) & (!sk[27]) & (text_inx88x) & (!g1706)) + ((!ld) & (!sk[27]) & (text_inx88x) & (g1706)) + ((!ld) & (sk[27]) & (!text_inx88x) & (g1706)) + ((!ld) & (sk[27]) & (text_inx88x) & (g1706)) + ((ld) & (!sk[27]) & (!text_inx88x) & (g1706)) + ((ld) & (!sk[27]) & (text_inx88x) & (!g1706)) + ((ld) & (!sk[27]) & (text_inx88x) & (g1706)) + ((ld) & (sk[27]) & (text_inx88x) & (!g1706)) + ((ld) & (sk[27]) & (text_inx88x) & (g1706)));
	assign g1707 = (((!sk[28]) & (!g787) & (g836) & (!g900)) + ((!sk[28]) & (!g787) & (g836) & (g900)) + ((!sk[28]) & (g787) & (!g836) & (g900)) + ((!sk[28]) & (g787) & (g836) & (!g900)) + ((!sk[28]) & (g787) & (g836) & (g900)) + ((sk[28]) & (!g787) & (!g836) & (g900)) + ((sk[28]) & (!g787) & (g836) & (!g900)) + ((sk[28]) & (g787) & (!g836) & (!g900)) + ((sk[28]) & (g787) & (g836) & (g900)));
	assign g1708 = (((!g659) & (!g723) & (!g852) & (!g1163) & (!g1706) & (g1707)) + ((!g659) & (!g723) & (!g852) & (!g1163) & (g1706) & (g1707)) + ((!g659) & (!g723) & (!g852) & (g1163) & (g1706) & (!g1707)) + ((!g659) & (!g723) & (!g852) & (g1163) & (g1706) & (g1707)) + ((!g659) & (!g723) & (g852) & (!g1163) & (!g1706) & (!g1707)) + ((!g659) & (!g723) & (g852) & (!g1163) & (g1706) & (!g1707)) + ((!g659) & (!g723) & (g852) & (g1163) & (!g1706) & (!g1707)) + ((!g659) & (!g723) & (g852) & (g1163) & (!g1706) & (g1707)) + ((!g659) & (g723) & (!g852) & (!g1163) & (!g1706) & (!g1707)) + ((!g659) & (g723) & (!g852) & (!g1163) & (g1706) & (!g1707)) + ((!g659) & (g723) & (!g852) & (g1163) & (g1706) & (!g1707)) + ((!g659) & (g723) & (!g852) & (g1163) & (g1706) & (g1707)) + ((!g659) & (g723) & (g852) & (!g1163) & (!g1706) & (g1707)) + ((!g659) & (g723) & (g852) & (!g1163) & (g1706) & (g1707)) + ((!g659) & (g723) & (g852) & (g1163) & (!g1706) & (!g1707)) + ((!g659) & (g723) & (g852) & (g1163) & (!g1706) & (g1707)) + ((g659) & (!g723) & (!g852) & (!g1163) & (!g1706) & (!g1707)) + ((g659) & (!g723) & (!g852) & (!g1163) & (g1706) & (!g1707)) + ((g659) & (!g723) & (!g852) & (g1163) & (g1706) & (!g1707)) + ((g659) & (!g723) & (!g852) & (g1163) & (g1706) & (g1707)) + ((g659) & (!g723) & (g852) & (!g1163) & (!g1706) & (g1707)) + ((g659) & (!g723) & (g852) & (!g1163) & (g1706) & (g1707)) + ((g659) & (!g723) & (g852) & (g1163) & (!g1706) & (!g1707)) + ((g659) & (!g723) & (g852) & (g1163) & (!g1706) & (g1707)) + ((g659) & (g723) & (!g852) & (!g1163) & (!g1706) & (g1707)) + ((g659) & (g723) & (!g852) & (!g1163) & (g1706) & (g1707)) + ((g659) & (g723) & (!g852) & (g1163) & (g1706) & (!g1707)) + ((g659) & (g723) & (!g852) & (g1163) & (g1706) & (g1707)) + ((g659) & (g723) & (g852) & (!g1163) & (!g1706) & (!g1707)) + ((g659) & (g723) & (g852) & (!g1163) & (g1706) & (!g1707)) + ((g659) & (g723) & (g852) & (g1163) & (!g1706) & (!g1707)) + ((g659) & (g723) & (g852) & (g1163) & (!g1706) & (g1707)));
	assign g2171 = (((!ld) & (!text_inx89x) & (sk[30]) & (g1709)) + ((!ld) & (text_inx89x) & (!sk[30]) & (!g1709)) + ((!ld) & (text_inx89x) & (!sk[30]) & (g1709)) + ((!ld) & (text_inx89x) & (sk[30]) & (g1709)) + ((ld) & (!text_inx89x) & (!sk[30]) & (g1709)) + ((ld) & (text_inx89x) & (!sk[30]) & (!g1709)) + ((ld) & (text_inx89x) & (!sk[30]) & (g1709)) + ((ld) & (text_inx89x) & (sk[30]) & (!g1709)) + ((ld) & (text_inx89x) & (sk[30]) & (g1709)));
	assign g1710 = (((!sk[31]) & (!g666) & (g730) & (!g794) & (!g851) & (!g859)) + ((!sk[31]) & (!g666) & (g730) & (!g794) & (!g851) & (g859)) + ((!sk[31]) & (!g666) & (g730) & (!g794) & (g851) & (!g859)) + ((!sk[31]) & (!g666) & (g730) & (!g794) & (g851) & (g859)) + ((!sk[31]) & (!g666) & (g730) & (g794) & (!g851) & (!g859)) + ((!sk[31]) & (!g666) & (g730) & (g794) & (!g851) & (g859)) + ((!sk[31]) & (!g666) & (g730) & (g794) & (g851) & (!g859)) + ((!sk[31]) & (!g666) & (g730) & (g794) & (g851) & (g859)) + ((!sk[31]) & (g666) & (!g730) & (!g794) & (!g851) & (!g859)) + ((!sk[31]) & (g666) & (!g730) & (!g794) & (!g851) & (g859)) + ((!sk[31]) & (g666) & (!g730) & (!g794) & (g851) & (!g859)) + ((!sk[31]) & (g666) & (!g730) & (!g794) & (g851) & (g859)) + ((!sk[31]) & (g666) & (!g730) & (g794) & (!g851) & (!g859)) + ((!sk[31]) & (g666) & (!g730) & (g794) & (!g851) & (g859)) + ((!sk[31]) & (g666) & (!g730) & (g794) & (g851) & (!g859)) + ((!sk[31]) & (g666) & (!g730) & (g794) & (g851) & (g859)) + ((!sk[31]) & (g666) & (g730) & (!g794) & (!g851) & (!g859)) + ((!sk[31]) & (g666) & (g730) & (!g794) & (!g851) & (g859)) + ((!sk[31]) & (g666) & (g730) & (!g794) & (g851) & (!g859)) + ((!sk[31]) & (g666) & (g730) & (!g794) & (g851) & (g859)) + ((!sk[31]) & (g666) & (g730) & (g794) & (!g851) & (!g859)) + ((!sk[31]) & (g666) & (g730) & (g794) & (!g851) & (g859)) + ((!sk[31]) & (g666) & (g730) & (g794) & (g851) & (!g859)) + ((!sk[31]) & (g666) & (g730) & (g794) & (g851) & (g859)) + ((sk[31]) & (!g666) & (!g730) & (!g794) & (!g851) & (g859)) + ((sk[31]) & (!g666) & (!g730) & (!g794) & (g851) & (!g859)) + ((sk[31]) & (!g666) & (!g730) & (g794) & (!g851) & (!g859)) + ((sk[31]) & (!g666) & (!g730) & (g794) & (g851) & (g859)) + ((sk[31]) & (!g666) & (g730) & (!g794) & (!g851) & (!g859)) + ((sk[31]) & (!g666) & (g730) & (!g794) & (g851) & (g859)) + ((sk[31]) & (!g666) & (g730) & (g794) & (!g851) & (g859)) + ((sk[31]) & (!g666) & (g730) & (g794) & (g851) & (!g859)) + ((sk[31]) & (g666) & (!g730) & (!g794) & (!g851) & (!g859)) + ((sk[31]) & (g666) & (!g730) & (!g794) & (g851) & (g859)) + ((sk[31]) & (g666) & (!g730) & (g794) & (!g851) & (g859)) + ((sk[31]) & (g666) & (!g730) & (g794) & (g851) & (!g859)) + ((sk[31]) & (g666) & (g730) & (!g794) & (!g851) & (g859)) + ((sk[31]) & (g666) & (g730) & (!g794) & (g851) & (!g859)) + ((sk[31]) & (g666) & (g730) & (g794) & (!g851) & (!g859)) + ((sk[31]) & (g666) & (g730) & (g794) & (g851) & (g859)));
	assign g1711 = (((!g859) & (!g1163) & (!g1707) & (!g1709) & (sk[32]) & (g1710)) + ((!g859) & (!g1163) & (!g1707) & (g1709) & (sk[32]) & (g1710)) + ((!g859) & (!g1163) & (g1707) & (!g1709) & (sk[32]) & (!g1710)) + ((!g859) & (!g1163) & (g1707) & (g1709) & (sk[32]) & (!g1710)) + ((!g859) & (g1163) & (!g1707) & (!g1709) & (!sk[32]) & (!g1710)) + ((!g859) & (g1163) & (!g1707) & (!g1709) & (!sk[32]) & (g1710)) + ((!g859) & (g1163) & (!g1707) & (g1709) & (!sk[32]) & (!g1710)) + ((!g859) & (g1163) & (!g1707) & (g1709) & (!sk[32]) & (g1710)) + ((!g859) & (g1163) & (!g1707) & (g1709) & (sk[32]) & (!g1710)) + ((!g859) & (g1163) & (!g1707) & (g1709) & (sk[32]) & (g1710)) + ((!g859) & (g1163) & (g1707) & (!g1709) & (!sk[32]) & (!g1710)) + ((!g859) & (g1163) & (g1707) & (!g1709) & (!sk[32]) & (g1710)) + ((!g859) & (g1163) & (g1707) & (g1709) & (!sk[32]) & (!g1710)) + ((!g859) & (g1163) & (g1707) & (g1709) & (!sk[32]) & (g1710)) + ((!g859) & (g1163) & (g1707) & (g1709) & (sk[32]) & (!g1710)) + ((!g859) & (g1163) & (g1707) & (g1709) & (sk[32]) & (g1710)) + ((g859) & (!g1163) & (!g1707) & (!g1709) & (!sk[32]) & (!g1710)) + ((g859) & (!g1163) & (!g1707) & (!g1709) & (!sk[32]) & (g1710)) + ((g859) & (!g1163) & (!g1707) & (!g1709) & (sk[32]) & (g1710)) + ((g859) & (!g1163) & (!g1707) & (g1709) & (!sk[32]) & (!g1710)) + ((g859) & (!g1163) & (!g1707) & (g1709) & (!sk[32]) & (g1710)) + ((g859) & (!g1163) & (!g1707) & (g1709) & (sk[32]) & (g1710)) + ((g859) & (!g1163) & (g1707) & (!g1709) & (!sk[32]) & (!g1710)) + ((g859) & (!g1163) & (g1707) & (!g1709) & (!sk[32]) & (g1710)) + ((g859) & (!g1163) & (g1707) & (!g1709) & (sk[32]) & (!g1710)) + ((g859) & (!g1163) & (g1707) & (g1709) & (!sk[32]) & (!g1710)) + ((g859) & (!g1163) & (g1707) & (g1709) & (!sk[32]) & (g1710)) + ((g859) & (!g1163) & (g1707) & (g1709) & (sk[32]) & (!g1710)) + ((g859) & (g1163) & (!g1707) & (!g1709) & (!sk[32]) & (!g1710)) + ((g859) & (g1163) & (!g1707) & (!g1709) & (!sk[32]) & (g1710)) + ((g859) & (g1163) & (!g1707) & (!g1709) & (sk[32]) & (!g1710)) + ((g859) & (g1163) & (!g1707) & (!g1709) & (sk[32]) & (g1710)) + ((g859) & (g1163) & (!g1707) & (g1709) & (!sk[32]) & (!g1710)) + ((g859) & (g1163) & (!g1707) & (g1709) & (!sk[32]) & (g1710)) + ((g859) & (g1163) & (g1707) & (!g1709) & (!sk[32]) & (!g1710)) + ((g859) & (g1163) & (g1707) & (!g1709) & (!sk[32]) & (g1710)) + ((g859) & (g1163) & (g1707) & (!g1709) & (sk[32]) & (!g1710)) + ((g859) & (g1163) & (g1707) & (!g1709) & (sk[32]) & (g1710)) + ((g859) & (g1163) & (g1707) & (g1709) & (!sk[32]) & (!g1710)) + ((g859) & (g1163) & (g1707) & (g1709) & (!sk[32]) & (g1710)));
	assign g2172 = (((!sk[33]) & (!ld) & (text_inx90x) & (!g1712)) + ((!sk[33]) & (!ld) & (text_inx90x) & (g1712)) + ((!sk[33]) & (ld) & (!text_inx90x) & (g1712)) + ((!sk[33]) & (ld) & (text_inx90x) & (!g1712)) + ((!sk[33]) & (ld) & (text_inx90x) & (g1712)) + ((sk[33]) & (!ld) & (!text_inx90x) & (g1712)) + ((sk[33]) & (!ld) & (text_inx90x) & (g1712)) + ((sk[33]) & (ld) & (text_inx90x) & (!g1712)) + ((sk[33]) & (ld) & (text_inx90x) & (g1712)));
	assign g1713 = (((!g673) & (!g737) & (sk[34]) & (g794)) + ((!g673) & (g737) & (!sk[34]) & (!g794)) + ((!g673) & (g737) & (!sk[34]) & (g794)) + ((!g673) & (g737) & (sk[34]) & (!g794)) + ((g673) & (!g737) & (!sk[34]) & (g794)) + ((g673) & (!g737) & (sk[34]) & (!g794)) + ((g673) & (g737) & (!sk[34]) & (!g794)) + ((g673) & (g737) & (!sk[34]) & (g794)) + ((g673) & (g737) & (sk[34]) & (g794)));
	assign g1714 = (((!g801) & (!g858) & (!g866) & (!g1163) & (!g1712) & (g1713)) + ((!g801) & (!g858) & (!g866) & (!g1163) & (g1712) & (g1713)) + ((!g801) & (!g858) & (!g866) & (g1163) & (g1712) & (!g1713)) + ((!g801) & (!g858) & (!g866) & (g1163) & (g1712) & (g1713)) + ((!g801) & (!g858) & (g866) & (!g1163) & (!g1712) & (!g1713)) + ((!g801) & (!g858) & (g866) & (!g1163) & (g1712) & (!g1713)) + ((!g801) & (!g858) & (g866) & (g1163) & (!g1712) & (!g1713)) + ((!g801) & (!g858) & (g866) & (g1163) & (!g1712) & (g1713)) + ((!g801) & (g858) & (!g866) & (!g1163) & (!g1712) & (!g1713)) + ((!g801) & (g858) & (!g866) & (!g1163) & (g1712) & (!g1713)) + ((!g801) & (g858) & (!g866) & (g1163) & (g1712) & (!g1713)) + ((!g801) & (g858) & (!g866) & (g1163) & (g1712) & (g1713)) + ((!g801) & (g858) & (g866) & (!g1163) & (!g1712) & (g1713)) + ((!g801) & (g858) & (g866) & (!g1163) & (g1712) & (g1713)) + ((!g801) & (g858) & (g866) & (g1163) & (!g1712) & (!g1713)) + ((!g801) & (g858) & (g866) & (g1163) & (!g1712) & (g1713)) + ((g801) & (!g858) & (!g866) & (!g1163) & (!g1712) & (!g1713)) + ((g801) & (!g858) & (!g866) & (!g1163) & (g1712) & (!g1713)) + ((g801) & (!g858) & (!g866) & (g1163) & (g1712) & (!g1713)) + ((g801) & (!g858) & (!g866) & (g1163) & (g1712) & (g1713)) + ((g801) & (!g858) & (g866) & (!g1163) & (!g1712) & (g1713)) + ((g801) & (!g858) & (g866) & (!g1163) & (g1712) & (g1713)) + ((g801) & (!g858) & (g866) & (g1163) & (!g1712) & (!g1713)) + ((g801) & (!g858) & (g866) & (g1163) & (!g1712) & (g1713)) + ((g801) & (g858) & (!g866) & (!g1163) & (!g1712) & (g1713)) + ((g801) & (g858) & (!g866) & (!g1163) & (g1712) & (g1713)) + ((g801) & (g858) & (!g866) & (g1163) & (g1712) & (!g1713)) + ((g801) & (g858) & (!g866) & (g1163) & (g1712) & (g1713)) + ((g801) & (g858) & (g866) & (!g1163) & (!g1712) & (!g1713)) + ((g801) & (g858) & (g866) & (!g1163) & (g1712) & (!g1713)) + ((g801) & (g858) & (g866) & (g1163) & (!g1712) & (!g1713)) + ((g801) & (g858) & (g866) & (g1163) & (!g1712) & (g1713)));
	assign g2173 = (((!ld) & (!sk[36]) & (text_inx91x) & (!g1715)) + ((!ld) & (!sk[36]) & (text_inx91x) & (g1715)) + ((!ld) & (sk[36]) & (!text_inx91x) & (g1715)) + ((!ld) & (sk[36]) & (text_inx91x) & (g1715)) + ((ld) & (!sk[36]) & (!text_inx91x) & (g1715)) + ((ld) & (!sk[36]) & (text_inx91x) & (!g1715)) + ((ld) & (!sk[36]) & (text_inx91x) & (g1715)) + ((ld) & (sk[36]) & (text_inx91x) & (!g1715)) + ((ld) & (sk[36]) & (text_inx91x) & (g1715)));
	assign g1716 = (((!g801) & (!sk[37]) & (g836)) + ((!g801) & (sk[37]) & (g836)) + ((g801) & (!sk[37]) & (g836)) + ((g801) & (sk[37]) & (!g836)));
	assign g1717 = (((!g680) & (!g873) & (!g1163) & (!g1514) & (!g1715) & (g1716)) + ((!g680) & (!g873) & (!g1163) & (!g1514) & (g1715) & (g1716)) + ((!g680) & (!g873) & (!g1163) & (g1514) & (!g1715) & (!g1716)) + ((!g680) & (!g873) & (!g1163) & (g1514) & (g1715) & (!g1716)) + ((!g680) & (!g873) & (g1163) & (!g1514) & (g1715) & (!g1716)) + ((!g680) & (!g873) & (g1163) & (!g1514) & (g1715) & (g1716)) + ((!g680) & (!g873) & (g1163) & (g1514) & (g1715) & (!g1716)) + ((!g680) & (!g873) & (g1163) & (g1514) & (g1715) & (g1716)) + ((!g680) & (g873) & (!g1163) & (!g1514) & (!g1715) & (!g1716)) + ((!g680) & (g873) & (!g1163) & (!g1514) & (g1715) & (!g1716)) + ((!g680) & (g873) & (!g1163) & (g1514) & (!g1715) & (g1716)) + ((!g680) & (g873) & (!g1163) & (g1514) & (g1715) & (g1716)) + ((!g680) & (g873) & (g1163) & (!g1514) & (!g1715) & (!g1716)) + ((!g680) & (g873) & (g1163) & (!g1514) & (!g1715) & (g1716)) + ((!g680) & (g873) & (g1163) & (g1514) & (!g1715) & (!g1716)) + ((!g680) & (g873) & (g1163) & (g1514) & (!g1715) & (g1716)) + ((g680) & (!g873) & (!g1163) & (!g1514) & (!g1715) & (!g1716)) + ((g680) & (!g873) & (!g1163) & (!g1514) & (g1715) & (!g1716)) + ((g680) & (!g873) & (!g1163) & (g1514) & (!g1715) & (g1716)) + ((g680) & (!g873) & (!g1163) & (g1514) & (g1715) & (g1716)) + ((g680) & (!g873) & (g1163) & (!g1514) & (g1715) & (!g1716)) + ((g680) & (!g873) & (g1163) & (!g1514) & (g1715) & (g1716)) + ((g680) & (!g873) & (g1163) & (g1514) & (g1715) & (!g1716)) + ((g680) & (!g873) & (g1163) & (g1514) & (g1715) & (g1716)) + ((g680) & (g873) & (!g1163) & (!g1514) & (!g1715) & (g1716)) + ((g680) & (g873) & (!g1163) & (!g1514) & (g1715) & (g1716)) + ((g680) & (g873) & (!g1163) & (g1514) & (!g1715) & (!g1716)) + ((g680) & (g873) & (!g1163) & (g1514) & (g1715) & (!g1716)) + ((g680) & (g873) & (g1163) & (!g1514) & (!g1715) & (!g1716)) + ((g680) & (g873) & (g1163) & (!g1514) & (!g1715) & (g1716)) + ((g680) & (g873) & (g1163) & (g1514) & (!g1715) & (!g1716)) + ((g680) & (g873) & (g1163) & (g1514) & (!g1715) & (g1716)));
	assign g2174 = (((!ld) & (!sk[39]) & (text_inx94x) & (!g1718)) + ((!ld) & (!sk[39]) & (text_inx94x) & (g1718)) + ((!ld) & (sk[39]) & (!text_inx94x) & (g1718)) + ((!ld) & (sk[39]) & (text_inx94x) & (g1718)) + ((ld) & (!sk[39]) & (!text_inx94x) & (g1718)) + ((ld) & (!sk[39]) & (text_inx94x) & (!g1718)) + ((ld) & (!sk[39]) & (text_inx94x) & (g1718)) + ((ld) & (sk[39]) & (text_inx94x) & (!g1718)) + ((ld) & (sk[39]) & (text_inx94x) & (g1718)));
	assign g1719 = (((!sk[40]) & (!g701) & (g765) & (!g822)) + ((!sk[40]) & (!g701) & (g765) & (g822)) + ((!sk[40]) & (g701) & (!g765) & (g822)) + ((!sk[40]) & (g701) & (g765) & (!g822)) + ((!sk[40]) & (g701) & (g765) & (g822)) + ((sk[40]) & (!g701) & (!g765) & (g822)) + ((sk[40]) & (!g701) & (g765) & (!g822)) + ((sk[40]) & (g701) & (!g765) & (!g822)) + ((sk[40]) & (g701) & (g765) & (g822)));
	assign g1720 = (((!g829) & (!g886) & (!g894) & (!g1163) & (!g1718) & (g1719)) + ((!g829) & (!g886) & (!g894) & (!g1163) & (g1718) & (g1719)) + ((!g829) & (!g886) & (!g894) & (g1163) & (g1718) & (!g1719)) + ((!g829) & (!g886) & (!g894) & (g1163) & (g1718) & (g1719)) + ((!g829) & (!g886) & (g894) & (!g1163) & (!g1718) & (!g1719)) + ((!g829) & (!g886) & (g894) & (!g1163) & (g1718) & (!g1719)) + ((!g829) & (!g886) & (g894) & (g1163) & (!g1718) & (!g1719)) + ((!g829) & (!g886) & (g894) & (g1163) & (!g1718) & (g1719)) + ((!g829) & (g886) & (!g894) & (!g1163) & (!g1718) & (!g1719)) + ((!g829) & (g886) & (!g894) & (!g1163) & (g1718) & (!g1719)) + ((!g829) & (g886) & (!g894) & (g1163) & (g1718) & (!g1719)) + ((!g829) & (g886) & (!g894) & (g1163) & (g1718) & (g1719)) + ((!g829) & (g886) & (g894) & (!g1163) & (!g1718) & (g1719)) + ((!g829) & (g886) & (g894) & (!g1163) & (g1718) & (g1719)) + ((!g829) & (g886) & (g894) & (g1163) & (!g1718) & (!g1719)) + ((!g829) & (g886) & (g894) & (g1163) & (!g1718) & (g1719)) + ((g829) & (!g886) & (!g894) & (!g1163) & (!g1718) & (!g1719)) + ((g829) & (!g886) & (!g894) & (!g1163) & (g1718) & (!g1719)) + ((g829) & (!g886) & (!g894) & (g1163) & (g1718) & (!g1719)) + ((g829) & (!g886) & (!g894) & (g1163) & (g1718) & (g1719)) + ((g829) & (!g886) & (g894) & (!g1163) & (!g1718) & (g1719)) + ((g829) & (!g886) & (g894) & (!g1163) & (g1718) & (g1719)) + ((g829) & (!g886) & (g894) & (g1163) & (!g1718) & (!g1719)) + ((g829) & (!g886) & (g894) & (g1163) & (!g1718) & (g1719)) + ((g829) & (g886) & (!g894) & (!g1163) & (!g1718) & (g1719)) + ((g829) & (g886) & (!g894) & (!g1163) & (g1718) & (g1719)) + ((g829) & (g886) & (!g894) & (g1163) & (g1718) & (!g1719)) + ((g829) & (g886) & (!g894) & (g1163) & (g1718) & (g1719)) + ((g829) & (g886) & (g894) & (!g1163) & (!g1718) & (!g1719)) + ((g829) & (g886) & (g894) & (!g1163) & (g1718) & (!g1719)) + ((g829) & (g886) & (g894) & (g1163) & (!g1718) & (!g1719)) + ((g829) & (g886) & (g894) & (g1163) & (!g1718) & (g1719)));
	assign g2175 = (((!ld) & (!text_inx93x) & (sk[42]) & (g1721)) + ((!ld) & (text_inx93x) & (!sk[42]) & (!g1721)) + ((!ld) & (text_inx93x) & (!sk[42]) & (g1721)) + ((!ld) & (text_inx93x) & (sk[42]) & (g1721)) + ((ld) & (!text_inx93x) & (!sk[42]) & (g1721)) + ((ld) & (text_inx93x) & (!sk[42]) & (!g1721)) + ((ld) & (text_inx93x) & (!sk[42]) & (g1721)) + ((ld) & (text_inx93x) & (sk[42]) & (!g1721)) + ((ld) & (text_inx93x) & (sk[42]) & (g1721)));
	assign g1722 = (((!g694) & (!sk[43]) & (g758) & (!g815)) + ((!g694) & (!sk[43]) & (g758) & (g815)) + ((!g694) & (sk[43]) & (!g758) & (g815)) + ((!g694) & (sk[43]) & (g758) & (!g815)) + ((g694) & (!sk[43]) & (!g758) & (g815)) + ((g694) & (!sk[43]) & (g758) & (!g815)) + ((g694) & (!sk[43]) & (g758) & (g815)) + ((g694) & (sk[43]) & (!g758) & (!g815)) + ((g694) & (sk[43]) & (g758) & (g815)));
	assign g1723 = (((!g822) & (!g879) & (!g887) & (!g1163) & (!g1721) & (g1722)) + ((!g822) & (!g879) & (!g887) & (!g1163) & (g1721) & (g1722)) + ((!g822) & (!g879) & (!g887) & (g1163) & (g1721) & (!g1722)) + ((!g822) & (!g879) & (!g887) & (g1163) & (g1721) & (g1722)) + ((!g822) & (!g879) & (g887) & (!g1163) & (!g1721) & (!g1722)) + ((!g822) & (!g879) & (g887) & (!g1163) & (g1721) & (!g1722)) + ((!g822) & (!g879) & (g887) & (g1163) & (!g1721) & (!g1722)) + ((!g822) & (!g879) & (g887) & (g1163) & (!g1721) & (g1722)) + ((!g822) & (g879) & (!g887) & (!g1163) & (!g1721) & (!g1722)) + ((!g822) & (g879) & (!g887) & (!g1163) & (g1721) & (!g1722)) + ((!g822) & (g879) & (!g887) & (g1163) & (g1721) & (!g1722)) + ((!g822) & (g879) & (!g887) & (g1163) & (g1721) & (g1722)) + ((!g822) & (g879) & (g887) & (!g1163) & (!g1721) & (g1722)) + ((!g822) & (g879) & (g887) & (!g1163) & (g1721) & (g1722)) + ((!g822) & (g879) & (g887) & (g1163) & (!g1721) & (!g1722)) + ((!g822) & (g879) & (g887) & (g1163) & (!g1721) & (g1722)) + ((g822) & (!g879) & (!g887) & (!g1163) & (!g1721) & (!g1722)) + ((g822) & (!g879) & (!g887) & (!g1163) & (g1721) & (!g1722)) + ((g822) & (!g879) & (!g887) & (g1163) & (g1721) & (!g1722)) + ((g822) & (!g879) & (!g887) & (g1163) & (g1721) & (g1722)) + ((g822) & (!g879) & (g887) & (!g1163) & (!g1721) & (g1722)) + ((g822) & (!g879) & (g887) & (!g1163) & (g1721) & (g1722)) + ((g822) & (!g879) & (g887) & (g1163) & (!g1721) & (!g1722)) + ((g822) & (!g879) & (g887) & (g1163) & (!g1721) & (g1722)) + ((g822) & (g879) & (!g887) & (!g1163) & (!g1721) & (g1722)) + ((g822) & (g879) & (!g887) & (!g1163) & (g1721) & (g1722)) + ((g822) & (g879) & (!g887) & (g1163) & (g1721) & (!g1722)) + ((g822) & (g879) & (!g887) & (g1163) & (g1721) & (g1722)) + ((g822) & (g879) & (g887) & (!g1163) & (!g1721) & (!g1722)) + ((g822) & (g879) & (g887) & (!g1163) & (g1721) & (!g1722)) + ((g822) & (g879) & (g887) & (g1163) & (!g1721) & (!g1722)) + ((g822) & (g879) & (g887) & (g1163) & (!g1721) & (g1722)));
	assign g2176 = (((!sk[45]) & (!ld) & (text_inx92x) & (!g1724)) + ((!sk[45]) & (!ld) & (text_inx92x) & (g1724)) + ((!sk[45]) & (ld) & (!text_inx92x) & (g1724)) + ((!sk[45]) & (ld) & (text_inx92x) & (!g1724)) + ((!sk[45]) & (ld) & (text_inx92x) & (g1724)) + ((sk[45]) & (!ld) & (!text_inx92x) & (g1724)) + ((sk[45]) & (!ld) & (text_inx92x) & (g1724)) + ((sk[45]) & (ld) & (text_inx92x) & (!g1724)) + ((sk[45]) & (ld) & (text_inx92x) & (g1724)));
	assign g1725 = (((!sk[46]) & (!g687) & (g751) & (!g808)) + ((!sk[46]) & (!g687) & (g751) & (g808)) + ((!sk[46]) & (g687) & (!g751) & (g808)) + ((!sk[46]) & (g687) & (g751) & (!g808)) + ((!sk[46]) & (g687) & (g751) & (g808)) + ((sk[46]) & (!g687) & (!g751) & (g808)) + ((sk[46]) & (!g687) & (g751) & (!g808)) + ((sk[46]) & (g687) & (!g751) & (!g808)) + ((sk[46]) & (g687) & (g751) & (g808)));
	assign g1726 = (((!g815) & (!g836) & (!g872) & (sk[47]) & (!g880) & (g900)) + ((!g815) & (!g836) & (!g872) & (sk[47]) & (g880) & (!g900)) + ((!g815) & (!g836) & (g872) & (sk[47]) & (!g880) & (!g900)) + ((!g815) & (!g836) & (g872) & (sk[47]) & (g880) & (g900)) + ((!g815) & (g836) & (!g872) & (!sk[47]) & (!g880) & (!g900)) + ((!g815) & (g836) & (!g872) & (!sk[47]) & (!g880) & (g900)) + ((!g815) & (g836) & (!g872) & (!sk[47]) & (g880) & (!g900)) + ((!g815) & (g836) & (!g872) & (!sk[47]) & (g880) & (g900)) + ((!g815) & (g836) & (!g872) & (sk[47]) & (!g880) & (!g900)) + ((!g815) & (g836) & (!g872) & (sk[47]) & (g880) & (g900)) + ((!g815) & (g836) & (g872) & (!sk[47]) & (!g880) & (!g900)) + ((!g815) & (g836) & (g872) & (!sk[47]) & (!g880) & (g900)) + ((!g815) & (g836) & (g872) & (!sk[47]) & (g880) & (!g900)) + ((!g815) & (g836) & (g872) & (!sk[47]) & (g880) & (g900)) + ((!g815) & (g836) & (g872) & (sk[47]) & (!g880) & (g900)) + ((!g815) & (g836) & (g872) & (sk[47]) & (g880) & (!g900)) + ((g815) & (!g836) & (!g872) & (!sk[47]) & (!g880) & (!g900)) + ((g815) & (!g836) & (!g872) & (!sk[47]) & (!g880) & (g900)) + ((g815) & (!g836) & (!g872) & (!sk[47]) & (g880) & (!g900)) + ((g815) & (!g836) & (!g872) & (!sk[47]) & (g880) & (g900)) + ((g815) & (!g836) & (!g872) & (sk[47]) & (!g880) & (!g900)) + ((g815) & (!g836) & (!g872) & (sk[47]) & (g880) & (g900)) + ((g815) & (!g836) & (g872) & (!sk[47]) & (!g880) & (!g900)) + ((g815) & (!g836) & (g872) & (!sk[47]) & (!g880) & (g900)) + ((g815) & (!g836) & (g872) & (!sk[47]) & (g880) & (!g900)) + ((g815) & (!g836) & (g872) & (!sk[47]) & (g880) & (g900)) + ((g815) & (!g836) & (g872) & (sk[47]) & (!g880) & (g900)) + ((g815) & (!g836) & (g872) & (sk[47]) & (g880) & (!g900)) + ((g815) & (g836) & (!g872) & (!sk[47]) & (!g880) & (!g900)) + ((g815) & (g836) & (!g872) & (!sk[47]) & (!g880) & (g900)) + ((g815) & (g836) & (!g872) & (!sk[47]) & (g880) & (!g900)) + ((g815) & (g836) & (!g872) & (!sk[47]) & (g880) & (g900)) + ((g815) & (g836) & (!g872) & (sk[47]) & (!g880) & (g900)) + ((g815) & (g836) & (!g872) & (sk[47]) & (g880) & (!g900)) + ((g815) & (g836) & (g872) & (!sk[47]) & (!g880) & (!g900)) + ((g815) & (g836) & (g872) & (!sk[47]) & (!g880) & (g900)) + ((g815) & (g836) & (g872) & (!sk[47]) & (g880) & (!g900)) + ((g815) & (g836) & (g872) & (!sk[47]) & (g880) & (g900)) + ((g815) & (g836) & (g872) & (sk[47]) & (!g880) & (!g900)) + ((g815) & (g836) & (g872) & (sk[47]) & (g880) & (g900)));
	assign g1727 = (((!g880) & (!sk[48]) & (g1163) & (!g1724) & (!g1725) & (!g1726)) + ((!g880) & (!sk[48]) & (g1163) & (!g1724) & (!g1725) & (g1726)) + ((!g880) & (!sk[48]) & (g1163) & (!g1724) & (g1725) & (!g1726)) + ((!g880) & (!sk[48]) & (g1163) & (!g1724) & (g1725) & (g1726)) + ((!g880) & (!sk[48]) & (g1163) & (g1724) & (!g1725) & (!g1726)) + ((!g880) & (!sk[48]) & (g1163) & (g1724) & (!g1725) & (g1726)) + ((!g880) & (!sk[48]) & (g1163) & (g1724) & (g1725) & (!g1726)) + ((!g880) & (!sk[48]) & (g1163) & (g1724) & (g1725) & (g1726)) + ((!g880) & (sk[48]) & (!g1163) & (!g1724) & (!g1725) & (g1726)) + ((!g880) & (sk[48]) & (!g1163) & (!g1724) & (g1725) & (!g1726)) + ((!g880) & (sk[48]) & (!g1163) & (g1724) & (!g1725) & (g1726)) + ((!g880) & (sk[48]) & (!g1163) & (g1724) & (g1725) & (!g1726)) + ((!g880) & (sk[48]) & (g1163) & (g1724) & (!g1725) & (!g1726)) + ((!g880) & (sk[48]) & (g1163) & (g1724) & (!g1725) & (g1726)) + ((!g880) & (sk[48]) & (g1163) & (g1724) & (g1725) & (!g1726)) + ((!g880) & (sk[48]) & (g1163) & (g1724) & (g1725) & (g1726)) + ((g880) & (!sk[48]) & (!g1163) & (!g1724) & (!g1725) & (!g1726)) + ((g880) & (!sk[48]) & (!g1163) & (!g1724) & (!g1725) & (g1726)) + ((g880) & (!sk[48]) & (!g1163) & (!g1724) & (g1725) & (!g1726)) + ((g880) & (!sk[48]) & (!g1163) & (!g1724) & (g1725) & (g1726)) + ((g880) & (!sk[48]) & (!g1163) & (g1724) & (!g1725) & (!g1726)) + ((g880) & (!sk[48]) & (!g1163) & (g1724) & (!g1725) & (g1726)) + ((g880) & (!sk[48]) & (!g1163) & (g1724) & (g1725) & (!g1726)) + ((g880) & (!sk[48]) & (!g1163) & (g1724) & (g1725) & (g1726)) + ((g880) & (!sk[48]) & (g1163) & (!g1724) & (!g1725) & (!g1726)) + ((g880) & (!sk[48]) & (g1163) & (!g1724) & (!g1725) & (g1726)) + ((g880) & (!sk[48]) & (g1163) & (!g1724) & (g1725) & (!g1726)) + ((g880) & (!sk[48]) & (g1163) & (!g1724) & (g1725) & (g1726)) + ((g880) & (!sk[48]) & (g1163) & (g1724) & (!g1725) & (!g1726)) + ((g880) & (!sk[48]) & (g1163) & (g1724) & (!g1725) & (g1726)) + ((g880) & (!sk[48]) & (g1163) & (g1724) & (g1725) & (!g1726)) + ((g880) & (!sk[48]) & (g1163) & (g1724) & (g1725) & (g1726)) + ((g880) & (sk[48]) & (!g1163) & (!g1724) & (!g1725) & (g1726)) + ((g880) & (sk[48]) & (!g1163) & (!g1724) & (g1725) & (!g1726)) + ((g880) & (sk[48]) & (!g1163) & (g1724) & (!g1725) & (g1726)) + ((g880) & (sk[48]) & (!g1163) & (g1724) & (g1725) & (!g1726)) + ((g880) & (sk[48]) & (g1163) & (!g1724) & (!g1725) & (!g1726)) + ((g880) & (sk[48]) & (g1163) & (!g1724) & (!g1725) & (g1726)) + ((g880) & (sk[48]) & (g1163) & (!g1724) & (g1725) & (!g1726)) + ((g880) & (sk[48]) & (g1163) & (!g1724) & (g1725) & (g1726)));
	assign g1728 = (((!g829) & (!sk[49]) & (g893)) + ((!g829) & (sk[49]) & (g893)) + ((g829) & (!sk[49]) & (g893)) + ((g829) & (sk[49]) & (!g893)));
	assign g2177 = (((!ld) & (!text_inx95x) & (sk[50]) & (g1729)) + ((!ld) & (text_inx95x) & (!sk[50]) & (!g1729)) + ((!ld) & (text_inx95x) & (!sk[50]) & (g1729)) + ((!ld) & (text_inx95x) & (sk[50]) & (g1729)) + ((ld) & (!text_inx95x) & (!sk[50]) & (g1729)) + ((ld) & (text_inx95x) & (!sk[50]) & (!g1729)) + ((ld) & (text_inx95x) & (!sk[50]) & (g1729)) + ((ld) & (text_inx95x) & (sk[50]) & (!g1729)) + ((ld) & (text_inx95x) & (sk[50]) & (g1729)));
	assign g1730 = (((!g836) & (!g901) & (!g1163) & (!g1246) & (g1728) & (!g1729)) + ((!g836) & (!g901) & (!g1163) & (!g1246) & (g1728) & (g1729)) + ((!g836) & (!g901) & (!g1163) & (g1246) & (!g1728) & (!g1729)) + ((!g836) & (!g901) & (!g1163) & (g1246) & (!g1728) & (g1729)) + ((!g836) & (!g901) & (g1163) & (!g1246) & (!g1728) & (g1729)) + ((!g836) & (!g901) & (g1163) & (!g1246) & (g1728) & (g1729)) + ((!g836) & (!g901) & (g1163) & (g1246) & (!g1728) & (g1729)) + ((!g836) & (!g901) & (g1163) & (g1246) & (g1728) & (g1729)) + ((!g836) & (g901) & (!g1163) & (!g1246) & (!g1728) & (!g1729)) + ((!g836) & (g901) & (!g1163) & (!g1246) & (!g1728) & (g1729)) + ((!g836) & (g901) & (!g1163) & (g1246) & (g1728) & (!g1729)) + ((!g836) & (g901) & (!g1163) & (g1246) & (g1728) & (g1729)) + ((!g836) & (g901) & (g1163) & (!g1246) & (!g1728) & (!g1729)) + ((!g836) & (g901) & (g1163) & (!g1246) & (g1728) & (!g1729)) + ((!g836) & (g901) & (g1163) & (g1246) & (!g1728) & (!g1729)) + ((!g836) & (g901) & (g1163) & (g1246) & (g1728) & (!g1729)) + ((g836) & (!g901) & (!g1163) & (!g1246) & (!g1728) & (!g1729)) + ((g836) & (!g901) & (!g1163) & (!g1246) & (!g1728) & (g1729)) + ((g836) & (!g901) & (!g1163) & (g1246) & (g1728) & (!g1729)) + ((g836) & (!g901) & (!g1163) & (g1246) & (g1728) & (g1729)) + ((g836) & (!g901) & (g1163) & (!g1246) & (!g1728) & (g1729)) + ((g836) & (!g901) & (g1163) & (!g1246) & (g1728) & (g1729)) + ((g836) & (!g901) & (g1163) & (g1246) & (!g1728) & (g1729)) + ((g836) & (!g901) & (g1163) & (g1246) & (g1728) & (g1729)) + ((g836) & (g901) & (!g1163) & (!g1246) & (g1728) & (!g1729)) + ((g836) & (g901) & (!g1163) & (!g1246) & (g1728) & (g1729)) + ((g836) & (g901) & (!g1163) & (g1246) & (!g1728) & (!g1729)) + ((g836) & (g901) & (!g1163) & (g1246) & (!g1728) & (g1729)) + ((g836) & (g901) & (g1163) & (!g1246) & (!g1728) & (!g1729)) + ((g836) & (g901) & (g1163) & (!g1246) & (g1728) & (!g1729)) + ((g836) & (g901) & (g1163) & (g1246) & (!g1728) & (!g1729)) + ((g836) & (g901) & (g1163) & (g1246) & (g1728) & (!g1729)));
	assign g1731 = (((!ld) & (!g852) & (!g1438) & (g1440) & (sk[52]) & (!keyx88x)) + ((!ld) & (!g852) & (!g1438) & (g1440) & (sk[52]) & (keyx88x)) + ((!ld) & (!g852) & (g1438) & (!g1440) & (sk[52]) & (!keyx88x)) + ((!ld) & (!g852) & (g1438) & (!g1440) & (sk[52]) & (keyx88x)) + ((!ld) & (g852) & (!g1438) & (!g1440) & (!sk[52]) & (!keyx88x)) + ((!ld) & (g852) & (!g1438) & (!g1440) & (!sk[52]) & (keyx88x)) + ((!ld) & (g852) & (!g1438) & (!g1440) & (sk[52]) & (!keyx88x)) + ((!ld) & (g852) & (!g1438) & (!g1440) & (sk[52]) & (keyx88x)) + ((!ld) & (g852) & (!g1438) & (g1440) & (!sk[52]) & (!keyx88x)) + ((!ld) & (g852) & (!g1438) & (g1440) & (!sk[52]) & (keyx88x)) + ((!ld) & (g852) & (g1438) & (!g1440) & (!sk[52]) & (!keyx88x)) + ((!ld) & (g852) & (g1438) & (!g1440) & (!sk[52]) & (keyx88x)) + ((!ld) & (g852) & (g1438) & (g1440) & (!sk[52]) & (!keyx88x)) + ((!ld) & (g852) & (g1438) & (g1440) & (!sk[52]) & (keyx88x)) + ((!ld) & (g852) & (g1438) & (g1440) & (sk[52]) & (!keyx88x)) + ((!ld) & (g852) & (g1438) & (g1440) & (sk[52]) & (keyx88x)) + ((ld) & (!g852) & (!g1438) & (!g1440) & (!sk[52]) & (!keyx88x)) + ((ld) & (!g852) & (!g1438) & (!g1440) & (!sk[52]) & (keyx88x)) + ((ld) & (!g852) & (!g1438) & (!g1440) & (sk[52]) & (keyx88x)) + ((ld) & (!g852) & (!g1438) & (g1440) & (!sk[52]) & (!keyx88x)) + ((ld) & (!g852) & (!g1438) & (g1440) & (!sk[52]) & (keyx88x)) + ((ld) & (!g852) & (!g1438) & (g1440) & (sk[52]) & (keyx88x)) + ((ld) & (!g852) & (g1438) & (!g1440) & (!sk[52]) & (!keyx88x)) + ((ld) & (!g852) & (g1438) & (!g1440) & (!sk[52]) & (keyx88x)) + ((ld) & (!g852) & (g1438) & (!g1440) & (sk[52]) & (keyx88x)) + ((ld) & (!g852) & (g1438) & (g1440) & (!sk[52]) & (!keyx88x)) + ((ld) & (!g852) & (g1438) & (g1440) & (!sk[52]) & (keyx88x)) + ((ld) & (!g852) & (g1438) & (g1440) & (sk[52]) & (keyx88x)) + ((ld) & (g852) & (!g1438) & (!g1440) & (!sk[52]) & (!keyx88x)) + ((ld) & (g852) & (!g1438) & (!g1440) & (!sk[52]) & (keyx88x)) + ((ld) & (g852) & (!g1438) & (!g1440) & (sk[52]) & (keyx88x)) + ((ld) & (g852) & (!g1438) & (g1440) & (!sk[52]) & (!keyx88x)) + ((ld) & (g852) & (!g1438) & (g1440) & (!sk[52]) & (keyx88x)) + ((ld) & (g852) & (!g1438) & (g1440) & (sk[52]) & (keyx88x)) + ((ld) & (g852) & (g1438) & (!g1440) & (!sk[52]) & (!keyx88x)) + ((ld) & (g852) & (g1438) & (!g1440) & (!sk[52]) & (keyx88x)) + ((ld) & (g852) & (g1438) & (!g1440) & (sk[52]) & (keyx88x)) + ((ld) & (g852) & (g1438) & (g1440) & (!sk[52]) & (!keyx88x)) + ((ld) & (g852) & (g1438) & (g1440) & (!sk[52]) & (keyx88x)) + ((ld) & (g852) & (g1438) & (g1440) & (sk[52]) & (keyx88x)));
	assign g1732 = (((!ld) & (!g859) & (!g1447) & (sk[53]) & (g1449) & (!keyx89x)) + ((!ld) & (!g859) & (!g1447) & (sk[53]) & (g1449) & (keyx89x)) + ((!ld) & (!g859) & (g1447) & (sk[53]) & (!g1449) & (!keyx89x)) + ((!ld) & (!g859) & (g1447) & (sk[53]) & (!g1449) & (keyx89x)) + ((!ld) & (g859) & (!g1447) & (!sk[53]) & (!g1449) & (!keyx89x)) + ((!ld) & (g859) & (!g1447) & (!sk[53]) & (!g1449) & (keyx89x)) + ((!ld) & (g859) & (!g1447) & (!sk[53]) & (g1449) & (!keyx89x)) + ((!ld) & (g859) & (!g1447) & (!sk[53]) & (g1449) & (keyx89x)) + ((!ld) & (g859) & (!g1447) & (sk[53]) & (!g1449) & (!keyx89x)) + ((!ld) & (g859) & (!g1447) & (sk[53]) & (!g1449) & (keyx89x)) + ((!ld) & (g859) & (g1447) & (!sk[53]) & (!g1449) & (!keyx89x)) + ((!ld) & (g859) & (g1447) & (!sk[53]) & (!g1449) & (keyx89x)) + ((!ld) & (g859) & (g1447) & (!sk[53]) & (g1449) & (!keyx89x)) + ((!ld) & (g859) & (g1447) & (!sk[53]) & (g1449) & (keyx89x)) + ((!ld) & (g859) & (g1447) & (sk[53]) & (g1449) & (!keyx89x)) + ((!ld) & (g859) & (g1447) & (sk[53]) & (g1449) & (keyx89x)) + ((ld) & (!g859) & (!g1447) & (!sk[53]) & (!g1449) & (!keyx89x)) + ((ld) & (!g859) & (!g1447) & (!sk[53]) & (!g1449) & (keyx89x)) + ((ld) & (!g859) & (!g1447) & (!sk[53]) & (g1449) & (!keyx89x)) + ((ld) & (!g859) & (!g1447) & (!sk[53]) & (g1449) & (keyx89x)) + ((ld) & (!g859) & (!g1447) & (sk[53]) & (!g1449) & (keyx89x)) + ((ld) & (!g859) & (!g1447) & (sk[53]) & (g1449) & (keyx89x)) + ((ld) & (!g859) & (g1447) & (!sk[53]) & (!g1449) & (!keyx89x)) + ((ld) & (!g859) & (g1447) & (!sk[53]) & (!g1449) & (keyx89x)) + ((ld) & (!g859) & (g1447) & (!sk[53]) & (g1449) & (!keyx89x)) + ((ld) & (!g859) & (g1447) & (!sk[53]) & (g1449) & (keyx89x)) + ((ld) & (!g859) & (g1447) & (sk[53]) & (!g1449) & (keyx89x)) + ((ld) & (!g859) & (g1447) & (sk[53]) & (g1449) & (keyx89x)) + ((ld) & (g859) & (!g1447) & (!sk[53]) & (!g1449) & (!keyx89x)) + ((ld) & (g859) & (!g1447) & (!sk[53]) & (!g1449) & (keyx89x)) + ((ld) & (g859) & (!g1447) & (!sk[53]) & (g1449) & (!keyx89x)) + ((ld) & (g859) & (!g1447) & (!sk[53]) & (g1449) & (keyx89x)) + ((ld) & (g859) & (!g1447) & (sk[53]) & (!g1449) & (keyx89x)) + ((ld) & (g859) & (!g1447) & (sk[53]) & (g1449) & (keyx89x)) + ((ld) & (g859) & (g1447) & (!sk[53]) & (!g1449) & (!keyx89x)) + ((ld) & (g859) & (g1447) & (!sk[53]) & (!g1449) & (keyx89x)) + ((ld) & (g859) & (g1447) & (!sk[53]) & (g1449) & (!keyx89x)) + ((ld) & (g859) & (g1447) & (!sk[53]) & (g1449) & (keyx89x)) + ((ld) & (g859) & (g1447) & (sk[53]) & (!g1449) & (keyx89x)) + ((ld) & (g859) & (g1447) & (sk[53]) & (g1449) & (keyx89x)));
	assign g1733 = (((!ld) & (!g866) & (sk[54]) & (!g1456) & (g1458) & (!keyx90x)) + ((!ld) & (!g866) & (sk[54]) & (!g1456) & (g1458) & (keyx90x)) + ((!ld) & (!g866) & (sk[54]) & (g1456) & (!g1458) & (!keyx90x)) + ((!ld) & (!g866) & (sk[54]) & (g1456) & (!g1458) & (keyx90x)) + ((!ld) & (g866) & (!sk[54]) & (!g1456) & (!g1458) & (!keyx90x)) + ((!ld) & (g866) & (!sk[54]) & (!g1456) & (!g1458) & (keyx90x)) + ((!ld) & (g866) & (!sk[54]) & (!g1456) & (g1458) & (!keyx90x)) + ((!ld) & (g866) & (!sk[54]) & (!g1456) & (g1458) & (keyx90x)) + ((!ld) & (g866) & (!sk[54]) & (g1456) & (!g1458) & (!keyx90x)) + ((!ld) & (g866) & (!sk[54]) & (g1456) & (!g1458) & (keyx90x)) + ((!ld) & (g866) & (!sk[54]) & (g1456) & (g1458) & (!keyx90x)) + ((!ld) & (g866) & (!sk[54]) & (g1456) & (g1458) & (keyx90x)) + ((!ld) & (g866) & (sk[54]) & (!g1456) & (!g1458) & (!keyx90x)) + ((!ld) & (g866) & (sk[54]) & (!g1456) & (!g1458) & (keyx90x)) + ((!ld) & (g866) & (sk[54]) & (g1456) & (g1458) & (!keyx90x)) + ((!ld) & (g866) & (sk[54]) & (g1456) & (g1458) & (keyx90x)) + ((ld) & (!g866) & (!sk[54]) & (!g1456) & (!g1458) & (!keyx90x)) + ((ld) & (!g866) & (!sk[54]) & (!g1456) & (!g1458) & (keyx90x)) + ((ld) & (!g866) & (!sk[54]) & (!g1456) & (g1458) & (!keyx90x)) + ((ld) & (!g866) & (!sk[54]) & (!g1456) & (g1458) & (keyx90x)) + ((ld) & (!g866) & (!sk[54]) & (g1456) & (!g1458) & (!keyx90x)) + ((ld) & (!g866) & (!sk[54]) & (g1456) & (!g1458) & (keyx90x)) + ((ld) & (!g866) & (!sk[54]) & (g1456) & (g1458) & (!keyx90x)) + ((ld) & (!g866) & (!sk[54]) & (g1456) & (g1458) & (keyx90x)) + ((ld) & (!g866) & (sk[54]) & (!g1456) & (!g1458) & (keyx90x)) + ((ld) & (!g866) & (sk[54]) & (!g1456) & (g1458) & (keyx90x)) + ((ld) & (!g866) & (sk[54]) & (g1456) & (!g1458) & (keyx90x)) + ((ld) & (!g866) & (sk[54]) & (g1456) & (g1458) & (keyx90x)) + ((ld) & (g866) & (!sk[54]) & (!g1456) & (!g1458) & (!keyx90x)) + ((ld) & (g866) & (!sk[54]) & (!g1456) & (!g1458) & (keyx90x)) + ((ld) & (g866) & (!sk[54]) & (!g1456) & (g1458) & (!keyx90x)) + ((ld) & (g866) & (!sk[54]) & (!g1456) & (g1458) & (keyx90x)) + ((ld) & (g866) & (!sk[54]) & (g1456) & (!g1458) & (!keyx90x)) + ((ld) & (g866) & (!sk[54]) & (g1456) & (!g1458) & (keyx90x)) + ((ld) & (g866) & (!sk[54]) & (g1456) & (g1458) & (!keyx90x)) + ((ld) & (g866) & (!sk[54]) & (g1456) & (g1458) & (keyx90x)) + ((ld) & (g866) & (sk[54]) & (!g1456) & (!g1458) & (keyx90x)) + ((ld) & (g866) & (sk[54]) & (!g1456) & (g1458) & (keyx90x)) + ((ld) & (g866) & (sk[54]) & (g1456) & (!g1458) & (keyx90x)) + ((ld) & (g866) & (sk[54]) & (g1456) & (g1458) & (keyx90x)));
	assign g1734 = (((!ld) & (!g873) & (!g1465) & (sk[55]) & (g1467) & (!keyx91x)) + ((!ld) & (!g873) & (!g1465) & (sk[55]) & (g1467) & (keyx91x)) + ((!ld) & (!g873) & (g1465) & (sk[55]) & (!g1467) & (!keyx91x)) + ((!ld) & (!g873) & (g1465) & (sk[55]) & (!g1467) & (keyx91x)) + ((!ld) & (g873) & (!g1465) & (!sk[55]) & (!g1467) & (!keyx91x)) + ((!ld) & (g873) & (!g1465) & (!sk[55]) & (!g1467) & (keyx91x)) + ((!ld) & (g873) & (!g1465) & (!sk[55]) & (g1467) & (!keyx91x)) + ((!ld) & (g873) & (!g1465) & (!sk[55]) & (g1467) & (keyx91x)) + ((!ld) & (g873) & (!g1465) & (sk[55]) & (!g1467) & (!keyx91x)) + ((!ld) & (g873) & (!g1465) & (sk[55]) & (!g1467) & (keyx91x)) + ((!ld) & (g873) & (g1465) & (!sk[55]) & (!g1467) & (!keyx91x)) + ((!ld) & (g873) & (g1465) & (!sk[55]) & (!g1467) & (keyx91x)) + ((!ld) & (g873) & (g1465) & (!sk[55]) & (g1467) & (!keyx91x)) + ((!ld) & (g873) & (g1465) & (!sk[55]) & (g1467) & (keyx91x)) + ((!ld) & (g873) & (g1465) & (sk[55]) & (g1467) & (!keyx91x)) + ((!ld) & (g873) & (g1465) & (sk[55]) & (g1467) & (keyx91x)) + ((ld) & (!g873) & (!g1465) & (!sk[55]) & (!g1467) & (!keyx91x)) + ((ld) & (!g873) & (!g1465) & (!sk[55]) & (!g1467) & (keyx91x)) + ((ld) & (!g873) & (!g1465) & (!sk[55]) & (g1467) & (!keyx91x)) + ((ld) & (!g873) & (!g1465) & (!sk[55]) & (g1467) & (keyx91x)) + ((ld) & (!g873) & (!g1465) & (sk[55]) & (!g1467) & (keyx91x)) + ((ld) & (!g873) & (!g1465) & (sk[55]) & (g1467) & (keyx91x)) + ((ld) & (!g873) & (g1465) & (!sk[55]) & (!g1467) & (!keyx91x)) + ((ld) & (!g873) & (g1465) & (!sk[55]) & (!g1467) & (keyx91x)) + ((ld) & (!g873) & (g1465) & (!sk[55]) & (g1467) & (!keyx91x)) + ((ld) & (!g873) & (g1465) & (!sk[55]) & (g1467) & (keyx91x)) + ((ld) & (!g873) & (g1465) & (sk[55]) & (!g1467) & (keyx91x)) + ((ld) & (!g873) & (g1465) & (sk[55]) & (g1467) & (keyx91x)) + ((ld) & (g873) & (!g1465) & (!sk[55]) & (!g1467) & (!keyx91x)) + ((ld) & (g873) & (!g1465) & (!sk[55]) & (!g1467) & (keyx91x)) + ((ld) & (g873) & (!g1465) & (!sk[55]) & (g1467) & (!keyx91x)) + ((ld) & (g873) & (!g1465) & (!sk[55]) & (g1467) & (keyx91x)) + ((ld) & (g873) & (!g1465) & (sk[55]) & (!g1467) & (keyx91x)) + ((ld) & (g873) & (!g1465) & (sk[55]) & (g1467) & (keyx91x)) + ((ld) & (g873) & (g1465) & (!sk[55]) & (!g1467) & (!keyx91x)) + ((ld) & (g873) & (g1465) & (!sk[55]) & (!g1467) & (keyx91x)) + ((ld) & (g873) & (g1465) & (!sk[55]) & (g1467) & (!keyx91x)) + ((ld) & (g873) & (g1465) & (!sk[55]) & (g1467) & (keyx91x)) + ((ld) & (g873) & (g1465) & (sk[55]) & (!g1467) & (keyx91x)) + ((ld) & (g873) & (g1465) & (sk[55]) & (g1467) & (keyx91x)));
	assign g1735 = (((!ld) & (!g880) & (!g1474) & (g1476) & (sk[56]) & (!keyx92x)) + ((!ld) & (!g880) & (!g1474) & (g1476) & (sk[56]) & (keyx92x)) + ((!ld) & (!g880) & (g1474) & (!g1476) & (sk[56]) & (!keyx92x)) + ((!ld) & (!g880) & (g1474) & (!g1476) & (sk[56]) & (keyx92x)) + ((!ld) & (g880) & (!g1474) & (!g1476) & (!sk[56]) & (!keyx92x)) + ((!ld) & (g880) & (!g1474) & (!g1476) & (!sk[56]) & (keyx92x)) + ((!ld) & (g880) & (!g1474) & (!g1476) & (sk[56]) & (!keyx92x)) + ((!ld) & (g880) & (!g1474) & (!g1476) & (sk[56]) & (keyx92x)) + ((!ld) & (g880) & (!g1474) & (g1476) & (!sk[56]) & (!keyx92x)) + ((!ld) & (g880) & (!g1474) & (g1476) & (!sk[56]) & (keyx92x)) + ((!ld) & (g880) & (g1474) & (!g1476) & (!sk[56]) & (!keyx92x)) + ((!ld) & (g880) & (g1474) & (!g1476) & (!sk[56]) & (keyx92x)) + ((!ld) & (g880) & (g1474) & (g1476) & (!sk[56]) & (!keyx92x)) + ((!ld) & (g880) & (g1474) & (g1476) & (!sk[56]) & (keyx92x)) + ((!ld) & (g880) & (g1474) & (g1476) & (sk[56]) & (!keyx92x)) + ((!ld) & (g880) & (g1474) & (g1476) & (sk[56]) & (keyx92x)) + ((ld) & (!g880) & (!g1474) & (!g1476) & (!sk[56]) & (!keyx92x)) + ((ld) & (!g880) & (!g1474) & (!g1476) & (!sk[56]) & (keyx92x)) + ((ld) & (!g880) & (!g1474) & (!g1476) & (sk[56]) & (keyx92x)) + ((ld) & (!g880) & (!g1474) & (g1476) & (!sk[56]) & (!keyx92x)) + ((ld) & (!g880) & (!g1474) & (g1476) & (!sk[56]) & (keyx92x)) + ((ld) & (!g880) & (!g1474) & (g1476) & (sk[56]) & (keyx92x)) + ((ld) & (!g880) & (g1474) & (!g1476) & (!sk[56]) & (!keyx92x)) + ((ld) & (!g880) & (g1474) & (!g1476) & (!sk[56]) & (keyx92x)) + ((ld) & (!g880) & (g1474) & (!g1476) & (sk[56]) & (keyx92x)) + ((ld) & (!g880) & (g1474) & (g1476) & (!sk[56]) & (!keyx92x)) + ((ld) & (!g880) & (g1474) & (g1476) & (!sk[56]) & (keyx92x)) + ((ld) & (!g880) & (g1474) & (g1476) & (sk[56]) & (keyx92x)) + ((ld) & (g880) & (!g1474) & (!g1476) & (!sk[56]) & (!keyx92x)) + ((ld) & (g880) & (!g1474) & (!g1476) & (!sk[56]) & (keyx92x)) + ((ld) & (g880) & (!g1474) & (!g1476) & (sk[56]) & (keyx92x)) + ((ld) & (g880) & (!g1474) & (g1476) & (!sk[56]) & (!keyx92x)) + ((ld) & (g880) & (!g1474) & (g1476) & (!sk[56]) & (keyx92x)) + ((ld) & (g880) & (!g1474) & (g1476) & (sk[56]) & (keyx92x)) + ((ld) & (g880) & (g1474) & (!g1476) & (!sk[56]) & (!keyx92x)) + ((ld) & (g880) & (g1474) & (!g1476) & (!sk[56]) & (keyx92x)) + ((ld) & (g880) & (g1474) & (!g1476) & (sk[56]) & (keyx92x)) + ((ld) & (g880) & (g1474) & (g1476) & (!sk[56]) & (!keyx92x)) + ((ld) & (g880) & (g1474) & (g1476) & (!sk[56]) & (keyx92x)) + ((ld) & (g880) & (g1474) & (g1476) & (sk[56]) & (keyx92x)));
	assign g1736 = (((!sk[57]) & (!ld) & (g887) & (!g1483) & (!g1485) & (!keyx93x)) + ((!sk[57]) & (!ld) & (g887) & (!g1483) & (!g1485) & (keyx93x)) + ((!sk[57]) & (!ld) & (g887) & (!g1483) & (g1485) & (!keyx93x)) + ((!sk[57]) & (!ld) & (g887) & (!g1483) & (g1485) & (keyx93x)) + ((!sk[57]) & (!ld) & (g887) & (g1483) & (!g1485) & (!keyx93x)) + ((!sk[57]) & (!ld) & (g887) & (g1483) & (!g1485) & (keyx93x)) + ((!sk[57]) & (!ld) & (g887) & (g1483) & (g1485) & (!keyx93x)) + ((!sk[57]) & (!ld) & (g887) & (g1483) & (g1485) & (keyx93x)) + ((!sk[57]) & (ld) & (!g887) & (!g1483) & (!g1485) & (!keyx93x)) + ((!sk[57]) & (ld) & (!g887) & (!g1483) & (!g1485) & (keyx93x)) + ((!sk[57]) & (ld) & (!g887) & (!g1483) & (g1485) & (!keyx93x)) + ((!sk[57]) & (ld) & (!g887) & (!g1483) & (g1485) & (keyx93x)) + ((!sk[57]) & (ld) & (!g887) & (g1483) & (!g1485) & (!keyx93x)) + ((!sk[57]) & (ld) & (!g887) & (g1483) & (!g1485) & (keyx93x)) + ((!sk[57]) & (ld) & (!g887) & (g1483) & (g1485) & (!keyx93x)) + ((!sk[57]) & (ld) & (!g887) & (g1483) & (g1485) & (keyx93x)) + ((!sk[57]) & (ld) & (g887) & (!g1483) & (!g1485) & (!keyx93x)) + ((!sk[57]) & (ld) & (g887) & (!g1483) & (!g1485) & (keyx93x)) + ((!sk[57]) & (ld) & (g887) & (!g1483) & (g1485) & (!keyx93x)) + ((!sk[57]) & (ld) & (g887) & (!g1483) & (g1485) & (keyx93x)) + ((!sk[57]) & (ld) & (g887) & (g1483) & (!g1485) & (!keyx93x)) + ((!sk[57]) & (ld) & (g887) & (g1483) & (!g1485) & (keyx93x)) + ((!sk[57]) & (ld) & (g887) & (g1483) & (g1485) & (!keyx93x)) + ((!sk[57]) & (ld) & (g887) & (g1483) & (g1485) & (keyx93x)) + ((sk[57]) & (!ld) & (!g887) & (!g1483) & (g1485) & (!keyx93x)) + ((sk[57]) & (!ld) & (!g887) & (!g1483) & (g1485) & (keyx93x)) + ((sk[57]) & (!ld) & (!g887) & (g1483) & (!g1485) & (!keyx93x)) + ((sk[57]) & (!ld) & (!g887) & (g1483) & (!g1485) & (keyx93x)) + ((sk[57]) & (!ld) & (g887) & (!g1483) & (!g1485) & (!keyx93x)) + ((sk[57]) & (!ld) & (g887) & (!g1483) & (!g1485) & (keyx93x)) + ((sk[57]) & (!ld) & (g887) & (g1483) & (g1485) & (!keyx93x)) + ((sk[57]) & (!ld) & (g887) & (g1483) & (g1485) & (keyx93x)) + ((sk[57]) & (ld) & (!g887) & (!g1483) & (!g1485) & (keyx93x)) + ((sk[57]) & (ld) & (!g887) & (!g1483) & (g1485) & (keyx93x)) + ((sk[57]) & (ld) & (!g887) & (g1483) & (!g1485) & (keyx93x)) + ((sk[57]) & (ld) & (!g887) & (g1483) & (g1485) & (keyx93x)) + ((sk[57]) & (ld) & (g887) & (!g1483) & (!g1485) & (keyx93x)) + ((sk[57]) & (ld) & (g887) & (!g1483) & (g1485) & (keyx93x)) + ((sk[57]) & (ld) & (g887) & (g1483) & (!g1485) & (keyx93x)) + ((sk[57]) & (ld) & (g887) & (g1483) & (g1485) & (keyx93x)));
	assign g1737 = (((!ld) & (!g894) & (!g1492) & (g1494) & (sk[58]) & (!keyx94x)) + ((!ld) & (!g894) & (!g1492) & (g1494) & (sk[58]) & (keyx94x)) + ((!ld) & (!g894) & (g1492) & (!g1494) & (sk[58]) & (!keyx94x)) + ((!ld) & (!g894) & (g1492) & (!g1494) & (sk[58]) & (keyx94x)) + ((!ld) & (g894) & (!g1492) & (!g1494) & (!sk[58]) & (!keyx94x)) + ((!ld) & (g894) & (!g1492) & (!g1494) & (!sk[58]) & (keyx94x)) + ((!ld) & (g894) & (!g1492) & (!g1494) & (sk[58]) & (!keyx94x)) + ((!ld) & (g894) & (!g1492) & (!g1494) & (sk[58]) & (keyx94x)) + ((!ld) & (g894) & (!g1492) & (g1494) & (!sk[58]) & (!keyx94x)) + ((!ld) & (g894) & (!g1492) & (g1494) & (!sk[58]) & (keyx94x)) + ((!ld) & (g894) & (g1492) & (!g1494) & (!sk[58]) & (!keyx94x)) + ((!ld) & (g894) & (g1492) & (!g1494) & (!sk[58]) & (keyx94x)) + ((!ld) & (g894) & (g1492) & (g1494) & (!sk[58]) & (!keyx94x)) + ((!ld) & (g894) & (g1492) & (g1494) & (!sk[58]) & (keyx94x)) + ((!ld) & (g894) & (g1492) & (g1494) & (sk[58]) & (!keyx94x)) + ((!ld) & (g894) & (g1492) & (g1494) & (sk[58]) & (keyx94x)) + ((ld) & (!g894) & (!g1492) & (!g1494) & (!sk[58]) & (!keyx94x)) + ((ld) & (!g894) & (!g1492) & (!g1494) & (!sk[58]) & (keyx94x)) + ((ld) & (!g894) & (!g1492) & (!g1494) & (sk[58]) & (keyx94x)) + ((ld) & (!g894) & (!g1492) & (g1494) & (!sk[58]) & (!keyx94x)) + ((ld) & (!g894) & (!g1492) & (g1494) & (!sk[58]) & (keyx94x)) + ((ld) & (!g894) & (!g1492) & (g1494) & (sk[58]) & (keyx94x)) + ((ld) & (!g894) & (g1492) & (!g1494) & (!sk[58]) & (!keyx94x)) + ((ld) & (!g894) & (g1492) & (!g1494) & (!sk[58]) & (keyx94x)) + ((ld) & (!g894) & (g1492) & (!g1494) & (sk[58]) & (keyx94x)) + ((ld) & (!g894) & (g1492) & (g1494) & (!sk[58]) & (!keyx94x)) + ((ld) & (!g894) & (g1492) & (g1494) & (!sk[58]) & (keyx94x)) + ((ld) & (!g894) & (g1492) & (g1494) & (sk[58]) & (keyx94x)) + ((ld) & (g894) & (!g1492) & (!g1494) & (!sk[58]) & (!keyx94x)) + ((ld) & (g894) & (!g1492) & (!g1494) & (!sk[58]) & (keyx94x)) + ((ld) & (g894) & (!g1492) & (!g1494) & (sk[58]) & (keyx94x)) + ((ld) & (g894) & (!g1492) & (g1494) & (!sk[58]) & (!keyx94x)) + ((ld) & (g894) & (!g1492) & (g1494) & (!sk[58]) & (keyx94x)) + ((ld) & (g894) & (!g1492) & (g1494) & (sk[58]) & (keyx94x)) + ((ld) & (g894) & (g1492) & (!g1494) & (!sk[58]) & (!keyx94x)) + ((ld) & (g894) & (g1492) & (!g1494) & (!sk[58]) & (keyx94x)) + ((ld) & (g894) & (g1492) & (!g1494) & (sk[58]) & (keyx94x)) + ((ld) & (g894) & (g1492) & (g1494) & (!sk[58]) & (!keyx94x)) + ((ld) & (g894) & (g1492) & (g1494) & (!sk[58]) & (keyx94x)) + ((ld) & (g894) & (g1492) & (g1494) & (sk[58]) & (keyx94x)));
	assign g1738 = (((!ld) & (!g901) & (!g1501) & (g1503) & (sk[59]) & (!keyx95x)) + ((!ld) & (!g901) & (!g1501) & (g1503) & (sk[59]) & (keyx95x)) + ((!ld) & (!g901) & (g1501) & (!g1503) & (sk[59]) & (!keyx95x)) + ((!ld) & (!g901) & (g1501) & (!g1503) & (sk[59]) & (keyx95x)) + ((!ld) & (g901) & (!g1501) & (!g1503) & (!sk[59]) & (!keyx95x)) + ((!ld) & (g901) & (!g1501) & (!g1503) & (!sk[59]) & (keyx95x)) + ((!ld) & (g901) & (!g1501) & (!g1503) & (sk[59]) & (!keyx95x)) + ((!ld) & (g901) & (!g1501) & (!g1503) & (sk[59]) & (keyx95x)) + ((!ld) & (g901) & (!g1501) & (g1503) & (!sk[59]) & (!keyx95x)) + ((!ld) & (g901) & (!g1501) & (g1503) & (!sk[59]) & (keyx95x)) + ((!ld) & (g901) & (g1501) & (!g1503) & (!sk[59]) & (!keyx95x)) + ((!ld) & (g901) & (g1501) & (!g1503) & (!sk[59]) & (keyx95x)) + ((!ld) & (g901) & (g1501) & (g1503) & (!sk[59]) & (!keyx95x)) + ((!ld) & (g901) & (g1501) & (g1503) & (!sk[59]) & (keyx95x)) + ((!ld) & (g901) & (g1501) & (g1503) & (sk[59]) & (!keyx95x)) + ((!ld) & (g901) & (g1501) & (g1503) & (sk[59]) & (keyx95x)) + ((ld) & (!g901) & (!g1501) & (!g1503) & (!sk[59]) & (!keyx95x)) + ((ld) & (!g901) & (!g1501) & (!g1503) & (!sk[59]) & (keyx95x)) + ((ld) & (!g901) & (!g1501) & (!g1503) & (sk[59]) & (keyx95x)) + ((ld) & (!g901) & (!g1501) & (g1503) & (!sk[59]) & (!keyx95x)) + ((ld) & (!g901) & (!g1501) & (g1503) & (!sk[59]) & (keyx95x)) + ((ld) & (!g901) & (!g1501) & (g1503) & (sk[59]) & (keyx95x)) + ((ld) & (!g901) & (g1501) & (!g1503) & (!sk[59]) & (!keyx95x)) + ((ld) & (!g901) & (g1501) & (!g1503) & (!sk[59]) & (keyx95x)) + ((ld) & (!g901) & (g1501) & (!g1503) & (sk[59]) & (keyx95x)) + ((ld) & (!g901) & (g1501) & (g1503) & (!sk[59]) & (!keyx95x)) + ((ld) & (!g901) & (g1501) & (g1503) & (!sk[59]) & (keyx95x)) + ((ld) & (!g901) & (g1501) & (g1503) & (sk[59]) & (keyx95x)) + ((ld) & (g901) & (!g1501) & (!g1503) & (!sk[59]) & (!keyx95x)) + ((ld) & (g901) & (!g1501) & (!g1503) & (!sk[59]) & (keyx95x)) + ((ld) & (g901) & (!g1501) & (!g1503) & (sk[59]) & (keyx95x)) + ((ld) & (g901) & (!g1501) & (g1503) & (!sk[59]) & (!keyx95x)) + ((ld) & (g901) & (!g1501) & (g1503) & (!sk[59]) & (keyx95x)) + ((ld) & (g901) & (!g1501) & (g1503) & (sk[59]) & (keyx95x)) + ((ld) & (g901) & (g1501) & (!g1503) & (!sk[59]) & (!keyx95x)) + ((ld) & (g901) & (g1501) & (!g1503) & (!sk[59]) & (keyx95x)) + ((ld) & (g901) & (g1501) & (!g1503) & (sk[59]) & (keyx95x)) + ((ld) & (g901) & (g1501) & (g1503) & (!sk[59]) & (!keyx95x)) + ((ld) & (g901) & (g1501) & (g1503) & (!sk[59]) & (keyx95x)) + ((ld) & (g901) & (g1501) & (g1503) & (sk[59]) & (keyx95x)));
	assign g2178 = (((!ld) & (!sk[60]) & (text_inx0x) & (!g1739)) + ((!ld) & (!sk[60]) & (text_inx0x) & (g1739)) + ((!ld) & (sk[60]) & (!text_inx0x) & (g1739)) + ((!ld) & (sk[60]) & (text_inx0x) & (g1739)) + ((ld) & (!sk[60]) & (!text_inx0x) & (g1739)) + ((ld) & (!sk[60]) & (text_inx0x) & (!g1739)) + ((ld) & (!sk[60]) & (text_inx0x) & (g1739)) + ((ld) & (sk[60]) & (text_inx0x) & (!g1739)) + ((ld) & (sk[60]) & (text_inx0x) & (g1739)));
	assign g1740 = (((!g196) & (!g339) & (sk[61]) & (g388)) + ((!g196) & (g339) & (!sk[61]) & (!g388)) + ((!g196) & (g339) & (!sk[61]) & (g388)) + ((!g196) & (g339) & (sk[61]) & (!g388)) + ((g196) & (!g339) & (!sk[61]) & (g388)) + ((g196) & (!g339) & (sk[61]) & (!g388)) + ((g196) & (g339) & (!sk[61]) & (!g388)) + ((g196) & (g339) & (!sk[61]) & (g388)) + ((g196) & (g339) & (sk[61]) & (g388)));
	assign g1741 = (((!g148) & (!g211) & (!g275) & (!g1163) & (!g1739) & (g1740)) + ((!g148) & (!g211) & (!g275) & (!g1163) & (g1739) & (g1740)) + ((!g148) & (!g211) & (!g275) & (g1163) & (g1739) & (!g1740)) + ((!g148) & (!g211) & (!g275) & (g1163) & (g1739) & (g1740)) + ((!g148) & (!g211) & (g275) & (!g1163) & (!g1739) & (!g1740)) + ((!g148) & (!g211) & (g275) & (!g1163) & (g1739) & (!g1740)) + ((!g148) & (!g211) & (g275) & (g1163) & (g1739) & (!g1740)) + ((!g148) & (!g211) & (g275) & (g1163) & (g1739) & (g1740)) + ((!g148) & (g211) & (!g275) & (!g1163) & (!g1739) & (!g1740)) + ((!g148) & (g211) & (!g275) & (!g1163) & (g1739) & (!g1740)) + ((!g148) & (g211) & (!g275) & (g1163) & (g1739) & (!g1740)) + ((!g148) & (g211) & (!g275) & (g1163) & (g1739) & (g1740)) + ((!g148) & (g211) & (g275) & (!g1163) & (!g1739) & (g1740)) + ((!g148) & (g211) & (g275) & (!g1163) & (g1739) & (g1740)) + ((!g148) & (g211) & (g275) & (g1163) & (g1739) & (!g1740)) + ((!g148) & (g211) & (g275) & (g1163) & (g1739) & (g1740)) + ((g148) & (!g211) & (!g275) & (!g1163) & (!g1739) & (!g1740)) + ((g148) & (!g211) & (!g275) & (!g1163) & (g1739) & (!g1740)) + ((g148) & (!g211) & (!g275) & (g1163) & (!g1739) & (!g1740)) + ((g148) & (!g211) & (!g275) & (g1163) & (!g1739) & (g1740)) + ((g148) & (!g211) & (g275) & (!g1163) & (!g1739) & (g1740)) + ((g148) & (!g211) & (g275) & (!g1163) & (g1739) & (g1740)) + ((g148) & (!g211) & (g275) & (g1163) & (!g1739) & (!g1740)) + ((g148) & (!g211) & (g275) & (g1163) & (!g1739) & (g1740)) + ((g148) & (g211) & (!g275) & (!g1163) & (!g1739) & (g1740)) + ((g148) & (g211) & (!g275) & (!g1163) & (g1739) & (g1740)) + ((g148) & (g211) & (!g275) & (g1163) & (!g1739) & (!g1740)) + ((g148) & (g211) & (!g275) & (g1163) & (!g1739) & (g1740)) + ((g148) & (g211) & (g275) & (!g1163) & (!g1739) & (!g1740)) + ((g148) & (g211) & (g275) & (!g1163) & (g1739) & (!g1740)) + ((g148) & (g211) & (g275) & (g1163) & (!g1739) & (!g1740)) + ((g148) & (g211) & (g275) & (g1163) & (!g1739) & (g1740)));
	assign g2179 = (((!ld) & (!text_inx1x) & (sk[63]) & (g1742)) + ((!ld) & (text_inx1x) & (!sk[63]) & (!g1742)) + ((!ld) & (text_inx1x) & (!sk[63]) & (g1742)) + ((!ld) & (text_inx1x) & (sk[63]) & (g1742)) + ((ld) & (!text_inx1x) & (!sk[63]) & (g1742)) + ((ld) & (text_inx1x) & (!sk[63]) & (!g1742)) + ((ld) & (text_inx1x) & (!sk[63]) & (g1742)) + ((ld) & (text_inx1x) & (sk[63]) & (!g1742)) + ((ld) & (text_inx1x) & (sk[63]) & (g1742)));
	assign g1743 = (((!g155) & (!g218) & (!g1163) & (!g1647) & (g1740) & (!g1742)) + ((!g155) & (!g218) & (!g1163) & (!g1647) & (g1740) & (g1742)) + ((!g155) & (!g218) & (!g1163) & (g1647) & (!g1740) & (!g1742)) + ((!g155) & (!g218) & (!g1163) & (g1647) & (!g1740) & (g1742)) + ((!g155) & (!g218) & (g1163) & (!g1647) & (!g1740) & (g1742)) + ((!g155) & (!g218) & (g1163) & (!g1647) & (g1740) & (g1742)) + ((!g155) & (!g218) & (g1163) & (g1647) & (!g1740) & (g1742)) + ((!g155) & (!g218) & (g1163) & (g1647) & (g1740) & (g1742)) + ((!g155) & (g218) & (!g1163) & (!g1647) & (!g1740) & (!g1742)) + ((!g155) & (g218) & (!g1163) & (!g1647) & (!g1740) & (g1742)) + ((!g155) & (g218) & (!g1163) & (g1647) & (g1740) & (!g1742)) + ((!g155) & (g218) & (!g1163) & (g1647) & (g1740) & (g1742)) + ((!g155) & (g218) & (g1163) & (!g1647) & (!g1740) & (g1742)) + ((!g155) & (g218) & (g1163) & (!g1647) & (g1740) & (g1742)) + ((!g155) & (g218) & (g1163) & (g1647) & (!g1740) & (g1742)) + ((!g155) & (g218) & (g1163) & (g1647) & (g1740) & (g1742)) + ((g155) & (!g218) & (!g1163) & (!g1647) & (!g1740) & (!g1742)) + ((g155) & (!g218) & (!g1163) & (!g1647) & (!g1740) & (g1742)) + ((g155) & (!g218) & (!g1163) & (g1647) & (g1740) & (!g1742)) + ((g155) & (!g218) & (!g1163) & (g1647) & (g1740) & (g1742)) + ((g155) & (!g218) & (g1163) & (!g1647) & (!g1740) & (!g1742)) + ((g155) & (!g218) & (g1163) & (!g1647) & (g1740) & (!g1742)) + ((g155) & (!g218) & (g1163) & (g1647) & (!g1740) & (!g1742)) + ((g155) & (!g218) & (g1163) & (g1647) & (g1740) & (!g1742)) + ((g155) & (g218) & (!g1163) & (!g1647) & (g1740) & (!g1742)) + ((g155) & (g218) & (!g1163) & (!g1647) & (g1740) & (g1742)) + ((g155) & (g218) & (!g1163) & (g1647) & (!g1740) & (!g1742)) + ((g155) & (g218) & (!g1163) & (g1647) & (!g1740) & (g1742)) + ((g155) & (g218) & (g1163) & (!g1647) & (!g1740) & (!g1742)) + ((g155) & (g218) & (g1163) & (!g1647) & (g1740) & (!g1742)) + ((g155) & (g218) & (g1163) & (g1647) & (!g1740) & (!g1742)) + ((g155) & (g218) & (g1163) & (g1647) & (g1740) & (!g1742)));
	assign g2180 = (((!sk[65]) & (!ld) & (text_inx2x) & (!g1744)) + ((!sk[65]) & (!ld) & (text_inx2x) & (g1744)) + ((!sk[65]) & (ld) & (!text_inx2x) & (g1744)) + ((!sk[65]) & (ld) & (text_inx2x) & (!g1744)) + ((!sk[65]) & (ld) & (text_inx2x) & (g1744)) + ((sk[65]) & (!ld) & (!text_inx2x) & (g1744)) + ((sk[65]) & (!ld) & (text_inx2x) & (g1744)) + ((sk[65]) & (ld) & (text_inx2x) & (!g1744)) + ((sk[65]) & (ld) & (text_inx2x) & (g1744)));
	assign g1745 = (((!g162) & (!g225) & (!g346) & (!g1163) & (g1651) & (!g1744)) + ((!g162) & (!g225) & (!g346) & (!g1163) & (g1651) & (g1744)) + ((!g162) & (!g225) & (!g346) & (g1163) & (!g1651) & (g1744)) + ((!g162) & (!g225) & (!g346) & (g1163) & (g1651) & (g1744)) + ((!g162) & (!g225) & (g346) & (!g1163) & (!g1651) & (!g1744)) + ((!g162) & (!g225) & (g346) & (!g1163) & (!g1651) & (g1744)) + ((!g162) & (!g225) & (g346) & (g1163) & (!g1651) & (g1744)) + ((!g162) & (!g225) & (g346) & (g1163) & (g1651) & (g1744)) + ((!g162) & (g225) & (!g346) & (!g1163) & (!g1651) & (!g1744)) + ((!g162) & (g225) & (!g346) & (!g1163) & (!g1651) & (g1744)) + ((!g162) & (g225) & (!g346) & (g1163) & (!g1651) & (g1744)) + ((!g162) & (g225) & (!g346) & (g1163) & (g1651) & (g1744)) + ((!g162) & (g225) & (g346) & (!g1163) & (g1651) & (!g1744)) + ((!g162) & (g225) & (g346) & (!g1163) & (g1651) & (g1744)) + ((!g162) & (g225) & (g346) & (g1163) & (!g1651) & (g1744)) + ((!g162) & (g225) & (g346) & (g1163) & (g1651) & (g1744)) + ((g162) & (!g225) & (!g346) & (!g1163) & (!g1651) & (!g1744)) + ((g162) & (!g225) & (!g346) & (!g1163) & (!g1651) & (g1744)) + ((g162) & (!g225) & (!g346) & (g1163) & (!g1651) & (!g1744)) + ((g162) & (!g225) & (!g346) & (g1163) & (g1651) & (!g1744)) + ((g162) & (!g225) & (g346) & (!g1163) & (g1651) & (!g1744)) + ((g162) & (!g225) & (g346) & (!g1163) & (g1651) & (g1744)) + ((g162) & (!g225) & (g346) & (g1163) & (!g1651) & (!g1744)) + ((g162) & (!g225) & (g346) & (g1163) & (g1651) & (!g1744)) + ((g162) & (g225) & (!g346) & (!g1163) & (g1651) & (!g1744)) + ((g162) & (g225) & (!g346) & (!g1163) & (g1651) & (g1744)) + ((g162) & (g225) & (!g346) & (g1163) & (!g1651) & (!g1744)) + ((g162) & (g225) & (!g346) & (g1163) & (g1651) & (!g1744)) + ((g162) & (g225) & (g346) & (!g1163) & (!g1651) & (!g1744)) + ((g162) & (g225) & (g346) & (!g1163) & (!g1651) & (g1744)) + ((g162) & (g225) & (g346) & (g1163) & (!g1651) & (!g1744)) + ((g162) & (g225) & (g346) & (g1163) & (g1651) & (!g1744)));
	assign g2181 = (((!ld) & (!sk[67]) & (text_inx3x) & (!g1746)) + ((!ld) & (!sk[67]) & (text_inx3x) & (g1746)) + ((!ld) & (sk[67]) & (!text_inx3x) & (g1746)) + ((!ld) & (sk[67]) & (text_inx3x) & (g1746)) + ((ld) & (!sk[67]) & (!text_inx3x) & (g1746)) + ((ld) & (!sk[67]) & (text_inx3x) & (!g1746)) + ((ld) & (!sk[67]) & (text_inx3x) & (g1746)) + ((ld) & (sk[67]) & (text_inx3x) & (!g1746)) + ((ld) & (sk[67]) & (text_inx3x) & (g1746)));
	assign g1747 = (((!g169) & (!sk[68]) & (g196) & (!g232) & (!g353) & (!g388)) + ((!g169) & (!sk[68]) & (g196) & (!g232) & (!g353) & (g388)) + ((!g169) & (!sk[68]) & (g196) & (!g232) & (g353) & (!g388)) + ((!g169) & (!sk[68]) & (g196) & (!g232) & (g353) & (g388)) + ((!g169) & (!sk[68]) & (g196) & (g232) & (!g353) & (!g388)) + ((!g169) & (!sk[68]) & (g196) & (g232) & (!g353) & (g388)) + ((!g169) & (!sk[68]) & (g196) & (g232) & (g353) & (!g388)) + ((!g169) & (!sk[68]) & (g196) & (g232) & (g353) & (g388)) + ((!g169) & (sk[68]) & (!g196) & (!g232) & (!g353) & (g388)) + ((!g169) & (sk[68]) & (!g196) & (!g232) & (g353) & (!g388)) + ((!g169) & (sk[68]) & (!g196) & (g232) & (!g353) & (!g388)) + ((!g169) & (sk[68]) & (!g196) & (g232) & (g353) & (g388)) + ((!g169) & (sk[68]) & (g196) & (!g232) & (!g353) & (!g388)) + ((!g169) & (sk[68]) & (g196) & (!g232) & (g353) & (g388)) + ((!g169) & (sk[68]) & (g196) & (g232) & (!g353) & (g388)) + ((!g169) & (sk[68]) & (g196) & (g232) & (g353) & (!g388)) + ((g169) & (!sk[68]) & (!g196) & (!g232) & (!g353) & (!g388)) + ((g169) & (!sk[68]) & (!g196) & (!g232) & (!g353) & (g388)) + ((g169) & (!sk[68]) & (!g196) & (!g232) & (g353) & (!g388)) + ((g169) & (!sk[68]) & (!g196) & (!g232) & (g353) & (g388)) + ((g169) & (!sk[68]) & (!g196) & (g232) & (!g353) & (!g388)) + ((g169) & (!sk[68]) & (!g196) & (g232) & (!g353) & (g388)) + ((g169) & (!sk[68]) & (!g196) & (g232) & (g353) & (!g388)) + ((g169) & (!sk[68]) & (!g196) & (g232) & (g353) & (g388)) + ((g169) & (!sk[68]) & (g196) & (!g232) & (!g353) & (!g388)) + ((g169) & (!sk[68]) & (g196) & (!g232) & (!g353) & (g388)) + ((g169) & (!sk[68]) & (g196) & (!g232) & (g353) & (!g388)) + ((g169) & (!sk[68]) & (g196) & (!g232) & (g353) & (g388)) + ((g169) & (!sk[68]) & (g196) & (g232) & (!g353) & (!g388)) + ((g169) & (!sk[68]) & (g196) & (g232) & (!g353) & (g388)) + ((g169) & (!sk[68]) & (g196) & (g232) & (g353) & (!g388)) + ((g169) & (!sk[68]) & (g196) & (g232) & (g353) & (g388)) + ((g169) & (sk[68]) & (!g196) & (!g232) & (!g353) & (!g388)) + ((g169) & (sk[68]) & (!g196) & (!g232) & (g353) & (g388)) + ((g169) & (sk[68]) & (!g196) & (g232) & (!g353) & (g388)) + ((g169) & (sk[68]) & (!g196) & (g232) & (g353) & (!g388)) + ((g169) & (sk[68]) & (g196) & (!g232) & (!g353) & (g388)) + ((g169) & (sk[68]) & (g196) & (!g232) & (g353) & (!g388)) + ((g169) & (sk[68]) & (g196) & (g232) & (!g353) & (!g388)) + ((g169) & (sk[68]) & (g196) & (g232) & (g353) & (g388)));
	assign g1748 = (((!g169) & (!g1163) & (!g1654) & (!g1746) & (sk[69]) & (g1747)) + ((!g169) & (!g1163) & (!g1654) & (g1746) & (sk[69]) & (g1747)) + ((!g169) & (!g1163) & (g1654) & (!g1746) & (sk[69]) & (!g1747)) + ((!g169) & (!g1163) & (g1654) & (g1746) & (sk[69]) & (!g1747)) + ((!g169) & (g1163) & (!g1654) & (!g1746) & (!sk[69]) & (!g1747)) + ((!g169) & (g1163) & (!g1654) & (!g1746) & (!sk[69]) & (g1747)) + ((!g169) & (g1163) & (!g1654) & (g1746) & (!sk[69]) & (!g1747)) + ((!g169) & (g1163) & (!g1654) & (g1746) & (!sk[69]) & (g1747)) + ((!g169) & (g1163) & (!g1654) & (g1746) & (sk[69]) & (!g1747)) + ((!g169) & (g1163) & (!g1654) & (g1746) & (sk[69]) & (g1747)) + ((!g169) & (g1163) & (g1654) & (!g1746) & (!sk[69]) & (!g1747)) + ((!g169) & (g1163) & (g1654) & (!g1746) & (!sk[69]) & (g1747)) + ((!g169) & (g1163) & (g1654) & (g1746) & (!sk[69]) & (!g1747)) + ((!g169) & (g1163) & (g1654) & (g1746) & (!sk[69]) & (g1747)) + ((!g169) & (g1163) & (g1654) & (g1746) & (sk[69]) & (!g1747)) + ((!g169) & (g1163) & (g1654) & (g1746) & (sk[69]) & (g1747)) + ((g169) & (!g1163) & (!g1654) & (!g1746) & (!sk[69]) & (!g1747)) + ((g169) & (!g1163) & (!g1654) & (!g1746) & (!sk[69]) & (g1747)) + ((g169) & (!g1163) & (!g1654) & (!g1746) & (sk[69]) & (g1747)) + ((g169) & (!g1163) & (!g1654) & (g1746) & (!sk[69]) & (!g1747)) + ((g169) & (!g1163) & (!g1654) & (g1746) & (!sk[69]) & (g1747)) + ((g169) & (!g1163) & (!g1654) & (g1746) & (sk[69]) & (g1747)) + ((g169) & (!g1163) & (g1654) & (!g1746) & (!sk[69]) & (!g1747)) + ((g169) & (!g1163) & (g1654) & (!g1746) & (!sk[69]) & (g1747)) + ((g169) & (!g1163) & (g1654) & (!g1746) & (sk[69]) & (!g1747)) + ((g169) & (!g1163) & (g1654) & (g1746) & (!sk[69]) & (!g1747)) + ((g169) & (!g1163) & (g1654) & (g1746) & (!sk[69]) & (g1747)) + ((g169) & (!g1163) & (g1654) & (g1746) & (sk[69]) & (!g1747)) + ((g169) & (g1163) & (!g1654) & (!g1746) & (!sk[69]) & (!g1747)) + ((g169) & (g1163) & (!g1654) & (!g1746) & (!sk[69]) & (g1747)) + ((g169) & (g1163) & (!g1654) & (!g1746) & (sk[69]) & (!g1747)) + ((g169) & (g1163) & (!g1654) & (!g1746) & (sk[69]) & (g1747)) + ((g169) & (g1163) & (!g1654) & (g1746) & (!sk[69]) & (!g1747)) + ((g169) & (g1163) & (!g1654) & (g1746) & (!sk[69]) & (g1747)) + ((g169) & (g1163) & (g1654) & (!g1746) & (!sk[69]) & (!g1747)) + ((g169) & (g1163) & (g1654) & (!g1746) & (!sk[69]) & (g1747)) + ((g169) & (g1163) & (g1654) & (!g1746) & (sk[69]) & (!g1747)) + ((g169) & (g1163) & (g1654) & (!g1746) & (sk[69]) & (g1747)) + ((g169) & (g1163) & (g1654) & (g1746) & (!sk[69]) & (!g1747)) + ((g169) & (g1163) & (g1654) & (g1746) & (!sk[69]) & (g1747)));
	assign g2182 = (((!sk[70]) & (!ld) & (text_inx6x) & (!g1749)) + ((!sk[70]) & (!ld) & (text_inx6x) & (g1749)) + ((!sk[70]) & (ld) & (!text_inx6x) & (g1749)) + ((!sk[70]) & (ld) & (text_inx6x) & (!g1749)) + ((!sk[70]) & (ld) & (text_inx6x) & (g1749)) + ((sk[70]) & (!ld) & (!text_inx6x) & (g1749)) + ((sk[70]) & (!ld) & (text_inx6x) & (g1749)) + ((sk[70]) & (ld) & (text_inx6x) & (!g1749)) + ((sk[70]) & (ld) & (text_inx6x) & (g1749)));
	assign g1750 = (((!g190) & (!g253) & (!g374) & (!g1163) & (g1658) & (!g1749)) + ((!g190) & (!g253) & (!g374) & (!g1163) & (g1658) & (g1749)) + ((!g190) & (!g253) & (!g374) & (g1163) & (!g1658) & (g1749)) + ((!g190) & (!g253) & (!g374) & (g1163) & (g1658) & (g1749)) + ((!g190) & (!g253) & (g374) & (!g1163) & (!g1658) & (!g1749)) + ((!g190) & (!g253) & (g374) & (!g1163) & (!g1658) & (g1749)) + ((!g190) & (!g253) & (g374) & (g1163) & (!g1658) & (g1749)) + ((!g190) & (!g253) & (g374) & (g1163) & (g1658) & (g1749)) + ((!g190) & (g253) & (!g374) & (!g1163) & (!g1658) & (!g1749)) + ((!g190) & (g253) & (!g374) & (!g1163) & (!g1658) & (g1749)) + ((!g190) & (g253) & (!g374) & (g1163) & (!g1658) & (g1749)) + ((!g190) & (g253) & (!g374) & (g1163) & (g1658) & (g1749)) + ((!g190) & (g253) & (g374) & (!g1163) & (g1658) & (!g1749)) + ((!g190) & (g253) & (g374) & (!g1163) & (g1658) & (g1749)) + ((!g190) & (g253) & (g374) & (g1163) & (!g1658) & (g1749)) + ((!g190) & (g253) & (g374) & (g1163) & (g1658) & (g1749)) + ((g190) & (!g253) & (!g374) & (!g1163) & (!g1658) & (!g1749)) + ((g190) & (!g253) & (!g374) & (!g1163) & (!g1658) & (g1749)) + ((g190) & (!g253) & (!g374) & (g1163) & (!g1658) & (!g1749)) + ((g190) & (!g253) & (!g374) & (g1163) & (g1658) & (!g1749)) + ((g190) & (!g253) & (g374) & (!g1163) & (g1658) & (!g1749)) + ((g190) & (!g253) & (g374) & (!g1163) & (g1658) & (g1749)) + ((g190) & (!g253) & (g374) & (g1163) & (!g1658) & (!g1749)) + ((g190) & (!g253) & (g374) & (g1163) & (g1658) & (!g1749)) + ((g190) & (g253) & (!g374) & (!g1163) & (g1658) & (!g1749)) + ((g190) & (g253) & (!g374) & (!g1163) & (g1658) & (g1749)) + ((g190) & (g253) & (!g374) & (g1163) & (!g1658) & (!g1749)) + ((g190) & (g253) & (!g374) & (g1163) & (g1658) & (!g1749)) + ((g190) & (g253) & (g374) & (!g1163) & (!g1658) & (!g1749)) + ((g190) & (g253) & (g374) & (!g1163) & (!g1658) & (g1749)) + ((g190) & (g253) & (g374) & (g1163) & (!g1658) & (!g1749)) + ((g190) & (g253) & (g374) & (g1163) & (g1658) & (!g1749)));
	assign g2183 = (((!sk[72]) & (!ld) & (text_inx5x) & (!g1751)) + ((!sk[72]) & (!ld) & (text_inx5x) & (g1751)) + ((!sk[72]) & (ld) & (!text_inx5x) & (g1751)) + ((!sk[72]) & (ld) & (text_inx5x) & (!g1751)) + ((!sk[72]) & (ld) & (text_inx5x) & (g1751)) + ((sk[72]) & (!ld) & (!text_inx5x) & (g1751)) + ((sk[72]) & (!ld) & (text_inx5x) & (g1751)) + ((sk[72]) & (ld) & (text_inx5x) & (!g1751)) + ((sk[72]) & (ld) & (text_inx5x) & (g1751)));
	assign g1752 = (((!g183) & (!g246) & (!g367) & (!g1163) & (g1661) & (!g1751)) + ((!g183) & (!g246) & (!g367) & (!g1163) & (g1661) & (g1751)) + ((!g183) & (!g246) & (!g367) & (g1163) & (!g1661) & (g1751)) + ((!g183) & (!g246) & (!g367) & (g1163) & (g1661) & (g1751)) + ((!g183) & (!g246) & (g367) & (!g1163) & (!g1661) & (!g1751)) + ((!g183) & (!g246) & (g367) & (!g1163) & (!g1661) & (g1751)) + ((!g183) & (!g246) & (g367) & (g1163) & (!g1661) & (g1751)) + ((!g183) & (!g246) & (g367) & (g1163) & (g1661) & (g1751)) + ((!g183) & (g246) & (!g367) & (!g1163) & (!g1661) & (!g1751)) + ((!g183) & (g246) & (!g367) & (!g1163) & (!g1661) & (g1751)) + ((!g183) & (g246) & (!g367) & (g1163) & (!g1661) & (g1751)) + ((!g183) & (g246) & (!g367) & (g1163) & (g1661) & (g1751)) + ((!g183) & (g246) & (g367) & (!g1163) & (g1661) & (!g1751)) + ((!g183) & (g246) & (g367) & (!g1163) & (g1661) & (g1751)) + ((!g183) & (g246) & (g367) & (g1163) & (!g1661) & (g1751)) + ((!g183) & (g246) & (g367) & (g1163) & (g1661) & (g1751)) + ((g183) & (!g246) & (!g367) & (!g1163) & (!g1661) & (!g1751)) + ((g183) & (!g246) & (!g367) & (!g1163) & (!g1661) & (g1751)) + ((g183) & (!g246) & (!g367) & (g1163) & (!g1661) & (!g1751)) + ((g183) & (!g246) & (!g367) & (g1163) & (g1661) & (!g1751)) + ((g183) & (!g246) & (g367) & (!g1163) & (g1661) & (!g1751)) + ((g183) & (!g246) & (g367) & (!g1163) & (g1661) & (g1751)) + ((g183) & (!g246) & (g367) & (g1163) & (!g1661) & (!g1751)) + ((g183) & (!g246) & (g367) & (g1163) & (g1661) & (!g1751)) + ((g183) & (g246) & (!g367) & (!g1163) & (g1661) & (!g1751)) + ((g183) & (g246) & (!g367) & (!g1163) & (g1661) & (g1751)) + ((g183) & (g246) & (!g367) & (g1163) & (!g1661) & (!g1751)) + ((g183) & (g246) & (!g367) & (g1163) & (g1661) & (!g1751)) + ((g183) & (g246) & (g367) & (!g1163) & (!g1661) & (!g1751)) + ((g183) & (g246) & (g367) & (!g1163) & (!g1661) & (g1751)) + ((g183) & (g246) & (g367) & (g1163) & (!g1661) & (!g1751)) + ((g183) & (g246) & (g367) & (g1163) & (g1661) & (!g1751)));
	assign g2184 = (((!ld) & (!text_inx4x) & (sk[74]) & (g1753)) + ((!ld) & (text_inx4x) & (!sk[74]) & (!g1753)) + ((!ld) & (text_inx4x) & (!sk[74]) & (g1753)) + ((!ld) & (text_inx4x) & (sk[74]) & (g1753)) + ((ld) & (!text_inx4x) & (!sk[74]) & (g1753)) + ((ld) & (text_inx4x) & (!sk[74]) & (!g1753)) + ((ld) & (text_inx4x) & (!sk[74]) & (g1753)) + ((ld) & (text_inx4x) & (sk[74]) & (!g1753)) + ((ld) & (text_inx4x) & (sk[74]) & (g1753)));
	assign g1754 = (((!g168) & (!g176) & (!g196) & (!g239) & (!g360) & (g388)) + ((!g168) & (!g176) & (!g196) & (!g239) & (g360) & (!g388)) + ((!g168) & (!g176) & (!g196) & (g239) & (!g360) & (!g388)) + ((!g168) & (!g176) & (!g196) & (g239) & (g360) & (g388)) + ((!g168) & (!g176) & (g196) & (!g239) & (!g360) & (!g388)) + ((!g168) & (!g176) & (g196) & (!g239) & (g360) & (g388)) + ((!g168) & (!g176) & (g196) & (g239) & (!g360) & (g388)) + ((!g168) & (!g176) & (g196) & (g239) & (g360) & (!g388)) + ((!g168) & (g176) & (!g196) & (!g239) & (!g360) & (!g388)) + ((!g168) & (g176) & (!g196) & (!g239) & (g360) & (g388)) + ((!g168) & (g176) & (!g196) & (g239) & (!g360) & (g388)) + ((!g168) & (g176) & (!g196) & (g239) & (g360) & (!g388)) + ((!g168) & (g176) & (g196) & (!g239) & (!g360) & (g388)) + ((!g168) & (g176) & (g196) & (!g239) & (g360) & (!g388)) + ((!g168) & (g176) & (g196) & (g239) & (!g360) & (!g388)) + ((!g168) & (g176) & (g196) & (g239) & (g360) & (g388)) + ((g168) & (!g176) & (!g196) & (!g239) & (!g360) & (!g388)) + ((g168) & (!g176) & (!g196) & (!g239) & (g360) & (g388)) + ((g168) & (!g176) & (!g196) & (g239) & (!g360) & (g388)) + ((g168) & (!g176) & (!g196) & (g239) & (g360) & (!g388)) + ((g168) & (!g176) & (g196) & (!g239) & (!g360) & (g388)) + ((g168) & (!g176) & (g196) & (!g239) & (g360) & (!g388)) + ((g168) & (!g176) & (g196) & (g239) & (!g360) & (!g388)) + ((g168) & (!g176) & (g196) & (g239) & (g360) & (g388)) + ((g168) & (g176) & (!g196) & (!g239) & (!g360) & (g388)) + ((g168) & (g176) & (!g196) & (!g239) & (g360) & (!g388)) + ((g168) & (g176) & (!g196) & (g239) & (!g360) & (!g388)) + ((g168) & (g176) & (!g196) & (g239) & (g360) & (g388)) + ((g168) & (g176) & (g196) & (!g239) & (!g360) & (!g388)) + ((g168) & (g176) & (g196) & (!g239) & (g360) & (g388)) + ((g168) & (g176) & (g196) & (g239) & (!g360) & (g388)) + ((g168) & (g176) & (g196) & (g239) & (g360) & (!g388)));
	assign g1755 = (((!g176) & (!g1163) & (sk[76]) & (!g1664) & (!g1753) & (g1754)) + ((!g176) & (!g1163) & (sk[76]) & (!g1664) & (g1753) & (g1754)) + ((!g176) & (!g1163) & (sk[76]) & (g1664) & (!g1753) & (!g1754)) + ((!g176) & (!g1163) & (sk[76]) & (g1664) & (g1753) & (!g1754)) + ((!g176) & (g1163) & (!sk[76]) & (!g1664) & (!g1753) & (!g1754)) + ((!g176) & (g1163) & (!sk[76]) & (!g1664) & (!g1753) & (g1754)) + ((!g176) & (g1163) & (!sk[76]) & (!g1664) & (g1753) & (!g1754)) + ((!g176) & (g1163) & (!sk[76]) & (!g1664) & (g1753) & (g1754)) + ((!g176) & (g1163) & (!sk[76]) & (g1664) & (!g1753) & (!g1754)) + ((!g176) & (g1163) & (!sk[76]) & (g1664) & (!g1753) & (g1754)) + ((!g176) & (g1163) & (!sk[76]) & (g1664) & (g1753) & (!g1754)) + ((!g176) & (g1163) & (!sk[76]) & (g1664) & (g1753) & (g1754)) + ((!g176) & (g1163) & (sk[76]) & (!g1664) & (g1753) & (!g1754)) + ((!g176) & (g1163) & (sk[76]) & (!g1664) & (g1753) & (g1754)) + ((!g176) & (g1163) & (sk[76]) & (g1664) & (g1753) & (!g1754)) + ((!g176) & (g1163) & (sk[76]) & (g1664) & (g1753) & (g1754)) + ((g176) & (!g1163) & (!sk[76]) & (!g1664) & (!g1753) & (!g1754)) + ((g176) & (!g1163) & (!sk[76]) & (!g1664) & (!g1753) & (g1754)) + ((g176) & (!g1163) & (!sk[76]) & (!g1664) & (g1753) & (!g1754)) + ((g176) & (!g1163) & (!sk[76]) & (!g1664) & (g1753) & (g1754)) + ((g176) & (!g1163) & (!sk[76]) & (g1664) & (!g1753) & (!g1754)) + ((g176) & (!g1163) & (!sk[76]) & (g1664) & (!g1753) & (g1754)) + ((g176) & (!g1163) & (!sk[76]) & (g1664) & (g1753) & (!g1754)) + ((g176) & (!g1163) & (!sk[76]) & (g1664) & (g1753) & (g1754)) + ((g176) & (!g1163) & (sk[76]) & (!g1664) & (!g1753) & (g1754)) + ((g176) & (!g1163) & (sk[76]) & (!g1664) & (g1753) & (g1754)) + ((g176) & (!g1163) & (sk[76]) & (g1664) & (!g1753) & (!g1754)) + ((g176) & (!g1163) & (sk[76]) & (g1664) & (g1753) & (!g1754)) + ((g176) & (g1163) & (!sk[76]) & (!g1664) & (!g1753) & (!g1754)) + ((g176) & (g1163) & (!sk[76]) & (!g1664) & (!g1753) & (g1754)) + ((g176) & (g1163) & (!sk[76]) & (!g1664) & (g1753) & (!g1754)) + ((g176) & (g1163) & (!sk[76]) & (!g1664) & (g1753) & (g1754)) + ((g176) & (g1163) & (!sk[76]) & (g1664) & (!g1753) & (!g1754)) + ((g176) & (g1163) & (!sk[76]) & (g1664) & (!g1753) & (g1754)) + ((g176) & (g1163) & (!sk[76]) & (g1664) & (g1753) & (!g1754)) + ((g176) & (g1163) & (!sk[76]) & (g1664) & (g1753) & (g1754)) + ((g176) & (g1163) & (sk[76]) & (!g1664) & (!g1753) & (!g1754)) + ((g176) & (g1163) & (sk[76]) & (!g1664) & (!g1753) & (g1754)) + ((g176) & (g1163) & (sk[76]) & (g1664) & (!g1753) & (!g1754)) + ((g176) & (g1163) & (sk[76]) & (g1664) & (!g1753) & (g1754)));
	assign g2185 = (((!ld) & (!sk[77]) & (text_inx7x) & (!g1756)) + ((!ld) & (!sk[77]) & (text_inx7x) & (g1756)) + ((!ld) & (sk[77]) & (!text_inx7x) & (g1756)) + ((!ld) & (sk[77]) & (text_inx7x) & (g1756)) + ((ld) & (!sk[77]) & (!text_inx7x) & (g1756)) + ((ld) & (!sk[77]) & (text_inx7x) & (!g1756)) + ((ld) & (!sk[77]) & (text_inx7x) & (g1756)) + ((ld) & (sk[77]) & (text_inx7x) & (!g1756)) + ((ld) & (sk[77]) & (text_inx7x) & (g1756)));
	assign g1757 = (((!ld) & (!g916) & (g1193) & (!sk[78]) & (!keyx96x)) + ((!ld) & (!g916) & (g1193) & (!sk[78]) & (keyx96x)) + ((!ld) & (!g916) & (g1193) & (sk[78]) & (!keyx96x)) + ((!ld) & (!g916) & (g1193) & (sk[78]) & (keyx96x)) + ((!ld) & (g916) & (!g1193) & (!sk[78]) & (!keyx96x)) + ((!ld) & (g916) & (!g1193) & (!sk[78]) & (keyx96x)) + ((!ld) & (g916) & (!g1193) & (sk[78]) & (!keyx96x)) + ((!ld) & (g916) & (!g1193) & (sk[78]) & (keyx96x)) + ((!ld) & (g916) & (g1193) & (!sk[78]) & (!keyx96x)) + ((!ld) & (g916) & (g1193) & (!sk[78]) & (keyx96x)) + ((ld) & (!g916) & (!g1193) & (sk[78]) & (keyx96x)) + ((ld) & (!g916) & (g1193) & (!sk[78]) & (!keyx96x)) + ((ld) & (!g916) & (g1193) & (!sk[78]) & (keyx96x)) + ((ld) & (!g916) & (g1193) & (sk[78]) & (keyx96x)) + ((ld) & (g916) & (!g1193) & (!sk[78]) & (!keyx96x)) + ((ld) & (g916) & (!g1193) & (!sk[78]) & (keyx96x)) + ((ld) & (g916) & (!g1193) & (sk[78]) & (keyx96x)) + ((ld) & (g916) & (g1193) & (!sk[78]) & (!keyx96x)) + ((ld) & (g916) & (g1193) & (!sk[78]) & (keyx96x)) + ((ld) & (g916) & (g1193) & (sk[78]) & (keyx96x)));
	assign g1758 = (((!ld) & (!g923) & (!sk[79]) & (g1200) & (!keyx97x)) + ((!ld) & (!g923) & (!sk[79]) & (g1200) & (keyx97x)) + ((!ld) & (!g923) & (sk[79]) & (g1200) & (!keyx97x)) + ((!ld) & (!g923) & (sk[79]) & (g1200) & (keyx97x)) + ((!ld) & (g923) & (!sk[79]) & (!g1200) & (!keyx97x)) + ((!ld) & (g923) & (!sk[79]) & (!g1200) & (keyx97x)) + ((!ld) & (g923) & (!sk[79]) & (g1200) & (!keyx97x)) + ((!ld) & (g923) & (!sk[79]) & (g1200) & (keyx97x)) + ((!ld) & (g923) & (sk[79]) & (!g1200) & (!keyx97x)) + ((!ld) & (g923) & (sk[79]) & (!g1200) & (keyx97x)) + ((ld) & (!g923) & (!sk[79]) & (g1200) & (!keyx97x)) + ((ld) & (!g923) & (!sk[79]) & (g1200) & (keyx97x)) + ((ld) & (!g923) & (sk[79]) & (!g1200) & (keyx97x)) + ((ld) & (!g923) & (sk[79]) & (g1200) & (keyx97x)) + ((ld) & (g923) & (!sk[79]) & (!g1200) & (!keyx97x)) + ((ld) & (g923) & (!sk[79]) & (!g1200) & (keyx97x)) + ((ld) & (g923) & (!sk[79]) & (g1200) & (!keyx97x)) + ((ld) & (g923) & (!sk[79]) & (g1200) & (keyx97x)) + ((ld) & (g923) & (sk[79]) & (!g1200) & (keyx97x)) + ((ld) & (g923) & (sk[79]) & (g1200) & (keyx97x)));
	assign g1759 = (((!ld) & (!g930) & (!sk[80]) & (g1207) & (!keyx98x)) + ((!ld) & (!g930) & (!sk[80]) & (g1207) & (keyx98x)) + ((!ld) & (!g930) & (sk[80]) & (g1207) & (!keyx98x)) + ((!ld) & (!g930) & (sk[80]) & (g1207) & (keyx98x)) + ((!ld) & (g930) & (!sk[80]) & (!g1207) & (!keyx98x)) + ((!ld) & (g930) & (!sk[80]) & (!g1207) & (keyx98x)) + ((!ld) & (g930) & (!sk[80]) & (g1207) & (!keyx98x)) + ((!ld) & (g930) & (!sk[80]) & (g1207) & (keyx98x)) + ((!ld) & (g930) & (sk[80]) & (!g1207) & (!keyx98x)) + ((!ld) & (g930) & (sk[80]) & (!g1207) & (keyx98x)) + ((ld) & (!g930) & (!sk[80]) & (g1207) & (!keyx98x)) + ((ld) & (!g930) & (!sk[80]) & (g1207) & (keyx98x)) + ((ld) & (!g930) & (sk[80]) & (!g1207) & (keyx98x)) + ((ld) & (!g930) & (sk[80]) & (g1207) & (keyx98x)) + ((ld) & (g930) & (!sk[80]) & (!g1207) & (!keyx98x)) + ((ld) & (g930) & (!sk[80]) & (!g1207) & (keyx98x)) + ((ld) & (g930) & (!sk[80]) & (g1207) & (!keyx98x)) + ((ld) & (g930) & (!sk[80]) & (g1207) & (keyx98x)) + ((ld) & (g930) & (sk[80]) & (!g1207) & (keyx98x)) + ((ld) & (g930) & (sk[80]) & (g1207) & (keyx98x)));
	assign g1760 = (((!sk[81]) & (!ld) & (!g937) & (g1214) & (!keyx99x)) + ((!sk[81]) & (!ld) & (!g937) & (g1214) & (keyx99x)) + ((!sk[81]) & (!ld) & (g937) & (!g1214) & (!keyx99x)) + ((!sk[81]) & (!ld) & (g937) & (!g1214) & (keyx99x)) + ((!sk[81]) & (!ld) & (g937) & (g1214) & (!keyx99x)) + ((!sk[81]) & (!ld) & (g937) & (g1214) & (keyx99x)) + ((!sk[81]) & (ld) & (!g937) & (g1214) & (!keyx99x)) + ((!sk[81]) & (ld) & (!g937) & (g1214) & (keyx99x)) + ((!sk[81]) & (ld) & (g937) & (!g1214) & (!keyx99x)) + ((!sk[81]) & (ld) & (g937) & (!g1214) & (keyx99x)) + ((!sk[81]) & (ld) & (g937) & (g1214) & (!keyx99x)) + ((!sk[81]) & (ld) & (g937) & (g1214) & (keyx99x)) + ((sk[81]) & (!ld) & (!g937) & (g1214) & (!keyx99x)) + ((sk[81]) & (!ld) & (!g937) & (g1214) & (keyx99x)) + ((sk[81]) & (!ld) & (g937) & (!g1214) & (!keyx99x)) + ((sk[81]) & (!ld) & (g937) & (!g1214) & (keyx99x)) + ((sk[81]) & (ld) & (!g937) & (!g1214) & (keyx99x)) + ((sk[81]) & (ld) & (!g937) & (g1214) & (keyx99x)) + ((sk[81]) & (ld) & (g937) & (!g1214) & (keyx99x)) + ((sk[81]) & (ld) & (g937) & (g1214) & (keyx99x)));
	assign g1761 = (((!ld) & (!g944) & (!sk[82]) & (g1221) & (!keyx100x)) + ((!ld) & (!g944) & (!sk[82]) & (g1221) & (keyx100x)) + ((!ld) & (!g944) & (sk[82]) & (g1221) & (!keyx100x)) + ((!ld) & (!g944) & (sk[82]) & (g1221) & (keyx100x)) + ((!ld) & (g944) & (!sk[82]) & (!g1221) & (!keyx100x)) + ((!ld) & (g944) & (!sk[82]) & (!g1221) & (keyx100x)) + ((!ld) & (g944) & (!sk[82]) & (g1221) & (!keyx100x)) + ((!ld) & (g944) & (!sk[82]) & (g1221) & (keyx100x)) + ((!ld) & (g944) & (sk[82]) & (!g1221) & (!keyx100x)) + ((!ld) & (g944) & (sk[82]) & (!g1221) & (keyx100x)) + ((ld) & (!g944) & (!sk[82]) & (g1221) & (!keyx100x)) + ((ld) & (!g944) & (!sk[82]) & (g1221) & (keyx100x)) + ((ld) & (!g944) & (sk[82]) & (!g1221) & (keyx100x)) + ((ld) & (!g944) & (sk[82]) & (g1221) & (keyx100x)) + ((ld) & (g944) & (!sk[82]) & (!g1221) & (!keyx100x)) + ((ld) & (g944) & (!sk[82]) & (!g1221) & (keyx100x)) + ((ld) & (g944) & (!sk[82]) & (g1221) & (!keyx100x)) + ((ld) & (g944) & (!sk[82]) & (g1221) & (keyx100x)) + ((ld) & (g944) & (sk[82]) & (!g1221) & (keyx100x)) + ((ld) & (g944) & (sk[82]) & (g1221) & (keyx100x)));
	assign g1762 = (((!sk[83]) & (!ld) & (!g951) & (g1228) & (!keyx101x)) + ((!sk[83]) & (!ld) & (!g951) & (g1228) & (keyx101x)) + ((!sk[83]) & (!ld) & (g951) & (!g1228) & (!keyx101x)) + ((!sk[83]) & (!ld) & (g951) & (!g1228) & (keyx101x)) + ((!sk[83]) & (!ld) & (g951) & (g1228) & (!keyx101x)) + ((!sk[83]) & (!ld) & (g951) & (g1228) & (keyx101x)) + ((!sk[83]) & (ld) & (!g951) & (g1228) & (!keyx101x)) + ((!sk[83]) & (ld) & (!g951) & (g1228) & (keyx101x)) + ((!sk[83]) & (ld) & (g951) & (!g1228) & (!keyx101x)) + ((!sk[83]) & (ld) & (g951) & (!g1228) & (keyx101x)) + ((!sk[83]) & (ld) & (g951) & (g1228) & (!keyx101x)) + ((!sk[83]) & (ld) & (g951) & (g1228) & (keyx101x)) + ((sk[83]) & (!ld) & (!g951) & (g1228) & (!keyx101x)) + ((sk[83]) & (!ld) & (!g951) & (g1228) & (keyx101x)) + ((sk[83]) & (!ld) & (g951) & (!g1228) & (!keyx101x)) + ((sk[83]) & (!ld) & (g951) & (!g1228) & (keyx101x)) + ((sk[83]) & (ld) & (!g951) & (!g1228) & (keyx101x)) + ((sk[83]) & (ld) & (!g951) & (g1228) & (keyx101x)) + ((sk[83]) & (ld) & (g951) & (!g1228) & (keyx101x)) + ((sk[83]) & (ld) & (g951) & (g1228) & (keyx101x)));
	assign g1763 = (((!ld) & (!g958) & (g1235) & (!sk[84]) & (!keyx102x)) + ((!ld) & (!g958) & (g1235) & (!sk[84]) & (keyx102x)) + ((!ld) & (!g958) & (g1235) & (sk[84]) & (!keyx102x)) + ((!ld) & (!g958) & (g1235) & (sk[84]) & (keyx102x)) + ((!ld) & (g958) & (!g1235) & (!sk[84]) & (!keyx102x)) + ((!ld) & (g958) & (!g1235) & (!sk[84]) & (keyx102x)) + ((!ld) & (g958) & (!g1235) & (sk[84]) & (!keyx102x)) + ((!ld) & (g958) & (!g1235) & (sk[84]) & (keyx102x)) + ((!ld) & (g958) & (g1235) & (!sk[84]) & (!keyx102x)) + ((!ld) & (g958) & (g1235) & (!sk[84]) & (keyx102x)) + ((ld) & (!g958) & (!g1235) & (sk[84]) & (keyx102x)) + ((ld) & (!g958) & (g1235) & (!sk[84]) & (!keyx102x)) + ((ld) & (!g958) & (g1235) & (!sk[84]) & (keyx102x)) + ((ld) & (!g958) & (g1235) & (sk[84]) & (keyx102x)) + ((ld) & (g958) & (!g1235) & (!sk[84]) & (!keyx102x)) + ((ld) & (g958) & (!g1235) & (!sk[84]) & (keyx102x)) + ((ld) & (g958) & (!g1235) & (sk[84]) & (keyx102x)) + ((ld) & (g958) & (g1235) & (!sk[84]) & (!keyx102x)) + ((ld) & (g958) & (g1235) & (!sk[84]) & (keyx102x)) + ((ld) & (g958) & (g1235) & (sk[84]) & (keyx102x)));
	assign g1764 = (((!ld) & (!sk[85]) & (!g965) & (g1242) & (!keyx103x)) + ((!ld) & (!sk[85]) & (!g965) & (g1242) & (keyx103x)) + ((!ld) & (!sk[85]) & (g965) & (!g1242) & (!keyx103x)) + ((!ld) & (!sk[85]) & (g965) & (!g1242) & (keyx103x)) + ((!ld) & (!sk[85]) & (g965) & (g1242) & (!keyx103x)) + ((!ld) & (!sk[85]) & (g965) & (g1242) & (keyx103x)) + ((!ld) & (sk[85]) & (!g965) & (g1242) & (!keyx103x)) + ((!ld) & (sk[85]) & (!g965) & (g1242) & (keyx103x)) + ((!ld) & (sk[85]) & (g965) & (!g1242) & (!keyx103x)) + ((!ld) & (sk[85]) & (g965) & (!g1242) & (keyx103x)) + ((ld) & (!sk[85]) & (!g965) & (g1242) & (!keyx103x)) + ((ld) & (!sk[85]) & (!g965) & (g1242) & (keyx103x)) + ((ld) & (!sk[85]) & (g965) & (!g1242) & (!keyx103x)) + ((ld) & (!sk[85]) & (g965) & (!g1242) & (keyx103x)) + ((ld) & (!sk[85]) & (g965) & (g1242) & (!keyx103x)) + ((ld) & (!sk[85]) & (g965) & (g1242) & (keyx103x)) + ((ld) & (sk[85]) & (!g965) & (!g1242) & (keyx103x)) + ((ld) & (sk[85]) & (!g965) & (g1242) & (keyx103x)) + ((ld) & (sk[85]) & (g965) & (!g1242) & (keyx103x)) + ((ld) & (sk[85]) & (g965) & (g1242) & (keyx103x)));
	assign g2186 = (((!ld) & (!sk[86]) & (text_inx40x) & (!g1765)) + ((!ld) & (!sk[86]) & (text_inx40x) & (g1765)) + ((!ld) & (sk[86]) & (!text_inx40x) & (g1765)) + ((!ld) & (sk[86]) & (text_inx40x) & (g1765)) + ((ld) & (!sk[86]) & (!text_inx40x) & (g1765)) + ((ld) & (!sk[86]) & (text_inx40x) & (!g1765)) + ((ld) & (!sk[86]) & (text_inx40x) & (g1765)) + ((ld) & (sk[86]) & (text_inx40x) & (!g1765)) + ((ld) & (sk[86]) & (text_inx40x) & (g1765)));
	assign g1766 = (((!sk[87]) & (!g403) & (!g452) & (g468) & (!g516)) + ((!sk[87]) & (!g403) & (!g452) & (g468) & (g516)) + ((!sk[87]) & (!g403) & (g452) & (!g468) & (!g516)) + ((!sk[87]) & (!g403) & (g452) & (!g468) & (g516)) + ((!sk[87]) & (!g403) & (g452) & (g468) & (!g516)) + ((!sk[87]) & (!g403) & (g452) & (g468) & (g516)) + ((!sk[87]) & (g403) & (!g452) & (g468) & (!g516)) + ((!sk[87]) & (g403) & (!g452) & (g468) & (g516)) + ((!sk[87]) & (g403) & (g452) & (!g468) & (!g516)) + ((!sk[87]) & (g403) & (g452) & (!g468) & (g516)) + ((!sk[87]) & (g403) & (g452) & (g468) & (!g516)) + ((!sk[87]) & (g403) & (g452) & (g468) & (g516)) + ((sk[87]) & (!g403) & (!g452) & (!g468) & (g516)) + ((sk[87]) & (!g403) & (!g452) & (g468) & (!g516)) + ((sk[87]) & (!g403) & (g452) & (!g468) & (!g516)) + ((sk[87]) & (!g403) & (g452) & (g468) & (g516)) + ((sk[87]) & (g403) & (!g452) & (!g468) & (!g516)) + ((sk[87]) & (g403) & (!g452) & (g468) & (g516)) + ((sk[87]) & (g403) & (g452) & (!g468) & (g516)) + ((sk[87]) & (g403) & (g452) & (g468) & (!g516)));
	assign g1767 = (((!g468) & (!g531) & (!g595) & (!g1163) & (!g1765) & (g1766)) + ((!g468) & (!g531) & (!g595) & (!g1163) & (g1765) & (g1766)) + ((!g468) & (!g531) & (!g595) & (g1163) & (g1765) & (!g1766)) + ((!g468) & (!g531) & (!g595) & (g1163) & (g1765) & (g1766)) + ((!g468) & (!g531) & (g595) & (!g1163) & (!g1765) & (!g1766)) + ((!g468) & (!g531) & (g595) & (!g1163) & (g1765) & (!g1766)) + ((!g468) & (!g531) & (g595) & (g1163) & (g1765) & (!g1766)) + ((!g468) & (!g531) & (g595) & (g1163) & (g1765) & (g1766)) + ((!g468) & (g531) & (!g595) & (!g1163) & (!g1765) & (!g1766)) + ((!g468) & (g531) & (!g595) & (!g1163) & (g1765) & (!g1766)) + ((!g468) & (g531) & (!g595) & (g1163) & (g1765) & (!g1766)) + ((!g468) & (g531) & (!g595) & (g1163) & (g1765) & (g1766)) + ((!g468) & (g531) & (g595) & (!g1163) & (!g1765) & (g1766)) + ((!g468) & (g531) & (g595) & (!g1163) & (g1765) & (g1766)) + ((!g468) & (g531) & (g595) & (g1163) & (g1765) & (!g1766)) + ((!g468) & (g531) & (g595) & (g1163) & (g1765) & (g1766)) + ((g468) & (!g531) & (!g595) & (!g1163) & (!g1765) & (g1766)) + ((g468) & (!g531) & (!g595) & (!g1163) & (g1765) & (g1766)) + ((g468) & (!g531) & (!g595) & (g1163) & (!g1765) & (!g1766)) + ((g468) & (!g531) & (!g595) & (g1163) & (!g1765) & (g1766)) + ((g468) & (!g531) & (g595) & (!g1163) & (!g1765) & (!g1766)) + ((g468) & (!g531) & (g595) & (!g1163) & (g1765) & (!g1766)) + ((g468) & (!g531) & (g595) & (g1163) & (!g1765) & (!g1766)) + ((g468) & (!g531) & (g595) & (g1163) & (!g1765) & (g1766)) + ((g468) & (g531) & (!g595) & (!g1163) & (!g1765) & (!g1766)) + ((g468) & (g531) & (!g595) & (!g1163) & (g1765) & (!g1766)) + ((g468) & (g531) & (!g595) & (g1163) & (!g1765) & (!g1766)) + ((g468) & (g531) & (!g595) & (g1163) & (!g1765) & (g1766)) + ((g468) & (g531) & (g595) & (!g1163) & (!g1765) & (g1766)) + ((g468) & (g531) & (g595) & (!g1163) & (g1765) & (g1766)) + ((g468) & (g531) & (g595) & (g1163) & (!g1765) & (!g1766)) + ((g468) & (g531) & (g595) & (g1163) & (!g1765) & (g1766)));
	assign g2187 = (((!ld) & (!sk[89]) & (text_inx41x) & (!g1768)) + ((!ld) & (!sk[89]) & (text_inx41x) & (g1768)) + ((!ld) & (sk[89]) & (!text_inx41x) & (g1768)) + ((!ld) & (sk[89]) & (text_inx41x) & (g1768)) + ((ld) & (!sk[89]) & (!text_inx41x) & (g1768)) + ((ld) & (!sk[89]) & (text_inx41x) & (!g1768)) + ((ld) & (!sk[89]) & (text_inx41x) & (g1768)) + ((ld) & (sk[89]) & (text_inx41x) & (!g1768)) + ((ld) & (sk[89]) & (text_inx41x) & (g1768)));
	assign g2188 = (((!ld) & (!sk[90]) & (text_inx42x) & (!g1769)) + ((!ld) & (!sk[90]) & (text_inx42x) & (g1769)) + ((!ld) & (sk[90]) & (!text_inx42x) & (g1769)) + ((!ld) & (sk[90]) & (text_inx42x) & (g1769)) + ((ld) & (!sk[90]) & (!text_inx42x) & (g1769)) + ((ld) & (!sk[90]) & (text_inx42x) & (!g1769)) + ((ld) & (!sk[90]) & (text_inx42x) & (g1769)) + ((ld) & (sk[90]) & (text_inx42x) & (!g1769)) + ((ld) & (sk[90]) & (text_inx42x) & (g1769)));
	assign g1770 = (((!g417) & (!g474) & (!g482) & (!g1163) & (g1172) & (!g1769)) + ((!g417) & (!g474) & (!g482) & (!g1163) & (g1172) & (g1769)) + ((!g417) & (!g474) & (!g482) & (g1163) & (!g1172) & (g1769)) + ((!g417) & (!g474) & (!g482) & (g1163) & (g1172) & (g1769)) + ((!g417) & (!g474) & (g482) & (!g1163) & (!g1172) & (!g1769)) + ((!g417) & (!g474) & (g482) & (!g1163) & (!g1172) & (g1769)) + ((!g417) & (!g474) & (g482) & (g1163) & (!g1172) & (!g1769)) + ((!g417) & (!g474) & (g482) & (g1163) & (g1172) & (!g1769)) + ((!g417) & (g474) & (!g482) & (!g1163) & (!g1172) & (!g1769)) + ((!g417) & (g474) & (!g482) & (!g1163) & (!g1172) & (g1769)) + ((!g417) & (g474) & (!g482) & (g1163) & (!g1172) & (g1769)) + ((!g417) & (g474) & (!g482) & (g1163) & (g1172) & (g1769)) + ((!g417) & (g474) & (g482) & (!g1163) & (g1172) & (!g1769)) + ((!g417) & (g474) & (g482) & (!g1163) & (g1172) & (g1769)) + ((!g417) & (g474) & (g482) & (g1163) & (!g1172) & (!g1769)) + ((!g417) & (g474) & (g482) & (g1163) & (g1172) & (!g1769)) + ((g417) & (!g474) & (!g482) & (!g1163) & (!g1172) & (!g1769)) + ((g417) & (!g474) & (!g482) & (!g1163) & (!g1172) & (g1769)) + ((g417) & (!g474) & (!g482) & (g1163) & (!g1172) & (g1769)) + ((g417) & (!g474) & (!g482) & (g1163) & (g1172) & (g1769)) + ((g417) & (!g474) & (g482) & (!g1163) & (g1172) & (!g1769)) + ((g417) & (!g474) & (g482) & (!g1163) & (g1172) & (g1769)) + ((g417) & (!g474) & (g482) & (g1163) & (!g1172) & (!g1769)) + ((g417) & (!g474) & (g482) & (g1163) & (g1172) & (!g1769)) + ((g417) & (g474) & (!g482) & (!g1163) & (g1172) & (!g1769)) + ((g417) & (g474) & (!g482) & (!g1163) & (g1172) & (g1769)) + ((g417) & (g474) & (!g482) & (g1163) & (!g1172) & (g1769)) + ((g417) & (g474) & (!g482) & (g1163) & (g1172) & (g1769)) + ((g417) & (g474) & (g482) & (!g1163) & (!g1172) & (!g1769)) + ((g417) & (g474) & (g482) & (!g1163) & (!g1172) & (g1769)) + ((g417) & (g474) & (g482) & (g1163) & (!g1172) & (!g1769)) + ((g417) & (g474) & (g482) & (g1163) & (g1172) & (!g1769)));
	assign g2189 = (((!sk[92]) & (!ld) & (text_inx43x) & (!g1771)) + ((!sk[92]) & (!ld) & (text_inx43x) & (g1771)) + ((!sk[92]) & (ld) & (!text_inx43x) & (g1771)) + ((!sk[92]) & (ld) & (text_inx43x) & (!g1771)) + ((!sk[92]) & (ld) & (text_inx43x) & (g1771)) + ((sk[92]) & (!ld) & (!text_inx43x) & (g1771)) + ((sk[92]) & (!ld) & (text_inx43x) & (g1771)) + ((sk[92]) & (ld) & (text_inx43x) & (!g1771)) + ((sk[92]) & (ld) & (text_inx43x) & (g1771)));
	assign g1772 = (((!sk[93]) & (!g417) & (g452) & (!g489) & (!g516) & (!g552)) + ((!sk[93]) & (!g417) & (g452) & (!g489) & (!g516) & (g552)) + ((!sk[93]) & (!g417) & (g452) & (!g489) & (g516) & (!g552)) + ((!sk[93]) & (!g417) & (g452) & (!g489) & (g516) & (g552)) + ((!sk[93]) & (!g417) & (g452) & (g489) & (!g516) & (!g552)) + ((!sk[93]) & (!g417) & (g452) & (g489) & (!g516) & (g552)) + ((!sk[93]) & (!g417) & (g452) & (g489) & (g516) & (!g552)) + ((!sk[93]) & (!g417) & (g452) & (g489) & (g516) & (g552)) + ((!sk[93]) & (g417) & (!g452) & (!g489) & (!g516) & (!g552)) + ((!sk[93]) & (g417) & (!g452) & (!g489) & (!g516) & (g552)) + ((!sk[93]) & (g417) & (!g452) & (!g489) & (g516) & (!g552)) + ((!sk[93]) & (g417) & (!g452) & (!g489) & (g516) & (g552)) + ((!sk[93]) & (g417) & (!g452) & (g489) & (!g516) & (!g552)) + ((!sk[93]) & (g417) & (!g452) & (g489) & (!g516) & (g552)) + ((!sk[93]) & (g417) & (!g452) & (g489) & (g516) & (!g552)) + ((!sk[93]) & (g417) & (!g452) & (g489) & (g516) & (g552)) + ((!sk[93]) & (g417) & (g452) & (!g489) & (!g516) & (!g552)) + ((!sk[93]) & (g417) & (g452) & (!g489) & (!g516) & (g552)) + ((!sk[93]) & (g417) & (g452) & (!g489) & (g516) & (!g552)) + ((!sk[93]) & (g417) & (g452) & (!g489) & (g516) & (g552)) + ((!sk[93]) & (g417) & (g452) & (g489) & (!g516) & (!g552)) + ((!sk[93]) & (g417) & (g452) & (g489) & (!g516) & (g552)) + ((!sk[93]) & (g417) & (g452) & (g489) & (g516) & (!g552)) + ((!sk[93]) & (g417) & (g452) & (g489) & (g516) & (g552)) + ((sk[93]) & (!g417) & (!g452) & (!g489) & (!g516) & (g552)) + ((sk[93]) & (!g417) & (!g452) & (!g489) & (g516) & (!g552)) + ((sk[93]) & (!g417) & (!g452) & (g489) & (!g516) & (!g552)) + ((sk[93]) & (!g417) & (!g452) & (g489) & (g516) & (g552)) + ((sk[93]) & (!g417) & (g452) & (!g489) & (!g516) & (!g552)) + ((sk[93]) & (!g417) & (g452) & (!g489) & (g516) & (g552)) + ((sk[93]) & (!g417) & (g452) & (g489) & (!g516) & (g552)) + ((sk[93]) & (!g417) & (g452) & (g489) & (g516) & (!g552)) + ((sk[93]) & (g417) & (!g452) & (!g489) & (!g516) & (!g552)) + ((sk[93]) & (g417) & (!g452) & (!g489) & (g516) & (g552)) + ((sk[93]) & (g417) & (!g452) & (g489) & (!g516) & (g552)) + ((sk[93]) & (g417) & (!g452) & (g489) & (g516) & (!g552)) + ((sk[93]) & (g417) & (g452) & (!g489) & (!g516) & (g552)) + ((sk[93]) & (g417) & (g452) & (!g489) & (g516) & (!g552)) + ((sk[93]) & (g417) & (g452) & (g489) & (!g516) & (!g552)) + ((sk[93]) & (g417) & (g452) & (g489) & (g516) & (g552)));
	assign g1773 = (((!sk[94]) & (!g489) & (g1163) & (!g1686) & (!g1771) & (!g1772)) + ((!sk[94]) & (!g489) & (g1163) & (!g1686) & (!g1771) & (g1772)) + ((!sk[94]) & (!g489) & (g1163) & (!g1686) & (g1771) & (!g1772)) + ((!sk[94]) & (!g489) & (g1163) & (!g1686) & (g1771) & (g1772)) + ((!sk[94]) & (!g489) & (g1163) & (g1686) & (!g1771) & (!g1772)) + ((!sk[94]) & (!g489) & (g1163) & (g1686) & (!g1771) & (g1772)) + ((!sk[94]) & (!g489) & (g1163) & (g1686) & (g1771) & (!g1772)) + ((!sk[94]) & (!g489) & (g1163) & (g1686) & (g1771) & (g1772)) + ((!sk[94]) & (g489) & (!g1163) & (!g1686) & (!g1771) & (!g1772)) + ((!sk[94]) & (g489) & (!g1163) & (!g1686) & (!g1771) & (g1772)) + ((!sk[94]) & (g489) & (!g1163) & (!g1686) & (g1771) & (!g1772)) + ((!sk[94]) & (g489) & (!g1163) & (!g1686) & (g1771) & (g1772)) + ((!sk[94]) & (g489) & (!g1163) & (g1686) & (!g1771) & (!g1772)) + ((!sk[94]) & (g489) & (!g1163) & (g1686) & (!g1771) & (g1772)) + ((!sk[94]) & (g489) & (!g1163) & (g1686) & (g1771) & (!g1772)) + ((!sk[94]) & (g489) & (!g1163) & (g1686) & (g1771) & (g1772)) + ((!sk[94]) & (g489) & (g1163) & (!g1686) & (!g1771) & (!g1772)) + ((!sk[94]) & (g489) & (g1163) & (!g1686) & (!g1771) & (g1772)) + ((!sk[94]) & (g489) & (g1163) & (!g1686) & (g1771) & (!g1772)) + ((!sk[94]) & (g489) & (g1163) & (!g1686) & (g1771) & (g1772)) + ((!sk[94]) & (g489) & (g1163) & (g1686) & (!g1771) & (!g1772)) + ((!sk[94]) & (g489) & (g1163) & (g1686) & (!g1771) & (g1772)) + ((!sk[94]) & (g489) & (g1163) & (g1686) & (g1771) & (!g1772)) + ((!sk[94]) & (g489) & (g1163) & (g1686) & (g1771) & (g1772)) + ((sk[94]) & (!g489) & (!g1163) & (!g1686) & (!g1771) & (g1772)) + ((sk[94]) & (!g489) & (!g1163) & (!g1686) & (g1771) & (g1772)) + ((sk[94]) & (!g489) & (!g1163) & (g1686) & (!g1771) & (!g1772)) + ((sk[94]) & (!g489) & (!g1163) & (g1686) & (g1771) & (!g1772)) + ((sk[94]) & (!g489) & (g1163) & (!g1686) & (g1771) & (!g1772)) + ((sk[94]) & (!g489) & (g1163) & (!g1686) & (g1771) & (g1772)) + ((sk[94]) & (!g489) & (g1163) & (g1686) & (g1771) & (!g1772)) + ((sk[94]) & (!g489) & (g1163) & (g1686) & (g1771) & (g1772)) + ((sk[94]) & (g489) & (!g1163) & (!g1686) & (!g1771) & (g1772)) + ((sk[94]) & (g489) & (!g1163) & (!g1686) & (g1771) & (g1772)) + ((sk[94]) & (g489) & (!g1163) & (g1686) & (!g1771) & (!g1772)) + ((sk[94]) & (g489) & (!g1163) & (g1686) & (g1771) & (!g1772)) + ((sk[94]) & (g489) & (g1163) & (!g1686) & (!g1771) & (!g1772)) + ((sk[94]) & (g489) & (g1163) & (!g1686) & (!g1771) & (g1772)) + ((sk[94]) & (g489) & (g1163) & (g1686) & (!g1771) & (!g1772)) + ((sk[94]) & (g489) & (g1163) & (g1686) & (!g1771) & (g1772)));
	assign g2190 = (((!sk[95]) & (!ld) & (text_inx46x) & (!g1774)) + ((!sk[95]) & (!ld) & (text_inx46x) & (g1774)) + ((!sk[95]) & (ld) & (!text_inx46x) & (g1774)) + ((!sk[95]) & (ld) & (text_inx46x) & (!g1774)) + ((!sk[95]) & (ld) & (text_inx46x) & (g1774)) + ((sk[95]) & (!ld) & (!text_inx46x) & (g1774)) + ((sk[95]) & (!ld) & (text_inx46x) & (g1774)) + ((sk[95]) & (ld) & (text_inx46x) & (!g1774)) + ((sk[95]) & (ld) & (text_inx46x) & (g1774)));
	assign g1775 = (((!g445) & (!g502) & (!g510) & (!g1163) & (g1177) & (!g1774)) + ((!g445) & (!g502) & (!g510) & (!g1163) & (g1177) & (g1774)) + ((!g445) & (!g502) & (!g510) & (g1163) & (!g1177) & (g1774)) + ((!g445) & (!g502) & (!g510) & (g1163) & (g1177) & (g1774)) + ((!g445) & (!g502) & (g510) & (!g1163) & (!g1177) & (!g1774)) + ((!g445) & (!g502) & (g510) & (!g1163) & (!g1177) & (g1774)) + ((!g445) & (!g502) & (g510) & (g1163) & (!g1177) & (!g1774)) + ((!g445) & (!g502) & (g510) & (g1163) & (g1177) & (!g1774)) + ((!g445) & (g502) & (!g510) & (!g1163) & (!g1177) & (!g1774)) + ((!g445) & (g502) & (!g510) & (!g1163) & (!g1177) & (g1774)) + ((!g445) & (g502) & (!g510) & (g1163) & (!g1177) & (g1774)) + ((!g445) & (g502) & (!g510) & (g1163) & (g1177) & (g1774)) + ((!g445) & (g502) & (g510) & (!g1163) & (g1177) & (!g1774)) + ((!g445) & (g502) & (g510) & (!g1163) & (g1177) & (g1774)) + ((!g445) & (g502) & (g510) & (g1163) & (!g1177) & (!g1774)) + ((!g445) & (g502) & (g510) & (g1163) & (g1177) & (!g1774)) + ((g445) & (!g502) & (!g510) & (!g1163) & (!g1177) & (!g1774)) + ((g445) & (!g502) & (!g510) & (!g1163) & (!g1177) & (g1774)) + ((g445) & (!g502) & (!g510) & (g1163) & (!g1177) & (g1774)) + ((g445) & (!g502) & (!g510) & (g1163) & (g1177) & (g1774)) + ((g445) & (!g502) & (g510) & (!g1163) & (g1177) & (!g1774)) + ((g445) & (!g502) & (g510) & (!g1163) & (g1177) & (g1774)) + ((g445) & (!g502) & (g510) & (g1163) & (!g1177) & (!g1774)) + ((g445) & (!g502) & (g510) & (g1163) & (g1177) & (!g1774)) + ((g445) & (g502) & (!g510) & (!g1163) & (g1177) & (!g1774)) + ((g445) & (g502) & (!g510) & (!g1163) & (g1177) & (g1774)) + ((g445) & (g502) & (!g510) & (g1163) & (!g1177) & (g1774)) + ((g445) & (g502) & (!g510) & (g1163) & (g1177) & (g1774)) + ((g445) & (g502) & (g510) & (!g1163) & (!g1177) & (!g1774)) + ((g445) & (g502) & (g510) & (!g1163) & (!g1177) & (g1774)) + ((g445) & (g502) & (g510) & (g1163) & (!g1177) & (!g1774)) + ((g445) & (g502) & (g510) & (g1163) & (g1177) & (!g1774)));
	assign g2191 = (((!sk[97]) & (!ld) & (text_inx45x) & (!g1776)) + ((!sk[97]) & (!ld) & (text_inx45x) & (g1776)) + ((!sk[97]) & (ld) & (!text_inx45x) & (g1776)) + ((!sk[97]) & (ld) & (text_inx45x) & (!g1776)) + ((!sk[97]) & (ld) & (text_inx45x) & (g1776)) + ((sk[97]) & (!ld) & (!text_inx45x) & (g1776)) + ((sk[97]) & (!ld) & (text_inx45x) & (g1776)) + ((sk[97]) & (ld) & (text_inx45x) & (!g1776)) + ((sk[97]) & (ld) & (text_inx45x) & (g1776)));
	assign g1777 = (((!g438) & (!g495) & (!g503) & (!g1163) & (g1180) & (!g1776)) + ((!g438) & (!g495) & (!g503) & (!g1163) & (g1180) & (g1776)) + ((!g438) & (!g495) & (!g503) & (g1163) & (!g1180) & (g1776)) + ((!g438) & (!g495) & (!g503) & (g1163) & (g1180) & (g1776)) + ((!g438) & (!g495) & (g503) & (!g1163) & (!g1180) & (!g1776)) + ((!g438) & (!g495) & (g503) & (!g1163) & (!g1180) & (g1776)) + ((!g438) & (!g495) & (g503) & (g1163) & (!g1180) & (!g1776)) + ((!g438) & (!g495) & (g503) & (g1163) & (g1180) & (!g1776)) + ((!g438) & (g495) & (!g503) & (!g1163) & (!g1180) & (!g1776)) + ((!g438) & (g495) & (!g503) & (!g1163) & (!g1180) & (g1776)) + ((!g438) & (g495) & (!g503) & (g1163) & (!g1180) & (g1776)) + ((!g438) & (g495) & (!g503) & (g1163) & (g1180) & (g1776)) + ((!g438) & (g495) & (g503) & (!g1163) & (g1180) & (!g1776)) + ((!g438) & (g495) & (g503) & (!g1163) & (g1180) & (g1776)) + ((!g438) & (g495) & (g503) & (g1163) & (!g1180) & (!g1776)) + ((!g438) & (g495) & (g503) & (g1163) & (g1180) & (!g1776)) + ((g438) & (!g495) & (!g503) & (!g1163) & (!g1180) & (!g1776)) + ((g438) & (!g495) & (!g503) & (!g1163) & (!g1180) & (g1776)) + ((g438) & (!g495) & (!g503) & (g1163) & (!g1180) & (g1776)) + ((g438) & (!g495) & (!g503) & (g1163) & (g1180) & (g1776)) + ((g438) & (!g495) & (g503) & (!g1163) & (g1180) & (!g1776)) + ((g438) & (!g495) & (g503) & (!g1163) & (g1180) & (g1776)) + ((g438) & (!g495) & (g503) & (g1163) & (!g1180) & (!g1776)) + ((g438) & (!g495) & (g503) & (g1163) & (g1180) & (!g1776)) + ((g438) & (g495) & (!g503) & (!g1163) & (g1180) & (!g1776)) + ((g438) & (g495) & (!g503) & (!g1163) & (g1180) & (g1776)) + ((g438) & (g495) & (!g503) & (g1163) & (!g1180) & (g1776)) + ((g438) & (g495) & (!g503) & (g1163) & (g1180) & (g1776)) + ((g438) & (g495) & (g503) & (!g1163) & (!g1180) & (!g1776)) + ((g438) & (g495) & (g503) & (!g1163) & (!g1180) & (g1776)) + ((g438) & (g495) & (g503) & (g1163) & (!g1180) & (!g1776)) + ((g438) & (g495) & (g503) & (g1163) & (g1180) & (!g1776)));
	assign g2192 = (((!sk[99]) & (!ld) & (text_inx44x) & (!g1778)) + ((!sk[99]) & (!ld) & (text_inx44x) & (g1778)) + ((!sk[99]) & (ld) & (!text_inx44x) & (g1778)) + ((!sk[99]) & (ld) & (text_inx44x) & (!g1778)) + ((!sk[99]) & (ld) & (text_inx44x) & (g1778)) + ((sk[99]) & (!ld) & (!text_inx44x) & (g1778)) + ((sk[99]) & (!ld) & (text_inx44x) & (g1778)) + ((sk[99]) & (ld) & (text_inx44x) & (!g1778)) + ((sk[99]) & (ld) & (text_inx44x) & (g1778)));
	assign g1779 = (((!g431) & (!g452) & (!g488) & (!g496) & (sk[100]) & (g516)) + ((!g431) & (!g452) & (!g488) & (g496) & (sk[100]) & (!g516)) + ((!g431) & (!g452) & (g488) & (!g496) & (sk[100]) & (!g516)) + ((!g431) & (!g452) & (g488) & (g496) & (sk[100]) & (g516)) + ((!g431) & (g452) & (!g488) & (!g496) & (!sk[100]) & (!g516)) + ((!g431) & (g452) & (!g488) & (!g496) & (!sk[100]) & (g516)) + ((!g431) & (g452) & (!g488) & (!g496) & (sk[100]) & (!g516)) + ((!g431) & (g452) & (!g488) & (g496) & (!sk[100]) & (!g516)) + ((!g431) & (g452) & (!g488) & (g496) & (!sk[100]) & (g516)) + ((!g431) & (g452) & (!g488) & (g496) & (sk[100]) & (g516)) + ((!g431) & (g452) & (g488) & (!g496) & (!sk[100]) & (!g516)) + ((!g431) & (g452) & (g488) & (!g496) & (!sk[100]) & (g516)) + ((!g431) & (g452) & (g488) & (!g496) & (sk[100]) & (g516)) + ((!g431) & (g452) & (g488) & (g496) & (!sk[100]) & (!g516)) + ((!g431) & (g452) & (g488) & (g496) & (!sk[100]) & (g516)) + ((!g431) & (g452) & (g488) & (g496) & (sk[100]) & (!g516)) + ((g431) & (!g452) & (!g488) & (!g496) & (!sk[100]) & (!g516)) + ((g431) & (!g452) & (!g488) & (!g496) & (!sk[100]) & (g516)) + ((g431) & (!g452) & (!g488) & (!g496) & (sk[100]) & (!g516)) + ((g431) & (!g452) & (!g488) & (g496) & (!sk[100]) & (!g516)) + ((g431) & (!g452) & (!g488) & (g496) & (!sk[100]) & (g516)) + ((g431) & (!g452) & (!g488) & (g496) & (sk[100]) & (g516)) + ((g431) & (!g452) & (g488) & (!g496) & (!sk[100]) & (!g516)) + ((g431) & (!g452) & (g488) & (!g496) & (!sk[100]) & (g516)) + ((g431) & (!g452) & (g488) & (!g496) & (sk[100]) & (g516)) + ((g431) & (!g452) & (g488) & (g496) & (!sk[100]) & (!g516)) + ((g431) & (!g452) & (g488) & (g496) & (!sk[100]) & (g516)) + ((g431) & (!g452) & (g488) & (g496) & (sk[100]) & (!g516)) + ((g431) & (g452) & (!g488) & (!g496) & (!sk[100]) & (!g516)) + ((g431) & (g452) & (!g488) & (!g496) & (!sk[100]) & (g516)) + ((g431) & (g452) & (!g488) & (!g496) & (sk[100]) & (g516)) + ((g431) & (g452) & (!g488) & (g496) & (!sk[100]) & (!g516)) + ((g431) & (g452) & (!g488) & (g496) & (!sk[100]) & (g516)) + ((g431) & (g452) & (!g488) & (g496) & (sk[100]) & (!g516)) + ((g431) & (g452) & (g488) & (!g496) & (!sk[100]) & (!g516)) + ((g431) & (g452) & (g488) & (!g496) & (!sk[100]) & (g516)) + ((g431) & (g452) & (g488) & (!g496) & (sk[100]) & (!g516)) + ((g431) & (g452) & (g488) & (g496) & (!sk[100]) & (!g516)) + ((g431) & (g452) & (g488) & (g496) & (!sk[100]) & (g516)) + ((g431) & (g452) & (g488) & (g496) & (sk[100]) & (g516)));
	assign g1780 = (((!g496) & (!g1163) & (!g1183) & (!g1778) & (sk[101]) & (g1779)) + ((!g496) & (!g1163) & (!g1183) & (g1778) & (sk[101]) & (g1779)) + ((!g496) & (!g1163) & (g1183) & (!g1778) & (sk[101]) & (!g1779)) + ((!g496) & (!g1163) & (g1183) & (g1778) & (sk[101]) & (!g1779)) + ((!g496) & (g1163) & (!g1183) & (!g1778) & (!sk[101]) & (!g1779)) + ((!g496) & (g1163) & (!g1183) & (!g1778) & (!sk[101]) & (g1779)) + ((!g496) & (g1163) & (!g1183) & (g1778) & (!sk[101]) & (!g1779)) + ((!g496) & (g1163) & (!g1183) & (g1778) & (!sk[101]) & (g1779)) + ((!g496) & (g1163) & (!g1183) & (g1778) & (sk[101]) & (!g1779)) + ((!g496) & (g1163) & (!g1183) & (g1778) & (sk[101]) & (g1779)) + ((!g496) & (g1163) & (g1183) & (!g1778) & (!sk[101]) & (!g1779)) + ((!g496) & (g1163) & (g1183) & (!g1778) & (!sk[101]) & (g1779)) + ((!g496) & (g1163) & (g1183) & (g1778) & (!sk[101]) & (!g1779)) + ((!g496) & (g1163) & (g1183) & (g1778) & (!sk[101]) & (g1779)) + ((!g496) & (g1163) & (g1183) & (g1778) & (sk[101]) & (!g1779)) + ((!g496) & (g1163) & (g1183) & (g1778) & (sk[101]) & (g1779)) + ((g496) & (!g1163) & (!g1183) & (!g1778) & (!sk[101]) & (!g1779)) + ((g496) & (!g1163) & (!g1183) & (!g1778) & (!sk[101]) & (g1779)) + ((g496) & (!g1163) & (!g1183) & (!g1778) & (sk[101]) & (g1779)) + ((g496) & (!g1163) & (!g1183) & (g1778) & (!sk[101]) & (!g1779)) + ((g496) & (!g1163) & (!g1183) & (g1778) & (!sk[101]) & (g1779)) + ((g496) & (!g1163) & (!g1183) & (g1778) & (sk[101]) & (g1779)) + ((g496) & (!g1163) & (g1183) & (!g1778) & (!sk[101]) & (!g1779)) + ((g496) & (!g1163) & (g1183) & (!g1778) & (!sk[101]) & (g1779)) + ((g496) & (!g1163) & (g1183) & (!g1778) & (sk[101]) & (!g1779)) + ((g496) & (!g1163) & (g1183) & (g1778) & (!sk[101]) & (!g1779)) + ((g496) & (!g1163) & (g1183) & (g1778) & (!sk[101]) & (g1779)) + ((g496) & (!g1163) & (g1183) & (g1778) & (sk[101]) & (!g1779)) + ((g496) & (g1163) & (!g1183) & (!g1778) & (!sk[101]) & (!g1779)) + ((g496) & (g1163) & (!g1183) & (!g1778) & (!sk[101]) & (g1779)) + ((g496) & (g1163) & (!g1183) & (!g1778) & (sk[101]) & (!g1779)) + ((g496) & (g1163) & (!g1183) & (!g1778) & (sk[101]) & (g1779)) + ((g496) & (g1163) & (!g1183) & (g1778) & (!sk[101]) & (!g1779)) + ((g496) & (g1163) & (!g1183) & (g1778) & (!sk[101]) & (g1779)) + ((g496) & (g1163) & (g1183) & (!g1778) & (!sk[101]) & (!g1779)) + ((g496) & (g1163) & (g1183) & (!g1778) & (!sk[101]) & (g1779)) + ((g496) & (g1163) & (g1183) & (!g1778) & (sk[101]) & (!g1779)) + ((g496) & (g1163) & (g1183) & (!g1778) & (sk[101]) & (g1779)) + ((g496) & (g1163) & (g1183) & (g1778) & (!sk[101]) & (!g1779)) + ((g496) & (g1163) & (g1183) & (g1778) & (!sk[101]) & (g1779)));
	assign g2193 = (((!ld) & (!text_inx47x) & (sk[102]) & (g1781)) + ((!ld) & (text_inx47x) & (!sk[102]) & (!g1781)) + ((!ld) & (text_inx47x) & (!sk[102]) & (g1781)) + ((!ld) & (text_inx47x) & (sk[102]) & (g1781)) + ((ld) & (!text_inx47x) & (!sk[102]) & (g1781)) + ((ld) & (text_inx47x) & (!sk[102]) & (!g1781)) + ((ld) & (text_inx47x) & (!sk[102]) & (g1781)) + ((ld) & (text_inx47x) & (sk[102]) & (!g1781)) + ((ld) & (text_inx47x) & (sk[102]) & (g1781)));
	assign g1782 = (((!g452) & (!g509) & (!g517) & (!g1163) & (g1187) & (!g1781)) + ((!g452) & (!g509) & (!g517) & (!g1163) & (g1187) & (g1781)) + ((!g452) & (!g509) & (!g517) & (g1163) & (!g1187) & (g1781)) + ((!g452) & (!g509) & (!g517) & (g1163) & (g1187) & (g1781)) + ((!g452) & (!g509) & (g517) & (!g1163) & (!g1187) & (!g1781)) + ((!g452) & (!g509) & (g517) & (!g1163) & (!g1187) & (g1781)) + ((!g452) & (!g509) & (g517) & (g1163) & (!g1187) & (!g1781)) + ((!g452) & (!g509) & (g517) & (g1163) & (g1187) & (!g1781)) + ((!g452) & (g509) & (!g517) & (!g1163) & (!g1187) & (!g1781)) + ((!g452) & (g509) & (!g517) & (!g1163) & (!g1187) & (g1781)) + ((!g452) & (g509) & (!g517) & (g1163) & (!g1187) & (g1781)) + ((!g452) & (g509) & (!g517) & (g1163) & (g1187) & (g1781)) + ((!g452) & (g509) & (g517) & (!g1163) & (g1187) & (!g1781)) + ((!g452) & (g509) & (g517) & (!g1163) & (g1187) & (g1781)) + ((!g452) & (g509) & (g517) & (g1163) & (!g1187) & (!g1781)) + ((!g452) & (g509) & (g517) & (g1163) & (g1187) & (!g1781)) + ((g452) & (!g509) & (!g517) & (!g1163) & (!g1187) & (!g1781)) + ((g452) & (!g509) & (!g517) & (!g1163) & (!g1187) & (g1781)) + ((g452) & (!g509) & (!g517) & (g1163) & (!g1187) & (g1781)) + ((g452) & (!g509) & (!g517) & (g1163) & (g1187) & (g1781)) + ((g452) & (!g509) & (g517) & (!g1163) & (g1187) & (!g1781)) + ((g452) & (!g509) & (g517) & (!g1163) & (g1187) & (g1781)) + ((g452) & (!g509) & (g517) & (g1163) & (!g1187) & (!g1781)) + ((g452) & (!g509) & (g517) & (g1163) & (g1187) & (!g1781)) + ((g452) & (g509) & (!g517) & (!g1163) & (g1187) & (!g1781)) + ((g452) & (g509) & (!g517) & (!g1163) & (g1187) & (g1781)) + ((g452) & (g509) & (!g517) & (g1163) & (!g1187) & (g1781)) + ((g452) & (g509) & (!g517) & (g1163) & (g1187) & (g1781)) + ((g452) & (g509) & (g517) & (!g1163) & (!g1187) & (!g1781)) + ((g452) & (g509) & (g517) & (!g1163) & (!g1187) & (g1781)) + ((g452) & (g509) & (g517) & (g1163) & (!g1187) & (!g1781)) + ((g452) & (g509) & (g517) & (g1163) & (g1187) & (!g1781)));
	assign g1783 = (((!sk[104]) & (!ld) & (!g980) & (g1276) & (!keyx104x)) + ((!sk[104]) & (!ld) & (!g980) & (g1276) & (keyx104x)) + ((!sk[104]) & (!ld) & (g980) & (!g1276) & (!keyx104x)) + ((!sk[104]) & (!ld) & (g980) & (!g1276) & (keyx104x)) + ((!sk[104]) & (!ld) & (g980) & (g1276) & (!keyx104x)) + ((!sk[104]) & (!ld) & (g980) & (g1276) & (keyx104x)) + ((!sk[104]) & (ld) & (!g980) & (g1276) & (!keyx104x)) + ((!sk[104]) & (ld) & (!g980) & (g1276) & (keyx104x)) + ((!sk[104]) & (ld) & (g980) & (!g1276) & (!keyx104x)) + ((!sk[104]) & (ld) & (g980) & (!g1276) & (keyx104x)) + ((!sk[104]) & (ld) & (g980) & (g1276) & (!keyx104x)) + ((!sk[104]) & (ld) & (g980) & (g1276) & (keyx104x)) + ((sk[104]) & (!ld) & (!g980) & (g1276) & (!keyx104x)) + ((sk[104]) & (!ld) & (!g980) & (g1276) & (keyx104x)) + ((sk[104]) & (!ld) & (g980) & (!g1276) & (!keyx104x)) + ((sk[104]) & (!ld) & (g980) & (!g1276) & (keyx104x)) + ((sk[104]) & (ld) & (!g980) & (!g1276) & (keyx104x)) + ((sk[104]) & (ld) & (!g980) & (g1276) & (keyx104x)) + ((sk[104]) & (ld) & (g980) & (!g1276) & (keyx104x)) + ((sk[104]) & (ld) & (g980) & (g1276) & (keyx104x)));
	assign g1784 = (((!ld) & (!sk[105]) & (!g987) & (g1283) & (!keyx105x)) + ((!ld) & (!sk[105]) & (!g987) & (g1283) & (keyx105x)) + ((!ld) & (!sk[105]) & (g987) & (!g1283) & (!keyx105x)) + ((!ld) & (!sk[105]) & (g987) & (!g1283) & (keyx105x)) + ((!ld) & (!sk[105]) & (g987) & (g1283) & (!keyx105x)) + ((!ld) & (!sk[105]) & (g987) & (g1283) & (keyx105x)) + ((!ld) & (sk[105]) & (!g987) & (g1283) & (!keyx105x)) + ((!ld) & (sk[105]) & (!g987) & (g1283) & (keyx105x)) + ((!ld) & (sk[105]) & (g987) & (!g1283) & (!keyx105x)) + ((!ld) & (sk[105]) & (g987) & (!g1283) & (keyx105x)) + ((ld) & (!sk[105]) & (!g987) & (g1283) & (!keyx105x)) + ((ld) & (!sk[105]) & (!g987) & (g1283) & (keyx105x)) + ((ld) & (!sk[105]) & (g987) & (!g1283) & (!keyx105x)) + ((ld) & (!sk[105]) & (g987) & (!g1283) & (keyx105x)) + ((ld) & (!sk[105]) & (g987) & (g1283) & (!keyx105x)) + ((ld) & (!sk[105]) & (g987) & (g1283) & (keyx105x)) + ((ld) & (sk[105]) & (!g987) & (!g1283) & (keyx105x)) + ((ld) & (sk[105]) & (!g987) & (g1283) & (keyx105x)) + ((ld) & (sk[105]) & (g987) & (!g1283) & (keyx105x)) + ((ld) & (sk[105]) & (g987) & (g1283) & (keyx105x)));
	assign g1785 = (((!ld) & (!sk[106]) & (!g994) & (g1290) & (!keyx106x)) + ((!ld) & (!sk[106]) & (!g994) & (g1290) & (keyx106x)) + ((!ld) & (!sk[106]) & (g994) & (!g1290) & (!keyx106x)) + ((!ld) & (!sk[106]) & (g994) & (!g1290) & (keyx106x)) + ((!ld) & (!sk[106]) & (g994) & (g1290) & (!keyx106x)) + ((!ld) & (!sk[106]) & (g994) & (g1290) & (keyx106x)) + ((!ld) & (sk[106]) & (!g994) & (g1290) & (!keyx106x)) + ((!ld) & (sk[106]) & (!g994) & (g1290) & (keyx106x)) + ((!ld) & (sk[106]) & (g994) & (!g1290) & (!keyx106x)) + ((!ld) & (sk[106]) & (g994) & (!g1290) & (keyx106x)) + ((ld) & (!sk[106]) & (!g994) & (g1290) & (!keyx106x)) + ((ld) & (!sk[106]) & (!g994) & (g1290) & (keyx106x)) + ((ld) & (!sk[106]) & (g994) & (!g1290) & (!keyx106x)) + ((ld) & (!sk[106]) & (g994) & (!g1290) & (keyx106x)) + ((ld) & (!sk[106]) & (g994) & (g1290) & (!keyx106x)) + ((ld) & (!sk[106]) & (g994) & (g1290) & (keyx106x)) + ((ld) & (sk[106]) & (!g994) & (!g1290) & (keyx106x)) + ((ld) & (sk[106]) & (!g994) & (g1290) & (keyx106x)) + ((ld) & (sk[106]) & (g994) & (!g1290) & (keyx106x)) + ((ld) & (sk[106]) & (g994) & (g1290) & (keyx106x)));
	assign g1786 = (((!ld) & (!g1001) & (g1297) & (!sk[107]) & (!keyx107x)) + ((!ld) & (!g1001) & (g1297) & (!sk[107]) & (keyx107x)) + ((!ld) & (!g1001) & (g1297) & (sk[107]) & (!keyx107x)) + ((!ld) & (!g1001) & (g1297) & (sk[107]) & (keyx107x)) + ((!ld) & (g1001) & (!g1297) & (!sk[107]) & (!keyx107x)) + ((!ld) & (g1001) & (!g1297) & (!sk[107]) & (keyx107x)) + ((!ld) & (g1001) & (!g1297) & (sk[107]) & (!keyx107x)) + ((!ld) & (g1001) & (!g1297) & (sk[107]) & (keyx107x)) + ((!ld) & (g1001) & (g1297) & (!sk[107]) & (!keyx107x)) + ((!ld) & (g1001) & (g1297) & (!sk[107]) & (keyx107x)) + ((ld) & (!g1001) & (!g1297) & (sk[107]) & (keyx107x)) + ((ld) & (!g1001) & (g1297) & (!sk[107]) & (!keyx107x)) + ((ld) & (!g1001) & (g1297) & (!sk[107]) & (keyx107x)) + ((ld) & (!g1001) & (g1297) & (sk[107]) & (keyx107x)) + ((ld) & (g1001) & (!g1297) & (!sk[107]) & (!keyx107x)) + ((ld) & (g1001) & (!g1297) & (!sk[107]) & (keyx107x)) + ((ld) & (g1001) & (!g1297) & (sk[107]) & (keyx107x)) + ((ld) & (g1001) & (g1297) & (!sk[107]) & (!keyx107x)) + ((ld) & (g1001) & (g1297) & (!sk[107]) & (keyx107x)) + ((ld) & (g1001) & (g1297) & (sk[107]) & (keyx107x)));
	assign g1787 = (((!ld) & (!sk[108]) & (!g1008) & (g1304) & (!keyx108x)) + ((!ld) & (!sk[108]) & (!g1008) & (g1304) & (keyx108x)) + ((!ld) & (!sk[108]) & (g1008) & (!g1304) & (!keyx108x)) + ((!ld) & (!sk[108]) & (g1008) & (!g1304) & (keyx108x)) + ((!ld) & (!sk[108]) & (g1008) & (g1304) & (!keyx108x)) + ((!ld) & (!sk[108]) & (g1008) & (g1304) & (keyx108x)) + ((!ld) & (sk[108]) & (!g1008) & (g1304) & (!keyx108x)) + ((!ld) & (sk[108]) & (!g1008) & (g1304) & (keyx108x)) + ((!ld) & (sk[108]) & (g1008) & (!g1304) & (!keyx108x)) + ((!ld) & (sk[108]) & (g1008) & (!g1304) & (keyx108x)) + ((ld) & (!sk[108]) & (!g1008) & (g1304) & (!keyx108x)) + ((ld) & (!sk[108]) & (!g1008) & (g1304) & (keyx108x)) + ((ld) & (!sk[108]) & (g1008) & (!g1304) & (!keyx108x)) + ((ld) & (!sk[108]) & (g1008) & (!g1304) & (keyx108x)) + ((ld) & (!sk[108]) & (g1008) & (g1304) & (!keyx108x)) + ((ld) & (!sk[108]) & (g1008) & (g1304) & (keyx108x)) + ((ld) & (sk[108]) & (!g1008) & (!g1304) & (keyx108x)) + ((ld) & (sk[108]) & (!g1008) & (g1304) & (keyx108x)) + ((ld) & (sk[108]) & (g1008) & (!g1304) & (keyx108x)) + ((ld) & (sk[108]) & (g1008) & (g1304) & (keyx108x)));
	assign g1788 = (((!ld) & (!g1015) & (!sk[109]) & (g1311) & (!keyx109x)) + ((!ld) & (!g1015) & (!sk[109]) & (g1311) & (keyx109x)) + ((!ld) & (!g1015) & (sk[109]) & (g1311) & (!keyx109x)) + ((!ld) & (!g1015) & (sk[109]) & (g1311) & (keyx109x)) + ((!ld) & (g1015) & (!sk[109]) & (!g1311) & (!keyx109x)) + ((!ld) & (g1015) & (!sk[109]) & (!g1311) & (keyx109x)) + ((!ld) & (g1015) & (!sk[109]) & (g1311) & (!keyx109x)) + ((!ld) & (g1015) & (!sk[109]) & (g1311) & (keyx109x)) + ((!ld) & (g1015) & (sk[109]) & (!g1311) & (!keyx109x)) + ((!ld) & (g1015) & (sk[109]) & (!g1311) & (keyx109x)) + ((ld) & (!g1015) & (!sk[109]) & (g1311) & (!keyx109x)) + ((ld) & (!g1015) & (!sk[109]) & (g1311) & (keyx109x)) + ((ld) & (!g1015) & (sk[109]) & (!g1311) & (keyx109x)) + ((ld) & (!g1015) & (sk[109]) & (g1311) & (keyx109x)) + ((ld) & (g1015) & (!sk[109]) & (!g1311) & (!keyx109x)) + ((ld) & (g1015) & (!sk[109]) & (!g1311) & (keyx109x)) + ((ld) & (g1015) & (!sk[109]) & (g1311) & (!keyx109x)) + ((ld) & (g1015) & (!sk[109]) & (g1311) & (keyx109x)) + ((ld) & (g1015) & (sk[109]) & (!g1311) & (keyx109x)) + ((ld) & (g1015) & (sk[109]) & (g1311) & (keyx109x)));
	assign g1789 = (((!ld) & (!sk[110]) & (!g1022) & (g1318) & (!keyx110x)) + ((!ld) & (!sk[110]) & (!g1022) & (g1318) & (keyx110x)) + ((!ld) & (!sk[110]) & (g1022) & (!g1318) & (!keyx110x)) + ((!ld) & (!sk[110]) & (g1022) & (!g1318) & (keyx110x)) + ((!ld) & (!sk[110]) & (g1022) & (g1318) & (!keyx110x)) + ((!ld) & (!sk[110]) & (g1022) & (g1318) & (keyx110x)) + ((!ld) & (sk[110]) & (!g1022) & (g1318) & (!keyx110x)) + ((!ld) & (sk[110]) & (!g1022) & (g1318) & (keyx110x)) + ((!ld) & (sk[110]) & (g1022) & (!g1318) & (!keyx110x)) + ((!ld) & (sk[110]) & (g1022) & (!g1318) & (keyx110x)) + ((ld) & (!sk[110]) & (!g1022) & (g1318) & (!keyx110x)) + ((ld) & (!sk[110]) & (!g1022) & (g1318) & (keyx110x)) + ((ld) & (!sk[110]) & (g1022) & (!g1318) & (!keyx110x)) + ((ld) & (!sk[110]) & (g1022) & (!g1318) & (keyx110x)) + ((ld) & (!sk[110]) & (g1022) & (g1318) & (!keyx110x)) + ((ld) & (!sk[110]) & (g1022) & (g1318) & (keyx110x)) + ((ld) & (sk[110]) & (!g1022) & (!g1318) & (keyx110x)) + ((ld) & (sk[110]) & (!g1022) & (g1318) & (keyx110x)) + ((ld) & (sk[110]) & (g1022) & (!g1318) & (keyx110x)) + ((ld) & (sk[110]) & (g1022) & (g1318) & (keyx110x)));
	assign g1790 = (((!ld) & (!g1029) & (!sk[111]) & (g1325) & (!keyx111x)) + ((!ld) & (!g1029) & (!sk[111]) & (g1325) & (keyx111x)) + ((!ld) & (!g1029) & (sk[111]) & (g1325) & (!keyx111x)) + ((!ld) & (!g1029) & (sk[111]) & (g1325) & (keyx111x)) + ((!ld) & (g1029) & (!sk[111]) & (!g1325) & (!keyx111x)) + ((!ld) & (g1029) & (!sk[111]) & (!g1325) & (keyx111x)) + ((!ld) & (g1029) & (!sk[111]) & (g1325) & (!keyx111x)) + ((!ld) & (g1029) & (!sk[111]) & (g1325) & (keyx111x)) + ((!ld) & (g1029) & (sk[111]) & (!g1325) & (!keyx111x)) + ((!ld) & (g1029) & (sk[111]) & (!g1325) & (keyx111x)) + ((ld) & (!g1029) & (!sk[111]) & (g1325) & (!keyx111x)) + ((ld) & (!g1029) & (!sk[111]) & (g1325) & (keyx111x)) + ((ld) & (!g1029) & (sk[111]) & (!g1325) & (keyx111x)) + ((ld) & (!g1029) & (sk[111]) & (g1325) & (keyx111x)) + ((ld) & (g1029) & (!sk[111]) & (!g1325) & (!keyx111x)) + ((ld) & (g1029) & (!sk[111]) & (!g1325) & (keyx111x)) + ((ld) & (g1029) & (!sk[111]) & (g1325) & (!keyx111x)) + ((ld) & (g1029) & (!sk[111]) & (g1325) & (keyx111x)) + ((ld) & (g1029) & (sk[111]) & (!g1325) & (keyx111x)) + ((ld) & (g1029) & (sk[111]) & (g1325) & (keyx111x)));
	assign g2194 = (((!sk[112]) & (!ld) & (text_inx80x) & (!g1791)) + ((!sk[112]) & (!ld) & (text_inx80x) & (g1791)) + ((!sk[112]) & (ld) & (!text_inx80x) & (g1791)) + ((!sk[112]) & (ld) & (text_inx80x) & (!g1791)) + ((!sk[112]) & (ld) & (text_inx80x) & (g1791)) + ((sk[112]) & (!ld) & (!text_inx80x) & (g1791)) + ((sk[112]) & (!ld) & (text_inx80x) & (g1791)) + ((sk[112]) & (ld) & (text_inx80x) & (!g1791)) + ((sk[112]) & (ld) & (text_inx80x) & (g1791)));
	assign g1792 = (((!g772) & (!g788) & (!g836) & (sk[113]) & (g851)) + ((!g772) & (!g788) & (g836) & (!sk[113]) & (!g851)) + ((!g772) & (!g788) & (g836) & (!sk[113]) & (g851)) + ((!g772) & (!g788) & (g836) & (sk[113]) & (!g851)) + ((!g772) & (g788) & (!g836) & (!sk[113]) & (!g851)) + ((!g772) & (g788) & (!g836) & (!sk[113]) & (g851)) + ((!g772) & (g788) & (!g836) & (sk[113]) & (!g851)) + ((!g772) & (g788) & (g836) & (!sk[113]) & (!g851)) + ((!g772) & (g788) & (g836) & (!sk[113]) & (g851)) + ((!g772) & (g788) & (g836) & (sk[113]) & (g851)) + ((g772) & (!g788) & (!g836) & (sk[113]) & (!g851)) + ((g772) & (!g788) & (g836) & (!sk[113]) & (!g851)) + ((g772) & (!g788) & (g836) & (!sk[113]) & (g851)) + ((g772) & (!g788) & (g836) & (sk[113]) & (g851)) + ((g772) & (g788) & (!g836) & (!sk[113]) & (!g851)) + ((g772) & (g788) & (!g836) & (!sk[113]) & (g851)) + ((g772) & (g788) & (!g836) & (sk[113]) & (g851)) + ((g772) & (g788) & (g836) & (!sk[113]) & (!g851)) + ((g772) & (g788) & (g836) & (!sk[113]) & (g851)) + ((g772) & (g788) & (g836) & (sk[113]) & (!g851)));
	assign g1793 = (((!g659) & (!g723) & (!g788) & (!g1163) & (!g1791) & (g1792)) + ((!g659) & (!g723) & (!g788) & (!g1163) & (g1791) & (g1792)) + ((!g659) & (!g723) & (!g788) & (g1163) & (g1791) & (!g1792)) + ((!g659) & (!g723) & (!g788) & (g1163) & (g1791) & (g1792)) + ((!g659) & (!g723) & (g788) & (!g1163) & (!g1791) & (g1792)) + ((!g659) & (!g723) & (g788) & (!g1163) & (g1791) & (g1792)) + ((!g659) & (!g723) & (g788) & (g1163) & (!g1791) & (!g1792)) + ((!g659) & (!g723) & (g788) & (g1163) & (!g1791) & (g1792)) + ((!g659) & (g723) & (!g788) & (!g1163) & (!g1791) & (!g1792)) + ((!g659) & (g723) & (!g788) & (!g1163) & (g1791) & (!g1792)) + ((!g659) & (g723) & (!g788) & (g1163) & (g1791) & (!g1792)) + ((!g659) & (g723) & (!g788) & (g1163) & (g1791) & (g1792)) + ((!g659) & (g723) & (g788) & (!g1163) & (!g1791) & (!g1792)) + ((!g659) & (g723) & (g788) & (!g1163) & (g1791) & (!g1792)) + ((!g659) & (g723) & (g788) & (g1163) & (!g1791) & (!g1792)) + ((!g659) & (g723) & (g788) & (g1163) & (!g1791) & (g1792)) + ((g659) & (!g723) & (!g788) & (!g1163) & (!g1791) & (!g1792)) + ((g659) & (!g723) & (!g788) & (!g1163) & (g1791) & (!g1792)) + ((g659) & (!g723) & (!g788) & (g1163) & (g1791) & (!g1792)) + ((g659) & (!g723) & (!g788) & (g1163) & (g1791) & (g1792)) + ((g659) & (!g723) & (g788) & (!g1163) & (!g1791) & (!g1792)) + ((g659) & (!g723) & (g788) & (!g1163) & (g1791) & (!g1792)) + ((g659) & (!g723) & (g788) & (g1163) & (!g1791) & (!g1792)) + ((g659) & (!g723) & (g788) & (g1163) & (!g1791) & (g1792)) + ((g659) & (g723) & (!g788) & (!g1163) & (!g1791) & (g1792)) + ((g659) & (g723) & (!g788) & (!g1163) & (g1791) & (g1792)) + ((g659) & (g723) & (!g788) & (g1163) & (g1791) & (!g1792)) + ((g659) & (g723) & (!g788) & (g1163) & (g1791) & (g1792)) + ((g659) & (g723) & (g788) & (!g1163) & (!g1791) & (g1792)) + ((g659) & (g723) & (g788) & (!g1163) & (g1791) & (g1792)) + ((g659) & (g723) & (g788) & (g1163) & (!g1791) & (!g1792)) + ((g659) & (g723) & (g788) & (g1163) & (!g1791) & (g1792)));
	assign g2195 = (((!ld) & (!text_inx81x) & (sk[115]) & (g1794)) + ((!ld) & (text_inx81x) & (!sk[115]) & (!g1794)) + ((!ld) & (text_inx81x) & (!sk[115]) & (g1794)) + ((!ld) & (text_inx81x) & (sk[115]) & (g1794)) + ((ld) & (!text_inx81x) & (!sk[115]) & (g1794)) + ((ld) & (text_inx81x) & (!sk[115]) & (!g1794)) + ((ld) & (text_inx81x) & (!sk[115]) & (g1794)) + ((ld) & (text_inx81x) & (sk[115]) & (!g1794)) + ((ld) & (text_inx81x) & (sk[115]) & (g1794)));
	assign g1795 = (((!g723) & (!g730) & (!g772) & (!g787) & (!g795) & (g836)) + ((!g723) & (!g730) & (!g772) & (!g787) & (g795) & (!g836)) + ((!g723) & (!g730) & (!g772) & (g787) & (!g795) & (!g836)) + ((!g723) & (!g730) & (!g772) & (g787) & (g795) & (g836)) + ((!g723) & (!g730) & (g772) & (!g787) & (!g795) & (!g836)) + ((!g723) & (!g730) & (g772) & (!g787) & (g795) & (g836)) + ((!g723) & (!g730) & (g772) & (g787) & (!g795) & (g836)) + ((!g723) & (!g730) & (g772) & (g787) & (g795) & (!g836)) + ((!g723) & (g730) & (!g772) & (!g787) & (!g795) & (!g836)) + ((!g723) & (g730) & (!g772) & (!g787) & (g795) & (g836)) + ((!g723) & (g730) & (!g772) & (g787) & (!g795) & (g836)) + ((!g723) & (g730) & (!g772) & (g787) & (g795) & (!g836)) + ((!g723) & (g730) & (g772) & (!g787) & (!g795) & (g836)) + ((!g723) & (g730) & (g772) & (!g787) & (g795) & (!g836)) + ((!g723) & (g730) & (g772) & (g787) & (!g795) & (!g836)) + ((!g723) & (g730) & (g772) & (g787) & (g795) & (g836)) + ((g723) & (!g730) & (!g772) & (!g787) & (!g795) & (!g836)) + ((g723) & (!g730) & (!g772) & (!g787) & (g795) & (g836)) + ((g723) & (!g730) & (!g772) & (g787) & (!g795) & (g836)) + ((g723) & (!g730) & (!g772) & (g787) & (g795) & (!g836)) + ((g723) & (!g730) & (g772) & (!g787) & (!g795) & (g836)) + ((g723) & (!g730) & (g772) & (!g787) & (g795) & (!g836)) + ((g723) & (!g730) & (g772) & (g787) & (!g795) & (!g836)) + ((g723) & (!g730) & (g772) & (g787) & (g795) & (g836)) + ((g723) & (g730) & (!g772) & (!g787) & (!g795) & (g836)) + ((g723) & (g730) & (!g772) & (!g787) & (g795) & (!g836)) + ((g723) & (g730) & (!g772) & (g787) & (!g795) & (!g836)) + ((g723) & (g730) & (!g772) & (g787) & (g795) & (g836)) + ((g723) & (g730) & (g772) & (!g787) & (!g795) & (!g836)) + ((g723) & (g730) & (g772) & (!g787) & (g795) & (g836)) + ((g723) & (g730) & (g772) & (g787) & (!g795) & (g836)) + ((g723) & (g730) & (g772) & (g787) & (g795) & (!g836)));
	assign g1796 = (((!g795) & (!g1163) & (!g1250) & (!g1794) & (sk[117]) & (g1795)) + ((!g795) & (!g1163) & (!g1250) & (g1794) & (sk[117]) & (g1795)) + ((!g795) & (!g1163) & (g1250) & (!g1794) & (sk[117]) & (!g1795)) + ((!g795) & (!g1163) & (g1250) & (g1794) & (sk[117]) & (!g1795)) + ((!g795) & (g1163) & (!g1250) & (!g1794) & (!sk[117]) & (!g1795)) + ((!g795) & (g1163) & (!g1250) & (!g1794) & (!sk[117]) & (g1795)) + ((!g795) & (g1163) & (!g1250) & (g1794) & (!sk[117]) & (!g1795)) + ((!g795) & (g1163) & (!g1250) & (g1794) & (!sk[117]) & (g1795)) + ((!g795) & (g1163) & (!g1250) & (g1794) & (sk[117]) & (!g1795)) + ((!g795) & (g1163) & (!g1250) & (g1794) & (sk[117]) & (g1795)) + ((!g795) & (g1163) & (g1250) & (!g1794) & (!sk[117]) & (!g1795)) + ((!g795) & (g1163) & (g1250) & (!g1794) & (!sk[117]) & (g1795)) + ((!g795) & (g1163) & (g1250) & (g1794) & (!sk[117]) & (!g1795)) + ((!g795) & (g1163) & (g1250) & (g1794) & (!sk[117]) & (g1795)) + ((!g795) & (g1163) & (g1250) & (g1794) & (sk[117]) & (!g1795)) + ((!g795) & (g1163) & (g1250) & (g1794) & (sk[117]) & (g1795)) + ((g795) & (!g1163) & (!g1250) & (!g1794) & (!sk[117]) & (!g1795)) + ((g795) & (!g1163) & (!g1250) & (!g1794) & (!sk[117]) & (g1795)) + ((g795) & (!g1163) & (!g1250) & (!g1794) & (sk[117]) & (g1795)) + ((g795) & (!g1163) & (!g1250) & (g1794) & (!sk[117]) & (!g1795)) + ((g795) & (!g1163) & (!g1250) & (g1794) & (!sk[117]) & (g1795)) + ((g795) & (!g1163) & (!g1250) & (g1794) & (sk[117]) & (g1795)) + ((g795) & (!g1163) & (g1250) & (!g1794) & (!sk[117]) & (!g1795)) + ((g795) & (!g1163) & (g1250) & (!g1794) & (!sk[117]) & (g1795)) + ((g795) & (!g1163) & (g1250) & (!g1794) & (sk[117]) & (!g1795)) + ((g795) & (!g1163) & (g1250) & (g1794) & (!sk[117]) & (!g1795)) + ((g795) & (!g1163) & (g1250) & (g1794) & (!sk[117]) & (g1795)) + ((g795) & (!g1163) & (g1250) & (g1794) & (sk[117]) & (!g1795)) + ((g795) & (g1163) & (!g1250) & (!g1794) & (!sk[117]) & (!g1795)) + ((g795) & (g1163) & (!g1250) & (!g1794) & (!sk[117]) & (g1795)) + ((g795) & (g1163) & (!g1250) & (!g1794) & (sk[117]) & (!g1795)) + ((g795) & (g1163) & (!g1250) & (!g1794) & (sk[117]) & (g1795)) + ((g795) & (g1163) & (!g1250) & (g1794) & (!sk[117]) & (!g1795)) + ((g795) & (g1163) & (!g1250) & (g1794) & (!sk[117]) & (g1795)) + ((g795) & (g1163) & (g1250) & (!g1794) & (!sk[117]) & (!g1795)) + ((g795) & (g1163) & (g1250) & (!g1794) & (!sk[117]) & (g1795)) + ((g795) & (g1163) & (g1250) & (!g1794) & (sk[117]) & (!g1795)) + ((g795) & (g1163) & (g1250) & (!g1794) & (sk[117]) & (g1795)) + ((g795) & (g1163) & (g1250) & (g1794) & (!sk[117]) & (!g1795)) + ((g795) & (g1163) & (g1250) & (g1794) & (!sk[117]) & (g1795)));
	assign g2196 = (((!ld) & (!sk[118]) & (text_inx82x) & (!g1797)) + ((!ld) & (!sk[118]) & (text_inx82x) & (g1797)) + ((!ld) & (sk[118]) & (!text_inx82x) & (g1797)) + ((!ld) & (sk[118]) & (text_inx82x) & (g1797)) + ((ld) & (!sk[118]) & (!text_inx82x) & (g1797)) + ((ld) & (!sk[118]) & (text_inx82x) & (!g1797)) + ((ld) & (!sk[118]) & (text_inx82x) & (g1797)) + ((ld) & (sk[118]) & (text_inx82x) & (!g1797)) + ((ld) & (sk[118]) & (text_inx82x) & (g1797)));
	assign g1798 = (((!g730) & (!g802) & (!g865) & (!g1163) & (g1713) & (!g1797)) + ((!g730) & (!g802) & (!g865) & (!g1163) & (g1713) & (g1797)) + ((!g730) & (!g802) & (!g865) & (g1163) & (!g1713) & (g1797)) + ((!g730) & (!g802) & (!g865) & (g1163) & (g1713) & (g1797)) + ((!g730) & (!g802) & (g865) & (!g1163) & (!g1713) & (!g1797)) + ((!g730) & (!g802) & (g865) & (!g1163) & (!g1713) & (g1797)) + ((!g730) & (!g802) & (g865) & (g1163) & (!g1713) & (g1797)) + ((!g730) & (!g802) & (g865) & (g1163) & (g1713) & (g1797)) + ((!g730) & (g802) & (!g865) & (!g1163) & (!g1713) & (!g1797)) + ((!g730) & (g802) & (!g865) & (!g1163) & (!g1713) & (g1797)) + ((!g730) & (g802) & (!g865) & (g1163) & (!g1713) & (!g1797)) + ((!g730) & (g802) & (!g865) & (g1163) & (g1713) & (!g1797)) + ((!g730) & (g802) & (g865) & (!g1163) & (g1713) & (!g1797)) + ((!g730) & (g802) & (g865) & (!g1163) & (g1713) & (g1797)) + ((!g730) & (g802) & (g865) & (g1163) & (!g1713) & (!g1797)) + ((!g730) & (g802) & (g865) & (g1163) & (g1713) & (!g1797)) + ((g730) & (!g802) & (!g865) & (!g1163) & (!g1713) & (!g1797)) + ((g730) & (!g802) & (!g865) & (!g1163) & (!g1713) & (g1797)) + ((g730) & (!g802) & (!g865) & (g1163) & (!g1713) & (g1797)) + ((g730) & (!g802) & (!g865) & (g1163) & (g1713) & (g1797)) + ((g730) & (!g802) & (g865) & (!g1163) & (g1713) & (!g1797)) + ((g730) & (!g802) & (g865) & (!g1163) & (g1713) & (g1797)) + ((g730) & (!g802) & (g865) & (g1163) & (!g1713) & (g1797)) + ((g730) & (!g802) & (g865) & (g1163) & (g1713) & (g1797)) + ((g730) & (g802) & (!g865) & (!g1163) & (g1713) & (!g1797)) + ((g730) & (g802) & (!g865) & (!g1163) & (g1713) & (g1797)) + ((g730) & (g802) & (!g865) & (g1163) & (!g1713) & (!g1797)) + ((g730) & (g802) & (!g865) & (g1163) & (g1713) & (!g1797)) + ((g730) & (g802) & (g865) & (!g1163) & (!g1713) & (!g1797)) + ((g730) & (g802) & (g865) & (!g1163) & (!g1713) & (g1797)) + ((g730) & (g802) & (g865) & (g1163) & (!g1713) & (!g1797)) + ((g730) & (g802) & (g865) & (g1163) & (g1713) & (!g1797)));
	assign g2197 = (((!sk[120]) & (!ld) & (text_inx83x) & (!g1799)) + ((!sk[120]) & (!ld) & (text_inx83x) & (g1799)) + ((!sk[120]) & (ld) & (!text_inx83x) & (g1799)) + ((!sk[120]) & (ld) & (text_inx83x) & (!g1799)) + ((!sk[120]) & (ld) & (text_inx83x) & (g1799)) + ((sk[120]) & (!ld) & (!text_inx83x) & (g1799)) + ((sk[120]) & (!ld) & (text_inx83x) & (g1799)) + ((sk[120]) & (ld) & (text_inx83x) & (!g1799)) + ((sk[120]) & (ld) & (text_inx83x) & (g1799)));
	assign g1800 = (((!g680) & (!sk[121]) & (g737) & (!g744) & (!g772) & (!g809)) + ((!g680) & (!sk[121]) & (g737) & (!g744) & (!g772) & (g809)) + ((!g680) & (!sk[121]) & (g737) & (!g744) & (g772) & (!g809)) + ((!g680) & (!sk[121]) & (g737) & (!g744) & (g772) & (g809)) + ((!g680) & (!sk[121]) & (g737) & (g744) & (!g772) & (!g809)) + ((!g680) & (!sk[121]) & (g737) & (g744) & (!g772) & (g809)) + ((!g680) & (!sk[121]) & (g737) & (g744) & (g772) & (!g809)) + ((!g680) & (!sk[121]) & (g737) & (g744) & (g772) & (g809)) + ((!g680) & (sk[121]) & (!g737) & (!g744) & (!g772) & (g809)) + ((!g680) & (sk[121]) & (!g737) & (!g744) & (g772) & (!g809)) + ((!g680) & (sk[121]) & (!g737) & (g744) & (!g772) & (!g809)) + ((!g680) & (sk[121]) & (!g737) & (g744) & (g772) & (g809)) + ((!g680) & (sk[121]) & (g737) & (!g744) & (!g772) & (!g809)) + ((!g680) & (sk[121]) & (g737) & (!g744) & (g772) & (g809)) + ((!g680) & (sk[121]) & (g737) & (g744) & (!g772) & (g809)) + ((!g680) & (sk[121]) & (g737) & (g744) & (g772) & (!g809)) + ((g680) & (!sk[121]) & (!g737) & (!g744) & (!g772) & (!g809)) + ((g680) & (!sk[121]) & (!g737) & (!g744) & (!g772) & (g809)) + ((g680) & (!sk[121]) & (!g737) & (!g744) & (g772) & (!g809)) + ((g680) & (!sk[121]) & (!g737) & (!g744) & (g772) & (g809)) + ((g680) & (!sk[121]) & (!g737) & (g744) & (!g772) & (!g809)) + ((g680) & (!sk[121]) & (!g737) & (g744) & (!g772) & (g809)) + ((g680) & (!sk[121]) & (!g737) & (g744) & (g772) & (!g809)) + ((g680) & (!sk[121]) & (!g737) & (g744) & (g772) & (g809)) + ((g680) & (!sk[121]) & (g737) & (!g744) & (!g772) & (!g809)) + ((g680) & (!sk[121]) & (g737) & (!g744) & (!g772) & (g809)) + ((g680) & (!sk[121]) & (g737) & (!g744) & (g772) & (!g809)) + ((g680) & (!sk[121]) & (g737) & (!g744) & (g772) & (g809)) + ((g680) & (!sk[121]) & (g737) & (g744) & (!g772) & (!g809)) + ((g680) & (!sk[121]) & (g737) & (g744) & (!g772) & (g809)) + ((g680) & (!sk[121]) & (g737) & (g744) & (g772) & (!g809)) + ((g680) & (!sk[121]) & (g737) & (g744) & (g772) & (g809)) + ((g680) & (sk[121]) & (!g737) & (!g744) & (!g772) & (!g809)) + ((g680) & (sk[121]) & (!g737) & (!g744) & (g772) & (g809)) + ((g680) & (sk[121]) & (!g737) & (g744) & (!g772) & (g809)) + ((g680) & (sk[121]) & (!g737) & (g744) & (g772) & (!g809)) + ((g680) & (sk[121]) & (g737) & (!g744) & (!g772) & (g809)) + ((g680) & (sk[121]) & (g737) & (!g744) & (g772) & (!g809)) + ((g680) & (sk[121]) & (g737) & (g744) & (!g772) & (!g809)) + ((g680) & (sk[121]) & (g737) & (g744) & (g772) & (g809)));
	assign g1801 = (((!g809) & (!g872) & (!g1163) & (!g1716) & (!g1799) & (g1800)) + ((!g809) & (!g872) & (!g1163) & (!g1716) & (g1799) & (g1800)) + ((!g809) & (!g872) & (!g1163) & (g1716) & (!g1799) & (!g1800)) + ((!g809) & (!g872) & (!g1163) & (g1716) & (g1799) & (!g1800)) + ((!g809) & (!g872) & (g1163) & (!g1716) & (g1799) & (!g1800)) + ((!g809) & (!g872) & (g1163) & (!g1716) & (g1799) & (g1800)) + ((!g809) & (!g872) & (g1163) & (g1716) & (g1799) & (!g1800)) + ((!g809) & (!g872) & (g1163) & (g1716) & (g1799) & (g1800)) + ((!g809) & (g872) & (!g1163) & (!g1716) & (!g1799) & (!g1800)) + ((!g809) & (g872) & (!g1163) & (!g1716) & (g1799) & (!g1800)) + ((!g809) & (g872) & (!g1163) & (g1716) & (!g1799) & (g1800)) + ((!g809) & (g872) & (!g1163) & (g1716) & (g1799) & (g1800)) + ((!g809) & (g872) & (g1163) & (!g1716) & (g1799) & (!g1800)) + ((!g809) & (g872) & (g1163) & (!g1716) & (g1799) & (g1800)) + ((!g809) & (g872) & (g1163) & (g1716) & (g1799) & (!g1800)) + ((!g809) & (g872) & (g1163) & (g1716) & (g1799) & (g1800)) + ((g809) & (!g872) & (!g1163) & (!g1716) & (!g1799) & (g1800)) + ((g809) & (!g872) & (!g1163) & (!g1716) & (g1799) & (g1800)) + ((g809) & (!g872) & (!g1163) & (g1716) & (!g1799) & (!g1800)) + ((g809) & (!g872) & (!g1163) & (g1716) & (g1799) & (!g1800)) + ((g809) & (!g872) & (g1163) & (!g1716) & (!g1799) & (!g1800)) + ((g809) & (!g872) & (g1163) & (!g1716) & (!g1799) & (g1800)) + ((g809) & (!g872) & (g1163) & (g1716) & (!g1799) & (!g1800)) + ((g809) & (!g872) & (g1163) & (g1716) & (!g1799) & (g1800)) + ((g809) & (g872) & (!g1163) & (!g1716) & (!g1799) & (!g1800)) + ((g809) & (g872) & (!g1163) & (!g1716) & (g1799) & (!g1800)) + ((g809) & (g872) & (!g1163) & (g1716) & (!g1799) & (g1800)) + ((g809) & (g872) & (!g1163) & (g1716) & (g1799) & (g1800)) + ((g809) & (g872) & (g1163) & (!g1716) & (!g1799) & (!g1800)) + ((g809) & (g872) & (g1163) & (!g1716) & (!g1799) & (g1800)) + ((g809) & (g872) & (g1163) & (g1716) & (!g1799) & (!g1800)) + ((g809) & (g872) & (g1163) & (g1716) & (!g1799) & (g1800)));
	assign g2198 = (((!ld) & (!text_inx86x) & (sk[123]) & (g1802)) + ((!ld) & (text_inx86x) & (!sk[123]) & (!g1802)) + ((!ld) & (text_inx86x) & (!sk[123]) & (g1802)) + ((!ld) & (text_inx86x) & (sk[123]) & (g1802)) + ((ld) & (!text_inx86x) & (!sk[123]) & (g1802)) + ((ld) & (text_inx86x) & (!sk[123]) & (!g1802)) + ((ld) & (text_inx86x) & (!sk[123]) & (g1802)) + ((ld) & (text_inx86x) & (sk[123]) & (!g1802)) + ((ld) & (text_inx86x) & (sk[123]) & (g1802)));
	assign g1803 = (((!g758) & (!g830) & (!g893) & (!g1163) & (g1719) & (!g1802)) + ((!g758) & (!g830) & (!g893) & (!g1163) & (g1719) & (g1802)) + ((!g758) & (!g830) & (!g893) & (g1163) & (!g1719) & (g1802)) + ((!g758) & (!g830) & (!g893) & (g1163) & (g1719) & (g1802)) + ((!g758) & (!g830) & (g893) & (!g1163) & (!g1719) & (!g1802)) + ((!g758) & (!g830) & (g893) & (!g1163) & (!g1719) & (g1802)) + ((!g758) & (!g830) & (g893) & (g1163) & (!g1719) & (g1802)) + ((!g758) & (!g830) & (g893) & (g1163) & (g1719) & (g1802)) + ((!g758) & (g830) & (!g893) & (!g1163) & (!g1719) & (!g1802)) + ((!g758) & (g830) & (!g893) & (!g1163) & (!g1719) & (g1802)) + ((!g758) & (g830) & (!g893) & (g1163) & (!g1719) & (!g1802)) + ((!g758) & (g830) & (!g893) & (g1163) & (g1719) & (!g1802)) + ((!g758) & (g830) & (g893) & (!g1163) & (g1719) & (!g1802)) + ((!g758) & (g830) & (g893) & (!g1163) & (g1719) & (g1802)) + ((!g758) & (g830) & (g893) & (g1163) & (!g1719) & (!g1802)) + ((!g758) & (g830) & (g893) & (g1163) & (g1719) & (!g1802)) + ((g758) & (!g830) & (!g893) & (!g1163) & (!g1719) & (!g1802)) + ((g758) & (!g830) & (!g893) & (!g1163) & (!g1719) & (g1802)) + ((g758) & (!g830) & (!g893) & (g1163) & (!g1719) & (g1802)) + ((g758) & (!g830) & (!g893) & (g1163) & (g1719) & (g1802)) + ((g758) & (!g830) & (g893) & (!g1163) & (g1719) & (!g1802)) + ((g758) & (!g830) & (g893) & (!g1163) & (g1719) & (g1802)) + ((g758) & (!g830) & (g893) & (g1163) & (!g1719) & (g1802)) + ((g758) & (!g830) & (g893) & (g1163) & (g1719) & (g1802)) + ((g758) & (g830) & (!g893) & (!g1163) & (g1719) & (!g1802)) + ((g758) & (g830) & (!g893) & (!g1163) & (g1719) & (g1802)) + ((g758) & (g830) & (!g893) & (g1163) & (!g1719) & (!g1802)) + ((g758) & (g830) & (!g893) & (g1163) & (g1719) & (!g1802)) + ((g758) & (g830) & (g893) & (!g1163) & (!g1719) & (!g1802)) + ((g758) & (g830) & (g893) & (!g1163) & (!g1719) & (g1802)) + ((g758) & (g830) & (g893) & (g1163) & (!g1719) & (!g1802)) + ((g758) & (g830) & (g893) & (g1163) & (g1719) & (!g1802)));
	assign g2199 = (((!ld) & (!sk[125]) & (text_inx85x) & (!g1804)) + ((!ld) & (!sk[125]) & (text_inx85x) & (g1804)) + ((!ld) & (sk[125]) & (!text_inx85x) & (g1804)) + ((!ld) & (sk[125]) & (text_inx85x) & (g1804)) + ((ld) & (!sk[125]) & (!text_inx85x) & (g1804)) + ((ld) & (!sk[125]) & (text_inx85x) & (!g1804)) + ((ld) & (!sk[125]) & (text_inx85x) & (g1804)) + ((ld) & (sk[125]) & (text_inx85x) & (!g1804)) + ((ld) & (sk[125]) & (text_inx85x) & (g1804)));
	assign g1805 = (((!g751) & (!g823) & (!g886) & (!g1163) & (g1722) & (!g1804)) + ((!g751) & (!g823) & (!g886) & (!g1163) & (g1722) & (g1804)) + ((!g751) & (!g823) & (!g886) & (g1163) & (!g1722) & (g1804)) + ((!g751) & (!g823) & (!g886) & (g1163) & (g1722) & (g1804)) + ((!g751) & (!g823) & (g886) & (!g1163) & (!g1722) & (!g1804)) + ((!g751) & (!g823) & (g886) & (!g1163) & (!g1722) & (g1804)) + ((!g751) & (!g823) & (g886) & (g1163) & (!g1722) & (g1804)) + ((!g751) & (!g823) & (g886) & (g1163) & (g1722) & (g1804)) + ((!g751) & (g823) & (!g886) & (!g1163) & (!g1722) & (!g1804)) + ((!g751) & (g823) & (!g886) & (!g1163) & (!g1722) & (g1804)) + ((!g751) & (g823) & (!g886) & (g1163) & (!g1722) & (!g1804)) + ((!g751) & (g823) & (!g886) & (g1163) & (g1722) & (!g1804)) + ((!g751) & (g823) & (g886) & (!g1163) & (g1722) & (!g1804)) + ((!g751) & (g823) & (g886) & (!g1163) & (g1722) & (g1804)) + ((!g751) & (g823) & (g886) & (g1163) & (!g1722) & (!g1804)) + ((!g751) & (g823) & (g886) & (g1163) & (g1722) & (!g1804)) + ((g751) & (!g823) & (!g886) & (!g1163) & (!g1722) & (!g1804)) + ((g751) & (!g823) & (!g886) & (!g1163) & (!g1722) & (g1804)) + ((g751) & (!g823) & (!g886) & (g1163) & (!g1722) & (g1804)) + ((g751) & (!g823) & (!g886) & (g1163) & (g1722) & (g1804)) + ((g751) & (!g823) & (g886) & (!g1163) & (g1722) & (!g1804)) + ((g751) & (!g823) & (g886) & (!g1163) & (g1722) & (g1804)) + ((g751) & (!g823) & (g886) & (g1163) & (!g1722) & (g1804)) + ((g751) & (!g823) & (g886) & (g1163) & (g1722) & (g1804)) + ((g751) & (g823) & (!g886) & (!g1163) & (g1722) & (!g1804)) + ((g751) & (g823) & (!g886) & (!g1163) & (g1722) & (g1804)) + ((g751) & (g823) & (!g886) & (g1163) & (!g1722) & (!g1804)) + ((g751) & (g823) & (!g886) & (g1163) & (g1722) & (!g1804)) + ((g751) & (g823) & (g886) & (!g1163) & (!g1722) & (!g1804)) + ((g751) & (g823) & (g886) & (!g1163) & (!g1722) & (g1804)) + ((g751) & (g823) & (g886) & (g1163) & (!g1722) & (!g1804)) + ((g751) & (g823) & (g886) & (g1163) & (g1722) & (!g1804)));
	assign g2200 = (((!sk[127]) & (!ld) & (text_inx84x) & (!g1806)) + ((!sk[127]) & (!ld) & (text_inx84x) & (g1806)) + ((!sk[127]) & (ld) & (!text_inx84x) & (g1806)) + ((!sk[127]) & (ld) & (text_inx84x) & (!g1806)) + ((!sk[127]) & (ld) & (text_inx84x) & (g1806)) + ((sk[127]) & (!ld) & (!text_inx84x) & (g1806)) + ((sk[127]) & (!ld) & (text_inx84x) & (g1806)) + ((sk[127]) & (ld) & (text_inx84x) & (!g1806)) + ((sk[127]) & (ld) & (text_inx84x) & (g1806)));
	assign g1807 = (((!g744) & (!g772) & (!g816) & (sk[0]) & (!g836) & (g879)) + ((!g744) & (!g772) & (!g816) & (sk[0]) & (g836) & (!g879)) + ((!g744) & (!g772) & (g816) & (sk[0]) & (!g836) & (!g879)) + ((!g744) & (!g772) & (g816) & (sk[0]) & (g836) & (g879)) + ((!g744) & (g772) & (!g816) & (!sk[0]) & (!g836) & (!g879)) + ((!g744) & (g772) & (!g816) & (!sk[0]) & (!g836) & (g879)) + ((!g744) & (g772) & (!g816) & (!sk[0]) & (g836) & (!g879)) + ((!g744) & (g772) & (!g816) & (!sk[0]) & (g836) & (g879)) + ((!g744) & (g772) & (!g816) & (sk[0]) & (!g836) & (!g879)) + ((!g744) & (g772) & (!g816) & (sk[0]) & (g836) & (g879)) + ((!g744) & (g772) & (g816) & (!sk[0]) & (!g836) & (!g879)) + ((!g744) & (g772) & (g816) & (!sk[0]) & (!g836) & (g879)) + ((!g744) & (g772) & (g816) & (!sk[0]) & (g836) & (!g879)) + ((!g744) & (g772) & (g816) & (!sk[0]) & (g836) & (g879)) + ((!g744) & (g772) & (g816) & (sk[0]) & (!g836) & (g879)) + ((!g744) & (g772) & (g816) & (sk[0]) & (g836) & (!g879)) + ((g744) & (!g772) & (!g816) & (!sk[0]) & (!g836) & (!g879)) + ((g744) & (!g772) & (!g816) & (!sk[0]) & (!g836) & (g879)) + ((g744) & (!g772) & (!g816) & (!sk[0]) & (g836) & (!g879)) + ((g744) & (!g772) & (!g816) & (!sk[0]) & (g836) & (g879)) + ((g744) & (!g772) & (!g816) & (sk[0]) & (!g836) & (!g879)) + ((g744) & (!g772) & (!g816) & (sk[0]) & (g836) & (g879)) + ((g744) & (!g772) & (g816) & (!sk[0]) & (!g836) & (!g879)) + ((g744) & (!g772) & (g816) & (!sk[0]) & (!g836) & (g879)) + ((g744) & (!g772) & (g816) & (!sk[0]) & (g836) & (!g879)) + ((g744) & (!g772) & (g816) & (!sk[0]) & (g836) & (g879)) + ((g744) & (!g772) & (g816) & (sk[0]) & (!g836) & (g879)) + ((g744) & (!g772) & (g816) & (sk[0]) & (g836) & (!g879)) + ((g744) & (g772) & (!g816) & (!sk[0]) & (!g836) & (!g879)) + ((g744) & (g772) & (!g816) & (!sk[0]) & (!g836) & (g879)) + ((g744) & (g772) & (!g816) & (!sk[0]) & (g836) & (!g879)) + ((g744) & (g772) & (!g816) & (!sk[0]) & (g836) & (g879)) + ((g744) & (g772) & (!g816) & (sk[0]) & (!g836) & (g879)) + ((g744) & (g772) & (!g816) & (sk[0]) & (g836) & (!g879)) + ((g744) & (g772) & (g816) & (!sk[0]) & (!g836) & (!g879)) + ((g744) & (g772) & (g816) & (!sk[0]) & (!g836) & (g879)) + ((g744) & (g772) & (g816) & (!sk[0]) & (g836) & (!g879)) + ((g744) & (g772) & (g816) & (!sk[0]) & (g836) & (g879)) + ((g744) & (g772) & (g816) & (sk[0]) & (!g836) & (!g879)) + ((g744) & (g772) & (g816) & (sk[0]) & (g836) & (g879)));
	assign g1808 = (((!sk[1]) & (!g816) & (g1163) & (!g1725) & (!g1806) & (!g1807)) + ((!sk[1]) & (!g816) & (g1163) & (!g1725) & (!g1806) & (g1807)) + ((!sk[1]) & (!g816) & (g1163) & (!g1725) & (g1806) & (!g1807)) + ((!sk[1]) & (!g816) & (g1163) & (!g1725) & (g1806) & (g1807)) + ((!sk[1]) & (!g816) & (g1163) & (g1725) & (!g1806) & (!g1807)) + ((!sk[1]) & (!g816) & (g1163) & (g1725) & (!g1806) & (g1807)) + ((!sk[1]) & (!g816) & (g1163) & (g1725) & (g1806) & (!g1807)) + ((!sk[1]) & (!g816) & (g1163) & (g1725) & (g1806) & (g1807)) + ((!sk[1]) & (g816) & (!g1163) & (!g1725) & (!g1806) & (!g1807)) + ((!sk[1]) & (g816) & (!g1163) & (!g1725) & (!g1806) & (g1807)) + ((!sk[1]) & (g816) & (!g1163) & (!g1725) & (g1806) & (!g1807)) + ((!sk[1]) & (g816) & (!g1163) & (!g1725) & (g1806) & (g1807)) + ((!sk[1]) & (g816) & (!g1163) & (g1725) & (!g1806) & (!g1807)) + ((!sk[1]) & (g816) & (!g1163) & (g1725) & (!g1806) & (g1807)) + ((!sk[1]) & (g816) & (!g1163) & (g1725) & (g1806) & (!g1807)) + ((!sk[1]) & (g816) & (!g1163) & (g1725) & (g1806) & (g1807)) + ((!sk[1]) & (g816) & (g1163) & (!g1725) & (!g1806) & (!g1807)) + ((!sk[1]) & (g816) & (g1163) & (!g1725) & (!g1806) & (g1807)) + ((!sk[1]) & (g816) & (g1163) & (!g1725) & (g1806) & (!g1807)) + ((!sk[1]) & (g816) & (g1163) & (!g1725) & (g1806) & (g1807)) + ((!sk[1]) & (g816) & (g1163) & (g1725) & (!g1806) & (!g1807)) + ((!sk[1]) & (g816) & (g1163) & (g1725) & (!g1806) & (g1807)) + ((!sk[1]) & (g816) & (g1163) & (g1725) & (g1806) & (!g1807)) + ((!sk[1]) & (g816) & (g1163) & (g1725) & (g1806) & (g1807)) + ((sk[1]) & (!g816) & (!g1163) & (!g1725) & (!g1806) & (g1807)) + ((sk[1]) & (!g816) & (!g1163) & (!g1725) & (g1806) & (g1807)) + ((sk[1]) & (!g816) & (!g1163) & (g1725) & (!g1806) & (!g1807)) + ((sk[1]) & (!g816) & (!g1163) & (g1725) & (g1806) & (!g1807)) + ((sk[1]) & (!g816) & (g1163) & (!g1725) & (g1806) & (!g1807)) + ((sk[1]) & (!g816) & (g1163) & (!g1725) & (g1806) & (g1807)) + ((sk[1]) & (!g816) & (g1163) & (g1725) & (g1806) & (!g1807)) + ((sk[1]) & (!g816) & (g1163) & (g1725) & (g1806) & (g1807)) + ((sk[1]) & (g816) & (!g1163) & (!g1725) & (!g1806) & (g1807)) + ((sk[1]) & (g816) & (!g1163) & (!g1725) & (g1806) & (g1807)) + ((sk[1]) & (g816) & (!g1163) & (g1725) & (!g1806) & (!g1807)) + ((sk[1]) & (g816) & (!g1163) & (g1725) & (g1806) & (!g1807)) + ((sk[1]) & (g816) & (g1163) & (!g1725) & (!g1806) & (!g1807)) + ((sk[1]) & (g816) & (g1163) & (!g1725) & (!g1806) & (g1807)) + ((sk[1]) & (g816) & (g1163) & (g1725) & (!g1806) & (!g1807)) + ((sk[1]) & (g816) & (g1163) & (g1725) & (!g1806) & (g1807)));
	assign g2201 = (((!ld) & (!sk[2]) & (text_inx87x) & (!g1809)) + ((!ld) & (!sk[2]) & (text_inx87x) & (g1809)) + ((!ld) & (sk[2]) & (!text_inx87x) & (g1809)) + ((!ld) & (sk[2]) & (text_inx87x) & (g1809)) + ((ld) & (!sk[2]) & (!text_inx87x) & (g1809)) + ((ld) & (!sk[2]) & (text_inx87x) & (!g1809)) + ((ld) & (!sk[2]) & (text_inx87x) & (g1809)) + ((ld) & (sk[2]) & (text_inx87x) & (!g1809)) + ((ld) & (sk[2]) & (text_inx87x) & (g1809)));
	assign g1810 = (((!ld) & (!sk[3]) & (!g1044) & (g1358) & (!keyx112x)) + ((!ld) & (!sk[3]) & (!g1044) & (g1358) & (keyx112x)) + ((!ld) & (!sk[3]) & (g1044) & (!g1358) & (!keyx112x)) + ((!ld) & (!sk[3]) & (g1044) & (!g1358) & (keyx112x)) + ((!ld) & (!sk[3]) & (g1044) & (g1358) & (!keyx112x)) + ((!ld) & (!sk[3]) & (g1044) & (g1358) & (keyx112x)) + ((!ld) & (sk[3]) & (!g1044) & (g1358) & (!keyx112x)) + ((!ld) & (sk[3]) & (!g1044) & (g1358) & (keyx112x)) + ((!ld) & (sk[3]) & (g1044) & (!g1358) & (!keyx112x)) + ((!ld) & (sk[3]) & (g1044) & (!g1358) & (keyx112x)) + ((ld) & (!sk[3]) & (!g1044) & (g1358) & (!keyx112x)) + ((ld) & (!sk[3]) & (!g1044) & (g1358) & (keyx112x)) + ((ld) & (!sk[3]) & (g1044) & (!g1358) & (!keyx112x)) + ((ld) & (!sk[3]) & (g1044) & (!g1358) & (keyx112x)) + ((ld) & (!sk[3]) & (g1044) & (g1358) & (!keyx112x)) + ((ld) & (!sk[3]) & (g1044) & (g1358) & (keyx112x)) + ((ld) & (sk[3]) & (!g1044) & (!g1358) & (keyx112x)) + ((ld) & (sk[3]) & (!g1044) & (g1358) & (keyx112x)) + ((ld) & (sk[3]) & (g1044) & (!g1358) & (keyx112x)) + ((ld) & (sk[3]) & (g1044) & (g1358) & (keyx112x)));
	assign g1811 = (((!ld) & (!sk[4]) & (!g1051) & (g1365) & (!keyx113x)) + ((!ld) & (!sk[4]) & (!g1051) & (g1365) & (keyx113x)) + ((!ld) & (!sk[4]) & (g1051) & (!g1365) & (!keyx113x)) + ((!ld) & (!sk[4]) & (g1051) & (!g1365) & (keyx113x)) + ((!ld) & (!sk[4]) & (g1051) & (g1365) & (!keyx113x)) + ((!ld) & (!sk[4]) & (g1051) & (g1365) & (keyx113x)) + ((!ld) & (sk[4]) & (!g1051) & (g1365) & (!keyx113x)) + ((!ld) & (sk[4]) & (!g1051) & (g1365) & (keyx113x)) + ((!ld) & (sk[4]) & (g1051) & (!g1365) & (!keyx113x)) + ((!ld) & (sk[4]) & (g1051) & (!g1365) & (keyx113x)) + ((ld) & (!sk[4]) & (!g1051) & (g1365) & (!keyx113x)) + ((ld) & (!sk[4]) & (!g1051) & (g1365) & (keyx113x)) + ((ld) & (!sk[4]) & (g1051) & (!g1365) & (!keyx113x)) + ((ld) & (!sk[4]) & (g1051) & (!g1365) & (keyx113x)) + ((ld) & (!sk[4]) & (g1051) & (g1365) & (!keyx113x)) + ((ld) & (!sk[4]) & (g1051) & (g1365) & (keyx113x)) + ((ld) & (sk[4]) & (!g1051) & (!g1365) & (keyx113x)) + ((ld) & (sk[4]) & (!g1051) & (g1365) & (keyx113x)) + ((ld) & (sk[4]) & (g1051) & (!g1365) & (keyx113x)) + ((ld) & (sk[4]) & (g1051) & (g1365) & (keyx113x)));
	assign g1812 = (((!ld) & (!sk[5]) & (!g1058) & (g1372) & (!keyx114x)) + ((!ld) & (!sk[5]) & (!g1058) & (g1372) & (keyx114x)) + ((!ld) & (!sk[5]) & (g1058) & (!g1372) & (!keyx114x)) + ((!ld) & (!sk[5]) & (g1058) & (!g1372) & (keyx114x)) + ((!ld) & (!sk[5]) & (g1058) & (g1372) & (!keyx114x)) + ((!ld) & (!sk[5]) & (g1058) & (g1372) & (keyx114x)) + ((!ld) & (sk[5]) & (!g1058) & (g1372) & (!keyx114x)) + ((!ld) & (sk[5]) & (!g1058) & (g1372) & (keyx114x)) + ((!ld) & (sk[5]) & (g1058) & (!g1372) & (!keyx114x)) + ((!ld) & (sk[5]) & (g1058) & (!g1372) & (keyx114x)) + ((ld) & (!sk[5]) & (!g1058) & (g1372) & (!keyx114x)) + ((ld) & (!sk[5]) & (!g1058) & (g1372) & (keyx114x)) + ((ld) & (!sk[5]) & (g1058) & (!g1372) & (!keyx114x)) + ((ld) & (!sk[5]) & (g1058) & (!g1372) & (keyx114x)) + ((ld) & (!sk[5]) & (g1058) & (g1372) & (!keyx114x)) + ((ld) & (!sk[5]) & (g1058) & (g1372) & (keyx114x)) + ((ld) & (sk[5]) & (!g1058) & (!g1372) & (keyx114x)) + ((ld) & (sk[5]) & (!g1058) & (g1372) & (keyx114x)) + ((ld) & (sk[5]) & (g1058) & (!g1372) & (keyx114x)) + ((ld) & (sk[5]) & (g1058) & (g1372) & (keyx114x)));
	assign g1813 = (((!ld) & (!sk[6]) & (!g1065) & (g1379) & (!keyx115x)) + ((!ld) & (!sk[6]) & (!g1065) & (g1379) & (keyx115x)) + ((!ld) & (!sk[6]) & (g1065) & (!g1379) & (!keyx115x)) + ((!ld) & (!sk[6]) & (g1065) & (!g1379) & (keyx115x)) + ((!ld) & (!sk[6]) & (g1065) & (g1379) & (!keyx115x)) + ((!ld) & (!sk[6]) & (g1065) & (g1379) & (keyx115x)) + ((!ld) & (sk[6]) & (!g1065) & (g1379) & (!keyx115x)) + ((!ld) & (sk[6]) & (!g1065) & (g1379) & (keyx115x)) + ((!ld) & (sk[6]) & (g1065) & (!g1379) & (!keyx115x)) + ((!ld) & (sk[6]) & (g1065) & (!g1379) & (keyx115x)) + ((ld) & (!sk[6]) & (!g1065) & (g1379) & (!keyx115x)) + ((ld) & (!sk[6]) & (!g1065) & (g1379) & (keyx115x)) + ((ld) & (!sk[6]) & (g1065) & (!g1379) & (!keyx115x)) + ((ld) & (!sk[6]) & (g1065) & (!g1379) & (keyx115x)) + ((ld) & (!sk[6]) & (g1065) & (g1379) & (!keyx115x)) + ((ld) & (!sk[6]) & (g1065) & (g1379) & (keyx115x)) + ((ld) & (sk[6]) & (!g1065) & (!g1379) & (keyx115x)) + ((ld) & (sk[6]) & (!g1065) & (g1379) & (keyx115x)) + ((ld) & (sk[6]) & (g1065) & (!g1379) & (keyx115x)) + ((ld) & (sk[6]) & (g1065) & (g1379) & (keyx115x)));
	assign g1814 = (((!ld) & (!g1072) & (g1386) & (!sk[7]) & (!keyx116x)) + ((!ld) & (!g1072) & (g1386) & (!sk[7]) & (keyx116x)) + ((!ld) & (!g1072) & (g1386) & (sk[7]) & (!keyx116x)) + ((!ld) & (!g1072) & (g1386) & (sk[7]) & (keyx116x)) + ((!ld) & (g1072) & (!g1386) & (!sk[7]) & (!keyx116x)) + ((!ld) & (g1072) & (!g1386) & (!sk[7]) & (keyx116x)) + ((!ld) & (g1072) & (!g1386) & (sk[7]) & (!keyx116x)) + ((!ld) & (g1072) & (!g1386) & (sk[7]) & (keyx116x)) + ((!ld) & (g1072) & (g1386) & (!sk[7]) & (!keyx116x)) + ((!ld) & (g1072) & (g1386) & (!sk[7]) & (keyx116x)) + ((ld) & (!g1072) & (!g1386) & (sk[7]) & (keyx116x)) + ((ld) & (!g1072) & (g1386) & (!sk[7]) & (!keyx116x)) + ((ld) & (!g1072) & (g1386) & (!sk[7]) & (keyx116x)) + ((ld) & (!g1072) & (g1386) & (sk[7]) & (keyx116x)) + ((ld) & (g1072) & (!g1386) & (!sk[7]) & (!keyx116x)) + ((ld) & (g1072) & (!g1386) & (!sk[7]) & (keyx116x)) + ((ld) & (g1072) & (!g1386) & (sk[7]) & (keyx116x)) + ((ld) & (g1072) & (g1386) & (!sk[7]) & (!keyx116x)) + ((ld) & (g1072) & (g1386) & (!sk[7]) & (keyx116x)) + ((ld) & (g1072) & (g1386) & (sk[7]) & (keyx116x)));
	assign g1815 = (((!ld) & (!sk[8]) & (!g1079) & (g1393) & (!keyx117x)) + ((!ld) & (!sk[8]) & (!g1079) & (g1393) & (keyx117x)) + ((!ld) & (!sk[8]) & (g1079) & (!g1393) & (!keyx117x)) + ((!ld) & (!sk[8]) & (g1079) & (!g1393) & (keyx117x)) + ((!ld) & (!sk[8]) & (g1079) & (g1393) & (!keyx117x)) + ((!ld) & (!sk[8]) & (g1079) & (g1393) & (keyx117x)) + ((!ld) & (sk[8]) & (!g1079) & (g1393) & (!keyx117x)) + ((!ld) & (sk[8]) & (!g1079) & (g1393) & (keyx117x)) + ((!ld) & (sk[8]) & (g1079) & (!g1393) & (!keyx117x)) + ((!ld) & (sk[8]) & (g1079) & (!g1393) & (keyx117x)) + ((ld) & (!sk[8]) & (!g1079) & (g1393) & (!keyx117x)) + ((ld) & (!sk[8]) & (!g1079) & (g1393) & (keyx117x)) + ((ld) & (!sk[8]) & (g1079) & (!g1393) & (!keyx117x)) + ((ld) & (!sk[8]) & (g1079) & (!g1393) & (keyx117x)) + ((ld) & (!sk[8]) & (g1079) & (g1393) & (!keyx117x)) + ((ld) & (!sk[8]) & (g1079) & (g1393) & (keyx117x)) + ((ld) & (sk[8]) & (!g1079) & (!g1393) & (keyx117x)) + ((ld) & (sk[8]) & (!g1079) & (g1393) & (keyx117x)) + ((ld) & (sk[8]) & (g1079) & (!g1393) & (keyx117x)) + ((ld) & (sk[8]) & (g1079) & (g1393) & (keyx117x)));
	assign g1816 = (((!ld) & (!sk[9]) & (!g1086) & (g1400) & (!keyx118x)) + ((!ld) & (!sk[9]) & (!g1086) & (g1400) & (keyx118x)) + ((!ld) & (!sk[9]) & (g1086) & (!g1400) & (!keyx118x)) + ((!ld) & (!sk[9]) & (g1086) & (!g1400) & (keyx118x)) + ((!ld) & (!sk[9]) & (g1086) & (g1400) & (!keyx118x)) + ((!ld) & (!sk[9]) & (g1086) & (g1400) & (keyx118x)) + ((!ld) & (sk[9]) & (!g1086) & (g1400) & (!keyx118x)) + ((!ld) & (sk[9]) & (!g1086) & (g1400) & (keyx118x)) + ((!ld) & (sk[9]) & (g1086) & (!g1400) & (!keyx118x)) + ((!ld) & (sk[9]) & (g1086) & (!g1400) & (keyx118x)) + ((ld) & (!sk[9]) & (!g1086) & (g1400) & (!keyx118x)) + ((ld) & (!sk[9]) & (!g1086) & (g1400) & (keyx118x)) + ((ld) & (!sk[9]) & (g1086) & (!g1400) & (!keyx118x)) + ((ld) & (!sk[9]) & (g1086) & (!g1400) & (keyx118x)) + ((ld) & (!sk[9]) & (g1086) & (g1400) & (!keyx118x)) + ((ld) & (!sk[9]) & (g1086) & (g1400) & (keyx118x)) + ((ld) & (sk[9]) & (!g1086) & (!g1400) & (keyx118x)) + ((ld) & (sk[9]) & (!g1086) & (g1400) & (keyx118x)) + ((ld) & (sk[9]) & (g1086) & (!g1400) & (keyx118x)) + ((ld) & (sk[9]) & (g1086) & (g1400) & (keyx118x)));
	assign g1817 = (((!ld) & (!g1093) & (!sk[10]) & (g1407) & (!keyx119x)) + ((!ld) & (!g1093) & (!sk[10]) & (g1407) & (keyx119x)) + ((!ld) & (!g1093) & (sk[10]) & (g1407) & (!keyx119x)) + ((!ld) & (!g1093) & (sk[10]) & (g1407) & (keyx119x)) + ((!ld) & (g1093) & (!sk[10]) & (!g1407) & (!keyx119x)) + ((!ld) & (g1093) & (!sk[10]) & (!g1407) & (keyx119x)) + ((!ld) & (g1093) & (!sk[10]) & (g1407) & (!keyx119x)) + ((!ld) & (g1093) & (!sk[10]) & (g1407) & (keyx119x)) + ((!ld) & (g1093) & (sk[10]) & (!g1407) & (!keyx119x)) + ((!ld) & (g1093) & (sk[10]) & (!g1407) & (keyx119x)) + ((ld) & (!g1093) & (!sk[10]) & (g1407) & (!keyx119x)) + ((ld) & (!g1093) & (!sk[10]) & (g1407) & (keyx119x)) + ((ld) & (!g1093) & (sk[10]) & (!g1407) & (keyx119x)) + ((ld) & (!g1093) & (sk[10]) & (g1407) & (keyx119x)) + ((ld) & (g1093) & (!sk[10]) & (!g1407) & (!keyx119x)) + ((ld) & (g1093) & (!sk[10]) & (!g1407) & (keyx119x)) + ((ld) & (g1093) & (!sk[10]) & (g1407) & (!keyx119x)) + ((ld) & (g1093) & (!sk[10]) & (g1407) & (keyx119x)) + ((ld) & (g1093) & (sk[10]) & (!g1407) & (keyx119x)) + ((ld) & (g1093) & (sk[10]) & (g1407) & (keyx119x)));
	assign g2202 = (((!sk[11]) & (!ld) & (text_inx120x) & (!g1818)) + ((!sk[11]) & (!ld) & (text_inx120x) & (g1818)) + ((!sk[11]) & (ld) & (!text_inx120x) & (g1818)) + ((!sk[11]) & (ld) & (text_inx120x) & (!g1818)) + ((!sk[11]) & (ld) & (text_inx120x) & (g1818)) + ((sk[11]) & (!ld) & (!text_inx120x) & (g1818)) + ((sk[11]) & (!ld) & (text_inx120x) & (g1818)) + ((sk[11]) & (ld) & (text_inx120x) & (!g1818)) + ((sk[11]) & (ld) & (text_inx120x) & (g1818)));
	assign g1819 = (((!sk[12]) & (!g1043) & (g1092) & (!g1156)) + ((!sk[12]) & (!g1043) & (g1092) & (g1156)) + ((!sk[12]) & (g1043) & (!g1092) & (g1156)) + ((!sk[12]) & (g1043) & (g1092) & (!g1156)) + ((!sk[12]) & (g1043) & (g1092) & (g1156)) + ((sk[12]) & (!g1043) & (!g1092) & (g1156)) + ((sk[12]) & (!g1043) & (g1092) & (!g1156)) + ((sk[12]) & (g1043) & (!g1092) & (!g1156)) + ((sk[12]) & (g1043) & (g1092) & (g1156)));
	assign g1820 = (((!g1108) & (!g1163) & (!g1330) & (!g1818) & (sk[13]) & (g1819)) + ((!g1108) & (!g1163) & (!g1330) & (g1818) & (sk[13]) & (g1819)) + ((!g1108) & (!g1163) & (g1330) & (!g1818) & (sk[13]) & (!g1819)) + ((!g1108) & (!g1163) & (g1330) & (g1818) & (sk[13]) & (!g1819)) + ((!g1108) & (g1163) & (!g1330) & (!g1818) & (!sk[13]) & (!g1819)) + ((!g1108) & (g1163) & (!g1330) & (!g1818) & (!sk[13]) & (g1819)) + ((!g1108) & (g1163) & (!g1330) & (g1818) & (!sk[13]) & (!g1819)) + ((!g1108) & (g1163) & (!g1330) & (g1818) & (!sk[13]) & (g1819)) + ((!g1108) & (g1163) & (!g1330) & (g1818) & (sk[13]) & (!g1819)) + ((!g1108) & (g1163) & (!g1330) & (g1818) & (sk[13]) & (g1819)) + ((!g1108) & (g1163) & (g1330) & (!g1818) & (!sk[13]) & (!g1819)) + ((!g1108) & (g1163) & (g1330) & (!g1818) & (!sk[13]) & (g1819)) + ((!g1108) & (g1163) & (g1330) & (g1818) & (!sk[13]) & (!g1819)) + ((!g1108) & (g1163) & (g1330) & (g1818) & (!sk[13]) & (g1819)) + ((!g1108) & (g1163) & (g1330) & (g1818) & (sk[13]) & (!g1819)) + ((!g1108) & (g1163) & (g1330) & (g1818) & (sk[13]) & (g1819)) + ((g1108) & (!g1163) & (!g1330) & (!g1818) & (!sk[13]) & (!g1819)) + ((g1108) & (!g1163) & (!g1330) & (!g1818) & (!sk[13]) & (g1819)) + ((g1108) & (!g1163) & (!g1330) & (!g1818) & (sk[13]) & (!g1819)) + ((g1108) & (!g1163) & (!g1330) & (g1818) & (!sk[13]) & (!g1819)) + ((g1108) & (!g1163) & (!g1330) & (g1818) & (!sk[13]) & (g1819)) + ((g1108) & (!g1163) & (!g1330) & (g1818) & (sk[13]) & (!g1819)) + ((g1108) & (!g1163) & (g1330) & (!g1818) & (!sk[13]) & (!g1819)) + ((g1108) & (!g1163) & (g1330) & (!g1818) & (!sk[13]) & (g1819)) + ((g1108) & (!g1163) & (g1330) & (!g1818) & (sk[13]) & (g1819)) + ((g1108) & (!g1163) & (g1330) & (g1818) & (!sk[13]) & (!g1819)) + ((g1108) & (!g1163) & (g1330) & (g1818) & (!sk[13]) & (g1819)) + ((g1108) & (!g1163) & (g1330) & (g1818) & (sk[13]) & (g1819)) + ((g1108) & (g1163) & (!g1330) & (!g1818) & (!sk[13]) & (!g1819)) + ((g1108) & (g1163) & (!g1330) & (!g1818) & (!sk[13]) & (g1819)) + ((g1108) & (g1163) & (!g1330) & (!g1818) & (sk[13]) & (!g1819)) + ((g1108) & (g1163) & (!g1330) & (!g1818) & (sk[13]) & (g1819)) + ((g1108) & (g1163) & (!g1330) & (g1818) & (!sk[13]) & (!g1819)) + ((g1108) & (g1163) & (!g1330) & (g1818) & (!sk[13]) & (g1819)) + ((g1108) & (g1163) & (g1330) & (!g1818) & (!sk[13]) & (!g1819)) + ((g1108) & (g1163) & (g1330) & (!g1818) & (!sk[13]) & (g1819)) + ((g1108) & (g1163) & (g1330) & (!g1818) & (sk[13]) & (!g1819)) + ((g1108) & (g1163) & (g1330) & (!g1818) & (sk[13]) & (g1819)) + ((g1108) & (g1163) & (g1330) & (g1818) & (!sk[13]) & (!g1819)) + ((g1108) & (g1163) & (g1330) & (g1818) & (!sk[13]) & (g1819)));
	assign g2203 = (((!ld) & (!sk[14]) & (text_inx121x) & (!g1821)) + ((!ld) & (!sk[14]) & (text_inx121x) & (g1821)) + ((!ld) & (sk[14]) & (!text_inx121x) & (g1821)) + ((!ld) & (sk[14]) & (text_inx121x) & (g1821)) + ((ld) & (!sk[14]) & (!text_inx121x) & (g1821)) + ((ld) & (!sk[14]) & (text_inx121x) & (!g1821)) + ((ld) & (!sk[14]) & (text_inx121x) & (g1821)) + ((ld) & (sk[14]) & (text_inx121x) & (!g1821)) + ((ld) & (sk[14]) & (text_inx121x) & (g1821)));
	assign g1822 = (((!g922) & (!g1115) & (!g1163) & (!g1622) & (g1819) & (!g1821)) + ((!g922) & (!g1115) & (!g1163) & (!g1622) & (g1819) & (g1821)) + ((!g922) & (!g1115) & (!g1163) & (g1622) & (!g1819) & (!g1821)) + ((!g922) & (!g1115) & (!g1163) & (g1622) & (!g1819) & (g1821)) + ((!g922) & (!g1115) & (g1163) & (!g1622) & (!g1819) & (g1821)) + ((!g922) & (!g1115) & (g1163) & (!g1622) & (g1819) & (g1821)) + ((!g922) & (!g1115) & (g1163) & (g1622) & (!g1819) & (g1821)) + ((!g922) & (!g1115) & (g1163) & (g1622) & (g1819) & (g1821)) + ((!g922) & (g1115) & (!g1163) & (!g1622) & (!g1819) & (!g1821)) + ((!g922) & (g1115) & (!g1163) & (!g1622) & (!g1819) & (g1821)) + ((!g922) & (g1115) & (!g1163) & (g1622) & (g1819) & (!g1821)) + ((!g922) & (g1115) & (!g1163) & (g1622) & (g1819) & (g1821)) + ((!g922) & (g1115) & (g1163) & (!g1622) & (!g1819) & (!g1821)) + ((!g922) & (g1115) & (g1163) & (!g1622) & (g1819) & (!g1821)) + ((!g922) & (g1115) & (g1163) & (g1622) & (!g1819) & (!g1821)) + ((!g922) & (g1115) & (g1163) & (g1622) & (g1819) & (!g1821)) + ((g922) & (!g1115) & (!g1163) & (!g1622) & (!g1819) & (!g1821)) + ((g922) & (!g1115) & (!g1163) & (!g1622) & (!g1819) & (g1821)) + ((g922) & (!g1115) & (!g1163) & (g1622) & (g1819) & (!g1821)) + ((g922) & (!g1115) & (!g1163) & (g1622) & (g1819) & (g1821)) + ((g922) & (!g1115) & (g1163) & (!g1622) & (!g1819) & (g1821)) + ((g922) & (!g1115) & (g1163) & (!g1622) & (g1819) & (g1821)) + ((g922) & (!g1115) & (g1163) & (g1622) & (!g1819) & (g1821)) + ((g922) & (!g1115) & (g1163) & (g1622) & (g1819) & (g1821)) + ((g922) & (g1115) & (!g1163) & (!g1622) & (g1819) & (!g1821)) + ((g922) & (g1115) & (!g1163) & (!g1622) & (g1819) & (g1821)) + ((g922) & (g1115) & (!g1163) & (g1622) & (!g1819) & (!g1821)) + ((g922) & (g1115) & (!g1163) & (g1622) & (!g1819) & (g1821)) + ((g922) & (g1115) & (g1163) & (!g1622) & (!g1819) & (!g1821)) + ((g922) & (g1115) & (g1163) & (!g1622) & (g1819) & (!g1821)) + ((g922) & (g1115) & (g1163) & (g1622) & (!g1819) & (!g1821)) + ((g922) & (g1115) & (g1163) & (g1622) & (g1819) & (!g1821)));
	assign g2204 = (((!ld) & (!sk[16]) & (text_inx122x) & (!g1823)) + ((!ld) & (!sk[16]) & (text_inx122x) & (g1823)) + ((!ld) & (sk[16]) & (!text_inx122x) & (g1823)) + ((!ld) & (sk[16]) & (text_inx122x) & (g1823)) + ((ld) & (!sk[16]) & (!text_inx122x) & (g1823)) + ((ld) & (!sk[16]) & (text_inx122x) & (!g1823)) + ((ld) & (!sk[16]) & (text_inx122x) & (g1823)) + ((ld) & (sk[16]) & (text_inx122x) & (!g1823)) + ((ld) & (sk[16]) & (text_inx122x) & (g1823)));
	assign g1824 = (((!g1057) & (!g1114) & (!g1122) & (!g1163) & (g1337) & (!g1823)) + ((!g1057) & (!g1114) & (!g1122) & (!g1163) & (g1337) & (g1823)) + ((!g1057) & (!g1114) & (!g1122) & (g1163) & (!g1337) & (g1823)) + ((!g1057) & (!g1114) & (!g1122) & (g1163) & (g1337) & (g1823)) + ((!g1057) & (!g1114) & (g1122) & (!g1163) & (!g1337) & (!g1823)) + ((!g1057) & (!g1114) & (g1122) & (!g1163) & (!g1337) & (g1823)) + ((!g1057) & (!g1114) & (g1122) & (g1163) & (!g1337) & (!g1823)) + ((!g1057) & (!g1114) & (g1122) & (g1163) & (g1337) & (!g1823)) + ((!g1057) & (g1114) & (!g1122) & (!g1163) & (!g1337) & (!g1823)) + ((!g1057) & (g1114) & (!g1122) & (!g1163) & (!g1337) & (g1823)) + ((!g1057) & (g1114) & (!g1122) & (g1163) & (!g1337) & (g1823)) + ((!g1057) & (g1114) & (!g1122) & (g1163) & (g1337) & (g1823)) + ((!g1057) & (g1114) & (g1122) & (!g1163) & (g1337) & (!g1823)) + ((!g1057) & (g1114) & (g1122) & (!g1163) & (g1337) & (g1823)) + ((!g1057) & (g1114) & (g1122) & (g1163) & (!g1337) & (!g1823)) + ((!g1057) & (g1114) & (g1122) & (g1163) & (g1337) & (!g1823)) + ((g1057) & (!g1114) & (!g1122) & (!g1163) & (!g1337) & (!g1823)) + ((g1057) & (!g1114) & (!g1122) & (!g1163) & (!g1337) & (g1823)) + ((g1057) & (!g1114) & (!g1122) & (g1163) & (!g1337) & (g1823)) + ((g1057) & (!g1114) & (!g1122) & (g1163) & (g1337) & (g1823)) + ((g1057) & (!g1114) & (g1122) & (!g1163) & (g1337) & (!g1823)) + ((g1057) & (!g1114) & (g1122) & (!g1163) & (g1337) & (g1823)) + ((g1057) & (!g1114) & (g1122) & (g1163) & (!g1337) & (!g1823)) + ((g1057) & (!g1114) & (g1122) & (g1163) & (g1337) & (!g1823)) + ((g1057) & (g1114) & (!g1122) & (!g1163) & (g1337) & (!g1823)) + ((g1057) & (g1114) & (!g1122) & (!g1163) & (g1337) & (g1823)) + ((g1057) & (g1114) & (!g1122) & (g1163) & (!g1337) & (g1823)) + ((g1057) & (g1114) & (!g1122) & (g1163) & (g1337) & (g1823)) + ((g1057) & (g1114) & (g1122) & (!g1163) & (!g1337) & (!g1823)) + ((g1057) & (g1114) & (g1122) & (!g1163) & (!g1337) & (g1823)) + ((g1057) & (g1114) & (g1122) & (g1163) & (!g1337) & (!g1823)) + ((g1057) & (g1114) & (g1122) & (g1163) & (g1337) & (!g1823)));
	assign g2205 = (((!ld) & (!text_inx123x) & (sk[18]) & (g1825)) + ((!ld) & (text_inx123x) & (!sk[18]) & (!g1825)) + ((!ld) & (text_inx123x) & (!sk[18]) & (g1825)) + ((!ld) & (text_inx123x) & (sk[18]) & (g1825)) + ((ld) & (!text_inx123x) & (!sk[18]) & (g1825)) + ((ld) & (text_inx123x) & (!sk[18]) & (!g1825)) + ((ld) & (text_inx123x) & (!sk[18]) & (g1825)) + ((ld) & (text_inx123x) & (sk[18]) & (!g1825)) + ((ld) & (text_inx123x) & (sk[18]) & (g1825)));
	assign g2206 = (((!sk[19]) & (!ld) & (text_inx126x) & (!g1826)) + ((!sk[19]) & (!ld) & (text_inx126x) & (g1826)) + ((!sk[19]) & (ld) & (!text_inx126x) & (g1826)) + ((!sk[19]) & (ld) & (text_inx126x) & (!g1826)) + ((!sk[19]) & (ld) & (text_inx126x) & (g1826)) + ((sk[19]) & (!ld) & (!text_inx126x) & (g1826)) + ((sk[19]) & (!ld) & (text_inx126x) & (g1826)) + ((sk[19]) & (ld) & (text_inx126x) & (!g1826)) + ((sk[19]) & (ld) & (text_inx126x) & (g1826)));
	assign g1827 = (((!g1085) & (!g1142) & (!g1150) & (!g1163) & (g1342) & (!g1826)) + ((!g1085) & (!g1142) & (!g1150) & (!g1163) & (g1342) & (g1826)) + ((!g1085) & (!g1142) & (!g1150) & (g1163) & (!g1342) & (g1826)) + ((!g1085) & (!g1142) & (!g1150) & (g1163) & (g1342) & (g1826)) + ((!g1085) & (!g1142) & (g1150) & (!g1163) & (!g1342) & (!g1826)) + ((!g1085) & (!g1142) & (g1150) & (!g1163) & (!g1342) & (g1826)) + ((!g1085) & (!g1142) & (g1150) & (g1163) & (!g1342) & (!g1826)) + ((!g1085) & (!g1142) & (g1150) & (g1163) & (g1342) & (!g1826)) + ((!g1085) & (g1142) & (!g1150) & (!g1163) & (!g1342) & (!g1826)) + ((!g1085) & (g1142) & (!g1150) & (!g1163) & (!g1342) & (g1826)) + ((!g1085) & (g1142) & (!g1150) & (g1163) & (!g1342) & (g1826)) + ((!g1085) & (g1142) & (!g1150) & (g1163) & (g1342) & (g1826)) + ((!g1085) & (g1142) & (g1150) & (!g1163) & (g1342) & (!g1826)) + ((!g1085) & (g1142) & (g1150) & (!g1163) & (g1342) & (g1826)) + ((!g1085) & (g1142) & (g1150) & (g1163) & (!g1342) & (!g1826)) + ((!g1085) & (g1142) & (g1150) & (g1163) & (g1342) & (!g1826)) + ((g1085) & (!g1142) & (!g1150) & (!g1163) & (!g1342) & (!g1826)) + ((g1085) & (!g1142) & (!g1150) & (!g1163) & (!g1342) & (g1826)) + ((g1085) & (!g1142) & (!g1150) & (g1163) & (!g1342) & (g1826)) + ((g1085) & (!g1142) & (!g1150) & (g1163) & (g1342) & (g1826)) + ((g1085) & (!g1142) & (g1150) & (!g1163) & (g1342) & (!g1826)) + ((g1085) & (!g1142) & (g1150) & (!g1163) & (g1342) & (g1826)) + ((g1085) & (!g1142) & (g1150) & (g1163) & (!g1342) & (!g1826)) + ((g1085) & (!g1142) & (g1150) & (g1163) & (g1342) & (!g1826)) + ((g1085) & (g1142) & (!g1150) & (!g1163) & (g1342) & (!g1826)) + ((g1085) & (g1142) & (!g1150) & (!g1163) & (g1342) & (g1826)) + ((g1085) & (g1142) & (!g1150) & (g1163) & (!g1342) & (g1826)) + ((g1085) & (g1142) & (!g1150) & (g1163) & (g1342) & (g1826)) + ((g1085) & (g1142) & (g1150) & (!g1163) & (!g1342) & (!g1826)) + ((g1085) & (g1142) & (g1150) & (!g1163) & (!g1342) & (g1826)) + ((g1085) & (g1142) & (g1150) & (g1163) & (!g1342) & (!g1826)) + ((g1085) & (g1142) & (g1150) & (g1163) & (g1342) & (!g1826)));
	assign g2207 = (((!sk[21]) & (!ld) & (text_inx125x) & (!g1828)) + ((!sk[21]) & (!ld) & (text_inx125x) & (g1828)) + ((!sk[21]) & (ld) & (!text_inx125x) & (g1828)) + ((!sk[21]) & (ld) & (text_inx125x) & (!g1828)) + ((!sk[21]) & (ld) & (text_inx125x) & (g1828)) + ((sk[21]) & (!ld) & (!text_inx125x) & (g1828)) + ((sk[21]) & (!ld) & (text_inx125x) & (g1828)) + ((sk[21]) & (ld) & (text_inx125x) & (!g1828)) + ((sk[21]) & (ld) & (text_inx125x) & (g1828)));
	assign g1829 = (((!g1078) & (!g1135) & (!g1143) & (!g1163) & (g1345) & (!g1828)) + ((!g1078) & (!g1135) & (!g1143) & (!g1163) & (g1345) & (g1828)) + ((!g1078) & (!g1135) & (!g1143) & (g1163) & (!g1345) & (g1828)) + ((!g1078) & (!g1135) & (!g1143) & (g1163) & (g1345) & (g1828)) + ((!g1078) & (!g1135) & (g1143) & (!g1163) & (!g1345) & (!g1828)) + ((!g1078) & (!g1135) & (g1143) & (!g1163) & (!g1345) & (g1828)) + ((!g1078) & (!g1135) & (g1143) & (g1163) & (!g1345) & (!g1828)) + ((!g1078) & (!g1135) & (g1143) & (g1163) & (g1345) & (!g1828)) + ((!g1078) & (g1135) & (!g1143) & (!g1163) & (!g1345) & (!g1828)) + ((!g1078) & (g1135) & (!g1143) & (!g1163) & (!g1345) & (g1828)) + ((!g1078) & (g1135) & (!g1143) & (g1163) & (!g1345) & (g1828)) + ((!g1078) & (g1135) & (!g1143) & (g1163) & (g1345) & (g1828)) + ((!g1078) & (g1135) & (g1143) & (!g1163) & (g1345) & (!g1828)) + ((!g1078) & (g1135) & (g1143) & (!g1163) & (g1345) & (g1828)) + ((!g1078) & (g1135) & (g1143) & (g1163) & (!g1345) & (!g1828)) + ((!g1078) & (g1135) & (g1143) & (g1163) & (g1345) & (!g1828)) + ((g1078) & (!g1135) & (!g1143) & (!g1163) & (!g1345) & (!g1828)) + ((g1078) & (!g1135) & (!g1143) & (!g1163) & (!g1345) & (g1828)) + ((g1078) & (!g1135) & (!g1143) & (g1163) & (!g1345) & (g1828)) + ((g1078) & (!g1135) & (!g1143) & (g1163) & (g1345) & (g1828)) + ((g1078) & (!g1135) & (g1143) & (!g1163) & (g1345) & (!g1828)) + ((g1078) & (!g1135) & (g1143) & (!g1163) & (g1345) & (g1828)) + ((g1078) & (!g1135) & (g1143) & (g1163) & (!g1345) & (!g1828)) + ((g1078) & (!g1135) & (g1143) & (g1163) & (g1345) & (!g1828)) + ((g1078) & (g1135) & (!g1143) & (!g1163) & (g1345) & (!g1828)) + ((g1078) & (g1135) & (!g1143) & (!g1163) & (g1345) & (g1828)) + ((g1078) & (g1135) & (!g1143) & (g1163) & (!g1345) & (g1828)) + ((g1078) & (g1135) & (!g1143) & (g1163) & (g1345) & (g1828)) + ((g1078) & (g1135) & (g1143) & (!g1163) & (!g1345) & (!g1828)) + ((g1078) & (g1135) & (g1143) & (!g1163) & (!g1345) & (g1828)) + ((g1078) & (g1135) & (g1143) & (g1163) & (!g1345) & (!g1828)) + ((g1078) & (g1135) & (g1143) & (g1163) & (g1345) & (!g1828)));
	assign g2208 = (((!sk[23]) & (!ld) & (text_inx124x) & (!g1830)) + ((!sk[23]) & (!ld) & (text_inx124x) & (g1830)) + ((!sk[23]) & (ld) & (!text_inx124x) & (g1830)) + ((!sk[23]) & (ld) & (text_inx124x) & (!g1830)) + ((!sk[23]) & (ld) & (text_inx124x) & (g1830)) + ((sk[23]) & (!ld) & (!text_inx124x) & (g1830)) + ((sk[23]) & (!ld) & (text_inx124x) & (g1830)) + ((sk[23]) & (ld) & (text_inx124x) & (!g1830)) + ((sk[23]) & (ld) & (text_inx124x) & (g1830)));
	assign g1831 = (((!sk[24]) & (!g1085) & (g1149)) + ((!sk[24]) & (g1085) & (g1149)) + ((sk[24]) & (!g1085) & (g1149)) + ((sk[24]) & (g1085) & (!g1149)));
	assign g2209 = (((!ld) & (!sk[25]) & (text_inx127x) & (!g1832)) + ((!ld) & (!sk[25]) & (text_inx127x) & (g1832)) + ((!ld) & (sk[25]) & (!text_inx127x) & (g1832)) + ((!ld) & (sk[25]) & (text_inx127x) & (g1832)) + ((ld) & (!sk[25]) & (!text_inx127x) & (g1832)) + ((ld) & (!sk[25]) & (text_inx127x) & (!g1832)) + ((ld) & (!sk[25]) & (text_inx127x) & (g1832)) + ((ld) & (sk[25]) & (text_inx127x) & (!g1832)) + ((ld) & (sk[25]) & (text_inx127x) & (g1832)));
	assign g1833 = (((!g964) & (!g1157) & (!g1163) & (!g1329) & (g1831) & (!g1832)) + ((!g964) & (!g1157) & (!g1163) & (!g1329) & (g1831) & (g1832)) + ((!g964) & (!g1157) & (!g1163) & (g1329) & (!g1831) & (!g1832)) + ((!g964) & (!g1157) & (!g1163) & (g1329) & (!g1831) & (g1832)) + ((!g964) & (!g1157) & (g1163) & (!g1329) & (!g1831) & (g1832)) + ((!g964) & (!g1157) & (g1163) & (!g1329) & (g1831) & (g1832)) + ((!g964) & (!g1157) & (g1163) & (g1329) & (!g1831) & (g1832)) + ((!g964) & (!g1157) & (g1163) & (g1329) & (g1831) & (g1832)) + ((!g964) & (g1157) & (!g1163) & (!g1329) & (!g1831) & (!g1832)) + ((!g964) & (g1157) & (!g1163) & (!g1329) & (!g1831) & (g1832)) + ((!g964) & (g1157) & (!g1163) & (g1329) & (g1831) & (!g1832)) + ((!g964) & (g1157) & (!g1163) & (g1329) & (g1831) & (g1832)) + ((!g964) & (g1157) & (g1163) & (!g1329) & (!g1831) & (!g1832)) + ((!g964) & (g1157) & (g1163) & (!g1329) & (g1831) & (!g1832)) + ((!g964) & (g1157) & (g1163) & (g1329) & (!g1831) & (!g1832)) + ((!g964) & (g1157) & (g1163) & (g1329) & (g1831) & (!g1832)) + ((g964) & (!g1157) & (!g1163) & (!g1329) & (!g1831) & (!g1832)) + ((g964) & (!g1157) & (!g1163) & (!g1329) & (!g1831) & (g1832)) + ((g964) & (!g1157) & (!g1163) & (g1329) & (g1831) & (!g1832)) + ((g964) & (!g1157) & (!g1163) & (g1329) & (g1831) & (g1832)) + ((g964) & (!g1157) & (g1163) & (!g1329) & (!g1831) & (g1832)) + ((g964) & (!g1157) & (g1163) & (!g1329) & (g1831) & (g1832)) + ((g964) & (!g1157) & (g1163) & (g1329) & (!g1831) & (g1832)) + ((g964) & (!g1157) & (g1163) & (g1329) & (g1831) & (g1832)) + ((g964) & (g1157) & (!g1163) & (!g1329) & (g1831) & (!g1832)) + ((g964) & (g1157) & (!g1163) & (!g1329) & (g1831) & (g1832)) + ((g964) & (g1157) & (!g1163) & (g1329) & (!g1831) & (!g1832)) + ((g964) & (g1157) & (!g1163) & (g1329) & (!g1831) & (g1832)) + ((g964) & (g1157) & (g1163) & (!g1329) & (!g1831) & (!g1832)) + ((g964) & (g1157) & (g1163) & (!g1329) & (g1831) & (!g1832)) + ((g964) & (g1157) & (g1163) & (g1329) & (!g1831) & (!g1832)) + ((g964) & (g1157) & (g1163) & (g1329) & (g1831) & (!g1832)));
	assign g1834 = (((!ld) & (!g1438) & (!sk[27]) & (g1440) & (!keyx120x)) + ((!ld) & (!g1438) & (!sk[27]) & (g1440) & (keyx120x)) + ((!ld) & (!g1438) & (sk[27]) & (g1440) & (!keyx120x)) + ((!ld) & (!g1438) & (sk[27]) & (g1440) & (keyx120x)) + ((!ld) & (g1438) & (!sk[27]) & (!g1440) & (!keyx120x)) + ((!ld) & (g1438) & (!sk[27]) & (!g1440) & (keyx120x)) + ((!ld) & (g1438) & (!sk[27]) & (g1440) & (!keyx120x)) + ((!ld) & (g1438) & (!sk[27]) & (g1440) & (keyx120x)) + ((!ld) & (g1438) & (sk[27]) & (!g1440) & (!keyx120x)) + ((!ld) & (g1438) & (sk[27]) & (!g1440) & (keyx120x)) + ((ld) & (!g1438) & (!sk[27]) & (g1440) & (!keyx120x)) + ((ld) & (!g1438) & (!sk[27]) & (g1440) & (keyx120x)) + ((ld) & (!g1438) & (sk[27]) & (!g1440) & (keyx120x)) + ((ld) & (!g1438) & (sk[27]) & (g1440) & (keyx120x)) + ((ld) & (g1438) & (!sk[27]) & (!g1440) & (!keyx120x)) + ((ld) & (g1438) & (!sk[27]) & (!g1440) & (keyx120x)) + ((ld) & (g1438) & (!sk[27]) & (g1440) & (!keyx120x)) + ((ld) & (g1438) & (!sk[27]) & (g1440) & (keyx120x)) + ((ld) & (g1438) & (sk[27]) & (!g1440) & (keyx120x)) + ((ld) & (g1438) & (sk[27]) & (g1440) & (keyx120x)));
	assign g1835 = (((!ld) & (!g1447) & (!sk[28]) & (g1449) & (!keyx121x)) + ((!ld) & (!g1447) & (!sk[28]) & (g1449) & (keyx121x)) + ((!ld) & (!g1447) & (sk[28]) & (g1449) & (!keyx121x)) + ((!ld) & (!g1447) & (sk[28]) & (g1449) & (keyx121x)) + ((!ld) & (g1447) & (!sk[28]) & (!g1449) & (!keyx121x)) + ((!ld) & (g1447) & (!sk[28]) & (!g1449) & (keyx121x)) + ((!ld) & (g1447) & (!sk[28]) & (g1449) & (!keyx121x)) + ((!ld) & (g1447) & (!sk[28]) & (g1449) & (keyx121x)) + ((!ld) & (g1447) & (sk[28]) & (!g1449) & (!keyx121x)) + ((!ld) & (g1447) & (sk[28]) & (!g1449) & (keyx121x)) + ((ld) & (!g1447) & (!sk[28]) & (g1449) & (!keyx121x)) + ((ld) & (!g1447) & (!sk[28]) & (g1449) & (keyx121x)) + ((ld) & (!g1447) & (sk[28]) & (!g1449) & (keyx121x)) + ((ld) & (!g1447) & (sk[28]) & (g1449) & (keyx121x)) + ((ld) & (g1447) & (!sk[28]) & (!g1449) & (!keyx121x)) + ((ld) & (g1447) & (!sk[28]) & (!g1449) & (keyx121x)) + ((ld) & (g1447) & (!sk[28]) & (g1449) & (!keyx121x)) + ((ld) & (g1447) & (!sk[28]) & (g1449) & (keyx121x)) + ((ld) & (g1447) & (sk[28]) & (!g1449) & (keyx121x)) + ((ld) & (g1447) & (sk[28]) & (g1449) & (keyx121x)));
	assign g1836 = (((!ld) & (!sk[29]) & (!g1456) & (g1458) & (!keyx122x)) + ((!ld) & (!sk[29]) & (!g1456) & (g1458) & (keyx122x)) + ((!ld) & (!sk[29]) & (g1456) & (!g1458) & (!keyx122x)) + ((!ld) & (!sk[29]) & (g1456) & (!g1458) & (keyx122x)) + ((!ld) & (!sk[29]) & (g1456) & (g1458) & (!keyx122x)) + ((!ld) & (!sk[29]) & (g1456) & (g1458) & (keyx122x)) + ((!ld) & (sk[29]) & (!g1456) & (g1458) & (!keyx122x)) + ((!ld) & (sk[29]) & (!g1456) & (g1458) & (keyx122x)) + ((!ld) & (sk[29]) & (g1456) & (!g1458) & (!keyx122x)) + ((!ld) & (sk[29]) & (g1456) & (!g1458) & (keyx122x)) + ((ld) & (!sk[29]) & (!g1456) & (g1458) & (!keyx122x)) + ((ld) & (!sk[29]) & (!g1456) & (g1458) & (keyx122x)) + ((ld) & (!sk[29]) & (g1456) & (!g1458) & (!keyx122x)) + ((ld) & (!sk[29]) & (g1456) & (!g1458) & (keyx122x)) + ((ld) & (!sk[29]) & (g1456) & (g1458) & (!keyx122x)) + ((ld) & (!sk[29]) & (g1456) & (g1458) & (keyx122x)) + ((ld) & (sk[29]) & (!g1456) & (!g1458) & (keyx122x)) + ((ld) & (sk[29]) & (!g1456) & (g1458) & (keyx122x)) + ((ld) & (sk[29]) & (g1456) & (!g1458) & (keyx122x)) + ((ld) & (sk[29]) & (g1456) & (g1458) & (keyx122x)));
	assign g1837 = (((!sk[30]) & (!ld) & (!g1465) & (g1467) & (!keyx123x)) + ((!sk[30]) & (!ld) & (!g1465) & (g1467) & (keyx123x)) + ((!sk[30]) & (!ld) & (g1465) & (!g1467) & (!keyx123x)) + ((!sk[30]) & (!ld) & (g1465) & (!g1467) & (keyx123x)) + ((!sk[30]) & (!ld) & (g1465) & (g1467) & (!keyx123x)) + ((!sk[30]) & (!ld) & (g1465) & (g1467) & (keyx123x)) + ((!sk[30]) & (ld) & (!g1465) & (g1467) & (!keyx123x)) + ((!sk[30]) & (ld) & (!g1465) & (g1467) & (keyx123x)) + ((!sk[30]) & (ld) & (g1465) & (!g1467) & (!keyx123x)) + ((!sk[30]) & (ld) & (g1465) & (!g1467) & (keyx123x)) + ((!sk[30]) & (ld) & (g1465) & (g1467) & (!keyx123x)) + ((!sk[30]) & (ld) & (g1465) & (g1467) & (keyx123x)) + ((sk[30]) & (!ld) & (!g1465) & (g1467) & (!keyx123x)) + ((sk[30]) & (!ld) & (!g1465) & (g1467) & (keyx123x)) + ((sk[30]) & (!ld) & (g1465) & (!g1467) & (!keyx123x)) + ((sk[30]) & (!ld) & (g1465) & (!g1467) & (keyx123x)) + ((sk[30]) & (ld) & (!g1465) & (!g1467) & (keyx123x)) + ((sk[30]) & (ld) & (!g1465) & (g1467) & (keyx123x)) + ((sk[30]) & (ld) & (g1465) & (!g1467) & (keyx123x)) + ((sk[30]) & (ld) & (g1465) & (g1467) & (keyx123x)));
	assign g1838 = (((!ld) & (!g1474) & (!sk[31]) & (g1476) & (!keyx124x)) + ((!ld) & (!g1474) & (!sk[31]) & (g1476) & (keyx124x)) + ((!ld) & (!g1474) & (sk[31]) & (g1476) & (!keyx124x)) + ((!ld) & (!g1474) & (sk[31]) & (g1476) & (keyx124x)) + ((!ld) & (g1474) & (!sk[31]) & (!g1476) & (!keyx124x)) + ((!ld) & (g1474) & (!sk[31]) & (!g1476) & (keyx124x)) + ((!ld) & (g1474) & (!sk[31]) & (g1476) & (!keyx124x)) + ((!ld) & (g1474) & (!sk[31]) & (g1476) & (keyx124x)) + ((!ld) & (g1474) & (sk[31]) & (!g1476) & (!keyx124x)) + ((!ld) & (g1474) & (sk[31]) & (!g1476) & (keyx124x)) + ((ld) & (!g1474) & (!sk[31]) & (g1476) & (!keyx124x)) + ((ld) & (!g1474) & (!sk[31]) & (g1476) & (keyx124x)) + ((ld) & (!g1474) & (sk[31]) & (!g1476) & (keyx124x)) + ((ld) & (!g1474) & (sk[31]) & (g1476) & (keyx124x)) + ((ld) & (g1474) & (!sk[31]) & (!g1476) & (!keyx124x)) + ((ld) & (g1474) & (!sk[31]) & (!g1476) & (keyx124x)) + ((ld) & (g1474) & (!sk[31]) & (g1476) & (!keyx124x)) + ((ld) & (g1474) & (!sk[31]) & (g1476) & (keyx124x)) + ((ld) & (g1474) & (sk[31]) & (!g1476) & (keyx124x)) + ((ld) & (g1474) & (sk[31]) & (g1476) & (keyx124x)));
	assign g1839 = (((!ld) & (!g1483) & (g1485) & (!sk[32]) & (!keyx125x)) + ((!ld) & (!g1483) & (g1485) & (!sk[32]) & (keyx125x)) + ((!ld) & (!g1483) & (g1485) & (sk[32]) & (!keyx125x)) + ((!ld) & (!g1483) & (g1485) & (sk[32]) & (keyx125x)) + ((!ld) & (g1483) & (!g1485) & (!sk[32]) & (!keyx125x)) + ((!ld) & (g1483) & (!g1485) & (!sk[32]) & (keyx125x)) + ((!ld) & (g1483) & (!g1485) & (sk[32]) & (!keyx125x)) + ((!ld) & (g1483) & (!g1485) & (sk[32]) & (keyx125x)) + ((!ld) & (g1483) & (g1485) & (!sk[32]) & (!keyx125x)) + ((!ld) & (g1483) & (g1485) & (!sk[32]) & (keyx125x)) + ((ld) & (!g1483) & (!g1485) & (sk[32]) & (keyx125x)) + ((ld) & (!g1483) & (g1485) & (!sk[32]) & (!keyx125x)) + ((ld) & (!g1483) & (g1485) & (!sk[32]) & (keyx125x)) + ((ld) & (!g1483) & (g1485) & (sk[32]) & (keyx125x)) + ((ld) & (g1483) & (!g1485) & (!sk[32]) & (!keyx125x)) + ((ld) & (g1483) & (!g1485) & (!sk[32]) & (keyx125x)) + ((ld) & (g1483) & (!g1485) & (sk[32]) & (keyx125x)) + ((ld) & (g1483) & (g1485) & (!sk[32]) & (!keyx125x)) + ((ld) & (g1483) & (g1485) & (!sk[32]) & (keyx125x)) + ((ld) & (g1483) & (g1485) & (sk[32]) & (keyx125x)));
	assign g1840 = (((!ld) & (!g1492) & (!sk[33]) & (g1494) & (!keyx126x)) + ((!ld) & (!g1492) & (!sk[33]) & (g1494) & (keyx126x)) + ((!ld) & (!g1492) & (sk[33]) & (g1494) & (!keyx126x)) + ((!ld) & (!g1492) & (sk[33]) & (g1494) & (keyx126x)) + ((!ld) & (g1492) & (!sk[33]) & (!g1494) & (!keyx126x)) + ((!ld) & (g1492) & (!sk[33]) & (!g1494) & (keyx126x)) + ((!ld) & (g1492) & (!sk[33]) & (g1494) & (!keyx126x)) + ((!ld) & (g1492) & (!sk[33]) & (g1494) & (keyx126x)) + ((!ld) & (g1492) & (sk[33]) & (!g1494) & (!keyx126x)) + ((!ld) & (g1492) & (sk[33]) & (!g1494) & (keyx126x)) + ((ld) & (!g1492) & (!sk[33]) & (g1494) & (!keyx126x)) + ((ld) & (!g1492) & (!sk[33]) & (g1494) & (keyx126x)) + ((ld) & (!g1492) & (sk[33]) & (!g1494) & (keyx126x)) + ((ld) & (!g1492) & (sk[33]) & (g1494) & (keyx126x)) + ((ld) & (g1492) & (!sk[33]) & (!g1494) & (!keyx126x)) + ((ld) & (g1492) & (!sk[33]) & (!g1494) & (keyx126x)) + ((ld) & (g1492) & (!sk[33]) & (g1494) & (!keyx126x)) + ((ld) & (g1492) & (!sk[33]) & (g1494) & (keyx126x)) + ((ld) & (g1492) & (sk[33]) & (!g1494) & (keyx126x)) + ((ld) & (g1492) & (sk[33]) & (g1494) & (keyx126x)));
	assign g1841 = (((!sk[34]) & (!ld) & (!g1501) & (g1503) & (!keyx127x)) + ((!sk[34]) & (!ld) & (!g1501) & (g1503) & (keyx127x)) + ((!sk[34]) & (!ld) & (g1501) & (!g1503) & (!keyx127x)) + ((!sk[34]) & (!ld) & (g1501) & (!g1503) & (keyx127x)) + ((!sk[34]) & (!ld) & (g1501) & (g1503) & (!keyx127x)) + ((!sk[34]) & (!ld) & (g1501) & (g1503) & (keyx127x)) + ((!sk[34]) & (ld) & (!g1501) & (g1503) & (!keyx127x)) + ((!sk[34]) & (ld) & (!g1501) & (g1503) & (keyx127x)) + ((!sk[34]) & (ld) & (g1501) & (!g1503) & (!keyx127x)) + ((!sk[34]) & (ld) & (g1501) & (!g1503) & (keyx127x)) + ((!sk[34]) & (ld) & (g1501) & (g1503) & (!keyx127x)) + ((!sk[34]) & (ld) & (g1501) & (g1503) & (keyx127x)) + ((sk[34]) & (!ld) & (!g1501) & (g1503) & (!keyx127x)) + ((sk[34]) & (!ld) & (!g1501) & (g1503) & (keyx127x)) + ((sk[34]) & (!ld) & (g1501) & (!g1503) & (!keyx127x)) + ((sk[34]) & (!ld) & (g1501) & (!g1503) & (keyx127x)) + ((sk[34]) & (ld) & (!g1501) & (!g1503) & (keyx127x)) + ((sk[34]) & (ld) & (!g1501) & (g1503) & (keyx127x)) + ((sk[34]) & (ld) & (g1501) & (!g1503) & (keyx127x)) + ((sk[34]) & (ld) & (g1501) & (g1503) & (keyx127x)));
	assign g1845 = (((!ld) & (!g1842) & (!sk[35]) & (g1843) & (!g1844)) + ((!ld) & (!g1842) & (!sk[35]) & (g1843) & (g1844)) + ((!ld) & (g1842) & (!sk[35]) & (!g1843) & (!g1844)) + ((!ld) & (g1842) & (!sk[35]) & (!g1843) & (g1844)) + ((!ld) & (g1842) & (!sk[35]) & (g1843) & (!g1844)) + ((!ld) & (g1842) & (!sk[35]) & (g1843) & (g1844)) + ((!ld) & (g1842) & (sk[35]) & (g1843) & (g1844)) + ((ld) & (!g1842) & (!sk[35]) & (g1843) & (!g1844)) + ((ld) & (!g1842) & (!sk[35]) & (g1843) & (g1844)) + ((ld) & (!g1842) & (sk[35]) & (!g1843) & (!g1844)) + ((ld) & (!g1842) & (sk[35]) & (!g1843) & (g1844)) + ((ld) & (!g1842) & (sk[35]) & (g1843) & (!g1844)) + ((ld) & (!g1842) & (sk[35]) & (g1843) & (g1844)) + ((ld) & (g1842) & (!sk[35]) & (!g1843) & (!g1844)) + ((ld) & (g1842) & (!sk[35]) & (!g1843) & (g1844)) + ((ld) & (g1842) & (!sk[35]) & (g1843) & (!g1844)) + ((ld) & (g1842) & (!sk[35]) & (g1843) & (g1844)) + ((ld) & (g1842) & (sk[35]) & (!g1843) & (!g1844)) + ((ld) & (g1842) & (sk[35]) & (!g1843) & (g1844)) + ((ld) & (g1842) & (sk[35]) & (g1843) & (!g1844)) + ((ld) & (g1842) & (sk[35]) & (g1843) & (g1844)));
	assign g1847 = (((!ld) & (!sk[36]) & (g1842) & (!g1843) & (!g1844) & (!g1846)) + ((!ld) & (!sk[36]) & (g1842) & (!g1843) & (!g1844) & (g1846)) + ((!ld) & (!sk[36]) & (g1842) & (!g1843) & (g1844) & (!g1846)) + ((!ld) & (!sk[36]) & (g1842) & (!g1843) & (g1844) & (g1846)) + ((!ld) & (!sk[36]) & (g1842) & (g1843) & (!g1844) & (!g1846)) + ((!ld) & (!sk[36]) & (g1842) & (g1843) & (!g1844) & (g1846)) + ((!ld) & (!sk[36]) & (g1842) & (g1843) & (g1844) & (!g1846)) + ((!ld) & (!sk[36]) & (g1842) & (g1843) & (g1844) & (g1846)) + ((!ld) & (sk[36]) & (g1842) & (!g1843) & (g1844) & (!g1846)) + ((ld) & (!sk[36]) & (!g1842) & (!g1843) & (!g1844) & (!g1846)) + ((ld) & (!sk[36]) & (!g1842) & (!g1843) & (!g1844) & (g1846)) + ((ld) & (!sk[36]) & (!g1842) & (!g1843) & (g1844) & (!g1846)) + ((ld) & (!sk[36]) & (!g1842) & (!g1843) & (g1844) & (g1846)) + ((ld) & (!sk[36]) & (!g1842) & (g1843) & (!g1844) & (!g1846)) + ((ld) & (!sk[36]) & (!g1842) & (g1843) & (!g1844) & (g1846)) + ((ld) & (!sk[36]) & (!g1842) & (g1843) & (g1844) & (!g1846)) + ((ld) & (!sk[36]) & (!g1842) & (g1843) & (g1844) & (g1846)) + ((ld) & (!sk[36]) & (g1842) & (!g1843) & (!g1844) & (!g1846)) + ((ld) & (!sk[36]) & (g1842) & (!g1843) & (!g1844) & (g1846)) + ((ld) & (!sk[36]) & (g1842) & (!g1843) & (g1844) & (!g1846)) + ((ld) & (!sk[36]) & (g1842) & (!g1843) & (g1844) & (g1846)) + ((ld) & (!sk[36]) & (g1842) & (g1843) & (!g1844) & (!g1846)) + ((ld) & (!sk[36]) & (g1842) & (g1843) & (!g1844) & (g1846)) + ((ld) & (!sk[36]) & (g1842) & (g1843) & (g1844) & (!g1846)) + ((ld) & (!sk[36]) & (g1842) & (g1843) & (g1844) & (g1846)));
	assign g1848 = (((!ld) & (!g1842) & (sk[37]) & (g1843) & (g1844) & (!g1846)) + ((!ld) & (g1842) & (!sk[37]) & (!g1843) & (!g1844) & (!g1846)) + ((!ld) & (g1842) & (!sk[37]) & (!g1843) & (!g1844) & (g1846)) + ((!ld) & (g1842) & (!sk[37]) & (!g1843) & (g1844) & (!g1846)) + ((!ld) & (g1842) & (!sk[37]) & (!g1843) & (g1844) & (g1846)) + ((!ld) & (g1842) & (!sk[37]) & (g1843) & (!g1844) & (!g1846)) + ((!ld) & (g1842) & (!sk[37]) & (g1843) & (!g1844) & (g1846)) + ((!ld) & (g1842) & (!sk[37]) & (g1843) & (g1844) & (!g1846)) + ((!ld) & (g1842) & (!sk[37]) & (g1843) & (g1844) & (g1846)) + ((ld) & (!g1842) & (!sk[37]) & (!g1843) & (!g1844) & (!g1846)) + ((ld) & (!g1842) & (!sk[37]) & (!g1843) & (!g1844) & (g1846)) + ((ld) & (!g1842) & (!sk[37]) & (!g1843) & (g1844) & (!g1846)) + ((ld) & (!g1842) & (!sk[37]) & (!g1843) & (g1844) & (g1846)) + ((ld) & (!g1842) & (!sk[37]) & (g1843) & (!g1844) & (!g1846)) + ((ld) & (!g1842) & (!sk[37]) & (g1843) & (!g1844) & (g1846)) + ((ld) & (!g1842) & (!sk[37]) & (g1843) & (g1844) & (!g1846)) + ((ld) & (!g1842) & (!sk[37]) & (g1843) & (g1844) & (g1846)) + ((ld) & (g1842) & (!sk[37]) & (!g1843) & (!g1844) & (!g1846)) + ((ld) & (g1842) & (!sk[37]) & (!g1843) & (!g1844) & (g1846)) + ((ld) & (g1842) & (!sk[37]) & (!g1843) & (g1844) & (!g1846)) + ((ld) & (g1842) & (!sk[37]) & (!g1843) & (g1844) & (g1846)) + ((ld) & (g1842) & (!sk[37]) & (g1843) & (!g1844) & (!g1846)) + ((ld) & (g1842) & (!sk[37]) & (g1843) & (!g1844) & (g1846)) + ((ld) & (g1842) & (!sk[37]) & (g1843) & (g1844) & (!g1846)) + ((ld) & (g1842) & (!sk[37]) & (g1843) & (g1844) & (g1846)));
	assign g1849 = (((!sk[38]) & (!ld) & (g1842)) + ((!sk[38]) & (ld) & (g1842)) + ((sk[38]) & (!ld) & (!g1842)));
	assign g1850 = (((!sk[39]) & (!ld) & (g1842) & (!g1843)) + ((!sk[39]) & (!ld) & (g1842) & (g1843)) + ((!sk[39]) & (ld) & (!g1842) & (g1843)) + ((!sk[39]) & (ld) & (g1842) & (!g1843)) + ((!sk[39]) & (ld) & (g1842) & (g1843)) + ((sk[39]) & (!ld) & (!g1842) & (g1843)) + ((sk[39]) & (!ld) & (g1842) & (!g1843)));
	assign g1851 = (((!ld) & (!g1842) & (!g1843) & (sk[40]) & (g1844)) + ((!ld) & (!g1842) & (g1843) & (!sk[40]) & (!g1844)) + ((!ld) & (!g1842) & (g1843) & (!sk[40]) & (g1844)) + ((!ld) & (!g1842) & (g1843) & (sk[40]) & (g1844)) + ((!ld) & (g1842) & (!g1843) & (!sk[40]) & (!g1844)) + ((!ld) & (g1842) & (!g1843) & (!sk[40]) & (g1844)) + ((!ld) & (g1842) & (!g1843) & (sk[40]) & (g1844)) + ((!ld) & (g1842) & (g1843) & (!sk[40]) & (!g1844)) + ((!ld) & (g1842) & (g1843) & (!sk[40]) & (g1844)) + ((!ld) & (g1842) & (g1843) & (sk[40]) & (!g1844)) + ((ld) & (!g1842) & (g1843) & (!sk[40]) & (!g1844)) + ((ld) & (!g1842) & (g1843) & (!sk[40]) & (g1844)) + ((ld) & (g1842) & (!g1843) & (!sk[40]) & (!g1844)) + ((ld) & (g1842) & (!g1843) & (!sk[40]) & (g1844)) + ((ld) & (g1842) & (g1843) & (!sk[40]) & (!g1844)) + ((ld) & (g1842) & (g1843) & (!sk[40]) & (g1844)));
	assign g1852 = (((!ld) & (!sk[41]) & (g1842) & (!g1843) & (!g1844) & (!g1846)) + ((!ld) & (!sk[41]) & (g1842) & (!g1843) & (!g1844) & (g1846)) + ((!ld) & (!sk[41]) & (g1842) & (!g1843) & (g1844) & (!g1846)) + ((!ld) & (!sk[41]) & (g1842) & (!g1843) & (g1844) & (g1846)) + ((!ld) & (!sk[41]) & (g1842) & (g1843) & (!g1844) & (!g1846)) + ((!ld) & (!sk[41]) & (g1842) & (g1843) & (!g1844) & (g1846)) + ((!ld) & (!sk[41]) & (g1842) & (g1843) & (g1844) & (!g1846)) + ((!ld) & (!sk[41]) & (g1842) & (g1843) & (g1844) & (g1846)) + ((!ld) & (sk[41]) & (!g1842) & (!g1843) & (!g1844) & (g1846)) + ((!ld) & (sk[41]) & (!g1842) & (!g1843) & (g1844) & (g1846)) + ((!ld) & (sk[41]) & (!g1842) & (g1843) & (!g1844) & (g1846)) + ((!ld) & (sk[41]) & (!g1842) & (g1843) & (g1844) & (g1846)) + ((!ld) & (sk[41]) & (g1842) & (!g1843) & (!g1844) & (g1846)) + ((!ld) & (sk[41]) & (g1842) & (!g1843) & (g1844) & (g1846)) + ((!ld) & (sk[41]) & (g1842) & (g1843) & (!g1844) & (g1846)) + ((!ld) & (sk[41]) & (g1842) & (g1843) & (g1844) & (!g1846)) + ((ld) & (!sk[41]) & (!g1842) & (!g1843) & (!g1844) & (!g1846)) + ((ld) & (!sk[41]) & (!g1842) & (!g1843) & (!g1844) & (g1846)) + ((ld) & (!sk[41]) & (!g1842) & (!g1843) & (g1844) & (!g1846)) + ((ld) & (!sk[41]) & (!g1842) & (!g1843) & (g1844) & (g1846)) + ((ld) & (!sk[41]) & (!g1842) & (g1843) & (!g1844) & (!g1846)) + ((ld) & (!sk[41]) & (!g1842) & (g1843) & (!g1844) & (g1846)) + ((ld) & (!sk[41]) & (!g1842) & (g1843) & (g1844) & (!g1846)) + ((ld) & (!sk[41]) & (!g1842) & (g1843) & (g1844) & (g1846)) + ((ld) & (!sk[41]) & (g1842) & (!g1843) & (!g1844) & (!g1846)) + ((ld) & (!sk[41]) & (g1842) & (!g1843) & (!g1844) & (g1846)) + ((ld) & (!sk[41]) & (g1842) & (!g1843) & (g1844) & (!g1846)) + ((ld) & (!sk[41]) & (g1842) & (!g1843) & (g1844) & (g1846)) + ((ld) & (!sk[41]) & (g1842) & (g1843) & (!g1844) & (!g1846)) + ((ld) & (!sk[41]) & (g1842) & (g1843) & (!g1844) & (g1846)) + ((ld) & (!sk[41]) & (g1842) & (g1843) & (g1844) & (!g1846)) + ((ld) & (!sk[41]) & (g1842) & (g1843) & (g1844) & (g1846)));
	assign g1853 = (((!g1846) & (g1844) & (!g1843) & (!sk[42]) & (!g1842) & (!ld)) + ((!g1846) & (g1844) & (!g1843) & (!sk[42]) & (!g1842) & (ld)) + ((!g1846) & (g1844) & (!g1843) & (!sk[42]) & (g1842) & (!ld)) + ((!g1846) & (g1844) & (!g1843) & (!sk[42]) & (g1842) & (ld)) + ((!g1846) & (g1844) & (!g1843) & (sk[42]) & (!g1842) & (!ld)) + ((!g1846) & (g1844) & (g1843) & (!sk[42]) & (!g1842) & (!ld)) + ((!g1846) & (g1844) & (g1843) & (!sk[42]) & (!g1842) & (ld)) + ((!g1846) & (g1844) & (g1843) & (!sk[42]) & (g1842) & (!ld)) + ((!g1846) & (g1844) & (g1843) & (!sk[42]) & (g1842) & (ld)) + ((g1846) & (!g1844) & (!g1843) & (!sk[42]) & (!g1842) & (!ld)) + ((g1846) & (!g1844) & (!g1843) & (!sk[42]) & (!g1842) & (ld)) + ((g1846) & (!g1844) & (!g1843) & (!sk[42]) & (g1842) & (!ld)) + ((g1846) & (!g1844) & (!g1843) & (!sk[42]) & (g1842) & (ld)) + ((g1846) & (!g1844) & (!g1843) & (sk[42]) & (!g1842) & (!ld)) + ((g1846) & (!g1844) & (g1843) & (!sk[42]) & (!g1842) & (!ld)) + ((g1846) & (!g1844) & (g1843) & (!sk[42]) & (!g1842) & (ld)) + ((g1846) & (!g1844) & (g1843) & (!sk[42]) & (g1842) & (!ld)) + ((g1846) & (!g1844) & (g1843) & (!sk[42]) & (g1842) & (ld)) + ((g1846) & (g1844) & (!g1843) & (!sk[42]) & (!g1842) & (!ld)) + ((g1846) & (g1844) & (!g1843) & (!sk[42]) & (!g1842) & (ld)) + ((g1846) & (g1844) & (!g1843) & (!sk[42]) & (g1842) & (!ld)) + ((g1846) & (g1844) & (!g1843) & (!sk[42]) & (g1842) & (ld)) + ((g1846) & (g1844) & (g1843) & (!sk[42]) & (!g1842) & (!ld)) + ((g1846) & (g1844) & (g1843) & (!sk[42]) & (!g1842) & (ld)) + ((g1846) & (g1844) & (g1843) & (!sk[42]) & (g1842) & (!ld)) + ((g1846) & (g1844) & (g1843) & (!sk[42]) & (g1842) & (ld)));
	assign g1854 = (((!g1846) & (!g1844) & (g1843) & (g1842) & (sk[43]) & (!ld)) + ((!g1846) & (g1844) & (!g1843) & (!g1842) & (!sk[43]) & (!ld)) + ((!g1846) & (g1844) & (!g1843) & (!g1842) & (!sk[43]) & (ld)) + ((!g1846) & (g1844) & (!g1843) & (g1842) & (!sk[43]) & (!ld)) + ((!g1846) & (g1844) & (!g1843) & (g1842) & (!sk[43]) & (ld)) + ((!g1846) & (g1844) & (g1843) & (!g1842) & (!sk[43]) & (!ld)) + ((!g1846) & (g1844) & (g1843) & (!g1842) & (!sk[43]) & (ld)) + ((!g1846) & (g1844) & (g1843) & (g1842) & (!sk[43]) & (!ld)) + ((!g1846) & (g1844) & (g1843) & (g1842) & (!sk[43]) & (ld)) + ((!g1846) & (g1844) & (g1843) & (g1842) & (sk[43]) & (!ld)) + ((g1846) & (!g1844) & (!g1843) & (!g1842) & (!sk[43]) & (!ld)) + ((g1846) & (!g1844) & (!g1843) & (!g1842) & (!sk[43]) & (ld)) + ((g1846) & (!g1844) & (!g1843) & (!g1842) & (sk[43]) & (!ld)) + ((g1846) & (!g1844) & (!g1843) & (g1842) & (!sk[43]) & (!ld)) + ((g1846) & (!g1844) & (!g1843) & (g1842) & (!sk[43]) & (ld)) + ((g1846) & (!g1844) & (g1843) & (!g1842) & (!sk[43]) & (!ld)) + ((g1846) & (!g1844) & (g1843) & (!g1842) & (!sk[43]) & (ld)) + ((g1846) & (!g1844) & (g1843) & (g1842) & (!sk[43]) & (!ld)) + ((g1846) & (!g1844) & (g1843) & (g1842) & (!sk[43]) & (ld)) + ((g1846) & (g1844) & (!g1843) & (!g1842) & (!sk[43]) & (!ld)) + ((g1846) & (g1844) & (!g1843) & (!g1842) & (!sk[43]) & (ld)) + ((g1846) & (g1844) & (!g1843) & (g1842) & (!sk[43]) & (!ld)) + ((g1846) & (g1844) & (!g1843) & (g1842) & (!sk[43]) & (ld)) + ((g1846) & (g1844) & (g1843) & (!g1842) & (!sk[43]) & (!ld)) + ((g1846) & (g1844) & (g1843) & (!g1842) & (!sk[43]) & (ld)) + ((g1846) & (g1844) & (g1843) & (g1842) & (!sk[43]) & (!ld)) + ((g1846) & (g1844) & (g1843) & (g1842) & (!sk[43]) & (ld)));
	assign g1855 = (((!g1846) & (!g1844) & (g1843) & (!g1842) & (sk[44]) & (!ld)) + ((!g1846) & (g1844) & (!g1843) & (!g1842) & (!sk[44]) & (!ld)) + ((!g1846) & (g1844) & (!g1843) & (!g1842) & (!sk[44]) & (ld)) + ((!g1846) & (g1844) & (!g1843) & (g1842) & (!sk[44]) & (!ld)) + ((!g1846) & (g1844) & (!g1843) & (g1842) & (!sk[44]) & (ld)) + ((!g1846) & (g1844) & (g1843) & (!g1842) & (!sk[44]) & (!ld)) + ((!g1846) & (g1844) & (g1843) & (!g1842) & (!sk[44]) & (ld)) + ((!g1846) & (g1844) & (g1843) & (g1842) & (!sk[44]) & (!ld)) + ((!g1846) & (g1844) & (g1843) & (g1842) & (!sk[44]) & (ld)) + ((!g1846) & (g1844) & (g1843) & (g1842) & (sk[44]) & (!ld)) + ((g1846) & (!g1844) & (!g1843) & (!g1842) & (!sk[44]) & (!ld)) + ((g1846) & (!g1844) & (!g1843) & (!g1842) & (!sk[44]) & (ld)) + ((g1846) & (!g1844) & (!g1843) & (g1842) & (!sk[44]) & (!ld)) + ((g1846) & (!g1844) & (!g1843) & (g1842) & (!sk[44]) & (ld)) + ((g1846) & (!g1844) & (g1843) & (!g1842) & (!sk[44]) & (!ld)) + ((g1846) & (!g1844) & (g1843) & (!g1842) & (!sk[44]) & (ld)) + ((g1846) & (!g1844) & (g1843) & (g1842) & (!sk[44]) & (!ld)) + ((g1846) & (!g1844) & (g1843) & (g1842) & (!sk[44]) & (ld)) + ((g1846) & (g1844) & (!g1843) & (!g1842) & (!sk[44]) & (!ld)) + ((g1846) & (g1844) & (!g1843) & (!g1842) & (!sk[44]) & (ld)) + ((g1846) & (g1844) & (!g1843) & (g1842) & (!sk[44]) & (!ld)) + ((g1846) & (g1844) & (!g1843) & (g1842) & (!sk[44]) & (ld)) + ((g1846) & (g1844) & (g1843) & (!g1842) & (!sk[44]) & (!ld)) + ((g1846) & (g1844) & (g1843) & (!g1842) & (!sk[44]) & (ld)) + ((g1846) & (g1844) & (g1843) & (g1842) & (!sk[44]) & (!ld)) + ((g1846) & (g1844) & (g1843) & (g1842) & (!sk[44]) & (ld)));
	assign g1856 = (((!g1846) & (!g1844) & (sk[45]) & (!g1843) & (g1842) & (!ld)) + ((!g1846) & (g1844) & (!sk[45]) & (!g1843) & (!g1842) & (!ld)) + ((!g1846) & (g1844) & (!sk[45]) & (!g1843) & (!g1842) & (ld)) + ((!g1846) & (g1844) & (!sk[45]) & (!g1843) & (g1842) & (!ld)) + ((!g1846) & (g1844) & (!sk[45]) & (!g1843) & (g1842) & (ld)) + ((!g1846) & (g1844) & (!sk[45]) & (g1843) & (!g1842) & (!ld)) + ((!g1846) & (g1844) & (!sk[45]) & (g1843) & (!g1842) & (ld)) + ((!g1846) & (g1844) & (!sk[45]) & (g1843) & (g1842) & (!ld)) + ((!g1846) & (g1844) & (!sk[45]) & (g1843) & (g1842) & (ld)) + ((g1846) & (!g1844) & (!sk[45]) & (!g1843) & (!g1842) & (!ld)) + ((g1846) & (!g1844) & (!sk[45]) & (!g1843) & (!g1842) & (ld)) + ((g1846) & (!g1844) & (!sk[45]) & (!g1843) & (g1842) & (!ld)) + ((g1846) & (!g1844) & (!sk[45]) & (!g1843) & (g1842) & (ld)) + ((g1846) & (!g1844) & (!sk[45]) & (g1843) & (!g1842) & (!ld)) + ((g1846) & (!g1844) & (!sk[45]) & (g1843) & (!g1842) & (ld)) + ((g1846) & (!g1844) & (!sk[45]) & (g1843) & (g1842) & (!ld)) + ((g1846) & (!g1844) & (!sk[45]) & (g1843) & (g1842) & (ld)) + ((g1846) & (!g1844) & (sk[45]) & (!g1843) & (!g1842) & (!ld)) + ((g1846) & (g1844) & (!sk[45]) & (!g1843) & (!g1842) & (!ld)) + ((g1846) & (g1844) & (!sk[45]) & (!g1843) & (!g1842) & (ld)) + ((g1846) & (g1844) & (!sk[45]) & (!g1843) & (g1842) & (!ld)) + ((g1846) & (g1844) & (!sk[45]) & (!g1843) & (g1842) & (ld)) + ((g1846) & (g1844) & (!sk[45]) & (g1843) & (!g1842) & (!ld)) + ((g1846) & (g1844) & (!sk[45]) & (g1843) & (!g1842) & (ld)) + ((g1846) & (g1844) & (!sk[45]) & (g1843) & (g1842) & (!ld)) + ((g1846) & (g1844) & (!sk[45]) & (g1843) & (g1842) & (ld)));
	assign g1857 = (((!g1846) & (!g1844) & (sk[46]) & (!g1843) & (!g1842) & (!ld)) + ((!g1846) & (g1844) & (!sk[46]) & (!g1843) & (!g1842) & (!ld)) + ((!g1846) & (g1844) & (!sk[46]) & (!g1843) & (!g1842) & (ld)) + ((!g1846) & (g1844) & (!sk[46]) & (!g1843) & (g1842) & (!ld)) + ((!g1846) & (g1844) & (!sk[46]) & (!g1843) & (g1842) & (ld)) + ((!g1846) & (g1844) & (!sk[46]) & (g1843) & (!g1842) & (!ld)) + ((!g1846) & (g1844) & (!sk[46]) & (g1843) & (!g1842) & (ld)) + ((!g1846) & (g1844) & (!sk[46]) & (g1843) & (g1842) & (!ld)) + ((!g1846) & (g1844) & (!sk[46]) & (g1843) & (g1842) & (ld)) + ((!g1846) & (g1844) & (sk[46]) & (g1843) & (g1842) & (!ld)) + ((g1846) & (!g1844) & (!sk[46]) & (!g1843) & (!g1842) & (!ld)) + ((g1846) & (!g1844) & (!sk[46]) & (!g1843) & (!g1842) & (ld)) + ((g1846) & (!g1844) & (!sk[46]) & (!g1843) & (g1842) & (!ld)) + ((g1846) & (!g1844) & (!sk[46]) & (!g1843) & (g1842) & (ld)) + ((g1846) & (!g1844) & (!sk[46]) & (g1843) & (!g1842) & (!ld)) + ((g1846) & (!g1844) & (!sk[46]) & (g1843) & (!g1842) & (ld)) + ((g1846) & (!g1844) & (!sk[46]) & (g1843) & (g1842) & (!ld)) + ((g1846) & (!g1844) & (!sk[46]) & (g1843) & (g1842) & (ld)) + ((g1846) & (!g1844) & (sk[46]) & (!g1843) & (!g1842) & (!ld)) + ((g1846) & (g1844) & (!sk[46]) & (!g1843) & (!g1842) & (!ld)) + ((g1846) & (g1844) & (!sk[46]) & (!g1843) & (!g1842) & (ld)) + ((g1846) & (g1844) & (!sk[46]) & (!g1843) & (g1842) & (!ld)) + ((g1846) & (g1844) & (!sk[46]) & (!g1843) & (g1842) & (ld)) + ((g1846) & (g1844) & (!sk[46]) & (g1843) & (!g1842) & (!ld)) + ((g1846) & (g1844) & (!sk[46]) & (g1843) & (!g1842) & (ld)) + ((g1846) & (g1844) & (!sk[46]) & (g1843) & (g1842) & (!ld)) + ((g1846) & (g1844) & (!sk[46]) & (g1843) & (g1842) & (ld)));
	assign g1858 = (((!sk[47]) & (!g1859) & (g1860)) + ((!sk[47]) & (g1859) & (g1860)) + ((sk[47]) & (!g1859) & (!g1860)));
	assign g1859 = (((!sk[48]) & (!g943) & (g1861)) + ((!sk[48]) & (g943) & (g1861)) + ((sk[48]) & (!g943) & (g1861)));
	assign g1860 = (((!g943) & (!sk[49]) & (g1864)) + ((g943) & (!sk[49]) & (g1864)) + ((g943) & (sk[49]) & (g1864)));
	assign g1861 = (((!sk[50]) & (!g1862) & (g1863)) + ((!sk[50]) & (g1862) & (g1863)) + ((sk[50]) & (!g1862) & (!g1863)));
	assign g1862 = (((!g1163) & (!sk[51]) & (g1867)) + ((!g1163) & (sk[51]) & (g1867)) + ((g1163) & (!sk[51]) & (g1867)));
	assign g1863 = (((!sk[52]) & (!g1163) & (g1868)) + ((!sk[52]) & (g1163) & (g1868)) + ((sk[52]) & (g1163) & (g1868)));
	assign g1864 = (((!sk[53]) & (!g1865) & (g1866)) + ((!sk[53]) & (g1865) & (g1866)) + ((sk[53]) & (!g1865) & (!g1866)));
	assign g1865 = (((!sk[54]) & (!g1163) & (g1869)) + ((!sk[54]) & (g1163) & (g1869)) + ((sk[54]) & (!g1163) & (g1869)));
	assign g1866 = (((!sk[55]) & (!g1163) & (g1870)) + ((!sk[55]) & (g1163) & (g1870)) + ((sk[55]) & (g1163) & (g1870)));
	assign g1867 = (((!sk[56]) & (!g1092) & (!g1064) & (g1635) & (!g1136)) + ((!sk[56]) & (!g1092) & (!g1064) & (g1635) & (g1136)) + ((!sk[56]) & (!g1092) & (g1064) & (!g1635) & (!g1136)) + ((!sk[56]) & (!g1092) & (g1064) & (!g1635) & (g1136)) + ((!sk[56]) & (!g1092) & (g1064) & (g1635) & (!g1136)) + ((!sk[56]) & (!g1092) & (g1064) & (g1635) & (g1136)) + ((!sk[56]) & (g1092) & (!g1064) & (g1635) & (!g1136)) + ((!sk[56]) & (g1092) & (!g1064) & (g1635) & (g1136)) + ((!sk[56]) & (g1092) & (g1064) & (!g1635) & (!g1136)) + ((!sk[56]) & (g1092) & (g1064) & (!g1635) & (g1136)) + ((!sk[56]) & (g1092) & (g1064) & (g1635) & (!g1136)) + ((!sk[56]) & (g1092) & (g1064) & (g1635) & (g1136)) + ((sk[56]) & (!g1092) & (!g1064) & (!g1635) & (g1136)) + ((sk[56]) & (!g1092) & (!g1064) & (g1635) & (!g1136)) + ((sk[56]) & (!g1092) & (g1064) & (!g1635) & (!g1136)) + ((sk[56]) & (!g1092) & (g1064) & (g1635) & (g1136)) + ((sk[56]) & (g1092) & (!g1064) & (!g1635) & (!g1136)) + ((sk[56]) & (g1092) & (!g1064) & (g1635) & (g1136)) + ((sk[56]) & (g1092) & (g1064) & (!g1635) & (g1136)) + ((sk[56]) & (g1092) & (g1064) & (g1635) & (!g1136)));
	assign g1868 = (((!g1830) & (!sk[57]) & (g1136)) + ((!g1830) & (sk[57]) & (g1136)) + ((g1830) & (!sk[57]) & (g1136)) + ((g1830) & (sk[57]) & (!g1136)));
	assign g1869 = (((!g1092) & (!sk[58]) & (!g1064) & (g1635) & (!g1136)) + ((!g1092) & (!sk[58]) & (!g1064) & (g1635) & (g1136)) + ((!g1092) & (!sk[58]) & (g1064) & (!g1635) & (!g1136)) + ((!g1092) & (!sk[58]) & (g1064) & (!g1635) & (g1136)) + ((!g1092) & (!sk[58]) & (g1064) & (g1635) & (!g1136)) + ((!g1092) & (!sk[58]) & (g1064) & (g1635) & (g1136)) + ((!g1092) & (sk[58]) & (!g1064) & (!g1635) & (!g1136)) + ((!g1092) & (sk[58]) & (!g1064) & (g1635) & (g1136)) + ((!g1092) & (sk[58]) & (g1064) & (!g1635) & (g1136)) + ((!g1092) & (sk[58]) & (g1064) & (g1635) & (!g1136)) + ((g1092) & (!sk[58]) & (!g1064) & (g1635) & (!g1136)) + ((g1092) & (!sk[58]) & (!g1064) & (g1635) & (g1136)) + ((g1092) & (!sk[58]) & (g1064) & (!g1635) & (!g1136)) + ((g1092) & (!sk[58]) & (g1064) & (!g1635) & (g1136)) + ((g1092) & (!sk[58]) & (g1064) & (g1635) & (!g1136)) + ((g1092) & (!sk[58]) & (g1064) & (g1635) & (g1136)) + ((g1092) & (sk[58]) & (!g1064) & (!g1635) & (g1136)) + ((g1092) & (sk[58]) & (!g1064) & (g1635) & (!g1136)) + ((g1092) & (sk[58]) & (g1064) & (!g1635) & (!g1136)) + ((g1092) & (sk[58]) & (g1064) & (g1635) & (g1136)));
	assign g1870 = (((!g1830) & (!sk[59]) & (g1136)) + ((!g1830) & (sk[59]) & (g1136)) + ((g1830) & (!sk[59]) & (g1136)) + ((g1830) & (sk[59]) & (!g1136)));
	assign g1871 = (((!sk[60]) & (!g1872) & (g1873)) + ((!sk[60]) & (g1872) & (g1873)) + ((sk[60]) & (!g1872) & (!g1873)));
	assign g1872 = (((!g1064) & (!sk[61]) & (g1874)) + ((!g1064) & (sk[61]) & (g1874)) + ((g1064) & (!sk[61]) & (g1874)));
	assign g1873 = (((!sk[62]) & (!g1064) & (g1877)) + ((!sk[62]) & (g1064) & (g1877)) + ((sk[62]) & (g1064) & (g1877)));
	assign g1874 = (((!sk[63]) & (!g1875) & (g1876)) + ((!sk[63]) & (g1875) & (g1876)) + ((sk[63]) & (!g1875) & (!g1876)));
	assign g1875 = (((!sk[64]) & (!g1163) & (g1880)) + ((!sk[64]) & (g1163) & (g1880)) + ((sk[64]) & (!g1163) & (g1880)));
	assign g1876 = (((!g1163) & (!sk[65]) & (g1881)) + ((g1163) & (!sk[65]) & (g1881)) + ((g1163) & (sk[65]) & (g1881)));
	assign g1877 = (((!g1878) & (!sk[66]) & (g1879)) + ((!g1878) & (sk[66]) & (!g1879)) + ((g1878) & (!sk[66]) & (g1879)));
	assign g1878 = (((!sk[67]) & (!g1163) & (g1882)) + ((!sk[67]) & (g1163) & (g1882)) + ((sk[67]) & (!g1163) & (g1882)));
	assign g1879 = (((!sk[68]) & (!g1163) & (g1883)) + ((!sk[68]) & (g1163) & (g1883)) + ((sk[68]) & (g1163) & (g1883)));
	assign g1880 = (((!g1156) & (!g1121) & (!sk[69]) & (g1340) & (!g1129)) + ((!g1156) & (!g1121) & (!sk[69]) & (g1340) & (g1129)) + ((!g1156) & (!g1121) & (sk[69]) & (!g1340) & (g1129)) + ((!g1156) & (!g1121) & (sk[69]) & (g1340) & (!g1129)) + ((!g1156) & (g1121) & (!sk[69]) & (!g1340) & (!g1129)) + ((!g1156) & (g1121) & (!sk[69]) & (!g1340) & (g1129)) + ((!g1156) & (g1121) & (!sk[69]) & (g1340) & (!g1129)) + ((!g1156) & (g1121) & (!sk[69]) & (g1340) & (g1129)) + ((!g1156) & (g1121) & (sk[69]) & (!g1340) & (!g1129)) + ((!g1156) & (g1121) & (sk[69]) & (g1340) & (g1129)) + ((g1156) & (!g1121) & (!sk[69]) & (g1340) & (!g1129)) + ((g1156) & (!g1121) & (!sk[69]) & (g1340) & (g1129)) + ((g1156) & (!g1121) & (sk[69]) & (!g1340) & (!g1129)) + ((g1156) & (!g1121) & (sk[69]) & (g1340) & (g1129)) + ((g1156) & (g1121) & (!sk[69]) & (!g1340) & (!g1129)) + ((g1156) & (g1121) & (!sk[69]) & (!g1340) & (g1129)) + ((g1156) & (g1121) & (!sk[69]) & (g1340) & (!g1129)) + ((g1156) & (g1121) & (!sk[69]) & (g1340) & (g1129)) + ((g1156) & (g1121) & (sk[69]) & (!g1340) & (g1129)) + ((g1156) & (g1121) & (sk[69]) & (g1340) & (!g1129)));
	assign g1881 = (((!sk[70]) & (!g1825) & (g1129)) + ((!sk[70]) & (g1825) & (g1129)) + ((sk[70]) & (!g1825) & (g1129)) + ((sk[70]) & (g1825) & (!g1129)));
	assign g1882 = (((!g1156) & (!g1121) & (!sk[71]) & (g1340) & (!g1129)) + ((!g1156) & (!g1121) & (!sk[71]) & (g1340) & (g1129)) + ((!g1156) & (!g1121) & (sk[71]) & (!g1340) & (!g1129)) + ((!g1156) & (!g1121) & (sk[71]) & (g1340) & (g1129)) + ((!g1156) & (g1121) & (!sk[71]) & (!g1340) & (!g1129)) + ((!g1156) & (g1121) & (!sk[71]) & (!g1340) & (g1129)) + ((!g1156) & (g1121) & (!sk[71]) & (g1340) & (!g1129)) + ((!g1156) & (g1121) & (!sk[71]) & (g1340) & (g1129)) + ((!g1156) & (g1121) & (sk[71]) & (!g1340) & (g1129)) + ((!g1156) & (g1121) & (sk[71]) & (g1340) & (!g1129)) + ((g1156) & (!g1121) & (!sk[71]) & (g1340) & (!g1129)) + ((g1156) & (!g1121) & (!sk[71]) & (g1340) & (g1129)) + ((g1156) & (!g1121) & (sk[71]) & (!g1340) & (g1129)) + ((g1156) & (!g1121) & (sk[71]) & (g1340) & (!g1129)) + ((g1156) & (g1121) & (!sk[71]) & (!g1340) & (!g1129)) + ((g1156) & (g1121) & (!sk[71]) & (!g1340) & (g1129)) + ((g1156) & (g1121) & (!sk[71]) & (g1340) & (!g1129)) + ((g1156) & (g1121) & (!sk[71]) & (g1340) & (g1129)) + ((g1156) & (g1121) & (sk[71]) & (!g1340) & (!g1129)) + ((g1156) & (g1121) & (sk[71]) & (g1340) & (g1129)));
	assign g1883 = (((!g1825) & (!sk[72]) & (g1129)) + ((!g1825) & (sk[72]) & (g1129)) + ((g1825) & (!sk[72]) & (g1129)) + ((g1825) & (sk[72]) & (!g1129)));
	assign g1884 = (((!g1885) & (!sk[73]) & (g1886)) + ((!g1885) & (sk[73]) & (!g1886)) + ((g1885) & (!sk[73]) & (g1886)));
	assign g1885 = (((!g837) & (!sk[74]) & (g1887)) + ((!g837) & (sk[74]) & (g1887)) + ((g837) & (!sk[74]) & (g1887)));
	assign g1886 = (((!sk[75]) & (!g837) & (g1890)) + ((!sk[75]) & (g837) & (g1890)) + ((sk[75]) & (g837) & (g1890)));
	assign g1887 = (((!g1888) & (!sk[76]) & (g1889)) + ((!g1888) & (sk[76]) & (!g1889)) + ((g1888) & (!sk[76]) & (g1889)));
	assign g1888 = (((!sk[77]) & (!g1163) & (g1893)) + ((!sk[77]) & (g1163) & (g1893)) + ((sk[77]) & (!g1163) & (g1893)));
	assign g1889 = (((!sk[78]) & (!g1163) & (g1809)) + ((!sk[78]) & (g1163) & (g1809)) + ((sk[78]) & (g1163) & (g1809)));
	assign g1890 = (((!g1891) & (!sk[79]) & (g1892)) + ((!g1891) & (sk[79]) & (!g1892)) + ((g1891) & (!sk[79]) & (g1892)));
	assign g1891 = (((!g1163) & (!sk[80]) & (g1894)) + ((!g1163) & (sk[80]) & (g1894)) + ((g1163) & (!sk[80]) & (g1894)));
	assign g1892 = (((!sk[81]) & (!g1163) & (g1809)) + ((!sk[81]) & (g1163) & (g1809)) + ((sk[81]) & (g1163) & (!g1809)));
	assign g1893 = (((!g900) & (!g829) & (!sk[82]) & (g1246) & (!g765)) + ((!g900) & (!g829) & (!sk[82]) & (g1246) & (g765)) + ((!g900) & (!g829) & (sk[82]) & (!g1246) & (g765)) + ((!g900) & (!g829) & (sk[82]) & (g1246) & (!g765)) + ((!g900) & (g829) & (!sk[82]) & (!g1246) & (!g765)) + ((!g900) & (g829) & (!sk[82]) & (!g1246) & (g765)) + ((!g900) & (g829) & (!sk[82]) & (g1246) & (!g765)) + ((!g900) & (g829) & (!sk[82]) & (g1246) & (g765)) + ((!g900) & (g829) & (sk[82]) & (!g1246) & (!g765)) + ((!g900) & (g829) & (sk[82]) & (g1246) & (g765)) + ((g900) & (!g829) & (!sk[82]) & (g1246) & (!g765)) + ((g900) & (!g829) & (!sk[82]) & (g1246) & (g765)) + ((g900) & (!g829) & (sk[82]) & (!g1246) & (!g765)) + ((g900) & (!g829) & (sk[82]) & (g1246) & (g765)) + ((g900) & (g829) & (!sk[82]) & (!g1246) & (!g765)) + ((g900) & (g829) & (!sk[82]) & (!g1246) & (g765)) + ((g900) & (g829) & (!sk[82]) & (g1246) & (!g765)) + ((g900) & (g829) & (!sk[82]) & (g1246) & (g765)) + ((g900) & (g829) & (sk[82]) & (!g1246) & (g765)) + ((g900) & (g829) & (sk[82]) & (g1246) & (!g765)));
	assign g1894 = (((!g900) & (!g829) & (!sk[83]) & (g1246) & (!g765)) + ((!g900) & (!g829) & (!sk[83]) & (g1246) & (g765)) + ((!g900) & (!g829) & (sk[83]) & (!g1246) & (!g765)) + ((!g900) & (!g829) & (sk[83]) & (g1246) & (g765)) + ((!g900) & (g829) & (!sk[83]) & (!g1246) & (!g765)) + ((!g900) & (g829) & (!sk[83]) & (!g1246) & (g765)) + ((!g900) & (g829) & (!sk[83]) & (g1246) & (!g765)) + ((!g900) & (g829) & (!sk[83]) & (g1246) & (g765)) + ((!g900) & (g829) & (sk[83]) & (!g1246) & (g765)) + ((!g900) & (g829) & (sk[83]) & (g1246) & (!g765)) + ((g900) & (!g829) & (!sk[83]) & (g1246) & (!g765)) + ((g900) & (!g829) & (!sk[83]) & (g1246) & (g765)) + ((g900) & (!g829) & (sk[83]) & (!g1246) & (g765)) + ((g900) & (!g829) & (sk[83]) & (g1246) & (!g765)) + ((g900) & (g829) & (!sk[83]) & (!g1246) & (!g765)) + ((g900) & (g829) & (!sk[83]) & (!g1246) & (g765)) + ((g900) & (g829) & (!sk[83]) & (g1246) & (!g765)) + ((g900) & (g829) & (!sk[83]) & (g1246) & (g765)) + ((g900) & (g829) & (sk[83]) & (!g1246) & (!g765)) + ((g900) & (g829) & (sk[83]) & (g1246) & (g765)));
	assign g1895 = (((!sk[84]) & (!g1896) & (g1897)) + ((!sk[84]) & (g1896) & (g1897)) + ((sk[84]) & (!g1896) & (!g1897)));
	assign g1896 = (((!sk[85]) & (!g403) & (g1898)) + ((!sk[85]) & (g403) & (g1898)) + ((sk[85]) & (!g403) & (g1898)));
	assign g1897 = (((!sk[86]) & (!g403) & (g1901)) + ((!sk[86]) & (g403) & (g1901)) + ((sk[86]) & (g403) & (g1901)));
	assign g1898 = (((!g1899) & (!sk[87]) & (g1900)) + ((!g1899) & (sk[87]) & (!g1900)) + ((g1899) & (!sk[87]) & (g1900)));
	assign g1899 = (((!sk[88]) & (!g1163) & (g1904)) + ((!sk[88]) & (g1163) & (g1904)) + ((sk[88]) & (!g1163) & (g1904)));
	assign g1900 = (((!g1163) & (!sk[89]) & (g1905)) + ((g1163) & (!sk[89]) & (g1905)) + ((g1163) & (sk[89]) & (g1905)));
	assign g1901 = (((!g1902) & (!sk[90]) & (g1903)) + ((!g1902) & (sk[90]) & (!g1903)) + ((g1902) & (!sk[90]) & (g1903)));
	assign g1902 = (((!g1163) & (!sk[91]) & (g1906)) + ((!g1163) & (sk[91]) & (g1906)) + ((g1163) & (!sk[91]) & (g1906)));
	assign g1903 = (((!sk[92]) & (!g1163) & (g1907)) + ((!sk[92]) & (g1163) & (g1907)) + ((sk[92]) & (g1163) & (g1907)));
	assign g1904 = (((!sk[93]) & (!g538) & (!g452) & (g1682) & (!g475)) + ((!sk[93]) & (!g538) & (!g452) & (g1682) & (g475)) + ((!sk[93]) & (!g538) & (g452) & (!g1682) & (!g475)) + ((!sk[93]) & (!g538) & (g452) & (!g1682) & (g475)) + ((!sk[93]) & (!g538) & (g452) & (g1682) & (!g475)) + ((!sk[93]) & (!g538) & (g452) & (g1682) & (g475)) + ((!sk[93]) & (g538) & (!g452) & (g1682) & (!g475)) + ((!sk[93]) & (g538) & (!g452) & (g1682) & (g475)) + ((!sk[93]) & (g538) & (g452) & (!g1682) & (!g475)) + ((!sk[93]) & (g538) & (g452) & (!g1682) & (g475)) + ((!sk[93]) & (g538) & (g452) & (g1682) & (!g475)) + ((!sk[93]) & (g538) & (g452) & (g1682) & (g475)) + ((sk[93]) & (!g538) & (!g452) & (!g1682) & (g475)) + ((sk[93]) & (!g538) & (!g452) & (g1682) & (!g475)) + ((sk[93]) & (!g538) & (g452) & (!g1682) & (!g475)) + ((sk[93]) & (!g538) & (g452) & (g1682) & (g475)) + ((sk[93]) & (g538) & (!g452) & (!g1682) & (!g475)) + ((sk[93]) & (g538) & (!g452) & (g1682) & (g475)) + ((sk[93]) & (g538) & (g452) & (!g1682) & (g475)) + ((sk[93]) & (g538) & (g452) & (g1682) & (!g475)));
	assign g1905 = (((!g1768) & (!sk[94]) & (g475)) + ((!g1768) & (sk[94]) & (g475)) + ((g1768) & (!sk[94]) & (g475)) + ((g1768) & (sk[94]) & (!g475)));
	assign g1906 = (((!g538) & (!sk[95]) & (!g452) & (g1682) & (!g475)) + ((!g538) & (!sk[95]) & (!g452) & (g1682) & (g475)) + ((!g538) & (!sk[95]) & (g452) & (!g1682) & (!g475)) + ((!g538) & (!sk[95]) & (g452) & (!g1682) & (g475)) + ((!g538) & (!sk[95]) & (g452) & (g1682) & (!g475)) + ((!g538) & (!sk[95]) & (g452) & (g1682) & (g475)) + ((!g538) & (sk[95]) & (!g452) & (!g1682) & (!g475)) + ((!g538) & (sk[95]) & (!g452) & (g1682) & (g475)) + ((!g538) & (sk[95]) & (g452) & (!g1682) & (g475)) + ((!g538) & (sk[95]) & (g452) & (g1682) & (!g475)) + ((g538) & (!sk[95]) & (!g452) & (g1682) & (!g475)) + ((g538) & (!sk[95]) & (!g452) & (g1682) & (g475)) + ((g538) & (!sk[95]) & (g452) & (!g1682) & (!g475)) + ((g538) & (!sk[95]) & (g452) & (!g1682) & (g475)) + ((g538) & (!sk[95]) & (g452) & (g1682) & (!g475)) + ((g538) & (!sk[95]) & (g452) & (g1682) & (g475)) + ((g538) & (sk[95]) & (!g452) & (!g1682) & (g475)) + ((g538) & (sk[95]) & (!g452) & (g1682) & (!g475)) + ((g538) & (sk[95]) & (g452) & (!g1682) & (!g475)) + ((g538) & (sk[95]) & (g452) & (g1682) & (g475)));
	assign g1907 = (((!sk[96]) & (!g1768) & (g475)) + ((!sk[96]) & (g1768) & (g475)) + ((sk[96]) & (!g1768) & (g475)) + ((sk[96]) & (g1768) & (!g475)));
	assign g1908 = (((!g1909) & (!sk[97]) & (g1910)) + ((!g1909) & (sk[97]) & (!g1910)) + ((g1909) & (!sk[97]) & (g1910)));
	assign g1909 = (((!g197) & (!sk[98]) & (g1911)) + ((!g197) & (sk[98]) & (g1911)) + ((g197) & (!sk[98]) & (g1911)));
	assign g1910 = (((!sk[99]) & (!g197) & (g1914)) + ((!sk[99]) & (g197) & (g1914)) + ((sk[99]) & (g197) & (g1914)));
	assign g1911 = (((!sk[100]) & (!g1912) & (g1913)) + ((!sk[100]) & (g1912) & (g1913)) + ((sk[100]) & (!g1912) & (!g1913)));
	assign g1912 = (((!sk[101]) & (!g1163) & (g1917)) + ((!sk[101]) & (g1163) & (g1917)) + ((sk[101]) & (!g1163) & (g1917)));
	assign g1913 = (((!g1163) & (!sk[102]) & (g1756)) + ((g1163) & (!sk[102]) & (g1756)) + ((g1163) & (sk[102]) & (g1756)));
	assign g1914 = (((!sk[103]) & (!g1915) & (g1916)) + ((!sk[103]) & (g1915) & (g1916)) + ((sk[103]) & (!g1915) & (!g1916)));
	assign g1915 = (((!g1163) & (!sk[104]) & (g1918)) + ((!g1163) & (sk[104]) & (g1918)) + ((g1163) & (!sk[104]) & (g1918)));
	assign g1916 = (((!g1163) & (!sk[105]) & (g1756)) + ((g1163) & (!sk[105]) & (g1756)) + ((g1163) & (sk[105]) & (!g1756)));
	assign g1917 = (((!sk[106]) & (!g388) & (!g381) & (g1566) & (!g189)) + ((!sk[106]) & (!g388) & (!g381) & (g1566) & (g189)) + ((!sk[106]) & (!g388) & (g381) & (!g1566) & (!g189)) + ((!sk[106]) & (!g388) & (g381) & (!g1566) & (g189)) + ((!sk[106]) & (!g388) & (g381) & (g1566) & (!g189)) + ((!sk[106]) & (!g388) & (g381) & (g1566) & (g189)) + ((!sk[106]) & (g388) & (!g381) & (g1566) & (!g189)) + ((!sk[106]) & (g388) & (!g381) & (g1566) & (g189)) + ((!sk[106]) & (g388) & (g381) & (!g1566) & (!g189)) + ((!sk[106]) & (g388) & (g381) & (!g1566) & (g189)) + ((!sk[106]) & (g388) & (g381) & (g1566) & (!g189)) + ((!sk[106]) & (g388) & (g381) & (g1566) & (g189)) + ((sk[106]) & (!g388) & (!g381) & (!g1566) & (g189)) + ((sk[106]) & (!g388) & (!g381) & (g1566) & (!g189)) + ((sk[106]) & (!g388) & (g381) & (!g1566) & (!g189)) + ((sk[106]) & (!g388) & (g381) & (g1566) & (g189)) + ((sk[106]) & (g388) & (!g381) & (!g1566) & (!g189)) + ((sk[106]) & (g388) & (!g381) & (g1566) & (g189)) + ((sk[106]) & (g388) & (g381) & (!g1566) & (g189)) + ((sk[106]) & (g388) & (g381) & (g1566) & (!g189)));
	assign g1918 = (((!g388) & (!g381) & (!sk[107]) & (g1566) & (!g189)) + ((!g388) & (!g381) & (!sk[107]) & (g1566) & (g189)) + ((!g388) & (!g381) & (sk[107]) & (!g1566) & (!g189)) + ((!g388) & (!g381) & (sk[107]) & (g1566) & (g189)) + ((!g388) & (g381) & (!sk[107]) & (!g1566) & (!g189)) + ((!g388) & (g381) & (!sk[107]) & (!g1566) & (g189)) + ((!g388) & (g381) & (!sk[107]) & (g1566) & (!g189)) + ((!g388) & (g381) & (!sk[107]) & (g1566) & (g189)) + ((!g388) & (g381) & (sk[107]) & (!g1566) & (g189)) + ((!g388) & (g381) & (sk[107]) & (g1566) & (!g189)) + ((g388) & (!g381) & (!sk[107]) & (g1566) & (!g189)) + ((g388) & (!g381) & (!sk[107]) & (g1566) & (g189)) + ((g388) & (!g381) & (sk[107]) & (!g1566) & (g189)) + ((g388) & (!g381) & (sk[107]) & (g1566) & (!g189)) + ((g388) & (g381) & (!sk[107]) & (!g1566) & (!g189)) + ((g388) & (g381) & (!sk[107]) & (!g1566) & (g189)) + ((g388) & (g381) & (!sk[107]) & (g1566) & (!g189)) + ((g388) & (g381) & (!sk[107]) & (g1566) & (g189)) + ((g388) & (g381) & (sk[107]) & (!g1566) & (!g189)) + ((g388) & (g381) & (sk[107]) & (g1566) & (g189)));
	assign g1919 = (((!g1920) & (!sk[108]) & (g1921)) + ((!g1920) & (sk[108]) & (!g1921)) + ((g1920) & (!sk[108]) & (g1921)));
	assign g1920 = (((!sk[109]) & (!g474) & (g1922)) + ((!sk[109]) & (g474) & (g1922)) + ((sk[109]) & (!g474) & (g1922)));
	assign g1921 = (((!sk[110]) & (!g474) & (g1925)) + ((!sk[110]) & (g474) & (g1925)) + ((sk[110]) & (g474) & (g1925)));
	assign g1922 = (((!g1923) & (!sk[111]) & (g1924)) + ((!g1923) & (sk[111]) & (!g1924)) + ((g1923) & (!sk[111]) & (g1924)));
	assign g1923 = (((!sk[112]) & (!g1163) & (g1928)) + ((!sk[112]) & (g1163) & (g1928)) + ((sk[112]) & (!g1163) & (g1928)));
	assign g1924 = (((!g1163) & (!sk[113]) & (g1929)) + ((g1163) & (!sk[113]) & (g1929)) + ((g1163) & (sk[113]) & (g1929)));
	assign g1925 = (((!sk[114]) & (!g1926) & (g1927)) + ((!sk[114]) & (g1926) & (g1927)) + ((sk[114]) & (!g1926) & (!g1927)));
	assign g1926 = (((!sk[115]) & (!g1163) & (g1930)) + ((!sk[115]) & (g1163) & (g1930)) + ((sk[115]) & (!g1163) & (g1930)));
	assign g1927 = (((!g1163) & (!sk[116]) & (g1931)) + ((g1163) & (!sk[116]) & (g1931)) + ((g1163) & (sk[116]) & (g1931)));
	assign g1928 = (((!g580) & (!sk[117]) & (!g531) & (g1682) & (!g539)) + ((!g580) & (!sk[117]) & (!g531) & (g1682) & (g539)) + ((!g580) & (!sk[117]) & (g531) & (!g1682) & (!g539)) + ((!g580) & (!sk[117]) & (g531) & (!g1682) & (g539)) + ((!g580) & (!sk[117]) & (g531) & (g1682) & (!g539)) + ((!g580) & (!sk[117]) & (g531) & (g1682) & (g539)) + ((!g580) & (sk[117]) & (!g531) & (!g1682) & (g539)) + ((!g580) & (sk[117]) & (!g531) & (g1682) & (!g539)) + ((!g580) & (sk[117]) & (g531) & (!g1682) & (!g539)) + ((!g580) & (sk[117]) & (g531) & (g1682) & (g539)) + ((g580) & (!sk[117]) & (!g531) & (g1682) & (!g539)) + ((g580) & (!sk[117]) & (!g531) & (g1682) & (g539)) + ((g580) & (!sk[117]) & (g531) & (!g1682) & (!g539)) + ((g580) & (!sk[117]) & (g531) & (!g1682) & (g539)) + ((g580) & (!sk[117]) & (g531) & (g1682) & (!g539)) + ((g580) & (!sk[117]) & (g531) & (g1682) & (g539)) + ((g580) & (sk[117]) & (!g531) & (!g1682) & (!g539)) + ((g580) & (sk[117]) & (!g531) & (g1682) & (g539)) + ((g580) & (sk[117]) & (g531) & (!g1682) & (g539)) + ((g580) & (sk[117]) & (g531) & (g1682) & (!g539)));
	assign g1929 = (((!g1681) & (!sk[118]) & (g539)) + ((!g1681) & (sk[118]) & (g539)) + ((g1681) & (!sk[118]) & (g539)) + ((g1681) & (sk[118]) & (!g539)));
	assign g1930 = (((!sk[119]) & (!g580) & (!g531) & (g1682) & (!g539)) + ((!sk[119]) & (!g580) & (!g531) & (g1682) & (g539)) + ((!sk[119]) & (!g580) & (g531) & (!g1682) & (!g539)) + ((!sk[119]) & (!g580) & (g531) & (!g1682) & (g539)) + ((!sk[119]) & (!g580) & (g531) & (g1682) & (!g539)) + ((!sk[119]) & (!g580) & (g531) & (g1682) & (g539)) + ((!sk[119]) & (g580) & (!g531) & (g1682) & (!g539)) + ((!sk[119]) & (g580) & (!g531) & (g1682) & (g539)) + ((!sk[119]) & (g580) & (g531) & (!g1682) & (!g539)) + ((!sk[119]) & (g580) & (g531) & (!g1682) & (g539)) + ((!sk[119]) & (g580) & (g531) & (g1682) & (!g539)) + ((!sk[119]) & (g580) & (g531) & (g1682) & (g539)) + ((sk[119]) & (!g580) & (!g531) & (!g1682) & (!g539)) + ((sk[119]) & (!g580) & (!g531) & (g1682) & (g539)) + ((sk[119]) & (!g580) & (g531) & (!g1682) & (g539)) + ((sk[119]) & (!g580) & (g531) & (g1682) & (!g539)) + ((sk[119]) & (g580) & (!g531) & (!g1682) & (g539)) + ((sk[119]) & (g580) & (!g531) & (g1682) & (!g539)) + ((sk[119]) & (g580) & (g531) & (!g1682) & (!g539)) + ((sk[119]) & (g580) & (g531) & (g1682) & (g539)));
	assign g1931 = (((!sk[120]) & (!g1681) & (g539)) + ((!sk[120]) & (g1681) & (g539)) + ((sk[120]) & (!g1681) & (g539)) + ((sk[120]) & (g1681) & (!g539)));
	assign g1932 = (((!sk[121]) & (!g1933) & (g1934)) + ((!sk[121]) & (g1933) & (g1934)) + ((sk[121]) & (!g1933) & (!g1934)));
	assign g1933 = (((!g212) & (!sk[122]) & (g1935)) + ((!g212) & (sk[122]) & (g1935)) + ((g212) & (!sk[122]) & (g1935)));
	assign g1934 = (((!g212) & (!sk[123]) & (g1938)) + ((g212) & (!sk[123]) & (g1938)) + ((g212) & (sk[123]) & (g1938)));
	assign g1935 = (((!sk[124]) & (!g1936) & (g1937)) + ((!sk[124]) & (g1936) & (g1937)) + ((sk[124]) & (!g1936) & (!g1937)));
	assign g1936 = (((!g1163) & (!sk[125]) & (g1941)) + ((!g1163) & (sk[125]) & (g1941)) + ((g1163) & (!sk[125]) & (g1941)));
	assign g1937 = (((!sk[126]) & (!g1163) & (g1645)) + ((!sk[126]) & (g1163) & (g1645)) + ((sk[126]) & (g1163) & (g1645)));
	assign g1938 = (((!g1939) & (!sk[127]) & (g1940)) + ((!g1939) & (sk[127]) & (!g1940)) + ((g1939) & (!sk[127]) & (g1940)));
	assign g1939 = (((!g1163) & (!sk[0]) & (g1942)) + ((!g1163) & (sk[0]) & (g1942)) + ((g1163) & (!sk[0]) & (g1942)));
	assign g1940 = (((!sk[1]) & (!g1163) & (g1645)) + ((!sk[1]) & (g1163) & (g1645)) + ((sk[1]) & (g1163) & (!g1645)));
	assign g1941 = (((!g339) & (!g275) & (!g1431) & (sk[2]) & (g147)) + ((!g339) & (!g275) & (g1431) & (!sk[2]) & (!g147)) + ((!g339) & (!g275) & (g1431) & (!sk[2]) & (g147)) + ((!g339) & (!g275) & (g1431) & (sk[2]) & (!g147)) + ((!g339) & (g275) & (!g1431) & (!sk[2]) & (!g147)) + ((!g339) & (g275) & (!g1431) & (!sk[2]) & (g147)) + ((!g339) & (g275) & (!g1431) & (sk[2]) & (!g147)) + ((!g339) & (g275) & (g1431) & (!sk[2]) & (!g147)) + ((!g339) & (g275) & (g1431) & (!sk[2]) & (g147)) + ((!g339) & (g275) & (g1431) & (sk[2]) & (g147)) + ((g339) & (!g275) & (!g1431) & (sk[2]) & (!g147)) + ((g339) & (!g275) & (g1431) & (!sk[2]) & (!g147)) + ((g339) & (!g275) & (g1431) & (!sk[2]) & (g147)) + ((g339) & (!g275) & (g1431) & (sk[2]) & (g147)) + ((g339) & (g275) & (!g1431) & (!sk[2]) & (!g147)) + ((g339) & (g275) & (!g1431) & (!sk[2]) & (g147)) + ((g339) & (g275) & (!g1431) & (sk[2]) & (g147)) + ((g339) & (g275) & (g1431) & (!sk[2]) & (!g147)) + ((g339) & (g275) & (g1431) & (!sk[2]) & (g147)) + ((g339) & (g275) & (g1431) & (sk[2]) & (!g147)));
	assign g1942 = (((!g339) & (!sk[3]) & (!g275) & (g1431) & (!g147)) + ((!g339) & (!sk[3]) & (!g275) & (g1431) & (g147)) + ((!g339) & (!sk[3]) & (g275) & (!g1431) & (!g147)) + ((!g339) & (!sk[3]) & (g275) & (!g1431) & (g147)) + ((!g339) & (!sk[3]) & (g275) & (g1431) & (!g147)) + ((!g339) & (!sk[3]) & (g275) & (g1431) & (g147)) + ((!g339) & (sk[3]) & (!g275) & (!g1431) & (!g147)) + ((!g339) & (sk[3]) & (!g275) & (g1431) & (g147)) + ((!g339) & (sk[3]) & (g275) & (!g1431) & (g147)) + ((!g339) & (sk[3]) & (g275) & (g1431) & (!g147)) + ((g339) & (!sk[3]) & (!g275) & (g1431) & (!g147)) + ((g339) & (!sk[3]) & (!g275) & (g1431) & (g147)) + ((g339) & (!sk[3]) & (g275) & (!g1431) & (!g147)) + ((g339) & (!sk[3]) & (g275) & (!g1431) & (g147)) + ((g339) & (!sk[3]) & (g275) & (g1431) & (!g147)) + ((g339) & (!sk[3]) & (g275) & (g1431) & (g147)) + ((g339) & (sk[3]) & (!g275) & (!g1431) & (g147)) + ((g339) & (sk[3]) & (!g275) & (g1431) & (!g147)) + ((g339) & (sk[3]) & (g275) & (!g1431) & (!g147)) + ((g339) & (sk[3]) & (g275) & (g1431) & (g147)));
	assign g1943 = (((!g1944) & (!sk[4]) & (g1945)) + ((!g1944) & (sk[4]) & (!g1945)) + ((g1944) & (!sk[4]) & (g1945)));
	assign g1944 = (((!sk[5]) & (!g965) & (g1946)) + ((!sk[5]) & (g965) & (g1946)) + ((sk[5]) & (!g965) & (g1946)));
	assign g1945 = (((!g965) & (!sk[6]) & (g1949)) + ((g965) & (!sk[6]) & (g1949)) + ((g965) & (sk[6]) & (g1949)));
	assign g1946 = (((!g1947) & (!sk[7]) & (g1948)) + ((!g1947) & (sk[7]) & (!g1948)) + ((g1947) & (!sk[7]) & (g1948)));
	assign g1947 = (((!sk[8]) & (!g1163) & (g1952)) + ((!sk[8]) & (g1163) & (g1952)) + ((sk[8]) & (!g1163) & (g1952)));
	assign g1948 = (((!sk[9]) & (!g1163) & (g1636)) + ((!sk[9]) & (g1163) & (g1636)) + ((sk[9]) & (g1163) & (g1636)));
	assign g1949 = (((!sk[10]) & (!g1950) & (g1951)) + ((!sk[10]) & (g1950) & (g1951)) + ((sk[10]) & (!g1950) & (!g1951)));
	assign g1950 = (((!g1163) & (!sk[11]) & (g1953)) + ((!g1163) & (sk[11]) & (g1953)) + ((g1163) & (!sk[11]) & (g1953)));
	assign g1951 = (((!sk[12]) & (!g1163) & (g1636)) + ((!sk[12]) & (g1163) & (g1636)) + ((sk[12]) & (g1163) & (!g1636)));
	assign g1952 = (((!g1156) & (!g1149) & (!g1329) & (sk[13]) & (g957)) + ((!g1156) & (!g1149) & (g1329) & (!sk[13]) & (!g957)) + ((!g1156) & (!g1149) & (g1329) & (!sk[13]) & (g957)) + ((!g1156) & (!g1149) & (g1329) & (sk[13]) & (!g957)) + ((!g1156) & (g1149) & (!g1329) & (!sk[13]) & (!g957)) + ((!g1156) & (g1149) & (!g1329) & (!sk[13]) & (g957)) + ((!g1156) & (g1149) & (!g1329) & (sk[13]) & (!g957)) + ((!g1156) & (g1149) & (g1329) & (!sk[13]) & (!g957)) + ((!g1156) & (g1149) & (g1329) & (!sk[13]) & (g957)) + ((!g1156) & (g1149) & (g1329) & (sk[13]) & (g957)) + ((g1156) & (!g1149) & (!g1329) & (sk[13]) & (!g957)) + ((g1156) & (!g1149) & (g1329) & (!sk[13]) & (!g957)) + ((g1156) & (!g1149) & (g1329) & (!sk[13]) & (g957)) + ((g1156) & (!g1149) & (g1329) & (sk[13]) & (g957)) + ((g1156) & (g1149) & (!g1329) & (!sk[13]) & (!g957)) + ((g1156) & (g1149) & (!g1329) & (!sk[13]) & (g957)) + ((g1156) & (g1149) & (!g1329) & (sk[13]) & (g957)) + ((g1156) & (g1149) & (g1329) & (!sk[13]) & (!g957)) + ((g1156) & (g1149) & (g1329) & (!sk[13]) & (g957)) + ((g1156) & (g1149) & (g1329) & (sk[13]) & (!g957)));
	assign g1953 = (((!g1156) & (!g1149) & (!g1329) & (sk[14]) & (!g957)) + ((!g1156) & (!g1149) & (g1329) & (!sk[14]) & (!g957)) + ((!g1156) & (!g1149) & (g1329) & (!sk[14]) & (g957)) + ((!g1156) & (!g1149) & (g1329) & (sk[14]) & (g957)) + ((!g1156) & (g1149) & (!g1329) & (!sk[14]) & (!g957)) + ((!g1156) & (g1149) & (!g1329) & (!sk[14]) & (g957)) + ((!g1156) & (g1149) & (!g1329) & (sk[14]) & (g957)) + ((!g1156) & (g1149) & (g1329) & (!sk[14]) & (!g957)) + ((!g1156) & (g1149) & (g1329) & (!sk[14]) & (g957)) + ((!g1156) & (g1149) & (g1329) & (sk[14]) & (!g957)) + ((g1156) & (!g1149) & (!g1329) & (sk[14]) & (g957)) + ((g1156) & (!g1149) & (g1329) & (!sk[14]) & (!g957)) + ((g1156) & (!g1149) & (g1329) & (!sk[14]) & (g957)) + ((g1156) & (!g1149) & (g1329) & (sk[14]) & (!g957)) + ((g1156) & (g1149) & (!g1329) & (!sk[14]) & (!g957)) + ((g1156) & (g1149) & (!g1329) & (!sk[14]) & (g957)) + ((g1156) & (g1149) & (!g1329) & (sk[14]) & (!g957)) + ((g1156) & (g1149) & (g1329) & (!sk[14]) & (!g957)) + ((g1156) & (g1149) & (g1329) & (!sk[14]) & (g957)) + ((g1156) & (g1149) & (g1329) & (sk[14]) & (g957)));
	assign g1954 = (((!sk[15]) & (!g1955) & (g1956)) + ((!sk[15]) & (g1955) & (g1956)) + ((sk[15]) & (!g1955) & (!g1956)));
	assign g1955 = (((!sk[16]) & (!g936) & (g1957)) + ((!sk[16]) & (g936) & (g1957)) + ((sk[16]) & (!g936) & (g1957)));
	assign g1956 = (((!g936) & (!sk[17]) & (g1960)) + ((g936) & (!sk[17]) & (g1960)) + ((g936) & (sk[17]) & (g1960)));
	assign g1957 = (((!g1958) & (!sk[18]) & (g1959)) + ((!g1958) & (sk[18]) & (!g1959)) + ((g1958) & (!sk[18]) & (g1959)));
	assign g1958 = (((!g1163) & (!sk[19]) & (g1963)) + ((!g1163) & (sk[19]) & (g1963)) + ((g1163) & (!sk[19]) & (g1963)));
	assign g1959 = (((!sk[20]) & (!g1163) & (g1964)) + ((!sk[20]) & (g1163) & (g1964)) + ((sk[20]) & (g1163) & (g1964)));
	assign g1960 = (((!g1961) & (!sk[21]) & (g1962)) + ((!g1961) & (sk[21]) & (!g1962)) + ((g1961) & (!sk[21]) & (g1962)));
	assign g1961 = (((!sk[22]) & (!g1163) & (g1965)) + ((!sk[22]) & (g1163) & (g1965)) + ((sk[22]) & (!g1163) & (g1965)));
	assign g1962 = (((!g1163) & (!sk[23]) & (g1966)) + ((g1163) & (!sk[23]) & (g1966)) + ((g1163) & (sk[23]) & (g1966)));
	assign g1963 = (((!g1135) & (!g964) & (!g1635) & (sk[24]) & (g944)) + ((!g1135) & (!g964) & (g1635) & (!sk[24]) & (!g944)) + ((!g1135) & (!g964) & (g1635) & (!sk[24]) & (g944)) + ((!g1135) & (!g964) & (g1635) & (sk[24]) & (!g944)) + ((!g1135) & (g964) & (!g1635) & (!sk[24]) & (!g944)) + ((!g1135) & (g964) & (!g1635) & (!sk[24]) & (g944)) + ((!g1135) & (g964) & (!g1635) & (sk[24]) & (!g944)) + ((!g1135) & (g964) & (g1635) & (!sk[24]) & (!g944)) + ((!g1135) & (g964) & (g1635) & (!sk[24]) & (g944)) + ((!g1135) & (g964) & (g1635) & (sk[24]) & (g944)) + ((g1135) & (!g964) & (!g1635) & (sk[24]) & (!g944)) + ((g1135) & (!g964) & (g1635) & (!sk[24]) & (!g944)) + ((g1135) & (!g964) & (g1635) & (!sk[24]) & (g944)) + ((g1135) & (!g964) & (g1635) & (sk[24]) & (g944)) + ((g1135) & (g964) & (!g1635) & (!sk[24]) & (!g944)) + ((g1135) & (g964) & (!g1635) & (!sk[24]) & (g944)) + ((g1135) & (g964) & (!g1635) & (sk[24]) & (g944)) + ((g1135) & (g964) & (g1635) & (!sk[24]) & (!g944)) + ((g1135) & (g964) & (g1635) & (!sk[24]) & (g944)) + ((g1135) & (g964) & (g1635) & (sk[24]) & (!g944)));
	assign g1964 = (((!sk[25]) & (!g1634) & (g944)) + ((!sk[25]) & (g1634) & (g944)) + ((sk[25]) & (!g1634) & (g944)) + ((sk[25]) & (g1634) & (!g944)));
	assign g1965 = (((!g1135) & (!g964) & (!g1635) & (sk[26]) & (!g944)) + ((!g1135) & (!g964) & (g1635) & (!sk[26]) & (!g944)) + ((!g1135) & (!g964) & (g1635) & (!sk[26]) & (g944)) + ((!g1135) & (!g964) & (g1635) & (sk[26]) & (g944)) + ((!g1135) & (g964) & (!g1635) & (!sk[26]) & (!g944)) + ((!g1135) & (g964) & (!g1635) & (!sk[26]) & (g944)) + ((!g1135) & (g964) & (!g1635) & (sk[26]) & (g944)) + ((!g1135) & (g964) & (g1635) & (!sk[26]) & (!g944)) + ((!g1135) & (g964) & (g1635) & (!sk[26]) & (g944)) + ((!g1135) & (g964) & (g1635) & (sk[26]) & (!g944)) + ((g1135) & (!g964) & (!g1635) & (sk[26]) & (g944)) + ((g1135) & (!g964) & (g1635) & (!sk[26]) & (!g944)) + ((g1135) & (!g964) & (g1635) & (!sk[26]) & (g944)) + ((g1135) & (!g964) & (g1635) & (sk[26]) & (!g944)) + ((g1135) & (g964) & (!g1635) & (!sk[26]) & (!g944)) + ((g1135) & (g964) & (!g1635) & (!sk[26]) & (g944)) + ((g1135) & (g964) & (!g1635) & (sk[26]) & (!g944)) + ((g1135) & (g964) & (g1635) & (!sk[26]) & (!g944)) + ((g1135) & (g964) & (g1635) & (!sk[26]) & (g944)) + ((g1135) & (g964) & (g1635) & (sk[26]) & (g944)));
	assign g1966 = (((!sk[27]) & (!g1634) & (g944)) + ((!sk[27]) & (g1634) & (g944)) + ((sk[27]) & (!g1634) & (g944)) + ((sk[27]) & (g1634) & (!g944)));
	assign g1967 = (((!sk[28]) & (!g1968) & (g1969)) + ((!sk[28]) & (g1968) & (g1969)) + ((sk[28]) & (!g1968) & (!g1969)));
	assign g1968 = (((!sk[29]) & (!g424) & (g1970)) + ((!sk[29]) & (g424) & (g1970)) + ((sk[29]) & (!g424) & (g1970)));
	assign g1969 = (((!sk[30]) & (!g424) & (g1973)) + ((!sk[30]) & (g424) & (g1973)) + ((sk[30]) & (g424) & (g1973)));
	assign g1970 = (((!g1971) & (!sk[31]) & (g1972)) + ((!g1971) & (sk[31]) & (!g1972)) + ((g1971) & (!sk[31]) & (g1972)));
	assign g1971 = (((!sk[32]) & (!g1163) & (g1976)) + ((!sk[32]) & (g1163) & (g1976)) + ((sk[32]) & (!g1163) & (g1976)));
	assign g1972 = (((!sk[33]) & (!g1163) & (g1977)) + ((!sk[33]) & (g1163) & (g1977)) + ((sk[33]) & (g1163) & (g1977)));
	assign g1973 = (((!g1974) & (!sk[34]) & (g1975)) + ((!g1974) & (sk[34]) & (!g1975)) + ((g1974) & (!sk[34]) & (g1975)));
	assign g1974 = (((!sk[35]) & (!g1163) & (g1978)) + ((!sk[35]) & (g1163) & (g1978)) + ((sk[35]) & (!g1163) & (g1978)));
	assign g1975 = (((!sk[36]) & (!g1163) & (g1979)) + ((!sk[36]) & (g1163) & (g1979)) + ((sk[36]) & (g1163) & (g1979)));
	assign g1976 = (((!sk[37]) & (!g580) & (!g545) & (g1175) & (!g617)) + ((!sk[37]) & (!g580) & (!g545) & (g1175) & (g617)) + ((!sk[37]) & (!g580) & (g545) & (!g1175) & (!g617)) + ((!sk[37]) & (!g580) & (g545) & (!g1175) & (g617)) + ((!sk[37]) & (!g580) & (g545) & (g1175) & (!g617)) + ((!sk[37]) & (!g580) & (g545) & (g1175) & (g617)) + ((!sk[37]) & (g580) & (!g545) & (g1175) & (!g617)) + ((!sk[37]) & (g580) & (!g545) & (g1175) & (g617)) + ((!sk[37]) & (g580) & (g545) & (!g1175) & (!g617)) + ((!sk[37]) & (g580) & (g545) & (!g1175) & (g617)) + ((!sk[37]) & (g580) & (g545) & (g1175) & (!g617)) + ((!sk[37]) & (g580) & (g545) & (g1175) & (g617)) + ((sk[37]) & (!g580) & (!g545) & (!g1175) & (g617)) + ((sk[37]) & (!g580) & (!g545) & (g1175) & (!g617)) + ((sk[37]) & (!g580) & (g545) & (!g1175) & (!g617)) + ((sk[37]) & (!g580) & (g545) & (g1175) & (g617)) + ((sk[37]) & (g580) & (!g545) & (!g1175) & (!g617)) + ((sk[37]) & (g580) & (!g545) & (g1175) & (g617)) + ((sk[37]) & (g580) & (g545) & (!g1175) & (g617)) + ((sk[37]) & (g580) & (g545) & (g1175) & (!g617)));
	assign g1977 = (((!sk[38]) & (!g1596) & (g617)) + ((!sk[38]) & (g1596) & (g617)) + ((sk[38]) & (!g1596) & (g617)) + ((sk[38]) & (g1596) & (!g617)));
	assign g1978 = (((!sk[39]) & (!g580) & (!g545) & (g1175) & (!g617)) + ((!sk[39]) & (!g580) & (!g545) & (g1175) & (g617)) + ((!sk[39]) & (!g580) & (g545) & (!g1175) & (!g617)) + ((!sk[39]) & (!g580) & (g545) & (!g1175) & (g617)) + ((!sk[39]) & (!g580) & (g545) & (g1175) & (!g617)) + ((!sk[39]) & (!g580) & (g545) & (g1175) & (g617)) + ((!sk[39]) & (g580) & (!g545) & (g1175) & (!g617)) + ((!sk[39]) & (g580) & (!g545) & (g1175) & (g617)) + ((!sk[39]) & (g580) & (g545) & (!g1175) & (!g617)) + ((!sk[39]) & (g580) & (g545) & (!g1175) & (g617)) + ((!sk[39]) & (g580) & (g545) & (g1175) & (!g617)) + ((!sk[39]) & (g580) & (g545) & (g1175) & (g617)) + ((sk[39]) & (!g580) & (!g545) & (!g1175) & (!g617)) + ((sk[39]) & (!g580) & (!g545) & (g1175) & (g617)) + ((sk[39]) & (!g580) & (g545) & (!g1175) & (g617)) + ((sk[39]) & (!g580) & (g545) & (g1175) & (!g617)) + ((sk[39]) & (g580) & (!g545) & (!g1175) & (g617)) + ((sk[39]) & (g580) & (!g545) & (g1175) & (!g617)) + ((sk[39]) & (g580) & (g545) & (!g1175) & (!g617)) + ((sk[39]) & (g580) & (g545) & (g1175) & (g617)));
	assign g1979 = (((!sk[40]) & (!g1596) & (g617)) + ((!sk[40]) & (g1596) & (g617)) + ((sk[40]) & (!g1596) & (g617)) + ((sk[40]) & (g1596) & (!g617)));
	assign g1980 = (((!sk[41]) & (!g1981) & (g1982)) + ((!sk[41]) & (g1981) & (g1982)) + ((sk[41]) & (!g1981) & (!g1982)));
	assign g1981 = (((!sk[42]) & (!g325) & (g1983)) + ((!sk[42]) & (g325) & (g1983)) + ((sk[42]) & (!g325) & (g1983)));
	assign g1982 = (((!g325) & (!sk[43]) & (g1986)) + ((g325) & (!sk[43]) & (g1986)) + ((g325) & (sk[43]) & (g1986)));
	assign g1983 = (((!sk[44]) & (!g1984) & (g1985)) + ((!sk[44]) & (g1984) & (g1985)) + ((sk[44]) & (!g1984) & (!g1985)));
	assign g1984 = (((!g1163) & (!sk[45]) & (g1989)) + ((!g1163) & (sk[45]) & (g1989)) + ((g1163) & (!sk[45]) & (g1989)));
	assign g1985 = (((!g1163) & (!sk[46]) & (g1579)) + ((g1163) & (!sk[46]) & (g1579)) + ((g1163) & (sk[46]) & (g1579)));
	assign g1986 = (((!sk[47]) & (!g1987) & (g1988)) + ((!sk[47]) & (g1987) & (g1988)) + ((sk[47]) & (!g1987) & (!g1988)));
	assign g1987 = (((!sk[48]) & (!g1163) & (g1990)) + ((!sk[48]) & (g1163) & (g1990)) + ((sk[48]) & (!g1163) & (g1990)));
	assign g1988 = (((!g1163) & (!sk[49]) & (g1579)) + ((g1163) & (!sk[49]) & (g1579)) + ((g1163) & (sk[49]) & (!g1579)));
	assign g1989 = (((!g388) & (!sk[50]) & (!g317) & (g1431) & (!g253)) + ((!g388) & (!sk[50]) & (!g317) & (g1431) & (g253)) + ((!g388) & (!sk[50]) & (g317) & (!g1431) & (!g253)) + ((!g388) & (!sk[50]) & (g317) & (!g1431) & (g253)) + ((!g388) & (!sk[50]) & (g317) & (g1431) & (!g253)) + ((!g388) & (!sk[50]) & (g317) & (g1431) & (g253)) + ((!g388) & (sk[50]) & (!g317) & (!g1431) & (g253)) + ((!g388) & (sk[50]) & (!g317) & (g1431) & (!g253)) + ((!g388) & (sk[50]) & (g317) & (!g1431) & (!g253)) + ((!g388) & (sk[50]) & (g317) & (g1431) & (g253)) + ((g388) & (!sk[50]) & (!g317) & (g1431) & (!g253)) + ((g388) & (!sk[50]) & (!g317) & (g1431) & (g253)) + ((g388) & (!sk[50]) & (g317) & (!g1431) & (!g253)) + ((g388) & (!sk[50]) & (g317) & (!g1431) & (g253)) + ((g388) & (!sk[50]) & (g317) & (g1431) & (!g253)) + ((g388) & (!sk[50]) & (g317) & (g1431) & (g253)) + ((g388) & (sk[50]) & (!g317) & (!g1431) & (!g253)) + ((g388) & (sk[50]) & (!g317) & (g1431) & (g253)) + ((g388) & (sk[50]) & (g317) & (!g1431) & (g253)) + ((g388) & (sk[50]) & (g317) & (g1431) & (!g253)));
	assign g1990 = (((!sk[51]) & (!g388) & (!g317) & (g1431) & (!g253)) + ((!sk[51]) & (!g388) & (!g317) & (g1431) & (g253)) + ((!sk[51]) & (!g388) & (g317) & (!g1431) & (!g253)) + ((!sk[51]) & (!g388) & (g317) & (!g1431) & (g253)) + ((!sk[51]) & (!g388) & (g317) & (g1431) & (!g253)) + ((!sk[51]) & (!g388) & (g317) & (g1431) & (g253)) + ((!sk[51]) & (g388) & (!g317) & (g1431) & (!g253)) + ((!sk[51]) & (g388) & (!g317) & (g1431) & (g253)) + ((!sk[51]) & (g388) & (g317) & (!g1431) & (!g253)) + ((!sk[51]) & (g388) & (g317) & (!g1431) & (g253)) + ((!sk[51]) & (g388) & (g317) & (g1431) & (!g253)) + ((!sk[51]) & (g388) & (g317) & (g1431) & (g253)) + ((sk[51]) & (!g388) & (!g317) & (!g1431) & (!g253)) + ((sk[51]) & (!g388) & (!g317) & (g1431) & (g253)) + ((sk[51]) & (!g388) & (g317) & (!g1431) & (g253)) + ((sk[51]) & (!g388) & (g317) & (g1431) & (!g253)) + ((sk[51]) & (g388) & (!g317) & (!g1431) & (g253)) + ((sk[51]) & (g388) & (!g317) & (g1431) & (!g253)) + ((sk[51]) & (g388) & (g317) & (!g1431) & (!g253)) + ((sk[51]) & (g388) & (g317) & (g1431) & (g253)));
	assign g1991 = (((!sk[52]) & (!g1992) & (g1993)) + ((!sk[52]) & (g1992) & (g1993)) + ((sk[52]) & (!g1992) & (!g1993)));
	assign g1992 = (((!g232) & (!sk[53]) & (g1994)) + ((!g232) & (sk[53]) & (g1994)) + ((g232) & (!sk[53]) & (g1994)));
	assign g1993 = (((!g232) & (!sk[54]) & (g1997)) + ((g232) & (!sk[54]) & (g1997)) + ((g232) & (sk[54]) & (g1997)));
	assign g1994 = (((!g1995) & (!sk[55]) & (g1996)) + ((!g1995) & (sk[55]) & (!g1996)) + ((g1995) & (!sk[55]) & (g1996)));
	assign g1995 = (((!sk[56]) & (!g1163) & (g2000)) + ((!sk[56]) & (g1163) & (g2000)) + ((sk[56]) & (!g1163) & (g2000)));
	assign g1996 = (((!g1163) & (!sk[57]) & (g2001)) + ((g1163) & (!sk[57]) & (g2001)) + ((g1163) & (sk[57]) & (g2001)));
	assign g1997 = (((!sk[58]) & (!g1998) & (g1999)) + ((!sk[58]) & (g1998) & (g1999)) + ((sk[58]) & (!g1998) & (!g1999)));
	assign g1998 = (((!sk[59]) & (!g1163) & (g2002)) + ((!sk[59]) & (g1163) & (g2002)) + ((sk[59]) & (!g1163) & (g2002)));
	assign g1999 = (((!sk[60]) & (!g1163) & (g2003)) + ((!sk[60]) & (g1163) & (g2003)) + ((sk[60]) & (g1163) & (g2003)));
	assign g2000 = (((!g367) & (!sk[61]) & (!g260) & (g1429) & (!g304)) + ((!g367) & (!sk[61]) & (!g260) & (g1429) & (g304)) + ((!g367) & (!sk[61]) & (g260) & (!g1429) & (!g304)) + ((!g367) & (!sk[61]) & (g260) & (!g1429) & (g304)) + ((!g367) & (!sk[61]) & (g260) & (g1429) & (!g304)) + ((!g367) & (!sk[61]) & (g260) & (g1429) & (g304)) + ((!g367) & (sk[61]) & (!g260) & (!g1429) & (g304)) + ((!g367) & (sk[61]) & (!g260) & (g1429) & (!g304)) + ((!g367) & (sk[61]) & (g260) & (!g1429) & (!g304)) + ((!g367) & (sk[61]) & (g260) & (g1429) & (g304)) + ((g367) & (!sk[61]) & (!g260) & (g1429) & (!g304)) + ((g367) & (!sk[61]) & (!g260) & (g1429) & (g304)) + ((g367) & (!sk[61]) & (g260) & (!g1429) & (!g304)) + ((g367) & (!sk[61]) & (g260) & (!g1429) & (g304)) + ((g367) & (!sk[61]) & (g260) & (g1429) & (!g304)) + ((g367) & (!sk[61]) & (g260) & (g1429) & (g304)) + ((g367) & (sk[61]) & (!g260) & (!g1429) & (!g304)) + ((g367) & (sk[61]) & (!g260) & (g1429) & (g304)) + ((g367) & (sk[61]) & (g260) & (!g1429) & (g304)) + ((g367) & (sk[61]) & (g260) & (g1429) & (!g304)));
	assign g2001 = (((!sk[62]) & (!g1578) & (g304)) + ((!sk[62]) & (g1578) & (g304)) + ((sk[62]) & (!g1578) & (g304)) + ((sk[62]) & (g1578) & (!g304)));
	assign g2002 = (((!g367) & (!g260) & (!g1429) & (sk[63]) & (!g304)) + ((!g367) & (!g260) & (g1429) & (!sk[63]) & (!g304)) + ((!g367) & (!g260) & (g1429) & (!sk[63]) & (g304)) + ((!g367) & (!g260) & (g1429) & (sk[63]) & (g304)) + ((!g367) & (g260) & (!g1429) & (!sk[63]) & (!g304)) + ((!g367) & (g260) & (!g1429) & (!sk[63]) & (g304)) + ((!g367) & (g260) & (!g1429) & (sk[63]) & (g304)) + ((!g367) & (g260) & (g1429) & (!sk[63]) & (!g304)) + ((!g367) & (g260) & (g1429) & (!sk[63]) & (g304)) + ((!g367) & (g260) & (g1429) & (sk[63]) & (!g304)) + ((g367) & (!g260) & (!g1429) & (sk[63]) & (g304)) + ((g367) & (!g260) & (g1429) & (!sk[63]) & (!g304)) + ((g367) & (!g260) & (g1429) & (!sk[63]) & (g304)) + ((g367) & (!g260) & (g1429) & (sk[63]) & (!g304)) + ((g367) & (g260) & (!g1429) & (!sk[63]) & (!g304)) + ((g367) & (g260) & (!g1429) & (!sk[63]) & (g304)) + ((g367) & (g260) & (!g1429) & (sk[63]) & (!g304)) + ((g367) & (g260) & (g1429) & (!sk[63]) & (!g304)) + ((g367) & (g260) & (g1429) & (!sk[63]) & (g304)) + ((g367) & (g260) & (g1429) & (sk[63]) & (g304)));
	assign g2003 = (((!g1578) & (!sk[64]) & (g304)) + ((!g1578) & (sk[64]) & (g304)) + ((g1578) & (!sk[64]) & (g304)) + ((g1578) & (sk[64]) & (!g304)));
	assign g2004 = (((!sk[65]) & (!g2005) & (g2006)) + ((!sk[65]) & (g2005) & (g2006)) + ((sk[65]) & (!g2005) & (!g2006)));
	assign g2005 = (((!sk[66]) & (!g211) & (g2007)) + ((!sk[66]) & (g211) & (g2007)) + ((sk[66]) & (!g211) & (g2007)));
	assign g2006 = (((!g211) & (!sk[67]) & (g2010)) + ((g211) & (!sk[67]) & (g2010)) + ((g211) & (sk[67]) & (g2010)));
	assign g2007 = (((!sk[68]) & (!g2008) & (g2009)) + ((!sk[68]) & (g2008) & (g2009)) + ((sk[68]) & (!g2008) & (!g2009)));
	assign g2008 = (((!g1163) & (!sk[69]) & (g2013)) + ((!g1163) & (sk[69]) & (g2013)) + ((g1163) & (!sk[69]) & (g2013)));
	assign g2009 = (((!g1163) & (!sk[70]) & (g2014)) + ((g1163) & (!sk[70]) & (g2014)) + ((g1163) & (sk[70]) & (g2014)));
	assign g2010 = (((!sk[71]) & (!g2011) & (g2012)) + ((!sk[71]) & (g2011) & (g2012)) + ((sk[71]) & (!g2011) & (!g2012)));
	assign g2011 = (((!g1163) & (!sk[72]) & (g2015)) + ((!g1163) & (sk[72]) & (g2015)) + ((g1163) & (!sk[72]) & (g2015)));
	assign g2012 = (((!sk[73]) & (!g1163) & (g2016)) + ((!sk[73]) & (g1163) & (g2016)) + ((sk[73]) & (g1163) & (g2016)));
	assign g2013 = (((!g346) & (!sk[74]) & (!g260) & (g1415) & (!g283)) + ((!g346) & (!sk[74]) & (!g260) & (g1415) & (g283)) + ((!g346) & (!sk[74]) & (g260) & (!g1415) & (!g283)) + ((!g346) & (!sk[74]) & (g260) & (!g1415) & (g283)) + ((!g346) & (!sk[74]) & (g260) & (g1415) & (!g283)) + ((!g346) & (!sk[74]) & (g260) & (g1415) & (g283)) + ((!g346) & (sk[74]) & (!g260) & (!g1415) & (g283)) + ((!g346) & (sk[74]) & (!g260) & (g1415) & (!g283)) + ((!g346) & (sk[74]) & (g260) & (!g1415) & (!g283)) + ((!g346) & (sk[74]) & (g260) & (g1415) & (g283)) + ((g346) & (!sk[74]) & (!g260) & (g1415) & (!g283)) + ((g346) & (!sk[74]) & (!g260) & (g1415) & (g283)) + ((g346) & (!sk[74]) & (g260) & (!g1415) & (!g283)) + ((g346) & (!sk[74]) & (g260) & (!g1415) & (g283)) + ((g346) & (!sk[74]) & (g260) & (g1415) & (!g283)) + ((g346) & (!sk[74]) & (g260) & (g1415) & (g283)) + ((g346) & (sk[74]) & (!g260) & (!g1415) & (!g283)) + ((g346) & (sk[74]) & (!g260) & (g1415) & (g283)) + ((g346) & (sk[74]) & (g260) & (!g1415) & (g283)) + ((g346) & (sk[74]) & (g260) & (g1415) & (!g283)));
	assign g2014 = (((!g1568) & (!sk[75]) & (g283)) + ((!g1568) & (sk[75]) & (g283)) + ((g1568) & (!sk[75]) & (g283)) + ((g1568) & (sk[75]) & (!g283)));
	assign g2015 = (((!g346) & (!g260) & (!sk[76]) & (g1415) & (!g283)) + ((!g346) & (!g260) & (!sk[76]) & (g1415) & (g283)) + ((!g346) & (!g260) & (sk[76]) & (!g1415) & (!g283)) + ((!g346) & (!g260) & (sk[76]) & (g1415) & (g283)) + ((!g346) & (g260) & (!sk[76]) & (!g1415) & (!g283)) + ((!g346) & (g260) & (!sk[76]) & (!g1415) & (g283)) + ((!g346) & (g260) & (!sk[76]) & (g1415) & (!g283)) + ((!g346) & (g260) & (!sk[76]) & (g1415) & (g283)) + ((!g346) & (g260) & (sk[76]) & (!g1415) & (g283)) + ((!g346) & (g260) & (sk[76]) & (g1415) & (!g283)) + ((g346) & (!g260) & (!sk[76]) & (g1415) & (!g283)) + ((g346) & (!g260) & (!sk[76]) & (g1415) & (g283)) + ((g346) & (!g260) & (sk[76]) & (!g1415) & (g283)) + ((g346) & (!g260) & (sk[76]) & (g1415) & (!g283)) + ((g346) & (g260) & (!sk[76]) & (!g1415) & (!g283)) + ((g346) & (g260) & (!sk[76]) & (!g1415) & (g283)) + ((g346) & (g260) & (!sk[76]) & (g1415) & (!g283)) + ((g346) & (g260) & (!sk[76]) & (g1415) & (g283)) + ((g346) & (g260) & (sk[76]) & (!g1415) & (!g283)) + ((g346) & (g260) & (sk[76]) & (g1415) & (g283)));
	assign g2016 = (((!g1568) & (!sk[77]) & (g283)) + ((!g1568) & (sk[77]) & (g283)) + ((g1568) & (!sk[77]) & (g283)) + ((g1568) & (sk[77]) & (!g283)));
	assign g2017 = (((!g2018) & (!sk[78]) & (g2019)) + ((!g2018) & (sk[78]) & (!g2019)) + ((g2018) & (!sk[78]) & (g2019)));
	assign g2018 = (((!g673) & (!sk[79]) & (g2020)) + ((!g673) & (sk[79]) & (g2020)) + ((g673) & (!sk[79]) & (g2020)));
	assign g2019 = (((!g673) & (!sk[80]) & (g2023)) + ((g673) & (!sk[80]) & (g2023)) + ((g673) & (sk[80]) & (g2023)));
	assign g2020 = (((!sk[81]) & (!g2021) & (g2022)) + ((!sk[81]) & (g2021) & (g2022)) + ((sk[81]) & (!g2021) & (!g2022)));
	assign g2021 = (((!g1163) & (!sk[82]) & (g2026)) + ((!g1163) & (sk[82]) & (g2026)) + ((g1163) & (!sk[82]) & (g2026)));
	assign g2022 = (((!g1163) & (!sk[83]) & (g2027)) + ((g1163) & (!sk[83]) & (g2027)) + ((g1163) & (sk[83]) & (g2027)));
	assign g2023 = (((!g2024) & (!sk[84]) & (g2025)) + ((!g2024) & (sk[84]) & (!g2025)) + ((g2024) & (!sk[84]) & (g2025)));
	assign g2024 = (((!sk[85]) & (!g1163) & (g2028)) + ((!sk[85]) & (g1163) & (g2028)) + ((sk[85]) & (!g1163) & (g2028)));
	assign g2025 = (((!g1163) & (!sk[86]) & (g2029)) + ((g1163) & (!sk[86]) & (g2029)) + ((g1163) & (sk[86]) & (g2029)));
	assign g2026 = (((!g872) & (!g708) & (!g1514) & (sk[87]) & (g681)) + ((!g872) & (!g708) & (g1514) & (!sk[87]) & (!g681)) + ((!g872) & (!g708) & (g1514) & (!sk[87]) & (g681)) + ((!g872) & (!g708) & (g1514) & (sk[87]) & (!g681)) + ((!g872) & (g708) & (!g1514) & (!sk[87]) & (!g681)) + ((!g872) & (g708) & (!g1514) & (!sk[87]) & (g681)) + ((!g872) & (g708) & (!g1514) & (sk[87]) & (!g681)) + ((!g872) & (g708) & (g1514) & (!sk[87]) & (!g681)) + ((!g872) & (g708) & (g1514) & (!sk[87]) & (g681)) + ((!g872) & (g708) & (g1514) & (sk[87]) & (g681)) + ((g872) & (!g708) & (!g1514) & (sk[87]) & (!g681)) + ((g872) & (!g708) & (g1514) & (!sk[87]) & (!g681)) + ((g872) & (!g708) & (g1514) & (!sk[87]) & (g681)) + ((g872) & (!g708) & (g1514) & (sk[87]) & (g681)) + ((g872) & (g708) & (!g1514) & (!sk[87]) & (!g681)) + ((g872) & (g708) & (!g1514) & (!sk[87]) & (g681)) + ((g872) & (g708) & (!g1514) & (sk[87]) & (g681)) + ((g872) & (g708) & (g1514) & (!sk[87]) & (!g681)) + ((g872) & (g708) & (g1514) & (!sk[87]) & (g681)) + ((g872) & (g708) & (g1514) & (sk[87]) & (!g681)));
	assign g2027 = (((!g1513) & (!sk[88]) & (g681)) + ((!g1513) & (sk[88]) & (g681)) + ((g1513) & (!sk[88]) & (g681)) + ((g1513) & (sk[88]) & (!g681)));
	assign g2028 = (((!g872) & (!g708) & (!g1514) & (sk[89]) & (!g681)) + ((!g872) & (!g708) & (g1514) & (!sk[89]) & (!g681)) + ((!g872) & (!g708) & (g1514) & (!sk[89]) & (g681)) + ((!g872) & (!g708) & (g1514) & (sk[89]) & (g681)) + ((!g872) & (g708) & (!g1514) & (!sk[89]) & (!g681)) + ((!g872) & (g708) & (!g1514) & (!sk[89]) & (g681)) + ((!g872) & (g708) & (!g1514) & (sk[89]) & (g681)) + ((!g872) & (g708) & (g1514) & (!sk[89]) & (!g681)) + ((!g872) & (g708) & (g1514) & (!sk[89]) & (g681)) + ((!g872) & (g708) & (g1514) & (sk[89]) & (!g681)) + ((g872) & (!g708) & (!g1514) & (sk[89]) & (g681)) + ((g872) & (!g708) & (g1514) & (!sk[89]) & (!g681)) + ((g872) & (!g708) & (g1514) & (!sk[89]) & (g681)) + ((g872) & (!g708) & (g1514) & (sk[89]) & (!g681)) + ((g872) & (g708) & (!g1514) & (!sk[89]) & (!g681)) + ((g872) & (g708) & (!g1514) & (!sk[89]) & (g681)) + ((g872) & (g708) & (!g1514) & (sk[89]) & (!g681)) + ((g872) & (g708) & (g1514) & (!sk[89]) & (!g681)) + ((g872) & (g708) & (g1514) & (!sk[89]) & (g681)) + ((g872) & (g708) & (g1514) & (sk[89]) & (g681)));
	assign g2029 = (((!g1513) & (!sk[90]) & (g681)) + ((!g1513) & (sk[90]) & (g681)) + ((g1513) & (!sk[90]) & (g681)) + ((g1513) & (sk[90]) & (!g681)));
	assign g2030 = (((!sk[91]) & (!g2031) & (g2032)) + ((!sk[91]) & (g2031) & (g2032)) + ((sk[91]) & (!g2031) & (!g2032)));
	assign g2031 = (((!g303) & (!sk[92]) & (g2033)) + ((!g303) & (sk[92]) & (g2033)) + ((g303) & (!sk[92]) & (g2033)));
	assign g2032 = (((!g303) & (!sk[93]) & (g2036)) + ((g303) & (!sk[93]) & (g2036)) + ((g303) & (sk[93]) & (g2036)));
	assign g2033 = (((!g2034) & (!sk[94]) & (g2035)) + ((!g2034) & (sk[94]) & (!g2035)) + ((g2034) & (!sk[94]) & (g2035)));
	assign g2034 = (((!g1163) & (!sk[95]) & (g2039)) + ((!g1163) & (sk[95]) & (g2039)) + ((g1163) & (!sk[95]) & (g2039)));
	assign g2035 = (((!g1163) & (!sk[96]) & (g2040)) + ((g1163) & (!sk[96]) & (g2040)) + ((g1163) & (sk[96]) & (g2040)));
	assign g2036 = (((!sk[97]) & (!g2037) & (g2038)) + ((!sk[97]) & (g2037) & (g2038)) + ((sk[97]) & (!g2037) & (!g2038)));
	assign g2037 = (((!g1163) & (!sk[98]) & (g2041)) + ((!g1163) & (sk[98]) & (g2041)) + ((g1163) & (!sk[98]) & (g2041)));
	assign g2038 = (((!g1163) & (!sk[99]) & (g2042)) + ((g1163) & (!sk[99]) & (g2042)) + ((g1163) & (sk[99]) & (g2042)));
	assign g2039 = (((!g388) & (!g360) & (!sk[100]) & (g1429) & (!g368)) + ((!g388) & (!g360) & (!sk[100]) & (g1429) & (g368)) + ((!g388) & (!g360) & (sk[100]) & (!g1429) & (g368)) + ((!g388) & (!g360) & (sk[100]) & (g1429) & (!g368)) + ((!g388) & (g360) & (!sk[100]) & (!g1429) & (!g368)) + ((!g388) & (g360) & (!sk[100]) & (!g1429) & (g368)) + ((!g388) & (g360) & (!sk[100]) & (g1429) & (!g368)) + ((!g388) & (g360) & (!sk[100]) & (g1429) & (g368)) + ((!g388) & (g360) & (sk[100]) & (!g1429) & (!g368)) + ((!g388) & (g360) & (sk[100]) & (g1429) & (g368)) + ((g388) & (!g360) & (!sk[100]) & (g1429) & (!g368)) + ((g388) & (!g360) & (!sk[100]) & (g1429) & (g368)) + ((g388) & (!g360) & (sk[100]) & (!g1429) & (!g368)) + ((g388) & (!g360) & (sk[100]) & (g1429) & (g368)) + ((g388) & (g360) & (!sk[100]) & (!g1429) & (!g368)) + ((g388) & (g360) & (!sk[100]) & (!g1429) & (g368)) + ((g388) & (g360) & (!sk[100]) & (g1429) & (!g368)) + ((g388) & (g360) & (!sk[100]) & (g1429) & (g368)) + ((g388) & (g360) & (sk[100]) & (!g1429) & (g368)) + ((g388) & (g360) & (sk[100]) & (g1429) & (!g368)));
	assign g2040 = (((!sk[101]) & (!g1428) & (g368)) + ((!sk[101]) & (g1428) & (g368)) + ((sk[101]) & (!g1428) & (g368)) + ((sk[101]) & (g1428) & (!g368)));
	assign g2041 = (((!g388) & (!sk[102]) & (!g360) & (g1429) & (!g368)) + ((!g388) & (!sk[102]) & (!g360) & (g1429) & (g368)) + ((!g388) & (!sk[102]) & (g360) & (!g1429) & (!g368)) + ((!g388) & (!sk[102]) & (g360) & (!g1429) & (g368)) + ((!g388) & (!sk[102]) & (g360) & (g1429) & (!g368)) + ((!g388) & (!sk[102]) & (g360) & (g1429) & (g368)) + ((!g388) & (sk[102]) & (!g360) & (!g1429) & (!g368)) + ((!g388) & (sk[102]) & (!g360) & (g1429) & (g368)) + ((!g388) & (sk[102]) & (g360) & (!g1429) & (g368)) + ((!g388) & (sk[102]) & (g360) & (g1429) & (!g368)) + ((g388) & (!sk[102]) & (!g360) & (g1429) & (!g368)) + ((g388) & (!sk[102]) & (!g360) & (g1429) & (g368)) + ((g388) & (!sk[102]) & (g360) & (!g1429) & (!g368)) + ((g388) & (!sk[102]) & (g360) & (!g1429) & (g368)) + ((g388) & (!sk[102]) & (g360) & (g1429) & (!g368)) + ((g388) & (!sk[102]) & (g360) & (g1429) & (g368)) + ((g388) & (sk[102]) & (!g360) & (!g1429) & (g368)) + ((g388) & (sk[102]) & (!g360) & (g1429) & (!g368)) + ((g388) & (sk[102]) & (g360) & (!g1429) & (!g368)) + ((g388) & (sk[102]) & (g360) & (g1429) & (g368)));
	assign g2042 = (((!sk[103]) & (!g1428) & (g368)) + ((!sk[103]) & (g1428) & (g368)) + ((sk[103]) & (!g1428) & (g368)) + ((sk[103]) & (g1428) & (!g368)));
	assign g2043 = (((!g2044) & (!sk[104]) & (g2045)) + ((!g2044) & (sk[104]) & (!g2045)) + ((g2044) & (!sk[104]) & (g2045)));
	assign g2044 = (((!sk[105]) & (!g282) & (g2046)) + ((!sk[105]) & (g282) & (g2046)) + ((sk[105]) & (!g282) & (g2046)));
	assign g2045 = (((!sk[106]) & (!g282) & (g2049)) + ((!sk[106]) & (g282) & (g2049)) + ((sk[106]) & (g282) & (g2049)));
	assign g2046 = (((!g2047) & (!sk[107]) & (g2048)) + ((!g2047) & (sk[107]) & (!g2048)) + ((g2047) & (!sk[107]) & (g2048)));
	assign g2047 = (((!sk[108]) & (!g1163) & (g2052)) + ((!sk[108]) & (g1163) & (g2052)) + ((sk[108]) & (!g1163) & (g2052)));
	assign g2048 = (((!g1163) & (!sk[109]) & (g2053)) + ((g1163) & (!sk[109]) & (g2053)) + ((g1163) & (sk[109]) & (g2053)));
	assign g2049 = (((!sk[110]) & (!g2050) & (g2051)) + ((!sk[110]) & (g2050) & (g2051)) + ((sk[110]) & (!g2050) & (!g2051)));
	assign g2050 = (((!sk[111]) & (!g1163) & (g2054)) + ((!sk[111]) & (g1163) & (g2054)) + ((sk[111]) & (!g1163) & (g2054)));
	assign g2051 = (((!sk[112]) & (!g1163) & (g2055)) + ((!sk[112]) & (g1163) & (g2055)) + ((sk[112]) & (g1163) & (g2055)));
	assign g2052 = (((!g388) & (!sk[113]) & (!g339) & (g1415) & (!g347)) + ((!g388) & (!sk[113]) & (!g339) & (g1415) & (g347)) + ((!g388) & (!sk[113]) & (g339) & (!g1415) & (!g347)) + ((!g388) & (!sk[113]) & (g339) & (!g1415) & (g347)) + ((!g388) & (!sk[113]) & (g339) & (g1415) & (!g347)) + ((!g388) & (!sk[113]) & (g339) & (g1415) & (g347)) + ((!g388) & (sk[113]) & (!g339) & (!g1415) & (g347)) + ((!g388) & (sk[113]) & (!g339) & (g1415) & (!g347)) + ((!g388) & (sk[113]) & (g339) & (!g1415) & (!g347)) + ((!g388) & (sk[113]) & (g339) & (g1415) & (g347)) + ((g388) & (!sk[113]) & (!g339) & (g1415) & (!g347)) + ((g388) & (!sk[113]) & (!g339) & (g1415) & (g347)) + ((g388) & (!sk[113]) & (g339) & (!g1415) & (!g347)) + ((g388) & (!sk[113]) & (g339) & (!g1415) & (g347)) + ((g388) & (!sk[113]) & (g339) & (g1415) & (!g347)) + ((g388) & (!sk[113]) & (g339) & (g1415) & (g347)) + ((g388) & (sk[113]) & (!g339) & (!g1415) & (!g347)) + ((g388) & (sk[113]) & (!g339) & (g1415) & (g347)) + ((g388) & (sk[113]) & (g339) & (!g1415) & (g347)) + ((g388) & (sk[113]) & (g339) & (g1415) & (!g347)));
	assign g2053 = (((!g1414) & (!sk[114]) & (g347)) + ((!g1414) & (sk[114]) & (g347)) + ((g1414) & (!sk[114]) & (g347)) + ((g1414) & (sk[114]) & (!g347)));
	assign g2054 = (((!g388) & (!g339) & (!g1415) & (sk[115]) & (!g347)) + ((!g388) & (!g339) & (g1415) & (!sk[115]) & (!g347)) + ((!g388) & (!g339) & (g1415) & (!sk[115]) & (g347)) + ((!g388) & (!g339) & (g1415) & (sk[115]) & (g347)) + ((!g388) & (g339) & (!g1415) & (!sk[115]) & (!g347)) + ((!g388) & (g339) & (!g1415) & (!sk[115]) & (g347)) + ((!g388) & (g339) & (!g1415) & (sk[115]) & (g347)) + ((!g388) & (g339) & (g1415) & (!sk[115]) & (!g347)) + ((!g388) & (g339) & (g1415) & (!sk[115]) & (g347)) + ((!g388) & (g339) & (g1415) & (sk[115]) & (!g347)) + ((g388) & (!g339) & (!g1415) & (sk[115]) & (g347)) + ((g388) & (!g339) & (g1415) & (!sk[115]) & (!g347)) + ((g388) & (!g339) & (g1415) & (!sk[115]) & (g347)) + ((g388) & (!g339) & (g1415) & (sk[115]) & (!g347)) + ((g388) & (g339) & (!g1415) & (!sk[115]) & (!g347)) + ((g388) & (g339) & (!g1415) & (!sk[115]) & (g347)) + ((g388) & (g339) & (!g1415) & (sk[115]) & (!g347)) + ((g388) & (g339) & (g1415) & (!sk[115]) & (!g347)) + ((g388) & (g339) & (g1415) & (!sk[115]) & (g347)) + ((g388) & (g339) & (g1415) & (sk[115]) & (g347)));
	assign g2055 = (((!g1414) & (!sk[116]) & (g347)) + ((!g1414) & (sk[116]) & (g347)) + ((g1414) & (!sk[116]) & (g347)) + ((g1414) & (sk[116]) & (!g347)));
	assign g2056 = (((!g2057) & (!sk[117]) & (g2058)) + ((!g2057) & (sk[117]) & (!g2058)) + ((g2057) & (!sk[117]) & (g2058)));
	assign g2057 = (((!sk[118]) & (!g993) & (g2059)) + ((!sk[118]) & (g993) & (g2059)) + ((sk[118]) & (!g993) & (g2059)));
	assign g2058 = (((!g993) & (!sk[119]) & (g2062)) + ((g993) & (!sk[119]) & (g2062)) + ((g993) & (sk[119]) & (g2062)));
	assign g2059 = (((!g2060) & (!sk[120]) & (g2061)) + ((!g2060) & (sk[120]) & (!g2061)) + ((g2060) & (!sk[120]) & (g2061)));
	assign g2060 = (((!g1163) & (!sk[121]) & (g2065)) + ((!g1163) & (sk[121]) & (g2065)) + ((g1163) & (!sk[121]) & (g2065)));
	assign g2061 = (((!g1163) & (!sk[122]) & (g2066)) + ((g1163) & (!sk[122]) & (g2066)) + ((g1163) & (sk[122]) & (g2066)));
	assign g2062 = (((!sk[123]) & (!g2063) & (g2064)) + ((!sk[123]) & (g2063) & (g2064)) + ((sk[123]) & (!g2063) & (!g2064)));
	assign g2063 = (((!g1163) & (!sk[124]) & (g2067)) + ((!g1163) & (sk[124]) & (g2067)) + ((g1163) & (!sk[124]) & (g2067)));
	assign g2064 = (((!g1163) & (!sk[125]) & (g2068)) + ((g1163) & (!sk[125]) & (g2068)) + ((g1163) & (sk[125]) & (g2068)));
	assign g2065 = (((!g1128) & (!g1028) & (!sk[126]) & (g1340) & (!g1065)) + ((!g1128) & (!g1028) & (!sk[126]) & (g1340) & (g1065)) + ((!g1128) & (!g1028) & (sk[126]) & (!g1340) & (g1065)) + ((!g1128) & (!g1028) & (sk[126]) & (g1340) & (!g1065)) + ((!g1128) & (g1028) & (!sk[126]) & (!g1340) & (!g1065)) + ((!g1128) & (g1028) & (!sk[126]) & (!g1340) & (g1065)) + ((!g1128) & (g1028) & (!sk[126]) & (g1340) & (!g1065)) + ((!g1128) & (g1028) & (!sk[126]) & (g1340) & (g1065)) + ((!g1128) & (g1028) & (sk[126]) & (!g1340) & (!g1065)) + ((!g1128) & (g1028) & (sk[126]) & (g1340) & (g1065)) + ((g1128) & (!g1028) & (!sk[126]) & (g1340) & (!g1065)) + ((g1128) & (!g1028) & (!sk[126]) & (g1340) & (g1065)) + ((g1128) & (!g1028) & (sk[126]) & (!g1340) & (!g1065)) + ((g1128) & (!g1028) & (sk[126]) & (g1340) & (g1065)) + ((g1128) & (g1028) & (!sk[126]) & (!g1340) & (!g1065)) + ((g1128) & (g1028) & (!sk[126]) & (!g1340) & (g1065)) + ((g1128) & (g1028) & (!sk[126]) & (g1340) & (!g1065)) + ((g1128) & (g1028) & (!sk[126]) & (g1340) & (g1065)) + ((g1128) & (g1028) & (sk[126]) & (!g1340) & (g1065)) + ((g1128) & (g1028) & (sk[126]) & (g1340) & (!g1065)));
	assign g2066 = (((!g1339) & (!sk[127]) & (g1065)) + ((!g1339) & (sk[127]) & (g1065)) + ((g1339) & (!sk[127]) & (g1065)) + ((g1339) & (sk[127]) & (!g1065)));
	assign g2067 = (((!g1128) & (!g1028) & (!g1340) & (sk[0]) & (!g1065)) + ((!g1128) & (!g1028) & (g1340) & (!sk[0]) & (!g1065)) + ((!g1128) & (!g1028) & (g1340) & (!sk[0]) & (g1065)) + ((!g1128) & (!g1028) & (g1340) & (sk[0]) & (g1065)) + ((!g1128) & (g1028) & (!g1340) & (!sk[0]) & (!g1065)) + ((!g1128) & (g1028) & (!g1340) & (!sk[0]) & (g1065)) + ((!g1128) & (g1028) & (!g1340) & (sk[0]) & (g1065)) + ((!g1128) & (g1028) & (g1340) & (!sk[0]) & (!g1065)) + ((!g1128) & (g1028) & (g1340) & (!sk[0]) & (g1065)) + ((!g1128) & (g1028) & (g1340) & (sk[0]) & (!g1065)) + ((g1128) & (!g1028) & (!g1340) & (sk[0]) & (g1065)) + ((g1128) & (!g1028) & (g1340) & (!sk[0]) & (!g1065)) + ((g1128) & (!g1028) & (g1340) & (!sk[0]) & (g1065)) + ((g1128) & (!g1028) & (g1340) & (sk[0]) & (!g1065)) + ((g1128) & (g1028) & (!g1340) & (!sk[0]) & (!g1065)) + ((g1128) & (g1028) & (!g1340) & (!sk[0]) & (g1065)) + ((g1128) & (g1028) & (!g1340) & (sk[0]) & (!g1065)) + ((g1128) & (g1028) & (g1340) & (!sk[0]) & (!g1065)) + ((g1128) & (g1028) & (g1340) & (!sk[0]) & (g1065)) + ((g1128) & (g1028) & (g1340) & (sk[0]) & (g1065)));
	assign g2068 = (((!g1339) & (!sk[1]) & (g1065)) + ((!g1339) & (sk[1]) & (g1065)) + ((g1339) & (!sk[1]) & (g1065)) + ((g1339) & (sk[1]) & (!g1065)));
	assign g2069 = (((!g2070) & (!sk[2]) & (g2071)) + ((!g2070) & (sk[2]) & (!g2071)) + ((g2070) & (!sk[2]) & (g2071)));
	assign g2070 = (((!g417) & (!sk[3]) & (g2072)) + ((!g417) & (sk[3]) & (g2072)) + ((g417) & (!sk[3]) & (g2072)));
	assign g2071 = (((!sk[4]) & (!g417) & (g2075)) + ((!sk[4]) & (g417) & (g2075)) + ((sk[4]) & (g417) & (g2075)));
	assign g2072 = (((!g2073) & (!sk[5]) & (g2074)) + ((!g2073) & (sk[5]) & (!g2074)) + ((g2073) & (!sk[5]) & (g2074)));
	assign g2073 = (((!sk[6]) & (!g1163) & (g2078)) + ((!sk[6]) & (g1163) & (g2078)) + ((sk[6]) & (!g1163) & (g2078)));
	assign g2074 = (((!sk[7]) & (!g1163) & (g2079)) + ((!sk[7]) & (g1163) & (g2079)) + ((sk[7]) & (g1163) & (g2079)));
	assign g2075 = (((!sk[8]) & (!g2076) & (g2077)) + ((!sk[8]) & (g2076) & (g2077)) + ((sk[8]) & (!g2076) & (!g2077)));
	assign g2076 = (((!g1163) & (!sk[9]) & (g2080)) + ((!g1163) & (sk[9]) & (g2080)) + ((g1163) & (!sk[9]) & (g2080)));
	assign g2077 = (((!sk[10]) & (!g1163) & (g2081)) + ((!sk[10]) & (g1163) & (g2081)) + ((sk[10]) & (g1163) & (g2081)));
	assign g2078 = (((!g616) & (!g452) & (!g1175) & (sk[11]) & (g425)) + ((!g616) & (!g452) & (g1175) & (!sk[11]) & (!g425)) + ((!g616) & (!g452) & (g1175) & (!sk[11]) & (g425)) + ((!g616) & (!g452) & (g1175) & (sk[11]) & (!g425)) + ((!g616) & (g452) & (!g1175) & (!sk[11]) & (!g425)) + ((!g616) & (g452) & (!g1175) & (!sk[11]) & (g425)) + ((!g616) & (g452) & (!g1175) & (sk[11]) & (!g425)) + ((!g616) & (g452) & (g1175) & (!sk[11]) & (!g425)) + ((!g616) & (g452) & (g1175) & (!sk[11]) & (g425)) + ((!g616) & (g452) & (g1175) & (sk[11]) & (g425)) + ((g616) & (!g452) & (!g1175) & (sk[11]) & (!g425)) + ((g616) & (!g452) & (g1175) & (!sk[11]) & (!g425)) + ((g616) & (!g452) & (g1175) & (!sk[11]) & (g425)) + ((g616) & (!g452) & (g1175) & (sk[11]) & (g425)) + ((g616) & (g452) & (!g1175) & (!sk[11]) & (!g425)) + ((g616) & (g452) & (!g1175) & (!sk[11]) & (g425)) + ((g616) & (g452) & (!g1175) & (sk[11]) & (g425)) + ((g616) & (g452) & (g1175) & (!sk[11]) & (!g425)) + ((g616) & (g452) & (g1175) & (!sk[11]) & (g425)) + ((g616) & (g452) & (g1175) & (sk[11]) & (!g425)));
	assign g2079 = (((!g1174) & (!sk[12]) & (g425)) + ((!g1174) & (sk[12]) & (g425)) + ((g1174) & (!sk[12]) & (g425)) + ((g1174) & (sk[12]) & (!g425)));
	assign g2080 = (((!g616) & (!g452) & (!g1175) & (sk[13]) & (!g425)) + ((!g616) & (!g452) & (g1175) & (!sk[13]) & (!g425)) + ((!g616) & (!g452) & (g1175) & (!sk[13]) & (g425)) + ((!g616) & (!g452) & (g1175) & (sk[13]) & (g425)) + ((!g616) & (g452) & (!g1175) & (!sk[13]) & (!g425)) + ((!g616) & (g452) & (!g1175) & (!sk[13]) & (g425)) + ((!g616) & (g452) & (!g1175) & (sk[13]) & (g425)) + ((!g616) & (g452) & (g1175) & (!sk[13]) & (!g425)) + ((!g616) & (g452) & (g1175) & (!sk[13]) & (g425)) + ((!g616) & (g452) & (g1175) & (sk[13]) & (!g425)) + ((g616) & (!g452) & (!g1175) & (sk[13]) & (g425)) + ((g616) & (!g452) & (g1175) & (!sk[13]) & (!g425)) + ((g616) & (!g452) & (g1175) & (!sk[13]) & (g425)) + ((g616) & (!g452) & (g1175) & (sk[13]) & (!g425)) + ((g616) & (g452) & (!g1175) & (!sk[13]) & (!g425)) + ((g616) & (g452) & (!g1175) & (!sk[13]) & (g425)) + ((g616) & (g452) & (!g1175) & (sk[13]) & (!g425)) + ((g616) & (g452) & (g1175) & (!sk[13]) & (!g425)) + ((g616) & (g452) & (g1175) & (!sk[13]) & (g425)) + ((g616) & (g452) & (g1175) & (sk[13]) & (g425)));
	assign g2081 = (((!g1174) & (!sk[14]) & (g425)) + ((!g1174) & (sk[14]) & (g425)) + ((g1174) & (!sk[14]) & (g425)) + ((g1174) & (sk[14]) & (!g425)));

endmodule