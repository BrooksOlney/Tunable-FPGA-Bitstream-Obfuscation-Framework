module pdc (
	i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, 
	i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, o_0_, o_1_, 
	o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, 
	o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, 
	o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, 
	o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_);

input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, i_14_, i_15_;

output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_;

wire n10, n247, n6, n5, n3, n7, n13, n11, n17, n16, n14, n21, n18, n24, n22, n25, n28, n34, n31, n35, n39, n37, n40, n45, n43, n46, n47, n49, n50, n51, n54, n55, n53, n61, n62, n63, n64, n66, n65, n70, n71, n73, n74, n75, n76, n77, n72, n79, n78, n80, n82, n81, n83, n86, n88, n87, n103, n105, n104, n108, n109, n112, n118, n119, n122, n124, n125, n131, n128, n135, n132, n139, n136, n140, n143, n146, n152, n150, n151, n154, n157, n158, n159, n160, n156, n164, n161, n166, n165, n167, n170, n172, n173, n178, n175, n176, n174, n181, n182, n180, n179, n185, n184, n183, n188, n187, n186, n191, n190, n189, n193, n192, n196, n195, n194, n200, n198, n197, n202, n201, n204, n203, n207, n206, n205, n209, n208, n211, n210, n216, n213, n214, n212, n217, n220, n224, n225, n226, n227, n228, n229, n230, n231, n223, n233, n234, n235, n236, n237, n238, n239, n240, n232, n244, n245, n243, n241, n248, n246, n251, n252, n254, n255, n256, n257, n258, n250, n260, n261, n262, n263, n259, n266, n264, n269, n270, n272, n273, n274, n275, n276, n268, n280, n277, n281, n283, n286, n284, n288, n289, n287, n291, n292, n293, n290, n295, n296, n294, n300, n301, n299, n304, n305, n306, n307, n308, n309, n303, n311, n312, n313, n310, n315, n316, n314, n319, n320, n318, n317, n321, n323, n324, n322, n327, n325, n332, n328, n334, n333, n337, n338, n336, n335, n340, n341, n342, n339, n344, n345, n343, n347, n346, n350, n348, n354, n351, n355, n357, n358, n356, n360, n359, n363, n364, n362, n367, n366, n370, n371, n369, n373, n374, n372, n378, n375, n380, n381, n379, n383, n384, n385, n386, n387, n388, n389, n390, n382, n392, n393, n394, n395, n396, n397, n398, n391, n400, n401, n399, n404, n405, n406, n407, n408, n409, n410, n403, n412, n413, n411, n415, n416, n417, n418, n419, n420, n421, n422, n414, n426, n423, n429, n430, n431, n432, n433, n434, n427, n436, n437, n438, n439, n440, n441, n442, n443, n435, n446, n445, n444, n449, n448, n447, n450, n452, n453, n451, n456, n457, n458, n459, n460, n461, n462, n454, n464, n465, n466, n467, n468, n463, n471, n470, n469, n472, n476, n474, n477, n479, n478, n481, n484, n486, n492, n491, n489, n495, n494, n493, n497, n496, n499, n501, n502, n503, n504, n505, n506, n507, n508, n500, n509, n511, n512, n513, n510, n516, n514, n518, n517, n521, n519, n525, n526, n524, n522, n528, n527, n531, n532, n530, n529, n534, n533, n536, n537, n535, n538, n542, n541, n540, n546, n547, n544, n545, n543, n549, n550, n551, n552, n553, n554, n548, n556, n557, n558, n559, n560, n561, n555, n563, n564, n565, n566, n567, n568, n562, n569, n573, n572, n578, n576, n575, n582, n580, n581, n579, n583, n588, n589, n590, n591, n592, n593, n587, n595, n596, n597, n598, n599, n600, n601, n602, n594, n604, n603, n606, n605, n609, n608, n607, n611, n612, n610, n613, n614, n616, n615, n619, n620, n621, n622, n623, n624, n625, n626, n618, n627, n630, n634, n635, n636, n637, n638, n639, n633, n642, n641, n640, n643, n646, n647, n645, n644, n649, n650, n648, n653, n654, n652, n651, n656, n657, n655, n660, n659, n658, n662, n663, n661, n666, n667, n665, n664, n669, n670, n668, n672, n673, n671, n675, n674, n678, n679, n677, n676, n681, n680, n683, n682, n686, n687, n688, n689, n690, n691, n692, n693, n685, n695, n696, n694, n700, n697, n702, n701, n704, n705, n706, n707, n703, n709, n710, n711, n708, n712, n714, n715, n713, n716, n718, n719, n720, n721, n722, n723, n724, n717, n728, n726, n727, n725, n730, n729, n732, n734, n733, n737, n736, n739, n740, n738, n742, n743, n741, n744, n747, n748, n750, n753, n754, n755, n752, n757, n758, n759, n760, n761, n762, n763, n764, n756, n766, n765, n768, n767, n772, n773, n771, n769, n776, n775, n774, n779, n780, n778, n777, n782, n783, n784, n785, n786, n781, n789, n788, n787, n791, n790, n793, n794, n792, n795, n796, n799, n800, n797, n802, n803, n804, n805, n806, n807, n808, n801, n810, n809, n813, n812, n811, n816, n815, n814, n819, n817, n821, n820, n823, n824, n822, n826, n827, n828, n829, n830, n825, n832, n833, n831, n834, n837, n836, n840, n839, n838, n842, n841, n844, n845, n846, n847, n843, n849, n850, n848, n852, n851, n855, n856, n854, n853, n857, n859, n862, n864, n863, n866, n869, n870, n871, n872, n873, n868, n875, n876, n877, n878, n874, n879, n882, n884, n889, n887, n886, n893, n892, n890, n894, n897, n896, n901, n900, n899, n903, n904, n905, n906, n902, n908, n907, n910, n911, n912, n913, n909, n915, n916, n914, n918, n917, n919, n921, n920, n923, n924, n922, n926, n927, n928, n929, n925, n931, n932, n933, n934, n935, n936, n937, n930, n939, n940, n941, n938, n945, n942, n947, n948, n946, n951, n950, n949, n953, n952, n954, n955, n959, n960, n958, n962, n963, n961, n965, n964, n968, n967, n966, n970, n969, n972, n973, n971, n976, n977, n978, n979, n982, n980, n981, n984, n983, n987, n988, n985, n990, n991, n989, n993, n994, n992, n995, n996, n997, n1002, n1003, n1001, n1004, n1005, n1007, n1006, n1010, n1009, n1013, n1012, n1011, n1016, n1019, n1021, n1020, n1023, n1024, n1025, n1026, n1027, n1028, n1022, n1030, n1029, n1033, n1031, n1035, n1034, n1037, n1038, n1039, n1040, n1036, n1041, n1043, n1044, n1045, n1042, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1046, n1056, n1057, n1055, n1059, n1060, n1061, n1062, n1058, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1071, n1070, n1073, n1075, n1076, n1077, n1074, n1080, n1078, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1081, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1089, n1099, n1100, n1101, n1102, n1103, n1104, n1098, n1106, n1105, n1108, n1109, n1110, n1111, n1112, n1113, n1107, n1115, n1114, n1117, n1118, n1116, n1120, n1121, n1122, n1123, n1119, n1125, n1126, n1127, n1128, n1129, n1124, n1130, n1136, n1133, n1138, n1139, n1137, n1141, n1140, n1142, n1145, n1144, n1148, n1149, n1150, n1146, n1151, n1153, n1154, n1155, n1156, n1157, n1158, n1152, n1159, n1163, n1164, n1162, n1165, n1168, n1169, n1172, n1174, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1176, n1184, n1187, n1188, n1186, n1185, n1191, n1189, n1193, n1194, n1195, n1196, n1192, n1198, n1199, n1200, n1201, n1202, n1197, n1204, n1203, n1206, n1205, n1207, n1208, n1212, n1210, n1209, n1214, n1215, n1213, n1217, n1218, n1219, n1220, n1216, n1222, n1221, n1226, n1224, n1227, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1228, n1237, n1236, n1239, n1238, n1240, n1242, n1243, n1244, n1245, n1246, n1241, n1248, n1247, n1250, n1251, n1249, n1253, n1252, n1254, n1257, n1258, n1256, n1260, n1259, n1262, n1261, n1264, n1265, n1263, n1266, n1269, n1270, n1271, n1272, n1268, n1274, n1275, n1276, n1277, n1273, n1279, n1280, n1278, n1282, n1283, n1284, n1285, n1286, n1287, n1281, n1289, n1290, n1291, n1292, n1288, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1293, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1301, n1311, n1314, n1315, n1316, n1319, n1321, n1323, n1322, n1325, n1326, n1327, n1329, n1330, n1331, n1332, n1328, n1336, n1337, n1339, n1341, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1351, n1352, n1353, n1354, n1350, n1355, n1356, n1357, n1359, n1361, n1362, n1364, n1363, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1384, n1385, n1388, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1400, n1401, n1402, n1403, n1404, n1399, n1406, n1407, n1405, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1411, n1420, n1421, n1422, n1419, n1423, n1424, n1425, n1426, n1427, n1428, n1431, n1432, n1433, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1452, n1453, n1454, n1455, n1451, n1457, n1459, n1460, n1461, n1462, n1464, n1465, n1466, n1463, n1468, n1469, n1470, n1467, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1482, n1483, n1481, n1484, n1485, n1486, n1487, n1488, n1490, n1491, n1492, n1493, n1495, n1496, n1498, n1499, n1500, n1502, n1503, n1504, n1505, n1501, n1506, n1507, n1508, n1509, n1510, n1511, n1513, n1514, n1515, n1516, n1512, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1531, n1532, n1533, n1530, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1543, n1542, n1545, n1544, n1547, n1546, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1556, n1558, n1555, n1560, n1561, n1559, n1562, n1563, n1564, n1565, n1567, n1566, n1569, n1568, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1578, n1579, n1581, n1577, n1583, n1584, n1585, n1586, n1582, n1588, n1587, n1589, n1592, n1593, n1594, n1591, n1596, n1598, n1599, n1600, n1597, n1601, n1602, n1603, n1604, n1605, n1608, n1606, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1630, n1631, n1632, n1633, n1634, n1629, n1635, n1637, n1638, n1639, n1640, n1641, n1642, n1644, n1645, n1646, n1647, n1648, n1643, n1649, n1650, n1651, n1653, n1654, n1655, n1656, n1657, n1652, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1666, n1667, n1668, n1665, n1671, n1669, n1673, n1674, n1672, n1677, n1678, n1679, n1680, n1676, n1682, n1683, n1684, n1685, n1686, n1681, n1688, n1689, n1690, n1691, n1687, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1709, n1710, n1708, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1719, n1720, n1721, n1722, n1723, n1718, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1724, n1733, n1734, n1735, n1736, n1738, n1739, n1740, n1741, n1742, n1737, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1743, n1752, n1751, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1753, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1771, n1770, n1772, n1774, n1776, n1777, n1775, n1779, n1780, n1778, n1783, n1781, n1784, n1786, n1785, n1788, n1787, n1790, n1791, n1792, n1789, n1793, n1794, n1796, n1795, n1797, n1799, n1798, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1809, n1810, n1811, n1812, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1826, n1827, n1828, n1825, n1830, n1831, n1832, n1833, n1829, n1834, n1835, n1836, n1838, n1839, n1840, n1841, n1842, n1837, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1873, n1874, n1876, n1877, n1878, n1879, n1880, n1872, n1881, n1883, n1884, n1885, n1882, n1887, n1888, n1889, n1886, n1890, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1916, n1915, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1917, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1925, n1934, n1935, n1936, n1937, n1938, n1939, n1933, n1941, n1942, n1943, n1940, n1945, n1947, n1948, n1944, n1950, n1951, n1949, n1953, n1954, n1955, n1952, n1956, n1957, n1958, n1960, n1962, n1964, n1965, n1959, n1967, n1966, n1969, n1970, n1971, n1968, n1975, n1976, n1977, n1972, n1978, n1979, n1980, n1981, n1983, n1984, n1986, n1987, n1989, n1991, n1985, n1992, n1994, n1995, n1996, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2009, n2010, n2011, n2012, n2014, n2015, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2028, n2027, n2030, n2031, n2032, n2029, n2034, n2035, n2033, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2064, n2065, n2067, n2066, n2068, n2070, n2071, n2069, n2072, n2073, n2075, n2076, n2077, n2078, n2079, n2074, n2080, n2081, n2082, n2083, n2084, n2085, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2103, n2102, n2105, n2106, n2108, n2107, n2109, n2110, n2112, n2113, n2114, n2115, n2116, n2111, n2118, n2119, n2117, n2121, n2120, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2139, n2138, n2141, n2140, n2143, n2142, n2144, n2145, n2146, n2148, n2150, n2151, n2149, n2152, n2157, n2159, n2161, n2163, n2164, n2168, n2169, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2182, n2184, n2185, n2183, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2197, n2196, n2198, n2199, n2200, n2201, n2203, n2204, n2205, n2202, n2207, n2208, n2206, n2209, n2210, n2215, n2216, n2217, n2218, n2221, n2224, n2225, n2226, n2228, n2227, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2239, n2240, n2238, n2242, n2243, n2241, n2244, n2245, n2247, n2248, n2246, n2249, n2251, n2250, n2252, n2253, n2254, n2256, n2257, n2255, n2259, n2260, n2261, n2258, n2263, n2264, n2265, n2262, n2266, n2268, n2269, n2267, n2270, n2271, n2274, n2272, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2284, n2285, n2286, n2283, n2287, n2288, n2290, n2291, n2292, n2289, n2293, n2294, n2295, n2297, n2298, n2296, n2299, n2300, n2301, n2302, n2304, n2303, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2313, n2314, n2315, n2317, n2318, n2319, n2320, n2321, n2323, n2324, n2322, n2325, n2326, n2327, n2329, n2330, n2331, n2328, n2332, n2334, n2335, n2336, n2337, n2333, n2338, n2339, n2340, n2341, n2343, n2347, n2344, n2348, n2349, n2350, n2351, n2353, n2352, n2355, n2356, n2357, n2354, n2359, n2360, n2361, n2358, n2363, n2364, n2365, n2362, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2378, n2379, n2380, n2381, n2383, n2384, n2385, n2382, n2386, n2387, n2388, n2389, n2390, n2392, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2403, n2404, n2402, n2406, n2405, n2407, n2408, n2410, n2411, n2412, n2413, n2415, n2416, n2417, n2418, n2420, n2422, n2423, n2424, n2425, n2426, n2427, n2429, n2431, n2432, n2433, n2434, n2435, n2436, n2438, n2439, n2441, n2437, n2442, n2443, n2445, n2444, n2448, n2449, n2447, n2450, n2451, n2453, n2455, n2457, n2460, n2459, n2461, n2462, n2463, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2479, n2478, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2494, n2495, n2496, n2497, n2500, n2502, n2501, n2504, n2505, n2506, n2509, n2510, n2512, n2511, n2513, n2515, n2514, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2526, n2525, n2528, n2529, n2530, n2531, n2534, n2535, n2536, n2539, n2540, n2541, n2543, n2544, n2547, n2546, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2562, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2591, n2590, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618;

assign o_0_ = ( n50  &  (~ n54) ) | ( (~ n54)  &  n124 ) ;
 assign o_1_ = ( (~ n54)  &  n122 ) | ( (~ n54)  &  (~ n1137) ) | ( (~ n54)  &  (~ n1766) ) ;
 assign o_2_ = ( (~ n54)  &  n118 ) | ( (~ n54)  &  n119 ) | ( (~ n54)  &  (~ n769) ) ;
 assign o_3_ = ( (~ n54)  &  (~ n2483) ) | ( (~ n54)  &  (~ n2488) ) ;
 assign o_4_ = ( (~ n54)  &  (~ n2462) ) | ( (~ n54)  &  (~ n2472) ) | ( (~ n54)  &  (~ n2474) ) ;
 assign o_5_ = ( (~ n2617) ) ;
 assign o_6_ = ( (~ n112) ) ;
 assign o_7_ = ( (~ n54)  &  n109 ) | ( (~ n54)  &  (~ n1511) ) | ( (~ n54)  &  (~ n1512) ) ;
 assign o_8_ = ( (~ n2616) ) ;
 assign o_9_ = ( (~ n54)  &  n108 ) | ( (~ n54)  &  (~ n2175) ) | ( (~ n54)  &  (~ n2177) ) ;
 assign o_10_ = ( (~ n104) ) ;
 assign o_11_ = ( (~ n1081) ) ;
 assign o_12_ = ( (~ n1293) ) ;
 assign o_13_ = ( (~ n1281) ) ;
 assign o_14_ = ( (~ n1499) ) ;
 assign o_15_ = ( (~ n103) ) ;
 assign o_16_ = ( (~ n54)  &  (~ n2596) ) | ( (~ n54)  &  (~ n2598) ) | ( (~ n54)  &  (~ n2600) ) ;
 assign o_17_ = ( (~ n54)  &  (~ n2584) ) | ( (~ n54)  &  (~ n2586) ) | ( (~ n54)  &  (~ n2588) ) ;
 assign o_18_ = ( (~ n54)  &  (~ n2569) ) | ( (~ n54)  &  (~ n2571) ) | ( (~ n54)  &  (~ n2573) ) ;
 assign o_19_ = ( (~ n54)  &  (~ n2553) ) | ( (~ n54)  &  (~ n2554) ) | ( (~ n54)  &  (~ n2555) ) ;
 assign o_20_ = ( (~ n54)  &  (~ n2531) ) | ( (~ n54)  &  (~ n2535) ) ;
 assign o_21_ = ( (~ n87) ) ;
 assign o_22_ = ( n83 ) | ( n86 ) | ( (~ n1011) ) | ( (~ n1579) ) ;
 assign o_23_ = ( (~ n81) ) ;
 assign o_24_ = ( (~ n80) ) ;
 assign o_25_ = ( (~ n78) ) ;
 assign o_26_ = ( (~ n72) ) ;
 assign o_27_ = ( (~ n54)  &  n70  &  n71 ) ;
 assign o_28_ = ( (~ n2615) ) ;
 assign o_29_ = ( (~ n54)  &  (~ n938) ) | ( (~ n54)  &  (~ n2511) ) | ( (~ n54)  &  (~ n2513) ) ;
 assign o_30_ = ( (~ n65) ) ;
 assign o_31_ = ( n62 ) | ( n63 ) | ( n64 ) ;
 assign o_32_ = ( (~ n61) ) ;
 assign o_33_ = ( (~ n2614) ) ;
 assign o_34_ = ( (~ n54)  &  (~ n2506) ) | ( (~ n54)  &  (~ n2510) ) ;
 assign o_35_ = ( (~ n54)  &  (~ n1775) ) | ( (~ n54)  &  (~ n1778) ) | ( (~ n54)  &  (~ n2504) ) ;
 assign o_36_ = ( (~ n53) ) ;
 assign o_37_ = ( n49  &  (~ n54) ) | ( n50  &  (~ n54) ) | ( n51  &  (~ n54) ) ;
 assign o_38_ = ( n46  &  (~ n1380) ) ;
 assign o_39_ = ( n46  &  n47 ) ;
 assign n10 = ( n1368  &  n1397 ) ;
 assign n247 = ( n1368  &  n158 ) ;
 assign n6 = ( n1355  &  n1368 ) ;
 assign n5 = ( (~ n380) ) | ( (~ n1519) ) ;
 assign n3 = ( n6  &  n5 ) | ( n6  &  (~ n665) ) ;
 assign n7 = ( n10  &  (~ n608) ) | ( n10  &  (~ n1012) ) ;
 assign n13 = ( (~ n665) ) | ( (~ n1290) ) ;
 assign n11 = ( n10  &  n13 ) | ( n10  &  (~ n380) ) ;
 assign n17 = ( n1381  &  n1388 ) ;
 assign n16 = ( (~ n645) ) | ( (~ n1523) ) ;
 assign n14 = ( n17  &  n16 ) | ( n17  &  (~ n537) ) ;
 assign n21 = ( n1388  &  n1397 ) ;
 assign n18 = ( n21  &  (~ n347) ) | ( n21  &  (~ n1477) ) ;
 assign n24 = ( (~ n312) ) | ( (~ n706) ) ;
 assign n22 = ( n21  &  n24 ) | ( n21  &  (~ n740) ) ;
 assign n25 = ( n21  &  (~ n448) ) | ( n21  &  (~ n1524) ) ;
 assign n28 = ( n21  &  (~ n839) ) | ( n21  &  (~ n1956) ) ;
 assign n34 = ( (~ n1339)  &  n1388 ) ;
 assign n31 = ( n34  &  (~ n1473) ) | ( n34  &  (~ n1565) ) ;
 assign n35 = ( n34  &  (~ n837) ) | ( n34  &  (~ n1956) ) ;
 assign n39 = ( n1355  &  n1359 ) ;
 assign n37 = ( n39  &  (~ n706) ) | ( n39  &  (~ n1524) ) ;
 assign n40 = ( n34  &  (~ n263) ) | ( n34  &  (~ n1289) ) ;
 assign n45 = ( (~ n213) ) | ( (~ n921) ) ;
 assign n43 = ( n39  &  n45 ) | ( n39  &  (~ n506) ) ;
 assign n46 = ( n152  &  n150 ) | ( n152  &  n151 ) ;
 assign n47 = ( i_6_  &  (~ i_7_) ) ;
 assign n49 = ( n159  &  n1355 ) ;
 assign n50 = ( n119 ) | ( (~ n769) ) | ( (~ n1511) ) | ( (~ n1512) ) ;
 assign n51 = ( n1803 ) | ( n774 ) | ( n2489 ) ;
 assign n54 = ( (~ n112) ) | ( n154 ) | ( n156 ) | ( n161 ) | ( n165 ) | ( n167 ) | ( (~ n2179) ) | ( (~ n2180) ) ;
 assign n55 = ( n801  &  n886  &  n1010  &  n1770  &  n1772  &  (~ n2501) ) ;
 assign n53 = ( n54 ) | ( n55 ) ;
 assign n61 = ( (~ n71)  &  n976  &  n977 ) | ( n976  &  n977  &  (~ n1366) ) ;
 assign n62 = ( (~ n516)  &  n978 ) | ( (~ n516)  &  n979 ) ;
 assign n63 = ( n982  &  n980 ) | ( n982  &  n981 ) ;
 assign n64 = ( n1802 ) | ( n1803 ) ;
 assign n66 = ( (~ n119)  &  n489  &  n939  &  n976  &  n987  &  n1511  &  n1804  &  n2182 ) ;
 assign n65 = ( n54 ) | ( n66 ) ;
 assign n70 = ( i_0_  &  i_1_  &  (~ i_2_) ) ;
 assign n71 = ( i_6_  &  i_7_ ) ;
 assign n73 = ( n990 ) | ( n839 ) ;
 assign n74 = ( n1002  &  n1003  &  n1001 ) | ( n1002  &  n1003  &  n994 ) ;
 assign n75 = ( (~ n997)  &  n1806  &  n1807  &  n1809  &  n1810  &  n1811 ) ;
 assign n76 = ( (~ n995)  &  n996  &  n1812  &  n1814  &  n1815  &  n1816 ) ;
 assign n77 = ( (~ n146)  &  n989  &  n992  &  n1817  &  n1818  &  n1819 ) ;
 assign n72 = ( n73  &  n74  &  n75  &  n76  &  n77 ) ;
 assign n79 = ( n808  &  n807  &  n1606  &  n797  &  n889  &  n1770  &  n1004  &  n2516 ) ;
 assign n78 = ( n54 ) | ( n79 ) ;
 assign n80 = ( (~ n124)  &  n1010 ) | ( n1010  &  n1009 ) ;
 assign n82 = ( n1775  &  n930  &  n966  &  n781  &  n886  &  n801 ) ;
 assign n81 = ( n54 ) | ( n82 ) ;
 assign n83 = ( n1019  &  (~ n1077) ) | ( n1019  &  (~ n1253) ) ;
 assign n86 = ( (~ n730)  &  n1016 ) | ( n1016  &  (~ n1821) ) ;
 assign n88 = ( n1063  &  n1064  &  n1065  &  n1066  &  n1022  &  n1067  &  n1068  &  n1069 ) ;
 assign n87 = ( n54 ) | ( n88 ) ;
 assign n103 = ( (~ i_0_)  &  n172 ) | ( i_1_  &  n172 ) | ( i_2_  &  n172 ) ;
 assign n105 = ( n1770  &  n1772  &  n1687  &  n825  &  n1800  &  n1011  &  n2029 ) ;
 assign n104 = ( n54 ) | ( n105 ) ;
 assign n108 = ( n359 ) | ( n362 ) | ( n366 ) | ( n369 ) | ( (~ n372) ) | ( n2152 ) | ( (~ n2157) ) | ( (~ n2164) ) ;
 assign n109 = ( n1337  &  (~ n1339) ) ;
 assign n112 = ( (~ i_3_)  &  n172 ) | ( n170  &  n172 ) | ( (~ i_3_)  &  n173 ) | ( n170  &  n173 ) ;
 assign n118 = ( n1337  &  n157 ) ;
 assign n119 = ( n1341  &  (~ n1499) ) ;
 assign n122 = ( (~ n516)  &  (~ n1363) ) ;
 assign n124 = ( n118 ) | ( n109 ) ;
 assign n125 = ( n6  &  (~ n381) ) | ( n6  &  (~ n530) ) ;
 assign n131 = ( n1368  &  n1381 ) ;
 assign n128 = ( n131  &  (~ n204) ) | ( n131  &  (~ n323) ) ;
 assign n135 = ( (~ n1362)  &  n1382 ) ;
 assign n132 = ( n135  &  (~ n707) ) | ( n135  &  (~ n1106) ) ;
 assign n139 = ( n157  &  n1359 ) ;
 assign n136 = ( n139  &  (~ n1290) ) | ( n139  &  (~ n1519) ) ;
 assign n140 = ( n21  &  (~ n340) ) | ( n21  &  (~ n1563) ) ;
 assign n143 = ( n139  &  (~ n768) ) | ( n139  &  (~ n1478) ) ;
 assign n146 = ( (~ n959)  &  (~ n990) ) | ( (~ n990)  &  (~ n1071) ) ;
 assign n152 = ( (~ i_0_)  &  i_1_  &  (~ i_2_) ) ;
 assign n150 = ( i_5_  &  i_4_  &  i_3_ ) ;
 assign n151 = ( i_3_  &  i_4_  &  (~ i_5_) ) ;
 assign n154 = ( n109  &  (~ n2618) ) | ( n118  &  (~ n2618) ) ;
 assign n157 = ( n47  &  i_8_ ) ;
 assign n158 = ( i_8_  &  n71 ) ;
 assign n159 = ( n152  &  n1341 ) ;
 assign n160 = ( n152  &  n1343 ) ;
 assign n156 = ( n157  &  n159 ) | ( n158  &  n159 ) | ( n157  &  n160 ) | ( n158  &  n160 ) ;
 assign n164 = ( n1355  &  n160 ) ;
 assign n161 = ( n49  &  (~ n1350) ) | ( n164  &  (~ n1350) ) | ( n49  &  (~ n2178) ) | ( n164  &  (~ n2178) ) ;
 assign n166 = ( i_3_ ) | ( (~ n1336) ) | ( n1343 ) | ( (~ n1356) ) ;
 assign n165 = ( n70  &  n166 ) ;
 assign n167 = ( (~ n1350)  &  (~ n1363) ) | ( i_12_  &  (~ n1035)  &  (~ n1363) ) ;
 assign n170 = ( i_1_ ) | ( i_2_ ) | ( i_0_ ) ;
 assign n172 = ( i_0_ ) | ( (~ i_2_) ) ;
 assign n173 = ( i_1_ ) | ( (~ i_3_) ) ;
 assign n178 = ( (~ n6) ) | ( n323 ) ;
 assign n175 = ( n1369 ) | ( n1374 ) ;
 assign n176 = ( n1369 ) | ( n1372 ) ;
 assign n174 = ( (~ n6)  &  n178 ) | ( n178  &  n175  &  n176 ) ;
 assign n181 = ( (~ n6) ) | ( n324 ) ;
 assign n182 = ( (~ n6) ) | ( n291 ) ;
 assign n180 = ( n1374 ) | ( n1393 ) ;
 assign n179 = ( (~ n6)  &  n181  &  n182 ) | ( n181  &  n182  &  n180 ) ;
 assign n185 = ( (~ n6) ) | ( n1071 ) ;
 assign n184 = ( n261  &  n1329 ) ;
 assign n183 = ( (~ n6)  &  n185 ) | ( n185  &  n184 ) ;
 assign n188 = ( (~ n6) ) | ( n1215 ) ;
 assign n187 = ( n340  &  n468 ) ;
 assign n186 = ( (~ n6)  &  n188 ) | ( n188  &  n187 ) ;
 assign n191 = ( (~ n6) ) | ( n1395 ) ;
 assign n190 = ( n1367 ) | ( n1374 ) ;
 assign n189 = ( (~ n6)  &  n191 ) | ( n191  &  n190 ) ;
 assign n193 = ( n1315 ) | ( n1396 ) ;
 assign n192 = ( (~ n6)  &  n189 ) | ( n189  &  n193 ) ;
 assign n196 = ( (~ n6) ) | ( n565 ) ;
 assign n195 = ( n341  &  n466 ) ;
 assign n194 = ( (~ n6)  &  n196 ) | ( n196  &  n195 ) ;
 assign n200 = ( (~ n247) ) | ( n288 ) ;
 assign n198 = ( n318  &  n213 ) ;
 assign n197 = ( (~ n247)  &  n200 ) | ( n200  &  n198 ) ;
 assign n202 = ( (~ n247) ) | ( n176 ) ;
 assign n201 = ( (~ n247)  &  n202 ) | ( n175  &  n202 ) ;
 assign n204 = ( n1315 ) | ( n1327 ) ;
 assign n203 = ( (~ n247)  &  n201 ) | ( n201  &  n204 ) ;
 assign n207 = ( (~ n247) ) | ( n291 ) ;
 assign n206 = ( n180  &  n373 ) ;
 assign n205 = ( (~ n247)  &  n207 ) | ( n207  &  n206 ) ;
 assign n209 = ( (~ n247) ) | ( n1215 ) ;
 assign n208 = ( (~ n247)  &  n209 ) | ( n187  &  n209 ) ;
 assign n211 = ( (~ n247) ) | ( n565 ) ;
 assign n210 = ( (~ n247)  &  n211 ) | ( n195  &  n211 ) ;
 assign n216 = ( (~ n139) ) | ( n468 ) ;
 assign n213 = ( n1315 ) | ( n1321 ) ;
 assign n214 = ( n1344 ) | ( n1347 ) ;
 assign n212 = ( (~ n139)  &  n216 ) | ( n216  &  n213  &  n214 ) ;
 assign n217 = ( n34  &  (~ n342) ) | ( n34  &  (~ n345) ) ;
 assign n220 = ( n21  &  (~ n508) ) | ( n21  &  (~ n1329) ) ;
 assign n224 = ( (~ n10) ) | ( n204 ) ;
 assign n225 = ( (~ n10) ) | ( n243 ) ;
 assign n226 = ( (~ n10) ) | ( n323 ) ;
 assign n227 = ( (~ n10) ) | ( n1271 ) ;
 assign n228 = ( (~ n10) ) | ( n1377 ) ;
 assign n229 = ( n936  &  n903  &  n1700  &  n2106  &  n1626  &  n910 ) ;
 assign n230 = ( n1047  &  n2109  &  n1874  &  n1025  &  n1024  &  n1840  &  n2110  &  n2107 ) ;
 assign n231 = ( n2123  &  n2124  &  n2009  &  n2125  &  n2126  &  n2122  &  n2120  &  n2117 ) ;
 assign n223 = ( n224  &  n225  &  n226  &  n227  &  n228  &  n229  &  n230  &  n231 ) ;
 assign n233 = ( (~ n10) ) | ( n1376 ) ;
 assign n234 = ( (~ n10) ) | ( n190 ) ;
 assign n235 = ( (~ n10) ) | ( n180 ) ;
 assign n236 = ( (~ n280) ) | ( n665 ) ;
 assign n237 = ( (~ n10) ) | ( n261 ) ;
 assign n238 = ( (~ n280)  &  n2105 ) | ( n190  &  n313  &  n2105 ) ;
 assign n239 = ( (~ n266) ) | ( n2236 ) ;
 assign n240 = ( (~ n21)  &  n260 ) | ( n180  &  n260 ) | ( (~ n21)  &  n990 ) | ( n180  &  n990 ) ;
 assign n232 = ( n233  &  n234  &  n235  &  n236  &  n237  &  n238  &  n239  &  n240 ) ;
 assign n244 = ( (~ n139) ) | ( n323 ) ;
 assign n245 = ( (~ n10) ) | ( n324 ) ;
 assign n243 = ( n1347 ) | ( n1367 ) ;
 assign n241 = ( (~ n21)  &  n244  &  n245 ) | ( n244  &  n245  &  n243 ) ;
 assign n248 = ( n280 ) | ( n21 ) ;
 assign n246 = ( n247  &  (~ n815) ) | ( n248  &  (~ n815) ) ;
 assign n251 = ( (~ n10) ) | ( n342 ) ;
 assign n252 = ( (~ n34) ) | ( n1379 ) ;
 assign n254 = ( (~ n21)  &  (~ n683) ) | ( (~ n683)  &  n1433 ) | ( (~ n21)  &  n2039 ) | ( n1433  &  n2039 ) ;
 assign n255 = ( (~ n10)  &  (~ n247) ) | ( (~ n247)  &  n175 ) | ( (~ n10)  &  n810 ) | ( n175  &  n810 ) ;
 assign n256 = ( (~ n139)  &  n1009 ) | ( (~ n266)  &  n1009 ) | ( (~ n139)  &  n2148 ) | ( (~ n266)  &  n2148 ) ;
 assign n257 = ( n203  &  n205  &  n1154  &  n1419  &  n1411  &  n223  &  n232  &  n241 ) ;
 assign n258 = ( n2014  &  n1984  &  n1964  &  n2144  &  n2145  &  n2146  &  n2142  &  n2140 ) ;
 assign n250 = ( (~ n246)  &  n251  &  n252  &  n254  &  n255  &  n256  &  n257  &  n258 ) ;
 assign n260 = ( n180  &  n312 ) ;
 assign n261 = ( n1346 ) | ( n1374 ) ;
 assign n262 = ( (~ i_15_) ) | ( n1345 ) ;
 assign n263 = ( n1314 ) | ( n1325 ) ;
 assign n259 = ( n260  &  n261  &  n262  &  n263 ) ;
 assign n266 = ( (~ n175) ) | ( (~ n665) ) ;
 assign n264 = ( (~ n260)  &  (~ n336) ) | ( n266  &  (~ n336) ) ;
 assign n269 = ( (~ n139) ) | ( n652 ) ;
 assign n270 = ( (~ n139) ) | ( n190 ) ;
 assign n272 = ( n2100  &  n2101 ) | ( n2100  &  n318 ) ;
 assign n273 = ( (~ n21)  &  (~ n139) ) | ( (~ n21)  &  n341 ) | ( (~ n139)  &  n645 ) | ( n341  &  n645 ) ;
 assign n274 = ( (~ n363)  &  n2102 ) | ( n652  &  n2102 ) ;
 assign n275 = ( n1833  &  n1839  &  n1910  &  n1864  &  n1655  &  n1870 ) ;
 assign n276 = ( n1723  &  n1728  &  n1757  &  n1702  &  n2034  &  n1749 ) ;
 assign n268 = ( (~ n264)  &  n269  &  n270  &  n272  &  n273  &  n274  &  n275  &  n276 ) ;
 assign n280 = ( (~ n1339)  &  n1382 ) ;
 assign n277 = ( n280  &  (~ n288) ) | ( n280  &  (~ n291) ) ;
 assign n281 = ( n176 ) | ( (~ n370) ) ;
 assign n283 = ( n39  &  (~ n291) ) | ( n39  &  (~ n1071) ) ;
 assign n286 = ( n1215  &  n316 ) ;
 assign n284 = ( (~ n17) ) | ( n286 ) ;
 assign n288 = ( n1344 ) | ( n1372 ) ;
 assign n289 = ( (~ n17)  &  (~ n39) ) ;
 assign n287 = ( n288 ) | ( n289 ) ;
 assign n291 = ( n1372 ) | ( n1393 ) ;
 assign n292 = ( n1325 ) | ( n1367 ) ;
 assign n293 = ( n576  &  n1012  &  n176 ) ;
 assign n290 = ( n291  &  n292  &  n293 ) ;
 assign n295 = ( (~ n616)  &  n1428 ) ;
 assign n296 = ( (~ n400)  &  n1427 ) ;
 assign n294 = ( (~ n34)  &  (~ n131)  &  n295  &  n296 ) ;
 assign n300 = ( n34 ) | ( n616 ) ;
 assign n301 = ( n135 ) | ( n21 ) ;
 assign n299 = ( n139  &  (~ n726) ) | ( n300  &  (~ n726) ) | ( n301  &  (~ n726) ) ;
 assign n304 = ( (~ n283)  &  n284  &  n287  &  n1435  &  n1436  &  n1437  &  n1438  &  n1439 ) ;
 assign n305 = ( n606  &  n534  &  n609 ) ;
 assign n306 = ( (~ n21)  &  (~ n280) ) | ( (~ n21)  &  n292 ) | ( (~ n280)  &  n544 ) | ( n292  &  n544 ) ;
 assign n307 = ( (~ n10)  &  n296 ) | ( (~ n10)  &  n959 ) | ( n296  &  n1012 ) | ( n959  &  n1012 ) ;
 assign n308 = ( (~ n248)  &  n290 ) | ( (~ n248)  &  (~ n426) ) | ( n290  &  n1431 ) | ( (~ n426)  &  n1431 ) ;
 assign n309 = ( (~ n299)  &  n518  &  n604  &  n1543  &  n1545  &  n1547  &  n2084  &  n2085 ) ;
 assign n303 = ( n304  &  n305  &  n306  &  n307  &  n308  &  n309 ) ;
 assign n311 = ( n659  &  n652 ) ;
 assign n312 = ( n1325 ) | ( n1398 ) ;
 assign n313 = ( n1325 ) | ( n1396 ) ;
 assign n310 = ( n311  &  n312  &  n313  &  n263 ) ;
 assign n315 = ( n1329  &  n213 ) ;
 assign n316 = ( n1370 ) | ( n1372 ) ;
 assign n314 = ( n315  &  n316  &  n288  &  n193 ) ;
 assign n319 = ( (~ n6) ) | ( n214 ) ;
 assign n320 = ( (~ n6) ) | ( n288 ) ;
 assign n318 = ( n1344 ) | ( n1374 ) ;
 assign n317 = ( (~ n6)  &  n319  &  n320 ) | ( n319  &  n320  &  n318 ) ;
 assign n321 = ( (~ n6)  &  n317 ) | ( n213  &  n317 ) ;
 assign n323 = ( n1347 ) | ( n1369 ) ;
 assign n324 = ( n1347 ) | ( n1393 ) ;
 assign n322 = ( n323  &  n204  &  n324 ) ;
 assign n327 = ( n323  &  n508 ) ;
 assign n325 = ( (~ n135) ) | ( n327 ) ;
 assign n332 = ( n616 ) | ( n17 ) ;
 assign n328 = ( (~ n214)  &  n332 ) | ( n332  &  (~ n897) ) | ( n332  &  (~ n1271) ) ;
 assign n334 = ( (~ n135)  &  (~ n616) ) ;
 assign n333 = ( n324 ) | ( n334 ) ;
 assign n337 = ( n1440  &  n1441  &  n1442  &  n1443  &  n1444  &  n1445  &  n1446  &  n1447 ) ;
 assign n338 = ( n322  &  n525  &  n532 ) | ( (~ n426)  &  n525  &  n532 ) ;
 assign n336 = ( (~ n300)  &  n1426 ) ;
 assign n335 = ( n337  &  n338  &  n336 ) | ( n337  &  n338  &  n243 ) ;
 assign n340 = ( n1374 ) | ( n1378 ) ;
 assign n341 = ( n1374 ) | ( n1385 ) ;
 assign n342 = ( n1315 ) | ( n1385 ) ;
 assign n339 = ( n340  &  n341  &  n342 ) ;
 assign n344 = ( n1379  &  n345 ) ;
 assign n345 = ( n1315 ) | ( n1344 ) ;
 assign n343 = ( (~ n6)  &  n295 ) | ( (~ n6)  &  n344 ) | ( n295  &  n345 ) | ( n344  &  n345 ) ;
 assign n347 = ( n1376  &  n1377 ) ;
 assign n346 = ( n323  &  n190  &  n347 ) ;
 assign n350 = ( n357 ) | ( n371 ) ;
 assign n348 = ( n350  &  (~ n815) ) | ( n350  &  (~ n1009) ) ;
 assign n354 = ( n135 ) | ( (~ n295) ) ;
 assign n351 = ( n354  &  (~ n1007) ) | ( n354  &  (~ n1395) ) ;
 assign n355 = ( (~ n291)  &  n300 ) | ( n300  &  (~ n508) ) ;
 assign n357 = ( n426 ) | ( n131 ) ;
 assign n358 = ( (~ n336) ) | ( n363 ) ;
 assign n356 = ( n357  &  (~ n837) ) | ( n358  &  (~ n837) ) ;
 assign n360 = ( n426 ) | ( n135 ) ;
 assign n359 = ( n10  &  (~ n1379) ) | ( n360  &  (~ n1379) ) ;
 assign n363 = ( n6 ) | ( n247 ) ;
 assign n364 = ( n34 ) | ( (~ n295) ) ;
 assign n362 = ( (~ n262)  &  n363 ) | ( (~ n262)  &  n364 ) ;
 assign n367 = ( n400 ) | ( n358 ) | ( n378 ) ;
 assign n366 = ( n280  &  (~ n645) ) | ( n367  &  (~ n645) ) ;
 assign n370 = ( n1359  &  n158 ) ;
 assign n371 = ( n6 ) | ( (~ n336) ) ;
 assign n369 = ( (~ n204)  &  n370 ) | ( (~ n204)  &  n371 ) ;
 assign n373 = ( n1315 ) | ( n1398 ) ;
 assign n374 = ( (~ n6)  &  n1448 ) ;
 assign n372 = ( n373 ) | ( n374 ) ;
 assign n378 = ( n131 ) | ( n10 ) ;
 assign n375 = ( (~ n262)  &  n378 ) | ( n378  &  (~ n652) ) | ( n378  &  (~ n1450) ) ;
 assign n380 = ( n1327 ) | ( n1348 ) ;
 assign n381 = ( n1314 ) | ( n1374 ) ;
 assign n379 = ( n380  &  n381 ) ;
 assign n383 = ( (~ n247) ) | ( n530 ) ;
 assign n384 = ( (~ n247) ) | ( n611 ) ;
 assign n385 = ( (~ n10) ) | ( n470 ) ;
 assign n386 = ( (~ n10) ) | ( n448 ) ;
 assign n387 = ( (~ n10) ) | ( n743 ) ;
 assign n388 = ( n2276  &  n2277  &  n1859  &  n1759 ) ;
 assign n389 = ( n2278  &  n2279  &  n1092  &  n2280  &  n2281  &  n1879  &  n1039  &  n2282 ) ;
 assign n390 = ( n2037  &  n2288  &  n1101  &  n1110  &  n2019  &  n1198  &  n2287  &  n2283 ) ;
 assign n382 = ( n383  &  n384  &  n385  &  n386  &  n387  &  n388  &  n389  &  n390 ) ;
 assign n392 = ( (~ n39)  &  (~ n426) ) | ( (~ n39)  &  n470 ) | ( (~ n426)  &  n1250 ) | ( n470  &  n1250 ) ;
 assign n393 = ( n380  &  n2310 ) | ( (~ n400)  &  n2310 ) ;
 assign n394 = ( (~ n135)  &  n2309 ) | ( n448  &  n1474  &  n2309 ) ;
 assign n395 = ( n1187  &  n2308  &  n1244  &  n1243 ) ;
 assign n396 = ( n2305  &  n2306  &  n1991  &  n1947  &  n1976  &  n1002  &  n2307  &  n2303 ) ;
 assign n397 = ( n2299  &  n1845  &  n1855  &  n2300  &  n2301  &  n2302  &  n1867  &  n2296 ) ;
 assign n398 = ( n2293  &  n1720  &  n1729  &  n2294  &  n1680  &  n2295  &  n1635  &  n2289 ) ;
 assign n391 = ( n392  &  n382  &  n393  &  n394  &  n395  &  n396  &  n397  &  n398 ) ;
 assign n400 = ( n426 ) | ( n139 ) ;
 assign n401 = ( n131 ) | ( n21 ) ;
 assign n399 = ( n400  &  (~ n921) ) | ( n401  &  (~ n921) ) ;
 assign n404 = ( (~ n139) ) | ( n1474 ) ;
 assign n405 = ( (~ n139) ) | ( n743 ) ;
 assign n406 = ( (~ n280) ) | ( n1474 ) ;
 assign n407 = ( (~ n10) ) | ( n921 ) ;
 assign n408 = ( (~ n21)  &  n2311 ) | ( n448  &  n743  &  n2311 ) ;
 assign n409 = ( (~ n131)  &  (~ n139) ) | ( (~ n139)  &  n380 ) | ( (~ n131)  &  n448 ) | ( n380  &  n448 ) ;
 assign n410 = ( (~ n363)  &  n2313 ) | ( n1474  &  n2313 ) ;
 assign n403 = ( n404  &  n405  &  n406  &  n407  &  n408  &  n409  &  n391  &  n410 ) ;
 assign n412 = ( i_15_ ) | ( n1475 ) ;
 assign n413 = ( n1372 ) | ( n1390 ) ;
 assign n411 = ( n412  &  n413 ) ;
 assign n415 = ( (~ n17) ) | ( n465 ) ;
 assign n416 = ( (~ n17) ) | ( n413 ) ;
 assign n417 = ( (~ n248)  &  n411 ) | ( (~ n248)  &  n994 ) | ( n411  &  n1479 ) | ( n994  &  n1479 ) ;
 assign n418 = ( (~ n39)  &  n1481  &  n2271 ) | ( n465  &  n1481  &  n2271 ) ;
 assign n419 = ( n1907  &  n2270  &  n1906  &  n1969  &  n1094  &  n2267 ) ;
 assign n420 = ( n1912  &  n2000  &  n2266  &  n1986  &  n1948  &  n1937  &  n2262  &  n2258 ) ;
 assign n421 = ( n1868  &  n1843  &  n2252  &  n1852  &  n2253  &  n2254  &  n2250  &  n2249 ) ;
 assign n422 = ( n1662  &  n782  &  n793  &  n2244  &  n2245  &  n832  &  n2237  &  n2241 ) ;
 assign n414 = ( n415  &  n416  &  n417  &  n418  &  n419  &  n420  &  n421  &  n422 ) ;
 assign n426 = ( n1359  &  (~ n1361) ) ;
 assign n423 = ( n426  &  (~ n453) ) | ( n426  &  (~ n567) ) | ( n426  &  (~ n768) ) ;
 assign n429 = ( (~ n139) ) | ( n1477 ) ;
 assign n430 = ( (~ n280) ) | ( n413 ) ;
 assign n431 = ( (~ n10) ) | ( n465 ) ;
 assign n432 = ( (~ n280)  &  n2272 ) | ( n452  &  n2272 ) ;
 assign n433 = ( (~ n21)  &  (~ n139) ) | ( (~ n21)  &  n505 ) | ( (~ n139)  &  n1477 ) | ( n505  &  n1477 ) ;
 assign n434 = ( (~ n363)  &  n2275 ) | ( n413  &  n2275 ) ;
 assign n427 = ( n414  &  (~ n423)  &  n429  &  n430  &  n431  &  n432  &  n433  &  n434 ) ;
 assign n436 = ( (~ n21) ) | ( n1352 ) ;
 assign n437 = ( (~ n34) ) | ( n1265 ) ;
 assign n438 = ( (~ n34) ) | ( n1264 ) ;
 assign n439 = ( (~ n21) ) | ( n1484 ) ;
 assign n440 = ( n1084  &  n2236 ) | ( n1084  &  n1258 ) ;
 assign n441 = ( n1485  &  n1486  &  n1487  &  n1488 ) ;
 assign n442 = ( n2230  &  n2231  &  n2232  &  n2233  &  n2234  &  n1588  &  n2235  &  n1050 ) ;
 assign n443 = ( n1889  &  n845  &  n1651  &  n1622  &  n1885  &  n1567  &  n2229  &  n2227 ) ;
 assign n435 = ( n436  &  n437  &  n438  &  n439  &  n440  &  n441  &  n442  &  n443 ) ;
 assign n446 = ( (~ n10) ) | ( n1473 ) ;
 assign n445 = ( n1478  &  n1473 ) ;
 assign n444 = ( (~ n21)  &  n435  &  n446 ) | ( n435  &  n446  &  n445 ) ;
 assign n449 = ( (~ n247) ) | ( n505 ) ;
 assign n448 = ( n1374 ) | ( n1398 ) ;
 assign n447 = ( (~ n247)  &  n449 ) | ( n449  &  n448 ) ;
 assign n450 = ( (~ n247)  &  n447 ) | ( n373  &  n447 ) ;
 assign n452 = ( n768  &  n507 ) ;
 assign n453 = ( n1348 ) | ( n1369 ) ;
 assign n451 = ( n452  &  n453 ) ;
 assign n456 = ( (~ n21) ) | ( n505 ) ;
 assign n457 = ( (~ n21) ) | ( n1480 ) ;
 assign n458 = ( (~ n21) ) | ( n506 ) ;
 assign n459 = ( (~ n21)  &  n990 ) | ( n451  &  n990 ) | ( (~ n21)  &  n991 ) | ( n451  &  n991 ) ;
 assign n460 = ( (~ n280) ) | ( n465 ) ;
 assign n461 = ( n2189  &  n1083  &  n2190  &  n2191  &  n2192  &  n2193  &  n2194 ) ;
 assign n462 = ( n2186  &  n1709  &  n1760  &  n1755  &  n1873  &  n2187  &  n2188  &  n2183 ) ;
 assign n454 = ( (~ n143)  &  n456  &  n457  &  n458  &  n459  &  n460  &  n461  &  n462 ) ;
 assign n464 = ( n1347 ) | ( n1375 ) ;
 assign n465 = ( i_15_ ) | ( n1353 ) ;
 assign n466 = ( n1315 ) | ( n1391 ) ;
 assign n467 = ( n1352  &  n1191 ) ;
 assign n468 = ( n1315 ) | ( n1390 ) ;
 assign n463 = ( n315  &  n464  &  n373  &  n465  &  n193  &  n466  &  n467  &  n468 ) ;
 assign n471 = ( (~ n6) ) | ( n507 ) ;
 assign n470 = ( n1374 ) | ( n1396 ) ;
 assign n469 = ( (~ n6)  &  n471 ) | ( n471  &  n470 ) ;
 assign n472 = ( n247  &  n45 ) | ( n6  &  n45 ) | ( n247  &  (~ n193) ) | ( n6  &  (~ n193) ) ;
 assign n476 = ( (~ n204) ) | ( (~ n608) ) ;
 assign n474 = ( (~ n336)  &  n476 ) | ( (~ n336)  &  (~ n1491) ) ;
 assign n477 = ( n10  &  (~ n380) ) | ( n371  &  (~ n380) ) ;
 assign n479 = ( n131 ) | ( (~ n296) ) ;
 assign n478 = ( n17  &  (~ n1352) ) | ( n479  &  (~ n1352) ) ;
 assign n481 = ( (~ n295)  &  (~ n323) ) | ( (~ n295)  &  (~ n740) ) | ( (~ n295)  &  (~ n1492) ) ;
 assign n484 = ( (~ n336)  &  (~ n1258) ) | ( n378  &  (~ n1258) ) | ( n400  &  (~ n1258) ) ;
 assign n486 = ( (~ n296)  &  (~ n1265) ) | ( n354  &  (~ n1265) ) | ( n378  &  (~ n1265) ) ;
 assign n492 = ( n1357 ) | ( n1380 ) ;
 assign n491 = ( n1357 ) | ( n1362 ) ;
 assign n489 = ( n492  &  n491 ) | ( n492  &  (~ n892) ) ;
 assign n495 = ( n1780  &  n1776  &  n2182 ) ;
 assign n494 = ( n468  &  n544 ) ;
 assign n493 = ( n489  &  n495  &  n494 ) | ( n489  &  n495  &  n491 ) ;
 assign n497 = ( n466  &  n503 ) ;
 assign n496 = ( (~ n476)  &  n497 ) ;
 assign n499 = ( (~ n247)  &  (~ n6) ) | ( (~ n247)  &  n497 ) | ( (~ n6)  &  n496 ) | ( n497  &  n496 ) ;
 assign n501 = ( n413  &  n1474 ) ;
 assign n502 = ( n448  &  n921 ) ;
 assign n503 = ( n766  &  n709 ) ;
 assign n504 = ( n768  &  n381 ) ;
 assign n505 = ( n1372 ) | ( n1398 ) ;
 assign n506 = ( n1321 ) | ( n1372 ) ;
 assign n507 = ( n1372 ) | ( n1396 ) ;
 assign n508 = ( n1346 ) | ( n1347 ) ;
 assign n500 = ( n501  &  n502  &  n503  &  n504  &  n505  &  n506  &  n507  &  n508 ) ;
 assign n509 = ( n280  &  (~ n381) ) | ( (~ n381)  &  n400 ) ;
 assign n511 = ( n454  &  n450  &  n223  &  n828  &  n1506  &  n1507  &  n1508  &  n1509 ) ;
 assign n512 = ( n335  &  n241  &  n1501  &  n2320 ) ;
 assign n513 = ( n1532  &  n947  &  n915  &  n2314  &  n2317  &  n1139  &  n2315  &  n2318 ) ;
 assign n510 = ( n427  &  n444  &  n403  &  n493  &  n499  &  n511  &  n512  &  n513 ) ;
 assign n516 = ( i_10_ ) | ( i_9_ ) ;
 assign n514 = ( n516 ) | ( (~ n978) ) ;
 assign n518 = ( (~ n6) ) | ( n544 ) ;
 assign n517 = ( (~ n6)  &  n518 ) | ( n501  &  n518 ) ;
 assign n521 = ( (~ n10) ) | ( n214 ) ;
 assign n519 = ( (~ n5)  &  n521 ) | ( (~ n131)  &  n521 ) ;
 assign n525 = ( (~ n131) ) | ( n214 ) ;
 assign n526 = ( (~ n10) ) | ( n1518 ) ;
 assign n524 = ( n1348 ) | ( n1375 ) ;
 assign n522 = ( (~ n10)  &  n525  &  n526 ) | ( n525  &  n526  &  n524 ) ;
 assign n528 = ( (~ n131) ) | ( n1518 ) ;
 assign n527 = ( (~ n131)  &  n245  &  n528 ) | ( n245  &  n524  &  n528 ) ;
 assign n531 = ( (~ n10) ) | ( n1237 ) ;
 assign n532 = ( (~ n131) ) | ( n508 ) ;
 assign n530 = ( (~ i_15_) ) | ( n1351 ) ;
 assign n529 = ( (~ n10)  &  n531  &  n532 ) | ( n531  &  n532  &  n530 ) ;
 assign n534 = ( (~ n6) ) | ( n1431 ) ;
 assign n533 = ( (~ n6)  &  n534 ) | ( n503  &  n534 ) ;
 assign n536 = ( n1391 ) | ( n1517 ) ;
 assign n537 = ( n1348 ) | ( n1391 ) ;
 assign n535 = ( n536  &  n537 ) ;
 assign n538 = ( (~ n34)  &  n535 ) | ( n243  &  n535 ) | ( (~ n34)  &  (~ n616) ) | ( n243  &  (~ n616) ) ;
 assign n542 = ( (~ n10) ) | ( n292 ) ;
 assign n541 = ( n1367 ) | ( n1522 ) ;
 assign n540 = ( (~ n10)  &  n446  &  n542 ) | ( n446  &  n542  &  n541 ) ;
 assign n546 = ( n959 ) | ( n727 ) ;
 assign n547 = ( (~ n21) ) | ( n536 ) ;
 assign n544 = ( n1325 ) | ( n1378 ) ;
 assign n545 = ( n1362 ) | ( (~ n1368) ) ;
 assign n543 = ( n546  &  n547  &  n544 ) | ( n546  &  n547  &  n545 ) ;
 assign n549 = ( (~ n131) ) | ( n1521 ) ;
 assign n550 = ( (~ n131) ) | ( n568 ) ;
 assign n551 = ( (~ n6) ) | ( n1520 ) ;
 assign n552 = ( (~ n6) ) | ( n1043 ) ;
 assign n553 = ( (~ n1019)  &  n2394 ) | ( n1077  &  n2394 ) ;
 assign n554 = ( n953 ) | ( n545 ) ;
 assign n548 = ( n549  &  n550  &  n551  &  n552  &  n553  &  n554 ) ;
 assign n556 = ( n737  &  n541 ) ;
 assign n557 = ( n1523  &  n706 ) ;
 assign n558 = ( n1071  &  n1395 ) ;
 assign n559 = ( n1369 ) | ( n1517 ) ;
 assign n560 = ( n1367 ) | ( n1517 ) ;
 assign n561 = ( n1378 ) | ( n1522 ) ;
 assign n555 = ( n556  &  n557  &  n558  &  n559  &  n560  &  n561 ) ;
 assign n563 = ( n1012  &  n1290  &  n453 ) ;
 assign n564 = ( n1344 ) | ( n1522 ) ;
 assign n565 = ( n1372 ) | ( n1385 ) ;
 assign n566 = ( n1370 ) | ( n1522 ) ;
 assign n567 = ( n1348 ) | ( n1370 ) ;
 assign n568 = ( n1370 ) | ( n1517 ) ;
 assign n562 = ( n286  &  n563  &  n288  &  n564  &  n565  &  n566  &  n567  &  n568 ) ;
 assign n569 = ( n21  &  (~ n1289) ) | ( n21  &  (~ n1527) ) | ( n21  &  (~ n2392) ) ;
 assign n573 = ( n566  &  n1526 ) ;
 assign n572 = ( (~ n17)  &  (~ n569) ) | ( n563  &  (~ n569)  &  n573 ) ;
 assign n578 = ( (~ n280) ) | ( n567 ) ;
 assign n576 = ( n1325 ) | ( n1370 ) ;
 assign n575 = ( (~ n280)  &  n578 ) | ( n578  &  n576 ) ;
 assign n582 = ( (~ n280) ) | ( n566 ) ;
 assign n580 = ( (~ n479)  &  n1493 ) ;
 assign n581 = ( n1393 ) | ( n1517 ) ;
 assign n579 = ( n582  &  n575  &  n580 ) | ( n582  &  n575  &  n581 ) ;
 assign n583 = ( n21  &  (~ n561) ) | ( n21  &  (~ n568) ) | ( n21  &  (~ n1528) ) ;
 assign n588 = ( (~ n6)  &  n612 ) | ( n612  &  n641 ) | ( (~ n6)  &  (~ n1019) ) | ( n641  &  (~ n1019) ) ;
 assign n589 = ( (~ n10)  &  (~ n426) ) | ( (~ n10)  &  n560 ) | ( (~ n426)  &  n737 ) | ( n560  &  n737 ) ;
 assign n590 = ( (~ n360)  &  n2413  &  n2415 ) | ( n1521  &  n2413  &  n2415 ) ;
 assign n591 = ( n1530  &  n540  &  n543  &  n548  &  n572  &  n579  &  n827  &  n1034 ) ;
 assign n592 = ( n2412  &  n1420  &  n2402  &  n2405  &  n2411  &  n2410  &  n2408  &  n2407 ) ;
 assign n593 = ( n209  &  n207  &  n185  &  n2401  &  n188  &  n2397  &  n2396  &  n2400 ) ;
 assign n587 = ( n588  &  n589  &  n590  &  n591  &  n592  &  n593 ) ;
 assign n595 = ( n1535  &  n1536  &  n1199  &  n1537  &  n1538  &  n1539  &  n1540  &  n1541 ) ;
 assign n596 = ( (~ n146)  &  (~ n277)  &  n281  &  n1457  &  n1459  &  n1460  &  n1461  &  n1462 ) ;
 assign n597 = ( n1311  &  n2390 ) | ( (~ n1534)  &  n2390 ) ;
 assign n598 = ( (~ n34)  &  n559 ) | ( n559  &  n1520 ) | ( (~ n34)  &  n2236 ) | ( n1520  &  n2236 ) ;
 assign n599 = ( (~ n21)  &  n2015  &  n2389 ) | ( n558  &  n2015  &  n2389 ) ;
 assign n600 = ( n1204  &  n2386  &  n2387  &  n2006  &  n1163  &  n1922  &  n2388  &  n2382 ) ;
 assign n601 = ( n2380  &  n1888  &  n1841  &  n1051  &  n2381  &  n1817  &  n1809  &  n2379 ) ;
 assign n602 = ( n1689  &  n1599  &  n1615  &  n1619  &  n1631  &  n1603  &  n1575  &  n2378 ) ;
 assign n594 = ( n595  &  n596  &  n597  &  n598  &  n599  &  n600  &  n601  &  n602 ) ;
 assign n604 = ( (~ n247) ) | ( n544 ) ;
 assign n603 = ( (~ n247)  &  n604 ) | ( n501  &  n604 ) ;
 assign n606 = ( (~ n247) ) | ( n1431 ) ;
 assign n605 = ( (~ n247)  &  n606 ) | ( n503  &  n606 ) ;
 assign n609 = ( (~ n247) ) | ( n1012 ) ;
 assign n608 = ( n1480  &  n1476 ) ;
 assign n607 = ( (~ n247)  &  n609 ) | ( n609  &  n608 ) ;
 assign n611 = ( (~ i_15_) ) | ( n1475 ) ;
 assign n612 = ( n1390 ) | ( n1517 ) ;
 assign n610 = ( n611  &  n612 ) ;
 assign n613 = ( (~ n34)  &  n610 ) | ( n508  &  n610 ) | ( (~ n34)  &  (~ n616) ) | ( n508  &  (~ n616) ) ;
 assign n614 = ( n39  &  (~ n959) ) | ( n135  &  (~ n959) ) | ( n400  &  (~ n959) ) ;
 assign n616 = ( (~ n1362)  &  n1388 ) ;
 assign n615 = ( n360  &  (~ n1122) ) | ( n616  &  (~ n1122) ) ;
 assign n619 = ( (~ n39)  &  (~ n135) ) | ( (~ n39)  &  n566 ) | ( (~ n135)  &  n1077 ) | ( n566  &  n1077 ) ;
 assign n620 = ( n927  &  n1548  &  n924  &  n1549 ) ;
 assign n621 = ( (~ n332)  &  (~ n426) ) | ( (~ n332)  &  n541 ) | ( (~ n426)  &  n641 ) | ( n541  &  n641 ) ;
 assign n622 = ( (~ n248)  &  n334 ) | ( (~ n248)  &  n1237 ) | ( n334  &  n1523 ) | ( n1237  &  n1523 ) ;
 assign n623 = ( (~ n615)  &  n1188  &  n1242  &  n1903  &  n2339  &  n2340  &  n2341 ) ;
 assign n624 = ( n1992  &  n1911  &  n1975  &  n2338  &  n1811  &  n2025  &  n1806  &  n2333 ) ;
 assign n625 = ( n1865  &  n1866  &  n1846  &  n2332  &  n1893  &  n1231  &  n1901  &  n2328 ) ;
 assign n626 = ( n2325  &  n2326  &  n783  &  n785  &  n1682  &  n1696  &  n2327  &  n2322 ) ;
 assign n618 = ( n619  &  n620  &  n621  &  n622  &  n623  &  n624  &  n625  &  n626 ) ;
 assign n627 = ( (~ n295)  &  (~ n788) ) | ( (~ n295)  &  (~ n1551) ) ;
 assign n630 = ( (~ n323)  &  n400 ) | ( n400  &  (~ n1523) ) | ( n400  &  (~ n1552) ) ;
 assign n634 = ( n291  &  (~ n363) ) | ( (~ n300)  &  (~ n363) ) | ( n291  &  n466 ) | ( (~ n300)  &  n466 ) ;
 assign n635 = ( (~ n426)  &  n2424 ) | ( n1915  &  n2424 ) ;
 assign n636 = ( (~ n34)  &  n2420  &  n2422 ) | ( n2420  &  n2422  &  n2423 ) ;
 assign n637 = ( n1954  &  n1981  &  n2004  &  n1849  &  n1686  &  n1179  &  n2418  &  n2417 ) ;
 assign n638 = ( n594  &  n1559  &  n587  &  n533  &  n538  &  n517  &  n519  &  n2427 ) ;
 assign n639 = ( n435  &  n414  &  n511  &  n1555  &  n618  &  n2426 ) ;
 assign n633 = ( n634  &  n635  &  n636  &  n637  &  n638  &  n639 ) ;
 assign n642 = ( (~ n6) ) | ( n740 ) ;
 assign n641 = ( n1398 ) | ( n1517 ) ;
 assign n640 = ( (~ n6)  &  n642 ) | ( n642  &  n641 ) ;
 assign n643 = ( (~ n6)  &  n640 ) | ( n312  &  n640 ) ;
 assign n646 = ( (~ n10) ) | ( n1523 ) ;
 assign n647 = ( (~ n10) ) | ( n537 ) ;
 assign n645 = ( n1325 ) | ( n1391 ) ;
 assign n644 = ( (~ n10)  &  n646  &  n647 ) | ( n646  &  n647  &  n645 ) ;
 assign n649 = ( (~ n131) ) | ( n1523 ) ;
 assign n650 = ( (~ n131) ) | ( n537 ) ;
 assign n648 = ( (~ n131)  &  n649  &  n650 ) | ( n645  &  n649  &  n650 ) ;
 assign n653 = ( (~ n10) ) | ( n561 ) ;
 assign n654 = ( (~ n10) ) | ( n611 ) ;
 assign n652 = ( n1325 ) | ( n1390 ) ;
 assign n651 = ( (~ n10)  &  n653  &  n654 ) | ( n653  &  n654  &  n652 ) ;
 assign n656 = ( (~ n131) ) | ( n561 ) ;
 assign n657 = ( (~ n131) ) | ( n611 ) ;
 assign n655 = ( (~ n131)  &  n656  &  n657 ) | ( n652  &  n656  &  n657 ) ;
 assign n660 = ( (~ n139) ) | ( n566 ) ;
 assign n659 = ( n1325 ) | ( n1375 ) ;
 assign n658 = ( (~ n139)  &  n660 ) | ( n660  &  n659 ) ;
 assign n662 = ( (~ n139)  &  (~ n616) ) | ( (~ n139)  &  n1253 ) | ( (~ n616)  &  n1523 ) | ( n1253  &  n1523 ) ;
 assign n663 = ( (~ n357)  &  n2443 ) | ( n705  &  n2443 ) ;
 assign n661 = ( n662  &  n618  &  n663 ) ;
 assign n666 = ( (~ n247) ) | ( n380 ) ;
 assign n667 = ( (~ n247) ) | ( n1519 ) ;
 assign n665 = ( n1325 ) | ( n1327 ) ;
 assign n664 = ( (~ n247)  &  n666  &  n667 ) | ( n666  &  n667  &  n665 ) ;
 assign n669 = ( (~ n247) ) | ( n740 ) ;
 assign n670 = ( (~ n247) ) | ( n641 ) ;
 assign n668 = ( (~ n247)  &  n669  &  n670 ) | ( n312  &  n669  &  n670 ) ;
 assign n672 = ( (~ n10) ) | ( n564 ) ;
 assign n673 = ( (~ n10) ) | ( n1250 ) ;
 assign n671 = ( (~ n10)  &  n672  &  n673 ) | ( n262  &  n672  &  n673 ) ;
 assign n675 = ( (~ n10) ) | ( n706 ) ;
 assign n674 = ( (~ n10)  &  n675 ) | ( n312  &  n675 ) ;
 assign n678 = ( (~ n34) ) | ( n839 ) ;
 assign n679 = ( n1612  &  n1602  &  n73 ) ;
 assign n677 = ( n524  &  n1562 ) ;
 assign n676 = ( (~ n21)  &  n678  &  n679 ) | ( n678  &  n679  &  n677 ) ;
 assign n681 = ( n707  &  n812  &  n864 ) ;
 assign n680 = ( n261  &  n190  &  n681 ) ;
 assign n683 = ( n10 ) | ( n21 ) ;
 assign n682 = ( n683  &  (~ n799) ) | ( (~ n799)  &  (~ n990) ) ;
 assign n686 = ( (~ n10) ) | ( n2609 ) ;
 assign n687 = ( (~ n10) ) | ( n677 ) ;
 assign n688 = ( (~ n280) ) | ( n707 ) ;
 assign n689 = ( n1331 ) | ( (~ n1534) ) ;
 assign n690 = ( (~ n280) ) | ( n839 ) ;
 assign n691 = ( n2432  &  n2433  &  n2434  &  n2435 ) ;
 assign n692 = ( (~ n11)  &  n1618  &  n1630  &  n1649  &  n1666  &  n1673  &  n2429  &  n2431 ) ;
 assign n693 = ( n664  &  n668  &  n671  &  n1568  &  n1566  &  n676  &  n2442  &  n2437 ) ;
 assign n685 = ( n686  &  n687  &  n688  &  n689  &  n690  &  n691  &  n692  &  n693 ) ;
 assign n695 = ( (~ n6) ) | ( n1250 ) ;
 assign n696 = ( (~ n6) ) | ( n1077 ) ;
 assign n694 = ( (~ n6)  &  n695  &  n696 ) | ( n262  &  n695  &  n696 ) ;
 assign n700 = ( (~ n426) ) | ( n537 ) ;
 assign n697 = ( (~ n16)  &  n700 ) | ( (~ n426)  &  n700 ) ;
 assign n702 = ( n537  &  n611 ) ;
 assign n701 = ( (~ n616) ) | ( n702 ) ;
 assign n704 = ( n1391 ) | ( n1522 ) ;
 assign n705 = ( n1290  &  n1519 ) ;
 assign n706 = ( n1393 ) | ( n1522 ) ;
 assign n707 = ( n1390 ) | ( n1522 ) ;
 assign n703 = ( n556  &  n704  &  n705  &  n706  &  n707  &  n380 ) ;
 assign n709 = ( n1374 ) | ( n1391 ) ;
 assign n710 = ( (~ n1226)  &  n1474  &  n1562 ) ;
 assign n711 = ( n564  &  n262 ) ;
 assign n708 = ( (~ n16)  &  n381  &  n709  &  n710  &  n711 ) ;
 assign n712 = ( n180  &  n175  &  n502  &  n470  &  n709  &  n318 ) ;
 assign n714 = ( (~ n6) ) | ( n739 ) ;
 assign n715 = ( (~ n6) ) | ( n1122 ) ;
 assign n713 = ( (~ n6)  &  n714  &  n715 ) | ( n313  &  n714  &  n715 ) ;
 assign n716 = ( n313  &  n262  &  n659  &  n645 ) ;
 assign n718 = ( (~ n247) ) | ( n739 ) ;
 assign n719 = ( (~ n247) ) | ( n1122 ) ;
 assign n720 = ( (~ n247) ) | ( n1077 ) ;
 assign n721 = ( (~ n247)  &  n2228 ) | ( n716  &  n2228 ) ;
 assign n722 = ( n1574  &  n1575 ) ;
 assign n723 = ( n1570  &  n1571  &  n1572  &  n1573 ) ;
 assign n724 = ( (~ n6) ) | ( n645 ) ;
 assign n717 = ( n718  &  n719  &  n720  &  n721  &  n713  &  n722  &  n723  &  n724 ) ;
 assign n728 = ( n292 ) | ( n727 ) ;
 assign n726 = ( n1325 ) | ( n1393 ) ;
 assign n727 = ( n1339 ) | ( (~ n1368) ) ;
 assign n725 = ( n728  &  n726 ) | ( n728  &  n727 ) ;
 assign n730 = ( n641  &  n1122 ) ;
 assign n729 = ( n547  &  n725  &  n730 ) | ( n547  &  n725  &  (~ n1016) ) ;
 assign n732 = ( n358  &  (~ n799) ) | ( n479  &  (~ n799) ) ;
 assign n734 = ( (~ n378)  &  n994 ) ;
 assign n733 = ( (~ n6)  &  n295  &  (~ n360)  &  n734 ) ;
 assign n737 = ( n1346 ) | ( n1522 ) ;
 assign n736 = ( (~ n139)  &  n526  &  n531 ) | ( n526  &  n531  &  n737 ) ;
 assign n739 = ( n1348 ) | ( n1396 ) ;
 assign n740 = ( n1348 ) | ( n1398 ) ;
 assign n738 = ( n739  &  n740 ) ;
 assign n742 = ( n190  &  n1376  &  n340 ) ;
 assign n743 = ( n1374 ) | ( n1375 ) ;
 assign n741 = ( n742  &  n261  &  n743  &  n341 ) ;
 assign n744 = ( (~ n175)  &  n378 ) | ( n378  &  (~ n1576) ) ;
 assign n747 = ( n135  &  (~ n561) ) | ( n135  &  (~ n1523) ) ;
 assign n748 = ( n21  &  (~ n537) ) | ( n21  &  (~ n1376) ) ;
 assign n750 = ( (~ n296)  &  (~ n381) ) | ( (~ n296)  &  (~ n812) ) | ( (~ n296)  &  (~ n1528) ) ;
 assign n753 = ( (~ n10)  &  (~ n248) ) | ( (~ n248)  &  n559 ) | ( (~ n10)  &  n993 ) | ( n559  &  n993 ) ;
 assign n754 = ( (~ n280)  &  n2475 ) | ( n1524  &  n2475 ) ;
 assign n755 = ( (~ n34)  &  n449  &  n1099 ) | ( n449  &  n1099  &  n1195 ) ;
 assign n752 = ( n736  &  n594  &  n753  &  n454  &  n754  &  n755 ) ;
 assign n757 = ( n214 ) | ( n1364 ) ;
 assign n758 = ( n897 ) | ( n1364 ) ;
 assign n759 = ( n508 ) | ( n1364 ) ;
 assign n760 = ( n959 ) | ( n1364 ) ;
 assign n761 = ( n953 ) | ( n1364 ) ;
 assign n762 = ( n1329 ) | ( n1364 ) ;
 assign n763 = ( n213 ) | ( n1364 ) ;
 assign n764 = ( n1801  &  n494 ) | ( n1801  &  n1364 ) ;
 assign n756 = ( n757  &  n758  &  n759  &  n760  &  n761  &  n762  &  n763  &  n764 ) ;
 assign n766 = ( n1372 ) | ( n1391 ) ;
 assign n765 = ( n766  &  n576  &  n507  &  n413  &  n465 ) ;
 assign n768 = ( n1314 ) | ( n1372 ) ;
 assign n767 = ( n506  &  n768 ) ;
 assign n772 = ( n214 ) | ( n771 ) ;
 assign n773 = ( (~ n71) ) | ( (~ n1337) ) ;
 assign n771 = ( (~ n1337) ) | ( n1361 ) ;
 assign n769 = ( n772  &  n773  &  n771 ) | ( n772  &  n773  &  (~ n775) ) ;
 assign n776 = ( n159  &  (~ n1361) ) ;
 assign n775 = ( (~ n516) ) | ( (~ n819) ) | ( n892 ) ;
 assign n774 = ( (~ n214)  &  n776 ) | ( n776  &  n775 ) ;
 assign n779 = ( (~ n6) ) | ( n1484 ) ;
 assign n780 = ( n1413  &  n1487  &  n2401 ) ;
 assign n778 = ( n815  &  n854 ) ;
 assign n777 = ( (~ n6)  &  n779  &  n780 ) | ( n779  &  n780  &  n778 ) ;
 assign n782 = ( (~ n6) ) | ( n412 ) ;
 assign n783 = ( (~ n6) ) | ( n561 ) ;
 assign n784 = ( (~ n6) ) | ( n611 ) ;
 assign n785 = ( (~ n6) ) | ( n612 ) ;
 assign n786 = ( (~ n6)  &  n186 ) | ( n186  &  n652 ) ;
 assign n781 = ( n782  &  n783  &  n784  &  n785  &  n786  &  n517 ) ;
 assign n789 = ( (~ n6) ) | ( n576 ) ;
 assign n788 = ( n1477  &  n743 ) ;
 assign n787 = ( (~ n6)  &  n789 ) | ( n789  &  n788 ) ;
 assign n791 = ( (~ n247) ) | ( n959 ) ;
 assign n790 = ( (~ n247)  &  n791 ) | ( n504  &  n791 ) ;
 assign n793 = ( (~ n247) ) | ( n1478 ) ;
 assign n794 = ( (~ n247) ) | ( n737 ) ;
 assign n792 = ( (~ n247)  &  n793  &  n794 ) | ( n263  &  n793  &  n794 ) ;
 assign n795 = ( (~ n6) ) | ( n263 ) ;
 assign n796 = ( (~ n6) ) | ( n345 ) ;
 assign n799 = ( n1398 ) | ( n1522 ) ;
 assign n800 = ( n1315 ) | ( n1393 ) ;
 assign n797 = ( (~ n6)  &  (~ n363) ) | ( (~ n6)  &  n799 ) | ( (~ n363)  &  n800 ) | ( n799  &  n800 ) ;
 assign n802 = ( (~ n247) ) | ( n568 ) ;
 assign n803 = ( (~ n6) ) | ( n1958 ) ;
 assign n804 = ( (~ n247) ) | ( n464 ) ;
 assign n805 = ( (~ n247)  &  n797 ) | ( n797  &  n837 ) ;
 assign n806 = ( n1606  &  n790 ) ;
 assign n807 = ( n1613  &  n1614  &  n1615  &  n1616  &  n1617 ) ;
 assign n808 = ( n1583  &  n551  &  n1609  &  n1610  &  n1611  &  n1612  &  n796 ) ;
 assign n801 = ( n802  &  n803  &  n804  &  n805  &  n787  &  n806  &  n807  &  n808 ) ;
 assign n810 = ( n1315 ) | ( n1346 ) ;
 assign n809 = ( (~ n363) ) | ( n810 ) ;
 assign n813 = ( n1618  &  n1619  &  n1620  &  n1621  &  n1622  &  n1584  &  n809 ) ;
 assign n812 = ( n1314 ) | ( n1522 ) ;
 assign n811 = ( (~ n6)  &  n813 ) | ( n813  &  n812 ) ;
 assign n816 = ( (~ n6) ) | ( n704 ) ;
 assign n815 = ( n1315 ) | ( n1367 ) ;
 assign n814 = ( (~ n247)  &  n552  &  n816 ) | ( n552  &  n816  &  n815 ) ;
 assign n819 = ( n897  &  n494  &  n1596 ) ;
 assign n817 = ( n819 ) | ( (~ n1624) ) ;
 assign n821 = ( n1264  &  n1379 ) ;
 assign n820 = ( (~ n10)  &  (~ n131) ) | ( (~ n10)  &  n812 ) | ( (~ n131)  &  n821 ) | ( n812  &  n821 ) ;
 assign n823 = ( n316  &  n1376 ) ;
 assign n824 = ( n1395  &  n190 ) ;
 assign n822 = ( n823  &  n824  &  n318  &  n341 ) ;
 assign n826 = ( n1625  &  n1626  &  n1627  &  n1628 ) ;
 assign n827 = ( n211  &  n948  &  n947  &  n951  &  n196  &  n1529 ) ;
 assign n828 = ( (~ n472)  &  n1495  &  n1496  &  n1498 ) ;
 assign n829 = ( n317  &  n305  &  n1481 ) ;
 assign n830 = ( n1783  &  n928  &  n2133  &  n910  &  n2106  &  n201  &  n189  &  n2494 ) ;
 assign n825 = ( n826  &  n717  &  n620  &  n827  &  n499  &  n828  &  n829  &  n830 ) ;
 assign n832 = ( (~ n247) ) | ( n412 ) ;
 assign n833 = ( (~ n247) ) | ( n561 ) ;
 assign n831 = ( (~ n247)  &  n832  &  n833 ) | ( n652  &  n832  &  n833 ) ;
 assign n834 = ( n6  &  (~ n659) ) | ( n6  &  (~ n839) ) ;
 assign n837 = ( n1315 ) | ( n1370 ) ;
 assign n836 = ( (~ n6) ) | ( n837 ) ;
 assign n840 = ( (~ n10) ) | ( n568 ) ;
 assign n839 = ( n1375 ) | ( n1522 ) ;
 assign n838 = ( (~ n10)  &  n840 ) | ( n464  &  n840  &  n839 ) ;
 assign n842 = ( (~ n131) ) | ( n464 ) ;
 assign n841 = ( (~ n131)  &  n842 ) | ( n839  &  n842 ) ;
 assign n844 = ( (~ n378) ) | ( n800 ) ;
 assign n845 = ( (~ n10) ) | ( n1206 ) ;
 assign n846 = ( (~ n10) ) | ( n581 ) ;
 assign n847 = ( (~ n10)  &  (~ n131) ) | ( (~ n131)  &  n799 ) | ( (~ n10)  &  n1206 ) | ( n799  &  n1206 ) ;
 assign n843 = ( n844  &  n550  &  n845  &  n846  &  n847  &  n841 ) ;
 assign n849 = ( (~ n131) ) | ( n1269 ) ;
 assign n850 = ( (~ n131) ) | ( n1043 ) ;
 assign n848 = ( (~ n131)  &  n849  &  n850 ) | ( n704  &  n849  &  n850 ) ;
 assign n852 = ( n1564  &  n1009 ) ;
 assign n851 = ( (~ n6) ) | ( n852 ) ;
 assign n855 = ( (~ n10) ) | ( n1484 ) ;
 assign n856 = ( (~ n10) ) | ( n560 ) ;
 assign n854 = ( n1396 ) | ( n1522 ) ;
 assign n853 = ( (~ n10)  &  n855  &  n856 ) | ( n855  &  n856  &  n854 ) ;
 assign n857 = ( n131  &  (~ n1352) ) | ( n131  &  (~ n1658) ) ;
 assign n859 = ( n131  &  (~ n707) ) | ( n131  &  (~ n810) ) | ( n131  &  (~ n1659) ) ;
 assign n862 = ( (~ n10) ) | ( n810 ) ;
 assign n864 = ( n1321 ) | ( n1522 ) ;
 assign n863 = ( (~ n13)  &  n176  &  n318  &  n581  &  n799  &  n864 ) ;
 assign n866 = ( (~ n175)  &  n378 ) | ( n378  &  (~ n1280) ) ;
 assign n869 = ( n251  &  n1181  &  n1652 ) ;
 assign n870 = ( n1672  &  n1669  &  n1676  &  n1687  &  n1681 ) ;
 assign n871 = ( (~ n11)  &  (~ n128)  &  n1301  &  n1415  &  n1585  &  n1665  &  n2129  &  n2492 ) ;
 assign n872 = ( n1453  &  n1407  &  n1488  &  n2139  &  n1412  &  n2092  &  n237  &  n2491 ) ;
 assign n873 = ( (~ n7)  &  n224  &  n2067  &  n2184  &  n2239  &  n2291  &  n2361  &  n2490 ) ;
 assign n868 = ( n838  &  n869  &  n843  &  n848  &  n870  &  n871  &  n872  &  n873 ) ;
 assign n875 = ( n1701  &  n1702  &  n1703  &  n1704  &  n1705  &  n1706  &  n1707 ) ;
 assign n876 = ( n234  &  n1698  &  n225  &  n385  &  n1699  &  n1700 ) ;
 assign n877 = ( (~ n10)  &  n540 ) | ( n540  &  n2040 ) ;
 assign n878 = ( n1467  &  n648  &  n1692  &  n1693  &  n1694  &  n1695  &  n1696  &  n1697 ) ;
 assign n874 = ( n875  &  n876  &  n877  &  n878 ) ;
 assign n879 = ( n10  &  (~ n737) ) | ( n10  &  (~ n1562) ) ;
 assign n882 = ( n131  &  (~ n312) ) | ( n131  &  (~ n837) ) | ( n131  &  (~ n1562) ) ;
 assign n884 = ( n263 ) | ( (~ n378) ) ;
 assign n889 = ( n1724  &  n912  &  n1737  &  n868  &  n1743  &  n1763  &  n1764  &  n1765 ) ;
 assign n887 = ( i_7_ ) | ( i_6_ ) ;
 assign n886 = ( n889  &  n887 ) | ( n889  &  (~ n1762) ) ;
 assign n893 = ( n160  &  (~ n1361) ) ;
 assign n892 = ( (~ n959) ) | ( (~ n1329) ) ;
 assign n890 = ( (~ n214)  &  n893 ) | ( (~ n819)  &  n893 ) | ( n893  &  n892 ) ;
 assign n894 = ( n214 ) | ( (~ n1774) ) ;
 assign n897 = ( n1347 ) | ( n1378 ) ;
 assign n896 = ( n897 ) | ( (~ n1784) ) ;
 assign n901 = ( n508 ) | ( (~ n978) ) ;
 assign n900 = ( n984  &  (~ n1624) ) ;
 assign n899 = ( n759  &  n901  &  n900 ) | ( n759  &  n901  &  n508 ) ;
 assign n903 = ( (~ n247) ) | ( n324 ) ;
 assign n904 = ( (~ n6)  &  n205 ) | ( n205  &  n260 ) ;
 assign n905 = ( n1714  &  n1715  &  n1716  &  n1717 ) ;
 assign n906 = ( n1711  &  n668  &  n1712  &  n1713 ) ;
 assign n902 = ( n181  &  n182  &  n903  &  n904  &  n905  &  n906  &  n640  &  n447 ) ;
 assign n908 = ( (~ n247) ) | ( n576 ) ;
 assign n907 = ( (~ n247)  &  n908 ) | ( n788  &  n908 ) ;
 assign n910 = ( (~ n247) ) | ( n1271 ) ;
 assign n911 = ( (~ n247) ) | ( n1958 ) ;
 assign n912 = ( n1733  &  n227  &  n228  &  n233  &  n387  &  n1734  &  n1735  &  n1736 ) ;
 assign n913 = ( (~ n131)  &  n1724  &  n2445 ) | ( n837  &  n1724  &  n2445 ) ;
 assign n909 = ( n526  &  n910  &  n528  &  n687  &  n911  &  n907  &  n912  &  n913 ) ;
 assign n915 = ( (~ n247) ) | ( n567 ) ;
 assign n916 = ( (~ n247) ) | ( n566 ) ;
 assign n914 = ( (~ n247)  &  n915  &  n916 ) | ( n659  &  n915  &  n916 ) ;
 assign n918 = ( (~ n10) ) | ( n1521 ) ;
 assign n917 = ( (~ n10)  &  n918 ) | ( n821  &  n918 ) ;
 assign n919 = ( n247  &  (~ n262) ) | ( n247  &  (~ n921) ) ;
 assign n921 = ( n1321 ) | ( n1374 ) ;
 assign n920 = ( (~ n6) ) | ( n921 ) ;
 assign n923 = ( (~ n247) ) | ( n1479 ) ;
 assign n924 = ( (~ n247) ) | ( n1523 ) ;
 assign n922 = ( (~ n247)  &  n923  &  n924 ) | ( n645  &  n923  &  n924 ) ;
 assign n926 = ( (~ n6) ) | ( n1479 ) ;
 assign n927 = ( (~ n6) ) | ( n1523 ) ;
 assign n928 = ( (~ n6) ) | ( n1394 ) ;
 assign n929 = ( (~ n6)  &  n194 ) | ( n194  &  n645 ) ;
 assign n925 = ( n926  &  n927  &  n928  &  n929  &  n922  &  n723  &  n533  &  n605 ) ;
 assign n931 = ( n1601  &  n1602  &  n1603 ) ;
 assign n932 = ( n1623  &  n1452  &  n814 ) ;
 assign n933 = ( (~ n6)  &  n777  &  n1597 ) | ( n777  &  n812  &  n1597 ) ;
 assign n934 = ( (~ n247) ) | ( n2606 ) ;
 assign n935 = ( n544 ) | ( (~ n978) ) ;
 assign n936 = ( (~ n247) ) | ( n508 ) ;
 assign n937 = ( n2032  &  n1771  &  n967 ) | ( n2032  &  n1771  &  n544 ) ;
 assign n930 = ( n813  &  n931  &  n932  &  n933  &  n934  &  n935  &  n936  &  n937 ) ;
 assign n939 = ( (~ n71) ) | ( n1589 ) ;
 assign n940 = ( (~ n71) ) | ( n1510 ) ;
 assign n941 = ( (~ n71)  &  n491 ) | ( (~ n119)  &  n491 ) | ( (~ n71)  &  n953 ) | ( (~ n119)  &  n953 ) ;
 assign n938 = ( n939  &  n940  &  n941 ) ;
 assign n945 = ( (~ n47) ) | ( n1510 ) ;
 assign n942 = ( (~ n47)  &  n945 ) | ( (~ n119)  &  n945 ) ;
 assign n947 = ( (~ n247) ) | ( n1473 ) ;
 assign n948 = ( (~ n247) ) | ( n541 ) ;
 assign n946 = ( (~ n247)  &  n947  &  n948 ) | ( n313  &  n947  &  n948 ) ;
 assign n951 = ( (~ n247) ) | ( n292 ) ;
 assign n950 = ( n507  &  n470 ) ;
 assign n949 = ( (~ n247)  &  n951 ) | ( n951  &  n950 ) ;
 assign n953 = ( i_15_ ) | ( n1345 ) ;
 assign n952 = ( n953 ) | ( n900 ) ;
 assign n954 = ( n131  &  (~ n263) ) | ( n131  &  (~ n312) ) | ( n131  &  (~ n812) ) ;
 assign n955 = ( (~ n516)  &  n893 ) | ( (~ n516)  &  (~ n1364) ) ;
 assign n959 = ( n1325 ) | ( n1346 ) ;
 assign n960 = ( n491  &  n984 ) ;
 assign n958 = ( n959 ) | ( n960 ) ;
 assign n962 = ( (~ n119) ) | ( n1380 ) ;
 assign n963 = ( n1380 ) | ( n1510 ) ;
 assign n961 = ( n962  &  n963  &  n213 ) | ( n962  &  n963  &  n491 ) ;
 assign n965 = ( n887 ) | ( n1510 ) ;
 assign n964 = ( (~ n119)  &  n965 ) | ( n887  &  n965 ) ;
 assign n968 = ( n468 ) | ( (~ n978) ) ;
 assign n967 = ( n1363  &  (~ n1784) ) ;
 assign n966 = ( n968  &  n967 ) | ( n968  &  n468 ) ;
 assign n970 = ( n1592  &  n2321  &  n1502 ) ;
 assign n969 = ( n763  &  n970  &  n900 ) | ( n763  &  n970  &  n213 ) ;
 assign n972 = ( n1514  &  n1767  &  n1594  &  n1503  &  n762 ) ;
 assign n973 = ( n960  &  n1363 ) | ( n1329  &  n1363 ) | ( n960  &  n516 ) | ( n1329  &  n516 ) ;
 assign n971 = ( n972  &  n964  &  n961  &  n966  &  n969  &  n973 ) ;
 assign n976 = ( n773  &  n1515  &  n1801 ) ;
 assign n977 = ( n492  &  (~ n1762) ) | ( (~ n71)  &  n492  &  n887 ) ;
 assign n978 = ( n1337  &  (~ n1362) ) ;
 assign n979 = ( (~ n771) ) | ( n776 ) ;
 assign n982 = ( n2489 ) | ( n2502 ) ;
 assign n980 = ( i_9_  &  (~ i_10_) ) ;
 assign n981 = ( (~ i_9_)  &  i_10_ ) ;
 assign n984 = ( n771  &  (~ n1774) ) ;
 assign n983 = ( (~ n892) ) | ( n984 ) ;
 assign n987 = ( n1797  &  n972  &  n983  &  n899 ) ;
 assign n988 = ( n942  &  (~ n982)  &  n2514 ) | ( n942  &  (~ n981)  &  n2514 ) ;
 assign n985 = ( (~ n64)  &  n964  &  n987  &  n988 ) ;
 assign n990 = ( (~ n157) ) | ( (~ n1368) ) ;
 assign n991 = ( n768  &  n1478 ) ;
 assign n989 = ( n990 ) | ( n991 ) ;
 assign n993 = ( n1346 ) | ( n1517 ) ;
 assign n994 = ( n1361 ) | ( (~ n1368) ) ;
 assign n992 = ( n993 ) | ( n994 ) ;
 assign n995 = ( (~ n260)  &  (~ n990) ) | ( (~ n799)  &  (~ n990) ) ;
 assign n996 = ( n799 ) | ( n994 ) ;
 assign n997 = ( (~ n413)  &  (~ n994) ) | ( (~ n994)  &  (~ n1210) ) ;
 assign n1002 = ( n994 ) | ( n743 ) ;
 assign n1003 = ( n2305  &  n2337  &  n2338 ) ;
 assign n1001 = ( n839  &  n1805 ) ;
 assign n1004 = ( (~ n247)  &  n802  &  n804 ) | ( n802  &  n804  &  n837 ) ;
 assign n1005 = ( (~ n6) ) | ( n823 ) ;
 assign n1007 = ( n261  &  n1071 ) ;
 assign n1006 = ( (~ n247) ) | ( n1007 ) ;
 assign n1010 = ( n1767  &  n817  &  n1768  &  n1769 ) ;
 assign n1009 = ( n1315 ) | ( n1369 ) ;
 assign n1013 = ( n2517  &  n545 ) | ( n2517  &  n1820  &  n953 ) ;
 assign n1012 = ( n1325 ) | ( n1369 ) ;
 assign n1011 = ( n725  &  n1013  &  n1012 ) | ( n725  &  n1013  &  n727 ) ;
 assign n1016 = ( n158  &  n1388 ) ;
 assign n1019 = ( n1355  &  n1388 ) ;
 assign n1021 = ( n135 ) | ( n280 ) ;
 assign n1020 = ( (~ n740)  &  n1021 ) | ( n1021  &  (~ n1524) ) ;
 assign n1023 = ( (~ n280) ) | ( n1071 ) ;
 assign n1024 = ( (~ n280) ) | ( n1329 ) ;
 assign n1025 = ( (~ n280) ) | ( n508 ) ;
 assign n1026 = ( (~ n135)  &  n2349 ) | ( n508  &  n2349 ) ;
 assign n1027 = ( n1311 ) | ( (~ n1534) ) ;
 assign n1028 = ( n2050  &  n2252  &  n2188  &  n2276  &  n2364  &  n2301 ) ;
 assign n1022 = ( n1023  &  n1024  &  n1025  &  n1026  &  n1027  &  n1028 ) ;
 assign n1030 = ( n709  &  n1823 ) ;
 assign n1029 = ( (~ n135) ) | ( n1030 ) ;
 assign n1033 = ( (~ i_11_) ) | ( (~ n980) ) ;
 assign n1031 = ( n1033 ) | ( (~ n1525) ) ;
 assign n1035 = ( i_11_ ) | ( n1323 ) ;
 assign n1034 = ( n1035 ) | ( (~ n1525) ) ;
 assign n1037 = ( (~ n280) ) | ( n1077 ) ;
 assign n1038 = ( (~ n280) ) | ( n1075 ) ;
 assign n1039 = ( (~ n280) ) | ( n921 ) ;
 assign n1040 = ( (~ n280)  &  n2187 ) | ( n288  &  n1076  &  n2187 ) ;
 assign n1036 = ( n1037  &  n1038  &  n1039  &  n1040 ) ;
 assign n1041 = ( (~ n280) ) | ( n1030 ) ;
 assign n1043 = ( n1385 ) | ( n1517 ) ;
 assign n1044 = ( n1122  &  n1473  &  n1276 ) ;
 assign n1045 = ( n704  &  n1123 ) ;
 assign n1042 = ( n292  &  n1043  &  n739  &  n1044  &  n1045 ) ;
 assign n1047 = ( n243 ) | ( (~ n280) ) ;
 assign n1048 = ( (~ n280) ) | ( n1395 ) ;
 assign n1049 = ( (~ n135) ) | ( n536 ) ;
 assign n1050 = ( (~ n280) ) | ( n1484 ) ;
 assign n1051 = ( (~ n280) ) | ( n560 ) ;
 assign n1052 = ( (~ n135)  &  n1825 ) | ( n1042  &  n1825 ) ;
 assign n1053 = ( (~ n280)  &  n2519 ) | ( n190  &  n854  &  n2519 ) ;
 assign n1054 = ( n2251  &  n2299  &  n2047  &  n2109  &  n2186  &  n2127  &  n689  &  n2518 ) ;
 assign n1046 = ( n1047  &  n1048  &  n1049  &  n1050  &  n1051  &  n1052  &  n1053  &  n1054 ) ;
 assign n1056 = ( n318  &  n345 ) ;
 assign n1057 = ( n260  &  n1834  &  n706  &  n737 ) ;
 assign n1055 = ( n1056  &  n1057  &  n852  &  n800 ) ;
 assign n1059 = ( (~ n476)  &  n1071  &  n1237 ) ;
 assign n1060 = ( n342  &  n1210  &  n1836  &  n1519  &  n1376  &  n1478 ) ;
 assign n1061 = ( n837  &  n839 ) ;
 assign n1062 = ( n324  &  n530  &  n340 ) ;
 assign n1058 = ( n710  &  n563  &  n1059  &  n1060  &  n1061  &  n864  &  n854  &  n1062 ) ;
 assign n1063 = ( n1849  &  n1031  &  n1850  &  n1851  &  n1852  &  n1853  &  n1854  &  n1855 ) ;
 assign n1064 = ( n1843  &  n1844  &  n1845  &  n1846  &  n1847  &  n1848  &  n1034 ) ;
 assign n1065 = ( n1856  &  n1857  &  n1858  &  n1859  &  n1860  &  n1861  &  n1862  &  n1863 ) ;
 assign n1066 = ( n1864  &  n1865  &  n1866  &  n1867  &  n1868  &  n1869  &  n1870  &  n1871 ) ;
 assign n1067 = ( n1886  &  n1882  &  n1096  &  n1872 ) ;
 assign n1068 = ( (~ n132)  &  n1036  &  n1046  &  n1837  &  n2091  &  n2115  &  n2524  &  n2525 ) ;
 assign n1069 = ( n2105  &  n2116  &  n2190  &  n2280  &  n2090  &  n2191  &  n2523  &  n2522 ) ;
 assign n1071 = ( n1346 ) | ( n1372 ) ;
 assign n1070 = ( (~ n39) ) | ( n1071 ) ;
 assign n1073 = ( (~ n39) ) | ( n291 ) ;
 assign n1075 = ( n1520  &  n1352  &  n864 ) ;
 assign n1076 = ( n953  &  n465  &  n1824 ) ;
 assign n1077 = ( n1321 ) | ( n1517 ) ;
 assign n1074 = ( n1075  &  n1076  &  n288  &  n1077 ) ;
 assign n1080 = ( (~ n39) ) | ( n214 ) ;
 assign n1078 = ( (~ n39)  &  (~ n43)  &  n1080 ) | ( (~ n43)  &  n1074  &  n1080 ) ;
 assign n1082 = ( (~ n370) ) | ( n1012 ) ;
 assign n1083 = ( (~ n370) ) | ( n453 ) ;
 assign n1084 = ( (~ n370) ) | ( (~ n476) ) ;
 assign n1085 = ( n2278  &  n2367  &  n2368 ) ;
 assign n1086 = ( n1896  &  n1070  &  n1897  &  n1898  &  n1899  &  n1900  &  n1901  &  n1902 ) ;
 assign n1087 = ( (~ n37)  &  n1073  &  n1892  &  n1893  &  n1894  &  n1895 ) ;
 assign n1088 = ( (~ n39)  &  (~ n370) ) | ( (~ n370)  &  n1257 ) | ( (~ n39)  &  n1835 ) | ( n1257  &  n1835 ) ;
 assign n1081 = ( n1082  &  n1083  &  n1084  &  n1085  &  n1086  &  n1087  &  n1088  &  n1078 ) ;
 assign n1090 = ( (~ n139) ) | ( n612 ) ;
 assign n1091 = ( (~ n139) ) | ( n1271 ) ;
 assign n1092 = ( (~ n139) ) | ( n611 ) ;
 assign n1093 = ( (~ n139) ) | ( n544 ) ;
 assign n1094 = ( (~ n139) ) | ( n567 ) ;
 assign n1095 = ( n269  &  n1903  &  n1904 ) ;
 assign n1096 = ( n1881  &  n575 ) ;
 assign n1097 = ( (~ n139)  &  n404  &  n1587 ) | ( n404  &  n1075  &  n1587 ) ;
 assign n1089 = ( n1090  &  n1091  &  n1092  &  n1093  &  n1094  &  n1095  &  n1096  &  n1097 ) ;
 assign n1099 = ( (~ n139) ) | ( n413 ) ;
 assign n1100 = ( (~ n139) ) | ( n1251 ) ;
 assign n1101 = ( (~ n139) ) | ( n1250 ) ;
 assign n1102 = ( (~ n139) ) | ( n1077 ) ;
 assign n1103 = ( (~ n400)  &  (~ n426) ) | ( (~ n426)  &  n711 ) | ( (~ n400)  &  n1075 ) | ( n711  &  n1075 ) ;
 assign n1104 = ( n1229  &  n2052  &  n2077  &  n2051  &  n2260  &  n2096  &  n2189  &  n2150 ) ;
 assign n1098 = ( n1099  &  n1100  &  n1101  &  n1102  &  n1103  &  n1089  &  n1104 ) ;
 assign n1106 = ( n1379  &  n1214 ) ;
 assign n1105 = ( (~ n426) ) | ( n1106 ) ;
 assign n1108 = ( (~ n139) ) | ( n508 ) ;
 assign n1109 = ( (~ n139) ) | ( n1071 ) ;
 assign n1110 = ( (~ n139) ) | ( n530 ) ;
 assign n1111 = ( (~ n143)  &  (~ n400) ) | ( (~ n143)  &  n2526 ) ;
 assign n1112 = ( (~ n426) ) | ( n707 ) ;
 assign n1113 = ( n2371  &  n2055  &  n2118  &  n2057  &  n2263  &  n2075 ) ;
 assign n1107 = ( n1108  &  n1109  &  n1110  &  n1111  &  n1112  &  n1113 ) ;
 assign n1115 = ( (~ n139) ) | ( n466 ) ;
 assign n1114 = ( (~ n139)  &  n1115 ) | ( n341  &  n565  &  n1115 ) ;
 assign n1117 = ( (~ n139) ) | ( n766 ) ;
 assign n1118 = ( n2080  &  n2259  &  n2298 ) ;
 assign n1116 = ( (~ n16)  &  n1117  &  n1118 ) | ( (~ n139)  &  n1117  &  n1118 ) ;
 assign n1120 = ( n739  &  n1565 ) ;
 assign n1121 = ( n292  &  n950 ) ;
 assign n1122 = ( n1396 ) | ( n1517 ) ;
 assign n1123 = ( n1484  &  n560 ) ;
 assign n1119 = ( n1120  &  n778  &  n1121  &  n190  &  n1122  &  n1123 ) ;
 assign n1125 = ( n1905  &  n1906  &  n1907  &  n1908 ) ;
 assign n1126 = ( n1909  &  n1910  &  n1911  &  n1912  &  n1913  &  n1914 ) ;
 assign n1127 = ( (~ n426)  &  n2134  &  n2144 ) | ( n1119  &  n2134  &  n2144 ) ;
 assign n1128 = ( n1485  &  n2336  &  n1416 ) ;
 assign n1129 = ( n2053  &  n2261  &  n2081  &  n2112  &  n2054  &  n2528 ) ;
 assign n1124 = ( n1116  &  n697  &  n1125  &  n1126  &  n1114  &  n1127  &  n1128  &  n1129 ) ;
 assign n1130 = ( n400  &  (~ n1056) ) | ( n400  &  (~ n1836) ) ;
 assign n1136 = ( (~ n340) ) | ( (~ n652) ) | ( (~ n837) ) ;
 assign n1133 = ( n426  &  (~ n1001) ) | ( n426  &  n1136 ) | ( n426  &  (~ n1915) ) ;
 assign n1138 = ( (~ n157) ) | ( n1357 ) ;
 assign n1139 = ( n1339 ) | ( n1357 ) ;
 assign n1137 = ( n1138  &  n1139 ) ;
 assign n1141 = ( (~ n16)  &  n1479 ) ;
 assign n1140 = ( (~ n616) ) | ( n1141 ) ;
 assign n1142 = ( n21  &  (~ n537) ) | ( n21  &  (~ n1823) ) ;
 assign n1145 = ( n1043  &  n1269  &  n342 ) ;
 assign n1144 = ( (~ n17) ) | ( n1145 ) ;
 assign n1148 = ( (~ n34) ) | ( n1186 ) ;
 assign n1149 = ( (~ n280) ) | ( n659 ) ;
 assign n1150 = ( (~ n21)  &  n838 ) | ( n838  &  n2540 ) ;
 assign n1146 = ( (~ n35)  &  n582  &  n1004  &  n1148  &  n1149  &  n1150 ) ;
 assign n1151 = ( n360  &  (~ n1376) ) | ( n360  &  (~ n1562) ) ;
 assign n1153 = ( (~ n834)  &  n1635  &  n1637  &  n1638  &  n1639  &  n1640  &  n1641  &  n1642 ) ;
 assign n1154 = ( n1423  &  n1424  &  n1425 ) ;
 assign n1155 = ( (~ n426)  &  (~ n616) ) | ( (~ n426)  &  n1956 ) | ( (~ n616)  &  n2540 ) | ( n1956  &  n2540 ) ;
 assign n1156 = ( (~ n17)  &  n2543 ) | ( n567  &  n1248  &  n2543 ) ;
 assign n1157 = ( n1940  &  n1063  &  n74  &  n909  &  n1959  &  n1146  &  n1966 ) ;
 assign n1158 = ( n1091  &  (~ n1151)  &  n1838  &  n1881  &  n2285  &  n2373  &  n2449  &  n2541 ) ;
 assign n1152 = ( n1153  &  n787  &  n676  &  n1154  &  n1155  &  n1156  &  n1157  &  n1158 ) ;
 assign n1159 = ( n17  &  (~ n470) ) | ( n17  &  (~ n1120) ) | ( n17  &  (~ n1527) ) ;
 assign n1163 = ( (~ n21) ) | ( n560 ) ;
 assign n1164 = ( (~ n17)  &  n778 ) | ( n778  &  n1045 ) | ( (~ n17)  &  n1428 ) | ( n1045  &  n1428 ) ;
 assign n1162 = ( n439  &  n1163  &  n1164 ) ;
 assign n1165 = ( n17  &  (~ n1479) ) | ( n17  &  (~ n1822) ) ;
 assign n1168 = ( n34  &  (~ n342) ) | ( n34  &  (~ n815) ) ;
 assign n1169 = ( n616  &  (~ n704) ) | ( n616  &  (~ n815) ) | ( n616  &  (~ n1043) ) ;
 assign n1172 = ( (~ n193)  &  n616 ) | ( n616  &  (~ n1044) ) | ( n616  &  (~ n1120) ) ;
 assign n1174 = ( n21  &  (~ n193) ) | ( n21  &  (~ n1121) ) | ( n21  &  (~ n1473) ) ;
 assign n1177 = ( (~ n34) ) | ( n1141 ) ;
 assign n1178 = ( (~ n21) ) | ( n1120 ) ;
 assign n1179 = ( (~ n34) ) | ( n2611 ) ;
 assign n1180 = ( n2028  &  n251  &  n1428 ) | ( n2028  &  n251  &  n1276 ) ;
 assign n1181 = ( n1649  &  n1650  &  n1651 ) ;
 assign n1182 = ( (~ n135)  &  (~ n1172)  &  (~ n1174) ) | ( n854  &  (~ n1172)  &  (~ n1174) ) ;
 assign n1183 = ( n1294  &  n1972  &  n1985  &  n1283  &  n1162  &  n2539 ) ;
 assign n1176 = ( n1177  &  n1178  &  n1179  &  n1180  &  n1181  &  n814  &  n1182  &  n1183 ) ;
 assign n1184 = ( n799  &  n800 ) ;
 assign n1187 = ( n524 ) | ( (~ n616) ) ;
 assign n1188 = ( (~ n616) ) | ( n1518 ) ;
 assign n1186 = ( n567  &  n1562 ) ;
 assign n1185 = ( (~ n616)  &  n1187  &  n1188 ) | ( n1187  &  n1188  &  n1186 ) ;
 assign n1191 = ( n1348 ) | ( n1393 ) ;
 assign n1189 = ( (~ n24)  &  n206  &  n291  &  n1191 ) ;
 assign n1193 = ( n726  &  n448  &  n505 ) ;
 assign n1194 = ( n706  &  n373  &  n260 ) ;
 assign n1195 = ( n291  &  n1191 ) ;
 assign n1196 = ( n740  &  n641 ) ;
 assign n1192 = ( n1193  &  n324  &  n1194  &  n1195  &  n1196 ) ;
 assign n1198 = ( (~ n34) ) | ( n740 ) ;
 assign n1199 = ( (~ n34) ) | ( n641 ) ;
 assign n1200 = ( (~ n34) ) | ( n324 ) ;
 assign n1201 = ( (~ n34)  &  (~ n616) ) | ( (~ n616)  &  n1189 ) | ( (~ n34)  &  n1192 ) | ( n1189  &  n1192 ) ;
 assign n1202 = ( n2387  &  n2348  &  n2230  &  n1417  &  n2351  &  n2135 ) ;
 assign n1197 = ( n1198  &  n1199  &  n1200  &  n1201  &  n1185  &  n1202 ) ;
 assign n1204 = ( (~ n34) ) | ( n1043 ) ;
 assign n1203 = ( (~ n34)  &  n1204 ) | ( n704  &  n1204 ) ;
 assign n1206 = ( n1347 ) | ( n1398 ) ;
 assign n1205 = ( n1206  &  n180  &  n800 ) ;
 assign n1207 = ( n400  &  (~ n706) ) | ( (~ n706)  &  n1021 ) ;
 assign n1208 = ( (~ n21) ) | ( n504 ) ;
 assign n1212 = ( n2269  &  n2304  &  n2060 ) ;
 assign n1210 = ( n412  &  n544 ) ;
 assign n1209 = ( (~ n21)  &  (~ n140)  &  n1212 ) | ( (~ n140)  &  n1212  &  n1210 ) ;
 assign n1214 = ( n1264  &  n1521 ) ;
 assign n1215 = ( n1372 ) | ( n1378 ) ;
 assign n1213 = ( n897  &  n707  &  n340  &  n1214  &  n1215 ) ;
 assign n1217 = ( (~ n17) ) | ( n1474 ) ;
 assign n1218 = ( (~ n17) ) | ( n468 ) ;
 assign n1219 = ( (~ n17)  &  (~ n21) ) | ( (~ n17)  &  n707 ) | ( (~ n21)  &  n1213 ) | ( n707  &  n1213 ) ;
 assign n1220 = ( n2093  &  n2372  &  n2547  &  n2439  &  n2448  &  n2124  &  n2339 ) ;
 assign n1216 = ( n416  &  n1217  &  n1218  &  n1219  &  n1209  &  n1220 ) ;
 assign n1222 = ( n1215  &  n187 ) ;
 assign n1221 = ( n501  &  n1210  &  n1222  &  (~ n1226) ) ;
 assign n1226 = ( (~ n561) ) | ( (~ n652) ) ;
 assign n1224 = ( (~ n412)  &  n616 ) | ( n616  &  (~ n897) ) | ( n616  &  n1226 ) ;
 assign n1227 = ( n340  &  (~ n1226) ) ;
 assign n1229 = ( (~ n139) ) | ( n1215 ) ;
 assign n1230 = ( (~ n139) ) | ( n340 ) ;
 assign n1231 = ( (~ n280) ) | ( n561 ) ;
 assign n1232 = ( (~ n360)  &  n1210 ) | ( n1210  &  n1227 ) | ( (~ n360)  &  n1426 ) | ( n1227  &  n1426 ) ;
 assign n1233 = ( (~ n132)  &  n1214 ) | ( (~ n21)  &  (~ n132)  &  (~ n616) ) ;
 assign n1234 = ( n1839  &  n1092  &  n1090  &  n1840  &  n2282  &  n2363  &  n1578  &  n1771 ) ;
 assign n1235 = ( n1095  &  n1064  &  n1829  &  n75  &  n1295  &  n1933  &  n1216  &  n2558 ) ;
 assign n1228 = ( n216  &  n1229  &  n1230  &  n1231  &  n1232  &  n1233  &  n1234  &  n1235 ) ;
 assign n1237 = ( n1314 ) | ( n1517 ) ;
 assign n1236 = ( n1237  &  n1122 ) ;
 assign n1239 = ( n39 ) | ( n248 ) ;
 assign n1238 = ( (~ n336)  &  (~ n810) ) | ( (~ n336)  &  (~ n812) ) | ( (~ n810)  &  n1239 ) | ( (~ n812)  &  n1239 ) ;
 assign n1240 = ( n332  &  (~ n737) ) | ( (~ n737)  &  n1021 ) ;
 assign n1242 = ( (~ n17) ) | ( n564 ) ;
 assign n1243 = ( (~ n17) ) | ( n1250 ) ;
 assign n1244 = ( (~ n17) ) | ( n921 ) ;
 assign n1245 = ( (~ n17)  &  n1985 ) | ( n953  &  n1352  &  n1985 ) ;
 assign n1246 = ( n2064  &  n2268  &  n2340  &  n2099  &  n2350  &  n2441  &  n2374  &  n547 ) ;
 assign n1241 = ( n415  &  n1242  &  n1243  &  n436  &  n458  &  n1244  &  n1245  &  n1246 ) ;
 assign n1248 = ( n1271  &  n1957  &  n1958 ) ;
 assign n1247 = ( (~ n616) ) | ( n1248 ) ;
 assign n1250 = ( (~ i_15_) ) | ( n1353 ) ;
 assign n1251 = ( n953  &  n921  &  n506 ) ;
 assign n1249 = ( n1250  &  n1077  &  n1251 ) ;
 assign n1253 = ( n536  &  n612 ) ;
 assign n1252 = ( n1253  &  n465  &  n564  &  n213 ) ;
 assign n1254 = ( n176  &  (~ n266)  &  (~ n476)  &  n563 ) ;
 assign n1257 = ( n959  &  n1260 ) ;
 assign n1258 = ( n1327 ) | ( n1347 ) ;
 assign n1256 = ( n1257  &  n711  &  n1258  &  n380 ) ;
 assign n1260 = ( n260  &  n1834  &  n1890  &  n812  &  n1265  &  n318 ) ;
 assign n1259 = ( n711  &  n740  &  n1260 ) ;
 assign n1262 = ( (~ n5)  &  n681  &  n799  &  n1280  &  n1352  &  n2039 ) ;
 assign n1261 = ( n1194  &  n778  &  n1262  &  n243  &  n508  &  n1045 ) ;
 assign n1264 = ( n1347 ) | ( n1390 ) ;
 assign n1265 = ( n1314 ) | ( n1347 ) ;
 assign n1263 = ( n323  &  n318  &  n344  &  n1264  &  n1265  &  n470 ) ;
 assign n1266 = ( n448  &  n799 ) ;
 assign n1269 = ( n1347 ) | ( n1391 ) ;
 assign n1270 = ( n262  &  n214  &  n288 ) ;
 assign n1271 = ( n1347 ) | ( n1370 ) ;
 assign n1272 = ( n1477  &  n1043  &  n1377 ) ;
 assign n1268 = ( n316  &  (~ n476)  &  n1060  &  n1061  &  n1269  &  n1270  &  n1271  &  n1272 ) ;
 assign n1274 = ( n345  &  n810 ) ;
 assign n1275 = ( n812  &  n1659 ) ;
 assign n1276 = ( n243  &  n824 ) ;
 assign n1277 = ( n524  &  n318  &  n743  &  n659  &  n1520  &  n1379 ) ;
 assign n1273 = ( n864  &  n1071  &  n1274  &  n1275  &  n1276  &  n1277 ) ;
 assign n1279 = ( n184  &  n193  &  (~ n266)  &  n327  &  n453  &  n1214  &  n2040  &  n2041 ) ;
 assign n1280 = ( n559  &  n1258  &  n852 ) ;
 assign n1278 = ( n180  &  n380  &  n950  &  n1279  &  n1280 ) ;
 assign n1282 = ( (~ n22)  &  n1996  &  n1998  &  n1999  &  n2000  &  n2001  &  n2002  &  n2003 ) ;
 assign n1283 = ( (~ n1159)  &  n1992  &  n1994  &  n1995 ) ;
 assign n1284 = ( n2020  &  n1208  &  n2021  &  n2022  &  n2023  &  n2024  &  n2025  &  n2026 ) ;
 assign n1285 = ( n1968  &  n1959  &  n1162 ) ;
 assign n1286 = ( (~ n17)  &  n572  &  n1949 ) | ( n572  &  n1268  &  n1949 ) ;
 assign n1287 = ( n2288  &  n2098  &  n457  &  n1400  &  n1401  &  n2375  &  n2602  &  n2601 ) ;
 assign n1281 = ( n1282  &  n1283  &  n1216  &  n1241  &  n1284  &  n1285  &  n1286  &  n1287 ) ;
 assign n1289 = ( n1478  &  n737 ) ;
 assign n1290 = ( n1369 ) | ( n1522 ) ;
 assign n1291 = ( n1379  &  n581  &  n214 ) ;
 assign n1292 = ( n2043  &  n2042  &  n1279  &  n1956  &  n1061  &  n1059  &  n1044  &  n1659 ) ;
 assign n1288 = ( n1289  &  n1206  &  n176  &  n1290  &  n541  &  n1012  &  n1291  &  n1292 ) ;
 assign n1294 = ( (~ n31)  &  n1978  &  n1979  &  n1980  &  n1981  &  n1983  &  n1984 ) ;
 assign n1295 = ( n1203  &  (~ n1224)  &  n2004  &  n2005  &  n2006  &  n2007  &  n2009  &  n2010 ) ;
 assign n1296 = ( n2036  &  n1536  &  n2037  &  n1247  &  n2027  &  n2038 ) ;
 assign n1297 = ( (~ n40)  &  n437  &  n2014  &  n2015  &  n2017  &  n2018  &  n2019 ) ;
 assign n1298 = ( n1952  &  n613  &  n1972 ) ;
 assign n1299 = ( (~ n616)  &  n2604 ) | ( n1288  &  n2604 ) ;
 assign n1300 = ( (~ n35)  &  n1402  &  n1556  &  n2121  &  n2136  &  n2603 ) ;
 assign n1293 = ( n1197  &  n1294  &  n1295  &  n1296  &  n1297  &  n1298  &  n1299  &  n1300 ) ;
 assign n1302 = ( (~ n10) ) | ( n815 ) ;
 assign n1303 = ( (~ n131) ) | ( n1484 ) ;
 assign n1304 = ( (~ n131) ) | ( n560 ) ;
 assign n1305 = ( (~ n131) ) | ( n292 ) ;
 assign n1306 = ( n1660  &  n1661  &  n644  &  n1662  &  n1663  &  n1664 ) ;
 assign n1307 = ( (~ n131) ) | ( n313  &  n778 ) ;
 assign n1308 = ( n2242  &  n2325  &  n2290  &  n2326  &  n2132  &  n2089  &  n2034  &  n2356 ) ;
 assign n1301 = ( n1302  &  n1303  &  n1304  &  n1305  &  n1306  &  n853  &  n1307  &  n1308 ) ;
 assign n1311 = ( i_11_ ) | ( (~ n981) ) ;
 assign n1314 = ( (~ i_15_) ) | ( n1311 ) ;
 assign n1315 = ( i_14_ ) | ( i_13_ ) | ( i_12_ ) ;
 assign n1316 = ( i_12_ ) | ( (~ i_13_) ) ;
 assign n1319 = ( i_11_ ) | ( (~ n980) ) ;
 assign n1321 = ( (~ i_15_) ) | ( n1319 ) ;
 assign n1323 = ( (~ i_9_) ) | ( (~ i_10_) ) ;
 assign n1322 = ( n1323  &  n1033 ) ;
 assign n1325 = ( i_12_ ) | ( i_13_ ) | ( (~ i_14_) ) ;
 assign n1326 = ( i_11_ ) | ( n516 ) ;
 assign n1327 = ( (~ i_15_) ) | ( n1326 ) ;
 assign n1329 = ( n1314 ) | ( n1315 ) ;
 assign n1330 = ( (~ i_12_) ) | ( n1311 ) ;
 assign n1331 = ( (~ i_11_) ) | ( (~ n981) ) ;
 assign n1332 = ( (~ i_12_) ) | ( n1319 ) ;
 assign n1328 = ( n1329  &  n1322  &  n1330  &  n213  &  n1331  &  n1332  &  n1325  &  n1316 ) ;
 assign n1336 = ( i_5_ ) | ( i_4_ ) | ( i_3_ ) ;
 assign n1337 = ( n152  &  (~ n1336) ) ;
 assign n1339 = ( (~ i_8_) ) | ( n887 ) ;
 assign n1341 = ( (~ i_3_)  &  (~ i_4_)  &  i_5_ ) ;
 assign n1343 = ( (~ i_3_)  &  i_4_  &  i_5_ ) ;
 assign n1344 = ( i_15_ ) | ( n1319 ) ;
 assign n1345 = ( n1319 ) | ( n1325 ) ;
 assign n1346 = ( i_15_ ) | ( n1311 ) ;
 assign n1347 = ( i_14_ ) | ( n1316 ) ;
 assign n1348 = ( (~ i_14_) ) | ( n1316 ) ;
 assign n1349 = ( n516  &  n1323 ) ;
 assign n1351 = ( n1311 ) | ( n1348 ) ;
 assign n1352 = ( n1321 ) | ( n1347 ) ;
 assign n1353 = ( n1319 ) | ( n1348 ) ;
 assign n1354 = ( n262  &  n1332  &  n1330  &  n1033  &  n1331  &  n263 ) ;
 assign n1350 = ( n810  &  n1265  &  n1351  &  n1352  &  n1353  &  n1354 ) ;
 assign n1355 = ( (~ i_8_)  &  n71 ) ;
 assign n1356 = ( i_3_ ) | ( (~ i_4_) ) | ( i_5_ ) ;
 assign n1357 = ( (~ n152) ) | ( n1356 ) ;
 assign n1359 = ( (~ n170)  &  (~ n1336) ) ;
 assign n1361 = ( i_8_ ) | ( (~ n47) ) ;
 assign n1362 = ( i_8_ ) | ( n887 ) ;
 assign n1364 = ( n1357 ) | ( n1361 ) ;
 assign n1363 = ( n1364  &  n491 ) ;
 assign n1365 = ( i_3_  &  (~ i_4_)  &  (~ i_5_) ) ;
 assign n1366 = ( n152  &  n151 ) ;
 assign n1367 = ( i_15_ ) | ( n1331 ) ;
 assign n1368 = ( (~ n170)  &  n1343 ) ;
 assign n1369 = ( i_15_ ) | ( n1326 ) ;
 assign n1370 = ( i_15_ ) | ( n1033 ) ;
 assign n1371 = ( (~ i_12_) ) | ( i_13_ ) ;
 assign n1372 = ( i_14_ ) | ( n1371 ) ;
 assign n1373 = ( (~ i_12_) ) | ( (~ i_13_) ) ;
 assign n1374 = ( i_14_ ) | ( n1373 ) ;
 assign n1375 = ( (~ i_15_) ) | ( n1033 ) ;
 assign n1376 = ( n1370 ) | ( n1374 ) ;
 assign n1377 = ( n1315 ) | ( n1375 ) ;
 assign n1378 = ( i_15_ ) | ( n1035 ) ;
 assign n1379 = ( n1315 ) | ( n1378 ) ;
 assign n1380 = ( i_6_ ) | ( (~ i_7_) ) ;
 assign n1381 = ( (~ i_8_)  &  (~ n1380) ) ;
 assign n1382 = ( (~ n170)  &  n1341 ) ;
 assign n1384 = ( (~ i_11_) ) | ( n1323 ) ;
 assign n1385 = ( i_15_ ) | ( n1384 ) ;
 assign n1388 = ( (~ n170)  &  (~ n1356) ) ;
 assign n1390 = ( (~ i_15_) ) | ( n1035 ) ;
 assign n1391 = ( (~ i_15_) ) | ( n1384 ) ;
 assign n1392 = ( (~ i_11_) ) | ( n516 ) ;
 assign n1393 = ( i_15_ ) | ( n1392 ) ;
 assign n1394 = ( n1347 ) | ( n1385 ) ;
 assign n1395 = ( n1367 ) | ( n1372 ) ;
 assign n1396 = ( (~ i_15_) ) | ( n1331 ) ;
 assign n1397 = ( i_8_  &  (~ n1380) ) ;
 assign n1398 = ( (~ i_15_) ) | ( n1392 ) ;
 assign n1400 = ( (~ n21) ) | ( n213 ) ;
 assign n1401 = ( (~ n21) ) | ( n214 ) ;
 assign n1402 = ( (~ n34) ) | ( n214 ) ;
 assign n1403 = ( n1995  &  n2134  &  n1980  &  n2135 ) ;
 assign n1404 = ( n2127  &  n2128  &  n2129  &  n2130  &  n2131  &  n2132  &  n1627  &  n2133 ) ;
 assign n1399 = ( n1400  &  n212  &  n1401  &  n1402  &  n1403  &  n1404 ) ;
 assign n1406 = ( (~ n10) ) | ( n1329 ) ;
 assign n1407 = ( (~ n10) ) | ( n508 ) ;
 assign n1405 = ( (~ n220)  &  n1406  &  n1407 ) ;
 assign n1412 = ( (~ n10) ) | ( n345 ) ;
 assign n1413 = ( (~ n247) ) | ( n342 ) ;
 assign n1414 = ( (~ n247) ) | ( n345 ) ;
 assign n1415 = ( (~ n10) ) | ( n318 ) ;
 assign n1416 = ( (~ n139) ) | ( n342 ) ;
 assign n1417 = ( (~ n34) ) | ( n1958 ) ;
 assign n1418 = ( n208  &  n210  &  (~ n217)  &  n1230  &  n1399  &  n2136 ) ;
 assign n1411 = ( n521  &  n1412  &  n1413  &  n1414  &  n1415  &  n1416  &  n1417  &  n1418 ) ;
 assign n1420 = ( (~ n139) ) | ( n316 ) ;
 assign n1421 = ( (~ n139) ) | ( n1376 ) ;
 assign n1422 = ( (~ n139) ) | ( n1377 ) ;
 assign n1419 = ( n1420  &  n1421  &  n1422 ) ;
 assign n1423 = ( (~ n280) ) | ( n316 ) ;
 assign n1424 = ( (~ n280) ) | ( n1377 ) ;
 assign n1425 = ( (~ n280) ) | ( n1376 ) ;
 assign n1426 = ( (~ n17)  &  (~ n135) ) ;
 assign n1427 = ( (~ n39)  &  (~ n280) ) ;
 assign n1428 = ( (~ n17)  &  (~ n21) ) ;
 assign n1431 = ( n1325 ) | ( n1385 ) ;
 assign n1432 = ( n1431  &  n544 ) ;
 assign n1433 = ( n292  &  n959 ) ;
 assign n1435 = ( n2083  &  n994 ) | ( n2083  &  n544 ) ;
 assign n1436 = ( n1913  &  n1908  &  n1807  &  n1950  &  n2082  &  n1998 ) ;
 assign n1437 = ( n1830  &  n1847  &  n1877  &  n1850  &  n2080  &  n2081  &  n1909  &  n2074 ) ;
 assign n1438 = ( n1634  &  n1714  &  n1628  &  n1783  &  n789  &  n2068  &  n791  &  n2066 ) ;
 assign n1439 = ( n1732  &  n1725  &  n2072  &  n1744  &  n1719  &  n2073  &  n1754  &  n2069 ) ;
 assign n1440 = ( n1970  &  n2060  &  n1955  &  n2061  &  n2001  &  n1999  &  n1987  &  n1951 ) ;
 assign n1441 = ( (~ n128)  &  n325  &  (~ n328)  &  n333  &  n1218  &  n2023  &  n2024  &  n2064 ) ;
 assign n1442 = ( n2051  &  n2052  &  n2053  &  n2054  &  n1080  &  n1115  &  n1895  &  n1897 ) ;
 assign n1443 = ( n1938  &  n1945  &  n2055  &  n1934  &  n2056  &  n2057  &  n2058  &  n2059 ) ;
 assign n1444 = ( n2045  &  n2046  &  n2047  &  n1861  &  n2048  &  n1828  &  n1654  &  n1657 ) ;
 assign n1445 = ( n2049  &  n1832  &  n1848  &  n1869  &  n2050  &  n1844  &  n1853  &  n1851 ) ;
 assign n1446 = ( n1701  &  n1706  &  n1601  &  n1661  &  n1639  &  n2044  &  n1625  &  n928 ) ;
 assign n1447 = ( n1722  &  n1756  &  n1727  &  n1726  &  n1748  &  n1745  &  n1693  &  n1684 ) ;
 assign n1448 = ( (~ n39)  &  (~ n300) ) ;
 assign n1449 = ( n313  &  n312  &  n665 ) ;
 assign n1450 = ( n263  &  n1449 ) ;
 assign n1452 = ( (~ n6) ) | ( n342 ) ;
 assign n1453 = ( (~ n131) ) | ( n342 ) ;
 assign n1454 = ( (~ n616) ) | ( n2612 ) ;
 assign n1455 = ( (~ n135)  &  n2065 ) | ( n342  &  n2065 ) ;
 assign n1451 = ( n1452  &  n1453  &  n1454  &  n1455 ) ;
 assign n1457 = ( (~ n21) ) | ( n176 ) ;
 assign n1459 = ( n2097  &  n2098  &  n1229  &  n2099 ) ;
 assign n1460 = ( n1994  &  n2093  &  n1109  &  n2094  &  n2095  &  n1930  &  n1082  &  n2096 ) ;
 assign n1461 = ( n1740  &  n1742  &  n1736  &  n1733  &  n1698  &  n2088  &  n1711  &  n2089 ) ;
 assign n1462 = ( n2090  &  n2091  &  n1048  &  n1023  &  n2092  &  n1710  &  n1792  &  n1758 ) ;
 assign n1464 = ( (~ n426) ) | ( n466 ) ;
 assign n1465 = ( n341 ) | ( (~ n426) ) ;
 assign n1466 = ( (~ n426) ) | ( n565 ) ;
 assign n1463 = ( n1464  &  n1465  &  n1466 ) ;
 assign n1468 = ( (~ n131) ) | ( n341 ) ;
 assign n1469 = ( (~ n131) ) | ( n565 ) ;
 assign n1470 = ( (~ n131) ) | ( n1394 ) ;
 assign n1467 = ( n1468  &  n1469  &  n1470 ) ;
 assign n1473 = ( n1348 ) | ( n1367 ) ;
 assign n1474 = ( n1374 ) | ( n1390 ) ;
 assign n1475 = ( n1348 ) | ( n1035 ) ;
 assign n1476 = ( n1327 ) | ( n1374 ) ;
 assign n1477 = ( n1372 ) | ( n1375 ) ;
 assign n1478 = ( i_15_ ) | ( n1351 ) ;
 assign n1479 = ( n1348 ) | ( n1385 ) ;
 assign n1480 = ( n1327 ) | ( n1372 ) ;
 assign n1482 = ( (~ n247) ) | ( n465 ) ;
 assign n1483 = ( (~ n6) ) | ( n1473 ) ;
 assign n1481 = ( n926  &  n1482  &  n923  &  n1483 ) ;
 assign n1484 = ( n1347 ) | ( n1396 ) ;
 assign n1485 = ( (~ n139) ) | ( n1269 ) ;
 assign n1486 = ( (~ n34) ) | ( n1269 ) ;
 assign n1487 = ( (~ n247) ) | ( n1269 ) ;
 assign n1488 = ( (~ n10) ) | ( n1352 ) ;
 assign n1490 = ( n1377  &  n788 ) ;
 assign n1491 = ( n1479  &  n412  &  n445 ) ;
 assign n1492 = ( n739  &  n1264 ) ;
 assign n1493 = ( (~ n135)  &  (~ n332) ) ;
 assign n1495 = ( (~ n247) ) | ( n506 ) ;
 assign n1496 = ( (~ n6) ) | ( n506 ) ;
 assign n1498 = ( (~ n247)  &  n469 ) | ( n469  &  n950  &  n1490 ) ;
 assign n1499 = ( (~ i_0_) ) | ( i_1_ ) ;
 assign n1500 = ( n1356 ) | ( n1499 ) ;
 assign n1502 = ( n1380 ) | ( n1500 ) ;
 assign n1503 = ( n887 ) | ( n1500 ) ;
 assign n1504 = ( (~ n71) ) | ( n1500 ) ;
 assign n1505 = ( (~ n47) ) | ( n1500 ) ;
 assign n1501 = ( n1502  &  n1503  &  n1504  &  n1505 ) ;
 assign n1506 = ( (~ n21)  &  n1399  &  n2226 ) | ( n530  &  n1399  &  n2226 ) ;
 assign n1507 = ( (~ n484)  &  (~ n486)  &  n2217  &  n2218  &  n2221  &  n2224 ) ;
 assign n1508 = ( n1892  &  n1464  &  n2215  &  n1953  &  n1424  &  n2216  &  n2206  &  n2210 ) ;
 assign n1509 = ( n669  &  n779  &  n1623  &  n2031  &  n1691  &  n2198  &  n2196  &  n2202 ) ;
 assign n1510 = ( n1336 ) | ( n1499 ) ;
 assign n1511 = ( n945  &  n965  &  n940  &  n963 ) ;
 assign n1513 = ( n959 ) | ( (~ n978) ) ;
 assign n1514 = ( (~ n978) ) | ( n1329 ) ;
 assign n1515 = ( (~ n1337) ) | ( n1380 ) ;
 assign n1516 = ( n1779  &  n1788  &  n2321  &  n1777  &  n935  &  n968 ) ;
 assign n1512 = ( n901  &  n1513  &  n1514  &  n1515  &  n514  &  n1516 ) ;
 assign n1517 = ( (~ i_14_) ) | ( n1371 ) ;
 assign n1518 = ( n1375 ) | ( n1517 ) ;
 assign n1519 = ( n1327 ) | ( n1517 ) ;
 assign n1520 = ( n1344 ) | ( n1517 ) ;
 assign n1521 = ( n1378 ) | ( n1517 ) ;
 assign n1522 = ( (~ i_14_) ) | ( n1373 ) ;
 assign n1523 = ( n1385 ) | ( n1522 ) ;
 assign n1524 = ( n1191  &  n726 ) ;
 assign n1525 = ( n1381  &  n1382 ) ;
 assign n1526 = ( n567  &  n576 ) ;
 assign n1527 = ( n1473  &  n292 ) ;
 assign n1528 = ( n564  &  n706 ) ;
 assign n1529 = ( n915  &  n908  &  n200  &  n916 ) ;
 assign n1531 = ( (~ n6) ) | ( n1290 ) ;
 assign n1532 = ( (~ n6) ) | ( n453 ) ;
 assign n1533 = ( (~ n6) ) | ( n1012 ) ;
 assign n1530 = ( n1531  &  n1532  &  n1533 ) ;
 assign n1534 = ( n1382  &  n1397 ) ;
 assign n1535 = ( (~ n21) ) | ( n1290 ) ;
 assign n1536 = ( (~ n34) ) | ( n1077 ) ;
 assign n1537 = ( (~ n136)  &  (~ n280)  &  n2018 ) | ( (~ n136)  &  n556  &  n2018 ) ;
 assign n1538 = ( n2374  &  n1102  &  n2375  &  n1818  &  n1819  &  n2376 ) ;
 assign n1539 = ( n1996  &  n1814  &  n1816  &  n1923  &  n2371  &  n1960 ) ;
 assign n1540 = ( n1971  &  n2372  &  n2021  &  n1978  &  n2373  &  n1926 ) ;
 assign n1541 = ( n2366  &  n2367  &  n2368  &  n2369  &  n2370  &  n1090  &  n2362  &  n2358 ) ;
 assign n1543 = ( (~ n139) ) | ( n576 ) ;
 assign n1542 = ( n1543  &  n405  &  n429 ) ;
 assign n1545 = ( (~ n10) ) | ( n953 ) ;
 assign n1544 = ( n431  &  n1545  &  n407 ) ;
 assign n1547 = ( (~ n280) ) | ( n544 ) ;
 assign n1546 = ( n1547  &  n406  &  n430 ) ;
 assign n1548 = ( (~ n247) ) | ( n564 ) ;
 assign n1549 = ( (~ n6) ) | ( n541 ) ;
 assign n1550 = ( n470  &  n702 ) ;
 assign n1551 = ( n1520  &  n1521 ) ;
 assign n1552 = ( n706  &  n176  &  n993  &  n559 ) ;
 assign n1553 = ( n1237  &  n566  &  n1077  &  n641  &  n561 ) ;
 assign n1554 = ( n611  &  n530  &  n1250  &  n743  &  n740 ) ;
 assign n1556 = ( (~ n616) ) | ( n2613 ) ;
 assign n1558 = ( n508  &  n2343 ) | ( (~ n616)  &  n2343 ) ;
 assign n1555 = ( n404  &  n613  &  (~ n614)  &  n1093  &  n1099  &  n1546  &  n1556  &  n1558 ) ;
 assign n1560 = ( (~ n280)  &  n1542  &  n2352 ) | ( n953  &  n1542  &  n2352 ) ;
 assign n1561 = ( n2348  &  n1928  &  n2349  &  n2017  &  n2350  &  n1983  &  n2351  &  n2344 ) ;
 assign n1559 = ( n605  &  n603  &  n1544  &  n607  &  n1560  &  n1561 ) ;
 assign n1562 = ( n659  &  n566 ) ;
 assign n1563 = ( n611  &  (~ n1226) ) ;
 assign n1564 = ( n1327 ) | ( n1522 ) ;
 assign n1565 = ( n541  &  n313 ) ;
 assign n1567 = ( (~ n280) ) | ( n524 ) ;
 assign n1566 = ( n1567  &  n1149  &  n582 ) ;
 assign n1569 = ( (~ n10) ) | ( n740 ) ;
 assign n1568 = ( n1569  &  n674 ) ;
 assign n1570 = ( (~ n6) ) | ( n536 ) ;
 assign n1571 = ( (~ n6) ) | ( n537 ) ;
 assign n1572 = ( (~ n247) ) | ( n536 ) ;
 assign n1573 = ( (~ n247) ) | ( n537 ) ;
 assign n1574 = ( (~ n247) ) | ( n524 ) ;
 assign n1575 = ( (~ n247) ) | ( n1518 ) ;
 assign n1576 = ( n854  &  n812 ) ;
 assign n1578 = ( n1431 ) | ( n545 ) ;
 assign n1579 = ( (~ n1019) ) | ( n1518 ) ;
 assign n1581 = ( n536  &  n545 ) | ( n536  &  n576 ) | ( n545  &  (~ n1019) ) | ( n576  &  (~ n1019) ) ;
 assign n1577 = ( n729  &  (~ n732)  &  n1578  &  n1579  &  n1581 ) ;
 assign n1583 = ( (~ n6) ) | ( n864 ) ;
 assign n1584 = ( (~ n6) ) | ( n707 ) ;
 assign n1585 = ( (~ n131) ) | ( n1824 ) ;
 assign n1586 = ( n336  &  (~ n357) ) | ( n336  &  n707 ) | ( (~ n357)  &  n864 ) | ( n707  &  n864 ) ;
 assign n1582 = ( n816  &  n1583  &  n1584  &  n1585  &  n701  &  n697  &  n694  &  n1586 ) ;
 assign n1588 = ( (~ n139) ) | ( n524 ) ;
 assign n1587 = ( n1588  &  n658 ) ;
 assign n1589 = ( (~ n1343) ) | ( n1499 ) ;
 assign n1592 = ( n1380 ) | ( n1589 ) ;
 assign n1593 = ( (~ n47) ) | ( n1589 ) ;
 assign n1594 = ( n887 ) | ( n1589 ) ;
 assign n1591 = ( n1592  &  n1593  &  n1594 ) ;
 assign n1596 = ( n213  &  n953  &  n508 ) ;
 assign n1598 = ( (~ n247) ) | ( n854 ) ;
 assign n1599 = ( (~ n247) ) | ( n560 ) ;
 assign n1600 = ( (~ n247) ) | ( n1484 ) ;
 assign n1597 = ( n1598  &  n1599  &  n1600 ) ;
 assign n1601 = ( (~ n6) ) | ( n897 ) ;
 assign n1602 = ( (~ n247) ) | ( n704 ) ;
 assign n1603 = ( (~ n247) ) | ( n1043 ) ;
 assign n1604 = ( n1597  &  n777 ) ;
 assign n1605 = ( n781  &  n1604  &  n936  &  n931 ) ;
 assign n1608 = ( n2044  &  n2355  &  n2068  &  n2244  &  n2323  &  n2245  &  n2131  &  n2324 ) ;
 assign n1606 = ( (~ n125)  &  n183  &  n208  &  n383  &  n603  &  n792  &  n795  &  n1608 ) ;
 assign n1609 = ( (~ n247) ) | ( n1258 ) ;
 assign n1610 = ( (~ n247) ) | ( n1009 ) ;
 assign n1611 = ( (~ n6) ) | ( n1352 ) ;
 assign n1612 = ( (~ n247) ) | ( n839 ) ;
 assign n1613 = ( (~ n6) ) | ( n581 ) ;
 assign n1614 = ( (~ n6) ) | ( n1206 ) ;
 assign n1615 = ( (~ n247) ) | ( n581 ) ;
 assign n1616 = ( (~ n247) ) | ( n1206 ) ;
 assign n1617 = ( (~ n247) ) | ( n800 ) ;
 assign n1618 = ( (~ n247) ) | ( n812 ) ;
 assign n1619 = ( (~ n247) ) | ( n993 ) ;
 assign n1620 = ( (~ n6) ) | ( n993 ) ;
 assign n1621 = ( (~ n6) ) | ( n1265 ) ;
 assign n1622 = ( (~ n247) ) | ( n1265 ) ;
 assign n1623 = ( (~ n6) ) | ( n1269 ) ;
 assign n1624 = ( n160  &  (~ n1362) ) ;
 assign n1625 = ( (~ n6) ) | ( n243 ) ;
 assign n1626 = ( (~ n247) ) | ( n243 ) ;
 assign n1627 = ( (~ n247) ) | ( n1394 ) ;
 assign n1628 = ( (~ n6) ) | ( n292 ) ;
 assign n1630 = ( (~ n247) ) | ( n707 ) ;
 assign n1631 = ( (~ n247) ) | ( n1521 ) ;
 assign n1632 = ( (~ n6) ) | ( n564 ) ;
 assign n1633 = ( (~ n6) ) | ( n465 ) ;
 assign n1634 = ( (~ n6) ) | ( n953 ) ;
 assign n1629 = ( n1630  &  n1631  &  n836  &  n1632  &  n1633  &  n1634 ) ;
 assign n1635 = ( (~ n6) ) | ( n524 ) ;
 assign n1637 = ( (~ n6) ) | ( n464 ) ;
 assign n1638 = ( (~ n6) ) | ( n1518 ) ;
 assign n1639 = ( (~ n6) ) | ( n1271 ) ;
 assign n1640 = ( (~ n6) ) | ( n568 ) ;
 assign n1641 = ( (~ n6) ) | ( n566 ) ;
 assign n1642 = ( (~ n6) ) | ( n567 ) ;
 assign n1644 = ( (~ n247) ) | ( n1264 ) ;
 assign n1645 = ( (~ n247) ) | ( n1379 ) ;
 assign n1646 = ( (~ n247) ) | ( n612 ) ;
 assign n1647 = ( (~ n6) ) | ( n1264 ) ;
 assign n1648 = ( (~ n6) ) | ( n1379 ) ;
 assign n1643 = ( n1644  &  n1645  &  n1646  &  n384  &  n1647  &  n1648  &  n831 ) ;
 assign n1649 = ( (~ n10) ) | ( n704 ) ;
 assign n1650 = ( (~ n10) ) | ( n1043 ) ;
 assign n1651 = ( (~ n10) ) | ( n1269 ) ;
 assign n1653 = ( (~ n131) ) | ( n413 ) ;
 assign n1654 = ( (~ n131) ) | ( n468 ) ;
 assign n1655 = ( (~ n131) ) | ( n340 ) ;
 assign n1656 = ( (~ n131) ) | ( n1215 ) ;
 assign n1657 = ( (~ n131) ) | ( n897 ) ;
 assign n1652 = ( n1653  &  n1654  &  n1655  &  n1656  &  n1657 ) ;
 assign n1658 = ( n345  &  n1520 ) ;
 assign n1659 = ( n1265  &  n993 ) ;
 assign n1660 = ( (~ n10) ) | ( n766 ) ;
 assign n1661 = ( (~ n10) ) | ( n466 ) ;
 assign n1662 = ( (~ n10) ) | ( n1479 ) ;
 assign n1663 = ( (~ n10) ) | ( n1431 ) ;
 assign n1664 = ( (~ n10) ) | ( n709 ) ;
 assign n1666 = ( (~ n10) ) | ( n707 ) ;
 assign n1667 = ( (~ n131) ) | ( n1264 ) ;
 assign n1668 = ( (~ n131) ) | ( n1379 ) ;
 assign n1665 = ( n1666  &  n1667  &  n1668 ) ;
 assign n1671 = ( (~ n10) ) | ( n1275 ) ;
 assign n1669 = ( n549  &  (~ n859)  &  n862  &  n1671 ) ;
 assign n1673 = ( (~ n10) ) | ( n864 ) ;
 assign n1674 = ( (~ n10) ) | ( n1520 ) ;
 assign n1672 = ( (~ n857)  &  n1673  &  n1674 ) ;
 assign n1677 = ( (~ n131) ) | ( n612 ) ;
 assign n1678 = ( (~ n131) ) | ( n412 ) ;
 assign n1679 = ( (~ n131) ) | ( n544 ) ;
 assign n1680 = ( (~ n131) ) | ( n1474 ) ;
 assign n1676 = ( n1677  &  n1678  &  n1679  &  n1680  &  n655 ) ;
 assign n1682 = ( (~ n131) ) | ( n1077 ) ;
 assign n1683 = ( (~ n131) ) | ( n506 ) ;
 assign n1684 = ( (~ n131) ) | ( n213 ) ;
 assign n1685 = ( (~ n131) ) | ( n288 ) ;
 assign n1686 = ( (~ n131) ) | ( n2608 ) ;
 assign n1681 = ( n1682  &  n1683  &  n1684  &  n1685  &  n1686 ) ;
 assign n1688 = ( (~ n247) ) | ( n1564 ) ;
 assign n1689 = ( (~ n247) ) | ( n559 ) ;
 assign n1690 = ( (~ n6) ) | ( n559 ) ;
 assign n1691 = ( (~ n6) ) | ( n1258 ) ;
 assign n1687 = ( n1688  &  n1689  &  n851  &  n1414  &  n1690  &  n1691 ) ;
 assign n1692 = ( (~ n131) ) | ( n766 ) ;
 assign n1693 = ( (~ n131) ) | ( n466 ) ;
 assign n1694 = ( (~ n131) ) | ( n1431 ) ;
 assign n1695 = ( (~ n131) ) | ( n709 ) ;
 assign n1696 = ( (~ n131) ) | ( n536 ) ;
 assign n1697 = ( (~ n131) ) | ( n1479 ) ;
 assign n1698 = ( (~ n10) ) | ( n1395 ) ;
 assign n1699 = ( (~ n10) ) | ( n507 ) ;
 assign n1700 = ( (~ n10) ) | ( n193 ) ;
 assign n1701 = ( (~ n131) ) | ( n193 ) ;
 assign n1702 = ( (~ n131) ) | ( n190 ) ;
 assign n1703 = ( (~ n131) ) | ( n470 ) ;
 assign n1704 = ( (~ n131) ) | ( n507 ) ;
 assign n1705 = ( (~ n131) ) | ( n1395 ) ;
 assign n1706 = ( (~ n131) ) | ( n243 ) ;
 assign n1707 = ( (~ n10) ) | ( n1122 ) ;
 assign n1709 = ( (~ n10) ) | ( n506 ) ;
 assign n1710 = ( (~ n10) ) | ( n288 ) ;
 assign n1708 = ( n1709  &  n1710  &  n1544 ) ;
 assign n1711 = ( (~ n247) ) | ( n726 ) ;
 assign n1712 = ( (~ n247) ) | ( n706 ) ;
 assign n1713 = ( (~ n247) ) | ( n1191 ) ;
 assign n1714 = ( (~ n6) ) | ( n726 ) ;
 assign n1715 = ( (~ n6) ) | ( n2605 ) ;
 assign n1716 = ( (~ n6) ) | ( n706 ) ;
 assign n1717 = ( (~ n6) ) | ( n1191 ) ;
 assign n1719 = ( (~ n10) ) | ( n544 ) ;
 assign n1720 = ( (~ n10) ) | ( n1474 ) ;
 assign n1721 = ( (~ n10) ) | ( n413 ) ;
 assign n1722 = ( (~ n10) ) | ( n468 ) ;
 assign n1723 = ( (~ n10) ) | ( n340 ) ;
 assign n1718 = ( n1719  &  n1720  &  n1721  &  n1722  &  n1723 ) ;
 assign n1725 = ( (~ n131) ) | ( n316 ) ;
 assign n1726 = ( (~ n131) ) | ( n1271 ) ;
 assign n1727 = ( (~ n131) ) | ( n1377 ) ;
 assign n1728 = ( (~ n131) ) | ( n1376 ) ;
 assign n1729 = ( (~ n131) ) | ( n743 ) ;
 assign n1730 = ( (~ n131) ) | ( n1477 ) ;
 assign n1731 = ( (~ n131) ) | ( n567 ) ;
 assign n1732 = ( (~ n131) ) | ( n576 ) ;
 assign n1724 = ( n1725  &  n1726  &  n1727  &  n1728  &  n1729  &  n1730  &  n1731  &  n1732 ) ;
 assign n1733 = ( (~ n10) ) | ( n316 ) ;
 assign n1734 = ( (~ n10) ) | ( n1477 ) ;
 assign n1735 = ( (~ n10) ) | ( n567 ) ;
 assign n1736 = ( (~ n10) ) | ( n576 ) ;
 assign n1738 = ( (~ n10) ) | ( n505 ) ;
 assign n1739 = ( (~ n10) ) | ( n1191 ) ;
 assign n1740 = ( (~ n10) ) | ( n726 ) ;
 assign n1741 = ( (~ n10) ) | ( n373 ) ;
 assign n1742 = ( (~ n10) ) | ( n291 ) ;
 assign n1737 = ( n386  &  n1738  &  n1739  &  n1740  &  n1741  &  n235  &  n1742 ) ;
 assign n1744 = ( (~ n131) ) | ( n291 ) ;
 assign n1745 = ( (~ n131) ) | ( n324 ) ;
 assign n1746 = ( (~ n10) ) | ( n641 ) ;
 assign n1747 = ( (~ n131) ) | ( n505 ) ;
 assign n1748 = ( (~ n131) ) | ( n373 ) ;
 assign n1749 = ( (~ n131) ) | ( n180 ) ;
 assign n1750 = ( n2243  &  n2072  &  n2294  &  n2327  &  n2292  &  n2331 ) ;
 assign n1743 = ( n1744  &  n1745  &  n1746  &  n1747  &  n1748  &  n1749  &  n1750 ) ;
 assign n1752 = ( (~ n3)  &  n174  &  n1530  &  n2185  &  n2197  &  n2357 ) ;
 assign n1751 = ( n664  &  n694  &  n1629  &  n1153  &  n1643  &  n1752 ) ;
 assign n1754 = ( (~ n131) ) | ( n1071 ) ;
 assign n1755 = ( (~ n10) ) | ( n1478 ) ;
 assign n1756 = ( (~ n131) ) | ( n1329 ) ;
 assign n1757 = ( (~ n131) ) | ( n261 ) ;
 assign n1758 = ( (~ n10) ) | ( n959 ) ;
 assign n1759 = ( (~ n10) ) | ( n381 ) ;
 assign n1760 = ( (~ n10) ) | ( n768 ) ;
 assign n1761 = ( n2329  &  n2248  &  n2330  &  n2293  &  n2073  &  n2295  &  n2247 ) ;
 assign n1753 = ( n1754  &  n1755  &  n1756  &  n1757  &  n1758  &  n1759  &  n1760  &  n1761 ) ;
 assign n1762 = ( n152  &  n150 ) ;
 assign n1763 = ( n825  &  n820  &  n1751  &  n1753 ) ;
 assign n1764 = ( n905  &  n1718  &  n874  &  n906  &  n643  &  n1708  &  n651  &  n2500 ) ;
 assign n1765 = ( n918  &  n2359  &  n1792  &  n1790  &  n1791  &  n1786  &  n2495  &  n2497 ) ;
 assign n1766 = ( n939  &  n1501  &  n493  &  n1591  &  n756 ) ;
 assign n1767 = ( n1329 ) | ( (~ n1624) ) ;
 assign n1768 = ( n214 ) | ( (~ n1624) ) ;
 assign n1769 = ( n959 ) | ( (~ n1624) ) ;
 assign n1771 = ( (~ n6) ) | ( n1521 ) ;
 assign n1770 = ( n1771  &  n932  &  n811 ) ;
 assign n1772 = ( n934  &  n1605 ) ;
 assign n1774 = ( n776 ) | ( n49 ) | ( n893 ) | ( n164 ) ;
 assign n1776 = ( n897 ) | ( n491 ) ;
 assign n1777 = ( n897 ) | ( (~ n978) ) ;
 assign n1775 = ( n1776  &  n896  &  n1777  &  n758 ) ;
 assign n1779 = ( n214 ) | ( (~ n978) ) ;
 assign n1780 = ( n214 ) | ( n491 ) ;
 assign n1778 = ( n772  &  n757  &  n894  &  n1779  &  n1768  &  n1780 ) ;
 assign n1783 = ( (~ n247) ) | ( n953 ) ;
 assign n1781 = ( n197  &  (~ n919)  &  n1482  &  n1495  &  n1548  &  n1783 ) ;
 assign n1784 = ( n1624 ) | ( n893 ) | ( n979 ) ;
 assign n1786 = ( (~ n10) ) | ( n412 ) ;
 assign n1785 = ( n1786  &  n651  &  n1718 ) ;
 assign n1788 = ( n953 ) | ( (~ n978) ) ;
 assign n1787 = ( n761  &  n952  &  n1788  &  n1504 ) ;
 assign n1790 = ( (~ n10) ) | ( n897 ) ;
 assign n1791 = ( (~ n10) ) | ( n612 ) ;
 assign n1792 = ( (~ n10) ) | ( n1215 ) ;
 assign n1789 = ( n1790  &  n1785  &  n1791  &  n1792 ) ;
 assign n1793 = ( n686  &  n1753  &  n532  &  n531 ) ;
 assign n1794 = ( n1737  &  n1743  &  n245  &  n1568 ) ;
 assign n1796 = ( n718  &  n2141  &  n210  &  n1549  &  n1483  &  n719 ) ;
 assign n1795 = ( n826  &  n949  &  n946  &  n192  &  n469  &  n713  &  n1796 ) ;
 assign n1797 = ( n1513  &  n1593  &  n1769  &  n1505  &  n760 ) ;
 assign n1799 = ( n321  &  n671  &  n525  &  n920  &  n1496  &  n2359  &  n720  &  n2228 ) ;
 assign n1798 = ( n878  &  n1708  &  n722  &  n781  &  n1781  &  n917  &  n914  &  n1799 ) ;
 assign n1800 = ( n1751  &  n801  &  n902 ) ;
 assign n1801 = ( (~ n71) ) | ( n1357 ) ;
 assign n1802 = ( (~ n516)  &  (~ n1339)  &  n1366 ) ;
 assign n1803 = ( n152  &  (~ n516)  &  (~ n1339)  &  n1365 ) ;
 assign n1804 = ( n1778  &  n1787  &  n969 ) ;
 assign n1805 = ( n1376  &  n659 ) ;
 assign n1806 = ( n994 ) | ( n561 ) ;
 assign n1807 = ( n1215 ) | ( n994 ) ;
 assign n1809 = ( n990 ) | ( n1521 ) ;
 assign n1810 = ( n994 ) | ( n1521 ) ;
 assign n1811 = ( n994 ) | ( n612 ) ;
 assign n1812 = ( n990 ) | ( n448 ) ;
 assign n1814 = ( n990 ) | ( n641 ) ;
 assign n1815 = ( n990 ) | ( n740 ) ;
 assign n1816 = ( n990 ) | ( n706 ) ;
 assign n1817 = ( n990 ) | ( n993 ) ;
 assign n1818 = ( n990 ) | ( n1237 ) ;
 assign n1819 = ( n990 ) | ( n737 ) ;
 assign n1820 = ( n544  &  n576 ) ;
 assign n1821 = ( n1519  &  n1237 ) ;
 assign n1822 = ( n341  &  n1431 ) ;
 assign n1823 = ( n1822  &  n1141 ) ;
 assign n1824 = ( n1250  &  n711 ) ;
 assign n1826 = ( (~ n280) ) | ( n565 ) ;
 assign n1827 = ( (~ n280) ) | ( n766 ) ;
 assign n1828 = ( (~ n280) ) | ( n466 ) ;
 assign n1825 = ( n1826  &  n1041  &  n1827  &  n1828 ) ;
 assign n1830 = ( (~ n280) ) | ( n1215 ) ;
 assign n1831 = ( (~ n280) ) | ( n412 ) ;
 assign n1832 = ( (~ n280) ) | ( n468 ) ;
 assign n1833 = ( (~ n280) ) | ( n340 ) ;
 assign n1829 = ( n1830  &  n1831  &  n1832  &  n1833  &  n1546 ) ;
 assign n1834 = ( n581  &  n263  &  n261  &  n799  &  n1206 ) ;
 assign n1835 = ( n176  &  (~ n266)  &  n323  &  n1280 ) ;
 assign n1836 = ( n959  &  n380  &  n800  &  n1835  &  n1057 ) ;
 assign n1838 = ( (~ n280) ) | ( n1477 ) ;
 assign n1839 = ( (~ n280) ) | ( n652 ) ;
 assign n1840 = ( (~ n280) ) | ( n897 ) ;
 assign n1841 = ( (~ n280) ) | ( n568 ) ;
 assign n1842 = ( n2110  &  n2363  &  n2282 ) ;
 assign n1837 = ( n1838  &  n1839  &  n1231  &  n1154  &  n1829  &  n1840  &  n1841  &  n1842 ) ;
 assign n1843 = ( (~ n135) ) | ( n413 ) ;
 assign n1844 = ( (~ n135) ) | ( n468 ) ;
 assign n1845 = ( (~ n135) ) | ( n611 ) ;
 assign n1846 = ( (~ n135) ) | ( n612 ) ;
 assign n1847 = ( (~ n135) ) | ( n1215 ) ;
 assign n1848 = ( (~ n135) ) | ( n897 ) ;
 assign n1849 = ( (~ n135) ) | ( n1957 ) ;
 assign n1850 = ( (~ n135) ) | ( n316 ) ;
 assign n1851 = ( (~ n135) ) | ( n1271 ) ;
 assign n1852 = ( (~ n135) ) | ( n567 ) ;
 assign n1853 = ( (~ n135) ) | ( n1377 ) ;
 assign n1854 = ( (~ n135) ) | ( n1518 ) ;
 assign n1855 = ( (~ n135) ) | ( n524 ) ;
 assign n1856 = ( (~ n135) ) | ( n1269 ) ;
 assign n1857 = ( n1384 ) | ( (~ n1525) ) ;
 assign n1858 = ( (~ n280) ) | ( n536 ) ;
 assign n1859 = ( (~ n280) ) | ( n537 ) ;
 assign n1860 = ( (~ n135) ) | ( n766 ) ;
 assign n1861 = ( (~ n135) ) | ( n466 ) ;
 assign n1862 = ( (~ n135) ) | ( n565 ) ;
 assign n1863 = ( n2229  &  n2143  &  n1029  &  n2045  &  n2435  &  n2381 ) ;
 assign n1864 = ( (~ n135) ) | ( n262 ) ;
 assign n1865 = ( (~ n135) ) | ( n564 ) ;
 assign n1866 = ( (~ n135) ) | ( n1077 ) ;
 assign n1867 = ( (~ n135) ) | ( n1250 ) ;
 assign n1868 = ( (~ n135) ) | ( n506 ) ;
 assign n1869 = ( (~ n135) ) | ( n213 ) ;
 assign n1870 = ( (~ n135) ) | ( n318 ) ;
 assign n1871 = ( n2254  &  n2070  &  n2071  &  n2048  &  n2302  &  n2404  &  n2203 ) ;
 assign n1873 = ( (~ n280) ) | ( n505 ) ;
 assign n1874 = ( (~ n280) ) | ( n373 ) ;
 assign n1876 = ( n1392  &  n2520 ) | ( (~ n1534)  &  n2520 ) ;
 assign n1877 = ( (~ n135) ) | ( n291 ) ;
 assign n1878 = ( (~ n280) ) | ( n641 ) ;
 assign n1879 = ( (~ n280) ) | ( n448 ) ;
 assign n1880 = ( n2253  &  n2046  &  n2108  &  n2332 ) ;
 assign n1872 = ( (~ n1020)  &  n1873  &  n1874  &  n1876  &  n1877  &  n1878  &  n1879  &  n1880 ) ;
 assign n1881 = ( (~ n280) ) | ( n743 ) ;
 assign n1883 = ( (~ n280) ) | ( n837 ) ;
 assign n1884 = ( (~ n280) ) | ( n1518 ) ;
 assign n1885 = ( (~ n280) ) | ( n464 ) ;
 assign n1882 = ( n1883  &  n690  &  n1884  &  n1885 ) ;
 assign n1887 = ( (~ n280) ) | ( n1379 ) ;
 assign n1888 = ( (~ n280) ) | ( n1521 ) ;
 assign n1889 = ( (~ n280) ) | ( n1264 ) ;
 assign n1886 = ( n1887  &  n688  &  n1888  &  n1889 ) ;
 assign n1890 = ( n800  &  n1274 ) ;
 assign n1892 = ( (~ n39) ) | ( n2605 ) ;
 assign n1893 = ( (~ n39) ) | ( n641 ) ;
 assign n1894 = ( (~ n39) ) | ( n740 ) ;
 assign n1895 = ( (~ n39) ) | ( n324 ) ;
 assign n1896 = ( (~ n39) ) | ( n2610 ) ;
 assign n1897 = ( (~ n39) ) | ( n508 ) ;
 assign n1898 = ( (~ n39) ) | ( n993 ) ;
 assign n1899 = ( (~ n39) ) | ( n737 ) ;
 assign n1900 = ( (~ n39) ) | ( n1478 ) ;
 assign n1901 = ( (~ n39) ) | ( n1237 ) ;
 assign n1902 = ( (~ n39) ) | ( n530 ) ;
 assign n1903 = ( (~ n139) ) | ( n561 ) ;
 assign n1904 = ( (~ n139) ) | ( n412 ) ;
 assign n1905 = ( (~ n426) ) | ( n709 ) ;
 assign n1906 = ( (~ n426) ) | ( n766 ) ;
 assign n1907 = ( (~ n426) ) | ( n1479 ) ;
 assign n1908 = ( (~ n426) ) | ( n1431 ) ;
 assign n1909 = ( (~ n139) ) | ( n1395 ) ;
 assign n1910 = ( (~ n139) ) | ( n313 ) ;
 assign n1911 = ( (~ n139) ) | ( n541 ) ;
 assign n1912 = ( (~ n139) ) | ( n1473 ) ;
 assign n1913 = ( (~ n139) ) | ( n292 ) ;
 assign n1914 = ( n2061  &  n270  &  n2307  &  n2270 ) ;
 assign n1916 = ( n1519  &  n291  &  n324 ) ;
 assign n1915 = ( (~ n476)  &  n504  &  n563  &  n1251  &  n1526  &  n1553  &  n1554  &  n1916 ) ;
 assign n1918 = ( (~ n426) ) | ( n1043 ) ;
 assign n1919 = ( (~ n426) ) | ( n704 ) ;
 assign n1920 = ( (~ n139) ) | ( n537 ) ;
 assign n1921 = ( (~ n139) ) | ( n704 ) ;
 assign n1922 = ( (~ n139) ) | ( n1043 ) ;
 assign n1923 = ( (~ n139) ) | ( n536 ) ;
 assign n1924 = ( n2208  &  n2151 ) ;
 assign n1917 = ( n1918  &  n1463  &  n1919  &  n1920  &  n1921  &  n1922  &  n1923  &  n1924 ) ;
 assign n1926 = ( (~ n139) ) | ( n641 ) ;
 assign n1927 = ( (~ n139) ) | ( n740 ) ;
 assign n1928 = ( (~ n139) ) | ( n1193 ) ;
 assign n1929 = ( (~ n139) ) | ( n373 ) ;
 assign n1930 = ( (~ n139) ) | ( n291 ) ;
 assign n1931 = ( (~ n139) ) | ( n324 ) ;
 assign n1932 = ( n2256  &  n2058  &  n2194  &  n2257  &  n2078  &  n2297 ) ;
 assign n1925 = ( n1926  &  n1927  &  n1928  &  n1929  &  n1930  &  n1931  &  n1932 ) ;
 assign n1934 = ( (~ n426) ) | ( n468 ) ;
 assign n1935 = ( (~ n426) ) | ( n1215 ) ;
 assign n1936 = ( (~ n426) ) | ( n1474 ) ;
 assign n1937 = ( n413 ) | ( (~ n426) ) ;
 assign n1938 = ( (~ n426) ) | ( n897 ) ;
 assign n1939 = ( n2265  &  n2076  &  n2388  &  n2334  &  n2233  &  n2145  &  n2113  &  n2434 ) ;
 assign n1933 = ( n1934  &  n1935  &  n1936  &  n1937  &  n1938  &  n1105  &  n1886  &  n1939 ) ;
 assign n1941 = ( (~ n426) ) | ( n524 ) ;
 assign n1942 = ( n2056  &  n2412  &  n2216 ) ;
 assign n1943 = ( n2432  &  n2335  &  n2264  &  n2059  &  n2079  &  n2234  &  n2146  &  n2529 ) ;
 assign n1940 = ( n658  &  n1882  &  n1419  &  n1542  &  n1094  &  n1941  &  n1942  &  n1943 ) ;
 assign n1945 = ( (~ n21) ) | ( n466 ) ;
 assign n1947 = ( (~ n21) ) | ( n709 ) ;
 assign n1948 = ( (~ n21) ) | ( n766 ) ;
 assign n1944 = ( (~ n1142)  &  n1945  &  n1947  &  n1948 ) ;
 assign n1950 = ( (~ n17) ) | ( n565 ) ;
 assign n1951 = ( (~ n17) ) | ( n1394 ) ;
 assign n1949 = ( n1950  &  n1951  &  n1944 ) ;
 assign n1953 = ( (~ n616) ) | ( n1269 ) ;
 assign n1954 = ( (~ n616) ) | ( n2611 ) ;
 assign n1955 = ( (~ n616) ) | ( n1394 ) ;
 assign n1952 = ( n1953  &  n1140  &  n1954  &  n1955 ) ;
 assign n1956 = ( n464  &  n568 ) ;
 assign n1957 = ( n576  &  n788 ) ;
 assign n1958 = ( n316  &  n347 ) ;
 assign n1960 = ( (~ n21) ) | ( n1518 ) ;
 assign n1962 = ( (~ n17) ) | ( n1518 ) ;
 assign n1964 = ( (~ n21) ) | ( n837 ) ;
 assign n1965 = ( n2097  &  n2123  &  n2406  &  n2215 ) ;
 assign n1959 = ( (~ n18)  &  (~ n28)  &  n1960  &  n1962  &  n1964  &  n1965 ) ;
 assign n1967 = ( n1451  &  n848  &  n925  &  n1623  &  n2049  &  n1144 ) ;
 assign n1966 = ( n1065  &  n1125  &  n1917  &  n1949  &  n1952  &  n1967 ) ;
 assign n1969 = ( (~ n17) ) | ( n507 ) ;
 assign n1970 = ( (~ n17) ) | ( n193 ) ;
 assign n1971 = ( (~ n21) ) | ( n1122 ) ;
 assign n1968 = ( n1969  &  n1970  &  n1971 ) ;
 assign n1975 = ( (~ n34) ) | ( n536 ) ;
 assign n1976 = ( (~ n34) ) | ( n537 ) ;
 assign n1977 = ( (~ n300)  &  n1486 ) | ( n854  &  n1123  &  n1486 ) ;
 assign n1972 = ( n538  &  (~ n1168)  &  (~ n1169)  &  n1975  &  n1976  &  n1977 ) ;
 assign n1978 = ( (~ n34) ) | ( n1122 ) ;
 assign n1979 = ( (~ n34) ) | ( n739 ) ;
 assign n1980 = ( (~ n34) ) | ( n1394 ) ;
 assign n1981 = ( (~ n616) ) | ( n1121 ) ;
 assign n1983 = ( (~ n34) ) | ( n1121 ) ;
 assign n1984 = ( (~ n34) ) | ( n2607 ) ;
 assign n1986 = ( (~ n17) ) | ( n766 ) ;
 assign n1987 = ( (~ n17) ) | ( n466 ) ;
 assign n1989 = ( (~ n17) ) | ( n536 ) ;
 assign n1991 = ( (~ n17) ) | ( n709 ) ;
 assign n1985 = ( (~ n14)  &  (~ n1165)  &  n1986  &  n1987  &  n1989  &  n1991 ) ;
 assign n1992 = ( (~ n17) ) | ( n1122 ) ;
 assign n1994 = ( (~ n21) ) | ( n565 ) ;
 assign n1995 = ( (~ n21) ) | ( n1394 ) ;
 assign n1996 = ( (~ n21) ) | ( n641 ) ;
 assign n1998 = ( (~ n17) ) | ( n291 ) ;
 assign n1999 = ( (~ n17) ) | ( n324 ) ;
 assign n2000 = ( (~ n17) ) | ( n505 ) ;
 assign n2001 = ( (~ n17) ) | ( n373 ) ;
 assign n2002 = ( n2266  &  n2082  &  n2306 ) ;
 assign n2003 = ( (~ n25)  &  n456  &  n2094  &  n2119  &  n2125  &  n2231  &  n2386  &  n2536 ) ;
 assign n2004 = ( (~ n616) ) | ( n2423 ) ;
 assign n2005 = ( (~ n616) ) | ( n1222 ) ;
 assign n2006 = ( (~ n34) ) | ( n1521 ) ;
 assign n2007 = ( n438  &  n252 ) ;
 assign n2009 = ( (~ n34) ) | ( n897 ) ;
 assign n2010 = ( (~ n34) ) | ( n1221 ) ;
 assign n2011 = ( n530  &  n1237 ) ;
 assign n2012 = ( n295  &  (~ n1021) ) ;
 assign n2014 = ( (~ n34) ) | ( n2606 ) ;
 assign n2015 = ( (~ n34) ) | ( n993 ) ;
 assign n2017 = ( (~ n34) ) | ( n2613 ) ;
 assign n2018 = ( (~ n34) ) | ( n1237 ) ;
 assign n2019 = ( (~ n34) ) | ( n530 ) ;
 assign n2020 = ( (~ n17) ) | ( n381 ) ;
 assign n2021 = ( (~ n21) ) | ( n1237 ) ;
 assign n2022 = ( (~ n17) ) | ( n530 ) ;
 assign n2023 = ( (~ n17) ) | ( n1329 ) ;
 assign n2024 = ( (~ n17) ) | ( n508 ) ;
 assign n2025 = ( (~ n17) ) | ( n1237 ) ;
 assign n2026 = ( (~ n17) ) | ( n768 ) ;
 assign n2028 = ( (~ n34) ) | ( n2612 ) ;
 assign n2027 = ( n1177  &  n1179  &  n2028 ) ;
 assign n2030 = ( (~ n247) ) | ( n1520 ) ;
 assign n2031 = ( (~ n247) ) | ( n1352 ) ;
 assign n2032 = ( (~ n247) ) | ( n864 ) ;
 assign n2029 = ( n2030  &  n2031  &  n2032 ) ;
 assign n2034 = ( (~ n10) ) | ( n341 ) ;
 assign n2035 = ( n1114  &  n2029  &  n1837  &  n1116 ) ;
 assign n2033 = ( n2034  &  n1975  &  n1976  &  n1306  &  n1825  &  n2035 ) ;
 assign n2036 = ( (~ n616) ) | ( n1251 ) ;
 assign n2037 = ( (~ n34) ) | ( n1250 ) ;
 assign n2038 = ( n2353  &  n2341  &  n2308  &  n2376  &  n2284  &  n2574 ) ;
 assign n2039 = ( n800  &  n810 ) ;
 assign n2040 = ( n739  &  n313 ) ;
 assign n2041 = ( n263  &  n530 ) ;
 assign n2042 = ( n465  &  n711 ) ;
 assign n2043 = ( n288  &  n198 ) ;
 assign n2044 = ( (~ n6) ) | ( n508 ) ;
 assign n2045 = ( (~ n135) ) | ( n1394 ) ;
 assign n2046 = ( (~ n135) ) | ( n373 ) ;
 assign n2047 = ( (~ n135) ) | ( n193 ) ;
 assign n2048 = ( (~ n135) ) | ( n214 ) ;
 assign n2049 = ( (~ n426) ) | ( n1394 ) ;
 assign n2050 = ( (~ n135) ) | ( n1329 ) ;
 assign n2051 = ( n213 ) | ( (~ n426) ) ;
 assign n2052 = ( n214 ) | ( (~ n426) ) ;
 assign n2053 = ( n193 ) | ( (~ n426) ) ;
 assign n2054 = ( n243 ) | ( (~ n426) ) ;
 assign n2055 = ( (~ n426) ) | ( n508 ) ;
 assign n2056 = ( (~ n426) ) | ( n1271 ) ;
 assign n2057 = ( (~ n426) ) | ( n1329 ) ;
 assign n2058 = ( n373 ) | ( (~ n426) ) ;
 assign n2059 = ( (~ n426) ) | ( n1377 ) ;
 assign n2060 = ( (~ n21) ) | ( n468 ) ;
 assign n2061 = ( (~ n139) ) | ( n193 ) ;
 assign n2064 = ( (~ n17) ) | ( n213 ) ;
 assign n2065 = ( n342 ) | ( (~ n616) ) ;
 assign n2067 = ( (~ n131) ) | ( n1012 ) ;
 assign n2066 = ( n1694  &  n2067  &  n1685  &  n1663  &  n1305  &  n1705 ) ;
 assign n2068 = ( (~ n6) ) | ( n959 ) ;
 assign n2070 = ( (~ n135) ) | ( n953 ) ;
 assign n2071 = ( (~ n135) ) | ( n288 ) ;
 assign n2069 = ( n1826  &  n1862  &  n2070  &  n1679  &  n1656  &  n2071 ) ;
 assign n2072 = ( (~ n131) ) | ( n726 ) ;
 assign n2073 = ( (~ n131) ) | ( n959 ) ;
 assign n2075 = ( (~ n426) ) | ( n1071 ) ;
 assign n2076 = ( (~ n426) ) | ( n544 ) ;
 assign n2077 = ( n288 ) | ( (~ n426) ) ;
 assign n2078 = ( (~ n426) ) | ( n726 ) ;
 assign n2079 = ( n316 ) | ( (~ n426) ) ;
 assign n2074 = ( n2075  &  n2076  &  n1935  &  n2077  &  n2078  &  n2079 ) ;
 assign n2080 = ( (~ n139) ) | ( n1431 ) ;
 assign n2081 = ( (~ n426) ) | ( n1395 ) ;
 assign n2082 = ( (~ n17) ) | ( n726 ) ;
 assign n2083 = ( (~ n131)  &  (~ n139) ) | ( (~ n139)  &  n176 ) | ( (~ n131)  &  n565 ) | ( n176  &  n565 ) ;
 assign n2084 = ( n1093  &  n336 ) | ( n1093  &  n1433  &  n1432 ) ;
 assign n2085 = ( n294 ) | ( n953 ) ;
 assign n2088 = ( (~ n10) ) | ( n176 ) ;
 assign n2089 = ( (~ n10) ) | ( n565 ) ;
 assign n2090 = ( (~ n280) ) | ( n1012 ) ;
 assign n2091 = ( n176 ) | ( (~ n280) ) ;
 assign n2092 = ( (~ n10) ) | ( n1071 ) ;
 assign n2093 = ( (~ n21) ) | ( n1215 ) ;
 assign n2094 = ( (~ n21) ) | ( n291 ) ;
 assign n2095 = ( (~ n139) ) | ( n1012 ) ;
 assign n2096 = ( (~ n139) ) | ( n288 ) ;
 assign n2097 = ( (~ n21) ) | ( n316 ) ;
 assign n2098 = ( (~ n21) ) | ( n1012 ) ;
 assign n2099 = ( (~ n21) ) | ( n288 ) ;
 assign n2100 = ( n1805  &  n296 ) | ( n994  &  n296 ) | ( n1805  &  n259 ) | ( n994  &  n259 ) ;
 assign n2101 = ( n295  &  (~ n479) ) ;
 assign n2103 = ( n336  &  (~ n426) ) ;
 assign n2102 = ( n263  &  n313 ) | ( n313  &  (~ n358) ) | ( n263  &  n2103 ) | ( (~ n358)  &  n2103 ) ;
 assign n2105 = ( n175 ) | ( (~ n280) ) ;
 assign n2106 = ( (~ n247) ) | ( n323 ) ;
 assign n2108 = ( (~ n280) ) | ( n324 ) ;
 assign n2107 = ( n1790  &  n1741  &  n2108 ) ;
 assign n2109 = ( n193 ) | ( (~ n280) ) ;
 assign n2110 = ( (~ n280) ) | ( n1271 ) ;
 assign n2112 = ( (~ n139) ) | ( n243 ) ;
 assign n2113 = ( (~ n139) ) | ( n897 ) ;
 assign n2114 = ( (~ n139) ) | ( n204 ) ;
 assign n2115 = ( (~ n280) ) | ( n323 ) ;
 assign n2116 = ( n204 ) | ( (~ n280) ) ;
 assign n2111 = ( n2112  &  n2113  &  n2114  &  n2115  &  n2116  &  n1091 ) ;
 assign n2118 = ( (~ n139) ) | ( n1329 ) ;
 assign n2119 = ( (~ n21) ) | ( n324 ) ;
 assign n2117 = ( n1931  &  n1929  &  n2118  &  n2119  &  n1108  &  n2111 ) ;
 assign n2121 = ( (~ n34) ) | ( n323 ) ;
 assign n2120 = ( n323  &  n1200  &  n2121 ) | ( (~ n370)  &  n1200  &  n2121 ) ;
 assign n2122 = ( (~ n21)  &  n1405 ) | ( n193  &  n1405 ) ;
 assign n2123 = ( (~ n21) ) | ( n1271 ) ;
 assign n2124 = ( (~ n21) ) | ( n897 ) ;
 assign n2125 = ( (~ n21) ) | ( n373 ) ;
 assign n2126 = ( (~ n21) ) | ( n204 ) ;
 assign n2127 = ( (~ n280) ) | ( n1394 ) ;
 assign n2128 = ( n213 ) | ( (~ n280) ) ;
 assign n2129 = ( (~ n10) ) | ( n213 ) ;
 assign n2130 = ( n214 ) | ( (~ n280) ) ;
 assign n2131 = ( (~ n247) ) | ( n897 ) ;
 assign n2132 = ( (~ n10) ) | ( n1394 ) ;
 assign n2133 = ( (~ n247) ) | ( n214 ) ;
 assign n2134 = ( (~ n139) ) | ( n1394 ) ;
 assign n2135 = ( (~ n34) ) | ( n1271 ) ;
 assign n2136 = ( (~ n34) ) | ( n2043 ) ;
 assign n2139 = ( (~ n10) ) | ( n837 ) ;
 assign n2138 = ( n2139  &  n1302 ) ;
 assign n2141 = ( (~ n247) ) | ( n2607 ) ;
 assign n2140 = ( n1610  &  n934  &  n1617  &  n542  &  n1645  &  n911  &  n2141  &  n2138 ) ;
 assign n2143 = ( (~ n280) ) | ( n342 ) ;
 assign n2142 = ( n1883  &  n1887  &  n2143 ) ;
 assign n2144 = ( (~ n139) ) | ( n815 ) ;
 assign n2145 = ( (~ n139) ) | ( n1379 ) ;
 assign n2146 = ( (~ n139) ) | ( n837 ) ;
 assign n2148 = ( (~ n10)  &  (~ n139)  &  (~ n248)  &  (~ n370) ) ;
 assign n2150 = ( (~ n135) ) | ( n345 ) ;
 assign n2151 = ( n342 ) | ( (~ n426) ) ;
 assign n2149 = ( n2150  &  n2151  &  n1648  &  n1668  &  n908  &  n803  &  n951  &  n1533 ) ;
 assign n2152 = ( n348 ) | ( n351 ) | ( n355 ) | ( n356 ) | ( (~ n1149) ) | ( (~ n2005) ) | ( (~ n2028) ) | ( (~ n2149) ) ;
 assign n2157 = ( n295  &  (~ n371) ) | ( n346  &  (~ n371) ) | ( n295  &  n2039 ) | ( n346  &  n2039 ) ;
 assign n2159 = ( n339  &  (~ n479) ) | ( (~ n479)  &  n1428 ) | ( n339  &  n1890 ) | ( n1428  &  n1890 ) ;
 assign n2161 = ( (~ n39)  &  (~ n375)  &  n2159 ) | ( n315  &  (~ n375)  &  n2159 ) ;
 assign n2163 = ( (~ n21)  &  n314 ) | ( n310  &  n314 ) | ( (~ n21)  &  (~ n616) ) | ( n310  &  (~ n616) ) ;
 assign n2164 = ( (~ n363)  &  n2161  &  n2163 ) | ( n1449  &  n2161  &  n2163 ) ;
 assign n2168 = ( n1427  &  n2103 ) | ( n726  &  n2103 ) | ( n1427  &  n652 ) | ( n726  &  n652 ) ;
 assign n2169 = ( n293  &  (~ n367) ) | ( n336  &  (~ n367) ) | ( n293  &  n659 ) | ( n336  &  n659 ) ;
 assign n2171 = ( (~ n34)  &  (~ n360) ) | ( (~ n34)  &  n742 ) | ( (~ n360)  &  n1222 ) | ( n742  &  n1222 ) ;
 assign n2172 = ( (~ n266)  &  n2171 ) | ( (~ n426)  &  n2171 ) ;
 assign n2173 = ( (~ n248)  &  n341 ) | ( n341  &  n576 ) | ( (~ n248)  &  (~ n1021) ) | ( n576  &  (~ n1021) ) ;
 assign n2174 = ( (~ n131)  &  (~ n139) ) | ( (~ n139)  &  n175 ) | ( (~ n131)  &  n176 ) | ( n175  &  n176 ) ;
 assign n2175 = ( n335  &  n343  &  n321  &  n2174  &  n2173  &  n2169  &  n2168  &  n2172 ) ;
 assign n2176 = ( n1467  &  n186  &  n194  &  n192  &  n183  &  n179  &  n174 ) ;
 assign n2177 = ( n596  &  n268  &  n1451  &  n303  &  n250  &  n1463  &  n197  &  n2176 ) ;
 assign n2178 = ( n345  &  n1349 ) ;
 assign n2179 = ( (~ n39)  &  n516 ) | ( (~ n39)  &  n1137 ) | ( n516  &  n1322 ) | ( n1137  &  n1322 ) ;
 assign n2180 = ( (~ n982)  &  n1137 ) | ( (~ n982)  &  n1328 ) | ( n1137  &  n1349 ) | ( n1328  &  n1349 ) ;
 assign n2182 = ( n1596 ) | ( n491 ) ;
 assign n2184 = ( (~ n10) ) | ( n453 ) ;
 assign n2185 = ( (~ n247) ) | ( n453 ) ;
 assign n2183 = ( n1738  &  n1739  &  n1734  &  n1735  &  n2184  &  n1699  &  n1713  &  n2185 ) ;
 assign n2186 = ( (~ n280) ) | ( n1473 ) ;
 assign n2187 = ( (~ n280) ) | ( n506 ) ;
 assign n2188 = ( (~ n280) ) | ( n1478 ) ;
 assign n2189 = ( (~ n139) ) | ( n465 ) ;
 assign n2190 = ( (~ n280) ) | ( n1480 ) ;
 assign n2191 = ( (~ n280) ) | ( n453 ) ;
 assign n2192 = ( (~ n139) ) | ( n1480 ) ;
 assign n2193 = ( (~ n139) ) | ( n453 ) ;
 assign n2194 = ( (~ n139) ) | ( n1191 ) ;
 assign n2195 = ( n695  &  n319  &  n642 ) ;
 assign n2197 = ( (~ n6) ) | ( (~ n476) ) ;
 assign n2196 = ( n714  &  n1571  &  n2197  &  n178  &  n666  &  n1715  &  n181  &  n2195 ) ;
 assign n2198 = ( n1614  &  n1637  &  n1611  &  n804 ) ;
 assign n2199 = ( n1303  &  n855  &  n654  &  n657 ) ;
 assign n2200 = ( n1621  &  n647  &  n650  &  n1470  &  n1569  &  n2199 ) ;
 assign n2201 = ( n849  &  n842  &  n1647 ) ;
 assign n2203 = ( (~ n135) ) | ( n1352 ) ;
 assign n2204 = ( (~ n6) ) | ( n1490 ) ;
 assign n2205 = ( (~ n247) ) | ( n2610 ) ;
 assign n2202 = ( n1856  &  n2203  &  n2204  &  n2205  &  n673  &  n1667  &  n2201  &  n2200 ) ;
 assign n2207 = ( (~ n135) ) | ( n464 ) ;
 assign n2208 = ( (~ n426) ) | ( n1269 ) ;
 assign n2206 = ( n2207  &  n2208  &  n578 ) ;
 assign n2209 = ( (~ n43)  &  n1428 ) | ( (~ n43)  &  n524  &  n1269 ) ;
 assign n2210 = ( (~ n474)  &  (~ n477)  &  (~ n478)  &  (~ n481)  &  n700  &  n1422  &  n1896  &  n2209 ) ;
 assign n2215 = ( (~ n17) ) | ( n464 ) ;
 assign n2216 = ( (~ n426) ) | ( n464 ) ;
 assign n2217 = ( n464  &  n1484 ) | ( (~ n683)  &  n1484 ) | ( n464  &  n2103 ) | ( (~ n683)  &  n2103 ) ;
 assign n2218 = ( (~ n364)  &  (~ n401) ) | ( (~ n364)  &  n1250 ) | ( (~ n401)  &  n1377 ) | ( n1250  &  n1377 ) ;
 assign n2221 = ( (~ n300)  &  n580 ) | ( n463  &  n580 ) | ( (~ n300)  &  n1206 ) | ( n463  &  n1206 ) ;
 assign n2224 = ( (~ n10) ) | ( n1492 ) ;
 assign n2225 = ( (~ n360)  &  (~ n363) ) | ( (~ n360)  &  n468 ) | ( (~ n363)  &  n1264 ) | ( n468  &  n1264 ) ;
 assign n2226 = ( (~ n6)  &  n2225 ) | ( n1329  &  n2225 ) ;
 assign n2228 = ( (~ n247) ) | ( n1250 ) ;
 assign n2227 = ( n1644  &  n1616  &  n1609  &  n1600  &  n1574  &  n2228  &  n718  &  n1573 ) ;
 assign n2229 = ( (~ n280) ) | ( n1269 ) ;
 assign n2230 = ( (~ n34) ) | ( n1206 ) ;
 assign n2231 = ( (~ n21) ) | ( n1206 ) ;
 assign n2232 = ( (~ n139) ) | ( n1484 ) ;
 assign n2233 = ( (~ n139) ) | ( n1264 ) ;
 assign n2234 = ( (~ n139) ) | ( n464 ) ;
 assign n2235 = ( (~ n280) ) | ( n1258 ) ;
 assign n2236 = ( (~ n21)  &  (~ n370) ) ;
 assign n2237 = ( n1717  &  n1633  &  n1642 ) ;
 assign n2239 = ( (~ n131) ) | ( n1480 ) ;
 assign n2240 = ( (~ n131) ) | ( n453 ) ;
 assign n2238 = ( n2239  &  n2240 ) ;
 assign n2242 = ( (~ n131) ) | ( n1473 ) ;
 assign n2243 = ( (~ n131) ) | ( n1191 ) ;
 assign n2241 = ( n2242  &  n1660  &  n1704  &  n1692  &  n1697  &  n2243  &  n1683  &  n2238 ) ;
 assign n2244 = ( (~ n6) ) | ( n768 ) ;
 assign n2245 = ( (~ n6) ) | ( n1478 ) ;
 assign n2247 = ( (~ n131) ) | ( n768 ) ;
 assign n2248 = ( (~ n131) ) | ( n1478 ) ;
 assign n2246 = ( n1653  &  n1678  &  n2247  &  n2248 ) ;
 assign n2249 = ( n1731  &  n1747  &  n1730  &  n1721  &  n1786  &  n2246 ) ;
 assign n2251 = ( (~ n135) ) | ( n507 ) ;
 assign n2250 = ( n2251  &  n1827  &  n1860 ) ;
 assign n2252 = ( (~ n135) ) | ( n768 ) ;
 assign n2253 = ( (~ n135) ) | ( n505 ) ;
 assign n2254 = ( (~ n135) ) | ( n465 ) ;
 assign n2256 = ( (~ n426) ) | ( n505 ) ;
 assign n2257 = ( (~ n426) ) | ( n1191 ) ;
 assign n2255 = ( n2256  &  n2257 ) ;
 assign n2259 = ( (~ n139) ) | ( n1479 ) ;
 assign n2260 = ( (~ n426) ) | ( n465 ) ;
 assign n2261 = ( (~ n426) ) | ( n1473 ) ;
 assign n2258 = ( n1831  &  n1838  &  n1900  &  n1117  &  n2259  &  n2260  &  n2261  &  n2255 ) ;
 assign n2263 = ( (~ n426) ) | ( n1478 ) ;
 assign n2264 = ( (~ n426) ) | ( n1477 ) ;
 assign n2265 = ( n412 ) | ( (~ n426) ) ;
 assign n2262 = ( n2263  &  n2264  &  n2265 ) ;
 assign n2266 = ( (~ n17) ) | ( n1191 ) ;
 assign n2268 = ( (~ n17) ) | ( n506 ) ;
 assign n2269 = ( (~ n21) ) | ( n413 ) ;
 assign n2267 = ( n2268  &  n1904  &  n2026  &  n2269 ) ;
 assign n2270 = ( (~ n139) ) | ( n507 ) ;
 assign n2271 = ( (~ n21)  &  (~ n426) ) | ( n412  &  (~ n426) ) | ( (~ n21)  &  n507 ) | ( n412  &  n507 ) ;
 assign n2274 = ( (~ n10)  &  (~ n426) ) ;
 assign n2272 = ( (~ n301)  &  n1480 ) | ( n1191  &  n1480 ) | ( (~ n301)  &  n2274 ) | ( n1191  &  n2274 ) ;
 assign n2275 = ( (~ n400)  &  (~ n401) ) | ( (~ n400)  &  n465 ) | ( (~ n401)  &  n506 ) | ( n465  &  n506 ) ;
 assign n2276 = ( (~ n280) ) | ( n530 ) ;
 assign n2277 = ( (~ n280) ) | ( n739 ) ;
 assign n2278 = ( (~ n370) ) | ( n380 ) ;
 assign n2279 = ( (~ n139) ) | ( n739 ) ;
 assign n2280 = ( (~ n280) ) | ( n1476 ) ;
 assign n2281 = ( (~ n280) ) | ( n380 ) ;
 assign n2282 = ( (~ n280) ) | ( n611 ) ;
 assign n2284 = ( (~ n34) ) | ( n611 ) ;
 assign n2285 = ( (~ n34) ) | ( n524 ) ;
 assign n2286 = ( (~ n139) ) | ( n1476 ) ;
 assign n2283 = ( n2284  &  n1927  &  n1920  &  n2285  &  n1979  &  n1812  &  n1815  &  n2286 ) ;
 assign n2287 = ( (~ n21)  &  (~ n280) ) | ( (~ n280)  &  n379 ) | ( (~ n21)  &  n1250 ) | ( n379  &  n1250 ) ;
 assign n2288 = ( (~ n21) ) | ( n1476 ) ;
 assign n2290 = ( (~ n131) ) | ( n739 ) ;
 assign n2291 = ( (~ n131) ) | ( n1476 ) ;
 assign n2292 = ( (~ n131) ) | ( n740 ) ;
 assign n2289 = ( n1703  &  n2290  &  n1664  &  n784  &  n2291  &  n1695  &  n2292 ) ;
 assign n2293 = ( (~ n131) ) | ( n530 ) ;
 assign n2294 = ( (~ n131) ) | ( n448 ) ;
 assign n2295 = ( (~ n131) ) | ( n381 ) ;
 assign n2297 = ( (~ n426) ) | ( n448 ) ;
 assign n2298 = ( (~ n139) ) | ( n709 ) ;
 assign n2296 = ( n2297  &  n2298  &  n1936  &  n1894  &  n1881  &  n1902 ) ;
 assign n2299 = ( (~ n135) ) | ( n470 ) ;
 assign n2300 = ( (~ n135) ) | ( n537 ) ;
 assign n2301 = ( (~ n135) ) | ( n381 ) ;
 assign n2302 = ( (~ n135) ) | ( n921 ) ;
 assign n2304 = ( (~ n21) ) | ( n1474 ) ;
 assign n2303 = ( n2020  &  n2022  &  n1217  &  n1941  &  n1905  &  n2304 ) ;
 assign n2305 = ( n994 ) | ( n524 ) ;
 assign n2306 = ( (~ n17) ) | ( n448 ) ;
 assign n2307 = ( (~ n139) ) | ( n470 ) ;
 assign n2308 = ( (~ n616) ) | ( n1250 ) ;
 assign n2309 = ( (~ n125)  &  (~ n1021) ) | ( (~ n125)  &  n709  &  n740 ) ;
 assign n2310 = ( n334  &  (~ n360) ) | ( (~ n360)  &  n530 ) | ( n334  &  n739 ) | ( n530  &  n739 ) ;
 assign n2311 = ( (~ n399)  &  n470 ) | ( (~ n34)  &  (~ n280)  &  (~ n399) ) ;
 assign n2313 = ( (~ n426)  &  n1476 ) | ( n1476  &  n1554 ) | ( (~ n426)  &  n2274 ) | ( n1554  &  n2274 ) ;
 assign n2314 = ( (~ n300)  &  n521  &  n1099 ) | ( n500  &  n521  &  n1099 ) ;
 assign n2315 = ( n336  &  (~ n509) ) | ( n453  &  (~ n509)  &  n788 ) ;
 assign n2317 = ( n295  &  (~ n364) ) | ( n295  &  n567 ) | ( (~ n364)  &  n1550 ) | ( n567  &  n1550 ) ;
 assign n2318 = ( n1427 ) | ( n1191 ) ;
 assign n2319 = ( (~ n10)  &  (~ n378) ) | ( (~ n10)  &  n524 ) | ( (~ n378)  &  n530 ) | ( n524  &  n530 ) ;
 assign n2320 = ( n2319  &  n516 ) | ( n2319  &  n491 ) ;
 assign n2321 = ( n213 ) | ( (~ n978) ) ;
 assign n2323 = ( (~ n6) ) | ( n737 ) ;
 assign n2324 = ( (~ n6) ) | ( n1237 ) ;
 assign n2322 = ( n833  &  n1641  &  n1716  &  n1632  &  n2323  &  n2324  &  n794 ) ;
 assign n2325 = ( (~ n131) ) | ( n541 ) ;
 assign n2326 = ( (~ n131) ) | ( n1122 ) ;
 assign n2327 = ( (~ n131) ) | ( n641 ) ;
 assign n2329 = ( (~ n131) ) | ( n737 ) ;
 assign n2330 = ( (~ n131) ) | ( n1237 ) ;
 assign n2331 = ( (~ n131) ) | ( n706 ) ;
 assign n2328 = ( n1677  &  n2329  &  n2330  &  n2331  &  n1854  &  n1638  &  n1049 ) ;
 assign n2332 = ( (~ n135) ) | ( n641 ) ;
 assign n2334 = ( (~ n426) ) | ( n612 ) ;
 assign n2335 = ( (~ n426) ) | ( n1518 ) ;
 assign n2336 = ( (~ n426) ) | ( n536 ) ;
 assign n2337 = ( n994 ) | ( n1518 ) ;
 assign n2333 = ( n2334  &  n2335  &  n2336  &  n1899  &  n1962  &  n1989  &  n2337 ) ;
 assign n2338 = ( n994 ) | ( n566 ) ;
 assign n2339 = ( (~ n17) ) | ( n612 ) ;
 assign n2340 = ( (~ n17) ) | ( n1077 ) ;
 assign n2341 = ( (~ n616) ) | ( n1077 ) ;
 assign n2343 = ( (~ n400)  &  n993 ) | ( n737  &  n993 ) | ( (~ n400)  &  n2012 ) | ( n737  &  n2012 ) ;
 assign n2347 = ( (~ n280) ) | ( n1121 ) ;
 assign n2344 = ( (~ n7)  &  (~ n25)  &  n2347 ) ;
 assign n2348 = ( (~ n34) ) | ( n1193 ) ;
 assign n2349 = ( (~ n280) ) | ( n2613 ) ;
 assign n2350 = ( (~ n21) ) | ( n2608 ) ;
 assign n2351 = ( (~ n34) ) | ( n1957 ) ;
 assign n2353 = ( (~ n34) ) | ( n1251 ) ;
 assign n2352 = ( (~ n139)  &  n1100  &  n2353 ) | ( n381  &  n1100  &  n2353 ) ;
 assign n2355 = ( (~ n247) ) | ( n1237 ) ;
 assign n2356 = ( (~ n10) ) | ( n536 ) ;
 assign n2357 = ( (~ n247) ) | ( n1290 ) ;
 assign n2354 = ( n2355  &  n2356  &  n1707  &  n2357  &  n1712  &  n1646 ) ;
 assign n2359 = ( (~ n10) ) | ( n1077 ) ;
 assign n2360 = ( (~ n280) ) | ( n1122 ) ;
 assign n2361 = ( (~ n10) ) | ( n1519 ) ;
 assign n2358 = ( n2359  &  n1858  &  n2360  &  n2361  &  n1746  &  n1791  &  n2354 ) ;
 assign n2363 = ( (~ n280) ) | ( n612 ) ;
 assign n2364 = ( (~ n280) ) | ( n1237 ) ;
 assign n2365 = ( (~ n280) ) | ( n1519 ) ;
 assign n2362 = ( n2363  &  n1037  &  n1878  &  n1884  &  n2364  &  n2365 ) ;
 assign n2366 = ( (~ n139) ) | ( n1122 ) ;
 assign n2367 = ( (~ n370) ) | ( n1519 ) ;
 assign n2368 = ( (~ n370) ) | ( n1290 ) ;
 assign n2369 = ( (~ n280) ) | ( n1290 ) ;
 assign n2370 = ( (~ n139) ) | ( n1518 ) ;
 assign n2371 = ( (~ n139) ) | ( n1237 ) ;
 assign n2372 = ( (~ n21) ) | ( n612 ) ;
 assign n2373 = ( (~ n34) ) | ( n1518 ) ;
 assign n2374 = ( (~ n21) ) | ( n1077 ) ;
 assign n2375 = ( (~ n21) ) | ( n1519 ) ;
 assign n2376 = ( (~ n34) ) | ( n612 ) ;
 assign n2378 = ( n719  &  n1572  &  n720 ) ;
 assign n2379 = ( n1674  &  n1650  &  n846 ) ;
 assign n2380 = ( n1326 ) | ( (~ n1534) ) ;
 assign n2381 = ( (~ n280) ) | ( n1043 ) ;
 assign n2383 = ( (~ n139) ) | ( n568 ) ;
 assign n2384 = ( (~ n280) ) | ( n559 ) ;
 assign n2385 = ( (~ n139) ) | ( n560 ) ;
 assign n2382 = ( n2383  &  n2384  &  n2385 ) ;
 assign n2386 = ( (~ n21) ) | ( n581 ) ;
 assign n2387 = ( (~ n34) ) | ( n581 ) ;
 assign n2388 = ( (~ n139) ) | ( n1521 ) ;
 assign n2389 = ( (~ n1016) ) | ( n1821 ) ;
 assign n2390 = ( (~ n280)  &  n727 ) | ( n706  &  n727 ) | ( (~ n280)  &  n1012 ) | ( n706  &  n1012 ) ;
 assign n2392 = ( n959  &  n541  &  n573 ) ;
 assign n2394 = ( n1319 ) | ( (~ n1525) ) ;
 assign n2395 = ( n670  &  n182 ) ;
 assign n2396 = ( n191  &  n715  &  n1570  &  n202  &  n667  &  n320  &  n696  &  n2395 ) ;
 assign n2397 = ( n1613  &  n802  &  n1690  &  n2030 ) ;
 assign n2398 = ( n1620  &  n1640  &  n1771 ) ;
 assign n2399 = ( n1423  &  n1810  &  n672  &  n918  &  n840  &  n850  &  n856  &  n1304 ) ;
 assign n2400 = ( n656  &  n653  &  n675  &  n1469  &  n649  &  n646  &  n2398  &  n2399 ) ;
 assign n2401 = ( (~ n6) ) | ( n560 ) ;
 assign n2403 = ( (~ n135) ) | ( n568 ) ;
 assign n2404 = ( (~ n135) ) | ( n1520 ) ;
 assign n2402 = ( n2403  &  n2404  &  n1898 ) ;
 assign n2406 = ( (~ n17) ) | ( n568 ) ;
 assign n2405 = ( (~ n37)  &  n660  &  n1466  &  n2406 ) ;
 assign n2407 = ( (~ n371)  &  n1918 ) | ( n176  &  n1519  &  n1918 ) ;
 assign n2408 = ( (~ n479)  &  (~ n583) ) | ( n564  &  (~ n583)  &  n1520 ) ;
 assign n2410 = ( (~ n247)  &  n734 ) | ( n558  &  n734 ) | ( (~ n247)  &  n993 ) | ( n558  &  n993 ) ;
 assign n2411 = ( (~ n300)  &  n336 ) | ( (~ n300)  &  n555 ) | ( n336  &  n562 ) | ( n555  &  n562 ) ;
 assign n2412 = ( (~ n426) ) | ( n568 ) ;
 assign n2413 = ( (~ n135)  &  (~ n354) ) | ( (~ n354)  &  n563 ) | ( (~ n135)  &  n1043 ) | ( n563  &  n1043 ) ;
 assign n2415 = ( n316  &  (~ n378) ) | ( (~ n363)  &  (~ n378) ) | ( n316  &  n566 ) | ( (~ n363)  &  n566 ) ;
 assign n2416 = ( (~ n1021)  &  n2036 ) | ( n1431  &  n1524  &  n2036 ) ;
 assign n2417 = ( (~ n378)  &  n2416 ) | ( n559  &  n1290  &  n2416 ) ;
 assign n2418 = ( (~ n627)  &  n1428 ) | ( (~ n627)  &  n1432  &  n1550 ) ;
 assign n2420 = ( (~ n616)  &  (~ n630) ) | ( n576  &  (~ n630)  &  n1193 ) ;
 assign n2422 = ( (~ n17)  &  n289 ) | ( (~ n17)  &  n953 ) | ( n289  &  n1433 ) | ( n953  &  n1433 ) ;
 assign n2423 = ( n544  &  n501 ) ;
 assign n2424 = ( n243  &  n292 ) | ( n292  &  (~ n354) ) | ( n243  &  (~ n360) ) | ( (~ n354)  &  (~ n360) ) ;
 assign n2425 = ( (~ n247)  &  (~ n135) ) | ( (~ n135)  &  n204 ) | ( (~ n247)  &  n544 ) | ( n204  &  n544 ) ;
 assign n2426 = ( n391  &  n337  &  n2425  &  n304 ) ;
 assign n2427 = ( n527  &  n529  &  n522 ) ;
 assign n2429 = ( n1688  &  n1598 ) ;
 assign n2431 = ( (~ n10) ) | ( n1120 ) ;
 assign n2432 = ( (~ n139) ) | ( n839 ) ;
 assign n2433 = ( (~ n139) ) | ( n854 ) ;
 assign n2434 = ( (~ n139) ) | ( n707 ) ;
 assign n2435 = ( (~ n280) ) | ( n704 ) ;
 assign n2436 = ( (~ n21)  &  n1564 ) | ( n680  &  n1564 ) | ( (~ n21)  &  n2148 ) | ( n680  &  n2148 ) ;
 assign n2438 = ( (~ n21) ) | ( n2609 ) ;
 assign n2439 = ( (~ n21) ) | ( n704 ) ;
 assign n2441 = ( (~ n21) ) | ( n1824 ) ;
 assign n2437 = ( (~ n22)  &  (~ n682)  &  n1178  &  n1921  &  n2436  &  n2438  &  n2439  &  n2441 ) ;
 assign n2442 = ( (~ n248)  &  n1392 ) | ( n854  &  n1392 ) | ( (~ n248)  &  (~ n1534) ) | ( n854  &  (~ n1534) ) ;
 assign n2443 = ( (~ n426)  &  n528 ) | ( n528  &  n737  &  n1553 ) ;
 assign n2445 = ( (~ n131) ) | ( n677 ) ;
 assign n2444 = ( (~ n3)  &  n916  &  n948  &  n1415  &  n1468  &  n1531  &  n1857  &  n2445 ) ;
 assign n2448 = ( (~ n17) ) | ( n1563 ) ;
 assign n2449 = ( (~ n17) ) | ( n677 ) ;
 assign n2447 = ( (~ n14)  &  n1230  &  n1421  &  n1425  &  n1465  &  n1919  &  n2448  &  n2449 ) ;
 assign n2450 = ( (~ n332)  &  (~ n358) ) | ( (~ n358)  &  n738 ) | ( (~ n332)  &  n741 ) | ( n738  &  n741 ) ;
 assign n2451 = ( (~ n426)  &  (~ n744) ) | ( n742  &  (~ n744)  &  n854 ) ;
 assign n2453 = ( (~ n131)  &  (~ n747) ) | ( n704  &  (~ n747)  &  n1450 ) ;
 assign n2455 = ( n645  &  (~ n748) ) | ( (~ n139)  &  (~ n748)  &  (~ n1021) ) ;
 assign n2457 = ( n502  &  (~ n750)  &  n2455 ) | ( (~ n750)  &  n1448  &  n2455 ) ;
 assign n2460 = ( (~ n358)  &  (~ n370) ) ;
 assign n2459 = ( n311  &  n1476 ) | ( (~ n360)  &  n1476 ) | ( n311  &  n2460 ) | ( (~ n360)  &  n2460 ) ;
 assign n2461 = ( (~ n371)  &  n2457  &  n2459 ) | ( n1576  &  n2457  &  n2459 ) ;
 assign n2462 = ( (~ n140)  &  n2032  &  n2444  &  n2447  &  n2450  &  n2451  &  n2453  &  n2461 ) ;
 assign n2463 = ( (~ n350)  &  n733 ) | ( (~ n350)  &  n839 ) | ( n733  &  n1564 ) | ( n839  &  n1564 ) ;
 assign n2465 = ( (~ n300)  &  (~ n363) ) | ( (~ n363)  &  n708 ) | ( (~ n300)  &  n712 ) | ( n708  &  n712 ) ;
 assign n2466 = ( (~ n266)  &  n336 ) | ( n336  &  (~ n400) ) | ( (~ n266)  &  n703 ) | ( (~ n400)  &  n703 ) ;
 assign n2467 = ( (~ n248)  &  (~ n479) ) | ( n341  &  (~ n479) ) | ( (~ n248)  &  n864 ) | ( n341  &  n864 ) ;
 assign n2468 = ( (~ n34)  &  n295 ) | ( n295  &  n318 ) | ( (~ n34)  &  n470 ) | ( n318  &  n470 ) ;
 assign n2469 = ( (~ n247)  &  (~ n6) ) | ( (~ n6)  &  n381 ) | ( (~ n247)  &  n659 ) | ( n381  &  n659 ) ;
 assign n2470 = ( (~ n17)  &  n799 ) | ( n262  &  n799 ) | ( (~ n17)  &  n994 ) | ( n262  &  n994 ) ;
 assign n2471 = ( n232  &  n1033 ) | ( n232  &  (~ n1525) ) ;
 assign n2472 = ( n2471  &  n2470  &  n2469  &  n2468  &  n2467  &  n2466  &  n2465  &  n2463 ) ;
 assign n2473 = ( n1582  &  n685  &  n1577  &  n717  &  n595  &  n736  &  n268  &  n403 ) ;
 assign n2474 = ( n655  &  n651  &  n661  &  n1587  &  n648  &  n644  &  n643  &  n2473 ) ;
 assign n2475 = ( (~ n21)  &  (~ n139) ) | ( (~ n139)  &  n1551 ) | ( (~ n21)  &  n1552 ) | ( n1551  &  n1552 ) ;
 assign n2476 = ( (~ n426)  &  n767 ) | ( n557  &  n767 ) | ( (~ n426)  &  n1448 ) | ( n557  &  n1448 ) ;
 assign n2477 = ( n2476  &  n374 ) | ( n2476  &  n505 ) ;
 assign n2479 = ( (~ n332)  &  (~ n360) ) ;
 assign n2478 = ( n2479  &  n2460 ) | ( n993  &  n2460 ) | ( n2479  &  n1480 ) | ( n993  &  n1480 ) ;
 assign n2480 = ( (~ n300)  &  (~ n616) ) | ( (~ n616)  &  n765 ) | ( (~ n300)  &  n1195 ) | ( n765  &  n1195 ) ;
 assign n2481 = ( (~ n247)  &  (~ n332) ) | ( (~ n332)  &  n452 ) | ( (~ n247)  &  n1551 ) | ( n452  &  n1551 ) ;
 assign n2482 = ( n2481  &  n336 ) | ( n2481  &  n1491 ) ;
 assign n2483 = ( n1496  &  n1495  &  n471  &  n939  &  n2477  &  n2480  &  n2478  &  n2482 ) ;
 assign n2484 = ( (~ n358)  &  (~ n363) ) | ( (~ n358)  &  n766 ) | ( (~ n363)  &  n1477 ) | ( n766  &  n1477 ) ;
 assign n2485 = ( (~ n357)  &  n1138  &  n2484 ) | ( n559  &  n1138  &  n2484 ) ;
 assign n2486 = ( (~ n10)  &  (~ n135) ) | ( (~ n10)  &  n576 ) | ( (~ n135)  &  n1290 ) | ( n576  &  n1290 ) ;
 assign n2487 = ( n2486  &  n2485  &  n516 ) | ( n2486  &  n2485  &  n1364 ) ;
 assign n2488 = ( n661  &  n587  &  n427  &  n303  &  n756  &  n1591  &  n752  &  n2487 ) ;
 assign n2489 = ( n152  &  (~ n1362)  &  n1365 ) ;
 assign n2490 = ( n2031  &  n2030  &  n2240 ) ;
 assign n2491 = ( n226  &  n2088  &  n1406 ) ;
 assign n2492 = ( (~ n131)  &  n519  &  (~ n866) ) | ( n519  &  n863  &  (~ n866) ) ;
 assign n2494 = ( (~ n247)  &  (~ n6) ) | ( (~ n247)  &  n341 ) | ( (~ n6)  &  n822 ) | ( n341  &  n822 ) ;
 assign n2495 = ( n207  &  n903  &  n1569 ) ;
 assign n2496 = ( (~ n247)  &  n179 ) | ( n180  &  n179 ) ;
 assign n2497 = ( n450  &  n522  &  n527  &  n529  &  (~ n879)  &  (~ n882)  &  n884  &  n2496 ) ;
 assign n2500 = ( n674  &  n671 ) ;
 assign n2502 = ( (~ n1362)  &  n1366 ) ;
 assign n2501 = ( n164 ) | ( n890 ) | ( (~ n1766) ) | ( n1802 ) | ( (~ n2032) ) | ( n2502 ) ;
 assign n2504 = ( n899  &  n491 ) | ( n899  &  n516  &  n508 ) ;
 assign n2505 = ( n876  &  n875  &  n868  &  n958  &  n203  &  n607 ) ;
 assign n2506 = ( n446  &  n542  &  (~ n954)  &  (~ n955)  &  n2106  &  n2133  &  n2431  &  n2505 ) ;
 assign n2509 = ( n1798  &  n909  &  n1800  &  n938  &  n930  &  n925 ) ;
 assign n2510 = ( n1793  &  n1794  &  n1787  &  n1789  &  n1795  &  n942  &  n1797  &  n2509 ) ;
 assign n2512 = ( (~ n47)  &  (~ n71)  &  n1380 ) ;
 assign n2511 = ( (~ n982)  &  (~ n1762) ) | ( (~ n980)  &  (~ n1762) ) | ( (~ n982)  &  n2512 ) | ( (~ n980)  &  n2512 ) ;
 assign n2513 = ( (~ n64)  &  n961  &  n1804 ) ;
 assign n2515 = ( (~ n1366) ) | ( n2512 ) ;
 assign n2514 = ( n491  &  n2515 ) | ( n508  &  (~ n892)  &  n2515 ) ;
 assign n2516 = ( n1006  &  n1605  &  n2032  &  n1005  &  n2204  &  n2205  &  n789  &  n791 ) ;
 assign n2517 = ( n546  &  n1578 ) ;
 assign n2518 = ( n2277  &  n2360  &  n2300 ) ;
 assign n2519 = ( (~ n1021)  &  n2347 ) | ( n815  &  n1565  &  n2347 ) ;
 assign n2520 = ( (~ n135)  &  (~ n280) ) | ( (~ n135)  &  n291 ) | ( (~ n280)  &  n448 ) | ( n291  &  n448 ) ;
 assign n2521 = ( n2380  &  n2130  &  n2394 ) ;
 assign n2522 = ( n2384  &  n2128  &  n2235  &  n2207  &  n2403  &  n2150  &  n2365  &  n2521 ) ;
 assign n2523 = ( n236  &  n2281  &  n2369 ) ;
 assign n2524 = ( (~ n135)  &  (~ n280) ) | ( (~ n135)  &  n1055 ) | ( (~ n280)  &  n1058 ) | ( n1055  &  n1058 ) ;
 assign n2526 = ( n810  &  n1275 ) ;
 assign n2525 = ( (~ n1021)  &  n1566 ) | ( n1566  &  n2526 ) ;
 assign n2528 = ( n2385  &  n2433  &  n2232  &  n2279  &  n2366  &  n2049 ) ;
 assign n2529 = ( n2370  &  n1588  &  n2383 ) ;
 assign n2530 = ( n2193  &  n2095  &  n2286 ) ;
 assign n2531 = ( (~ n136)  &  n1081  &  (~ n1130)  &  (~ n1133)  &  n1230  &  n2114  &  n2192  &  n2530 ) ;
 assign n2534 = ( n88  &  (~ n139)  &  n212 ) | ( n88  &  n212  &  n381 ) ;
 assign n2535 = ( n1107  &  n1925  &  n1933  &  n1098  &  n1940  &  n1124  &  n1917  &  n2534 ) ;
 assign n2536 = ( (~ n17)  &  (~ n21) ) | ( (~ n17)  &  n1184 ) | ( (~ n21)  &  n1196 ) | ( n1184  &  n1196 ) ;
 assign n2539 = ( n1124  &  n1046  &  n1968  &  n874  &  n1301  &  n1795 ) ;
 assign n2540 = ( n743  &  n1526 ) ;
 assign n2541 = ( n2207  &  n2403  &  n1841  &  n2110  &  n1567  &  n2139  &  n1603  &  n803 ) ;
 assign n2543 = ( n2479 ) | ( n1061 ) ;
 assign n2544 = ( (~ n426)  &  (~ n1207) ) | ( n291  &  n1196  &  (~ n1207) ) ;
 assign n2547 = ( (~ n21) ) | ( n1145 ) ;
 assign n2546 = ( n2547  &  n2439  &  n2544 ) ;
 assign n2548 = ( n296  &  n1493 ) | ( n1205  &  n1493 ) | ( n296  &  n1206 ) | ( n1205  &  n1206 ) ;
 assign n2549 = ( (~ n17)  &  (~ n371) ) | ( (~ n24)  &  (~ n371) ) | ( (~ n17)  &  n800 ) | ( (~ n24)  &  n800 ) ;
 assign n2550 = ( (~ n135)  &  (~ n616) ) | ( n260  &  (~ n616) ) | ( (~ n135)  &  n1248 ) | ( n260  &  n1248 ) ;
 assign n2551 = ( n312  &  n324 ) | ( n312  &  (~ n360) ) | ( n324  &  (~ n479) ) | ( (~ n360)  &  (~ n479) ) ;
 assign n2552 = ( (~ n6)  &  n180 ) | ( n180  &  n837 ) | ( (~ n6)  &  n1428 ) | ( n837  &  n1428 ) ;
 assign n2553 = ( n722  &  n579  &  n2552  &  n2551  &  n2550  &  n2549  &  n2548  &  n2546 ) ;
 assign n2554 = ( n1794  &  n76  &  n902  &  n914  &  n807  &  n843  &  n1577  &  n1604 ) ;
 assign n2555 = ( n1176  &  n1152  &  n1197  &  n1282  &  n1925  &  n1203  &  n1872  &  n1087 ) ;
 assign n2556 = ( (~ n300)  &  (~ n1019) ) | ( n707  &  (~ n1019) ) | ( (~ n300)  &  n1253 ) | ( n707  &  n1253 ) ;
 assign n2557 = ( (~ n135)  &  (~ n426) ) | ( (~ n135)  &  n611 ) | ( (~ n426)  &  n1474 ) | ( n611  &  n1474 ) ;
 assign n2558 = ( n1789  &  n1676  &  n1665  &  n1643  &  n2557  &  n2556 ) ;
 assign n2559 = ( n918  &  n2092  &  n728  &  n1631  &  n1630  &  n237 ) ;
 assign n2560 = ( (~ n354)  &  (~ n1238) ) | ( n1007  &  (~ n1238)  &  n1478 ) ;
 assign n2562 = ( (~ n616)  &  (~ n1240) ) | ( (~ n1240)  &  n1329  &  n2011 ) ;
 assign n2564 = ( n1265  &  n2562 ) | ( (~ n39)  &  n2012  &  n2562 ) ;
 assign n2565 = ( (~ n360)  &  (~ n1016) ) | ( (~ n360)  &  n1236 ) | ( (~ n1016)  &  n2011 ) | ( n1236  &  n2011 ) ;
 assign n2566 = ( n263  &  n381 ) | ( n263  &  (~ n400) ) | ( n381  &  n580 ) | ( (~ n400)  &  n580 ) ;
 assign n2567 = ( n295  &  n296 ) | ( n1379  &  n296 ) | ( n295  &  n261 ) | ( n1379  &  n261 ) ;
 assign n2568 = ( n2566  &  n2567  &  n1428 ) | ( n2566  &  n2567  &  n959 ) ;
 assign n2569 = ( n2376  &  n2438  &  n2284  &  n2560  &  n2559  &  n2565  &  n2564  &  n2568 ) ;
 assign n2570 = ( (~ n426)  &  n543  &  n1405 ) | ( n543  &  n768  &  n1405 ) ;
 assign n2571 = ( n1652  &  n811  &  n1669  &  n1772  &  n820  &  n806  &  n1555  &  n2570 ) ;
 assign n2572 = ( n1793  &  n77  &  n1022 ) ;
 assign n2573 = ( n1966  &  n1176  &  n1228  &  n1297  &  n1284  &  n1086  &  n1107  &  n2572 ) ;
 assign n2574 = ( (~ n34) ) | ( n2042 ) ;
 assign n2575 = ( n2300  &  n2089  &  n1049  &  n1611  &  n1601  &  n2356 ) ;
 assign n2576 = ( (~ n616)  &  n1579 ) | ( n1252  &  n1579 ) ;
 assign n2577 = ( n318  &  (~ n426) ) | ( n318  &  n1249 ) | ( (~ n426)  &  n2101 ) | ( n1249  &  n2101 ) ;
 assign n2578 = ( (~ n332)  &  n704 ) | ( n704  &  n1270 ) | ( (~ n332)  &  n1493 ) | ( n1270  &  n1493 ) ;
 assign n2579 = ( (~ n364)  &  n2578 ) | ( n1520  &  n2578 ) ;
 assign n2580 = ( n2577  &  n2579  &  n1820 ) | ( n2577  &  n2579  &  n545 ) ;
 assign n2581 = ( n334  &  (~ n401) ) | ( n334  &  n864 ) | ( (~ n401)  &  n1043 ) | ( n864  &  n1043 ) ;
 assign n2582 = ( (~ n300)  &  n2581 ) | ( n1352  &  n2581 ) ;
 assign n2583 = ( n1411  &  n296 ) | ( n1411  &  n345 ) ;
 assign n2584 = ( n2351  &  n2336  &  n1994  &  n2576  &  n2575  &  n2583  &  n2582  &  n2580 ) ;
 assign n2585 = ( n603  &  n1582  &  n1629  &  n343  &  n441  &  n548 ) ;
 assign n2586 = ( n841  &  n1672  &  n1681  &  n869  &  n1798  &  n2585 ) ;
 assign n2587 = ( n1036  &  n1066  &  n1078 ) ;
 assign n2588 = ( n1152  &  n1228  &  n2033  &  n1296  &  n1241  &  n1098  &  n1185  &  n2587 ) ;
 assign n2589 = ( (~ n18)  &  (~ n28)  &  (~ n31)  &  n1038  &  n1671  &  n2547 ) ;
 assign n2591 = ( (~ n34) ) | ( n1254 ) ;
 assign n2590 = ( (~ n40)  &  n546  &  n2010  &  n2574  &  n2589  &  n2591 ) ;
 assign n2592 = ( (~ n247)  &  (~ n21) ) | ( (~ n247)  &  n1263 ) | ( (~ n21)  &  n1266 ) | ( n1263  &  n1266 ) ;
 assign n2593 = ( (~ n34)  &  n2592 ) | ( n1261  &  n2592 ) ;
 assign n2594 = ( (~ n139)  &  (~ n280) ) | ( (~ n280)  &  n1256 ) | ( (~ n139)  &  n1259 ) | ( n1256  &  n1259 ) ;
 assign n2595 = ( (~ n10)  &  n2594 ) | ( n1258  &  n2594 ) ;
 assign n2596 = ( n382  &  n250  &  n444  &  n729  &  n1559  &  n2595  &  n2593  &  n2590 ) ;
 assign n2597 = ( n790  &  n831  &  n853  &  n685  &  n752  &  n792 ) ;
 assign n2598 = ( n907  &  n1781  &  n917  &  n914  &  n922  &  n2597 ) ;
 assign n2599 = ( n949  &  n946  &  n1785 ) ;
 assign n2600 = ( n1944  &  n1146  &  n1209  &  n2027  &  n2033  &  n1089  &  n1126  &  n2599 ) ;
 assign n2601 = ( n1457  &  n2126  &  n1535 ) ;
 assign n2602 = ( (~ n21)  &  n1273 ) | ( n1273  &  n1278 ) | ( (~ n21)  &  n1428 ) | ( n1278  &  n1428 ) ;
 assign n2603 = ( n2065  &  n1148  &  n678  &  n2373  &  n1454  &  n2285 ) ;
 assign n2604 = ( (~ n300)  &  n2591 ) | ( n1262  &  n1658  &  n2591 ) ;
 assign n2605 = ( n448  &  n373  &  n505 ) ;
 assign n2606 = ( n1329  &  n1007 ) ;
 assign n2607 = ( n193  &  n824 ) ;
 assign n2608 = ( n953  &  n465  &  n921 ) ;
 assign n2609 = ( n263  &  n530  &  n737 ) ;
 assign n2610 = ( n1329  &  n504 ) ;
 assign n2611 = ( n1431  &  n503 ) ;
 assign n2612 = ( n565  &  n195 ) ;
 assign n2613 = ( n959  &  n504 ) ;
 assign n2614 = ( n971 ) | ( n54 ) ;
 assign n2615 = ( n985 ) | ( n54 ) ;
 assign n2616 = ( n510 ) | ( n54 ) ;
 assign n2617 = ( n633 ) | ( n54 ) ;
 assign n2618 = ( (~ i_12_)  &  n204  &  n1328  &  n1392 ) ;


endmodule

