module ex1010x6xv (i_9_, i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_, o_1_, o_2_, o_0_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

	input i_9_;
	input i_7_;
	input i_8_;
	input i_5_;
	input i_6_;
	input i_3_;
	input i_4_;
	input i_1_;
	input i_2_;
	input i_0_;
	output o_1_;
	output o_2_;
	output o_0_;
	output o_9_;
	output o_7_;
	output o_8_;
	output o_5_;
	output o_6_;
	output o_3_;
	output o_4_;

	wire [2889 : 0] sk /* synthesis noprune */;

	lut_sub lut_3 ({sk[0], x12042x, n_n1004, x12041x}, o_1_);
	defparam lut_3.LUT_SIZE = 4;
	defparam lut_3.mask = 16'h0f7f;

	lut_sub lut_7 ({sk[1], n_n1390, n_n1392, x12587x, x12588x}, o_2_);
	defparam lut_7.LUT_SIZE = 5;
	defparam lut_7.mask = 32'h0fff7fff;

	lut_sub lut_12 ({sk[2], x13147x, n_n621, n_n620, n_n630, n_n631, n_n629}, o_0_);
	defparam lut_12.LUT_SIZE = 7;
	defparam lut_12.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_19 ({sk[3], x13684x, x13574x, n_n3990, n_n3992, n_n3988, n_n3987}, o_9_);
	defparam lut_19.LUT_SIZE = 7;
	defparam lut_19.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_26 ({sk[4], x14222x, n_n3257, n_n3259, n_n3251, n_n3253, x14214x}, o_7_);
	defparam lut_26.LUT_SIZE = 7;
	defparam lut_26.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_33 ({sk[5], x14780x, n_n3623, n_n3624, x14775x, x14778x}, o_8_);
	defparam lut_33.LUT_SIZE = 6;
	defparam lut_33.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_39 ({sk[6], x15301x, x15297x, n_n2526, n_n2528, x15300x}, o_5_);
	defparam lut_39.LUT_SIZE = 6;
	defparam lut_39.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_45 ({sk[7], n_n2897, n_n2898, x15815x, x15816x}, o_6_);
	defparam lut_45.LUT_SIZE = 5;
	defparam lut_45.mask = 32'h33ff7fff;

	lut_sub lut_50 ({sk[8], x16324x, x16242x, n_n1789, n_n1790, x16323x}, o_3_);
	defparam lut_50.LUT_SIZE = 6;
	defparam lut_50.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_56 ({sk[9], x16831x, n_n2159, x16744x, x16745x, x16763x, x16830x}, o_4_);
	defparam lut_56.LUT_SIZE = 7;
	defparam lut_56.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_63 ({sk[10], n_n1014, n_n1013, x11894x, n_n1010, n_n1012}, x12042x);
	defparam lut_63.LUT_SIZE = 6;
	defparam lut_63.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_69 ({sk[11], x12038x, n_n1007, n_n1023, n_n1022, x12026x, x12027x}, n_n1004);
	defparam lut_69.LUT_SIZE = 7;
	defparam lut_69.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_76 ({sk[12], n_n1015, x11746x, n_n957, n_n956, n_n937, x11743x}, x12041x);
	defparam lut_76.LUT_SIZE = 7;
	defparam lut_76.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_83 ({sk[13], n_n1394, n_n1393, x12387x, x12388x, x12390x}, n_n1390);
	defparam lut_83.LUT_SIZE = 6;
	defparam lut_83.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_89 ({sk[14], x12585x, n_n1400, x12567x, x12568x}, n_n1392);
	defparam lut_89.LUT_SIZE = 5;
	defparam lut_89.mask = 32'h33ff7fff;

	lut_sub lut_94 ({sk[15], n_n1396, x12248x, n_n1471, n_n1472, x12245x}, x12587x);
	defparam lut_94.LUT_SIZE = 6;
	defparam lut_94.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_100 ({sk[16], x12151x, n_n1398, n_n1321, x12148x, x12149x}, x12588x);
	defparam lut_100.LUT_SIZE = 6;
	defparam lut_100.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_106 ({sk[17], x12693x, x12694x, x13142x, x13143x, x13145x}, x13147x);
	defparam lut_106.LUT_SIZE = 6;
	defparam lut_106.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_112 ({sk[18], x12775x, x12776x, n_n628, x12867x}, n_n621);
	defparam lut_112.LUT_SIZE = 5;
	defparam lut_112.mask = 32'h33ff7fff;

	lut_sub lut_117 ({sk[19], n_n684, n_n683, x12948x, x13001x, x12945x, x13000x}, n_n620);
	defparam lut_117.LUT_SIZE = 7;
	defparam lut_117.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_124 ({sk[20], x13016x, x13017x, x13039x, x13040x, x13046x}, n_n630);
	defparam lut_124.LUT_SIZE = 6;
	defparam lut_124.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_130 ({sk[21], n_n657, x13080x, x13081x, x13086x, x13087x}, n_n631);
	defparam lut_130.LUT_SIZE = 6;
	defparam lut_130.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_136 ({sk[22], x13111x, x13112x, x13123x, x13124x, x13133x}, n_n629);
	defparam lut_136.LUT_SIZE = 6;
	defparam lut_136.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_142 ({sk[23], n_n3916, n_n3936, n_n3935, n_n3937, x13682x}, x13684x);
	defparam lut_142.LUT_SIZE = 6;
	defparam lut_142.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_148 ({sk[24], n_n3989, n_n3993, n_n3995, x13555x, x13569x}, x13574x);
	defparam lut_148.LUT_SIZE = 6;
	defparam lut_148.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_154 ({sk[25], x13213x, x13214x, x13228x, x13229x, x13233x, x13234x}, n_n3990);
	defparam lut_154.LUT_SIZE = 7;
	defparam lut_154.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_161 ({sk[26], x13254x, x13255x, x13269x, x13278x, n_n4078, n_n4077}, n_n3992);
	defparam lut_161.LUT_SIZE = 7;
	defparam lut_161.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_168 ({sk[27], n_n4000, x13318x, x144x, x13315x, x13324x, x13325x}, n_n3988);
	defparam lut_168.LUT_SIZE = 7;
	defparam lut_168.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_175 ({sk[28], x13348x, x13349x, x13364x, x13365x, x13372x, x13373x}, n_n3987);
	defparam lut_175.LUT_SIZE = 7;
	defparam lut_175.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_182 ({sk[29], n_n3207, n_n3187, n_n3206, n_n3205, x14220x}, x14222x);
	defparam lut_182.LUT_SIZE = 6;
	defparam lut_182.mask = 64'h0f7f0f7f7fffffff;

	lut_sub lut_188 ({sk[30], x13843x, x13844x, x13860x, x13861x, x13876x, x13877x}, n_n3257);
	defparam lut_188.LUT_SIZE = 7;
	defparam lut_188.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_195 ({sk[31], x192x, x13896x, x13910x, x13911x, x13919x, x13893x}, n_n3259);
	defparam lut_195.LUT_SIZE = 7;
	defparam lut_195.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_202 ({sk[32], x13976x, x13977x, x14025x, x14067x, x14022x, x14023x}, n_n3251);
	defparam lut_202.LUT_SIZE = 7;
	defparam lut_202.mask = 128'h5577557755ff55ff7fffffffffffffff;

	lut_sub lut_209 ({sk[33], x14117x, x14118x, n_n3262, x14211x}, n_n3253);
	defparam lut_209.LUT_SIZE = 5;
	defparam lut_209.mask = 32'h33ff7fff;

	lut_sub lut_214 ({sk[34], x13796x, x13797x, n_n3275, x13825x, x13826x, x14213x}, x14214x);
	defparam lut_214.LUT_SIZE = 7;
	defparam lut_214.mask = 128'h0fff0fff5fffffff7fffffffffffffff;

	lut_sub lut_221 ({sk[35], x14540x, n_n3625, n_n3627, n_n3629, n_n3631}, x14780x);
	defparam lut_221.LUT_SIZE = 6;
	defparam lut_221.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_227 ({sk[36], n_n3632, x14582x, x14583x, x14589x, x14590x}, n_n3623);
	defparam lut_227.LUT_SIZE = 6;
	defparam lut_227.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_233 ({sk[37], n_n3674, n_n3673, n_n3637, n_n3635, x14636x}, n_n3624);
	defparam lut_233.LUT_SIZE = 6;
	defparam lut_233.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_239 ({sk[38], x14388x, x14357x, x14358x, n_n3649, x14774x}, x14775x);
	defparam lut_239.LUT_SIZE = 6;
	defparam lut_239.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_245 ({sk[39], n_n3626, x14277x, x14278x, x14341x, x14342x}, x14778x);
	defparam lut_245.LUT_SIZE = 6;
	defparam lut_245.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_251 ({sk[40], n_n2530, n_n2529, x15169x, n_n2533, x15150x, x15151x}, x15301x);
	defparam lut_251.LUT_SIZE = 7;
	defparam lut_251.mask = 128'h0fff0fff5fffffff7fffffffffffffff;

	lut_sub lut_258 ({sk[41], x15221x, x15222x, x15278x, x15279x, x15295x}, x15297x);
	defparam lut_258.LUT_SIZE = 6;
	defparam lut_258.mask = 64'h3f3f3f3f7fffffff;

	lut_sub lut_264 ({sk[42], n_n2568, n_n2569, x15184x, n_n2535, x15204x, x15205x}, n_n2526);
	defparam lut_264.LUT_SIZE = 7;
	defparam lut_264.mask = 128'h0fff0fff5fffffff7fffffffffffffff;

	lut_sub lut_271 ({sk[43], x15234x, x15235x, x15249x, x15262x, x22136x}, n_n2528);
	defparam lut_271.LUT_SIZE = 6;
	defparam lut_271.mask = 64'h3f3f3f3fbfffffff;

	lut_sub lut_277 ({sk[44], n_n2449, n_n2531, x14888x, x14889x, x14891x}, x15300x);
	defparam lut_277.LUT_SIZE = 6;
	defparam lut_277.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_283 ({sk[45], x15594x, x15595x, x15642x, x15643x, x15674x, x15675x}, n_n2897);
	defparam lut_283.LUT_SIZE = 7;
	defparam lut_283.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_290 ({sk[46], x15808x, x15743x, n_n2905, x15740x, x15741x}, n_n2898);
	defparam lut_290.LUT_SIZE = 6;
	defparam lut_290.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_296 ({sk[47], x15504x, n_n2908, n_n2993, n_n2992, x15501x}, x15815x);
	defparam lut_296.LUT_SIZE = 6;
	defparam lut_296.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_302 ({sk[48], x15401x, n_n2907, x15812x, x22106x}, x15816x);
	defparam lut_302.LUT_SIZE = 5;
	defparam lut_302.mask = 32'h0fffbfff;

	lut_sub lut_307 ({sk[49], n_n1793, n_n1792, n_n1794, n_n1787}, x16324x);
	defparam lut_307.LUT_SIZE = 5;
	defparam lut_307.mask = 32'h0fff7fff;

	lut_sub lut_312 ({sk[50], n_n1810, n_n1870, x16144x, x16239x, x22094x}, x16242x);
	defparam lut_312.LUT_SIZE = 6;
	defparam lut_312.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_318 ({sk[51], x16157x, x16158x, x16168x, x16169x, x16180x}, n_n1789);
	defparam lut_318.LUT_SIZE = 6;
	defparam lut_318.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_324 ({sk[52], x16198x, x16199x, x16213x, x16214x, x16222x, x16223x}, n_n1790);
	defparam lut_324.LUT_SIZE = 7;
	defparam lut_324.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_331 ({sk[53], n_n1788, x15902x, x15903x, x15942x, x22083x}, x16323x);
	defparam lut_331.LUT_SIZE = 6;
	defparam lut_331.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_337 ({sk[54], n_n2165, n_n2164, n_n2162, n_n2163, x16468x, x16469x}, x16831x);
	defparam lut_337.LUT_SIZE = 7;
	defparam lut_337.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_344 ({sk[55], x16683x, x16697x, x16703x, x16704x, x22071x}, n_n2159);
	defparam lut_344.LUT_SIZE = 6;
	defparam lut_344.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_350 ({sk[56], n_n4161, x14661x, n_n2214, x253x, x16742x}, x16744x);
	defparam lut_350.LUT_SIZE = 6;
	defparam lut_350.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_356 ({sk[57], n_n2209, x16715x, x16730x, x16714x, x22068x}, x16745x);
	defparam lut_356.LUT_SIZE = 6;
	defparam lut_356.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_362 ({sk[58], x16662x, x16758x, x16759x, x22066x}, x16763x);
	defparam lut_362.LUT_SIZE = 5;
	defparam lut_362.mask = 32'h0fffbfff;

	lut_sub lut_367 ({sk[59], n_n2166, x16823x, x16826x, x22058x}, x16830x);
	defparam lut_367.LUT_SIZE = 5;
	defparam lut_367.mask = 32'h0fffbfff;

	lut_sub lut_372 ({sk[60], x11501x, x11502x, x11518x, x11519x, x11528x, x11529x}, n_n1014);
	defparam lut_372.LUT_SIZE = 7;
	defparam lut_372.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_379 ({sk[61], x11581x, n_n1099, x11558x, x11574x, x11575x, x11557x}, n_n1013);
	defparam lut_379.LUT_SIZE = 7;
	defparam lut_379.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_386 ({sk[62], n_n1029, x11781x, x11782x, x11890x, x11891x}, x11894x);
	defparam lut_386.LUT_SIZE = 6;
	defparam lut_386.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_392 ({sk[63], x11796x, x11797x, n_n1071, n_n1072, x11815x, x11832x}, n_n1010);
	defparam lut_392.LUT_SIZE = 7;
	defparam lut_392.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_399 ({sk[64], x11851x, x11852x, x11875x, x11876x, x11882x, x11883x}, n_n1012);
	defparam lut_399.LUT_SIZE = 7;
	defparam lut_399.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_406 ({sk[65], n_n553, n_n554, x12691x}, x12693x);
	defparam lut_406.LUT_SIZE = 4;
	defparam lut_406.mask = 16'h5f7f;

	lut_sub lut_410 ({sk[66], n_n546, n_n547, x12649x, x12672x, x12673x}, x12694x);
	defparam lut_410.LUT_SIZE = 6;
	defparam lut_410.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_416 ({sk[67], x12699x, x13140x, x22216x, x22341x}, x13142x);
	defparam lut_416.LUT_SIZE = 5;
	defparam lut_416.mask = 32'h0fffefff;

	lut_sub lut_421 ({sk[68], x12707x, x12714x, x12706x, x12713x, x22215x}, x13143x);
	defparam lut_421.LUT_SIZE = 6;
	defparam lut_421.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_427 ({sk[69], x12609x, x12629x, n_n555, n_n557, n_n559, n_n558}, x13145x);
	defparam lut_427.LUT_SIZE = 7;
	defparam lut_427.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_434 ({sk[70], n_n3923, n_n3928, n_n3927, x13613x, x13614x}, n_n3916);
	defparam lut_434.LUT_SIZE = 6;
	defparam lut_434.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_440 ({sk[71], x500x, x11x, x23x, x499x, x13622x, x22197x}, n_n3936);
	defparam lut_440.LUT_SIZE = 7;
	defparam lut_440.mask = 128'h777f777f777f777fbbbfbbbfbbbfffff;

	lut_sub lut_445 ({sk[72], x15x, x495x, x22196x, x22315x}, n_n3935);
	defparam lut_445.LUT_SIZE = 5;
	defparam lut_445.mask = 32'h0fffeeef;

	lut_sub lut_449 ({sk[73], x13678x, x16x, x474x, x478x, x536x, x124x}, n_n3937);
	defparam lut_449.LUT_SIZE = 7;
	defparam lut_449.mask = 128'h777f777f777f777f55557fffffffffff;

	lut_sub lut_455 ({sk[74], x13645x, x13665x, n_n3931, n_n3929, n_n3933, n_n3932}, x13682x);
	defparam lut_455.LUT_SIZE = 7;
	defparam lut_455.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_462 ({sk[75], x20x, x499x, x13687x, x13688x, x22323x}, n_n3207);
	defparam lut_462.LUT_SIZE = 6;
	defparam lut_462.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_467 ({sk[76], n_n3196, n_n3194, x13714x, n_n3197, x13728x}, n_n3187);
	defparam lut_467.LUT_SIZE = 6;
	defparam lut_467.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_473 ({sk[77], x13x, x472x, x559x, x13731x, x13732x, x13734x}, n_n3206);
	defparam lut_473.LUT_SIZE = 7;
	defparam lut_473.mask = 128'h777f777f777f777f7f7f7f7f7fffffff;

	lut_sub lut_479 ({sk[78], x22x, x504x, x471x, x13739x, x22179x}, n_n3205);
	defparam lut_479.LUT_SIZE = 6;
	defparam lut_479.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_484 ({sk[79], x13761x, x13782x, n_n3202, n_n3204, n_n3199, n_n3201}, x14220x);
	defparam lut_484.LUT_SIZE = 7;
	defparam lut_484.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_491 ({sk[80], x14458x, x14459x, x14530x, n_n3729, n_n3731, x14538x}, x14540x);
	defparam lut_491.LUT_SIZE = 7;
	defparam lut_491.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_498 ({sk[81], n_n3679, n_n3678, x14654x, x14668x, x22339x}, n_n3625);
	defparam lut_498.LUT_SIZE = 6;
	defparam lut_498.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_504 ({sk[82], x14730x, x14710x, x14711x, x14722x, x14723x}, n_n3627);
	defparam lut_504.LUT_SIZE = 6;
	defparam lut_504.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_510 ({sk[83], x14405x, x14406x, x14419x, x14420x, x14436x}, n_n3629);
	defparam lut_510.LUT_SIZE = 6;
	defparam lut_510.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_516 ({sk[84], n_n3737, n_n3736, n_n3658, x14507x, x14508x, x14511x}, n_n3631);
	defparam lut_516.LUT_SIZE = 7;
	defparam lut_516.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_523 ({sk[85], x14935x, x14928x, n_n2601, n_n2602, x22145x}, n_n2530);
	defparam lut_523.LUT_SIZE = 6;
	defparam lut_523.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_529 ({sk[86], x14960x, x14961x, x14974x, x14975x, x14979x, x14980x}, n_n2529);
	defparam lut_529.LUT_SIZE = 7;
	defparam lut_529.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_536 ({sk[87], n_n2637, n_n2638, n_n2559, x15038x, x15039x, x15167x}, x15169x);
	defparam lut_536.LUT_SIZE = 7;
	defparam lut_536.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_543 ({sk[88], x15075x, x15076x, n_n2557, x15101x, x15102x}, n_n2533);
	defparam lut_543.LUT_SIZE = 6;
	defparam lut_543.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_549 ({sk[89], x471x, x82x, x222x, x15149x, x22253x}, x15150x);
	defparam lut_549.LUT_SIZE = 6;
	defparam lut_549.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_555 ({sk[90], x15140x, x15141x, n_n2619, n_n2618, x15119x, x15120x}, x15151x);
	defparam lut_555.LUT_SIZE = 7;
	defparam lut_555.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_562 ({sk[91], x16027x, x16008x, x16018x, x16019x, x16004x, x16005x}, n_n1793);
	defparam lut_562.LUT_SIZE = 7;
	defparam lut_562.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_569 ({sk[92], n_n1813, x16065x, x16066x, x16070x, x16071x}, n_n1792);
	defparam lut_569.LUT_SIZE = 6;
	defparam lut_569.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_575 ({sk[93], x16114x, n_n1896, x16086x, x16105x, x16106x, x16085x}, n_n1794);
	defparam lut_575.LUT_SIZE = 7;
	defparam lut_575.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_582 ({sk[94], x16289x, x16262x, x16263x, n_n1828, n_n1829, x16280x}, n_n1787);
	defparam lut_582.LUT_SIZE = 7;
	defparam lut_582.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_589 ({sk[95], x16598x, x16570x, x16590x, n_n2253, x22081x}, n_n2165);
	defparam lut_589.LUT_SIZE = 6;
	defparam lut_589.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_595 ({sk[96], n_n2251, n_n2250, n_n2185, x16637x, x16638x, x16643x}, n_n2164);
	defparam lut_595.LUT_SIZE = 7;
	defparam lut_595.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_602 ({sk[97], x16342x, x16343x, x16364x, x16365x, x16374x, x16375x}, n_n2162);
	defparam lut_602.LUT_SIZE = 7;
	defparam lut_602.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_609 ({sk[98], x16399x, x16400x, x16415x, x16416x, x16423x, x16424x}, n_n2163);
	defparam lut_609.LUT_SIZE = 7;
	defparam lut_609.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_616 ({sk[99], n_n3803, n_n3805, x16327x, n_n2220, x16466x}, x16468x);
	defparam lut_616.LUT_SIZE = 6;
	defparam lut_616.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_622 ({sk[100], x16442x, x16443x, x16456x, x16457x}, x16469x);
	defparam lut_622.LUT_SIZE = 5;
	defparam lut_622.mask = 32'h0fff7fff;

	lut_sub lut_627 ({sk[101], x13x, x562x, x130x, n_n4246, x22249x}, x11501x);
	defparam lut_627.LUT_SIZE = 6;
	defparam lut_627.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_632 ({sk[102], x65x, n_n1107, x307x, x11497x}, x11502x);
	defparam lut_632.LUT_SIZE = 5;
	defparam lut_632.mask = 32'h0fff7fff;

	lut_sub lut_637 ({sk[103], x24x, x476x, x194x, n_n1285, x11516x}, x11518x);
	defparam lut_637.LUT_SIZE = 6;
	defparam lut_637.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_642 ({sk[104], x22x, x476x, x184x, n_n1111, x11511x, x11510x}, x11519x);
	defparam lut_642.LUT_SIZE = 7;
	defparam lut_642.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_648 ({sk[105], x20x, x23x, x495x, x11525x, x11526x}, x11528x);
	defparam lut_648.LUT_SIZE = 6;
	defparam lut_648.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_653 ({sk[106], n_n1112, x235x, x421x, x22248x}, x11529x);
	defparam lut_653.LUT_SIZE = 5;
	defparam lut_653.mask = 32'h0fffbfff;

	lut_sub lut_658 ({sk[107], x25x, x13x, x509x, x24x, x504x}, n_n4243);
	defparam lut_658.LUT_SIZE = 6;
	defparam lut_658.mask = 64'h77ff77ff111f555f;

	lut_sub lut_662 ({sk[108], i_9_, i_7_, i_8_, i_6_, n_n455, n_n473}, n_n1104);
	defparam lut_662.LUT_SIZE = 7;
	defparam lut_662.mask = 128'h777f777f777f777f1111101001010010;

	lut_sub lut_672 ({sk[109], i_9_, i_7_, i_8_, i_6_, n_n455, n_n464}, n_n1103);
	defparam lut_672.LUT_SIZE = 7;
	defparam lut_672.mask = 128'h777f777f777f777f0101011101010101;

	lut_sub lut_682 ({sk[110], x13x, x20x, x23x, x580x, x543x}, n_n3875);
	defparam lut_682.LUT_SIZE = 6;
	defparam lut_682.mask = 64'h77ff77ff05553777;

	lut_sub lut_686 ({sk[111], x15x, x538x, x22x, x13x, x543x}, x11577x);
	defparam lut_686.LUT_SIZE = 6;
	defparam lut_686.mask = 64'h77ff77ff05375577;

	lut_sub lut_690 ({sk[112], n_n4243, n_n1104, n_n1103, n_n3875, x11577x}, x11581x);
	defparam lut_690.LUT_SIZE = 6;
	defparam lut_690.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_696 ({sk[113], x10x, x472x, x563x, n_n4611, n_n4232, x22250x}, n_n1099);
	defparam lut_696.LUT_SIZE = 7;
	defparam lut_696.mask = 128'h777f777f777f777fbfbfbfbfbfffffff;

	lut_sub lut_702 ({sk[114], x10x, x518x, x309x, n_n3861, x11555x}, x11558x);
	defparam lut_702.LUT_SIZE = 6;
	defparam lut_702.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_707 ({sk[115], x13x, x516x, x525x, x471x, x222x, x22247x}, x11574x);
	defparam lut_707.LUT_SIZE = 7;
	defparam lut_707.mask = 128'h777f777f777f777fbfbfbfbfbfffffff;

	lut_sub lut_713 ({sk[116], x11562x, x11563x, x11570x, x11571x}, x11575x);
	defparam lut_713.LUT_SIZE = 5;
	defparam lut_713.mask = 32'h0fff7fff;

	lut_sub lut_718 ({sk[117], x11x, x10x, x519x, x571x, x119x, x11554x}, x11557x);
	defparam lut_718.LUT_SIZE = 7;
	defparam lut_718.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_723 ({sk[118], x25x, x15x, x500x, n_n4391, x93x, x11602x}, x11604x);
	defparam lut_723.LUT_SIZE = 7;
	defparam lut_723.mask = 128'h777f777f777f777f7f7f7fff7fff7fff;

	lut_sub lut_729 ({sk[119], x16x, x580x, n_n1117, x22242x, x22261x}, x11605x);
	defparam lut_729.LUT_SIZE = 6;
	defparam lut_729.mask = 64'h77ff77ffefefefff;

	lut_sub lut_734 ({sk[120], x300x, n_n1120, n_n3176, x11618x, x161x}, n_n1041);
	defparam lut_734.LUT_SIZE = 6;
	defparam lut_734.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_740 ({sk[121], x16x, x517x, x198x, x410x, x22241x}, x11632x);
	defparam lut_740.LUT_SIZE = 6;
	defparam lut_740.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_745 ({sk[122], x25x, x473x, n_n1123, x11626x, x22262x}, x11633x);
	defparam lut_745.LUT_SIZE = 6;
	defparam lut_745.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_750 ({sk[123], x11604x, x11605x, n_n1041, x11632x, x11633x}, n_n1015);
	defparam lut_750.LUT_SIZE = 6;
	defparam lut_750.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_756 ({sk[124], x25x, x15x, x571x, x479x, x11640x, x22240x}, n_n954);
	defparam lut_756.LUT_SIZE = 7;
	defparam lut_756.mask = 128'h777f777f777f777fbbbbbfbfbbffbfff;

	lut_sub lut_761 ({sk[125], x21x, x595x, x193x, x312x, x11644x, x11645x}, n_n953);
	defparam lut_761.LUT_SIZE = 7;
	defparam lut_761.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_767 ({sk[126], x11x, x543x, x99x, x11651x, x22239x}, x11655x);
	defparam lut_767.LUT_SIZE = 6;
	defparam lut_767.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_772 ({sk[127], x14x, x478x, x11675x, x22266x}, n_n952);
	defparam lut_772.LUT_SIZE = 5;
	defparam lut_772.mask = 32'h0fffbbbf;

	lut_sub lut_776 ({sk[128], x23x, x553x, x11685x, x11687x, x22267x}, x11690x);
	defparam lut_776.LUT_SIZE = 6;
	defparam lut_776.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_781 ({sk[129], x17x, x585x, x303x, x11678x, x22238x}, n_n951);
	defparam lut_781.LUT_SIZE = 6;
	defparam lut_781.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_786 ({sk[130], n_n954, n_n953, x11655x, n_n952, x11690x, n_n951}, x11746x);
	defparam lut_786.LUT_SIZE = 7;
	defparam lut_786.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_793 ({sk[131], n_n2003, x11756x, x11757x, n_n1082, x11763x, x11764x}, n_n1029);
	defparam lut_793.LUT_SIZE = 7;
	defparam lut_793.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_800 ({sk[132], x17x, x546x, n_n3460, x177x, x11778x}, x11781x);
	defparam lut_800.LUT_SIZE = 6;
	defparam lut_800.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_805 ({sk[133], x539x, x17x, x11772x, x185x, x11777x, x22246x}, x11782x);
	defparam lut_805.LUT_SIZE = 7;
	defparam lut_805.mask = 128'h777f777f777f777fbfffbfffbfffffff;

	lut_sub lut_811 ({sk[134], x14x, x558x, x520x, x11887x, x11888x}, x11890x);
	defparam lut_811.LUT_SIZE = 6;
	defparam lut_811.mask = 64'h77ff77ff77777fff;

	lut_sub lut_816 ({sk[135], n_n1086, x11836x, n_n4210, x11835x}, x11891x);
	defparam lut_816.LUT_SIZE = 5;
	defparam lut_816.mask = 32'h0fff7fff;

	lut_sub lut_821 ({sk[136], x510x, x12x, x508x, x114x, x44x, x11905x}, x11908x);
	defparam lut_821.LUT_SIZE = 7;
	defparam lut_821.mask = 128'h777f777f777f777f7f7f7fff7f7fffff;

	lut_sub lut_827 ({sk[137], x11899x, x11897x, x11898x, x11903x, x11904x}, x11909x);
	defparam lut_827.LUT_SIZE = 6;
	defparam lut_827.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_833 ({sk[138], x24x, x555x, x220x, x11973x, x11975x}, x11977x);
	defparam lut_833.LUT_SIZE = 6;
	defparam lut_833.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_838 ({sk[139], x11967x, n_n1927, x11970x, x11969x, x22245x}, x11978x);
	defparam lut_838.LUT_SIZE = 6;
	defparam lut_838.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_844 ({sk[140], x23x, x568x, x125x, x12030x, x12032x}, x12034x);
	defparam lut_844.LUT_SIZE = 6;
	defparam lut_844.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_849 ({sk[141], x11912x, x11913x, x11914x, x11915x, x11918x}, x12035x);
	defparam lut_849.LUT_SIZE = 6;
	defparam lut_849.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_855 ({sk[142], x11908x, x11909x, x11977x, x11978x, x12034x, x12035x}, x12038x);
	defparam lut_855.LUT_SIZE = 7;
	defparam lut_855.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_862 ({sk[143], n_n1017, n_n1045, x11953x, x11958x, x11959x, x11961x}, n_n1007);
	defparam lut_862.LUT_SIZE = 7;
	defparam lut_862.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_869 ({sk[144], x11993x, n_n1066, x12003x, x11988x, x11989x}, n_n1023);
	defparam lut_869.LUT_SIZE = 6;
	defparam lut_869.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_875 ({sk[145], n_n1061, x12014x, x12018x, x12019x, x22244x}, n_n1022);
	defparam lut_875.LUT_SIZE = 6;
	defparam lut_875.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_881 ({sk[146], x18x, x477x, x581x, x12023x, x12024x}, x12026x);
	defparam lut_881.LUT_SIZE = 6;
	defparam lut_881.mask = 64'h77ff77ff77777fff;

	lut_sub lut_886 ({sk[147], x248x, x299x, x11986x, x11987x, x22243x}, x12027x);
	defparam lut_886.LUT_SIZE = 6;
	defparam lut_886.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_892 ({sk[148], x10x, x572x, x172x, x12048x, x12046x}, n_n1338);
	defparam lut_892.LUT_SIZE = 6;
	defparam lut_892.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_897 ({sk[149], x16x, x489x, x184x, n_n4458, x12050x, x12052x}, n_n1340);
	defparam lut_897.LUT_SIZE = 7;
	defparam lut_897.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_903 ({sk[150], x13x, x562x, x12060x, x22270x}, x12062x);
	defparam lut_903.LUT_SIZE = 5;
	defparam lut_903.mask = 32'h0fffbbbf;

	lut_sub lut_907 ({sk[151], x11x, x565x, x350x, x12066x, x22225x}, n_n1336);
	defparam lut_907.LUT_SIZE = 6;
	defparam lut_907.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_912 ({sk[152], x14x, x517x, x594x, x12074x, x22255x}, n_n1337);
	defparam lut_912.LUT_SIZE = 6;
	defparam lut_912.mask = 64'h77ff77ffbbbbbfff;

	lut_sub lut_917 ({sk[153], x23x, x530x, x12081x, x22289x}, x12083x);
	defparam lut_917.LUT_SIZE = 5;
	defparam lut_917.mask = 32'h0fffbbbf;

	lut_sub lut_921 ({sk[154], n_n1338, n_n1340, x12062x, n_n1336, n_n1337, x12083x}, x12151x);
	defparam lut_921.LUT_SIZE = 7;
	defparam lut_921.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_928 ({sk[155], x210x, x12165x, x142x, x12161x, x12174x, x12175x}, n_n1412);
	defparam lut_928.LUT_SIZE = 7;
	defparam lut_928.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_935 ({sk[156], n_n3810, n_n1592, x12188x}, x12191x);
	defparam lut_935.LUT_SIZE = 4;
	defparam lut_935.mask = 16'h5f7f;

	lut_sub lut_939 ({sk[157], x353x, x306x, x12181x, x12182x, x12187x}, x12192x);
	defparam lut_939.LUT_SIZE = 6;
	defparam lut_939.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_945 ({sk[158], x15x, x597x, x342x, x362x, x22286x}, x12197x);
	defparam lut_945.LUT_SIZE = 6;
	defparam lut_945.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_950 ({sk[159], n_n1576, x12155x, x12159x, x12154x, x22227x}, x12198x);
	defparam lut_950.LUT_SIZE = 6;
	defparam lut_950.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_956 ({sk[160], n_n1412, x12191x, x12192x, x12197x, x12198x}, n_n1396);
	defparam lut_956.LUT_SIZE = 6;
	defparam lut_956.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_962 ({sk[161], x21x, x484x, x23x, x12216x, x12221x}, x12223x);
	defparam lut_962.LUT_SIZE = 6;
	defparam lut_962.mask = 64'h77ff77ff777f77ff;

	lut_sub lut_967 ({sk[162], x12213x, x12214x, x12218x, x12219x}, x12224x);
	defparam lut_967.LUT_SIZE = 5;
	defparam lut_967.mask = 32'h0fff7fff;

	lut_sub lut_972 ({sk[163], x22x, x530x, n_n4824, x185x, x186x, n_n4196}, x12240x);
	defparam lut_972.LUT_SIZE = 7;
	defparam lut_972.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_978 ({sk[164], x21x, x596x, x372x, n_n1468, x12235x, x12233x}, x12241x);
	defparam lut_978.LUT_SIZE = 7;
	defparam lut_978.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_984 ({sk[165], x12223x, x12224x, x12240x, x12241x}, x12248x);
	defparam lut_984.LUT_SIZE = 5;
	defparam lut_984.mask = 32'h0fff7fff;

	lut_sub lut_989 ({sk[166], x12282x, x12283x, n_n1406, x12303x, x12304x}, n_n1394);
	defparam lut_989.LUT_SIZE = 6;
	defparam lut_989.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_995 ({sk[167], n_n1435, n_n1436, x12359x, n_n1402, x12379x, x12380x}, n_n1393);
	defparam lut_995.LUT_SIZE = 7;
	defparam lut_995.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1002 ({sk[168], x23x, x577x, n_n1570, x253x, x22280x}, x12387x);
	defparam lut_1002.LUT_SIZE = 6;
	defparam lut_1002.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1007 ({sk[169], x519x, x18x, n_n5017, x12252x, n_n1454, x12251x}, x12388x);
	defparam lut_1007.LUT_SIZE = 7;
	defparam lut_1007.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_1013 ({sk[170], n_n1446, x12324x, x12325x, n_n1448, x12340x}, x12390x);
	defparam lut_1013.LUT_SIZE = 6;
	defparam lut_1013.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1019 ({sk[171], i_9_, i_7_, i_8_, i_6_, n_n325, n_n491}, n_n1473);
	defparam lut_1019.LUT_SIZE = 7;
	defparam lut_1019.mask = 128'h777f777f777f777f0011101001101110;

	lut_sub lut_1029 ({sk[172], i_9_, n_n524, n_n534, n_n509, n_n325, n_n500}, x12399x);
	defparam lut_1029.LUT_SIZE = 7;
	defparam lut_1029.mask = 128'h777f777f777f777f0011031300110313;

	lut_sub lut_1034 ({sk[173], i_9_, i_7_, i_8_, i_6_, n_n509, n_n325}, x12400x);
	defparam lut_1034.LUT_SIZE = 7;
	defparam lut_1034.mask = 128'h777f777f777f777f0110000001100010;

	lut_sub lut_1040 ({sk[174], x21x, x14x, x565x, x536x}, x12434x);
	defparam lut_1040.LUT_SIZE = 5;
	defparam lut_1040.mask = 32'h0fff0537;

	lut_sub lut_1043 ({sk[175], x25x, x24x, x14x, x565x, x562x, x575x}, x12435x);
	defparam lut_1043.LUT_SIZE = 7;
	defparam lut_1043.mask = 128'h777f777f777f777f00330f3f55775f7f;

	lut_sub lut_1047 ({sk[176], x15x, x14x, x20x, x518x, x565x, x574x}, x12436x);
	defparam lut_1047.LUT_SIZE = 7;
	defparam lut_1047.mask = 128'h777f777f777f777f00335f7f33337f7f;

	lut_sub lut_1052 ({sk[177], n_n1473, x12399x, x12400x, x12434x, x12435x, x12436x}, x12440x);
	defparam lut_1052.LUT_SIZE = 7;
	defparam lut_1052.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1059 ({sk[178], x12414x, x12415x}, x12416x);
	defparam lut_1059.LUT_SIZE = 3;
	defparam lut_1059.mask = 8'h17;

	lut_sub lut_1062 ({sk[179], i_9_, i_7_, i_8_, i_6_, n_n390, n_n464}, x12431x);
	defparam lut_1062.LUT_SIZE = 7;
	defparam lut_1062.mask = 128'h777f777f777f777f0111001010111010;

	lut_sub lut_1072 ({sk[180], n_n1636, x12420x, x12425x, x12424x, x22224x}, x12432x);
	defparam lut_1072.LUT_SIZE = 6;
	defparam lut_1072.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_1078 ({sk[181], x14x, x548x, x86x, x12404x, x12402x}, n_n1478);
	defparam lut_1078.LUT_SIZE = 6;
	defparam lut_1078.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_1083 ({sk[182], x22x, x595x, x101x, x12406x, x22223x}, n_n1476);
	defparam lut_1083.LUT_SIZE = 6;
	defparam lut_1083.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1088 ({sk[183], x12440x, x12416x, x12431x, x12432x, n_n1478, n_n1476}, n_n1398);
	defparam lut_1088.LUT_SIZE = 7;
	defparam lut_1088.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1095 ({sk[184], x25x, x498x, x12453x, x22283x}, x12455x);
	defparam lut_1095.LUT_SIZE = 5;
	defparam lut_1095.mask = 32'h0fffbbbf;

	lut_sub lut_1099 ({sk[185], x12445x, x27x, x12443x, x12444x, x12451x}, x12456x);
	defparam lut_1099.LUT_SIZE = 6;
	defparam lut_1099.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1105 ({sk[186], x15x, x22x, x11x, x496x, n_n2803, x12466x}, x12469x);
	defparam lut_1105.LUT_SIZE = 7;
	defparam lut_1105.mask = 128'h777f777f777f777f777f7f7f7f7f7f7f;

	lut_sub lut_1111 ({sk[187], x12459x, x12457x, x12458x, x12464x, x12465x}, x12470x);
	defparam lut_1111.LUT_SIZE = 6;
	defparam lut_1111.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1117 ({sk[188], x16x, x594x, x585x, x410x, x106x, n_n1703}, x12581x);
	defparam lut_1117.LUT_SIZE = 7;
	defparam lut_1117.mask = 128'h777f777f777f777f7f7f7f7f7fffffff;

	lut_sub lut_1123 ({sk[189], x16x, x482x, n_n4341, x12572x, n_n1508, x448x}, x12582x);
	defparam lut_1123.LUT_SIZE = 7;
	defparam lut_1123.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_1129 ({sk[190], x12455x, x12456x, x12469x, x12470x, x12581x, x12582x}, x12585x);
	defparam lut_1129.LUT_SIZE = 7;
	defparam lut_1129.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1136 ({sk[191], x12485x, x12486x, n_n1495, n_n1496, n_n1423, x12515x}, n_n1400);
	defparam lut_1136.LUT_SIZE = 7;
	defparam lut_1136.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1143 ({sk[192], x24x, x479x, n_n4599, n_n2036, x12563x, x12566x}, x12567x);
	defparam lut_1143.LUT_SIZE = 7;
	defparam lut_1143.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_1149 ({sk[193], n_n1489, x12534x, x12559x, x12560x, x12533x}, x12568x);
	defparam lut_1149.LUT_SIZE = 6;
	defparam lut_1149.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1155 ({sk[194], i_9_, i_7_, i_8_, i_6_}, x25x);
	defparam lut_1155.LUT_SIZE = 5;
	defparam lut_1155.mask = 32'h0fff0100;

	lut_sub lut_1157 ({sk[195], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x515x);
	defparam lut_1157.LUT_SIZE = 7;
	defparam lut_1157.mask = 128'h777f777f777f777f0000000080000000;

	lut_sub lut_1159 ({sk[196], i_9_, i_7_, i_8_, i_6_}, x15x);
	defparam lut_1159.LUT_SIZE = 5;
	defparam lut_1159.mask = 32'h0fff1000;

	lut_sub lut_1161 ({sk[197], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x592x);
	defparam lut_1161.LUT_SIZE = 7;
	defparam lut_1161.mask = 128'h777f777f777f777f0080000000000000;

	lut_sub lut_1163 ({sk[198], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x538x);
	defparam lut_1163.LUT_SIZE = 7;
	defparam lut_1163.mask = 128'h777f777f777f777f0000000000004000;

	lut_sub lut_1165 ({sk[199], i_9_, i_1_, i_2_, i_0_}, x19x);
	defparam lut_1165.LUT_SIZE = 5;
	defparam lut_1165.mask = 32'h0fff0080;

	lut_sub lut_1167 ({sk[200], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x492x);
	defparam lut_1167.LUT_SIZE = 7;
	defparam lut_1167.mask = 128'h777f777f777f777f0000004000000000;

	lut_sub lut_1169 ({sk[201], i_9_, i_1_, i_2_, i_0_}, x10x);
	defparam lut_1169.LUT_SIZE = 5;
	defparam lut_1169.mask = 32'h0fff0010;

	lut_sub lut_1171 ({sk[202], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x548x);
	defparam lut_1171.LUT_SIZE = 7;
	defparam lut_1171.mask = 128'h777f777f777f777f0000000100000000;

	lut_sub lut_1173 ({sk[203], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x523x);
	defparam lut_1173.LUT_SIZE = 7;
	defparam lut_1173.mask = 128'h777f777f777f777f0400000000000000;

	lut_sub lut_1175 ({sk[204], x538x, x13x, x20x, x504x}, x12605x);
	defparam lut_1175.LUT_SIZE = 5;
	defparam lut_1175.mask = 32'h0fff111f;

	lut_sub lut_1178 ({sk[205], x21x, x11x, x24x, x543x, x504x, x523x}, x22214x);
	defparam lut_1178.LUT_SIZE = 7;
	defparam lut_1178.mask = 128'h777f777f777f777fff80aa80f080a080;

	lut_sub lut_1184 ({sk[206], x15x, x10x, x548x, x523x, x12605x, x22214x}, x12609x);
	defparam lut_1184.LUT_SIZE = 7;
	defparam lut_1184.mask = 128'h777f777f777f777fbbbbbbffbfbfbfff;

	lut_sub lut_1189 ({sk[207], i_9_, i_1_, i_2_, i_0_}, x14x);
	defparam lut_1189.LUT_SIZE = 5;
	defparam lut_1189.mask = 32'h0fff0040;

	lut_sub lut_1191 ({sk[208], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x475x);
	defparam lut_1191.LUT_SIZE = 7;
	defparam lut_1191.mask = 128'h777f777f777f777f0000000000000020;

	lut_sub lut_1193 ({sk[209], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x556x);
	defparam lut_1193.LUT_SIZE = 7;
	defparam lut_1193.mask = 128'h777f777f777f777f0200000000000000;

	lut_sub lut_1195 ({sk[210], i_9_, i_7_, i_8_, i_6_, x483x, x595x}, x12623x);
	defparam lut_1195.LUT_SIZE = 7;
	defparam lut_1195.mask = 128'h777f777f777f777f5003000000000000;

	lut_sub lut_1198 ({sk[211], i_9_, i_1_, i_2_, i_0_, x481x, x559x}, x12624x);
	defparam lut_1198.LUT_SIZE = 7;
	defparam lut_1198.mask = 128'h777f777f777f777f0000000007000000;

	lut_sub lut_1201 ({sk[212], x15x, x11x, x483x, x14x, x472x, x565x}, x12626x);
	defparam lut_1201.LUT_SIZE = 7;
	defparam lut_1201.mask = 128'h777f777f777f777f030303ff575757ff;

	lut_sub lut_1205 ({sk[213], x14x, x475x, x556x, x12623x, x12624x, x12626x}, x12629x);
	defparam lut_1205.LUT_SIZE = 7;
	defparam lut_1205.mask = 128'h777f777f777f777f7f7f7f7f7fffffff;

	lut_sub lut_1211 ({sk[214], x17x, x573x, x560x, x12678x, x12677x}, n_n553);
	defparam lut_1211.LUT_SIZE = 6;
	defparam lut_1211.mask = 64'h77ff77ff77777fff;

	lut_sub lut_1216 ({sk[215], x11x, x530x, x38x, x395x, x12680x, x12681x}, n_n554);
	defparam lut_1216.LUT_SIZE = 7;
	defparam lut_1216.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_1222 ({sk[216], x18x, x549x, x369x, x12687x, x12689x}, x12691x);
	defparam lut_1222.LUT_SIZE = 6;
	defparam lut_1222.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_1227 ({sk[217], x21x, x20x, x23x, x599x, x12634x, x12632x}, n_n546);
	defparam lut_1227.LUT_SIZE = 7;
	defparam lut_1227.mask = 128'h777f777f777f777f777f7f7f7f7f7f7f;

	lut_sub lut_1233 ({sk[218], x24x, x114x, x555x, x12638x, x22218x}, n_n547);
	defparam lut_1233.LUT_SIZE = 6;
	defparam lut_1233.mask = 64'h77ff77ffbbffbfff;

	lut_sub lut_1238 ({sk[219], x11x, x568x, x12645x, x12646x, x22300x}, x12649x);
	defparam lut_1238.LUT_SIZE = 6;
	defparam lut_1238.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1243 ({sk[220], x18x, x522x, x12670x, x22302x}, x12672x);
	defparam lut_1243.LUT_SIZE = 5;
	defparam lut_1243.mask = 32'h0fffbbbf;

	lut_sub lut_1247 ({sk[221], x12656x, x12663x, x12655x, x12662x, x22217x}, x12673x);
	defparam lut_1247.LUT_SIZE = 6;
	defparam lut_1247.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_1253 ({sk[222], i_9_, i_1_, i_2_, i_0_}, x13x);
	defparam lut_1253.LUT_SIZE = 5;
	defparam lut_1253.mask = 32'h0fff0004;

	lut_sub lut_1255 ({sk[223], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x573x);
	defparam lut_1255.LUT_SIZE = 7;
	defparam lut_1255.mask = 128'h777f777f777f777f0000000000040000;

	lut_sub lut_1257 ({sk[224], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x517x);
	defparam lut_1257.LUT_SIZE = 7;
	defparam lut_1257.mask = 128'h777f777f777f777f0000000000100000;

	lut_sub lut_1259 ({sk[225], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x585x);
	defparam lut_1259.LUT_SIZE = 7;
	defparam lut_1259.mask = 128'h777f777f777f777f0000010000000000;

	lut_sub lut_1261 ({sk[226], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x476x);
	defparam lut_1261.LUT_SIZE = 7;
	defparam lut_1261.mask = 128'h777f777f777f777f0000000000000400;

	lut_sub lut_1263 ({sk[227], x25x, x13x, x573x, x517x, x585x, x476x}, x12707x);
	defparam lut_1263.LUT_SIZE = 7;
	defparam lut_1263.mask = 128'h777f777f777f777f00003fff55557fff;

	lut_sub lut_1268 ({sk[228], i_9_, i_1_, i_2_, i_0_}, x16x);
	defparam lut_1268.LUT_SIZE = 5;
	defparam lut_1268.mask = 32'h0fff0001;

	lut_sub lut_1270 ({sk[229], i_9_, i_7_, i_8_, i_6_}, x24x);
	defparam lut_1270.LUT_SIZE = 5;
	defparam lut_1270.mask = 32'h0fff0400;

	lut_sub lut_1272 ({sk[230], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x497x);
	defparam lut_1272.LUT_SIZE = 7;
	defparam lut_1272.mask = 128'h777f777f777f777f0000000000000001;

	lut_sub lut_1274 ({sk[231], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x498x);
	defparam lut_1274.LUT_SIZE = 7;
	defparam lut_1274.mask = 128'h777f777f777f777f0000010000000000;

	lut_sub lut_1276 ({sk[232], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x535x);
	defparam lut_1276.LUT_SIZE = 7;
	defparam lut_1276.mask = 128'h777f777f777f777f0000000000000010;

	lut_sub lut_1278 ({sk[233], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x473x);
	defparam lut_1278.LUT_SIZE = 7;
	defparam lut_1278.mask = 128'h777f777f777f777f0000000000000100;

	lut_sub lut_1280 ({sk[234], x16x, x24x, x497x, x498x, x535x, x473x}, x12714x);
	defparam lut_1280.LUT_SIZE = 7;
	defparam lut_1280.mask = 128'h777f777f777f777f00005fff33337fff;

	lut_sub lut_1285 ({sk[235], i_9_, i_7_, i_8_, i_6_}, x22x);
	defparam lut_1285.LUT_SIZE = 5;
	defparam lut_1285.mask = 32'h0fff0200;

	lut_sub lut_1287 ({sk[236], x13397x, x13398x, x13414x, x13415x, x13423x}, n_n3989);
	defparam lut_1287.LUT_SIZE = 6;
	defparam lut_1287.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1293 ({sk[237], n_n4016, x13467x, x13468x, x13480x, x13481x}, n_n3993);
	defparam lut_1293.LUT_SIZE = 6;
	defparam lut_1293.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1299 ({sk[238], n_n2446, x13547x, n_n4279, x13520x, n_n4021, x13516x}, n_n3995);
	defparam lut_1299.LUT_SIZE = 7;
	defparam lut_1299.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1306 ({sk[239], x13438x, x13439x, x13501x, x13502x, x13551x, x13552x}, x13555x);
	defparam lut_1306.LUT_SIZE = 7;
	defparam lut_1306.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1313 ({sk[240], x13166x, x13167x, n_n4009, x13188x, n_n3996}, x13569x);
	defparam lut_1313.LUT_SIZE = 6;
	defparam lut_1313.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1319 ({sk[241], x20x, x534x, x22199x, x22313x}, n_n3923);
	defparam lut_1319.LUT_SIZE = 5;
	defparam lut_1319.mask = 32'h0fffeeef;

	lut_sub lut_1323 ({sk[242], x474x, x18x, x13596x, x13598x, x22314x}, n_n3928);
	defparam lut_1323.LUT_SIZE = 6;
	defparam lut_1323.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1328 ({sk[243], x25x, x15x, x590x, x577x, x13605x, x22198x}, n_n3927);
	defparam lut_1328.LUT_SIZE = 7;
	defparam lut_1328.mask = 128'h777f777f777f777fbbbbbbffbfbfbfff;

	lut_sub lut_1333 ({sk[244], x15x, x555x, x107x, x13609x, x13611x}, x13613x);
	defparam lut_1333.LUT_SIZE = 6;
	defparam lut_1333.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_1338 ({sk[245], x13579x, x13586x, x13577x, x13578x, x13584x, x13585x}, x13614x);
	defparam lut_1338.LUT_SIZE = 7;
	defparam lut_1338.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1345 ({sk[246], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x500x);
	defparam lut_1345.LUT_SIZE = 7;
	defparam lut_1345.mask = 128'h777f777f777f777f0001000000000000;

	lut_sub lut_1347 ({sk[247], i_9_, i_7_, i_8_, i_6_}, x11x);
	defparam lut_1347.LUT_SIZE = 5;
	defparam lut_1347.mask = 32'h0fff4000;

	lut_sub lut_1349 ({sk[248], i_9_, i_7_, i_8_, i_6_}, x23x);
	defparam lut_1349.LUT_SIZE = 5;
	defparam lut_1349.mask = 32'h0fff8000;

	lut_sub lut_1351 ({sk[249], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x499x);
	defparam lut_1351.LUT_SIZE = 7;
	defparam lut_1351.mask = 128'h777f777f777f777f0000000000010000;

	lut_sub lut_1353 ({sk[250], x492x, x16x, x500x, x23x, x520x}, x13622x);
	defparam lut_1353.LUT_SIZE = 6;
	defparam lut_1353.mask = 64'h77ff77ff035703ff;

	lut_sub lut_1357 ({sk[251], x16x, x21x, x510x, x587x, x573x, x498x}, x22197x);
	defparam lut_1357.LUT_SIZE = 7;
	defparam lut_1357.mask = 128'h777f777f777f777fffffaaaac0008000;

	lut_sub lut_1362 ({sk[252], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x529x);
	defparam lut_1362.LUT_SIZE = 7;
	defparam lut_1362.mask = 128'h777f777f777f777f0000000000000800;

	lut_sub lut_1364 ({sk[253], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x575x);
	defparam lut_1364.LUT_SIZE = 7;
	defparam lut_1364.mask = 128'h777f777f777f777f0000000000400000;

	lut_sub lut_1366 ({sk[254], x15x, x483x, x14x, x588x, x478x}, x13642x);
	defparam lut_1366.LUT_SIZE = 6;
	defparam lut_1366.mask = 64'h77ff77ff050537ff;

	lut_sub lut_1370 ({sk[255], x14x, x20x, x502x, x595x, x562x, x493x}, x13643x);
	defparam lut_1370.LUT_SIZE = 7;
	defparam lut_1370.mask = 128'h777f777f777f777f00000f0f77ff7fff;

	lut_sub lut_1375 ({sk[256], x15x, x14x, x529x, x575x, x13642x, x13643x}, x13645x);
	defparam lut_1375.LUT_SIZE = 7;
	defparam lut_1375.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_1380 ({sk[257], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x542x);
	defparam lut_1380.LUT_SIZE = 7;
	defparam lut_1380.mask = 128'h777f777f777f777f0000000000040000;

	lut_sub lut_1382 ({sk[258], x25x, x13x, x587x, x503x, x543x}, x13662x);
	defparam lut_1382.LUT_SIZE = 6;
	defparam lut_1382.mask = 64'h77ff77ff003f557f;

	lut_sub lut_1386 ({sk[259], x13x, x23x, x508x, x518x, x574x, x543x}, x22195x);
	defparam lut_1386.LUT_SIZE = 7;
	defparam lut_1386.mask = 128'h777f777f777f777fffffaaaac0008000;

	lut_sub lut_1391 ({sk[260], x15x, x24x, x542x, x13662x, x22195x}, x13665x);
	defparam lut_1391.LUT_SIZE = 6;
	defparam lut_1391.mask = 64'h77ff77ffbbbfbfbf;

	lut_sub lut_1396 ({sk[261], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x495x);
	defparam lut_1396.LUT_SIZE = 7;
	defparam lut_1396.mask = 128'h777f777f777f777f0000000001000000;

	lut_sub lut_1398 ({sk[262], x25x, x13x, x482x, x475x, x581x, x476x}, x22196x);
	defparam lut_1398.LUT_SIZE = 7;
	defparam lut_1398.mask = 128'h777f777f777f777fffffc000aaaa8000;

	lut_sub lut_1403 ({sk[263], x25x, x16x, x544x, x509x, x24x, x488x}, x22315x);
	defparam lut_1403.LUT_SIZE = 7;
	defparam lut_1403.mask = 128'h777f777f777f777fffcca080ff00a000;

	lut_sub lut_1408 ({sk[264], i_9_, i_7_, i_8_, i_6_}, x20x);
	defparam lut_1408.LUT_SIZE = 5;
	defparam lut_1408.mask = 32'h0fff2000;

	lut_sub lut_1410 ({sk[265], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x550x);
	defparam lut_1410.LUT_SIZE = 7;
	defparam lut_1410.mask = 128'h777f777f777f777f0000000000000001;

	lut_sub lut_1412 ({sk[266], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x563x);
	defparam lut_1412.LUT_SIZE = 7;
	defparam lut_1412.mask = 128'h777f777f777f777f0000000002000000;

	lut_sub lut_1414 ({sk[267], x15x, x16x, x20x, x550x, x497x, x563x}, x13678x);
	defparam lut_1414.LUT_SIZE = 7;
	defparam lut_1414.mask = 128'h777f777f777f777f00335f7f33337f7f;

	lut_sub lut_1419 ({sk[268], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x474x);
	defparam lut_1419.LUT_SIZE = 7;
	defparam lut_1419.mask = 128'h777f777f777f777f0000000000200000;

	lut_sub lut_1421 ({sk[269], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x478x);
	defparam lut_1421.LUT_SIZE = 7;
	defparam lut_1421.mask = 128'h777f777f777f777f0020000000000000;

	lut_sub lut_1423 ({sk[270], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x536x);
	defparam lut_1423.LUT_SIZE = 7;
	defparam lut_1423.mask = 128'h777f777f777f777f0000000000002000;

	lut_sub lut_1425 ({sk[271], x16x, x501x, x20x, x494x}, x124x);
	defparam lut_1425.LUT_SIZE = 5;
	defparam lut_1425.mask = 32'h0fff0357;

	lut_sub lut_1428 ({sk[272], i_9_, i_7_, i_8_, i_6_, x499x, x498x}, x13687x);
	defparam lut_1428.LUT_SIZE = 7;
	defparam lut_1428.mask = 128'h777f777f777f777f0003005000000000;

	lut_sub lut_1431 ({sk[273], x16x, x24x, x499x, x573x, x494x}, x13688x);
	defparam lut_1431.LUT_SIZE = 6;
	defparam lut_1431.mask = 64'h77ff77ff000f777f;

	lut_sub lut_1435 ({sk[274], x22x, x16x, x21x, x501x, x500x, x549x}, x22323x);
	defparam lut_1435.LUT_SIZE = 7;
	defparam lut_1435.mask = 128'h777f777f777f777ffff0aaa0ccc08880;

	lut_sub lut_1444 ({sk[275], x25x, x568x, x578x, x13696x, x13695x}, n_n3196);
	defparam lut_1444.LUT_SIZE = 6;
	defparam lut_1444.mask = 64'h77ff77ff77777fff;

	lut_sub lut_1449 ({sk[276], x19x, x22x, x491x, x579x, x13710x, x13709x}, n_n3194);
	defparam lut_1449.LUT_SIZE = 7;
	defparam lut_1449.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_1454 ({sk[277], x13700x, x13702x, x13713x, x22181x}, x13714x);
	defparam lut_1454.LUT_SIZE = 5;
	defparam lut_1454.mask = 32'h0fffbfff;

	lut_sub lut_1459 ({sk[278], x23x, x513x, x532x, x13718x, x22180x}, n_n3197);
	defparam lut_1459.LUT_SIZE = 6;
	defparam lut_1459.mask = 64'h77ff77ffbbbbbfff;

	lut_sub lut_1464 ({sk[279], x25x, x24x, x590x, x513x, x13725x, x13726x}, x13728x);
	defparam lut_1464.LUT_SIZE = 7;
	defparam lut_1464.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_1469 ({sk[280], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x472x);
	defparam lut_1469.LUT_SIZE = 7;
	defparam lut_1469.mask = 128'h777f777f777f777f0000002000000000;

	lut_sub lut_1471 ({sk[281], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x559x);
	defparam lut_1471.LUT_SIZE = 7;
	defparam lut_1471.mask = 128'h777f777f777f777f0100000000000000;

	lut_sub lut_1473 ({sk[282], i_9_, i_7_, i_8_, i_6_, x496x, x476x}, x13731x);
	defparam lut_1473.LUT_SIZE = 7;
	defparam lut_1473.mask = 128'h777f777f777f777f5030000000000000;

	lut_sub lut_1476 ({sk[283], x25x, x13x, x482x, x495x}, x13732x);
	defparam lut_1476.LUT_SIZE = 5;
	defparam lut_1476.mask = 32'h0fff0357;

	lut_sub lut_1479 ({sk[284], x16x, x13x, x594x, x527x, x593x}, x13734x);
	defparam lut_1479.LUT_SIZE = 6;
	defparam lut_1479.mask = 64'h77ff77ff005f337f;

	lut_sub lut_1483 ({sk[285], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x504x);
	defparam lut_1483.LUT_SIZE = 7;
	defparam lut_1483.mask = 128'h777f777f777f777f0000000004000000;

	lut_sub lut_1485 ({sk[286], x13x, x20x, x489x, x523x}, x471x);
	defparam lut_1485.LUT_SIZE = 5;
	defparam lut_1485.mask = 32'h0fff0537;

	lut_sub lut_1488 ({sk[287], x21x, x13x, x541x, x493x}, x13739x);
	defparam lut_1488.LUT_SIZE = 5;
	defparam lut_1488.mask = 32'h0fff0537;

	lut_sub lut_1491 ({sk[288], x13x, x20x, x503x, x543x, n_n4539, n_n4507}, x22179x);
	defparam lut_1491.LUT_SIZE = 7;
	defparam lut_1491.mask = 128'h777f777f777f777f8888808088008000;

	lut_sub lut_1496 ({sk[289], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x582x);
	defparam lut_1496.LUT_SIZE = 7;
	defparam lut_1496.mask = 128'h777f777f777f777f0010000000000000;

	lut_sub lut_1498 ({sk[290], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x526x);
	defparam lut_1498.LUT_SIZE = 7;
	defparam lut_1498.mask = 128'h777f777f777f777f1000000000000000;

	lut_sub lut_1500 ({sk[291], x25x, x24x, x14x, x550x, x551x}, n_n3125);
	defparam lut_1500.LUT_SIZE = 6;
	defparam lut_1500.mask = 64'h77ff77ff03575757;

	lut_sub lut_1504 ({sk[292], x10x, x24x, x557x, x580x, x537x, x526x}, x13759x);
	defparam lut_1504.LUT_SIZE = 7;
	defparam lut_1504.mask = 128'h777f777f777f777f000055553fff7fff;

	lut_sub lut_1509 ({sk[293], x15x, x23x, x582x, x526x, n_n3125, x13759x}, x13761x);
	defparam lut_1509.LUT_SIZE = 7;
	defparam lut_1509.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_1514 ({sk[294], i_9_, i_1_, i_2_, i_0_}, x17x);
	defparam lut_1514.LUT_SIZE = 5;
	defparam lut_1514.mask = 32'h0fff0002;

	lut_sub lut_1516 ({sk[295], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x584x);
	defparam lut_1516.LUT_SIZE = 7;
	defparam lut_1516.mask = 128'h777f777f777f777f0000040000000000;

	lut_sub lut_1518 ({sk[296], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x576x);
	defparam lut_1518.LUT_SIZE = 7;
	defparam lut_1518.mask = 128'h777f777f777f777f0000000000020000;

	lut_sub lut_1520 ({sk[297], x492x, x22x, x17x, x596x, x537x}, x13779x);
	defparam lut_1520.LUT_SIZE = 6;
	defparam lut_1520.mask = 64'h77ff77ff05370f3f;

	lut_sub lut_1524 ({sk[298], x538x, x11x, x17x, x20x, x475x, x596x}, x13780x);
	defparam lut_1524.LUT_SIZE = 7;
	defparam lut_1524.mask = 128'h777f777f777f777f0537557705ff55ff;

	lut_sub lut_1529 ({sk[299], x24x, x17x, x584x, x576x, x13779x, x13780x}, x13782x);
	defparam lut_1529.LUT_SIZE = 7;
	defparam lut_1529.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_1534 ({sk[300], x21x, x14x, x20x, x565x, x491x}, n_n4210);
	defparam lut_1534.LUT_SIZE = 6;
	defparam lut_1534.mask = 64'h77ff77ff03573377;

	lut_sub lut_1538 ({sk[301], x24x, x14x, x572x, x574x, x560x, x575x}, x14375x);
	defparam lut_1538.LUT_SIZE = 7;
	defparam lut_1538.mask = 128'h777f777f777f777f00003fff55557fff;

	lut_sub lut_1543 ({sk[302], i_9_, i_7_, i_8_, i_6_, n_n325, n_n491}, x14376x);
	defparam lut_1543.LUT_SIZE = 7;
	defparam lut_1543.mask = 128'h777f777f777f777f0101000101000100;

	lut_sub lut_1549 ({sk[303], i_9_, i_7_, i_8_, i_6_, n_n509, n_n325}, n_n3707);
	defparam lut_1549.LUT_SIZE = 7;
	defparam lut_1549.mask = 128'h777f777f777f777f0100101011110101;

	lut_sub lut_1559 ({sk[304], i_9_, i_7_, i_8_, i_6_, x483x, x565x}, x14383x);
	defparam lut_1559.LUT_SIZE = 7;
	defparam lut_1559.mask = 128'h777f777f777f777f3000000500000000;

	lut_sub lut_1562 ({sk[305], i_9_, i_7_, i_8_, i_6_, n_n325, n_n500}, x14384x);
	defparam lut_1562.LUT_SIZE = 7;
	defparam lut_1562.mask = 128'h777f777f777f777f0101000001001000;

	lut_sub lut_1567 ({sk[306], n_n4210, x14375x, x14376x, n_n3707, x14383x, x14384x}, x14388x);
	defparam lut_1567.LUT_SIZE = 7;
	defparam lut_1567.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1574 ({sk[307], x22x, x543x, x189x, n_n3875, x22165x}, x14458x);
	defparam lut_1574.LUT_SIZE = 6;
	defparam lut_1574.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1579 ({sk[308], x130x, n_n3879, x14446x, x14447x, x14453x, x14454x}, x14459x);
	defparam lut_1579.LUT_SIZE = 7;
	defparam lut_1579.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1586 ({sk[309], x20x, x496x, x14529x, x22303x}, x14530x);
	defparam lut_1586.LUT_SIZE = 5;
	defparam lut_1586.mask = 32'h0fffbbbf;

	lut_sub lut_1590 ({sk[310], x15x, x544x, n_n3889, n_n4458, x14515x, x14516x}, n_n3729);
	defparam lut_1590.LUT_SIZE = 7;
	defparam lut_1590.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_1596 ({sk[311], x22x, x11x, x496x, x215x, x14522x}, n_n3731);
	defparam lut_1596.LUT_SIZE = 6;
	defparam lut_1596.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_1601 ({sk[312], n_n3727, n_n3726, x14534x, x22164x}, x14538x);
	defparam lut_1601.LUT_SIZE = 5;
	defparam lut_1601.mask = 32'h0fffbfff;

	lut_sub lut_1606 ({sk[313], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x525x);
	defparam lut_1606.LUT_SIZE = 7;
	defparam lut_1606.mask = 128'h777f777f777f777f8000000000000000;

	lut_sub lut_1608 ({sk[314], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x489x);
	defparam lut_1608.LUT_SIZE = 7;
	defparam lut_1608.mask = 128'h777f777f777f777f0000800000000000;

	lut_sub lut_1610 ({sk[315], i_9_, i_1_, i_2_, i_0_, x525x, x489x}, x149x);
	defparam lut_1610.LUT_SIZE = 7;
	defparam lut_1610.mask = 128'h777f777f777f777f0000000070000000;

	lut_sub lut_1613 ({sk[316], n_n3661, x14560x, x14564x, x14565x, x22156x}, n_n3632);
	defparam lut_1613.LUT_SIZE = 6;
	defparam lut_1613.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_1619 ({sk[317], x24x, x599x, x318x, n_n761, x22155x}, x14582x);
	defparam lut_1619.LUT_SIZE = 6;
	defparam lut_1619.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1624 ({sk[318], x383x, x14572x, x14571x, x14578x, x22154x}, x14583x);
	defparam lut_1624.LUT_SIZE = 6;
	defparam lut_1624.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_1630 ({sk[319], x592x, x24x, x14584x, x14586x, x22321x}, x14589x);
	defparam lut_1630.LUT_SIZE = 6;
	defparam lut_1630.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1635 ({sk[320], x19x, x560x, x217x, x14545x, n_n3665, x14543x}, x14590x);
	defparam lut_1635.LUT_SIZE = 7;
	defparam lut_1635.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_1641 ({sk[321], x12x, x574x, x76x, x126x, x22325x}, n_n3674);
	defparam lut_1641.LUT_SIZE = 6;
	defparam lut_1641.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1646 ({sk[322], x24x, x591x, x14598x, x22301x}, n_n3673);
	defparam lut_1646.LUT_SIZE = 5;
	defparam lut_1646.mask = 32'h0fffbbbf;

	lut_sub lut_1650 ({sk[323], n_n3412, n_n3051, n_n3676, x14608x, x14609x, x14611x}, n_n3637);
	defparam lut_1650.LUT_SIZE = 7;
	defparam lut_1650.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1657 ({sk[324], n_n3670, x14624x, x14625x, x14626x, x14627x}, n_n3635);
	defparam lut_1657.LUT_SIZE = 6;
	defparam lut_1657.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1663 ({sk[325], x12x, x114x, x520x, x14632x, x14634x}, x14636x);
	defparam lut_1663.LUT_SIZE = 6;
	defparam lut_1663.mask = 64'h77ff77ff77ff7fff;

	lut_sub lut_1668 ({sk[326], x24x, x554x, x123x, x14642x, x22162x}, n_n3679);
	defparam lut_1668.LUT_SIZE = 6;
	defparam lut_1668.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1673 ({sk[327], x11x, x598x, x34x, x122x, x232x, x14646x}, n_n3678);
	defparam lut_1673.LUT_SIZE = 7;
	defparam lut_1673.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_1679 ({sk[328], x18x, x488x, x524x, n_n4152, x22309x}, x14654x);
	defparam lut_1679.LUT_SIZE = 6;
	defparam lut_1679.mask = 64'h77ff77ffbbbbbfff;

	lut_sub lut_1684 ({sk[329], n_n4161, x14659x, x14661x, x253x, x14657x, x14658x}, x14668x);
	defparam lut_1684.LUT_SIZE = 7;
	defparam lut_1684.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1691 ({sk[330], n_n3685, n_n3686, x14665x, x14666x, x14680x, x22163x}, x22339x);
	defparam lut_1691.LUT_SIZE = 7;
	defparam lut_1691.mask = 128'h777f777f777f777f4000000000000000;

	lut_sub lut_1693 ({sk[331], x15x, x24x, x17x, x484x, x480x}, n_n2727);
	defparam lut_1693.LUT_SIZE = 6;
	defparam lut_1693.mask = 64'h77ff77ff05373737;

	lut_sub lut_1697 ({sk[332], i_9_, n_n534, x474x, n_n260, x472x, n_n500}, x14689x);
	defparam lut_1697.LUT_SIZE = 7;
	defparam lut_1697.mask = 128'h777f777f777f777f00000505030f070f;

	lut_sub lut_1702 ({sk[333], i_9_, i_7_, i_8_, i_6_, n_n509, n_n260}, x14690x);
	defparam lut_1702.LUT_SIZE = 7;
	defparam lut_1702.mask = 128'h777f777f777f777f1100101001000000;

	lut_sub lut_1708 ({sk[334], i_9_, i_7_, i_8_, i_6_, n_n518, n_n260}, n_n3698);
	defparam lut_1708.LUT_SIZE = 7;
	defparam lut_1708.mask = 128'h777f777f777f777f0101110001011110;

	lut_sub lut_1718 ({sk[335], x17x, x20x, x481x, x596x}, x14725x);
	defparam lut_1718.LUT_SIZE = 5;
	defparam lut_1718.mask = 32'h0fff0537;

	lut_sub lut_1721 ({sk[336], i_9_, n_n518, n_n534, n_n509, n_n260, n_n520}, x14726x);
	defparam lut_1721.LUT_SIZE = 7;
	defparam lut_1721.mask = 128'h777f777f777f777f0003111300031113;

	lut_sub lut_1726 ({sk[337], n_n2727, x14689x, x14690x, n_n3698, x14725x, x14726x}, x14730x);
	defparam lut_1726.LUT_SIZE = 7;
	defparam lut_1726.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1733 ({sk[338], x17x, x549x, x389x, x14706x, x22161x}, x14710x);
	defparam lut_1733.LUT_SIZE = 6;
	defparam lut_1733.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1738 ({sk[339], x14x, x529x, x395x, x14697x, x22160x, x22254x}, x14711x);
	defparam lut_1738.LUT_SIZE = 7;
	defparam lut_1738.mask = 128'h777f777f777f777fefffefffefffffff;

	lut_sub lut_1744 ({sk[340], x11x, x14x, x588x, x520x, n_n4204, x447x}, x14722x);
	defparam lut_1744.LUT_SIZE = 7;
	defparam lut_1744.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_1749 ({sk[341], x11x, x511x, x179x, x14714x, x14712x, x14721x}, x14723x);
	defparam lut_1749.LUT_SIZE = 7;
	defparam lut_1749.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_1755 ({sk[342], x105x, x42x, x142x, n_n3691, x14746x, x14748x}, n_n3642);
	defparam lut_1755.LUT_SIZE = 7;
	defparam lut_1755.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1762 ({sk[343], n_n4172, x13836x, x14762x}, x14764x);
	defparam lut_1762.LUT_SIZE = 4;
	defparam lut_1762.mask = 16'h5f7f;

	lut_sub lut_1766 ({sk[344], n_n3803, n_n3802, x14754x, x14757x, x22151x}, x14765x);
	defparam lut_1766.LUT_SIZE = 6;
	defparam lut_1766.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_1772 ({sk[345], i_9_, i_7_, i_8_, i_6_, n_n260, n_n500}, x14770x);
	defparam lut_1772.LUT_SIZE = 7;
	defparam lut_1772.mask = 128'h777f777f777f777f0001011001111110;

	lut_sub lut_1782 ({sk[346], n_n3810, n_n2718, x14733x, x14738x, x14732x, x14737x}, x14771x);
	defparam lut_1782.LUT_SIZE = 7;
	defparam lut_1782.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1789 ({sk[347], n_n3642, x14764x, x14765x, x14770x, x14771x}, n_n3626);
	defparam lut_1789.LUT_SIZE = 6;
	defparam lut_1789.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1795 ({sk[348], x21x, x18x, x573x, x513x, x14793x, x14794x}, x14796x);
	defparam lut_1795.LUT_SIZE = 7;
	defparam lut_1795.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_1800 ({sk[349], x14807x, x14801x, x14802x, x22135x}, n_n2451);
	defparam lut_1800.LUT_SIZE = 5;
	defparam lut_1800.mask = 32'h0fffbfff;

	lut_sub lut_1805 ({sk[350], x539x, x12x, x34x, x155x, x143x, x14782x}, n_n2460);
	defparam lut_1805.LUT_SIZE = 7;
	defparam lut_1805.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_1811 ({sk[351], x12x, x572x, x520x, n_n5234, x385x, x14790x}, n_n2459);
	defparam lut_1811.LUT_SIZE = 7;
	defparam lut_1811.mask = 128'h777f777f777f777f7f7f7f7f7fffffff;

	lut_sub lut_1817 ({sk[352], x17x, x506x, x31x, x353x, x22134x}, x14827x);
	defparam lut_1817.LUT_SIZE = 6;
	defparam lut_1817.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1822 ({sk[353], x14813x, x14820x, x14811x, x14812x, x14818x, x14819x}, x14828x);
	defparam lut_1822.LUT_SIZE = 7;
	defparam lut_1822.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1829 ({sk[354], x14796x, n_n2451, n_n2460, n_n2459, x14827x, x14828x}, n_n2449);
	defparam lut_1829.LUT_SIZE = 7;
	defparam lut_1829.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1836 ({sk[355], x17x, x20x, x23x, x566x, x574x}, n_n3450);
	defparam lut_1836.LUT_SIZE = 6;
	defparam lut_1836.mask = 64'h77ff77ff03335777;

	lut_sub lut_1840 ({sk[356], i_9_, i_7_, i_8_, i_6_, n_n260, n_n500}, n_n2598);
	defparam lut_1840.LUT_SIZE = 7;
	defparam lut_1840.mask = 128'h777f777f777f777f0100110100111110;

	lut_sub lut_1850 ({sk[357], x15x, x17x, x557x, x572x, x576x}, x14912x);
	defparam lut_1850.LUT_SIZE = 6;
	defparam lut_1850.mask = 64'h77ff77ff003f557f;

	lut_sub lut_1854 ({sk[358], x25x, x24x, x17x, x573x, x576x}, x48x);
	defparam lut_1854.LUT_SIZE = 6;
	defparam lut_1854.mask = 64'h77ff77ff03575757;

	lut_sub lut_1858 ({sk[359], x21x, x17x, x484x, x477x, x478x, x564x}, x14931x);
	defparam lut_1858.LUT_SIZE = 7;
	defparam lut_1858.mask = 128'h777f777f777f777f00007f7f00ff7fff;

	lut_sub lut_1863 ({sk[360], i_9_, i_7_, i_8_, i_6_, n_n509, n_n260}, x14932x);
	defparam lut_1863.LUT_SIZE = 7;
	defparam lut_1863.mask = 128'h777f777f777f777f0101010000011000;

	lut_sub lut_1869 ({sk[361], n_n3450, n_n2598, x14912x, x48x, x14931x, x14932x}, x14935x);
	defparam lut_1869.LUT_SIZE = 7;
	defparam lut_1869.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1876 ({sk[362], x14918x, x14922x, x14923x, x22147x}, x14928x);
	defparam lut_1876.LUT_SIZE = 5;
	defparam lut_1876.mask = 32'h0fffbfff;

	lut_sub lut_1881 ({sk[363], x25x, x552x, x20x, x596x, n_n3461, x14894x}, n_n2601);
	defparam lut_1881.LUT_SIZE = 7;
	defparam lut_1881.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_1886 ({sk[364], x14x, x516x, x38x, x389x, x22146x}, n_n2602);
	defparam lut_1886.LUT_SIZE = 6;
	defparam lut_1886.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1891 ({sk[365], x14904x, x14905x, x14924x, x14925x}, x22145x);
	defparam lut_1891.LUT_SIZE = 5;
	defparam lut_1891.mask = 32'h0fff8000;

	lut_sub lut_1893 ({sk[366], i_9_, i_7_, i_8_, i_6_, n_n482, n_n260}, x14960x);
	defparam lut_1893.LUT_SIZE = 7;
	defparam lut_1893.mask = 128'h777f777f777f777f0111100011101010;

	lut_sub lut_1903 ({sk[367], x14948x, x14954x, x14952x, x14953x, x22144x}, x14961x);
	defparam lut_1903.LUT_SIZE = 6;
	defparam lut_1903.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_1909 ({sk[368], x23x, x512x, x14972x, x22269x}, x14974x);
	defparam lut_1909.LUT_SIZE = 5;
	defparam lut_1909.mask = 32'h0fffbbbf;

	lut_sub lut_1913 ({sk[369], x24x, x531x, x382x, n_n2591, x22143x}, x14975x);
	defparam lut_1913.LUT_SIZE = 6;
	defparam lut_1913.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1918 ({sk[370], x521x, x18x, x20x, x553x, x29x, x14977x}, x14979x);
	defparam lut_1918.LUT_SIZE = 7;
	defparam lut_1918.mask = 128'h777f777f777f777f777f777f777fffff;

	lut_sub lut_1923 ({sk[371], x14938x, x14939x, x247x, x393x, x14943x}, x14980x);
	defparam lut_1923.LUT_SIZE = 6;
	defparam lut_1923.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1929 ({sk[372], x10x, x528x, x426x, x14997x, x14998x, x14999x}, x15005x);
	defparam lut_1929.LUT_SIZE = 7;
	defparam lut_1929.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_1935 ({sk[373], x219x, n_n2614, x417x, x445x, x442x}, x15006x);
	defparam lut_1935.LUT_SIZE = 6;
	defparam lut_1935.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1941 ({sk[374], x243x, n_n856, n_n2611, x15011x, x15012x, x15013x}, n_n2551);
	defparam lut_1941.LUT_SIZE = 7;
	defparam lut_1941.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_1948 ({sk[375], x14x, x586x, x20x, x575x, x15020x, x15021x}, x15023x);
	defparam lut_1948.LUT_SIZE = 7;
	defparam lut_1948.mask = 128'h777f777f777f777f777f777f777fffff;

	lut_sub lut_1953 ({sk[376], x14985x, x14991x, x350x, x14984x, x22133x}, x15024x);
	defparam lut_1953.LUT_SIZE = 6;
	defparam lut_1953.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_1959 ({sk[377], x15005x, x15006x, n_n2551, x15023x, x15024x}, n_n2531);
	defparam lut_1959.LUT_SIZE = 6;
	defparam lut_1959.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1965 ({sk[378], x16x, x573x, x560x, x537x, x423x, x22142x}, n_n2637);
	defparam lut_1965.LUT_SIZE = 7;
	defparam lut_1965.mask = 128'h777f777f777f777fbbbbbbbbbfffffff;

	lut_sub lut_1971 ({sk[379], x24x, x498x, x161x, x15032x, x22281x}, n_n2638);
	defparam lut_1971.LUT_SIZE = 6;
	defparam lut_1971.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_1976 ({sk[380], n_n2634, x15049x, x15055x, x15047x, x15048x}, n_n2559);
	defparam lut_1976.LUT_SIZE = 6;
	defparam lut_1976.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_1982 ({sk[381], i_9_, i_7_, i_8_, i_6_, n_n536, n_n491}, x15038x);
	defparam lut_1982.LUT_SIZE = 7;
	defparam lut_1982.mask = 128'h777f777f777f777f0010101000001000;

	lut_sub lut_1987 ({sk[382], i_9_, n_n536, n_n482, n_n532, n_n534, n_n4388}, x15039x);
	defparam lut_1987.LUT_SIZE = 7;
	defparam lut_1987.mask = 128'h777f777f777f777f5555557f5555557f;

	lut_sub lut_1993 ({sk[383], x156x, n_n2640, n_n2641, x337x, x15161x, x15162x}, x15167x);
	defparam lut_1993.LUT_SIZE = 7;
	defparam lut_1993.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_2000 ({sk[384], x19x, x545x, x15219x, x22327x}, x15221x);
	defparam lut_2000.LUT_SIZE = 5;
	defparam lut_2000.mask = 32'h0fffbbbf;

	lut_sub lut_2004 ({sk[385], n_n2570, x220x, x223x, x15217x}, x15222x);
	defparam lut_2004.LUT_SIZE = 5;
	defparam lut_2004.mask = 32'h0fff7fff;

	lut_sub lut_2009 ({sk[386], x510x, x12x, x22256x, x22274x}, x15278x);
	defparam lut_2009.LUT_SIZE = 5;
	defparam lut_2009.mask = 32'h0fffeeef;

	lut_sub lut_2013 ({sk[387], x15269x, x152x, x15268x, x15273x, x22138x}, x15279x);
	defparam lut_2013.LUT_SIZE = 6;
	defparam lut_2013.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2019 ({sk[388], x15283x, x15287x, x15288x, x15281x, x15282x, x15293x}, x15295x);
	defparam lut_2019.LUT_SIZE = 7;
	defparam lut_2019.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_2026 ({sk[389], x16x, x21x, x11x, x529x, x498x, x496x}, x15307x);
	defparam lut_2026.LUT_SIZE = 7;
	defparam lut_2026.mask = 128'h777f777f777f777f005533770f5f3f7f;

	lut_sub lut_2030 ({sk[390], x15x, x500x, x23x, x499x, x473x, n_n4384}, x22110x);
	defparam lut_2030.LUT_SIZE = 7;
	defparam lut_2030.mask = 128'h777f777f777f777faa80aa80aa800000;

	lut_sub lut_2035 ({sk[391], x22x, x16x, x489x, x495x, x15307x, x22110x}, n_n2845);
	defparam lut_2035.LUT_SIZE = 7;
	defparam lut_2035.mask = 128'h777f777f777f777fbbbbbbffbfbfbfff;

	lut_sub lut_2040 ({sk[392], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x477x);
	defparam lut_2040.LUT_SIZE = 7;
	defparam lut_2040.mask = 128'h777f777f777f777f0002000000000000;

	lut_sub lut_2042 ({sk[393], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x594x);
	defparam lut_2042.LUT_SIZE = 7;
	defparam lut_2042.mask = 128'h777f777f777f777f0000000000000100;

	lut_sub lut_2044 ({sk[394], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x593x);
	defparam lut_2044.LUT_SIZE = 7;
	defparam lut_2044.mask = 128'h777f777f777f777f0000000001000000;

	lut_sub lut_2046 ({sk[395], x13x, x477x, x23x, x594x, x476x, x593x}, x15315x);
	defparam lut_2046.LUT_SIZE = 7;
	defparam lut_2046.mask = 128'h777f777f777f777f003300335f7fffff;

	lut_sub lut_2051 ({sk[396], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x544x);
	defparam lut_2051.LUT_SIZE = 7;
	defparam lut_2051.mask = 128'h777f777f777f777f0000000400000000;

	lut_sub lut_2053 ({sk[397], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x564x);
	defparam lut_2053.LUT_SIZE = 7;
	defparam lut_2053.mask = 128'h777f777f777f777f0000000000000200;

	lut_sub lut_2055 ({sk[398], x21x, x13x, x20x, x540x, x480x}, x15314x);
	defparam lut_2055.LUT_SIZE = 6;
	defparam lut_2055.mask = 64'h77ff77ff03573377;

	lut_sub lut_2059 ({sk[399], x25x, x15315x, x13x, x544x, x564x, x15314x}, n_n2844);
	defparam lut_2059.LUT_SIZE = 7;
	defparam lut_2059.mask = 128'h777f777f777f777f5577ffff5f7fffff;

	lut_sub lut_2064 ({sk[400], i_9_, i_7_, i_8_, i_6_, x501x, x473x}, x15320x);
	defparam lut_2064.LUT_SIZE = 7;
	defparam lut_2064.mask = 128'h777f777f777f777f0300500000000000;

	lut_sub lut_2067 ({sk[401], x25x, x16x, x11x, x497x, x548x, x473x}, x15321x);
	defparam lut_2067.LUT_SIZE = 7;
	defparam lut_2067.mask = 128'h777f777f777f777f000f333f555f777f;

	lut_sub lut_2071 ({sk[402], x16x, x24x, x497x, x480x, x535x}, x22282x);
	defparam lut_2071.LUT_SIZE = 6;
	defparam lut_2071.mask = 64'h77ff77fffff08880;

	lut_sub lut_2076 ({sk[403], x20x, x473x, x15320x, x15321x, x22282x}, n_n2846);
	defparam lut_2076.LUT_SIZE = 6;
	defparam lut_2076.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_2081 ({sk[404], x13x, x11x, x505x, x504x}, x416x);
	defparam lut_2081.LUT_SIZE = 5;
	defparam lut_2081.mask = 32'h0fff0537;

	lut_sub lut_2084 ({sk[405], x15x, x538x, x13x, x543x}, x15337x);
	defparam lut_2084.LUT_SIZE = 5;
	defparam lut_2084.mask = 32'h0fff0357;

	lut_sub lut_2087 ({sk[406], x13x, x11x, x519x, x580x, x542x, x543x}, x22109x);
	defparam lut_2087.LUT_SIZE = 7;
	defparam lut_2087.mask = 128'h777f777f777f777fffff8888f0008000;

	lut_sub lut_2092 ({sk[407], x13x, x529x, x416x, x15337x, x22109x}, x15342x);
	defparam lut_2092.LUT_SIZE = 6;
	defparam lut_2092.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_2097 ({sk[408], x12x, x550x, x279x, x15365x, x22115x}, x15369x);
	defparam lut_2097.LUT_SIZE = 6;
	defparam lut_2097.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_2102 ({sk[409], x11x, x24x, x568x, x578x, x15354x, x22114x}, n_n2832);
	defparam lut_2102.LUT_SIZE = 7;
	defparam lut_2102.mask = 128'h777f777f777f777fbbbbbfbfbbffbfff;

	lut_sub lut_2107 ({sk[410], x25x, x120x, x567x, x15357x, x15358x, x15359x}, n_n2834);
	defparam lut_2107.LUT_SIZE = 7;
	defparam lut_2107.mask = 128'h777f777f777f777f7f7fffff7fffffff;

	lut_sub lut_2113 ({sk[411], x15348x, x15390x, x15347x, x15389x, x22113x}, x15399x);
	defparam lut_2113.LUT_SIZE = 6;
	defparam lut_2113.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2119 ({sk[412], x15369x, n_n2832, n_n2834, x15399x}, x15401x);
	defparam lut_2119.LUT_SIZE = 5;
	defparam lut_2119.mask = 32'h0fff7fff;

	lut_sub lut_2124 ({sk[413], x24x, x483x, x14x, x480x}, x73x);
	defparam lut_2124.LUT_SIZE = 5;
	defparam lut_2124.mask = 32'h0fff111f;

	lut_sub lut_2127 ({sk[414], x15x, x483x, x14x, x474x, x475x}, n_n1760);
	defparam lut_2127.LUT_SIZE = 6;
	defparam lut_2127.mask = 64'h77ff77ff070707ff;

	lut_sub lut_2131 ({sk[415], i_9_, i_7_, i_8_, i_6_, x483x, x551x}, x15414x);
	defparam lut_2131.LUT_SIZE = 7;
	defparam lut_2131.mask = 128'h777f777f777f777f5000000300000000;

	lut_sub lut_2134 ({sk[416], x14x, x548x, x559x, x73x, n_n1760, x15414x}, x15418x);
	defparam lut_2134.LUT_SIZE = 7;
	defparam lut_2134.mask = 128'h777f777f777f777f7f7f7f7f7fffffff;

	lut_sub lut_2140 ({sk[417], x13x, x563x, x189x, n_n3509, x162x, x15433x}, x15437x);
	defparam lut_2140.LUT_SIZE = 7;
	defparam lut_2140.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_2146 ({sk[418], x22x, x476x, x184x, n_n2999, x11511x, x11510x}, x15438x);
	defparam lut_2146.LUT_SIZE = 7;
	defparam lut_2146.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_2152 ({sk[419], i_9_, i_7_, i_8_, i_6_, n_n455, n_n473}, x15453x);
	defparam lut_2152.LUT_SIZE = 7;
	defparam lut_2152.mask = 128'h777f777f777f777f0011101010011110;

	lut_sub lut_2162 ({sk[420], n_n3152, x15440x, x15445x, x15439x, x15443x, x15444x}, x15454x);
	defparam lut_2162.LUT_SIZE = 7;
	defparam lut_2162.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_2169 ({sk[421], x13x, x546x, x559x, n_n4465, x291x, x22112x}, x15461x);
	defparam lut_2169.LUT_SIZE = 7;
	defparam lut_2169.mask = 128'h777f777f777f777fbfbfbfbfbfffffff;

	lut_sub lut_2175 ({sk[422], n_n3162, n_n3003, x15422x, x22111x}, x15462x);
	defparam lut_2175.LUT_SIZE = 5;
	defparam lut_2175.mask = 32'h0fffbfff;

	lut_sub lut_2180 ({sk[423], x15437x, x15438x, x15453x, x15454x, x15461x, x15462x}, n_n2907);
	defparam lut_2180.LUT_SIZE = 7;
	defparam lut_2180.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_2187 ({sk[424], x10x, x562x, n_n4232, x272x, x22326x}, n_n2990);
	defparam lut_2187.LUT_SIZE = 6;
	defparam lut_2187.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_2192 ({sk[425], x521x, x10x, x559x, x15487x, x22120x}, n_n2991);
	defparam lut_2192.LUT_SIZE = 6;
	defparam lut_2192.mask = 64'h77ff77ffbbbfbbff;

	lut_sub lut_2197 ({sk[426], x492x, x10x, x520x, n_n3132, x11856x, x11857x}, x15471x);
	defparam lut_2197.LUT_SIZE = 7;
	defparam lut_2197.mask = 128'h777f777f777f777f7f7f7fff7f7fffff;

	lut_sub lut_2203 ({sk[427], x21x, x20x, x571x, n_n2987, x157x, x15468x}, x15472x);
	defparam lut_2203.LUT_SIZE = 7;
	defparam lut_2203.mask = 128'h777f777f777f777f7f7f7fff7fff7fff;

	lut_sub lut_2209 ({sk[428], x15x, x10x, x561x, x574x, n_n1646, x15492x}, x15494x);
	defparam lut_2209.LUT_SIZE = 7;
	defparam lut_2209.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_2214 ({sk[429], n_n2990, n_n2991, x15471x, x15472x, x15494x}, x15504x);
	defparam lut_2214.LUT_SIZE = 6;
	defparam lut_2214.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2220 ({sk[430], x15517x, x15518x, x15521x, x15522x, x15527x}, n_n2934);
	defparam lut_2220.LUT_SIZE = 6;
	defparam lut_2220.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2226 ({sk[431], x427x, n_n3004, n_n3005, x15540x, x22119x}, n_n2932);
	defparam lut_2226.LUT_SIZE = 6;
	defparam lut_2226.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2232 ({sk[432], x22x, x16x, x20x, x498x, x560x, x15546x}, x15547x);
	defparam lut_2232.LUT_SIZE = 7;
	defparam lut_2232.mask = 128'h777f777f777f777f555f777f5f5f7f7f;

	lut_sub lut_2237 ({sk[433], x15507x, x15512x, x15506x, x15511x, x22118x}, x15548x);
	defparam lut_2237.LUT_SIZE = 6;
	defparam lut_2237.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2243 ({sk[434], n_n2934, n_n2932, x15547x, x15548x}, n_n2908);
	defparam lut_2243.LUT_SIZE = 5;
	defparam lut_2243.mask = 32'h0fff7fff;

	lut_sub lut_2248 ({sk[435], n_n2948, n_n2949, x15592x}, x15594x);
	defparam lut_2248.LUT_SIZE = 4;
	defparam lut_2248.mask = 16'h5f7f;

	lut_sub lut_2252 ({sk[436], n_n2945, x15564x, x15579x, x22127x}, x15595x);
	defparam lut_2252.LUT_SIZE = 5;
	defparam lut_2252.mask = 32'h0fffbfff;

	lut_sub lut_2257 ({sk[437], n_n2957, x15602x, x15600x, x15601x, x15640x}, x15642x);
	defparam lut_2257.LUT_SIZE = 6;
	defparam lut_2257.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2263 ({sk[438], n_n2953, n_n2955, x15618x, x15633x, x15634x}, x15643x);
	defparam lut_2263.LUT_SIZE = 6;
	defparam lut_2263.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2269 ({sk[439], n_n3019, x15663x, x15667x, x15666x, x22126x}, x15674x);
	defparam lut_2269.LUT_SIZE = 6;
	defparam lut_2269.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2275 ({sk[440], n_n2939, n_n2940, x15647x, x15648x, x22125x}, x15675x);
	defparam lut_2275.LUT_SIZE = 6;
	defparam lut_2275.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2281 ({sk[441], x17x, x546x, n_n3460, x177x, x15693x}, x15696x);
	defparam lut_2281.LUT_SIZE = 6;
	defparam lut_2281.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_2286 ({sk[442], n_n3461, x15686x, x15685x, x15691x, x15692x}, x15697x);
	defparam lut_2286.LUT_SIZE = 6;
	defparam lut_2286.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2292 ({sk[443], x14x, x20x, x506x, x511x, n_n4197, x390x}, x15798x);
	defparam lut_2292.LUT_SIZE = 7;
	defparam lut_2292.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_2297 ({sk[444], x15790x, x15794x, x15795x, x22124x}, x15799x);
	defparam lut_2297.LUT_SIZE = 5;
	defparam lut_2297.mask = 32'h0fffbfff;

	lut_sub lut_2302 ({sk[445], n_n3450, n_n2970, n_n2968, x15801x, x15802x}, x15806x);
	defparam lut_2302.LUT_SIZE = 6;
	defparam lut_2302.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2308 ({sk[446], x15696x, x15697x, x15798x, x15799x, x15806x}, x15808x);
	defparam lut_2308.LUT_SIZE = 6;
	defparam lut_2308.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2314 ({sk[447], x137x, x15714x, x15715x, n_n2962, x15726x, x15727x}, x15743x);
	defparam lut_2314.LUT_SIZE = 7;
	defparam lut_2314.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_2321 ({sk[448], x15766x, x15767x, x15778x, x15779x, x15784x, x15785x}, n_n2905);
	defparam lut_2321.LUT_SIZE = 7;
	defparam lut_2321.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_2328 ({sk[449], i_9_, i_7_, i_8_, i_6_, n_n482, n_n260}, x15740x);
	defparam lut_2328.LUT_SIZE = 7;
	defparam lut_2328.mask = 128'h777f777f777f777f0001001111111010;

	lut_sub lut_2338 ({sk[450], x132x, x105x, x15701x, x15733x, x22121x}, x15741x);
	defparam lut_2338.LUT_SIZE = 6;
	defparam lut_2338.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2344 ({sk[451], x18x, x505x, x488x, x15954x, x22308x}, x15957x);
	defparam lut_2344.LUT_SIZE = 6;
	defparam lut_2344.mask = 64'h77ff77ffbbbbbfff;

	lut_sub lut_2349 ({sk[452], x123x, n_n1952, x209x, x15950x, x15951x, x15944x}, x15958x);
	defparam lut_2349.LUT_SIZE = 7;
	defparam lut_2349.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_2356 ({sk[453], i_9_, i_7_, i_8_, i_6_, n_n130, n_n500}, x15973x);
	defparam lut_2356.LUT_SIZE = 7;
	defparam lut_2356.mask = 128'h777f777f777f777f0100101101110110;

	lut_sub lut_2366 ({sk[454], x15962x, x15967x, x15961x, x15966x, x22092x}, x15974x);
	defparam lut_2366.LUT_SIZE = 6;
	defparam lut_2366.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2372 ({sk[455], x18x, x587x, x111x, x15986x, x22279x}, x15989x);
	defparam lut_2372.LUT_SIZE = 6;
	defparam lut_2372.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_2377 ({sk[456], x15978x, x15982x, x15976x, x15981x, x22091x}, x15990x);
	defparam lut_2377.LUT_SIZE = 6;
	defparam lut_2377.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2383 ({sk[457], x15957x, x15958x, x15973x, x15974x, x15989x, x15990x}, n_n1788);
	defparam lut_2383.LUT_SIZE = 7;
	defparam lut_2383.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_2390 ({sk[458], i_9_, i_7_, i_8_, i_6_, n_n455, n_n500}, n_n1885);
	defparam lut_2390.LUT_SIZE = 7;
	defparam lut_2390.mask = 128'h777f777f777f777f0101100100011111;

	lut_sub lut_2400 ({sk[459], i_9_, i_7_, i_8_, i_6_, n_n455, n_n509}, n_n1886);
	defparam lut_2400.LUT_SIZE = 7;
	defparam lut_2400.mask = 128'h777f777f777f777f1101110000111010;

	lut_sub lut_2410 ({sk[460], x13x, x519x, x23x, x574x, x537x, x541x}, x16023x);
	defparam lut_2410.LUT_SIZE = 7;
	defparam lut_2410.mask = 128'h777f777f777f777f005500553f7fffff;

	lut_sub lut_2415 ({sk[461], x492x, x13x, x572x, x491x, x189x}, x22105x);
	defparam lut_2415.LUT_SIZE = 6;
	defparam lut_2415.mask = 64'h77ff77ffaa80aa00;

	lut_sub lut_2418 ({sk[462], n_n1885, n_n1886, x16023x, x22105x}, x16027x);
	defparam lut_2418.LUT_SIZE = 5;
	defparam lut_2418.mask = 32'h0fffbfff;

	lut_sub lut_2423 ({sk[463], x13x, x550x, x548x, n_n3889, x22104x, x22337x}, x16008x);
	defparam lut_2423.LUT_SIZE = 7;
	defparam lut_2423.mask = 128'h777f777f777f777fefefefefefffffff;

	lut_sub lut_2429 ({sk[464], x25x, x13x, x558x, x543x, n_n3504, x202x}, x16018x);
	defparam lut_2429.LUT_SIZE = 7;
	defparam lut_2429.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_2434 ({sk[465], n_n4243, x307x, x16011x, x16014x, x22103x}, x16019x);
	defparam lut_2434.LUT_SIZE = 6;
	defparam lut_2434.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2440 ({sk[466], i_9_, n_n524, n_n526, n_n455, n_n535, n_n1285}, x16004x);
	defparam lut_2440.LUT_SIZE = 7;
	defparam lut_2440.mask = 128'h777f777f777f777f5557555755575757;

	lut_sub lut_2445 ({sk[467], i_9_, i_7_, i_8_, i_6_, n_n518, n_n455}, x16005x);
	defparam lut_2445.LUT_SIZE = 7;
	defparam lut_2445.mask = 128'h777f777f777f777f0001010101010001;

	lut_sub lut_2452 ({sk[468], n_n2037, x16038x, x16048x, n_n1876, x16037x}, n_n1813);
	defparam lut_2452.LUT_SIZE = 6;
	defparam lut_2452.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2458 ({sk[469], i_9_, i_7_, i_8_, i_6_, n_n390, n_n491}, x16065x);
	defparam lut_2458.LUT_SIZE = 7;
	defparam lut_2458.mask = 128'h777f777f777f777f0101010101010111;

	lut_sub lut_2468 ({sk[470], x10x, x519x, x309x, x16059x, x22101x, x22102x}, x16066x);
	defparam lut_2468.LUT_SIZE = 7;
	defparam lut_2468.mask = 128'h777f777f777f777fefffefffefffffff;

	lut_sub lut_2474 ({sk[471], x13x, x522x, x23x, x504x, n_n4239, x16068x}, x16070x);
	defparam lut_2474.LUT_SIZE = 7;
	defparam lut_2474.mask = 128'h777f777f777f777f777f777f777fffff;

	lut_sub lut_2479 ({sk[472], x16031x, x22099x, x22100x}, x16071x);
	defparam lut_2479.LUT_SIZE = 4;
	defparam lut_2479.mask = 16'h5fef;

	lut_sub lut_2483 ({sk[473], i_9_, i_7_, i_8_, i_6_, x498x, x473x}, x161x);
	defparam lut_2483.LUT_SIZE = 7;
	defparam lut_2483.mask = 128'h777f777f777f777f5000000300000000;

	lut_sub lut_2486 ({sk[474], i_9_, i_7_, i_8_, i_6_, n_n536, n_n500}, n_n1894);
	defparam lut_2486.LUT_SIZE = 7;
	defparam lut_2486.mask = 128'h777f777f777f777f1101001011110010;

	lut_sub lut_2496 ({sk[475], i_9_, i_7_, i_8_, i_6_, n_n536, n_n491}, n_n1893);
	defparam lut_2496.LUT_SIZE = 7;
	defparam lut_2496.mask = 128'h777f777f777f777f0101011100011110;

	lut_sub lut_2506 ({sk[476], x16x, x24x, x472x, x498x}, x16107x);
	defparam lut_2506.LUT_SIZE = 5;
	defparam lut_2506.mask = 32'h0fff0537;

	lut_sub lut_2509 ({sk[477], i_9_, i_7_, i_8_, i_6_, n_n536, n_n509}, x16111x);
	defparam lut_2509.LUT_SIZE = 7;
	defparam lut_2509.mask = 128'h777f777f777f777f0010100011001000;

	lut_sub lut_2515 ({sk[478], x161x, n_n1894, n_n1893, x16107x, x16111x}, x16114x);
	defparam lut_2515.LUT_SIZE = 6;
	defparam lut_2515.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2521 ({sk[479], x501x, x11x, x53x, x124x, x22098x}, n_n1896);
	defparam lut_2521.LUT_SIZE = 6;
	defparam lut_2521.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_2526 ({sk[480], x16x, x594x, x546x, x410x, n_n1703, x22330x}, x16086x);
	defparam lut_2526.LUT_SIZE = 7;
	defparam lut_2526.mask = 128'h777f777f777f777fbfbfbfbfbfffffff;

	lut_sub lut_2532 ({sk[481], x93x, x427x, x16101x, x16102x}, x16105x);
	defparam lut_2532.LUT_SIZE = 5;
	defparam lut_2532.mask = 32'h0fff7fff;

	lut_sub lut_2537 ({sk[482], x285x, x16094x, x16095x, x16097x, x22097x}, x16106x);
	defparam lut_2537.LUT_SIZE = 6;
	defparam lut_2537.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2543 ({sk[483], x20x, x23x, x497x, x443x, x16081x}, x16085x);
	defparam lut_2543.LUT_SIZE = 6;
	defparam lut_2543.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_2548 ({sk[484], x16119x, x16120x, n_n1866, x16130x}, n_n1810);
	defparam lut_2548.LUT_SIZE = 5;
	defparam lut_2548.mask = 32'h0fff7fff;

	lut_sub lut_2553 ({sk[485], x10x, x489x, x86x, x221x, x445x, x16132x}, n_n1870);
	defparam lut_2553.LUT_SIZE = 7;
	defparam lut_2553.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_2559 ({sk[486], x10x, x529x, x426x, x464x, x16138x}, x16144x);
	defparam lut_2559.LUT_SIZE = 6;
	defparam lut_2559.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_2564 ({sk[487], n_n2003, x259x, x16228x, x16234x, x16227x, x16230x}, x16239x);
	defparam lut_2564.LUT_SIZE = 7;
	defparam lut_2564.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_2571 ({sk[488], n_n4204, n_n3469, x219x, x80x, x16141x, x16236x}, x22094x);
	defparam lut_2571.LUT_SIZE = 7;
	defparam lut_2571.mask = 128'h777f777f777f777f8000000000000000;

	lut_sub lut_2573 ({sk[489], x21x, x12x, x587x, x578x}, x15580x);
	defparam lut_2573.LUT_SIZE = 5;
	defparam lut_2573.mask = 32'h0fff0357;

	lut_sub lut_2576 ({sk[490], i_9_, x492x, n_n491, n_n520, n_n130, x20x}, x15581x);
	defparam lut_2576.LUT_SIZE = 7;
	defparam lut_2576.mask = 128'h777f777f777f777f0013001300133333;

	lut_sub lut_2581 ({sk[491], x25x, x24x, x586x, x12x, x591x}, x16245x);
	defparam lut_2581.LUT_SIZE = 6;
	defparam lut_2581.mask = 64'h77ff77ff03575757;

	lut_sub lut_2585 ({sk[492], i_9_, i_7_, i_8_, i_6_, n_n482, n_n130}, n_n1833);
	defparam lut_2585.LUT_SIZE = 7;
	defparam lut_2585.mask = 128'h777f777f777f777f0110001011111010;

	lut_sub lut_2595 ({sk[493], i_9_, x519x, n_n130, x573x, x288x}, x16285x);
	defparam lut_2595.LUT_SIZE = 6;
	defparam lut_2595.mask = 64'h77ff77ff5555575f;

	lut_sub lut_2599 ({sk[494], i_9_, i_7_, i_8_, i_6_, n_n491, n_n130}, x16286x);
	defparam lut_2599.LUT_SIZE = 7;
	defparam lut_2599.mask = 128'h777f777f777f777f0000011001010010;

	lut_sub lut_2605 ({sk[495], x15580x, x15581x, x16245x, n_n1833, x16285x, x16286x}, x16289x);
	defparam lut_2605.LUT_SIZE = 7;
	defparam lut_2605.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_2612 ({sk[496], x22x, x11x, x533x, n_n1927, x22311x}, x16262x);
	defparam lut_2612.LUT_SIZE = 6;
	defparam lut_2612.mask = 64'h77ff77ffbbbfbfbf;

	lut_sub lut_2617 ({sk[497], x220x, x454x, x152x, x16254x, x22096x}, x16263x);
	defparam lut_2617.LUT_SIZE = 6;
	defparam lut_2617.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2623 ({sk[498], x19x, x477x, x319x, x386x, x22095x}, n_n1828);
	defparam lut_2623.LUT_SIZE = 6;
	defparam lut_2623.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_2628 ({sk[499], x11x, x555x, x385x, x16272x, x16270x}, n_n1829);
	defparam lut_2628.LUT_SIZE = 6;
	defparam lut_2628.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_2633 ({sk[500], x11x, x24x, x487x, x569x, x16277x, x16278x}, x16280x);
	defparam lut_2633.LUT_SIZE = 7;
	defparam lut_2633.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_2638 ({sk[501], i_9_, i_7_, i_8_, i_6_, n_n473, n_n65}, x117x);
	defparam lut_2638.LUT_SIZE = 7;
	defparam lut_2638.mask = 128'h777f777f777f777f0010101000101010;

	lut_sub lut_2645 ({sk[502], x515x, x19x, x24x, x508x}, x377x);
	defparam lut_2645.LUT_SIZE = 5;
	defparam lut_2645.mask = 32'h0fff0537;

	lut_sub lut_2648 ({sk[503], x592x, x19x, x20x, x493x}, x63x);
	defparam lut_2648.LUT_SIZE = 5;
	defparam lut_2648.mask = 32'h0fff0537;

	lut_sub lut_2651 ({sk[504], i_9_, i_7_, i_8_, i_6_, n_n473, n_n65}, x16309x);
	defparam lut_2651.LUT_SIZE = 7;
	defparam lut_2651.mask = 128'h777f777f777f777f0101000101000001;

	lut_sub lut_2657 ({sk[505], x515x, x19x, x23x, x524x, x489x, n_n5329}, x22090x);
	defparam lut_2657.LUT_SIZE = 7;
	defparam lut_2657.mask = 128'h777f777f777f777faaaa8080aa008000;

	lut_sub lut_2662 ({sk[506], x117x, x377x, x63x, x16309x, x22090x}, x16318x);
	defparam lut_2662.LUT_SIZE = 6;
	defparam lut_2662.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2668 ({sk[507], i_9_, i_1_, i_2_, i_0_, x493x}, n_n4404);
	defparam lut_2668.LUT_SIZE = 6;
	defparam lut_2668.mask = 64'h77ff77ff00000001;

	lut_sub lut_2670 ({sk[508], x538x, x16x, x20x, x499x}, x16472x);
	defparam lut_2670.LUT_SIZE = 5;
	defparam lut_2670.mask = 32'h0fff111f;

	lut_sub lut_2673 ({sk[509], x16x, x500x, x23x, x488x}, x16473x);
	defparam lut_2673.LUT_SIZE = 5;
	defparam lut_2673.mask = 32'h0fff0357;

	lut_sub lut_2676 ({sk[510], x16x, x500x, x20x, x580x, x503x}, x16475x);
	defparam lut_2676.LUT_SIZE = 6;
	defparam lut_2676.mask = 64'h77ff77ff000f777f;

	lut_sub lut_2680 ({sk[511], x15x, n_n4404, x495x, x16472x, x16473x, x16475x}, n_n2104);
	defparam lut_2680.LUT_SIZE = 7;
	defparam lut_2680.mask = 128'h777f777f777f777f7f7fffff7fffffff;

	lut_sub lut_2686 ({sk[512], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x522x);
	defparam lut_2686.LUT_SIZE = 7;
	defparam lut_2686.mask = 128'h777f777f777f777f0000000000008000;

	lut_sub lut_2688 ({sk[513], x25x, x24x, x547x, x543x, x523x}, x16493x);
	defparam lut_2688.LUT_SIZE = 6;
	defparam lut_2688.mask = 64'h77ff77ff003f557f;

	lut_sub lut_2692 ({sk[514], x25x, x21x, x24x, x543x, x504x, n_n4544}, x22060x);
	defparam lut_2692.LUT_SIZE = 7;
	defparam lut_2692.mask = 128'h777f777f777f777faa888888a0808080;

	lut_sub lut_2697 ({sk[515], x15x, x13x, x522x, x523x, x16493x, x22060x}, x16496x);
	defparam lut_2697.LUT_SIZE = 7;
	defparam lut_2697.mask = 128'h777f777f777f777fbbbbbbffbfbfbfff;

	lut_sub lut_2702 ({sk[516], x22x, x13x, x570x, x542x, x562x, x536x}, x16482x);
	defparam lut_2702.LUT_SIZE = 7;
	defparam lut_2702.mask = 128'h777f777f777f777f000077ff0f0f7fff;

	lut_sub lut_2707 ({sk[517], i_9_, i_7_, i_8_, i_6_, n_n455, n_n509}, x16483x);
	defparam lut_2707.LUT_SIZE = 7;
	defparam lut_2707.mask = 128'h777f777f777f777f0100001010100100;

	lut_sub lut_2713 ({sk[518], x25x, x10x, x545x, x472x, x561x, x548x}, x16487x);
	defparam lut_2713.LUT_SIZE = 7;
	defparam lut_2713.mask = 128'h777f777f777f777f00005fff33337fff;

	lut_sub lut_2718 ({sk[519], x10x, x20x, x547x, x537x}, x16485x);
	defparam lut_2718.LUT_SIZE = 5;
	defparam lut_2718.mask = 32'h0fff0357;

	lut_sub lut_2721 ({sk[520], x11x, x10x, x561x, x481x, x480x}, x16486x);
	defparam lut_2721.LUT_SIZE = 6;
	defparam lut_2721.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_2725 ({sk[521], x16482x, x16483x, x16487x, x16485x, x16486x}, x16497x);
	defparam lut_2725.LUT_SIZE = 6;
	defparam lut_2725.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2731 ({sk[522], i_9_, i_7_, i_8_, i_6_}, x21x);
	defparam lut_2731.LUT_SIZE = 5;
	defparam lut_2731.mask = 32'h0fff0800;

	lut_sub lut_2733 ({sk[523], x25x, x14x, x588x, x586x, x584x}, n_n2130);
	defparam lut_2733.LUT_SIZE = 6;
	defparam lut_2733.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_2737 ({sk[524], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x511x);
	defparam lut_2737.LUT_SIZE = 7;
	defparam lut_2737.mask = 128'h777f777f777f777f0000000040000000;

	lut_sub lut_2739 ({sk[525], i_9_, i_7_, i_8_, i_6_, x588x, x530x}, x16513x);
	defparam lut_2739.LUT_SIZE = 7;
	defparam lut_2739.mask = 128'h777f777f777f777f0003050000000000;

	lut_sub lut_2742 ({sk[526], x11x, x14x, x588x, x503x, x527x}, x22317x);
	defparam lut_2742.LUT_SIZE = 6;
	defparam lut_2742.mask = 64'h77ff77ffff88f080;

	lut_sub lut_2747 ({sk[527], x21x, n_n2130, x511x, x16513x, x22317x}, x16516x);
	defparam lut_2747.LUT_SIZE = 6;
	defparam lut_2747.mask = 64'h77ff77ffbbffbfff;

	lut_sub lut_2752 ({sk[528], n_n2263, x16527x, x16533x, x215x, x16523x}, n_n2190);
	defparam lut_2752.LUT_SIZE = 6;
	defparam lut_2752.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2758 ({sk[529], x16537x, x16535x, x16536x, x16540x, x16541x}, x16546x);
	defparam lut_2758.LUT_SIZE = 6;
	defparam lut_2758.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2764 ({sk[530], i_9_, i_7_, i_8_, i_6_, n_n536, n_n535}, x16542x);
	defparam lut_2764.LUT_SIZE = 7;
	defparam lut_2764.mask = 128'h777f777f777f777f1001000010100001;

	lut_sub lut_2770 ({sk[531], i_9_, i_7_, i_8_, i_6_, n_n536, n_n518}, x16543x);
	defparam lut_2770.LUT_SIZE = 7;
	defparam lut_2770.mask = 128'h777f777f777f777f0000111000100101;

	lut_sub lut_2777 ({sk[532], n_n2435, x54x, x282x}, x16555x);
	defparam lut_2777.LUT_SIZE = 4;
	defparam lut_2777.mask = 16'h5f7f;

	lut_sub lut_2781 ({sk[533], x16548x, x423x, n_n4275, x16550x, x22065x}, x16556x);
	defparam lut_2781.LUT_SIZE = 6;
	defparam lut_2781.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2787 ({sk[534], n_n2190, x16546x, x16542x, x16543x, x16555x, x16556x}, n_n2166);
	defparam lut_2787.LUT_SIZE = 7;
	defparam lut_2787.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_2794 ({sk[535], i_9_, i_7_, i_8_, i_6_, n_n455, n_n500}, n_n2257);
	defparam lut_2794.LUT_SIZE = 7;
	defparam lut_2794.mask = 128'h777f777f777f777f0100111101001101;

	lut_sub lut_2804 ({sk[536], i_9_, i_7_, i_8_, i_6_, n_n455, n_n509}, n_n2258);
	defparam lut_2804.LUT_SIZE = 7;
	defparam lut_2804.mask = 128'h777f777f777f777f1011110001011010;

	lut_sub lut_2814 ({sk[537], x25x, x13x, x573x, x542x}, x189x);
	defparam lut_2814.LUT_SIZE = 5;
	defparam lut_2814.mask = 32'h0fff0357;

	lut_sub lut_2817 ({sk[538], x15x, x13x, x24x, x572x, x542x}, x387x);
	defparam lut_2817.LUT_SIZE = 6;
	defparam lut_2817.mask = 64'h77ff77ff05375577;

	lut_sub lut_2821 ({sk[539], x13x, x23x, x491x, x574x, x560x, x541x}, x22082x);
	defparam lut_2821.LUT_SIZE = 7;
	defparam lut_2821.mask = 128'h777f777f777f777fffffaaaac0008000;

	lut_sub lut_2826 ({sk[540], n_n2257, n_n2258, x189x, x387x, x22082x}, x16598x);
	defparam lut_2826.LUT_SIZE = 6;
	defparam lut_2826.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2832 ({sk[541], n_n3889, x14515x, x14516x, x16564x, x16565x}, x16570x);
	defparam lut_2832.LUT_SIZE = 6;
	defparam lut_2832.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_2838 ({sk[542], x21x, n_n4247, x543x, n_n4517, x16582x, x16584x}, x16590x);
	defparam lut_2838.LUT_SIZE = 7;
	defparam lut_2838.mask = 128'h777f777f777f777f7f7fffff7fffffff;

	lut_sub lut_2844 ({sk[543], x15x, x504x, n_n889, x416x, x22324x}, n_n2253);
	defparam lut_2844.LUT_SIZE = 6;
	defparam lut_2844.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_2849 ({sk[544], n_n2261, x178x, x307x, x16566x, x16567x, x16586x}, x22081x);
	defparam lut_2849.LUT_SIZE = 7;
	defparam lut_2849.mask = 128'h777f777f777f777f8000000000000000;

	lut_sub lut_2851 ({sk[545], x22x, x523x, n_n4568, x455x, x121x, n_n4239}, n_n2251);
	defparam lut_2851.LUT_SIZE = 7;
	defparam lut_2851.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_2857 ({sk[546], x22x, x10x, x547x, x535x, x16605x, x16604x}, n_n2250);
	defparam lut_2857.LUT_SIZE = 7;
	defparam lut_2857.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_2862 ({sk[547], x16622x, x16611x, x16612x, x16617x, x22080x}, n_n2185);
	defparam lut_2862.LUT_SIZE = 6;
	defparam lut_2862.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_2868 ({sk[548], x10x, x23x, x561x, x573x, x271x, x16636x}, x16637x);
	defparam lut_2868.LUT_SIZE = 7;
	defparam lut_2868.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_2873 ({sk[549], x25x, x309x, x582x, x16627x, n_n2246, x16625x}, x16638x);
	defparam lut_2873.LUT_SIZE = 7;
	defparam lut_2873.mask = 128'h777f777f777f777f7f7fffff7fffffff;

	lut_sub lut_2879 ({sk[550], x24x, x523x, x429x, x212x, x213x, x16639x}, x16643x);
	defparam lut_2879.LUT_SIZE = 7;
	defparam lut_2879.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_2885 ({sk[551], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x560x);
	defparam lut_2885.LUT_SIZE = 7;
	defparam lut_2885.mask = 128'h777f777f777f777f2000000000000000;

	lut_sub lut_2887 ({sk[552], x16x, x501x, x20x, x478x, x473x}, x16650x);
	defparam lut_2887.LUT_SIZE = 6;
	defparam lut_2887.mask = 64'h77ff77ff050f373f;

	lut_sub lut_2891 ({sk[553], x25x, n_n4338, x20x, x497x, n_n4380, x473x}, x22062x);
	defparam lut_2891.LUT_SIZE = 7;
	defparam lut_2891.mask = 128'h777f777f777f777fccc0000088800000;

	lut_sub lut_2896 ({sk[554], x16x, x11x, x498x, x560x, x16650x, x22062x}, n_n2105);
	defparam lut_2896.LUT_SIZE = 7;
	defparam lut_2896.mask = 128'h777f777f777f777fbbbbbbffbfbfbfff;

	lut_sub lut_2901 ({sk[555], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x540x);
	defparam lut_2901.LUT_SIZE = 7;
	defparam lut_2901.mask = 128'h777f777f777f777f0000000000000004;

	lut_sub lut_2903 ({sk[556], x15x, x16x, x24x, x496x, x528x}, x16768x);
	defparam lut_2903.LUT_SIZE = 6;
	defparam lut_2903.mask = 64'h77ff77ff03573377;

	lut_sub lut_2907 ({sk[557], x15x, x16x, x544x, x522x, x525x, n_n4421}, x22061x);
	defparam lut_2907.LUT_SIZE = 7;
	defparam lut_2907.mask = 128'h777f777f777f777faaaa8080aa008000;

	lut_sub lut_2912 ({sk[558], x22x, x544x, x24x, x540x, x16768x, x22061x}, n_n2103);
	defparam lut_2912.LUT_SIZE = 7;
	defparam lut_2912.mask = 128'h777f777f777f777fbbbfbbbfbbbfffff;

	lut_sub lut_2917 ({sk[559], x19x, x556x, x16777x, x22063x, x22299x}, n_n2083);
	defparam lut_2917.LUT_SIZE = 6;
	defparam lut_2917.mask = 64'h77ff77ffefefefff;

	lut_sub lut_2922 ({sk[560], x25x, x22x, x484x, x589x, x16784x, x16783x}, n_n2095);
	defparam lut_2922.LUT_SIZE = 7;
	defparam lut_2922.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_2927 ({sk[561], x22x, x552x, n_n4813, x16808x, x16810x, x16811x}, n_n2096);
	defparam lut_2927.LUT_SIZE = 7;
	defparam lut_2927.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_2933 ({sk[562], x538x, x558x, x17x, x488x, x16816x, x16818x}, x16820x);
	defparam lut_2933.LUT_SIZE = 7;
	defparam lut_2933.mask = 128'h777f777f777f777f777f77ff77ff77ff;

	lut_sub lut_2939 ({sk[563], n_n2083, n_n2095, n_n2096, x16820x}, x16823x);
	defparam lut_2939.LUT_SIZE = 5;
	defparam lut_2939.mask = 32'h0fff7fff;

	lut_sub lut_2944 ({sk[564], i_1_, i_2_, i_0_}, n_n536);
	defparam lut_2944.LUT_SIZE = 4;
	defparam lut_2944.mask = 16'h5f01;

	lut_sub lut_2946 ({sk[565], i_7_, i_8_, i_6_}, n_n524);
	defparam lut_2946.LUT_SIZE = 4;
	defparam lut_2946.mask = 16'h5f08;

	lut_sub lut_2948 ({sk[566], i_5_, i_3_, i_4_}, n_n518);
	defparam lut_2948.LUT_SIZE = 4;
	defparam lut_2948.mask = 16'h5f10;

	lut_sub lut_2950 ({sk[567], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x521x);
	defparam lut_2950.LUT_SIZE = 7;
	defparam lut_2950.mask = 128'h777f777f777f777f0000000010000000;

	lut_sub lut_2952 ({sk[568], i_9_, i_1_, i_2_, i_0_, x521x}, n_n4338);
	defparam lut_2952.LUT_SIZE = 6;
	defparam lut_2952.mask = 64'h77ff77ff00000001;

	lut_sub lut_2954 ({sk[569], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x501x);
	defparam lut_2954.LUT_SIZE = 7;
	defparam lut_2954.mask = 128'h777f777f777f777f0000000100000000;

	lut_sub lut_2956 ({sk[570], i_7_, i_8_, i_6_}, n_n526);
	defparam lut_2956.LUT_SIZE = 4;
	defparam lut_2956.mask = 16'h5f02;

	lut_sub lut_2958 ({sk[571], i_5_, i_3_, i_4_}, n_n482);
	defparam lut_2958.LUT_SIZE = 4;
	defparam lut_2958.mask = 16'h5f40;

	lut_sub lut_2960 ({sk[572], i_1_, i_2_, i_0_}, n_n455);
	defparam lut_2960.LUT_SIZE = 4;
	defparam lut_2960.mask = 16'h5f04;

	lut_sub lut_2962 ({sk[573], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x539x);
	defparam lut_2962.LUT_SIZE = 7;
	defparam lut_2962.mask = 128'h777f777f777f777f0000000000001000;

	lut_sub lut_2964 ({sk[574], i_7_, i_8_, i_6_}, n_n528);
	defparam lut_2964.LUT_SIZE = 4;
	defparam lut_2964.mask = 16'h5f40;

	lut_sub lut_2966 ({sk[575], i_1_, i_2_, i_0_}, n_n390);
	defparam lut_2966.LUT_SIZE = 4;
	defparam lut_2966.mask = 16'h5f10;

	lut_sub lut_2968 ({sk[576], i_5_, i_3_, i_4_}, n_n473);
	defparam lut_2968.LUT_SIZE = 4;
	defparam lut_2968.mask = 16'h5f08;

	lut_sub lut_2970 ({sk[577], i_7_, i_8_, i_6_}, n_n532);
	defparam lut_2970.LUT_SIZE = 4;
	defparam lut_2970.mask = 16'h5f04;

	lut_sub lut_2972 ({sk[578], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x509x);
	defparam lut_2972.LUT_SIZE = 7;
	defparam lut_2972.mask = 128'h777f777f777f777f0000000000080000;

	lut_sub lut_2974 ({sk[579], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x507x);
	defparam lut_2974.LUT_SIZE = 7;
	defparam lut_2974.mask = 128'h777f777f777f777f0000000010000000;

	lut_sub lut_2976 ({sk[580], i_7_, i_8_, i_6_}, n_n534);
	defparam lut_2976.LUT_SIZE = 4;
	defparam lut_2976.mask = 16'h5f01;

	lut_sub lut_2978 ({sk[581], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x510x);
	defparam lut_2978.LUT_SIZE = 7;
	defparam lut_2978.mask = 128'h777f777f777f777f0000000000000008;

	lut_sub lut_2980 ({sk[582], i_5_, i_3_, i_4_}, n_n509);
	defparam lut_2980.LUT_SIZE = 4;
	defparam lut_2980.mask = 16'h5f02;

	lut_sub lut_2982 ({sk[583], i_1_, i_2_, i_0_}, n_n325);
	defparam lut_2982.LUT_SIZE = 4;
	defparam lut_2982.mask = 16'h5f40;

	lut_sub lut_2984 ({sk[584], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x483x);
	defparam lut_2984.LUT_SIZE = 7;
	defparam lut_2984.mask = 128'h777f777f777f777f0000000000004000;

	lut_sub lut_2986 ({sk[585], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x558x);
	defparam lut_2986.LUT_SIZE = 7;
	defparam lut_2986.mask = 128'h777f777f777f777f0400000000000000;

	lut_sub lut_2988 ({sk[586], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x588x);
	defparam lut_2988.LUT_SIZE = 7;
	defparam lut_2988.mask = 128'h777f777f777f777f0040000000000000;

	lut_sub lut_2990 ({sk[587], i_1_, i_2_, i_0_}, n_n260);
	defparam lut_2990.LUT_SIZE = 4;
	defparam lut_2990.mask = 16'h5f02;

	lut_sub lut_2992 ({sk[588], i_5_, i_3_, i_4_}, n_n535);
	defparam lut_2992.LUT_SIZE = 4;
	defparam lut_2992.mask = 16'h5f01;

	lut_sub lut_2994 ({sk[589], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x545x);
	defparam lut_2994.LUT_SIZE = 7;
	defparam lut_2994.mask = 128'h777f777f777f777f0001000000000000;

	lut_sub lut_2996 ({sk[590], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x552x);
	defparam lut_2996.LUT_SIZE = 7;
	defparam lut_2996.mask = 128'h777f777f777f777f0000000000000002;

	lut_sub lut_2998 ({sk[591], i_7_, i_8_, i_6_}, n_n522);
	defparam lut_2998.LUT_SIZE = 4;
	defparam lut_2998.mask = 16'h5f20;

	lut_sub lut_3000 ({sk[592], i_5_, i_3_, i_4_}, n_n491);
	defparam lut_3000.LUT_SIZE = 4;
	defparam lut_3000.mask = 16'h5f04;

	lut_sub lut_3002 ({sk[593], i_7_, i_8_, i_6_}, n_n520);
	defparam lut_3002.LUT_SIZE = 4;
	defparam lut_3002.mask = 16'h5f80;

	lut_sub lut_3004 ({sk[594], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x570x);
	defparam lut_3004.LUT_SIZE = 7;
	defparam lut_3004.mask = 128'h777f777f777f777f0040000000000000;

	lut_sub lut_3006 ({sk[595], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x519x);
	defparam lut_3006.LUT_SIZE = 7;
	defparam lut_3006.mask = 128'h777f777f777f777f0000000000400000;

	lut_sub lut_3008 ({sk[596], i_1_, i_2_, i_0_}, n_n195);
	defparam lut_3008.LUT_SIZE = 4;
	defparam lut_3008.mask = 16'h5f08;

	lut_sub lut_3010 ({sk[597], i_9_, i_1_, i_2_, i_0_}, x18x);
	defparam lut_3010.LUT_SIZE = 5;
	defparam lut_3010.mask = 32'h0fff0008;

	lut_sub lut_3012 ({sk[598], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x597x);
	defparam lut_3012.LUT_SIZE = 7;
	defparam lut_3012.mask = 128'h777f777f777f777f0000000800000000;

	lut_sub lut_3014 ({sk[599], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x586x);
	defparam lut_3014.LUT_SIZE = 7;
	defparam lut_3014.mask = 128'h777f777f777f777f0000000004000000;

	lut_sub lut_3016 ({sk[600], i_1_, i_2_, i_0_}, n_n130);
	defparam lut_3016.LUT_SIZE = 4;
	defparam lut_3016.mask = 16'h5f20;

	lut_sub lut_3018 ({sk[601], i_9_, i_1_, i_2_, i_0_}, x12x);
	defparam lut_3018.LUT_SIZE = 5;
	defparam lut_3018.mask = 32'h0fff0020;

	lut_sub lut_3020 ({sk[602], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x490x);
	defparam lut_3020.LUT_SIZE = 7;
	defparam lut_3020.mask = 128'h777f777f777f777f0000001000000000;

	lut_sub lut_3022 ({sk[603], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x554x);
	defparam lut_3022.LUT_SIZE = 7;
	defparam lut_3022.mask = 128'h777f777f777f777f0000000000000020;

	lut_sub lut_3024 ({sk[604], x21x, x12x, x490x, x20x, x554x}, n_n4148);
	defparam lut_3024.LUT_SIZE = 6;
	defparam lut_3024.mask = 64'h77ff77ff111f555f;

	lut_sub lut_3028 ({sk[605], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x516x);
	defparam lut_3028.LUT_SIZE = 7;
	defparam lut_3028.mask = 128'h777f777f777f777f0000000080000000;

	lut_sub lut_3030 ({sk[606], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x496x);
	defparam lut_3030.LUT_SIZE = 7;
	defparam lut_3030.mask = 128'h777f777f777f777f0100000000000000;

	lut_sub lut_3032 ({sk[607], i_9_, i_7_, i_8_, i_6_, x496x}, n_n4433);
	defparam lut_3032.LUT_SIZE = 6;
	defparam lut_3032.mask = 64'h77ff77ff00040000;

	lut_sub lut_3034 ({sk[608], i_9_, i_7_, i_8_, i_6_, x496x}, x98x);
	defparam lut_3034.LUT_SIZE = 6;
	defparam lut_3034.mask = 64'h77ff77ff10040000;

	lut_sub lut_3037 ({sk[609], x16x, x23x, x496x, x525x}, x233x);
	defparam lut_3037.LUT_SIZE = 5;
	defparam lut_3037.mask = 32'h0fff0357;

	lut_sub lut_3040 ({sk[610], x16x, x20x, x496x, x489x}, x236x);
	defparam lut_3040.LUT_SIZE = 5;
	defparam lut_3040.mask = 32'h0fff0357;

	lut_sub lut_3043 ({sk[611], i_5_, i_3_, i_4_}, n_n464);
	defparam lut_3043.LUT_SIZE = 4;
	defparam lut_3043.mask = 16'h5f80;

	lut_sub lut_3045 ({sk[612], i_9_, n_n536, n_n520, x236x, n_n464}, x13428x);
	defparam lut_3045.LUT_SIZE = 6;
	defparam lut_3045.mask = 64'h77ff77ff33373337;

	lut_sub lut_3049 ({sk[613], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x595x);
	defparam lut_3049.LUT_SIZE = 7;
	defparam lut_3049.mask = 128'h777f777f777f777f0000004000000000;

	lut_sub lut_3051 ({sk[614], x15x, x14x, x595x, x559x}, x241x);
	defparam lut_3051.LUT_SIZE = 5;
	defparam lut_3051.mask = 32'h0fff0537;

	lut_sub lut_3054 ({sk[615], x15x, x539x, x14x, x595x, x559x}, n_n4216);
	defparam lut_3054.LUT_SIZE = 6;
	defparam lut_3054.mask = 64'h77ff77ff050f373f;

	lut_sub lut_3058 ({sk[616], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x484x);
	defparam lut_3058.LUT_SIZE = 7;
	defparam lut_3058.mask = 128'h777f777f777f777f0000000000000200;

	lut_sub lut_3060 ({sk[617], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x482x);
	defparam lut_3060.LUT_SIZE = 7;
	defparam lut_3060.mask = 128'h777f777f777f777f0000000000000002;

	lut_sub lut_3062 ({sk[618], i_9_, i_5_, i_3_, i_4_, n_n260, n_n520}, x102x);
	defparam lut_3062.LUT_SIZE = 7;
	defparam lut_3062.mask = 128'h777f777f777f777f0001000000010000;

	lut_sub lut_3065 ({sk[619], i_9_, n_n518, n_n532, n_n509, n_n260, n_n520}, x13170x);
	defparam lut_3065.LUT_SIZE = 7;
	defparam lut_3065.mask = 128'h777f777f777f777f0003111300031113;

	lut_sub lut_3070 ({sk[620], i_9_, i_7_, i_8_, i_6_, n_n509, n_n260}, x13171x);
	defparam lut_3070.LUT_SIZE = 7;
	defparam lut_3070.mask = 128'h777f777f777f777f0100001101000001;

	lut_sub lut_3076 ({sk[621], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x485x);
	defparam lut_3076.LUT_SIZE = 7;
	defparam lut_3076.mask = 128'h777f777f777f777f0000000000000800;

	lut_sub lut_3078 ({sk[622], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x567x);
	defparam lut_3078.LUT_SIZE = 7;
	defparam lut_3078.mask = 128'h777f777f777f777f0000080000000000;

	lut_sub lut_3080 ({sk[623], x25x, x18x, x564x, x567x}, x103x);
	defparam lut_3080.LUT_SIZE = 5;
	defparam lut_3080.mask = 32'h0fff0357;

	lut_sub lut_3083 ({sk[624], i_9_, i_7_, i_8_, i_6_, n_n509, n_n195}, x13380x);
	defparam lut_3083.LUT_SIZE = 7;
	defparam lut_3083.mask = 128'h777f777f777f777f0100100000100010;

	lut_sub lut_3088 ({sk[625], i_5_, i_3_, i_4_}, n_n500);
	defparam lut_3088.LUT_SIZE = 4;
	defparam lut_3088.mask = 16'h5f20;

	lut_sub lut_3090 ({sk[626], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x561x);
	defparam lut_3090.LUT_SIZE = 7;
	defparam lut_3090.mask = 128'h777f777f777f777f0000100000000000;

	lut_sub lut_3092 ({sk[627], i_7_, i_8_, i_6_}, n_n530);
	defparam lut_3092.LUT_SIZE = 4;
	defparam lut_3092.mask = 16'h5f10;

	lut_sub lut_3094 ({sk[628], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x571x);
	defparam lut_3094.LUT_SIZE = 7;
	defparam lut_3094.mask = 128'h777f777f777f777f0000000000100000;

	lut_sub lut_3096 ({sk[629], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x479x);
	defparam lut_3096.LUT_SIZE = 7;
	defparam lut_3096.mask = 128'h777f777f777f777f0000000000001000;

	lut_sub lut_3098 ({sk[630], i_9_, i_7_, i_8_, i_6_, x479x}, n_n4613);
	defparam lut_3098.LUT_SIZE = 6;
	defparam lut_3098.mask = 64'h77ff77ff04000000;

	lut_sub lut_3100 ({sk[631], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x512x);
	defparam lut_3100.LUT_SIZE = 7;
	defparam lut_3100.mask = 128'h777f777f777f777f0000000002000000;

	lut_sub lut_3102 ({sk[632], i_9_, i_1_, i_2_, i_0_, x510x}, n_n4920);
	defparam lut_3102.LUT_SIZE = 6;
	defparam lut_3102.mask = 64'h77ff77ff00000004;

	lut_sub lut_3104 ({sk[633], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x557x);
	defparam lut_3104.LUT_SIZE = 7;
	defparam lut_3104.mask = 128'h777f777f777f777f0004000000000000;

	lut_sub lut_3106 ({sk[634], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x572x);
	defparam lut_3106.LUT_SIZE = 7;
	defparam lut_3106.mask = 128'h777f777f777f777f0000000400000000;

	lut_sub lut_3108 ({sk[635], i_9_, i_1_, i_2_, i_0_, x572x}, n_n4380);
	defparam lut_3108.LUT_SIZE = 6;
	defparam lut_3108.mask = 64'h77ff77ff00000001;

	lut_sub lut_3110 ({sk[636], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x508x);
	defparam lut_3110.LUT_SIZE = 7;
	defparam lut_3110.mask = 128'h777f777f777f777f0000000800000000;

	lut_sub lut_3112 ({sk[637], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x581x);
	defparam lut_3112.LUT_SIZE = 7;
	defparam lut_3112.mask = 128'h777f777f777f777f1000000000000000;

	lut_sub lut_3114 ({sk[638], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x590x);
	defparam lut_3114.LUT_SIZE = 7;
	defparam lut_3114.mask = 128'h777f777f777f777f0008000000000000;

	lut_sub lut_3116 ({sk[639], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x587x);
	defparam lut_3116.LUT_SIZE = 7;
	defparam lut_3116.mask = 128'h777f777f777f777f0000000000000400;

	lut_sub lut_3118 ({sk[640], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x598x);
	defparam lut_3118.LUT_SIZE = 7;
	defparam lut_3118.mask = 128'h777f777f777f777f0000002000000000;

	lut_sub lut_3120 ({sk[641], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x591x);
	defparam lut_3120.LUT_SIZE = 7;
	defparam lut_3120.mask = 128'h777f777f777f777f0020000000000000;

	lut_sub lut_3122 ({sk[642], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x580x);
	defparam lut_3122.LUT_SIZE = 7;
	defparam lut_3122.mask = 128'h777f777f777f777f4000000000000000;

	lut_sub lut_3124 ({sk[643], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x583x);
	defparam lut_3124.LUT_SIZE = 7;
	defparam lut_3124.mask = 128'h777f777f777f777f0000001000000000;

	lut_sub lut_3126 ({sk[644], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x481x);
	defparam lut_3126.LUT_SIZE = 7;
	defparam lut_3126.mask = 128'h777f777f777f777f0000000000020000;

	lut_sub lut_3128 ({sk[645], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x518x);
	defparam lut_3128.LUT_SIZE = 7;
	defparam lut_3128.mask = 128'h777f777f777f777f0000000020000000;

	lut_sub lut_3130 ({sk[646], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x565x);
	defparam lut_3130.LUT_SIZE = 7;
	defparam lut_3130.mask = 128'h777f777f777f777f0000400000000000;

	lut_sub lut_3132 ({sk[647], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x491x);
	defparam lut_3132.LUT_SIZE = 7;
	defparam lut_3132.mask = 128'h777f777f777f777f0000200000000000;

	lut_sub lut_3134 ({sk[648], i_9_, i_7_, i_8_, i_6_, n_n325, n_n500}, n_n3336);
	defparam lut_3134.LUT_SIZE = 7;
	defparam lut_3134.mask = 128'h777f777f777f777f0111010001111001;

	lut_sub lut_3144 ({sk[649], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x566x);
	defparam lut_3144.LUT_SIZE = 7;
	defparam lut_3144.mask = 128'h777f777f777f777f0000020000000000;

	lut_sub lut_3146 ({sk[650], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x574x);
	defparam lut_3146.LUT_SIZE = 7;
	defparam lut_3146.mask = 128'h777f777f777f777f0000000000000004;

	lut_sub lut_3148 ({sk[651], x21x, x17x, x518x, x491x, x566x}, n_n3451);
	defparam lut_3148.LUT_SIZE = 6;
	defparam lut_3148.mask = 64'h77ff77ff003f557f;

	lut_sub lut_3152 ({sk[652], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x577x);
	defparam lut_3152.LUT_SIZE = 7;
	defparam lut_3152.mask = 128'h777f777f777f777f0000000000080000;

	lut_sub lut_3154 ({sk[653], x22x, x21x, x519x, x18x, x577x}, n_n3424);
	defparam lut_3154.LUT_SIZE = 6;
	defparam lut_3154.mask = 64'h77ff77ff03575757;

	lut_sub lut_3158 ({sk[654], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x514x);
	defparam lut_3158.LUT_SIZE = 7;
	defparam lut_3158.mask = 128'h777f777f777f777f0000000020000000;

	lut_sub lut_3160 ({sk[655], x509x, x24x, x12x, x514x}, x114x);
	defparam lut_3160.LUT_SIZE = 5;
	defparam lut_3160.mask = 32'h0fff0537;

	lut_sub lut_3163 ({sk[656], i_9_, i_7_, i_8_, i_6_, x514x}, n_n5181);
	defparam lut_3163.LUT_SIZE = 6;
	defparam lut_3163.mask = 64'h77ff77ff01000000;

	lut_sub lut_3165 ({sk[657], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x503x);
	defparam lut_3165.LUT_SIZE = 7;
	defparam lut_3165.mask = 128'h777f777f777f777f0000000000000080;

	lut_sub lut_3167 ({sk[658], i_9_, i_7_, i_8_, i_6_, n_n473, n_n130}, n_n3303);
	defparam lut_3167.LUT_SIZE = 7;
	defparam lut_3167.mask = 128'h777f777f777f777f0101111000011110;

	lut_sub lut_3177 ({sk[659], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x505x);
	defparam lut_3177.LUT_SIZE = 7;
	defparam lut_3177.mask = 128'h777f777f777f777f0008000000000000;

	lut_sub lut_3179 ({sk[660], i_9_, i_1_, i_2_, i_0_, x505x}, n_n5310);
	defparam lut_3179.LUT_SIZE = 6;
	defparam lut_3179.mask = 64'h77ff77ff00004000;

	lut_sub lut_3181 ({sk[661], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x506x);
	defparam lut_3181.LUT_SIZE = 7;
	defparam lut_3181.mask = 128'h777f777f777f777f0080000000000000;

	lut_sub lut_3183 ({sk[662], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x488x);
	defparam lut_3183.LUT_SIZE = 7;
	defparam lut_3183.mask = 128'h777f777f777f777f0000008000000000;

	lut_sub lut_3185 ({sk[663], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x502x);
	defparam lut_3185.LUT_SIZE = 7;
	defparam lut_3185.mask = 128'h777f777f777f777f0000000000800000;

	lut_sub lut_3187 ({sk[664], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x534x);
	defparam lut_3187.LUT_SIZE = 7;
	defparam lut_3187.mask = 128'h777f777f777f777f8000000000000000;

	lut_sub lut_3189 ({sk[665], i_9_, i_7_, i_8_, i_6_, x515x, x534x}, x268x);
	defparam lut_3189.LUT_SIZE = 7;
	defparam lut_3189.mask = 128'h777f777f777f777f3000000500000000;

	lut_sub lut_3192 ({sk[666], i_1_, i_2_, i_0_}, n_n65);
	defparam lut_3192.LUT_SIZE = 4;
	defparam lut_3192.mask = 16'h5f80;

	lut_sub lut_3194 ({sk[667], i_9_, i_7_, i_8_, i_6_, n_n473, n_n65}, x13934x);
	defparam lut_3194.LUT_SIZE = 7;
	defparam lut_3194.mask = 128'h777f777f777f777f0000001011000010;

	lut_sub lut_3199 ({sk[668], i_9_, n_n534, x268x, n_n464, n_n65}, x13933x);
	defparam lut_3199.LUT_SIZE = 6;
	defparam lut_3199.mask = 64'h77ff77ff0f0f0f1f;

	lut_sub lut_3202 ({sk[669], x19x, x488x, x502x, x13934x, x13933x}, n_n3292);
	defparam lut_3202.LUT_SIZE = 6;
	defparam lut_3202.mask = 64'h77ff77ff77777fff;

	lut_sub lut_3207 ({sk[670], i_9_, i_1_, i_2_, i_0_, x564x}, n_n4616);
	defparam lut_3207.LUT_SIZE = 6;
	defparam lut_3207.mask = 64'h77ff77ff00000100;

	lut_sub lut_3209 ({sk[671], i_9_, i_7_, i_8_, i_6_, x479x}, n_n4607);
	defparam lut_3209.LUT_SIZE = 6;
	defparam lut_3209.mask = 64'h77ff77ff10000000;

	lut_sub lut_3211 ({sk[672], x22x, x10x, x472x, x479x}, x273x);
	defparam lut_3211.LUT_SIZE = 5;
	defparam lut_3211.mask = 32'h0fff0357;

	lut_sub lut_3214 ({sk[673], i_9_, i_1_, i_2_, i_0_, x477x, x475x}, x396x);
	defparam lut_3214.LUT_SIZE = 7;
	defparam lut_3214.mask = 128'h777f777f777f777f0000000000070000;

	lut_sub lut_3217 ({sk[674], x25x, x20x, x23x, x561x, x479x, n_n4616}, x22170x);
	defparam lut_3217.LUT_SIZE = 7;
	defparam lut_3217.mask = 128'h777f777f777f777faa888888a0808080;

	lut_sub lut_3222 ({sk[675], x11x, x479x, x273x, x396x, x22170x}, n_n3346);
	defparam lut_3222.LUT_SIZE = 6;
	defparam lut_3222.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_3227 ({sk[676], x22x, x10x, x561x, x518x, x536x}, n_n1649);
	defparam lut_3227.LUT_SIZE = 6;
	defparam lut_3227.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_3231 ({sk[677], i_9_, i_7_, i_8_, i_6_, x561x}, x118x);
	defparam lut_3231.LUT_SIZE = 6;
	defparam lut_3231.mask = 64'h77ff77ff01100000;

	lut_sub lut_3234 ({sk[678], i_9_, i_7_, i_8_, i_6_, x571x}, x309x);
	defparam lut_3234.LUT_SIZE = 6;
	defparam lut_3234.mask = 64'h77ff77ff04400000;

	lut_sub lut_3237 ({sk[679], x11x, x10x, x519x, x571x}, x348x);
	defparam lut_3237.LUT_SIZE = 5;
	defparam lut_3237.mask = 32'h0fff0357;

	lut_sub lut_3240 ({sk[680], x10x, x23x, x561x, x574x}, x349x);
	defparam lut_3240.LUT_SIZE = 5;
	defparam lut_3240.mask = 32'h0fff0357;

	lut_sub lut_3243 ({sk[681], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x513x);
	defparam lut_3243.LUT_SIZE = 7;
	defparam lut_3243.mask = 128'h777f777f777f777f0000000008000000;

	lut_sub lut_3245 ({sk[682], i_9_, i_1_, i_2_, i_0_, x506x, x529x}, x120x);
	defparam lut_3245.LUT_SIZE = 7;
	defparam lut_3245.mask = 128'h777f777f777f777f0000000000007000;

	lut_sub lut_3248 ({sk[683], i_9_, i_7_, i_8_, i_6_, n_n473, n_n195}, x13981x);
	defparam lut_3248.LUT_SIZE = 7;
	defparam lut_3248.mask = 128'h777f777f777f777f0000001000101100;

	lut_sub lut_3253 ({sk[684], i_9_, i_7_, i_8_, i_6_, n_n482, n_n195}, x230x);
	defparam lut_3253.LUT_SIZE = 7;
	defparam lut_3253.mask = 128'h777f777f777f777f0100001001001010;

	lut_sub lut_3259 ({sk[685], i_9_, i_5_, i_3_, i_4_, n_n532, n_n195}, x231x);
	defparam lut_3259.LUT_SIZE = 7;
	defparam lut_3259.mask = 128'h777f777f777f777f0100000001000000;

	lut_sub lut_3262 ({sk[686], x492x, x18x, n_n3424, x584x, x230x}, x13991x);
	defparam lut_3262.LUT_SIZE = 6;
	defparam lut_3262.mask = 64'h77ff77ff5f7f5fff;

	lut_sub lut_3267 ({sk[687], x11x, x18x, x505x, x513x}, x13979x);
	defparam lut_3267.LUT_SIZE = 5;
	defparam lut_3267.mask = 32'h0fff0357;

	lut_sub lut_3270 ({sk[688], x21x, x18x, x506x, x529x, x513x}, x13980x);
	defparam lut_3270.LUT_SIZE = 6;
	defparam lut_3270.mask = 64'h77ff77ff003f557f;

	lut_sub lut_3274 ({sk[689], i_9_, n_n482, n_n532, n_n491, n_n520, n_n195}, x13987x);
	defparam lut_3274.LUT_SIZE = 7;
	defparam lut_3274.mask = 128'h777f777f777f777f0101015501010155;

	lut_sub lut_3279 ({sk[690], x510x, x18x, x587x, x580x, x493x}, x13988x);
	defparam lut_3279.LUT_SIZE = 6;
	defparam lut_3279.mask = 64'h77ff77ff007f00ff;

	lut_sub lut_3284 ({sk[691], x13981x, x13979x, x13980x, x13987x, x13988x}, x13992x);
	defparam lut_3284.LUT_SIZE = 6;
	defparam lut_3284.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_3290 ({sk[692], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x547x);
	defparam lut_3290.LUT_SIZE = 7;
	defparam lut_3290.mask = 128'h777f777f777f777f0000000000000010;

	lut_sub lut_3292 ({sk[693], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x549x);
	defparam lut_3292.LUT_SIZE = 7;
	defparam lut_3292.mask = 128'h777f777f777f777f0000000000010000;

	lut_sub lut_3294 ({sk[694], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x596x);
	defparam lut_3294.LUT_SIZE = 7;
	defparam lut_3294.mask = 128'h777f777f777f777f0000000200000000;

	lut_sub lut_3296 ({sk[695], i_9_, i_7_, i_8_, i_6_, x554x}, n_n5085);
	defparam lut_3296.LUT_SIZE = 6;
	defparam lut_3296.mask = 64'h77ff77ff01000000;

	lut_sub lut_3298 ({sk[696], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x494x);
	defparam lut_3298.LUT_SIZE = 7;
	defparam lut_3298.mask = 128'h777f777f777f777f0000100000000000;

	lut_sub lut_3300 ({sk[697], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x486x);
	defparam lut_3300.LUT_SIZE = 7;
	defparam lut_3300.mask = 128'h777f777f777f777f0000000000002000;

	lut_sub lut_3302 ({sk[698], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x568x);
	defparam lut_3302.LUT_SIZE = 7;
	defparam lut_3302.mask = 128'h777f777f777f777f0000200000000000;

	lut_sub lut_3304 ({sk[699], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x578x);
	defparam lut_3304.LUT_SIZE = 7;
	defparam lut_3304.mask = 128'h777f777f777f777f0000000000200000;

	lut_sub lut_3306 ({sk[700], x21x, x12x, x598x, x563x, x560x, x486x}, x13696x);
	defparam lut_3306.LUT_SIZE = 7;
	defparam lut_3306.mask = 128'h777f777f777f777f00003f3f55ff7fff;

	lut_sub lut_3311 ({sk[701], x15x, x492x, x12x, x581x, x598x}, x13695x);
	defparam lut_3311.LUT_SIZE = 6;
	defparam lut_3311.mask = 64'h77ff77ff030f575f;

	lut_sub lut_3315 ({sk[702], i_9_, i_1_, i_2_, i_0_, x492x}, n_n4388);
	defparam lut_3315.LUT_SIZE = 6;
	defparam lut_3315.mask = 64'h77ff77ff00000001;

	lut_sub lut_3317 ({sk[703], i_9_, i_7_, i_8_, i_6_, x540x}, n_n4455);
	defparam lut_3317.LUT_SIZE = 6;
	defparam lut_3317.mask = 64'h77ff77ff40000000;

	lut_sub lut_3319 ({sk[704], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x537x);
	defparam lut_3319.LUT_SIZE = 7;
	defparam lut_3319.mask = 128'h777f777f777f777f0000000000000040;

	lut_sub lut_3321 ({sk[705], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x480x);
	defparam lut_3321.LUT_SIZE = 7;
	defparam lut_3321.mask = 128'h777f777f777f777f0000000200000000;

	lut_sub lut_3323 ({sk[706], i_9_, i_7_, i_8_, i_6_, x512x}, n_n4925);
	defparam lut_3323.LUT_SIZE = 6;
	defparam lut_3323.mask = 64'h77ff77ff01000000;

	lut_sub lut_3325 ({sk[707], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x520x);
	defparam lut_3325.LUT_SIZE = 7;
	defparam lut_3325.mask = 128'h777f777f777f777f0000000040000000;

	lut_sub lut_3327 ({sk[708], i_9_, i_7_, i_8_, i_6_, x595x}, n_n4727);
	defparam lut_3327.LUT_SIZE = 6;
	defparam lut_3327.mask = 64'h77ff77ff40000000;

	lut_sub lut_3329 ({sk[709], x14x, x20x, x581x, x595x}, x101x);
	defparam lut_3329.LUT_SIZE = 5;
	defparam lut_3329.mask = 32'h0fff0537;

	lut_sub lut_3332 ({sk[710], x14x, x20x, x482x, x581x, x481x, x595x}, x15746x);
	defparam lut_3332.LUT_SIZE = 7;
	defparam lut_3332.mask = 128'h777f777f777f777f000055553fff7fff;

	lut_sub lut_3337 ({sk[711], i_9_, i_7_, i_8_, i_6_, n_n509, n_n260}, n_n2970);
	defparam lut_3337.LUT_SIZE = 7;
	defparam lut_3337.mask = 128'h777f777f777f777f0011010011110110;

	lut_sub lut_3347 ({sk[712], i_9_, i_1_, i_2_, i_0_, x557x}, n_n5022);
	defparam lut_3347.LUT_SIZE = 6;
	defparam lut_3347.mask = 64'h77ff77ff00000040;

	lut_sub lut_3349 ({sk[713], i_9_, i_7_, i_8_, i_6_, x577x}, n_n5017);
	defparam lut_3349.LUT_SIZE = 6;
	defparam lut_3349.mask = 64'h77ff77ff00010000;

	lut_sub lut_3351 ({sk[714], i_9_, i_7_, i_8_, i_6_, n_n195, n_n500}, x135x);
	defparam lut_3351.LUT_SIZE = 7;
	defparam lut_3351.mask = 128'h777f777f777f777f1000000010000000;

	lut_sub lut_3354 ({sk[715], x24x, x18x, x572x, x577x}, x298x);
	defparam lut_3354.LUT_SIZE = 5;
	defparam lut_3354.mask = 32'h0fff0357;

	lut_sub lut_3357 ({sk[716], i_9_, i_7_, i_8_, i_6_, n_n491, n_n195}, x15704x);
	defparam lut_3357.LUT_SIZE = 7;
	defparam lut_3357.mask = 128'h777f777f777f777f0101010000010000;

	lut_sub lut_3362 ({sk[717], x21x, x474x, x18x, x485x, x472x}, n_n1576);
	defparam lut_3362.LUT_SIZE = 6;
	defparam lut_3362.mask = 64'h77ff77ff050f373f;

	lut_sub lut_3366 ({sk[718], i_9_, n_n509, n_n195, n_n530, x581x, x494x}, x14938x);
	defparam lut_3366.LUT_SIZE = 7;
	defparam lut_3366.mask = 128'h777f777f777f777f0000000f0077007f;

	lut_sub lut_3371 ({sk[719], i_9_, i_7_, i_8_, i_6_, n_n509, n_n195}, x14939x);
	defparam lut_3371.LUT_SIZE = 7;
	defparam lut_3371.mask = 128'h777f777f777f777f0000111000101000;

	lut_sub lut_3377 ({sk[720], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x562x);
	defparam lut_3377.LUT_SIZE = 7;
	defparam lut_3377.mask = 128'h777f777f777f777f0000020000000000;

	lut_sub lut_3379 ({sk[721], x11x, x18x, x567x, x556x}, x136x);
	defparam lut_3379.LUT_SIZE = 5;
	defparam lut_3379.mask = 32'h0fff0537;

	lut_sub lut_3382 ({sk[722], x18x, x20x, x485x, x478x}, x247x);
	defparam lut_3382.LUT_SIZE = 5;
	defparam lut_3382.mask = 32'h0fff0357;

	lut_sub lut_3385 ({sk[723], x24x, x18x, x563x, x567x}, x393x);
	defparam lut_3385.LUT_SIZE = 5;
	defparam lut_3385.mask = 32'h0fff0357;

	lut_sub lut_3388 ({sk[724], i_9_, i_7_, i_8_, i_6_, n_n195, n_n500}, x14943x);
	defparam lut_3388.LUT_SIZE = 7;
	defparam lut_3388.mask = 128'h777f777f777f777f0101000001010001;

	lut_sub lut_3394 ({sk[725], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x589x);
	defparam lut_3394.LUT_SIZE = 7;
	defparam lut_3394.mask = 128'h777f777f777f777f0002000000000000;

	lut_sub lut_3396 ({sk[726], x24x, x18x, x586x, x20x, x590x}, x14793x);
	defparam lut_3396.LUT_SIZE = 6;
	defparam lut_3396.mask = 64'h77ff77ff111f555f;

	lut_sub lut_3400 ({sk[727], i_9_, n_n526, n_n482, x510x, n_n195, x23x}, x14794x);
	defparam lut_3400.LUT_SIZE = 7;
	defparam lut_3400.mask = 128'h777f777f777f777f0011003303130333;

	lut_sub lut_3405 ({sk[728], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x527x);
	defparam lut_3405.LUT_SIZE = 7;
	defparam lut_3405.mask = 128'h777f777f777f777f0000080000000000;

	lut_sub lut_3407 ({sk[729], x538x, x19x, x23x, x529x, x534x, x527x}, x14807x);
	defparam lut_3407.LUT_SIZE = 7;
	defparam lut_3407.mask = 128'h777f777f777f777f00335f7f0033ffff;

	lut_sub lut_3412 ({sk[730], x19x, x21x, x584x, x599x}, x14801x);
	defparam lut_3412.LUT_SIZE = 5;
	defparam lut_3412.mask = 32'h0fff0537;

	lut_sub lut_3415 ({sk[731], x19x, x492x, x482x, x475x}, x14802x);
	defparam lut_3415.LUT_SIZE = 5;
	defparam lut_3415.mask = 32'h0fff007f;

	lut_sub lut_3419 ({sk[732], x15x, x23x, x487x, x569x, x579x, n_n5278}, x22135x);
	defparam lut_3419.LUT_SIZE = 7;
	defparam lut_3419.mask = 128'h777f777f777f777faaaa8888a0008000;

	lut_sub lut_3424 ({sk[733], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x531x);
	defparam lut_3424.LUT_SIZE = 7;
	defparam lut_3424.mask = 128'h777f777f777f777f0200000000000000;

	lut_sub lut_3426 ({sk[734], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x553x);
	defparam lut_3426.LUT_SIZE = 7;
	defparam lut_3426.mask = 128'h777f777f777f777f0000000000000008;

	lut_sub lut_3428 ({sk[735], x18x, x23x, x518x, x567x, x531x, x553x}, x14813x);
	defparam lut_3428.LUT_SIZE = 7;
	defparam lut_3428.mask = 128'h777f777f777f777f00007f7f00ff7fff;

	lut_sub lut_3433 ({sk[736], x22x, x21x, x17x, x585x, x576x, x548x}, x14820x);
	defparam lut_3433.LUT_SIZE = 7;
	defparam lut_3433.mask = 128'h777f777f777f777f005f337f337f337f;

	lut_sub lut_3438 ({sk[737], x22x, x17x, x512x, x503x}, x31x);
	defparam lut_3438.LUT_SIZE = 5;
	defparam lut_3438.mask = 32'h0fff0537;

	lut_sub lut_3441 ({sk[738], x17x, x20x, x587x, x576x}, x353x);
	defparam lut_3441.LUT_SIZE = 5;
	defparam lut_3441.mask = 32'h0fff0537;

	lut_sub lut_3444 ({sk[739], i_9_, i_7_, i_8_, i_6_, x540x}, n_n4453);
	defparam lut_3444.LUT_SIZE = 6;
	defparam lut_3444.mask = 64'h77ff77ff04000000;

	lut_sub lut_3446 ({sk[740], x22x, x11x, x24x, x583x, x547x, x543x}, x14845x);
	defparam lut_3446.LUT_SIZE = 7;
	defparam lut_3446.mask = 128'h777f777f777f777f003355770f3f5f7f;

	lut_sub lut_3450 ({sk[741], x15x, x24x, x20x, x583x, x543x, x523x}, x14846x);
	defparam lut_3450.LUT_SIZE = 7;
	defparam lut_3450.mask = 128'h777f777f777f777f00330f3f5f7f5f7f;

	lut_sub lut_3455 ({sk[742], x13x, x539x, x10x, x527x, x14845x, x14846x}, x14848x);
	defparam lut_3455.LUT_SIZE = 7;
	defparam lut_3455.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_3460 ({sk[743], x15x, x10x, x24x, x23x, x561x, x574x}, x14833x);
	defparam lut_3460.LUT_SIZE = 7;
	defparam lut_3460.mask = 128'h777f777f777f777f0333577733337777;

	lut_sub lut_3465 ({sk[744], x13x, x544x, x11x, x581x, x585x, x556x}, x14839x);
	defparam lut_3465.LUT_SIZE = 7;
	defparam lut_3465.mask = 128'h777f777f777f777f000000ff7f7f7fff;

	lut_sub lut_3470 ({sk[745], x15x, x13x, x574x, x543x}, x14837x);
	defparam lut_3470.LUT_SIZE = 5;
	defparam lut_3470.mask = 32'h0fff0357;

	lut_sub lut_3473 ({sk[746], x25x, x13x, x544x, x24x, x480x, x476x}, x14838x);
	defparam lut_3473.LUT_SIZE = 7;
	defparam lut_3473.mask = 128'h777f777f777f777f0505373705ff37ff;

	lut_sub lut_3477 ({sk[747], x10x, x20x, x561x, x564x, x491x, x396x}, x22130x);
	defparam lut_3477.LUT_SIZE = 7;
	defparam lut_3477.mask = 128'h777f777f777f777faaaaaa0080808000;

	lut_sub lut_3482 ({sk[748], x14833x, x14839x, x14837x, x14838x, x22130x}, x14849x);
	defparam lut_3482.LUT_SIZE = 6;
	defparam lut_3482.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_3488 ({sk[749], i_9_, x492x, n_n524, n_n325, n_n491, x511x}, x14868x);
	defparam lut_3488.LUT_SIZE = 7;
	defparam lut_3488.mask = 128'h777f777f777f777f0057005700030f0f;

	lut_sub lut_3493 ({sk[750], x14x, x17x, x557x, x580x, x503x, x549x}, x22304x);
	defparam lut_3493.LUT_SIZE = 7;
	defparam lut_3493.mask = 128'h777f777f777f777fffffaaaac0008000;

	lut_sub lut_3498 ({sk[751], x20x, x511x, x14868x, x22304x}, x14870x);
	defparam lut_3498.LUT_SIZE = 5;
	defparam lut_3498.mask = 32'h0fffbbbf;

	lut_sub lut_3502 ({sk[752], x16x, x21x, x500x, x20x, x557x, x498x}, x14876x);
	defparam lut_3502.LUT_SIZE = 7;
	defparam lut_3502.mask = 128'h777f777f777f777f050555ff373777ff;

	lut_sub lut_3507 ({sk[753], x16x, x501x, x545x, x20x, x482x, x535x}, x14882x);
	defparam lut_3507.LUT_SIZE = 7;
	defparam lut_3507.mask = 128'h777f777f777f777f00000f0f77ff7fff;

	lut_sub lut_3512 ({sk[754], i_9_, i_1_, i_2_, i_0_, x550x, x548x}, x234x);
	defparam lut_3512.LUT_SIZE = 7;
	defparam lut_3512.mask = 128'h777f777f777f777f0000000000000700;

	lut_sub lut_3515 ({sk[755], i_9_, i_7_, i_8_, i_6_, x540x}, n_n4447);
	defparam lut_3515.LUT_SIZE = 6;
	defparam lut_3515.mask = 64'h77ff77ff10000000;

	lut_sub lut_3517 ({sk[756], x16x, x11x, x503x, x495x}, x327x);
	defparam lut_3517.LUT_SIZE = 5;
	defparam lut_3517.mask = 32'h0fff0537;

	lut_sub lut_3520 ({sk[757], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x524x);
	defparam lut_3520.LUT_SIZE = 7;
	defparam lut_3520.mask = 128'h777f777f777f777f0800000000000000;

	lut_sub lut_3522 ({sk[758], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x541x);
	defparam lut_3522.LUT_SIZE = 7;
	defparam lut_3522.mask = 128'h777f777f777f777f0000040000000000;

	lut_sub lut_3524 ({sk[759], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x599x);
	defparam lut_3524.LUT_SIZE = 7;
	defparam lut_3524.mask = 128'h777f777f777f777f0000008000000000;

	lut_sub lut_3526 ({sk[760], x492x, x21x, x13x, x542x}, x130x);
	defparam lut_3526.LUT_SIZE = 5;
	defparam lut_3526.mask = 32'h0fff0537;

	lut_sub lut_3529 ({sk[761], x492x, x21x, x13x, x519x, x542x}, n_n4247);
	defparam lut_3529.LUT_SIZE = 6;
	defparam lut_3529.mask = 64'h77ff77ff03570f5f;

	lut_sub lut_3533 ({sk[762], i_9_, n_n482, n_n390, x570x, n_n530, x587x}, x16627x);
	defparam lut_3533.LUT_SIZE = 7;
	defparam lut_3533.mask = 128'h777f777f777f777f00000033005f007f;

	lut_sub lut_3538 ({sk[763], i_9_, i_1_, i_2_, i_0_, x550x}, n_n4952);
	defparam lut_3538.LUT_SIZE = 6;
	defparam lut_3538.mask = 64'h77ff77ff00000040;

	lut_sub lut_3540 ({sk[764], i_9_, n_n260, n_n520, x18x, x550x, n_n464}, n_n3803);
	defparam lut_3540.LUT_SIZE = 7;
	defparam lut_3540.mask = 128'h777f777f777f777f0303035703030357;

	lut_sub lut_3544 ({sk[765], x15x, x11x, x17x, x524x, x531x}, n_n3805);
	defparam lut_3544.LUT_SIZE = 6;
	defparam lut_3544.mask = 64'h77ff77ff03575757;

	lut_sub lut_3548 ({sk[766], x22x, x17x, x20x, x516x, x531x}, x16327x);
	defparam lut_3548.LUT_SIZE = 6;
	defparam lut_3548.mask = 64'h77ff77ff05375577;

	lut_sub lut_3552 ({sk[767], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x487x);
	defparam lut_3552.LUT_SIZE = 7;
	defparam lut_3552.mask = 128'h777f777f777f777f0000000000008000;

	lut_sub lut_3554 ({sk[768], x19x, x11x, x477x, x487x}, x318x);
	defparam lut_3554.LUT_SIZE = 5;
	defparam lut_3554.mask = 32'h0fff0537;

	lut_sub lut_3557 ({sk[769], x19x, x482x, x23x, x599x}, x319x);
	defparam lut_3557.LUT_SIZE = 5;
	defparam lut_3557.mask = 32'h0fff111f;

	lut_sub lut_3560 ({sk[770], i_9_, i_7_, i_8_, i_6_, x540x}, n_n4441);
	defparam lut_3560.LUT_SIZE = 6;
	defparam lut_3560.mask = 64'h77ff77ff00010000;

	lut_sub lut_3562 ({sk[771], i_9_, i_7_, i_8_, i_6_, n_n455, n_n535}, n_n2261);
	defparam lut_3562.LUT_SIZE = 7;
	defparam lut_3562.mask = 128'h777f777f777f777f0101101100011110;

	lut_sub lut_3572 ({sk[772], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x546x);
	defparam lut_3572.LUT_SIZE = 7;
	defparam lut_3572.mask = 128'h777f777f777f777f0010000000000000;

	lut_sub lut_3574 ({sk[773], x13x, x490x, x20x, x540x, x546x}, n_n3889);
	defparam lut_3574.LUT_SIZE = 6;
	defparam lut_3574.mask = 64'h77ff77ff030357ff;

	lut_sub lut_3578 ({sk[774], i_9_, i_1_, i_2_, i_0_, x482x}, n_n4472);
	defparam lut_3578.LUT_SIZE = 6;
	defparam lut_3578.mask = 64'h77ff77ff00000010;

	lut_sub lut_3580 ({sk[775], x13x, x544x, x482x, x23x}, x413x);
	defparam lut_3580.LUT_SIZE = 5;
	defparam lut_3580.mask = 32'h0fff0537;

	lut_sub lut_3583 ({sk[776], x13x, x23x, x594x, x540x}, x14515x);
	defparam lut_3583.LUT_SIZE = 5;
	defparam lut_3583.mask = 32'h0fff0537;

	lut_sub lut_3586 ({sk[777], x25x, x13x, x544x, x559x}, x14516x);
	defparam lut_3586.LUT_SIZE = 5;
	defparam lut_3586.mask = 32'h0fff0537;

	lut_sub lut_3589 ({sk[778], x13x, x544x, x24x, x581x}, x16564x);
	defparam lut_3589.LUT_SIZE = 5;
	defparam lut_3589.mask = 32'h0fff0357;

	lut_sub lut_3592 ({sk[779], x25x, x13x, x585x, x476x}, x16565x);
	defparam lut_3592.LUT_SIZE = 5;
	defparam lut_3592.mask = 32'h0fff0357;

	lut_sub lut_3595 ({sk[780], i_9_, i_1_, i_2_, i_0_, x560x}, n_n4886);
	defparam lut_3595.LUT_SIZE = 6;
	defparam lut_3595.mask = 64'h77ff77ff00000004;

	lut_sub lut_3597 ({sk[781], i_9_, n_n260, n_n520, x20x, n_n500, x574x}, x16331x);
	defparam lut_3597.LUT_SIZE = 7;
	defparam lut_3597.mask = 128'h777f777f777f777f0000033300005777;

	lut_sub lut_3602 ({sk[782], i_9_, n_n518, x474x, n_n260, n_n522, x472x}, x16335x);
	defparam lut_3602.LUT_SIZE = 7;
	defparam lut_3602.mask = 128'h777f777f777f777f00000303050f070f;

	lut_sub lut_3607 ({sk[783], x15x, x17x, x478x, x564x, x566x}, x16339x);
	defparam lut_3607.LUT_SIZE = 6;
	defparam lut_3607.mask = 64'h77ff77ff003f557f;

	lut_sub lut_3611 ({sk[784], i_9_, i_7_, i_8_, i_6_, n_n260, n_n500}, x16340x);
	defparam lut_3611.LUT_SIZE = 7;
	defparam lut_3611.mask = 128'h777f777f777f777f0000011101000000;

	lut_sub lut_3616 ({sk[785], x17x, x20x, x484x, x536x, x16339x, x16340x}, x16342x);
	defparam lut_3616.LUT_SIZE = 7;
	defparam lut_3616.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_3621 ({sk[786], x11x, x17x, x573x, x576x}, x16330x);
	defparam lut_3621.LUT_SIZE = 5;
	defparam lut_3621.mask = 32'h0fff0357;

	lut_sub lut_3624 ({sk[787], x24x, x17x, x484x, x475x}, x16333x);
	defparam lut_3624.LUT_SIZE = 5;
	defparam lut_3624.mask = 32'h0fff0537;

	lut_sub lut_3627 ({sk[788], x15x, x521x, x17x, x484x, x477x}, x16334x);
	defparam lut_3627.LUT_SIZE = 6;
	defparam lut_3627.mask = 64'h77ff77ff050f373f;

	lut_sub lut_3631 ({sk[789], n_n3451, x16331x, x16335x, x16330x, x16333x, x16334x}, x16343x);
	defparam lut_3631.LUT_SIZE = 7;
	defparam lut_3631.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_3638 ({sk[790], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x528x);
	defparam lut_3638.LUT_SIZE = 7;
	defparam lut_3638.mask = 128'h777f777f777f777f0000000008000000;

	lut_sub lut_3640 ({sk[791], x19x, x24x, x534x, x527x, x528x}, n_n2274);
	defparam lut_3640.LUT_SIZE = 6;
	defparam lut_3640.mask = 64'h77ff77ff000f777f;

	lut_sub lut_3644 ({sk[792], i_9_, i_7_, i_8_, i_6_, x534x}, n_n5329);
	defparam lut_3644.LUT_SIZE = 6;
	defparam lut_3644.mask = 64'h77ff77ff00040000;

	lut_sub lut_3646 ({sk[793], i_9_, i_1_, i_2_, i_0_, x506x, x529x}, x116x);
	defparam lut_3646.LUT_SIZE = 7;
	defparam lut_3646.mask = 128'h777f777f777f777f0000000070000000;

	lut_sub lut_3649 ({sk[794], i_9_, i_1_, i_2_, i_0_, x509x, x580x}, x12968x);
	defparam lut_3649.LUT_SIZE = 7;
	defparam lut_3649.mask = 128'h777f777f777f777f0000000070000000;

	lut_sub lut_3652 ({sk[795], i_9_, n_n482, x510x, x23x, n_n65, x63x}, x12969x);
	defparam lut_3652.LUT_SIZE = 7;
	defparam lut_3652.mask = 128'h777f777f777f777f5555575755775777;

	lut_sub lut_3656 ({sk[796], i_9_, n_n524, n_n464, n_n65, x116x}, x16656x);
	defparam lut_3656.LUT_SIZE = 6;
	defparam lut_3656.mask = 64'h77ff77ff55575557;

	lut_sub lut_3660 ({sk[797], i_9_, i_7_, i_8_, i_6_, n_n464, n_n65}, x16658x);
	defparam lut_3660.LUT_SIZE = 7;
	defparam lut_3660.mask = 128'h777f777f777f777f0001001001100000;

	lut_sub lut_3665 ({sk[798], x25x, x515x, x11x, x24x, n_n5310, x534x}, x22067x);
	defparam lut_3665.LUT_SIZE = 7;
	defparam lut_3665.mask = 128'h777f777f777f777fccccc00088888000;

	lut_sub lut_3670 ({sk[799], n_n2274, x16656x, x16658x, x22067x}, x16662x);
	defparam lut_3670.LUT_SIZE = 5;
	defparam lut_3670.mask = 32'h0fffbfff;

	lut_sub lut_3675 ({sk[800], i_9_, i_7_, i_8_, i_6_, n_n473, n_n325}, x16349x);
	defparam lut_3675.LUT_SIZE = 7;
	defparam lut_3675.mask = 128'h777f777f777f777f0000010100100100;

	lut_sub lut_3680 ({sk[801], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x530x);
	defparam lut_3680.LUT_SIZE = 7;
	defparam lut_3680.mask = 128'h777f777f777f777f4000000000000000;

	lut_sub lut_3682 ({sk[802], i_9_, i_7_, i_8_, i_6_, n_n325, n_n464}, x16363x);
	defparam lut_3682.LUT_SIZE = 7;
	defparam lut_3682.mask = 128'h777f777f777f777f0010100000101100;

	lut_sub lut_3688 ({sk[803], x14x, x17x, x550x, x506x, x525x}, x22288x);
	defparam lut_3688.LUT_SIZE = 6;
	defparam lut_3688.mask = 64'h77ff77fffff08880;

	lut_sub lut_3693 ({sk[804], x23x, x530x, x16363x, x22288x}, x16364x);
	defparam lut_3693.LUT_SIZE = 5;
	defparam lut_3693.mask = 32'h0fffbbbf;

	lut_sub lut_3697 ({sk[805], x17x, x552x, x23x, x594x}, x177x);
	defparam lut_3697.LUT_SIZE = 5;
	defparam lut_3697.mask = 32'h0fff0357;

	lut_sub lut_3700 ({sk[806], i_9_, i_7_, i_8_, i_6_, n_n260, n_n535}, n_n2230);
	defparam lut_3700.LUT_SIZE = 7;
	defparam lut_3700.mask = 128'h777f777f777f777f0101100101011110;

	lut_sub lut_3710 ({sk[807], x15x, x17x, x596x, x585x}, x176x);
	defparam lut_3710.LUT_SIZE = 5;
	defparam lut_3710.mask = 32'h0fff0537;

	lut_sub lut_3713 ({sk[808], x24x, x552x, x20x, x596x, n_n4846, x372x}, x22079x);
	defparam lut_3713.LUT_SIZE = 7;
	defparam lut_3713.mask = 128'h777f777f777f777f8888880080808000;

	lut_sub lut_3718 ({sk[809], x177x, n_n2230, x176x, x22079x}, x16365x);
	defparam lut_3718.LUT_SIZE = 5;
	defparam lut_3718.mask = 32'h0fffbfff;

	lut_sub lut_3723 ({sk[810], i_9_, i_7_, i_8_, i_6_, n_n325, n_n491}, n_n2234);
	defparam lut_3723.LUT_SIZE = 7;
	defparam lut_3723.mask = 128'h777f777f777f777f0111111001001010;

	lut_sub lut_3733 ({sk[811], x14x, x587x, x16372x, x22306x}, x16374x);
	defparam lut_3733.LUT_SIZE = 5;
	defparam lut_3733.mask = 32'h0fffbbbf;

	lut_sub lut_3737 ({sk[812], x14x, x508x, x16349x, n_n2234, n_n4797, x16348x}, x16375x);
	defparam lut_3737.LUT_SIZE = 7;
	defparam lut_3737.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_3743 ({sk[813], i_9_, i_7_, i_8_, i_6_, n_n325, n_n500}, x16382x);
	defparam lut_3743.LUT_SIZE = 7;
	defparam lut_3743.mask = 128'h777f777f777f777f0001011000010000;

	lut_sub lut_3748 ({sk[814], i_9_, i_7_, i_8_, i_6_, n_n509, n_n325}, n_n2237);
	defparam lut_3748.LUT_SIZE = 7;
	defparam lut_3748.mask = 128'h777f777f777f777f0111110001011010;

	lut_sub lut_3758 ({sk[815], i_9_, i_7_, i_8_, i_6_, x565x}, n_n4759);
	defparam lut_3758.LUT_SIZE = 6;
	defparam lut_3758.mask = 64'h77ff77ff40000000;

	lut_sub lut_3760 ({sk[816], i_9_, i_1_, i_2_, i_0_, x535x}, n_n4704);
	defparam lut_3760.LUT_SIZE = 6;
	defparam lut_3760.mask = 64'h77ff77ff00001000;

	lut_sub lut_3762 ({sk[817], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x551x);
	defparam lut_3762.LUT_SIZE = 7;
	defparam lut_3762.mask = 128'h777f777f777f777f0000000000000040;

	lut_sub lut_3764 ({sk[818], i_9_, i_7_, i_8_, i_6_, n_n325, n_n535}, x16396x);
	defparam lut_3764.LUT_SIZE = 7;
	defparam lut_3764.mask = 128'h777f777f777f777f0010100001000100;

	lut_sub lut_3769 ({sk[819], x22x, x11x, n_n4216, n_n4704, x551x, x16396x}, x16399x);
	defparam lut_3769.LUT_SIZE = 7;
	defparam lut_3769.mask = 128'h777f777f777f777f5fff7fff7fff7fff;

	lut_sub lut_3775 ({sk[820], x14x, x550x, x23x, x526x}, x86x);
	defparam lut_3775.LUT_SIZE = 5;
	defparam lut_3775.mask = 32'h0fff111f;

	lut_sub lut_3778 ({sk[821], x24x, x14x, x595x, x593x}, x173x);
	defparam lut_3778.LUT_SIZE = 5;
	defparam lut_3778.mask = 32'h0fff0537;

	lut_sub lut_3781 ({sk[822], x25x, x483x, x14x, x20x, x581x, x595x}, x16388x);
	defparam lut_3781.LUT_SIZE = 7;
	defparam lut_3781.mask = 128'h777f777f777f777f053705370537ffff;

	lut_sub lut_3785 ({sk[823], i_9_, n_n325, n_n535, x23x, x594x, x442x}, x16395x);
	defparam lut_3785.LUT_SIZE = 7;
	defparam lut_3785.mask = 128'h777f777f777f777f5555555f5555777f;

	lut_sub lut_3789 ({sk[824], x14x, x482x, x481x, x494x, n_n4727, x39x}, x22078x);
	defparam lut_3789.LUT_SIZE = 7;
	defparam lut_3789.mask = 128'h777f777f777f777f8888888880000000;

	lut_sub lut_3792 ({sk[825], x86x, x173x, x16388x, x16395x, x22078x}, x16400x);
	defparam lut_3792.LUT_SIZE = 6;
	defparam lut_3792.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_3798 ({sk[826], x10x, x24x, x507x, x510x, x23x, x582x}, n_n1764);
	defparam lut_3798.LUT_SIZE = 7;
	defparam lut_3798.mask = 128'h777f777f777f777f111111ff1f1f1fff;

	lut_sub lut_3802 ({sk[827], i_9_, i_7_, i_8_, i_6_, n_n390, n_n464}, x16413x);
	defparam lut_3802.LUT_SIZE = 7;
	defparam lut_3802.mask = 128'h777f777f777f777f0010101010101000;

	lut_sub lut_3809 ({sk[828], x10x, x522x, x524x, n_n1764, x16413x}, x16415x);
	defparam lut_3809.LUT_SIZE = 6;
	defparam lut_3809.mask = 64'h77ff77ff77777fff;

	lut_sub lut_3814 ({sk[829], i_9_, i_7_, i_8_, i_6_, x507x}, n_n4679);
	defparam lut_3814.LUT_SIZE = 6;
	defparam lut_3814.mask = 64'h77ff77ff40000000;

	lut_sub lut_3816 ({sk[830], x10x, x24x, x580x, x520x, x493x, x526x}, x16411x);
	defparam lut_3816.LUT_SIZE = 7;
	defparam lut_3816.mask = 128'h777f777f777f777f000055553fff7fff;

	lut_sub lut_3821 ({sk[831], x22x, x10x, x507x, x20x, x506x, x488x}, x22076x);
	defparam lut_3821.LUT_SIZE = 7;
	defparam lut_3821.mask = 128'h777f777f777f777ffff08880ff008800;

	lut_sub lut_3826 ({sk[832], x22x, x10x, x582x, x528x, x338x, x431x}, x22077x);
	defparam lut_3826.LUT_SIZE = 7;
	defparam lut_3826.mask = 128'h777f777f777f777f8888808088008000;

	lut_sub lut_3831 ({sk[833], x25x, x526x, n_n4679, x16411x, x22076x, x22077x}, x16416x);
	defparam lut_3831.LUT_SIZE = 7;
	defparam lut_3831.mask = 128'h777f777f777f777fefffefffefffffff;

	lut_sub lut_3837 ({sk[834], x25x, x14x, x573x, x575x}, x69x);
	defparam lut_3837.LUT_SIZE = 5;
	defparam lut_3837.mask = 32'h0fff0357;

	lut_sub lut_3840 ({sk[835], x14x, x560x, x69x, x16419x, x16421x}, x16423x);
	defparam lut_3840.LUT_SIZE = 6;
	defparam lut_3840.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_3845 ({sk[836], x11x, x565x, x16382x, n_n2237, x22290x}, x16424x);
	defparam lut_3845.LUT_SIZE = 6;
	defparam lut_3845.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_3850 ({sk[837], i_9_, i_7_, i_8_, i_6_, x553x}, n_n4959);
	defparam lut_3850.LUT_SIZE = 6;
	defparam lut_3850.mask = 64'h77ff77ff10000000;

	lut_sub lut_3852 ({sk[838], x18x, x597x, x23x, x581x}, x251x);
	defparam lut_3852.LUT_SIZE = 5;
	defparam lut_3852.mask = 32'h0fff0357;

	lut_sub lut_3855 ({sk[839], x24x, x18x, x485x, x480x}, x133x);
	defparam lut_3855.LUT_SIZE = 5;
	defparam lut_3855.mask = 32'h0fff0537;

	lut_sub lut_3858 ({sk[840], x21x, x18x, x597x, x477x}, x16437x);
	defparam lut_3858.LUT_SIZE = 5;
	defparam lut_3858.mask = 32'h0fff0537;

	lut_sub lut_3861 ({sk[841], x25x, x18x, x482x, x485x}, x16438x);
	defparam lut_3861.LUT_SIZE = 5;
	defparam lut_3861.mask = 32'h0fff0357;

	lut_sub lut_3864 ({sk[842], x18x, x481x, x251x, x133x, x16437x, x16438x}, x16442x);
	defparam lut_3864.LUT_SIZE = 7;
	defparam lut_3864.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_3870 ({sk[843], i_9_, n_n509, n_n520, n_n195, x393x}, x16430x);
	defparam lut_3870.LUT_SIZE = 6;
	defparam lut_3870.mask = 64'h77ff77ff55575557;

	lut_sub lut_3874 ({sk[844], x18x, x23x, x518x, x491x, x573x, x567x}, x16435x);
	defparam lut_3874.LUT_SIZE = 7;
	defparam lut_3874.mask = 128'h777f777f777f777f000055553fff7fff;

	lut_sub lut_3879 ({sk[845], x25x, x474x, x18x, x567x, x562x, x136x}, x22075x);
	defparam lut_3879.LUT_SIZE = 7;
	defparam lut_3879.mask = 128'h777f777f777f777faa88aa00a080a000;

	lut_sub lut_3884 ({sk[846], x22x, x18x, x20x, x574x, x567x, x297x}, x22335x);
	defparam lut_3884.LUT_SIZE = 7;
	defparam lut_3884.mask = 128'h777f777f777f777faa88a08088888080;

	lut_sub lut_3889 ({sk[847], x16430x, x16435x, x22075x, x22335x}, x16443x);
	defparam lut_3889.LUT_SIZE = 5;
	defparam lut_3889.mask = 32'h0fffefff;

	lut_sub lut_3894 ({sk[848], x22x, x17x, x520x, x589x}, x351x);
	defparam lut_3894.LUT_SIZE = 5;
	defparam lut_3894.mask = 32'h0fff0357;

	lut_sub lut_3897 ({sk[849], x17x, x20x, x580x, x589x}, x369x);
	defparam lut_3897.LUT_SIZE = 5;
	defparam lut_3897.mask = 32'h0fff0537;

	lut_sub lut_3900 ({sk[850], x25x, x24x, x23x, x512x, n_n4920, x589x}, x22074x);
	defparam lut_3900.LUT_SIZE = 7;
	defparam lut_3900.mask = 128'h777f777f777f777fcc88c080c080c080;

	lut_sub lut_3905 ({sk[851], x21x, x589x, x351x, x369x, x22074x}, x16456x);
	defparam lut_3905.LUT_SIZE = 6;
	defparam lut_3905.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_3910 ({sk[852], i_9_, n_n528, n_n473, n_n260, x508x, x132x}, x249x);
	defparam lut_3910.LUT_SIZE = 7;
	defparam lut_3910.mask = 128'h777f777f777f777f5555555f57575757;

	lut_sub lut_3914 ({sk[853], x492x, x21x, x17x, x576x}, x226x);
	defparam lut_3914.LUT_SIZE = 5;
	defparam lut_3914.mask = 32'h0fff0537;

	lut_sub lut_3917 ({sk[854], i_9_, i_7_, i_8_, i_6_, n_n260, n_n491}, x16450x);
	defparam lut_3917.LUT_SIZE = 7;
	defparam lut_3917.mask = 128'h777f777f777f777f1010001000001010;

	lut_sub lut_3923 ({sk[855], i_9_, i_7_, i_8_, i_6_, x589x}, x16447x);
	defparam lut_3923.LUT_SIZE = 6;
	defparam lut_3923.mask = 64'h77ff77ff11000000;

	lut_sub lut_3926 ({sk[856], x25x, x20x, x23x, x512x, x31x, x531x}, x22073x);
	defparam lut_3926.LUT_SIZE = 7;
	defparam lut_3926.mask = 128'h777f777f777f777fccc0c0c088808080;

	lut_sub lut_3931 ({sk[857], x249x, x226x, x16450x, x16447x, x22073x}, x16457x);
	defparam lut_3931.LUT_SIZE = 6;
	defparam lut_3931.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_3937 ({sk[858], x25x, x18x, x597x, x594x}, x341x);
	defparam lut_3937.LUT_SIZE = 5;
	defparam lut_3937.mask = 32'h0fff0537;

	lut_sub lut_3940 ({sk[859], i_9_, i_7_, i_8_, i_6_, x553x}, x362x);
	defparam lut_3940.LUT_SIZE = 6;
	defparam lut_3940.mask = 64'h77ff77ff44000000;

	lut_sub lut_3943 ({sk[860], x22x, x521x, x539x, x18x, x597x, x546x}, x22285x);
	defparam lut_3943.LUT_SIZE = 7;
	defparam lut_3943.mask = 128'h777f777f777f777ffaf0f0f0c8c0c0c0;

	lut_sub lut_3948 ({sk[861], x18x, x585x, x341x, x362x, x22285x}, n_n2220);
	defparam lut_3948.LUT_SIZE = 6;
	defparam lut_3948.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_3953 ({sk[862], x25x, x24x, x18x, x549x, x553x}, n_n3802);
	defparam lut_3953.LUT_SIZE = 6;
	defparam lut_3953.mask = 64'h77ff77ff03575757;

	lut_sub lut_3957 ({sk[863], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x493x);
	defparam lut_3957.LUT_SIZE = 7;
	defparam lut_3957.mask = 128'h777f777f777f777f0000400000000000;

	lut_sub lut_3959 ({sk[864], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x543x);
	defparam lut_3959.LUT_SIZE = 7;
	defparam lut_3959.mask = 128'h777f777f777f777f0004000000000000;

	lut_sub lut_3961 ({sk[865], i_9_, i_7_, i_8_, i_6_, x504x}, n_n4539);
	defparam lut_3961.LUT_SIZE = 6;
	defparam lut_3961.mask = 64'h77ff77ff00100000;

	lut_sub lut_3963 ({sk[866], i_9_, i_1_, i_2_, i_0_, x503x}, n_n4544);
	defparam lut_3963.LUT_SIZE = 6;
	defparam lut_3963.mask = 64'h77ff77ff00000010;

	lut_sub lut_3965 ({sk[867], i_9_, i_1_, i_2_, i_0_, x522x}, n_n4560);
	defparam lut_3965.LUT_SIZE = 6;
	defparam lut_3965.mask = 64'h77ff77ff00000010;

	lut_sub lut_3967 ({sk[868], x11x, x14x, x490x, x472x, x595x, x546x}, x16503x);
	defparam lut_3967.LUT_SIZE = 7;
	defparam lut_3967.mask = 128'h777f777f777f777f00005fff33337fff;

	lut_sub lut_3972 ({sk[869], x492x, x11x, x14x, x572x, x526x}, x16502x);
	defparam lut_3972.LUT_SIZE = 6;
	defparam lut_3972.mask = 64'h77ff77ff03570f5f;

	lut_sub lut_3976 ({sk[870], x24x, x14x, x517x, x16503x, x551x, x16502x}, n_n2098);
	defparam lut_3976.LUT_SIZE = 7;
	defparam lut_3976.mask = 128'h777f777f777f777f5f5f5fff7f7f7fff;

	lut_sub lut_3981 ({sk[871], x11x, x10x, x507x, x503x}, x193x);
	defparam lut_3981.LUT_SIZE = 5;
	defparam lut_3981.mask = 32'h0fff0537;

	lut_sub lut_3984 ({sk[872], i_9_, i_7_, i_8_, i_6_, x507x, x582x}, x16506x);
	defparam lut_3984.LUT_SIZE = 7;
	defparam lut_3984.mask = 128'h777f777f777f777f0000700000000000;

	lut_sub lut_3987 ({sk[873], x538x, x10x, x23x, x571x, x502x, n_n4661}, x22059x);
	defparam lut_3987.LUT_SIZE = 7;
	defparam lut_3987.mask = 128'h777f777f777f777faaa08880aaa00000;

	lut_sub lut_3992 ({sk[874], x15x, x526x, x193x, x16506x, x22059x}, n_n2099);
	defparam lut_3992.LUT_SIZE = 6;
	defparam lut_3992.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_3997 ({sk[875], i_9_, i_1_, i_2_, i_0_, x550x}, n_n4824);
	defparam lut_3997.LUT_SIZE = 6;
	defparam lut_3997.mask = 64'h77ff77ff00000004;

	lut_sub lut_3999 ({sk[876], i_9_, i_1_, i_2_, i_0_, x528x}, n_n4938);
	defparam lut_3999.LUT_SIZE = 6;
	defparam lut_3999.mask = 64'h77ff77ff00000004;

	lut_sub lut_4001 ({sk[877], x15x, x24x, x558x, x18x, x590x}, n_n1570);
	defparam lut_4001.LUT_SIZE = 6;
	defparam lut_4001.mask = 64'h77ff77ff03575757;

	lut_sub lut_4005 ({sk[878], i_9_, i_7_, i_8_, i_6_, x590x}, n_n5043);
	defparam lut_4005.LUT_SIZE = 6;
	defparam lut_4005.mask = 64'h77ff77ff00400000;

	lut_sub lut_4007 ({sk[879], i_9_, i_1_, i_2_, i_0_, x580x}, n_n5302);
	defparam lut_4007.LUT_SIZE = 6;
	defparam lut_4007.mask = 64'h77ff77ff00004000;

	lut_sub lut_4009 ({sk[880], x24x, x510x, x17x, x557x, x589x, x525x}, x12089x);
	defparam lut_4009.LUT_SIZE = 7;
	defparam lut_4009.mask = 128'h777f777f777f777f005f00ff337f33ff;

	lut_sub lut_4014 ({sk[881], i_9_, i_7_, i_8_, i_6_, x568x}, n_n5131);
	defparam lut_4014.LUT_SIZE = 6;
	defparam lut_4014.mask = 64'h77ff77ff00100000;

	lut_sub lut_4016 ({sk[882], i_9_, i_1_, i_2_, i_0_, x489x}, n_n5204);
	defparam lut_4016.LUT_SIZE = 6;
	defparam lut_4016.mask = 64'h77ff77ff00000400;

	lut_sub lut_4018 ({sk[883], i_9_, n_n526, n_n130, x522x, n_n500, x525x}, x12096x);
	defparam lut_4018.LUT_SIZE = 7;
	defparam lut_4018.mask = 128'h777f777f777f777f00000033005f007f;

	lut_sub lut_4023 ({sk[884], i_9_, i_7_, i_8_, i_6_, x514x, x568x}, x12095x);
	defparam lut_4023.LUT_SIZE = 7;
	defparam lut_4023.mask = 128'h777f777f777f777f3000050500000000;

	lut_sub lut_4027 ({sk[885], x12x, x573x, x489x, x12096x, x12095x}, n_n1330);
	defparam lut_4027.LUT_SIZE = 6;
	defparam lut_4027.mask = 64'h77ff77ff77777fff;

	lut_sub lut_4032 ({sk[886], i_9_, i_7_, i_8_, i_6_, x486x}, n_n5113);
	defparam lut_4032.LUT_SIZE = 6;
	defparam lut_4032.mask = 64'h77ff77ff00010000;

	lut_sub lut_4034 ({sk[887], i_9_, i_7_, i_8_, i_6_, x554x}, n_n5081);
	defparam lut_4034.LUT_SIZE = 6;
	defparam lut_4034.mask = 64'h77ff77ff00010000;

	lut_sub lut_4036 ({sk[888], x18x, x23x, x513x, x528x}, x344x);
	defparam lut_4036.LUT_SIZE = 5;
	defparam lut_4036.mask = 32'h0fff0357;

	lut_sub lut_4039 ({sk[889], x12x, x472x, x481x, x594x, x480x, n_n5113}, x22222x);
	defparam lut_4039.LUT_SIZE = 7;
	defparam lut_4039.mask = 128'h777f777f777f777faaaaaaaa80000000;

	lut_sub lut_4042 ({sk[890], x25x, x22x, x554x, x344x, x22222x}, n_n1331);
	defparam lut_4042.LUT_SIZE = 6;
	defparam lut_4042.mask = 64'h77ff77ffbbbfbfbf;

	lut_sub lut_4047 ({sk[891], i_9_, i_1_, i_2_, i_0_, x539x}, n_n5232);
	defparam lut_4047.LUT_SIZE = 6;
	defparam lut_4047.mask = 64'h77ff77ff00004000;

	lut_sub lut_4049 ({sk[892], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x569x);
	defparam lut_4049.LUT_SIZE = 7;
	defparam lut_4049.mask = 128'h777f777f777f777f0000800000000000;

	lut_sub lut_4051 ({sk[893], i_9_, i_1_, i_2_, i_0_, x535x}, n_n5216);
	defparam lut_4051.LUT_SIZE = 6;
	defparam lut_4051.mask = 64'h77ff77ff00004000;

	lut_sub lut_4053 ({sk[894], x19x, x563x, x480x, x535x, x548x, x546x}, x12109x);
	defparam lut_4053.LUT_SIZE = 7;
	defparam lut_4053.mask = 128'h777f777f777f777f000000007fffffff;

	lut_sub lut_4059 ({sk[895], x19x, x539x, x23x, x573x, x487x}, x22259x);
	defparam lut_4059.LUT_SIZE = 6;
	defparam lut_4059.mask = 64'h77ff77fffafac800;

	lut_sub lut_4064 ({sk[896], x21x, x569x, x12109x, x22259x}, x12110x);
	defparam lut_4064.LUT_SIZE = 5;
	defparam lut_4064.mask = 32'h0fffbbbf;

	lut_sub lut_4068 ({sk[897], i_9_, i_1_, i_2_, i_0_, x482x}, n_n4344);
	defparam lut_4068.LUT_SIZE = 6;
	defparam lut_4068.mask = 64'h77ff77ff00000001;

	lut_sub lut_4070 ({sk[898], i_9_, i_7_, i_8_, i_6_, x499x}, n_n4391);
	defparam lut_4070.LUT_SIZE = 6;
	defparam lut_4070.mask = 64'h77ff77ff40000000;

	lut_sub lut_4072 ({sk[899], i_9_, i_7_, i_8_, i_6_, x479x}, n_n4611);
	defparam lut_4072.LUT_SIZE = 6;
	defparam lut_4072.mask = 64'h77ff77ff00400000;

	lut_sub lut_4074 ({sk[900], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x532x);
	defparam lut_4074.LUT_SIZE = 7;
	defparam lut_4074.mask = 128'h777f777f777f777f0800000000000000;

	lut_sub lut_4076 ({sk[901], i_9_, i_7_, i_8_, i_6_, x498x}, n_n4367);
	defparam lut_4076.LUT_SIZE = 6;
	defparam lut_4076.mask = 64'h77ff77ff10000000;

	lut_sub lut_4078 ({sk[902], i_9_, i_7_, i_8_, i_6_, x498x}, n_n4365);
	defparam lut_4078.LUT_SIZE = 6;
	defparam lut_4078.mask = 64'h77ff77ff01000000;

	lut_sub lut_4080 ({sk[903], x15x, x16x, x11x, x498x, x556x}, n_n1308);
	defparam lut_4080.LUT_SIZE = 6;
	defparam lut_4080.mask = 64'h77ff77ff03573377;

	lut_sub lut_4084 ({sk[904], x15x, x14x, x557x, x575x}, x165x);
	defparam lut_4084.LUT_SIZE = 5;
	defparam lut_4084.mask = 32'h0fff0357;

	lut_sub lut_4087 ({sk[905], i_9_, i_7_, i_8_, i_6_, n_n325, n_n491}, n_n1086);
	defparam lut_4087.LUT_SIZE = 7;
	defparam lut_4087.mask = 128'h777f777f777f777f0101101011111000;

	lut_sub lut_4097 ({sk[906], x538x, x11x, x17x, x589x}, x306x);
	defparam lut_4097.LUT_SIZE = 5;
	defparam lut_4097.mask = 32'h0fff0537;

	lut_sub lut_4100 ({sk[907], i_9_, i_7_, i_8_, i_6_, n_n482, n_n260}, n_n1075);
	defparam lut_4100.LUT_SIZE = 7;
	defparam lut_4100.mask = 128'h777f777f777f777f0100001100111111;

	lut_sub lut_4110 ({sk[908], i_9_, n_n526, n_n473, n_n195, n_n530, x580x}, x11993x);
	defparam lut_4110.LUT_SIZE = 7;
	defparam lut_4110.mask = 128'h777f777f777f777f0003000f0507050f;

	lut_sub lut_4116 ({sk[909], x509x, x24x, x14x, x511x}, x179x);
	defparam lut_4116.LUT_SIZE = 5;
	defparam lut_4116.mask = 32'h0fff0537;

	lut_sub lut_4119 ({sk[910], x25x, x509x, x24x, x14x, x511x}, n_n2003);
	defparam lut_4119.LUT_SIZE = 6;
	defparam lut_4119.mask = 64'h77ff77ff05375577;

	lut_sub lut_4123 ({sk[911], x25x, x14x, x503x, x505x, x530x, x528x}, x11756x);
	defparam lut_4123.LUT_SIZE = 7;
	defparam lut_4123.mask = 128'h777f777f777f777f00005fff33337fff;

	lut_sub lut_4128 ({sk[912], i_9_, i_7_, i_8_, i_6_, n_n473, n_n325}, x11757x);
	defparam lut_4128.LUT_SIZE = 7;
	defparam lut_4128.mask = 128'h777f777f777f777f1000100010101000;

	lut_sub lut_4134 ({sk[913], i_9_, i_7_, i_8_, i_6_, n_n325, n_n464}, n_n1082);
	defparam lut_4134.LUT_SIZE = 7;
	defparam lut_4134.mask = 128'h777f777f777f777f0110110011011010;

	lut_sub lut_4144 ({sk[914], i_9_, n_n482, n_n325, x23x, x580x}, x292x);
	defparam lut_4144.LUT_SIZE = 6;
	defparam lut_4144.mask = 64'h77ff77ff00030507;

	lut_sub lut_4147 ({sk[915], x21x, x510x, x14x, x588x}, x11763x);
	defparam lut_4147.LUT_SIZE = 5;
	defparam lut_4147.mask = 32'h0fff0357;

	lut_sub lut_4150 ({sk[916], i_9_, n_n482, n_n325, n_n522, x23x, x580x}, x11764x);
	defparam lut_4150.LUT_SIZE = 7;
	defparam lut_4150.mask = 128'h777f777f777f777f0000003f0055007f;

	lut_sub lut_4155 ({sk[917], i_9_, i_7_, i_8_, i_6_, x596x}, n_n4843);
	defparam lut_4155.LUT_SIZE = 6;
	defparam lut_4155.mask = 64'h77ff77ff00100000;

	lut_sub lut_4157 ({sk[918], i_9_, i_1_, i_2_, i_0_, x559x}, n_n4846);
	defparam lut_4157.LUT_SIZE = 6;
	defparam lut_4157.mask = 64'h77ff77ff00000004;

	lut_sub lut_4159 ({sk[919], x21x, x17x, x552x, x490x, x20x}, n_n3460);
	defparam lut_4159.LUT_SIZE = 6;
	defparam lut_4159.mask = 64'h77ff77ff05370f3f;

	lut_sub lut_4163 ({sk[920], i_9_, i_7_, i_8_, i_6_, n_n509, n_n260}, x11772x);
	defparam lut_4163.LUT_SIZE = 7;
	defparam lut_4163.mask = 128'h777f777f777f777f0001010001000100;

	lut_sub lut_4168 ({sk[921], x25x, x17x, x552x, x549x}, x185x);
	defparam lut_4168.LUT_SIZE = 5;
	defparam lut_4168.mask = 32'h0fff0537;

	lut_sub lut_4171 ({sk[922], i_9_, i_7_, i_8_, i_6_, n_n518, n_n260}, x372x);
	defparam lut_4171.LUT_SIZE = 7;
	defparam lut_4171.mask = 128'h777f777f777f777f0000000100000100;

	lut_sub lut_4174 ({sk[923], i_9_, i_7_, i_8_, i_6_, n_n518, n_n260}, x11778x);
	defparam lut_4174.LUT_SIZE = 7;
	defparam lut_4174.mask = 128'h777f777f777f777f0001101001100000;

	lut_sub lut_4180 ({sk[924], i_9_, x25x, n_n518, n_n532, n_n260, x552x}, x11777x);
	defparam lut_4180.LUT_SIZE = 7;
	defparam lut_4180.mask = 128'h777f777f777f777f0507053700030033;

	lut_sub lut_4185 ({sk[925], x17x, x20x, x482x, x102x, x596x, x480x}, x22246x);
	defparam lut_4185.LUT_SIZE = 7;
	defparam lut_4185.mask = 128'h777f777f777f777ff0f0c0c0a0008000;

	lut_sub lut_4190 ({sk[926], i_9_, i_1_, i_2_, i_0_, x537x}, n_n4384);
	defparam lut_4190.LUT_SIZE = 6;
	defparam lut_4190.mask = 64'h77ff77ff00000001;

	lut_sub lut_4192 ({sk[927], i_9_, i_7_, i_8_, i_6_, x571x}, n_n4633);
	defparam lut_4192.LUT_SIZE = 6;
	defparam lut_4192.mask = 64'h77ff77ff00010000;

	lut_sub lut_4194 ({sk[928], i_9_, i_7_, i_8_, i_6_, x541x}, n_n4489);
	defparam lut_4194.LUT_SIZE = 6;
	defparam lut_4194.mask = 64'h77ff77ff00010000;

	lut_sub lut_4196 ({sk[929], i_9_, i_1_, i_2_, i_0_, x574x}, n_n4504);
	defparam lut_4196.LUT_SIZE = 6;
	defparam lut_4196.mask = 64'h77ff77ff00000010;

	lut_sub lut_4198 ({sk[930], i_9_, i_1_, i_2_, i_0_, x550x}, n_n4568);
	defparam lut_4198.LUT_SIZE = 6;
	defparam lut_4198.mask = 64'h77ff77ff00000100;

	lut_sub lut_4200 ({sk[931], i_9_, i_1_, i_2_, i_0_, x537x}, n_n4640);
	defparam lut_4200.LUT_SIZE = 6;
	defparam lut_4200.mask = 64'h77ff77ff00000100;

	lut_sub lut_4202 ({sk[932], i_9_, i_7_, i_8_, i_6_, x486x}, n_n5127);
	defparam lut_4202.LUT_SIZE = 6;
	defparam lut_4202.mask = 64'h77ff77ff40000000;

	lut_sub lut_4204 ({sk[933], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x533x);
	defparam lut_4204.LUT_SIZE = 7;
	defparam lut_4204.mask = 128'h777f777f777f777f2000000000000000;

	lut_sub lut_4206 ({sk[934], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x579x);
	defparam lut_4206.LUT_SIZE = 7;
	defparam lut_4206.mask = 128'h777f777f777f777f0000000000800000;

	lut_sub lut_4208 ({sk[935], x13x, x24x, x586x, x584x, x543x}, n_n4246);
	defparam lut_4208.LUT_SIZE = 6;
	defparam lut_4208.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_4212 ({sk[936], i_9_, i_7_, i_8_, i_6_, x554x}, n_n5087);
	defparam lut_4212.LUT_SIZE = 6;
	defparam lut_4212.mask = 64'h77ff77ff10000000;

	lut_sub lut_4214 ({sk[937], x15x, x10x, x24x, x583x, x559x}, n_n881);
	defparam lut_4214.LUT_SIZE = 6;
	defparam lut_4214.mask = 64'h77ff77ff03573377;

	lut_sub lut_4218 ({sk[938], i_9_, i_1_, i_2_, i_0_, x539x}, n_n4592);
	defparam lut_4218.LUT_SIZE = 6;
	defparam lut_4218.mask = 64'h77ff77ff00000100;

	lut_sub lut_4220 ({sk[939], x539x, x11x, x10x, x583x}, x172x);
	defparam lut_4220.LUT_SIZE = 5;
	defparam lut_4220.mask = 32'h0fff0537;

	lut_sub lut_4223 ({sk[940], i_9_, i_7_, i_8_, i_6_, n_n518, n_n390}, n_n4083);
	defparam lut_4223.LUT_SIZE = 7;
	defparam lut_4223.mask = 128'h777f777f777f777f0101111001101010;

	lut_sub lut_4233 ({sk[941], x21x, x13x, x490x, x20x, x540x}, n_n3520);
	defparam lut_4233.LUT_SIZE = 6;
	defparam lut_4233.mask = 64'h77ff77ff111f555f;

	lut_sub lut_4237 ({sk[942], i_9_, i_1_, i_2_, i_0_, x594x}, n_n4584);
	defparam lut_4237.LUT_SIZE = 6;
	defparam lut_4237.mask = 64'h77ff77ff00000100;

	lut_sub lut_4239 ({sk[943], x17x, x484x, x478x, x23x, x564x}, x461x);
	defparam lut_4239.LUT_SIZE = 6;
	defparam lut_4239.mask = 64'h77ff77ff00335f7f;

	lut_sub lut_4243 ({sk[944], i_9_, i_7_, i_8_, i_6_, n_n260, n_n500}, x13850x);
	defparam lut_4243.LUT_SIZE = 7;
	defparam lut_4243.mask = 128'h777f777f777f777f0001001001000010;

	lut_sub lut_4248 ({sk[945], i_9_, i_1_, i_2_, i_0_, x548x}, n_n4572);
	defparam lut_4248.LUT_SIZE = 6;
	defparam lut_4248.mask = 64'h77ff77ff00000100;

	lut_sub lut_4250 ({sk[946], i_9_, i_7_, i_8_, i_6_, x547x}, n_n4573);
	defparam lut_4250.LUT_SIZE = 6;
	defparam lut_4250.mask = 64'h77ff77ff01000000;

	lut_sub lut_4252 ({sk[947], i_9_, i_7_, i_8_, i_6_, n_n390, n_n535}, x14101x);
	defparam lut_4252.LUT_SIZE = 7;
	defparam lut_4252.mask = 128'h777f777f777f777f0111101101010010;

	lut_sub lut_4262 ({sk[948], x22x, x10x, x583x, x481x}, x14085x);
	defparam lut_4262.LUT_SIZE = 5;
	defparam lut_4262.mask = 32'h0fff0537;

	lut_sub lut_4265 ({sk[949], x25x, x15x, x10x, x479x, x480x}, x14086x);
	defparam lut_4265.LUT_SIZE = 6;
	defparam lut_4265.mask = 64'h77ff77ff05373737;

	lut_sub lut_4269 ({sk[950], i_9_, i_7_, i_8_, n_n518, n_n390}, x22168x);
	defparam lut_4269.LUT_SIZE = 6;
	defparam lut_4269.mask = 64'h77ff77fffeefeeff;

	lut_sub lut_4275 ({sk[951], x10x, x594x, x546x, x593x, x172x}, x22169x);
	defparam lut_4275.LUT_SIZE = 6;
	defparam lut_4275.mask = 64'h77ff77ffaaaa8000;

	lut_sub lut_4278 ({sk[952], x14085x, x14086x, x22168x, x22169x}, x14102x);
	defparam lut_4278.LUT_SIZE = 5;
	defparam lut_4278.mask = 32'h0fffefff;

	lut_sub lut_4283 ({sk[953], x15x, x13x, x508x, x505x, x504x}, n_n3504);
	defparam lut_4283.LUT_SIZE = 6;
	defparam lut_4283.mask = 64'h77ff77ff003f557f;

	lut_sub lut_4287 ({sk[954], i_9_, i_7_, i_8_, i_6_, x543x}, n_n4531);
	defparam lut_4287.LUT_SIZE = 6;
	defparam lut_4287.mask = 64'h77ff77ff00400000;

	lut_sub lut_4289 ({sk[955], x13x, x23x, x529x, x504x}, x429x);
	defparam lut_4289.LUT_SIZE = 5;
	defparam lut_4289.mask = 32'h0fff0537;

	lut_sub lut_4292 ({sk[956], i_9_, n_n455, n_n534, n_n464, x429x}, n_n3871);
	defparam lut_4292.LUT_SIZE = 6;
	defparam lut_4292.mask = 64'h77ff77ff55575555;

	lut_sub lut_4295 ({sk[957], i_9_, i_7_, i_8_, i_6_, n_n455, n_n464}, x14106x);
	defparam lut_4295.LUT_SIZE = 7;
	defparam lut_4295.mask = 128'h777f777f777f777f0100001001010010;

	lut_sub lut_4301 ({sk[958], i_9_, i_7_, i_8_, i_6_, n_n455, n_n473}, x202x);
	defparam lut_4301.LUT_SIZE = 7;
	defparam lut_4301.mask = 128'h777f777f777f777f0110100010101000;

	lut_sub lut_4308 ({sk[959], x13x, x510x, x23x, x543x}, x415x);
	defparam lut_4308.LUT_SIZE = 5;
	defparam lut_4308.mask = 32'h0fff111f;

	lut_sub lut_4311 ({sk[960], x13x, x24x, x523x, x528x}, x430x);
	defparam lut_4311.LUT_SIZE = 5;
	defparam lut_4311.mask = 32'h0fff0357;

	lut_sub lut_4314 ({sk[961], x10x, x550x, x23x, x523x}, x222x);
	defparam lut_4314.LUT_SIZE = 5;
	defparam lut_4314.mask = 32'h0fff111f;

	lut_sub lut_4317 ({sk[962], x13x, x509x, x510x, x558x, x23x, x543x}, x14112x);
	defparam lut_4317.LUT_SIZE = 7;
	defparam lut_4317.mask = 128'h777f777f777f777f111111111fffffff;

	lut_sub lut_4322 ({sk[963], x15x, x21x, x543x, n_n3504, x202x}, x14115x);
	defparam lut_4322.LUT_SIZE = 6;
	defparam lut_4322.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_4327 ({sk[964], n_n3871, x14106x, x430x, x222x, x14112x, x14115x}, x14117x);
	defparam lut_4327.LUT_SIZE = 7;
	defparam lut_4327.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_4334 ({sk[965], n_n1649, x348x, x349x, x14076x, x14077x, x14079x}, x22167x);
	defparam lut_4334.LUT_SIZE = 7;
	defparam lut_4334.mask = 128'h777f777f777f777f8000000000000000;

	lut_sub lut_4336 ({sk[966], n_n3346, x14101x, x14102x, x22167x}, x14118x);
	defparam lut_4336.LUT_SIZE = 5;
	defparam lut_4336.mask = 32'h0fffbfff;

	lut_sub lut_4341 ({sk[967], i_9_, i_7_, i_8_, i_6_, x561x}, n_n4629);
	defparam lut_4341.LUT_SIZE = 6;
	defparam lut_4341.mask = 64'h77ff77ff04000000;

	lut_sub lut_4343 ({sk[968], i_9_, i_7_, i_8_, i_6_, x552x}, n_n4839);
	defparam lut_4343.LUT_SIZE = 6;
	defparam lut_4343.mask = 64'h77ff77ff40000000;

	lut_sub lut_4345 ({sk[969], i_9_, i_7_, i_8_, i_6_, x592x}, n_n5303);
	defparam lut_4345.LUT_SIZE = 6;
	defparam lut_4345.mask = 64'h77ff77ff40000000;

	lut_sub lut_4347 ({sk[970], i_9_, i_7_, i_8_, i_6_, x591x}, n_n5173);
	defparam lut_4347.LUT_SIZE = 6;
	defparam lut_4347.mask = 64'h77ff77ff04000000;

	lut_sub lut_4349 ({sk[971], x19x, x478x, x23x, x573x, x493x, x579x}, x13710x);
	defparam lut_4349.LUT_SIZE = 7;
	defparam lut_4349.mask = 128'h777f777f777f777f005500553f7fffff;

	lut_sub lut_4354 ({sk[972], x15x, x592x, x19x, x482x, x569x}, x13709x);
	defparam lut_4354.LUT_SIZE = 6;
	defparam lut_4354.mask = 64'h77ff77ff030357ff;

	lut_sub lut_4358 ({sk[973], x15x, x19x, x591x, x559x}, x13700x);
	defparam lut_4358.LUT_SIZE = 5;
	defparam lut_4358.mask = 32'h0fff0537;

	lut_sub lut_4361 ({sk[974], x19x, x545x, x23x, x581x, x599x}, x13702x);
	defparam lut_4361.LUT_SIZE = 6;
	defparam lut_4361.mask = 64'h77ff77ff050537ff;

	lut_sub lut_4365 ({sk[975], i_9_, x25x, x515x, n_n482, n_n520, n_n65}, x13713x);
	defparam lut_4365.LUT_SIZE = 7;
	defparam lut_4365.mask = 128'h777f777f777f777f010101ff010101ff;

	lut_sub lut_4369 ({sk[976], x24x, x558x, x12x, x20x, x591x, x505x}, x22181x);
	defparam lut_4369.LUT_SIZE = 7;
	defparam lut_4369.mask = 128'h777f777f777f777ffca8fc00cc88cc00;

	lut_sub lut_4374 ({sk[977], i_9_, n_n518, x24x, n_n534, n_n130, x532x}, x13718x);
	defparam lut_4374.LUT_SIZE = 7;
	defparam lut_4374.mask = 128'h777f777f777f777f0505053700000333;

	lut_sub lut_4378 ({sk[978], x21x, x18x, x522x, n_n5085, x532x, n_n5082}, x22180x);
	defparam lut_4378.LUT_SIZE = 7;
	defparam lut_4378.mask = 128'h777f777f777f777fa0a0a00080808000;

	lut_sub lut_4383 ({sk[979], i_9_, i_7_, i_8_, i_6_, x542x}, n_n4517);
	defparam lut_4383.LUT_SIZE = 6;
	defparam lut_4383.mask = 64'h77ff77ff04000000;

	lut_sub lut_4385 ({sk[980], x13x, x570x, x20x, x23x, x542x}, n_n3152);
	defparam lut_4385.LUT_SIZE = 6;
	defparam lut_4385.mask = 64'h77ff77ff151515ff;

	lut_sub lut_4389 ({sk[981], i_9_, i_1_, i_2_, i_0_, x539x}, n_n5104);
	defparam lut_4389.LUT_SIZE = 6;
	defparam lut_4389.mask = 64'h77ff77ff00000400;

	lut_sub lut_4391 ({sk[982], x25x, x16x, x499x, x574x}, x423x);
	defparam lut_4391.LUT_SIZE = 5;
	defparam lut_4391.mask = 32'h0fff0537;

	lut_sub lut_4394 ({sk[983], x16x, x24x, x499x, x572x, x536x, n_n4367}, x22142x);
	defparam lut_4394.LUT_SIZE = 7;
	defparam lut_4394.mask = 128'h777f777f777f777faaaaaa0080808000;

	lut_sub lut_4399 ({sk[984], x16x, x21x, x472x, x478x, x473x}, x15032x);
	defparam lut_4399.LUT_SIZE = 6;
	defparam lut_4399.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_4403 ({sk[985], x16x, x20x, x562x, x556x, x473x}, x22281x);
	defparam lut_4403.LUT_SIZE = 6;
	defparam lut_4403.mask = 64'h77ff77ffffaac080;

	lut_sub lut_4408 ({sk[986], i_9_, i_7_, i_8_, i_6_, n_n536, n_n473}, n_n2634);
	defparam lut_4408.LUT_SIZE = 7;
	defparam lut_4408.mask = 128'h777f777f777f777f1010111011010100;

	lut_sub lut_4418 ({sk[987], i_9_, i_7_, i_8_, i_6_, n_n536, n_n482}, x15049x);
	defparam lut_4418.LUT_SIZE = 7;
	defparam lut_4418.mask = 128'h777f777f777f777f0001001001000010;

	lut_sub lut_4423 ({sk[988], i_9_, i_7_, i_8_, i_6_, n_n536, n_n464}, x15055x);
	defparam lut_4423.LUT_SIZE = 7;
	defparam lut_4423.mask = 128'h777f777f777f777f0101010101010111;

	lut_sub lut_4433 ({sk[989], x25x, x16x, x493x, x495x}, x15047x);
	defparam lut_4433.LUT_SIZE = 5;
	defparam lut_4433.mask = 32'h0fff0357;

	lut_sub lut_4436 ({sk[990], x16x, x500x, x510x, x20x, x580x}, x15048x);
	defparam lut_4436.LUT_SIZE = 6;
	defparam lut_4436.mask = 64'h77ff77ff00335f7f;

	lut_sub lut_4440 ({sk[991], i_9_, i_7_, i_8_, i_6_, x552x}, n_n4837);
	defparam lut_4440.LUT_SIZE = 6;
	defparam lut_4440.mask = 64'h77ff77ff04000000;

	lut_sub lut_4442 ({sk[992], i_9_, i_7_, i_8_, i_6_, x511x}, n_n4797);
	defparam lut_4442.LUT_SIZE = 6;
	defparam lut_4442.mask = 64'h77ff77ff01000000;

	lut_sub lut_4444 ({sk[993], x15x, x17x, x512x, x505x}, x132x);
	defparam lut_4444.LUT_SIZE = 5;
	defparam lut_4444.mask = 32'h0fff0537;

	lut_sub lut_4447 ({sk[994], x21x, x12x, x20x, x598x, x494x}, n_n4144);
	defparam lut_4447.LUT_SIZE = 6;
	defparam lut_4447.mask = 64'h77ff77ff03573377;

	lut_sub lut_4451 ({sk[995], x12x, x554x, x23x, x593x}, x34x);
	defparam lut_4451.LUT_SIZE = 5;
	defparam lut_4451.mask = 32'h0fff0357;

	lut_sub lut_4454 ({sk[996], i_9_, i_7_, i_8_, i_6_, x598x}, x289x);
	defparam lut_4454.LUT_SIZE = 6;
	defparam lut_4454.mask = 64'h77ff77ff01040000;

	lut_sub lut_4457 ({sk[997], i_9_, i_7_, i_8_, i_6_, n_n518, n_n130}, x16719x);
	defparam lut_4457.LUT_SIZE = 7;
	defparam lut_4457.mask = 128'h777f777f777f777f0010100000110001;

	lut_sub lut_4463 ({sk[998], x21x, x13x, x518x, x541x}, x65x);
	defparam lut_4463.LUT_SIZE = 5;
	defparam lut_4463.mask = 32'h0fff0357;

	lut_sub lut_4466 ({sk[999], x15x, x13x, x24x, x480x, x476x}, n_n4254);
	defparam lut_4466.LUT_SIZE = 6;
	defparam lut_4466.mask = 64'h77ff77ff05375577;

	lut_sub lut_4470 ({sk[1000], i_9_, i_1_, i_2_, i_0_, x474x, x475x}, x184x);
	defparam lut_4470.LUT_SIZE = 7;
	defparam lut_4470.mask = 128'h777f777f777f777f0000000000000700;

	lut_sub lut_4473 ({sk[1001], x15x, x17x, x545x, x552x}, x38x);
	defparam lut_4473.LUT_SIZE = 5;
	defparam lut_4473.mask = 32'h0fff0357;

	lut_sub lut_4476 ({sk[1002], i_9_, n_n528, n_n260, n_n535, x548x, x38x}, x388x);
	defparam lut_4476.LUT_SIZE = 7;
	defparam lut_4476.mask = 128'h777f777f777f777f5555555f55775577;

	lut_sub lut_4480 ({sk[1003], i_9_, i_1_, i_2_, i_0_, x489x}, n_n4820);
	defparam lut_4480.LUT_SIZE = 6;
	defparam lut_4480.mask = 64'h77ff77ff00001000;

	lut_sub lut_4482 ({sk[1004], i_9_, i_7_, i_8_, i_6_, x530x}, x186x);
	defparam lut_4482.LUT_SIZE = 6;
	defparam lut_4482.mask = 64'h77ff77ff04400000;

	lut_sub lut_4485 ({sk[1005], i_9_, i_7_, i_8_, i_6_, n_n536, n_n473}, n_n2263);
	defparam lut_4485.LUT_SIZE = 7;
	defparam lut_4485.mask = 128'h777f777f777f777f0100111101010101;

	lut_sub lut_4495 ({sk[1006], i_9_, i_7_, i_8_, i_6_, n_n536, n_n464}, x16527x);
	defparam lut_4495.LUT_SIZE = 7;
	defparam lut_4495.mask = 128'h777f777f777f777f1100001001010000;

	lut_sub lut_4501 ({sk[1007], x22x, x16x, x500x, x520x}, x93x);
	defparam lut_4501.LUT_SIZE = 5;
	defparam lut_4501.mask = 32'h0fff0537;

	lut_sub lut_4504 ({sk[1008], i_9_, i_7_, i_8_, i_6_, x500x}, n_n4399);
	defparam lut_4504.LUT_SIZE = 6;
	defparam lut_4504.mask = 64'h77ff77ff10000000;

	lut_sub lut_4506 ({sk[1009], i_9_, i_7_, i_8_, i_6_, n_n536, n_n482}, x16533x);
	defparam lut_4506.LUT_SIZE = 7;
	defparam lut_4506.mask = 128'h777f777f777f777f0100111101011001;

	lut_sub lut_4516 ({sk[1010], x16x, x23x, x506x, x495x}, x215x);
	defparam lut_4516.LUT_SIZE = 5;
	defparam lut_4516.mask = 32'h0fff0537;

	lut_sub lut_4519 ({sk[1011], i_9_, i_1_, i_2_, i_0_, x550x, x516x}, x16523x);
	defparam lut_4519.LUT_SIZE = 7;
	defparam lut_4519.mask = 128'h777f777f777f777f0000000000000305;

	lut_sub lut_4522 ({sk[1012], x16x, x490x, x23x, x497x, x546x}, n_n2446);
	defparam lut_4522.LUT_SIZE = 6;
	defparam lut_4522.mask = 64'h77ff77ff030357ff;

	lut_sub lut_4526 ({sk[1013], i_9_, i_7_, i_8_, i_6_, n_n536, n_n509}, x16537x);
	defparam lut_4526.LUT_SIZE = 7;
	defparam lut_4526.mask = 128'h777f777f777f777f0100001001001000;

	lut_sub lut_4531 ({sk[1014], x15x, x16x, x501x, x585x}, x198x);
	defparam lut_4531.LUT_SIZE = 5;
	defparam lut_4531.mask = 32'h0fff0537;

	lut_sub lut_4534 ({sk[1015], x16x, x24x, x497x, x549x}, x283x);
	defparam lut_4534.LUT_SIZE = 5;
	defparam lut_4534.mask = 32'h0fff0357;

	lut_sub lut_4537 ({sk[1016], x16x, x501x, x475x, x23x}, x16535x);
	defparam lut_4537.LUT_SIZE = 5;
	defparam lut_4537.mask = 32'h0fff0537;

	lut_sub lut_4540 ({sk[1017], x15x, x16x, x24x, x481x, x473x}, x16536x);
	defparam lut_4540.LUT_SIZE = 6;
	defparam lut_4540.mask = 64'h77ff77ff05375577;

	lut_sub lut_4544 ({sk[1018], x22x, x16x, x539x, x11x, x497x}, x16540x);
	defparam lut_4544.LUT_SIZE = 6;
	defparam lut_4544.mask = 64'h77ff77ff111f555f;

	lut_sub lut_4548 ({sk[1019], i_9_, n_n536, n_n518, n_n530, x283x}, x16541x);
	defparam lut_4548.LUT_SIZE = 6;
	defparam lut_4548.mask = 64'h77ff77ff55575557;

	lut_sub lut_4552 ({sk[1020], x16x, x21x, x472x, x564x, x563x, x473x}, x16548x);
	defparam lut_4552.LUT_SIZE = 7;
	defparam lut_4552.mask = 128'h777f777f777f777f000055553fff7fff;

	lut_sub lut_4557 ({sk[1021], x492x, x16x, x570x, x23x, x499x}, n_n2435);
	defparam lut_4557.LUT_SIZE = 6;
	defparam lut_4557.mask = 64'h77ff77ff111f11ff;

	lut_sub lut_4561 ({sk[1022], i_9_, i_7_, i_8_, i_6_, n_n536, n_n491}, x54x);
	defparam lut_4561.LUT_SIZE = 7;
	defparam lut_4561.mask = 128'h777f777f777f777f0101001000001010;

	lut_sub lut_4567 ({sk[1023], x22x, x16x, x518x, x498x, x536x}, x282x);
	defparam lut_4567.LUT_SIZE = 6;
	defparam lut_4567.mask = 64'h77ff77ff005f337f;

	lut_sub lut_4571 ({sk[1024], x16x, x21x, x491x, x498x}, x300x);
	defparam lut_4571.LUT_SIZE = 5;
	defparam lut_4571.mask = 32'h0fff0537;

	lut_sub lut_4574 ({sk[1025], i_9_, i_7_, i_8_, i_6_, x541x}, n_n4503);
	defparam lut_4574.LUT_SIZE = 6;
	defparam lut_4574.mask = 64'h77ff77ff40000000;

	lut_sub lut_4576 ({sk[1026], i_9_, i_1_, i_2_, i_0_, x586x, x537x}, x16582x);
	defparam lut_4576.LUT_SIZE = 7;
	defparam lut_4576.mask = 128'h777f777f777f777f0000000000000700;

	lut_sub lut_4579 ({sk[1027], x538x, x13x, x11x, x557x, x542x}, x16584x);
	defparam lut_4579.LUT_SIZE = 6;
	defparam lut_4579.mask = 64'h77ff77ff053705ff;

	lut_sub lut_4583 ({sk[1028], x21x, x13x, x516x, x523x}, x455x);
	defparam lut_4583.LUT_SIZE = 5;
	defparam lut_4583.mask = 32'h0fff0357;

	lut_sub lut_4586 ({sk[1029], x25x, x10x, x547x, x549x}, x121x);
	defparam lut_4586.LUT_SIZE = 5;
	defparam lut_4586.mask = 32'h0fff0537;

	lut_sub lut_4589 ({sk[1030], x13x, x20x, x525x, x489x, x523x}, n_n4239);
	defparam lut_4589.LUT_SIZE = 6;
	defparam lut_4589.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_4593 ({sk[1031], i_9_, i_7_, i_8_, i_6_, n_n390, n_n535}, x16605x);
	defparam lut_4593.LUT_SIZE = 7;
	defparam lut_4593.mask = 128'h777f777f777f777f0101100000001000;

	lut_sub lut_4598 ({sk[1032], x10x, x490x, x23x, x547x, x594x}, x16604x);
	defparam lut_4598.LUT_SIZE = 6;
	defparam lut_4598.mask = 64'h77ff77ff030357ff;

	lut_sub lut_4602 ({sk[1033], i_9_, i_7_, i_8_, i_6_, n_n518, n_n390}, x16622x);
	defparam lut_4602.LUT_SIZE = 7;
	defparam lut_4602.mask = 128'h777f777f777f777f0101011101010110;

	lut_sub lut_4612 ({sk[1034], x21x, x11x, x10x, x479x, x564x, x563x}, x16611x);
	defparam lut_4612.LUT_SIZE = 7;
	defparam lut_4612.mask = 128'h777f777f777f777f00770f7f0f7f0f7f;

	lut_sub lut_4617 ({sk[1035], i_9_, i_7_, i_8_, i_6_, n_n390, n_n509}, x16612x);
	defparam lut_4617.LUT_SIZE = 7;
	defparam lut_4617.mask = 128'h777f777f777f777f0010001010001010;

	lut_sub lut_4623 ({sk[1036], x25x, x521x, x10x, x477x, x479x, x581x}, x16617x);
	defparam lut_4623.LUT_SIZE = 7;
	defparam lut_4623.mask = 128'h777f777f777f777f005f00ff337f33ff;

	lut_sub lut_4628 ({sk[1037], x15x, x10x, x24x, x482x, x479x, x255x}, x22080x);
	defparam lut_4628.LUT_SIZE = 7;
	defparam lut_4628.mask = 128'h777f777f777f777faa88a08088888080;

	lut_sub lut_4633 ({sk[1038], x15x, x10x, x571x, x557x}, x271x);
	defparam lut_4633.LUT_SIZE = 5;
	defparam lut_4633.mask = 32'h0fff0537;

	lut_sub lut_4636 ({sk[1039], i_9_, i_7_, i_8_, i_6_, n_n390, n_n491}, x16636x);
	defparam lut_4636.LUT_SIZE = 7;
	defparam lut_4636.mask = 128'h777f777f777f777f0100011100001000;

	lut_sub lut_4642 ({sk[1040], i_9_, i_7_, i_8_, i_6_, n_n390, n_n500}, n_n2246);
	defparam lut_4642.LUT_SIZE = 7;
	defparam lut_4642.mask = 128'h777f777f777f777f0011111010111000;

	lut_sub lut_4652 ({sk[1041], x492x, x10x, x24x, x582x}, x16625x);
	defparam lut_4652.LUT_SIZE = 5;
	defparam lut_4652.mask = 32'h0fff111f;

	lut_sub lut_4655 ({sk[1042], x13x, x20x, x488x, x504x}, x212x);
	defparam lut_4655.LUT_SIZE = 5;
	defparam lut_4655.mask = 32'h0fff0537;

	lut_sub lut_4658 ({sk[1043], x13x, x11x, x524x, x523x}, x213x);
	defparam lut_4658.LUT_SIZE = 5;
	defparam lut_4658.mask = 32'h0fff0537;

	lut_sub lut_4661 ({sk[1044], i_9_, i_7_, i_8_, i_6_, x501x}, n_n4341);
	defparam lut_4661.LUT_SIZE = 6;
	defparam lut_4661.mask = 64'h77ff77ff04000000;

	lut_sub lut_4663 ({sk[1045], x25x, x24x, x18x, x586x, x598x, x577x}, x16790x);
	defparam lut_4663.LUT_SIZE = 7;
	defparam lut_4663.mask = 128'h777f777f777f777f000f777f333f777f;

	lut_sub lut_4668 ({sk[1046], x15x, x22x, x474x, x12x, x486x}, x16789x);
	defparam lut_4668.LUT_SIZE = 6;
	defparam lut_4668.mask = 64'h77ff77ff03575757;

	lut_sub lut_4672 ({sk[1047], x521x, x539x, x12x, x16790x, x16789x}, n_n2092);
	defparam lut_4672.LUT_SIZE = 6;
	defparam lut_4672.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_4677 ({sk[1048], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x555x);
	defparam lut_4677.LUT_SIZE = 7;
	defparam lut_4677.mask = 128'h777f777f777f777f0000000000000080;

	lut_sub lut_4679 ({sk[1049], i_9_, i_7_, i_8_, i_6_, x555x}, n_n5223);
	defparam lut_4679.LUT_SIZE = 6;
	defparam lut_4679.mask = 64'h77ff77ff40000000;

	lut_sub lut_4681 ({sk[1050], i_9_, i_7_, i_8_, i_6_, x487x}, n_n5249);
	defparam lut_4681.LUT_SIZE = 6;
	defparam lut_4681.mask = 64'h77ff77ff00040000;

	lut_sub lut_4683 ({sk[1051], i_9_, i_1_, i_2_, i_0_, x557x}, n_n5278);
	defparam lut_4683.LUT_SIZE = 6;
	defparam lut_4683.mask = 64'h77ff77ff00004000;

	lut_sub lut_4685 ({sk[1052], i_9_, i_7_, i_8_, i_6_, x555x}, n_n5217);
	defparam lut_4685.LUT_SIZE = 6;
	defparam lut_4685.mask = 64'h77ff77ff00040000;

	lut_sub lut_4687 ({sk[1053], x19x, x22x, x522x, x478x, x599x, x487x}, x16777x);
	defparam lut_4687.LUT_SIZE = 7;
	defparam lut_4687.mask = 128'h777f777f777f777f000077770fff7fff;

	lut_sub lut_4692 ({sk[1054], x22x, x12x, x23x, x525x, n_n5216, x555x}, x22063x);
	defparam lut_4692.LUT_SIZE = 7;
	defparam lut_4692.mask = 128'h777f777f777f777fcc88c08088888080;

	lut_sub lut_4697 ({sk[1055], x25x, x592x, x19x, x586x, x557x, x494x}, x22299x);
	defparam lut_4697.LUT_SIZE = 7;
	defparam lut_4697.mask = 128'h777f777f777f777fff80ff80ff800000;

	lut_sub lut_4702 ({sk[1056], i_9_, x11x, n_n509, n_n325, n_n522, x564x}, x16119x);
	defparam lut_4702.LUT_SIZE = 7;
	defparam lut_4702.mask = 128'h777f777f777f777f0003000f0507050f;

	lut_sub lut_4707 ({sk[1057], i_9_, i_7_, i_8_, i_6_, n_n509, n_n325}, x16120x);
	defparam lut_4707.LUT_SIZE = 7;
	defparam lut_4707.mask = 128'h777f777f777f777f1000000111000001;

	lut_sub lut_4713 ({sk[1058], i_9_, i_1_, i_2_, i_0_, x574x}, n_n5016);
	defparam lut_4713.LUT_SIZE = 6;
	defparam lut_4713.mask = 64'h77ff77ff00000040;

	lut_sub lut_4715 ({sk[1059], i_9_, i_7_, i_8_, i_6_, n_n491, n_n195}, x12252x);
	defparam lut_4715.LUT_SIZE = 7;
	defparam lut_4715.mask = 128'h777f777f777f777f0101010000010000;

	lut_sub lut_4720 ({sk[1060], i_9_, i_1_, i_2_, i_0_, x509x}, n_n5306);
	defparam lut_4720.LUT_SIZE = 6;
	defparam lut_4720.mask = 64'h77ff77ff00004000;

	lut_sub lut_4722 ({sk[1061], x515x, x19x, x509x, x24x, x508x}, n_n3019);
	defparam lut_4722.LUT_SIZE = 6;
	defparam lut_4722.mask = 64'h77ff77ff005f337f;

	lut_sub lut_4726 ({sk[1062], i_9_, i_7_, i_8_, i_6_, x534x}, n_n5335);
	defparam lut_4726.LUT_SIZE = 6;
	defparam lut_4726.mask = 64'h77ff77ff40000000;

	lut_sub lut_4728 ({sk[1063], x25x, x10x, x561x, x563x, x547x, x535x}, x12048x);
	defparam lut_4728.LUT_SIZE = 7;
	defparam lut_4728.mask = 128'h777f777f777f777f00005f5f33ff7fff;

	lut_sub lut_4733 ({sk[1064], x10x, x24x, x490x, x571x}, x12046x);
	defparam lut_4733.LUT_SIZE = 5;
	defparam lut_4733.mask = 32'h0fff0537;

	lut_sub lut_4736 ({sk[1065], i_9_, i_1_, i_2_, i_0_, x593x}, n_n4458);
	defparam lut_4736.LUT_SIZE = 6;
	defparam lut_4736.mask = 64'h77ff77ff00000010;

	lut_sub lut_4738 ({sk[1066], x16x, x24x, x541x, x525x}, x12050x);
	defparam lut_4738.LUT_SIZE = 5;
	defparam lut_4738.mask = 32'h0fff0357;

	lut_sub lut_4741 ({sk[1067], x21x, x13x, x20x, x481x, x476x}, x12052x);
	defparam lut_4741.LUT_SIZE = 6;
	defparam lut_4741.mask = 64'h77ff77ff05375577;

	lut_sub lut_4745 ({sk[1068], x13x, x24x, x516x, x502x, x573x, x523x}, x12060x);
	defparam lut_4745.LUT_SIZE = 7;
	defparam lut_4745.mask = 128'h777f777f777f777f000055553fff7fff;

	lut_sub lut_4750 ({sk[1069], x13x, x558x, x23x, x537x, x536x, x543x}, x22270x);
	defparam lut_4750.LUT_SIZE = 7;
	defparam lut_4750.mask = 128'h777f777f777f777fffaaffaac0800000;

	lut_sub lut_4755 ({sk[1070], x24x, x14x, x572x, x575x}, x350x);
	defparam lut_4755.LUT_SIZE = 5;
	defparam lut_4755.mask = 32'h0fff0357;

	lut_sub lut_4758 ({sk[1071], x483x, x14x, x23x, x480x}, x12066x);
	defparam lut_4758.LUT_SIZE = 5;
	defparam lut_4758.mask = 32'h0fff0537;

	lut_sub lut_4761 ({sk[1072], x22x, x483x, x14x, x491x, x494x, n_n4759}, x22225x);
	defparam lut_4761.LUT_SIZE = 7;
	defparam lut_4761.mask = 128'h777f777f777f777faa80aa80aa800000;

	lut_sub lut_4766 ({sk[1073], x25x, x11x, x10x, x509x, x557x, x582x}, x12074x);
	defparam lut_4766.LUT_SIZE = 7;
	defparam lut_4766.mask = 128'h777f777f777f777f003f557f557f557f;

	lut_sub lut_4771 ({sk[1074], x10x, x14x, x490x, x520x, x593x}, x22255x);
	defparam lut_4771.LUT_SIZE = 6;
	defparam lut_4771.mask = 64'h77ff77ffffa0cc80;

	lut_sub lut_4776 ({sk[1075], x15x, x14x, x570x, x508x, x596x, x525x}, x12081x);
	defparam lut_4776.LUT_SIZE = 7;
	defparam lut_4776.mask = 128'h777f777f777f777f00005fff33337fff;

	lut_sub lut_4781 ({sk[1076], x21x, x14x, x552x, x580x, x506x, x493x}, x22289x);
	defparam lut_4781.LUT_SIZE = 7;
	defparam lut_4781.mask = 128'h777f777f777f777fffff8080ff008000;

	lut_sub lut_4786 ({sk[1077], i_9_, i_1_, i_2_, i_0_, x517x}, n_n4962);
	defparam lut_4786.LUT_SIZE = 6;
	defparam lut_4786.mask = 64'h77ff77ff00000040;

	lut_sub lut_4788 ({sk[1078], i_9_, i_7_, i_8_, i_6_, x514x}, n_n5189);
	defparam lut_4788.LUT_SIZE = 6;
	defparam lut_4788.mask = 64'h77ff77ff04000000;

	lut_sub lut_4790 ({sk[1079], i_9_, i_1_, i_2_, i_0_, x488x}, n_n5188);
	defparam lut_4790.LUT_SIZE = 6;
	defparam lut_4790.mask = 64'h77ff77ff00000400;

	lut_sub lut_4792 ({sk[1080], i_9_, i_7_, i_8_, i_6_, n_n536, n_n509}, n_n1120);
	defparam lut_4792.LUT_SIZE = 7;
	defparam lut_4792.mask = 128'h777f777f777f777f0110011010101110;

	lut_sub lut_4802 ({sk[1081], i_9_, i_7_, i_8_, i_6_, x542x}, n_n4507);
	defparam lut_4802.LUT_SIZE = 6;
	defparam lut_4802.mask = 64'h77ff77ff00100000;

	lut_sub lut_4804 ({sk[1082], x13x, x11x, x557x, x542x}, x308x);
	defparam lut_4804.LUT_SIZE = 5;
	defparam lut_4804.mask = 32'h0fff0537;

	lut_sub lut_4807 ({sk[1083], i_9_, i_7_, i_8_, i_6_, n_n455, n_n491}, n_n1107);
	defparam lut_4807.LUT_SIZE = 7;
	defparam lut_4807.mask = 128'h777f777f777f777f0101011001011110;

	lut_sub lut_4817 ({sk[1084], x15x, x10x, x561x, x556x, x536x}, n_n3861);
	defparam lut_4817.LUT_SIZE = 6;
	defparam lut_4817.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_4821 ({sk[1085], i_9_, i_1_, i_2_, i_0_, x516x}, n_n5074);
	defparam lut_4821.LUT_SIZE = 6;
	defparam lut_4821.mask = 64'h77ff77ff00000040;

	lut_sub lut_4823 ({sk[1086], x22x, x18x, x516x, x522x, x532x}, n_n4152);
	defparam lut_4823.LUT_SIZE = 6;
	defparam lut_4823.mask = 64'h77ff77ff003f557f;

	lut_sub lut_4827 ({sk[1087], i_9_, i_7_, i_8_, i_6_, n_n473, n_n260}, x11790x);
	defparam lut_4827.LUT_SIZE = 7;
	defparam lut_4827.mask = 128'h777f777f777f777f0001000101010000;

	lut_sub lut_4832 ({sk[1088], x17x, x23x, x512x, x506x}, x180x);
	defparam lut_4832.LUT_SIZE = 5;
	defparam lut_4832.mask = 32'h0fff0357;

	lut_sub lut_4835 ({sk[1089], x17x, x20x, x512x, x488x}, x382x);
	defparam lut_4835.LUT_SIZE = 5;
	defparam lut_4835.mask = 32'h0fff0357;

	lut_sub lut_4838 ({sk[1090], x24x, x17x, x531x, x527x}, x411x);
	defparam lut_4838.LUT_SIZE = 5;
	defparam lut_4838.mask = 32'h0fff0537;

	lut_sub lut_4841 ({sk[1091], x25x, x17x, x531x, x528x}, x11792x);
	defparam lut_4841.LUT_SIZE = 5;
	defparam lut_4841.mask = 32'h0fff0537;

	lut_sub lut_4844 ({sk[1092], x21x, x512x, x180x, x382x, x411x, x11792x}, x11796x);
	defparam lut_4844.LUT_SIZE = 7;
	defparam lut_4844.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_4850 ({sk[1093], x510x, x17x, x23x, x589x}, x105x);
	defparam lut_4850.LUT_SIZE = 5;
	defparam lut_4850.mask = 32'h0fff111f;

	lut_sub lut_4853 ({sk[1094], i_9_, i_1_, i_2_, i_0_, x509x, x502x}, x11788x);
	defparam lut_4853.LUT_SIZE = 7;
	defparam lut_4853.mask = 128'h777f777f777f777f0000000000000070;

	lut_sub lut_4856 ({sk[1095], x17x, x580x, n_n1075, x11790x, x105x, x11788x}, x11797x);
	defparam lut_4856.LUT_SIZE = 7;
	defparam lut_4856.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_4862 ({sk[1096], x25x, x18x, x597x, x593x}, x68x);
	defparam lut_4862.LUT_SIZE = 5;
	defparam lut_4862.mask = 32'h0fff0537;

	lut_sub lut_4865 ({sk[1097], x21x, x18x, x553x, x546x}, x11798x);
	defparam lut_4865.LUT_SIZE = 5;
	defparam lut_4865.mask = 32'h0fff0537;

	lut_sub lut_4868 ({sk[1098], x24x, x545x, x18x, x597x, x548x}, x11800x);
	defparam lut_4868.LUT_SIZE = 6;
	defparam lut_4868.mask = 64'h77ff77ff050f373f;

	lut_sub lut_4872 ({sk[1099], x18x, x517x, x594x, x68x, x11798x, x11800x}, n_n1071);
	defparam lut_4872.LUT_SIZE = 7;
	defparam lut_4872.mask = 128'h777f777f777f777f7f7f7f7f7fffffff;

	lut_sub lut_4878 ({sk[1100], i_9_, i_7_, i_8_, i_6_, n_n260, n_n464}, x11807x);
	defparam lut_4878.LUT_SIZE = 7;
	defparam lut_4878.mask = 128'h777f777f777f777f0100001011000000;

	lut_sub lut_4883 ({sk[1101], x24x, x18x, x550x, x549x, x553x}, x11806x);
	defparam lut_4883.LUT_SIZE = 6;
	defparam lut_4883.mask = 64'h77ff77ff003f557f;

	lut_sub lut_4887 ({sk[1102], x17x, x516x, x489x, x11807x, x11806x}, n_n1072);
	defparam lut_4887.LUT_SIZE = 6;
	defparam lut_4887.mask = 64'h77ff77ff77777fff;

	lut_sub lut_4892 ({sk[1103], x15x, x18x, x597x, x585x, x559x}, x29x);
	defparam lut_4892.LUT_SIZE = 6;
	defparam lut_4892.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_4896 ({sk[1104], i_9_, i_7_, i_8_, i_6_, n_n518, n_n195}, x11815x);
	defparam lut_4896.LUT_SIZE = 7;
	defparam lut_4896.mask = 128'h777f777f777f777f0111101001111000;

	lut_sub lut_4906 ({sk[1105], i_9_, i_7_, i_8_, i_6_, n_n260, n_n500}, n_n1077);
	defparam lut_4906.LUT_SIZE = 7;
	defparam lut_4906.mask = 128'h777f777f777f777f0011110000111110;

	lut_sub lut_4916 ({sk[1106], i_9_, i_7_, i_8_, i_6_, n_n509, n_n260}, x11823x);
	defparam lut_4916.LUT_SIZE = 7;
	defparam lut_4916.mask = 128'h777f777f777f777f0010000010101000;

	lut_sub lut_4921 ({sk[1107], x21x, x17x, x484x, x475x}, x11821x);
	defparam lut_4921.LUT_SIZE = 5;
	defparam lut_4921.mask = 32'h0fff0537;

	lut_sub lut_4924 ({sk[1108], i_9_, i_7_, i_8_, i_6_, x484x, x566x}, x11822x);
	defparam lut_4924.LUT_SIZE = 7;
	defparam lut_4924.mask = 128'h777f777f777f777f0300003500000000;

	lut_sub lut_4928 ({sk[1109], i_9_, i_7_, i_8_, i_6_, n_n260, n_n491}, x11830x);
	defparam lut_4928.LUT_SIZE = 7;
	defparam lut_4928.mask = 128'h777f777f777f777f1010101011111000;

	lut_sub lut_4938 ({sk[1110], n_n1077, x11823x, x11821x, x11822x, x11830x}, x11832x);
	defparam lut_4938.LUT_SIZE = 6;
	defparam lut_4938.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_4944 ({sk[1111], i_9_, i_1_, i_2_, i_0_, x477x}, n_n4350);
	defparam lut_4944.LUT_SIZE = 6;
	defparam lut_4944.mask = 64'h77ff77ff00000001;

	lut_sub lut_4946 ({sk[1112], x15x, x16x, x477x, x480x, x473x}, n_n1002);
	defparam lut_4946.LUT_SIZE = 6;
	defparam lut_4946.mask = 64'h77ff77ff003f557f;

	lut_sub lut_4950 ({sk[1113], i_9_, i_1_, i_2_, i_0_, x493x}, n_n5172);
	defparam lut_4950.LUT_SIZE = 6;
	defparam lut_4950.mask = 64'h77ff77ff00000400;

	lut_sub lut_4952 ({sk[1114], i_9_, i_7_, i_8_, i_6_, x582x}, n_n4661);
	defparam lut_4952.LUT_SIZE = 6;
	defparam lut_4952.mask = 64'h77ff77ff04000000;

	lut_sub lut_4954 ({sk[1115], i_9_, i_7_, i_8_, i_6_, x526x}, n_n4689);
	defparam lut_4954.LUT_SIZE = 6;
	defparam lut_4954.mask = 64'h77ff77ff00040000;

	lut_sub lut_4956 ({sk[1116], i_9_, i_7_, i_8_, i_6_, x551x}, n_n4697);
	defparam lut_4956.LUT_SIZE = 6;
	defparam lut_4956.mask = 64'h77ff77ff00010000;

	lut_sub lut_4958 ({sk[1117], i_9_, i_7_, i_8_, i_6_, x567x}, n_n5011);
	defparam lut_4958.LUT_SIZE = 6;
	defparam lut_4958.mask = 64'h77ff77ff00400000;

	lut_sub lut_4960 ({sk[1118], i_9_, i_7_, i_8_, i_6_, x568x}, n_n5135);
	defparam lut_4960.LUT_SIZE = 6;
	defparam lut_4960.mask = 64'h77ff77ff10000000;

	lut_sub lut_4962 ({sk[1119], i_9_, i_7_, i_8_, i_6_, x507x}, n_n4671);
	defparam lut_4962.LUT_SIZE = 6;
	defparam lut_4962.mask = 64'h77ff77ff10000000;

	lut_sub lut_4964 ({sk[1120], x492x, x21x, x14x, x20x, x575x}, n_n4205);
	defparam lut_4964.LUT_SIZE = 6;
	defparam lut_4964.mask = 64'h77ff77ff11551f5f;

	lut_sub lut_4968 ({sk[1121], x11x, x18x, x557x, x577x, x537x}, n_n4161);
	defparam lut_4968.LUT_SIZE = 6;
	defparam lut_4968.mask = 64'h77ff77ff005f337f;

	lut_sub lut_4972 ({sk[1122], i_9_, i_1_, i_2_, i_0_, x549x}, n_n5082);
	defparam lut_4972.LUT_SIZE = 6;
	defparam lut_4972.mask = 64'h77ff77ff00000400;

	lut_sub lut_4974 ({sk[1123], i_9_, i_7_, i_8_, i_6_, x583x}, n_n4599);
	defparam lut_4974.LUT_SIZE = 6;
	defparam lut_4974.mask = 64'h77ff77ff40000000;

	lut_sub lut_4976 ({sk[1124], x10x, x23x, x581x, x583x}, x45x);
	defparam lut_4976.LUT_SIZE = 5;
	defparam lut_4976.mask = 32'h0fff0537;

	lut_sub lut_4979 ({sk[1125], i_9_, i_7_, i_8_, i_6_, n_n390, n_n509}, x13446x);
	defparam lut_4979.LUT_SIZE = 7;
	defparam lut_4979.mask = 128'h777f777f777f777f0001000001011001;

	lut_sub lut_4985 ({sk[1126], x14x, x570x, x23x, x587x, x575x}, n_n4204);
	defparam lut_4985.LUT_SIZE = 6;
	defparam lut_4985.mask = 64'h77ff77ff050537ff;

	lut_sub lut_4989 ({sk[1127], i_9_, i_7_, i_8_, i_6_, n_n325, n_n491}, x447x);
	defparam lut_4989.LUT_SIZE = 7;
	defparam lut_4989.mask = 128'h777f777f777f777f0010101000101010;

	lut_sub lut_4996 ({sk[1128], i_9_, i_7_, i_8_, i_6_, n_n325, n_n491}, n_n4070);
	defparam lut_4996.LUT_SIZE = 7;
	defparam lut_4996.mask = 128'h777f777f777f777f0110101001111010;

	lut_sub lut_5006 ({sk[1129], x25x, x510x, x14x, x511x}, x158x);
	defparam lut_5006.LUT_SIZE = 5;
	defparam lut_5006.mask = 32'h0fff0357;

	lut_sub lut_5009 ({sk[1130], i_9_, n_n325, x580x, x505x, x158x}, x13153x);
	defparam lut_5009.LUT_SIZE = 6;
	defparam lut_5009.mask = 64'h77ff77ff5555557f;

	lut_sub lut_5013 ({sk[1131], i_9_, i_7_, i_8_, i_6_, n_n473, n_n325}, x13154x);
	defparam lut_5013.LUT_SIZE = 7;
	defparam lut_5013.mask = 128'h777f777f777f777f0101010000010100;

	lut_sub lut_5019 ({sk[1132], x25x, x24x, x14x, x530x, x528x}, n_n4197);
	defparam lut_5019.LUT_SIZE = 6;
	defparam lut_5019.mask = 64'h77ff77ff05373737;

	lut_sub lut_5023 ({sk[1133], i_9_, i_7_, i_8_, i_6_, n_n325, n_n464}, x390x);
	defparam lut_5023.LUT_SIZE = 7;
	defparam lut_5023.mask = 128'h777f777f777f777f0001100001110000;

	lut_sub lut_5029 ({sk[1134], x22x, x14x, x516x, x511x, n_n4197, x390x}, x13166x);
	defparam lut_5029.LUT_SIZE = 7;
	defparam lut_5029.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_5034 ({sk[1135], x14x, x20x, x506x, x511x}, x395x);
	defparam lut_5034.LUT_SIZE = 5;
	defparam lut_5034.mask = 32'h0fff0537;

	lut_sub lut_5037 ({sk[1136], x11x, x14x, x522x, x530x}, x151x);
	defparam lut_5037.LUT_SIZE = 5;
	defparam lut_5037.mask = 32'h0fff0357;

	lut_sub lut_5040 ({sk[1137], i_9_, i_7_, i_8_, i_6_, n_n260, n_n535}, x13157x);
	defparam lut_5040.LUT_SIZE = 7;
	defparam lut_5040.mask = 128'h777f777f777f777f0101010001010001;

	lut_sub lut_5047 ({sk[1138], x21x, x14x, x488x, x511x}, x13160x);
	defparam lut_5047.LUT_SIZE = 5;
	defparam lut_5047.mask = 32'h0fff0357;

	lut_sub lut_5050 ({sk[1139], x22x, x14x, x23x, x503x, x530x, x389x}, x22189x);
	defparam lut_5050.LUT_SIZE = 7;
	defparam lut_5050.mask = 128'h777f777f777f777faa88a08088888080;

	lut_sub lut_5055 ({sk[1140], x395x, x151x, x13157x, x13160x, x22189x}, x13167x);
	defparam lut_5055.LUT_SIZE = 6;
	defparam lut_5055.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_5061 ({sk[1141], i_9_, i_7_, i_8_, i_6_, n_n518, n_n260}, n_n4063);
	defparam lut_5061.LUT_SIZE = 7;
	defparam lut_5061.mask = 128'h777f777f777f777f0111101000111010;

	lut_sub lut_5071 ({sk[1142], i_9_, x22x, n_n524, n_n260, n_n535, x535x}, x13178x);
	defparam lut_5071.LUT_SIZE = 7;
	defparam lut_5071.mask = 128'h777f777f777f777f0003030305070707;

	lut_sub lut_5076 ({sk[1143], x24x, x17x, x596x, x546x, x177x, n_n4837}, x22188x);
	defparam lut_5076.LUT_SIZE = 7;
	defparam lut_5076.mask = 128'h777f777f777f777f8888808088008000;

	lut_sub lut_5081 ({sk[1144], x13170x, x13171x, n_n4063, x13178x, x22188x}, n_n4009);
	defparam lut_5081.LUT_SIZE = 6;
	defparam lut_5081.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_5087 ({sk[1145], i_9_, i_7_, i_8_, i_6_, x588x}, x13183x);
	defparam lut_5087.LUT_SIZE = 6;
	defparam lut_5087.mask = 64'h77ff77ff04100000;

	lut_sub lut_5090 ({sk[1146], i_9_, i_7_, i_8_, i_6_, n_n482, n_n325}, x13184x);
	defparam lut_5090.LUT_SIZE = 7;
	defparam lut_5090.mask = 128'h777f777f777f777f0000101001000010;

	lut_sub lut_5095 ({sk[1147], n_n4204, n_n4070, x13153x, x13154x, x13183x, x13184x}, x13188x);
	defparam lut_5095.LUT_SIZE = 7;
	defparam lut_5095.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_5102 ({sk[1148], i_9_, i_7_, i_8_, i_6_, n_n260, n_n500}, x13193x);
	defparam lut_5102.LUT_SIZE = 7;
	defparam lut_5102.mask = 128'h777f777f777f777f0110000001001000;

	lut_sub lut_5107 ({sk[1149], i_9_, i_7_, i_8_, i_6_, n_n260, n_n491}, n_n4059);
	defparam lut_5107.LUT_SIZE = 7;
	defparam lut_5107.mask = 128'h777f777f777f777f0101011011111000;

	lut_sub lut_5117 ({sk[1150], i_9_, x25x, n_n482, n_n260, n_n520, x512x}, n_n1592);
	defparam lut_5117.LUT_SIZE = 7;
	defparam lut_5117.mask = 128'h777f777f777f777f0003555700035557;

	lut_sub lut_5121 ({sk[1151], i_9_, n_n526, n_n473, n_n260, x42x}, x13211x);
	defparam lut_5121.LUT_SIZE = 6;
	defparam lut_5121.mask = 64'h77ff77ff55575557;

	lut_sub lut_5125 ({sk[1152], x15x, x17x, x512x, x505x, n_n1592, x13211x}, x13213x);
	defparam lut_5125.LUT_SIZE = 7;
	defparam lut_5125.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_5130 ({sk[1153], i_9_, i_7_, i_8_, i_6_, n_n482, n_n260}, n_n4058);
	defparam lut_5130.LUT_SIZE = 7;
	defparam lut_5130.mask = 128'h777f777f777f777f0111110000101110;

	lut_sub lut_5140 ({sk[1154], i_9_, i_7_, i_8_, i_6_, n_n260, n_n464}, x13208x);
	defparam lut_5140.LUT_SIZE = 7;
	defparam lut_5140.mask = 128'h777f777f777f777f0100000100000101;

	lut_sub lut_5145 ({sk[1155], x24x, x17x, x502x, x531x}, x13206x);
	defparam lut_5145.LUT_SIZE = 5;
	defparam lut_5145.mask = 32'h0fff0357;

	lut_sub lut_5148 ({sk[1156], x17x, x522x, x180x, n_n4058, x13208x, x13206x}, x13214x);
	defparam lut_5148.LUT_SIZE = 7;
	defparam lut_5148.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_5154 ({sk[1157], i_9_, i_7_, i_8_, i_6_, n_n518, n_n195}, x137x);
	defparam lut_5154.LUT_SIZE = 7;
	defparam lut_5154.mask = 128'h777f777f777f777f0101011000010010;

	lut_sub lut_5161 ({sk[1158], i_9_, i_7_, i_8_, i_6_, n_n535, n_n195}, x13225x);
	defparam lut_5161.LUT_SIZE = 7;
	defparam lut_5161.mask = 128'h777f777f777f777f0011010010110000;

	lut_sub lut_5168 ({sk[1159], x137x, x13225x}, x13228x);
	defparam lut_5168.LUT_SIZE = 3;
	defparam lut_5168.mask = 8'h17;

	lut_sub lut_5171 ({sk[1160], x11x, x18x, x535x, x553x}, x210x);
	defparam lut_5171.LUT_SIZE = 5;
	defparam lut_5171.mask = 32'h0fff0357;

	lut_sub lut_5174 ({sk[1161], x22x, x21x, x17x, x516x, x531x}, n_n814);
	defparam lut_5174.LUT_SIZE = 6;
	defparam lut_5174.mask = 64'h77ff77ff03575757;

	lut_sub lut_5178 ({sk[1162], x18x, x20x, x550x, x23x, x549x, x531x}, x13223x);
	defparam lut_5178.LUT_SIZE = 7;
	defparam lut_5178.mask = 128'h777f777f777f777f0505555537ff77ff;

	lut_sub lut_5183 ({sk[1163], x25x, x17x, x23x, x489x, x553x, n_n4962}, x22187x);
	defparam lut_5183.LUT_SIZE = 7;
	defparam lut_5183.mask = 128'h777f777f777f777faa88a08088888080;

	lut_sub lut_5188 ({sk[1164], x68x, x210x, n_n814, x13223x, x22187x}, x13229x);
	defparam lut_5188.LUT_SIZE = 6;
	defparam lut_5188.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_5194 ({sk[1165], x17x, x20x, x484x, x562x, x461x, x13231x}, x13233x);
	defparam lut_5194.LUT_SIZE = 7;
	defparam lut_5194.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_5199 ({sk[1166], x17x, x536x, x13193x, n_n4059, n_n4889, x13192x}, x13234x);
	defparam lut_5199.LUT_SIZE = 7;
	defparam lut_5199.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_5205 ({sk[1167], i_9_, i_7_, i_8_, i_6_, n_n509, n_n325}, n_n4072);
	defparam lut_5205.LUT_SIZE = 7;
	defparam lut_5205.mask = 128'h777f777f777f777f1110011001111000;

	lut_sub lut_5215 ({sk[1168], i_9_, n_n534, n_n325, n_n491, x560x, x69x}, x11836x);
	defparam lut_5215.LUT_SIZE = 7;
	defparam lut_5215.mask = 128'h777f777f777f777f555555555577557f;

	lut_sub lut_5219 ({sk[1169], x14x, x482x, x23x, x581x, x595x}, x243x);
	defparam lut_5219.LUT_SIZE = 6;
	defparam lut_5219.mask = 64'h77ff77ff050537ff;

	lut_sub lut_5223 ({sk[1170], x25x, x21x, x14x, x490x, x585x, x595x}, x13251x);
	defparam lut_5223.LUT_SIZE = 7;
	defparam lut_5223.mask = 128'h777f777f777f777f003f557f557f557f;

	lut_sub lut_5228 ({sk[1171], x539x, x14x, x241x, x243x, x13251x}, x13254x);
	defparam lut_5228.LUT_SIZE = 6;
	defparam lut_5228.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_5233 ({sk[1172], x11x, x14x, x545x, x535x, x551x}, n_n4219);
	defparam lut_5233.LUT_SIZE = 6;
	defparam lut_5233.mask = 64'h77ff77ff003f557f;

	lut_sub lut_5237 ({sk[1173], x24x, x14x, x549x, x551x}, x221x);
	defparam lut_5237.LUT_SIZE = 5;
	defparam lut_5237.mask = 32'h0fff0357;

	lut_sub lut_5240 ({sk[1174], i_9_, i_7_, i_8_, i_6_, n_n325, n_n535}, x13249x);
	defparam lut_5240.LUT_SIZE = 7;
	defparam lut_5240.mask = 128'h777f777f777f777f0010001010001000;

	lut_sub lut_5245 ({sk[1175], i_9_, i_7_, i_8_, i_6_, n_n518, n_n325}, x13250x);
	defparam lut_5245.LUT_SIZE = 7;
	defparam lut_5245.mask = 128'h777f777f777f777f0000011000001100;

	lut_sub lut_5250 ({sk[1176], x14x, x23x, x548x, x526x, n_n4697, n_n4694}, x22186x);
	defparam lut_5250.LUT_SIZE = 7;
	defparam lut_5250.mask = 128'h777f777f777f777f8888808088008000;

	lut_sub lut_5255 ({sk[1177], n_n4219, x221x, x13249x, x13250x, x22186x}, x13255x);
	defparam lut_5255.LUT_SIZE = 6;
	defparam lut_5255.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_5261 ({sk[1178], i_9_, i_7_, i_8_, i_6_, n_n390, n_n464}, x13269x);
	defparam lut_5261.LUT_SIZE = 7;
	defparam lut_5261.mask = 128'h777f777f777f777f0111110000011110;

	lut_sub lut_5271 ({sk[1179], i_9_, i_7_, i_8_, i_6_, x565x, x575x}, x11835x);
	defparam lut_5271.LUT_SIZE = 7;
	defparam lut_5271.mask = 128'h777f777f777f777f3000050000000000;

	lut_sub lut_5274 ({sk[1180], i_9_, i_7_, i_8_, i_6_, n_n325, n_n500}, x13276x);
	defparam lut_5274.LUT_SIZE = 7;
	defparam lut_5274.mask = 128'h777f777f777f777f0101011001001111;

	lut_sub lut_5284 ({sk[1181], n_n4072, x11836x, n_n4210, x11835x, x13276x}, x13278x);
	defparam lut_5284.LUT_SIZE = 6;
	defparam lut_5284.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_5290 ({sk[1182], x22x, x21x, x20x, x582x, x312x, x22185x}, n_n4078);
	defparam lut_5290.LUT_SIZE = 7;
	defparam lut_5290.mask = 128'h777f777f777f777fbbbfbfbfbfbfbfbf;

	lut_sub lut_5296 ({sk[1183], x10x, x505x, x529x, n_n4671, x80x, x13263x}, n_n4077);
	defparam lut_5296.LUT_SIZE = 7;
	defparam lut_5296.mask = 128'h777f777f777f777f7f7f7f7f7fffffff;

	lut_sub lut_5302 ({sk[1184], i_9_, i_7_, i_8_, i_6_, x532x}, n_n5079);
	defparam lut_5302.LUT_SIZE = 6;
	defparam lut_5302.mask = 64'h77ff77ff40000000;

	lut_sub lut_5304 ({sk[1185], i_9_, i_1_, i_2_, i_0_, x525x}, n_n5078);
	defparam lut_5304.LUT_SIZE = 6;
	defparam lut_5304.mask = 64'h77ff77ff00000040;

	lut_sub lut_5306 ({sk[1186], x15x, x12x, x554x, x548x}, x123x);
	defparam lut_5306.LUT_SIZE = 5;
	defparam lut_5306.mask = 32'h0fff0537;

	lut_sub lut_5309 ({sk[1187], i_9_, i_1_, i_2_, i_0_, x535x, x525x}, x14642x);
	defparam lut_5309.LUT_SIZE = 7;
	defparam lut_5309.mask = 128'h777f777f777f777f0000000000305000;

	lut_sub lut_5312 ({sk[1188], x21x, x18x, x23x, x489x, n_n5081, x532x}, x22162x);
	defparam lut_5312.LUT_SIZE = 7;
	defparam lut_5312.mask = 128'h777f777f777f777fcc88c08088888080;

	lut_sub lut_5317 ({sk[1189], i_9_, i_7_, i_8_, i_6_, x598x}, x122x);
	defparam lut_5317.LUT_SIZE = 6;
	defparam lut_5317.mask = 64'h77ff77ff01100000;

	lut_sub lut_5320 ({sk[1190], x21x, x12x, x554x, x517x}, x232x);
	defparam lut_5320.LUT_SIZE = 5;
	defparam lut_5320.mask = 32'h0fff0537;

	lut_sub lut_5323 ({sk[1191], i_9_, i_7_, i_8_, i_6_, x554x}, x14646x);
	defparam lut_5323.LUT_SIZE = 6;
	defparam lut_5323.mask = 64'h77ff77ff04040000;

	lut_sub lut_5326 ({sk[1192], x18x, x23x, x502x, x513x, x527x, x528x}, x22309x);
	defparam lut_5326.LUT_SIZE = 7;
	defparam lut_5326.mask = 128'h777f777f777f777ffffff0f088008000;

	lut_sub lut_5331 ({sk[1193], x25x, x19x, x564x, x569x}, x433x);
	defparam lut_5331.LUT_SIZE = 5;
	defparam lut_5331.mask = 32'h0fff0357;

	lut_sub lut_5334 ({sk[1194], x515x, x19x, x24x, x518x}, x14242x);
	defparam lut_5334.LUT_SIZE = 5;
	defparam lut_5334.mask = 32'h0fff0537;

	lut_sub lut_5337 ({sk[1195], x592x, x19x, x11x, x586x}, x14243x);
	defparam lut_5337.LUT_SIZE = 5;
	defparam lut_5337.mask = 32'h0fff0537;

	lut_sub lut_5340 ({sk[1196], x21x, x579x, x433x, x63x, x14242x, x14243x}, n_n3551);
	defparam lut_5340.LUT_SIZE = 7;
	defparam lut_5340.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_5346 ({sk[1197], i_5_, i_3_, i_4_, x25x, x11x, n_n260}, x14261x);
	defparam lut_5346.LUT_SIZE = 7;
	defparam lut_5346.mask = 128'h777f777f777f777f0000110500110005;

	lut_sub lut_5351 ({sk[1198], x21x, x17x, x20x, x484x, x478x, x566x}, x14260x);
	defparam lut_5351.LUT_SIZE = 7;
	defparam lut_5351.mask = 128'h777f777f777f777f000f333f555f777f;

	lut_sub lut_5355 ({sk[1199], x24x, x17x, x490x, x576x, x14261x, x14260x}, n_n3558);
	defparam lut_5355.LUT_SIZE = 7;
	defparam lut_5355.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_5360 ({sk[1200], x21x, x17x, x553x, x493x}, x14264x);
	defparam lut_5360.LUT_SIZE = 5;
	defparam lut_5360.mask = 32'h0fff0537;

	lut_sub lut_5363 ({sk[1201], x15x, x17x, x597x, x586x, x587x}, x14266x);
	defparam lut_5363.LUT_SIZE = 6;
	defparam lut_5363.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_5367 ({sk[1202], x25x, x17x, x545x, x18x, x512x, x489x}, x22298x);
	defparam lut_5367.LUT_SIZE = 7;
	defparam lut_5367.mask = 128'h777f777f777f777ffff0aaa0ccc08880;

	lut_sub lut_5376 ({sk[1203], x20x, x512x, x14264x, x14266x, x22298x}, n_n3557);
	defparam lut_5376.LUT_SIZE = 6;
	defparam lut_5376.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_5381 ({sk[1204], x15x, x19x, x474x, x472x, x529x, x534x}, x14252x);
	defparam lut_5381.LUT_SIZE = 7;
	defparam lut_5381.mask = 128'h777f777f777f777f00003fff55557fff;

	lut_sub lut_5386 ({sk[1205], x19x, x22x, x539x, x23x, x487x, x548x}, x14253x);
	defparam lut_5386.LUT_SIZE = 7;
	defparam lut_5386.mask = 128'h777f777f777f777f0303333357ff77ff;

	lut_sub lut_5391 ({sk[1206], x19x, x20x, x508x, x517x, x599x, x593x}, x14254x);
	defparam lut_5391.LUT_SIZE = 7;
	defparam lut_5391.mask = 128'h777f777f777f777f000033335fff7fff;

	lut_sub lut_5396 ({sk[1207], x22x, x18x, x513x, x559x, x14272x, x14273x}, x14275x);
	defparam lut_5396.LUT_SIZE = 7;
	defparam lut_5396.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_5401 ({sk[1208], n_n3551, x14252x, x14253x, x14254x, x14275x}, x14277x);
	defparam lut_5401.LUT_SIZE = 6;
	defparam lut_5401.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_5407 ({sk[1209], x25x, x22x, x24x, x578x, x168x, x22150x}, n_n3554);
	defparam lut_5407.LUT_SIZE = 7;
	defparam lut_5407.mask = 128'h777f777f777f777fbbbfbfbfbfbfbfbf;

	lut_sub lut_5413 ({sk[1210], x22x, x591x, x14230x, x14231x, x22273x}, n_n3553);
	defparam lut_5413.LUT_SIZE = 6;
	defparam lut_5413.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_5418 ({sk[1211], x25x, x12x, x490x, x581x, x598x, x585x}, x14238x);
	defparam lut_5418.LUT_SIZE = 7;
	defparam lut_5418.mask = 128'h777f777f777f777f00005fff33337fff;

	lut_sub lut_5423 ({sk[1212], i_9_, i_7_, i_8_, i_6_, x554x, x532x}, x14239x);
	defparam lut_5423.LUT_SIZE = 7;
	defparam lut_5423.mask = 128'h777f777f777f777f0750050500000000;

	lut_sub lut_5429 ({sk[1213], n_n3558, n_n3557, n_n3554, n_n3553, x14238x, x14239x}, x14278x);
	defparam lut_5429.LUT_SIZE = 7;
	defparam lut_5429.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_5436 ({sk[1214], i_9_, n_n518, x21x, n_n526, n_n455, x540x}, x14283x);
	defparam lut_5436.LUT_SIZE = 7;
	defparam lut_5436.mask = 128'h777f777f777f777f0555057700550377;

	lut_sub lut_5441 ({sk[1215], x15x, x16x, x539x, x11x, x497x, x563x}, x14290x);
	defparam lut_5441.LUT_SIZE = 7;
	defparam lut_5441.mask = 128'h777f777f777f777f030357ff333377ff;

	lut_sub lut_5446 ({sk[1216], x25x, x21x, x10x, x479x, x583x, x481x}, x14307x);
	defparam lut_5446.LUT_SIZE = 7;
	defparam lut_5446.mask = 128'h777f777f777f777f005533770f5f3f7f;

	lut_sub lut_5450 ({sk[1217], x10x, x20x, x550x, x547x, x546x, x559x}, x14308x);
	defparam lut_5450.LUT_SIZE = 7;
	defparam lut_5450.mask = 128'h777f777f777f777f00000f0f77ff7fff;

	lut_sub lut_5455 ({sk[1218], x21x, x10x, x475x, x547x, x14307x, x14308x}, x14310x);
	defparam lut_5455.LUT_SIZE = 7;
	defparam lut_5455.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_5460 ({sk[1219], x25x, x14x, x586x, x511x}, x14327x);
	defparam lut_5460.LUT_SIZE = 5;
	defparam lut_5460.mask = 32'h0fff0357;

	lut_sub lut_5463 ({sk[1220], x538x, x21x, x14x, x588x, x584x}, x14329x);
	defparam lut_5463.LUT_SIZE = 6;
	defparam lut_5463.mask = 64'h77ff77ff05370f3f;

	lut_sub lut_5467 ({sk[1221], x24x, x14x, x23x, x565x, x536x, x530x}, x22291x);
	defparam lut_5467.LUT_SIZE = 7;
	defparam lut_5467.mask = 128'h777f777f777f777ffff0ccc0aaa08880;

	lut_sub lut_5476 ({sk[1222], x24x, x565x, x14327x, x14329x, x22291x}, x14332x);
	defparam lut_5476.LUT_SIZE = 6;
	defparam lut_5476.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_5481 ({sk[1223], x21x, x14x, x519x, x20x, x575x}, n_n3469);
	defparam lut_5481.LUT_SIZE = 6;
	defparam lut_5481.mask = 64'h77ff77ff111f555f;

	lut_sub lut_5485 ({sk[1224], x18x, x20x, x491x, x560x, x567x}, n_n3427);
	defparam lut_5485.LUT_SIZE = 6;
	defparam lut_5485.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_5489 ({sk[1225], x15x, x12x, x572x, x578x}, x76x);
	defparam lut_5489.LUT_SIZE = 5;
	defparam lut_5489.mask = 32'h0fff0357;

	lut_sub lut_5492 ({sk[1226], i_9_, i_7_, i_8_, i_6_, n_n491, n_n130}, n_n3305);
	defparam lut_5492.LUT_SIZE = 7;
	defparam lut_5492.mask = 128'h777f777f777f777f0011011011011010;

	lut_sub lut_5502 ({sk[1227], x521x, x21x, x18x, x597x}, x57x);
	defparam lut_5502.LUT_SIZE = 5;
	defparam lut_5502.mask = 32'h0fff0537;

	lut_sub lut_5505 ({sk[1228], i_9_, i_7_, i_8_, i_6_, n_n518, n_n195}, x13833x);
	defparam lut_5505.LUT_SIZE = 7;
	defparam lut_5505.mask = 128'h777f777f777f777f1010000010000010;

	lut_sub lut_5510 ({sk[1229], x18x, x490x, x20x, x553x, x546x}, n_n4172);
	defparam lut_5510.LUT_SIZE = 6;
	defparam lut_5510.mask = 64'h77ff77ff030357ff;

	lut_sub lut_5514 ({sk[1230], i_9_, i_7_, i_8_, i_6_, n_n518, n_n195}, x13836x);
	defparam lut_5514.LUT_SIZE = 7;
	defparam lut_5514.mask = 128'h777f777f777f777f0100000100000101;

	lut_sub lut_5519 ({sk[1231], x21x, x18x, x517x, x553x}, x342x);
	defparam lut_5519.LUT_SIZE = 5;
	defparam lut_5519.mask = 32'h0fff0357;

	lut_sub lut_5522 ({sk[1232], x15x, x24x, x18x, x597x, x553x, x559x}, x22293x);
	defparam lut_5522.LUT_SIZE = 7;
	defparam lut_5522.mask = 128'h777f777f777f777fffaaf0a0cc88c080;

	lut_sub lut_5531 ({sk[1233], x17x, x489x, n_n4172, x13836x, x22293x}, x13843x);
	defparam lut_5531.LUT_SIZE = 6;
	defparam lut_5531.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_5536 ({sk[1234], i_9_, i_7_, i_8_, i_6_, x531x, x342x}, x13840x);
	defparam lut_5536.LUT_SIZE = 7;
	defparam lut_5536.mask = 128'h777f777f777f777f5575755555555555;

	lut_sub lut_5540 ({sk[1235], x25x, x18x, x482x, x485x, x480x, x57x}, x22176x);
	defparam lut_5540.LUT_SIZE = 7;
	defparam lut_5540.mask = 128'h777f777f777f777faaaa8800a0a08000;

	lut_sub lut_5545 ({sk[1236], n_n3803, x13833x, x13840x, x22176x}, x13844x);
	defparam lut_5545.LUT_SIZE = 5;
	defparam lut_5545.mask = 32'h0fffbfff;

	lut_sub lut_5550 ({sk[1237], i_9_, i_7_, i_8_, i_6_, n_n518, n_n455}, x14122x);
	defparam lut_5550.LUT_SIZE = 7;
	defparam lut_5550.mask = 128'h777f777f777f777f0100001100011000;

	lut_sub lut_5556 ({sk[1238], x13x, x544x, x20x, x581x}, x194x);
	defparam lut_5556.LUT_SIZE = 5;
	defparam lut_5556.mask = 32'h0fff0357;

	lut_sub lut_5559 ({sk[1239], x21x, x13x, x564x, x476x}, x14124x);
	defparam lut_5559.LUT_SIZE = 5;
	defparam lut_5559.mask = 32'h0fff0357;

	lut_sub lut_5562 ({sk[1240], i_9_, i_7_, i_8_, i_6_, n_n455, n_n509}, x14129x);
	defparam lut_5562.LUT_SIZE = 7;
	defparam lut_5562.mask = 128'h777f777f777f777f0101001001001010;

	lut_sub lut_5569 ({sk[1241], x13x, x544x, x23x, x563x, x14124x, x14129x}, x14131x);
	defparam lut_5569.LUT_SIZE = 7;
	defparam lut_5569.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_5574 ({sk[1242], x13x, x23x, x540x, x546x}, x128x);
	defparam lut_5574.LUT_SIZE = 5;
	defparam lut_5574.mask = 32'h0fff0357;

	lut_sub lut_5577 ({sk[1243], i_9_, i_7_, i_8_, i_6_, x544x}, x291x);
	defparam lut_5577.LUT_SIZE = 6;
	defparam lut_5577.mask = 64'h77ff77ff01100000;

	lut_sub lut_5580 ({sk[1244], i_9_, i_7_, i_8_, i_6_, x544x, x541x}, x14123x);
	defparam lut_5580.LUT_SIZE = 7;
	defparam lut_5580.mask = 128'h777f777f777f777f0000300500000000;

	lut_sub lut_5583 ({sk[1245], n_n455, x13x, x24x, n_n509, n_n500, n_n530}, x14126x);
	defparam lut_5583.LUT_SIZE = 7;
	defparam lut_5583.mask = 128'h777f777f777f777f00001515003f153f;

	lut_sub lut_5588 ({sk[1246], x14122x, x194x, x128x, x291x, x14123x, x14126x}, x14132x);
	defparam lut_5588.LUT_SIZE = 7;
	defparam lut_5588.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_5595 ({sk[1247], i_9_, i_7_, i_8_, i_6_, x495x}, n_n4421);
	defparam lut_5595.LUT_SIZE = 6;
	defparam lut_5595.mask = 64'h77ff77ff04000000;

	lut_sub lut_5597 ({sk[1248], i_9_, i_7_, i_8_, i_6_, n_n455, n_n535}, x14145x);
	defparam lut_5597.LUT_SIZE = 7;
	defparam lut_5597.mask = 128'h777f777f777f777f0001001001011010;

	lut_sub lut_5604 ({sk[1249], x20x, x23x, x495x, n_n3520, x14145x}, x14147x);
	defparam lut_5604.LUT_SIZE = 6;
	defparam lut_5604.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_5609 ({sk[1250], x25x, x16x, x506x, x529x, x496x}, x14142x);
	defparam lut_5609.LUT_SIZE = 6;
	defparam lut_5609.mask = 64'h77ff77ff003f557f;

	lut_sub lut_5613 ({sk[1251], i_9_, n_n536, n_n532, x488x, n_n464, x524x}, x14143x);
	defparam lut_5613.LUT_SIZE = 7;
	defparam lut_5613.mask = 128'h777f777f777f777f0000003300005f7f;

	lut_sub lut_5618 ({sk[1252], x16x, x11x, x516x, x522x, x496x, n_n4441}, x22166x);
	defparam lut_5618.LUT_SIZE = 7;
	defparam lut_5618.mask = 128'h777f777f777f777faaaa8888a0008000;

	lut_sub lut_5623 ({sk[1253], x16x, x21x, x23x, x496x, x489x, x421x}, x22340x);
	defparam lut_5623.LUT_SIZE = 7;
	defparam lut_5623.mask = 128'h777f777f777f777faaa0a0a088808080;

	lut_sub lut_5628 ({sk[1254], x14142x, x14143x, x22166x, x22340x}, x14148x);
	defparam lut_5628.LUT_SIZE = 5;
	defparam lut_5628.mask = 32'h0fffefff;

	lut_sub lut_5633 ({sk[1255], i_9_, i_7_, i_8_, i_6_, x501x}, n_n4331);
	defparam lut_5633.LUT_SIZE = 6;
	defparam lut_5633.mask = 64'h77ff77ff00100000;

	lut_sub lut_5635 ({sk[1256], x521x, x21x, x13x, x544x, x494x}, n_n3162);
	defparam lut_5635.LUT_SIZE = 6;
	defparam lut_5635.mask = 64'h77ff77ff05370f3f;

	lut_sub lut_5639 ({sk[1257], x10x, x478x, x23x, x479x, x564x}, n_n4232);
	defparam lut_5639.LUT_SIZE = 6;
	defparam lut_5639.mask = 64'h77ff77ff030357ff;

	lut_sub lut_5643 ({sk[1258], x10x, x474x, x20x, x479x}, x272x);
	defparam lut_5643.LUT_SIZE = 5;
	defparam lut_5643.mask = 32'h0fff111f;

	lut_sub lut_5646 ({sk[1259], x25x, x11x, x10x, x561x, x479x, x563x}, x22326x);
	defparam lut_5646.LUT_SIZE = 7;
	defparam lut_5646.mask = 128'h777f777f777f777fffaacc88f0a0c080;

	lut_sub lut_5655 ({sk[1260], i_9_, i_7_, i_8_, i_6_, n_n482, n_n195}, n_n2957);
	defparam lut_5655.LUT_SIZE = 7;
	defparam lut_5655.mask = 128'h777f777f777f777f0111101001101010;

	lut_sub lut_5665 ({sk[1261], i_9_, i_7_, i_8_, i_6_, n_n473, n_n325}, x14918x);
	defparam lut_5665.LUT_SIZE = 7;
	defparam lut_5665.mask = 128'h777f777f777f777f0000010101100000;

	lut_sub lut_5670 ({sk[1262], i_9_, i_7_, i_8_, i_6_, n_n482, n_n325}, x14922x);
	defparam lut_5670.LUT_SIZE = 7;
	defparam lut_5670.mask = 128'h777f777f777f777f0010101000100000;

	lut_sub lut_5675 ({sk[1263], n_n526, n_n482, x11x, n_n325, x14x, x151x}, x14923x);
	defparam lut_5675.LUT_SIZE = 7;
	defparam lut_5675.mask = 128'h777f777f777f777f5555555f5555777f;

	lut_sub lut_5679 ({sk[1264], x15x, x11x, x14x, x502x, x511x, x440x}, x22147x);
	defparam lut_5679.LUT_SIZE = 7;
	defparam lut_5679.mask = 128'h777f777f777f777faaa0888088808880;

	lut_sub lut_5684 ({sk[1265], i_9_, i_7_, i_8_, i_6_, n_n473, n_n260}, x14948x);
	defparam lut_5684.LUT_SIZE = 7;
	defparam lut_5684.mask = 128'h777f777f777f777f0100010100010000;

	lut_sub lut_5689 ({sk[1266], x11x, x17x, x519x, x23x, x584x, x576x}, x14954x);
	defparam lut_5689.LUT_SIZE = 7;
	defparam lut_5689.mask = 128'h777f777f777f777f050537ff555577ff;

	lut_sub lut_5694 ({sk[1267], x25x, x17x, x586x, x589x}, x14952x);
	defparam lut_5694.LUT_SIZE = 5;
	defparam lut_5694.mask = 32'h0fff0357;

	lut_sub lut_5697 ({sk[1268], x492x, x17x, x570x, x537x}, x14953x);
	defparam lut_5697.LUT_SIZE = 5;
	defparam lut_5697.mask = 32'h0fff070f;

	lut_sub lut_5701 ({sk[1269], x21x, x17x, x512x, x505x, x502x, x105x}, x22144x);
	defparam lut_5701.LUT_SIZE = 7;
	defparam lut_5701.mask = 128'h777f777f777f777faaaa8080aa008000;

	lut_sub lut_5706 ({sk[1270], i_9_, i_7_, i_8_, i_6_, n_n260, n_n464}, x14972x);
	defparam lut_5706.LUT_SIZE = 7;
	defparam lut_5706.mask = 128'h777f777f777f777f0101001001010010;

	lut_sub lut_5713 ({sk[1271], x21x, x17x, x516x, x529x, x531x, x489x}, x22269x);
	defparam lut_5713.LUT_SIZE = 7;
	defparam lut_5713.mask = 128'h777f777f777f777fffffa000cccc8000;

	lut_sub lut_5718 ({sk[1272], i_9_, i_7_, i_8_, i_6_, n_n535, n_n195}, n_n2591);
	defparam lut_5718.LUT_SIZE = 7;
	defparam lut_5718.mask = 128'h777f777f777f777f0101010101110110;

	lut_sub lut_5728 ({sk[1273], x25x, x17x, x20x, x531x, n_n4952, x525x}, x22143x);
	defparam lut_5728.LUT_SIZE = 7;
	defparam lut_5728.mask = 128'h777f777f777f777fccc08880c0c08080;

	lut_sub lut_5733 ({sk[1274], x21x, x483x, x14x, x20x, x564x, x563x}, x14985x);
	defparam lut_5733.LUT_SIZE = 7;
	defparam lut_5733.mask = 128'h777f777f777f777f00770f7f0077ffff;

	lut_sub lut_5738 ({sk[1275], i_9_, i_7_, i_8_, i_6_, n_n325, n_n491}, x14991x);
	defparam lut_5738.LUT_SIZE = 7;
	defparam lut_5738.mask = 128'h777f777f777f777f0101001100000010;

	lut_sub lut_5744 ({sk[1276], x10x, x24x, x527x, x526x}, x426x);
	defparam lut_5744.LUT_SIZE = 5;
	defparam lut_5744.mask = 32'h0fff0537;

	lut_sub lut_5747 ({sk[1277], i_9_, i_1_, i_2_, i_0_, x522x, x549x}, x14997x);
	defparam lut_5747.LUT_SIZE = 7;
	defparam lut_5747.mask = 128'h777f777f777f777f0000000005030000;

	lut_sub lut_5750 ({sk[1278], x11x, x10x, x529x, x526x}, x14998x);
	defparam lut_5750.LUT_SIZE = 5;
	defparam lut_5750.mask = 32'h0fff0357;

	lut_sub lut_5753 ({sk[1279], i_9_, n_n390, n_n520, n_n464, x86x}, x14999x);
	defparam lut_5753.LUT_SIZE = 6;
	defparam lut_5753.mask = 64'h77ff77ff55555557;

	lut_sub lut_5756 ({sk[1280], x15x, x10x, x524x, x526x}, x219x);
	defparam lut_5756.LUT_SIZE = 5;
	defparam lut_5756.mask = 32'h0fff0357;

	lut_sub lut_5759 ({sk[1281], i_9_, i_7_, i_8_, i_6_, n_n390, n_n473}, n_n2614);
	defparam lut_5759.LUT_SIZE = 7;
	defparam lut_5759.mask = 128'h777f777f777f777f0111100001111100;

	lut_sub lut_5769 ({sk[1282], x10x, x507x, x23x, x506x}, x417x);
	defparam lut_5769.LUT_SIZE = 5;
	defparam lut_5769.mask = 32'h0fff0357;

	lut_sub lut_5772 ({sk[1283], i_9_, i_7_, i_8_, i_6_, x526x}, x445x);
	defparam lut_5772.LUT_SIZE = 6;
	defparam lut_5772.mask = 64'h77ff77ff04400000;

	lut_sub lut_5775 ({sk[1284], x15x, x14x, x548x, x551x}, x442x);
	defparam lut_5775.LUT_SIZE = 5;
	defparam lut_5775.mask = 32'h0fff0357;

	lut_sub lut_5778 ({sk[1285], x25x, x24x, x483x, x14x, x477x}, n_n856);
	defparam lut_5778.LUT_SIZE = 6;
	defparam lut_5778.mask = 64'h77ff77ff111f1f1f;

	lut_sub lut_5782 ({sk[1286], i_9_, i_7_, i_8_, i_6_, n_n325, n_n535}, n_n2611);
	defparam lut_5782.LUT_SIZE = 7;
	defparam lut_5782.mask = 128'h777f777f777f777f1110101011001010;

	lut_sub lut_5792 ({sk[1287], i_9_, x22x, n_n524, n_n509, n_n325, x595x}, x15011x);
	defparam lut_5792.LUT_SIZE = 7;
	defparam lut_5792.mask = 128'h777f777f777f777f0055035700030303;

	lut_sub lut_5796 ({sk[1288], x22x, x521x, x14x, x475x, x594x, x595x}, x15012x);
	defparam lut_5796.LUT_SIZE = 7;
	defparam lut_5796.mask = 128'h777f777f777f777f003f00ff557f55ff;

	lut_sub lut_5801 ({sk[1289], i_9_, i_7_, i_8_, i_6_, n_n518, n_n325}, x15013x);
	defparam lut_5801.LUT_SIZE = 7;
	defparam lut_5801.mask = 128'h777f777f777f777f0001000101010010;

	lut_sub lut_5807 ({sk[1290], i_9_, i_1_, i_2_, i_0_, x585x}, n_n4972);
	defparam lut_5807.LUT_SIZE = 6;
	defparam lut_5807.mask = 64'h77ff77ff00000040;

	lut_sub lut_5809 ({sk[1291], i_9_, i_7_, i_8_, i_6_, x592x}, n_n5295);
	defparam lut_5809.LUT_SIZE = 6;
	defparam lut_5809.mask = 64'h77ff77ff10000000;

	lut_sub lut_5811 ({sk[1292], x13x, x509x, x510x, x508x}, n_n889);
	defparam lut_5811.LUT_SIZE = 5;
	defparam lut_5811.mask = 32'h0fff007f;

	lut_sub lut_5815 ({sk[1293], x13x, x20x, x23x, x493x, x543x}, x22324x);
	defparam lut_5815.LUT_SIZE = 6;
	defparam lut_5815.mask = 64'h77ff77fffaaac888;

	lut_sub lut_5820 ({sk[1294], i_9_, i_1_, i_2_, i_0_, x506x}, n_n4678);
	defparam lut_5820.LUT_SIZE = 6;
	defparam lut_5820.mask = 64'h77ff77ff00000100;

	lut_sub lut_5822 ({sk[1295], x15x, x10x, x507x, x505x}, x338x);
	defparam lut_5822.LUT_SIZE = 5;
	defparam lut_5822.mask = 32'h0fff0537;

	lut_sub lut_5825 ({sk[1296], x11x, x12x, x477x, x486x}, x414x);
	defparam lut_5825.LUT_SIZE = 5;
	defparam lut_5825.mask = 32'h0fff0357;

	lut_sub lut_5828 ({sk[1297], i_9_, i_7_, i_8_, i_6_, x598x, x486x}, x16720x);
	defparam lut_5828.LUT_SIZE = 7;
	defparam lut_5828.mask = 128'h777f777f777f777f3000000500000000;

	lut_sub lut_5831 ({sk[1298], x24x, x12x, x482x, x581x, x486x}, x16722x);
	defparam lut_5831.LUT_SIZE = 6;
	defparam lut_5831.mask = 64'h77ff77ff003f557f;

	lut_sub lut_5835 ({sk[1299], x12x, x481x, x480x, x414x, x16720x, x16722x}, n_n2209);
	defparam lut_5835.LUT_SIZE = 7;
	defparam lut_5835.mask = 128'h777f777f777f777f7f7f7f7f7fffffff;

	lut_sub lut_5841 ({sk[1300], x15x, x16x, x498x, x562x, x556x}, n_n4275);
	defparam lut_5841.LUT_SIZE = 6;
	defparam lut_5841.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_5845 ({sk[1301], i_9_, i_1_, i_2_, i_0_, x564x, x563x}, x345x);
	defparam lut_5845.LUT_SIZE = 7;
	defparam lut_5845.mask = 128'h777f777f777f777f0000000000000007;

	lut_sub lut_5848 ({sk[1302], i_9_, i_7_, i_8_, i_6_, x544x}, n_n4465);
	defparam lut_5848.LUT_SIZE = 6;
	defparam lut_5848.mask = 64'h77ff77ff00040000;

	lut_sub lut_5850 ({sk[1303], i_9_, i_7_, i_8_, i_6_, x476x}, x199x);
	defparam lut_5850.LUT_SIZE = 6;
	defparam lut_5850.mask = 64'h77ff77ff10040000;

	lut_sub lut_5853 ({sk[1304], x17x, x570x, x482x, x557x, x581x}, x16784x);
	defparam lut_5853.LUT_SIZE = 6;
	defparam lut_5853.mask = 64'h77ff77ff00007fff;

	lut_sub lut_5858 ({sk[1305], i_9_, x15x, n_n482, n_n532, n_n260, x576x}, x16783x);
	defparam lut_5858.LUT_SIZE = 7;
	defparam lut_5858.mask = 128'h777f777f777f777f0003555700035557;

	lut_sub lut_5862 ({sk[1306], x12x, x20x, x560x, x568x}, x126x);
	defparam lut_5862.LUT_SIZE = 5;
	defparam lut_5862.mask = 32'h0fff0537;

	lut_sub lut_5865 ({sk[1307], x22x, x12x, x573x, x568x}, x16793x);
	defparam lut_5865.LUT_SIZE = 5;
	defparam lut_5865.mask = 32'h0fff0357;

	lut_sub lut_5868 ({sk[1308], x538x, x12x, x20x, x560x, x568x}, x16795x);
	defparam lut_5868.LUT_SIZE = 6;
	defparam lut_5868.mask = 64'h77ff77ff053705ff;

	lut_sub lut_5872 ({sk[1309], x21x, x24x, x12x, x505x, x486x, x568x}, x22328x);
	defparam lut_5872.LUT_SIZE = 7;
	defparam lut_5872.mask = 128'h777f777f777f777ffff0aaa0ccc08880;

	lut_sub lut_5881 ({sk[1310], x25x, x533x, x16793x, x16795x, x22328x}, n_n2091);
	defparam lut_5881.LUT_SIZE = 6;
	defparam lut_5881.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_5886 ({sk[1311], x15x, x11x, x597x, x20x, x485x, x567x}, x22064x);
	defparam lut_5886.LUT_SIZE = 7;
	defparam lut_5886.mask = 128'h777f777f777f777ffff0cc00aa008800;

	lut_sub lut_5892 ({sk[1312], x18x, x472x, x475x, x564x}, x22332x);
	defparam lut_5892.LUT_SIZE = 5;
	defparam lut_5892.mask = 32'h0fffff80;

	lut_sub lut_5895 ({sk[1313], x15x, x553x, x22064x, x22332x}, x16805x);
	defparam lut_5895.LUT_SIZE = 5;
	defparam lut_5895.mask = 32'h0fffeeef;

	lut_sub lut_5899 ({sk[1314], i_9_, i_7_, i_8_, i_6_, x479x}, n_n4603);
	defparam lut_5899.LUT_SIZE = 6;
	defparam lut_5899.mask = 64'h77ff77ff00100000;

	lut_sub lut_5901 ({sk[1315], x10x, x24x, x482x, x479x, x480x}, n_n2037);
	defparam lut_5901.LUT_SIZE = 6;
	defparam lut_5901.mask = 64'h77ff77ff00335f7f;

	lut_sub lut_5905 ({sk[1316], i_9_, i_7_, i_8_, i_6_, n_n518, n_n390}, x16038x);
	defparam lut_5905.LUT_SIZE = 7;
	defparam lut_5905.mask = 128'h777f777f777f777f1100000010000010;

	lut_sub lut_5910 ({sk[1317], i_9_, i_7_, i_8_, i_6_, n_n473, n_n195}, x12310x);
	defparam lut_5910.LUT_SIZE = 7;
	defparam lut_5910.mask = 128'h777f777f777f777f0100100000100010;

	lut_sub lut_5915 ({sk[1318], i_9_, i_7_, i_8_, i_6_, n_n491, n_n130}, n_n1443);
	defparam lut_5915.LUT_SIZE = 7;
	defparam lut_5915.mask = 128'h777f777f777f777f1111100011001010;

	lut_sub lut_5925 ({sk[1319], x592x, x19x, x22x, x520x}, x424x);
	defparam lut_5925.LUT_SIZE = 5;
	defparam lut_5925.mask = 32'h0fff0537;

	lut_sub lut_5928 ({sk[1320], i_9_, i_7_, i_8_, i_6_, n_n482, n_n65}, n_n1432);
	defparam lut_5928.LUT_SIZE = 7;
	defparam lut_5928.mask = 128'h777f777f777f777f0101011100011101;

	lut_sub lut_5938 ({sk[1321], x492x, x21x, x18x, x20x, x557x, x590x}, x12117x);
	defparam lut_5938.LUT_SIZE = 7;
	defparam lut_5938.mask = 128'h777f777f777f777f0537557705ff55ff;

	lut_sub lut_5943 ({sk[1322], x22x, x510x, x18x, x577x, x567x}, x12116x);
	defparam lut_5943.LUT_SIZE = 6;
	defparam lut_5943.mask = 64'h77ff77ff000f777f;

	lut_sub lut_5947 ({sk[1323], x15x, x22x, x513x, x12117x, x12116x}, n_n1332);
	defparam lut_5947.LUT_SIZE = 6;
	defparam lut_5947.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_5952 ({sk[1324], x15x, x24x, x597x, x485x, x567x, n_n4972}, x22221x);
	defparam lut_5952.LUT_SIZE = 7;
	defparam lut_5952.mask = 128'h777f777f777f777faaaaa00088888000;

	lut_sub lut_5957 ({sk[1325], x18x, x549x, x494x, x559x, x68x, x22221x}, n_n1333);
	defparam lut_5957.LUT_SIZE = 7;
	defparam lut_5957.mask = 128'h777f777f777f777fbbbbbbbbbfffffff;

	lut_sub lut_5963 ({sk[1326], x12089x, x12088x, x12127x, x22220x}, x12129x);
	defparam lut_5963.LUT_SIZE = 5;
	defparam lut_5963.mask = 32'h0fffbfff;

	lut_sub lut_5968 ({sk[1327], n_n1330, n_n1331, x12110x, n_n1332, n_n1333, x12129x}, n_n1321);
	defparam lut_5968.LUT_SIZE = 7;
	defparam lut_5968.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_5975 ({sk[1328], i_9_, i_7_, i_8_, i_6_, x568x}, n_n5139);
	defparam lut_5975.LUT_SIZE = 6;
	defparam lut_5975.mask = 64'h77ff77ff00400000;

	lut_sub lut_5977 ({sk[1329], x515x, x15x, x19x, x508x, x505x}, n_n1128);
	defparam lut_5977.LUT_SIZE = 6;
	defparam lut_5977.mask = 64'h77ff77ff070707ff;

	lut_sub lut_5981 ({sk[1330], i_9_, i_7_, i_8_, i_6_, n_n536, n_n491}, n_n1117);
	defparam lut_5981.LUT_SIZE = 7;
	defparam lut_5981.mask = 128'h777f777f777f777f0111111000111000;

	lut_sub lut_5991 ({sk[1331], x22x, x521x, x21x, x13x, x544x}, n_n1285);
	defparam lut_5991.LUT_SIZE = 6;
	defparam lut_5991.mask = 64'h77ff77ff05375577;

	lut_sub lut_5995 ({sk[1332], i_9_, i_7_, i_8_, i_6_, x561x, x479x}, x22250x);
	defparam lut_5995.LUT_SIZE = 7;
	defparam lut_5995.mask = 128'h777f777f777f777fffaffcfcffffffff;

	lut_sub lut_6007 ({sk[1333], x492x, x21x, x18x, x577x}, x111x);
	defparam lut_6007.LUT_SIZE = 5;
	defparam lut_6007.mask = 32'h0fff0537;

	lut_sub lut_6010 ({sk[1334], x570x, x18x, x20x, x23x, x577x}, x458x);
	defparam lut_6010.LUT_SIZE = 6;
	defparam lut_6010.mask = 64'h77ff77ff151515ff;

	lut_sub lut_6014 ({sk[1335], i_9_, i_7_, i_8_, i_6_, n_n491, n_n195}, n_n1066);
	defparam lut_6014.LUT_SIZE = 7;
	defparam lut_6014.mask = 128'h777f777f777f777f1111100011101000;

	lut_sub lut_6024 ({sk[1336], i_9_, i_7_, i_8_, i_6_, n_n325, n_n500}, n_n1088);
	defparam lut_6024.LUT_SIZE = 7;
	defparam lut_6024.mask = 128'h777f777f777f777f0100011101011101;

	lut_sub lut_6034 ({sk[1337], x22x, x521x, x14x, x595x}, x39x);
	defparam lut_6034.LUT_SIZE = 5;
	defparam lut_6034.mask = 32'h0fff0357;

	lut_sub lut_6037 ({sk[1338], x22x, x521x, x539x, x14x, x595x}, x457x);
	defparam lut_6037.LUT_SIZE = 6;
	defparam lut_6037.mask = 64'h77ff77ff03335777;

	lut_sub lut_6041 ({sk[1339], x11x, x483x, x14x, x477x, x475x}, x11845x);
	defparam lut_6041.LUT_SIZE = 6;
	defparam lut_6041.mask = 64'h77ff77ff070707ff;

	lut_sub lut_6045 ({sk[1340], i_9_, i_7_, i_8_, i_6_, n_n509, n_n325}, x11848x);
	defparam lut_6045.LUT_SIZE = 7;
	defparam lut_6045.mask = 128'h777f777f777f777f1001000000000101;

	lut_sub lut_6050 ({sk[1341], x539x, x14x, x39x, x11845x, x11848x}, x11851x);
	defparam lut_6050.LUT_SIZE = 6;
	defparam lut_6050.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_6055 ({sk[1342], i_9_, i_7_, i_8_, i_6_, n_n509, n_n325}, x11847x);
	defparam lut_6055.LUT_SIZE = 7;
	defparam lut_6055.mask = 128'h777f777f777f777f0010101000001000;

	lut_sub lut_6060 ({sk[1343], x101x, n_n1088, x73x, x11847x}, x11852x);
	defparam lut_6060.LUT_SIZE = 5;
	defparam lut_6060.mask = 32'h0fff7fff;

	lut_sub lut_6065 ({sk[1344], i_9_, x492x, n_n491, n_n130, x20x}, x287x);
	defparam lut_6065.LUT_SIZE = 6;
	defparam lut_6065.mask = 64'h77ff77ff01010133;

	lut_sub lut_6068 ({sk[1345], i_9_, n_n522, n_n491, x519x, x586x, n_n130}, x11899x);
	defparam lut_6068.LUT_SIZE = 7;
	defparam lut_6068.mask = 128'h777f777f777f777f0000005515151555;

	lut_sub lut_6073 ({sk[1346], x21x, x12x, x591x, x520x}, x107x);
	defparam lut_6073.LUT_SIZE = 5;
	defparam lut_6073.mask = 32'h0fff0537;

	lut_sub lut_6076 ({sk[1347], i_9_, x22x, n_n473, n_n130, x503x}, x113x);
	defparam lut_6076.LUT_SIZE = 6;
	defparam lut_6076.mask = 64'h77ff77ff00031113;

	lut_sub lut_6079 ({sk[1348], x12x, x23x, x591x, x580x}, x44x);
	defparam lut_6079.LUT_SIZE = 5;
	defparam lut_6079.mask = 32'h0fff0357;

	lut_sub lut_6082 ({sk[1349], i_9_, i_7_, i_8_, i_6_, x591x, x514x}, x11905x);
	defparam lut_6082.LUT_SIZE = 7;
	defparam lut_6082.mask = 128'h777f777f777f777f0035033000000000;

	lut_sub lut_6087 ({sk[1350], x12x, x23x, x578x, x537x}, x11897x);
	defparam lut_6087.LUT_SIZE = 5;
	defparam lut_6087.mask = 32'h0fff0357;

	lut_sub lut_6090 ({sk[1351], x11x, x12x, x557x, x587x, x578x}, x11898x);
	defparam lut_6090.LUT_SIZE = 6;
	defparam lut_6090.mask = 64'h77ff77ff003f557f;

	lut_sub lut_6094 ({sk[1352], i_9_, n_n482, n_n130, n_n530, x107x}, x11903x);
	defparam lut_6094.LUT_SIZE = 6;
	defparam lut_6094.mask = 64'h77ff77ff55575557;

	lut_sub lut_6098 ({sk[1353], i_9_, n_n482, n_n528, n_n130, x113x}, x11904x);
	defparam lut_6098.LUT_SIZE = 6;
	defparam lut_6098.mask = 64'h77ff77ff55575557;

	lut_sub lut_6102 ({sk[1354], x22x, x14x, x565x, x491x}, x258x);
	defparam lut_6102.LUT_SIZE = 5;
	defparam lut_6102.mask = 32'h0fff0537;

	lut_sub lut_6105 ({sk[1355], i_9_, i_7_, i_8_, i_6_, x588x, x575x}, x12612x);
	defparam lut_6105.LUT_SIZE = 7;
	defparam lut_6105.mask = 128'h777f777f777f777f0000353000000000;

	lut_sub lut_6109 ({sk[1356], x510x, x14x, x572x, x165x, x258x, x12612x}, n_n555);
	defparam lut_6109.LUT_SIZE = 7;
	defparam lut_6109.mask = 128'h777f777f777f777f7f7f7fff7f7fffff;

	lut_sub lut_6115 ({sk[1357], i_9_, i_7_, i_8_, i_6_, x541x}, n_n4501);
	defparam lut_6115.LUT_SIZE = 6;
	defparam lut_6115.mask = 64'h77ff77ff04000000;

	lut_sub lut_6117 ({sk[1358], x22x, x521x, x539x, x17x, x596x}, n_n834);
	defparam lut_6117.LUT_SIZE = 6;
	defparam lut_6117.mask = 64'h77ff77ff03335777;

	lut_sub lut_6121 ({sk[1359], i_9_, n_n524, n_n482, n_n534, n_n491, n_n130}, x13287x);
	defparam lut_6121.LUT_SIZE = 7;
	defparam lut_6121.mask = 128'h777f777f777f777f0005111500051115;

	lut_sub lut_6126 ({sk[1360], i_9_, i_7_, i_8_, i_6_, n_n491, n_n130}, x13288x);
	defparam lut_6126.LUT_SIZE = 7;
	defparam lut_6126.mask = 128'h777f777f777f777f1110001000000010;

	lut_sub lut_6132 ({sk[1361], i_9_, x11x, n_n473, n_n130, x580x, x113x}, x13292x);
	defparam lut_6132.LUT_SIZE = 7;
	defparam lut_6132.mask = 128'h777f777f777f777f5555555f5757575f;

	lut_sub lut_6136 ({sk[1362], i_9_, i_7_, i_8_, i_6_, n_n473, n_n130}, x13293x);
	defparam lut_6136.LUT_SIZE = 7;
	defparam lut_6136.mask = 128'h777f777f777f777f0001000001010101;

	lut_sub lut_6142 ({sk[1363], i_9_, i_7_, i_8_, i_6_, n_n482, n_n130}, n_n4037);
	defparam lut_6142.LUT_SIZE = 7;
	defparam lut_6142.mask = 128'h777f777f777f777f0111001001110110;

	lut_sub lut_6152 ({sk[1364], i_9_, x21x, n_n473, n_n522, n_n130, x527x}, x13301x);
	defparam lut_6152.LUT_SIZE = 7;
	defparam lut_6152.mask = 128'h777f777f777f777f0003003311131133;

	lut_sub lut_6157 ({sk[1365], i_9_, i_7_, i_8_, i_6_, n_n130, n_n464}, x13302x);
	defparam lut_6157.LUT_SIZE = 7;
	defparam lut_6157.mask = 128'h777f777f777f777f0100010001000011;

	lut_sub lut_6163 ({sk[1366], x13292x, x13293x, n_n4037, x13301x, x13302x}, n_n4000);
	defparam lut_6163.LUT_SIZE = 6;
	defparam lut_6163.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_6169 ({sk[1367], x12x, x23x, x581x, x598x}, x11914x);
	defparam lut_6169.LUT_SIZE = 5;
	defparam lut_6169.mask = 32'h0fff0537;

	lut_sub lut_6172 ({sk[1368], x24x, x12x, x481x, x486x, x480x}, x11915x);
	defparam lut_6172.LUT_SIZE = 6;
	defparam lut_6172.mask = 64'h77ff77ff005f337f;

	lut_sub lut_6176 ({sk[1369], i_9_, i_7_, i_8_, i_6_, n_n518, n_n130}, x13313x);
	defparam lut_6176.LUT_SIZE = 7;
	defparam lut_6176.mask = 128'h777f777f777f777f0001001100000001;

	lut_sub lut_6181 ({sk[1370], i_9_, n_n518, n_n532, n_n130, x554x, n_n530}, x13314x);
	defparam lut_6181.LUT_SIZE = 7;
	defparam lut_6181.mask = 128'h777f777f777f777f1111111f0000050f;

	lut_sub lut_6186 ({sk[1371], n_n5113, n_n4144, x11914x, x11915x, x13313x, x13314x}, x13318x);
	defparam lut_6186.LUT_SIZE = 7;
	defparam lut_6186.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_6193 ({sk[1372], i_9_, i_7_, i_8_, i_6_, n_n535, n_n130}, x144x);
	defparam lut_6193.LUT_SIZE = 7;
	defparam lut_6193.mask = 128'h777f777f777f777f0010101000101010;

	lut_sub lut_6200 ({sk[1373], i_9_, x521x, n_n528, n_n535, n_n130, x23x}, x13315x);
	defparam lut_6200.LUT_SIZE = 7;
	defparam lut_6200.mask = 128'h777f777f777f777f0103010301033333;

	lut_sub lut_6205 ({sk[1374], x12x, x556x, x13322x, x22275x}, x13324x);
	defparam lut_6205.LUT_SIZE = 5;
	defparam lut_6205.mask = 32'h0fffbbbf;

	lut_sub lut_6209 ({sk[1375], x13287x, x13288x, x407x, x13282x, x22184x}, x13325x);
	defparam lut_6209.LUT_SIZE = 6;
	defparam lut_6209.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_6215 ({sk[1376], i_9_, i_7_, i_8_, i_6_, n_n491, n_n65}, n_n4028);
	defparam lut_6215.LUT_SIZE = 7;
	defparam lut_6215.mask = 128'h777f777f777f777f0101111000011110;

	lut_sub lut_6225 ({sk[1377], i_9_, i_7_, i_8_, i_6_, n_n500, n_n65}, x205x);
	defparam lut_6225.LUT_SIZE = 7;
	defparam lut_6225.mask = 128'h777f777f777f777f0000001000000010;

	lut_sub lut_6228 ({sk[1378], i_9_, i_7_, i_8_, i_6_, n_n500, n_n65}, x13347x);
	defparam lut_6228.LUT_SIZE = 7;
	defparam lut_6228.mask = 128'h777f777f777f777f1010000010101000;

	lut_sub lut_6234 ({sk[1379], i_9_, n_n534, n_n491, n_n65, x205x, x13347x}, x13348x);
	defparam lut_6234.LUT_SIZE = 7;
	defparam lut_6234.mask = 128'h777f777f777f777f7777777f7777777f;

	lut_sub lut_6239 ({sk[1380], x19x, x21x, x20x, x478x, x563x, x487x}, x13338x);
	defparam lut_6239.LUT_SIZE = 7;
	defparam lut_6239.mask = 128'h777f777f777f777f005555553f7f7f7f;

	lut_sub lut_6244 ({sk[1381], i_9_, i_7_, i_8_, i_6_, n_n509, n_n65}, x13342x);
	defparam lut_6244.LUT_SIZE = 7;
	defparam lut_6244.mask = 128'h777f777f777f777f0100010001010000;

	lut_sub lut_6249 ({sk[1382], x15x, x19x, x472x, x569x}, x13336x);
	defparam lut_6249.LUT_SIZE = 5;
	defparam lut_6249.mask = 32'h0fff0357;

	lut_sub lut_6252 ({sk[1383], x19x, x24x, x564x, x556x, x569x}, x13337x);
	defparam lut_6252.LUT_SIZE = 6;
	defparam lut_6252.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_6256 ({sk[1384], i_9_, i_7_, i_8_, i_6_, x599x, x487x}, x13340x);
	defparam lut_6256.LUT_SIZE = 7;
	defparam lut_6256.mask = 128'h777f777f777f777f3005000000000000;

	lut_sub lut_6259 ({sk[1385], x25x, x19x, x22x, x481x, x487x}, x13341x);
	defparam lut_6259.LUT_SIZE = 6;
	defparam lut_6259.mask = 64'h77ff77ff05375577;

	lut_sub lut_6263 ({sk[1386], x13338x, x13342x, x13336x, x13337x, x13340x, x13341x}, x13349x);
	defparam lut_6263.LUT_SIZE = 7;
	defparam lut_6263.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_6270 ({sk[1387], x25x, x19x, x594x, x599x, x593x}, n_n1530);
	defparam lut_6270.LUT_SIZE = 6;
	defparam lut_6270.mask = 64'h77ff77ff005f337f;

	lut_sub lut_6274 ({sk[1388], x19x, x11x, x545x, x517x, x555x}, n_n2290);
	defparam lut_6274.LUT_SIZE = 6;
	defparam lut_6274.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_6278 ({sk[1389], x19x, x21x, x490x, x20x, x533x}, x22319x);
	defparam lut_6278.LUT_SIZE = 6;
	defparam lut_6278.mask = 64'h77ff77ffeeaae0a0;

	lut_sub lut_6283 ({sk[1390], x24x, x555x, n_n1530, n_n2290, x22319x}, x13364x);
	defparam lut_6283.LUT_SIZE = 6;
	defparam lut_6283.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_6288 ({sk[1391], x19x, x550x, x23x, x533x}, x450x);
	defparam lut_6288.LUT_SIZE = 5;
	defparam lut_6288.mask = 32'h0fff111f;

	lut_sub lut_6291 ({sk[1392], i_9_, i_7_, i_8_, i_6_, n_n518, n_n65}, n_n4032);
	defparam lut_6291.LUT_SIZE = 7;
	defparam lut_6291.mask = 128'h777f777f777f777f0111101011010010;

	lut_sub lut_6301 ({sk[1393], i_9_, i_7_, i_8_, i_6_, n_n535, n_n65}, x13359x);
	defparam lut_6301.LUT_SIZE = 7;
	defparam lut_6301.mask = 128'h777f777f777f777f1010000100000100;

	lut_sub lut_6306 ({sk[1394], x22x, n_n5204, x533x, x450x, n_n4032, x13359x}, x13365x);
	defparam lut_6306.LUT_SIZE = 7;
	defparam lut_6306.mask = 128'h777f777f777f777f7f7fffff7fffffff;

	lut_sub lut_6312 ({sk[1395], x23x, x579x, x22183x, x22322x}, x13372x);
	defparam lut_6312.LUT_SIZE = 5;
	defparam lut_6312.mask = 32'h0fffeeef;

	lut_sub lut_6316 ({sk[1396], n_n1128, n_n4028, x63x, x22182x}, x13373x);
	defparam lut_6316.LUT_SIZE = 5;
	defparam lut_6316.mask = 32'h0fffbfff;

	lut_sub lut_6321 ({sk[1397], i_9_, i_7_, i_8_, i_6_, n_n195, n_n500}, n_n4050);
	defparam lut_6321.LUT_SIZE = 7;
	defparam lut_6321.mask = 128'h777f777f777f777f0110010001111110;

	lut_sub lut_6331 ({sk[1398], x15x, x11x, x18x, x524x, x532x}, n_n1952);
	defparam lut_6331.LUT_SIZE = 6;
	defparam lut_6331.mask = 64'h77ff77ff03575757;

	lut_sub lut_6335 ({sk[1399], i_9_, n_n534, n_n195, x23x, x513x, n_n464}, n_n789);
	defparam lut_6335.LUT_SIZE = 7;
	defparam lut_6335.mask = 128'h777f777f777f777f0303035703030357;

	lut_sub lut_6339 ({sk[1400], x21x, x11x, x513x, n_n4152, n_n1952, n_n789}, x13397x);
	defparam lut_6339.LUT_SIZE = 7;
	defparam lut_6339.mask = 128'h777f777f777f777f7f7f7fff7fff7fff;

	lut_sub lut_6345 ({sk[1401], x21x, x18x, x525x, x532x}, x13387x);
	defparam lut_6345.LUT_SIZE = 5;
	defparam lut_6345.mask = 32'h0fff0357;

	lut_sub lut_6348 ({sk[1402], i_9_, i_1_, i_2_, i_0_, x550x, x209x}, x13388x);
	defparam lut_6348.LUT_SIZE = 7;
	defparam lut_6348.mask = 128'h777f777f777f777f5555555555755555;

	lut_sub lut_6351 ({sk[1403], x25x, x12x, x554x, x549x}, x404x);
	defparam lut_6351.LUT_SIZE = 5;
	defparam lut_6351.mask = 32'h0fff0537;

	lut_sub lut_6354 ({sk[1404], x12x, x23x, x548x, x532x}, x13389x);
	defparam lut_6354.LUT_SIZE = 5;
	defparam lut_6354.mask = 32'h0fff0537;

	lut_sub lut_6357 ({sk[1405], x22x, x24x, x18x, x502x, x513x, x532x}, x13392x);
	defparam lut_6357.LUT_SIZE = 7;
	defparam lut_6357.mask = 128'h777f777f777f777f000f555f333f777f;

	lut_sub lut_6361 ({sk[1406], x18x, x20x, x506x, x513x, x527x, x528x}, x13393x);
	defparam lut_6361.LUT_SIZE = 7;
	defparam lut_6361.mask = 128'h777f777f777f777f00000f0f77ff7fff;

	lut_sub lut_6366 ({sk[1407], x13387x, x13388x, x404x, x13389x, x13392x, x13393x}, x13398x);
	defparam lut_6366.LUT_SIZE = 7;
	defparam lut_6366.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_6373 ({sk[1408], i_9_, i_7_, i_8_, i_6_, n_n491, n_n195}, x13413x);
	defparam lut_6373.LUT_SIZE = 7;
	defparam lut_6373.mask = 128'h777f777f777f777f0100101001001010;

	lut_sub lut_6380 ({sk[1409], x24x, x18x, x577x, x573x, x560x, x13413x}, x13414x);
	defparam lut_6380.LUT_SIZE = 7;
	defparam lut_6380.mask = 128'h777f777f777f777f55557f7f55ff7fff;

	lut_sub lut_6385 ({sk[1410], i_9_, i_7_, i_8_, i_6_, n_n473, n_n195}, x13404x);
	defparam lut_6385.LUT_SIZE = 7;
	defparam lut_6385.mask = 128'h777f777f777f777f0000000101000101;

	lut_sub lut_6390 ({sk[1411], i_9_, i_7_, i_8_, i_6_, n_n482, n_n195}, x13409x);
	defparam lut_6390.LUT_SIZE = 7;
	defparam lut_6390.mask = 128'h777f777f777f777f0000001001000110;

	lut_sub lut_6395 ({sk[1412], i_9_, i_7_, i_8_, i_6_, x590x, x513x}, x13402x);
	defparam lut_6395.LUT_SIZE = 7;
	defparam lut_6395.mask = 128'h777f777f777f777f0030050000000000;

	lut_sub lut_6398 ({sk[1413], x15x, x18x, x508x, x513x, x493x}, x13403x);
	defparam lut_6398.LUT_SIZE = 6;
	defparam lut_6398.mask = 64'h77ff77ff005f337f;

	lut_sub lut_6402 ({sk[1414], x21x, x18x, x590x, x520x}, x13408x);
	defparam lut_6402.LUT_SIZE = 5;
	defparam lut_6402.mask = 32'h0fff0537;

	lut_sub lut_6405 ({sk[1415], x458x, x13404x, x13409x, x13402x, x13403x, x13408x}, x13415x);
	defparam lut_6405.LUT_SIZE = 7;
	defparam lut_6405.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_6412 ({sk[1416], i_9_, i_7_, i_8_, i_6_, n_n518, n_n195}, x13419x);
	defparam lut_6412.LUT_SIZE = 7;
	defparam lut_6412.mask = 128'h777f777f777f777f0010100010001000;

	lut_sub lut_6417 ({sk[1417], i_9_, n_n534, n_n509, n_n195, n_n530, x494x}, x13420x);
	defparam lut_6417.LUT_SIZE = 7;
	defparam lut_6417.mask = 128'h777f777f777f777f0003000f0507050f;

	lut_sub lut_6423 ({sk[1418], x18x, x477x, x485x, x478x, x23x, x103x}, x22192x);
	defparam lut_6423.LUT_SIZE = 7;
	defparam lut_6423.mask = 128'h777f777f777f777faa88aa88a0800000;

	lut_sub lut_6428 ({sk[1419], x13380x, n_n4050, x13419x, x13420x, x22192x}, x13423x);
	defparam lut_6428.LUT_SIZE = 6;
	defparam lut_6428.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_6434 ({sk[1420], i_9_, n_n482, x510x, n_n195, x23x}, x371x);
	defparam lut_6434.LUT_SIZE = 6;
	defparam lut_6434.mask = 64'h77ff77ff00110313;

	lut_sub lut_6437 ({sk[1421], x509x, x18x, x505x, x371x}, x14659x);
	defparam lut_6437.LUT_SIZE = 5;
	defparam lut_6437.mask = 32'h0fff575f;

	lut_sub lut_6441 ({sk[1422], x492x, x21x, x18x, x23x, x577x}, x14661x);
	defparam lut_6441.LUT_SIZE = 6;
	defparam lut_6441.mask = 64'h77ff77ff11551f5f;

	lut_sub lut_6445 ({sk[1423], x25x, x18x, x590x, x587x}, x253x);
	defparam lut_6445.LUT_SIZE = 5;
	defparam lut_6445.mask = 32'h0fff0537;

	lut_sub lut_6448 ({sk[1424], i_9_, i_7_, i_8_, i_6_, x590x, x513x}, x14657x);
	defparam lut_6448.LUT_SIZE = 7;
	defparam lut_6448.mask = 128'h777f777f777f777f0035000000000000;

	lut_sub lut_6451 ({sk[1425], x11x, x24x, x18x, x503x, x513x}, x14658x);
	defparam lut_6451.LUT_SIZE = 6;
	defparam lut_6451.mask = 64'h77ff77ff03575757;

	lut_sub lut_6455 ({sk[1426], i_9_, i_5_, i_3_, i_4_, n_n534, n_n130}, x168x);
	defparam lut_6455.LUT_SIZE = 7;
	defparam lut_6455.mask = 128'h777f777f777f777f0100000001000000;

	lut_sub lut_6458 ({sk[1427], x15x, x12x, x472x, x486x, x537x, n_n5135}, x22150x);
	defparam lut_6458.LUT_SIZE = 7;
	defparam lut_6458.mask = 128'h777f777f777f777faaaa8800a0a08000;

	lut_sub lut_6463 ({sk[1428], x24x, x510x, x12x, x555x}, x14230x);
	defparam lut_6463.LUT_SIZE = 5;
	defparam lut_6463.mask = 32'h0fff0357;

	lut_sub lut_6466 ({sk[1429], i_9_, n_n482, n_n528, n_n130, x20x, x533x}, x14231x);
	defparam lut_6466.LUT_SIZE = 7;
	defparam lut_6466.mask = 128'h777f777f777f777f1111111f1111111f;

	lut_sub lut_6470 ({sk[1430], x15x, x12x, x23x, x493x, x533x}, x22273x);
	defparam lut_6470.LUT_SIZE = 6;
	defparam lut_6470.mask = 64'h77ff77fffac8aa88;

	lut_sub lut_6475 ({sk[1431], i_9_, i_7_, i_8_, i_6_, x532x}, x159x);
	defparam lut_6475.LUT_SIZE = 6;
	defparam lut_6475.mask = 64'h77ff77ff10100000;

	lut_sub lut_6478 ({sk[1432], i_9_, i_1_, i_2_, i_0_, x593x}, n_n5226);
	defparam lut_6478.LUT_SIZE = 6;
	defparam lut_6478.mask = 64'h77ff77ff00004000;

	lut_sub lut_6480 ({sk[1433], x22x, x521x, x539x, x12x, x598x}, n_n3412);
	defparam lut_6480.LUT_SIZE = 6;
	defparam lut_6480.mask = 64'h77ff77ff03335777;

	lut_sub lut_6484 ({sk[1434], i_9_, i_7_, i_8_, i_6_, n_n482, n_n325}, n_n3333);
	defparam lut_6484.LUT_SIZE = 7;
	defparam lut_6484.mask = 128'h777f777f777f777f1110101011100010;

	lut_sub lut_6494 ({sk[1435], i_9_, i_7_, i_8_, i_6_, n_n491, n_n195}, x13996x);
	defparam lut_6494.LUT_SIZE = 7;
	defparam lut_6494.mask = 128'h777f777f777f777f0101000001000011;

	lut_sub lut_6500 ({sk[1436], x15x, x22x, x12x, x568x, x536x}, n_n3771);
	defparam lut_6500.LUT_SIZE = 6;
	defparam lut_6500.mask = 64'h77ff77ff05373737;

	lut_sub lut_6504 ({sk[1437], i_9_, i_7_, i_8_, i_6_, n_n482, n_n390}, n_n2987);
	defparam lut_6504.LUT_SIZE = 7;
	defparam lut_6504.mask = 128'h777f777f777f777f0101011101010110;

	lut_sub lut_6514 ({sk[1438], i_9_, i_7_, i_8_, i_6_, x582x}, x72x);
	defparam lut_6514.LUT_SIZE = 6;
	defparam lut_6514.mask = 64'h77ff77ff04400000;

	lut_sub lut_6517 ({sk[1439], i_9_, i_7_, i_8_, i_6_, n_n390, n_n473}, x192x);
	defparam lut_6517.LUT_SIZE = 7;
	defparam lut_6517.mask = 128'h777f777f777f777f1010100010101000;

	lut_sub lut_6524 ({sk[1440], x25x, x10x, x529x, x526x}, x418x);
	defparam lut_6524.LUT_SIZE = 5;
	defparam lut_6524.mask = 32'h0fff0357;

	lut_sub lut_6527 ({sk[1441], x338x, n_n2987, x72x, x193x, x418x}, x13896x);
	defparam lut_6527.LUT_SIZE = 6;
	defparam lut_6527.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_6533 ({sk[1442], i_9_, i_7_, i_8_, i_6_, x485x}, x248x);
	defparam lut_6533.LUT_SIZE = 6;
	defparam lut_6533.mask = 64'h77ff77ff04400000;

	lut_sub lut_6536 ({sk[1443], i_9_, i_7_, i_8_, i_6_, n_n509, n_n195}, x14000x);
	defparam lut_6536.LUT_SIZE = 7;
	defparam lut_6536.mask = 128'h777f777f777f777f0101001011000000;

	lut_sub lut_6542 ({sk[1444], i_9_, n_n536, n_n534, n_n509, n_n522, n_n500}, x14153x);
	defparam lut_6542.LUT_SIZE = 7;
	defparam lut_6542.mask = 128'h777f777f777f777f0000035700000357;

	lut_sub lut_6547 ({sk[1445], i_9_, i_7_, i_8_, i_6_, n_n536, n_n509}, x14154x);
	defparam lut_6547.LUT_SIZE = 7;
	defparam lut_6547.mask = 128'h777f777f777f777f0100001011001000;

	lut_sub lut_6553 ({sk[1446], x16x, x20x, x498x, x560x}, x301x);
	defparam lut_6553.LUT_SIZE = 5;
	defparam lut_6553.mask = 32'h0fff0357;

	lut_sub lut_6556 ({sk[1447], i_9_, i_7_, i_8_, i_6_, n_n536, n_n500}, x14160x);
	defparam lut_6556.LUT_SIZE = 7;
	defparam lut_6556.mask = 128'h777f777f777f777f0000110000011100;

	lut_sub lut_6562 ({sk[1448], x23x, x498x, n_n1308, x423x, x14160x}, x14163x);
	defparam lut_6562.LUT_SIZE = 6;
	defparam lut_6562.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_6567 ({sk[1449], i_9_, n_n536, n_n528, n_n491, x572x, x491x}, x14159x);
	defparam lut_6567.LUT_SIZE = 7;
	defparam lut_6567.mask = 128'h777f777f777f777f0000000f0000777f;

	lut_sub lut_6572 ({sk[1450], x16x, x536x, x14153x, x14154x, x301x, x14159x}, x14164x);
	defparam lut_6572.LUT_SIZE = 7;
	defparam lut_6572.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_6578 ({sk[1451], i_9_, i_7_, i_8_, i_6_, n_n536, n_n482}, n_n3363);
	defparam lut_6578.LUT_SIZE = 7;
	defparam lut_6578.mask = 128'h777f777f777f777f1110100011110010;

	lut_sub lut_6588 ({sk[1452], i_9_, i_7_, i_8_, i_6_, n_n536, n_n473}, n_n3362);
	defparam lut_6588.LUT_SIZE = 7;
	defparam lut_6588.mask = 128'h777f777f777f777f0101111001011001;

	lut_sub lut_6598 ({sk[1453], x16x, x500x, x24x, x586x}, x14177x);
	defparam lut_6598.LUT_SIZE = 5;
	defparam lut_6598.mask = 32'h0fff0357;

	lut_sub lut_6601 ({sk[1454], i_9_, n_n536, n_n524, n_n491, x587x, x537x}, x14178x);
	defparam lut_6601.LUT_SIZE = 7;
	defparam lut_6601.mask = 128'h777f777f777f777f0000000f0000777f;

	lut_sub lut_6606 ({sk[1455], n_n2435, n_n3363, n_n3362, x14177x, x14178x}, n_n3287);
	defparam lut_6606.LUT_SIZE = 6;
	defparam lut_6606.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_6612 ({sk[1456], i_9_, i_7_, i_8_, i_6_, n_n536, n_n535}, n_n3370);
	defparam lut_6612.LUT_SIZE = 7;
	defparam lut_6612.mask = 128'h777f777f777f777f0101111001011010;

	lut_sub lut_6622 ({sk[1457], x16x, x501x, x23x, x581x}, x156x);
	defparam lut_6622.LUT_SIZE = 5;
	defparam lut_6622.mask = 32'h0fff0357;

	lut_sub lut_6625 ({sk[1458], x25x, x501x, x20x, x473x, x14190x, x14191x}, x14193x);
	defparam lut_6625.LUT_SIZE = 7;
	defparam lut_6625.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_6630 ({sk[1459], x198x, n_n3370, n_n4279, x106x, x14182x}, x14194x);
	defparam lut_6630.LUT_SIZE = 6;
	defparam lut_6630.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_6636 ({sk[1460], x14163x, x14164x, n_n3287, x14193x, x14194x}, n_n3262);
	defparam lut_6636.LUT_SIZE = 6;
	defparam lut_6636.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_6642 ({sk[1461], i_9_, i_1_, i_2_, i_0_, x527x}, n_n4428);
	defparam lut_6642.LUT_SIZE = 6;
	defparam lut_6642.mask = 64'h77ff77ff00000001;

	lut_sub lut_6644 ({sk[1462], x25x, x16x, x499x, x574x, x573x}, n_n3176);
	defparam lut_6644.LUT_SIZE = 6;
	defparam lut_6644.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_6648 ({sk[1463], x15x, x539x, x10x, x479x, x480x}, x15487x);
	defparam lut_6648.LUT_SIZE = 6;
	defparam lut_6648.mask = 64'h77ff77ff050f373f;

	lut_sub lut_6652 ({sk[1464], i_9_, i_7_, i_6_, x479x, x583x}, x22120x);
	defparam lut_6652.LUT_SIZE = 6;
	defparam lut_6652.mask = 64'h77ff77ffffacffff;

	lut_sub lut_6658 ({sk[1465], x25x, x509x, x18x, x580x, x505x, x513x}, x15602x);
	defparam lut_6658.LUT_SIZE = 7;
	defparam lut_6658.mask = 128'h777f777f777f777f003f00ff557f55ff;

	lut_sub lut_6663 ({sk[1466], i_9_, i_1_, i_2_, i_0_, x521x}, n_n5234);
	defparam lut_6663.LUT_SIZE = 6;
	defparam lut_6663.mask = 64'h77ff77ff00004000;

	lut_sub lut_6665 ({sk[1467], i_9_, i_1_, i_2_, i_0_, x570x}, n_n5286);
	defparam lut_6665.LUT_SIZE = 6;
	defparam lut_6665.mask = 64'h77ff77ff00004000;

	lut_sub lut_6667 ({sk[1468], x22x, x17x, x519x, x537x, x576x}, n_n3810);
	defparam lut_6667.LUT_SIZE = 6;
	defparam lut_6667.mask = 64'h77ff77ff003f557f;

	lut_sub lut_6671 ({sk[1469], x15x, x12x, x563x, x568x, x556x}, n_n2304);
	defparam lut_6671.LUT_SIZE = 6;
	defparam lut_6671.mask = 64'h77ff77ff005f337f;

	lut_sub lut_6675 ({sk[1470], x19x, x20x, x23x, x564x, x487x}, n_n1139);
	defparam lut_6675.LUT_SIZE = 6;
	defparam lut_6675.mask = 64'h77ff77ff05553777;

	lut_sub lut_6679 ({sk[1471], x19x, x21x, x474x, x472x, x487x}, n_n3031);
	defparam lut_6679.LUT_SIZE = 6;
	defparam lut_6679.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_6683 ({sk[1472], x25x, x16x, x509x, x495x}, x427x);
	defparam lut_6683.LUT_SIZE = 5;
	defparam lut_6683.mask = 32'h0fff0357;

	lut_sub lut_6686 ({sk[1473], x11x, x483x, x14x, x477x, x475x}, n_n3475);
	defparam lut_6686.LUT_SIZE = 6;
	defparam lut_6686.mask = 64'h77ff77ff070707ff;

	lut_sub lut_6690 ({sk[1474], i_9_, i_7_, i_8_, i_6_, n_n491, n_n130}, x16665x);
	defparam lut_6690.LUT_SIZE = 7;
	defparam lut_6690.mask = 128'h777f777f777f777f0000110100001000;

	lut_sub lut_6695 ({sk[1475], i_9_, n_n482, n_n130, x20x, x493x, x44x}, x16669x);
	defparam lut_6695.LUT_SIZE = 7;
	defparam lut_6695.mask = 128'h777f777f777f777f5555555f5577557f;

	lut_sub lut_6699 ({sk[1476], x12x, x20x, x489x, x533x}, x220x);
	defparam lut_6699.LUT_SIZE = 5;
	defparam lut_6699.mask = 32'h0fff0537;

	lut_sub lut_6702 ({sk[1477], i_9_, i_7_, i_8_, i_6_, x555x}, x454x);
	defparam lut_6702.LUT_SIZE = 6;
	defparam lut_6702.mask = 64'h77ff77ff01100000;

	lut_sub lut_6705 ({sk[1478], i_9_, n_n526, n_n473, n_n130, x89x}, x16673x);
	defparam lut_6705.LUT_SIZE = 6;
	defparam lut_6705.mask = 64'h77ff77ff55575557;

	lut_sub lut_6709 ({sk[1479], i_9_, i_7_, i_8_, i_6_, n_n473, n_n130}, x16674x);
	defparam lut_6709.LUT_SIZE = 7;
	defparam lut_6709.mask = 128'h777f777f777f777f0100100010101000;

	lut_sub lut_6715 ({sk[1480], i_9_, i_7_, i_8_, i_6_, n_n130, n_n464}, x16678x);
	defparam lut_6715.LUT_SIZE = 7;
	defparam lut_6715.mask = 128'h777f777f777f777f0000001000011100;

	lut_sub lut_6720 ({sk[1481], x220x, x454x, x16673x, x16674x, x16678x}, x16683x);
	defparam lut_6720.LUT_SIZE = 6;
	defparam lut_6720.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_6726 ({sk[1482], i_9_, i_1_, i_2_, i_0_, x581x, x480x}, x16684x);
	defparam lut_6726.LUT_SIZE = 7;
	defparam lut_6726.mask = 128'h777f777f777f777f0000000070000000;

	lut_sub lut_6729 ({sk[1483], x25x, x15x, x19x, x481x, x487x}, x16685x);
	defparam lut_6729.LUT_SIZE = 6;
	defparam lut_6729.mask = 64'h77ff77ff03575757;

	lut_sub lut_6733 ({sk[1484], i_9_, n_n532, n_n500, n_n65, x181x}, x16691x);
	defparam lut_6733.LUT_SIZE = 6;
	defparam lut_6733.mask = 64'h77ff77ff55575557;

	lut_sub lut_6737 ({sk[1485], x19x, x21x, x539x, x20x, x599x, x555x}, x16692x);
	defparam lut_6737.LUT_SIZE = 7;
	defparam lut_6737.mask = 128'h777f777f777f777f0707575707ff57ff;

	lut_sub lut_6742 ({sk[1486], x318x, x319x, x16684x, x16685x, x16691x, x16692x}, x16697x);
	defparam lut_6742.LUT_SIZE = 7;
	defparam lut_6742.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_6749 ({sk[1487], i_9_, i_7_, i_8_, i_6_, n_n482, n_n130}, x16703x);
	defparam lut_6749.LUT_SIZE = 7;
	defparam lut_6749.mask = 128'h777f777f777f777f0001011101011101;

	lut_sub lut_6759 ({sk[1488], x16665x, x16669x, x22072x, x22334x}, x16704x);
	defparam lut_6759.LUT_SIZE = 5;
	defparam lut_6759.mask = 32'h0fffefff;

	lut_sub lut_6764 ({sk[1489], n_n1139, n_n3031, x16679x, x16680x, x16693x}, x22071x);
	defparam lut_6764.LUT_SIZE = 6;
	defparam lut_6764.mask = 64'h77ff77ff80000000;

	lut_sub lut_6766 ({sk[1490], x24x, x554x, x23x, x532x, n_n4152, x144x}, x16715x);
	defparam lut_6766.LUT_SIZE = 7;
	defparam lut_6766.mask = 128'h777f777f777f777f777f777f777fffff;

	lut_sub lut_6771 ({sk[1491], x11x, x12x, x564x, x568x, x536x, n_n5127}, x22069x);
	defparam lut_6771.LUT_SIZE = 7;
	defparam lut_6771.mask = 128'h777f777f777f777faaaa8800a0a08000;

	lut_sub lut_6776 ({sk[1492], x21x, x20x, x486x, x568x, n_n2304, x22069x}, x16730x);
	defparam lut_6776.LUT_SIZE = 7;
	defparam lut_6776.mask = 128'h777f777f777f777fbbbbbbffbfbfbfff;

	lut_sub lut_6781 ({sk[1493], i_9_, i_7_, i_8_, i_6_, n_n473, n_n195}, n_n2214);
	defparam lut_6781.LUT_SIZE = 7;
	defparam lut_6781.mask = 128'h777f777f777f777f0111101010111000;

	lut_sub lut_6791 ({sk[1494], x11x, x20x, x590x, x577x, x16740x, x22070x}, x16742x);
	defparam lut_6791.LUT_SIZE = 7;
	defparam lut_6791.mask = 128'h777f777f777f777fbbbbbfbfbbffbfff;

	lut_sub lut_6796 ({sk[1495], x18x, x529x, n_n5087, x13387x, x13388x, x404x}, x16714x);
	defparam lut_6796.LUT_SIZE = 7;
	defparam lut_6796.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_6802 ({sk[1496], x34x, x289x, x16719x, x123x, x159x, x16709x}, x22068x);
	defparam lut_6802.LUT_SIZE = 7;
	defparam lut_6802.mask = 128'h777f777f777f777f8000000000000000;

	lut_sub lut_6804 ({sk[1497], i_9_, i_7_, i_8_, i_6_, n_n491, n_n65}, x16756x);
	defparam lut_6804.LUT_SIZE = 7;
	defparam lut_6804.mask = 128'h777f777f777f777f1110001010000010;

	lut_sub lut_6811 ({sk[1498], x15x, x19x, x518x, x573x, x569x}, x22318x);
	defparam lut_6811.LUT_SIZE = 6;
	defparam lut_6811.mask = 64'h77ff77ffffc0aa80;

	lut_sub lut_6816 ({sk[1499], x24x, x579x, x16756x, x22318x}, x16758x);
	defparam lut_6816.LUT_SIZE = 5;
	defparam lut_6816.mask = 32'h0fffbbbf;

	lut_sub lut_6820 ({sk[1500], i_9_, i_7_, i_8_, i_6_, n_n482, n_n65}, n_n2196);
	defparam lut_6820.LUT_SIZE = 7;
	defparam lut_6820.mask = 128'h777f777f777f777f0101111001011010;

	lut_sub lut_6830 ({sk[1501], x19x, x20x, x560x, x569x}, x419x);
	defparam lut_6830.LUT_SIZE = 5;
	defparam lut_6830.mask = 32'h0fff0537;

	lut_sub lut_6833 ({sk[1502], x15x, x19x, x572x, x579x}, x438x);
	defparam lut_6833.LUT_SIZE = 5;
	defparam lut_6833.mask = 32'h0fff0357;

	lut_sub lut_6836 ({sk[1503], i_9_, n_n526, n_n534, n_n491, n_n500, n_n65}, x16753x);
	defparam lut_6836.LUT_SIZE = 7;
	defparam lut_6836.mask = 128'h777f777f777f777f0005111500051115;

	lut_sub lut_6841 ({sk[1504], n_n2196, x419x, x438x, x16753x}, x16759x);
	defparam lut_6841.LUT_SIZE = 5;
	defparam lut_6841.mask = 32'h0fff7fff;

	lut_sub lut_6846 ({sk[1505], i_9_, i_1_, i_2_, i_0_, x525x}, n_n5334);
	defparam lut_6846.LUT_SIZE = 6;
	defparam lut_6846.mask = 64'h77ff77ff00004000;

	lut_sub lut_6848 ({sk[1506], i_9_, i_7_, i_8_, i_6_, x534x}, n_n5333);
	defparam lut_6848.LUT_SIZE = 6;
	defparam lut_6848.mask = 64'h77ff77ff04000000;

	lut_sub lut_6850 ({sk[1507], i_9_, i_7_, i_8_, i_6_, x530x}, n_n4813);
	defparam lut_6850.LUT_SIZE = 6;
	defparam lut_6850.mask = 64'h77ff77ff01000000;

	lut_sub lut_6852 ({sk[1508], x24x, x14x, x552x, x522x}, x16808x);
	defparam lut_6852.LUT_SIZE = 5;
	defparam lut_6852.mask = 32'h0fff0537;

	lut_sub lut_6855 ({sk[1509], x11x, x17x, x530x, x546x}, x16810x);
	defparam lut_6855.LUT_SIZE = 5;
	defparam lut_6855.mask = 32'h0fff0537;

	lut_sub lut_6858 ({sk[1510], i_9_, x22x, n_n528, n_n325, x596x, n_n464}, x16811x);
	defparam lut_6858.LUT_SIZE = 7;
	defparam lut_6858.mask = 128'h777f777f777f777f0033053700050505;

	lut_sub lut_6862 ({sk[1511], i_9_, n_n526, n_n482, n_n195, x505x, x520x}, x12315x);
	defparam lut_6862.LUT_SIZE = 7;
	defparam lut_6862.mask = 128'h777f777f777f777f0000000f0707070f;

	lut_sub lut_6867 ({sk[1512], i_9_, i_7_, i_8_, i_6_, n_n482, n_n130}, n_n1442);
	defparam lut_6867.LUT_SIZE = 7;
	defparam lut_6867.mask = 128'h777f777f777f777f0101011101010011;

	lut_sub lut_6877 ({sk[1513], i_9_, i_7_, i_8_, i_6_, x511x}, n_n4807);
	defparam lut_6877.LUT_SIZE = 6;
	defparam lut_6877.mask = 64'h77ff77ff40000000;

	lut_sub lut_6879 ({sk[1514], i_9_, n_n390, x481x, x480x, x45x}, x11562x);
	defparam lut_6879.LUT_SIZE = 6;
	defparam lut_6879.mask = 64'h77ff77ff5555557f;

	lut_sub lut_6883 ({sk[1515], i_7_, i_8_, i_6_, x10x, n_n509, x494x}, x11563x);
	defparam lut_6883.LUT_SIZE = 7;
	defparam lut_6883.mask = 128'h777f777f777f777f0507050507050707;

	lut_sub lut_6889 ({sk[1516], x21x, x14x, x488x, x511x}, x71x);
	defparam lut_6889.LUT_SIZE = 5;
	defparam lut_6889.mask = 32'h0fff0357;

	lut_sub lut_6892 ({sk[1517], x25x, x14x, x530x, x528x}, x439x);
	defparam lut_6892.LUT_SIZE = 5;
	defparam lut_6892.mask = 32'h0fff0537;

	lut_sub lut_6895 ({sk[1518], i_9_, i_1_, i_2_, i_0_, x574x, x560x}, x370x);
	defparam lut_6895.LUT_SIZE = 7;
	defparam lut_6895.mask = 128'h777f777f777f777f0000000007000000;

	lut_sub lut_6898 ({sk[1519], x24x, x12x, x568x, x562x}, x155x);
	defparam lut_6898.LUT_SIZE = 5;
	defparam lut_6898.mask = 32'h0fff0537;

	lut_sub lut_6901 ({sk[1520], x24x, x12x, x472x, x478x, x568x, x562x}, x11912x);
	defparam lut_6901.LUT_SIZE = 7;
	defparam lut_6901.mask = 128'h777f777f777f777f00005fff33337fff;

	lut_sub lut_6906 ({sk[1521], i_9_, i_7_, i_8_, i_6_, n_n130, n_n500}, x11913x);
	defparam lut_6906.LUT_SIZE = 7;
	defparam lut_6906.mask = 128'h777f777f777f777f0101000001000011;

	lut_sub lut_6912 ({sk[1522], i_9_, i_7_, i_8_, i_6_, n_n509, n_n130}, x11918x);
	defparam lut_6912.LUT_SIZE = 7;
	defparam lut_6912.mask = 128'h777f777f777f777f0001001000000011;

	lut_sub lut_6917 ({sk[1523], i_9_, i_7_, i_8_, i_6_, x569x}, n_n5259);
	defparam lut_6917.LUT_SIZE = 6;
	defparam lut_6917.mask = 64'h77ff77ff00100000;

	lut_sub lut_6919 ({sk[1524], x21x, x10x, x20x, x561x, x491x}, n_n1648);
	defparam lut_6919.LUT_SIZE = 6;
	defparam lut_6919.mask = 64'h77ff77ff03573377;

	lut_sub lut_6923 ({sk[1525], x15x, x16x, x496x, x524x}, x302x);
	defparam lut_6923.LUT_SIZE = 5;
	defparam lut_6923.mask = 32'h0fff0537;

	lut_sub lut_6926 ({sk[1526], i_9_, i_7_, i_8_, i_6_, x496x, x495x}, x13433x);
	defparam lut_6926.LUT_SIZE = 7;
	defparam lut_6926.mask = 128'h777f777f777f777f5000000300000000;

	lut_sub lut_6929 ({sk[1527], x16x, x24x, x496x, x527x, x528x}, x13435x);
	defparam lut_6929.LUT_SIZE = 6;
	defparam lut_6929.mask = 64'h77ff77ff000f777f;

	lut_sub lut_6933 ({sk[1528], x16x, x529x, n_n4421, x302x, x13433x, x13435x}, x13438x);
	defparam lut_6933.LUT_SIZE = 7;
	defparam lut_6933.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_6939 ({sk[1529], i_9_, i_7_, i_8_, i_6_, n_n455, n_n535}, n_n4094);
	defparam lut_6939.LUT_SIZE = 7;
	defparam lut_6939.mask = 128'h777f777f777f777f0101011101010110;

	lut_sub lut_6949 ({sk[1530], i_9_, i_1_, i_2_, i_0_, x550x, x516x}, x13426x);
	defparam lut_6949.LUT_SIZE = 7;
	defparam lut_6949.mask = 128'h777f777f777f777f0000000000000305;

	lut_sub lut_6952 ({sk[1531], x16x, x522x, x98x, x13428x, n_n4094, x13426x}, x13439x);
	defparam lut_6952.LUT_SIZE = 7;
	defparam lut_6952.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_6958 ({sk[1532], x273x, n_n4083, x45x, x13446x, x13450x, x13451x}, n_n4016);
	defparam lut_6958.LUT_SIZE = 7;
	defparam lut_6958.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_6965 ({sk[1533], x22x, x23x, x561x, n_n4232, n_n1648, x13460x}, x13467x);
	defparam lut_6965.LUT_SIZE = 7;
	defparam lut_6965.mask = 128'h777f777f777f777f7f7f7fff7fff7fff;

	lut_sub lut_6971 ({sk[1534], x118x, x357x, x13457x, x13458x, x13463x}, x13468x);
	defparam lut_6971.LUT_SIZE = 6;
	defparam lut_6971.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_6977 ({sk[1535], x13x, x11x, x580x, x543x, n_n4243, x13478x}, x13480x);
	defparam lut_6977.LUT_SIZE = 7;
	defparam lut_6977.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_6982 ({sk[1536], x455x, n_n4239, x13474x, x13475x, x222x, x13469x}, x13481x);
	defparam lut_6982.LUT_SIZE = 7;
	defparam lut_6982.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_6989 ({sk[1537], i_9_, i_7_, i_8_, i_6_, n_n455, n_n509}, x13488x);
	defparam lut_6989.LUT_SIZE = 7;
	defparam lut_6989.mask = 128'h777f777f777f777f1010100011000000;

	lut_sub lut_6995 ({sk[1538], x13x, x537x, n_n4247, n_n4246, n_n3152, n_n4503}, x13501x);
	defparam lut_6995.LUT_SIZE = 7;
	defparam lut_6995.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_7001 ({sk[1539], x13x, x20x, x560x, x541x}, x162x);
	defparam lut_7001.LUT_SIZE = 5;
	defparam lut_7001.mask = 32'h0fff0537;

	lut_sub lut_7004 ({sk[1540], i_9_, i_7_, i_8_, i_6_, n_n455, n_n500}, n_n4090);
	defparam lut_7004.LUT_SIZE = 7;
	defparam lut_7004.mask = 128'h777f777f777f777f0101111001110010;

	lut_sub lut_7014 ({sk[1541], x13x, x572x, x189x, x308x, x162x, n_n4090}, x13502x);
	defparam lut_7014.LUT_SIZE = 7;
	defparam lut_7014.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_7020 ({sk[1542], i_9_, i_7_, i_8_, i_6_, n_n518, n_n455}, x13505x);
	defparam lut_7020.LUT_SIZE = 7;
	defparam lut_7020.mask = 128'h777f777f777f777f1100100000000010;

	lut_sub lut_7025 ({sk[1543], x15x, x16x, x557x, x499x, x572x}, x27x);
	defparam lut_7025.LUT_SIZE = 6;
	defparam lut_7025.mask = 64'h77ff77ff005f337f;

	lut_sub lut_7029 ({sk[1544], i_9_, i_7_, i_8_, i_6_, n_n536, n_n509}, n_n4102);
	defparam lut_7029.LUT_SIZE = 7;
	defparam lut_7029.mask = 128'h777f777f777f777f0111101001110010;

	lut_sub lut_7039 ({sk[1545], i_9_, i_7_, i_8_, i_6_, x498x, x473x}, x13543x);
	defparam lut_7039.LUT_SIZE = 7;
	defparam lut_7039.mask = 128'h777f777f777f777f5300003300000000;

	lut_sub lut_7044 ({sk[1546], i_9_, i_7_, i_8_, i_6_, n_n536, n_n500}, x13544x);
	defparam lut_7044.LUT_SIZE = 7;
	defparam lut_7044.mask = 128'h777f777f777f777f0001000001011001;

	lut_sub lut_7050 ({sk[1547], x16x, x23x, x491x, x498x, x423x, x301x}, x22295x);
	defparam lut_7050.LUT_SIZE = 7;
	defparam lut_7050.mask = 128'h777f777f777f777f8888808088008000;

	lut_sub lut_7055 ({sk[1548], x27x, n_n4102, x13543x, x13544x, x22295x}, x13547x);
	defparam lut_7055.LUT_SIZE = 6;
	defparam lut_7055.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_7061 ({sk[1549], x25x, x16x, x501x, x594x, x593x}, n_n4279);
	defparam lut_7061.LUT_SIZE = 6;
	defparam lut_7061.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_7065 ({sk[1550], x283x, x13509x, x363x, x443x, x22191x}, x13520x);
	defparam lut_7065.LUT_SIZE = 6;
	defparam lut_7065.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_7071 ({sk[1551], n_n4097, x13532x, x13539x, x13530x, x13531x}, n_n4021);
	defparam lut_7071.LUT_SIZE = 6;
	defparam lut_7071.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_7077 ({sk[1552], x25x, x16x, x539x, x497x, x535x, x548x}, x13516x);
	defparam lut_7077.LUT_SIZE = 7;
	defparam lut_7077.mask = 128'h777f777f777f777f000077ff0f0f7fff;

	lut_sub lut_7082 ({sk[1553], x15x, x13x, x544x, x585x, x559x}, x55x);
	defparam lut_7082.LUT_SIZE = 6;
	defparam lut_7082.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_7086 ({sk[1554], n_n3520, x55x, x13549x}, x13551x);
	defparam lut_7086.LUT_SIZE = 4;
	defparam lut_7086.mask = 16'h5f7f;

	lut_sub lut_7090 ({sk[1555], n_n4254, x199x, x13488x, x13505x, x22190x}, x13552x);
	defparam lut_7090.LUT_SIZE = 6;
	defparam lut_7090.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_7096 ({sk[1556], i_9_, i_7_, i_8_, i_6_, n_n390, n_n500}, x14394x);
	defparam lut_7096.LUT_SIZE = 7;
	defparam lut_7096.mask = 128'h777f777f777f777f0001001001010010;

	lut_sub lut_7102 ({sk[1557], i_9_, n_n482, x11x, n_n390, n_n532, x558x}, x14397x);
	defparam lut_7102.LUT_SIZE = 7;
	defparam lut_7102.mask = 128'h777f777f777f777f0000030f0505070f;

	lut_sub lut_7107 ({sk[1558], x10x, x23x, x561x, x573x}, x119x);
	defparam lut_7107.LUT_SIZE = 5;
	defparam lut_7107.mask = 32'h0fff0357;

	lut_sub lut_7110 ({sk[1559], i_9_, i_7_, i_8_, i_6_, x571x}, x14401x);
	defparam lut_7110.LUT_SIZE = 6;
	defparam lut_7110.mask = 64'h77ff77ff00500000;

	lut_sub lut_7113 ({sk[1560], i_9_, i_7_, i_8_, i_6_, n_n390, n_n491}, x14403x);
	defparam lut_7113.LUT_SIZE = 7;
	defparam lut_7113.mask = 128'h777f777f777f777f0100001000100010;

	lut_sub lut_7118 ({sk[1561], x10x, x519x, x119x, x14401x, x14403x}, x14405x);
	defparam lut_7118.LUT_SIZE = 6;
	defparam lut_7118.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_7123 ({sk[1562], x10x, x20x, x23x, x571x, x587x}, n_n2761);
	defparam lut_7123.LUT_SIZE = 6;
	defparam lut_7123.mask = 64'h77ff77ff03335777;

	lut_sub lut_7127 ({sk[1563], i_7_, i_8_, i_6_, n_n482, x10x, x584x}, x14396x);
	defparam lut_7127.LUT_SIZE = 7;
	defparam lut_7127.mask = 128'h777f777f777f777f1111111111111311;

	lut_sub lut_7130 ({sk[1564], x10x, x23x, x479x, x563x, x560x, n_n4629}, x22159x);
	defparam lut_7130.LUT_SIZE = 7;
	defparam lut_7130.mask = 128'h777f777f777f777faaaaaa0080808000;

	lut_sub lut_7135 ({sk[1565], x14394x, x14397x, n_n2761, x14396x, x22159x}, x14406x);
	defparam lut_7135.LUT_SIZE = 6;
	defparam lut_7135.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_7141 ({sk[1566], x21x, x13x, x516x, x489x, x523x}, n_n3870);
	defparam lut_7141.LUT_SIZE = 6;
	defparam lut_7141.mask = 64'h77ff77ff003f557f;

	lut_sub lut_7145 ({sk[1567], i_9_, i_7_, i_8_, i_6_, n_n455, n_n473}, n_n3722);
	defparam lut_7145.LUT_SIZE = 7;
	defparam lut_7145.mask = 128'h777f777f777f777f0101111100011001;

	lut_sub lut_7155 ({sk[1568], x15x, x13x, x524x, x523x}, x214x);
	defparam lut_7155.LUT_SIZE = 5;
	defparam lut_7155.mask = 32'h0fff0357;

	lut_sub lut_7158 ({sk[1569], x25x, x13x, x506x, x547x, x525x, x527x}, x14416x);
	defparam lut_7158.LUT_SIZE = 7;
	defparam lut_7158.mask = 128'h777f777f777f777f000077ff0f0f7fff;

	lut_sub lut_7163 ({sk[1570], x13x, x489x, n_n3871, x455x, x14416x}, x14419x);
	defparam lut_7163.LUT_SIZE = 6;
	defparam lut_7163.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_7168 ({sk[1571], i_9_, n_n455, n_n532, x522x, x547x, x430x}, x14415x);
	defparam lut_7168.LUT_SIZE = 7;
	defparam lut_7168.mask = 128'h777f777f777f777f5577557755555f5f;

	lut_sub lut_7172 ({sk[1572], x212x, n_n3722, x214x, x14415x}, x14420x);
	defparam lut_7172.LUT_SIZE = 5;
	defparam lut_7172.mask = 32'h0fff7fff;

	lut_sub lut_7177 ({sk[1573], i_9_, i_7_, i_8_, i_6_, n_n518, n_n390}, n_n3718);
	defparam lut_7177.LUT_SIZE = 7;
	defparam lut_7177.mask = 128'h777f777f777f777f1110001010111010;

	lut_sub lut_7187 ({sk[1574], i_9_, i_7_, i_8_, i_6_, n_n390, n_n535}, x14428x);
	defparam lut_7187.LUT_SIZE = 7;
	defparam lut_7187.mask = 128'h777f777f777f777f0100001000001010;

	lut_sub lut_7192 ({sk[1575], x10x, x24x, x583x, x593x}, x14426x);
	defparam lut_7192.LUT_SIZE = 5;
	defparam lut_7192.mask = 32'h0fff0357;

	lut_sub lut_7195 ({sk[1576], x10x, x545x, x23x, x547x, x548x}, x14427x);
	defparam lut_7195.LUT_SIZE = 6;
	defparam lut_7195.mask = 64'h77ff77ff030357ff;

	lut_sub lut_7199 ({sk[1577], i_9_, i_7_, i_8_, i_6_, n_n390, n_n509}, x14434x);
	defparam lut_7199.LUT_SIZE = 7;
	defparam lut_7199.mask = 128'h777f777f777f777f0100111011110001;

	lut_sub lut_7209 ({sk[1578], n_n3718, x14428x, x14426x, x14427x, x14434x}, x14436x);
	defparam lut_7209.LUT_SIZE = 6;
	defparam lut_7209.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_7215 ({sk[1579], x22x, x11x, x17x, x552x, x535x}, n_n3461);
	defparam lut_7215.LUT_SIZE = 6;
	defparam lut_7215.mask = 64'h77ff77ff05373737;

	lut_sub lut_7219 ({sk[1580], x25x, x17x, x596x, x594x, x546x}, x13808x);
	defparam lut_7219.LUT_SIZE = 6;
	defparam lut_7219.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_7223 ({sk[1581], i_9_, i_7_, i_8_, i_6_, n_n260, n_n535}, x13809x);
	defparam lut_7223.LUT_SIZE = 7;
	defparam lut_7223.mask = 128'h777f777f777f777f0110101000100010;

	lut_sub lut_7230 ({sk[1582], x22x, x474x, x12x, x478x, x486x}, x13923x);
	defparam lut_7230.LUT_SIZE = 6;
	defparam lut_7230.mask = 64'h77ff77ff030f575f;

	lut_sub lut_7234 ({sk[1583], x12x, x472x, x23x, x564x, x486x}, x22276x);
	defparam lut_7234.LUT_SIZE = 6;
	defparam lut_7234.mask = 64'h77ff77fffafac800;

	lut_sub lut_7239 ({sk[1584], x20x, x486x, x155x, x13923x, x22276x}, n_n3307);
	defparam lut_7239.LUT_SIZE = 6;
	defparam lut_7239.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_7244 ({sk[1585], x14x, x572x, n_n4759, n_n2130, n_n4204, n_n3469}, x13796x);
	defparam lut_7244.LUT_SIZE = 7;
	defparam lut_7244.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_7250 ({sk[1586], i_9_, n_n526, n_n325, n_n491, x574x, x560x}, x13792x);
	defparam lut_7250.LUT_SIZE = 7;
	defparam lut_7250.mask = 128'h777f777f777f777f0000000f0077007f;

	lut_sub lut_7255 ({sk[1587], x15x, x69x, x575x, n_n3333, x13792x}, x13797x);
	defparam lut_7255.LUT_SIZE = 6;
	defparam lut_7255.mask = 64'h77ff77ff77ff7fff;

	lut_sub lut_7260 ({sk[1588], x15x, x14x, x524x, x530x, x527x}, n_n4196);
	defparam lut_7260.LUT_SIZE = 6;
	defparam lut_7260.mask = 64'h77ff77ff005f337f;

	lut_sub lut_7264 ({sk[1589], i_9_, i_7_, i_8_, i_6_, n_n473, n_n325}, n_n3332);
	defparam lut_7264.LUT_SIZE = 7;
	defparam lut_7264.mask = 128'h777f777f777f777f0000011101011111;

	lut_sub lut_7274 ({sk[1590], i_9_, i_7_, i_8_, i_6_, n_n509, n_n260}, n_n3327);
	defparam lut_7274.LUT_SIZE = 7;
	defparam lut_7274.mask = 128'h777f777f777f777f0110111100011100;

	lut_sub lut_7284 ({sk[1591], x15x, x521x, x24x, x17x, x482x, x596x}, x13818x);
	defparam lut_7284.LUT_SIZE = 7;
	defparam lut_7284.mask = 128'h777f777f777f777f03570f5f57575f5f;

	lut_sub lut_7289 ({sk[1592], i_9_, i_7_, i_8_, i_6_, n_n518, n_n260}, x13819x);
	defparam lut_7289.LUT_SIZE = 7;
	defparam lut_7289.mask = 128'h777f777f777f777f1000000011100010;

	lut_sub lut_7295 ({sk[1593], x13808x, x13809x, n_n3327, x13818x, x13819x}, n_n3275);
	defparam lut_7295.LUT_SIZE = 6;
	defparam lut_7295.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_7301 ({sk[1594], x15x, x17x, x524x, x531x, x527x}, n_n2710);
	defparam lut_7301.LUT_SIZE = 6;
	defparam lut_7301.mask = 64'h77ff77ff005f337f;

	lut_sub lut_7305 ({sk[1595], x25x, x15x, x17x, x557x, x589x, x576x}, x13857x);
	defparam lut_7305.LUT_SIZE = 7;
	defparam lut_7305.mask = 128'h777f777f777f777f000f333f777f777f;

	lut_sub lut_7310 ({sk[1596], n_n3450, n_n3451, x13857x}, x13860x);
	defparam lut_7310.LUT_SIZE = 4;
	defparam lut_7310.mask = 16'h5f7f;

	lut_sub lut_7314 ({sk[1597], x15x, x17x, x572x, x576x}, x49x);
	defparam lut_7314.LUT_SIZE = 5;
	defparam lut_7314.mask = 32'h0fff0357;

	lut_sub lut_7317 ({sk[1598], x11x, x17x, x566x, x562x}, x13849x);
	defparam lut_7317.LUT_SIZE = 5;
	defparam lut_7317.mask = 32'h0fff0537;

	lut_sub lut_7320 ({sk[1599], x24x, x17x, x570x, x589x}, x13852x);
	defparam lut_7320.LUT_SIZE = 5;
	defparam lut_7320.mask = 32'h0fff0357;

	lut_sub lut_7323 ({sk[1600], x22x, x17x, x519x, x20x, x587x, x576x}, x13855x);
	defparam lut_7323.LUT_SIZE = 7;
	defparam lut_7323.mask = 128'h777f777f777f777f050537ff555577ff;

	lut_sub lut_7328 ({sk[1601], x461x, x13850x, x49x, x13849x, x13852x, x13855x}, x13861x);
	defparam lut_7328.LUT_SIZE = 7;
	defparam lut_7328.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_7335 ({sk[1602], i_9_, i_7_, i_8_, i_6_, n_n473, n_n260}, n_n3322);
	defparam lut_7335.LUT_SIZE = 7;
	defparam lut_7335.mask = 128'h777f777f777f777f0111101011001010;

	lut_sub lut_7345 ({sk[1603], x22x, x11x, x17x, x522x, x531x}, x58x);
	defparam lut_7345.LUT_SIZE = 6;
	defparam lut_7345.mask = 64'h77ff77ff03575757;

	lut_sub lut_7349 ({sk[1604], i_9_, i_7_, i_8_, i_6_, n_n482, n_n260}, x138x);
	defparam lut_7349.LUT_SIZE = 7;
	defparam lut_7349.mask = 128'h777f777f777f777f1110000011100000;

	lut_sub lut_7356 ({sk[1605], x25x, x17x, x531x, x528x}, x331x);
	defparam lut_7356.LUT_SIZE = 5;
	defparam lut_7356.mask = 32'h0fff0537;

	lut_sub lut_7359 ({sk[1606], x25x, x23x, x512x, n_n2710, x138x}, x13876x);
	defparam lut_7359.LUT_SIZE = 6;
	defparam lut_7359.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_7364 ({sk[1607], x25x, x531x, n_n4938, n_n3322, x58x, x13871x}, x13877x);
	defparam lut_7364.LUT_SIZE = 7;
	defparam lut_7364.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_7370 ({sk[1608], i_9_, i_7_, i_8_, i_6_, n_n325, n_n535}, x13908x);
	defparam lut_7370.LUT_SIZE = 7;
	defparam lut_7370.mask = 128'h777f777f777f777f0100101000101010;

	lut_sub lut_7377 ({sk[1609], x11x, x23x, x595x, x551x, x457x, x13908x}, x13910x);
	defparam lut_7377.LUT_SIZE = 7;
	defparam lut_7377.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_7382 ({sk[1610], i_9_, i_7_, i_8_, i_6_, n_n390, n_n464}, x13903x);
	defparam lut_7382.LUT_SIZE = 7;
	defparam lut_7382.mask = 128'h777f777f777f777f0010100011000010;

	lut_sub lut_7388 ({sk[1611], x14x, x20x, x594x, x546x, x551x, x593x}, x13906x);
	defparam lut_7388.LUT_SIZE = 7;
	defparam lut_7388.mask = 128'h777f777f777f777f000033335fff7fff;

	lut_sub lut_7393 ({sk[1612], x10x, x14x, x516x, x241x, x585x, n_n4689}, x22175x);
	defparam lut_7393.LUT_SIZE = 7;
	defparam lut_7393.mask = 128'h777f777f777f777fa0a08080a0008000;

	lut_sub lut_7398 ({sk[1613], x442x, x13903x, x13906x, x22175x}, x13911x);
	defparam lut_7398.LUT_SIZE = 5;
	defparam lut_7398.mask = 32'h0fffbfff;

	lut_sub lut_7403 ({sk[1614], i_9_, i_7_, i_8_, i_6_, n_n509, n_n325}, x456x);
	defparam lut_7403.LUT_SIZE = 7;
	defparam lut_7403.mask = 128'h777f777f777f777f1010101010001000;

	lut_sub lut_7410 ({sk[1615], i_9_, i_7_, i_8_, i_6_, n_n509, n_n325}, x13914x);
	defparam lut_7410.LUT_SIZE = 7;
	defparam lut_7410.mask = 128'h777f777f777f777f0000010000010101;

	lut_sub lut_7415 ({sk[1616], x25x, x15x, x483x, x23x, x595x, x101x}, x22174x);
	defparam lut_7415.LUT_SIZE = 7;
	defparam lut_7415.mask = 128'h777f777f777f777fa8a8a800a800a800;

	lut_sub lut_7420 ({sk[1617], n_n3336, n_n3475, x456x, x13914x, x22174x}, x13919x);
	defparam lut_7420.LUT_SIZE = 6;
	defparam lut_7420.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_7426 ({sk[1618], x25x, x22x, x10x, x507x, x520x, x527x}, x13893x);
	defparam lut_7426.LUT_SIZE = 7;
	defparam lut_7426.mask = 128'h777f777f777f777f00770f7f0f7f0f7f;

	lut_sub lut_7431 ({sk[1619], i_9_, i_7_, i_8_, i_6_, x588x, x565x}, x13744x);
	defparam lut_7431.LUT_SIZE = 7;
	defparam lut_7431.mask = 128'h777f777f777f777f0003500000000000;

	lut_sub lut_7434 ({sk[1620], x21x, x11x, x14x, x494x, x595x, x511x}, x13746x);
	defparam lut_7434.LUT_SIZE = 7;
	defparam lut_7434.mask = 128'h777f777f777f777f000f555f333f777f;

	lut_sub lut_7438 ({sk[1621], x24x, x14x, x588x, x520x, x536x}, x22292x);
	defparam lut_7438.LUT_SIZE = 6;
	defparam lut_7438.mask = 64'h77ff77ffff88f080;

	lut_sub lut_7443 ({sk[1622], x11x, x575x, x13744x, x13746x, x22292x}, n_n3202);
	defparam lut_7443.LUT_SIZE = 6;
	defparam lut_7443.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_7448 ({sk[1623], x25x, x10x, x571x, x560x}, x357x);
	defparam lut_7448.LUT_SIZE = 5;
	defparam lut_7448.mask = 32'h0fff0537;

	lut_sub lut_7451 ({sk[1624], i_9_, x521x, n_n390, n_n532, n_n535, x517x}, x13753x);
	defparam lut_7451.LUT_SIZE = 7;
	defparam lut_7451.mask = 128'h777f777f777f777f00030003005700ff;

	lut_sub lut_7456 ({sk[1625], i_9_, i_7_, i_8_, i_6_, x561x, x547x}, x13751x);
	defparam lut_7456.LUT_SIZE = 7;
	defparam lut_7456.mask = 128'h777f777f777f777f5030000000000000;

	lut_sub lut_7459 ({sk[1626], x24x, x571x, x357x, x13753x, x13751x}, n_n3204);
	defparam lut_7459.LUT_SIZE = 6;
	defparam lut_7459.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_7464 ({sk[1627], i_9_, i_7_, i_8_, i_6_, n_n455, n_n500}, n_n2999);
	defparam lut_7464.LUT_SIZE = 7;
	defparam lut_7464.mask = 128'h777f777f777f777f0100111001111010;

	lut_sub lut_7474 ({sk[1628], x22x, x10x, x519x, x571x, x537x}, n_n3132);
	defparam lut_7474.LUT_SIZE = 6;
	defparam lut_7474.mask = 64'h77ff77ff005f337f;

	lut_sub lut_7478 ({sk[1629], i_9_, i_7_, i_8_, i_6_, n_n482, n_n325}, x15756x);
	defparam lut_7478.LUT_SIZE = 7;
	defparam lut_7478.mask = 128'h777f777f777f777f0100010000001010;

	lut_sub lut_7483 ({sk[1630], i_9_, i_7_, i_8_, i_6_, n_n473, n_n260}, x15701x);
	defparam lut_7483.LUT_SIZE = 7;
	defparam lut_7483.mask = 128'h777f777f777f777f0010000000101110;

	lut_sub lut_7489 ({sk[1631], x16x, x20x, x23x, x506x, x495x}, n_n2803);
	defparam lut_7489.LUT_SIZE = 6;
	defparam lut_7489.mask = 64'h77ff77ff05553777;

	lut_sub lut_7493 ({sk[1632], x17x, x552x, x490x, x23x, x517x, x594x}, x14894x);
	defparam lut_7493.LUT_SIZE = 7;
	defparam lut_7493.mask = 128'h777f777f777f777f00000f0f77ff7fff;

	lut_sub lut_7498 ({sk[1633], x14x, x20x, x525x, x530x}, x389x);
	defparam lut_7498.LUT_SIZE = 5;
	defparam lut_7498.mask = 32'h0fff0537;

	lut_sub lut_7501 ({sk[1634], x25x, x24x, x552x, x23x, x530x, n_n4824}, x22146x);
	defparam lut_7501.LUT_SIZE = 7;
	defparam lut_7501.mask = 128'h777f777f777f777fa8a8a800a800a800;

	lut_sub lut_7506 ({sk[1635], i_9_, i_7_, i_8_, i_6_, x569x}, n_n5257);
	defparam lut_7506.LUT_SIZE = 6;
	defparam lut_7506.mask = 64'h77ff77ff00010000;

	lut_sub lut_7508 ({sk[1636], i_9_, i_7_, i_8_, i_6_, n_n509, n_n65}, x15175x);
	defparam lut_7508.LUT_SIZE = 7;
	defparam lut_7508.mask = 128'h777f777f777f777f0010100010101000;

	lut_sub lut_7514 ({sk[1637], x19x, x23x, x563x, x487x, x433x, x15175x}, n_n2568);
	defparam lut_7514.LUT_SIZE = 7;
	defparam lut_7514.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_7519 ({sk[1638], x19x, x24x, x480x, x487x}, x146x);
	defparam lut_7519.LUT_SIZE = 5;
	defparam lut_7519.mask = 32'h0fff0537;

	lut_sub lut_7522 ({sk[1639], i_9_, i_7_, i_8_, i_6_, x599x}, x320x);
	defparam lut_7522.LUT_SIZE = 6;
	defparam lut_7522.mask = 64'h77ff77ff44000000;

	lut_sub lut_7525 ({sk[1640], x19x, x22x, x581x, x487x}, x15176x);
	defparam lut_7525.LUT_SIZE = 5;
	defparam lut_7525.mask = 32'h0fff0537;

	lut_sub lut_7528 ({sk[1641], x19x, x481x, x318x, x146x, x320x, x15176x}, n_n2569);
	defparam lut_7528.LUT_SIZE = 7;
	defparam lut_7528.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_7534 ({sk[1642], i_9_, i_7_, i_8_, i_6_, n_n500, n_n65}, x15184x);
	defparam lut_7534.LUT_SIZE = 7;
	defparam lut_7534.mask = 128'h777f777f777f777f0010111011101010;

	lut_sub lut_7544 ({sk[1643], i_9_, i_7_, i_8_, i_6_, n_n473, n_n65}, x267x);
	defparam lut_7544.LUT_SIZE = 7;
	defparam lut_7544.mask = 128'h777f777f777f777f0010100010101000;

	lut_sub lut_7550 ({sk[1644], x19x, x21x, x516x, x503x, x534x}, x15187x);
	defparam lut_7550.LUT_SIZE = 6;
	defparam lut_7550.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_7554 ({sk[1645], i_9_, i_7_, i_8_, i_6_, n_n464, n_n65}, x15189x);
	defparam lut_7554.LUT_SIZE = 7;
	defparam lut_7554.mask = 128'h777f777f777f777f0101000001000110;

	lut_sub lut_7560 ({sk[1646], x149x, x268x, n_n3019, x267x, x15187x, x15189x}, n_n2535);
	defparam lut_7560.LUT_SIZE = 7;
	defparam lut_7560.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_7567 ({sk[1647], i_9_, n_n482, x510x, x23x, n_n65, x63x}, x15195x);
	defparam lut_7567.LUT_SIZE = 7;
	defparam lut_7567.mask = 128'h777f777f777f777f5555575755775777;

	lut_sub lut_7571 ({sk[1648], i_9_, n_n534, n_n491, n_n65, x438x}, x15198x);
	defparam lut_7571.LUT_SIZE = 6;
	defparam lut_7571.mask = 64'h77ff77ff55575557;

	lut_sub lut_7575 ({sk[1649], i_9_, i_1_, i_2_, i_0_, x570x, x587x}, x207x);
	defparam lut_7575.LUT_SIZE = 7;
	defparam lut_7575.mask = 128'h777f777f777f777f0000000070000000;

	lut_sub lut_7578 ({sk[1650], x592x, x19x, x24x, x586x, x15201x, x15202x}, x15204x);
	defparam lut_7578.LUT_SIZE = 7;
	defparam lut_7578.mask = 128'h777f777f777f777f77777f7f77ff7fff;

	lut_sub lut_7583 ({sk[1651], x15195x, x15198x, x15194x, x15197x, x22137x}, x15205x);
	defparam lut_7583.LUT_SIZE = 6;
	defparam lut_7583.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_7589 ({sk[1652], x11x, x12x, x554x, x535x}, x143x);
	defparam lut_7589.LUT_SIZE = 5;
	defparam lut_7589.mask = 32'h0fff0537;

	lut_sub lut_7592 ({sk[1653], i_9_, i_7_, i_8_, i_6_, x554x, x486x}, x14782x);
	defparam lut_7592.LUT_SIZE = 7;
	defparam lut_7592.mask = 128'h777f777f777f777f0000000700000000;

	lut_sub lut_7595 ({sk[1654], i_9_, i_5_, i_3_, i_4_, n_n532, n_n65}, x385x);
	defparam lut_7595.LUT_SIZE = 7;
	defparam lut_7595.mask = 128'h777f777f777f777f0001000000010000;

	lut_sub lut_7598 ({sk[1655], x19x, x12x, x580x, x503x, x548x, x493x}, x14790x);
	defparam lut_7598.LUT_SIZE = 7;
	defparam lut_7598.mask = 128'h777f777f777f777f00005fff33337fff;

	lut_sub lut_7603 ({sk[1656], i_9_, i_7_, i_8_, i_6_, x578x}, x125x);
	defparam lut_7603.LUT_SIZE = 6;
	defparam lut_7603.mask = 64'h77ff77ff00110000;

	lut_sub lut_7606 ({sk[1657], x18x, x20x, x489x, x532x}, x209x);
	defparam lut_7606.LUT_SIZE = 5;
	defparam lut_7606.mask = 32'h0fff0537;

	lut_sub lut_7609 ({sk[1658], x25x, x16x, x501x, x593x}, x410x);
	defparam lut_7609.LUT_SIZE = 5;
	defparam lut_7609.mask = 32'h0fff0537;

	lut_sub lut_7612 ({sk[1659], x18x, x597x, x482x, x23x}, x43x);
	defparam lut_7612.LUT_SIZE = 5;
	defparam lut_7612.mask = 32'h0fff0537;

	lut_sub lut_7615 ({sk[1660], i_9_, n_n524, n_n518, n_n195, x43x}, x12155x);
	defparam lut_7615.LUT_SIZE = 6;
	defparam lut_7615.mask = 64'h77ff77ff55575557;

	lut_sub lut_7619 ({sk[1661], x19x, x23x, x574x, x560x, x569x}, n_n1521);
	defparam lut_7619.LUT_SIZE = 6;
	defparam lut_7619.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_7623 ({sk[1662], x22x, x21x, x10x, x516x, x526x}, n_n3849);
	defparam lut_7623.LUT_SIZE = 6;
	defparam lut_7623.mask = 64'h77ff77ff03575757;

	lut_sub lut_7627 ({sk[1663], i_9_, i_7_, i_8_, i_6_, n_n390, n_n464}, x11863x);
	defparam lut_7627.LUT_SIZE = 7;
	defparam lut_7627.mask = 128'h777f777f777f777f0000111000101000;

	lut_sub lut_7633 ({sk[1664], x15x, x18x, x567x, x562x}, x299x);
	defparam lut_7633.LUT_SIZE = 5;
	defparam lut_7633.mask = 32'h0fff0537;

	lut_sub lut_7636 ({sk[1665], i_9_, i_7_, i_8_, i_6_, n_n509, n_n65}, x11921x);
	defparam lut_7636.LUT_SIZE = 7;
	defparam lut_7636.mask = 128'h777f777f777f777f0100000001101000;

	lut_sub lut_7641 ({sk[1666], i_9_, i_7_, i_8_, i_6_, n_n500, n_n65}, n_n1049);
	defparam lut_7641.LUT_SIZE = 7;
	defparam lut_7641.mask = 128'h777f777f777f777f0111010100011110;

	lut_sub lut_7651 ({sk[1667], i_9_, n_n522, n_n491, x570x, x587x, n_n65}, x11929x);
	defparam lut_7651.LUT_SIZE = 7;
	defparam lut_7651.mask = 128'h777f777f777f777f0000005515151555;

	lut_sub lut_7656 ({sk[1668], i_9_, i_7_, i_8_, i_6_, n_n491, n_n65}, x11930x);
	defparam lut_7656.LUT_SIZE = 7;
	defparam lut_7656.mask = 128'h777f777f777f777f1100101000000010;

	lut_sub lut_7662 ({sk[1669], i_9_, x24x, n_n491, x573x, n_n65, x438x}, x11933x);
	defparam lut_7662.LUT_SIZE = 7;
	defparam lut_7662.mask = 128'h777f777f777f777f5555557757575777;

	lut_sub lut_7666 ({sk[1670], i_9_, i_7_, i_8_, i_6_, n_n482, n_n65}, x11940x);
	defparam lut_7666.LUT_SIZE = 7;
	defparam lut_7666.mask = 128'h777f777f777f777f0011110001101110;

	lut_sub lut_7676 ({sk[1671], x25x, x19x, x557x, x579x}, x11932x);
	defparam lut_7676.LUT_SIZE = 5;
	defparam lut_7676.mask = 32'h0fff0357;

	lut_sub lut_7679 ({sk[1672], n_n1521, x11929x, x11930x, x11933x, x11940x, x11932x}, n_n1017);
	defparam lut_7679.LUT_SIZE = 7;
	defparam lut_7679.mask = 128'h777f777f777f777f7fffffffffffffff;

	lut_sub lut_7686 ({sk[1673], i_9_, i_7_, i_8_, i_6_, n_n473, n_n65}, x11944x);
	defparam lut_7686.LUT_SIZE = 7;
	defparam lut_7686.mask = 128'h777f777f777f777f0000001100000110;

	lut_sub lut_7691 ({sk[1674], x515x, x11x, n_n5303, n_n1128, x11944x}, n_n1045);
	defparam lut_7691.LUT_SIZE = 6;
	defparam lut_7691.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_7696 ({sk[1675], x25x, x19x, x24x, x534x, x528x}, n_n1900);
	defparam lut_7696.LUT_SIZE = 6;
	defparam lut_7696.mask = 64'h77ff77ff03573377;

	lut_sub lut_7700 ({sk[1676], i_9_, n_n524, n_n473, n_n522, n_n464, n_n65}, x11949x);
	defparam lut_7700.LUT_SIZE = 7;
	defparam lut_7700.mask = 128'h777f777f777f777f0005111500051115;

	lut_sub lut_7705 ({sk[1677], i_9_, i_7_, i_8_, i_6_, n_n464, n_n65}, x11950x);
	defparam lut_7705.LUT_SIZE = 7;
	defparam lut_7705.mask = 128'h777f777f777f777f0101000001010000;

	lut_sub lut_7710 ({sk[1678], x515x, x23x, n_n5333, n_n1900, x11949x, x11950x}, x11953x);
	defparam lut_7710.LUT_SIZE = 7;
	defparam lut_7710.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_7716 ({sk[1679], i_9_, x24x, n_n534, n_n509, x581x, n_n65}, x11958x);
	defparam lut_7716.LUT_SIZE = 7;
	defparam lut_7716.mask = 128'h777f777f777f777f0005050511151515;

	lut_sub lut_7721 ({sk[1680], i_9_, i_7_, i_8_, i_6_, n_n518, n_n65}, x11959x);
	defparam lut_7721.LUT_SIZE = 7;
	defparam lut_7721.mask = 128'h777f777f777f777f1010001001100000;

	lut_sub lut_7727 ({sk[1681], x19x, x480x, n_n5249, n_n1139, x11921x, n_n1049}, x11961x);
	defparam lut_7727.LUT_SIZE = 7;
	defparam lut_7727.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_7733 ({sk[1682], i_7_, i_8_, i_6_, x10x, n_n473, n_n464}, x12621x);
	defparam lut_7733.LUT_SIZE = 7;
	defparam lut_7733.mask = 128'h777f777f777f777f0007050300000300;

	lut_sub lut_7739 ({sk[1683], x538x, x11x, x10x, x488x, x551x}, x22264x);
	defparam lut_7739.LUT_SIZE = 6;
	defparam lut_7739.mask = 64'h77ff77fffca8f0a0;

	lut_sub lut_7744 ({sk[1684], x14x, x549x, x12621x, x22264x}, n_n557);
	defparam lut_7744.LUT_SIZE = 5;
	defparam lut_7744.mask = 32'h0fffbbbf;

	lut_sub lut_7748 ({sk[1685], i_9_, n_n532, n_n500, x556x, n_n65, x548x}, x12634x);
	defparam lut_7748.LUT_SIZE = 7;
	defparam lut_7748.mask = 128'h777f777f777f777f0000003313131333;

	lut_sub lut_7753 ({sk[1686], i_9_, i_1_, i_2_, i_0_, x518x, x494x}, x12632x);
	defparam lut_7753.LUT_SIZE = 7;
	defparam lut_7753.mask = 128'h777f777f777f777f0000000070000000;

	lut_sub lut_7756 ({sk[1687], i_9_, i_7_, i_8_, i_6_, x576x}, n_n4889);
	defparam lut_7756.LUT_SIZE = 6;
	defparam lut_7756.mask = 64'h77ff77ff00010000;

	lut_sub lut_7758 ({sk[1688], i_9_, i_7_, i_8_, i_6_, n_n464, n_n65}, x13567x);
	defparam lut_7758.LUT_SIZE = 7;
	defparam lut_7758.mask = 128'h777f777f777f777f0101001001010111;

	lut_sub lut_7767 ({sk[1689], x19x, x23x, x525x, x534x}, x13562x);
	defparam lut_7767.LUT_SIZE = 5;
	defparam lut_7767.mask = 32'h0fff0537;

	lut_sub lut_7770 ({sk[1690], x515x, x22x, x268x, x267x, x13567x, x13562x}, n_n3996);
	defparam lut_7770.LUT_SIZE = 7;
	defparam lut_7770.mask = 128'h777f777f777f777f7fff7fff7fffffff;

	lut_sub lut_7776 ({sk[1691], i_9_, x25x, n_n482, n_n390, n_n532, x587x}, x13457x);
	defparam lut_7776.LUT_SIZE = 7;
	defparam lut_7776.mask = 128'h777f777f777f777f0003000f0507050f;

	lut_sub lut_7781 ({sk[1692], i_9_, n_n524, n_n390, n_n491, x584x, n_n3132}, x13458x);
	defparam lut_7781.LUT_SIZE = 7;
	defparam lut_7781.mask = 128'h777f777f777f777f5555555f55775577;

	lut_sub lut_7785 ({sk[1693], i_9_, i_7_, i_8_, i_6_, n_n518, n_n325}, n_n3708);
	defparam lut_7785.LUT_SIZE = 7;
	defparam lut_7785.mask = 128'h777f777f777f777f0100110011111010;

	lut_sub lut_7795 ({sk[1694], i_9_, n_n532, n_n325, n_n535, x442x}, x14350x);
	defparam lut_7795.LUT_SIZE = 6;
	defparam lut_7795.mask = 64'h77ff77ff55575557;

	lut_sub lut_7799 ({sk[1695], x25x, x14x, x594x, x595x, x593x}, x14354x);
	defparam lut_7799.LUT_SIZE = 6;
	defparam lut_7799.mask = 64'h77ff77ff005f337f;

	lut_sub lut_7803 ({sk[1696], i_9_, i_7_, i_8_, i_6_, n_n325, n_n535}, x14355x);
	defparam lut_7803.LUT_SIZE = 7;
	defparam lut_7803.mask = 128'h777f777f777f777f1000001000001010;

	lut_sub lut_7808 ({sk[1697], x21x, x14x, x546x, x551x, x14354x, x14355x}, x14357x);
	defparam lut_7808.LUT_SIZE = 7;
	defparam lut_7808.mask = 128'h777f777f777f777f777777ff7f7f7fff;

	lut_sub lut_7813 ({sk[1698], x10x, x20x, x525x, x489x, x526x}, n_n3848);
	defparam lut_7813.LUT_SIZE = 6;
	defparam lut_7813.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_7817 ({sk[1699], x14x, x545x, x550x, n_n3708, x14350x, n_n3848}, x14358x);
	defparam lut_7817.LUT_SIZE = 7;
	defparam lut_7817.mask = 128'h777f777f777f777f7f7f7f7f7fffffff;

	lut_sub lut_7823 ({sk[1700], i_9_, i_7_, i_8_, i_6_, n_n390, n_n464}, n_n3711);
	defparam lut_7823.LUT_SIZE = 7;
	defparam lut_7823.mask = 128'h0fff0fff3fff3fff0001111001011110;

	lut_sub lut_7833 ({sk[1701], i_9_, i_7_, i_8_, i_6_, n_n482, n_n390}, x14370x);
	defparam lut_7833.LUT_SIZE = 7;
	defparam lut_7833.mask = 128'h0fff0fff3fff3fff1010101010000000;

	lut_sub lut_7839 ({sk[1702], i_9_, i_7_, i_8_, i_6_, n_n390, n_n473}, x22152x);
	defparam lut_7839.LUT_SIZE = 7;
	defparam lut_7839.mask = 128'h0fff0fff3fff3fffffeeeeefffffeefe;

	lut_sub lut_7847 ({sk[1703], x10x, x507x, x23x, x503x, x488x, x418x}, x22153x);
	defparam lut_7847.LUT_SIZE = 7;
	defparam lut_7847.mask = 128'h0fff0fff3fff3fffaaaaaa0080808000;

	lut_sub lut_7852 ({sk[1704], n_n3711, x14370x, x22152x, x22153x}, n_n3649);
	defparam lut_7852.LUT_SIZE = 5;
	defparam lut_7852.mask = 32'h00ffefff;

	lut_sub lut_7857 ({sk[1705], i_9_, i_7_, i_8_, i_6_, n_n455, n_n509}, n_n3727);
	defparam lut_7857.LUT_SIZE = 7;
	defparam lut_7857.mask = 128'h0fff0fff3fff3fff1100111001111000;

	lut_sub lut_7867 ({sk[1706], i_9_, i_7_, i_8_, i_6_, n_n455, n_n500}, n_n3726);
	defparam lut_7867.LUT_SIZE = 7;
	defparam lut_7867.mask = 128'h0fff0fff3fff3fff0100010101110111;

	lut_sub lut_7877 ({sk[1707], x13x, x24x, x557x, x542x, n_n4531, n_n4501}, x22165x);
	defparam lut_7877.LUT_SIZE = 7;
	defparam lut_7877.mask = 128'h0fff0fff3fff3fff8888808088008000;

	lut_sub lut_7882 ({sk[1708], x13x, x570x, x23x, x587x, x542x}, n_n3879);
	defparam lut_7882.LUT_SIZE = 6;
	defparam lut_7882.mask = 64'h00ff55ff050537ff;

	lut_sub lut_7886 ({sk[1709], i_9_, i_7_, i_8_, i_6_, x543x}, x14446x);
	defparam lut_7886.LUT_SIZE = 6;
	defparam lut_7886.mask = 64'h00ff55ff00110000;

	lut_sub lut_7889 ({sk[1710], x13x, x20x, x584x, x542x}, x14447x);
	defparam lut_7889.LUT_SIZE = 5;
	defparam lut_7889.mask = 32'h00ff0537;

	lut_sub lut_7892 ({sk[1711], i_9_, n_n526, n_n455, n_n491, x378x}, x14453x);
	defparam lut_7892.LUT_SIZE = 6;
	defparam lut_7892.mask = 64'h00ff55ff55575557;

	lut_sub lut_7896 ({sk[1712], x13x, x23x, x574x, x520x, x541x, x493x}, x14454x);
	defparam lut_7896.LUT_SIZE = 7;
	defparam lut_7896.mask = 128'h0fff0fff3fff3fff000033335fff7fff;

	lut_sub lut_7901 ({sk[1713], x16x, x472x, x478x, x14465x, x22158x}, n_n3737);
	defparam lut_7901.LUT_SIZE = 6;
	defparam lut_7901.mask = 64'h5fffffffbbbbbfff;

	lut_sub lut_7906 ({sk[1714], x16x, x574x, x300x, x14471x, x14469x}, n_n3736);
	defparam lut_7906.LUT_SIZE = 6;
	defparam lut_7906.mask = 64'h5fffffff7f7f7fff;

	lut_sub lut_7911 ({sk[1715], n_n3740, x14484x, x14485x, x14487x, x22157x}, n_n3658);
	defparam lut_7911.LUT_SIZE = 6;
	defparam lut_7911.mask = 64'h5fffffffbfffffff;

	lut_sub lut_7917 ({sk[1716], x24x, x495x, x14505x, x22297x}, x14507x);
	defparam lut_7917.LUT_SIZE = 5;
	defparam lut_7917.mask = 32'h77ffbbbf;

	lut_sub lut_7921 ({sk[1717], x15x, x500x, n_n4391, n_n1693, n_n3732, x14498x}, x14508x);
	defparam lut_7921.LUT_SIZE = 7;
	defparam lut_7921.mask = 128'h33ff77ff33ff77ff7fff7fff7fffffff;

	lut_sub lut_7927 ({sk[1718], i_9_, i_7_, i_8_, i_6_, n_n536, n_n491}, x14511x);
	defparam lut_7927.LUT_SIZE = 7;
	defparam lut_7927.mask = 128'h33ff77ff33ff77ff0101011101011010;

	lut_sub lut_7937 ({sk[1719], i_9_, i_7_, i_8_, i_6_, n_n455, n_n535}, x14529x);
	defparam lut_7937.LUT_SIZE = 7;
	defparam lut_7937.mask = 128'h33ff33ffffffffff0100010001001001;

	lut_sub lut_7943 ({sk[1720], x15x, x13x, x549x, x540x, x548x}, x22303x);
	defparam lut_7943.LUT_SIZE = 6;
	defparam lut_7943.mask = 64'h77ff77ffffa0cc80;

	lut_sub lut_7948 ({sk[1721], x15x, x11x, x12x, x475x, x486x}, n_n2685);
	defparam lut_7948.LUT_SIZE = 6;
	defparam lut_7948.mask = 64'h77ff77ff03575757;

	lut_sub lut_7952 ({sk[1722], x12x, x482x, x23x, x598x, x481x, x480x}, x13929x);
	defparam lut_7952.LUT_SIZE = 7;
	defparam lut_7952.mask = 128'h33ff33ffffffffff000f000f777fffff;

	lut_sub lut_7957 ({sk[1723], x25x, x20x, x598x, x486x, n_n2685, x13929x}, n_n3308);
	defparam lut_7957.LUT_SIZE = 7;
	defparam lut_7957.mask = 128'h33ff33ffffffffff777777ff7f7f7fff;

	lut_sub lut_7962 ({sk[1724], i_9_, i_7_, i_8_, i_6_, n_n464, n_n65}, x13947x);
	defparam lut_7962.LUT_SIZE = 7;
	defparam lut_7962.mask = 128'h33ff33ffffffffff0101011001011110;

	lut_sub lut_7972 ({sk[1725], x19x, x20x, x494x, x599x}, x386x);
	defparam lut_7972.LUT_SIZE = 5;
	defparam lut_7972.mask = 32'h33330537;

	lut_sub lut_7975 ({sk[1726], x25x, x21x, x599x, x487x, n_n5232, n_n5234}, x22173x);
	defparam lut_7975.LUT_SIZE = 7;
	defparam lut_7975.mask = 128'h33ff33ffffffffff8888880080808000;

	lut_sub lut_7980 ({sk[1727], x19x, x477x, x146x, x386x, x22173x}, x13961x);
	defparam lut_7980.LUT_SIZE = 6;
	defparam lut_7980.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_7985 ({sk[1728], i_9_, i_7_, i_8_, i_6_, n_n500, n_n65}, n_n3296);
	defparam lut_7985.LUT_SIZE = 7;
	defparam lut_7985.mask = 128'h33ff33ffffffffff0110110011011100;

	lut_sub lut_7995 ({sk[1729], i_9_, i_7_, i_8_, i_6_, n_n491, n_n65}, x204x);
	defparam lut_7995.LUT_SIZE = 7;
	defparam lut_7995.mask = 128'h33ff33ffffffffff0101010101010000;

	lut_sub lut_8002 ({sk[1730], i_9_, i_7_, i_8_, i_6_, n_n491, n_n65}, n_n3295);
	defparam lut_8002.LUT_SIZE = 7;
	defparam lut_8002.mask = 128'h33ff33ffffffffff0101110101011010;

	lut_sub lut_8012 ({sk[1731], x19x, x492x, x558x, x20x, x579x, n_n5295}, x13972x);
	defparam lut_8012.LUT_SIZE = 7;
	defparam lut_8012.mask = 128'h33ff33ffffffffff5757575757ffffff;

	lut_sub lut_8017 ({sk[1732], i_9_, n_n482, n_n532, n_n534, n_n65, n_n5286}, x13973x);
	defparam lut_8017.LUT_SIZE = 7;
	defparam lut_8017.mask = 128'h33ff33ffffffffff5555577755555777;

	lut_sub lut_8023 ({sk[1733], n_n3296, n_n3295, x13972x, x13973x}, x13976x);
	defparam lut_8023.LUT_SIZE = 5;
	defparam lut_8023.mask = 32'h33337fff;

	lut_sub lut_8028 ({sk[1734], x25x, x599x, x384x, x181x, x22312x}, n_n3299);
	defparam lut_8028.LUT_SIZE = 6;
	defparam lut_8028.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_8033 ({sk[1735], x19x, x508x, x22172x, x22272x}, n_n3293);
	defparam lut_8033.LUT_SIZE = 5;
	defparam lut_8033.mask = 32'h3333eeef;

	lut_sub lut_8037 ({sk[1736], x19x, x11x, x474x, x487x, n_n3385, x13954x}, n_n3297);
	defparam lut_8037.LUT_SIZE = 7;
	defparam lut_8037.mask = 128'h33ff33ffffffffff77777f7f77ff7fff;

	lut_sub lut_8042 ({sk[1737], n_n3292, x13947x, x13961x, n_n3299, n_n3293, n_n3297}, x13977x);
	defparam lut_8042.LUT_SIZE = 7;
	defparam lut_8042.mask = 128'h33ff33ffffffffff7fffffffffffffff;

	lut_sub lut_8049 ({sk[1738], x11x, x12x, x598x, x585x, x559x}, n_n1167);
	defparam lut_8049.LUT_SIZE = 6;
	defparam lut_8049.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_8053 ({sk[1739], x12x, x490x, x20x, x554x, x546x}, n_n783);
	defparam lut_8053.LUT_SIZE = 6;
	defparam lut_8053.mask = 64'h77ff77ff030357ff;

	lut_sub lut_8057 ({sk[1740], x545x, x12x, n_n5087, n_n3412, n_n1167, n_n783}, x14015x);
	defparam lut_8057.LUT_SIZE = 7;
	defparam lut_8057.mask = 128'h0077ffffffffffff7fff7fff7fffffff;

	lut_sub lut_8063 ({sk[1741], x18x, x516x, x489x, x14005x, x22171x}, n_n3311);
	defparam lut_8063.LUT_SIZE = 6;
	defparam lut_8063.mask = 64'h0f0fffffbbbbbfff;

	lut_sub lut_8068 ({sk[1742], x12x, x548x, x34x, x232x, x14008x}, x14014x);
	defparam lut_8068.LUT_SIZE = 6;
	defparam lut_8068.mask = 64'h00ff05ff7f7f7fff;

	lut_sub lut_8073 ({sk[1743], x13991x, x13992x, x14015x, n_n3311, x14014x}, x14025x);
	defparam lut_8073.LUT_SIZE = 6;
	defparam lut_8073.mask = 64'h00ff05ff7fffffff;

	lut_sub lut_8079 ({sk[1744], i_5_, i_3_, i_4_, n_n532, x12x, n_n530}, x14037x);
	defparam lut_8079.LUT_SIZE = 7;
	defparam lut_8079.mask = 128'h0033ffffffffffff0013000000000000;

	lut_sub lut_8082 ({sk[1745], i_9_, n_n473, n_n534, n_n130, x152x}, x14038x);
	defparam lut_8082.LUT_SIZE = 6;
	defparam lut_8082.mask = 64'h00ff05ff55555557;

	lut_sub lut_8085 ({sk[1746], i_9_, i_7_, i_8_, i_6_, n_n482, n_n130}, x14039x);
	defparam lut_8085.LUT_SIZE = 7;
	defparam lut_8085.mask = 128'h0033ffffffffffff0100100110000000;

	lut_sub lut_8090 ({sk[1747], n_n3303, n_n3305, x14037x, x14038x, x14039x}, n_n3267);
	defparam lut_8090.LUT_SIZE = 6;
	defparam lut_8090.mask = 64'h00ff05ff7fffffff;

	lut_sub lut_8096 ({sk[1748], i_9_, i_7_, i_8_, i_6_, n_n130, n_n464}, x14056x);
	defparam lut_8096.LUT_SIZE = 7;
	defparam lut_8096.mask = 128'h0033ffffffffffff0001000001010101;

	lut_sub lut_8102 ({sk[1749], x25x, x11x, x533x, n_n5189, n_n5188, x14056x}, x14057x);
	defparam lut_8102.LUT_SIZE = 7;
	defparam lut_8102.mask = 128'h0033ffffffffffff7f7f7fff7fff7fff;

	lut_sub lut_8108 ({sk[1750], x22x, x12x, x516x, x533x}, x36x);
	defparam lut_8108.LUT_SIZE = 5;
	defparam lut_8108.mask = 32'h1f1f0357;

	lut_sub lut_8111 ({sk[1751], i_9_, i_7_, i_8_, i_6_, n_n535, n_n65}, n_n3300);
	defparam lut_8111.LUT_SIZE = 7;
	defparam lut_8111.mask = 128'h0000ffffffffffff0000111100111110;

	lut_sub lut_8121 ({sk[1752], i_9_, i_7_, i_8_, i_6_, n_n130, n_n464}, x14050x);
	defparam lut_8121.LUT_SIZE = 7;
	defparam lut_8121.mask = 128'h0000ffffffffffff0010100010100010;

	lut_sub lut_8127 ({sk[1753], x36x, x450x, n_n3300, x14050x}, x14058x);
	defparam lut_8127.LUT_SIZE = 5;
	defparam lut_8127.mask = 32'h55ff7fff;

	lut_sub lut_8132 ({sk[1754], x12x, x23x, x574x, x568x, n_n3771, x14061x}, x14063x);
	defparam lut_8132.LUT_SIZE = 7;
	defparam lut_8132.mask = 128'h0000ffffffffffff77777f7f77ff7fff;

	lut_sub lut_8137 ({sk[1755], n_n3307, n_n3308, n_n3267, x14057x, x14058x, x14063x}, x14067x);
	defparam lut_8137.LUT_SIZE = 7;
	defparam lut_8137.mask = 128'h0000ffffffffffff7fffffffffffffff;

	lut_sub lut_8144 ({sk[1756], i_9_, i_7_, i_8_, i_6_, n_n195, n_n500}, x14022x);
	defparam lut_8144.LUT_SIZE = 7;
	defparam lut_8144.mask = 128'h0000ffffffffffff0111110010101010;

	lut_sub lut_8154 ({sk[1757], x103x, x298x, x13996x, x248x, x14000x, x13993x}, x14023x);
	defparam lut_8154.LUT_SIZE = 7;
	defparam lut_8154.mask = 128'h0000ffffffffffff7fffffffffffffff;

	lut_sub lut_8161 ({sk[1758], i_9_, i_1_, i_2_, i_0_, x494x, x585x}, x13765x);
	defparam lut_8161.LUT_SIZE = 7;
	defparam lut_8161.mask = 128'h0000ffffffffffff0000000000007000;

	lut_sub lut_8164 ({sk[1759], x22x, x509x, x510x, x17x, x597x, n_n4959}, x22178x);
	defparam lut_8164.LUT_SIZE = 7;
	defparam lut_8164.mask = 128'h0000ffffffffffffaaa0a0a088808080;

	lut_sub lut_8169 ({sk[1760], x25x, x553x, x351x, x13765x, x22178x}, n_n3199);
	defparam lut_8169.LUT_SIZE = 6;
	defparam lut_8169.mask = 64'h5f5f7f7fbfbfbfff;

	lut_sub lut_8174 ({sk[1761], x24x, x14x, x516x, x522x, x530x, x71x}, x22177x);
	defparam lut_8174.LUT_SIZE = 7;
	defparam lut_8174.mask = 128'h0fffffff0fffffffaaaaa00088888000;

	lut_sub lut_8179 ({sk[1762], x17x, x585x, x548x, x593x, n_n4839, x22177x}, n_n3201);
	defparam lut_8179.LUT_SIZE = 7;
	defparam lut_8179.mask = 128'h0fffffff0fffffffbbbbbbbbbfffffff;

	lut_sub lut_8185 ({sk[1763], x15x, x13x, x557x, x572x, x542x}, n_n3509);
	defparam lut_8185.LUT_SIZE = 6;
	defparam lut_8185.mask = 64'h777777ff003f557f;

	lut_sub lut_8189 ({sk[1764], i_9_, i_7_, i_8_, i_6_, x571x}, n_n1646);
	defparam lut_8189.LUT_SIZE = 6;
	defparam lut_8189.mask = 64'h777777ff11010000;

	lut_sub lut_8193 ({sk[1765], i_9_, i_7_, i_8_, i_6_, n_n473, n_n325}, x15790x);
	defparam lut_8193.LUT_SIZE = 7;
	defparam lut_8193.mask = 128'h0fffffff0fffffff0000000101010001;

	lut_sub lut_8198 ({sk[1766], x15x, x16x, x500x, x558x}, x359x);
	defparam lut_8198.LUT_SIZE = 5;
	defparam lut_8198.mask = 32'h0f0f0537;

	lut_sub lut_8201 ({sk[1767], x19x, x22x, x539x, x599x}, x182x);
	defparam lut_8201.LUT_SIZE = 5;
	defparam lut_8201.mask = 32'h0f0f0537;

	lut_sub lut_8204 ({sk[1768], x25x, x19x, x585x, x599x}, x383x);
	defparam lut_8204.LUT_SIZE = 5;
	defparam lut_8204.mask = 32'h0f0f0357;

	lut_sub lut_8207 ({sk[1769], i_9_, i_7_, i_8_, i_6_, n_n518, n_n65}, n_n2570);
	defparam lut_8207.LUT_SIZE = 7;
	defparam lut_8207.mask = 128'h0fffffff0fffffff0101001101110011;

	lut_sub lut_8217 ({sk[1770], x25x, x19x, x549x, x555x}, x223x);
	defparam lut_8217.LUT_SIZE = 5;
	defparam lut_8217.mask = 32'h0f0f0357;

	lut_sub lut_8220 ({sk[1771], i_9_, i_7_, i_8_, i_6_, x555x}, x384x);
	defparam lut_8220.LUT_SIZE = 6;
	defparam lut_8220.mask = 64'h1f5f1f5f44000000;

	lut_sub lut_8223 ({sk[1772], i_9_, i_7_, i_8_, i_6_, n_n535, n_n65}, x15219x);
	defparam lut_8223.LUT_SIZE = 7;
	defparam lut_8223.mask = 128'h55ff55ff5fff5fff0100101000101010;

	lut_sub lut_8230 ({sk[1773], x19x, x12x, x23x, x525x, x546x, x533x}, x22327x);
	defparam lut_8230.LUT_SIZE = 7;
	defparam lut_8230.mask = 128'h55ff55ff5fff5fffffaaf0a0cc88c080;

	lut_sub lut_8239 ({sk[1774], i_9_, i_7_, i_8_, i_6_, x555x}, x15217x);
	defparam lut_8239.LUT_SIZE = 6;
	defparam lut_8239.mask = 64'h1f5f1f5f45100000;

	lut_sub lut_8244 ({sk[1775], i_9_, i_7_, i_8_, i_6_, n_n455, n_n473}, x15061x);
	defparam lut_8244.LUT_SIZE = 7;
	defparam lut_8244.mask = 128'h55ff55ff5fff5fff0000110000000110;

	lut_sub lut_8249 ({sk[1776], x22x, x16x, x21x, x516x, x496x}, n_n910);
	defparam lut_8249.LUT_SIZE = 6;
	defparam lut_8249.mask = 64'h1f5f1f5f05375577;

	lut_sub lut_8253 ({sk[1777], i_9_, i_7_, i_8_, i_6_, x540x, x496x}, x15072x);
	defparam lut_8253.LUT_SIZE = 7;
	defparam lut_8253.mask = 128'h55ff55ff5fff5fff5000030000000000;

	lut_sub lut_8256 ({sk[1778], x25x, x15x, x236x, x540x, n_n910, x15072x}, x15075x);
	defparam lut_8256.LUT_SIZE = 7;
	defparam lut_8256.mask = 128'h55ff55ff5fff5fff77ff7fff7fff7fff;

	lut_sub lut_8262 ({sk[1779], x13x, x539x, x544x, x20x, x482x, x23x}, x15069x);
	defparam lut_8262.LUT_SIZE = 7;
	defparam lut_8262.mask = 128'h55ff55ff5fff5fff005f005f337fffff;

	lut_sub lut_8267 ({sk[1780], i_9_, i_7_, i_8_, i_6_, n_n518, n_n455}, x15070x);
	defparam lut_8267.LUT_SIZE = 7;
	defparam lut_8267.mask = 128'h55ff55ff5fff5fff0000101001101000;

	lut_sub lut_8273 ({sk[1781], i_9_, i_1_, i_2_, i_0_, x594x, x593x}, x15063x);
	defparam lut_8273.LUT_SIZE = 7;
	defparam lut_8273.mask = 128'h0055ffffffffffff0000000000000700;

	lut_sub lut_8276 ({sk[1782], x22x, x21x, x13x, x545x, x540x}, x15064x);
	defparam lut_8276.LUT_SIZE = 6;
	defparam lut_8276.mask = 64'h1f1fffff03575757;

	lut_sub lut_8280 ({sk[1783], x128x, x291x, x15069x, x15070x, x15063x, x15064x}, x15076x);
	defparam lut_8280.LUT_SIZE = 7;
	defparam lut_8280.mask = 128'h0055ffffffffffff7fffffffffffffff;

	lut_sub lut_8287 ({sk[1784], x13x, x478x, x23x, x564x, x476x}, n_n1677);
	defparam lut_8287.LUT_SIZE = 6;
	defparam lut_8287.mask = 64'h1f1fffff050537ff;

	lut_sub lut_8291 ({sk[1785], i_9_, i_7_, i_8_, i_6_, n_n455, n_n509}, n_n2629);
	defparam lut_8291.LUT_SIZE = 7;
	defparam lut_8291.mask = 128'h0055ffffffffffff0011101100101110;

	lut_sub lut_8301 ({sk[1786], i_9_, i_7_, i_8_, i_6_, n_n455, n_n500}, x15093x);
	defparam lut_8301.LUT_SIZE = 7;
	defparam lut_8301.mask = 128'h0055ffffffffffff0101101110001100;

	lut_sub lut_8310 ({sk[1787], x25x, x13x, x24x, x542x, x562x, n_n4501}, x22141x);
	defparam lut_8310.LUT_SIZE = 7;
	defparam lut_8310.mask = 128'h0055ffffffffffffaaa08880a0a08080;

	lut_sub lut_8315 ({sk[1788], n_n3509, n_n1677, n_n2629, x15093x, x22141x}, n_n2557);
	defparam lut_8315.LUT_SIZE = 6;
	defparam lut_8315.mask = 64'h1f1fffffbfffffff;

	lut_sub lut_8321 ({sk[1789], x22x, x13x, x520x, x543x}, x178x);
	defparam lut_8321.LUT_SIZE = 5;
	defparam lut_8321.mask = 32'h1f1f0357;

	lut_sub lut_8324 ({sk[1790], i_9_, i_7_, i_8_, i_6_, n_n482, n_n455}, x15101x);
	defparam lut_8324.LUT_SIZE = 7;
	defparam lut_8324.mask = 128'h5577ffff5577ffff0000111011101110;

	lut_sub lut_8334 ({sk[1791], x25x, x15x, x504x, x15061x, x22139x, x22140x}, x15102x);
	defparam lut_8334.LUT_SIZE = 7;
	defparam lut_8334.mask = 128'h5577ffff5577ffffefefefffefffefff;

	lut_sub lut_8340 ({sk[1792], i_9_, i_7_, i_8_, i_6_, n_n390, n_n535}, n_n2621);
	defparam lut_8340.LUT_SIZE = 7;
	defparam lut_8340.mask = 128'h5577ffff5577ffff0111001011101010;

	lut_sub lut_8350 ({sk[1793], x11x, x10x, x519x, x561x}, x15134x);
	defparam lut_8350.LUT_SIZE = 5;
	defparam lut_8350.mask = 32'h1f1f0357;

	lut_sub lut_8353 ({sk[1794], x11x, x10x, x24x, x571x, x557x, x537x}, x22305x);
	defparam lut_8353.LUT_SIZE = 7;
	defparam lut_8353.mask = 128'h5577ffff5577fffffff08880f0f08080;

	lut_sub lut_8358 ({sk[1795], x10x, x573x, n_n2761, x15134x, x22305x}, x15140x);
	defparam lut_8358.LUT_SIZE = 6;
	defparam lut_8358.mask = 64'h555f555fbfbfbfff;

	lut_sub lut_8363 ({sk[1796], i_9_, i_7_, i_8_, i_6_, n_n482, n_n390}, n_n2615);
	defparam lut_8363.LUT_SIZE = 7;
	defparam lut_8363.mask = 128'h5577ffff5577ffff1110111101010000;

	lut_sub lut_8373 ({sk[1797], i_9_, n_n390, n_n491, n_n530, x357x}, x15135x);
	defparam lut_8373.LUT_SIZE = 6;
	defparam lut_8373.mask = 64'h555f555f55575557;

	lut_sub lut_8377 ({sk[1798], x22x, x21x, x561x, x571x, n_n2615, x15135x}, x15141x);
	defparam lut_8377.LUT_SIZE = 7;
	defparam lut_8377.mask = 128'h5577ffff5577ffff77777fff7fff7fff;

	lut_sub lut_8384 ({sk[1799], x25x, x13x, x529x, x523x, x528x}, x82x);
	defparam lut_8384.LUT_SIZE = 6;
	defparam lut_8384.mask = 64'h0fff0fff005f337f;

	lut_sub lut_8388 ({sk[1800], x23x, x504x, x212x, n_n2621, x121x, x15142x}, x15149x);
	defparam lut_8388.LUT_SIZE = 7;
	defparam lut_8388.mask = 128'h33ff3fffffffffff7fff7fff7fffffff;

	lut_sub lut_8394 ({sk[1801], x13x, x24x, x516x, x525x, x523x, n_n4572}, x22253x);
	defparam lut_8394.LUT_SIZE = 7;
	defparam lut_8394.mask = 128'h33ff3fffffffffffaaaa8888a0008000;

	lut_sub lut_8399 ({sk[1802], x25x, x10x, x479x, x481x, x45x, x15109x}, n_n2619);
	defparam lut_8399.LUT_SIZE = 7;
	defparam lut_8399.mask = 128'h33ff3fffffffffff77777f7f77ff7fff;

	lut_sub lut_8404 ({sk[1803], x10x, x562x, x22251x, x22252x}, n_n2618);
	defparam lut_8404.LUT_SIZE = 5;
	defparam lut_8404.mask = 32'h3333eeef;

	lut_sub lut_8408 ({sk[1804], x521x, x10x, x23x, x547x, x585x, x593x}, x15119x);
	defparam lut_8408.LUT_SIZE = 7;
	defparam lut_8408.mask = 128'h55555f5f555f5f5f000f777f000fffff;

	lut_sub lut_8413 ({sk[1805], i_9_, i_7_, i_8_, i_6_, n_n518, n_n390}, x15120x);
	defparam lut_8413.LUT_SIZE = 7;
	defparam lut_8413.mask = 128'h55555f5f555f5f5f0110100101000000;

	lut_sub lut_8419 ({sk[1806], i_9_, i_7_, i_8_, i_6_, n_n536, n_n518}, n_n2640);
	defparam lut_8419.LUT_SIZE = 7;
	defparam lut_8419.mask = 128'h55555f5f555f5f5f0101101101011010;

	lut_sub lut_8429 ({sk[1807], i_9_, i_7_, i_8_, i_6_, n_n536, n_n535}, n_n2641);
	defparam lut_8429.LUT_SIZE = 7;
	defparam lut_8429.mask = 128'h55555f5f555f5f5f1110011010101100;

	lut_sub lut_8439 ({sk[1808], x25x, x16x, x481x, x473x}, x337x);
	defparam lut_8439.LUT_SIZE = 5;
	defparam lut_8439.mask = 32'h0f5f0357;

	lut_sub lut_8442 ({sk[1809], x19x, x11x, x537x, x579x}, x217x);
	defparam lut_8442.LUT_SIZE = 5;
	defparam lut_8442.mask = 32'h0f5f0537;

	lut_sub lut_8445 ({sk[1810], x12x, x23x, x514x, x529x}, x89x);
	defparam lut_8445.LUT_SIZE = 5;
	defparam lut_8445.mask = 32'h0f5f0357;

	lut_sub lut_8448 ({sk[1811], i_9_, n_n130, x23x, n_n500, x560x}, x288x);
	defparam lut_8448.LUT_SIZE = 6;
	defparam lut_8448.mask = 64'h00ff77ff00030057;

	lut_sub lut_8451 ({sk[1812], i_9_, n_n522, n_n130, x23x, n_n500, x560x}, x12265x);
	defparam lut_8451.LUT_SIZE = 7;
	defparam lut_8451.mask = 128'h55555f5f555f5f5f0003003300570077;

	lut_sub lut_8456 ({sk[1813], x19x, x22x, x475x, x487x}, x446x);
	defparam lut_8456.LUT_SIZE = 5;
	defparam lut_8456.mask = 32'h0f5f0537;

	lut_sub lut_8459 ({sk[1814], x19x, x24x, x478x, x569x}, x12346x);
	defparam lut_8459.LUT_SIZE = 5;
	defparam lut_8459.mask = 32'h0f5f0537;

	lut_sub lut_8462 ({sk[1815], x11x, x487x, n_n3031, n_n5257, x446x, x12346x}, n_n1435);
	defparam lut_8462.LUT_SIZE = 7;
	defparam lut_8462.mask = 128'h55555f5f555f5f5f7fff7fff7fffffff;

	lut_sub lut_8468 ({sk[1816], x25x, x10x, x529x, x528x, x526x}, n_n1636);
	defparam lut_8468.LUT_SIZE = 6;
	defparam lut_8468.mask = 64'h00ff77ff003f557f;

	lut_sub lut_8472 ({sk[1817], x25x, x24x, x18x, x572x, x518x, x577x}, x11986x);
	defparam lut_8472.LUT_SIZE = 7;
	defparam lut_8472.mask = 128'h55555f5f555f5f5f003f557f557f557f;

	lut_sub lut_8477 ({sk[1818], i_9_, i_7_, i_8_, i_6_, n_n195, n_n500}, x11987x);
	defparam lut_8477.LUT_SIZE = 7;
	defparam lut_8477.mask = 128'h55555f5f555f5f5f1100001010100000;

	lut_sub lut_8483 ({sk[1819], x15x, x19x, x585x, x599x}, x181x);
	defparam lut_8483.LUT_SIZE = 5;
	defparam lut_8483.mask = 32'h0f5f0357;

	lut_sub lut_8486 ({sk[1820], i_9_, x490x, n_n65, x548x, x181x}, x11967x);
	defparam lut_8486.LUT_SIZE = 6;
	defparam lut_8486.mask = 64'h00ff77ff5555575f;

	lut_sub lut_8490 ({sk[1821], x25x, x24x, x12x, x528x, x533x}, n_n1927);
	defparam lut_8490.LUT_SIZE = 6;
	defparam lut_8490.mask = 64'h00ff77ff03575757;

	lut_sub lut_8494 ({sk[1822], i_9_, n_n522, n_n130, x514x, x506x}, x188x);
	defparam lut_8494.LUT_SIZE = 6;
	defparam lut_8494.mask = 64'h00ff77ff00330505;

	lut_sub lut_8497 ({sk[1823], x12x, x20x, x514x, x506x, x524x, x527x}, x11970x);
	defparam lut_8497.LUT_SIZE = 7;
	defparam lut_8497.mask = 128'h55555f5f555f5f5f000000ff7f7f7fff;

	lut_sub lut_8502 ({sk[1824], i_9_, i_1_, i_2_, i_0_, x550x, x549x}, x11973x);
	defparam lut_8502.LUT_SIZE = 7;
	defparam lut_8502.mask = 128'h55555f5f555f5f5f0000000070000000;

	lut_sub lut_8505 ({sk[1825], i_9_, i_7_, i_8_, i_6_, n_n130, n_n464}, x11975x);
	defparam lut_8505.LUT_SIZE = 7;
	defparam lut_8505.mask = 128'h55555f5f555f5f5f1000101000001000;

	lut_sub lut_8510 ({sk[1826], i_9_, i_1_, i_2_, i_0_, x522x, x488x}, x11969x);
	defparam lut_8510.LUT_SIZE = 7;
	defparam lut_8510.mask = 128'h55555f5f555f5f5f0000000000700000;

	lut_sub lut_8513 ({sk[1827], x25x, x11x, x599x, x555x, n_n5226, x384x}, x22245x);
	defparam lut_8513.LUT_SIZE = 7;
	defparam lut_8513.mask = 128'h55555f5f555f5f5f8888808088008000;

	lut_sub lut_8518 ({sk[1828], x25x, x22x, x541x, x543x, n_n4504, n_n4517}, x22249x);
	defparam lut_8518.LUT_SIZE = 7;
	defparam lut_8518.mask = 128'h55555f5f555f5f5f8888880080808000;

	lut_sub lut_8523 ({sk[1829], x13x, x23x, x587x, x542x}, x307x);
	defparam lut_8523.LUT_SIZE = 5;
	defparam lut_8523.mask = 32'h0f5f0537;

	lut_sub lut_8526 ({sk[1830], i_9_, i_7_, i_8_, i_6_, n_n455, n_n500}, x11497x);
	defparam lut_8526.LUT_SIZE = 7;
	defparam lut_8526.mask = 128'h33337777777777770111000010000000;

	lut_sub lut_8531 ({sk[1831], i_9_, n_n455, x544x, n_n534, n_n509, x23x}, x11516x);
	defparam lut_8531.LUT_SIZE = 7;
	defparam lut_8531.mask = 128'h33337777777777770055135700551357;

	lut_sub lut_8536 ({sk[1832], i_9_, i_7_, i_8_, i_6_, n_n518, n_n455}, n_n1111);
	defparam lut_8536.LUT_SIZE = 7;
	defparam lut_8536.mask = 128'h33337777777777770101010101010111;

	lut_sub lut_8546 ({sk[1833], x21x, x13x, x20x, x472x, x476x}, x11511x);
	defparam lut_8546.LUT_SIZE = 6;
	defparam lut_8546.mask = 64'h0000ffff05375577;

	lut_sub lut_8550 ({sk[1834], x25x, x13x, x478x, x541x}, x11510x);
	defparam lut_8550.LUT_SIZE = 5;
	defparam lut_8550.mask = 32'h03ff0357;

	lut_sub lut_8553 ({sk[1835], i_9_, i_7_, i_8_, i_6_, n_n455, n_n535}, n_n1112);
	defparam lut_8553.LUT_SIZE = 7;
	defparam lut_8553.mask = 128'h33337777777777770011101011101010;

	lut_sub lut_8563 ({sk[1836], x15x, x10x, x24x, x571x, x587x, x491x}, x11555x);
	defparam lut_8563.LUT_SIZE = 7;
	defparam lut_8563.mask = 128'h3333777777777777000f777f0f0f7f7f;

	lut_sub lut_8568 ({sk[1837], x21x, x11x, x23x, x583x, x547x, n_n4592}, x22247x);
	defparam lut_8568.LUT_SIZE = 7;
	defparam lut_8568.mask = 128'h3333777777777777aa88a08088888080;

	lut_sub lut_8573 ({sk[1838], i_9_, i_7_, i_8_, i_6_, n_n518, n_n390}, x11570x);
	defparam lut_8573.LUT_SIZE = 7;
	defparam lut_8573.mask = 128'h33337777777777770001001000011000;

	lut_sub lut_8578 ({sk[1839], i_9_, i_7_, i_8_, i_6_, n_n390, n_n535}, x11571x);
	defparam lut_8578.LUT_SIZE = 7;
	defparam lut_8578.mask = 128'h33337777777777770001000110001000;

	lut_sub lut_8583 ({sk[1840], i_9_, i_7_, i_8_, i_6_, n_n536, n_n535}, n_n1123);
	defparam lut_8583.LUT_SIZE = 7;
	defparam lut_8583.mask = 128'h33337777777777770001011101010111;

	lut_sub lut_8593 ({sk[1841], i_9_, i_7_, i_8_, i_6_, n_n536, n_n482}, x11602x);
	defparam lut_8593.LUT_SIZE = 7;
	defparam lut_8593.mask = 128'h33337777777777770100000000010011;

	lut_sub lut_8598 ({sk[1842], x21x, x500x, x11x, x23x, n_n4404, x495x}, x22242x);
	defparam lut_8598.LUT_SIZE = 7;
	defparam lut_8598.mask = 128'h3333777777777777cc88c080cc880000;

	lut_sub lut_8603 ({sk[1843], x15x, x16x, x24x, x510x, x508x, x495x}, x22261x);
	defparam lut_8603.LUT_SIZE = 7;
	defparam lut_8603.mask = 128'h3333777777777777ffaac080aaaa8080;

	lut_sub lut_8608 ({sk[1844], i_9_, i_7_, i_8_, i_6_, n_n536, n_n500}, x11618x);
	defparam lut_8608.LUT_SIZE = 7;
	defparam lut_8608.mask = 128'h33337777777777771101011001011111;

	lut_sub lut_8620 ({sk[1845], i_9_, i_7_, i_8_, i_6_, n_n536, n_n518}, x11626x);
	defparam lut_8620.LUT_SIZE = 7;
	defparam lut_8620.mask = 128'h33337777777777770110100010001000;

	lut_sub lut_8626 ({sk[1846], i_9_, i_1_, i_2_, i_0_, x538x, x558x}, x12638x);
	defparam lut_8626.LUT_SIZE = 7;
	defparam lut_8626.mask = 128'h33337777777777770000000000700000;

	lut_sub lut_8629 ({sk[1847], x11x, x12x, x514x, x505x, x489x, n_n5173}, x22218x);
	defparam lut_8629.LUT_SIZE = 7;
	defparam lut_8629.mask = 128'h3333777777777777aaaa8080aa008000;

	lut_sub lut_8634 ({sk[1848], x15x, x10x, x520x, x582x}, x312x);
	defparam lut_8634.LUT_SIZE = 5;
	defparam lut_8634.mask = 32'h03ff0357;

	lut_sub lut_8637 ({sk[1849], x10x, x509x, x24x, x507x, x510x, x580x}, x22185x);
	defparam lut_8637.LUT_SIZE = 7;
	defparam lut_8637.mask = 128'h3333777777777777fff0fff088800000;

	lut_sub lut_8642 ({sk[1850], x11x, x17x, x566x, x556x}, x330x);
	defparam lut_8642.LUT_SIZE = 5;
	defparam lut_8642.mask = 32'h03ff0537;

	lut_sub lut_8645 ({sk[1851], i_9_, i_7_, i_8_, i_6_, n_n455, n_n500}, n_n3355);
	defparam lut_8645.LUT_SIZE = 7;
	defparam lut_8645.mask = 128'h33337777777777770111001011101010;

	lut_sub lut_8655 ({sk[1852], i_9_, i_7_, i_8_, i_6_, n_n455, n_n491}, x14202x);
	defparam lut_8655.LUT_SIZE = 7;
	defparam lut_8655.mask = 128'h33337777777777770000001100000110;

	lut_sub lut_8660 ({sk[1853], x13x, x519x, x130x, n_n4246, x14205x}, x14207x);
	defparam lut_8660.LUT_SIZE = 6;
	defparam lut_8660.mask = 64'h0000ffff7f7f7fff;

	lut_sub lut_8665 ({sk[1854], x11x, x542x, n_n4503, n_n3509, n_n3355, x14202x}, x14208x);
	defparam lut_8665.LUT_SIZE = 7;
	defparam lut_8665.mask = 128'h33337777777777777fff7fff7fffffff;

	lut_sub lut_8671 ({sk[1855], x14131x, x14132x, x14147x, x14148x, x14207x, x14208x}, x14211x);
	defparam lut_8671.LUT_SIZE = 7;
	defparam lut_8671.mask = 128'h33337777777777777fffffffffffffff;

	lut_sub lut_8678 ({sk[1856], i_9_, n_n526, n_n482, n_n455, n_n532, n_n491}, x15440x);
	defparam lut_8678.LUT_SIZE = 7;
	defparam lut_8678.mask = 128'h33337777777777770003050700030507;

	lut_sub lut_8683 ({sk[1857], i_9_, i_7_, i_8_, i_6_, n_n325, n_n500}, x15761x);
	defparam lut_8683.LUT_SIZE = 7;
	defparam lut_8683.mask = 128'h33337777777777771100000011000010;

	lut_sub lut_8689 ({sk[1858], i_9_, i_7_, i_8_, i_6_, n_n260, n_n491}, n_n2968);
	defparam lut_8689.LUT_SIZE = 7;
	defparam lut_8689.mask = 128'h33337777777777771001010110110110;

	lut_sub lut_8699 ({sk[1859], x19x, x11x, x545x, x535x, x555x}, n_n3037);
	defparam lut_8699.LUT_SIZE = 6;
	defparam lut_8699.mask = 64'h0000ffff00553f7f;

	lut_sub lut_8703 ({sk[1860], i_9_, i_1_, i_2_, i_0_, x522x, x525x}, x15551x);
	defparam lut_8703.LUT_SIZE = 7;
	defparam lut_8703.mask = 128'h33337777777777770000000000700000;

	lut_sub lut_8706 ({sk[1861], i_9_, i_7_, i_8_, i_6_, x533x, x555x}, x15552x);
	defparam lut_8706.LUT_SIZE = 7;
	defparam lut_8706.mask = 128'h33337777777777770300000500000000;

	lut_sub lut_8709 ({sk[1862], x12x, x516x, x220x, x450x, x15551x, x15552x}, n_n2945);
	defparam lut_8709.LUT_SIZE = 7;
	defparam lut_8709.mask = 128'h33337777777777777fff7fff7fffffff;

	lut_sub lut_8715 ({sk[1863], i_9_, i_7_, i_8_, i_6_, x555x}, x183x);
	defparam lut_8715.LUT_SIZE = 6;
	defparam lut_8715.mask = 64'h0000ffff04400000;

	lut_sub lut_8718 ({sk[1864], x11x, x12x, x514x, x488x}, x15556x);
	defparam lut_8718.LUT_SIZE = 5;
	defparam lut_8718.mask = 32'h03ff0537;

	lut_sub lut_8721 ({sk[1865], x21x, x12x, x514x, x502x, x524x}, x15558x);
	defparam lut_8721.LUT_SIZE = 6;
	defparam lut_8721.mask = 64'h0000ffff00770f7f;

	lut_sub lut_8725 ({sk[1866], x19x, x490x, x549x, n_n3037, x15556x, x15558x}, x15564x);
	defparam lut_8725.LUT_SIZE = 7;
	defparam lut_8725.mask = 128'h33337777777777777f7f7f7f7fffffff;

	lut_sub lut_8731 ({sk[1867], i_9_, i_7_, i_8_, i_6_, n_n518, n_n65}, x15570x);
	defparam lut_8731.LUT_SIZE = 7;
	defparam lut_8731.mask = 128'h33337777777777770000010100010101;

	lut_sub lut_8737 ({sk[1868], i_9_, i_7_, i_8_, i_6_, x487x, x433x}, n_n3385);
	defparam lut_8737.LUT_SIZE = 7;
	defparam lut_8737.mask = 128'h33337777777777777555555555555555;

	lut_sub lut_8740 ({sk[1869], i_9_, i_7_, i_8_, i_6_, x599x, x555x}, x15566x);
	defparam lut_8740.LUT_SIZE = 7;
	defparam lut_8740.mask = 128'h33337777777777775003000000000000;

	lut_sub lut_8743 ({sk[1870], i_9_, n_n532, n_n500, n_n65, x446x}, x15574x);
	defparam lut_8743.LUT_SIZE = 6;
	defparam lut_8743.mask = 64'h0000ffff55575557;

	lut_sub lut_8747 ({sk[1871], x319x, x146x, x182x, x15570x, x15566x, x15574x}, x15579x);
	defparam lut_8747.LUT_SIZE = 7;
	defparam lut_8747.mask = 128'h33337777777777777fffffffffffffff;

	lut_sub lut_8754 ({sk[1872], x11x, x24x, x591x, n_n5172, x15580x, x15581x}, n_n2948);
	defparam lut_8754.LUT_SIZE = 7;
	defparam lut_8754.mask = 128'h33337777777777777f7f7fff7fff7fff;

	lut_sub lut_8760 ({sk[1873], x22x, x12x, x573x, x578x, x537x, n_n5139}, x22128x);
	defparam lut_8760.LUT_SIZE = 7;
	defparam lut_8760.mask = 128'h3333777777777777aaaa8800a0a08000;

	lut_sub lut_8765 ({sk[1874], x11x, x578x, x76x, x126x, x22128x}, n_n2949);
	defparam lut_8765.LUT_SIZE = 6;
	defparam lut_8765.mask = 64'h0000ffffbfbfbfff;

	lut_sub lut_8770 ({sk[1875], x24x, x20x, x591x, x514x, x44x, x15591x}, x15592x);
	defparam lut_8770.LUT_SIZE = 7;
	defparam lut_8770.mask = 128'h3333777777777777777777ff7f7f7fff;

	lut_sub lut_8775 ({sk[1876], n_n3031, x454x, x89x, n_n3385, x15560x, x15575x}, x22127x);
	defparam lut_8775.LUT_SIZE = 7;
	defparam lut_8775.mask = 128'h33337777777777778000000000000000;

	lut_sub lut_8777 ({sk[1877], i_9_, i_7_, i_8_, i_6_, x507x}, x80x);
	defparam lut_8777.LUT_SIZE = 6;
	defparam lut_8777.mask = 64'h0000ffff04400000;

	lut_sub lut_8780 ({sk[1878], x15x, x10x, x507x, x508x}, x157x);
	defparam lut_8780.LUT_SIZE = 5;
	defparam lut_8780.mask = 32'h03ff0537;

	lut_sub lut_8783 ({sk[1879], x15x, x11x, x558x, x17x, x589x}, n_n2718);
	defparam lut_8783.LUT_SIZE = 6;
	defparam lut_8783.mask = 64'h0000ffff03575757;

	lut_sub lut_8787 ({sk[1880], i_9_, i_7_, i_8_, i_6_, n_n473, n_n195}, n_n2584);
	defparam lut_8787.LUT_SIZE = 7;
	defparam lut_8787.mask = 128'h7777ffff7777ffff0111001000111110;

	lut_sub lut_8797 ({sk[1881], x25x, x12x, x517x, x532x}, x15229x);
	defparam lut_8797.LUT_SIZE = 5;
	defparam lut_8797.mask = 32'h3f3f0357;

	lut_sub lut_8800 ({sk[1882], x12x, x550x, n_n4152, x13387x, x209x, x15229x}, x15234x);
	defparam lut_8800.LUT_SIZE = 7;
	defparam lut_8800.mask = 128'h7777ffff7777ffff7fff7fff7fffffff;

	lut_sub lut_8806 ({sk[1883], i_9_, i_1_, i_2_, i_0_, x549x, x524x}, x15228x);
	defparam lut_8806.LUT_SIZE = 7;
	defparam lut_8806.mask = 128'h7777ffff7777ffff0000000000305000;

	lut_sub lut_8809 ({sk[1884], x344x, x123x, x159x, n_n2584, x15228x}, x15235x);
	defparam lut_8809.LUT_SIZE = 6;
	defparam lut_8809.mask = 64'h5557ffff7fffffff;

	lut_sub lut_8815 ({sk[1885], i_9_, n_n534, x474x, n_n130, x472x, n_n500}, x15239x);
	defparam lut_8815.LUT_SIZE = 7;
	defparam lut_8815.mask = 128'h7777ffff7777ffff00000505030f070f;

	lut_sub lut_8820 ({sk[1886], i_9_, i_7_, i_8_, i_6_, n_n509, n_n130}, x15240x);
	defparam lut_8820.LUT_SIZE = 7;
	defparam lut_8820.mask = 128'h7777ffff7777ffff0111000010000010;

	lut_sub lut_8826 ({sk[1887], x12x, n_n4148, x494x, x546x, x11914x, x11915x}, x15249x);
	defparam lut_8826.LUT_SIZE = 7;
	defparam lut_8826.mask = 128'h7777ffff7777ffff7777ffff7fffffff;

	lut_sub lut_8832 ({sk[1888], i_9_, n_n534, n_n195, x513x, x584x, x253x}, x15254x);
	defparam lut_8832.LUT_SIZE = 7;
	defparam lut_8832.mask = 128'h7777ffff7777ffff55555f5f55775577;

	lut_sub lut_8836 ({sk[1889], i_9_, i_7_, i_8_, i_6_, n_n482, n_n195}, x15255x);
	defparam lut_8836.LUT_SIZE = 7;
	defparam lut_8836.mask = 128'h7777ffff7777ffff0101100010100000;

	lut_sub lut_8842 ({sk[1890], i_9_, i_7_, i_8_, i_6_, n_n491, n_n195}, n_n2586);
	defparam lut_8842.LUT_SIZE = 7;
	defparam lut_8842.mask = 128'h7777ffff7777ffff1110101010101010;

	lut_sub lut_8852 ({sk[1891], i_9_, i_7_, i_8_, i_6_, x577x}, x297x);
	defparam lut_8852.LUT_SIZE = 6;
	defparam lut_8852.mask = 64'h5557ffff01010000;

	lut_sub lut_8855 ({sk[1892], x22x, x18x, x567x, x536x}, x394x);
	defparam lut_8855.LUT_SIZE = 5;
	defparam lut_8855.mask = 32'h3f3f0537;

	lut_sub lut_8858 ({sk[1893], x21x, n_n5022, x567x, n_n3427, x297x, x394x}, x15262x);
	defparam lut_8858.LUT_SIZE = 7;
	defparam lut_8858.mask = 128'h7777ffff7777ffff7f7fffff7fffffff;

	lut_sub lut_8864 ({sk[1894], x15239x, x15240x, x15254x, x15255x, n_n2586, x15248x}, x22136x);
	defparam lut_8864.LUT_SIZE = 7;
	defparam lut_8864.mask = 128'h7777ffff7777ffff8000000000000000;

	lut_sub lut_8866 ({sk[1895], x25x, x538x, x10x, x493x, x551x, x526x}, x14855x);
	defparam lut_8866.LUT_SIZE = 7;
	defparam lut_8866.mask = 128'h7777ffff7777ffff000f00ff777f77ff;

	lut_sub lut_8871 ({sk[1896], x22x, x10x, x507x, x516x, x489x}, x14854x);
	defparam lut_8871.LUT_SIZE = 6;
	defparam lut_8871.mask = 64'h5557ffff00770f7f;

	lut_sub lut_8875 ({sk[1897], x25x, x507x, x14x, x490x, x14855x, x14854x}, n_n2467);
	defparam lut_8875.LUT_SIZE = 7;
	defparam lut_8875.mask = 128'h7777ffff7777ffff777f777f777fffff;

	lut_sub lut_8880 ({sk[1898], i_9_, i_7_, i_8_, i_6_, x483x, x595x}, x14858x);
	defparam lut_8880.LUT_SIZE = 7;
	defparam lut_8880.mask = 128'h7777ffff7777ffff0053000000000000;

	lut_sub lut_8883 ({sk[1899], x11x, x483x, x14x, x494x, x593x, x370x}, x22129x);
	defparam lut_8883.LUT_SIZE = 7;
	defparam lut_8883.mask = 128'h7777ffff7777ffffaa80aa80aa800000;

	lut_sub lut_8888 ({sk[1900], x25x, x24x, x565x, x14858x, x22129x}, n_n2466);
	defparam lut_8888.LUT_SIZE = 6;
	defparam lut_8888.mask = 64'h5557ffffbbbfbfbf;

	lut_sub lut_8893 ({sk[1901], x13x, x11x, x558x, x543x}, x378x);
	defparam lut_8893.LUT_SIZE = 5;
	defparam lut_8893.mask = 32'h3f3f0537;

	lut_sub lut_8896 ({sk[1902], x24x, x18x, x567x, x562x, x556x}, n_n801);
	defparam lut_8896.LUT_SIZE = 6;
	defparam lut_8896.mask = 64'h5557ffff00770f7f;

	lut_sub lut_8900 ({sk[1903], i_9_, n_n524, n_n195, x20x, n_n500, x491x}, x405x);
	defparam lut_8900.LUT_SIZE = 7;
	defparam lut_8900.mask = 128'h5555ffff5555ffff0003003300570077;

	lut_sub lut_8905 ({sk[1904], i_9_, i_7_, i_8_, i_6_, n_n195, n_n500}, n_n1454);
	defparam lut_8905.LUT_SIZE = 7;
	defparam lut_8905.mask = 128'h5555ffff5555ffff0110110001111010;

	lut_sub lut_8915 ({sk[1905], x25x, x19x, x477x, x481x, x487x}, x12352x);
	defparam lut_8915.LUT_SIZE = 6;
	defparam lut_8915.mask = 64'h3333ffff003f557f;

	lut_sub lut_8919 ({sk[1906], x15x, x19x, x21x, x482x, x599x, x487x}, x22278x);
	defparam lut_8919.LUT_SIZE = 7;
	defparam lut_8919.mask = 128'h5555ffff5555ffffffccf0c0aa88a080;

	lut_sub lut_8928 ({sk[1907], x24x, x487x, x320x, x12352x, x22278x}, n_n1436);
	defparam lut_8928.LUT_SIZE = 6;
	defparam lut_8928.mask = 64'h3333ffffbfbfbfff;

	lut_sub lut_8933 ({sk[1908], x16x, x21x, x522x, x496x}, x235x);
	defparam lut_8933.LUT_SIZE = 5;
	defparam lut_8933.mask = 32'h3f3f0537;

	lut_sub lut_8936 ({sk[1909], x13x, x24x, x549x, x540x}, x421x);
	defparam lut_8936.LUT_SIZE = 5;
	defparam lut_8936.mask = 32'h5f5f0537;

	lut_sub lut_8939 ({sk[1910], x10x, x20x, x582x, x493x}, x11856x);
	defparam lut_8939.LUT_SIZE = 5;
	defparam lut_8939.mask = 32'h5f5f0357;

	lut_sub lut_8942 ({sk[1911], i_9_, n_n390, n_n473, n_n534, x23x, x582x}, x11857x);
	defparam lut_8942.LUT_SIZE = 7;
	defparam lut_8942.mask = 128'h37ff37ff3fff3fff1111111f1111111f;

	lut_sub lut_8946 ({sk[1912], i_9_, x22x, n_n390, n_n473, x580x, x157x}, x11859x);
	defparam lut_8946.LUT_SIZE = 7;
	defparam lut_8946.mask = 128'h37ff37ff3fff3fff5555555f5577557f;

	lut_sub lut_8950 ({sk[1913], x21x, x17x, x20x, x491x, x566x}, n_n1985);
	defparam lut_8950.LUT_SIZE = 6;
	defparam lut_8950.mask = 64'h77ff77ff05375577;

	lut_sub lut_8954 ({sk[1914], i_9_, i_7_, i_8_, i_6_, n_n482, n_n195}, x12003x);
	defparam lut_8954.LUT_SIZE = 7;
	defparam lut_8954.mask = 128'h37ff37ff3fff3fff0100111101010101;

	lut_sub lut_8964 ({sk[1915], x11x, x509x, x18x, x513x}, x11988x);
	defparam lut_8964.LUT_SIZE = 5;
	defparam lut_8964.mask = 32'h5f5f0357;

	lut_sub lut_8967 ({sk[1916], i_9_, i_7_, i_8_, i_6_, x590x, x513x}, x11989x);
	defparam lut_8967.LUT_SIZE = 7;
	defparam lut_8967.mask = 128'h37ff37ff3fff3fff0030500000000000;

	lut_sub lut_8970 ({sk[1917], i_9_, i_7_, i_8_, i_6_, n_n518, n_n130}, n_n1061);
	defparam lut_8970.LUT_SIZE = 7;
	defparam lut_8970.mask = 128'h37ff37ff3fff3fff0110111001010101;

	lut_sub lut_8980 ({sk[1918], i_9_, i_7_, i_8_, i_6_, n_n535, n_n130}, x12014x);
	defparam lut_8980.LUT_SIZE = 7;
	defparam lut_8980.mask = 128'h37ff37ff3fff3fff0000001100010100;

	lut_sub lut_8985 ({sk[1919], x24x, x18x, x506x, x488x, x529x, x532x}, x12018x);
	defparam lut_8985.LUT_SIZE = 7;
	defparam lut_8985.mask = 128'h37ff37ff3fff3fff00003fff55557fff;

	lut_sub lut_8990 ({sk[1920], i_9_, i_7_, i_8_, i_6_, n_n195, n_n464}, x12019x);
	defparam lut_8990.LUT_SIZE = 7;
	defparam lut_8990.mask = 128'h37ff37ff3fff3fff0001001000001110;

	lut_sub lut_8996 ({sk[1921], x24x, x18x, x554x, x23x, x525x, x232x}, x22244x);
	defparam lut_8996.LUT_SIZE = 7;
	defparam lut_8996.mask = 128'h37ff37ff3fff3fffaaa08880aa008800;

	lut_sub lut_9001 ({sk[1922], i_9_, i_7_, i_8_, i_6_, n_n455, n_n535}, n_n727);
	defparam lut_9001.LUT_SIZE = 7;
	defparam lut_9001.mask = 128'h37ff37ff3fff3fff1101101011100010;

	lut_sub lut_9011 ({sk[1923], x16x, x24x, x540x, x496x, x489x, x527x}, x13013x);
	defparam lut_9011.LUT_SIZE = 7;
	defparam lut_9011.mask = 128'h37ff37ff3fff3fff00000fff77777fff;

	lut_sub lut_9016 ({sk[1924], x20x, x495x, x215x, n_n910, x13013x}, x13016x);
	defparam lut_9016.LUT_SIZE = 6;
	defparam lut_9016.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_9021 ({sk[1925], i_9_, i_7_, i_8_, i_6_, n_n536, n_n464}, x13012x);
	defparam lut_9021.LUT_SIZE = 7;
	defparam lut_9021.mask = 128'h37ff37ff3fff3fff0000000101000101;

	lut_sub lut_9026 ({sk[1926], x13x, x550x, x233x, x548x, n_n727, x13012x}, x13017x);
	defparam lut_9026.LUT_SIZE = 7;
	defparam lut_9026.mask = 128'h37ff37ff3fff3fff77ff77ff7fffffff;

	lut_sub lut_9032 ({sk[1927], i_9_, i_7_, i_8_, i_6_, n_n509, n_n260}, x12735x);
	defparam lut_9032.LUT_SIZE = 7;
	defparam lut_9032.mask = 128'h37ff37ff3fff3fff0000000101010010;

	lut_sub lut_9037 ({sk[1928], i_9_, n_n518, x11x, n_n260, n_n522, x484x}, x12734x);
	defparam lut_9037.LUT_SIZE = 7;
	defparam lut_9037.mask = 128'h37ff37ff3fff3fff0055035700550357;

	lut_sub lut_9041 ({sk[1929], x15x, x21x, x484x, x596x, x12735x, x12734x}, n_n696);
	defparam lut_9041.LUT_SIZE = 7;
	defparam lut_9041.mask = 128'h37ff37ff3fff3fff77777f7f77ff7fff;

	lut_sub lut_9046 ({sk[1930], x25x, x20x, x23x, x561x, x479x, x583x}, x12595x);
	defparam lut_9046.LUT_SIZE = 7;
	defparam lut_9046.mask = 128'h37ff37ff3fff3fff000f555f333f777f;

	lut_sub lut_9050 ({sk[1931], x10x, x20x, x547x, x517x, n_n4611, n_n4633}, x22213x);
	defparam lut_9050.LUT_SIZE = 7;
	defparam lut_9050.mask = 128'h37ff37ff3fff3fff8888880080808000;

	lut_sub lut_9055 ({sk[1932], x25x, x539x, x10x, x583x, x12595x, x22213x}, n_n559);
	defparam lut_9055.LUT_SIZE = 7;
	defparam lut_9055.mask = 128'h37ff37ff3fff3fffbbbbbbffbfbfbfff;

	lut_sub lut_9060 ({sk[1933], i_9_, i_7_, i_8_, i_6_, n_n390, n_n473}, x13263x);
	defparam lut_9060.LUT_SIZE = 7;
	defparam lut_9060.mask = 128'h37ff37ff3fff3fff0001001000011000;

	lut_sub lut_9065 ({sk[1934], i_9_, i_1_, i_2_, i_0_, x518x, x491x}, x343x);
	defparam lut_9065.LUT_SIZE = 7;
	defparam lut_9065.mask = 128'h37ff37ff3fff3fff0000000000007000;

	lut_sub lut_9068 ({sk[1935], i_9_, i_7_, i_8_, i_6_, n_n482, n_n455}, x15445x);
	defparam lut_9068.LUT_SIZE = 7;
	defparam lut_9068.mask = 128'h37ff37ff3fff3fff0010000001101000;

	lut_sub lut_9073 ({sk[1936], i_9_, n_n482, x11x, n_n390, x558x}, x431x);
	defparam lut_9073.LUT_SIZE = 6;
	defparam lut_9073.mask = 64'h77ff77ff00031113;

	lut_sub lut_9076 ({sk[1937], i_9_, i_7_, i_8_, i_6_, x514x, x89x}, x15269x);
	defparam lut_9076.LUT_SIZE = 7;
	defparam lut_9076.mask = 128'h37ff37ff3fff3fff5557557555555555;

	lut_sub lut_9080 ({sk[1938], i_9_, i_7_, i_8_, i_6_, x591x, x514x}, x152x);
	defparam lut_9080.LUT_SIZE = 7;
	defparam lut_9080.mask = 128'h37ff37ff3fff3fff3000000500000000;

	lut_sub lut_9083 ({sk[1939], x21x, x12x, x508x, x114x, x533x, n_n5173}, x22256x);
	defparam lut_9083.LUT_SIZE = 7;
	defparam lut_9083.mask = 128'h37ff37ff3fff3fffa0a0a00080808000;

	lut_sub lut_9088 ({sk[1940], x15x, x11x, x12x, x522x, x524x, x533x}, x22274x);
	defparam lut_9088.LUT_SIZE = 7;
	defparam lut_9088.mask = 128'h37ff37ff3fff3fffffc0aa80aa80aa80;

	lut_sub lut_9093 ({sk[1941], x21x, x12x, x514x, x506x, x502x}, x15268x);
	defparam lut_9093.LUT_SIZE = 6;
	defparam lut_9093.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_9097 ({sk[1942], i_9_, n_n526, n_n482, n_n130, x36x}, x15273x);
	defparam lut_9097.LUT_SIZE = 6;
	defparam lut_9097.mask = 64'h77ff77ff55575557;

	lut_sub lut_9101 ({sk[1943], x25x, x12x, x505x, x527x, x528x, x533x}, x22138x);
	defparam lut_9101.LUT_SIZE = 7;
	defparam lut_9101.mask = 128'h37ff37ff3fff3fffffffc000aaaa8000;

	lut_sub lut_9106 ({sk[1944], x10x, x23x, x547x, x594x}, x100x);
	defparam lut_9106.LUT_SIZE = 5;
	defparam lut_9106.mask = 32'h5f5f0357;

	lut_sub lut_9109 ({sk[1945], x21x, x10x, x547x, x517x}, x276x);
	defparam lut_9109.LUT_SIZE = 5;
	defparam lut_9109.mask = 32'h5f5f0537;

	lut_sub lut_9112 ({sk[1946], i_9_, i_7_, i_8_, i_6_, n_n509, n_n195}, x12159x);
	defparam lut_9112.LUT_SIZE = 7;
	defparam lut_9112.mask = 128'h37ff37ff3fff3fff0010001010000010;

	lut_sub lut_9117 ({sk[1947], i_9_, n_n130, x482x, x581x, x414x}, x12327x);
	defparam lut_9117.LUT_SIZE = 6;
	defparam lut_9117.mask = 64'h77ff77ff5555557f;

	lut_sub lut_9121 ({sk[1948], x15x, x24x, x486x, n_n4144, x12327x}, n_n1446);
	defparam lut_9121.LUT_SIZE = 6;
	defparam lut_9121.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_9126 ({sk[1949], i_9_, i_1_, i_2_, i_0_, n_n491, n_n520}, x139x);
	defparam lut_9126.LUT_SIZE = 7;
	defparam lut_9126.mask = 128'h37ff37ff3fff3fff0001000000010000;

	lut_sub lut_9129 ({sk[1950], i_9_, i_1_, i_2_, i_0_, x574x, x139x}, x11640x);
	defparam lut_9129.LUT_SIZE = 7;
	defparam lut_9129.mask = 128'h37ff37ff3fff3fff5555555555575555;

	lut_sub lut_9132 ({sk[1951], x492x, x22x, x10x, x571x, x557x, n_n4607}, x22240x);
	defparam lut_9132.LUT_SIZE = 7;
	defparam lut_9132.mask = 128'h37ff37ff3fff3fffaa88a080aa00a000;

	lut_sub lut_9137 ({sk[1952], i_9_, i_7_, i_8_, i_6_, x507x, x551x}, x11644x);
	defparam lut_9137.LUT_SIZE = 7;
	defparam lut_9137.mask = 128'h37ff37ff3fff3fff0500030000000000;

	lut_sub lut_9140 ({sk[1953], i_9_, i_1_, i_2_, i_0_, x490x, x527x}, x11645x);
	defparam lut_9140.LUT_SIZE = 7;
	defparam lut_9140.mask = 128'h37ff37ff3fff3fff0000000003050000;

	lut_sub lut_9143 ({sk[1954], x22x, x10x, x547x, x535x}, x99x);
	defparam lut_9143.LUT_SIZE = 5;
	defparam lut_9143.mask = 32'h5f5f0537;

	lut_sub lut_9146 ({sk[1955], i_9_, i_1_, i_2_, i_0_, x545x, x506x}, x11651x);
	defparam lut_9146.LUT_SIZE = 7;
	defparam lut_9146.mask = 128'h37ff37ff3fff3fff0000000000030500;

	lut_sub lut_9149 ({sk[1956], x25x, x24x, x479x, x583x, x547x, n_n4584}, x22239x);
	defparam lut_9149.LUT_SIZE = 7;
	defparam lut_9149.mask = 128'h37ff37ff3fff3fffaaaa8080aa008000;

	lut_sub lut_9154 ({sk[1957], x13x, x482x, x581x, x480x}, x13020x);
	defparam lut_9154.LUT_SIZE = 5;
	defparam lut_9154.mask = 32'h5f5f007f;

	lut_sub lut_9158 ({sk[1958], i_9_, i_7_, i_8_, i_6_, n_n455, n_n509}, x13021x);
	defparam lut_9158.LUT_SIZE = 7;
	defparam lut_9158.mask = 128'h37ff37ff3fff3fff0101001001001010;

	lut_sub lut_9165 ({sk[1959], i_9_, i_7_, i_8_, i_6_, x541x, x476x}, x13025x);
	defparam lut_9165.LUT_SIZE = 7;
	defparam lut_9165.mask = 128'h37ff37ff3fff3fff0050530300000000;

	lut_sub lut_9170 ({sk[1960], i_9_, i_7_, i_8_, i_6_, n_n260, n_n535}, n_n698);
	defparam lut_9170.LUT_SIZE = 7;
	defparam lut_9170.mask = 128'h37ff37ff3fff3fff1010101010111010;

	lut_sub lut_9180 ({sk[1961], x11x, x17x, x596x, x559x}, x52x);
	defparam lut_9180.LUT_SIZE = 5;
	defparam lut_9180.mask = 32'h5f5f0537;

	lut_sub lut_9183 ({sk[1962], x15x, x24x, x17x, x552x, x550x, x596x}, x12748x);
	defparam lut_9183.LUT_SIZE = 7;
	defparam lut_9183.mask = 128'h37ff37ff3fff3fff00335f7f55775f7f;

	lut_sub lut_9188 ({sk[1963], x22x, x23x, x530x, n_n698, x52x, x12748x}, x12753x);
	defparam lut_9188.LUT_SIZE = 7;
	defparam lut_9188.mask = 128'h37ff37ff3fff3fff7f7f7fff7fff7fff;

	lut_sub lut_9194 ({sk[1964], i_9_, i_7_, i_8_, i_6_, n_n390, n_n491}, x12600x);
	defparam lut_9194.LUT_SIZE = 7;
	defparam lut_9194.mask = 128'h37ff37ff3fff3fff1000101010000000;

	lut_sub lut_9199 ({sk[1965], i_9_, n_n482, n_n390, n_n532, x20x, x571x}, x12599x);
	defparam lut_9199.LUT_SIZE = 7;
	defparam lut_9199.mask = 128'h37ff37ff3fff3fff1111111f1111111f;

	lut_sub lut_9203 ({sk[1966], x10x, x24x, x571x, x587x, x12600x, x12599x}, n_n558);
	defparam lut_9203.LUT_SIZE = 7;
	defparam lut_9203.mask = 128'h37ff37ff3fff3fff777777ff7f7f7fff;

	lut_sub lut_9208 ({sk[1967], x22x, x11x, x12x, x554x, x598x, x593x}, x12656x);
	defparam lut_9208.LUT_SIZE = 7;
	defparam lut_9208.mask = 128'h37ff37ff3fff3fff005533773f7f3f7f;

	lut_sub lut_9213 ({sk[1968], x16x, x521x, x21x, x501x}, x53x);
	defparam lut_9213.LUT_SIZE = 5;
	defparam lut_9213.mask = 32'h5f5f111f;

	lut_sub lut_9216 ({sk[1969], i_9_, n_n536, n_n532, n_n509, x156x}, x13509x);
	defparam lut_9216.LUT_SIZE = 6;
	defparam lut_9216.mask = 64'h77ff77ff55575557;

	lut_sub lut_9220 ({sk[1970], i_9_, i_7_, i_8_, i_6_, n_n536, n_n535}, x363x);
	defparam lut_9220.LUT_SIZE = 7;
	defparam lut_9220.mask = 128'h37ff37ff3fff3fff0000101001001000;

	lut_sub lut_9225 ({sk[1971], x15x, x16x, x501x, x559x}, x443x);
	defparam lut_9225.LUT_SIZE = 5;
	defparam lut_9225.mask = 32'h5f5f0537;

	lut_sub lut_9228 ({sk[1972], x25x, x22x, x501x, x473x, n_n4344, x53x}, x22191x);
	defparam lut_9228.LUT_SIZE = 7;
	defparam lut_9228.mask = 128'h37ff37ff3fff3fff8888880080808000;

	lut_sub lut_9233 ({sk[1973], x24x, x12x, x573x, x578x}, x407x);
	defparam lut_9233.LUT_SIZE = 5;
	defparam lut_9233.mask = 32'h5f5f0357;

	lut_sub lut_9236 ({sk[1974], x509x, x24x, x17x, x512x}, x42x);
	defparam lut_9236.LUT_SIZE = 5;
	defparam lut_9236.mask = 32'h5f5f0537;

	lut_sub lut_9239 ({sk[1975], i_9_, i_7_, i_8_, i_6_, x497x}, x106x);
	defparam lut_9239.LUT_SIZE = 6;
	defparam lut_9239.mask = 64'h77ff77ff44000000;

	lut_sub lut_9242 ({sk[1976], x11x, x18x, x527x, x528x, x532x}, x14005x);
	defparam lut_9242.LUT_SIZE = 6;
	defparam lut_9242.mask = 64'h77ff77ff003f557f;

	lut_sub lut_9246 ({sk[1977], i_9_, i_7_, i_8_, i_6_, x554x, x532x}, x22171x);
	defparam lut_9246.LUT_SIZE = 7;
	defparam lut_9246.mask = 128'h37ff37ff3fff3fffffaafcfcffffffff;

	lut_sub lut_9256 ({sk[1978], i_9_, i_7_, i_8_, i_6_, n_n260, n_n535}, x15686x);
	defparam lut_9256.LUT_SIZE = 7;
	defparam lut_9256.mask = 128'h37ff37ff3fff3fff0001010001000001;

	lut_sub lut_9261 ({sk[1979], x521x, x21x, x17x, x596x}, x375x);
	defparam lut_9261.LUT_SIZE = 5;
	defparam lut_9261.mask = 32'h5f5f0537;

	lut_sub lut_9264 ({sk[1980], i_9_, i_7_, i_8_, i_6_, n_n518, n_n260}, x15693x);
	defparam lut_9264.LUT_SIZE = 7;
	defparam lut_9264.mask = 128'h37ff37ff3fff3fff1010001000000100;

	lut_sub lut_9269 ({sk[1981], x17x, x20x, x548x, x530x}, x15685x);
	defparam lut_9269.LUT_SIZE = 5;
	defparam lut_9269.mask = 32'h5f5f0537;

	lut_sub lut_9272 ({sk[1982], i_9_, n_n518, n_n260, n_n530, x52x}, x15691x);
	defparam lut_9272.LUT_SIZE = 6;
	defparam lut_9272.mask = 64'h77ff77ff55575557;

	lut_sub lut_9276 ({sk[1983], i_9_, n_n534, n_n509, n_n260, x375x}, x15692x);
	defparam lut_9276.LUT_SIZE = 6;
	defparam lut_9276.mask = 64'h77ff77ff55575557;

	lut_sub lut_9280 ({sk[1984], x25x, x10x, x24x, x583x, x593x}, n_n2401);
	defparam lut_9280.LUT_SIZE = 6;
	defparam lut_9280.mask = 64'h77ff77ff03573377;

	lut_sub lut_9284 ({sk[1985], i_9_, i_7_, i_8_, i_6_, n_n455, n_n473}, n_n1491);
	defparam lut_9284.LUT_SIZE = 7;
	defparam lut_9284.mask = 128'h37ff37ff3fff3fff0111101001110100;

	lut_sub lut_9294 ({sk[1986], i_9_, i_7_, i_8_, i_6_, n_n390, n_n473}, x12420x);
	defparam lut_9294.LUT_SIZE = 7;
	defparam lut_9294.mask = 128'h37ff37ff3fff3fff1000001011000000;

	lut_sub lut_9299 ({sk[1987], i_9_, i_7_, i_8_, i_6_, n_n536, n_n500}, x12445x);
	defparam lut_9299.LUT_SIZE = 7;
	defparam lut_9299.mask = 128'h37ff37ff3fff3fff0110100000000010;

	lut_sub lut_9304 ({sk[1988], x492x, x16x, x21x, x570x, x499x}, n_n1693);
	defparam lut_9304.LUT_SIZE = 6;
	defparam lut_9304.mask = 64'h77ff77ff053705ff;

	lut_sub lut_9308 ({sk[1989], i_9_, i_7_, i_8_, i_6_, n_n536, n_n491}, x12453x);
	defparam lut_9308.LUT_SIZE = 7;
	defparam lut_9308.mask = 128'h37ff37ff3fff3fff0000101010101010;

	lut_sub lut_9315 ({sk[1990], x16x, x24x, x563x, x498x, x480x, x562x}, x22283x);
	defparam lut_9315.LUT_SIZE = 7;
	defparam lut_9315.mask = 128'h37ff37ff3fff3ffffffff0f088008000;

	lut_sub lut_9320 ({sk[1991], x15x, x16x, x498x, x560x}, x12443x);
	defparam lut_9320.LUT_SIZE = 5;
	defparam lut_9320.mask = 32'h5f5f0537;

	lut_sub lut_9323 ({sk[1992], x16x, x24x, x499x, x518x, x573x}, x12444x);
	defparam lut_9323.LUT_SIZE = 6;
	defparam lut_9323.mask = 64'h77ff77ff000f777f;

	lut_sub lut_9327 ({sk[1993], i_9_, i_7_, i_8_, i_6_, n_n536, n_n509}, x12451x);
	defparam lut_9327.LUT_SIZE = 7;
	defparam lut_9327.mask = 128'h37ff37ff3fff3fff0010100010100000;

	lut_sub lut_9332 ({sk[1994], x538x, x21x, x14x, x588x, x20x, x23x}, x22226x);
	defparam lut_9332.LUT_SIZE = 7;
	defparam lut_9332.mask = 128'h37ff37ff3fff3ffff8f8f0f0f800f000;

	lut_sub lut_9337 ({sk[1995], x11x, x511x, x179x, x158x, x22226x}, n_n1471);
	defparam lut_9337.LUT_SIZE = 6;
	defparam lut_9337.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_9342 ({sk[1996], i_9_, i_7_, i_8_, i_6_, n_n482, n_n325}, x12208x);
	defparam lut_9342.LUT_SIZE = 7;
	defparam lut_9342.mask = 128'h37ff37ff3fff3fff0001000101000001;

	lut_sub lut_9347 ({sk[1997], x24x, x14x, x588x, x23x, x584x, x575x}, x12207x);
	defparam lut_9347.LUT_SIZE = 7;
	defparam lut_9347.mask = 128'h37ff37ff3fff3fff0505373705ff37ff;

	lut_sub lut_9351 ({sk[1998], x11x, x14x, x588x, x586x, x12208x, x12207x}, n_n1472);
	defparam lut_9351.LUT_SIZE = 7;
	defparam lut_9351.mask = 128'h37ff37ff3fff3fff77777f7f77ff7fff;

	lut_sub lut_9356 ({sk[1999], i_9_, i_7_, i_8_, i_6_, n_n130, n_n464}, n_n1439);
	defparam lut_9356.LUT_SIZE = 7;
	defparam lut_9356.mask = 128'h37ff37ff3fff3fff0101111101010001;

	lut_sub lut_9366 ({sk[2000], x19x, x22x, x11x, x517x, x555x}, n_n763);
	defparam lut_9366.LUT_SIZE = 6;
	defparam lut_9366.mask = 64'h77ff77ff05553777;

	lut_sub lut_9370 ({sk[2001], i_9_, i_7_, i_8_, i_6_, n_n535, n_n65}, x12280x);
	defparam lut_9370.LUT_SIZE = 7;
	defparam lut_9370.mask = 128'h37ff37ff3fff3fff0101001100001100;

	lut_sub lut_9377 ({sk[2002], x19x, x521x, x21x, x555x, n_n1530, x12280x}, x12282x);
	defparam lut_9377.LUT_SIZE = 7;
	defparam lut_9377.mask = 128'h37ff37ff3fff3fff777f777f777fffff;

	lut_sub lut_9382 ({sk[2003], x19x, x22x, x490x, x599x, x559x, n_n5223}, x22233x);
	defparam lut_9382.LUT_SIZE = 7;
	defparam lut_9382.mask = 128'h37ff37ff3fff3fffaaaaa0a088008000;

	lut_sub lut_9387 ({sk[2004], x20x, x533x, n_n1439, x450x, x22233x}, x12283x);
	defparam lut_9387.LUT_SIZE = 6;
	defparam lut_9387.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_9392 ({sk[2005], i_9_, x22x, n_n473, n_n532, n_n130, x503x}, x12291x);
	defparam lut_9392.LUT_SIZE = 7;
	defparam lut_9392.mask = 128'h37ff37ff3fff3fff0003003311131133;

	lut_sub lut_9397 ({sk[2006], i_9_, n_n482, n_n522, n_n130, x514x, x506x}, x12292x);
	defparam lut_9397.LUT_SIZE = 7;
	defparam lut_9397.mask = 128'h37ff37ff3fff3fff0033003f0505050f;

	lut_sub lut_9402 ({sk[2007], i_9_, x25x, n_n524, n_n473, n_n130, x591x}, x12293x);
	defparam lut_9402.LUT_SIZE = 7;
	defparam lut_9402.mask = 128'h37ff37ff3fff3fff0057035700030303;

	lut_sub lut_9407 ({sk[2008], x510x, x12x, x508x, n_n5181, x505x, x44x}, x22257x);
	defparam lut_9407.LUT_SIZE = 7;
	defparam lut_9407.mask = 128'h37ff37ff3fff3fffa0a08000a0a00000;

	lut_sub lut_9410 ({sk[2009], n_n1442, x12291x, x12292x, x12293x, x22257x}, n_n1406);
	defparam lut_9410.LUT_SIZE = 6;
	defparam lut_9410.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_9416 ({sk[2010], i_9_, i_7_, i_8_, i_6_, x486x}, x286x);
	defparam lut_9416.LUT_SIZE = 6;
	defparam lut_9416.mask = 64'h77ff77ff04400000;

	lut_sub lut_9419 ({sk[2011], x12x, x475x, x563x, x286x, x12299x, x12300x}, x12303x);
	defparam lut_9419.LUT_SIZE = 7;
	defparam lut_9419.mask = 128'h37ff37ff3fff3fff7f7f7f7f7fffffff;

	lut_sub lut_9425 ({sk[2012], x12x, x574x, n_n1443, x125x, x12265x, x12263x}, x12304x);
	defparam lut_9425.LUT_SIZE = 7;
	defparam lut_9425.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_9431 ({sk[2013], x16x, x500x, x23x, x488x, x524x, x493x}, x12136x);
	defparam lut_9431.LUT_SIZE = 7;
	defparam lut_9431.mask = 128'h37ff37ff3fff3fff000000ff7f7f7fff;

	lut_sub lut_9436 ({sk[2014], i_9_, x25x, n_n536, n_n528, n_n509, x494x}, x12141x);
	defparam lut_9436.LUT_SIZE = 7;
	defparam lut_9436.mask = 128'h37ff37ff3fff3fff0003003300570077;

	lut_sub lut_9441 ({sk[2015], x15x, x22x, x14x, x588x, x586x, x511x}, x11675x);
	defparam lut_9441.LUT_SIZE = 7;
	defparam lut_9441.mask = 128'h37ff37ff3fff3fff003355775f7f5f7f;

	lut_sub lut_9446 ({sk[2016], i_9_, i_7_, i_8_, i_6_, x530x, x575x}, x22266x);
	defparam lut_9446.LUT_SIZE = 7;
	defparam lut_9446.mask = 128'h37ff37ff3fff3fffcfacffcfffffffff;

	lut_sub lut_9456 ({sk[2017], i_9_, x482x, x581x, n_n65, x318x}, x12872x);
	defparam lut_9456.LUT_SIZE = 6;
	defparam lut_9456.mask = 64'h77ff77ff55555777;

	lut_sub lut_9460 ({sk[2018], x19x, x23x, x594x, x546x, x555x}, n_n761);
	defparam lut_9460.LUT_SIZE = 6;
	defparam lut_9460.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_9464 ({sk[2019], x15x, x19x, x490x, x550x, x599x, x223x}, x22310x);
	defparam lut_9464.LUT_SIZE = 7;
	defparam lut_9464.mask = 128'h37ff37ff3fff3fffaaaaa00088888000;

	lut_sub lut_9469 ({sk[2020], n_n763, n_n761, x22310x}, x12881x);
	defparam lut_9469.LUT_SIZE = 4;
	defparam lut_9469.mask = 16'h0fbf;

	lut_sub lut_9473 ({sk[2021], x25x, x19x, x521x, x481x, x487x}, x12871x);
	defparam lut_9473.LUT_SIZE = 6;
	defparam lut_9473.mask = 64'h77ff77ff003f557f;

	lut_sub lut_9477 ({sk[2022], x19x, x24x, x480x, x487x, x593x, x182x}, x22205x);
	defparam lut_9477.LUT_SIZE = 7;
	defparam lut_9477.mask = 128'h37ff37ff3fff3fffaaaaa0a088008000;

	lut_sub lut_9482 ({sk[2023], x383x, x183x, x12872x, x12871x, x22205x}, x12882x);
	defparam lut_9482.LUT_SIZE = 6;
	defparam lut_9482.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_9488 ({sk[2024], i_9_, i_7_, i_8_, i_6_, n_n482, n_n130}, x12888x);
	defparam lut_9488.LUT_SIZE = 7;
	defparam lut_9488.mask = 128'h37ff37ff3fff3fff0100000100000101;

	lut_sub lut_9493 ({sk[2025], i_9_, i_7_, i_8_, i_6_, n_n491, n_n130}, x12893x);
	defparam lut_9493.LUT_SIZE = 7;
	defparam lut_9493.mask = 128'h37ff37ff3fff3fff0001010001000100;

	lut_sub lut_9498 ({sk[2026], x22x, x24x, x23x, x591x, x578x, x287x}, x22204x);
	defparam lut_9498.LUT_SIZE = 7;
	defparam lut_9498.mask = 128'h37ff37ff3fff3fffaa88a080a080a080;

	lut_sub lut_9503 ({sk[2027], x12x, x574x, x126x, x12888x, x12893x, x22204x}, x12898x);
	defparam lut_9503.LUT_SIZE = 7;
	defparam lut_9503.mask = 128'h37ff37ff3fff3fffbfffbfffbfffffff;

	lut_sub lut_9509 ({sk[2028], x22x, x12x, x486x, x556x}, x12645x);
	defparam lut_9509.LUT_SIZE = 5;
	defparam lut_9509.mask = 32'h5f5f0537;

	lut_sub lut_9512 ({sk[2029], i_9_, i_7_, i_8_, i_6_, x486x, x578x}, x12646x);
	defparam lut_9512.LUT_SIZE = 7;
	defparam lut_9512.mask = 128'h37ff37ff3fff3fff0500700000000000;

	lut_sub lut_9516 ({sk[2030], x15x, x570x, x12x, x591x, x486x}, x22300x);
	defparam lut_9516.LUT_SIZE = 6;
	defparam lut_9516.mask = 64'h77ff77fffff08880;

	lut_sub lut_9521 ({sk[2031], i_9_, i_7_, i_8_, i_6_, n_n536, n_n473}, n_n4097);
	defparam lut_9521.LUT_SIZE = 7;
	defparam lut_9521.mask = 128'h37ff37ff3fff3fff0100111101011010;

	lut_sub lut_9531 ({sk[2032], i_9_, i_1_, i_2_, i_0_, x525x}, n_n4694);
	defparam lut_9531.LUT_SIZE = 6;
	defparam lut_9531.mask = 64'h77ff77ff00000100;

	lut_sub lut_9533 ({sk[2033], i_9_, i_1_, i_2_, i_0_, x548x}, n_n4700);
	defparam lut_9533.LUT_SIZE = 6;
	defparam lut_9533.mask = 64'h77ff77ff00001000;

	lut_sub lut_9535 ({sk[2034], x14x, x20x, x546x, x551x}, x30x);
	defparam lut_9535.LUT_SIZE = 5;
	defparam lut_9535.mask = 32'h5f5f0537;

	lut_sub lut_9538 ({sk[2035], i_9_, i_7_, i_8_, i_6_, n_n260, n_n535}, x303x);
	defparam lut_9538.LUT_SIZE = 7;
	defparam lut_9538.mask = 128'h37ff37ff3fff3fff0000001000001000;

	lut_sub lut_9541 ({sk[2036], x21x, x539x, x12x, x482x, x486x, x536x}, x13579x);
	defparam lut_9541.LUT_SIZE = 7;
	defparam lut_9541.mask = 128'h37ff37ff3fff3fff005f00ff337f33ff;

	lut_sub lut_9546 ({sk[2037], x19x, x570x, x557x, x494x, x562x}, x13586x);
	defparam lut_9546.LUT_SIZE = 6;
	defparam lut_9546.mask = 64'h77ff77ff00007fff;

	lut_sub lut_9551 ({sk[2038], x25x, x15x, x592x, x538x, x19x, x424x}, x22199x);
	defparam lut_9551.LUT_SIZE = 7;
	defparam lut_9551.mask = 128'h37ff37ff3fff3fffa8a8a800a800a800;

	lut_sub lut_9556 ({sk[2039], x515x, x19x, x11x, x24x, x503x, x534x}, x22313x);
	defparam lut_9556.LUT_SIZE = 7;
	defparam lut_9556.mask = 128'h37ff37ff3fff3ffffafac8c8fa00c800;

	lut_sub lut_9565 ({sk[2040], x21x, x18x, x553x, x559x}, x13596x);
	defparam lut_9565.LUT_SIZE = 5;
	defparam lut_9565.mask = 32'h5f5f0537;

	lut_sub lut_9568 ({sk[2041], i_9_, x22x, n_n528, n_n535, n_n195, x512x}, x13598x);
	defparam lut_9568.LUT_SIZE = 7;
	defparam lut_9568.mask = 128'h37ff37ff3fff3fff0055035700030303;

	lut_sub lut_9572 ({sk[2042], x22x, x24x, x510x, x17x, x485x, x567x}, x22314x);
	defparam lut_9572.LUT_SIZE = 7;
	defparam lut_9572.mask = 128'h37ff37ff3fff3ffffff0ccc0aaa08880;

	lut_sub lut_9581 ({sk[2043], x15x, x18x, x587x, x577x, x584x}, x13605x);
	defparam lut_9581.LUT_SIZE = 6;
	defparam lut_9581.mask = 64'h77ff77ff005f337f;

	lut_sub lut_9585 ({sk[2044], x18x, x23x, x572x, x590x, x503x, x567x}, x22198x);
	defparam lut_9585.LUT_SIZE = 7;
	defparam lut_9585.mask = 128'h37ff37ff3fff3fffffffa0a0cc008000;

	lut_sub lut_9590 ({sk[2045], x19x, x11x, x24x, x599x, x546x, x593x}, x22312x);
	defparam lut_9590.LUT_SIZE = 7;
	defparam lut_9590.mask = 128'h37ff37ff3fff3ffffff0f0f088808080;

	lut_sub lut_9595 ({sk[2046], i_9_, x25x, n_n509, n_n520, n_n130, x568x}, n_n3051);
	defparam lut_9595.LUT_SIZE = 7;
	defparam lut_9595.mask = 128'h37ff37ff3fff3fff0003555700035557;

	lut_sub lut_9599 ({sk[2047], x16x, x570x, x20x, x499x}, x285x);
	defparam lut_9599.LUT_SIZE = 5;
	defparam lut_9599.mask = 32'h5f5f111f;

	lut_sub lut_9602 ({sk[2048], i_9_, i_7_, i_8_, i_6_, n_n536, n_n491}, x15507x);
	defparam lut_9602.LUT_SIZE = 7;
	defparam lut_9602.mask = 128'h37ff37ff3fff3fff0110001010000000;

	lut_sub lut_9607 ({sk[2049], i_9_, i_7_, i_8_, i_6_, n_n455, n_n535}, n_n3003);
	defparam lut_9607.LUT_SIZE = 7;
	defparam lut_9607.mask = 128'h37ff37ff3fff3fff0101011001010111;

	lut_sub lut_9617 ({sk[2050], x14x, x23x, x529x, x511x}, x440x);
	defparam lut_9617.LUT_SIZE = 5;
	defparam lut_9617.mask = 32'h5f5f0537;

	lut_sub lut_9620 ({sk[2051], i_9_, i_7_, i_8_, i_6_, n_n536, n_n473}, x12459x);
	defparam lut_9620.LUT_SIZE = 7;
	defparam lut_9620.mask = 128'h37ff37ff3fff3fff0000110000011000;

	lut_sub lut_9625 ({sk[2052], i_9_, n_n536, n_n482, n_n528, x587x, n_n4428}, x12466x);
	defparam lut_9625.LUT_SIZE = 7;
	defparam lut_9625.mask = 128'h37ff37ff3fff3fff5555555f5555777f;

	lut_sub lut_9630 ({sk[2053], i_9_, i_7_, i_8_, i_6_, x500x, x495x}, x12457x);
	defparam lut_9630.LUT_SIZE = 7;
	defparam lut_9630.mask = 128'h37ff37ff3fff3fff0500300000000000;

	lut_sub lut_9633 ({sk[2054], x16x, x500x, x510x, x20x, x580x}, x12458x);
	defparam lut_9633.LUT_SIZE = 6;
	defparam lut_9633.mask = 64'h77ff77ff00335f7f;

	lut_sub lut_9637 ({sk[2055], i_9_, n_n536, x500x, n_n534, x586x, n_n464}, x12464x);
	defparam lut_9637.LUT_SIZE = 7;
	defparam lut_9637.mask = 128'h37ff37ff3fff3fff000f050f00003737;

	lut_sub lut_9642 ({sk[2056], i_9_, i_7_, i_8_, i_6_, n_n536, n_n482}, x12465x);
	defparam lut_9642.LUT_SIZE = 7;
	defparam lut_9642.mask = 128'h37ff37ff3fff3fff0000011000011000;

	lut_sub lut_9647 ({sk[2057], i_9_, i_7_, i_8_, i_6_, n_n500, n_n65}, x12357x);
	defparam lut_9647.LUT_SIZE = 7;
	defparam lut_9647.mask = 128'h37ff37ff3fff3fff0010000001110000;

	lut_sub lut_9652 ({sk[2058], i_9_, n_n526, n_n500, n_n65, n_n1521, x12357x}, x12359x);
	defparam lut_9652.LUT_SIZE = 7;
	defparam lut_9652.mask = 128'h37ff37ff3fff3fff7777777f7777777f;

	lut_sub lut_9657 ({sk[2059], i_9_, i_7_, i_8_, i_6_, n_n195, n_n464}, x12324x);
	defparam lut_9657.LUT_SIZE = 7;
	defparam lut_9657.mask = 128'h37ff37ff3fff3fff0101101001111010;

	lut_sub lut_9667 ({sk[2060], i_9_, i_7_, i_8_, i_6_, x513x, x532x}, x12308x);
	defparam lut_9667.LUT_SIZE = 7;
	defparam lut_9667.mask = 128'h37ff37ff3fff3fff0030050000000000;

	lut_sub lut_9670 ({sk[2061], i_9_, i_7_, i_8_, i_6_, x590x, x513x}, x12313x);
	defparam lut_9670.LUT_SIZE = 7;
	defparam lut_9670.mask = 128'h37ff37ff3fff3fff0300000500000000;

	lut_sub lut_9673 ({sk[2062], x18x, x508x, x580x, x502x, x120x, x493x}, x22232x);
	defparam lut_9673.LUT_SIZE = 7;
	defparam lut_9673.mask = 128'h37ff37ff3fff3fffcccccccc80000000;

	lut_sub lut_9676 ({sk[2063], x12310x, x12315x, x12308x, x12313x, x22232x}, x12325x);
	defparam lut_9676.LUT_SIZE = 6;
	defparam lut_9676.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_9682 ({sk[2064], x24x, x18x, x554x, x525x}, x12331x);
	defparam lut_9682.LUT_SIZE = 5;
	defparam lut_9682.mask = 32'h5f5f0537;

	lut_sub lut_9685 ({sk[2065], x15x, x12x, x554x, x549x, x548x, n_n5079}, x22231x);
	defparam lut_9685.LUT_SIZE = 7;
	defparam lut_9685.mask = 128'h37ff37ff3fff3fffaaaa8080aa008000;

	lut_sub lut_9690 ({sk[2066], x20x, x532x, x143x, x12331x, x22231x}, n_n1448);
	defparam lut_9690.LUT_SIZE = 6;
	defparam lut_9690.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_9695 ({sk[2067], x11x, x12x, x598x, x585x}, x12336x);
	defparam lut_9695.LUT_SIZE = 5;
	defparam lut_9695.mask = 32'h5f5f0537;

	lut_sub lut_9698 ({sk[2068], i_9_, i_7_, i_8_, i_6_, x554x, x598x}, x12338x);
	defparam lut_9698.LUT_SIZE = 7;
	defparam lut_9698.mask = 128'h37ff37ff3fff3fff0035305000000000;

	lut_sub lut_9703 ({sk[2069], x12x, x546x, x34x, x12336x, x12338x}, x12340x);
	defparam lut_9703.LUT_SIZE = 6;
	defparam lut_9703.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_9708 ({sk[2070], i_9_, i_7_, i_8_, i_6_, n_n491, n_n65}, n_n664);
	defparam lut_9708.LUT_SIZE = 7;
	defparam lut_9708.mask = 128'h37ff37ff3fff3fff0111110101000110;

	lut_sub lut_9718 ({sk[2071], i_9_, n_n522, n_n500, n_n65, x446x}, x12956x);
	defparam lut_9718.LUT_SIZE = 6;
	defparam lut_9718.mask = 64'h77ff77ff55575557;

	lut_sub lut_9722 ({sk[2072], i_9_, x21x, n_n526, n_n500, n_n65, x487x}, x12957x);
	defparam lut_9722.LUT_SIZE = 7;
	defparam lut_9722.mask = 128'h37ff37ff3fff3fff0003575700035757;

	lut_sub lut_9727 ({sk[2073], i_9_, n_n509, n_n522, x478x, x562x, n_n65}, x12958x);
	defparam lut_9727.LUT_SIZE = 7;
	defparam lut_9727.mask = 128'h37ff37ff3fff3fff0000005515151555;

	lut_sub lut_9732 ({sk[2074], n_n1521, n_n3385, n_n664, x12956x, x12957x, x12958x}, n_n634);
	defparam lut_9732.LUT_SIZE = 7;
	defparam lut_9732.mask = 128'h37ff37ff3fff3fff7fffffffffffffff;

	lut_sub lut_9739 ({sk[2075], x18x, x20x, x502x, x513x, x527x, x528x}, x22307x);
	defparam lut_9739.LUT_SIZE = 7;
	defparam lut_9739.mask = 128'h37ff37ff3fff3ffffffff0f088008000;

	lut_sub lut_9744 ({sk[2076], x22x, x21x, x513x, x532x, n_n789, x22307x}, n_n680);
	defparam lut_9744.LUT_SIZE = 7;
	defparam lut_9744.mask = 128'h37ff37ff3fff3fffbbbbbbffbfbfbfff;

	lut_sub lut_9749 ({sk[2077], i_9_, i_7_, i_8_, i_6_, n_n473, n_n195}, x12907x);
	defparam lut_9749.LUT_SIZE = 7;
	defparam lut_9749.mask = 128'h37ff37ff3fff3fff0100000101000100;

	lut_sub lut_9754 ({sk[2078], x15x, x24x, x18x, x508x, x513x}, x12906x);
	defparam lut_9754.LUT_SIZE = 6;
	defparam lut_9754.mask = 64'h77ff77ff03575757;

	lut_sub lut_9758 ({sk[2079], x22x, x23x, x590x, x513x, x12907x, x12906x}, n_n681);
	defparam lut_9758.LUT_SIZE = 7;
	defparam lut_9758.mask = 128'h37ff37ff3fff3fff777777ff7f7f7fff;

	lut_sub lut_9763 ({sk[2080], x25x, x15x, x12x, x554x, x549x, n_n5074}, x22208x);
	defparam lut_9763.LUT_SIZE = 7;
	defparam lut_9763.mask = 128'h37ff37ff3fff3fffaa88a080a080a080;

	lut_sub lut_9768 ({sk[2081], x24x, x12x, x554x, x550x, x209x}, x22260x);
	defparam lut_9768.LUT_SIZE = 6;
	defparam lut_9768.mask = 64'h77ff77ffaa88a080;

	lut_sub lut_9773 ({sk[2082], x23x, x532x, x22208x, x22260x}, x12915x);
	defparam lut_9773.LUT_SIZE = 5;
	defparam lut_9773.mask = 32'h5f5feeef;

	lut_sub lut_9777 ({sk[2083], x25x, x12x, x472x, x475x, x478x, x568x}, x12921x);
	defparam lut_9777.LUT_SIZE = 7;
	defparam lut_9777.mask = 128'h37ff37ff3fff3fff00003fff55557fff;

	lut_sub lut_9782 ({sk[2084], x521x, x12x, x559x, x11914x, x11915x, n_n783}, x12929x);
	defparam lut_9782.LUT_SIZE = 7;
	defparam lut_9782.mask = 128'h37ff37ff3fff3fff7f7f7fff7f7fffff;

	lut_sub lut_9788 ({sk[2085], i_9_, i_7_, i_8_, i_6_, n_n518, n_n130}, x12925x);
	defparam lut_9788.LUT_SIZE = 7;
	defparam lut_9788.mask = 128'h37ff37ff3fff3fff0001110000100000;

	lut_sub lut_9793 ({sk[2086], i_9_, n_n528, n_n535, n_n130, x482x, x143x}, x12926x);
	defparam lut_9793.LUT_SIZE = 7;
	defparam lut_9793.mask = 128'h37ff37ff3fff3fff555555555757575f;

	lut_sub lut_9797 ({sk[2087], x474x, x12x, x23x, x564x, x486x, x414x}, x22207x);
	defparam lut_9797.LUT_SIZE = 7;
	defparam lut_9797.mask = 128'h37ff37ff3fff3fffaa88a080aa880000;

	lut_sub lut_9802 ({sk[2088], x12921x, x12925x, x12926x, x22207x}, x12930x);
	defparam lut_9802.LUT_SIZE = 5;
	defparam lut_9802.mask = 32'h5f5fbfff;

	lut_sub lut_9807 ({sk[2089], x11x, x567x, n_n5016, n_n3427, x297x, x394x}, n_n684);
	defparam lut_9807.LUT_SIZE = 7;
	defparam lut_9807.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_9813 ({sk[2090], i_9_, i_7_, i_8_, i_6_, n_n491, n_n195}, x12938x);
	defparam lut_9813.LUT_SIZE = 7;
	defparam lut_9813.mask = 128'h37ff37ff3fff3fff0000001000101010;

	lut_sub lut_9818 ({sk[2091], x11x, x20x, x23x, x577x, x253x, x12938x}, n_n683);
	defparam lut_9818.LUT_SIZE = 7;
	defparam lut_9818.mask = 128'h37ff37ff3fff3fff777f7f7f7f7f7f7f;

	lut_sub lut_9824 ({sk[2092], n_n680, n_n681, x12915x, x12929x, x12930x}, x12948x);
	defparam lut_9824.LUT_SIZE = 6;
	defparam lut_9824.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_9830 ({sk[2093], i_9_, i_7_, i_8_, i_6_, n_n536, n_n491}, x13532x);
	defparam lut_9830.LUT_SIZE = 7;
	defparam lut_9830.mask = 128'h37ff37ff3fff3fff0100101000001000;

	lut_sub lut_9835 ({sk[2094], i_9_, i_7_, i_8_, i_6_, n_n536, n_n482}, x13539x);
	defparam lut_9835.LUT_SIZE = 7;
	defparam lut_9835.mask = 128'h37ff37ff3fff3fff0011101011110010;

	lut_sub lut_9845 ({sk[2095], x16x, x20x, x499x, x537x}, x13530x);
	defparam lut_9845.LUT_SIZE = 5;
	defparam lut_9845.mask = 32'h5f5f0357;

	lut_sub lut_9848 ({sk[2096], x25x, x16x, x500x, x570x, x586x}, x13531x);
	defparam lut_9848.LUT_SIZE = 6;
	defparam lut_9848.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_9852 ({sk[2097], x515x, x15x, x592x, x22x, x21x, n_n5306}, x22172x);
	defparam lut_9852.LUT_SIZE = 7;
	defparam lut_9852.mask = 128'h37ff37ff3fff3fffaa80aa80aa800000;

	lut_sub lut_9857 ({sk[2098], x592x, x538x, x19x, x510x, x20x, x520x}, x22272x);
	defparam lut_9857.LUT_SIZE = 7;
	defparam lut_9857.mask = 128'h37ff37ff3fff3fffffa0ff00cc80cc00;

	lut_sub lut_9862 ({sk[2099], i_9_, i_7_, i_8_, i_6_, n_n509, n_n65}, x13954x);
	defparam lut_9862.LUT_SIZE = 7;
	defparam lut_9862.mask = 128'h37ff37ff3fff3fff0010101000000010;

	lut_sub lut_9867 ({sk[2100], i_9_, i_7_, i_8_, i_6_, n_n455, n_n535}, x12475x);
	defparam lut_9867.LUT_SIZE = 7;
	defparam lut_9867.mask = 128'h37ff37ff3fff3fff0001000001010001;

	lut_sub lut_9872 ({sk[2101], i_9_, i_7_, i_8_, i_6_, n_n518, n_n455}, x12483x);
	defparam lut_9872.LUT_SIZE = 7;
	defparam lut_9872.mask = 128'h37ff37ff3fff3fff0001010101010001;

	lut_sub lut_9879 ({sk[2102], x21x, x13x, x540x, x535x, n_n3162, x12483x}, x12485x);
	defparam lut_9879.LUT_SIZE = 7;
	defparam lut_9879.mask = 128'h37ff37ff3fff3fff77777f7f77ff7fff;

	lut_sub lut_9884 ({sk[2103], x22x, x13x, x539x, x544x, x11x}, x12480x);
	defparam lut_9884.LUT_SIZE = 6;
	defparam lut_9884.mask = 64'h77ff77ff111f333f;

	lut_sub lut_9888 ({sk[2104], i_9_, n_n455, n_n535, x490x, x20x, x128x}, x12481x);
	defparam lut_9888.LUT_SIZE = 7;
	defparam lut_9888.mask = 128'h37ff37ff3fff3fff5555557755555f7f;

	lut_sub lut_9892 ({sk[2105], x21x, x11x, x20x, x540x, x496x, x421x}, x22230x);
	defparam lut_9892.LUT_SIZE = 7;
	defparam lut_9892.mask = 128'h37ff37ff3fff3fffaa88a08088888080;

	lut_sub lut_9897 ({sk[2106], x12475x, x12480x, x12481x, x22230x}, x12486x);
	defparam lut_9897.LUT_SIZE = 5;
	defparam lut_9897.mask = 32'h5f5fbfff;

	lut_sub lut_9902 ({sk[2107], i_9_, n_n518, n_n260, n_n522, x482x, x480x}, x12213x);
	defparam lut_9902.LUT_SIZE = 7;
	defparam lut_9902.mask = 128'h37ff37ff3fff3fff0000000f0077007f;

	lut_sub lut_9907 ({sk[2108], i_9_, n_n526, n_n532, n_n509, n_n260, x581x}, x12214x);
	defparam lut_9907.LUT_SIZE = 7;
	defparam lut_9907.mask = 128'h37ff37ff3fff3fff0003030311131313;

	lut_sub lut_9913 ({sk[2109], x15x, x17x, x478x, x566x}, x12216x);
	defparam lut_9913.LUT_SIZE = 5;
	defparam lut_9913.mask = 32'h5f5f0357;

	lut_sub lut_9916 ({sk[2110], i_9_, i_7_, i_8_, i_6_, n_n260, n_n500}, x12221x);
	defparam lut_9916.LUT_SIZE = 7;
	defparam lut_9916.mask = 128'h37ff37ff3fff3fff0010110000110100;

	lut_sub lut_9923 ({sk[2111], i_9_, i_7_, i_8_, i_6_, n_n260, n_n500}, x12218x);
	defparam lut_9923.LUT_SIZE = 7;
	defparam lut_9923.mask = 128'h37ff37ff3fff3fff0100001001001000;

	lut_sub lut_9928 ({sk[2112], i_9_, n_n534, n_n260, x472x, n_n500, x536x}, x12219x);
	defparam lut_9928.LUT_SIZE = 7;
	defparam lut_9928.mask = 128'h37ff37ff3fff3fff00000033005f007f;

	lut_sub lut_9933 ({sk[2113], i_9_, i_7_, i_8_, i_6_, n_n535, n_n195}, x12165x);
	defparam lut_9933.LUT_SIZE = 7;
	defparam lut_9933.mask = 128'h37ff37ff3fff3fff0001001101010000;

	lut_sub lut_9939 ({sk[2114], i_9_, i_7_, i_8_, i_6_, n_n260, n_n464}, x142x);
	defparam lut_9939.LUT_SIZE = 7;
	defparam lut_9939.mask = 128'h37ff37ff3fff3fff0111010101000110;

	lut_sub lut_9948 ({sk[2115], x18x, x550x, x23x, x531x}, x12161x);
	defparam lut_9948.LUT_SIZE = 5;
	defparam lut_9948.mask = 32'h5f5f111f;

	lut_sub lut_9951 ({sk[2116], x17x, x516x, x505x, x506x, x529x}, x12174x);
	defparam lut_9951.LUT_SIZE = 6;
	defparam lut_9951.mask = 64'h77ff77ff00007fff;

	lut_sub lut_9956 ({sk[2117], i_9_, i_7_, i_8_, i_6_, n_n473, n_n260}, x12175x);
	defparam lut_9956.LUT_SIZE = 7;
	defparam lut_9956.mask = 128'h37ff37ff3fff3fff0010111000000110;

	lut_sub lut_9963 ({sk[2118], i_9_, n_n260, n_n520, n_n500, x49x}, x12181x);
	defparam lut_9963.LUT_SIZE = 6;
	defparam lut_9963.mask = 64'h77ff77ff55575557;

	lut_sub lut_9967 ({sk[2119], i_9_, i_7_, i_8_, i_6_, n_n260, n_n491}, x12182x);
	defparam lut_9967.LUT_SIZE = 7;
	defparam lut_9967.mask = 128'h37ff37ff3fff3fff0100010100000101;

	lut_sub lut_9973 ({sk[2120], x15x, x17x, x584x, x589x}, x305x);
	defparam lut_9973.LUT_SIZE = 5;
	defparam lut_9973.mask = 32'h5f5f0357;

	lut_sub lut_9976 ({sk[2121], i_9_, i_7_, i_8_, i_6_, n_n482, n_n260}, x12188x);
	defparam lut_9976.LUT_SIZE = 7;
	defparam lut_9976.mask = 128'h37ff37ff3fff3fff0010100001001000;

	lut_sub lut_9981 ({sk[2122], i_9_, i_7_, i_8_, i_6_, n_n482, n_n260}, x12187x);
	defparam lut_9981.LUT_SIZE = 7;
	defparam lut_9981.mask = 128'h37ff37ff3fff3fff0001001100010000;

	lut_sub lut_9986 ({sk[2123], x24x, x18x, x485x, x518x, x577x, x546x}, x12663x);
	defparam lut_9986.LUT_SIZE = 7;
	defparam lut_9986.mask = 128'h37ff37ff3fff3fff00005f5f33ff7fff;

	lut_sub lut_9991 ({sk[2124], x24x, x18x, x557x, x572x, x520x, x532x}, x12670x);
	defparam lut_9991.LUT_SIZE = 7;
	defparam lut_9991.mask = 128'h37ff37ff3fff3fff00003fff55557fff;

	lut_sub lut_9996 ({sk[2125], x21x, x510x, x570x, x18x, x577x, x532x}, x22302x);
	defparam lut_9996.LUT_SIZE = 7;
	defparam lut_9996.mask = 128'h37ff37ff3fff3ffffff0f0f088808080;

	lut_sub lut_10001 ({sk[2126], x12x, x517x, x594x, x585x}, x12655x);
	defparam lut_10001.LUT_SIZE = 5;
	defparam lut_10001.mask = 32'h5f5f007f;

	lut_sub lut_10005 ({sk[2127], x539x, x18x, x475x, x593x}, x12662x);
	defparam lut_10005.LUT_SIZE = 5;
	defparam lut_10005.mask = 32'h5f5f070f;

	lut_sub lut_10009 ({sk[2128], x22x, x18x, x525x, x553x, n_n5104, n_n5011}, x22217x);
	defparam lut_10009.LUT_SIZE = 7;
	defparam lut_10009.mask = 128'h37ff37ff3fff3fff8888880080808000;

	lut_sub lut_10014 ({sk[2129], x11x, x20x, x23x, x566x, x589x, x576x}, x12678x);
	defparam lut_10014.LUT_SIZE = 7;
	defparam lut_10014.mask = 128'h37ff37ff3fff3fff00550f5f77777f7f;

	lut_sub lut_10019 ({sk[2130], x25x, x17x, x572x, x564x, x566x}, x12677x);
	defparam lut_10019.LUT_SIZE = 6;
	defparam lut_10019.mask = 64'h77ff77ff003f557f;

	lut_sub lut_10023 ({sk[2131], x25x, x14x, x552x, x503x}, x12680x);
	defparam lut_10023.LUT_SIZE = 5;
	defparam lut_10023.mask = 32'h5f5f0537;

	lut_sub lut_10026 ({sk[2132], x21x, x17x, x478x, x530x}, x12681x);
	defparam lut_10026.LUT_SIZE = 5;
	defparam lut_10026.mask = 32'h5f5f0357;

	lut_sub lut_10029 ({sk[2133], i_9_, i_5_, i_3_, i_4_, n_n534, n_n130}, x279x);
	defparam lut_10029.LUT_SIZE = 7;
	defparam lut_10029.mask = 128'h37ff37ff3fff3fff0001000000010000;

	lut_sub lut_10032 ({sk[2134], x11x, x10x, x23x, x547x, x594x, x593x}, x13450x);
	defparam lut_10032.LUT_SIZE = 7;
	defparam lut_10032.mask = 128'h37ff37ff3fff3fff000f777f0f0f7f7f;

	lut_sub lut_10037 ({sk[2135], i_9_, i_7_, i_8_, i_6_, n_n390, n_n535}, x13451x);
	defparam lut_10037.LUT_SIZE = 7;
	defparam lut_10037.mask = 128'h37ff37ff3fff3fff0011001001010000;

	lut_sub lut_10043 ({sk[2136], x11x, x10x, x561x, x556x}, x401x);
	defparam lut_10043.LUT_SIZE = 5;
	defparam lut_10043.mask = 32'h5f5f0537;

	lut_sub lut_10046 ({sk[2137], x10x, x24x, x571x, x562x}, x13460x);
	defparam lut_10046.LUT_SIZE = 5;
	defparam lut_10046.mask = 32'h5f5f0357;

	lut_sub lut_10049 ({sk[2138], i_9_, n_n390, x557x, x573x, x401x}, x13463x);
	defparam lut_10049.LUT_SIZE = 6;
	defparam lut_10049.mask = 64'h77ff77ff5555557f;

	lut_sub lut_10053 ({sk[2139], i_9_, x15x, n_n455, n_n473, x528x, x416x}, x13474x);
	defparam lut_10053.LUT_SIZE = 7;
	defparam lut_10053.mask = 128'h37ff37ff3fff3fff5555555f5577557f;

	lut_sub lut_10057 ({sk[2140], i_9_, i_7_, i_8_, i_6_, n_n455, n_n473}, x13475x);
	defparam lut_10057.LUT_SIZE = 7;
	defparam lut_10057.mask = 128'h37ff37ff3fff3fff0000101010101000;

	lut_sub lut_10063 ({sk[2141], x14x, x490x, x23x, x526x}, x14315x);
	defparam lut_10063.LUT_SIZE = 5;
	defparam lut_10063.mask = 32'h5f5f111f;

	lut_sub lut_10066 ({sk[2142], x25x, x22x, x14x, x564x, x595x, x551x}, x14316x);
	defparam lut_10066.LUT_SIZE = 7;
	defparam lut_10066.mask = 128'h37ff37ff3fff3fff000f333f555f777f;

	lut_sub lut_10070 ({sk[2143], x11x, x483x, x14x, x20x, x475x, x551x}, x22263x);
	defparam lut_10070.LUT_SIZE = 7;
	defparam lut_10070.mask = 128'h37ff37ff3fff3fffffccf0c0aa88a080;

	lut_sub lut_10079 ({sk[2144], x15x, x595x, x14315x, x14316x, x22263x}, n_n3560);
	defparam lut_10079.LUT_SIZE = 6;
	defparam lut_10079.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_10084 ({sk[2145], i_9_, i_7_, i_8_, i_6_, n_n536, n_n500}, x15512x);
	defparam lut_10084.LUT_SIZE = 7;
	defparam lut_10084.mask = 128'h37ff37ff3fff3fff0100000001000110;

	lut_sub lut_10089 ({sk[2146], i_9_, i_7_, i_8_, i_6_, n_n455, n_n500}, x12489x);
	defparam lut_10089.LUT_SIZE = 7;
	defparam lut_10089.mask = 128'h37ff37ff3fff3fff0100000101000100;

	lut_sub lut_10094 ({sk[2147], x15x, x22x, x541x, n_n1677, x12489x}, n_n1495);
	defparam lut_10094.LUT_SIZE = 6;
	defparam lut_10094.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_10099 ({sk[2148], x15x, x13x, x24x, x480x, x476x}, x12492x);
	defparam lut_10099.LUT_SIZE = 6;
	defparam lut_10099.mask = 64'h77ff77ff05375577;

	lut_sub lut_10103 ({sk[2149], x544x, x23x, n_n4472, x194x, x199x, x12492x}, n_n1496);
	defparam lut_10103.LUT_SIZE = 7;
	defparam lut_10103.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_10109 ({sk[2150], i_9_, i_7_, i_8_, i_6_, n_n260, n_n535}, n_n1468);
	defparam lut_10109.LUT_SIZE = 7;
	defparam lut_10109.mask = 128'h37ff37ff3fff3fff0101011011111000;

	lut_sub lut_10119 ({sk[2151], i_9_, i_7_, i_8_, i_6_, n_n518, n_n260}, x12235x);
	defparam lut_10119.LUT_SIZE = 7;
	defparam lut_10119.mask = 128'h37ff37ff3fff3fff0100011001000000;

	lut_sub lut_10124 ({sk[2152], x539x, x17x, x552x, x23x}, x12233x);
	defparam lut_10124.LUT_SIZE = 5;
	defparam lut_10124.mask = 32'h5f5f111f;

	lut_sub lut_10127 ({sk[2153], i_9_, n_n518, n_n528, n_n325, n_n530, x546x}, x11868x);
	defparam lut_10127.LUT_SIZE = 7;
	defparam lut_10127.mask = 128'h37ff37ff3fff3fff0000030f0505070f;

	lut_sub lut_10133 ({sk[2154], x22x, x14x, x502x, x511x}, x381x);
	defparam lut_10133.LUT_SIZE = 5;
	defparam lut_10133.mask = 32'h5f5f0357;

	lut_sub lut_10136 ({sk[2155], i_9_, n_n536, x482x, x581x, x124x}, x15517x);
	defparam lut_10136.LUT_SIZE = 6;
	defparam lut_10136.mask = 64'h77ff77ff5555557f;

	lut_sub lut_10140 ({sk[2156], i_9_, i_7_, i_8_, i_6_, n_n536, n_n509}, x15518x);
	defparam lut_10140.LUT_SIZE = 7;
	defparam lut_10140.mask = 128'h37ff37ff3fff3fff0001010001000110;

	lut_sub lut_10146 ({sk[2157], i_9_, i_7_, i_8_, i_6_, n_n390, n_n509}, x15109x);
	defparam lut_10146.LUT_SIZE = 7;
	defparam lut_10146.mask = 128'h37ff37ff3fff3fff0101010000010001;

	lut_sub lut_10152 ({sk[2158], x25x, x10x, x474x, x472x, x561x, n_n4611}, x22251x);
	defparam lut_10152.LUT_SIZE = 7;
	defparam lut_10152.mask = 128'h37ff37ff3fff3fffaaaaa00088888000;

	lut_sub lut_10157 ({sk[2159], x10x, x20x, x478x, x23x, x479x, x556x}, x22252x);
	defparam lut_10157.LUT_SIZE = 7;
	defparam lut_10157.mask = 128'h37ff37ff3fff3ffffcfccccca8008800;

	lut_sub lut_10162 ({sk[2160], i_9_, x538x, n_n455, n_n473, n_n534, x580x}, x12504x);
	defparam lut_10162.LUT_SIZE = 7;
	defparam lut_10162.mask = 128'h37ff37ff3fff3fff00030003005700ff;

	lut_sub lut_10167 ({sk[2161], i_9_, i_7_, i_8_, i_6_, n_n482, n_n455}, x12506x);
	defparam lut_10167.LUT_SIZE = 7;
	defparam lut_10167.mask = 128'h37ff37ff3fff3fff0001111100011100;

	lut_sub lut_10176 ({sk[2162], n_n4247, n_n1491, n_n3879, x12504x, x12506x}, n_n1423);
	defparam lut_10176.LUT_SIZE = 6;
	defparam lut_10176.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_10182 ({sk[2163], i_9_, i_7_, i_8_, i_6_, n_n464, n_n65}, n_n1429);
	defparam lut_10182.LUT_SIZE = 7;
	defparam lut_10182.mask = 128'h37ff37ff3fff3fff0111010010111000;

	lut_sub lut_10191 ({sk[2164], i_9_, i_7_, i_8_, i_6_, x515x}, x12366x);
	defparam lut_10191.LUT_SIZE = 6;
	defparam lut_10191.mask = 64'h77ff77ff11000000;

	lut_sub lut_10194 ({sk[2165], i_9_, n_n473, n_n522, x502x, n_n65, x528x}, x12368x);
	defparam lut_10194.LUT_SIZE = 7;
	defparam lut_10194.mask = 128'h37ff37ff3fff3fff0000003313131333;

	lut_sub lut_10199 ({sk[2166], x19x, x503x, x116x, n_n1429, x12366x, x12368x}, n_n1402);
	defparam lut_10199.LUT_SIZE = 7;
	defparam lut_10199.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_10205 ({sk[2167], x25x, x515x, x592x, x21x, n_n3019, x204x}, x12379x);
	defparam lut_10205.LUT_SIZE = 7;
	defparam lut_10205.mask = 128'h37ff37ff3fff3fff777f777f777fffff;

	lut_sub lut_10210 ({sk[2168], n_n1432, x12375x, x12376x}, x12380x);
	defparam lut_10210.LUT_SIZE = 4;
	defparam lut_10210.mask = 16'h0f7f;

	lut_sub lut_10214 ({sk[2169], x22x, x16x, x23x, x488x, x540x, x496x}, x22237x);
	defparam lut_10214.LUT_SIZE = 7;
	defparam lut_10214.mask = 128'h37ff37ff3fff3fffff88f080aa88a080;

	lut_sub lut_10221 ({sk[2170], x16x, x586x, x427x, x302x, x22237x}, n_n957);
	defparam lut_10221.LUT_SIZE = 6;
	defparam lut_10221.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_10226 ({sk[2171], x15x, x13x, x11x, x563x, x494x, x476x}, x22236x);
	defparam lut_10226.LUT_SIZE = 7;
	defparam lut_10226.mask = 128'h37ff37ff3fff3fffffaac080aaaa8080;

	lut_sub lut_10231 ({sk[2172], x13x, x570x, x491x, x480x, x536x}, x22271x);
	defparam lut_10231.LUT_SIZE = 6;
	defparam lut_10231.mask = 64'h77ff77ffffff8000;

	lut_sub lut_10234 ({sk[2173], x25x, x542x, x22236x, x22271x}, n_n956);
	defparam lut_10234.LUT_SIZE = 5;
	defparam lut_10234.mask = 32'h5f5feeef;

	lut_sub lut_10238 ({sk[2174], x21x, x17x, x529x, x531x}, x11685x);
	defparam lut_10238.LUT_SIZE = 5;
	defparam lut_10238.mask = 32'h5f5f0357;

	lut_sub lut_10241 ({sk[2175], x21x, x18x, x478x, x23x, x566x, x589x}, x11687x);
	defparam lut_10241.LUT_SIZE = 7;
	defparam lut_10241.mask = 128'h37ff37ff3fff3fff030303ff575757ff;

	lut_sub lut_10245 ({sk[2176], x11x, x24x, x18x, x481x, x566x, x589x}, x22267x);
	defparam lut_10245.LUT_SIZE = 7;
	defparam lut_10245.mask = 128'h37ff37ff3fff3ffffff0aaa0ccc08880;

	lut_sub lut_10254 ({sk[2177], x15x, x19x, x475x, x555x, x11698x, x11697x}, n_n945);
	defparam lut_10254.LUT_SIZE = 7;
	defparam lut_10254.mask = 128'h37ff37ff3fff3fff777777ff7f7f7fff;

	lut_sub lut_10259 ({sk[2178], x15x, x554x, n_n5087, x11716x, x11717x, x11718x}, n_n948);
	defparam lut_10259.LUT_SIZE = 7;
	defparam lut_10259.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_10265 ({sk[2179], x18x, x493x, n_n5011, x11722x, x11723x, x11725x}, n_n949);
	defparam lut_10265.LUT_SIZE = 7;
	defparam lut_10265.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_10271 ({sk[2180], x25x, x592x, x19x, x510x, x116x, x22235x}, x11733x);
	defparam lut_10271.LUT_SIZE = 7;
	defparam lut_10271.mask = 128'h37ff37ff3fff3fffbbbfbbbfbbbfffff;

	lut_sub lut_10276 ({sk[2181], x11705x, x11712x, x11710x, x11711x, x22234x}, x11735x);
	defparam lut_10276.LUT_SIZE = 6;
	defparam lut_10276.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_10282 ({sk[2182], n_n945, n_n948, n_n949, x11733x, x11735x}, n_n937);
	defparam lut_10282.LUT_SIZE = 6;
	defparam lut_10282.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_10288 ({sk[2183], x25x, x21x, x10x, x24x, x561x, x518x}, x22148x);
	defparam lut_10288.LUT_SIZE = 7;
	defparam lut_10288.mask = 128'h37ff37ff3fff3ffffca8cc88cc88cc88;

	lut_sub lut_10293 ({sk[2184], x10x, x574x, x272x, x271x, x22148x}, n_n3562);
	defparam lut_10293.LUT_SIZE = 6;
	defparam lut_10293.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_10298 ({sk[2185], x22x, x13x, x519x, x586x, x503x, x523x}, x14301x);
	defparam lut_10298.LUT_SIZE = 7;
	defparam lut_10298.mask = 128'h37ff37ff3fff3fff00003fff55557fff;

	lut_sub lut_10303 ({sk[2186], x15x, x13x, x505x, x543x}, x14299x);
	defparam lut_10303.LUT_SIZE = 5;
	defparam lut_10303.mask = 32'h5f5f0357;

	lut_sub lut_10306 ({sk[2187], x11x, x523x, x65x, x14301x, x14299x}, n_n3564);
	defparam lut_10306.LUT_SIZE = 6;
	defparam lut_10306.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_10311 ({sk[2188], x10x, x20x, x547x, x546x}, x237x);
	defparam lut_10311.LUT_SIZE = 5;
	defparam lut_10311.mask = 32'h5f5f0357;

	lut_sub lut_10314 ({sk[2189], x15x, x11x, x10x, x477x, x479x}, n_n2036);
	defparam lut_10314.LUT_SIZE = 6;
	defparam lut_10314.mask = 64'h77ff77ff03575757;

	lut_sub lut_10318 ({sk[2190], i_9_, i_7_, i_8_, i_6_}, x600x);
	defparam lut_10318.LUT_SIZE = 5;
	defparam lut_10318.mask = 32'h5f5f2800;

	lut_sub lut_10321 ({sk[2191], i_9_, n_n390, n_n532, n_n535, x523x, x600x}, x12524x);
	defparam lut_10321.LUT_SIZE = 7;
	defparam lut_10321.mask = 128'h37ff37ff3fff3fff1111111f1111111f;

	lut_sub lut_10325 ({sk[2192], x15x, x11x, x10x, x547x, x548x}, x12523x);
	defparam lut_10325.LUT_SIZE = 6;
	defparam lut_10325.mask = 64'h77ff77ff05373737;

	lut_sub lut_10329 ({sk[2193], x22x, x10x, x550x, x523x, x12524x, x12523x}, n_n1489);
	defparam lut_10329.LUT_SIZE = 7;
	defparam lut_10329.mask = 128'h37ff37ff3fff3fff777777ff7f7f7fff;

	lut_sub lut_10334 ({sk[2194], x22x, x13x, x547x, x527x, x528x}, x22284x);
	defparam lut_10334.LUT_SIZE = 6;
	defparam lut_10334.mask = 64'h77ff77ffff88f080;

	lut_sub lut_10339 ({sk[2195], x10x, x594x, n_n3871, n_n2401, x22284x}, x12534x);
	defparam lut_10339.LUT_SIZE = 6;
	defparam lut_10339.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_10344 ({sk[2196], x25x, x20x, x542x, x541x, x12512x, x22229x}, x12515x);
	defparam lut_10344.LUT_SIZE = 7;
	defparam lut_10344.mask = 128'h37ff37ff3fff3fffbbbbbfbfbbffbfff;

	lut_sub lut_10349 ({sk[2197], i_9_, i_7_, i_8_, i_6_, n_n325, n_n535}, x12414x);
	defparam lut_10349.LUT_SIZE = 7;
	defparam lut_10349.mask = 128'h37ff37ff3fff3fff1010000010000010;

	lut_sub lut_10354 ({sk[2198], i_9_, i_7_, i_8_, i_6_, n_n518, n_n325}, x12415x);
	defparam lut_10354.LUT_SIZE = 7;
	defparam lut_10354.mask = 128'h37ff37ff3fff3fff0001010101010000;

	lut_sub lut_10360 ({sk[2199], i_9_, x25x, n_n390, n_n473, x510x, x157x}, x12425x);
	defparam lut_10360.LUT_SIZE = 7;
	defparam lut_10360.mask = 128'h37ff37ff3fff3fff5555555f5577557f;

	lut_sub lut_10364 ({sk[2200], x21x, x10x, x20x, x582x, x493x}, x12424x);
	defparam lut_10364.LUT_SIZE = 6;
	defparam lut_10364.mask = 64'h77ff77ff03573377;

	lut_sub lut_10368 ({sk[2201], x11x, x10x, x24x, x507x, x580x, x502x}, x22224x);
	defparam lut_10368.LUT_SIZE = 7;
	defparam lut_10368.mask = 128'h37ff37ff3fff3ffffff08880f0f08080;

	lut_sub lut_10373 ({sk[2202], x14x, x20x, x565x, x574x}, x259x);
	defparam lut_10373.LUT_SIZE = 5;
	defparam lut_10373.mask = 32'h5f5f0357;

	lut_sub lut_10376 ({sk[2203], x22x, x13x, x518x, x541x, x536x}, n_n897);
	defparam lut_10376.LUT_SIZE = 6;
	defparam lut_10376.mask = 64'h77ff77ff005f337f;

	lut_sub lut_10380 ({sk[2204], i_9_, n_n526, n_n482, n_n390, x570x, x587x}, x12551x);
	defparam lut_10380.LUT_SIZE = 7;
	defparam lut_10380.mask = 128'h37ff37ff3fff3fff0000000f0707070f;

	lut_sub lut_10385 ({sk[2205], x10x, x24x, x561x, x564x}, x270x);
	defparam lut_10385.LUT_SIZE = 5;
	defparam lut_10385.mask = 32'h5f5f0357;

	lut_sub lut_10388 ({sk[2206], i_9_, n_n526, n_n390, n_n509, n_n520, x562x}, x12540x);
	defparam lut_10388.LUT_SIZE = 7;
	defparam lut_10388.mask = 128'h37ff37ff3fff3fff0003000f0057005f;

	lut_sub lut_10394 ({sk[2207], x22x, x521x, x10x, x583x}, x46x);
	defparam lut_10394.LUT_SIZE = 5;
	defparam lut_10394.mask = 32'h5f5f0357;

	lut_sub lut_10397 ({sk[2208], i_9_, i_5_, i_3_, i_4_, n_n390, n_n522}, x255x);
	defparam lut_10397.LUT_SIZE = 7;
	defparam lut_10397.mask = 128'h37ff37ff3fff3fff0001000000010000;

	lut_sub lut_10400 ({sk[2209], i_9_, i_7_, i_8_, i_6_, n_n518, n_n390}, n_n1487);
	defparam lut_10400.LUT_SIZE = 7;
	defparam lut_10400.mask = 128'h37ff37ff3fff3fff0011101011111000;

	lut_sub lut_10410 ({sk[2210], x15x, x561x, n_n1649, n_n4640, n_n1648, n_n1646}, x12559x);
	defparam lut_10410.LUT_SIZE = 7;
	defparam lut_10410.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_10416 ({sk[2211], x15x, x10x, x558x, x584x, x582x}, x12550x);
	defparam lut_10416.LUT_SIZE = 6;
	defparam lut_10416.mask = 64'h77ff77ff003f557f;

	lut_sub lut_10420 ({sk[2212], x10x, x23x, x561x, x574x, x560x}, x12554x);
	defparam lut_10420.LUT_SIZE = 6;
	defparam lut_10420.mask = 64'h77ff77ff000f777f;

	lut_sub lut_10424 ({sk[2213], x492x, x22x, x21x, x10x, x586x, x571x}, x22228x);
	defparam lut_10424.LUT_SIZE = 7;
	defparam lut_10424.mask = 128'h37ff37ff3fff3ffffca8a8a8f0a0a0a0;

	lut_sub lut_10429 ({sk[2214], x401x, x12551x, x12550x, x12554x, x22228x}, x12560x);
	defparam lut_10429.LUT_SIZE = 6;
	defparam lut_10429.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_10435 ({sk[2215], i_9_, i_7_, i_8_, i_6_, n_n390, n_n509}, x12563x);
	defparam lut_10435.LUT_SIZE = 7;
	defparam lut_10435.mask = 128'h37ff37ff3fff3fff0000000100010101;

	lut_sub lut_10440 ({sk[2216], x10x, x472x, n_n4611, x270x, x12540x, n_n1487}, x12566x);
	defparam lut_10440.LUT_SIZE = 7;
	defparam lut_10440.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_10446 ({sk[2217], x15x, x523x, n_n4560, x213x, x276x, x237x}, x12533x);
	defparam lut_10446.LUT_SIZE = 7;
	defparam lut_10446.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_10452 ({sk[2218], x16x, x21x, x490x, x497x, x517x}, n_n1703);
	defparam lut_10452.LUT_SIZE = 6;
	defparam lut_10452.mask = 64'h77ff77ff00335f7f;

	lut_sub lut_10456 ({sk[2219], i_9_, n_n536, n_n532, n_n509, x53x}, x12572x);
	defparam lut_10456.LUT_SIZE = 6;
	defparam lut_10456.mask = 64'h77ff77ff55575557;

	lut_sub lut_10460 ({sk[2220], i_9_, i_7_, i_8_, i_6_, n_n536, n_n535}, n_n1508);
	defparam lut_10460.LUT_SIZE = 7;
	defparam lut_10460.mask = 128'h37ff37ff3fff3fff0101011101010110;

	lut_sub lut_10470 ({sk[2221], i_9_, i_7_, i_8_, i_6_, x541x, x476x}, x15835x);
	defparam lut_10470.LUT_SIZE = 7;
	defparam lut_10470.mask = 128'h37ff37ff3fff3fff0050003500000000;

	lut_sub lut_10474 ({sk[2222], x13x, x477x, x478x, x481x, x560x}, x22085x);
	defparam lut_10474.LUT_SIZE = 6;
	defparam lut_10474.mask = 64'h77ff77ffffff8000;

	lut_sub lut_10477 ({sk[2223], x15x, x544x, x23x, x542x, x15835x, x22085x}, x15838x);
	defparam lut_10477.LUT_SIZE = 7;
	defparam lut_10477.mask = 128'h37ff37ff3fff3fffbbbbbbffbfbfbfff;

	lut_sub lut_10482 ({sk[2224], x22x, x14x, x489x, x511x, x15852x, x15851x}, n_n1722);
	defparam lut_10482.LUT_SIZE = 7;
	defparam lut_10482.mask = 128'h37ff37ff3fff3fff777777ff7f7f7fff;

	lut_sub lut_10487 ({sk[2225], i_9_, i_1_, i_2_, i_0_, x538x, x594x}, x15855x);
	defparam lut_10487.LUT_SIZE = 7;
	defparam lut_10487.mask = 128'h37ff37ff3fff3fff0000000000005030;

	lut_sub lut_10490 ({sk[2226], x22x, x17x, x23x, x512x, x566x, x502x}, x15858x);
	defparam lut_10490.LUT_SIZE = 7;
	defparam lut_10490.mask = 128'h37ff37ff3fff3fff003355770f3f5f7f;

	lut_sub lut_10494 ({sk[2227], x20x, x487x, n_n5257, x15845x, x15844x, x15898x}, x15899x);
	defparam lut_10494.LUT_SIZE = 7;
	defparam lut_10494.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_10500 ({sk[2228], x22x, x21x, x23x, x589x, x576x, x553x}, x22089x);
	defparam lut_10500.LUT_SIZE = 7;
	defparam lut_10500.mask = 128'h37ff37ff3fff3fffffaac080aaaa8080;

	lut_sub lut_10505 ({sk[2229], n_n1722, x15855x, x15858x, x15899x, x22089x}, x15902x);
	defparam lut_10505.LUT_SIZE = 6;
	defparam lut_10505.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_10511 ({sk[2230], x25x, x567x, x136x, x15864x, x15862x}, n_n1720);
	defparam lut_10511.LUT_SIZE = 6;
	defparam lut_10511.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_10516 ({sk[2231], x509x, x18x, x586x, x508x, x15883x, x15885x}, x15887x);
	defparam lut_10516.LUT_SIZE = 7;
	defparam lut_10516.mask = 128'h37ff37ff3fff3fff77777fff7777ffff;

	lut_sub lut_10522 ({sk[2232], x21x, x555x, x15891x, x15893x, x22320x}, n_n1716);
	defparam lut_10522.LUT_SIZE = 6;
	defparam lut_10522.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_10527 ({sk[2233], x18x, x12x, x494x, x525x, x15871x, x15870x}, n_n1718);
	defparam lut_10527.LUT_SIZE = 7;
	defparam lut_10527.mask = 128'h37ff37ff3fff3fff777777ff7f7f7fff;

	lut_sub lut_10532 ({sk[2234], x15x, x568x, x578x, x15877x, x22088x}, n_n1717);
	defparam lut_10532.LUT_SIZE = 6;
	defparam lut_10532.mask = 64'h77ff77ffbbbbbfff;

	lut_sub lut_10537 ({sk[2235], n_n1720, x15887x, n_n1716, n_n1718, n_n1717}, x15903x);
	defparam lut_10537.LUT_SIZE = 6;
	defparam lut_10537.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_10543 ({sk[2236], x16x, x20x, x587x, x498x}, x15905x);
	defparam lut_10543.LUT_SIZE = 5;
	defparam lut_10543.mask = 32'h5f5f0537;

	lut_sub lut_10546 ({sk[2237], x16x, x21x, x495x, x528x}, x15906x);
	defparam lut_10546.LUT_SIZE = 5;
	defparam lut_10546.mask = 32'h5f5f0357;

	lut_sub lut_10549 ({sk[2238], x16x, x500x, x23x, x508x, x488x}, x15908x);
	defparam lut_10549.LUT_SIZE = 6;
	defparam lut_10549.mask = 64'h77ff77ff000f777f;

	lut_sub lut_10553 ({sk[2239], x16x, x586x, x574x, x15905x, x15906x, x15908x}, n_n1730);
	defparam lut_10553.LUT_SIZE = 7;
	defparam lut_10553.mask = 128'h37ff37ff3fff3fff7f7f7f7f7fffffff;

	lut_sub lut_10559 ({sk[2240], i_9_, i_1_, i_2_, i_0_, x494x, x235x}, x15914x);
	defparam lut_10559.LUT_SIZE = 7;
	defparam lut_10559.mask = 128'h37ff37ff3fff3fff5555555555555755;

	lut_sub lut_10562 ({sk[2241], x25x, x13x, x539x, n_n4433, x23x, x540x}, x22087x);
	defparam lut_10562.LUT_SIZE = 7;
	defparam lut_10562.mask = 128'h37ff37ff3fff3fffe0e0e000a0a0a000;

	lut_sub lut_10567 ({sk[2242], x21x, x13x, x540x, x593x, x15914x, x22087x}, n_n1729);
	defparam lut_10567.LUT_SIZE = 7;
	defparam lut_10567.mask = 128'h37ff37ff3fff3fffbbbbbfbfbbffbfff;

	lut_sub lut_10572 ({sk[2243], x15x, x538x, x21x, x14x, x588x, x518x}, x15930x);
	defparam lut_10572.LUT_SIZE = 7;
	defparam lut_10572.mask = 128'h37ff37ff3fff3fff05370f3f37373f3f;

	lut_sub lut_10577 ({sk[2244], x492x, x22x, x14x, x557x, x537x, x575x}, x22333x);
	defparam lut_10577.LUT_SIZE = 7;
	defparam lut_10577.mask = 128'h37ff37ff3fff3fffffc0aa80ff00aa00;

	lut_sub lut_10582 ({sk[2245], x14x, x562x, x15930x, x22333x}, x15932x);
	defparam lut_10582.LUT_SIZE = 5;
	defparam lut_10582.mask = 32'h5f5fbbbf;

	lut_sub lut_10586 ({sk[2246], i_9_, n_n526, n_n482, x11x, n_n390, x488x}, x15920x);
	defparam lut_10586.LUT_SIZE = 7;
	defparam lut_10586.mask = 128'h37ff37ff3fff3fff0003003311131133;

	lut_sub lut_10591 ({sk[2247], x10x, x516x, x522x, x23x, x595x, x551x}, x15924x);
	defparam lut_10591.LUT_SIZE = 7;
	defparam lut_10591.mask = 128'h37ff37ff3fff3fff0707070707ffffff;

	lut_sub lut_10596 ({sk[2248], x11x, x20x, x595x, x526x, n_n4678, n_n4700}, x22084x);
	defparam lut_10596.LUT_SIZE = 7;
	defparam lut_10596.mask = 128'h37ff37ff3fff3fff8888880080808000;

	lut_sub lut_10601 ({sk[2249], n_n1764, x15920x, n_n1760, x15924x, x22084x}, x15933x);
	defparam lut_10601.LUT_SIZE = 6;
	defparam lut_10601.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_10607 ({sk[2250], x15x, x10x, x489x, x551x}, x13628x);
	defparam lut_10607.LUT_SIZE = 5;
	defparam lut_10607.mask = 32'h5f5f0357;

	lut_sub lut_10610 ({sk[2251], x10x, x507x, x14x, x23x, x494x, x524x}, x13629x);
	defparam lut_10610.LUT_SIZE = 7;
	defparam lut_10610.mask = 128'h37ff37ff3fff3fff00330f3f55775f7f;

	lut_sub lut_10614 ({sk[2252], x25x, x21x, x507x, x23x, x582x, x551x}, x22316x);
	defparam lut_10614.LUT_SIZE = 7;
	defparam lut_10614.mask = 128'h37ff37ff3fff3ffffcfca8a8fc00a800;

	lut_sub lut_10623 ({sk[2253], x10x, x503x, x13628x, x13629x, x22316x}, n_n3931);
	defparam lut_10623.LUT_SIZE = 6;
	defparam lut_10623.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_10628 ({sk[2254], i_9_, i_7_, i_8_, i_6_, x589x, x576x}, x13632x);
	defparam lut_10628.LUT_SIZE = 7;
	defparam lut_10628.mask = 128'h37ff37ff3fff3fff5000003000000000;

	lut_sub lut_10631 ({sk[2255], x17x, x20x, x587x, x576x}, x13634x);
	defparam lut_10631.LUT_SIZE = 5;
	defparam lut_10631.mask = 32'h5f5f0537;

	lut_sub lut_10634 ({sk[2256], x25x, x21x, x17x, x484x, x596x, x593x}, x13635x);
	defparam lut_10634.LUT_SIZE = 7;
	defparam lut_10634.mask = 128'h37ff37ff3fff3fff00550f5f33773f7f;

	lut_sub lut_10638 ({sk[2257], x25x, x589x, n_n4846, x13632x, x13634x, x13635x}, n_n3929);
	defparam lut_10638.LUT_SIZE = 7;
	defparam lut_10638.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_10644 ({sk[2258], i_9_, i_7_, i_8_, i_6_, n_n260, n_n491}, x14733x);
	defparam lut_10644.LUT_SIZE = 7;
	defparam lut_10644.mask = 128'h37ff37ff3fff3fff0000000101010001;

	lut_sub lut_10649 ({sk[2259], i_9_, i_7_, i_8_, i_6_, n_n473, n_n65}, n_n3661);
	defparam lut_10649.LUT_SIZE = 7;
	defparam lut_10649.mask = 128'h37ff37ff3fff3fff0110101101001110;

	lut_sub lut_10659 ({sk[2260], i_9_, i_7_, i_8_, i_6_, n_n518, n_n325}, n_n2982);
	defparam lut_10659.LUT_SIZE = 7;
	defparam lut_10659.mask = 128'h37ff37ff3fff3fff0101011100011110;

	lut_sub lut_10669 ({sk[2261], x21x, x12x, x554x, x585x}, x15604x);
	defparam lut_10669.LUT_SIZE = 5;
	defparam lut_10669.mask = 32'h5f5f0537;

	lut_sub lut_10672 ({sk[2262], x22x, x554x, x34x, x122x, x143x, x15604x}, n_n2953);
	defparam lut_10672.LUT_SIZE = 7;
	defparam lut_10672.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_10678 ({sk[2263], x18x, x20x, x522x, x513x}, x15608x);
	defparam lut_10678.LUT_SIZE = 5;
	defparam lut_10678.mask = 32'h5f5f0537;

	lut_sub lut_10681 ({sk[2264], x25x, x22x, x18x, x502x, x513x, x532x}, x15609x);
	defparam lut_10681.LUT_SIZE = 7;
	defparam lut_10681.mask = 128'h37ff37ff3fff3fff000f333f555f777f;

	lut_sub lut_10685 ({sk[2265], x11x, x24x, x344x, x532x, x15608x, x15609x}, n_n2955);
	defparam lut_10685.LUT_SIZE = 7;
	defparam lut_10685.mask = 128'h37ff37ff3fff3fff77ff7fff7fff7fff;

	lut_sub lut_10691 ({sk[2266], x22x, x545x, x12x, x532x}, x15613x);
	defparam lut_10691.LUT_SIZE = 5;
	defparam lut_10691.mask = 32'h5f5f0357;

	lut_sub lut_10694 ({sk[2267], i_9_, i_7_, i_8_, i_6_, n_n195, n_n464}, x15617x);
	defparam lut_10694.LUT_SIZE = 7;
	defparam lut_10694.mask = 128'h37ff37ff3fff3fff1010100000101000;

	lut_sub lut_10700 ({sk[2268], x25x, x15x, x554x, x15613x, x15617x}, x15618x);
	defparam lut_10700.LUT_SIZE = 6;
	defparam lut_10700.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_10705 ({sk[2269], x11x, x12x, x20x, x482x, x581x, x598x}, x15623x);
	defparam lut_10705.LUT_SIZE = 7;
	defparam lut_10705.mask = 128'h37ff37ff3fff3fff00553f7f55557f7f;

	lut_sub lut_10710 ({sk[2270], i_9_, i_7_, i_8_, i_6_, n_n518, n_n130}, x15624x);
	defparam lut_10710.LUT_SIZE = 7;
	defparam lut_10710.mask = 128'h37ff37ff3fff3fff0000100001101010;

	lut_sub lut_10716 ({sk[2271], x11x, x24x, x12x, x518x, x486x, x556x}, x15630x);
	defparam lut_10716.LUT_SIZE = 7;
	defparam lut_10716.mask = 128'h37ff37ff3fff3fff005f337f337f337f;

	lut_sub lut_10721 ({sk[2272], x12x, x563x, x155x, n_n3051, x15630x}, x15633x);
	defparam lut_10721.LUT_SIZE = 6;
	defparam lut_10721.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_10726 ({sk[2273], i_9_, i_7_, i_8_, i_6_, n_n509, n_n130}, x15628x);
	defparam lut_10726.LUT_SIZE = 7;
	defparam lut_10726.mask = 128'h37ff37ff3fff3fff0000001000011100;

	lut_sub lut_10731 ({sk[2274], i_9_, n_n509, n_n522, n_n130, x536x, x286x}, x15629x);
	defparam lut_10731.LUT_SIZE = 7;
	defparam lut_10731.mask = 128'h37ff37ff3fff3fff555555555757575f;

	lut_sub lut_10735 ({sk[2275], x15623x, x15624x, x15628x, x15629x}, x15634x);
	defparam lut_10735.LUT_SIZE = 5;
	defparam lut_10735.mask = 32'h5f5f7fff;

	lut_sub lut_10740 ({sk[2276], i_9_, i_7_, i_8_, i_6_, x590x, x513x}, x15600x);
	defparam lut_10740.LUT_SIZE = 7;
	defparam lut_10740.mask = 128'h37ff37ff3fff3fff3000050000000000;

	lut_sub lut_10743 ({sk[2277], x11x, x18x, x508x, x503x, x513x}, x15601x);
	defparam lut_10743.LUT_SIZE = 6;
	defparam lut_10743.mask = 64'h77ff77ff003f557f;

	lut_sub lut_10747 ({sk[2278], x20x, x577x, x231x, x15636x, x15638x}, x15640x);
	defparam lut_10747.LUT_SIZE = 6;
	defparam lut_10747.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_10752 ({sk[2279], x25x, x14x, x586x, x565x}, x15404x);
	defparam lut_10752.LUT_SIZE = 5;
	defparam lut_10752.mask = 32'h5f5f0357;

	lut_sub lut_10755 ({sk[2280], x22x, x509x, x14x, x493x, x575x, n_n4797}, x22108x);
	defparam lut_10755.LUT_SIZE = 7;
	defparam lut_10755.mask = 128'h37ff37ff3fff3fffaaa0aa0088808800;

	lut_sub lut_10760 ({sk[2281], x11x, x530x, x259x, x15404x, x22108x}, n_n2839);
	defparam lut_10760.LUT_SIZE = 6;
	defparam lut_10760.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_10765 ({sk[2282], x22x, x17x, x519x, x586x, x587x, x576x}, x16184x);
	defparam lut_10765.LUT_SIZE = 7;
	defparam lut_10765.mask = 128'h37ff37ff3fff3fff00003fff55557fff;

	lut_sub lut_10770 ({sk[2283], i_9_, i_7_, i_8_, i_6_, n_n260, n_n491}, x16185x);
	defparam lut_10770.LUT_SIZE = 7;
	defparam lut_10770.mask = 128'h37ff37ff3fff3fff1110000010100000;

	lut_sub lut_10776 ({sk[2284], i_9_, i_7_, i_8_, i_6_, n_n473, n_n130}, x16254x);
	defparam lut_10776.LUT_SIZE = 7;
	defparam lut_10776.mask = 128'h37ff37ff3fff3fff0100101001001000;

	lut_sub lut_10782 ({sk[2285], i_9_, i_7_, i_8_, i_6_, n_n325, n_n500}, n_n1866);
	defparam lut_10782.LUT_SIZE = 7;
	defparam lut_10782.mask = 128'h37ff37ff3fff3fff0101111101100010;

	lut_sub lut_10792 ({sk[2286], i_9_, i_7_, i_8_, i_6_, n_n518, n_n325}, x16130x);
	defparam lut_10792.LUT_SIZE = 7;
	defparam lut_10792.mask = 128'h37ff37ff3fff3fff0101110001101110;

	lut_sub lut_10802 ({sk[2287], i_9_, n_n518, n_n534, n_n535, n_n522, n_n130}, x15950x);
	defparam lut_10802.LUT_SIZE = 7;
	defparam lut_10802.mask = 128'h37ff37ff3fff3fff0101015501010155;

	lut_sub lut_10807 ({sk[2288], i_9_, i_7_, i_8_, i_6_, n_n535, n_n130}, x15951x);
	defparam lut_10807.LUT_SIZE = 7;
	defparam lut_10807.mask = 128'h37ff37ff3fff3fff0000101001001010;

	lut_sub lut_10813 ({sk[2289], x25x, x22x, x18x, x502x, x513x, x532x}, x15954x);
	defparam lut_10813.LUT_SIZE = 7;
	defparam lut_10813.mask = 128'h37ff37ff3fff3fff000f333f555f777f;

	lut_sub lut_10817 ({sk[2290], x24x, x18x, x529x, x527x, x528x, x532x}, x22308x);
	defparam lut_10817.LUT_SIZE = 7;
	defparam lut_10817.mask = 128'h37ff37ff3fff3fffffffc000aaaa8000;

	lut_sub lut_10822 ({sk[2291], x12x, x23x, x549x, x532x}, x15944x);
	defparam lut_10822.LUT_SIZE = 5;
	defparam lut_10822.mask = 32'h5f5f0537;

	lut_sub lut_10825 ({sk[2292], i_9_, i_7_, i_8_, i_6_, n_n509, n_n130}, x15962x);
	defparam lut_10825.LUT_SIZE = 7;
	defparam lut_10825.mask = 128'h37ff37ff3fff3fff0000100010100100;

	lut_sub lut_10830 ({sk[2293], x21x, x12x, x20x, x482x, x581x, x598x}, x15967x);
	defparam lut_10830.LUT_SIZE = 7;
	defparam lut_10830.mask = 128'h37ff37ff3fff3fff00553f7f55557f7f;

	lut_sub lut_10835 ({sk[2294], x22x, x474x, x12x, x477x, x486x}, x15961x);
	defparam lut_10835.LUT_SIZE = 6;
	defparam lut_10835.mask = 64'h77ff77ff030f575f;

	lut_sub lut_10839 ({sk[2295], x15x, x521x, x24x, x12x, x598x}, x15966x);
	defparam lut_10839.LUT_SIZE = 6;
	defparam lut_10839.mask = 64'h77ff77ff05375577;

	lut_sub lut_10843 ({sk[2296], x25x, x539x, x24x, x12x, x564x, x486x}, x22092x);
	defparam lut_10843.LUT_SIZE = 7;
	defparam lut_10843.mask = 128'h37ff37ff3fff3ffffca8f0a0a8a8a0a0;

	lut_sub lut_10848 ({sk[2297], i_9_, i_7_, i_8_, i_6_, n_n482, n_n195}, x15978x);
	defparam lut_10848.LUT_SIZE = 7;
	defparam lut_10848.mask = 128'h37ff37ff3fff3fff0000001001001010;

	lut_sub lut_10853 ({sk[2298], i_9_, i_7_, i_8_, i_6_, n_n491, n_n195}, x15982x);
	defparam lut_10853.LUT_SIZE = 7;
	defparam lut_10853.mask = 128'h37ff37ff3fff3fff0101001000000010;

	lut_sub lut_10858 ({sk[2299], i_9_, n_n325, n_n535, n_n520, x594x, x30x}, x12784x);
	defparam lut_10858.LUT_SIZE = 7;
	defparam lut_10858.mask = 128'h37ff37ff3fff3fff5555555f55557777;

	lut_sub lut_10862 ({sk[2300], i_9_, i_7_, i_8_, i_6_, n_n473, n_n260}, n_n691);
	defparam lut_10862.LUT_SIZE = 7;
	defparam lut_10862.mask = 128'h37ff37ff3fff3fff0101011101110100;

	lut_sub lut_10872 ({sk[2301], i_9_, n_n524, n_n260, n_n491, x20x, x587x}, x12724x);
	defparam lut_10872.LUT_SIZE = 7;
	defparam lut_10872.mask = 128'h37ff37ff3fff3fff0003000f0057005f;

	lut_sub lut_10877 ({sk[2302], i_9_, i_7_, i_8_, i_6_, n_n464, n_n65}, n_n632);
	defparam lut_10877.LUT_SIZE = 7;
	defparam lut_10877.mask = 128'h37ff37ff3fff3fff1111110110111110;

	lut_sub lut_10891 ({sk[2303], i_9_, n_n325, x508x, x505x, x292x}, x12765x);
	defparam lut_10891.LUT_SIZE = 6;
	defparam lut_10891.mask = 64'h77ff77ff5555557f;

	lut_sub lut_10895 ({sk[2304], x15x, x588x, x20x, x511x, n_n2003, x12765x}, x12767x);
	defparam lut_10895.LUT_SIZE = 7;
	defparam lut_10895.mask = 128'h37ff37ff3fff3fff777777ff7f7f7fff;

	lut_sub lut_10900 ({sk[2305], i_9_, i_7_, i_8_, i_6_, n_n482, n_n325}, n_n702);
	defparam lut_10900.LUT_SIZE = 7;
	defparam lut_10900.mask = 128'h37ff37ff3fff3fff0101010101110110;

	lut_sub lut_10910 ({sk[2306], x11x, x14x, x529x, x511x}, x12755x);
	defparam lut_10910.LUT_SIZE = 5;
	defparam lut_10910.mask = 32'h5f5f0357;

	lut_sub lut_10913 ({sk[2307], x25x, x24x, x23x, x530x, x511x, x71x}, x22211x);
	defparam lut_10913.LUT_SIZE = 7;
	defparam lut_10913.mask = 128'h37ff37ff3fff3fffaa88a080a080a080;

	lut_sub lut_10918 ({sk[2308], x381x, n_n702, x12755x, x22211x}, x12768x);
	defparam lut_10918.LUT_SIZE = 5;
	defparam lut_10918.mask = 32'h5f5fbfff;

	lut_sub lut_10923 ({sk[2309], x17x, x20x, x484x, x562x}, x12726x);
	defparam lut_10923.LUT_SIZE = 5;
	defparam lut_10923.mask = 32'h5f5f0357;

	lut_sub lut_10926 ({sk[2310], i_9_, i_7_, i_8_, i_6_, x484x, x566x}, x12727x);
	defparam lut_10926.LUT_SIZE = 7;
	defparam lut_10926.mask = 128'h37ff37ff3fff3fff3000050000000000;

	lut_sub lut_10929 ({sk[2311], x474x, x17x, x472x, x563x}, x12728x);
	defparam lut_10929.LUT_SIZE = 5;
	defparam lut_10929.mask = 32'h5f5f070f;

	lut_sub lut_10933 ({sk[2312], x25x, x17x, x574x, x576x, x12770x, x22212x}, x12773x);
	defparam lut_10933.LUT_SIZE = 7;
	defparam lut_10933.mask = 128'h37ff37ff3fff3fffbbbbbbffbfbfbfff;

	lut_sub lut_10938 ({sk[2313], x330x, n_n696, x12726x, x12727x, x12728x, x12773x}, x12775x);
	defparam lut_10938.LUT_SIZE = 7;
	defparam lut_10938.mask = 128'h37ff37ff3fff3fff7fffffffffffffff;

	lut_sub lut_10945 ({sk[2314], x14x, x17x, x549x, x594x, x585x, x525x}, x12749x);
	defparam lut_10945.LUT_SIZE = 7;
	defparam lut_10945.mask = 128'h37ff37ff3fff3fff00003fff55557fff;

	lut_sub lut_10950 ({sk[2315], n_n834, n_n4196, x12753x, x12767x, x12768x, x12749x}, x12776x);
	defparam lut_10950.LUT_SIZE = 7;
	defparam lut_10950.mask = 128'h37ff37ff3fff3fff7fffffffffffffff;

	lut_sub lut_10957 ({sk[2316], i_9_, i_7_, i_8_, i_6_, x551x}, x12792x);
	defparam lut_10957.LUT_SIZE = 6;
	defparam lut_10957.mask = 64'h77ff77ff00110000;

	lut_sub lut_10960 ({sk[2317], x14x, x545x, n_n3849, x86x, n_n4694, x12792x}, x12796x);
	defparam lut_10960.LUT_SIZE = 7;
	defparam lut_10960.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_10966 ({sk[2318], x15x, x539x, x11x, x14x, x482x, x595x}, x12790x);
	defparam lut_10966.LUT_SIZE = 7;
	defparam lut_10966.mask = 128'h37ff37ff3fff3fff03570f5f57575f5f;

	lut_sub lut_10971 ({sk[2319], i_9_, i_7_, i_8_, i_6_, n_n518, n_n325}, x12791x);
	defparam lut_10971.LUT_SIZE = 7;
	defparam lut_10971.mask = 128'h37ff37ff3fff3fff0010111010000000;

	lut_sub lut_10977 ({sk[2320], x21x, x14x, x490x, x551x}, x12782x);
	defparam lut_10977.LUT_SIZE = 5;
	defparam lut_10977.mask = 32'h5f5f0357;

	lut_sub lut_10980 ({sk[2321], x25x, x22x, x14x, x517x, x595x, x551x}, x12783x);
	defparam lut_10980.LUT_SIZE = 7;
	defparam lut_10980.mask = 128'h37ff37ff3fff3fff000f555f333f777f;

	lut_sub lut_10984 ({sk[2322], x12784x, x12790x, x12791x, x12782x, x12783x}, x12797x);
	defparam lut_10984.LUT_SIZE = 6;
	defparam lut_10984.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_10990 ({sk[2323], x25x, x492x, x22x, x10x, x582x}, x12810x);
	defparam lut_10990.LUT_SIZE = 6;
	defparam lut_10990.mask = 64'h77ff77ff05375577;

	lut_sub lut_10994 ({sk[2324], i_9_, i_7_, i_8_, i_6_, n_n482, n_n390}, x12811x);
	defparam lut_10994.LUT_SIZE = 7;
	defparam lut_10994.mask = 128'h37ff37ff3fff3fff0100100010001000;

	lut_sub lut_10999 ({sk[2325], x10x, x23x, x584x, x582x, x12810x, x12811x}, x12813x);
	defparam lut_10999.LUT_SIZE = 7;
	defparam lut_10999.mask = 128'h37ff37ff3fff3fff77777f7f77ff7fff;

	lut_sub lut_11004 ({sk[2326], i_9_, i_7_, i_8_, i_6_, n_n390, n_n473}, n_n710);
	defparam lut_11004.LUT_SIZE = 7;
	defparam lut_11004.mask = 128'h37ff37ff3fff3fff0101111100001101;

	lut_sub lut_11014 ({sk[2327], i_9_, i_7_, i_8_, i_6_, x507x, x526x}, x12798x);
	defparam lut_11014.LUT_SIZE = 7;
	defparam lut_11014.mask = 128'h37ff37ff3fff3fff0035000000000000;

	lut_sub lut_11017 ({sk[2328], x426x, n_n1636, x417x, n_n710, x12798x}, x12814x);
	defparam lut_11017.LUT_SIZE = 6;
	defparam lut_11017.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_11023 ({sk[2329], i_9_, i_7_, i_8_, i_6_, n_n325, n_n500}, n_n704);
	defparam lut_11023.LUT_SIZE = 7;
	defparam lut_11023.mask = 128'h37ff37ff3fff3fff0110110110000111;

	lut_sub lut_11033 ({sk[2330], x22x, x14x, x574x, x573x, x575x}, x12822x);
	defparam lut_11033.LUT_SIZE = 6;
	defparam lut_11033.mask = 64'h77ff77ff003f557f;

	lut_sub lut_11037 ({sk[2331], n_n4205, n_n4204, x456x, n_n856, n_n704, x12822x}, x12827x);
	defparam lut_11037.LUT_SIZE = 7;
	defparam lut_11037.mask = 128'h37ff37ff3fff3fff7fffffffffffffff;

	lut_sub lut_11044 ({sk[2332], x12796x, x12797x, x12813x, x12814x, x12827x}, n_n628);
	defparam lut_11044.LUT_SIZE = 6;
	defparam lut_11044.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_11050 ({sk[2333], x18x, x490x, x20x, x512x, x535x, n_n4938}, x22210x);
	defparam lut_11050.LUT_SIZE = 7;
	defparam lut_11050.mask = 128'h37ff37ff3fff3fffaaa0aaa088800000;

	lut_sub lut_11055 ({sk[2334], x24x, x597x, n_n3805, x180x, x22210x}, x12843x);
	defparam lut_11055.LUT_SIZE = 6;
	defparam lut_11055.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_11060 ({sk[2335], i_9_, i_7_, i_8_, i_6_, x597x, x485x}, x12850x);
	defparam lut_11060.LUT_SIZE = 7;
	defparam lut_11060.mask = 128'h37ff37ff3fff3fff5300000000000000;

	lut_sub lut_11063 ({sk[2336], x18x, x597x, x20x, x563x}, x12851x);
	defparam lut_11063.LUT_SIZE = 5;
	defparam lut_11063.mask = 32'h5f5f0357;

	lut_sub lut_11066 ({sk[2337], x29x, n_n801, x12850x, x12851x}, x12857x);
	defparam lut_11066.LUT_SIZE = 5;
	defparam lut_11066.mask = 32'h5f5f7fff;

	lut_sub lut_11071 ({sk[2338], i_9_, i_7_, i_8_, i_6_, n_n509, n_n195}, x12849x);
	defparam lut_11071.LUT_SIZE = 7;
	defparam lut_11071.mask = 128'h37ff37ff3fff3fff0001001000011100;

	lut_sub lut_11077 ({sk[2339], i_9_, i_7_, i_8_, i_6_, x485x}, x12845x);
	defparam lut_11077.LUT_SIZE = 6;
	defparam lut_11077.mask = 64'h77ff77ff10400000;

	lut_sub lut_11080 ({sk[2340], i_9_, n_n195, x103x, x581x, x494x}, x12852x);
	defparam lut_11080.LUT_SIZE = 6;
	defparam lut_11080.mask = 64'h77ff77ff0f0f0f7f;

	lut_sub lut_11084 ({sk[2341], x247x, x57x, x43x, x12849x, x12845x, x12852x}, x12858x);
	defparam lut_11084.LUT_SIZE = 7;
	defparam lut_11084.mask = 128'h37ff37ff3fff3fff7fffffffffffffff;

	lut_sub lut_11091 ({sk[2342], x25x, x24x, x553x, n_n814, x22209x}, n_n689);
	defparam lut_11091.LUT_SIZE = 6;
	defparam lut_11091.mask = 64'h77ff77ffbbbfbfbf;

	lut_sub lut_11096 ({sk[2343], x20x, x23x, x553x, x411x, x342x, x341x}, x12842x);
	defparam lut_11096.LUT_SIZE = 7;
	defparam lut_11096.mask = 128'h37ff37ff3fff3fff7f7f7fff7fff7fff;

	lut_sub lut_11102 ({sk[2344], n_n691, x12724x, x12722x, x12723x, x12861x, x12862x}, x12865x);
	defparam lut_11102.LUT_SIZE = 7;
	defparam lut_11102.mask = 128'h37ff37ff3fff3fff7fffffffffffffff;

	lut_sub lut_11109 ({sk[2345], x12843x, x12857x, x12858x, n_n689, x12842x, x12865x}, x12867x);
	defparam lut_11109.LUT_SIZE = 7;
	defparam lut_11109.mask = 128'h37ff37ff3fff3fff7fffffffffffffff;

	lut_sub lut_11116 ({sk[2346], x25x, x10x, x490x, x549x, x535x, x523x}, x22194x);
	defparam lut_11116.LUT_SIZE = 7;
	defparam lut_11116.mask = 128'h37ff37ff3fff3fffffffc000aaaa8000;

	lut_sub lut_11121 ({sk[2347], x20x, x504x, x429x, x214x, x22194x}, n_n3933);
	defparam lut_11121.LUT_SIZE = 6;
	defparam lut_11121.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_11126 ({sk[2348], x25x, x15x, x11x, x561x, x571x, n_n4611}, x22193x);
	defparam lut_11126.LUT_SIZE = 7;
	defparam lut_11126.mask = 128'h37ff37ff3fff3fffaa888888a0808080;

	lut_sub lut_11131 ({sk[2349], x10x, x475x, n_n4613, x481x, x139x, x22193x}, n_n3932);
	defparam lut_11131.LUT_SIZE = 7;
	defparam lut_11131.mask = 128'h37ff37ff3fff3fffbbffbbffbfffffff;

	lut_sub lut_11137 ({sk[2350], x25x, x16x, x24x, x474x, x498x}, x14465x);
	defparam lut_11137.LUT_SIZE = 6;
	defparam lut_11137.mask = 64'h77ff77ff05375577;

	lut_sub lut_11141 ({sk[2351], x16x, x475x, x23x, x564x, x473x, n_n4365}, x22158x);
	defparam lut_11141.LUT_SIZE = 7;
	defparam lut_11141.mask = 128'h37ff37ff3fff3fffaa88aa88a0800000;

	lut_sub lut_11146 ({sk[2352], x492x, x21x, x17x, x23x, x584x, x576x}, x14738x);
	defparam lut_11146.LUT_SIZE = 7;
	defparam lut_11146.mask = 128'h37ff37ff3fff3fff0537557705ff55ff;

	lut_sub lut_11151 ({sk[2353], i_9_, i_7_, i_8_, i_6_, n_n325, n_n491}, x15766x);
	defparam lut_11151.LUT_SIZE = 7;
	defparam lut_11151.mask = 128'h37ff37ff3fff3fff0001110011111010;

	lut_sub lut_11161 ({sk[2354], i_9_, i_7_, i_8_, i_6_, x588x}, x15754x);
	defparam lut_11161.LUT_SIZE = 6;
	defparam lut_11161.mask = 64'h77ff77ff00050000;

	lut_sub lut_11164 ({sk[2355], x15x, x14x, x558x, x588x, x23x, x575x}, x15755x);
	defparam lut_11164.LUT_SIZE = 7;
	defparam lut_11164.mask = 128'h37ff37ff3fff3fff111111ff1f1f1fff;

	lut_sub lut_11168 ({sk[2356], x69x, x258x, x15756x, x15761x, x15754x, x15755x}, x15767x);
	defparam lut_11168.LUT_SIZE = 7;
	defparam lut_11168.mask = 128'h37ff37ff3fff3fff7fffffffffffffff;

	lut_sub lut_11175 ({sk[2357], x10x, x472x, x581x, x549x, x548x}, x15328x);
	defparam lut_11175.LUT_SIZE = 6;
	defparam lut_11175.mask = 64'h77ff77ff00007fff;

	lut_sub lut_11180 ({sk[2358], i_9_, i_1_, i_2_, i_0_, x477x, x482x}, x15326x);
	defparam lut_11180.LUT_SIZE = 7;
	defparam lut_11180.mask = 128'h37ff37ff3fff3fff0000000000070000;

	lut_sub lut_11183 ({sk[2359], x22x, x479x, x401x, x15328x, x15326x}, n_n2842);
	defparam lut_11183.LUT_SIZE = 6;
	defparam lut_11183.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_11188 ({sk[2360], x22x, x14x, x549x, x526x}, x15331x);
	defparam lut_11188.LUT_SIZE = 5;
	defparam lut_11188.mask = 32'h5f5f0357;

	lut_sub lut_11191 ({sk[2361], x21x, x10x, x524x, x582x, x536x, x526x}, x22107x);
	defparam lut_11191.LUT_SIZE = 7;
	defparam lut_11191.mask = 128'h37ff37ff3fff3fffffffcc00a0a08000;

	lut_sub lut_11196 ({sk[2362], x11x, x526x, x119x, x15331x, x22107x}, n_n2841);
	defparam lut_11196.LUT_SIZE = 6;
	defparam lut_11196.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_11201 ({sk[2363], x15x, x16x, x24x, x482x, x480x, x473x}, x22098x);
	defparam lut_11201.LUT_SIZE = 7;
	defparam lut_11201.mask = 128'h37ff37ff3fff3fffffaac080aaaa8080;

	lut_sub lut_11206 ({sk[2364], x25x, x16x, x501x, x24x, x545x, x497x}, x22330x);
	defparam lut_11206.LUT_SIZE = 7;
	defparam lut_11206.mask = 128'h37ff37ff3fff3ffffff0ccc0aaa08880;

	lut_sub lut_11215 ({sk[2365], i_9_, i_7_, i_8_, i_6_, x551x}, x16132x);
	defparam lut_11215.LUT_SIZE = 6;
	defparam lut_11215.mask = 64'h77ff77ff01010000;

	lut_sub lut_11218 ({sk[2366], i_9_, i_7_, i_8_, i_6_, n_n325, n_n535}, x464x);
	defparam lut_11218.LUT_SIZE = 7;
	defparam lut_11218.mask = 128'h37ff37ff3fff3fff0110000011000010;

	lut_sub lut_11224 ({sk[2367], x21x, x14x, x490x, x551x}, x16138x);
	defparam lut_11224.LUT_SIZE = 5;
	defparam lut_11224.mask = 32'h5f5f0357;

	lut_sub lut_11227 ({sk[2368], x19x, x20x, x550x, x514x, x548x, x223x}, x22311x);
	defparam lut_11227.LUT_SIZE = 7;
	defparam lut_11227.mask = 128'h37ff37ff3fff3fffaaaaa0a088008000;

	lut_sub lut_11232 ({sk[2369], x12x, n_n5181, x503x, x524x, x527x, x89x}, x22096x);
	defparam lut_11232.LUT_SIZE = 7;
	defparam lut_11232.mask = 128'h37ff37ff3fff3fffaaaa000080000000;

	lut_sub lut_11235 ({sk[2370], i_9_, i_7_, i_8_, i_6_, n_n509, n_n195}, n_n1846);
	defparam lut_11235.LUT_SIZE = 7;
	defparam lut_11235.mask = 128'h37ff37ff3fff3fff1101010001110110;

	lut_sub lut_11245 ({sk[2371], x25x, x21x, x18x, x597x, x485x, x564x}, x22331x);
	defparam lut_11245.LUT_SIZE = 7;
	defparam lut_11245.mask = 128'h37ff37ff3fff3fffffaaf0a0cc88c080;

	lut_sub lut_11254 ({sk[2372], x11x, x597x, x299x, x405x, x22331x}, x16157x);
	defparam lut_11254.LUT_SIZE = 6;
	defparam lut_11254.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_11259 ({sk[2373], i_9_, n_n195, x581x, x494x, x393x}, x16152x);
	defparam lut_11259.LUT_SIZE = 6;
	defparam lut_11259.mask = 64'h77ff77ff5555557f;

	lut_sub lut_11263 ({sk[2374], i_9_, n_n518, n_n526, n_n195, x43x}, x16153x);
	defparam lut_11263.LUT_SIZE = 6;
	defparam lut_11263.mask = 64'h77ff77ff55575557;

	lut_sub lut_11267 ({sk[2375], n_n1846, x16152x, x16153x}, x16158x);
	defparam lut_11267.LUT_SIZE = 4;
	defparam lut_11267.mask = 16'h0f7f;

	lut_sub lut_11271 ({sk[2376], i_9_, i_7_, i_8_, i_6_, n_n473, n_n260}, n_n1852);
	defparam lut_11271.LUT_SIZE = 7;
	defparam lut_11271.mask = 128'h37ff37ff3fff3fff0101010001110111;

	lut_sub lut_11281 ({sk[2377], x24x, x17x, x529x, x589x, x524x}, x22268x);
	defparam lut_11281.LUT_SIZE = 6;
	defparam lut_11281.mask = 64'h77ff77ffffa0cc80;

	lut_sub lut_11286 ({sk[2378], x20x, x512x, x138x, x22268x}, x16168x);
	defparam lut_11286.LUT_SIZE = 5;
	defparam lut_11286.mask = 32'h5f5fbbbf;

	lut_sub lut_11290 ({sk[2379], x180x, x411x, x331x, x305x, n_n1852}, x16169x);
	defparam lut_11290.LUT_SIZE = 6;
	defparam lut_11290.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_11296 ({sk[2380], i_9_, i_7_, i_8_, i_6_, n_n260, n_n464}, n_n1850);
	defparam lut_11296.LUT_SIZE = 7;
	defparam lut_11296.mask = 128'h37ff37ff3fff3fff1110101010101010;

	lut_sub lut_11306 ({sk[2381], x25x, x24x, x597x, x553x, n_n4962, x68x}, x22093x);
	defparam lut_11306.LUT_SIZE = 7;
	defparam lut_11306.mask = 128'h37ff37ff3fff3fff8888880080808000;

	lut_sub lut_11311 ({sk[2382], i_9_, i_7_, i_8_, i_6_, n_n535, n_n195}, x22336x);
	defparam lut_11311.LUT_SIZE = 7;
	defparam lut_11311.mask = 128'h37ff37ff3fff3ffffeeefeffefeefeee;

	lut_sub lut_11319 ({sk[2383], x29x, n_n1850, x22093x, x22336x}, x16180x);
	defparam lut_11319.LUT_SIZE = 5;
	defparam lut_11319.mask = 32'h5f5fefff;

	lut_sub lut_11324 ({sk[2384], x592x, x19x, x11x, x24x, x478x, x580x}, x15845x);
	defparam lut_11324.LUT_SIZE = 7;
	defparam lut_11324.mask = 128'h37ff37ff3fff3fff000077770fff7fff;

	lut_sub lut_11329 ({sk[2385], i_9_, i_7_, i_8_, i_6_, n_n325, n_n535}, x12404x);
	defparam lut_11329.LUT_SIZE = 7;
	defparam lut_11329.mask = 128'h37ff37ff3fff3fff0100010100000100;

	lut_sub lut_11334 ({sk[2386], x15x, x14x, x545x, x551x}, x12402x);
	defparam lut_11334.LUT_SIZE = 5;
	defparam lut_11334.mask = 32'h5f5f0357;

	lut_sub lut_11337 ({sk[2387], x19x, x545x, x478x, x517x, x546x}, x11698x);
	defparam lut_11337.LUT_SIZE = 6;
	defparam lut_11337.mask = 64'h77ff77ff00007fff;

	lut_sub lut_11342 ({sk[2388], x19x, x539x, x24x, x535x, x599x}, x11697x);
	defparam lut_11342.LUT_SIZE = 6;
	defparam lut_11342.mask = 64'h77ff77ff050537ff;

	lut_sub lut_11346 ({sk[2389], i_9_, i_7_, i_8_, i_6_, n_n536, n_n473}, n_n730);
	defparam lut_11346.LUT_SIZE = 7;
	defparam lut_11346.mask = 128'h37ff37ff3fff3fff0101100001111110;

	lut_sub lut_11356 ({sk[2390], x15x, x11x, x20x, x531x, n_n4952, x553x}, x22209x);
	defparam lut_11356.LUT_SIZE = 7;
	defparam lut_11356.mask = 128'h37ff37ff3fff3fffccc0888088808880;

	lut_sub lut_11361 ({sk[2391], i_9_, i_7_, i_8_, i_6_, n_n473, n_n65}, x12974x);
	defparam lut_11361.LUT_SIZE = 7;
	defparam lut_11361.mask = 128'h37ff37ff3fff3fff0100000001100010;

	lut_sub lut_11366 ({sk[2392], i_9_, i_7_, i_8_, i_6_, n_n130, n_n464}, n_n670);
	defparam lut_11366.LUT_SIZE = 7;
	defparam lut_11366.mask = 128'h37ff37ff3fff3fff1111101001011000;

	lut_sub lut_11376 ({sk[2393], i_9_, i_7_, i_8_, i_6_, n_n473, n_n130}, x12991x);
	defparam lut_11376.LUT_SIZE = 7;
	defparam lut_11376.mask = 128'h37ff37ff3fff3fff0010100010001000;

	lut_sub lut_11381 ({sk[2394], i_9_, n_n534, n_n130, x488x, n_n464, n_n1927}, x12992x);
	defparam lut_11381.LUT_SIZE = 7;
	defparam lut_11381.mask = 128'h37ff37ff3fff3fff55555555555f557f;

	lut_sub lut_11385 ({sk[2395], x515x, x15x, x12968x, x12969x, x377x, n_n632}, x12982x);
	defparam lut_11385.LUT_SIZE = 7;
	defparam lut_11385.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_11391 ({sk[2396], x12974x, x12979x, x12980x, x22206x}, x12983x);
	defparam lut_11391.LUT_SIZE = 5;
	defparam lut_11391.mask = 32'h5f5fbfff;

	lut_sub lut_11396 ({sk[2397], x25x, x12x, x514x, x493x, x107x, x22258x}, x12997x);
	defparam lut_11396.LUT_SIZE = 7;
	defparam lut_11396.mask = 128'h37ff37ff3fff3fffbbbbbfbfbbffbfff;

	lut_sub lut_11401 ({sk[2398], n_n670, x12991x, x12992x}, x12998x);
	defparam lut_11401.LUT_SIZE = 4;
	defparam lut_11401.mask = 16'h0f7f;

	lut_sub lut_11405 ({sk[2399], n_n634, x12982x, x12983x, x12997x, x12998x}, x13001x);
	defparam lut_11405.LUT_SIZE = 6;
	defparam lut_11405.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_11411 ({sk[2400], i_9_, i_7_, i_8_, i_6_, n_n482, n_n195}, x12945x);
	defparam lut_11411.LUT_SIZE = 7;
	defparam lut_11411.mask = 128'h37ff37ff3fff3fff0101111000110110;

	lut_sub lut_11421 ({sk[2401], x12881x, x12882x, x12898x, x12894x, x12895x}, x13000x);
	defparam lut_11421.LUT_SIZE = 6;
	defparam lut_11421.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_11427 ({sk[2402], i_9_, i_7_, i_8_, i_6_, n_n536, n_n500}, x14471x);
	defparam lut_11427.LUT_SIZE = 7;
	defparam lut_11427.mask = 128'h37ff37ff3fff3fff0110001000000010;

	lut_sub lut_11432 ({sk[2403], x16x, x23x, x498x, x556x}, x14469x);
	defparam lut_11432.LUT_SIZE = 5;
	defparam lut_11432.mask = 32'h5f5f0357;

	lut_sub lut_11435 ({sk[2404], x21x, x12x, x23x, x518x, x491x, x568x}, x22325x);
	defparam lut_11435.LUT_SIZE = 7;
	defparam lut_11435.mask = 128'h37ff37ff3fff3fffffaac080aaaa8080;

	lut_sub lut_11440 ({sk[2405], i_9_, n_n390, x509x, n_n491, n_n520, x587x}, x15468x);
	defparam lut_11440.LUT_SIZE = 7;
	defparam lut_11440.mask = 128'h37ff37ff3fff3fff00000303000057ff;

	lut_sub lut_11445 ({sk[2406], i_9_, n_n524, n_n260, n_n491, n_n500, n_n530}, x15348x);
	defparam lut_11445.LUT_SIZE = 7;
	defparam lut_11445.mask = 128'h37ff37ff3fff3fff0011001f0011001f;

	lut_sub lut_11450 ({sk[2407], i_9_, n_n473, n_n325, n_n520, x503x, x440x}, x16189x);
	defparam lut_11450.LUT_SIZE = 7;
	defparam lut_11450.mask = 128'h37ff37ff3fff3fff555555555577557f;

	lut_sub lut_11454 ({sk[2408], i_9_, i_7_, i_8_, i_6_, n_n473, n_n325}, x16190x);
	defparam lut_11454.LUT_SIZE = 7;
	defparam lut_11454.mask = 128'h37ff37ff3fff3fff0110100000101000;

	lut_sub lut_11460 ({sk[2409], i_9_, i_1_, i_2_, i_0_, x535x, x527x}, x16191x);
	defparam lut_11460.LUT_SIZE = 7;
	defparam lut_11460.mask = 128'h37ff37ff3fff3fff0000000005000030;

	lut_sub lut_11463 ({sk[2410], x25x, x552x, n_n4824, x388x, n_n4197, x16191x}, x16198x);
	defparam lut_11463.LUT_SIZE = 7;
	defparam lut_11463.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_11469 ({sk[2411], x22x, x17x, x552x, x23x, x517x, x530x}, x16194x);
	defparam lut_11469.LUT_SIZE = 7;
	defparam lut_11469.mask = 128'h37ff37ff3fff3fff0505373755ff77ff;

	lut_sub lut_11474 ({sk[2412], x14x, x516x, x151x, x16189x, x16190x, x16194x}, x16199x);
	defparam lut_11474.LUT_SIZE = 7;
	defparam lut_11474.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_11480 ({sk[2413], i_9_, i_7_, i_8_, i_6_, n_n518, n_n260}, x16204x);
	defparam lut_11480.LUT_SIZE = 7;
	defparam lut_11480.mask = 128'h37ff37ff3fff3fff1100000011000010;

	lut_sub lut_11486 ({sk[2414], i_9_, i_7_, i_8_, i_6_, n_n509, n_n260}, n_n1857);
	defparam lut_11486.LUT_SIZE = 7;
	defparam lut_11486.mask = 128'h37ff37ff3fff3fff0111111001001010;

	lut_sub lut_11496 ({sk[2415], i_9_, i_7_, i_8_, i_6_, x552x, x596x}, x16208x);
	defparam lut_11496.LUT_SIZE = 7;
	defparam lut_11496.mask = 128'h37ff37ff3fff3fff0000350000000000;

	lut_sub lut_11499 ({sk[2416], x25x, x17x, x596x, x546x}, x16209x);
	defparam lut_11499.LUT_SIZE = 5;
	defparam lut_11499.mask = 32'h5f5f0537;

	lut_sub lut_11502 ({sk[2417], x17x, x490x, x177x, x176x, x16208x, x16209x}, x16213x);
	defparam lut_11502.LUT_SIZE = 7;
	defparam lut_11502.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_11508 ({sk[2418], x25x, x17x, x484x, x481x}, x16200x);
	defparam lut_11508.LUT_SIZE = 5;
	defparam lut_11508.mask = 32'h5f5f0537;

	lut_sub lut_11511 ({sk[2419], x375x, x16204x, n_n1857, x16200x}, x16214x);
	defparam lut_11511.LUT_SIZE = 5;
	defparam lut_11511.mask = 32'h5f5f7fff;

	lut_sub lut_11516 ({sk[2420], i_9_, i_7_, i_8_, i_6_, n_n260, n_n500}, x16217x);
	defparam lut_11516.LUT_SIZE = 7;
	defparam lut_11516.mask = 128'h37ff37ff3fff3fff0100001001001000;

	lut_sub lut_11521 ({sk[2421], x24x, x17x, x560x, x576x, n_n1985, x16220x}, x16222x);
	defparam lut_11521.LUT_SIZE = 7;
	defparam lut_11521.mask = 128'h37ff37ff3fff3fff777777ff7f7f7fff;

	lut_sub lut_11526 ({sk[2422], x461x, x16184x, x16185x, x16217x, x16216x}, x16223x);
	defparam lut_11526.LUT_SIZE = 6;
	defparam lut_11526.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_11532 ({sk[2423], x22x, x21x, x11x, x10x, x542x, x559x}, x15823x);
	defparam lut_11532.LUT_SIZE = 7;
	defparam lut_11532.mask = 128'h37ff37ff3fff3fff0537373737373737;

	lut_sub lut_11537 ({sk[2424], x13x, x570x, x529x, n_n4572, x46x, x15823x}, n_n1727);
	defparam lut_11537.LUT_SIZE = 7;
	defparam lut_11537.mask = 128'h37ff37ff3fff3fff7f7f7f7f7fffffff;

	lut_sub lut_11543 ({sk[2425], x22x, x10x, x571x, x587x}, x15825x);
	defparam lut_11543.LUT_SIZE = 5;
	defparam lut_11543.mask = 32'h5f5f0537;

	lut_sub lut_11546 ({sk[2426], x10x, x24x, x556x, x582x}, x15826x);
	defparam lut_11546.LUT_SIZE = 5;
	defparam lut_11546.mask = 32'h5f5f0537;

	lut_sub lut_11549 ({sk[2427], x21x, x10x, x561x, x562x}, x15827x);
	defparam lut_11549.LUT_SIZE = 5;
	defparam lut_11549.mask = 32'h5f5f0537;

	lut_sub lut_11552 ({sk[2428], x23x, x561x, x255x, x15825x, x15826x, x15827x}, n_n1726);
	defparam lut_11552.LUT_SIZE = 7;
	defparam lut_11552.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_11558 ({sk[2429], x17x, x20x, x472x, x480x, x530x, x593x}, x15852x);
	defparam lut_11558.LUT_SIZE = 7;
	defparam lut_11558.mask = 128'h37ff37ff3fff3fff000033335fff7fff;

	lut_sub lut_11563 ({sk[2430], x15x, x22x, x14x, x580x, x596x, x530x}, x15851x);
	defparam lut_11563.LUT_SIZE = 7;
	defparam lut_11563.mask = 128'h37ff37ff3fff3fff000f333f555f777f;

	lut_sub lut_11567 ({sk[2431], i_9_, i_7_, i_8_, i_6_, n_n509, n_n195}, x15864x);
	defparam lut_11567.LUT_SIZE = 7;
	defparam lut_11567.mask = 128'h37ff37ff3fff3fff0010101000001000;

	lut_sub lut_11572 ({sk[2432], x22x, x521x, x18x, x567x}, x15862x);
	defparam lut_11572.LUT_SIZE = 5;
	defparam lut_11572.mask = 32'h5f5f0357;

	lut_sub lut_11575 ({sk[2433], i_9_, i_7_, i_8_, i_6_, x590x, x513x}, x15883x);
	defparam lut_11575.LUT_SIZE = 7;
	defparam lut_11575.mask = 128'h37ff37ff3fff3fff5000000300000000;

	lut_sub lut_11578 ({sk[2434], x21x, x18x, x557x, x580x, x573x, x513x}, x15885x);
	defparam lut_11578.LUT_SIZE = 7;
	defparam lut_11578.mask = 128'h37ff37ff3fff3fff00003fff55557fff;

	lut_sub lut_11583 ({sk[2435], i_9_, i_7_, i_8_, i_6_, x599x, x555x}, x15891x);
	defparam lut_11583.LUT_SIZE = 7;
	defparam lut_11583.mask = 128'h37ff37ff3fff3fff0053000000000000;

	lut_sub lut_11586 ({sk[2436], x19x, x21x, x12x, x522x, x546x, x533x}, x15893x);
	defparam lut_11586.LUT_SIZE = 7;
	defparam lut_11586.mask = 128'h37ff37ff3fff3fff000f555f333f777f;

	lut_sub lut_11590 ({sk[2437], x19x, x545x, x23x, x517x, x533x}, x22320x);
	defparam lut_11590.LUT_SIZE = 6;
	defparam lut_11590.mask = 64'h77ff77fffafac800;

	lut_sub lut_11595 ({sk[2438], x12x, x505x, x502x, x525x, x493x}, x11705x);
	defparam lut_11595.LUT_SIZE = 6;
	defparam lut_11595.mask = 64'h77ff77ff00007fff;

	lut_sub lut_11600 ({sk[2439], i_9_, i_7_, i_8_, i_6_, n_n536, n_n535}, n_n738);
	defparam lut_11600.LUT_SIZE = 7;
	defparam lut_11600.mask = 128'h37ff37ff3fff3fff0101001101011101;

	lut_sub lut_11610 ({sk[2440], i_9_, i_7_, i_8_, i_6_, n_n455, n_n491}, n_n722);
	defparam lut_11610.LUT_SIZE = 7;
	defparam lut_11610.mask = 128'h37ff37ff3fff3fff0101111001111000;

	lut_sub lut_11620 ({sk[2441], x13x, x23x, x574x, x541x}, x346x);
	defparam lut_11620.LUT_SIZE = 5;
	defparam lut_11620.mask = 32'h5f5f0537;

	lut_sub lut_11623 ({sk[2442], x15x, x13x, x586x, x543x}, x13032x);
	defparam lut_11623.LUT_SIZE = 5;
	defparam lut_11623.mask = 32'h5f5f0357;

	lut_sub lut_11626 ({sk[2443], i_9_, i_7_, i_8_, i_6_, x542x, x541x}, x13033x);
	defparam lut_11626.LUT_SIZE = 7;
	defparam lut_11626.mask = 128'h37ff37ff3fff3fff0000500300000000;

	lut_sub lut_11629 ({sk[2444], x13x, x570x, x307x, n_n897, x13032x, x13033x}, x13039x);
	defparam lut_11629.LUT_SIZE = 7;
	defparam lut_11629.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_11635 ({sk[2445], x25x, x13x, x584x, x543x}, x13031x);
	defparam lut_11635.LUT_SIZE = 5;
	defparam lut_11635.mask = 32'h5f5f0357;

	lut_sub lut_11638 ({sk[2446], x378x, x162x, n_n722, x346x, x13031x}, x13040x);
	defparam lut_11638.LUT_SIZE = 6;
	defparam lut_11638.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_11644 ({sk[2447], x13x, x23x, x562x, x476x}, x13023x);
	defparam lut_11644.LUT_SIZE = 5;
	defparam lut_11644.mask = 32'h5f5f0537;

	lut_sub lut_11647 ({sk[2448], x13x, x11x, x478x, x556x, x541x}, x13024x);
	defparam lut_11647.LUT_SIZE = 6;
	defparam lut_11647.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_11651 ({sk[2449], i_9_, i_7_, i_8_, i_6_, n_n518, n_n455}, x13044x);
	defparam lut_11651.LUT_SIZE = 7;
	defparam lut_11651.mask = 128'h37ff37ff3fff3fff0110110101101001;

	lut_sub lut_11661 ({sk[2450], x13020x, x13021x, x13025x, x13023x, x13024x, x13044x}, x13046x);
	defparam lut_11661.LUT_SIZE = 7;
	defparam lut_11661.mask = 128'h37ff37ff3fff3fff7fffffffffffffff;

	lut_sub lut_11668 ({sk[2451], i_9_, i_7_, i_8_, i_6_, n_n473, n_n260}, n_n3691);
	defparam lut_11668.LUT_SIZE = 7;
	defparam lut_11668.mask = 128'h37ff37ff3fff3fff1101101011100010;

	lut_sub lut_11678 ({sk[2452], i_9_, x492x, n_n528, n_n491, n_n130, x20x}, x14598x);
	defparam lut_11678.LUT_SIZE = 7;
	defparam lut_11678.mask = 128'h37ff37ff3fff3fff0103010301033333;

	lut_sub lut_11683 ({sk[2453], x21x, x570x, x519x, x12x, x23x, x578x}, x22301x);
	defparam lut_11683.LUT_SIZE = 7;
	defparam lut_11683.mask = 128'h37ff37ff3fff3fffeee0e0e0aaa0a0a0;

	lut_sub lut_11688 ({sk[2454], i_9_, n_n534, n_n491, n_n65, x438x}, x14545x);
	defparam lut_11688.LUT_SIZE = 6;
	defparam lut_11688.mask = 64'h77ff77ff55575557;

	lut_sub lut_11692 ({sk[2455], x16x, x20x, x497x, x549x, x594x}, x15521x);
	defparam lut_11692.LUT_SIZE = 6;
	defparam lut_11692.mask = 64'h77ff77ff000f777f;

	lut_sub lut_11696 ({sk[2456], i_9_, i_7_, i_8_, i_6_, n_n536, n_n535}, x15522x);
	defparam lut_11696.LUT_SIZE = 7;
	defparam lut_11696.mask = 128'h37ff37ff3fff3fff0001101011001000;

	lut_sub lut_11703 ({sk[2457], i_9_, i_7_, i_8_, i_6_, n_n536, n_n518}, x15527x);
	defparam lut_11703.LUT_SIZE = 7;
	defparam lut_11703.mask = 128'h37ff37ff3fff3fff0001111101011010;

	lut_sub lut_11713 ({sk[2458], i_9_, i_7_, i_8_, i_6_, n_n390, n_n473}, x15770x);
	defparam lut_11713.LUT_SIZE = 7;
	defparam lut_11713.mask = 128'h37ff37ff3fff3fff0110100000000010;

	lut_sub lut_11718 ({sk[2459], i_9_, i_7_, i_8_, i_6_, n_n325, n_n535}, x15778x);
	defparam lut_11718.LUT_SIZE = 7;
	defparam lut_11718.mask = 128'h37ff37ff3fff3fff0110110111101011;

	lut_sub lut_11730 ({sk[2460], x10x, x20x, x516x, x522x, x526x}, x15774x);
	defparam lut_11730.LUT_SIZE = 6;
	defparam lut_11730.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_11734 ({sk[2461], x25x, x10x, x506x, x502x, x526x, x426x}, x22122x);
	defparam lut_11734.LUT_SIZE = 7;
	defparam lut_11734.mask = 128'h37ff37ff3fff3fffaaaaa00088888000;

	lut_sub lut_11739 ({sk[2462], x15x, x14x, x23x, x594x, x526x, n_n4694}, x22338x);
	defparam lut_11739.LUT_SIZE = 7;
	defparam lut_11739.mask = 128'h37ff37ff3fff3fffaa88a08088888080;

	lut_sub lut_11744 ({sk[2463], x15770x, x15774x, x22122x, x22338x}, x15779x);
	defparam lut_11744.LUT_SIZE = 5;
	defparam lut_11744.mask = 32'h5f5fefff;

	lut_sub lut_11749 ({sk[2464], x22x, x11x, x17x, x484x, x564x}, x15411x);
	defparam lut_11749.LUT_SIZE = 6;
	defparam lut_11749.mask = 64'h77ff77ff05373737;

	lut_sub lut_11753 ({sk[2465], x22x, x17x, x23x, x581x, x530x, n_n4843}, x22265x);
	defparam lut_11753.LUT_SIZE = 7;
	defparam lut_11753.mask = 128'h37ff37ff3fff3fffaa88a08088888080;

	lut_sub lut_11758 ({sk[2466], x17x, x549x, x494x, x15411x, x22265x}, n_n2838);
	defparam lut_11758.LUT_SIZE = 6;
	defparam lut_11758.mask = 64'h77ff77ffbbbbbfff;

	lut_sub lut_11763 ({sk[2467], i_9_, i_1_, i_2_, i_0_, x517x, x527x}, x15365x);
	defparam lut_11763.LUT_SIZE = 7;
	defparam lut_11763.mask = 128'h37ff37ff3fff3fff0000000000305000;

	lut_sub lut_11766 ({sk[2468], x15x, x12x, x490x, x548x, x532x, n_n5078}, x22115x);
	defparam lut_11766.LUT_SIZE = 7;
	defparam lut_11766.mask = 128'h37ff37ff3fff3fffaaaaa00088888000;

	lut_sub lut_11771 ({sk[2469], i_9_, x22x, n_n482, n_n130, n_n530, x555x}, x15373x);
	defparam lut_11771.LUT_SIZE = 7;
	defparam lut_11771.mask = 128'h37ff37ff3fff3fff0003555700035557;

	lut_sub lut_11775 ({sk[2470], x538x, x19x, x21x, x12x, x599x, x559x}, x22277x);
	defparam lut_11775.LUT_SIZE = 7;
	defparam lut_11775.mask = 128'h37ff37ff3fff3fffffccaa88f0c0a080;

	lut_sub lut_11784 ({sk[2471], x22x, x591x, x107x, x15373x, x22277x}, n_n2831);
	defparam lut_11784.LUT_SIZE = 6;
	defparam lut_11784.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_11789 ({sk[2472], x19x, x11x, x478x, x534x}, x15378x);
	defparam lut_11789.LUT_SIZE = 5;
	defparam lut_11789.mask = 32'h5f5f0537;

	lut_sub lut_11792 ({sk[2473], x515x, x19x, x23x, x557x}, x15379x);
	defparam lut_11792.LUT_SIZE = 5;
	defparam lut_11792.mask = 32'h5f5f0537;

	lut_sub lut_11795 ({sk[2474], x538x, x19x, x519x, x520x}, x15380x);
	defparam lut_11795.LUT_SIZE = 5;
	defparam lut_11795.mask = 32'h5f5f070f;

	lut_sub lut_11799 ({sk[2475], x25x, x15x, x22x, x534x, n_n5302, x579x}, x22117x);
	defparam lut_11799.LUT_SIZE = 7;
	defparam lut_11799.mask = 128'h37ff37ff3fff3fffccc0c0c088808080;

	lut_sub lut_11804 ({sk[2476], x386x, x15378x, x15379x, x15380x, x22117x}, x15385x);
	defparam lut_11804.LUT_SIZE = 6;
	defparam lut_11804.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_11810 ({sk[2477], x21x, x18x, x490x, x23x, x553x, x559x}, x15390x);
	defparam lut_11810.LUT_SIZE = 7;
	defparam lut_11810.mask = 128'h37ff37ff3fff3fff030357ff333377ff;

	lut_sub lut_11815 ({sk[2478], i_9_, n_n536, n_n534, x503x, n_n464, x524x}, x16094x);
	defparam lut_11815.LUT_SIZE = 7;
	defparam lut_11815.mask = 128'h37ff37ff3fff3fff0000003300005f7f;

	lut_sub lut_11820 ({sk[2479], i_9_, i_7_, i_8_, i_6_, n_n536, n_n473}, x16095x);
	defparam lut_11820.LUT_SIZE = 7;
	defparam lut_11820.mask = 128'h37ff37ff3fff3fff1010000011001000;

	lut_sub lut_11826 ({sk[2480], x538x, x16x, x21x, x500x}, x16101x);
	defparam lut_11826.LUT_SIZE = 5;
	defparam lut_11826.mask = 32'h5f5f111f;

	lut_sub lut_11829 ({sk[2481], x16x, x500x, x24x, x20x, x580x, x495x}, x16102x);
	defparam lut_11829.LUT_SIZE = 7;
	defparam lut_11829.mask = 128'h37ff37ff3fff3fff00550f5f33773f7f;

	lut_sub lut_11833 ({sk[2482], x16x, x23x, x499x, x584x}, x16097x);
	defparam lut_11833.LUT_SIZE = 5;
	defparam lut_11833.mask = 32'h5f5f0357;

	lut_sub lut_11836 ({sk[2483], x25x, x492x, x16x, x500x, x11x, x359x}, x22097x);
	defparam lut_11836.LUT_SIZE = 7;
	defparam lut_11836.mask = 128'h37ff37ff3fff3fffa8a8a800a0a0a000;

	lut_sub lut_11841 ({sk[2484], x510x, x14x, x588x, x23x, x508x, x505x}, x16228x);
	defparam lut_11841.LUT_SIZE = 7;
	defparam lut_11841.mask = 128'h37ff37ff3fff3fff000f777f000fffff;

	lut_sub lut_11846 ({sk[2485], i_9_, i_7_, i_8_, i_6_, n_n325, n_n491}, x16234x);
	defparam lut_11846.LUT_SIZE = 7;
	defparam lut_11846.mask = 128'h37ff37ff3fff3fff0001010100010100;

	lut_sub lut_11852 ({sk[2486], i_9_, i_7_, i_8_, i_6_, x483x, x595x}, x12406x);
	defparam lut_11852.LUT_SIZE = 7;
	defparam lut_11852.mask = 128'h37ff37ff3fff3fff5000000300000000;

	lut_sub lut_11855 ({sk[2487], x521x, x539x, x11x, x14x, x481x, x595x}, x22223x);
	defparam lut_11855.LUT_SIZE = 7;
	defparam lut_11855.mask = 128'h37ff37ff3fff3ffffca8f0a0f0a0f0a0;

	lut_sub lut_11860 ({sk[2488], x25x, x21x, x23x, x591x, x486x, x578x}, x11712x);
	defparam lut_11860.LUT_SIZE = 7;
	defparam lut_11860.mask = 128'h37ff37ff3fff3fff003355773f3f7f7f;

	lut_sub lut_11865 ({sk[2489], x22x, x16x, x501x, x539x, x11x}, x448x);
	defparam lut_11865.LUT_SIZE = 6;
	defparam lut_11865.mask = 64'h77ff77ff05370f3f;

	lut_sub lut_11869 ({sk[2490], i_9_, i_7_, i_8_, i_6_, n_n455, n_n473}, n_n719);
	defparam lut_11869.LUT_SIZE = 7;
	defparam lut_11869.mask = 128'h37ff37ff3fff3fff1001101011101010;

	lut_sub lut_11879 ({sk[2491], i_9_, i_7_, i_8_, i_6_, n_n536, n_n509}, n_n735);
	defparam lut_11879.LUT_SIZE = 7;
	defparam lut_11879.mask = 128'h37ff37ff3fff3fff1111100010101010;

	lut_sub lut_11889 ({sk[2492], x25x, x16x, x518x, x498x}, x13061x);
	defparam lut_11889.LUT_SIZE = 5;
	defparam lut_11889.mask = 32'h5f5f0357;

	lut_sub lut_11892 ({sk[2493], i_9_, i_7_, i_8_, i_6_, n_n536, n_n500}, x22203x);
	defparam lut_11892.LUT_SIZE = 7;
	defparam lut_11892.mask = 128'h37ff37ff3fff3ffffeeeffefeefefeee;

	lut_sub lut_11900 ({sk[2494], n_n3176, x27x, n_n735, x13061x, x22203x}, n_n657);
	defparam lut_11900.LUT_SIZE = 6;
	defparam lut_11900.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_11906 ({sk[2495], i_9_, i_7_, i_8_, i_6_, n_n536, n_n482}, x13079x);
	defparam lut_11906.LUT_SIZE = 7;
	defparam lut_11906.mask = 128'h37ff37ff3fff3fff1010001000001010;

	lut_sub lut_11912 ({sk[2496], x16x, x510x, x580x, x359x, x13079x}, x13080x);
	defparam lut_11912.LUT_SIZE = 6;
	defparam lut_11912.mask = 64'h77ff77ff77777fff;

	lut_sub lut_11917 ({sk[2497], x25x, x16x, x500x, x24x, x519x, x584x}, x22201x);
	defparam lut_11917.LUT_SIZE = 7;
	defparam lut_11917.mask = 128'h37ff37ff3fff3ffffff08880ff008800;

	lut_sub lut_11922 ({sk[2498], x492x, x16x, x11x, x586x, x499x, x285x}, x22202x);
	defparam lut_11922.LUT_SIZE = 7;
	defparam lut_11922.mask = 128'h37ff37ff3fff3fffaa88a080aa880000;

	lut_sub lut_11927 ({sk[2499], n_n730, x22201x, x22202x}, x13081x);
	defparam lut_11927.LUT_SIZE = 4;
	defparam lut_11927.mask = 16'h0fef;

	lut_sub lut_11931 ({sk[2500], x16x, x480x, x156x, x337x, x124x, x13082x}, x13086x);
	defparam lut_11931.LUT_SIZE = 7;
	defparam lut_11931.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_11937 ({sk[2501], x443x, n_n738, x448x, x13051x, x13052x}, x13087x);
	defparam lut_11937.LUT_SIZE = 6;
	defparam lut_11937.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_11943 ({sk[2502], i_9_, i_7_, i_8_, i_6_, n_n390, n_n535}, x13108x);
	defparam lut_11943.LUT_SIZE = 7;
	defparam lut_11943.mask = 128'h37ff37ff3fff3fff0000010011100000;

	lut_sub lut_11948 ({sk[2503], x13x, x525x, n_n881, x121x, x13108x}, x13111x);
	defparam lut_11948.LUT_SIZE = 6;
	defparam lut_11948.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_11953 ({sk[2504], x22x, x521x, x10x, x482x, x581x, x583x}, x13101x);
	defparam lut_11953.LUT_SIZE = 7;
	defparam lut_11953.mask = 128'h37ff37ff3fff3fff003f00ff557f55ff;

	lut_sub lut_11958 ({sk[2505], x21x, x10x, x23x, x583x, x494x}, x13100x);
	defparam lut_11958.LUT_SIZE = 6;
	defparam lut_11958.mask = 64'h77ff77ff03573377;

	lut_sub lut_11962 ({sk[2506], x15x, x11x, x583x, x547x, n_n4603, x100x}, x22200x);
	defparam lut_11962.LUT_SIZE = 7;
	defparam lut_11962.mask = 128'h37ff37ff3fff3fff8888800080808000;

	lut_sub lut_11966 ({sk[2507], x99x, x222x, x13101x, x13100x, x22200x}, x13112x);
	defparam lut_11966.LUT_SIZE = 6;
	defparam lut_11966.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_11972 ({sk[2508], x25x, x10x, x561x, x491x, x573x, x537x}, x13120x);
	defparam lut_11972.LUT_SIZE = 7;
	defparam lut_11972.mask = 128'h37ff37ff3fff3fff00007f7f00ff7fff;

	lut_sub lut_11977 ({sk[2509], x10x, x574x, x348x, n_n3861, x13120x}, x13123x);
	defparam lut_11977.LUT_SIZE = 6;
	defparam lut_11977.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_11982 ({sk[2510], i_9_, i_7_, i_8_, i_6_, n_n390, n_n509}, n_n714);
	defparam lut_11982.LUT_SIZE = 7;
	defparam lut_11982.mask = 128'h37ff37ff3fff3fff1111001011101000;

	lut_sub lut_11992 ({sk[2511], i_9_, i_7_, i_8_, i_6_, n_n390, n_n500}, x13119x);
	defparam lut_11992.LUT_SIZE = 7;
	defparam lut_11992.mask = 128'h37ff37ff3fff3fff0010010010000001;

	lut_sub lut_11997 ({sk[2512], x22x, x21x, x561x, x271x, n_n714, x13119x}, x13124x);
	defparam lut_11997.LUT_SIZE = 7;
	defparam lut_11997.mask = 128'h37ff37ff3fff3fff7f7f7fff7fff7fff;

	lut_sub lut_12003 ({sk[2513], x22x, x13x, x520x, x493x, x543x, x523x}, x13127x);
	defparam lut_12003.LUT_SIZE = 7;
	defparam lut_12003.mask = 128'h37ff37ff3fff3fff00000fff77777fff;

	lut_sub lut_12008 ({sk[2514], i_7_, i_8_, i_6_, x13x, n_n464, n_n889}, x13128x);
	defparam lut_12008.LUT_SIZE = 7;
	defparam lut_12008.mask = 128'h37ff37ff3fff3fff5557555755555555;

	lut_sub lut_12012 ({sk[2515], i_9_, i_7_, i_8_, i_6_, n_n455, n_n464}, x13129x);
	defparam lut_12012.LUT_SIZE = 7;
	defparam lut_12012.mask = 128'h37ff37ff3fff3fff0000100100101101;

	lut_sub lut_12019 ({sk[2516], n_n3875, n_n719, x13127x, x13128x, x13129x}, x13133x);
	defparam lut_12019.LUT_SIZE = 6;
	defparam lut_12019.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_12025 ({sk[2517], x10x, x570x, x508x, x505x, x506x}, x14323x);
	defparam lut_12025.LUT_SIZE = 6;
	defparam lut_12025.mask = 64'h77ff77ff00007fff;

	lut_sub lut_12030 ({sk[2518], x25x, x10x, x507x, x493x}, x14321x);
	defparam lut_12030.LUT_SIZE = 5;
	defparam lut_12030.mask = 32'h5f5f0537;

	lut_sub lut_12033 ({sk[2519], x11x, x526x, x312x, x14323x, x14321x}, n_n3561);
	defparam lut_12033.LUT_SIZE = 6;
	defparam lut_12033.mask = 64'h77ff77ff7f7f7fff;

	lut_sub lut_12038 ({sk[2520], i_9_, i_7_, i_8_, i_6_, n_n491, n_n65}, n_n2939);
	defparam lut_12038.LUT_SIZE = 7;
	defparam lut_12038.mask = 128'h37ff37ff3fff3fff0100111000110111;

	lut_sub lut_12048 ({sk[2521], x10x, x545x, n_n4573, n_n3870, x276x, x222x}, n_n2993);
	defparam lut_12048.LUT_SIZE = 7;
	defparam lut_12048.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_12054 ({sk[2522], i_9_, n_n390, n_n535, n_n520, x594x, x237x}, x15478x);
	defparam lut_12054.LUT_SIZE = 7;
	defparam lut_12054.mask = 128'h37ff37ff3fff3fff5555555f55557777;

	lut_sub lut_12058 ({sk[2523], x25x, x15x, x10x, x583x, x585x}, x15477x);
	defparam lut_12058.LUT_SIZE = 6;
	defparam lut_12058.mask = 64'h77ff77ff05373737;

	lut_sub lut_12062 ({sk[2524], x10x, x24x, x490x, x583x, x15478x, x15477x}, n_n2992);
	defparam lut_12062.LUT_SIZE = 7;
	defparam lut_12062.mask = 128'h37ff37ff3fff3fff77777f7f77ff7fff;

	lut_sub lut_12067 ({sk[2525], x18x, x485x, x472x, x23x, x564x, x562x}, x15711x);
	defparam lut_12067.LUT_SIZE = 7;
	defparam lut_12067.mask = 128'h37ff37ff3fff3fff00000f0f77ff7fff;

	lut_sub lut_12072 ({sk[2526], x24x, x474x, x18x, x567x, x405x, x15711x}, x15714x);
	defparam lut_12072.LUT_SIZE = 7;
	defparam lut_12072.mask = 128'h37ff37ff3fff3fff777777ff7f7f7fff;

	lut_sub lut_12077 ({sk[2527], i_9_, n_n526, n_n195, x485x, x475x, x394x}, x15710x);
	defparam lut_12077.LUT_SIZE = 7;
	defparam lut_12077.mask = 128'h37ff37ff3fff3fff55555f5f55775577;

	lut_sub lut_12081 ({sk[2528], x25x, x18x, x557x, x577x, x573x, x135x}, x22123x);
	defparam lut_12081.LUT_SIZE = 7;
	defparam lut_12081.mask = 128'h37ff37ff3fff3fffaaaa8800a0a08000;

	lut_sub lut_12086 ({sk[2529], x15704x, x136x, x247x, x15710x, x22123x}, x15715x);
	defparam lut_12086.LUT_SIZE = 6;
	defparam lut_12086.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_12092 ({sk[2530], x25x, x23x, x598x, x486x, x568x}, x15354x);
	defparam lut_12092.LUT_SIZE = 6;
	defparam lut_12092.mask = 64'h77ff77ff005f337f;

	lut_sub lut_12096 ({sk[2531], x25x, x12x, x475x, x591x, x491x, x574x}, x22114x);
	defparam lut_12096.LUT_SIZE = 7;
	defparam lut_12096.mask = 128'h37ff37ff3fff3fffffff8800f0f08000;

	lut_sub lut_12101 ({sk[2532], x21x, x18x, x477x, x577x}, x15357x);
	defparam lut_12101.LUT_SIZE = 5;
	defparam lut_12101.mask = 32'h5f5f0357;

	lut_sub lut_12104 ({sk[2533], x15x, x510x, x18x, x513x}, x15358x);
	defparam lut_12104.LUT_SIZE = 5;
	defparam lut_12104.mask = 32'h5f5f0357;

	lut_sub lut_12107 ({sk[2534], i_9_, i_7_, i_8_, i_6_, x485x, x590x}, x15359x);
	defparam lut_12107.LUT_SIZE = 7;
	defparam lut_12107.mask = 128'h37ff37ff3fff3fff0003000500000000;

	lut_sub lut_12110 ({sk[2535], i_9_, i_7_, i_8_, i_6_, n_n482, n_n130}, x15283x);
	defparam lut_12110.LUT_SIZE = 7;
	defparam lut_12110.mask = 128'h37ff37ff3fff3fff0100000001010100;

	lut_sub lut_12115 ({sk[2536], i_9_, n_n518, n_n390, n_n534, x490x, n_n2401}, x16031x);
	defparam lut_12115.LUT_SIZE = 7;
	defparam lut_12115.mask = 128'h37ff37ff3fff3fff555555555577557f;

	lut_sub lut_12119 ({sk[2537], i_9_, i_7_, i_8_, i_6_, n_n325, n_n535}, x11875x);
	defparam lut_12119.LUT_SIZE = 7;
	defparam lut_12119.mask = 128'h37ff37ff3fff3fff0010111101010110;

	lut_sub lut_12129 ({sk[2538], x14x, x23x, x594x, x551x}, x11864x);
	defparam lut_12129.LUT_SIZE = 5;
	defparam lut_12129.mask = 32'h5f5f0537;

	lut_sub lut_12132 ({sk[2539], x86x, x219x, x11863x, x173x, x11868x, x11864x}, x11876x);
	defparam lut_12132.LUT_SIZE = 7;
	defparam lut_12132.mask = 128'h37ff37ff3fff3fff7fffffffffffffff;

	lut_sub lut_12139 ({sk[2540], i_9_, i_1_, i_2_, i_0_, x521x, x524x}, x11716x);
	defparam lut_12139.LUT_SIZE = 7;
	defparam lut_12139.mask = 128'h37ff37ff3fff3fff0000000000305000;

	lut_sub lut_12142 ({sk[2541], i_9_, i_7_, i_8_, i_6_, x513x, x532x}, x11717x);
	defparam lut_12142.LUT_SIZE = 7;
	defparam lut_12142.mask = 128'h37ff37ff3fff3fff3000500000000000;

	lut_sub lut_12145 ({sk[2542], x18x, x20x, x554x, x505x, x527x}, x11718x);
	defparam lut_12145.LUT_SIZE = 6;
	defparam lut_12145.mask = 64'h77ff77ff000f777f;

	lut_sub lut_12149 ({sk[2543], x22x, x11x, x18x, x517x, x553x}, x14754x);
	defparam lut_12149.LUT_SIZE = 6;
	defparam lut_12149.mask = 64'h77ff77ff03575757;

	lut_sub lut_12153 ({sk[2544], i_9_, i_7_, i_8_, i_6_, n_n536, n_n535}, n_n3740);
	defparam lut_12153.LUT_SIZE = 7;
	defparam lut_12153.mask = 128'h37ff37ff3fff3fff1010110100011011;

	lut_sub lut_12163 ({sk[2545], i_9_, n_n536, n_n518, n_n530, x156x}, x14484x);
	defparam lut_12163.LUT_SIZE = 6;
	defparam lut_12163.mask = 64'h77ff77ff55575557;

	lut_sub lut_12167 ({sk[2546], i_9_, n_n536, x24x, n_n534, n_n509, x337x}, x14485x);
	defparam lut_12167.LUT_SIZE = 7;
	defparam lut_12167.mask = 128'h37ff37ff3fff3fff5555557755555777;

	lut_sub lut_12171 ({sk[2547], i_9_, i_7_, i_8_, i_6_, n_n536, n_n518}, x14487x);
	defparam lut_12171.LUT_SIZE = 7;
	defparam lut_12171.mask = 128'h37ff37ff3fff3fff0000111000100101;

	lut_sub lut_12178 ({sk[2548], x15x, x16x, x11x, x473x, x559x, n_n4341}, x22157x);
	defparam lut_12178.LUT_SIZE = 7;
	defparam lut_12178.mask = 128'h37ff37ff3fff3fffaaa08880a0a08080;

	lut_sub lut_12183 ({sk[2549], i_9_, i_7_, i_8_, i_6_, n_n500, n_n65}, n_n2940);
	defparam lut_12183.LUT_SIZE = 7;
	defparam lut_12183.mask = 128'h37ff37ff3fff3fff1110101010101010;

	lut_sub lut_12193 ({sk[2550], i_9_, i_7_, i_8_, i_6_, n_n390, n_n500}, x15492x);
	defparam lut_12193.LUT_SIZE = 7;
	defparam lut_12193.mask = 128'h37ff37ff3fff3fff0010101000100000;

	lut_sub lut_12198 ({sk[2551], i_9_, i_7_, i_8_, i_6_, x597x, x485x}, x15716x);
	defparam lut_12198.LUT_SIZE = 7;
	defparam lut_12198.mask = 128'h37ff37ff3fff3fff0530000000000000;

	lut_sub lut_12201 ({sk[2552], x25x, x485x, x57x, x251x, x133x, x15716x}, n_n2962);
	defparam lut_12201.LUT_SIZE = 7;
	defparam lut_12201.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_12207 ({sk[2553], i_9_, n_n520, n_n130, n_n500, x407x}, x15287x);
	defparam lut_12207.LUT_SIZE = 6;
	defparam lut_12207.mask = 64'h77ff77ff55575557;

	lut_sub lut_12211 ({sk[2554], i_9_, i_7_, i_8_, i_6_, n_n491, n_n130}, x15288x);
	defparam lut_12211.LUT_SIZE = 7;
	defparam lut_12211.mask = 128'h37ff37ff3fff3fff0001101100000010;

	lut_sub lut_12217 ({sk[2555], i_9_, i_7_, i_8_, i_6_, x577x, x513x}, x11722x);
	defparam lut_12217.LUT_SIZE = 7;
	defparam lut_12217.mask = 128'h37ff37ff3fff3fff0000003500000000;

	lut_sub lut_12220 ({sk[2556], i_9_, i_7_, i_8_, i_6_, x590x, x513x}, x11723x);
	defparam lut_12220.LUT_SIZE = 7;
	defparam lut_12220.mask = 128'h37ff37ff3fff3fff3000050000000000;

	lut_sub lut_12223 ({sk[2557], x538x, x18x, x485x, x23x, x537x}, x11725x);
	defparam lut_12223.LUT_SIZE = 6;
	defparam lut_12223.mask = 64'h77ff77ff035703ff;

	lut_sub lut_12227 ({sk[2558], i_9_, i_7_, i_8_, i_6_, n_n130, n_n464}, n_n3670);
	defparam lut_12227.LUT_SIZE = 7;
	defparam lut_12227.mask = 128'h37ff37ff3fff3fff0100001101011111;

	lut_sub lut_12237 ({sk[2559], i_9_, i_7_, i_8_, i_6_, n_n536, n_n464}, n_n3004);
	defparam lut_12237.LUT_SIZE = 7;
	defparam lut_12237.mask = 128'h37ff37ff3fff3fff0001011111001110;

	lut_sub lut_12247 ({sk[2560], x592x, x19x, x21x, x505x, x502x, x493x}, x15663x);
	defparam lut_12247.LUT_SIZE = 7;
	defparam lut_12247.mask = 128'h37ff37ff3fff3fff00007f7f00ff7fff;

	lut_sub lut_12252 ({sk[2561], x13x, x24x, x574x, x542x}, x15433x);
	defparam lut_12252.LUT_SIZE = 5;
	defparam lut_12252.mask = 32'h5f5f0537;

	lut_sub lut_12255 ({sk[2562], i_9_, i_7_, i_8_, i_6_, n_n260, n_n464}, x15733x);
	defparam lut_12255.LUT_SIZE = 7;
	defparam lut_12255.mask = 128'h37ff37ff3fff3fff0001010001010000;

	lut_sub lut_12260 ({sk[2563], i_9_, x22x, n_n528, x506x, n_n464, n_n65}, x14560x);
	defparam lut_12260.LUT_SIZE = 7;
	defparam lut_12260.mask = 128'h37ff37ff3fff3fff0011111105151515;

	lut_sub lut_12265 ({sk[2564], i_9_, i_7_, i_8_, i_6_, n_n536, n_n473}, n_n3005);
	defparam lut_12265.LUT_SIZE = 7;
	defparam lut_12265.mask = 128'h37ff37ff3fff3fff1000110011111010;

	lut_sub lut_12275 ({sk[2565], x15x, x592x, x19x, x558x, x207x}, x15667x);
	defparam lut_12275.LUT_SIZE = 6;
	defparam lut_12275.mask = 64'h77ff77ff575757ff;

	lut_sub lut_12279 ({sk[2566], x21x, x13x, x587x, x542x}, x15439x);
	defparam lut_12279.LUT_SIZE = 5;
	defparam lut_12279.mask = 32'h5f5f0357;

	lut_sub lut_12282 ({sk[2567], x25x, x13x, x584x, x504x}, x15443x);
	defparam lut_12282.LUT_SIZE = 5;
	defparam lut_12282.mask = 32'h5f5f0357;

	lut_sub lut_12285 ({sk[2568], x22x, x13x, x510x, x23x, x543x}, x15444x);
	defparam lut_12285.LUT_SIZE = 6;
	defparam lut_12285.mask = 64'h77ff77ff111f555f;

	lut_sub lut_12289 ({sk[2569], x12x, x480x, x559x, x593x, n_n5087}, x15871x);
	defparam lut_12289.LUT_SIZE = 6;
	defparam lut_12289.mask = 64'h77ff77ff55557fff;

	lut_sub lut_12294 ({sk[2570], i_9_, n_n534, n_n535, n_n130, x23x, x598x}, x15870x);
	defparam lut_12294.LUT_SIZE = 7;
	defparam lut_12294.mask = 128'h37ff37ff3fff3fff1111111f1111111f;

	lut_sub lut_12298 ({sk[2571], x509x, x24x, x12x, x518x, x514x}, x15877x);
	defparam lut_12298.LUT_SIZE = 6;
	defparam lut_12298.mask = 64'h77ff77ff03570f5f;

	lut_sub lut_12302 ({sk[2572], x12x, x23x, x506x, x488x, x486x, n_n5131}, x22088x);
	defparam lut_12302.LUT_SIZE = 7;
	defparam lut_12302.mask = 128'h37ff37ff3fff3fffaaaa8888a0008000;

	lut_sub lut_12307 ({sk[2573], i_9_, i_7_, i_8_, i_6_, x484x, x596x}, x11678x);
	defparam lut_12307.LUT_SIZE = 7;
	defparam lut_12307.mask = 128'h37ff37ff3fff3fff0500000300000000;

	lut_sub lut_12310 ({sk[2574], x521x, x11x, x17x, x545x, x552x, x535x}, x22238x);
	defparam lut_12310.LUT_SIZE = 7;
	defparam lut_12310.mask = 128'h37ff37ff3fff3fffffa0cc80ff00cc00;

	lut_sub lut_12315 ({sk[2575], i_9_, i_7_, i_8_, i_6_, n_n500, n_n65}, n_n3665);
	defparam lut_12315.LUT_SIZE = 7;
	defparam lut_12315.mask = 128'h37ff37ff3fff3fff0111101001110010;

	lut_sub lut_12325 ({sk[2576], i_9_, i_7_, i_8_, i_6_, n_n536, n_n482}, x14505x);
	defparam lut_12325.LUT_SIZE = 7;
	defparam lut_12325.mask = 128'h37ff37ff3fff3fff1010000001000010;

	lut_sub lut_12330 ({sk[2577], x22x, x16x, x21x, x500x, x509x, x520x}, x22297x);
	defparam lut_12330.LUT_SIZE = 7;
	defparam lut_12330.mask = 128'h37ff37ff3fff3ffffff08880f0f08080;

	lut_sub lut_12335 ({sk[2578], i_9_, i_7_, i_8_, i_6_, n_n536, n_n473}, n_n3732);
	defparam lut_12335.LUT_SIZE = 7;
	defparam lut_12335.mask = 128'h37ff37ff3fff3fff0111101001111000;

	lut_sub lut_12345 ({sk[2579], i_9_, i_7_, i_8_, i_6_, n_n536, n_n482}, x14498x);
	defparam lut_12345.LUT_SIZE = 7;
	defparam lut_12345.mask = 128'h37ff37ff3fff3fff0000010100010100;

	lut_sub lut_12350 ({sk[2580], x22x, x16x, x500x, x510x, x520x}, x15540x);
	defparam lut_12350.LUT_SIZE = 6;
	defparam lut_12350.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_12354 ({sk[2581], x16x, x21x, x500x, x23x, x580x, x493x}, x22119x);
	defparam lut_12354.LUT_SIZE = 7;
	defparam lut_12354.mask = 128'h37ff37ff3fff3ffffff0ff0088808800;

	lut_sub lut_12359 ({sk[2582], i_9_, i_7_, i_8_, i_6_, x543x, x415x}, x16011x);
	defparam lut_12359.LUT_SIZE = 7;
	defparam lut_12359.mask = 128'h37ff37ff3fff3fff5575755555555555;

	lut_sub lut_12363 ({sk[2583], i_9_, i_7_, i_8_, i_6_, n_n491, n_n65}, n_n1825);
	defparam lut_12363.LUT_SIZE = 7;
	defparam lut_12363.mask = 128'h37ff37ff3fff3fff1110101001111000;

	lut_sub lut_12373 ({sk[2584], i_9_, i_7_, i_8_, i_6_, n_n482, n_n65}, n_n1824);
	defparam lut_12373.LUT_SIZE = 7;
	defparam lut_12373.mask = 128'h37ff37ff3fff3fff0001101101011110;

	lut_sub lut_12383 ({sk[2585], i_9_, n_n524, n_n534, n_n491, n_n500, n_n65}, x16304x);
	defparam lut_12383.LUT_SIZE = 7;
	defparam lut_12383.mask = 128'h37ff37ff3fff3fff0005111500051115;

	lut_sub lut_12388 ({sk[2586], x16x, x11x, x20x, x516x, x496x, x489x}, x22104x);
	defparam lut_12388.LUT_SIZE = 7;
	defparam lut_12388.mask = 128'h37ff37ff3fff3fffffcccccca0808080;

	lut_sub lut_12393 ({sk[2587], x13x, x11x, x233x, x482x, x540x, x194x}, x22337x);
	defparam lut_12393.LUT_SIZE = 7;
	defparam lut_12393.mask = 128'h37ff37ff3fff3fffaa008800a0008000;

	lut_sub lut_12398 ({sk[2588], i_9_, n_n482, n_n455, n_n532, x20x, x542x}, x16014x);
	defparam lut_12398.LUT_SIZE = 7;
	defparam lut_12398.mask = 128'h37ff37ff3fff3fff1111111f1111111f;

	lut_sub lut_12402 ({sk[2589], x15x, x22x, x13x, x584x, x493x, x543x}, x22103x);
	defparam lut_12402.LUT_SIZE = 7;
	defparam lut_12402.mask = 128'h37ff37ff3fff3fffffc0aa80aa80aa80;

	lut_sub lut_12407 ({sk[2590], i_9_, i_7_, i_8_, i_6_, n_n390, n_n500}, x16048x);
	defparam lut_12407.LUT_SIZE = 7;
	defparam lut_12407.mask = 128'h37ff37ff3fff3fff0101011110101001;

	lut_sub lut_12417 ({sk[2591], i_9_, i_7_, i_8_, i_6_, n_n390, n_n509}, n_n1876);
	defparam lut_12417.LUT_SIZE = 7;
	defparam lut_12417.mask = 128'h37ff37ff3fff3fff1111001011100010;

	lut_sub lut_12427 ({sk[2592], x21x, x10x, x583x, x585x}, x16037x);
	defparam lut_12427.LUT_SIZE = 5;
	defparam lut_12427.mask = 32'h5f5f0537;

	lut_sub lut_12430 ({sk[2593], x21x, x10x, x570x, x584x, x582x, x493x}, x16059x);
	defparam lut_12430.LUT_SIZE = 7;
	defparam lut_12430.mask = 128'h37ff37ff3fff3fff00005fff33337fff;

	lut_sub lut_12435 ({sk[2594], x10x, x509x, x580x, x502x, n_n4661, x193x}, x22101x);
	defparam lut_12435.LUT_SIZE = 7;
	defparam lut_12435.mask = 128'h37ff37ff3fff3fff8888888880000000;

	lut_sub lut_12438 ({sk[2595], x25x, x10x, x507x, x558x, x586x, x338x}, x22102x);
	defparam lut_12438.LUT_SIZE = 7;
	defparam lut_12438.mask = 128'h37ff37ff3fff3fffaaaa8080aa008000;

	lut_sub lut_12443 ({sk[2596], x25x, x21x, x582x, x192x, n_n1636}, x11882x);
	defparam lut_12443.LUT_SIZE = 6;
	defparam lut_12443.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_12448 ({sk[2597], x11856x, x11857x, x11859x, x11881x}, x11883x);
	defparam lut_12448.LUT_SIZE = 5;
	defparam lut_12448.mask = 32'h5f5f7fff;

	lut_sub lut_12453 ({sk[2598], i_9_, i_7_, i_8_, i_6_, n_n260, n_n535}, x14697x);
	defparam lut_12453.LUT_SIZE = 7;
	defparam lut_12453.mask = 128'h37ff37ff3fff3fff0001001001001000;

	lut_sub lut_12458 ({sk[2599], x21x, x14x, x516x, x530x}, x14706x);
	defparam lut_12458.LUT_SIZE = 5;
	defparam lut_12458.mask = 32'h5f5f0357;

	lut_sub lut_12461 ({sk[2600], x22x, x17x, x23x, x548x, x530x, n_n4820}, x22161x);
	defparam lut_12461.LUT_SIZE = 7;
	defparam lut_12461.mask = 128'h37ff37ff3fff3fffaa88a08088888080;

	lut_sub lut_12466 ({sk[2601], x14x, x488x, x527x, x528x, n_n4813, x151x}, x22160x);
	defparam lut_12466.LUT_SIZE = 7;
	defparam lut_12466.mask = 128'h37ff37ff3fff3fff8888888880000000;

	lut_sub lut_12469 ({sk[2602], x17x, x552x, x20x, x535x, x546x, x177x}, x22254x);
	defparam lut_12469.LUT_SIZE = 7;
	defparam lut_12469.mask = 128'h37ff37ff3fff3fffaaaaaa0080808000;

	lut_sub lut_12474 ({sk[2603], x592x, x538x, x19x, x510x, x23x, x520x}, x14564x);
	defparam lut_12474.LUT_SIZE = 7;
	defparam lut_12474.mask = 128'h37ff37ff3fff3fff005f00ff337f33ff;

	lut_sub lut_12479 ({sk[2604], i_9_, i_7_, i_8_, i_6_, n_n482, n_n65}, x14565x);
	defparam lut_12479.LUT_SIZE = 7;
	defparam lut_12479.mask = 128'h37ff37ff3fff3fff0001100011010000;

	lut_sub lut_12485 ({sk[2605], x19x, x522x, x268x, x527x, x528x}, x22156x);
	defparam lut_12485.LUT_SIZE = 6;
	defparam lut_12485.mask = 64'h77ff77fff0f08000;

	lut_sub lut_12488 ({sk[2606], x19x, x22x, x482x, x581x, x480x, x599x}, x14572x);
	defparam lut_12488.LUT_SIZE = 7;
	defparam lut_12488.mask = 128'h37ff37ff3fff3fff000055553fff7fff;

	lut_sub lut_12493 ({sk[2607], x15x, x19x, x475x, x478x, x487x, n_n5217}, x22155x);
	defparam lut_12493.LUT_SIZE = 7;
	defparam lut_12493.mask = 128'h37ff37ff3fff3fffaaaaa00088888000;

	lut_sub lut_12498 ({sk[2608], x25x, x19x, x521x, x481x, x487x}, x14571x);
	defparam lut_12498.LUT_SIZE = 6;
	defparam lut_12498.mask = 64'h77ff77ff003f557f;

	lut_sub lut_12502 ({sk[2609], i_9_, i_7_, i_8_, i_6_, x487x, x555x}, x14578x);
	defparam lut_12502.LUT_SIZE = 7;
	defparam lut_12502.mask = 128'h37ff37ff3fff3fff0070700000000000;

	lut_sub lut_12507 ({sk[2610], x15x, x19x, x21x, x563x, x599x, n_n5259}, x22154x);
	defparam lut_12507.LUT_SIZE = 7;
	defparam lut_12507.mask = 128'h37ff37ff3fff3fffaa88a08088888080;

	lut_sub lut_12512 ({sk[2611], x25x, x19x, x521x, x481x, x480x, x487x}, x22095x);
	defparam lut_12512.LUT_SIZE = 7;
	defparam lut_12512.mask = 128'h37ff37ff3fff3fffffffc000aaaa8000;

	lut_sub lut_12517 ({sk[2612], i_9_, x490x, x585x, n_n65, x182x}, x16272x);
	defparam lut_12517.LUT_SIZE = 6;
	defparam lut_12517.mask = 64'h77ff77ff55555777;

	lut_sub lut_12521 ({sk[2613], x25x, x19x, x594x, x599x}, x16270x);
	defparam lut_12521.LUT_SIZE = 5;
	defparam lut_12521.mask = 32'h5f5f0357;

	lut_sub lut_12524 ({sk[2614], x15x, x19x, x474x, x562x, x569x}, x16277x);
	defparam lut_12524.LUT_SIZE = 6;
	defparam lut_12524.mask = 64'h77ff77ff003f557f;

	lut_sub lut_12528 ({sk[2615], x19x, x22x, x21x, x472x, x563x, x487x}, x16278x);
	defparam lut_12528.LUT_SIZE = 7;
	defparam lut_12528.mask = 128'h37ff37ff3fff3fff005555553f7f7f7f;

	lut_sub lut_12533 ({sk[2616], i_9_, i_7_, i_8_, i_6_, n_n473, n_n325}, x14714x);
	defparam lut_12533.LUT_SIZE = 7;
	defparam lut_12533.mask = 128'h37ff37ff3fff3fff0000001001011000;

	lut_sub lut_12538 ({sk[2617], i_9_, i_7_, i_8_, i_6_, x588x, x511x}, x14712x);
	defparam lut_12538.LUT_SIZE = 7;
	defparam lut_12538.mask = 128'h37ff37ff3fff3fff3000500000000000;

	lut_sub lut_12541 ({sk[2618], i_9_, i_7_, i_8_, i_6_, n_n482, n_n325}, x14721x);
	defparam lut_12541.LUT_SIZE = 7;
	defparam lut_12541.mask = 128'h37ff37ff3fff3fff0011011011100000;

	lut_sub lut_12549 ({sk[2619], i_9_, i_7_, i_8_, i_6_, n_n509, n_n130}, n_n3676);
	defparam lut_12549.LUT_SIZE = 7;
	defparam lut_12549.mask = 128'h37ff37ff3fff3fff0110111001011010;

	lut_sub lut_12559 ({sk[2620], x25x, x12x, x481x, x486x}, x14608x);
	defparam lut_12559.LUT_SIZE = 5;
	defparam lut_12559.mask = 32'h5f5f0357;

	lut_sub lut_12562 ({sk[2621], x21x, x12x, x482x, x23x, x598x, x494x}, x14609x);
	defparam lut_12562.LUT_SIZE = 7;
	defparam lut_12562.mask = 128'h37ff37ff3fff3fff030357ff333377ff;

	lut_sub lut_12567 ({sk[2622], i_9_, i_7_, i_8_, i_6_, n_n130, n_n500}, x14611x);
	defparam lut_12567.LUT_SIZE = 7;
	defparam lut_12567.mask = 128'h37ff37ff3fff3fff0001011000010110;

	lut_sub lut_12574 ({sk[2623], i_9_, i_7_, i_8_, i_6_, x533x, x188x}, x14624x);
	defparam lut_12574.LUT_SIZE = 7;
	defparam lut_12574.mask = 128'h37ff37ff3fff3fff5555755555555555;

	lut_sub lut_12577 ({sk[2624], x22x, x11x, x12x, x514x, x525x, x489x}, x14625x);
	defparam lut_12577.LUT_SIZE = 7;
	defparam lut_12577.mask = 128'h37ff37ff3fff3fff00770f7f0f7f0f7f;

	lut_sub lut_12582 ({sk[2625], i_9_, i_7_, i_8_, i_6_, n_n473, n_n130}, x14626x);
	defparam lut_12582.LUT_SIZE = 7;
	defparam lut_12582.mask = 128'h37ff37ff3fff3fff1001000001110000;

	lut_sub lut_12588 ({sk[2626], i_9_, i_7_, i_8_, i_6_, n_n535, n_n65}, x14627x);
	defparam lut_12588.LUT_SIZE = 7;
	defparam lut_12588.mask = 128'h37ff37ff3fff3fff0101000101000110;

	lut_sub lut_12595 ({sk[2627], i_9_, i_7_, i_8_, i_6_, n_n195, n_n500}, n_n3685);
	defparam lut_12595.LUT_SIZE = 7;
	defparam lut_12595.mask = 128'h37ff37ff3fff3fff0101010101010111;

	lut_sub lut_12605 ({sk[2628], i_9_, i_7_, i_8_, i_6_, n_n509, n_n195}, n_n3686);
	defparam lut_12605.LUT_SIZE = 7;
	defparam lut_12605.mask = 128'h37ff37ff3fff3fff1111101011000010;

	lut_sub lut_12615 ({sk[2629], i_9_, i_7_, i_8_, i_6_, n_n536, n_n464}, x14522x);
	defparam lut_12615.LUT_SIZE = 7;
	defparam lut_12615.mask = 128'h37ff37ff3fff3fff0001010000011100;

	lut_sub lut_12621 ({sk[2630], x17x, x20x, x520x, x589x}, x14746x);
	defparam lut_12621.LUT_SIZE = 5;
	defparam lut_12621.mask = 32'h5f5f0537;

	lut_sub lut_12624 ({sk[2631], x538x, x21x, x17x, x508x, x580x, x531x}, x14748x);
	defparam lut_12624.LUT_SIZE = 7;
	defparam lut_12624.mask = 128'h37ff37ff3fff3fff003f557f00ff55ff;

	lut_sub lut_12629 ({sk[2632], x25x, x521x, x18x, x485x, x481x, x494x}, x14762x);
	defparam lut_12629.LUT_SIZE = 7;
	defparam lut_12629.mask = 128'h37ff37ff3fff3fff007700ff0f7f0fff;

	lut_sub lut_12634 ({sk[2633], i_9_, i_7_, i_8_, i_6_, x597x, x485x}, x14757x);
	defparam lut_12634.LUT_SIZE = 7;
	defparam lut_12634.mask = 128'h37ff37ff3fff3fff0030050000000000;

	lut_sub lut_12637 ({sk[2634], x22x, x539x, x18x, x597x, x585x, x43x}, x22151x);
	defparam lut_12637.LUT_SIZE = 7;
	defparam lut_12637.mask = 128'h37ff37ff3fff3fffaa88aa00a080a000;

	lut_sub lut_12642 ({sk[2635], i_9_, i_7_, i_8_, i_6_, n_n535, n_n195}, x15726x);
	defparam lut_12642.LUT_SIZE = 7;
	defparam lut_12642.mask = 128'h37ff37ff3fff3fff0010010100010000;

	lut_sub lut_12647 ({sk[2636], x20x, x23x, x531x, x341x, x15725x}, x15727x);
	defparam lut_12647.LUT_SIZE = 6;
	defparam lut_12647.mask = 64'h77ff77ff777f7f7f;

	lut_sub lut_12652 ({sk[2637], x15x, x483x, x23x, x565x, x15781x, x15782x}, x15784x);
	defparam lut_12652.LUT_SIZE = 7;
	defparam lut_12652.mask = 128'h37ff37ff3fff3fff777777ff7f7f7fff;

	lut_sub lut_12657 ({sk[2638], x14x, x494x, n_n4727, x15746x, n_n2982, x15745x}, x15785x);
	defparam lut_12657.LUT_SIZE = 7;
	defparam lut_12657.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_12663 ({sk[2639], x21x, x14x, x23x, x488x, x529x, x511x}, x15794x);
	defparam lut_12663.LUT_SIZE = 7;
	defparam lut_12663.mask = 128'h37ff37ff3fff3fff00553f7f55557f7f;

	lut_sub lut_12668 ({sk[2640], i_9_, n_n526, n_n473, n_n325, x522x, x381x}, x15795x);
	defparam lut_12668.LUT_SIZE = 7;
	defparam lut_12668.mask = 128'h37ff37ff3fff3fff555555555757575f;

	lut_sub lut_12672 ({sk[2641], x21x, x11x, x24x, x588x, x511x, x292x}, x22124x);
	defparam lut_12672.LUT_SIZE = 7;
	defparam lut_12672.mask = 128'h37ff37ff3fff3fffaa888888a0808080;

	lut_sub lut_12677 ({sk[2642], x25x, x16x, x529x, x496x, x527x}, x11525x);
	defparam lut_12677.LUT_SIZE = 6;
	defparam lut_12677.mask = 64'h77ff77ff005f337f;

	lut_sub lut_12681 ({sk[2643], i_9_, n_n536, n_n524, n_n473, n_n532, n_n464}, x11526x);
	defparam lut_12681.LUT_SIZE = 7;
	defparam lut_12681.mask = 128'h37ff37ff3fff3fff0000111f0000111f;

	lut_sub lut_12686 ({sk[2644], x16x, x13x, x550x, x516x, x236x, x525x}, x22248x);
	defparam lut_12686.LUT_SIZE = 7;
	defparam lut_12686.mask = 128'h37ff37ff3fff3fffcccccc0080808000;

	lut_sub lut_12691 ({sk[2645], i_9_, i_7_, i_8_, i_6_, n_n390, n_n500}, x11554x);
	defparam lut_12691.LUT_SIZE = 7;
	defparam lut_12691.mask = 128'h37ff37ff3fff3fff0010101010000000;

	lut_sub lut_12696 ({sk[2646], x16x, x23x, x497x, x594x, x559x, n_n4331}, x22241x);
	defparam lut_12696.LUT_SIZE = 7;
	defparam lut_12696.mask = 128'h37ff37ff3fff3fffaaaaaa0080808000;

	lut_sub lut_12701 ({sk[2647], x22x, x16x, x501x, x482x, x23x}, x22262x);
	defparam lut_12701.LUT_SIZE = 6;
	defparam lut_12701.mask = 64'h77ff77fffac8f0c0;

	lut_sub lut_12706 ({sk[2648], x11x, x12x, x477x, x486x}, x11710x);
	defparam lut_12706.LUT_SIZE = 5;
	defparam lut_12706.mask = 32'h5f5f0357;

	lut_sub lut_12709 ({sk[2649], x12x, x563x, x494x, x560x}, x11711x);
	defparam lut_12709.LUT_SIZE = 5;
	defparam lut_12709.mask = 32'h5f5f007f;

	lut_sub lut_12713 ({sk[2650], x515x, x19x, x24x, x580x, n_n5329, n_n5335}, x22235x);
	defparam lut_12713.LUT_SIZE = 7;
	defparam lut_12713.mask = 128'h37ff37ff3fff3fff8888808088008000;

	lut_sub lut_12718 ({sk[2651], x25x, x15x, x11x, x533x, x555x, x89x}, x22234x);
	defparam lut_12718.LUT_SIZE = 7;
	defparam lut_12718.mask = 128'h37ff37ff3fff3fffaaa0a0a088808080;

	lut_sub lut_12723 ({sk[2652], x16x, x570x, x490x, x494x, x537x}, x11741x);
	defparam lut_12723.LUT_SIZE = 6;
	defparam lut_12723.mask = 64'h77ff77ff00007fff;

	lut_sub lut_12728 ({sk[2653], x16x, x21x, x497x, x560x, n_n1002, x11741x}, x11743x);
	defparam lut_12728.LUT_SIZE = 7;
	defparam lut_12728.mask = 128'h37ff37ff3fff3fff777777ff7f7f7fff;

	lut_sub lut_12733 ({sk[2654], i_9_, i_7_, i_8_, i_6_, n_n482, n_n390}, x11881x);
	defparam lut_12733.LUT_SIZE = 7;
	defparam lut_12733.mask = 128'h37ff37ff3fff3fff0100011001010110;

	lut_sub lut_12741 ({sk[2655], x24x, x14x, x588x, x23x, x584x, x575x}, x11887x);
	defparam lut_12741.LUT_SIZE = 7;
	defparam lut_12741.mask = 128'h37ff37ff3fff3fff0505373705ff37ff;

	lut_sub lut_12745 ({sk[2656], i_9_, i_7_, i_8_, i_6_, n_n482, n_n325}, x11888x);
	defparam lut_12745.LUT_SIZE = 7;
	defparam lut_12745.mask = 128'h37ff37ff3fff3fff0100000100000011;

	lut_sub lut_12750 ({sk[2657], i_9_, n_n534, n_n509, n_n195, x43x}, x12023x);
	defparam lut_12750.LUT_SIZE = 6;
	defparam lut_12750.mask = 64'h77ff77ff55575555;

	lut_sub lut_12753 ({sk[2658], i_9_, i_7_, i_8_, i_6_, n_n509, n_n195}, x12024x);
	defparam lut_12753.LUT_SIZE = 7;
	defparam lut_12753.mask = 128'h37ff37ff3fff3fff0000011000010010;

	lut_sub lut_12758 ({sk[2659], x24x, x474x, x18x, x103x, x567x, x556x}, x22243x);
	defparam lut_12758.LUT_SIZE = 7;
	defparam lut_12758.mask = 128'h37ff37ff3fff3ffff0a0f000c080c000;

	lut_sub lut_12763 ({sk[2660], x15x, x12x, x518x, x578x}, x12030x);
	defparam lut_12763.LUT_SIZE = 5;
	defparam lut_12763.mask = 32'h5f5f0357;

	lut_sub lut_12766 ({sk[2661], i_9_, i_7_, i_8_, i_6_, n_n130, n_n500}, x12032x);
	defparam lut_12766.LUT_SIZE = 7;
	defparam lut_12766.mask = 128'h37ff37ff3fff3fff0010101000100000;

	lut_sub lut_12771 ({sk[2662], x492x, x21x, x17x, x570x, x531x}, x12088x);
	defparam lut_12771.LUT_SIZE = 6;
	defparam lut_12771.mask = 64'h77ff77ff03570f5f;

	lut_sub lut_12775 ({sk[2663], x25x, x19x, x23x, x524x, x534x}, x12127x);
	defparam lut_12775.LUT_SIZE = 6;
	defparam lut_12775.mask = 64'h77ff77ff05375577;

	lut_sub lut_12779 ({sk[2664], x19x, x558x, x17x, x580x, x502x, x493x}, x22220x);
	defparam lut_12779.LUT_SIZE = 7;
	defparam lut_12779.mask = 128'h37ff37ff3fff3fffff88ff88f0800000;

	lut_sub lut_12784 ({sk[2665], x16x, x509x, x24x, x496x, x528x}, x12135x);
	defparam lut_12784.LUT_SIZE = 6;
	defparam lut_12784.mask = 64'h77ff77ff030357ff;

	lut_sub lut_12788 ({sk[2666], x16x, x501x, x23x, x581x, x546x}, x12140x);
	defparam lut_12788.LUT_SIZE = 6;
	defparam lut_12788.mask = 64'h77ff77ff000f777f;

	lut_sub lut_12792 ({sk[2667], x538x, x16x, x11x, x499x, x564x}, x22294x);
	defparam lut_12792.LUT_SIZE = 6;
	defparam lut_12792.mask = 64'h77ff77fffca8fc00;

	lut_sub lut_12797 ({sk[2668], x22x, x16x, x23x, x491x, x498x, x423x}, x22296x);
	defparam lut_12797.LUT_SIZE = 7;
	defparam lut_12797.mask = 128'h37ff37ff3fff3fffaa88a08088888080;

	lut_sub lut_12802 ({sk[2669], x15x, x500x, x22294x, x22296x}, x12148x);
	defparam lut_12802.LUT_SIZE = 5;
	defparam lut_12802.mask = 32'h5f5feeef;

	lut_sub lut_12806 ({sk[2670], x25x, x22x, x16x, x550x, x495x, n_n4331}, x22219x);
	defparam lut_12806.LUT_SIZE = 7;
	defparam lut_12806.mask = 128'h37ff37ff3fff3fffaaa0888088808880;

	lut_sub lut_12811 ({sk[2671], x12136x, x12141x, x12135x, x12140x, x22219x}, x12149x);
	defparam lut_12811.LUT_SIZE = 6;
	defparam lut_12811.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_12817 ({sk[2672], x15x, x18x, x485x, x481x, x480x}, x12154x);
	defparam lut_12817.LUT_SIZE = 6;
	defparam lut_12817.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_12821 ({sk[2673], x22x, x539x, x18x, x597x, x490x, x594x}, x22286x);
	defparam lut_12821.LUT_SIZE = 7;
	defparam lut_12821.mask = 128'h37ff37ff3fff3fffff88ff00f080f000;

	lut_sub lut_12826 ({sk[2674], x25x, x11x, x18x, x485x, x581x, x564x}, x22227x);
	defparam lut_12826.LUT_SIZE = 7;
	defparam lut_12826.mask = 128'h37ff37ff3fff3fffff88f080f080f080;

	lut_sub lut_12831 ({sk[2675], x21x, x14x, x20x, x488x, x511x, x440x}, x22287x);
	defparam lut_12831.LUT_SIZE = 7;
	defparam lut_12831.mask = 128'h37ff37ff3fff3fffaa88a08088888080;

	lut_sub lut_12836 ({sk[2676], x24x, x14x, x502x, x530x, x439x, x22287x}, x12245x);
	defparam lut_12836.LUT_SIZE = 7;
	defparam lut_12836.mask = 128'h37ff37ff3fff3fffbbbbbbffbfbfbfff;

	lut_sub lut_12841 ({sk[2677], x18x, x23x, x574x, x560x, x567x}, x12251x);
	defparam lut_12841.LUT_SIZE = 6;
	defparam lut_12841.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_12845 ({sk[2678], x11x, x12x, x572x, x568x}, x12263x);
	defparam lut_12845.LUT_SIZE = 5;
	defparam lut_12845.mask = 32'h5f5f0357;

	lut_sub lut_12848 ({sk[2679], x12x, x23x, x486x, x562x}, x12299x);
	defparam lut_12848.LUT_SIZE = 5;
	defparam lut_12848.mask = 32'h5f5f0357;

	lut_sub lut_12851 ({sk[2680], x22x, x474x, x12x, x564x, x486x}, x12300x);
	defparam lut_12851.LUT_SIZE = 6;
	defparam lut_12851.mask = 64'h77ff77ff030f575f;

	lut_sub lut_12855 ({sk[2681], x19x, x21x, x570x, x519x, x579x}, x12375x);
	defparam lut_12855.LUT_SIZE = 6;
	defparam lut_12855.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_12859 ({sk[2682], i_9_, n_n482, x510x, x23x, n_n65, x63x}, x12376x);
	defparam lut_12859.LUT_SIZE = 7;
	defparam lut_12859.mask = 128'h37ff37ff3fff3fff5555575755775777;

	lut_sub lut_12863 ({sk[2683], x21x, x18x, x586x, x20x, x577x}, x22280x);
	defparam lut_12863.LUT_SIZE = 6;
	defparam lut_12863.mask = 64'h77ff77ffeee0aaa0;

	lut_sub lut_12868 ({sk[2684], i_9_, i_7_, i_8_, i_6_, x541x, x308x}, x12512x);
	defparam lut_12868.LUT_SIZE = 7;
	defparam lut_12868.mask = 128'h37ff37ff3fff3fff5555755555555555;

	lut_sub lut_12871 ({sk[2685], x15x, x24x, x23x, x542x, x541x, n_n4504}, x22229x);
	defparam lut_12871.LUT_SIZE = 7;
	defparam lut_12871.mask = 128'h37ff37ff3fff3fffaa88a080a080a080;

	lut_sub lut_12876 ({sk[2686], x21x, x17x, x512x, x489x}, x12687x);
	defparam lut_12876.LUT_SIZE = 5;
	defparam lut_12876.mask = 32'h5f5f0537;

	lut_sub lut_12879 ({sk[2687], x17x, x18x, x503x, x529x, x525x, x548x}, x12689x);
	defparam lut_12879.LUT_SIZE = 7;
	defparam lut_12879.mask = 128'h37ff37ff3fff3fff000055553fff7fff;

	lut_sub lut_12884 ({sk[2688], x22x, x21x, x13x, x549x, x498x, x495x}, x12699x);
	defparam lut_12884.LUT_SIZE = 7;
	defparam lut_12884.mask = 128'h37ff37ff3fff3fff000f333f555f777f;

	lut_sub lut_12888 ({sk[2689], x13x, x544x, x20x, x23x, x540x, x537x}, x12706x);
	defparam lut_12888.LUT_SIZE = 7;
	defparam lut_12888.mask = 128'h37ff37ff3fff3fff00330f3f55775f7f;

	lut_sub lut_12892 ({sk[2690], x16x, x521x, x23x, x497x, x546x}, x12713x);
	defparam lut_12892.LUT_SIZE = 6;
	defparam lut_12892.mask = 64'h77ff77ff030357ff;

	lut_sub lut_12896 ({sk[2691], i_9_, i_7_, i_8_, i_6_, x576x}, x12722x);
	defparam lut_12896.LUT_SIZE = 6;
	defparam lut_12896.mask = 64'h77ff77ff01040000;

	lut_sub lut_12899 ({sk[2692], x24x, x17x, x586x, x537x, x589x}, x12723x);
	defparam lut_12899.LUT_SIZE = 6;
	defparam lut_12899.mask = 64'h77ff77ff003f557f;

	lut_sub lut_12903 ({sk[2693], x21x, x24x, x17x, x491x, x566x, x576x}, x12770x);
	defparam lut_12903.LUT_SIZE = 7;
	defparam lut_12903.mask = 128'h37ff37ff3fff3fff000f555f333f777f;

	lut_sub lut_12907 ({sk[2694], x22x, x17x, x23x, x518x, x566x, x536x}, x22212x);
	defparam lut_12907.LUT_SIZE = 7;
	defparam lut_12907.mask = 128'h37ff37ff3fff3fffffcca080cccc8080;

	lut_sub lut_12912 ({sk[2695], x538x, x510x, x558x, x17x, x23x, x589x}, x12861x);
	defparam lut_12912.LUT_SIZE = 7;
	defparam lut_12912.mask = 128'h37ff37ff3fff3fff111f1f1f1f1f1f1f;

	lut_sub lut_12917 ({sk[2696], i_9_, i_7_, i_8_, i_6_, n_n482, n_n260}, x12862x);
	defparam lut_12917.LUT_SIZE = 7;
	defparam lut_12917.mask = 128'h37ff37ff3fff3fff0000101000111000;

	lut_sub lut_12923 ({sk[2697], i_9_, n_n526, n_n491, n_n130, n_n530, n_n3771}, x12894x);
	defparam lut_12923.LUT_SIZE = 7;
	defparam lut_12923.mask = 128'h37ff37ff3fff3fff5555555f55575557;

	lut_sub lut_12927 ({sk[2698], i_9_, i_7_, i_8_, i_6_, n_n130, n_n500}, x12895x);
	defparam lut_12927.LUT_SIZE = 7;
	defparam lut_12927.mask = 128'h37ff37ff3fff3fff0000110000111100;

	lut_sub lut_12934 ({sk[2699], i_9_, i_7_, i_8_, i_6_, x592x, x207x}, x12979x);
	defparam lut_12934.LUT_SIZE = 7;
	defparam lut_12934.mask = 128'h37ff37ff3fff3fff5755755555555555;

	lut_sub lut_12938 ({sk[2700], i_9_, i_7_, i_8_, i_6_, n_n482, n_n65}, x12980x);
	defparam lut_12938.LUT_SIZE = 7;
	defparam lut_12938.mask = 128'h37ff37ff3fff3fff0000010100011100;

	lut_sub lut_12944 ({sk[2701], i_9_, i_7_, i_8_, i_6_, x515x, x116x}, x22206x);
	defparam lut_12944.LUT_SIZE = 7;
	defparam lut_12944.mask = 128'h37ff37ff3fff3fff8aaa8a8aaaaaaaaa;

	lut_sub lut_12949 ({sk[2702], x510x, x12x, n_n5181, x503x, x44x}, x22258x);
	defparam lut_12949.LUT_SIZE = 6;
	defparam lut_12949.mask = 64'h77ff77ffa080a000;

	lut_sub lut_12952 ({sk[2703], i_9_, i_7_, i_8_, i_6_, x501x, x497x}, x13051x);
	defparam lut_12952.LUT_SIZE = 7;
	defparam lut_12952.mask = 128'h37ff37ff3fff3fff0050000300000000;

	lut_sub lut_12955 ({sk[2704], x16x, x21x, x497x, x593x}, x13052x);
	defparam lut_12955.LUT_SIZE = 5;
	defparam lut_12955.mask = 32'h5f5f0357;

	lut_sub lut_12958 ({sk[2705], x16x, x21x, x501x, x482x}, x13082x);
	defparam lut_12958.LUT_SIZE = 5;
	defparam lut_12958.mask = 32'h5f5f0357;

	lut_sub lut_12961 ({sk[2706], i_9_, i_7_, i_8_, i_6_, x515x, x592x}, x13140x);
	defparam lut_12961.LUT_SIZE = 7;
	defparam lut_12961.mask = 128'h37ff37ff3fff3fff0005005300000000;

	lut_sub lut_12965 ({sk[2707], x25x, x20x, x540x, x496x, n_n4404, n_n4384}, x22216x);
	defparam lut_12965.LUT_SIZE = 7;
	defparam lut_12965.mask = 128'h37ff37ff3fff3fff8888808088008000;

	lut_sub lut_12970 ({sk[2708], x538x, x19x, x492x, x24x, x499x, n_n4399}, x22341x);
	defparam lut_12970.LUT_SIZE = 7;
	defparam lut_12970.mask = 128'h37ff37ff3fff3fffa8a8a800a8a80000;

	lut_sub lut_12975 ({sk[2709], x501x, x13x, x24x, x564x, x593x, n_n4350}, x22215x);
	defparam lut_12975.LUT_SIZE = 7;
	defparam lut_12975.mask = 128'h37ff37ff3fff3fffaaaa8080aa008000;

	lut_sub lut_12980 ({sk[2710], x21x, x17x, x23x, x566x, x560x}, x13192x);
	defparam lut_12980.LUT_SIZE = 6;
	defparam lut_12980.mask = 64'h77ff77ff03573377;

	lut_sub lut_12984 ({sk[2711], x25x, x24x, x474x, x17x, x472x, x566x}, x13231x);
	defparam lut_12984.LUT_SIZE = 7;
	defparam lut_12984.mask = 128'h37ff37ff3fff3fff030f575f575f575f;

	lut_sub lut_12989 ({sk[2712], i_9_, i_7_, i_8_, i_6_, x568x, x76x}, x13282x);
	defparam lut_12989.LUT_SIZE = 7;
	defparam lut_12989.mask = 128'h37ff37ff3fff3fff7555555555555555;

	lut_sub lut_12992 ({sk[2713], i_9_, n_n509, n_n520, n_n130, x472x, x563x}, x13322x);
	defparam lut_12992.LUT_SIZE = 7;
	defparam lut_12992.mask = 128'h37ff37ff3fff3fff0000000f0707070f;

	lut_sub lut_12997 ({sk[2714], x22x, x474x, x12x, x20x, x477x, x486x}, x22275x);
	defparam lut_12997.LUT_SIZE = 7;
	defparam lut_12997.mask = 128'h37ff37ff3fff3ffffac8fa00aa88aa00;

	lut_sub lut_13002 ({sk[2715], x11x, x12x, x557x, x491x, x560x, x568x}, x22184x);
	defparam lut_13002.LUT_SIZE = 7;
	defparam lut_13002.mask = 128'h37ff37ff3fff3fffffffc000aaaa8000;

	lut_sub lut_13007 ({sk[2716], x592x, x19x, x21x, x24x, x558x, x586x}, x22183x);
	defparam lut_13007.LUT_SIZE = 7;
	defparam lut_13007.mask = 128'h37ff37ff3fff3fffffff8888f0008000;

	lut_sub lut_13012 ({sk[2717], x19x, x492x, x20x, x587x, x584x, x579x}, x22322x);
	defparam lut_13012.LUT_SIZE = 7;
	defparam lut_13012.mask = 128'h37ff37ff3fff3fffffaaffaac0800000;

	lut_sub lut_13017 ({sk[2718], x25x, x515x, x19x, x509x, x510x, n_n5303}, x22182x);
	defparam lut_13017.LUT_SIZE = 7;
	defparam lut_13017.mask = 128'h37ff37ff3fff3fffaa80aa80aa800000;

	lut_sub lut_13022 ({sk[2719], x25x, x13x, x522x, x547x}, x13469x);
	defparam lut_13022.LUT_SIZE = 5;
	defparam lut_13022.mask = 32'h5f5f0357;

	lut_sub lut_13025 ({sk[2720], i_9_, n_n482, n_n455, x510x, n_n522, x520x}, x13478x);
	defparam lut_13025.LUT_SIZE = 7;
	defparam lut_13025.mask = 128'h37ff37ff3fff3fff00000033005f007f;

	lut_sub lut_13030 ({sk[2721], x13x, x23x, x594x, x540x, x593x}, x13549x);
	defparam lut_13030.LUT_SIZE = 6;
	defparam lut_13030.mask = 64'h77ff77ff00335f7f;

	lut_sub lut_13034 ({sk[2722], x13x, x544x, x474x, x20x, x494x, n_n4489}, x22190x);
	defparam lut_13034.LUT_SIZE = 7;
	defparam lut_13034.mask = 128'h37ff37ff3fff3fffaaaaa0a088008000;

	lut_sub lut_13039 ({sk[2723], i_9_, i_7_, i_8_, i_6_, x486x}, x13577x);
	defparam lut_13039.LUT_SIZE = 6;
	defparam lut_13039.mask = 64'h77ff77ff11000000;

	lut_sub lut_13042 ({sk[2724], x22x, x21x, x12x, x574x, x568x}, x13578x);
	defparam lut_13042.LUT_SIZE = 6;
	defparam lut_13042.mask = 64'h77ff77ff03575757;

	lut_sub lut_13046 ({sk[2725], x19x, x21x, x474x, x555x}, x13584x);
	defparam lut_13046.LUT_SIZE = 5;
	defparam lut_13046.mask = 32'h5f5f0537;

	lut_sub lut_13049 ({sk[2726], x19x, x24x, x482x, x599x, x546x}, x13585x);
	defparam lut_13049.LUT_SIZE = 6;
	defparam lut_13049.mask = 64'h77ff77ff00335f7f;

	lut_sub lut_13053 ({sk[2727], i_9_, i_1_, i_2_, i_0_, x506x, x528x}, x13609x);
	defparam lut_13053.LUT_SIZE = 7;
	defparam lut_13053.mask = 128'h37ff37ff3fff3fff0000000000700000;

	lut_sub lut_13056 ({sk[2728], x25x, x492x, x12x, x23x, x591x, x514x}, x13611x);
	defparam lut_13056.LUT_SIZE = 7;
	defparam lut_13056.mask = 128'h37ff37ff3fff3fff070707ff575757ff;

	lut_sub lut_13061 ({sk[2729], x24x, x18x, x485x, x472x, x556x}, x13725x);
	defparam lut_13061.LUT_SIZE = 6;
	defparam lut_13061.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_13065 ({sk[2730], x15x, x474x, x18x, x503x, x563x, x513x}, x13726x);
	defparam lut_13065.LUT_SIZE = 7;
	defparam lut_13065.mask = 128'h37ff37ff3fff3fff003f00ff557f55ff;

	lut_sub lut_13070 ({sk[2731], x24x, x14x, x552x, x525x}, x13802x);
	defparam lut_13070.LUT_SIZE = 5;
	defparam lut_13070.mask = 32'h5f5f0537;

	lut_sub lut_13073 ({sk[2732], i_9_, i_7_, i_8_, i_6_, x530x, x185x}, x13803x);
	defparam lut_13073.LUT_SIZE = 7;
	defparam lut_13073.mask = 128'h37ff37ff3fff3fff5755555555555555;

	lut_sub lut_13076 ({sk[2733], x14x, x529x, n_n4807, x439x, n_n4196, x395x}, x13825x);
	defparam lut_13076.LUT_SIZE = 7;
	defparam lut_13076.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_13082 ({sk[2734], x38x, x186x, n_n3332, x13802x, x13803x}, x13826x);
	defparam lut_13082.LUT_SIZE = 6;
	defparam lut_13082.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_13088 ({sk[2735], x24x, x17x, x512x, x508x}, x13871x);
	defparam lut_13088.LUT_SIZE = 5;
	defparam lut_13088.mask = 32'h5f5f0537;

	lut_sub lut_13091 ({sk[2736], x18x, x23x, x573x, x567x}, x13993x);
	defparam lut_13091.LUT_SIZE = 5;
	defparam lut_13091.mask = 32'h5f5f0537;

	lut_sub lut_13094 ({sk[2737], i_9_, i_7_, i_8_, i_6_, x554x, x598x}, x14008x);
	defparam lut_13094.LUT_SIZE = 7;
	defparam lut_13094.mask = 128'h37ff37ff3fff3fff0000003500000000;

	lut_sub lut_13097 ({sk[2738], i_9_, n_n522, n_n130, n_n500, x518x, x573x}, x14061x);
	defparam lut_13097.LUT_SIZE = 7;
	defparam lut_13097.mask = 128'h37ff37ff3fff3fff0000000f0077007f;

	lut_sub lut_13102 ({sk[2739], x15x, x10x, x571x, x572x, x491x}, x14076x);
	defparam lut_13102.LUT_SIZE = 6;
	defparam lut_13102.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_13106 ({sk[2740], i_9_, i_7_, i_8_, i_6_, x561x, x571x}, x14077x);
	defparam lut_13106.LUT_SIZE = 7;
	defparam lut_13106.mask = 128'h37ff37ff3fff3fff0053530000000000;

	lut_sub lut_13111 ({sk[2741], x22x, x10x, x571x, x587x, x573x, x563x}, x14079x);
	defparam lut_13111.LUT_SIZE = 7;
	defparam lut_13111.mask = 128'h37ff37ff3fff3fff00007f7f00ff7fff;

	lut_sub lut_13116 ({sk[2742], x16x, x501x, x11x, x490x}, x14182x);
	defparam lut_13116.LUT_SIZE = 5;
	defparam lut_13116.mask = 32'h5f5f0357;

	lut_sub lut_13119 ({sk[2743], x16x, x24x, x481x, x480x, x473x}, x14190x);
	defparam lut_13119.LUT_SIZE = 6;
	defparam lut_13119.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_13123 ({sk[2744], i_9_, i_7_, i_8_, i_6_, n_n536, n_n518}, x14191x);
	defparam lut_13123.LUT_SIZE = 7;
	defparam lut_13123.mask = 128'h37ff37ff3fff3fff1000001010001000;

	lut_sub lut_13128 ({sk[2745], i_9_, n_n482, n_n455, n_n534, x20x, x542x}, x14205x);
	defparam lut_13128.LUT_SIZE = 7;
	defparam lut_13128.mask = 128'h37ff37ff3fff3fff1111111f1111111f;

	lut_sub lut_13132 ({sk[2746], i_9_, i_7_, i_8_, i_6_, n_n464, n_n65}, x14213x);
	defparam lut_13132.LUT_SIZE = 7;
	defparam lut_13132.mask = 128'h37ff37ff3fff3fff1010100010100000;

	lut_sub lut_13138 ({sk[2747], x474x, x18x, x20x, x506x, x513x}, x14272x);
	defparam lut_13138.LUT_SIZE = 6;
	defparam lut_13138.mask = 64'h77ff77ff053705ff;

	lut_sub lut_13142 ({sk[2748], x519x, x18x, x586x, x472x, x480x}, x14273x);
	defparam lut_13142.LUT_SIZE = 6;
	defparam lut_13142.mask = 64'h77ff77ff007f00ff;

	lut_sub lut_13147 ({sk[2749], x22x, x16x, x497x, x480x}, x14288x);
	defparam lut_13147.LUT_SIZE = 5;
	defparam lut_13147.mask = 32'h5f5f0537;

	lut_sub lut_13150 ({sk[2750], x16x, x21x, x490x, x549x, x473x}, x14289x);
	defparam lut_13150.LUT_SIZE = 6;
	defparam lut_13150.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_13154 ({sk[2751], x25x, x16x, x518x, x529x, x496x}, x14336x);
	defparam lut_13154.LUT_SIZE = 6;
	defparam lut_13154.mask = 64'h77ff77ff003f557f;

	lut_sub lut_13158 ({sk[2752], x16x, x510x, x580x, x560x, x562x}, x14337x);
	defparam lut_13158.LUT_SIZE = 6;
	defparam lut_13158.mask = 64'h77ff77ff00007fff;

	lut_sub lut_13163 ({sk[2753], x15x, x13x, x475x, x478x, x541x, x235x}, x22149x);
	defparam lut_13163.LUT_SIZE = 7;
	defparam lut_13163.mask = 128'h37ff37ff3fff3fffaaaaa00088888000;

	lut_sub lut_13168 ({sk[2754], x14283x, x14290x, x14288x, x14289x, x22149x}, x14340x);
	defparam lut_13168.LUT_SIZE = 6;
	defparam lut_13168.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_13174 ({sk[2755], x25x, x495x, n_n4399, x14336x, x14337x, x14340x}, x14341x);
	defparam lut_13174.LUT_SIZE = 7;
	defparam lut_13174.mask = 128'h37ff37ff3fff3fff7fff7fff7fffffff;

	lut_sub lut_13180 ({sk[2756], x14310x, x14332x, n_n3560, n_n3562, n_n3564, n_n3561}, x14342x);
	defparam lut_13180.LUT_SIZE = 7;
	defparam lut_13180.mask = 128'h37ff37ff3fff3fff7fffffffffffffff;

	lut_sub lut_13187 ({sk[2757], i_9_, i_7_, i_8_, i_6_, n_n518, n_n455}, x14534x);
	defparam lut_13187.LUT_SIZE = 7;
	defparam lut_13187.mask = 128'h37ff37ff3fff3fff0110000010001000;

	lut_sub lut_13192 ({sk[2758], x22x, x13x, x544x, x481x, x494x, x413x}, x22164x);
	defparam lut_13192.LUT_SIZE = 7;
	defparam lut_13192.mask = 128'h37ff37ff3fff3fffaaaa8080aa008000;

	lut_sub lut_13197 ({sk[2759], x19x, x24x, x557x, x579x}, x14543x);
	defparam lut_13197.LUT_SIZE = 5;
	defparam lut_13197.mask = 32'h5f5f0537;

	lut_sub lut_13200 ({sk[2760], x19x, x492x, x22x, x579x}, x14584x);
	defparam lut_13200.LUT_SIZE = 5;
	defparam lut_13200.mask = 32'h5f5f111f;

	lut_sub lut_13203 ({sk[2761], x25x, x592x, x19x, x519x}, x14586x);
	defparam lut_13203.LUT_SIZE = 5;
	defparam lut_13203.mask = 32'h5f5f111f;

	lut_sub lut_13206 ({sk[2762], x19x, x570x, x20x, x23x, x587x, x579x}, x22321x);
	defparam lut_13206.LUT_SIZE = 7;
	defparam lut_13206.mask = 128'h37ff37ff3fff3ffffaaafaaac8880000;

	lut_sub lut_13211 ({sk[2763], i_9_, i_7_, i_8_, i_6_, x591x, x514x}, x14632x);
	defparam lut_13211.LUT_SIZE = 7;
	defparam lut_13211.mask = 128'h37ff37ff3fff3fff3000000500000000;

	lut_sub lut_13214 ({sk[2764], i_9_, i_7_, i_8_, i_6_, n_n482, n_n130}, x14634x);
	defparam lut_13214.LUT_SIZE = 7;
	defparam lut_13214.mask = 128'h37ff37ff3fff3fff0011100000010000;

	lut_sub lut_13219 ({sk[2765], i_9_, n_n526, n_n482, n_n195, x577x, x520x}, x14665x);
	defparam lut_13219.LUT_SIZE = 7;
	defparam lut_13219.mask = 128'h37ff37ff3fff3fff0000333f0505050f;

	lut_sub lut_13224 ({sk[2766], i_9_, i_7_, i_8_, i_6_, n_n482, n_n195}, x14666x);
	defparam lut_13224.LUT_SIZE = 7;
	defparam lut_13224.mask = 128'h37ff37ff3fff3fff0101110001100000;

	lut_sub lut_13231 ({sk[2767], x25x, x18x, x572x, x577x, x573x, x560x}, x14680x);
	defparam lut_13231.LUT_SIZE = 7;
	defparam lut_13231.mask = 128'h37ff37ff3fff3fff000077ff0f0f7fff;

	lut_sub lut_13236 ({sk[2768], x17x, x20x, x566x, x573x}, x14732x);
	defparam lut_13236.LUT_SIZE = 5;
	defparam lut_13236.mask = 32'h5f5f0357;

	lut_sub lut_13239 ({sk[2769], i_9_, i_7_, i_8_, i_6_, x589x, x576x}, x14737x);
	defparam lut_13239.LUT_SIZE = 7;
	defparam lut_13239.mask = 128'h37ff37ff3fff3fff0050000300000000;

	lut_sub lut_13242 ({sk[2770], i_9_, i_7_, i_8_, i_6_, n_n464, n_n65}, x14774x);
	defparam lut_13242.LUT_SIZE = 7;
	defparam lut_13242.mask = 128'h37ff37ff3fff3fff1010100010101000;

	lut_sub lut_13249 ({sk[2771], x25x, x18x, x485x, x481x}, x14811x);
	defparam lut_13249.LUT_SIZE = 5;
	defparam lut_13249.mask = 32'h5f5f0537;

	lut_sub lut_13252 ({sk[2772], x11x, x18x, x597x, x23x, x517x}, x14812x);
	defparam lut_13252.LUT_SIZE = 6;
	defparam lut_13252.mask = 64'h77ff77ff03570f5f;

	lut_sub lut_13256 ({sk[2773], x22x, x17x, x484x, x560x}, x14818x);
	defparam lut_13256.LUT_SIZE = 5;
	defparam lut_13256.mask = 32'h5f5f0537;

	lut_sub lut_13259 ({sk[2774], x11x, x17x, x484x, x472x, x23x, x596x}, x14819x);
	defparam lut_13259.LUT_SIZE = 7;
	defparam lut_13259.mask = 128'h37ff37ff3fff3fff00330f3f55775f7f;

	lut_sub lut_13263 ({sk[2775], x22x, x509x, x24x, x17x, n_n4925, x589x}, x22134x);
	defparam lut_13263.LUT_SIZE = 7;
	defparam lut_13263.mask = 128'h37ff37ff3fff3fffcc88c08088888080;

	lut_sub lut_13268 ({sk[2776], x16x, x500x, x11x, x23x, x584x, x498x}, x14875x);
	defparam lut_13268.LUT_SIZE = 7;
	defparam lut_13268.mask = 128'h37ff37ff3fff3fff050505ff373737ff;

	lut_sub lut_13272 ({sk[2777], x16x, x11x, x475x, x473x, x593x}, x14881x);
	defparam lut_13272.LUT_SIZE = 6;
	defparam lut_13272.mask = 64'h77ff77ff00335f7f;

	lut_sub lut_13276 ({sk[2778], x16x, x13x, x488x, n_n4453, n_n4447, x535x}, x22132x);
	defparam lut_13276.LUT_SIZE = 7;
	defparam lut_13276.mask = 128'h37ff37ff3fff3fffc0c08080c0008000;

	lut_sub lut_13281 ({sk[2779], x500x, x23x, x234x, x327x, x22132x}, x14888x);
	defparam lut_13281.LUT_SIZE = 6;
	defparam lut_13281.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_13286 ({sk[2780], x25x, x16x, x497x, x563x, x548x, n_n4391}, x22131x);
	defparam lut_13286.LUT_SIZE = 7;
	defparam lut_13286.mask = 128'h37ff37ff3fff3fffaaaa8080aa008000;

	lut_sub lut_13291 ({sk[2781], x14876x, x14882x, x14875x, x14881x, x22131x}, x14889x);
	defparam lut_13291.LUT_SIZE = 6;
	defparam lut_13291.mask = 64'h77ff77ffbfffffff;

	lut_sub lut_13297 ({sk[2782], x14848x, x14849x, x14870x, n_n2467, n_n2466}, x14891x);
	defparam lut_13297.LUT_SIZE = 6;
	defparam lut_13297.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_13303 ({sk[2783], x15x, x17x, x20x, x482x, x481x, x596x}, x14904x);
	defparam lut_13303.LUT_SIZE = 7;
	defparam lut_13303.mask = 128'h37ff37ff3fff3fff00553f7f55557f7f;

	lut_sub lut_13308 ({sk[2784], i_9_, i_7_, i_8_, i_6_, n_n518, n_n260}, x14905x);
	defparam lut_13308.LUT_SIZE = 7;
	defparam lut_13308.mask = 128'h37ff37ff3fff3fff0000101000100110;

	lut_sub lut_13314 ({sk[2785], x22x, x510x, x14x, x558x, x520x, x530x}, x14924x);
	defparam lut_13314.LUT_SIZE = 7;
	defparam lut_13314.mask = 128'h37ff37ff3fff3fff003f00ff557f55ff;

	lut_sub lut_13319 ({sk[2786], i_9_, i_7_, i_8_, i_6_, n_n325, n_n464}, x14925x);
	defparam lut_13319.LUT_SIZE = 7;
	defparam lut_13319.mask = 128'h37ff37ff3fff3fff0001010101010100;

	lut_sub lut_13326 ({sk[2787], i_9_, i_7_, i_8_, i_6_, n_n518, n_n195}, x14977x);
	defparam lut_13326.LUT_SIZE = 7;
	defparam lut_13326.mask = 128'h37ff37ff3fff3fff0000001100000110;

	lut_sub lut_13331 ({sk[2788], x11x, x14x, x478x, x565x, x556x}, x14984x);
	defparam lut_13331.LUT_SIZE = 6;
	defparam lut_13331.mask = 64'h77ff77ff005f337f;

	lut_sub lut_13335 ({sk[2789], x24x, x14x, x588x, x23x, x584x, x575x}, x15020x);
	defparam lut_13335.LUT_SIZE = 7;
	defparam lut_13335.mask = 128'h37ff37ff3fff3fff0505373705ff37ff;

	lut_sub lut_13339 ({sk[2790], i_9_, x15x, n_n482, n_n534, n_n325, x570x}, x15021x);
	defparam lut_13339.LUT_SIZE = 7;
	defparam lut_13339.mask = 128'h37ff37ff3fff3fff0003003311131133;

	lut_sub lut_13344 ({sk[2791], i_9_, i_7_, i_8_, i_6_, x565x}, x22133x);
	defparam lut_13344.LUT_SIZE = 6;
	defparam lut_13344.mask = 64'h77ff77ffbebbffff;

	lut_sub lut_13350 ({sk[2792], x13x, x570x, x519x, x537x, x130x, x307x}, x22139x);
	defparam lut_13350.LUT_SIZE = 7;
	defparam lut_13350.mask = 128'h37ff37ff3fff3fff8888888880000000;

	lut_sub lut_13353 ({sk[2793], x25x, x11x, x542x, x543x, x504x, x415x}, x22140x);
	defparam lut_13353.LUT_SIZE = 7;
	defparam lut_13353.mask = 128'h37ff37ff3fff3fffaaaa8800a0a08000;

	lut_sub lut_13358 ({sk[2794], x22x, x13x, x522x, x523x}, x15142x);
	defparam lut_13358.LUT_SIZE = 5;
	defparam lut_13358.mask = 32'h5f5f0357;

	lut_sub lut_13361 ({sk[2795], i_9_, i_1_, i_2_, i_0_, x477x, x494x}, x15161x);
	defparam lut_13361.LUT_SIZE = 7;
	defparam lut_13361.mask = 128'h37ff37ff3fff3fff0000000000000007;

	lut_sub lut_13364 ({sk[2796], x22x, x16x, x474x, x480x, x473x}, x15162x);
	defparam lut_13364.LUT_SIZE = 6;
	defparam lut_13364.mask = 64'h77ff77ff003f557f;

	lut_sub lut_13368 ({sk[2797], x592x, x19x, x22x, x11x, x520x}, x15194x);
	defparam lut_13368.LUT_SIZE = 6;
	defparam lut_13368.mask = 64'h77ff77ff00553f7f;

	lut_sub lut_13372 ({sk[2798], x19x, x23x, x573x, x569x}, x15197x);
	defparam lut_13372.LUT_SIZE = 5;
	defparam lut_13372.mask = 32'h5f5f0537;

	lut_sub lut_13375 ({sk[2799], x15x, x592x, x19x, x558x, x20x, x579x}, x15201x);
	defparam lut_13375.LUT_SIZE = 7;
	defparam lut_13375.mask = 128'h37ff37ff3fff3fff111f111f111fffff;

	lut_sub lut_13379 ({sk[2800], i_9_, n_n524, n_n491, x570x, x587x, n_n65}, x15202x);
	defparam lut_13379.LUT_SIZE = 7;
	defparam lut_13379.mask = 128'h37ff37ff3fff3fff0000005515151555;

	lut_sub lut_13384 ({sk[2801], x25x, x515x, x22x, n_n5302, x579x, x217x}, x22137x);
	defparam lut_13384.LUT_SIZE = 7;
	defparam lut_13384.mask = 128'h37ff37ff3fff3fffa080a080a0800000;

	lut_sub lut_13389 ({sk[2802], i_9_, i_7_, i_8_, i_6_, n_n518, n_n130}, x15248x);
	defparam lut_13389.LUT_SIZE = 7;
	defparam lut_13389.mask = 128'h37ff37ff3fff3fff0101110001011001;

	lut_sub lut_13398 ({sk[2803], i_9_, i_7_, i_8_, i_6_, x591x, x578x}, x15281x);
	defparam lut_13398.LUT_SIZE = 7;
	defparam lut_13398.mask = 128'h37ff37ff3fff3fff0050030000000000;

	lut_sub lut_13401 ({sk[2804], x570x, x12x, x23x, x587x, x578x}, x15282x);
	defparam lut_13401.LUT_SIZE = 6;
	defparam lut_13401.mask = 64'h77ff77ff053705ff;

	lut_sub lut_13405 ({sk[2805], i_9_, i_7_, i_8_, i_6_, n_n130, n_n500}, x15293x);
	defparam lut_13405.LUT_SIZE = 7;
	defparam lut_13405.mask = 128'h37ff37ff3fff3fff0111101001101100;

	lut_sub lut_13415 ({sk[2806], x24x, x17x, x586x, x563x, x589x}, x15347x);
	defparam lut_13415.LUT_SIZE = 6;
	defparam lut_13415.mask = 64'h77ff77ff003f557f;

	lut_sub lut_13419 ({sk[2807], x22x, x11x, x18x, x535x, x553x}, x15389x);
	defparam lut_13419.LUT_SIZE = 6;
	defparam lut_13419.mask = 64'h77ff77ff03575757;

	lut_sub lut_13423 ({sk[2808], x15x, x18x, x550x, x549x, x553x}, x15395x);
	defparam lut_13423.LUT_SIZE = 6;
	defparam lut_13423.mask = 64'h77ff77ff003f557f;

	lut_sub lut_13427 ({sk[2809], x25x, x21x, x17x, x512x, x489x, x528x}, x22116x);
	defparam lut_13427.LUT_SIZE = 7;
	defparam lut_13427.mask = 128'h37ff37ff3fff3fffff88f080f080f080;

	lut_sub lut_13432 ({sk[2810], x17x, x20x, x529x, x589x, x15395x, x22116x}, x15398x);
	defparam lut_13432.LUT_SIZE = 7;
	defparam lut_13432.mask = 128'h37ff37ff3fff3fffbbbbbfbfbbffbfff;

	lut_sub lut_13437 ({sk[2811], x21x, x18x, x481x, x494x, x589x, n_n4886}, x22113x);
	defparam lut_13437.LUT_SIZE = 7;
	defparam lut_13437.mask = 128'h37ff37ff3fff3fffaaaaa00088888000;

	lut_sub lut_13442 ({sk[2812], x13x, x11x, x481x, x476x}, x15422x);
	defparam lut_13442.LUT_SIZE = 5;
	defparam lut_13442.mask = 32'h5f5f0537;

	lut_sub lut_13445 ({sk[2813], x13x, x544x, x11x, x490x, x517x, n_n4455}, x22112x);
	defparam lut_13445.LUT_SIZE = 7;
	defparam lut_13445.mask = 128'h37ff37ff3fff3fffaaaaaa0080808000;

	lut_sub lut_13450 ({sk[2814], x15x, x544x, x24x, x20x, x476x, n_n4472}, x22111x);
	defparam lut_13450.LUT_SIZE = 7;
	defparam lut_13450.mask = 128'h37ff37ff3fff3fffaa88a08088888080;

	lut_sub lut_13455 ({sk[2815], i_9_, i_7_, i_8_, i_6_, n_n455, n_n464}, x15501x);
	defparam lut_13455.LUT_SIZE = 7;
	defparam lut_13455.mask = 128'h37ff37ff3fff3fff0101011101010110;

	lut_sub lut_13465 ({sk[2816], x25x, x16x, x500x, x11x, x584x}, x15506x);
	defparam lut_13465.LUT_SIZE = 6;
	defparam lut_13465.mask = 64'h77ff77ff03570f5f;

	lut_sub lut_13469 ({sk[2817], x22x, x16x, x474x, x478x, x473x}, x15511x);
	defparam lut_13469.LUT_SIZE = 6;
	defparam lut_13469.mask = 64'h77ff77ff003f557f;

	lut_sub lut_13473 ({sk[2818], i_9_, i_7_, i_8_, i_6_, n_n536, n_n491}, x15546x);
	defparam lut_13473.LUT_SIZE = 7;
	defparam lut_13473.mask = 128'h37ff37ff3fff3fff0001000101010101;

	lut_sub lut_13480 ({sk[2819], x15x, x492x, x16x, x472x, x587x, x498x}, x22118x);
	defparam lut_13480.LUT_SIZE = 7;
	defparam lut_13480.mask = 128'h37ff37ff3fff3fffffc0ff00aa80aa00;

	lut_sub lut_13485 ({sk[2820], i_9_, i_7_, i_8_, i_6_, x533x, x555x}, x15560x);
	defparam lut_13485.LUT_SIZE = 7;
	defparam lut_13485.mask = 128'h37ff37ff3fff3fff0050530300000000;

	lut_sub lut_13490 ({sk[2821], x25x, x19x, x521x, x477x, x556x, x487x}, x15575x);
	defparam lut_13490.LUT_SIZE = 7;
	defparam lut_13490.mask = 128'h37ff37ff3fff3fff00003fff55557fff;

	lut_sub lut_13495 ({sk[2822], i_9_, i_7_, i_8_, i_6_, n_n473, n_n130}, x15591x);
	defparam lut_13495.LUT_SIZE = 7;
	defparam lut_13495.mask = 128'h37ff37ff3fff3fff0001000101010001;

	lut_sub lut_13501 ({sk[2823], x18x, x23x, x577x, x584x}, x15636x);
	defparam lut_13501.LUT_SIZE = 5;
	defparam lut_13501.mask = 32'h5f5f0357;

	lut_sub lut_13504 ({sk[2824], i_9_, x492x, n_n526, n_n491, n_n195, x587x}, x15638x);
	defparam lut_13504.LUT_SIZE = 7;
	defparam lut_13504.mask = 128'h37ff37ff3fff3fff0003000311133333;

	lut_sub lut_13509 ({sk[2825], x515x, x19x, x20x, x528x}, x15647x);
	defparam lut_13509.LUT_SIZE = 5;
	defparam lut_13509.mask = 32'h5f5f0537;

	lut_sub lut_13512 ({sk[2826], x515x, x19x, x21x, x506x, x529x}, x15648x);
	defparam lut_13512.LUT_SIZE = 6;
	defparam lut_13512.mask = 64'h77ff77ff00770f7f;

	lut_sub lut_13516 ({sk[2827], x25x, x592x, x19x, x24x, x584x}, x15666x);
	defparam lut_13516.LUT_SIZE = 6;
	defparam lut_13516.mask = 64'h77ff77ff053705ff;

	lut_sub lut_13520 ({sk[2828], x515x, x22x, x20x, x579x, n_n5303, n_n5295}, x22126x);
	defparam lut_13520.LUT_SIZE = 7;
	defparam lut_13520.mask = 128'h37ff37ff3fff3fff8880888088800000;

	lut_sub lut_13525 ({sk[2829], i_9_, i_7_, i_8_, i_6_, n_n464, n_n65}, x22125x);
	defparam lut_13525.LUT_SIZE = 7;
	defparam lut_13525.mask = 128'h37ff37ff3fff3fffefffeefeeeeeffef;

	lut_sub lut_13533 ({sk[2830], x21x, x545x, x18x, x517x, x531x, x546x}, x15725x);
	defparam lut_13533.LUT_SIZE = 7;
	defparam lut_13533.mask = 128'h37ff37ff3fff3fff005f00ff337f33ff;

	lut_sub lut_13538 ({sk[2831], x25x, x17x, x516x, x522x, x531x, x180x}, x22121x);
	defparam lut_13538.LUT_SIZE = 7;
	defparam lut_13538.mask = 128'h37ff37ff3fff3fffaaaaa00088888000;

	lut_sub lut_13543 ({sk[2832], x21x, x11x, x483x, x14x, x477x}, x15745x);
	defparam lut_13543.LUT_SIZE = 6;
	defparam lut_13543.mask = 64'h77ff77ff111f1f1f;

	lut_sub lut_13547 ({sk[2833], x24x, x14x, x478x, x565x, x562x}, x15781x);
	defparam lut_13547.LUT_SIZE = 6;
	defparam lut_13547.mask = 64'h77ff77ff005f337f;

	lut_sub lut_13551 ({sk[2834], i_9_, n_n509, n_n325, n_n522, x564x, x563x}, x15782x);
	defparam lut_13551.LUT_SIZE = 7;
	defparam lut_13551.mask = 128'h37ff37ff3fff3fff0000000f0077007f;

	lut_sub lut_13556 ({sk[2835], x11x, x17x, x491x, x566x}, x15801x);
	defparam lut_13556.LUT_SIZE = 5;
	defparam lut_13556.mask = 32'h5f5f0357;

	lut_sub lut_13559 ({sk[2836], i_9_, i_7_, i_8_, i_6_, n_n260, n_n500}, x15802x);
	defparam lut_13559.LUT_SIZE = 7;
	defparam lut_13559.mask = 128'h37ff37ff3fff3fff0000010101001000;

	lut_sub lut_13564 ({sk[2837], x15342x, x15418x, n_n2839, n_n2842, n_n2841, n_n2838}, x15812x);
	defparam lut_13564.LUT_SIZE = 7;
	defparam lut_13564.mask = 128'h37ff37ff3fff3fff7fffffffffffffff;

	lut_sub lut_13571 ({sk[2838], n_n2845, n_n2844, n_n2846, n_n2831, x15385x, x15398x}, x22106x);
	defparam lut_13571.LUT_SIZE = 7;
	defparam lut_13571.mask = 128'h37ff37ff3fff3fff8000000000000000;

	lut_sub lut_13573 ({sk[2839], x15x, x19x, x581x, x537x, x487x}, x15844x);
	defparam lut_13573.LUT_SIZE = 6;
	defparam lut_13573.mask = 64'h77ff77ff003f557f;

	lut_sub lut_13577 ({sk[2840], i_9_, i_7_, i_8_, i_6_, x592x, x534x}, x15898x);
	defparam lut_13577.LUT_SIZE = 7;
	defparam lut_13577.mask = 128'h37ff37ff3fff3fff3055500000000000;

	lut_sub lut_13582 ({sk[2841], x22x, x16x, x501x, x549x, x535x, x345x}, x22086x);
	defparam lut_13582.LUT_SIZE = 7;
	defparam lut_13582.mask = 128'h37ff37ff3fff3fffaaaa8080aa008000;

	lut_sub lut_13587 ({sk[2842], x21x, x501x, x23x, x498x, x337x, x22086x}, x15939x);
	defparam lut_13587.LUT_SIZE = 7;
	defparam lut_13587.mask = 128'h37ff37ff3fff3fffbbbbbbffbfbfbfff;

	lut_sub lut_13592 ({sk[2843], x15838x, x15932x, x15933x, n_n1727, n_n1726}, x15942x);
	defparam lut_13592.LUT_SIZE = 6;
	defparam lut_13592.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_13598 ({sk[2844], i_9_, i_7_, i_8_, i_6_, x590x, x513x}, x15976x);
	defparam lut_13598.LUT_SIZE = 7;
	defparam lut_13598.mask = 128'h37ff37ff3fff3fff0035000000000000;

	lut_sub lut_13601 ({sk[2845], i_9_, i_1_, i_2_, i_0_, x572x, x135x}, x15981x);
	defparam lut_13601.LUT_SIZE = 7;
	defparam lut_13601.mask = 128'h37ff37ff3fff3fff5555555555557555;

	lut_sub lut_13604 ({sk[2846], x570x, x18x, x20x, x23x, x577x}, x15986x);
	defparam lut_13604.LUT_SIZE = 6;
	defparam lut_13604.mask = 64'h77ff77ff151515ff;

	lut_sub lut_13608 ({sk[2847], x15x, x24x, x18x, x590x, x584x}, x22279x);
	defparam lut_13608.LUT_SIZE = 6;
	defparam lut_13608.mask = 64'h77ff77fffac8c8c8;

	lut_sub lut_13613 ({sk[2848], x519x, x18x, x574x, x493x, x371x}, x22091x);
	defparam lut_13613.LUT_SIZE = 6;
	defparam lut_13613.mask = 64'h77ff77ffaa80aa00;

	lut_sub lut_13616 ({sk[2849], i_9_, i_7_, i_8_, i_6_, n_n455, n_n464}, x16068x);
	defparam lut_13616.LUT_SIZE = 7;
	defparam lut_13616.mask = 128'h37ff37ff3fff3fff0001010001000100;

	lut_sub lut_13621 ({sk[2850], i_9_, i_7_, i_8_, i_6_, n_n390, n_n535}, x22099x);
	defparam lut_13621.LUT_SIZE = 7;
	defparam lut_13621.mask = 128'h37ff37ff3fff3ffffeefeeefefffefef;

	lut_sub lut_13628 ({sk[2851], x10x, x545x, x23x, x523x, n_n4573, x121x}, x22100x);
	defparam lut_13628.LUT_SIZE = 7;
	defparam lut_13628.mask = 128'h37ff37ff3fff3fff8880888088800000;

	lut_sub lut_13633 ({sk[2852], i_9_, i_7_, i_8_, i_6_, n_n536, n_n535}, x16081x);
	defparam lut_13633.LUT_SIZE = 7;
	defparam lut_13633.mask = 128'h37ff37ff3fff3fff0101001000010000;

	lut_sub lut_13638 ({sk[2853], x25x, x22x, x14x, x594x, x551x, x526x}, x16141x);
	defparam lut_13638.LUT_SIZE = 7;
	defparam lut_13638.mask = 128'h37ff37ff3fff3fff000f777f555f777f;

	lut_sub lut_13643 ({sk[2854], x24x, x17x, x566x, x562x}, x16216x);
	defparam lut_13643.LUT_SIZE = 5;
	defparam lut_13643.mask = 32'h5f5f0537;

	lut_sub lut_13646 ({sk[2855], i_9_, i_7_, i_8_, i_6_, n_n260, n_n491}, x16220x);
	defparam lut_13646.LUT_SIZE = 7;
	defparam lut_13646.mask = 128'h37ff37ff3fff3fff0000000101010001;

	lut_sub lut_13651 ({sk[2856], i_9_, i_7_, i_8_, i_6_, x588x, x511x}, x16227x);
	defparam lut_13651.LUT_SIZE = 7;
	defparam lut_13651.mask = 128'h37ff37ff3fff3fff0035000000000000;

	lut_sub lut_13654 ({sk[2857], i_9_, i_7_, i_8_, i_6_, x565x, x575x}, x16230x);
	defparam lut_13654.LUT_SIZE = 7;
	defparam lut_13654.mask = 128'h37ff37ff3fff3fff3500000000000000;

	lut_sub lut_13657 ({sk[2858], x25x, x14x, x558x, x588x, x493x}, x16236x);
	defparam lut_13657.LUT_SIZE = 6;
	defparam lut_13657.mask = 64'h77ff77ff005f337f;

	lut_sub lut_13661 ({sk[2859], x19x, x516x, x506x, x529x, n_n1900, n_n1825}, x16316x);
	defparam lut_13661.LUT_SIZE = 7;
	defparam lut_13661.mask = 128'h37ff37ff3fff3fff777777777fffffff;

	lut_sub lut_13667 ({sk[2860], x19x, x20x, x23x, x491x, x536x, x569x}, x22329x);
	defparam lut_13667.LUT_SIZE = 7;
	defparam lut_13667.mask = 128'h37ff37ff3fff3fffffaaaaaac0808080;

	lut_sub lut_13672 ({sk[2861], x24x, x579x, n_n1824, x16304x, x22329x}, x16317x);
	defparam lut_13672.LUT_SIZE = 6;
	defparam lut_13672.mask = 64'h77ff77ffbfbfbfff;

	lut_sub lut_13677 ({sk[2862], x16318x, n_n1730, n_n1729, x15939x, x16316x, x16317x}, x22083x);
	defparam lut_13677.LUT_SIZE = 7;
	defparam lut_13677.mask = 128'h37ff37ff3fff3fff8000000000000000;

	lut_sub lut_13679 ({sk[2863], x22x, x14x, x588x, x23x, x505x, x511x}, x16348x);
	defparam lut_13679.LUT_SIZE = 7;
	defparam lut_13679.mask = 128'h37ff37ff3fff3fff000f333f555f777f;

	lut_sub lut_13683 ({sk[2864], i_9_, i_7_, i_8_, i_6_, n_n482, n_n325}, x16372x);
	defparam lut_13683.LUT_SIZE = 7;
	defparam lut_13683.mask = 128'h37ff37ff3fff3fff0010010010100000;

	lut_sub lut_13688 ({sk[2865], x22x, x21x, x14x, x588x, x570x, x520x}, x22306x);
	defparam lut_13688.LUT_SIZE = 7;
	defparam lut_13688.mask = 128'h37ff37ff3fff3fffff88f080f080f080;

	lut_sub lut_13693 ({sk[2866], x14x, x23x, x565x, x574x}, x16419x);
	defparam lut_13693.LUT_SIZE = 5;
	defparam lut_13693.mask = 32'h5f5f0357;

	lut_sub lut_13696 ({sk[2867], i_9_, x21x, n_n325, n_n522, n_n500, x518x}, x16421x);
	defparam lut_13696.LUT_SIZE = 7;
	defparam lut_13696.mask = 128'h37ff37ff3fff3fff0003003300570077;

	lut_sub lut_13701 ({sk[2868], x483x, x14x, x478x, x23x, x556x, x536x}, x22290x);
	defparam lut_13701.LUT_SIZE = 7;
	defparam lut_13701.mask = 128'h37ff37ff3fff3fffffff8800f0f08000;

	lut_sub lut_13706 ({sk[2869], i_9_, i_7_, i_8_, i_6_, n_n535, n_n195}, x16466x);
	defparam lut_13706.LUT_SIZE = 7;
	defparam lut_13706.mask = 128'h37ff37ff3fff3fff0100110101110110;

	lut_sub lut_13716 ({sk[2870], x16x, x20x, x557x, x498x}, x16550x);
	defparam lut_13716.LUT_SIZE = 5;
	defparam lut_13716.mask = 32'h5f5f0537;

	lut_sub lut_13719 ({sk[2871], x24x, x23x, x499x, x498x, x473x, x300x}, x22065x);
	defparam lut_13719.LUT_SIZE = 7;
	defparam lut_13719.mask = 128'h37ff37ff3fff3fffaaaa8888a0008000;

	lut_sub lut_13724 ({sk[2872], x521x, x13x, x539x, x544x, x11x}, x16566x);
	defparam lut_13724.LUT_SIZE = 6;
	defparam lut_13724.mask = 64'h77ff77ff111f11ff;

	lut_sub lut_13728 ({sk[2873], x21x, x13x, x544x, x482x, x23x, x494x}, x16567x);
	defparam lut_13728.LUT_SIZE = 7;
	defparam lut_13728.mask = 128'h37ff37ff3fff3fff00335f7f00ff5fff;

	lut_sub lut_13733 ({sk[2874], i_9_, n_n482, n_n455, n_n530, x378x}, x16586x);
	defparam lut_13733.LUT_SIZE = 6;
	defparam lut_13733.mask = 64'h77ff77ff55575557;

	lut_sub lut_13737 ({sk[2875], i_9_, i_1_, i_2_, i_0_, x502x, x528x}, x16639x);
	defparam lut_13737.LUT_SIZE = 7;
	defparam lut_13737.mask = 128'h37ff37ff3fff3fff0000000000000700;

	lut_sub lut_13740 ({sk[2876], x15x, x19x, x21x, x24x, x548x, x533x}, x16679x);
	defparam lut_13740.LUT_SIZE = 7;
	defparam lut_13740.mask = 128'h37ff37ff3fff3fff0555377755557777;

	lut_sub lut_13745 ({sk[2877], i_9_, i_7_, i_8_, i_6_, n_n535, n_n65}, x16680x);
	defparam lut_13745.LUT_SIZE = 7;
	defparam lut_13745.mask = 128'h37ff37ff3fff3fff0100000101001101;

	lut_sub lut_13752 ({sk[2878], i_9_, n_n524, n_n518, x562x, n_n65, x593x}, x16693x);
	defparam lut_13752.LUT_SIZE = 7;
	defparam lut_13752.mask = 128'h37ff37ff3fff3fff0000003313131333;

	lut_sub lut_13757 ({sk[2879], x570x, x12x, x491x, x537x, x76x}, x22072x);
	defparam lut_13757.LUT_SIZE = 6;
	defparam lut_13757.mask = 64'h77ff77ffaa80aa00;

	lut_sub lut_13760 ({sk[2880], x25x, x21x, x591x, x114x, x514x, n_n5181}, x22334x);
	defparam lut_13760.LUT_SIZE = 7;
	defparam lut_13760.mask = 128'h37ff37ff3fff3fffa0a0a00080808000;

	lut_sub lut_13765 ({sk[2881], x18x, x23x, x513x, x527x, x528x}, x16709x);
	defparam lut_13765.LUT_SIZE = 6;
	defparam lut_13765.mask = 64'h77ff77ff000f777f;

	lut_sub lut_13769 ({sk[2882], x538x, x510x, x18x, x23x, x590x, x584x}, x16740x);
	defparam lut_13769.LUT_SIZE = 7;
	defparam lut_13769.mask = 128'h37ff37ff3fff3fff035703ff03ff03ff;

	lut_sub lut_13774 ({sk[2883], x25x, x509x, x18x, x513x, x493x, n_n5043}, x22070x);
	defparam lut_13774.LUT_SIZE = 7;
	defparam lut_13774.mask = 128'h37ff37ff3fff3fffaa88aa00a080a000;

	lut_sub lut_13779 ({sk[2884], x117x, x12968x, x12969x, n_n5335, n_n5334, n_n5333}, x22066x);
	defparam lut_13779.LUT_SIZE = 7;
	defparam lut_13779.mask = 128'h37ff37ff3fff3fff8000000000000000;

	lut_sub lut_13781 ({sk[2885], x21x, x17x, x522x, x512x}, x16816x);
	defparam lut_13781.LUT_SIZE = 5;
	defparam lut_13781.mask = 32'h5f5f0357;

	lut_sub lut_13784 ({sk[2886], x21x, x17x, x506x, x531x, x527x, x528x}, x16818x);
	defparam lut_13784.LUT_SIZE = 7;
	defparam lut_13784.mask = 128'h37ff37ff3fff3fff000077ff0f0f7fff;

	lut_sub lut_13789 ({sk[2887], x16496x, x16497x, x16516x, n_n2098, n_n2099}, x16826x);
	defparam lut_13789.LUT_SIZE = 6;
	defparam lut_13789.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_13795 ({sk[2888], n_n2104, n_n2105, n_n2103, n_n2092, n_n2091, x16805x}, x22058x);
	defparam lut_13795.LUT_SIZE = 7;
	defparam lut_13795.mask = 128'h37ff37ff3fff3fff8000000000000000;

	lut_sub lut_13797 ({sk[2889], x15x, x21x, x20x, x577x, x567x, x343x}, x22163x);
	defparam lut_13797.LUT_SIZE = 7;
	defparam lut_13797.mask = 128'h37ff37ff3fff3fffaa888888a0808080;


endmodule