module bigkey (
	Pstart_0_, Pkey_255_, Pkey_254_, Pkey_253_, Pkey_252_, Pkey_251_, Pkey_250_, Pkey_249_, 
	Pkey_248_, Pkey_247_, Pkey_246_, Pkey_245_, Pkey_244_, Pkey_243_, Pkey_242_, Pkey_241_, Pkey_240_, Pkey_239_, 
	Pkey_238_, Pkey_237_, Pkey_236_, Pkey_235_, Pkey_234_, Pkey_233_, Pkey_232_, Pkey_231_, Pkey_230_, Pkey_229_, 
	Pkey_228_, Pkey_227_, Pkey_226_, Pkey_225_, Pkey_224_, Pkey_223_, Pkey_222_, Pkey_221_, Pkey_220_, Pkey_219_, 
	Pkey_218_, Pkey_217_, Pkey_216_, Pkey_215_, Pkey_214_, Pkey_213_, Pkey_212_, Pkey_211_, Pkey_210_, Pkey_209_, 
	Pkey_208_, Pkey_207_, Pkey_206_, Pkey_205_, Pkey_204_, Pkey_203_, Pkey_202_, Pkey_201_, Pkey_200_, Pkey_199_, 
	Pkey_198_, Pkey_197_, Pkey_196_, Pkey_195_, Pkey_194_, Pkey_193_, Pkey_192_, Pkey_191_, Pkey_190_, Pkey_189_, 
	Pkey_188_, Pkey_187_, Pkey_186_, Pkey_185_, Pkey_184_, Pkey_183_, Pkey_182_, Pkey_181_, Pkey_180_, Pkey_179_, 
	Pkey_178_, Pkey_177_, Pkey_176_, Pkey_175_, Pkey_174_, Pkey_173_, Pkey_172_, Pkey_171_, Pkey_170_, Pkey_169_, 
	Pkey_168_, Pkey_167_, Pkey_166_, Pkey_165_, Pkey_164_, Pkey_163_, Pkey_162_, Pkey_161_, Pkey_160_, Pkey_159_, 
	Pkey_158_, Pkey_157_, Pkey_156_, Pkey_155_, Pkey_154_, Pkey_153_, Pkey_152_, Pkey_151_, Pkey_150_, Pkey_149_, 
	Pkey_148_, Pkey_147_, Pkey_146_, Pkey_145_, Pkey_144_, Pkey_143_, Pkey_142_, Pkey_141_, Pkey_140_, Pkey_139_, 
	Pkey_138_, Pkey_137_, Pkey_136_, Pkey_135_, Pkey_134_, Pkey_133_, Pkey_132_, Pkey_131_, Pkey_130_, Pkey_129_, 
	Pkey_128_, Pkey_127_, Pkey_126_, Pkey_125_, Pkey_124_, Pkey_123_, Pkey_122_, Pkey_121_, Pkey_120_, Pkey_119_, 
	Pkey_118_, Pkey_117_, Pkey_116_, Pkey_115_, Pkey_114_, Pkey_113_, Pkey_112_, Pkey_111_, Pkey_110_, Pkey_109_, 
	Pkey_108_, Pkey_107_, Pkey_106_, Pkey_105_, Pkey_104_, Pkey_103_, Pkey_102_, Pkey_101_, Pkey_100_, Pkey_99_, 
	Pkey_98_, Pkey_97_, Pkey_96_, Pkey_95_, Pkey_94_, Pkey_93_, Pkey_92_, Pkey_91_, Pkey_90_, Pkey_89_, 
	Pkey_88_, Pkey_87_, Pkey_86_, Pkey_85_, Pkey_84_, Pkey_83_, Pkey_82_, Pkey_81_, Pkey_80_, Pkey_79_, 
	Pkey_78_, Pkey_77_, Pkey_76_, Pkey_75_, Pkey_74_, Pkey_73_, Pkey_72_, Pkey_71_, Pkey_70_, Pkey_69_, 
	Pkey_68_, Pkey_67_, Pkey_66_, Pkey_65_, Pkey_64_, Pkey_63_, Pkey_62_, Pkey_61_, Pkey_60_, Pkey_59_, 
	Pkey_58_, Pkey_57_, Pkey_56_, Pkey_55_, Pkey_54_, Pkey_53_, Pkey_52_, Pkey_51_, Pkey_50_, Pkey_49_, 
	Pkey_48_, Pkey_47_, Pkey_46_, Pkey_45_, Pkey_44_, Pkey_43_, Pkey_42_, Pkey_41_, Pkey_40_, Pkey_39_, 
	Pkey_38_, Pkey_37_, Pkey_36_, Pkey_35_, Pkey_34_, Pkey_33_, Pkey_32_, Pkey_31_, Pkey_30_, Pkey_29_, 
	Pkey_28_, Pkey_27_, Pkey_26_, Pkey_25_, Pkey_24_, Pkey_23_, Pkey_22_, Pkey_21_, Pkey_20_, Pkey_19_, 
	Pkey_18_, Pkey_17_, Pkey_16_, Pkey_15_, Pkey_14_, Pkey_13_, Pkey_12_, Pkey_11_, Pkey_10_, Pkey_9_, 
	Pkey_8_, Pkey_7_, Pkey_6_, Pkey_5_, Pkey_4_, Pkey_3_, Pkey_2_, Pkey_1_, Pkey_0_, Pencrypt_0_, 
	Pcount_3_, Pcount_2_, Pcount_1_, Pcount_0_, PCLK, Pnew_count_3_, Pnew_count_2_, Pnew_count_1_, Pnew_count_0_, Pdata_ready_0_, 
	PKSi_191_, PKSi_190_, PKSi_189_, PKSi_188_, PKSi_187_, PKSi_186_, PKSi_185_, PKSi_184_, PKSi_183_, PKSi_182_, 
	PKSi_181_, PKSi_180_, PKSi_179_, PKSi_178_, PKSi_177_, PKSi_176_, PKSi_175_, PKSi_174_, PKSi_173_, PKSi_172_, 
	PKSi_171_, PKSi_170_, PKSi_169_, PKSi_168_, PKSi_167_, PKSi_166_, PKSi_165_, PKSi_164_, PKSi_163_, PKSi_162_, 
	PKSi_161_, PKSi_160_, PKSi_159_, PKSi_158_, PKSi_157_, PKSi_156_, PKSi_155_, PKSi_154_, PKSi_153_, PKSi_152_, 
	PKSi_151_, PKSi_150_, PKSi_149_, PKSi_148_, PKSi_147_, PKSi_146_, PKSi_145_, PKSi_144_, PKSi_143_, PKSi_142_, 
	PKSi_141_, PKSi_140_, PKSi_139_, PKSi_138_, PKSi_137_, PKSi_136_, PKSi_135_, PKSi_134_, PKSi_133_, PKSi_132_, 
	PKSi_131_, PKSi_130_, PKSi_129_, PKSi_128_, PKSi_127_, PKSi_126_, PKSi_125_, PKSi_124_, PKSi_123_, PKSi_122_, 
	PKSi_121_, PKSi_120_, PKSi_119_, PKSi_118_, PKSi_117_, PKSi_116_, PKSi_115_, PKSi_114_, PKSi_113_, PKSi_112_, 
	PKSi_111_, PKSi_110_, PKSi_109_, PKSi_108_, PKSi_107_, PKSi_106_, PKSi_105_, PKSi_104_, PKSi_103_, PKSi_102_, 
	PKSi_101_, PKSi_100_, PKSi_99_, PKSi_98_, PKSi_97_, PKSi_96_, PKSi_95_, PKSi_94_, PKSi_93_, PKSi_92_, 
	PKSi_91_, PKSi_90_, PKSi_89_, PKSi_88_, PKSi_87_, PKSi_86_, PKSi_85_, PKSi_84_, PKSi_83_, PKSi_82_, 
	PKSi_81_, PKSi_80_, PKSi_79_, PKSi_78_, PKSi_77_, PKSi_76_, PKSi_75_, PKSi_74_, PKSi_73_, PKSi_72_, 
	PKSi_71_, PKSi_70_, PKSi_69_, PKSi_68_, PKSi_67_, PKSi_66_, PKSi_65_, PKSi_64_, PKSi_63_, PKSi_62_, 
	PKSi_61_, PKSi_60_, PKSi_59_, PKSi_58_, PKSi_57_, PKSi_56_, PKSi_55_, PKSi_54_, PKSi_53_, PKSi_52_, 
	PKSi_51_, PKSi_50_, PKSi_49_, PKSi_48_, PKSi_47_, PKSi_46_, PKSi_45_, PKSi_44_, PKSi_43_, PKSi_42_, 
	PKSi_41_, PKSi_40_, PKSi_39_, PKSi_38_, PKSi_37_, PKSi_36_, PKSi_35_, PKSi_34_, PKSi_33_, PKSi_32_, 
	PKSi_31_, PKSi_30_, PKSi_29_, PKSi_28_, PKSi_27_, PKSi_26_, PKSi_25_, PKSi_24_, PKSi_23_, PKSi_22_, 
	PKSi_21_, PKSi_20_, PKSi_19_, PKSi_18_, PKSi_17_, PKSi_16_, PKSi_15_, PKSi_14_, PKSi_13_, PKSi_12_, 
	PKSi_11_, PKSi_10_, PKSi_9_, PKSi_8_, PKSi_7_, PKSi_6_, PKSi_5_, PKSi_4_, PKSi_3_, PKSi_2_, 
	PKSi_1_, PKSi_0_);

input Pstart_0_, Pkey_255_, Pkey_254_, Pkey_253_, Pkey_252_, Pkey_251_, Pkey_250_, Pkey_249_, Pkey_248_, Pkey_247_, Pkey_246_, Pkey_245_, Pkey_244_, Pkey_243_, Pkey_242_, Pkey_241_, Pkey_240_, Pkey_239_, Pkey_238_, Pkey_237_, Pkey_236_, Pkey_235_, Pkey_234_, Pkey_233_, Pkey_232_, Pkey_231_, Pkey_230_, Pkey_229_, Pkey_228_, Pkey_227_, Pkey_226_, Pkey_225_, Pkey_224_, Pkey_223_, Pkey_222_, Pkey_221_, Pkey_220_, Pkey_219_, Pkey_218_, Pkey_217_, Pkey_216_, Pkey_215_, Pkey_214_, Pkey_213_, Pkey_212_, Pkey_211_, Pkey_210_, Pkey_209_, Pkey_208_, Pkey_207_, Pkey_206_, Pkey_205_, Pkey_204_, Pkey_203_, Pkey_202_, Pkey_201_, Pkey_200_, Pkey_199_, Pkey_198_, Pkey_197_, Pkey_196_, Pkey_195_, Pkey_194_, Pkey_193_, Pkey_192_, Pkey_191_, Pkey_190_, Pkey_189_, Pkey_188_, Pkey_187_, Pkey_186_, Pkey_185_, Pkey_184_, Pkey_183_, Pkey_182_, Pkey_181_, Pkey_180_, Pkey_179_, Pkey_178_, Pkey_177_, Pkey_176_, Pkey_175_, Pkey_174_, Pkey_173_, Pkey_172_, Pkey_171_, Pkey_170_, Pkey_169_, Pkey_168_, Pkey_167_, Pkey_166_, Pkey_165_, Pkey_164_, Pkey_163_, Pkey_162_, Pkey_161_, Pkey_160_, Pkey_159_, Pkey_158_, Pkey_157_, Pkey_156_, Pkey_155_, Pkey_154_, Pkey_153_, Pkey_152_, Pkey_151_, Pkey_150_, Pkey_149_, Pkey_148_, Pkey_147_, Pkey_146_, Pkey_145_, Pkey_144_, Pkey_143_, Pkey_142_, Pkey_141_, Pkey_140_, Pkey_139_, Pkey_138_, Pkey_137_, Pkey_136_, Pkey_135_, Pkey_134_, Pkey_133_, Pkey_132_, Pkey_131_, Pkey_130_, Pkey_129_, Pkey_128_, Pkey_127_, Pkey_126_, Pkey_125_, Pkey_124_, Pkey_123_, Pkey_122_, Pkey_121_, Pkey_120_, Pkey_119_, Pkey_118_, Pkey_117_, Pkey_116_, Pkey_115_, Pkey_114_, Pkey_113_, Pkey_112_, Pkey_111_, Pkey_110_, Pkey_109_, Pkey_108_, Pkey_107_, Pkey_106_, Pkey_105_, Pkey_104_, Pkey_103_, Pkey_102_, Pkey_101_, Pkey_100_, Pkey_99_, Pkey_98_, Pkey_97_, Pkey_96_, Pkey_95_, Pkey_94_, Pkey_93_, Pkey_92_, Pkey_91_, Pkey_90_, Pkey_89_, Pkey_88_, Pkey_87_, Pkey_86_, Pkey_85_, Pkey_84_, Pkey_83_, Pkey_82_, Pkey_81_, Pkey_80_, Pkey_79_, Pkey_78_, Pkey_77_, Pkey_76_, Pkey_75_, Pkey_74_, Pkey_73_, Pkey_72_, Pkey_71_, Pkey_70_, Pkey_69_, Pkey_68_, Pkey_67_, Pkey_66_, Pkey_65_, Pkey_64_, Pkey_63_, Pkey_62_, Pkey_61_, Pkey_60_, Pkey_59_, Pkey_58_, Pkey_57_, Pkey_56_, Pkey_55_, Pkey_54_, Pkey_53_, Pkey_52_, Pkey_51_, Pkey_50_, Pkey_49_, Pkey_48_, Pkey_47_, Pkey_46_, Pkey_45_, Pkey_44_, Pkey_43_, Pkey_42_, Pkey_41_, Pkey_40_, Pkey_39_, Pkey_38_, Pkey_37_, Pkey_36_, Pkey_35_, Pkey_34_, Pkey_33_, Pkey_32_, Pkey_31_, Pkey_30_, Pkey_29_, Pkey_28_, Pkey_27_, Pkey_26_, Pkey_25_, Pkey_24_, Pkey_23_, Pkey_22_, Pkey_21_, Pkey_20_, Pkey_19_, Pkey_18_, Pkey_17_, Pkey_16_, Pkey_15_, Pkey_14_, Pkey_13_, Pkey_12_, Pkey_11_, Pkey_10_, Pkey_9_, Pkey_8_, Pkey_7_, Pkey_6_, Pkey_5_, Pkey_4_, Pkey_3_, Pkey_2_, Pkey_1_, Pkey_0_, Pencrypt_0_, Pcount_3_, Pcount_2_, Pcount_1_, Pcount_0_, PCLK;

output Pnew_count_3_, Pnew_count_2_, Pnew_count_1_, Pnew_count_0_, Pdata_ready_0_, PKSi_191_, PKSi_190_, PKSi_189_, PKSi_188_, PKSi_187_, PKSi_186_, PKSi_185_, PKSi_184_, PKSi_183_, PKSi_182_, PKSi_181_, PKSi_180_, PKSi_179_, PKSi_178_, PKSi_177_, PKSi_176_, PKSi_175_, PKSi_174_, PKSi_173_, PKSi_172_, PKSi_171_, PKSi_170_, PKSi_169_, PKSi_168_, PKSi_167_, PKSi_166_, PKSi_165_, PKSi_164_, PKSi_163_, PKSi_162_, PKSi_161_, PKSi_160_, PKSi_159_, PKSi_158_, PKSi_157_, PKSi_156_, PKSi_155_, PKSi_154_, PKSi_153_, PKSi_152_, PKSi_151_, PKSi_150_, PKSi_149_, PKSi_148_, PKSi_147_, PKSi_146_, PKSi_145_, PKSi_144_, PKSi_143_, PKSi_142_, PKSi_141_, PKSi_140_, PKSi_139_, PKSi_138_, PKSi_137_, PKSi_136_, PKSi_135_, PKSi_134_, PKSi_133_, PKSi_132_, PKSi_131_, PKSi_130_, PKSi_129_, PKSi_128_, PKSi_127_, PKSi_126_, PKSi_125_, PKSi_124_, PKSi_123_, PKSi_122_, PKSi_121_, PKSi_120_, PKSi_119_, PKSi_118_, PKSi_117_, PKSi_116_, PKSi_115_, PKSi_114_, PKSi_113_, PKSi_112_, PKSi_111_, PKSi_110_, PKSi_109_, PKSi_108_, PKSi_107_, PKSi_106_, PKSi_105_, PKSi_104_, PKSi_103_, PKSi_102_, PKSi_101_, PKSi_100_, PKSi_99_, PKSi_98_, PKSi_97_, PKSi_96_, PKSi_95_, PKSi_94_, PKSi_93_, PKSi_92_, PKSi_91_, PKSi_90_, PKSi_89_, PKSi_88_, PKSi_87_, PKSi_86_, PKSi_85_, PKSi_84_, PKSi_83_, PKSi_82_, PKSi_81_, PKSi_80_, PKSi_79_, PKSi_78_, PKSi_77_, PKSi_76_, PKSi_75_, PKSi_74_, PKSi_73_, PKSi_72_, PKSi_71_, PKSi_70_, PKSi_69_, PKSi_68_, PKSi_67_, PKSi_66_, PKSi_65_, PKSi_64_, PKSi_63_, PKSi_62_, PKSi_61_, PKSi_60_, PKSi_59_, PKSi_58_, PKSi_57_, PKSi_56_, PKSi_55_, PKSi_54_, PKSi_53_, PKSi_52_, PKSi_51_, PKSi_50_, PKSi_49_, PKSi_48_, PKSi_47_, PKSi_46_, PKSi_45_, PKSi_44_, PKSi_43_, PKSi_42_, PKSi_41_, PKSi_40_, PKSi_39_, PKSi_38_, PKSi_37_, PKSi_36_, PKSi_35_, PKSi_34_, PKSi_33_, PKSi_32_, PKSi_31_, PKSi_30_, PKSi_29_, PKSi_28_, PKSi_27_, PKSi_26_, PKSi_25_, PKSi_24_, PKSi_23_, PKSi_22_, PKSi_21_, PKSi_20_, PKSi_19_, PKSi_18_, PKSi_17_, PKSi_16_, PKSi_15_, PKSi_14_, PKSi_13_, PKSi_12_, PKSi_11_, PKSi_10_, PKSi_9_, PKSi_8_, PKSi_7_, PKSi_6_, PKSi_5_, PKSi_4_, PKSi_3_, PKSi_2_, PKSi_1_, PKSi_0_;

wire n15, n13, n11, n1741, n16, n17, n18, n19, n20, n21, N_N2862, n22, N_N2863, n23, N_N2864, n24, N_N2866, n25, N_N2867, n26, N_N2868, n27, N_N2869, n28, N_N2870, n29, N_N2871, n30, N_N2872, n31, N_N2873, n32, N_N2874, n33, N_N2875, n34, N_N2876, n35, N_N2878, n36, N_N2880, n37, N_N2882, n38, N_N2883, n39, N_N2884, n40, N_N2886, n41, N_N2887, n42, N_N2888, n43, N_N2890, n44, N_N2891, n45, N_N2892, n46, N_N2893, n47, N_N2894, n48, N_N2895, n49, N_N2896, n50, N_N2897, n51, N_N2898, n52, N_N2900, n53, N_N2901, n54, N_N2902, n55, N_N2903, n56, N_N2904, n57, N_N2905, n58, N_N2906, n59, N_N2907, n60, N_N2908, n61, N_N2910, n62, N_N2911, n63, N_N2912, n64, N_N2913, n65, N_N2914, n66, N_N2915, n67, N_N2916, n68, N_N2918, n69, N_N2919, n70, N_N2920, n71, N_N2922, n72, N_N2923, n73, N_N2924, n74, N_N2925, n75, N_N2926, n76, N_N2927, n77, N_N2928, n78, N_N2929, n79, N_N2930, n80, N_N2932, n81, N_N2933, n82, N_N2934, n83, N_N2935, n84, N_N2936, n85, N_N2937, n86, N_N2938, n87, N_N2939, n88, N_N2940, n89, N_N2941, n90, N_N2942, n91, N_N2944, n92, N_N2946, n93, N_N2947, n94, N_N2948, n95, N_N2949, n96, N_N2951, n97, N_N2952, n98, N_N2953, n99, N_N2955, n100, N_N2956, n101, N_N2957, n102, N_N2958, n103, N_N2959, n104, N_N2960, n105, N_N2961, n106, N_N2962, n107, N_N2963, n108, N_N2965, n109, N_N2966, n110, N_N2967, n111, N_N2968, n112, N_N2969, n113, N_N2970, n114, N_N2971, n115, N_N2972, n116, N_N2973, n117, N_N2974, n118, N_N2975, n119, N_N2977, n120, N_N2978, n121, N_N2979, n122, N_N2980, n123, N_N2981, n124, N_N2983, n125, N_N2984, n126, N_N2985, n127, N_N2987, n128, N_N2988, n129, N_N2989, n130, N_N2990, n131, N_N2991, n132, N_N2992, n133, N_N2733, n134, N_N2734, n135, N_N2735, n136, N_N2736, n137, N_N2738, n138, N_N2739, n139, N_N2740, n140, N_N2742, n141, N_N2743, n142, N_N2744, n143, N_N2745, n144, N_N2747, n145, N_N2748, n146, N_N2750, n147, N_N2751, n148, N_N2752, n149, N_N2753, n150, N_N2754, n151, N_N2755, n152, N_N2756, n153, N_N2758, n154, N_N2759, n155, N_N2760, n156, N_N2761, n157, N_N2762, n158, N_N2763, n159, N_N2764, n160, N_N2765, n161, N_N2766, n162, N_N2767, n163, N_N2768, n164, N_N2769, n165, N_N2771, n166, N_N2772, n167, N_N2773, n168, N_N2775, n169, N_N2776, n170, N_N2777, n171, N_N2778, n172, N_N2780, n173, N_N2781, n174, N_N2782, n175, N_N2783, n176, N_N2784, n177, N_N2785, n178, N_N2786, n179, N_N2787, n180, N_N2788, n181, N_N2790, n182, N_N2791, n183, N_N2792, n184, N_N2793, n185, N_N2794, n186, N_N2795, n187, N_N2796, n188, N_N2797, n189, N_N2798, n190, N_N2799, n191, N_N2800, n192, N_N2801, n193, N_N2803, n194, N_N2804, n195, N_N2805, n196, N_N2807, n197, N_N2808, n198, N_N2809, n199, N_N2810, n200, N_N2812, n201, N_N2813, n202, N_N2814, n203, N_N2815, n204, N_N2816, n205, N_N2817, n206, N_N2818, n207, N_N2819, n208, N_N2820, n209, N_N2822, n210, N_N2823, n211, N_N2824, n212, N_N2825, n213, N_N2826, n214, N_N2827, n215, N_N2828, n216, N_N2829, n217, N_N2830, n218, N_N2831, n219, N_N2832, n220, N_N2833, n221, N_N2835, n222, N_N2836, n223, N_N2837, n224, N_N2839, n225, N_N2840, n226, N_N2841, n227, N_N2842, n228, N_N2844, n229, N_N2845, n230, N_N2846, n231, N_N2847, n232, N_N2848, n233, N_N2849, n234, N_N2850, n235, N_N2851, n236, N_N2852, n237, N_N2854, n238, N_N2855, n239, N_N2856, n240, N_N2857, n241, N_N2858, n242, N_N2859, n243, N_N2860, n244, N_N2861, n248, n249, n246, n245, n251, n252, n250, n255, n256, n258, n259, n261, n262, n264, n265, n267, n268, n270, n271, n273, n274, n276, n277, n279, n280, n282, n283, n285, n286, n288, n289, n291, n292, n294, n295, n297, n298, n300, n301, n303, n304, n306, n307, n309, n310, n312, n313, n315, n316, n318, n319, n321, n322, n324, n325, n327, n328, n330, n331, n333, n334, n336, n337, n339, n340, n342, n343, n345, n346, n348, n349, n351, n352, n354, n355, n357, n358, n360, n361, n363, n364, n366, n367, n369, n370, n372, n373, n375, n376, n378, n379, n381, n382, n384, n385, n387, n388, n389, n390, n392, n393, n395, n396, n398, n399, n401, n402, n404, n405, n407, n408, n410, n411, n413, n414, n416, n417, n419, n420, n422, n423, n425, n426, n428, n429, n431, n432, n434, n435, n437, n438, n440, n441, n443, n444, n446, n447, n449, n450, n452, n453, n455, n456, n458, n459, n461, n462, n464, n465, n467, n468, n470, n471, n473, n474, n476, n477, n479, n480, n482, n483, n485, n486, n488, n489, n491, n492, n494, n495, n497, n498, n500, n501, n503, n504, n506, n507, n509, n510, n512, n513, n515, n516, n518, n519, n521, n522, n524, n525, n527, n528, n530, n531, n533, n534, n536, n537, n539, n540, n542, n543, n545, n546, n548, n549, n551, n552, n554, n555, n556, n557, n559, n560, n562, n563, n565, n566, n568, n569, n571, n572, n574, n575, n577, n578, n580, n581, n583, n584, n586, n587, n589, n590, n592, n593, n595, n596, n598, n599, n601, n602, n604, n605, n607, n608, n610, n611, n613, n614, n616, n617, n619, n620, n622, n623, n625, n626, n628, n629, n631, n632, n634, n635, n637, n638, n640, n641, n643, n644, n646, n647, n649, n650, n652, n653, n655, n656, n658, n659, n661, n662, n664, n665, n667, n668, n670, n671, n673, n674, n676, n677, n679, n680, n682, n683, n685, n686, n688, n689, n691, n692, n694, n695, n697, n698, n700, n701, n703, n704, n706, n707, n709, n710, n712, n713, n715, n716, n718, n719, n721, n722, n724, n725, n727, n728, n730, n731, n733, n734, n736, n737, n739, n740, n742, n743, n745, n746, n748, n749, n751, n752, n754, n755, n757, n758, n760, n761, n763, n764, n766, n767, n769, n770, n772, n773, n775, n776, n778, n779, n781, n782, n784, n785, n787, n788, n790, n791, n793, n794, n796, n797, n799, n800, n802, n803, n805, n806, n808, n809, n811, n812, n814, n815, n817, n818, n820, n821, n823, n824, n826, n827, n829, n830, n832, n833, n835, n836, n838, n839, n841, n842, n844, n845, n847, n848, n850, n851, n853, n854, n856, n857, n859, n860, n862, n863, n865, n866, n868, n869, n871, n872, n874, n875, n877, n878, n880, n881, n883, n884, n886, n887, n889, n890, n892, n893, n895, n896, n898, n899, n901, n902, n904, n905, n907, n908, n910, n911, n913, n914, n916, n917, n919, n920, n922, n923, n925, n924, n929, n928, n930, n934, n935, n939, n938, n937, n940, n942, n944, n946, n948, n950, n952, n954, n956, n958, n960, n962, n964, n966, n968, n970, n972, n974, n976, n978, n980, n982, n984, n986, n988, n990, n992, n994, n996, n998, n1000, n1002, n1004, n1006, n1008, n1010, n1012, n1014, n1016, n1018, n1020, n1022, n1024, n1026, n1028, n1030, n1032, n1034, n1036, n1038, n1040, n1042, n1044, n1046, n1048, n1050, n1052, n1054, n1056, n1058, n1060, n1062, n1064, n1066, n1068, n1070, n1072, n1074, n1076, n1078, n1080, n1082, n1084, n1086, n1088, n1090, n1092, n1094, n1096, n1098, n1100, n1102, n1104, n1106, n1108, n1110, n1112, n1114, n1116, n1118, n1120, n1122, n1124, n1126, n1128, n1130, n1132, n1134, n1136, n1138, n1140, n1142, n1144, n1146, n1148, n1150, n1152, n1154, n1156, n1158, n1160, n1162, n1167, n1166, n1170, n1285, n1284, n1286, n1287, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1740, n1744, n1746, n1748, n1750, n1752, n1754, n1756, n1758, n1760, n1762, n1764, n1766, n1768, n1770, n1772, n1774, n1776, n1778, n1780, n1782, n1784, n1786, n1788, n1790, n1792, n1794, n1796, n1798, n1800, n1802, n1804, n1806, n1808, n1810, n1812, n1814, n1816, n1818, n1820, n1822, n1824, n1826, n1828, n1830, n1832, n1834, n1836, n1838, n1840, n1842, n1844, n1846, n1848, n1850, n1852, n1854, n1856, n1858, n1860, n1862, n1864, n1866, n1868, n1870, n1872, n1874, n1876, n1878, n1880, n1882, n1884, n1886, n1888, n1890, n1892, n1894, n1896, n1898, n1900, n1902, n1904, n1906, n1908, n1910, n1912, n1914, n1916, n1918, n1920, n1922, n1924, n1926, n1928, n1930, n1932, n1934, n1936, n1938, n1940, n1942, n1944, n1946, n1948, n1950, n1952, n1954, n1956, n1958, n1960, n1962, n1964, n1966, n1967, n1968;

reg PKSi_79_, PKSi_92_, wire333, N_N2737, PKSi_75_, PKSi_84_, N_N2741, PKSi_82_, PKSi_93_, PKSi_85_, N_N2746, PKSi_73_, N_N2749, PKSi_80_, PKSi_72_, PKSi_94_, PKSi_86_, PKSi_74_, PKSi_83_, N_N2757, PKSi_89_, PKSi_91_, PKSi_81_, PKSi_77_, PKSi_87_, PKSi_78_, PKSi_95_, PKSi_76_, PKSi_55_, PKSi_68_, PKSi_64_, N_N2770, PKSi_51_, PKSi_60_, N_N2774, PKSi_58_, PKSi_69_, PKSi_61_, N_N2779, PKSi_49_, PKSi_66_, PKSi_56_, PKSi_48_, PKSi_70_, PKSi_62_, PKSi_50_, PKSi_59_, N_N2789, PKSi_65_, PKSi_67_, PKSi_57_, PKSi_53_, PKSi_63_, PKSi_54_, PKSi_71_, PKSi_52_, PKSi_31_, PKSi_44_, PKSi_40_, N_N2802, PKSi_27_, PKSi_36_, N_N2806, PKSi_34_, PKSi_45_, PKSi_37_, N_N2811, PKSi_25_, PKSi_42_, PKSi_32_, PKSi_24_, PKSi_46_, PKSi_38_, PKSi_26_, PKSi_35_, N_N2821, PKSi_41_, PKSi_43_, PKSi_33_, PKSi_29_, PKSi_39_, PKSi_30_, PKSi_47_, PKSi_28_, PKSi_7_, PKSi_20_, PKSi_16_, N_N2834, PKSi_3_, PKSi_12_, N_N2838, PKSi_10_, PKSi_21_, PKSi_13_, N_N2843, PKSi_1_, PKSi_18_, PKSi_8_, PKSi_0_, PKSi_22_, PKSi_14_, PKSi_2_, PKSi_11_, N_N2853, PKSi_17_, PKSi_19_, PKSi_9_, PKSi_5_, PKSi_15_, PKSi_6_, PKSi_23_, PKSi_4_, PKSi_183_, PKSi_173_, N_N2865, PKSi_185_, PKSi_169_, PKSi_176_, PKSi_188_, wire253, PKSi_179_, PKSi_172_, PKSi_186_, PKSi_177_, PKSi_180_, N_N2877, N_N2879, N_N2881, PKSi_175_, PKSi_182_, N_N2885, PKSi_171_, PKSi_189_, N_N2889, PKSi_184_, PKSi_178_, wire234, PKSi_170_, PKSi_174_, PKSi_190_, PKSi_159_, PKSi_149_, N_N2899, PKSi_161_, PKSi_145_, PKSi_152_, PKSi_164_, PKSi_157_, PKSi_155_, PKSi_148_, PKSi_162_, N_N2909, PKSi_156_, PKSi_153_, PKSi_163_, PKSi_144_, PKSi_151_, PKSi_158_, N_N2917, PKSi_147_, PKSi_165_, N_N2921, PKSi_160_, PKSi_154_, PKSi_167_, PKSi_146_, PKSi_150_, PKSi_166_, PKSi_135_, PKSi_125_, N_N2931, PKSi_137_, PKSi_121_, PKSi_128_, PKSi_140_, PKSi_133_, PKSi_131_, PKSi_124_, PKSi_138_, PKSi_129_, PKSi_132_, N_N2943, N_N2945, PKSi_120_, PKSi_127_, PKSi_134_, N_N2950, PKSi_123_, PKSi_141_, N_N2954, PKSi_136_, PKSi_130_, wire282, PKSi_122_, PKSi_126_, PKSi_142_, PKSi_111_, PKSi_101_, N_N2964, PKSi_113_, PKSi_97_, PKSi_104_, PKSi_116_, PKSi_109_, PKSi_107_, PKSi_100_, PKSi_114_, PKSi_105_, PKSi_108_, N_N2976, PKSi_115_, PKSi_96_, PKSi_103_, PKSi_110_, N_N2982, PKSi_99_, PKSi_117_, N_N2986, PKSi_112_, PKSi_106_, PKSi_119_, PKSi_98_, PKSi_102_, PKSi_118_;

always  @(posedge PCLK)
	PKSi_79_<=N_N2733;

 always  @(posedge PCLK)
	PKSi_92_<=N_N2734;

 always  @(posedge PCLK)
	wire333<=N_N2735;

 always  @(posedge PCLK)
	N_N2737<=N_N2736;

 always  @(posedge PCLK)
	PKSi_75_<=N_N2738;

 always  @(posedge PCLK)
	PKSi_84_<=N_N2739;

 always  @(posedge PCLK)
	N_N2741<=N_N2740;

 always  @(posedge PCLK)
	PKSi_82_<=N_N2742;

 always  @(posedge PCLK)
	PKSi_93_<=N_N2743;

 always  @(posedge PCLK)
	PKSi_85_<=N_N2744;

 always  @(posedge PCLK)
	N_N2746<=N_N2745;

 always  @(posedge PCLK)
	PKSi_73_<=N_N2747;

 always  @(posedge PCLK)
	N_N2749<=N_N2748;

 always  @(posedge PCLK)
	PKSi_80_<=N_N2750;

 always  @(posedge PCLK)
	PKSi_72_<=N_N2751;

 always  @(posedge PCLK)
	PKSi_94_<=N_N2752;

 always  @(posedge PCLK)
	PKSi_86_<=N_N2753;

 always  @(posedge PCLK)
	PKSi_74_<=N_N2754;

 always  @(posedge PCLK)
	PKSi_83_<=N_N2755;

 always  @(posedge PCLK)
	N_N2757<=N_N2756;

 always  @(posedge PCLK)
	PKSi_89_<=N_N2758;

 always  @(posedge PCLK)
	PKSi_91_<=N_N2759;

 always  @(posedge PCLK)
	PKSi_81_<=N_N2760;

 always  @(posedge PCLK)
	PKSi_77_<=N_N2761;

 always  @(posedge PCLK)
	PKSi_87_<=N_N2762;

 always  @(posedge PCLK)
	PKSi_78_<=N_N2763;

 always  @(posedge PCLK)
	PKSi_95_<=N_N2764;

 always  @(posedge PCLK)
	PKSi_76_<=N_N2765;

 always  @(posedge PCLK)
	PKSi_55_<=N_N2766;

 always  @(posedge PCLK)
	PKSi_68_<=N_N2767;

 always  @(posedge PCLK)
	PKSi_64_<=N_N2768;

 always  @(posedge PCLK)
	N_N2770<=N_N2769;

 always  @(posedge PCLK)
	PKSi_51_<=N_N2771;

 always  @(posedge PCLK)
	PKSi_60_<=N_N2772;

 always  @(posedge PCLK)
	N_N2774<=N_N2773;

 always  @(posedge PCLK)
	PKSi_58_<=N_N2775;

 always  @(posedge PCLK)
	PKSi_69_<=N_N2776;

 always  @(posedge PCLK)
	PKSi_61_<=N_N2777;

 always  @(posedge PCLK)
	N_N2779<=N_N2778;

 always  @(posedge PCLK)
	PKSi_49_<=N_N2780;

 always  @(posedge PCLK)
	PKSi_66_<=N_N2781;

 always  @(posedge PCLK)
	PKSi_56_<=N_N2782;

 always  @(posedge PCLK)
	PKSi_48_<=N_N2783;

 always  @(posedge PCLK)
	PKSi_70_<=N_N2784;

 always  @(posedge PCLK)
	PKSi_62_<=N_N2785;

 always  @(posedge PCLK)
	PKSi_50_<=N_N2786;

 always  @(posedge PCLK)
	PKSi_59_<=N_N2787;

 always  @(posedge PCLK)
	N_N2789<=N_N2788;

 always  @(posedge PCLK)
	PKSi_65_<=N_N2790;

 always  @(posedge PCLK)
	PKSi_67_<=N_N2791;

 always  @(posedge PCLK)
	PKSi_57_<=N_N2792;

 always  @(posedge PCLK)
	PKSi_53_<=N_N2793;

 always  @(posedge PCLK)
	PKSi_63_<=N_N2794;

 always  @(posedge PCLK)
	PKSi_54_<=N_N2795;

 always  @(posedge PCLK)
	PKSi_71_<=N_N2796;

 always  @(posedge PCLK)
	PKSi_52_<=N_N2797;

 always  @(posedge PCLK)
	PKSi_31_<=N_N2798;

 always  @(posedge PCLK)
	PKSi_44_<=N_N2799;

 always  @(posedge PCLK)
	PKSi_40_<=N_N2800;

 always  @(posedge PCLK)
	N_N2802<=N_N2801;

 always  @(posedge PCLK)
	PKSi_27_<=N_N2803;

 always  @(posedge PCLK)
	PKSi_36_<=N_N2804;

 always  @(posedge PCLK)
	N_N2806<=N_N2805;

 always  @(posedge PCLK)
	PKSi_34_<=N_N2807;

 always  @(posedge PCLK)
	PKSi_45_<=N_N2808;

 always  @(posedge PCLK)
	PKSi_37_<=N_N2809;

 always  @(posedge PCLK)
	N_N2811<=N_N2810;

 always  @(posedge PCLK)
	PKSi_25_<=N_N2812;

 always  @(posedge PCLK)
	PKSi_42_<=N_N2813;

 always  @(posedge PCLK)
	PKSi_32_<=N_N2814;

 always  @(posedge PCLK)
	PKSi_24_<=N_N2815;

 always  @(posedge PCLK)
	PKSi_46_<=N_N2816;

 always  @(posedge PCLK)
	PKSi_38_<=N_N2817;

 always  @(posedge PCLK)
	PKSi_26_<=N_N2818;

 always  @(posedge PCLK)
	PKSi_35_<=N_N2819;

 always  @(posedge PCLK)
	N_N2821<=N_N2820;

 always  @(posedge PCLK)
	PKSi_41_<=N_N2822;

 always  @(posedge PCLK)
	PKSi_43_<=N_N2823;

 always  @(posedge PCLK)
	PKSi_33_<=N_N2824;

 always  @(posedge PCLK)
	PKSi_29_<=N_N2825;

 always  @(posedge PCLK)
	PKSi_39_<=N_N2826;

 always  @(posedge PCLK)
	PKSi_30_<=N_N2827;

 always  @(posedge PCLK)
	PKSi_47_<=N_N2828;

 always  @(posedge PCLK)
	PKSi_28_<=N_N2829;

 always  @(posedge PCLK)
	PKSi_7_<=N_N2830;

 always  @(posedge PCLK)
	PKSi_20_<=N_N2831;

 always  @(posedge PCLK)
	PKSi_16_<=N_N2832;

 always  @(posedge PCLK)
	N_N2834<=N_N2833;

 always  @(posedge PCLK)
	PKSi_3_<=N_N2835;

 always  @(posedge PCLK)
	PKSi_12_<=N_N2836;

 always  @(posedge PCLK)
	N_N2838<=N_N2837;

 always  @(posedge PCLK)
	PKSi_10_<=N_N2839;

 always  @(posedge PCLK)
	PKSi_21_<=N_N2840;

 always  @(posedge PCLK)
	PKSi_13_<=N_N2841;

 always  @(posedge PCLK)
	N_N2843<=N_N2842;

 always  @(posedge PCLK)
	PKSi_1_<=N_N2844;

 always  @(posedge PCLK)
	PKSi_18_<=N_N2845;

 always  @(posedge PCLK)
	PKSi_8_<=N_N2846;

 always  @(posedge PCLK)
	PKSi_0_<=N_N2847;

 always  @(posedge PCLK)
	PKSi_22_<=N_N2848;

 always  @(posedge PCLK)
	PKSi_14_<=N_N2849;

 always  @(posedge PCLK)
	PKSi_2_<=N_N2850;

 always  @(posedge PCLK)
	PKSi_11_<=N_N2851;

 always  @(posedge PCLK)
	N_N2853<=N_N2852;

 always  @(posedge PCLK)
	PKSi_17_<=N_N2854;

 always  @(posedge PCLK)
	PKSi_19_<=N_N2855;

 always  @(posedge PCLK)
	PKSi_9_<=N_N2856;

 always  @(posedge PCLK)
	PKSi_5_<=N_N2857;

 always  @(posedge PCLK)
	PKSi_15_<=N_N2858;

 always  @(posedge PCLK)
	PKSi_6_<=N_N2859;

 always  @(posedge PCLK)
	PKSi_23_<=N_N2860;

 always  @(posedge PCLK)
	PKSi_4_<=N_N2861;

 always  @(posedge PCLK)
	PKSi_183_<=N_N2862;

 always  @(posedge PCLK)
	PKSi_173_<=N_N2863;

 always  @(posedge PCLK)
	N_N2865<=N_N2864;

 always  @(posedge PCLK)
	PKSi_185_<=N_N2866;

 always  @(posedge PCLK)
	PKSi_169_<=N_N2867;

 always  @(posedge PCLK)
	PKSi_176_<=N_N2868;

 always  @(posedge PCLK)
	PKSi_188_<=N_N2869;

 always  @(posedge PCLK)
	wire253<=N_N2870;

 always  @(posedge PCLK)
	PKSi_179_<=N_N2871;

 always  @(posedge PCLK)
	PKSi_172_<=N_N2872;

 always  @(posedge PCLK)
	PKSi_186_<=N_N2873;

 always  @(posedge PCLK)
	PKSi_177_<=N_N2874;

 always  @(posedge PCLK)
	PKSi_180_<=N_N2875;

 always  @(posedge PCLK)
	N_N2877<=N_N2876;

 always  @(posedge PCLK)
	N_N2879<=N_N2878;

 always  @(posedge PCLK)
	N_N2881<=N_N2880;

 always  @(posedge PCLK)
	PKSi_175_<=N_N2882;

 always  @(posedge PCLK)
	PKSi_182_<=N_N2883;

 always  @(posedge PCLK)
	N_N2885<=N_N2884;

 always  @(posedge PCLK)
	PKSi_171_<=N_N2886;

 always  @(posedge PCLK)
	PKSi_189_<=N_N2887;

 always  @(posedge PCLK)
	N_N2889<=N_N2888;

 always  @(posedge PCLK)
	PKSi_184_<=N_N2890;

 always  @(posedge PCLK)
	PKSi_178_<=N_N2891;

 always  @(posedge PCLK)
	wire234<=N_N2892;

 always  @(posedge PCLK)
	PKSi_170_<=N_N2893;

 always  @(posedge PCLK)
	PKSi_174_<=N_N2894;

 always  @(posedge PCLK)
	PKSi_190_<=N_N2895;

 always  @(posedge PCLK)
	PKSi_159_<=N_N2896;

 always  @(posedge PCLK)
	PKSi_149_<=N_N2897;

 always  @(posedge PCLK)
	N_N2899<=N_N2898;

 always  @(posedge PCLK)
	PKSi_161_<=N_N2900;

 always  @(posedge PCLK)
	PKSi_145_<=N_N2901;

 always  @(posedge PCLK)
	PKSi_152_<=N_N2902;

 always  @(posedge PCLK)
	PKSi_164_<=N_N2903;

 always  @(posedge PCLK)
	PKSi_157_<=N_N2904;

 always  @(posedge PCLK)
	PKSi_155_<=N_N2905;

 always  @(posedge PCLK)
	PKSi_148_<=N_N2906;

 always  @(posedge PCLK)
	PKSi_162_<=N_N2907;

 always  @(posedge PCLK)
	N_N2909<=N_N2908;

 always  @(posedge PCLK)
	PKSi_156_<=N_N2910;

 always  @(posedge PCLK)
	PKSi_153_<=N_N2911;

 always  @(posedge PCLK)
	PKSi_163_<=N_N2912;

 always  @(posedge PCLK)
	PKSi_144_<=N_N2913;

 always  @(posedge PCLK)
	PKSi_151_<=N_N2914;

 always  @(posedge PCLK)
	PKSi_158_<=N_N2915;

 always  @(posedge PCLK)
	N_N2917<=N_N2916;

 always  @(posedge PCLK)
	PKSi_147_<=N_N2918;

 always  @(posedge PCLK)
	PKSi_165_<=N_N2919;

 always  @(posedge PCLK)
	N_N2921<=N_N2920;

 always  @(posedge PCLK)
	PKSi_160_<=N_N2922;

 always  @(posedge PCLK)
	PKSi_154_<=N_N2923;

 always  @(posedge PCLK)
	PKSi_167_<=N_N2924;

 always  @(posedge PCLK)
	PKSi_146_<=N_N2925;

 always  @(posedge PCLK)
	PKSi_150_<=N_N2926;

 always  @(posedge PCLK)
	PKSi_166_<=N_N2927;

 always  @(posedge PCLK)
	PKSi_135_<=N_N2928;

 always  @(posedge PCLK)
	PKSi_125_<=N_N2929;

 always  @(posedge PCLK)
	N_N2931<=N_N2930;

 always  @(posedge PCLK)
	PKSi_137_<=N_N2932;

 always  @(posedge PCLK)
	PKSi_121_<=N_N2933;

 always  @(posedge PCLK)
	PKSi_128_<=N_N2934;

 always  @(posedge PCLK)
	PKSi_140_<=N_N2935;

 always  @(posedge PCLK)
	PKSi_133_<=N_N2936;

 always  @(posedge PCLK)
	PKSi_131_<=N_N2937;

 always  @(posedge PCLK)
	PKSi_124_<=N_N2938;

 always  @(posedge PCLK)
	PKSi_138_<=N_N2939;

 always  @(posedge PCLK)
	PKSi_129_<=N_N2940;

 always  @(posedge PCLK)
	PKSi_132_<=N_N2941;

 always  @(posedge PCLK)
	N_N2943<=N_N2942;

 always  @(posedge PCLK)
	N_N2945<=N_N2944;

 always  @(posedge PCLK)
	PKSi_120_<=N_N2946;

 always  @(posedge PCLK)
	PKSi_127_<=N_N2947;

 always  @(posedge PCLK)
	PKSi_134_<=N_N2948;

 always  @(posedge PCLK)
	N_N2950<=N_N2949;

 always  @(posedge PCLK)
	PKSi_123_<=N_N2951;

 always  @(posedge PCLK)
	PKSi_141_<=N_N2952;

 always  @(posedge PCLK)
	N_N2954<=N_N2953;

 always  @(posedge PCLK)
	PKSi_136_<=N_N2955;

 always  @(posedge PCLK)
	PKSi_130_<=N_N2956;

 always  @(posedge PCLK)
	wire282<=N_N2957;

 always  @(posedge PCLK)
	PKSi_122_<=N_N2958;

 always  @(posedge PCLK)
	PKSi_126_<=N_N2959;

 always  @(posedge PCLK)
	PKSi_142_<=N_N2960;

 always  @(posedge PCLK)
	PKSi_111_<=N_N2961;

 always  @(posedge PCLK)
	PKSi_101_<=N_N2962;

 always  @(posedge PCLK)
	N_N2964<=N_N2963;

 always  @(posedge PCLK)
	PKSi_113_<=N_N2965;

 always  @(posedge PCLK)
	PKSi_97_<=N_N2966;

 always  @(posedge PCLK)
	PKSi_104_<=N_N2967;

 always  @(posedge PCLK)
	PKSi_116_<=N_N2968;

 always  @(posedge PCLK)
	PKSi_109_<=N_N2969;

 always  @(posedge PCLK)
	PKSi_107_<=N_N2970;

 always  @(posedge PCLK)
	PKSi_100_<=N_N2971;

 always  @(posedge PCLK)
	PKSi_114_<=N_N2972;

 always  @(posedge PCLK)
	PKSi_105_<=N_N2973;

 always  @(posedge PCLK)
	PKSi_108_<=N_N2974;

 always  @(posedge PCLK)
	N_N2976<=N_N2975;

 always  @(posedge PCLK)
	PKSi_115_<=N_N2977;

 always  @(posedge PCLK)
	PKSi_96_<=N_N2978;

 always  @(posedge PCLK)
	PKSi_103_<=N_N2979;

 always  @(posedge PCLK)
	PKSi_110_<=N_N2980;

 always  @(posedge PCLK)
	N_N2982<=N_N2981;

 always  @(posedge PCLK)
	PKSi_99_<=N_N2983;

 always  @(posedge PCLK)
	PKSi_117_<=N_N2984;

 always  @(posedge PCLK)
	N_N2986<=N_N2985;

 always  @(posedge PCLK)
	PKSi_112_<=N_N2987;

 always  @(posedge PCLK)
	PKSi_106_<=N_N2988;

 always  @(posedge PCLK)
	PKSi_119_<=N_N2989;

 always  @(posedge PCLK)
	PKSi_98_<=N_N2990;

 always  @(posedge PCLK)
	PKSi_102_<=N_N2991;

 always  @(posedge PCLK)
	PKSi_118_<=N_N2992;

 assign Pnew_count_3_ = ( (~ n17) ) ;
 assign Pnew_count_2_ = ( (~ n18) ) ;
 assign Pnew_count_1_ = ( (~ n19) ) ;
 assign Pnew_count_0_ = ( (~ n20) ) ;
 assign Pdata_ready_0_ = ( (~ n16) ) ;
 assign n15 = ( (~ Pstart_0_) ) | ( Pencrypt_0_ ) ;
 assign n13 = ( (~ Pstart_0_) ) | ( (~ Pencrypt_0_) ) ;
 assign n11 = ( Pstart_0_ ) | ( Pencrypt_0_ ) | ( n245 ) ;
 assign n1741 = ( (~ Pstart_0_)  &  (~ Pencrypt_0_)  &  n245 ) ;
 assign n16 = ( n925  &  Pstart_0_ ) | ( n925  &  n924 ) ;
 assign n17 = ( Pstart_0_  &  n15 ) | ( n15  &  n937 ) ;
 assign n18 = ( Pencrypt_0_  &  (~ n930)  &  n934 ) | ( n249  &  (~ n930)  &  n934 ) ;
 assign n19 = ( (~ Pcount_0_)  &  n15  &  n929 ) | ( n15  &  n929  &  n928 ) ;
 assign n20 = ( Pstart_0_  &  n15 ) | ( Pcount_0_  &  n15 ) ;
 assign n21 = ( (~ Pkey_62_)  &  n586  &  n587 ) | ( n13  &  n586  &  n587 ) ;
 assign N_N2862 = ( (~ n21) ) ;
 assign n22 = ( (~ Pkey_195_)  &  n583  &  n584 ) | ( n13  &  n583  &  n584 ) ;
 assign N_N2863 = ( (~ n22) ) ;
 assign n23 = ( (~ Pkey_203_)  &  n580  &  n581 ) | ( n13  &  n580  &  n581 ) ;
 assign N_N2864 = ( (~ n23) ) ;
 assign n24 = ( (~ Pkey_211_)  &  n577  &  n578 ) | ( n13  &  n577  &  n578 ) ;
 assign N_N2866 = ( (~ n24) ) ;
 assign n25 = ( (~ Pkey_219_)  &  n574  &  n575 ) | ( n13  &  n574  &  n575 ) ;
 assign N_N2867 = ( (~ n25) ) ;
 assign n26 = ( (~ Pkey_196_)  &  n571  &  n572 ) | ( n13  &  n571  &  n572 ) ;
 assign N_N2868 = ( (~ n26) ) ;
 assign n27 = ( (~ Pkey_204_)  &  n568  &  n569 ) | ( n13  &  n568  &  n569 ) ;
 assign N_N2869 = ( (~ n27) ) ;
 assign n28 = ( (~ Pkey_212_)  &  n565  &  n566 ) | ( n13  &  n565  &  n566 ) ;
 assign N_N2870 = ( (~ n28) ) ;
 assign n29 = ( (~ Pkey_220_)  &  n562  &  n563 ) | ( n13  &  n562  &  n563 ) ;
 assign N_N2871 = ( (~ n29) ) ;
 assign n30 = ( (~ Pkey_228_)  &  n559  &  n560 ) | ( n13  &  n559  &  n560 ) ;
 assign N_N2872 = ( (~ n30) ) ;
 assign n31 = ( (~ Pkey_172_)  &  n556  &  n557 ) | ( n13  &  n556  &  n557 ) ;
 assign N_N2873 = ( (~ n31) ) ;
 assign n32 = ( (~ Pkey_244_)  &  n554  &  n555 ) | ( n13  &  n554  &  n555 ) ;
 assign N_N2874 = ( (~ n32) ) ;
 assign n33 = ( (~ Pkey_252_)  &  n551  &  n552 ) | ( n13  &  n551  &  n552 ) ;
 assign N_N2875 = ( (~ n33) ) ;
 assign n34 = ( (~ Pkey_197_)  &  n548  &  n549 ) | ( n13  &  n548  &  n549 ) ;
 assign N_N2876 = ( (~ n34) ) ;
 assign n35 = ( (~ Pkey_205_)  &  n545  &  n546 ) | ( n13  &  n545  &  n546 ) ;
 assign N_N2878 = ( (~ n35) ) ;
 assign n36 = ( (~ Pkey_213_)  &  n542  &  n543 ) | ( n13  &  n542  &  n543 ) ;
 assign N_N2880 = ( (~ n36) ) ;
 assign n37 = ( (~ Pkey_221_)  &  n539  &  n540 ) | ( n13  &  n539  &  n540 ) ;
 assign N_N2882 = ( (~ n37) ) ;
 assign n38 = ( (~ Pkey_229_)  &  n536  &  n537 ) | ( n13  &  n536  &  n537 ) ;
 assign N_N2883 = ( (~ n38) ) ;
 assign n39 = ( (~ Pkey_237_)  &  n533  &  n534 ) | ( n13  &  n533  &  n534 ) ;
 assign N_N2884 = ( (~ n39) ) ;
 assign n40 = ( (~ Pkey_245_)  &  n530  &  n531 ) | ( n13  &  n530  &  n531 ) ;
 assign N_N2886 = ( (~ n40) ) ;
 assign n41 = ( (~ Pkey_253_)  &  n527  &  n528 ) | ( n13  &  n527  &  n528 ) ;
 assign N_N2887 = ( (~ n41) ) ;
 assign n42 = ( (~ Pkey_198_)  &  n524  &  n525 ) | ( n13  &  n524  &  n525 ) ;
 assign N_N2888 = ( (~ n42) ) ;
 assign n43 = ( (~ Pkey_206_)  &  n521  &  n522 ) | ( n13  &  n521  &  n522 ) ;
 assign N_N2890 = ( (~ n43) ) ;
 assign n44 = ( (~ Pkey_214_)  &  n518  &  n519 ) | ( n13  &  n518  &  n519 ) ;
 assign N_N2891 = ( (~ n44) ) ;
 assign n45 = ( (~ Pkey_222_)  &  n515  &  n516 ) | ( n13  &  n515  &  n516 ) ;
 assign N_N2892 = ( (~ n45) ) ;
 assign n46 = ( (~ Pkey_230_)  &  n512  &  n513 ) | ( n13  &  n512  &  n513 ) ;
 assign N_N2893 = ( (~ n46) ) ;
 assign n47 = ( (~ Pkey_238_)  &  n509  &  n510 ) | ( n13  &  n509  &  n510 ) ;
 assign N_N2894 = ( (~ n47) ) ;
 assign n48 = ( (~ Pkey_246_)  &  n506  &  n507 ) | ( n13  &  n506  &  n507 ) ;
 assign N_N2895 = ( (~ n48) ) ;
 assign n49 = ( (~ Pkey_254_)  &  n503  &  n504 ) | ( n13  &  n503  &  n504 ) ;
 assign N_N2896 = ( (~ n49) ) ;
 assign n50 = ( (~ Pkey_131_)  &  n500  &  n501 ) | ( n13  &  n500  &  n501 ) ;
 assign N_N2897 = ( (~ n50) ) ;
 assign n51 = ( (~ Pkey_139_)  &  n497  &  n498 ) | ( n13  &  n497  &  n498 ) ;
 assign N_N2898 = ( (~ n51) ) ;
 assign n52 = ( (~ Pkey_147_)  &  n494  &  n495 ) | ( n13  &  n494  &  n495 ) ;
 assign N_N2900 = ( (~ n52) ) ;
 assign n53 = ( (~ Pkey_155_)  &  n491  &  n492 ) | ( n13  &  n491  &  n492 ) ;
 assign N_N2901 = ( (~ n53) ) ;
 assign n54 = ( (~ Pkey_132_)  &  n488  &  n489 ) | ( n13  &  n488  &  n489 ) ;
 assign N_N2902 = ( (~ n54) ) ;
 assign n55 = ( (~ Pkey_140_)  &  n485  &  n486 ) | ( n13  &  n485  &  n486 ) ;
 assign N_N2903 = ( (~ n55) ) ;
 assign n56 = ( (~ Pkey_148_)  &  n482  &  n483 ) | ( n13  &  n482  &  n483 ) ;
 assign N_N2904 = ( (~ n56) ) ;
 assign n57 = ( (~ Pkey_156_)  &  n479  &  n480 ) | ( n13  &  n479  &  n480 ) ;
 assign N_N2905 = ( (~ n57) ) ;
 assign n58 = ( (~ Pkey_164_)  &  n476  &  n477 ) | ( n13  &  n476  &  n477 ) ;
 assign N_N2906 = ( (~ n58) ) ;
 assign n59 = ( (~ Pkey_172_)  &  n473  &  n474 ) | ( n13  &  n473  &  n474 ) ;
 assign N_N2907 = ( (~ n59) ) ;
 assign n60 = ( (~ Pkey_180_)  &  n470  &  n471 ) | ( n13  &  n470  &  n471 ) ;
 assign N_N2908 = ( (~ n60) ) ;
 assign n61 = ( (~ Pkey_188_)  &  n467  &  n468 ) | ( n13  &  n467  &  n468 ) ;
 assign N_N2910 = ( (~ n61) ) ;
 assign n62 = ( (~ Pkey_133_)  &  n464  &  n465 ) | ( n13  &  n464  &  n465 ) ;
 assign N_N2911 = ( (~ n62) ) ;
 assign n63 = ( (~ Pkey_141_)  &  n461  &  n462 ) | ( n13  &  n461  &  n462 ) ;
 assign N_N2912 = ( (~ n63) ) ;
 assign n64 = ( (~ Pkey_149_)  &  n458  &  n459 ) | ( n13  &  n458  &  n459 ) ;
 assign N_N2913 = ( (~ n64) ) ;
 assign n65 = ( (~ Pkey_157_)  &  n455  &  n456 ) | ( n13  &  n455  &  n456 ) ;
 assign N_N2914 = ( (~ n65) ) ;
 assign n66 = ( (~ Pkey_165_)  &  n452  &  n453 ) | ( n13  &  n452  &  n453 ) ;
 assign N_N2915 = ( (~ n66) ) ;
 assign n67 = ( (~ Pkey_173_)  &  n449  &  n450 ) | ( n13  &  n449  &  n450 ) ;
 assign N_N2916 = ( (~ n67) ) ;
 assign n68 = ( (~ Pkey_181_)  &  n446  &  n447 ) | ( n13  &  n446  &  n447 ) ;
 assign N_N2918 = ( (~ n68) ) ;
 assign n69 = ( (~ Pkey_189_)  &  n443  &  n444 ) | ( n13  &  n443  &  n444 ) ;
 assign N_N2919 = ( (~ n69) ) ;
 assign n70 = ( (~ Pkey_134_)  &  n440  &  n441 ) | ( n13  &  n440  &  n441 ) ;
 assign N_N2920 = ( (~ n70) ) ;
 assign n71 = ( (~ Pkey_142_)  &  n437  &  n438 ) | ( n13  &  n437  &  n438 ) ;
 assign N_N2922 = ( (~ n71) ) ;
 assign n72 = ( (~ Pkey_150_)  &  n434  &  n435 ) | ( n13  &  n434  &  n435 ) ;
 assign N_N2923 = ( (~ n72) ) ;
 assign n73 = ( (~ Pkey_158_)  &  n431  &  n432 ) | ( n13  &  n431  &  n432 ) ;
 assign N_N2924 = ( (~ n73) ) ;
 assign n74 = ( (~ Pkey_166_)  &  n428  &  n429 ) | ( n13  &  n428  &  n429 ) ;
 assign N_N2925 = ( (~ n74) ) ;
 assign n75 = ( (~ Pkey_174_)  &  n425  &  n426 ) | ( n13  &  n425  &  n426 ) ;
 assign N_N2926 = ( (~ n75) ) ;
 assign n76 = ( (~ Pkey_182_)  &  n422  &  n423 ) | ( n13  &  n422  &  n423 ) ;
 assign N_N2927 = ( (~ n76) ) ;
 assign n77 = ( (~ Pkey_190_)  &  n419  &  n420 ) | ( n13  &  n419  &  n420 ) ;
 assign N_N2928 = ( (~ n77) ) ;
 assign n78 = ( (~ Pkey_67_)  &  n416  &  n417 ) | ( n13  &  n416  &  n417 ) ;
 assign N_N2929 = ( (~ n78) ) ;
 assign n79 = ( (~ Pkey_75_)  &  n413  &  n414 ) | ( n13  &  n413  &  n414 ) ;
 assign N_N2930 = ( (~ n79) ) ;
 assign n80 = ( (~ Pkey_83_)  &  n410  &  n411 ) | ( n13  &  n410  &  n411 ) ;
 assign N_N2932 = ( (~ n80) ) ;
 assign n81 = ( (~ Pkey_91_)  &  n407  &  n408 ) | ( n13  &  n407  &  n408 ) ;
 assign N_N2933 = ( (~ n81) ) ;
 assign n82 = ( (~ Pkey_68_)  &  n404  &  n405 ) | ( n13  &  n404  &  n405 ) ;
 assign N_N2934 = ( (~ n82) ) ;
 assign n83 = ( (~ Pkey_76_)  &  n401  &  n402 ) | ( n13  &  n401  &  n402 ) ;
 assign N_N2935 = ( (~ n83) ) ;
 assign n84 = ( (~ Pkey_84_)  &  n398  &  n399 ) | ( n13  &  n398  &  n399 ) ;
 assign N_N2936 = ( (~ n84) ) ;
 assign n85 = ( (~ Pkey_92_)  &  n395  &  n396 ) | ( n13  &  n395  &  n396 ) ;
 assign N_N2937 = ( (~ n85) ) ;
 assign n86 = ( (~ Pkey_100_)  &  n392  &  n393 ) | ( n13  &  n392  &  n393 ) ;
 assign N_N2938 = ( (~ n86) ) ;
 assign n87 = ( (~ Pkey_44_)  &  n389  &  n390 ) | ( n13  &  n389  &  n390 ) ;
 assign N_N2939 = ( (~ n87) ) ;
 assign n88 = ( (~ Pkey_116_)  &  n387  &  n388 ) | ( n13  &  n387  &  n388 ) ;
 assign N_N2940 = ( (~ n88) ) ;
 assign n89 = ( (~ Pkey_124_)  &  n384  &  n385 ) | ( n13  &  n384  &  n385 ) ;
 assign N_N2941 = ( (~ n89) ) ;
 assign n90 = ( (~ Pkey_69_)  &  n381  &  n382 ) | ( n13  &  n381  &  n382 ) ;
 assign N_N2942 = ( (~ n90) ) ;
 assign n91 = ( (~ Pkey_77_)  &  n378  &  n379 ) | ( n13  &  n378  &  n379 ) ;
 assign N_N2944 = ( (~ n91) ) ;
 assign n92 = ( (~ Pkey_85_)  &  n375  &  n376 ) | ( n13  &  n375  &  n376 ) ;
 assign N_N2946 = ( (~ n92) ) ;
 assign n93 = ( (~ Pkey_93_)  &  n372  &  n373 ) | ( n13  &  n372  &  n373 ) ;
 assign N_N2947 = ( (~ n93) ) ;
 assign n94 = ( (~ Pkey_101_)  &  n369  &  n370 ) | ( n13  &  n369  &  n370 ) ;
 assign N_N2948 = ( (~ n94) ) ;
 assign n95 = ( (~ Pkey_109_)  &  n366  &  n367 ) | ( n13  &  n366  &  n367 ) ;
 assign N_N2949 = ( (~ n95) ) ;
 assign n96 = ( (~ Pkey_117_)  &  n363  &  n364 ) | ( n13  &  n363  &  n364 ) ;
 assign N_N2951 = ( (~ n96) ) ;
 assign n97 = ( (~ Pkey_125_)  &  n360  &  n361 ) | ( n13  &  n360  &  n361 ) ;
 assign N_N2952 = ( (~ n97) ) ;
 assign n98 = ( (~ Pkey_70_)  &  n357  &  n358 ) | ( n13  &  n357  &  n358 ) ;
 assign N_N2953 = ( (~ n98) ) ;
 assign n99 = ( (~ Pkey_78_)  &  n354  &  n355 ) | ( n13  &  n354  &  n355 ) ;
 assign N_N2955 = ( (~ n99) ) ;
 assign n100 = ( (~ Pkey_86_)  &  n351  &  n352 ) | ( n13  &  n351  &  n352 ) ;
 assign N_N2956 = ( (~ n100) ) ;
 assign n101 = ( (~ Pkey_94_)  &  n348  &  n349 ) | ( n13  &  n348  &  n349 ) ;
 assign N_N2957 = ( (~ n101) ) ;
 assign n102 = ( (~ Pkey_102_)  &  n345  &  n346 ) | ( n13  &  n345  &  n346 ) ;
 assign N_N2958 = ( (~ n102) ) ;
 assign n103 = ( (~ Pkey_110_)  &  n342  &  n343 ) | ( n13  &  n342  &  n343 ) ;
 assign N_N2959 = ( (~ n103) ) ;
 assign n104 = ( (~ Pkey_118_)  &  n339  &  n340 ) | ( n13  &  n339  &  n340 ) ;
 assign N_N2960 = ( (~ n104) ) ;
 assign n105 = ( (~ Pkey_126_)  &  n336  &  n337 ) | ( n13  &  n336  &  n337 ) ;
 assign N_N2961 = ( (~ n105) ) ;
 assign n106 = ( (~ Pkey_3_)  &  n333  &  n334 ) | ( n13  &  n333  &  n334 ) ;
 assign N_N2962 = ( (~ n106) ) ;
 assign n107 = ( (~ Pkey_11_)  &  n330  &  n331 ) | ( n13  &  n330  &  n331 ) ;
 assign N_N2963 = ( (~ n107) ) ;
 assign n108 = ( (~ Pkey_19_)  &  n327  &  n328 ) | ( n13  &  n327  &  n328 ) ;
 assign N_N2965 = ( (~ n108) ) ;
 assign n109 = ( (~ Pkey_27_)  &  n324  &  n325 ) | ( n13  &  n324  &  n325 ) ;
 assign N_N2966 = ( (~ n109) ) ;
 assign n110 = ( (~ Pkey_4_)  &  n321  &  n322 ) | ( n13  &  n321  &  n322 ) ;
 assign N_N2967 = ( (~ n110) ) ;
 assign n111 = ( (~ Pkey_12_)  &  n318  &  n319 ) | ( n13  &  n318  &  n319 ) ;
 assign N_N2968 = ( (~ n111) ) ;
 assign n112 = ( (~ Pkey_20_)  &  n315  &  n316 ) | ( n13  &  n315  &  n316 ) ;
 assign N_N2969 = ( (~ n112) ) ;
 assign n113 = ( (~ Pkey_28_)  &  n312  &  n313 ) | ( n13  &  n312  &  n313 ) ;
 assign N_N2970 = ( (~ n113) ) ;
 assign n114 = ( (~ Pkey_36_)  &  n309  &  n310 ) | ( n13  &  n309  &  n310 ) ;
 assign N_N2971 = ( (~ n114) ) ;
 assign n115 = ( (~ Pkey_44_)  &  n306  &  n307 ) | ( n13  &  n306  &  n307 ) ;
 assign N_N2972 = ( (~ n115) ) ;
 assign n116 = ( (~ Pkey_52_)  &  n303  &  n304 ) | ( n13  &  n303  &  n304 ) ;
 assign N_N2973 = ( (~ n116) ) ;
 assign n117 = ( (~ Pkey_60_)  &  n300  &  n301 ) | ( n13  &  n300  &  n301 ) ;
 assign N_N2974 = ( (~ n117) ) ;
 assign n118 = ( (~ Pkey_5_)  &  n297  &  n298 ) | ( n13  &  n297  &  n298 ) ;
 assign N_N2975 = ( (~ n118) ) ;
 assign n119 = ( (~ Pkey_13_)  &  n294  &  n295 ) | ( n13  &  n294  &  n295 ) ;
 assign N_N2977 = ( (~ n119) ) ;
 assign n120 = ( (~ Pkey_21_)  &  n291  &  n292 ) | ( n13  &  n291  &  n292 ) ;
 assign N_N2978 = ( (~ n120) ) ;
 assign n121 = ( (~ Pkey_29_)  &  n288  &  n289 ) | ( n13  &  n288  &  n289 ) ;
 assign N_N2979 = ( (~ n121) ) ;
 assign n122 = ( (~ Pkey_37_)  &  n285  &  n286 ) | ( n13  &  n285  &  n286 ) ;
 assign N_N2980 = ( (~ n122) ) ;
 assign n123 = ( (~ Pkey_45_)  &  n282  &  n283 ) | ( n13  &  n282  &  n283 ) ;
 assign N_N2981 = ( (~ n123) ) ;
 assign n124 = ( (~ Pkey_53_)  &  n279  &  n280 ) | ( n13  &  n279  &  n280 ) ;
 assign N_N2983 = ( (~ n124) ) ;
 assign n125 = ( (~ Pkey_61_)  &  n276  &  n277 ) | ( n13  &  n276  &  n277 ) ;
 assign N_N2984 = ( (~ n125) ) ;
 assign n126 = ( (~ Pkey_6_)  &  n273  &  n274 ) | ( n13  &  n273  &  n274 ) ;
 assign N_N2985 = ( (~ n126) ) ;
 assign n127 = ( (~ Pkey_14_)  &  n270  &  n271 ) | ( n13  &  n270  &  n271 ) ;
 assign N_N2987 = ( (~ n127) ) ;
 assign n128 = ( (~ Pkey_22_)  &  n267  &  n268 ) | ( n13  &  n267  &  n268 ) ;
 assign N_N2988 = ( (~ n128) ) ;
 assign n129 = ( (~ Pkey_30_)  &  n264  &  n265 ) | ( n13  &  n264  &  n265 ) ;
 assign N_N2989 = ( (~ n129) ) ;
 assign n130 = ( (~ Pkey_38_)  &  n261  &  n262 ) | ( n13  &  n261  &  n262 ) ;
 assign N_N2990 = ( (~ n130) ) ;
 assign n131 = ( (~ Pkey_46_)  &  n258  &  n259 ) | ( n13  &  n258  &  n259 ) ;
 assign N_N2991 = ( (~ n131) ) ;
 assign n132 = ( (~ Pkey_54_)  &  n255  &  n256 ) | ( n13  &  n255  &  n256 ) ;
 assign N_N2992 = ( (~ n132) ) ;
 assign n133 = ( (~ Pkey_56_)  &  n922  &  n923 ) | ( n13  &  n922  &  n923 ) ;
 assign N_N2733 = ( (~ n133) ) ;
 assign n134 = ( (~ Pkey_227_)  &  n919  &  n920 ) | ( n13  &  n919  &  n920 ) ;
 assign N_N2734 = ( (~ n134) ) ;
 assign n135 = ( (~ Pkey_235_)  &  n916  &  n917 ) | ( n13  &  n916  &  n917 ) ;
 assign N_N2735 = ( (~ n135) ) ;
 assign n136 = ( (~ Pkey_243_)  &  n913  &  n914 ) | ( n13  &  n913  &  n914 ) ;
 assign N_N2736 = ( (~ n136) ) ;
 assign n137 = ( (~ Pkey_251_)  &  n910  &  n911 ) | ( n13  &  n910  &  n911 ) ;
 assign N_N2738 = ( (~ n137) ) ;
 assign n138 = ( (~ Pkey_194_)  &  n907  &  n908 ) | ( n13  &  n907  &  n908 ) ;
 assign N_N2739 = ( (~ n138) ) ;
 assign n139 = ( (~ Pkey_202_)  &  n904  &  n905 ) | ( n13  &  n904  &  n905 ) ;
 assign N_N2740 = ( (~ n139) ) ;
 assign n140 = ( (~ Pkey_210_)  &  n901  &  n902 ) | ( n13  &  n901  &  n902 ) ;
 assign N_N2742 = ( (~ n140) ) ;
 assign n141 = ( (~ Pkey_218_)  &  n898  &  n899 ) | ( n13  &  n898  &  n899 ) ;
 assign N_N2743 = ( (~ n141) ) ;
 assign n142 = ( (~ Pkey_226_)  &  n895  &  n896 ) | ( n13  &  n895  &  n896 ) ;
 assign N_N2744 = ( (~ n142) ) ;
 assign n143 = ( (~ Pkey_234_)  &  n892  &  n893 ) | ( n13  &  n892  &  n893 ) ;
 assign N_N2745 = ( (~ n143) ) ;
 assign n144 = ( (~ Pkey_242_)  &  n889  &  n890 ) | ( n13  &  n889  &  n890 ) ;
 assign N_N2747 = ( (~ n144) ) ;
 assign n145 = ( (~ Pkey_250_)  &  n886  &  n887 ) | ( n13  &  n886  &  n887 ) ;
 assign N_N2748 = ( (~ n145) ) ;
 assign n146 = ( (~ Pkey_193_)  &  n883  &  n884 ) | ( n13  &  n883  &  n884 ) ;
 assign N_N2750 = ( (~ n146) ) ;
 assign n147 = ( (~ Pkey_201_)  &  n880  &  n881 ) | ( n13  &  n880  &  n881 ) ;
 assign N_N2751 = ( (~ n147) ) ;
 assign n148 = ( (~ Pkey_209_)  &  n877  &  n878 ) | ( n13  &  n877  &  n878 ) ;
 assign N_N2752 = ( (~ n148) ) ;
 assign n149 = ( (~ Pkey_217_)  &  n874  &  n875 ) | ( n13  &  n874  &  n875 ) ;
 assign N_N2753 = ( (~ n149) ) ;
 assign n150 = ( (~ Pkey_225_)  &  n871  &  n872 ) | ( n13  &  n871  &  n872 ) ;
 assign N_N2754 = ( (~ n150) ) ;
 assign n151 = ( (~ Pkey_233_)  &  n868  &  n869 ) | ( n13  &  n868  &  n869 ) ;
 assign N_N2755 = ( (~ n151) ) ;
 assign n152 = ( (~ Pkey_241_)  &  n865  &  n866 ) | ( n13  &  n865  &  n866 ) ;
 assign N_N2756 = ( (~ n152) ) ;
 assign n153 = ( (~ Pkey_249_)  &  n862  &  n863 ) | ( n13  &  n862  &  n863 ) ;
 assign N_N2758 = ( (~ n153) ) ;
 assign n154 = ( (~ Pkey_192_)  &  n859  &  n860 ) | ( n13  &  n859  &  n860 ) ;
 assign N_N2759 = ( (~ n154) ) ;
 assign n155 = ( (~ Pkey_200_)  &  n856  &  n857 ) | ( n13  &  n856  &  n857 ) ;
 assign N_N2760 = ( (~ n155) ) ;
 assign n156 = ( (~ Pkey_208_)  &  n853  &  n854 ) | ( n13  &  n853  &  n854 ) ;
 assign N_N2761 = ( (~ n156) ) ;
 assign n157 = ( (~ Pkey_216_)  &  n850  &  n851 ) | ( n13  &  n850  &  n851 ) ;
 assign N_N2762 = ( (~ n157) ) ;
 assign n158 = ( (~ Pkey_224_)  &  n847  &  n848 ) | ( n13  &  n847  &  n848 ) ;
 assign N_N2763 = ( (~ n158) ) ;
 assign n159 = ( (~ Pkey_232_)  &  n844  &  n845 ) | ( n13  &  n844  &  n845 ) ;
 assign N_N2764 = ( (~ n159) ) ;
 assign n160 = ( (~ Pkey_240_)  &  n841  &  n842 ) | ( n13  &  n841  &  n842 ) ;
 assign N_N2765 = ( (~ n160) ) ;
 assign n161 = ( (~ Pkey_248_)  &  n838  &  n839 ) | ( n13  &  n838  &  n839 ) ;
 assign N_N2766 = ( (~ n161) ) ;
 assign n162 = ( (~ Pkey_163_)  &  n835  &  n836 ) | ( n13  &  n835  &  n836 ) ;
 assign N_N2767 = ( (~ n162) ) ;
 assign n163 = ( (~ Pkey_171_)  &  n832  &  n833 ) | ( n13  &  n832  &  n833 ) ;
 assign N_N2768 = ( (~ n163) ) ;
 assign n164 = ( (~ Pkey_179_)  &  n829  &  n830 ) | ( n13  &  n829  &  n830 ) ;
 assign N_N2769 = ( (~ n164) ) ;
 assign n165 = ( (~ Pkey_187_)  &  n826  &  n827 ) | ( n13  &  n826  &  n827 ) ;
 assign N_N2771 = ( (~ n165) ) ;
 assign n166 = ( (~ Pkey_130_)  &  n823  &  n824 ) | ( n13  &  n823  &  n824 ) ;
 assign N_N2772 = ( (~ n166) ) ;
 assign n167 = ( (~ Pkey_138_)  &  n820  &  n821 ) | ( n13  &  n820  &  n821 ) ;
 assign N_N2773 = ( (~ n167) ) ;
 assign n168 = ( (~ Pkey_146_)  &  n817  &  n818 ) | ( n13  &  n817  &  n818 ) ;
 assign N_N2775 = ( (~ n168) ) ;
 assign n169 = ( (~ Pkey_154_)  &  n814  &  n815 ) | ( n13  &  n814  &  n815 ) ;
 assign N_N2776 = ( (~ n169) ) ;
 assign n170 = ( (~ Pkey_162_)  &  n811  &  n812 ) | ( n13  &  n811  &  n812 ) ;
 assign N_N2777 = ( (~ n170) ) ;
 assign n171 = ( (~ Pkey_170_)  &  n808  &  n809 ) | ( n13  &  n808  &  n809 ) ;
 assign N_N2778 = ( (~ n171) ) ;
 assign n172 = ( (~ Pkey_178_)  &  n805  &  n806 ) | ( n13  &  n805  &  n806 ) ;
 assign N_N2780 = ( (~ n172) ) ;
 assign n173 = ( (~ Pkey_186_)  &  n802  &  n803 ) | ( n13  &  n802  &  n803 ) ;
 assign N_N2781 = ( (~ n173) ) ;
 assign n174 = ( (~ Pkey_129_)  &  n799  &  n800 ) | ( n13  &  n799  &  n800 ) ;
 assign N_N2782 = ( (~ n174) ) ;
 assign n175 = ( (~ Pkey_137_)  &  n796  &  n797 ) | ( n13  &  n796  &  n797 ) ;
 assign N_N2783 = ( (~ n175) ) ;
 assign n176 = ( (~ Pkey_145_)  &  n793  &  n794 ) | ( n13  &  n793  &  n794 ) ;
 assign N_N2784 = ( (~ n176) ) ;
 assign n177 = ( (~ Pkey_153_)  &  n790  &  n791 ) | ( n13  &  n790  &  n791 ) ;
 assign N_N2785 = ( (~ n177) ) ;
 assign n178 = ( (~ Pkey_161_)  &  n787  &  n788 ) | ( n13  &  n787  &  n788 ) ;
 assign N_N2786 = ( (~ n178) ) ;
 assign n179 = ( (~ Pkey_169_)  &  n784  &  n785 ) | ( n13  &  n784  &  n785 ) ;
 assign N_N2787 = ( (~ n179) ) ;
 assign n180 = ( (~ Pkey_177_)  &  n781  &  n782 ) | ( n13  &  n781  &  n782 ) ;
 assign N_N2788 = ( (~ n180) ) ;
 assign n181 = ( (~ Pkey_185_)  &  n778  &  n779 ) | ( n13  &  n778  &  n779 ) ;
 assign N_N2790 = ( (~ n181) ) ;
 assign n182 = ( (~ Pkey_128_)  &  n775  &  n776 ) | ( n13  &  n775  &  n776 ) ;
 assign N_N2791 = ( (~ n182) ) ;
 assign n183 = ( (~ Pkey_136_)  &  n772  &  n773 ) | ( n13  &  n772  &  n773 ) ;
 assign N_N2792 = ( (~ n183) ) ;
 assign n184 = ( (~ Pkey_144_)  &  n769  &  n770 ) | ( n13  &  n769  &  n770 ) ;
 assign N_N2793 = ( (~ n184) ) ;
 assign n185 = ( (~ Pkey_152_)  &  n766  &  n767 ) | ( n13  &  n766  &  n767 ) ;
 assign N_N2794 = ( (~ n185) ) ;
 assign n186 = ( (~ Pkey_160_)  &  n763  &  n764 ) | ( n13  &  n763  &  n764 ) ;
 assign N_N2795 = ( (~ n186) ) ;
 assign n187 = ( (~ Pkey_168_)  &  n760  &  n761 ) | ( n13  &  n760  &  n761 ) ;
 assign N_N2796 = ( (~ n187) ) ;
 assign n188 = ( (~ Pkey_176_)  &  n757  &  n758 ) | ( n13  &  n757  &  n758 ) ;
 assign N_N2797 = ( (~ n188) ) ;
 assign n189 = ( (~ Pkey_184_)  &  n754  &  n755 ) | ( n13  &  n754  &  n755 ) ;
 assign N_N2798 = ( (~ n189) ) ;
 assign n190 = ( (~ Pkey_99_)  &  n751  &  n752 ) | ( n13  &  n751  &  n752 ) ;
 assign N_N2799 = ( (~ n190) ) ;
 assign n191 = ( (~ Pkey_107_)  &  n748  &  n749 ) | ( n13  &  n748  &  n749 ) ;
 assign N_N2800 = ( (~ n191) ) ;
 assign n192 = ( (~ Pkey_115_)  &  n745  &  n746 ) | ( n13  &  n745  &  n746 ) ;
 assign N_N2801 = ( (~ n192) ) ;
 assign n193 = ( (~ Pkey_123_)  &  n742  &  n743 ) | ( n13  &  n742  &  n743 ) ;
 assign N_N2803 = ( (~ n193) ) ;
 assign n194 = ( (~ Pkey_66_)  &  n739  &  n740 ) | ( n13  &  n739  &  n740 ) ;
 assign N_N2804 = ( (~ n194) ) ;
 assign n195 = ( (~ Pkey_74_)  &  n736  &  n737 ) | ( n13  &  n736  &  n737 ) ;
 assign N_N2805 = ( (~ n195) ) ;
 assign n196 = ( (~ Pkey_82_)  &  n733  &  n734 ) | ( n13  &  n733  &  n734 ) ;
 assign N_N2807 = ( (~ n196) ) ;
 assign n197 = ( (~ Pkey_90_)  &  n730  &  n731 ) | ( n13  &  n730  &  n731 ) ;
 assign N_N2808 = ( (~ n197) ) ;
 assign n198 = ( (~ Pkey_98_)  &  n727  &  n728 ) | ( n13  &  n727  &  n728 ) ;
 assign N_N2809 = ( (~ n198) ) ;
 assign n199 = ( (~ Pkey_106_)  &  n724  &  n725 ) | ( n13  &  n724  &  n725 ) ;
 assign N_N2810 = ( (~ n199) ) ;
 assign n200 = ( (~ Pkey_114_)  &  n721  &  n722 ) | ( n13  &  n721  &  n722 ) ;
 assign N_N2812 = ( (~ n200) ) ;
 assign n201 = ( (~ Pkey_122_)  &  n718  &  n719 ) | ( n13  &  n718  &  n719 ) ;
 assign N_N2813 = ( (~ n201) ) ;
 assign n202 = ( (~ Pkey_65_)  &  n715  &  n716 ) | ( n13  &  n715  &  n716 ) ;
 assign N_N2814 = ( (~ n202) ) ;
 assign n203 = ( (~ Pkey_73_)  &  n712  &  n713 ) | ( n13  &  n712  &  n713 ) ;
 assign N_N2815 = ( (~ n203) ) ;
 assign n204 = ( (~ Pkey_81_)  &  n709  &  n710 ) | ( n13  &  n709  &  n710 ) ;
 assign N_N2816 = ( (~ n204) ) ;
 assign n205 = ( (~ Pkey_89_)  &  n706  &  n707 ) | ( n13  &  n706  &  n707 ) ;
 assign N_N2817 = ( (~ n205) ) ;
 assign n206 = ( (~ Pkey_97_)  &  n703  &  n704 ) | ( n13  &  n703  &  n704 ) ;
 assign N_N2818 = ( (~ n206) ) ;
 assign n207 = ( (~ Pkey_105_)  &  n700  &  n701 ) | ( n13  &  n700  &  n701 ) ;
 assign N_N2819 = ( (~ n207) ) ;
 assign n208 = ( (~ Pkey_113_)  &  n697  &  n698 ) | ( n13  &  n697  &  n698 ) ;
 assign N_N2820 = ( (~ n208) ) ;
 assign n209 = ( (~ Pkey_121_)  &  n694  &  n695 ) | ( n13  &  n694  &  n695 ) ;
 assign N_N2822 = ( (~ n209) ) ;
 assign n210 = ( (~ Pkey_64_)  &  n691  &  n692 ) | ( n13  &  n691  &  n692 ) ;
 assign N_N2823 = ( (~ n210) ) ;
 assign n211 = ( (~ Pkey_72_)  &  n688  &  n689 ) | ( n13  &  n688  &  n689 ) ;
 assign N_N2824 = ( (~ n211) ) ;
 assign n212 = ( (~ Pkey_80_)  &  n685  &  n686 ) | ( n13  &  n685  &  n686 ) ;
 assign N_N2825 = ( (~ n212) ) ;
 assign n213 = ( (~ Pkey_88_)  &  n682  &  n683 ) | ( n13  &  n682  &  n683 ) ;
 assign N_N2826 = ( (~ n213) ) ;
 assign n214 = ( (~ Pkey_96_)  &  n679  &  n680 ) | ( n13  &  n679  &  n680 ) ;
 assign N_N2827 = ( (~ n214) ) ;
 assign n215 = ( (~ Pkey_104_)  &  n676  &  n677 ) | ( n13  &  n676  &  n677 ) ;
 assign N_N2828 = ( (~ n215) ) ;
 assign n216 = ( (~ Pkey_112_)  &  n673  &  n674 ) | ( n13  &  n673  &  n674 ) ;
 assign N_N2829 = ( (~ n216) ) ;
 assign n217 = ( (~ Pkey_120_)  &  n670  &  n671 ) | ( n13  &  n670  &  n671 ) ;
 assign N_N2830 = ( (~ n217) ) ;
 assign n218 = ( (~ Pkey_35_)  &  n667  &  n668 ) | ( n13  &  n667  &  n668 ) ;
 assign N_N2831 = ( (~ n218) ) ;
 assign n219 = ( (~ Pkey_43_)  &  n664  &  n665 ) | ( n13  &  n664  &  n665 ) ;
 assign N_N2832 = ( (~ n219) ) ;
 assign n220 = ( (~ Pkey_51_)  &  n661  &  n662 ) | ( n13  &  n661  &  n662 ) ;
 assign N_N2833 = ( (~ n220) ) ;
 assign n221 = ( (~ Pkey_59_)  &  n658  &  n659 ) | ( n13  &  n658  &  n659 ) ;
 assign N_N2835 = ( (~ n221) ) ;
 assign n222 = ( (~ Pkey_2_)  &  n655  &  n656 ) | ( n13  &  n655  &  n656 ) ;
 assign N_N2836 = ( (~ n222) ) ;
 assign n223 = ( (~ Pkey_10_)  &  n652  &  n653 ) | ( n13  &  n652  &  n653 ) ;
 assign N_N2837 = ( (~ n223) ) ;
 assign n224 = ( (~ Pkey_18_)  &  n649  &  n650 ) | ( n13  &  n649  &  n650 ) ;
 assign N_N2839 = ( (~ n224) ) ;
 assign n225 = ( (~ Pkey_26_)  &  n646  &  n647 ) | ( n13  &  n646  &  n647 ) ;
 assign N_N2840 = ( (~ n225) ) ;
 assign n226 = ( (~ Pkey_34_)  &  n643  &  n644 ) | ( n13  &  n643  &  n644 ) ;
 assign N_N2841 = ( (~ n226) ) ;
 assign n227 = ( (~ Pkey_42_)  &  n640  &  n641 ) | ( n13  &  n640  &  n641 ) ;
 assign N_N2842 = ( (~ n227) ) ;
 assign n228 = ( (~ Pkey_50_)  &  n637  &  n638 ) | ( n13  &  n637  &  n638 ) ;
 assign N_N2844 = ( (~ n228) ) ;
 assign n229 = ( (~ Pkey_58_)  &  n634  &  n635 ) | ( n13  &  n634  &  n635 ) ;
 assign N_N2845 = ( (~ n229) ) ;
 assign n230 = ( (~ Pkey_1_)  &  n631  &  n632 ) | ( n13  &  n631  &  n632 ) ;
 assign N_N2846 = ( (~ n230) ) ;
 assign n231 = ( (~ Pkey_9_)  &  n628  &  n629 ) | ( n13  &  n628  &  n629 ) ;
 assign N_N2847 = ( (~ n231) ) ;
 assign n232 = ( (~ Pkey_17_)  &  n625  &  n626 ) | ( n13  &  n625  &  n626 ) ;
 assign N_N2848 = ( (~ n232) ) ;
 assign n233 = ( (~ Pkey_25_)  &  n622  &  n623 ) | ( n13  &  n622  &  n623 ) ;
 assign N_N2849 = ( (~ n233) ) ;
 assign n234 = ( (~ Pkey_33_)  &  n619  &  n620 ) | ( n13  &  n619  &  n620 ) ;
 assign N_N2850 = ( (~ n234) ) ;
 assign n235 = ( (~ Pkey_41_)  &  n616  &  n617 ) | ( n13  &  n616  &  n617 ) ;
 assign N_N2851 = ( (~ n235) ) ;
 assign n236 = ( (~ Pkey_49_)  &  n613  &  n614 ) | ( n13  &  n613  &  n614 ) ;
 assign N_N2852 = ( (~ n236) ) ;
 assign n237 = ( (~ Pkey_57_)  &  n610  &  n611 ) | ( n13  &  n610  &  n611 ) ;
 assign N_N2854 = ( (~ n237) ) ;
 assign n238 = ( (~ Pkey_0_)  &  n607  &  n608 ) | ( n13  &  n607  &  n608 ) ;
 assign N_N2855 = ( (~ n238) ) ;
 assign n239 = ( (~ Pkey_8_)  &  n604  &  n605 ) | ( n13  &  n604  &  n605 ) ;
 assign N_N2856 = ( (~ n239) ) ;
 assign n240 = ( (~ Pkey_16_)  &  n601  &  n602 ) | ( n13  &  n601  &  n602 ) ;
 assign N_N2857 = ( (~ n240) ) ;
 assign n241 = ( (~ Pkey_24_)  &  n598  &  n599 ) | ( n13  &  n598  &  n599 ) ;
 assign N_N2858 = ( (~ n241) ) ;
 assign n242 = ( (~ Pkey_32_)  &  n595  &  n596 ) | ( n13  &  n595  &  n596 ) ;
 assign N_N2859 = ( (~ n242) ) ;
 assign n243 = ( (~ Pkey_40_)  &  n592  &  n593 ) | ( n13  &  n592  &  n593 ) ;
 assign N_N2860 = ( (~ n243) ) ;
 assign n244 = ( (~ Pkey_48_)  &  n589  &  n590 ) | ( n13  &  n589  &  n590 ) ;
 assign N_N2861 = ( (~ n244) ) ;
 assign n248 = ( Pcount_1_ ) | ( Pcount_2_ ) | ( Pcount_3_ ) ;
 assign n249 = ( Pcount_1_ ) | ( Pcount_2_ ) | ( Pcount_0_ ) ;
 assign n246 = ( (~ Pcount_2_) ) | ( (~ Pcount_1_) ) | ( (~ Pcount_0_) ) ;
 assign n245 = ( (~ Pcount_3_)  &  n248  &  n249 ) | ( n248  &  n249  &  n246 ) ;
 assign n251 = ( (~ Pcount_3_) ) | ( (~ Pcount_2_) ) | ( (~ Pcount_1_) ) | ( Pcount_0_ ) ;
 assign n252 = ( Pcount_3_ ) | ( n246 ) ;
 assign n250 = ( n251  &  n252  &  Pcount_3_ ) | ( n251  &  n252  &  n249 ) ;
 assign n255 = ( (~ PKSi_118_)  &  n1290 ) | ( (~ PKSi_4_)  &  n1290 ) | ( n1166  &  n1290 ) ;
 assign n256 = ( (~ Pkey_62_)  &  n1291 ) | ( n15  &  n1291 ) ;
 assign n258 = ( (~ PKSi_102_)  &  n1292 ) | ( (~ PKSi_23_)  &  n1292 ) | ( n1166  &  n1292 ) ;
 assign n259 = ( (~ Pkey_54_)  &  n1293 ) | ( n15  &  n1293 ) ;
 assign n261 = ( (~ PKSi_98_)  &  n1294 ) | ( (~ PKSi_6_)  &  n1294 ) | ( n1166  &  n1294 ) ;
 assign n262 = ( (~ Pkey_46_)  &  n1295 ) | ( n15  &  n1295 ) ;
 assign n264 = ( (~ PKSi_119_)  &  n1296 ) | ( (~ PKSi_15_)  &  n1296 ) | ( n1166  &  n1296 ) ;
 assign n265 = ( (~ Pkey_38_)  &  n1297 ) | ( n15  &  n1297 ) ;
 assign n267 = ( (~ PKSi_106_)  &  n1298 ) | ( (~ PKSi_5_)  &  n1298 ) | ( n1166  &  n1298 ) ;
 assign n268 = ( (~ Pkey_30_)  &  n1299 ) | ( n15  &  n1299 ) ;
 assign n270 = ( (~ PKSi_112_)  &  n1300 ) | ( (~ PKSi_9_)  &  n1300 ) | ( n1166  &  n1300 ) ;
 assign n271 = ( (~ Pkey_22_)  &  n1301 ) | ( n15  &  n1301 ) ;
 assign n273 = ( (~ PKSi_19_)  &  n1302 ) | ( (~ N_N2986)  &  n1302 ) | ( n1166  &  n1302 ) ;
 assign n274 = ( (~ Pkey_14_)  &  n1303 ) | ( n15  &  n1303 ) ;
 assign n276 = ( (~ PKSi_117_)  &  n1304 ) | ( (~ PKSi_17_)  &  n1304 ) | ( n1166  &  n1304 ) ;
 assign n277 = ( (~ Pkey_6_)  &  n1305 ) | ( n15  &  n1305 ) ;
 assign n279 = ( (~ PKSi_99_)  &  n1306 ) | ( n1166  &  n1306 ) | ( (~ N_N2853)  &  n1306 ) ;
 assign n280 = ( (~ Pkey_61_)  &  n1307 ) | ( n15  &  n1307 ) ;
 assign n282 = ( (~ PKSi_11_)  &  n1308 ) | ( (~ N_N2982)  &  n1308 ) | ( n1166  &  n1308 ) ;
 assign n283 = ( (~ Pkey_53_)  &  n1309 ) | ( n15  &  n1309 ) ;
 assign n285 = ( (~ PKSi_110_)  &  n1310 ) | ( (~ PKSi_2_)  &  n1310 ) | ( n1166  &  n1310 ) ;
 assign n286 = ( (~ Pkey_45_)  &  n1311 ) | ( n15  &  n1311 ) ;
 assign n288 = ( (~ PKSi_103_)  &  n1312 ) | ( (~ PKSi_14_)  &  n1312 ) | ( n1166  &  n1312 ) ;
 assign n289 = ( (~ Pkey_37_)  &  n1313 ) | ( n15  &  n1313 ) ;
 assign n291 = ( (~ PKSi_96_)  &  n1314 ) | ( (~ PKSi_22_)  &  n1314 ) | ( n1166  &  n1314 ) ;
 assign n292 = ( (~ Pkey_29_)  &  n1315 ) | ( n15  &  n1315 ) ;
 assign n294 = ( (~ PKSi_115_)  &  n1316 ) | ( (~ PKSi_0_)  &  n1316 ) | ( n1166  &  n1316 ) ;
 assign n295 = ( (~ Pkey_21_)  &  n1317 ) | ( n15  &  n1317 ) ;
 assign n297 = ( (~ PKSi_8_)  &  n1318 ) | ( (~ N_N2976)  &  n1318 ) | ( n1166  &  n1318 ) ;
 assign n298 = ( (~ Pkey_13_)  &  n1319 ) | ( n15  &  n1319 ) ;
 assign n300 = ( (~ PKSi_108_)  &  n1320 ) | ( (~ PKSi_18_)  &  n1320 ) | ( n1166  &  n1320 ) ;
 assign n301 = ( (~ Pkey_5_)  &  n1321 ) | ( n15  &  n1321 ) ;
 assign n303 = ( (~ PKSi_105_)  &  n1322 ) | ( (~ PKSi_1_)  &  n1322 ) | ( n1166  &  n1322 ) ;
 assign n304 = ( (~ Pkey_60_)  &  n1323 ) | ( n15  &  n1323 ) ;
 assign n306 = ( (~ PKSi_114_)  &  n1324 ) | ( n1166  &  n1324 ) | ( (~ N_N2843)  &  n1324 ) ;
 assign n307 = ( (~ Pkey_52_)  &  n1325 ) | ( n15  &  n1325 ) ;
 assign n309 = ( (~ PKSi_100_)  &  n1326 ) | ( (~ PKSi_13_)  &  n1326 ) | ( n1166  &  n1326 ) ;
 assign n310 = ( (~ Pkey_44_)  &  n1327 ) | ( n15  &  n1327 ) ;
 assign n312 = ( (~ PKSi_107_)  &  n1328 ) | ( (~ PKSi_21_)  &  n1328 ) | ( n1166  &  n1328 ) ;
 assign n313 = ( (~ Pkey_36_)  &  n1329 ) | ( n15  &  n1329 ) ;
 assign n315 = ( (~ PKSi_109_)  &  n1330 ) | ( (~ PKSi_10_)  &  n1330 ) | ( n1166  &  n1330 ) ;
 assign n316 = ( (~ Pkey_28_)  &  n1331 ) | ( n15  &  n1331 ) ;
 assign n318 = ( (~ PKSi_116_)  &  n1332 ) | ( n1166  &  n1332 ) | ( (~ N_N2838)  &  n1332 ) ;
 assign n319 = ( (~ Pkey_20_)  &  n1333 ) | ( n15  &  n1333 ) ;
 assign n321 = ( (~ PKSi_104_)  &  n1334 ) | ( (~ PKSi_12_)  &  n1334 ) | ( n1166  &  n1334 ) ;
 assign n322 = ( (~ Pkey_12_)  &  n1335 ) | ( n15  &  n1335 ) ;
 assign n324 = ( (~ PKSi_97_)  &  n1336 ) | ( (~ PKSi_3_)  &  n1336 ) | ( n1166  &  n1336 ) ;
 assign n325 = ( (~ Pkey_4_)  &  n1337 ) | ( n15  &  n1337 ) ;
 assign n327 = ( (~ PKSi_113_)  &  n1338 ) | ( n1166  &  n1338 ) | ( (~ N_N2834)  &  n1338 ) ;
 assign n328 = ( (~ Pkey_27_)  &  n1339 ) | ( n15  &  n1339 ) ;
 assign n330 = ( (~ PKSi_16_)  &  n1340 ) | ( (~ N_N2964)  &  n1340 ) | ( n1166  &  n1340 ) ;
 assign n331 = ( (~ Pkey_19_)  &  n1341 ) | ( n15  &  n1341 ) ;
 assign n333 = ( (~ PKSi_101_)  &  n1342 ) | ( (~ PKSi_20_)  &  n1342 ) | ( n1166  &  n1342 ) ;
 assign n334 = ( (~ Pkey_11_)  &  n1343 ) | ( n15  &  n1343 ) ;
 assign n336 = ( (~ PKSi_111_)  &  n1344 ) | ( (~ PKSi_7_)  &  n1344 ) | ( n1166  &  n1344 ) ;
 assign n337 = ( (~ Pkey_3_)  &  n1345 ) | ( n15  &  n1345 ) ;
 assign n339 = ( (~ PKSi_142_)  &  n1346 ) | ( (~ PKSi_28_)  &  n1346 ) | ( n1166  &  n1346 ) ;
 assign n340 = ( (~ Pkey_126_)  &  n1347 ) | ( n15  &  n1347 ) ;
 assign n342 = ( (~ PKSi_126_)  &  n1348 ) | ( (~ PKSi_47_)  &  n1348 ) | ( n1166  &  n1348 ) ;
 assign n343 = ( (~ Pkey_118_)  &  n1349 ) | ( n15  &  n1349 ) ;
 assign n345 = ( (~ PKSi_122_)  &  n1350 ) | ( (~ PKSi_30_)  &  n1350 ) | ( n1166  &  n1350 ) ;
 assign n346 = ( (~ Pkey_110_)  &  n1351 ) | ( n15  &  n1351 ) ;
 assign n348 = ( (~ wire282)  &  n1352 ) | ( (~ PKSi_39_)  &  n1352 ) | ( n1166  &  n1352 ) ;
 assign n349 = ( (~ Pkey_102_)  &  n1353 ) | ( n15  &  n1353 ) ;
 assign n351 = ( (~ PKSi_130_)  &  n1354 ) | ( (~ PKSi_29_)  &  n1354 ) | ( n1166  &  n1354 ) ;
 assign n352 = ( (~ Pkey_94_)  &  n1355 ) | ( n15  &  n1355 ) ;
 assign n354 = ( (~ PKSi_136_)  &  n1356 ) | ( (~ PKSi_33_)  &  n1356 ) | ( n1166  &  n1356 ) ;
 assign n355 = ( (~ Pkey_86_)  &  n1357 ) | ( n15  &  n1357 ) ;
 assign n357 = ( (~ PKSi_43_)  &  n1358 ) | ( (~ N_N2954)  &  n1358 ) | ( n1166  &  n1358 ) ;
 assign n358 = ( (~ Pkey_78_)  &  n1359 ) | ( n15  &  n1359 ) ;
 assign n360 = ( (~ PKSi_141_)  &  n1360 ) | ( (~ PKSi_41_)  &  n1360 ) | ( n1166  &  n1360 ) ;
 assign n361 = ( (~ Pkey_70_)  &  n1361 ) | ( n15  &  n1361 ) ;
 assign n363 = ( (~ PKSi_123_)  &  n1362 ) | ( n1166  &  n1362 ) | ( (~ N_N2821)  &  n1362 ) ;
 assign n364 = ( (~ Pkey_125_)  &  n1363 ) | ( n15  &  n1363 ) ;
 assign n366 = ( (~ PKSi_35_)  &  n1364 ) | ( (~ N_N2950)  &  n1364 ) | ( n1166  &  n1364 ) ;
 assign n367 = ( (~ Pkey_117_)  &  n1365 ) | ( n15  &  n1365 ) ;
 assign n369 = ( (~ PKSi_134_)  &  n1366 ) | ( (~ PKSi_26_)  &  n1366 ) | ( n1166  &  n1366 ) ;
 assign n370 = ( (~ Pkey_109_)  &  n1367 ) | ( n15  &  n1367 ) ;
 assign n372 = ( (~ PKSi_127_)  &  n1368 ) | ( (~ PKSi_38_)  &  n1368 ) | ( n1166  &  n1368 ) ;
 assign n373 = ( (~ Pkey_101_)  &  n1369 ) | ( n15  &  n1369 ) ;
 assign n375 = ( (~ PKSi_120_)  &  n1370 ) | ( (~ PKSi_46_)  &  n1370 ) | ( n1166  &  n1370 ) ;
 assign n376 = ( (~ Pkey_93_)  &  n1371 ) | ( n15  &  n1371 ) ;
 assign n378 = ( (~ PKSi_24_)  &  n1372 ) | ( (~ N_N2945)  &  n1372 ) | ( n1166  &  n1372 ) ;
 assign n379 = ( (~ Pkey_85_)  &  n1373 ) | ( n15  &  n1373 ) ;
 assign n381 = ( (~ PKSi_32_)  &  n1374 ) | ( (~ N_N2943)  &  n1374 ) | ( n1166  &  n1374 ) ;
 assign n382 = ( (~ Pkey_77_)  &  n1375 ) | ( n15  &  n1375 ) ;
 assign n384 = ( (~ PKSi_132_)  &  n1376 ) | ( (~ PKSi_42_)  &  n1376 ) | ( n1166  &  n1376 ) ;
 assign n385 = ( (~ Pkey_69_)  &  n1377 ) | ( n15  &  n1377 ) ;
 assign n387 = ( (~ PKSi_129_)  &  n1378 ) | ( (~ PKSi_25_)  &  n1378 ) | ( n1166  &  n1378 ) ;
 assign n388 = ( (~ Pkey_124_)  &  n1379 ) | ( n15  &  n1379 ) ;
 assign n389 = ( (~ PKSi_138_)  &  n1380 ) | ( n1166  &  n1380 ) | ( (~ N_N2811)  &  n1380 ) ;
 assign n390 = ( (~ Pkey_116_)  &  n1381 ) | ( n15  &  n1381 ) ;
 assign n392 = ( (~ PKSi_124_)  &  n1382 ) | ( (~ PKSi_37_)  &  n1382 ) | ( n1166  &  n1382 ) ;
 assign n393 = ( (~ Pkey_44_)  &  n1383 ) | ( n15  &  n1383 ) ;
 assign n395 = ( (~ PKSi_131_)  &  n1384 ) | ( (~ PKSi_45_)  &  n1384 ) | ( n1166  &  n1384 ) ;
 assign n396 = ( (~ Pkey_100_)  &  n1385 ) | ( n15  &  n1385 ) ;
 assign n398 = ( (~ PKSi_133_)  &  n1386 ) | ( (~ PKSi_34_)  &  n1386 ) | ( n1166  &  n1386 ) ;
 assign n399 = ( (~ Pkey_92_)  &  n1387 ) | ( n15  &  n1387 ) ;
 assign n401 = ( (~ PKSi_140_)  &  n1388 ) | ( n1166  &  n1388 ) | ( (~ N_N2806)  &  n1388 ) ;
 assign n402 = ( (~ Pkey_84_)  &  n1389 ) | ( n15  &  n1389 ) ;
 assign n404 = ( (~ PKSi_128_)  &  n1390 ) | ( (~ PKSi_36_)  &  n1390 ) | ( n1166  &  n1390 ) ;
 assign n405 = ( (~ Pkey_76_)  &  n1391 ) | ( n15  &  n1391 ) ;
 assign n407 = ( (~ PKSi_121_)  &  n1392 ) | ( (~ PKSi_27_)  &  n1392 ) | ( n1166  &  n1392 ) ;
 assign n408 = ( (~ Pkey_68_)  &  n1393 ) | ( n15  &  n1393 ) ;
 assign n410 = ( (~ PKSi_137_)  &  n1394 ) | ( n1166  &  n1394 ) | ( (~ N_N2802)  &  n1394 ) ;
 assign n411 = ( (~ Pkey_91_)  &  n1395 ) | ( n15  &  n1395 ) ;
 assign n413 = ( (~ PKSi_40_)  &  n1396 ) | ( (~ N_N2931)  &  n1396 ) | ( n1166  &  n1396 ) ;
 assign n414 = ( (~ Pkey_83_)  &  n1397 ) | ( n15  &  n1397 ) ;
 assign n416 = ( (~ PKSi_125_)  &  n1398 ) | ( (~ PKSi_44_)  &  n1398 ) | ( n1166  &  n1398 ) ;
 assign n417 = ( (~ Pkey_75_)  &  n1399 ) | ( n15  &  n1399 ) ;
 assign n419 = ( (~ PKSi_135_)  &  n1400 ) | ( (~ PKSi_31_)  &  n1400 ) | ( n1166  &  n1400 ) ;
 assign n420 = ( (~ Pkey_67_)  &  n1401 ) | ( n15  &  n1401 ) ;
 assign n422 = ( (~ PKSi_166_)  &  n1402 ) | ( (~ PKSi_52_)  &  n1402 ) | ( n1166  &  n1402 ) ;
 assign n423 = ( (~ Pkey_190_)  &  n1403 ) | ( n15  &  n1403 ) ;
 assign n425 = ( (~ PKSi_150_)  &  n1404 ) | ( (~ PKSi_71_)  &  n1404 ) | ( n1166  &  n1404 ) ;
 assign n426 = ( (~ Pkey_182_)  &  n1405 ) | ( n15  &  n1405 ) ;
 assign n428 = ( (~ PKSi_146_)  &  n1406 ) | ( (~ PKSi_54_)  &  n1406 ) | ( n1166  &  n1406 ) ;
 assign n429 = ( (~ Pkey_174_)  &  n1407 ) | ( n15  &  n1407 ) ;
 assign n431 = ( (~ PKSi_167_)  &  n1408 ) | ( (~ PKSi_63_)  &  n1408 ) | ( n1166  &  n1408 ) ;
 assign n432 = ( (~ Pkey_166_)  &  n1409 ) | ( n15  &  n1409 ) ;
 assign n434 = ( (~ PKSi_154_)  &  n1410 ) | ( (~ PKSi_53_)  &  n1410 ) | ( n1166  &  n1410 ) ;
 assign n435 = ( (~ Pkey_158_)  &  n1411 ) | ( n15  &  n1411 ) ;
 assign n437 = ( (~ PKSi_160_)  &  n1412 ) | ( (~ PKSi_57_)  &  n1412 ) | ( n1166  &  n1412 ) ;
 assign n438 = ( (~ Pkey_150_)  &  n1413 ) | ( n15  &  n1413 ) ;
 assign n440 = ( (~ PKSi_67_)  &  n1414 ) | ( (~ N_N2921)  &  n1414 ) | ( n1166  &  n1414 ) ;
 assign n441 = ( (~ Pkey_142_)  &  n1415 ) | ( n15  &  n1415 ) ;
 assign n443 = ( (~ PKSi_165_)  &  n1416 ) | ( (~ PKSi_65_)  &  n1416 ) | ( n1166  &  n1416 ) ;
 assign n444 = ( (~ Pkey_134_)  &  n1417 ) | ( n15  &  n1417 ) ;
 assign n446 = ( (~ PKSi_147_)  &  n1418 ) | ( n1166  &  n1418 ) | ( (~ N_N2789)  &  n1418 ) ;
 assign n447 = ( (~ Pkey_189_)  &  n1419 ) | ( n15  &  n1419 ) ;
 assign n449 = ( (~ PKSi_59_)  &  n1420 ) | ( (~ N_N2917)  &  n1420 ) | ( n1166  &  n1420 ) ;
 assign n450 = ( (~ Pkey_181_)  &  n1421 ) | ( n15  &  n1421 ) ;
 assign n452 = ( (~ PKSi_158_)  &  n1422 ) | ( (~ PKSi_50_)  &  n1422 ) | ( n1166  &  n1422 ) ;
 assign n453 = ( (~ Pkey_173_)  &  n1423 ) | ( n15  &  n1423 ) ;
 assign n455 = ( (~ PKSi_151_)  &  n1424 ) | ( (~ PKSi_62_)  &  n1424 ) | ( n1166  &  n1424 ) ;
 assign n456 = ( (~ Pkey_165_)  &  n1425 ) | ( n15  &  n1425 ) ;
 assign n458 = ( (~ PKSi_144_)  &  n1426 ) | ( (~ PKSi_70_)  &  n1426 ) | ( n1166  &  n1426 ) ;
 assign n459 = ( (~ Pkey_157_)  &  n1427 ) | ( n15  &  n1427 ) ;
 assign n461 = ( (~ PKSi_163_)  &  n1428 ) | ( (~ PKSi_48_)  &  n1428 ) | ( n1166  &  n1428 ) ;
 assign n462 = ( (~ Pkey_149_)  &  n1429 ) | ( n15  &  n1429 ) ;
 assign n464 = ( (~ PKSi_153_)  &  n1430 ) | ( (~ PKSi_56_)  &  n1430 ) | ( n1166  &  n1430 ) ;
 assign n465 = ( (~ Pkey_141_)  &  n1431 ) | ( n15  &  n1431 ) ;
 assign n467 = ( (~ PKSi_156_)  &  n1432 ) | ( (~ PKSi_66_)  &  n1432 ) | ( n1166  &  n1432 ) ;
 assign n468 = ( (~ Pkey_133_)  &  n1433 ) | ( n15  &  n1433 ) ;
 assign n470 = ( (~ PKSi_49_)  &  n1434 ) | ( (~ N_N2909)  &  n1434 ) | ( n1166  &  n1434 ) ;
 assign n471 = ( (~ Pkey_188_)  &  n1435 ) | ( n15  &  n1435 ) ;
 assign n473 = ( (~ PKSi_162_)  &  n1436 ) | ( n1166  &  n1436 ) | ( (~ N_N2779)  &  n1436 ) ;
 assign n474 = ( (~ Pkey_180_)  &  n1437 ) | ( n15  &  n1437 ) ;
 assign n476 = ( (~ PKSi_148_)  &  n1438 ) | ( (~ PKSi_61_)  &  n1438 ) | ( n1166  &  n1438 ) ;
 assign n477 = ( (~ Pkey_172_)  &  n1439 ) | ( n15  &  n1439 ) ;
 assign n479 = ( (~ PKSi_155_)  &  n1440 ) | ( (~ PKSi_69_)  &  n1440 ) | ( n1166  &  n1440 ) ;
 assign n480 = ( (~ Pkey_164_)  &  n1441 ) | ( n15  &  n1441 ) ;
 assign n482 = ( (~ PKSi_157_)  &  n1442 ) | ( (~ PKSi_58_)  &  n1442 ) | ( n1166  &  n1442 ) ;
 assign n483 = ( (~ Pkey_156_)  &  n1443 ) | ( n15  &  n1443 ) ;
 assign n485 = ( (~ PKSi_164_)  &  n1444 ) | ( n1166  &  n1444 ) | ( (~ N_N2774)  &  n1444 ) ;
 assign n486 = ( (~ Pkey_148_)  &  n1445 ) | ( n15  &  n1445 ) ;
 assign n488 = ( (~ PKSi_152_)  &  n1446 ) | ( (~ PKSi_60_)  &  n1446 ) | ( n1166  &  n1446 ) ;
 assign n489 = ( (~ Pkey_140_)  &  n1447 ) | ( n15  &  n1447 ) ;
 assign n491 = ( (~ PKSi_145_)  &  n1448 ) | ( (~ PKSi_51_)  &  n1448 ) | ( n1166  &  n1448 ) ;
 assign n492 = ( (~ Pkey_132_)  &  n1449 ) | ( n15  &  n1449 ) ;
 assign n494 = ( (~ PKSi_161_)  &  n1450 ) | ( n1166  &  n1450 ) | ( (~ N_N2770)  &  n1450 ) ;
 assign n495 = ( (~ Pkey_155_)  &  n1451 ) | ( n15  &  n1451 ) ;
 assign n497 = ( (~ PKSi_64_)  &  n1452 ) | ( (~ N_N2899)  &  n1452 ) | ( n1166  &  n1452 ) ;
 assign n498 = ( (~ Pkey_147_)  &  n1453 ) | ( n15  &  n1453 ) ;
 assign n500 = ( (~ PKSi_149_)  &  n1454 ) | ( (~ PKSi_68_)  &  n1454 ) | ( n1166  &  n1454 ) ;
 assign n501 = ( (~ Pkey_139_)  &  n1455 ) | ( n15  &  n1455 ) ;
 assign n503 = ( (~ PKSi_159_)  &  n1456 ) | ( (~ PKSi_55_)  &  n1456 ) | ( n1166  &  n1456 ) ;
 assign n504 = ( (~ Pkey_131_)  &  n1457 ) | ( n15  &  n1457 ) ;
 assign n506 = ( (~ PKSi_190_)  &  n1458 ) | ( (~ PKSi_76_)  &  n1458 ) | ( n1166  &  n1458 ) ;
 assign n507 = ( (~ Pkey_254_)  &  n1459 ) | ( n15  &  n1459 ) ;
 assign n509 = ( (~ PKSi_174_)  &  n1460 ) | ( (~ PKSi_95_)  &  n1460 ) | ( n1166  &  n1460 ) ;
 assign n510 = ( (~ Pkey_246_)  &  n1461 ) | ( n15  &  n1461 ) ;
 assign n512 = ( (~ PKSi_170_)  &  n1462 ) | ( (~ PKSi_78_)  &  n1462 ) | ( n1166  &  n1462 ) ;
 assign n513 = ( (~ Pkey_238_)  &  n1463 ) | ( n15  &  n1463 ) ;
 assign n515 = ( (~ wire234)  &  n1464 ) | ( (~ PKSi_87_)  &  n1464 ) | ( n1166  &  n1464 ) ;
 assign n516 = ( (~ Pkey_230_)  &  n1465 ) | ( n15  &  n1465 ) ;
 assign n518 = ( (~ PKSi_178_)  &  n1466 ) | ( (~ PKSi_77_)  &  n1466 ) | ( n1166  &  n1466 ) ;
 assign n519 = ( (~ Pkey_222_)  &  n1467 ) | ( n15  &  n1467 ) ;
 assign n521 = ( (~ PKSi_184_)  &  n1468 ) | ( (~ PKSi_81_)  &  n1468 ) | ( n1166  &  n1468 ) ;
 assign n522 = ( (~ Pkey_214_)  &  n1469 ) | ( n15  &  n1469 ) ;
 assign n524 = ( (~ PKSi_91_)  &  n1470 ) | ( (~ N_N2889)  &  n1470 ) | ( n1166  &  n1470 ) ;
 assign n525 = ( (~ Pkey_206_)  &  n1471 ) | ( n15  &  n1471 ) ;
 assign n527 = ( (~ PKSi_189_)  &  n1472 ) | ( (~ PKSi_89_)  &  n1472 ) | ( n1166  &  n1472 ) ;
 assign n528 = ( (~ Pkey_198_)  &  n1473 ) | ( n15  &  n1473 ) ;
 assign n530 = ( (~ PKSi_171_)  &  n1474 ) | ( n1166  &  n1474 ) | ( (~ N_N2757)  &  n1474 ) ;
 assign n531 = ( (~ Pkey_253_)  &  n1475 ) | ( n15  &  n1475 ) ;
 assign n533 = ( (~ PKSi_83_)  &  n1476 ) | ( (~ N_N2885)  &  n1476 ) | ( n1166  &  n1476 ) ;
 assign n534 = ( (~ Pkey_245_)  &  n1477 ) | ( n15  &  n1477 ) ;
 assign n536 = ( (~ PKSi_182_)  &  n1478 ) | ( (~ PKSi_74_)  &  n1478 ) | ( n1166  &  n1478 ) ;
 assign n537 = ( (~ Pkey_237_)  &  n1479 ) | ( n15  &  n1479 ) ;
 assign n539 = ( (~ PKSi_175_)  &  n1480 ) | ( (~ PKSi_86_)  &  n1480 ) | ( n1166  &  n1480 ) ;
 assign n540 = ( (~ Pkey_229_)  &  n1481 ) | ( n15  &  n1481 ) ;
 assign n542 = ( (~ PKSi_94_)  &  n1482 ) | ( (~ N_N2881)  &  n1482 ) | ( n1166  &  n1482 ) ;
 assign n543 = ( (~ Pkey_221_)  &  n1483 ) | ( n15  &  n1483 ) ;
 assign n545 = ( (~ PKSi_72_)  &  n1484 ) | ( (~ N_N2879)  &  n1484 ) | ( n1166  &  n1484 ) ;
 assign n546 = ( (~ Pkey_213_)  &  n1485 ) | ( n15  &  n1485 ) ;
 assign n548 = ( (~ PKSi_80_)  &  n1486 ) | ( (~ N_N2877)  &  n1486 ) | ( n1166  &  n1486 ) ;
 assign n549 = ( (~ Pkey_205_)  &  n1487 ) | ( n15  &  n1487 ) ;
 assign n551 = ( (~ PKSi_180_)  &  n1488 ) | ( n1166  &  n1488 ) | ( (~ N_N2749)  &  n1488 ) ;
 assign n552 = ( (~ Pkey_197_)  &  n1489 ) | ( n15  &  n1489 ) ;
 assign n554 = ( (~ PKSi_177_)  &  n1490 ) | ( (~ PKSi_73_)  &  n1490 ) | ( n1166  &  n1490 ) ;
 assign n555 = ( (~ Pkey_252_)  &  n1491 ) | ( n15  &  n1491 ) ;
 assign n556 = ( (~ PKSi_186_)  &  n1492 ) | ( n1166  &  n1492 ) | ( (~ N_N2746)  &  n1492 ) ;
 assign n557 = ( (~ Pkey_244_)  &  n1493 ) | ( n15  &  n1493 ) ;
 assign n559 = ( (~ PKSi_172_)  &  n1494 ) | ( (~ PKSi_85_)  &  n1494 ) | ( n1166  &  n1494 ) ;
 assign n560 = ( (~ Pkey_172_)  &  n1495 ) | ( n15  &  n1495 ) ;
 assign n562 = ( (~ PKSi_179_)  &  n1496 ) | ( (~ PKSi_93_)  &  n1496 ) | ( n1166  &  n1496 ) ;
 assign n563 = ( (~ Pkey_228_)  &  n1497 ) | ( n15  &  n1497 ) ;
 assign n565 = ( (~ wire253)  &  n1498 ) | ( (~ PKSi_82_)  &  n1498 ) | ( n1166  &  n1498 ) ;
 assign n566 = ( (~ Pkey_220_)  &  n1499 ) | ( n15  &  n1499 ) ;
 assign n568 = ( (~ PKSi_188_)  &  n1500 ) | ( n1166  &  n1500 ) | ( (~ N_N2741)  &  n1500 ) ;
 assign n569 = ( (~ Pkey_212_)  &  n1501 ) | ( n15  &  n1501 ) ;
 assign n571 = ( (~ PKSi_176_)  &  n1502 ) | ( (~ PKSi_84_)  &  n1502 ) | ( n1166  &  n1502 ) ;
 assign n572 = ( (~ Pkey_204_)  &  n1503 ) | ( n15  &  n1503 ) ;
 assign n574 = ( (~ PKSi_169_)  &  n1504 ) | ( (~ PKSi_75_)  &  n1504 ) | ( n1166  &  n1504 ) ;
 assign n575 = ( (~ Pkey_196_)  &  n1505 ) | ( n15  &  n1505 ) ;
 assign n577 = ( (~ PKSi_185_)  &  n1506 ) | ( n1166  &  n1506 ) | ( (~ N_N2737)  &  n1506 ) ;
 assign n578 = ( (~ Pkey_219_)  &  n1507 ) | ( n15  &  n1507 ) ;
 assign n580 = ( (~ wire333)  &  n1508 ) | ( (~ N_N2865)  &  n1508 ) | ( n1166  &  n1508 ) ;
 assign n581 = ( (~ Pkey_211_)  &  n1509 ) | ( n15  &  n1509 ) ;
 assign n583 = ( (~ PKSi_173_)  &  n1510 ) | ( (~ PKSi_92_)  &  n1510 ) | ( n1166  &  n1510 ) ;
 assign n584 = ( (~ Pkey_203_)  &  n1511 ) | ( n15  &  n1511 ) ;
 assign n586 = ( (~ PKSi_183_)  &  n1512 ) | ( (~ PKSi_79_)  &  n1512 ) | ( n1166  &  n1512 ) ;
 assign n587 = ( (~ Pkey_195_)  &  n1513 ) | ( n15  &  n1513 ) ;
 assign n589 = ( n940  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n940  &  n1514 ) | ( n1286  &  n1514 ) ;
 assign n590 = ( (~ Pkey_56_)  &  n1516 ) | ( n15  &  n1516 ) ;
 assign n592 = ( n942  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n942  &  n1517 ) | ( n1286  &  n1517 ) ;
 assign n593 = ( (~ Pkey_48_)  &  n1518 ) | ( n15  &  n1518 ) ;
 assign n595 = ( n944  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n944  &  n1519 ) | ( n1286  &  n1519 ) ;
 assign n596 = ( (~ Pkey_40_)  &  n1520 ) | ( n15  &  n1520 ) ;
 assign n598 = ( n946  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n946  &  n1521 ) | ( n1286  &  n1521 ) ;
 assign n599 = ( (~ Pkey_32_)  &  n1522 ) | ( n15  &  n1522 ) ;
 assign n601 = ( n948  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n948  &  n1523 ) | ( n1286  &  n1523 ) ;
 assign n602 = ( (~ Pkey_24_)  &  n1524 ) | ( n15  &  n1524 ) ;
 assign n604 = ( n950  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n950  &  n1525 ) | ( n1286  &  n1525 ) ;
 assign n605 = ( (~ Pkey_16_)  &  n1526 ) | ( n15  &  n1526 ) ;
 assign n607 = ( n952  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n952  &  n1527 ) | ( n1286  &  n1527 ) ;
 assign n608 = ( (~ Pkey_8_)  &  n1528 ) | ( n15  &  n1528 ) ;
 assign n610 = ( n954  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n954  &  n1529 ) | ( n1286  &  n1529 ) ;
 assign n611 = ( (~ Pkey_0_)  &  n1530 ) | ( n15  &  n1530 ) ;
 assign n613 = ( n956  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n956  &  n1531 ) | ( n1286  &  n1531 ) ;
 assign n614 = ( (~ Pkey_57_)  &  n1532 ) | ( n15  &  n1532 ) ;
 assign n616 = ( n958  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n958  &  n1533 ) | ( n1286  &  n1533 ) ;
 assign n617 = ( (~ Pkey_49_)  &  n1534 ) | ( n15  &  n1534 ) ;
 assign n619 = ( n960  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n960  &  n1535 ) | ( n1286  &  n1535 ) ;
 assign n620 = ( (~ Pkey_41_)  &  n1536 ) | ( n15  &  n1536 ) ;
 assign n622 = ( n962  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n962  &  n1537 ) | ( n1286  &  n1537 ) ;
 assign n623 = ( (~ Pkey_33_)  &  n1538 ) | ( n15  &  n1538 ) ;
 assign n625 = ( n964  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n964  &  n1539 ) | ( n1286  &  n1539 ) ;
 assign n626 = ( (~ Pkey_25_)  &  n1540 ) | ( n15  &  n1540 ) ;
 assign n628 = ( n966  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n966  &  n1541 ) | ( n1286  &  n1541 ) ;
 assign n629 = ( (~ Pkey_17_)  &  n1542 ) | ( n15  &  n1542 ) ;
 assign n631 = ( n968  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n968  &  n1543 ) | ( n1286  &  n1543 ) ;
 assign n632 = ( (~ Pkey_9_)  &  n1544 ) | ( n15  &  n1544 ) ;
 assign n634 = ( n970  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n970  &  n1545 ) | ( n1286  &  n1545 ) ;
 assign n635 = ( (~ Pkey_1_)  &  n1546 ) | ( n15  &  n1546 ) ;
 assign n637 = ( n972  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n972  &  n1547 ) | ( n1286  &  n1547 ) ;
 assign n638 = ( (~ Pkey_58_)  &  n1548 ) | ( n15  &  n1548 ) ;
 assign n640 = ( n974  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n974  &  n1549 ) | ( n1286  &  n1549 ) ;
 assign n641 = ( (~ Pkey_50_)  &  n1550 ) | ( n15  &  n1550 ) ;
 assign n643 = ( n976  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n976  &  n1551 ) | ( n1286  &  n1551 ) ;
 assign n644 = ( (~ Pkey_42_)  &  n1552 ) | ( n15  &  n1552 ) ;
 assign n646 = ( n978  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n978  &  n1553 ) | ( n1286  &  n1553 ) ;
 assign n647 = ( (~ Pkey_34_)  &  n1554 ) | ( n15  &  n1554 ) ;
 assign n649 = ( n980  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n980  &  n1555 ) | ( n1286  &  n1555 ) ;
 assign n650 = ( (~ Pkey_26_)  &  n1556 ) | ( n15  &  n1556 ) ;
 assign n652 = ( n982  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n982  &  n1557 ) | ( n1286  &  n1557 ) ;
 assign n653 = ( (~ Pkey_18_)  &  n1558 ) | ( n15  &  n1558 ) ;
 assign n655 = ( n984  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n984  &  n1559 ) | ( n1286  &  n1559 ) ;
 assign n656 = ( (~ Pkey_10_)  &  n1560 ) | ( n15  &  n1560 ) ;
 assign n658 = ( n986  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n986  &  n1561 ) | ( n1286  &  n1561 ) ;
 assign n659 = ( (~ Pkey_2_)  &  n1562 ) | ( n15  &  n1562 ) ;
 assign n661 = ( n988  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n988  &  n1563 ) | ( n1286  &  n1563 ) ;
 assign n662 = ( (~ Pkey_59_)  &  n1564 ) | ( n15  &  n1564 ) ;
 assign n664 = ( n990  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n990  &  n1565 ) | ( n1286  &  n1565 ) ;
 assign n665 = ( (~ Pkey_51_)  &  n1566 ) | ( n15  &  n1566 ) ;
 assign n667 = ( n992  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n992  &  n1567 ) | ( n1286  &  n1567 ) ;
 assign n668 = ( (~ Pkey_43_)  &  n1568 ) | ( n15  &  n1568 ) ;
 assign n670 = ( n994  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n994  &  n1569 ) | ( n1286  &  n1569 ) ;
 assign n671 = ( (~ Pkey_35_)  &  n1570 ) | ( n15  &  n1570 ) ;
 assign n673 = ( n996  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n996  &  n1571 ) | ( n1286  &  n1571 ) ;
 assign n674 = ( (~ Pkey_120_)  &  n1572 ) | ( n15  &  n1572 ) ;
 assign n676 = ( n998  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n998  &  n1573 ) | ( n1286  &  n1573 ) ;
 assign n677 = ( (~ Pkey_112_)  &  n1574 ) | ( n15  &  n1574 ) ;
 assign n679 = ( n1000  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1000  &  n1575 ) | ( n1286  &  n1575 ) ;
 assign n680 = ( (~ Pkey_104_)  &  n1576 ) | ( n15  &  n1576 ) ;
 assign n682 = ( n1002  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1002  &  n1577 ) | ( n1286  &  n1577 ) ;
 assign n683 = ( (~ Pkey_96_)  &  n1578 ) | ( n15  &  n1578 ) ;
 assign n685 = ( n1004  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1004  &  n1579 ) | ( n1286  &  n1579 ) ;
 assign n686 = ( (~ Pkey_88_)  &  n1580 ) | ( n15  &  n1580 ) ;
 assign n688 = ( n1006  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1006  &  n1581 ) | ( n1286  &  n1581 ) ;
 assign n689 = ( (~ Pkey_80_)  &  n1582 ) | ( n15  &  n1582 ) ;
 assign n691 = ( n1008  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1008  &  n1583 ) | ( n1286  &  n1583 ) ;
 assign n692 = ( (~ Pkey_72_)  &  n1584 ) | ( n15  &  n1584 ) ;
 assign n694 = ( n1010  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1010  &  n1585 ) | ( n1286  &  n1585 ) ;
 assign n695 = ( (~ Pkey_64_)  &  n1586 ) | ( n15  &  n1586 ) ;
 assign n697 = ( n1012  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1012  &  n1587 ) | ( n1286  &  n1587 ) ;
 assign n698 = ( (~ Pkey_121_)  &  n1588 ) | ( n15  &  n1588 ) ;
 assign n700 = ( n1014  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1014  &  n1589 ) | ( n1286  &  n1589 ) ;
 assign n701 = ( (~ Pkey_113_)  &  n1590 ) | ( n15  &  n1590 ) ;
 assign n703 = ( n1016  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1016  &  n1591 ) | ( n1286  &  n1591 ) ;
 assign n704 = ( (~ Pkey_105_)  &  n1592 ) | ( n15  &  n1592 ) ;
 assign n706 = ( n1018  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1018  &  n1593 ) | ( n1286  &  n1593 ) ;
 assign n707 = ( (~ Pkey_97_)  &  n1594 ) | ( n15  &  n1594 ) ;
 assign n709 = ( n1020  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1020  &  n1595 ) | ( n1286  &  n1595 ) ;
 assign n710 = ( (~ Pkey_89_)  &  n1596 ) | ( n15  &  n1596 ) ;
 assign n712 = ( n1022  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1022  &  n1597 ) | ( n1286  &  n1597 ) ;
 assign n713 = ( (~ Pkey_81_)  &  n1598 ) | ( n15  &  n1598 ) ;
 assign n715 = ( n1024  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1024  &  n1599 ) | ( n1286  &  n1599 ) ;
 assign n716 = ( (~ Pkey_73_)  &  n1600 ) | ( n15  &  n1600 ) ;
 assign n718 = ( n1026  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1026  &  n1601 ) | ( n1286  &  n1601 ) ;
 assign n719 = ( (~ Pkey_65_)  &  n1602 ) | ( n15  &  n1602 ) ;
 assign n721 = ( n1028  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1028  &  n1603 ) | ( n1286  &  n1603 ) ;
 assign n722 = ( (~ Pkey_122_)  &  n1604 ) | ( n15  &  n1604 ) ;
 assign n724 = ( n1030  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1030  &  n1605 ) | ( n1286  &  n1605 ) ;
 assign n725 = ( (~ Pkey_114_)  &  n1606 ) | ( n15  &  n1606 ) ;
 assign n727 = ( n1032  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1032  &  n1607 ) | ( n1286  &  n1607 ) ;
 assign n728 = ( (~ Pkey_106_)  &  n1608 ) | ( n15  &  n1608 ) ;
 assign n730 = ( n1034  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1034  &  n1609 ) | ( n1286  &  n1609 ) ;
 assign n731 = ( (~ Pkey_98_)  &  n1610 ) | ( n15  &  n1610 ) ;
 assign n733 = ( n1036  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1036  &  n1611 ) | ( n1286  &  n1611 ) ;
 assign n734 = ( (~ Pkey_90_)  &  n1612 ) | ( n15  &  n1612 ) ;
 assign n736 = ( n1038  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1038  &  n1613 ) | ( n1286  &  n1613 ) ;
 assign n737 = ( (~ Pkey_82_)  &  n1614 ) | ( n15  &  n1614 ) ;
 assign n739 = ( n1040  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1040  &  n1615 ) | ( n1286  &  n1615 ) ;
 assign n740 = ( (~ Pkey_74_)  &  n1616 ) | ( n15  &  n1616 ) ;
 assign n742 = ( n1042  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1042  &  n1617 ) | ( n1286  &  n1617 ) ;
 assign n743 = ( (~ Pkey_66_)  &  n1618 ) | ( n15  &  n1618 ) ;
 assign n745 = ( n1044  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1044  &  n1619 ) | ( n1286  &  n1619 ) ;
 assign n746 = ( (~ Pkey_123_)  &  n1620 ) | ( n15  &  n1620 ) ;
 assign n748 = ( n1046  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1046  &  n1621 ) | ( n1286  &  n1621 ) ;
 assign n749 = ( (~ Pkey_115_)  &  n1622 ) | ( n15  &  n1622 ) ;
 assign n751 = ( n1048  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1048  &  n1623 ) | ( n1286  &  n1623 ) ;
 assign n752 = ( (~ Pkey_107_)  &  n1624 ) | ( n15  &  n1624 ) ;
 assign n754 = ( n1050  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1050  &  n1625 ) | ( n1286  &  n1625 ) ;
 assign n755 = ( (~ Pkey_99_)  &  n1626 ) | ( n15  &  n1626 ) ;
 assign n757 = ( n1052  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1052  &  n1627 ) | ( n1286  &  n1627 ) ;
 assign n758 = ( (~ Pkey_184_)  &  n1628 ) | ( n15  &  n1628 ) ;
 assign n760 = ( n1054  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1054  &  n1629 ) | ( n1286  &  n1629 ) ;
 assign n761 = ( (~ Pkey_176_)  &  n1630 ) | ( n15  &  n1630 ) ;
 assign n763 = ( n1056  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1056  &  n1631 ) | ( n1286  &  n1631 ) ;
 assign n764 = ( (~ Pkey_168_)  &  n1632 ) | ( n15  &  n1632 ) ;
 assign n766 = ( n1058  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1058  &  n1633 ) | ( n1286  &  n1633 ) ;
 assign n767 = ( (~ Pkey_160_)  &  n1634 ) | ( n15  &  n1634 ) ;
 assign n769 = ( n1060  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1060  &  n1635 ) | ( n1286  &  n1635 ) ;
 assign n770 = ( (~ Pkey_152_)  &  n1636 ) | ( n15  &  n1636 ) ;
 assign n772 = ( n1062  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1062  &  n1637 ) | ( n1286  &  n1637 ) ;
 assign n773 = ( (~ Pkey_144_)  &  n1638 ) | ( n15  &  n1638 ) ;
 assign n775 = ( n1064  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1064  &  n1639 ) | ( n1286  &  n1639 ) ;
 assign n776 = ( (~ Pkey_136_)  &  n1640 ) | ( n15  &  n1640 ) ;
 assign n778 = ( n1066  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1066  &  n1641 ) | ( n1286  &  n1641 ) ;
 assign n779 = ( (~ Pkey_128_)  &  n1642 ) | ( n15  &  n1642 ) ;
 assign n781 = ( n1068  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1068  &  n1643 ) | ( n1286  &  n1643 ) ;
 assign n782 = ( (~ Pkey_185_)  &  n1644 ) | ( n15  &  n1644 ) ;
 assign n784 = ( n1070  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1070  &  n1645 ) | ( n1286  &  n1645 ) ;
 assign n785 = ( (~ Pkey_177_)  &  n1646 ) | ( n15  &  n1646 ) ;
 assign n787 = ( n1072  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1072  &  n1647 ) | ( n1286  &  n1647 ) ;
 assign n788 = ( (~ Pkey_169_)  &  n1648 ) | ( n15  &  n1648 ) ;
 assign n790 = ( n1074  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1074  &  n1649 ) | ( n1286  &  n1649 ) ;
 assign n791 = ( (~ Pkey_161_)  &  n1650 ) | ( n15  &  n1650 ) ;
 assign n793 = ( n1076  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1076  &  n1651 ) | ( n1286  &  n1651 ) ;
 assign n794 = ( (~ Pkey_153_)  &  n1652 ) | ( n15  &  n1652 ) ;
 assign n796 = ( n1078  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1078  &  n1653 ) | ( n1286  &  n1653 ) ;
 assign n797 = ( (~ Pkey_145_)  &  n1654 ) | ( n15  &  n1654 ) ;
 assign n799 = ( n1080  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1080  &  n1655 ) | ( n1286  &  n1655 ) ;
 assign n800 = ( (~ Pkey_137_)  &  n1656 ) | ( n15  &  n1656 ) ;
 assign n802 = ( n1082  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1082  &  n1657 ) | ( n1286  &  n1657 ) ;
 assign n803 = ( (~ Pkey_129_)  &  n1658 ) | ( n15  &  n1658 ) ;
 assign n805 = ( n1084  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1084  &  n1659 ) | ( n1286  &  n1659 ) ;
 assign n806 = ( (~ Pkey_186_)  &  n1660 ) | ( n15  &  n1660 ) ;
 assign n808 = ( n1086  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1086  &  n1661 ) | ( n1286  &  n1661 ) ;
 assign n809 = ( (~ Pkey_178_)  &  n1662 ) | ( n15  &  n1662 ) ;
 assign n811 = ( n1088  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1088  &  n1663 ) | ( n1286  &  n1663 ) ;
 assign n812 = ( (~ Pkey_170_)  &  n1664 ) | ( n15  &  n1664 ) ;
 assign n814 = ( n1090  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1090  &  n1665 ) | ( n1286  &  n1665 ) ;
 assign n815 = ( (~ Pkey_162_)  &  n1666 ) | ( n15  &  n1666 ) ;
 assign n817 = ( n1092  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1092  &  n1667 ) | ( n1286  &  n1667 ) ;
 assign n818 = ( (~ Pkey_154_)  &  n1668 ) | ( n15  &  n1668 ) ;
 assign n820 = ( n1094  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1094  &  n1669 ) | ( n1286  &  n1669 ) ;
 assign n821 = ( (~ Pkey_146_)  &  n1670 ) | ( n15  &  n1670 ) ;
 assign n823 = ( n1096  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1096  &  n1671 ) | ( n1286  &  n1671 ) ;
 assign n824 = ( (~ Pkey_138_)  &  n1672 ) | ( n15  &  n1672 ) ;
 assign n826 = ( n1098  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1098  &  n1673 ) | ( n1286  &  n1673 ) ;
 assign n827 = ( (~ Pkey_130_)  &  n1674 ) | ( n15  &  n1674 ) ;
 assign n829 = ( n1100  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1100  &  n1675 ) | ( n1286  &  n1675 ) ;
 assign n830 = ( (~ Pkey_187_)  &  n1676 ) | ( n15  &  n1676 ) ;
 assign n832 = ( n1102  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1102  &  n1677 ) | ( n1286  &  n1677 ) ;
 assign n833 = ( (~ Pkey_179_)  &  n1678 ) | ( n15  &  n1678 ) ;
 assign n835 = ( n1104  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1104  &  n1679 ) | ( n1286  &  n1679 ) ;
 assign n836 = ( (~ Pkey_171_)  &  n1680 ) | ( n15  &  n1680 ) ;
 assign n838 = ( n1106  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1106  &  n1681 ) | ( n1286  &  n1681 ) ;
 assign n839 = ( (~ Pkey_163_)  &  n1682 ) | ( n15  &  n1682 ) ;
 assign n841 = ( n1108  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1108  &  n1683 ) | ( n1286  &  n1683 ) ;
 assign n842 = ( (~ Pkey_248_)  &  n1684 ) | ( n15  &  n1684 ) ;
 assign n844 = ( n1110  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1110  &  n1685 ) | ( n1286  &  n1685 ) ;
 assign n845 = ( (~ Pkey_240_)  &  n1686 ) | ( n15  &  n1686 ) ;
 assign n847 = ( n1112  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1112  &  n1687 ) | ( n1286  &  n1687 ) ;
 assign n848 = ( (~ Pkey_232_)  &  n1688 ) | ( n15  &  n1688 ) ;
 assign n850 = ( n1114  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1114  &  n1689 ) | ( n1286  &  n1689 ) ;
 assign n851 = ( (~ Pkey_224_)  &  n1690 ) | ( n15  &  n1690 ) ;
 assign n853 = ( n1116  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1116  &  n1691 ) | ( n1286  &  n1691 ) ;
 assign n854 = ( (~ Pkey_216_)  &  n1692 ) | ( n15  &  n1692 ) ;
 assign n856 = ( n1118  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1118  &  n1693 ) | ( n1286  &  n1693 ) ;
 assign n857 = ( (~ Pkey_208_)  &  n1694 ) | ( n15  &  n1694 ) ;
 assign n859 = ( n1120  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1120  &  n1695 ) | ( n1286  &  n1695 ) ;
 assign n860 = ( (~ Pkey_200_)  &  n1696 ) | ( n15  &  n1696 ) ;
 assign n862 = ( n1122  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1122  &  n1697 ) | ( n1286  &  n1697 ) ;
 assign n863 = ( (~ Pkey_192_)  &  n1698 ) | ( n15  &  n1698 ) ;
 assign n865 = ( n1124  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1124  &  n1699 ) | ( n1286  &  n1699 ) ;
 assign n866 = ( (~ Pkey_249_)  &  n1700 ) | ( n15  &  n1700 ) ;
 assign n868 = ( n1126  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1126  &  n1701 ) | ( n1286  &  n1701 ) ;
 assign n869 = ( (~ Pkey_241_)  &  n1702 ) | ( n15  &  n1702 ) ;
 assign n871 = ( n1128  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1128  &  n1703 ) | ( n1286  &  n1703 ) ;
 assign n872 = ( (~ Pkey_233_)  &  n1704 ) | ( n15  &  n1704 ) ;
 assign n874 = ( n1130  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1130  &  n1705 ) | ( n1286  &  n1705 ) ;
 assign n875 = ( (~ Pkey_225_)  &  n1706 ) | ( n15  &  n1706 ) ;
 assign n877 = ( n1132  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1132  &  n1707 ) | ( n1286  &  n1707 ) ;
 assign n878 = ( (~ Pkey_217_)  &  n1708 ) | ( n15  &  n1708 ) ;
 assign n880 = ( n1134  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1134  &  n1709 ) | ( n1286  &  n1709 ) ;
 assign n881 = ( (~ Pkey_209_)  &  n1710 ) | ( n15  &  n1710 ) ;
 assign n883 = ( n1136  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1136  &  n1711 ) | ( n1286  &  n1711 ) ;
 assign n884 = ( (~ Pkey_201_)  &  n1712 ) | ( n15  &  n1712 ) ;
 assign n886 = ( n1138  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1138  &  n1713 ) | ( n1286  &  n1713 ) ;
 assign n887 = ( (~ Pkey_193_)  &  n1714 ) | ( n15  &  n1714 ) ;
 assign n889 = ( n1140  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1140  &  n1715 ) | ( n1286  &  n1715 ) ;
 assign n890 = ( (~ Pkey_250_)  &  n1716 ) | ( n15  &  n1716 ) ;
 assign n892 = ( n1142  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1142  &  n1717 ) | ( n1286  &  n1717 ) ;
 assign n893 = ( (~ Pkey_242_)  &  n1718 ) | ( n15  &  n1718 ) ;
 assign n895 = ( n1144  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1144  &  n1719 ) | ( n1286  &  n1719 ) ;
 assign n896 = ( (~ Pkey_234_)  &  n1720 ) | ( n15  &  n1720 ) ;
 assign n898 = ( n1146  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1146  &  n1721 ) | ( n1286  &  n1721 ) ;
 assign n899 = ( (~ Pkey_226_)  &  n1722 ) | ( n15  &  n1722 ) ;
 assign n901 = ( n1148  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1148  &  n1723 ) | ( n1286  &  n1723 ) ;
 assign n902 = ( (~ Pkey_218_)  &  n1724 ) | ( n15  &  n1724 ) ;
 assign n904 = ( n1150  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1150  &  n1725 ) | ( n1286  &  n1725 ) ;
 assign n905 = ( (~ Pkey_210_)  &  n1726 ) | ( n15  &  n1726 ) ;
 assign n907 = ( n1152  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1152  &  n1727 ) | ( n1286  &  n1727 ) ;
 assign n908 = ( (~ Pkey_202_)  &  n1728 ) | ( n15  &  n1728 ) ;
 assign n910 = ( n1154  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1154  &  n1729 ) | ( n1286  &  n1729 ) ;
 assign n911 = ( (~ Pkey_194_)  &  n1730 ) | ( n15  &  n1730 ) ;
 assign n913 = ( n1156  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1156  &  n1731 ) | ( n1286  &  n1731 ) ;
 assign n914 = ( (~ Pkey_251_)  &  n1732 ) | ( n15  &  n1732 ) ;
 assign n916 = ( n1158  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1158  &  n1733 ) | ( n1286  &  n1733 ) ;
 assign n917 = ( (~ Pkey_243_)  &  n1734 ) | ( n15  &  n1734 ) ;
 assign n919 = ( n1160  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1160  &  n1735 ) | ( n1286  &  n1735 ) ;
 assign n920 = ( (~ Pkey_235_)  &  n1736 ) | ( n15  &  n1736 ) ;
 assign n922 = ( n1162  &  (~ n1284) ) | ( (~ n1284)  &  n1286 ) | ( n1162  &  n1737 ) | ( n1286  &  n1737 ) ;
 assign n923 = ( (~ Pkey_227_)  &  n1738 ) | ( n15  &  n1738 ) ;
 assign n925 = ( (~ Pcount_3_) ) | ( n246 ) | ( n1287 ) ;
 assign n924 = ( Pcount_3_ ) | ( Pencrypt_0_ ) | ( n249 ) ;
 assign n929 = ( (~ Pcount_1_)  &  n1966 ) | ( Pcount_1_  &  n1967 ) | ( n1966  &  n1967 ) ;
 assign n928 = ( Pencrypt_0_ ) | ( (~ Pcount_1_) ) ;
 assign n930 = ( Pcount_2_  &  (~ n928) ) | ( Pcount_2_  &  (~ n1967) ) ;
 assign n934 = ( Pstart_0_  &  n15 ) | ( (~ Pcount_0_)  &  n15 ) | ( n15  &  (~ n1289) ) ;
 assign n935 = ( (~ Pcount_2_)  &  (~ Pcount_0_) ) ;
 assign n939 = ( (~ Pencrypt_0_)  &  n924 ) | ( n252  &  n924 ) ;
 assign n938 = ( Pencrypt_0_  &  (~ n246) ) | ( (~ Pencrypt_0_)  &  n935 ) | ( (~ n246)  &  n935 ) ;
 assign n937 = ( (~ Pcount_3_)  &  n939 ) | ( n928  &  n939  &  n938 ) ;
 assign n940 = ( PKSi_118_  &  PKSi_4_ ) | ( (~ PKSi_118_)  &  (~ PKSi_4_) ) ;
 assign n942 = ( PKSi_102_  &  PKSi_23_ ) | ( (~ PKSi_102_)  &  (~ PKSi_23_) ) ;
 assign n944 = ( PKSi_98_  &  PKSi_6_ ) | ( (~ PKSi_98_)  &  (~ PKSi_6_) ) ;
 assign n946 = ( PKSi_119_  &  PKSi_15_ ) | ( (~ PKSi_119_)  &  (~ PKSi_15_) ) ;
 assign n948 = ( PKSi_106_  &  PKSi_5_ ) | ( (~ PKSi_106_)  &  (~ PKSi_5_) ) ;
 assign n950 = ( PKSi_112_  &  PKSi_9_ ) | ( (~ PKSi_112_)  &  (~ PKSi_9_) ) ;
 assign n952 = ( PKSi_19_  &  N_N2986 ) | ( (~ PKSi_19_)  &  (~ N_N2986) ) ;
 assign n954 = ( PKSi_117_  &  PKSi_17_ ) | ( (~ PKSi_117_)  &  (~ PKSi_17_) ) ;
 assign n956 = ( PKSi_99_  &  N_N2853 ) | ( (~ PKSi_99_)  &  (~ N_N2853) ) ;
 assign n958 = ( PKSi_11_  &  N_N2982 ) | ( (~ PKSi_11_)  &  (~ N_N2982) ) ;
 assign n960 = ( PKSi_110_  &  PKSi_2_ ) | ( (~ PKSi_110_)  &  (~ PKSi_2_) ) ;
 assign n962 = ( PKSi_103_  &  PKSi_14_ ) | ( (~ PKSi_103_)  &  (~ PKSi_14_) ) ;
 assign n964 = ( PKSi_96_  &  PKSi_22_ ) | ( (~ PKSi_96_)  &  (~ PKSi_22_) ) ;
 assign n966 = ( PKSi_115_  &  PKSi_0_ ) | ( (~ PKSi_115_)  &  (~ PKSi_0_) ) ;
 assign n968 = ( PKSi_8_  &  N_N2976 ) | ( (~ PKSi_8_)  &  (~ N_N2976) ) ;
 assign n970 = ( PKSi_108_  &  PKSi_18_ ) | ( (~ PKSi_108_)  &  (~ PKSi_18_) ) ;
 assign n972 = ( PKSi_105_  &  PKSi_1_ ) | ( (~ PKSi_105_)  &  (~ PKSi_1_) ) ;
 assign n974 = ( PKSi_114_  &  N_N2843 ) | ( (~ PKSi_114_)  &  (~ N_N2843) ) ;
 assign n976 = ( PKSi_100_  &  PKSi_13_ ) | ( (~ PKSi_100_)  &  (~ PKSi_13_) ) ;
 assign n978 = ( PKSi_107_  &  PKSi_21_ ) | ( (~ PKSi_107_)  &  (~ PKSi_21_) ) ;
 assign n980 = ( PKSi_109_  &  PKSi_10_ ) | ( (~ PKSi_109_)  &  (~ PKSi_10_) ) ;
 assign n982 = ( PKSi_116_  &  N_N2838 ) | ( (~ PKSi_116_)  &  (~ N_N2838) ) ;
 assign n984 = ( PKSi_104_  &  PKSi_12_ ) | ( (~ PKSi_104_)  &  (~ PKSi_12_) ) ;
 assign n986 = ( PKSi_97_  &  PKSi_3_ ) | ( (~ PKSi_97_)  &  (~ PKSi_3_) ) ;
 assign n988 = ( PKSi_113_  &  N_N2834 ) | ( (~ PKSi_113_)  &  (~ N_N2834) ) ;
 assign n990 = ( PKSi_16_  &  N_N2964 ) | ( (~ PKSi_16_)  &  (~ N_N2964) ) ;
 assign n992 = ( PKSi_101_  &  PKSi_20_ ) | ( (~ PKSi_101_)  &  (~ PKSi_20_) ) ;
 assign n994 = ( PKSi_111_  &  PKSi_7_ ) | ( (~ PKSi_111_)  &  (~ PKSi_7_) ) ;
 assign n996 = ( PKSi_142_  &  PKSi_28_ ) | ( (~ PKSi_142_)  &  (~ PKSi_28_) ) ;
 assign n998 = ( PKSi_126_  &  PKSi_47_ ) | ( (~ PKSi_126_)  &  (~ PKSi_47_) ) ;
 assign n1000 = ( PKSi_122_  &  PKSi_30_ ) | ( (~ PKSi_122_)  &  (~ PKSi_30_) ) ;
 assign n1002 = ( wire282  &  PKSi_39_ ) | ( (~ wire282)  &  (~ PKSi_39_) ) ;
 assign n1004 = ( PKSi_130_  &  PKSi_29_ ) | ( (~ PKSi_130_)  &  (~ PKSi_29_) ) ;
 assign n1006 = ( PKSi_136_  &  PKSi_33_ ) | ( (~ PKSi_136_)  &  (~ PKSi_33_) ) ;
 assign n1008 = ( PKSi_43_  &  N_N2954 ) | ( (~ PKSi_43_)  &  (~ N_N2954) ) ;
 assign n1010 = ( PKSi_141_  &  PKSi_41_ ) | ( (~ PKSi_141_)  &  (~ PKSi_41_) ) ;
 assign n1012 = ( PKSi_123_  &  N_N2821 ) | ( (~ PKSi_123_)  &  (~ N_N2821) ) ;
 assign n1014 = ( PKSi_35_  &  N_N2950 ) | ( (~ PKSi_35_)  &  (~ N_N2950) ) ;
 assign n1016 = ( PKSi_134_  &  PKSi_26_ ) | ( (~ PKSi_134_)  &  (~ PKSi_26_) ) ;
 assign n1018 = ( PKSi_127_  &  PKSi_38_ ) | ( (~ PKSi_127_)  &  (~ PKSi_38_) ) ;
 assign n1020 = ( PKSi_120_  &  PKSi_46_ ) | ( (~ PKSi_120_)  &  (~ PKSi_46_) ) ;
 assign n1022 = ( PKSi_24_  &  N_N2945 ) | ( (~ PKSi_24_)  &  (~ N_N2945) ) ;
 assign n1024 = ( PKSi_32_  &  N_N2943 ) | ( (~ PKSi_32_)  &  (~ N_N2943) ) ;
 assign n1026 = ( PKSi_132_  &  PKSi_42_ ) | ( (~ PKSi_132_)  &  (~ PKSi_42_) ) ;
 assign n1028 = ( PKSi_129_  &  PKSi_25_ ) | ( (~ PKSi_129_)  &  (~ PKSi_25_) ) ;
 assign n1030 = ( PKSi_138_  &  N_N2811 ) | ( (~ PKSi_138_)  &  (~ N_N2811) ) ;
 assign n1032 = ( PKSi_124_  &  PKSi_37_ ) | ( (~ PKSi_124_)  &  (~ PKSi_37_) ) ;
 assign n1034 = ( PKSi_131_  &  PKSi_45_ ) | ( (~ PKSi_131_)  &  (~ PKSi_45_) ) ;
 assign n1036 = ( PKSi_133_  &  PKSi_34_ ) | ( (~ PKSi_133_)  &  (~ PKSi_34_) ) ;
 assign n1038 = ( PKSi_140_  &  N_N2806 ) | ( (~ PKSi_140_)  &  (~ N_N2806) ) ;
 assign n1040 = ( PKSi_128_  &  PKSi_36_ ) | ( (~ PKSi_128_)  &  (~ PKSi_36_) ) ;
 assign n1042 = ( PKSi_121_  &  PKSi_27_ ) | ( (~ PKSi_121_)  &  (~ PKSi_27_) ) ;
 assign n1044 = ( PKSi_137_  &  N_N2802 ) | ( (~ PKSi_137_)  &  (~ N_N2802) ) ;
 assign n1046 = ( PKSi_40_  &  N_N2931 ) | ( (~ PKSi_40_)  &  (~ N_N2931) ) ;
 assign n1048 = ( PKSi_125_  &  PKSi_44_ ) | ( (~ PKSi_125_)  &  (~ PKSi_44_) ) ;
 assign n1050 = ( PKSi_135_  &  PKSi_31_ ) | ( (~ PKSi_135_)  &  (~ PKSi_31_) ) ;
 assign n1052 = ( PKSi_166_  &  PKSi_52_ ) | ( (~ PKSi_166_)  &  (~ PKSi_52_) ) ;
 assign n1054 = ( PKSi_150_  &  PKSi_71_ ) | ( (~ PKSi_150_)  &  (~ PKSi_71_) ) ;
 assign n1056 = ( PKSi_146_  &  PKSi_54_ ) | ( (~ PKSi_146_)  &  (~ PKSi_54_) ) ;
 assign n1058 = ( PKSi_167_  &  PKSi_63_ ) | ( (~ PKSi_167_)  &  (~ PKSi_63_) ) ;
 assign n1060 = ( PKSi_154_  &  PKSi_53_ ) | ( (~ PKSi_154_)  &  (~ PKSi_53_) ) ;
 assign n1062 = ( PKSi_160_  &  PKSi_57_ ) | ( (~ PKSi_160_)  &  (~ PKSi_57_) ) ;
 assign n1064 = ( PKSi_67_  &  N_N2921 ) | ( (~ PKSi_67_)  &  (~ N_N2921) ) ;
 assign n1066 = ( PKSi_165_  &  PKSi_65_ ) | ( (~ PKSi_165_)  &  (~ PKSi_65_) ) ;
 assign n1068 = ( PKSi_147_  &  N_N2789 ) | ( (~ PKSi_147_)  &  (~ N_N2789) ) ;
 assign n1070 = ( PKSi_59_  &  N_N2917 ) | ( (~ PKSi_59_)  &  (~ N_N2917) ) ;
 assign n1072 = ( PKSi_158_  &  PKSi_50_ ) | ( (~ PKSi_158_)  &  (~ PKSi_50_) ) ;
 assign n1074 = ( PKSi_151_  &  PKSi_62_ ) | ( (~ PKSi_151_)  &  (~ PKSi_62_) ) ;
 assign n1076 = ( PKSi_144_  &  PKSi_70_ ) | ( (~ PKSi_144_)  &  (~ PKSi_70_) ) ;
 assign n1078 = ( PKSi_163_  &  PKSi_48_ ) | ( (~ PKSi_163_)  &  (~ PKSi_48_) ) ;
 assign n1080 = ( PKSi_153_  &  PKSi_56_ ) | ( (~ PKSi_153_)  &  (~ PKSi_56_) ) ;
 assign n1082 = ( PKSi_156_  &  PKSi_66_ ) | ( (~ PKSi_156_)  &  (~ PKSi_66_) ) ;
 assign n1084 = ( PKSi_49_  &  N_N2909 ) | ( (~ PKSi_49_)  &  (~ N_N2909) ) ;
 assign n1086 = ( PKSi_162_  &  N_N2779 ) | ( (~ PKSi_162_)  &  (~ N_N2779) ) ;
 assign n1088 = ( PKSi_148_  &  PKSi_61_ ) | ( (~ PKSi_148_)  &  (~ PKSi_61_) ) ;
 assign n1090 = ( PKSi_155_  &  PKSi_69_ ) | ( (~ PKSi_155_)  &  (~ PKSi_69_) ) ;
 assign n1092 = ( PKSi_157_  &  PKSi_58_ ) | ( (~ PKSi_157_)  &  (~ PKSi_58_) ) ;
 assign n1094 = ( PKSi_164_  &  N_N2774 ) | ( (~ PKSi_164_)  &  (~ N_N2774) ) ;
 assign n1096 = ( PKSi_152_  &  PKSi_60_ ) | ( (~ PKSi_152_)  &  (~ PKSi_60_) ) ;
 assign n1098 = ( PKSi_145_  &  PKSi_51_ ) | ( (~ PKSi_145_)  &  (~ PKSi_51_) ) ;
 assign n1100 = ( PKSi_161_  &  N_N2770 ) | ( (~ PKSi_161_)  &  (~ N_N2770) ) ;
 assign n1102 = ( PKSi_64_  &  N_N2899 ) | ( (~ PKSi_64_)  &  (~ N_N2899) ) ;
 assign n1104 = ( PKSi_149_  &  PKSi_68_ ) | ( (~ PKSi_149_)  &  (~ PKSi_68_) ) ;
 assign n1106 = ( PKSi_159_  &  PKSi_55_ ) | ( (~ PKSi_159_)  &  (~ PKSi_55_) ) ;
 assign n1108 = ( PKSi_190_  &  PKSi_76_ ) | ( (~ PKSi_190_)  &  (~ PKSi_76_) ) ;
 assign n1110 = ( PKSi_174_  &  PKSi_95_ ) | ( (~ PKSi_174_)  &  (~ PKSi_95_) ) ;
 assign n1112 = ( PKSi_170_  &  PKSi_78_ ) | ( (~ PKSi_170_)  &  (~ PKSi_78_) ) ;
 assign n1114 = ( wire234  &  PKSi_87_ ) | ( (~ wire234)  &  (~ PKSi_87_) ) ;
 assign n1116 = ( PKSi_178_  &  PKSi_77_ ) | ( (~ PKSi_178_)  &  (~ PKSi_77_) ) ;
 assign n1118 = ( PKSi_184_  &  PKSi_81_ ) | ( (~ PKSi_184_)  &  (~ PKSi_81_) ) ;
 assign n1120 = ( PKSi_91_  &  N_N2889 ) | ( (~ PKSi_91_)  &  (~ N_N2889) ) ;
 assign n1122 = ( PKSi_189_  &  PKSi_89_ ) | ( (~ PKSi_189_)  &  (~ PKSi_89_) ) ;
 assign n1124 = ( PKSi_171_  &  N_N2757 ) | ( (~ PKSi_171_)  &  (~ N_N2757) ) ;
 assign n1126 = ( PKSi_83_  &  N_N2885 ) | ( (~ PKSi_83_)  &  (~ N_N2885) ) ;
 assign n1128 = ( PKSi_182_  &  PKSi_74_ ) | ( (~ PKSi_182_)  &  (~ PKSi_74_) ) ;
 assign n1130 = ( PKSi_175_  &  PKSi_86_ ) | ( (~ PKSi_175_)  &  (~ PKSi_86_) ) ;
 assign n1132 = ( PKSi_94_  &  N_N2881 ) | ( (~ PKSi_94_)  &  (~ N_N2881) ) ;
 assign n1134 = ( PKSi_72_  &  N_N2879 ) | ( (~ PKSi_72_)  &  (~ N_N2879) ) ;
 assign n1136 = ( PKSi_80_  &  N_N2877 ) | ( (~ PKSi_80_)  &  (~ N_N2877) ) ;
 assign n1138 = ( PKSi_180_  &  N_N2749 ) | ( (~ PKSi_180_)  &  (~ N_N2749) ) ;
 assign n1140 = ( PKSi_177_  &  PKSi_73_ ) | ( (~ PKSi_177_)  &  (~ PKSi_73_) ) ;
 assign n1142 = ( PKSi_186_  &  N_N2746 ) | ( (~ PKSi_186_)  &  (~ N_N2746) ) ;
 assign n1144 = ( PKSi_172_  &  PKSi_85_ ) | ( (~ PKSi_172_)  &  (~ PKSi_85_) ) ;
 assign n1146 = ( PKSi_179_  &  PKSi_93_ ) | ( (~ PKSi_179_)  &  (~ PKSi_93_) ) ;
 assign n1148 = ( wire253  &  PKSi_82_ ) | ( (~ wire253)  &  (~ PKSi_82_) ) ;
 assign n1150 = ( PKSi_188_  &  N_N2741 ) | ( (~ PKSi_188_)  &  (~ N_N2741) ) ;
 assign n1152 = ( PKSi_176_  &  PKSi_84_ ) | ( (~ PKSi_176_)  &  (~ PKSi_84_) ) ;
 assign n1154 = ( PKSi_169_  &  PKSi_75_ ) | ( (~ PKSi_169_)  &  (~ PKSi_75_) ) ;
 assign n1156 = ( PKSi_185_  &  N_N2737 ) | ( (~ PKSi_185_)  &  (~ N_N2737) ) ;
 assign n1158 = ( wire333  &  N_N2865 ) | ( (~ wire333)  &  (~ N_N2865) ) ;
 assign n1160 = ( PKSi_173_  &  PKSi_92_ ) | ( (~ PKSi_173_)  &  (~ PKSi_92_) ) ;
 assign n1162 = ( PKSi_183_  &  PKSi_79_ ) | ( (~ PKSi_183_)  &  (~ PKSi_79_) ) ;
 assign n1167 = ( Pencrypt_0_  &  (~ n250) ) ;
 assign n1166 = ( Pstart_0_ ) | ( n1167 ) ;
 assign n1170 = ( Pstart_0_ ) | ( (~ n1167) ) ;
 assign n1285 = ( (~ Pencrypt_0_) ) | ( (~ n250) ) ;
 assign n1284 = ( (~ Pstart_0_)  &  n1285 ) ;
 assign n1286 = ( Pstart_0_ ) | ( n1285 ) ;
 assign n1287 = ( Pstart_0_ ) | ( (~ Pencrypt_0_) ) ;
 assign n1289 = ( (~ Pcount_1_)  &  n1968 ) | ( Pencrypt_0_  &  (~ Pcount_2_)  &  n1968 ) ;
 assign n1290 = ( n940 ) | ( n1170 ) ;
 assign n1291 = ( n11  &  (~ n1741) ) | ( n11  &  n1740 ) | ( (~ n1741)  &  (~ n1740) ) ;
 assign n1292 = ( n942 ) | ( n1170 ) ;
 assign n1293 = ( n11  &  (~ n1741) ) | ( n11  &  n1744 ) | ( (~ n1741)  &  (~ n1744) ) ;
 assign n1294 = ( n944 ) | ( n1170 ) ;
 assign n1295 = ( n11  &  (~ n1741) ) | ( n11  &  n1746 ) | ( (~ n1741)  &  (~ n1746) ) ;
 assign n1296 = ( n946 ) | ( n1170 ) ;
 assign n1297 = ( n11  &  (~ n1741) ) | ( n11  &  n1748 ) | ( (~ n1741)  &  (~ n1748) ) ;
 assign n1298 = ( n948 ) | ( n1170 ) ;
 assign n1299 = ( n11  &  (~ n1741) ) | ( n11  &  n1750 ) | ( (~ n1741)  &  (~ n1750) ) ;
 assign n1300 = ( n950 ) | ( n1170 ) ;
 assign n1301 = ( n11  &  (~ n1741) ) | ( n11  &  n1752 ) | ( (~ n1741)  &  (~ n1752) ) ;
 assign n1302 = ( n952 ) | ( n1170 ) ;
 assign n1303 = ( n11  &  (~ n1741) ) | ( n11  &  n1754 ) | ( (~ n1741)  &  (~ n1754) ) ;
 assign n1304 = ( n954 ) | ( n1170 ) ;
 assign n1305 = ( n11  &  (~ n1741) ) | ( n11  &  n1756 ) | ( (~ n1741)  &  (~ n1756) ) ;
 assign n1306 = ( n956 ) | ( n1170 ) ;
 assign n1307 = ( n11  &  (~ n1741) ) | ( n11  &  n1758 ) | ( (~ n1741)  &  (~ n1758) ) ;
 assign n1308 = ( n958 ) | ( n1170 ) ;
 assign n1309 = ( n11  &  (~ n1741) ) | ( n11  &  n1760 ) | ( (~ n1741)  &  (~ n1760) ) ;
 assign n1310 = ( n960 ) | ( n1170 ) ;
 assign n1311 = ( n11  &  (~ n1741) ) | ( n11  &  n1762 ) | ( (~ n1741)  &  (~ n1762) ) ;
 assign n1312 = ( n962 ) | ( n1170 ) ;
 assign n1313 = ( n11  &  (~ n1741) ) | ( n11  &  n1764 ) | ( (~ n1741)  &  (~ n1764) ) ;
 assign n1314 = ( n964 ) | ( n1170 ) ;
 assign n1315 = ( n11  &  (~ n1741) ) | ( n11  &  n1766 ) | ( (~ n1741)  &  (~ n1766) ) ;
 assign n1316 = ( n966 ) | ( n1170 ) ;
 assign n1317 = ( n11  &  (~ n1741) ) | ( n11  &  n1768 ) | ( (~ n1741)  &  (~ n1768) ) ;
 assign n1318 = ( n968 ) | ( n1170 ) ;
 assign n1319 = ( n11  &  (~ n1741) ) | ( n11  &  n1770 ) | ( (~ n1741)  &  (~ n1770) ) ;
 assign n1320 = ( n970 ) | ( n1170 ) ;
 assign n1321 = ( n11  &  (~ n1741) ) | ( n11  &  n1772 ) | ( (~ n1741)  &  (~ n1772) ) ;
 assign n1322 = ( n972 ) | ( n1170 ) ;
 assign n1323 = ( n11  &  (~ n1741) ) | ( n11  &  n1774 ) | ( (~ n1741)  &  (~ n1774) ) ;
 assign n1324 = ( n974 ) | ( n1170 ) ;
 assign n1325 = ( n11  &  (~ n1741) ) | ( n11  &  n1776 ) | ( (~ n1741)  &  (~ n1776) ) ;
 assign n1326 = ( n976 ) | ( n1170 ) ;
 assign n1327 = ( n11  &  (~ n1741) ) | ( n11  &  n1778 ) | ( (~ n1741)  &  (~ n1778) ) ;
 assign n1328 = ( n978 ) | ( n1170 ) ;
 assign n1329 = ( n11  &  (~ n1741) ) | ( n11  &  n1780 ) | ( (~ n1741)  &  (~ n1780) ) ;
 assign n1330 = ( n980 ) | ( n1170 ) ;
 assign n1331 = ( n11  &  (~ n1741) ) | ( n11  &  n1782 ) | ( (~ n1741)  &  (~ n1782) ) ;
 assign n1332 = ( n982 ) | ( n1170 ) ;
 assign n1333 = ( n11  &  (~ n1741) ) | ( n11  &  n1784 ) | ( (~ n1741)  &  (~ n1784) ) ;
 assign n1334 = ( n984 ) | ( n1170 ) ;
 assign n1335 = ( n11  &  (~ n1741) ) | ( n11  &  n1786 ) | ( (~ n1741)  &  (~ n1786) ) ;
 assign n1336 = ( n986 ) | ( n1170 ) ;
 assign n1337 = ( n11  &  (~ n1741) ) | ( n11  &  n1788 ) | ( (~ n1741)  &  (~ n1788) ) ;
 assign n1338 = ( n988 ) | ( n1170 ) ;
 assign n1339 = ( n11  &  (~ n1741) ) | ( n11  &  n1790 ) | ( (~ n1741)  &  (~ n1790) ) ;
 assign n1340 = ( n990 ) | ( n1170 ) ;
 assign n1341 = ( n11  &  (~ n1741) ) | ( n11  &  n1792 ) | ( (~ n1741)  &  (~ n1792) ) ;
 assign n1342 = ( n992 ) | ( n1170 ) ;
 assign n1343 = ( n11  &  (~ n1741) ) | ( n11  &  n1794 ) | ( (~ n1741)  &  (~ n1794) ) ;
 assign n1344 = ( n994 ) | ( n1170 ) ;
 assign n1345 = ( n11  &  (~ n1741) ) | ( n11  &  n1796 ) | ( (~ n1741)  &  (~ n1796) ) ;
 assign n1346 = ( n996 ) | ( n1170 ) ;
 assign n1347 = ( n11  &  (~ n1741) ) | ( n11  &  n1798 ) | ( (~ n1741)  &  (~ n1798) ) ;
 assign n1348 = ( n998 ) | ( n1170 ) ;
 assign n1349 = ( n11  &  (~ n1741) ) | ( n11  &  n1800 ) | ( (~ n1741)  &  (~ n1800) ) ;
 assign n1350 = ( n1000 ) | ( n1170 ) ;
 assign n1351 = ( n11  &  (~ n1741) ) | ( n11  &  n1802 ) | ( (~ n1741)  &  (~ n1802) ) ;
 assign n1352 = ( n1002 ) | ( n1170 ) ;
 assign n1353 = ( n11  &  (~ n1741) ) | ( n11  &  n1804 ) | ( (~ n1741)  &  (~ n1804) ) ;
 assign n1354 = ( n1004 ) | ( n1170 ) ;
 assign n1355 = ( n11  &  (~ n1741) ) | ( n11  &  n1806 ) | ( (~ n1741)  &  (~ n1806) ) ;
 assign n1356 = ( n1006 ) | ( n1170 ) ;
 assign n1357 = ( n11  &  (~ n1741) ) | ( n11  &  n1808 ) | ( (~ n1741)  &  (~ n1808) ) ;
 assign n1358 = ( n1008 ) | ( n1170 ) ;
 assign n1359 = ( n11  &  (~ n1741) ) | ( n11  &  n1810 ) | ( (~ n1741)  &  (~ n1810) ) ;
 assign n1360 = ( n1010 ) | ( n1170 ) ;
 assign n1361 = ( n11  &  (~ n1741) ) | ( n11  &  n1812 ) | ( (~ n1741)  &  (~ n1812) ) ;
 assign n1362 = ( n1012 ) | ( n1170 ) ;
 assign n1363 = ( n11  &  (~ n1741) ) | ( n11  &  n1814 ) | ( (~ n1741)  &  (~ n1814) ) ;
 assign n1364 = ( n1014 ) | ( n1170 ) ;
 assign n1365 = ( n11  &  (~ n1741) ) | ( n11  &  n1816 ) | ( (~ n1741)  &  (~ n1816) ) ;
 assign n1366 = ( n1016 ) | ( n1170 ) ;
 assign n1367 = ( n11  &  (~ n1741) ) | ( n11  &  n1818 ) | ( (~ n1741)  &  (~ n1818) ) ;
 assign n1368 = ( n1018 ) | ( n1170 ) ;
 assign n1369 = ( n11  &  (~ n1741) ) | ( n11  &  n1820 ) | ( (~ n1741)  &  (~ n1820) ) ;
 assign n1370 = ( n1020 ) | ( n1170 ) ;
 assign n1371 = ( n11  &  (~ n1741) ) | ( n11  &  n1822 ) | ( (~ n1741)  &  (~ n1822) ) ;
 assign n1372 = ( n1022 ) | ( n1170 ) ;
 assign n1373 = ( n11  &  (~ n1741) ) | ( n11  &  n1824 ) | ( (~ n1741)  &  (~ n1824) ) ;
 assign n1374 = ( n1024 ) | ( n1170 ) ;
 assign n1375 = ( n11  &  (~ n1741) ) | ( n11  &  n1826 ) | ( (~ n1741)  &  (~ n1826) ) ;
 assign n1376 = ( n1026 ) | ( n1170 ) ;
 assign n1377 = ( n11  &  (~ n1741) ) | ( n11  &  n1828 ) | ( (~ n1741)  &  (~ n1828) ) ;
 assign n1378 = ( n1028 ) | ( n1170 ) ;
 assign n1379 = ( n11  &  (~ n1741) ) | ( n11  &  n1830 ) | ( (~ n1741)  &  (~ n1830) ) ;
 assign n1380 = ( n1030 ) | ( n1170 ) ;
 assign n1381 = ( n11  &  (~ n1741) ) | ( n11  &  n1832 ) | ( (~ n1741)  &  (~ n1832) ) ;
 assign n1382 = ( n1032 ) | ( n1170 ) ;
 assign n1383 = ( n11  &  (~ n1741) ) | ( n11  &  n1834 ) | ( (~ n1741)  &  (~ n1834) ) ;
 assign n1384 = ( n1034 ) | ( n1170 ) ;
 assign n1385 = ( n11  &  (~ n1741) ) | ( n11  &  n1836 ) | ( (~ n1741)  &  (~ n1836) ) ;
 assign n1386 = ( n1036 ) | ( n1170 ) ;
 assign n1387 = ( n11  &  (~ n1741) ) | ( n11  &  n1838 ) | ( (~ n1741)  &  (~ n1838) ) ;
 assign n1388 = ( n1038 ) | ( n1170 ) ;
 assign n1389 = ( n11  &  (~ n1741) ) | ( n11  &  n1840 ) | ( (~ n1741)  &  (~ n1840) ) ;
 assign n1390 = ( n1040 ) | ( n1170 ) ;
 assign n1391 = ( n11  &  (~ n1741) ) | ( n11  &  n1842 ) | ( (~ n1741)  &  (~ n1842) ) ;
 assign n1392 = ( n1042 ) | ( n1170 ) ;
 assign n1393 = ( n11  &  (~ n1741) ) | ( n11  &  n1844 ) | ( (~ n1741)  &  (~ n1844) ) ;
 assign n1394 = ( n1044 ) | ( n1170 ) ;
 assign n1395 = ( n11  &  (~ n1741) ) | ( n11  &  n1846 ) | ( (~ n1741)  &  (~ n1846) ) ;
 assign n1396 = ( n1046 ) | ( n1170 ) ;
 assign n1397 = ( n11  &  (~ n1741) ) | ( n11  &  n1848 ) | ( (~ n1741)  &  (~ n1848) ) ;
 assign n1398 = ( n1048 ) | ( n1170 ) ;
 assign n1399 = ( n11  &  (~ n1741) ) | ( n11  &  n1850 ) | ( (~ n1741)  &  (~ n1850) ) ;
 assign n1400 = ( n1050 ) | ( n1170 ) ;
 assign n1401 = ( n11  &  (~ n1741) ) | ( n11  &  n1852 ) | ( (~ n1741)  &  (~ n1852) ) ;
 assign n1402 = ( n1052 ) | ( n1170 ) ;
 assign n1403 = ( n11  &  (~ n1741) ) | ( n11  &  n1854 ) | ( (~ n1741)  &  (~ n1854) ) ;
 assign n1404 = ( n1054 ) | ( n1170 ) ;
 assign n1405 = ( n11  &  (~ n1741) ) | ( n11  &  n1856 ) | ( (~ n1741)  &  (~ n1856) ) ;
 assign n1406 = ( n1056 ) | ( n1170 ) ;
 assign n1407 = ( n11  &  (~ n1741) ) | ( n11  &  n1858 ) | ( (~ n1741)  &  (~ n1858) ) ;
 assign n1408 = ( n1058 ) | ( n1170 ) ;
 assign n1409 = ( n11  &  (~ n1741) ) | ( n11  &  n1860 ) | ( (~ n1741)  &  (~ n1860) ) ;
 assign n1410 = ( n1060 ) | ( n1170 ) ;
 assign n1411 = ( n11  &  (~ n1741) ) | ( n11  &  n1862 ) | ( (~ n1741)  &  (~ n1862) ) ;
 assign n1412 = ( n1062 ) | ( n1170 ) ;
 assign n1413 = ( n11  &  (~ n1741) ) | ( n11  &  n1864 ) | ( (~ n1741)  &  (~ n1864) ) ;
 assign n1414 = ( n1064 ) | ( n1170 ) ;
 assign n1415 = ( n11  &  (~ n1741) ) | ( n11  &  n1866 ) | ( (~ n1741)  &  (~ n1866) ) ;
 assign n1416 = ( n1066 ) | ( n1170 ) ;
 assign n1417 = ( n11  &  (~ n1741) ) | ( n11  &  n1868 ) | ( (~ n1741)  &  (~ n1868) ) ;
 assign n1418 = ( n1068 ) | ( n1170 ) ;
 assign n1419 = ( n11  &  (~ n1741) ) | ( n11  &  n1870 ) | ( (~ n1741)  &  (~ n1870) ) ;
 assign n1420 = ( n1070 ) | ( n1170 ) ;
 assign n1421 = ( n11  &  (~ n1741) ) | ( n11  &  n1872 ) | ( (~ n1741)  &  (~ n1872) ) ;
 assign n1422 = ( n1072 ) | ( n1170 ) ;
 assign n1423 = ( n11  &  (~ n1741) ) | ( n11  &  n1874 ) | ( (~ n1741)  &  (~ n1874) ) ;
 assign n1424 = ( n1074 ) | ( n1170 ) ;
 assign n1425 = ( n11  &  (~ n1741) ) | ( n11  &  n1876 ) | ( (~ n1741)  &  (~ n1876) ) ;
 assign n1426 = ( n1076 ) | ( n1170 ) ;
 assign n1427 = ( n11  &  (~ n1741) ) | ( n11  &  n1878 ) | ( (~ n1741)  &  (~ n1878) ) ;
 assign n1428 = ( n1078 ) | ( n1170 ) ;
 assign n1429 = ( n11  &  (~ n1741) ) | ( n11  &  n1880 ) | ( (~ n1741)  &  (~ n1880) ) ;
 assign n1430 = ( n1080 ) | ( n1170 ) ;
 assign n1431 = ( n11  &  (~ n1741) ) | ( n11  &  n1882 ) | ( (~ n1741)  &  (~ n1882) ) ;
 assign n1432 = ( n1082 ) | ( n1170 ) ;
 assign n1433 = ( n11  &  (~ n1741) ) | ( n11  &  n1884 ) | ( (~ n1741)  &  (~ n1884) ) ;
 assign n1434 = ( n1084 ) | ( n1170 ) ;
 assign n1435 = ( n11  &  (~ n1741) ) | ( n11  &  n1886 ) | ( (~ n1741)  &  (~ n1886) ) ;
 assign n1436 = ( n1086 ) | ( n1170 ) ;
 assign n1437 = ( n11  &  (~ n1741) ) | ( n11  &  n1888 ) | ( (~ n1741)  &  (~ n1888) ) ;
 assign n1438 = ( n1088 ) | ( n1170 ) ;
 assign n1439 = ( n11  &  (~ n1741) ) | ( n11  &  n1890 ) | ( (~ n1741)  &  (~ n1890) ) ;
 assign n1440 = ( n1090 ) | ( n1170 ) ;
 assign n1441 = ( n11  &  (~ n1741) ) | ( n11  &  n1892 ) | ( (~ n1741)  &  (~ n1892) ) ;
 assign n1442 = ( n1092 ) | ( n1170 ) ;
 assign n1443 = ( n11  &  (~ n1741) ) | ( n11  &  n1894 ) | ( (~ n1741)  &  (~ n1894) ) ;
 assign n1444 = ( n1094 ) | ( n1170 ) ;
 assign n1445 = ( n11  &  (~ n1741) ) | ( n11  &  n1896 ) | ( (~ n1741)  &  (~ n1896) ) ;
 assign n1446 = ( n1096 ) | ( n1170 ) ;
 assign n1447 = ( n11  &  (~ n1741) ) | ( n11  &  n1898 ) | ( (~ n1741)  &  (~ n1898) ) ;
 assign n1448 = ( n1098 ) | ( n1170 ) ;
 assign n1449 = ( n11  &  (~ n1741) ) | ( n11  &  n1900 ) | ( (~ n1741)  &  (~ n1900) ) ;
 assign n1450 = ( n1100 ) | ( n1170 ) ;
 assign n1451 = ( n11  &  (~ n1741) ) | ( n11  &  n1902 ) | ( (~ n1741)  &  (~ n1902) ) ;
 assign n1452 = ( n1102 ) | ( n1170 ) ;
 assign n1453 = ( n11  &  (~ n1741) ) | ( n11  &  n1904 ) | ( (~ n1741)  &  (~ n1904) ) ;
 assign n1454 = ( n1104 ) | ( n1170 ) ;
 assign n1455 = ( n11  &  (~ n1741) ) | ( n11  &  n1906 ) | ( (~ n1741)  &  (~ n1906) ) ;
 assign n1456 = ( n1106 ) | ( n1170 ) ;
 assign n1457 = ( n11  &  (~ n1741) ) | ( n11  &  n1908 ) | ( (~ n1741)  &  (~ n1908) ) ;
 assign n1458 = ( n1108 ) | ( n1170 ) ;
 assign n1459 = ( n11  &  (~ n1741) ) | ( n11  &  n1910 ) | ( (~ n1741)  &  (~ n1910) ) ;
 assign n1460 = ( n1110 ) | ( n1170 ) ;
 assign n1461 = ( n11  &  (~ n1741) ) | ( n11  &  n1912 ) | ( (~ n1741)  &  (~ n1912) ) ;
 assign n1462 = ( n1112 ) | ( n1170 ) ;
 assign n1463 = ( n11  &  (~ n1741) ) | ( n11  &  n1914 ) | ( (~ n1741)  &  (~ n1914) ) ;
 assign n1464 = ( n1114 ) | ( n1170 ) ;
 assign n1465 = ( n11  &  (~ n1741) ) | ( n11  &  n1916 ) | ( (~ n1741)  &  (~ n1916) ) ;
 assign n1466 = ( n1116 ) | ( n1170 ) ;
 assign n1467 = ( n11  &  (~ n1741) ) | ( n11  &  n1918 ) | ( (~ n1741)  &  (~ n1918) ) ;
 assign n1468 = ( n1118 ) | ( n1170 ) ;
 assign n1469 = ( n11  &  (~ n1741) ) | ( n11  &  n1920 ) | ( (~ n1741)  &  (~ n1920) ) ;
 assign n1470 = ( n1120 ) | ( n1170 ) ;
 assign n1471 = ( n11  &  (~ n1741) ) | ( n11  &  n1922 ) | ( (~ n1741)  &  (~ n1922) ) ;
 assign n1472 = ( n1122 ) | ( n1170 ) ;
 assign n1473 = ( n11  &  (~ n1741) ) | ( n11  &  n1924 ) | ( (~ n1741)  &  (~ n1924) ) ;
 assign n1474 = ( n1124 ) | ( n1170 ) ;
 assign n1475 = ( n11  &  (~ n1741) ) | ( n11  &  n1926 ) | ( (~ n1741)  &  (~ n1926) ) ;
 assign n1476 = ( n1126 ) | ( n1170 ) ;
 assign n1477 = ( n11  &  (~ n1741) ) | ( n11  &  n1928 ) | ( (~ n1741)  &  (~ n1928) ) ;
 assign n1478 = ( n1128 ) | ( n1170 ) ;
 assign n1479 = ( n11  &  (~ n1741) ) | ( n11  &  n1930 ) | ( (~ n1741)  &  (~ n1930) ) ;
 assign n1480 = ( n1130 ) | ( n1170 ) ;
 assign n1481 = ( n11  &  (~ n1741) ) | ( n11  &  n1932 ) | ( (~ n1741)  &  (~ n1932) ) ;
 assign n1482 = ( n1132 ) | ( n1170 ) ;
 assign n1483 = ( n11  &  (~ n1741) ) | ( n11  &  n1934 ) | ( (~ n1741)  &  (~ n1934) ) ;
 assign n1484 = ( n1134 ) | ( n1170 ) ;
 assign n1485 = ( n11  &  (~ n1741) ) | ( n11  &  n1936 ) | ( (~ n1741)  &  (~ n1936) ) ;
 assign n1486 = ( n1136 ) | ( n1170 ) ;
 assign n1487 = ( n11  &  (~ n1741) ) | ( n11  &  n1938 ) | ( (~ n1741)  &  (~ n1938) ) ;
 assign n1488 = ( n1138 ) | ( n1170 ) ;
 assign n1489 = ( n11  &  (~ n1741) ) | ( n11  &  n1940 ) | ( (~ n1741)  &  (~ n1940) ) ;
 assign n1490 = ( n1140 ) | ( n1170 ) ;
 assign n1491 = ( n11  &  (~ n1741) ) | ( n11  &  n1942 ) | ( (~ n1741)  &  (~ n1942) ) ;
 assign n1492 = ( n1142 ) | ( n1170 ) ;
 assign n1493 = ( n11  &  (~ n1741) ) | ( n11  &  n1944 ) | ( (~ n1741)  &  (~ n1944) ) ;
 assign n1494 = ( n1144 ) | ( n1170 ) ;
 assign n1495 = ( n11  &  (~ n1741) ) | ( n11  &  n1946 ) | ( (~ n1741)  &  (~ n1946) ) ;
 assign n1496 = ( n1146 ) | ( n1170 ) ;
 assign n1497 = ( n11  &  (~ n1741) ) | ( n11  &  n1948 ) | ( (~ n1741)  &  (~ n1948) ) ;
 assign n1498 = ( n1148 ) | ( n1170 ) ;
 assign n1499 = ( n11  &  (~ n1741) ) | ( n11  &  n1950 ) | ( (~ n1741)  &  (~ n1950) ) ;
 assign n1500 = ( n1150 ) | ( n1170 ) ;
 assign n1501 = ( n11  &  (~ n1741) ) | ( n11  &  n1952 ) | ( (~ n1741)  &  (~ n1952) ) ;
 assign n1502 = ( n1152 ) | ( n1170 ) ;
 assign n1503 = ( n11  &  (~ n1741) ) | ( n11  &  n1954 ) | ( (~ n1741)  &  (~ n1954) ) ;
 assign n1504 = ( n1154 ) | ( n1170 ) ;
 assign n1505 = ( n11  &  (~ n1741) ) | ( n11  &  n1956 ) | ( (~ n1741)  &  (~ n1956) ) ;
 assign n1506 = ( n1156 ) | ( n1170 ) ;
 assign n1507 = ( n11  &  (~ n1741) ) | ( n11  &  n1958 ) | ( (~ n1741)  &  (~ n1958) ) ;
 assign n1508 = ( n1158 ) | ( n1170 ) ;
 assign n1509 = ( n11  &  (~ n1741) ) | ( n11  &  n1960 ) | ( (~ n1741)  &  (~ n1960) ) ;
 assign n1510 = ( n1160 ) | ( n1170 ) ;
 assign n1511 = ( n11  &  (~ n1741) ) | ( n11  &  n1962 ) | ( (~ n1741)  &  (~ n1962) ) ;
 assign n1512 = ( n1162 ) | ( n1170 ) ;
 assign n1513 = ( n11  &  (~ n1741) ) | ( n11  &  n1964 ) | ( (~ n1741)  &  (~ n1964) ) ;
 assign n1514 = ( (~ PKSi_118_) ) | ( (~ PKSi_4_) ) ;
 assign n1516 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1740 ) | ( n11  &  (~ n1740) ) ;
 assign n1517 = ( (~ PKSi_102_) ) | ( (~ PKSi_23_) ) ;
 assign n1518 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1744 ) | ( n11  &  (~ n1744) ) ;
 assign n1519 = ( (~ PKSi_98_) ) | ( (~ PKSi_6_) ) ;
 assign n1520 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1746 ) | ( n11  &  (~ n1746) ) ;
 assign n1521 = ( (~ PKSi_119_) ) | ( (~ PKSi_15_) ) ;
 assign n1522 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1748 ) | ( n11  &  (~ n1748) ) ;
 assign n1523 = ( (~ PKSi_106_) ) | ( (~ PKSi_5_) ) ;
 assign n1524 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1750 ) | ( n11  &  (~ n1750) ) ;
 assign n1525 = ( (~ PKSi_112_) ) | ( (~ PKSi_9_) ) ;
 assign n1526 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1752 ) | ( n11  &  (~ n1752) ) ;
 assign n1527 = ( (~ PKSi_19_) ) | ( (~ N_N2986) ) ;
 assign n1528 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1754 ) | ( n11  &  (~ n1754) ) ;
 assign n1529 = ( (~ PKSi_117_) ) | ( (~ PKSi_17_) ) ;
 assign n1530 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1756 ) | ( n11  &  (~ n1756) ) ;
 assign n1531 = ( (~ PKSi_99_) ) | ( (~ N_N2853) ) ;
 assign n1532 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1758 ) | ( n11  &  (~ n1758) ) ;
 assign n1533 = ( (~ PKSi_11_) ) | ( (~ N_N2982) ) ;
 assign n1534 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1760 ) | ( n11  &  (~ n1760) ) ;
 assign n1535 = ( (~ PKSi_110_) ) | ( (~ PKSi_2_) ) ;
 assign n1536 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1762 ) | ( n11  &  (~ n1762) ) ;
 assign n1537 = ( (~ PKSi_103_) ) | ( (~ PKSi_14_) ) ;
 assign n1538 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1764 ) | ( n11  &  (~ n1764) ) ;
 assign n1539 = ( (~ PKSi_96_) ) | ( (~ PKSi_22_) ) ;
 assign n1540 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1766 ) | ( n11  &  (~ n1766) ) ;
 assign n1541 = ( (~ PKSi_115_) ) | ( (~ PKSi_0_) ) ;
 assign n1542 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1768 ) | ( n11  &  (~ n1768) ) ;
 assign n1543 = ( (~ PKSi_8_) ) | ( (~ N_N2976) ) ;
 assign n1544 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1770 ) | ( n11  &  (~ n1770) ) ;
 assign n1545 = ( (~ PKSi_108_) ) | ( (~ PKSi_18_) ) ;
 assign n1546 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1772 ) | ( n11  &  (~ n1772) ) ;
 assign n1547 = ( (~ PKSi_105_) ) | ( (~ PKSi_1_) ) ;
 assign n1548 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1774 ) | ( n11  &  (~ n1774) ) ;
 assign n1549 = ( (~ PKSi_114_) ) | ( (~ N_N2843) ) ;
 assign n1550 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1776 ) | ( n11  &  (~ n1776) ) ;
 assign n1551 = ( (~ PKSi_100_) ) | ( (~ PKSi_13_) ) ;
 assign n1552 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1778 ) | ( n11  &  (~ n1778) ) ;
 assign n1553 = ( (~ PKSi_107_) ) | ( (~ PKSi_21_) ) ;
 assign n1554 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1780 ) | ( n11  &  (~ n1780) ) ;
 assign n1555 = ( (~ PKSi_109_) ) | ( (~ PKSi_10_) ) ;
 assign n1556 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1782 ) | ( n11  &  (~ n1782) ) ;
 assign n1557 = ( (~ PKSi_116_) ) | ( (~ N_N2838) ) ;
 assign n1558 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1784 ) | ( n11  &  (~ n1784) ) ;
 assign n1559 = ( (~ PKSi_104_) ) | ( (~ PKSi_12_) ) ;
 assign n1560 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1786 ) | ( n11  &  (~ n1786) ) ;
 assign n1561 = ( (~ PKSi_97_) ) | ( (~ PKSi_3_) ) ;
 assign n1562 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1788 ) | ( n11  &  (~ n1788) ) ;
 assign n1563 = ( (~ PKSi_113_) ) | ( (~ N_N2834) ) ;
 assign n1564 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1790 ) | ( n11  &  (~ n1790) ) ;
 assign n1565 = ( (~ PKSi_16_) ) | ( (~ N_N2964) ) ;
 assign n1566 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1792 ) | ( n11  &  (~ n1792) ) ;
 assign n1567 = ( (~ PKSi_101_) ) | ( (~ PKSi_20_) ) ;
 assign n1568 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1794 ) | ( n11  &  (~ n1794) ) ;
 assign n1569 = ( (~ PKSi_111_) ) | ( (~ PKSi_7_) ) ;
 assign n1570 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1796 ) | ( n11  &  (~ n1796) ) ;
 assign n1571 = ( (~ PKSi_142_) ) | ( (~ PKSi_28_) ) ;
 assign n1572 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1798 ) | ( n11  &  (~ n1798) ) ;
 assign n1573 = ( (~ PKSi_126_) ) | ( (~ PKSi_47_) ) ;
 assign n1574 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1800 ) | ( n11  &  (~ n1800) ) ;
 assign n1575 = ( (~ PKSi_122_) ) | ( (~ PKSi_30_) ) ;
 assign n1576 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1802 ) | ( n11  &  (~ n1802) ) ;
 assign n1577 = ( (~ wire282) ) | ( (~ PKSi_39_) ) ;
 assign n1578 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1804 ) | ( n11  &  (~ n1804) ) ;
 assign n1579 = ( (~ PKSi_130_) ) | ( (~ PKSi_29_) ) ;
 assign n1580 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1806 ) | ( n11  &  (~ n1806) ) ;
 assign n1581 = ( (~ PKSi_136_) ) | ( (~ PKSi_33_) ) ;
 assign n1582 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1808 ) | ( n11  &  (~ n1808) ) ;
 assign n1583 = ( (~ PKSi_43_) ) | ( (~ N_N2954) ) ;
 assign n1584 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1810 ) | ( n11  &  (~ n1810) ) ;
 assign n1585 = ( (~ PKSi_141_) ) | ( (~ PKSi_41_) ) ;
 assign n1586 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1812 ) | ( n11  &  (~ n1812) ) ;
 assign n1587 = ( (~ PKSi_123_) ) | ( (~ N_N2821) ) ;
 assign n1588 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1814 ) | ( n11  &  (~ n1814) ) ;
 assign n1589 = ( (~ PKSi_35_) ) | ( (~ N_N2950) ) ;
 assign n1590 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1816 ) | ( n11  &  (~ n1816) ) ;
 assign n1591 = ( (~ PKSi_134_) ) | ( (~ PKSi_26_) ) ;
 assign n1592 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1818 ) | ( n11  &  (~ n1818) ) ;
 assign n1593 = ( (~ PKSi_127_) ) | ( (~ PKSi_38_) ) ;
 assign n1594 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1820 ) | ( n11  &  (~ n1820) ) ;
 assign n1595 = ( (~ PKSi_120_) ) | ( (~ PKSi_46_) ) ;
 assign n1596 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1822 ) | ( n11  &  (~ n1822) ) ;
 assign n1597 = ( (~ PKSi_24_) ) | ( (~ N_N2945) ) ;
 assign n1598 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1824 ) | ( n11  &  (~ n1824) ) ;
 assign n1599 = ( (~ PKSi_32_) ) | ( (~ N_N2943) ) ;
 assign n1600 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1826 ) | ( n11  &  (~ n1826) ) ;
 assign n1601 = ( (~ PKSi_132_) ) | ( (~ PKSi_42_) ) ;
 assign n1602 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1828 ) | ( n11  &  (~ n1828) ) ;
 assign n1603 = ( (~ PKSi_129_) ) | ( (~ PKSi_25_) ) ;
 assign n1604 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1830 ) | ( n11  &  (~ n1830) ) ;
 assign n1605 = ( (~ PKSi_138_) ) | ( (~ N_N2811) ) ;
 assign n1606 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1832 ) | ( n11  &  (~ n1832) ) ;
 assign n1607 = ( (~ PKSi_124_) ) | ( (~ PKSi_37_) ) ;
 assign n1608 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1834 ) | ( n11  &  (~ n1834) ) ;
 assign n1609 = ( (~ PKSi_131_) ) | ( (~ PKSi_45_) ) ;
 assign n1610 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1836 ) | ( n11  &  (~ n1836) ) ;
 assign n1611 = ( (~ PKSi_133_) ) | ( (~ PKSi_34_) ) ;
 assign n1612 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1838 ) | ( n11  &  (~ n1838) ) ;
 assign n1613 = ( (~ PKSi_140_) ) | ( (~ N_N2806) ) ;
 assign n1614 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1840 ) | ( n11  &  (~ n1840) ) ;
 assign n1615 = ( (~ PKSi_128_) ) | ( (~ PKSi_36_) ) ;
 assign n1616 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1842 ) | ( n11  &  (~ n1842) ) ;
 assign n1617 = ( (~ PKSi_121_) ) | ( (~ PKSi_27_) ) ;
 assign n1618 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1844 ) | ( n11  &  (~ n1844) ) ;
 assign n1619 = ( (~ PKSi_137_) ) | ( (~ N_N2802) ) ;
 assign n1620 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1846 ) | ( n11  &  (~ n1846) ) ;
 assign n1621 = ( (~ PKSi_40_) ) | ( (~ N_N2931) ) ;
 assign n1622 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1848 ) | ( n11  &  (~ n1848) ) ;
 assign n1623 = ( (~ PKSi_125_) ) | ( (~ PKSi_44_) ) ;
 assign n1624 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1850 ) | ( n11  &  (~ n1850) ) ;
 assign n1625 = ( (~ PKSi_135_) ) | ( (~ PKSi_31_) ) ;
 assign n1626 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1852 ) | ( n11  &  (~ n1852) ) ;
 assign n1627 = ( (~ PKSi_166_) ) | ( (~ PKSi_52_) ) ;
 assign n1628 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1854 ) | ( n11  &  (~ n1854) ) ;
 assign n1629 = ( (~ PKSi_150_) ) | ( (~ PKSi_71_) ) ;
 assign n1630 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1856 ) | ( n11  &  (~ n1856) ) ;
 assign n1631 = ( (~ PKSi_146_) ) | ( (~ PKSi_54_) ) ;
 assign n1632 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1858 ) | ( n11  &  (~ n1858) ) ;
 assign n1633 = ( (~ PKSi_167_) ) | ( (~ PKSi_63_) ) ;
 assign n1634 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1860 ) | ( n11  &  (~ n1860) ) ;
 assign n1635 = ( (~ PKSi_154_) ) | ( (~ PKSi_53_) ) ;
 assign n1636 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1862 ) | ( n11  &  (~ n1862) ) ;
 assign n1637 = ( (~ PKSi_160_) ) | ( (~ PKSi_57_) ) ;
 assign n1638 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1864 ) | ( n11  &  (~ n1864) ) ;
 assign n1639 = ( (~ PKSi_67_) ) | ( (~ N_N2921) ) ;
 assign n1640 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1866 ) | ( n11  &  (~ n1866) ) ;
 assign n1641 = ( (~ PKSi_165_) ) | ( (~ PKSi_65_) ) ;
 assign n1642 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1868 ) | ( n11  &  (~ n1868) ) ;
 assign n1643 = ( (~ PKSi_147_) ) | ( (~ N_N2789) ) ;
 assign n1644 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1870 ) | ( n11  &  (~ n1870) ) ;
 assign n1645 = ( (~ PKSi_59_) ) | ( (~ N_N2917) ) ;
 assign n1646 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1872 ) | ( n11  &  (~ n1872) ) ;
 assign n1647 = ( (~ PKSi_158_) ) | ( (~ PKSi_50_) ) ;
 assign n1648 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1874 ) | ( n11  &  (~ n1874) ) ;
 assign n1649 = ( (~ PKSi_151_) ) | ( (~ PKSi_62_) ) ;
 assign n1650 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1876 ) | ( n11  &  (~ n1876) ) ;
 assign n1651 = ( (~ PKSi_144_) ) | ( (~ PKSi_70_) ) ;
 assign n1652 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1878 ) | ( n11  &  (~ n1878) ) ;
 assign n1653 = ( (~ PKSi_163_) ) | ( (~ PKSi_48_) ) ;
 assign n1654 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1880 ) | ( n11  &  (~ n1880) ) ;
 assign n1655 = ( (~ PKSi_153_) ) | ( (~ PKSi_56_) ) ;
 assign n1656 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1882 ) | ( n11  &  (~ n1882) ) ;
 assign n1657 = ( (~ PKSi_156_) ) | ( (~ PKSi_66_) ) ;
 assign n1658 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1884 ) | ( n11  &  (~ n1884) ) ;
 assign n1659 = ( (~ PKSi_49_) ) | ( (~ N_N2909) ) ;
 assign n1660 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1886 ) | ( n11  &  (~ n1886) ) ;
 assign n1661 = ( (~ PKSi_162_) ) | ( (~ N_N2779) ) ;
 assign n1662 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1888 ) | ( n11  &  (~ n1888) ) ;
 assign n1663 = ( (~ PKSi_148_) ) | ( (~ PKSi_61_) ) ;
 assign n1664 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1890 ) | ( n11  &  (~ n1890) ) ;
 assign n1665 = ( (~ PKSi_155_) ) | ( (~ PKSi_69_) ) ;
 assign n1666 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1892 ) | ( n11  &  (~ n1892) ) ;
 assign n1667 = ( (~ PKSi_157_) ) | ( (~ PKSi_58_) ) ;
 assign n1668 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1894 ) | ( n11  &  (~ n1894) ) ;
 assign n1669 = ( (~ PKSi_164_) ) | ( (~ N_N2774) ) ;
 assign n1670 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1896 ) | ( n11  &  (~ n1896) ) ;
 assign n1671 = ( (~ PKSi_152_) ) | ( (~ PKSi_60_) ) ;
 assign n1672 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1898 ) | ( n11  &  (~ n1898) ) ;
 assign n1673 = ( (~ PKSi_145_) ) | ( (~ PKSi_51_) ) ;
 assign n1674 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1900 ) | ( n11  &  (~ n1900) ) ;
 assign n1675 = ( (~ PKSi_161_) ) | ( (~ N_N2770) ) ;
 assign n1676 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1902 ) | ( n11  &  (~ n1902) ) ;
 assign n1677 = ( (~ PKSi_64_) ) | ( (~ N_N2899) ) ;
 assign n1678 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1904 ) | ( n11  &  (~ n1904) ) ;
 assign n1679 = ( (~ PKSi_149_) ) | ( (~ PKSi_68_) ) ;
 assign n1680 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1906 ) | ( n11  &  (~ n1906) ) ;
 assign n1681 = ( (~ PKSi_159_) ) | ( (~ PKSi_55_) ) ;
 assign n1682 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1908 ) | ( n11  &  (~ n1908) ) ;
 assign n1683 = ( (~ PKSi_190_) ) | ( (~ PKSi_76_) ) ;
 assign n1684 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1910 ) | ( n11  &  (~ n1910) ) ;
 assign n1685 = ( (~ PKSi_174_) ) | ( (~ PKSi_95_) ) ;
 assign n1686 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1912 ) | ( n11  &  (~ n1912) ) ;
 assign n1687 = ( (~ PKSi_170_) ) | ( (~ PKSi_78_) ) ;
 assign n1688 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1914 ) | ( n11  &  (~ n1914) ) ;
 assign n1689 = ( (~ wire234) ) | ( (~ PKSi_87_) ) ;
 assign n1690 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1916 ) | ( n11  &  (~ n1916) ) ;
 assign n1691 = ( (~ PKSi_178_) ) | ( (~ PKSi_77_) ) ;
 assign n1692 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1918 ) | ( n11  &  (~ n1918) ) ;
 assign n1693 = ( (~ PKSi_184_) ) | ( (~ PKSi_81_) ) ;
 assign n1694 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1920 ) | ( n11  &  (~ n1920) ) ;
 assign n1695 = ( (~ PKSi_91_) ) | ( (~ N_N2889) ) ;
 assign n1696 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1922 ) | ( n11  &  (~ n1922) ) ;
 assign n1697 = ( (~ PKSi_189_) ) | ( (~ PKSi_89_) ) ;
 assign n1698 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1924 ) | ( n11  &  (~ n1924) ) ;
 assign n1699 = ( (~ PKSi_171_) ) | ( (~ N_N2757) ) ;
 assign n1700 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1926 ) | ( n11  &  (~ n1926) ) ;
 assign n1701 = ( (~ PKSi_83_) ) | ( (~ N_N2885) ) ;
 assign n1702 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1928 ) | ( n11  &  (~ n1928) ) ;
 assign n1703 = ( (~ PKSi_182_) ) | ( (~ PKSi_74_) ) ;
 assign n1704 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1930 ) | ( n11  &  (~ n1930) ) ;
 assign n1705 = ( (~ PKSi_175_) ) | ( (~ PKSi_86_) ) ;
 assign n1706 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1932 ) | ( n11  &  (~ n1932) ) ;
 assign n1707 = ( (~ PKSi_94_) ) | ( (~ N_N2881) ) ;
 assign n1708 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1934 ) | ( n11  &  (~ n1934) ) ;
 assign n1709 = ( (~ PKSi_72_) ) | ( (~ N_N2879) ) ;
 assign n1710 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1936 ) | ( n11  &  (~ n1936) ) ;
 assign n1711 = ( (~ PKSi_80_) ) | ( (~ N_N2877) ) ;
 assign n1712 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1938 ) | ( n11  &  (~ n1938) ) ;
 assign n1713 = ( (~ PKSi_180_) ) | ( (~ N_N2749) ) ;
 assign n1714 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1940 ) | ( n11  &  (~ n1940) ) ;
 assign n1715 = ( (~ PKSi_177_) ) | ( (~ PKSi_73_) ) ;
 assign n1716 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1942 ) | ( n11  &  (~ n1942) ) ;
 assign n1717 = ( (~ PKSi_186_) ) | ( (~ N_N2746) ) ;
 assign n1718 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1944 ) | ( n11  &  (~ n1944) ) ;
 assign n1719 = ( (~ PKSi_172_) ) | ( (~ PKSi_85_) ) ;
 assign n1720 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1946 ) | ( n11  &  (~ n1946) ) ;
 assign n1721 = ( (~ PKSi_179_) ) | ( (~ PKSi_93_) ) ;
 assign n1722 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1948 ) | ( n11  &  (~ n1948) ) ;
 assign n1723 = ( (~ wire253) ) | ( (~ PKSi_82_) ) ;
 assign n1724 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1950 ) | ( n11  &  (~ n1950) ) ;
 assign n1725 = ( (~ PKSi_188_) ) | ( (~ N_N2741) ) ;
 assign n1726 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1952 ) | ( n11  &  (~ n1952) ) ;
 assign n1727 = ( (~ PKSi_176_) ) | ( (~ PKSi_84_) ) ;
 assign n1728 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1954 ) | ( n11  &  (~ n1954) ) ;
 assign n1729 = ( (~ PKSi_169_) ) | ( (~ PKSi_75_) ) ;
 assign n1730 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1956 ) | ( n11  &  (~ n1956) ) ;
 assign n1731 = ( (~ PKSi_185_) ) | ( (~ N_N2737) ) ;
 assign n1732 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1958 ) | ( n11  &  (~ n1958) ) ;
 assign n1733 = ( (~ wire333) ) | ( (~ N_N2865) ) ;
 assign n1734 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1960 ) | ( n11  &  (~ n1960) ) ;
 assign n1735 = ( (~ PKSi_173_) ) | ( (~ PKSi_92_) ) ;
 assign n1736 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1962 ) | ( n11  &  (~ n1962) ) ;
 assign n1737 = ( (~ PKSi_183_) ) | ( (~ PKSi_79_) ) ;
 assign n1738 = ( n11  &  (~ n1741) ) | ( (~ n1741)  &  n1964 ) | ( n11  &  (~ n1964) ) ;
 assign n1740 = ( PKSi_4_ ) | ( PKSi_118_ ) ;
 assign n1744 = ( PKSi_23_ ) | ( PKSi_102_ ) ;
 assign n1746 = ( PKSi_6_ ) | ( PKSi_98_ ) ;
 assign n1748 = ( PKSi_15_ ) | ( PKSi_119_ ) ;
 assign n1750 = ( PKSi_5_ ) | ( PKSi_106_ ) ;
 assign n1752 = ( PKSi_9_ ) | ( PKSi_112_ ) ;
 assign n1754 = ( PKSi_19_ ) | ( N_N2986 ) ;
 assign n1756 = ( PKSi_17_ ) | ( PKSi_117_ ) ;
 assign n1758 = ( N_N2853 ) | ( PKSi_99_ ) ;
 assign n1760 = ( PKSi_11_ ) | ( N_N2982 ) ;
 assign n1762 = ( PKSi_2_ ) | ( PKSi_110_ ) ;
 assign n1764 = ( PKSi_14_ ) | ( PKSi_103_ ) ;
 assign n1766 = ( PKSi_22_ ) | ( PKSi_96_ ) ;
 assign n1768 = ( PKSi_0_ ) | ( PKSi_115_ ) ;
 assign n1770 = ( PKSi_8_ ) | ( N_N2976 ) ;
 assign n1772 = ( PKSi_18_ ) | ( PKSi_108_ ) ;
 assign n1774 = ( PKSi_1_ ) | ( PKSi_105_ ) ;
 assign n1776 = ( N_N2843 ) | ( PKSi_114_ ) ;
 assign n1778 = ( PKSi_13_ ) | ( PKSi_100_ ) ;
 assign n1780 = ( PKSi_21_ ) | ( PKSi_107_ ) ;
 assign n1782 = ( PKSi_10_ ) | ( PKSi_109_ ) ;
 assign n1784 = ( N_N2838 ) | ( PKSi_116_ ) ;
 assign n1786 = ( PKSi_12_ ) | ( PKSi_104_ ) ;
 assign n1788 = ( PKSi_3_ ) | ( PKSi_97_ ) ;
 assign n1790 = ( N_N2834 ) | ( PKSi_113_ ) ;
 assign n1792 = ( PKSi_16_ ) | ( N_N2964 ) ;
 assign n1794 = ( PKSi_20_ ) | ( PKSi_101_ ) ;
 assign n1796 = ( PKSi_7_ ) | ( PKSi_111_ ) ;
 assign n1798 = ( PKSi_28_ ) | ( PKSi_142_ ) ;
 assign n1800 = ( PKSi_47_ ) | ( PKSi_126_ ) ;
 assign n1802 = ( PKSi_30_ ) | ( PKSi_122_ ) ;
 assign n1804 = ( PKSi_39_ ) | ( wire282 ) ;
 assign n1806 = ( PKSi_29_ ) | ( PKSi_130_ ) ;
 assign n1808 = ( PKSi_33_ ) | ( PKSi_136_ ) ;
 assign n1810 = ( PKSi_43_ ) | ( N_N2954 ) ;
 assign n1812 = ( PKSi_41_ ) | ( PKSi_141_ ) ;
 assign n1814 = ( N_N2821 ) | ( PKSi_123_ ) ;
 assign n1816 = ( PKSi_35_ ) | ( N_N2950 ) ;
 assign n1818 = ( PKSi_26_ ) | ( PKSi_134_ ) ;
 assign n1820 = ( PKSi_38_ ) | ( PKSi_127_ ) ;
 assign n1822 = ( PKSi_46_ ) | ( PKSi_120_ ) ;
 assign n1824 = ( PKSi_24_ ) | ( N_N2945 ) ;
 assign n1826 = ( PKSi_32_ ) | ( N_N2943 ) ;
 assign n1828 = ( PKSi_42_ ) | ( PKSi_132_ ) ;
 assign n1830 = ( PKSi_25_ ) | ( PKSi_129_ ) ;
 assign n1832 = ( N_N2811 ) | ( PKSi_138_ ) ;
 assign n1834 = ( PKSi_37_ ) | ( PKSi_124_ ) ;
 assign n1836 = ( PKSi_45_ ) | ( PKSi_131_ ) ;
 assign n1838 = ( PKSi_34_ ) | ( PKSi_133_ ) ;
 assign n1840 = ( N_N2806 ) | ( PKSi_140_ ) ;
 assign n1842 = ( PKSi_36_ ) | ( PKSi_128_ ) ;
 assign n1844 = ( PKSi_27_ ) | ( PKSi_121_ ) ;
 assign n1846 = ( N_N2802 ) | ( PKSi_137_ ) ;
 assign n1848 = ( PKSi_40_ ) | ( N_N2931 ) ;
 assign n1850 = ( PKSi_44_ ) | ( PKSi_125_ ) ;
 assign n1852 = ( PKSi_31_ ) | ( PKSi_135_ ) ;
 assign n1854 = ( PKSi_52_ ) | ( PKSi_166_ ) ;
 assign n1856 = ( PKSi_71_ ) | ( PKSi_150_ ) ;
 assign n1858 = ( PKSi_54_ ) | ( PKSi_146_ ) ;
 assign n1860 = ( PKSi_63_ ) | ( PKSi_167_ ) ;
 assign n1862 = ( PKSi_53_ ) | ( PKSi_154_ ) ;
 assign n1864 = ( PKSi_57_ ) | ( PKSi_160_ ) ;
 assign n1866 = ( PKSi_67_ ) | ( N_N2921 ) ;
 assign n1868 = ( PKSi_65_ ) | ( PKSi_165_ ) ;
 assign n1870 = ( N_N2789 ) | ( PKSi_147_ ) ;
 assign n1872 = ( PKSi_59_ ) | ( N_N2917 ) ;
 assign n1874 = ( PKSi_50_ ) | ( PKSi_158_ ) ;
 assign n1876 = ( PKSi_62_ ) | ( PKSi_151_ ) ;
 assign n1878 = ( PKSi_70_ ) | ( PKSi_144_ ) ;
 assign n1880 = ( PKSi_48_ ) | ( PKSi_163_ ) ;
 assign n1882 = ( PKSi_56_ ) | ( PKSi_153_ ) ;
 assign n1884 = ( PKSi_66_ ) | ( PKSi_156_ ) ;
 assign n1886 = ( PKSi_49_ ) | ( N_N2909 ) ;
 assign n1888 = ( N_N2779 ) | ( PKSi_162_ ) ;
 assign n1890 = ( PKSi_61_ ) | ( PKSi_148_ ) ;
 assign n1892 = ( PKSi_69_ ) | ( PKSi_155_ ) ;
 assign n1894 = ( PKSi_58_ ) | ( PKSi_157_ ) ;
 assign n1896 = ( N_N2774 ) | ( PKSi_164_ ) ;
 assign n1898 = ( PKSi_60_ ) | ( PKSi_152_ ) ;
 assign n1900 = ( PKSi_51_ ) | ( PKSi_145_ ) ;
 assign n1902 = ( N_N2770 ) | ( PKSi_161_ ) ;
 assign n1904 = ( PKSi_64_ ) | ( N_N2899 ) ;
 assign n1906 = ( PKSi_68_ ) | ( PKSi_149_ ) ;
 assign n1908 = ( PKSi_55_ ) | ( PKSi_159_ ) ;
 assign n1910 = ( PKSi_76_ ) | ( PKSi_190_ ) ;
 assign n1912 = ( PKSi_95_ ) | ( PKSi_174_ ) ;
 assign n1914 = ( PKSi_78_ ) | ( PKSi_170_ ) ;
 assign n1916 = ( PKSi_87_ ) | ( wire234 ) ;
 assign n1918 = ( PKSi_77_ ) | ( PKSi_178_ ) ;
 assign n1920 = ( PKSi_81_ ) | ( PKSi_184_ ) ;
 assign n1922 = ( PKSi_91_ ) | ( N_N2889 ) ;
 assign n1924 = ( PKSi_89_ ) | ( PKSi_189_ ) ;
 assign n1926 = ( N_N2757 ) | ( PKSi_171_ ) ;
 assign n1928 = ( PKSi_83_ ) | ( N_N2885 ) ;
 assign n1930 = ( PKSi_74_ ) | ( PKSi_182_ ) ;
 assign n1932 = ( PKSi_86_ ) | ( PKSi_175_ ) ;
 assign n1934 = ( PKSi_94_ ) | ( N_N2881 ) ;
 assign n1936 = ( PKSi_72_ ) | ( N_N2879 ) ;
 assign n1938 = ( PKSi_80_ ) | ( N_N2877 ) ;
 assign n1940 = ( N_N2749 ) | ( PKSi_180_ ) ;
 assign n1942 = ( PKSi_73_ ) | ( PKSi_177_ ) ;
 assign n1944 = ( N_N2746 ) | ( PKSi_186_ ) ;
 assign n1946 = ( PKSi_85_ ) | ( PKSi_172_ ) ;
 assign n1948 = ( PKSi_93_ ) | ( PKSi_179_ ) ;
 assign n1950 = ( PKSi_82_ ) | ( wire253 ) ;
 assign n1952 = ( N_N2741 ) | ( PKSi_188_ ) ;
 assign n1954 = ( PKSi_84_ ) | ( PKSi_176_ ) ;
 assign n1956 = ( PKSi_75_ ) | ( PKSi_169_ ) ;
 assign n1958 = ( N_N2737 ) | ( PKSi_185_ ) ;
 assign n1960 = ( wire333 ) | ( N_N2865 ) ;
 assign n1962 = ( PKSi_92_ ) | ( PKSi_173_ ) ;
 assign n1964 = ( PKSi_79_ ) | ( PKSi_183_ ) ;
 assign n1966 = ( Pencrypt_0_  &  (~ Pcount_0_) ) | ( Pencrypt_0_  &  n1287 ) | ( Pcount_0_  &  n1287 ) ;
 assign n1967 = ( Pcount_0_ ) | ( n1287 ) ;
 assign n1968 = ( Pcount_1_ ) | ( Pcount_2_ ) ;
 assign PKSi_191_ = ( wire234 ) ;
 assign PKSi_187_ = ( wire234 ) ;
 assign PKSi_181_ = ( wire253 ) ;
 assign PKSi_168_ = ( wire253 ) ;
 assign PKSi_143_ = ( wire282 ) ;
 assign PKSi_139_ = ( wire282 ) ;
 assign PKSi_90_ = ( wire333 ) ;
 assign PKSi_88_ = ( wire333 ) ;


endmodule

