module splax6xv (i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, i_13_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_, i_15_, o_1_, o_19_, o_2_, o_0_, o_29_, o_39_, o_38_, o_25_, o_12_, o_37_, o_26_, o_11_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_43_, o_30_, o_44_, o_41_, o_42_, o_20_, o_45_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

	input i_9_;
	input i_10_;
	input i_7_;
	input i_8_;
	input i_5_;
	input i_6_;
	input i_14_;
	input i_3_;
	input i_13_;
	input i_4_;
	input i_12_;
	input i_1_;
	input i_11_;
	input i_2_;
	input i_0_;
	input i_15_;
	output o_1_;
	output o_19_;
	output o_2_;
	output o_0_;
	output o_29_;
	output o_39_;
	output o_38_;
	output o_25_;
	output o_12_;
	output o_37_;
	output o_26_;
	output o_11_;
	output o_36_;
	output o_27_;
	output o_14_;
	output o_35_;
	output o_28_;
	output o_13_;
	output o_34_;
	output o_21_;
	output o_16_;
	output o_40_;
	output o_33_;
	output o_22_;
	output o_15_;
	output o_32_;
	output o_23_;
	output o_18_;
	output o_31_;
	output o_24_;
	output o_17_;
	output o_43_;
	output o_30_;
	output o_44_;
	output o_41_;
	output o_42_;
	output o_20_;
	output o_45_;
	output o_10_;
	output o_9_;
	output o_7_;
	output o_8_;
	output o_5_;
	output o_6_;
	output o_3_;
	output o_4_;

	wire [2491 : 0] sk /* synthesis noprune */;

	lut_sub lut_3 ({sk[0], i_3_, i_1_, i_2_, i_0_, n_n245, x428x}, o_1_);
	defparam lut_3.LUT_SIZE = 7;
	defparam lut_3.mask = 128'h3fffffffffffffff77f777f77ff777f7;

	lut_sub lut_8 ({sk[1], i_5_, i_3_, i_4_, n_n5144, x736x}, o_19_);
	defparam lut_8.LUT_SIZE = 6;
	defparam lut_8.mask = 64'h55ffffff33333373;

	lut_sub lut_11 ({sk[2], i_5_, i_3_, i_4_, n_n5144, x736x, x453x}, o_2_);
	defparam lut_11.LUT_SIZE = 7;
	defparam lut_11.mask = 128'h0fffffff0fffffff5f5f5f5f7f5f5f5f;

	lut_sub lut_15 ({sk[3], i_3_, i_1_, i_2_, i_0_, n_n222}, o_0_);
	defparam lut_15.LUT_SIZE = 6;
	defparam lut_15.mask = 64'h77ff77ff5d5dfd5d;

	lut_sub lut_20 ({sk[4], x16911x, x729x, n_n149, x763x, x398x, x5027x}, o_29_);
	defparam lut_20.LUT_SIZE = 7;
	defparam lut_20.mask = 128'h0fffffff0fffffff5555557fffffffff;

	lut_sub lut_25 ({sk[5], n_n4721, n_n373, n_n374, x16929x, x16930x}, o_39_);
	defparam lut_25.LUT_SIZE = 6;
	defparam lut_25.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_31 ({sk[6], x17175x, x17159x, n_n4397, n_n4399}, o_38_);
	defparam lut_31.LUT_SIZE = 5;
	defparam lut_31.mask = 32'h77777fff;

	lut_sub lut_36 ({sk[7], i_7_, i_6_, i_3_, i_4_, n_n5144, n_n159}, o_25_);
	defparam lut_36.LUT_SIZE = 7;
	defparam lut_36.mask = 128'h00ff55ffffffffff3333333333373333;

	lut_sub lut_39 ({sk[8], x17408x, n_n2225, x17249x, x17401x, x17402x, x17403x}, o_12_);
	defparam lut_39.LUT_SIZE = 7;
	defparam lut_39.mask = 128'h00ff55ffffffffff7fffffffffffffff;

	lut_sub lut_46 ({sk[9], x17586x, x17582x, n_n4103, n_n4102}, o_37_);
	defparam lut_46.LUT_SIZE = 5;
	defparam lut_46.mask = 32'h3f3f7fff;

	lut_sub lut_51 ({sk[10], n_n5144, x4221x, x17592x, n_n2953, x17600x, x17601x}, o_26_);
	defparam lut_51.LUT_SIZE = 7;
	defparam lut_51.mask = 128'h00ff55ffffffffff7fffffffffffffff;

	lut_sub lut_58 ({sk[11], n_n2213, n_n51, n_n13, x569x, x17609x, x17610x}, o_11_);
	defparam lut_58.LUT_SIZE = 7;
	defparam lut_58.mask = 128'h00ff55ffffffffff7f7f7fffffffffff;

	lut_sub lut_64 ({sk[12], n_n3783, n_n3785, x17846x, x17847x}, o_36_);
	defparam lut_64.LUT_SIZE = 5;
	defparam lut_64.mask = 32'h3f3f7fff;

	lut_sub lut_69 ({sk[13], n_n5144, n_n2977, n_n2976, n_n2974, n_n2975, x17860x}, o_27_);
	defparam lut_69.LUT_SIZE = 7;
	defparam lut_69.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_76 ({sk[14], n_n2621, n_n2622, x17908x, x21377x}, o_14_);
	defparam lut_76.LUT_SIZE = 5;
	defparam lut_76.mask = 32'h1f1fbfff;

	lut_sub lut_81 ({sk[15], x18148x, x18144x, n_n3458, x18026x, x18027x, x18141x}, o_35_);
	defparam lut_81.LUT_SIZE = 7;
	defparam lut_81.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_88 ({sk[16], x18167x, n_n157, n_n2998, x18155x, x746x, x1525x}, o_28_);
	defparam lut_88.LUT_SIZE = 7;
	defparam lut_88.mask = 128'h55ff55ff55ff55ff0fff7fffffffffff;

	lut_sub lut_94 ({sk[17], n_n3027, n_n4308, n_n3085, n_n6268, x512x, x18223x}, o_13_);
	defparam lut_94.LUT_SIZE = 7;
	defparam lut_94.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_101 ({sk[18], x18214x, x18292x, n_n3033, n_n3393, x18295x, x18296x}, o_34_);
	defparam lut_101.LUT_SIZE = 7;
	defparam lut_101.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_108 ({sk[19], n_n5144, n_n65, x77x, n_n10, x525x, x270x}, o_21_);
	defparam lut_108.LUT_SIZE = 7;
	defparam lut_108.mask = 128'h55ff55ff55ff55ff373f3f3fffffffff;

	lut_sub lut_114 ({sk[20], x18313x, n_n33, x18304x, x52x, x63x, x1887x}, o_16_);
	defparam lut_114.LUT_SIZE = 7;
	defparam lut_114.mask = 128'h55ff55ff55ff55ff00ff7fffffffffff;

	lut_sub lut_120 ({sk[21], n_n5144, x725x, n_n6, n_n184, x267x, x768x}, o_40_);
	defparam lut_120.LUT_SIZE = 7;
	defparam lut_120.mask = 128'h55ff55ff55ff55ff00550357ffffffff;

	lut_sub lut_124 ({sk[22], x18330x, x530x, n_n5, x370x, x404x, x18327x}, o_33_);
	defparam lut_124.LUT_SIZE = 7;
	defparam lut_124.mask = 128'h55ff55ff55ff55ff557fffffffffffff;

	lut_sub lut_130 ({sk[23], n_n5144, n_n51, n_n14, x185x, x270x, x267x}, o_22_);
	defparam lut_130.LUT_SIZE = 7;
	defparam lut_130.mask = 128'h55ff55ff55ff55ff003f557fffffffff;

	lut_sub lut_135 ({sk[24], n_n5144, x18355x, x18344x, x18347x, x18348x, x21368x}, o_15_);
	defparam lut_135.LUT_SIZE = 7;
	defparam lut_135.mask = 128'h55ff55ff55ff55ffbfffffffffffffff;

	lut_sub lut_142 ({sk[25], n_n3166, x421x}, o_32_);
	defparam lut_142.LUT_SIZE = 3;
	defparam lut_142.mask = 8'h57;

	lut_sub lut_145 ({sk[26], x18512x, n_n2927, x18495x, x18498x, x18499x, x18507x}, o_23_);
	defparam lut_145.LUT_SIZE = 7;
	defparam lut_145.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_152 ({sk[27], x18526x, n_n2803, n_n2805, n_n2812, x21454x}, o_18_);
	defparam lut_152.LUT_SIZE = 6;
	defparam lut_152.mask = 64'h11ffffffbfffffff;

	lut_sub lut_158 ({sk[28], i_7_, i_6_, n_n5144, x18572x, n_n7346, x748x}, o_31_);
	defparam lut_158.LUT_SIZE = 7;
	defparam lut_158.mask = 128'h55ff55ff55ff55ff3fff3fff3fff7fff;

	lut_sub lut_163 ({sk[29], i_7_, i_6_, i_3_, i_4_, n_n5144, n_n159}, o_24_);
	defparam lut_163.LUT_SIZE = 7;
	defparam lut_163.mask = 128'h55ff55ff55ff55ff3333333733333333;

	lut_sub lut_166 ({sk[30], x18622x, n_n2747, x18615x, x18616x}, o_17_);
	defparam lut_166.LUT_SIZE = 5;
	defparam lut_166.mask = 32'h1f1f7fff;

	lut_sub lut_171 ({sk[31], x18684x, x18655x, x18656x, n_n4753, x18693x, x18694x}, o_43_);
	defparam lut_171.LUT_SIZE = 7;
	defparam lut_171.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_178 ({sk[32], n_n3028, x18214x, x18292x, n_n3033, n_n3393}, o_30_);
	defparam lut_178.LUT_SIZE = 6;
	defparam lut_178.mask = 64'h11ffffff7fffffff;

	lut_sub lut_184 ({sk[33], x18795x, x18790x, x18791x, x18792x}, o_44_);
	defparam lut_184.LUT_SIZE = 5;
	defparam lut_184.mask = 32'h1f1f7fff;

	lut_sub lut_189 ({sk[34], i_8_, n_n5144, n_n162, n_n184, n_n18, n_n163}, o_41_);
	defparam lut_189.LUT_SIZE = 7;
	defparam lut_189.mask = 128'h55ff55ff55ff55ff0001ffff0000ffff;

	lut_sub lut_192 ({sk[35], x18802x, x18803x, x18804x, x18805x}, o_42_);
	defparam lut_192.LUT_SIZE = 5;
	defparam lut_192.mask = 32'h1f1f7fff;

	lut_sub lut_197 ({sk[36], i_5_, i_3_, i_4_, n_n5144, x736x}, o_20_);
	defparam lut_197.LUT_SIZE = 6;
	defparam lut_197.mask = 64'h11ffffff33373333;

	lut_sub lut_200 ({sk[37], x421x, x18818x}, o_45_);
	defparam lut_200.LUT_SIZE = 3;
	defparam lut_200.mask = 8'h57;

	lut_sub lut_203 ({sk[38], n_n5144, x19036x, x19029x, x19027x, x19028x}, o_10_);
	defparam lut_203.LUT_SIZE = 6;
	defparam lut_203.mask = 64'h11ffffff7fffffff;

	lut_sub lut_209 ({sk[39], n_n1139, x19348x, x19349x, x19457x, x19458x}, o_9_);
	defparam lut_209.LUT_SIZE = 6;
	defparam lut_209.mask = 64'h11ffffff7fffffff;

	lut_sub lut_215 ({sk[40], x19503x, x19504x, x19682x, x19683x, x19689x}, o_7_);
	defparam lut_215.LUT_SIZE = 6;
	defparam lut_215.mask = 64'h11ffffff7fffffff;

	lut_sub lut_221 ({sk[41], i_3_, i_1_, i_2_, i_0_}, o_8_);
	defparam lut_221.LUT_SIZE = 5;
	defparam lut_221.mask = 32'h1f1f00a0;

	lut_sub lut_224 ({sk[42], x19914x, x19870x, x19871x}, o_5_);
	defparam lut_224.LUT_SIZE = 4;
	defparam lut_224.mask = 16'h557f;

	lut_sub lut_228 ({sk[43], i_8_, n_n16, x288x, x780x, x19920x, x19921x}, o_6_);
	defparam lut_228.LUT_SIZE = 7;
	defparam lut_228.mask = 128'h55ff55ff55ff55ff7777777f77777777;

	lut_sub lut_232 ({sk[44], n_n5144, x530x, n_n7259, n_n3389, x468x, x19927x}, o_3_);
	defparam lut_232.LUT_SIZE = 7;
	defparam lut_232.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_239 ({sk[45], x19946x, n_n3, n_n275, x936x, x19941x}, o_4_);
	defparam lut_239.LUT_SIZE = 6;
	defparam lut_239.mask = 64'h11ffffff5f7fffff;

	lut_sub lut_244 ({sk[46], x16870x, x386x, n_n7259, x463x, x1369x, x16862x}, n_n245);
	defparam lut_244.LUT_SIZE = 7;
	defparam lut_244.mask = 128'h55ff55ff55ff55ff1fffffffffffffff;

	lut_sub lut_250 ({sk[47], i_7_, i_5_, i_6_, i_3_, i_4_, n_n219}, x428x);
	defparam lut_250.LUT_SIZE = 7;
	defparam lut_250.mask = 128'h55ff55ff55ff55ff1010000010000000;

	lut_sub lut_254 ({sk[48], i_3_, i_1_, i_2_, i_0_}, n_n5144);
	defparam lut_254.LUT_SIZE = 5;
	defparam lut_254.mask = 32'h1f1f22a2;

	lut_sub lut_257 ({sk[49], i_7_, i_8_, i_6_, x725x, n_n184, n_n163}, x736x);
	defparam lut_257.LUT_SIZE = 7;
	defparam lut_257.mask = 128'h55ff55ff55ff55ff0100000000000000;

	lut_sub lut_259 ({sk[50], i_7_, i_8_, i_6_, n_n135, n_n162, n_n163}, x453x);
	defparam lut_259.LUT_SIZE = 7;
	defparam lut_259.mask = 128'h55ff55ff55ff55ff0000000001000000;

	lut_sub lut_261 ({sk[51], x736x, n_n162, n_n231, x16886x, x16895x, x16896x}, n_n222);
	defparam lut_261.LUT_SIZE = 7;
	defparam lut_261.mask = 128'h55ff55ff55ff55ff7fff7fff7fffffff;

	lut_sub lut_267 ({sk[52], n_n65, n_n71, n_n89, n_n12, x1042x, x16910x}, x16911x);
	defparam lut_267.LUT_SIZE = 7;
	defparam lut_267.mask = 128'h55ff55ff55ff55ff55775f7f77777f7f;

	lut_sub lut_272 ({sk[53], i_14_, i_13_, i_12_, i_15_}, x729x);
	defparam lut_272.LUT_SIZE = 5;
	defparam lut_272.mask = 32'h1f1f0800;

	lut_sub lut_274 ({sk[54], i_9_, i_10_, i_11_}, n_n149);
	defparam lut_274.LUT_SIZE = 4;
	defparam lut_274.mask = 16'h5520;

	lut_sub lut_276 ({sk[55], i_7_, i_8_, i_6_, n_n159, n_n111, n_n48}, x763x);
	defparam lut_276.LUT_SIZE = 7;
	defparam lut_276.mask = 128'h55ff55ff55ff55ff0703000000000000;

	lut_sub lut_280 ({sk[56], i_5_, i_3_, i_4_, n_n159, n_n124, n_n2}, x398x);
	defparam lut_280.LUT_SIZE = 7;
	defparam lut_280.mask = 128'h55ff55ff55ff55ff5557555555555555;

	lut_sub lut_283 ({sk[57], x729x, n_n156, x763x, n_n3, n_n2, n_n191}, x5027x);
	defparam lut_283.LUT_SIZE = 7;
	defparam lut_283.mask = 128'h55ff55ff55ff55ff0000000015553fff;

	lut_sub lut_290 ({sk[58], i_7_, i_8_, i_6_, x740x, x244x, x1595x}, n_n4721);
	defparam lut_290.LUT_SIZE = 7;
	defparam lut_290.mask = 128'h55ff55ff55ff55ff0005000700000000;

	lut_sub lut_294 ({sk[59], n_n124, x740x, n_n126, x244x, x235x, x236x}, n_n373);
	defparam lut_294.LUT_SIZE = 7;
	defparam lut_294.mask = 128'h55ff55ff55ff55ff0000007700000f7f;

	lut_sub lut_298 ({sk[60], n_n124, x740x, x140x, n_n126, x235x, x236x}, n_n374);
	defparam lut_298.LUT_SIZE = 7;
	defparam lut_298.mask = 128'h55ff55ff55ff55ff0000000f0000777f;

	lut_sub lut_302 ({sk[61], n_n5144, n_n38, n_n134, n_n6642, x390x, x712x}, x16929x);
	defparam lut_302.LUT_SIZE = 7;
	defparam lut_302.mask = 128'h55ff55ff55ff55ff7f7f7fffffffffff;

	lut_sub lut_308 ({sk[62], n_n124, x740x, n_n969, n_n519, n_n4597, x140x}, x16930x);
	defparam lut_308.LUT_SIZE = 7;
	defparam lut_308.mask = 128'h55ff55ff55ff55ff3fff3fff3fff7fff;

	lut_sub lut_313 ({sk[63], x16961x, x16962x, n_n4400, x17173x}, x17175x);
	defparam lut_313.LUT_SIZE = 5;
	defparam lut_313.mask = 32'h1f1f7fff;

	lut_sub lut_318 ({sk[64], x543x, n_n4408, x17093x, x17155x, x17156x, x21405x}, x17159x);
	defparam lut_318.LUT_SIZE = 7;
	defparam lut_318.mask = 128'h55ff55ff55ff55ffbfffffffffffffff;

	lut_sub lut_325 ({sk[65], n_n4191, x549x, n_n4404, n_n4403, x17060x, x17063x}, n_n4397);
	defparam lut_325.LUT_SIZE = 7;
	defparam lut_325.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_332 ({sk[66], x17120x, x17121x, n_n4409, x17149x}, n_n4399);
	defparam lut_332.LUT_SIZE = 5;
	defparam lut_332.mask = 32'h1f1f7fff;

	lut_sub lut_337 ({sk[67], i_1_, i_2_, i_0_}, n_n159);
	defparam lut_337.LUT_SIZE = 4;
	defparam lut_337.mask = 16'h5508;

	lut_sub lut_339 ({sk[68], x17347x, x17348x, n_n2231, n_n2234, n_n2233}, x17408x);
	defparam lut_339.LUT_SIZE = 6;
	defparam lut_339.mask = 64'h11ffffff7fffffff;

	lut_sub lut_345 ({sk[69], x17218x, x17228x, x17229x, x21397x}, n_n2225);
	defparam lut_345.LUT_SIZE = 5;
	defparam lut_345.mask = 32'h1f1f7fff;

	lut_sub lut_350 ({sk[70], x4639x, x17241x, n_n2235, x17245x, x17247x}, x17249x);
	defparam lut_350.LUT_SIZE = 6;
	defparam lut_350.mask = 64'h11ffffff7fffffff;

	lut_sub lut_356 ({sk[71], n_n5144, x17192x, n_n2253, x17185x, x17186x}, x17401x);
	defparam lut_356.LUT_SIZE = 6;
	defparam lut_356.mask = 64'h11ffffff7fffffff;

	lut_sub lut_362 ({sk[72], x17213x, x17277x, x17278x, x21455x}, x17402x);
	defparam lut_362.LUT_SIZE = 5;
	defparam lut_362.mask = 32'h1f1fbfff;

	lut_sub lut_367 ({sk[73], x17304x, x17305x, x17328x, x17325x, x17326x}, x17403x);
	defparam lut_367.LUT_SIZE = 6;
	defparam lut_367.mask = 64'h11ffffff7fffffff;

	lut_sub lut_373 ({sk[74], n_n4105, x17453x, x17454x, x17584x}, x17586x);
	defparam lut_373.LUT_SIZE = 5;
	defparam lut_373.mask = 32'h1f1f7fff;

	lut_sub lut_378 ({sk[75], x17466x, x17467x, n_n4116, x17578x, x17579x}, x17582x);
	defparam lut_378.LUT_SIZE = 6;
	defparam lut_378.mask = 64'h11ffffff7fffffff;

	lut_sub lut_384 ({sk[76], n_n4136, x17486x, x17487x, x543x, x17514x, x17500x}, n_n4103);
	defparam lut_384.LUT_SIZE = 7;
	defparam lut_384.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_391 ({sk[77], x17539x, x17540x, x17552x, x17553x, x17564x, x17565x}, n_n4102);
	defparam lut_391.LUT_SIZE = 7;
	defparam lut_391.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_398 ({sk[78], n_n149, n_n4, x717x, n_n3, n_n2}, x4221x);
	defparam lut_398.LUT_SIZE = 6;
	defparam lut_398.mask = 64'h11ffffff0000070f;

	lut_sub lut_402 ({sk[79], i_5_, x286x, n_n3, n_n2, x231x, x170x}, x17592x);
	defparam lut_402.LUT_SIZE = 7;
	defparam lut_402.mask = 128'h55ff55ff55ff55ff0555377705550555;

	lut_sub lut_406 ({sk[80], n_n9, n_n4, n_n144, n_n6, n_n5, x170x}, n_n2953);
	defparam lut_406.LUT_SIZE = 7;
	defparam lut_406.mask = 128'h55ff55ff55ff55ff153f557f15ff55ff;

	lut_sub lut_413 ({sk[81], i_7_, i_6_, n_n7254, x746x, x17590x, x17598x}, x17600x);
	defparam lut_413.LUT_SIZE = 7;
	defparam lut_413.mask = 128'h55ff55ff55ff55ff7fff7fff77ff77ff;

	lut_sub lut_419 ({sk[82], x569x, n_n7263, n_n14, n_n7255, x170x, n_n2954}, x17601x);
	defparam lut_419.LUT_SIZE = 7;
	defparam lut_419.mask = 128'h55ff55ff55ff55ff5f7fffffffffffff;

	lut_sub lut_425 ({sk[83], n_n135, n_n71, n_n13, n_n4, n_n59, x1495x}, n_n2213);
	defparam lut_425.LUT_SIZE = 7;
	defparam lut_425.mask = 128'h55ff55ff55ff55ff05370f3f05ff0fff;

	lut_sub lut_430 ({sk[84], i_9_, i_10_, i_11_, x725x}, n_n51);
	defparam lut_430.LUT_SIZE = 5;
	defparam lut_430.mask = 32'h1f1f0400;

	lut_sub lut_432 ({sk[85], i_7_, i_8_, i_6_, n_n159, n_n111}, n_n13);
	defparam lut_432.LUT_SIZE = 6;
	defparam lut_432.mask = 64'h11ffffff00100000;

	lut_sub lut_434 ({sk[86], i_7_, i_6_, i_1_, i_2_, i_0_, n_n111}, x569x);
	defparam lut_434.LUT_SIZE = 7;
	defparam lut_434.mask = 128'h55ff55ff55ff55ff1000100000000000;

	lut_sub lut_437 ({sk[87], i_7_, i_6_, n_n5144, n_n111, n_n19}, x17609x);
	defparam lut_437.LUT_SIZE = 6;
	defparam lut_437.mask = 64'h11ffffff1f1f1f1f;

	lut_sub lut_443 ({sk[88], i_7_, i_8_, i_6_, x288x, x77x, x568x}, x17610x);
	defparam lut_443.LUT_SIZE = 7;
	defparam lut_443.mask = 128'h55ff55ff55ff55ff575555555f555f55;

	lut_sub lut_447 ({sk[89], x17697x, x17659x, x17660x, x17684x, x17685x}, n_n3783);
	defparam lut_447.LUT_SIZE = 6;
	defparam lut_447.mask = 64'h11ffffff7fffffff;

	lut_sub lut_453 ({sk[90], x17778x, n_n3796, x17764x, x17765x}, n_n3785);
	defparam lut_453.LUT_SIZE = 5;
	defparam lut_453.mask = 32'h1f1f7fff;

	lut_sub lut_458 ({sk[91], n_n3794, x17839x, x17835x, x17836x, x17842x}, x17846x);
	defparam lut_458.LUT_SIZE = 6;
	defparam lut_458.mask = 64'h11ffffff7fffffff;

	lut_sub lut_464 ({sk[92], n_n3793, n_n3795, n_n3787, x17820x, x17821x}, x17847x);
	defparam lut_464.LUT_SIZE = 6;
	defparam lut_464.mask = 64'h11ffffff7fffffff;

	lut_sub lut_470 ({sk[93], i_8_, x568x, x750x, x145x, n_n18, x21407x}, n_n2977);
	defparam lut_470.LUT_SIZE = 7;
	defparam lut_470.mask = 128'h55ff55ff55ff55ffaaabffffaaaaffff;

	lut_sub lut_474 ({sk[94], n_n9, n_n14, n_n186, n_n10, x145x, n_n12}, n_n2976);
	defparam lut_474.LUT_SIZE = 7;
	defparam lut_474.mask = 128'h55ff55ff55ff55ff135f13ff337f33ff;

	lut_sub lut_481 ({sk[95], n_n4, n_n186, x145x, x748x, x231x, x1044x}, n_n2974);
	defparam lut_481.LUT_SIZE = 7;
	defparam lut_481.mask = 128'h55ff55ff55ff55ff035757570357ffff;

	lut_sub lut_486 ({sk[96], n_n9, n_n4, n_n186, n_n6, n_n5, x145x}, n_n2975);
	defparam lut_486.LUT_SIZE = 7;
	defparam lut_486.mask = 128'h55ff55ff55ff55ff153f557f15ff55ff;

	lut_sub lut_493 ({sk[97], i_7_, i_6_, x816x, x17857x, x17858x}, x17860x);
	defparam lut_493.LUT_SIZE = 6;
	defparam lut_493.mask = 64'h11ffffff7777777f;

	lut_sub lut_497 ({sk[98], x17867x, x17868x, x17869x, x17870x, x17874x, x17875x}, n_n2621);
	defparam lut_497.LUT_SIZE = 7;
	defparam lut_497.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_504 ({sk[99], n_n4461, x597x, x620x, x17882x, x21378x}, n_n2622);
	defparam lut_504.LUT_SIZE = 6;
	defparam lut_504.mask = 64'h11ffffffbfffffff;

	lut_sub lut_510 ({sk[100], x17893x, x17894x, x17899x, x17900x}, x17908x);
	defparam lut_510.LUT_SIZE = 5;
	defparam lut_510.mask = 32'h1f1f7fff;

	lut_sub lut_515 ({sk[101], n_n34, x765x, n_n2635, x1813x, x3836x, x17912x}, x21377x);
	defparam lut_515.LUT_SIZE = 7;
	defparam lut_515.mask = 128'h55ff55ff55ff55ff8800880080000000;

	lut_sub lut_518 ({sk[102], n_n3454, n_n3455, n_n3456, x18145x}, x18148x);
	defparam lut_518.LUT_SIZE = 5;
	defparam lut_518.mask = 32'h1f1f7fff;

	lut_sub lut_523 ({sk[103], n_n3464, n_n3463, n_n3460, n_n3462, x18078x, x18134x}, x18144x);
	defparam lut_523.LUT_SIZE = 7;
	defparam lut_523.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_530 ({sk[104], x17987x, x17988x, n_n3480, x17998x, x17999x}, n_n3458);
	defparam lut_530.LUT_SIZE = 6;
	defparam lut_530.mask = 64'h11ffffff7fffffff;

	lut_sub lut_536 ({sk[105], n_n39, n_n6642, n_n132, x434x, n_n3532, x21440x}, x18026x);
	defparam lut_536.LUT_SIZE = 7;
	defparam lut_536.mask = 128'h55ff55ff55ff55ffbfbfffffbfffffff;

	lut_sub lut_542 ({sk[106], n_n41, x1824x, x1880x, x18012x, x18013x, x18019x}, x18027x);
	defparam lut_542.LUT_SIZE = 7;
	defparam lut_542.mask = 128'h55ff55ff55ff55ff7f7f7f7f7fffffff;

	lut_sub lut_548 ({sk[107], x3773x, x17978x, x17981x, x17982x, x18137x, x18138x}, x18141x);
	defparam lut_548.LUT_SIZE = 7;
	defparam lut_548.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_555 ({sk[108], x398x, x3622x, x253x, n_n6, x1550x, x18165x}, x18167x);
	defparam lut_555.LUT_SIZE = 7;
	defparam lut_555.mask = 128'h55ff55ff55ff55ff557fffff55ffffff;

	lut_sub lut_561 ({sk[109], i_7_, i_6_}, n_n157);
	defparam lut_561.LUT_SIZE = 3;
	defparam lut_561.mask = 8'h58;

	lut_sub lut_563 ({sk[110], x253x, n_n10, n_n151, n_n12, x1462x, x18150x}, n_n2998);
	defparam lut_563.LUT_SIZE = 7;
	defparam lut_563.mask = 128'h55ff55ff55ff55ff557755775f7fffff;

	lut_sub lut_568 ({sk[111], i_7_, i_6_, x733x, n_n7253, x746x, x1525x}, x18155x);
	defparam lut_568.LUT_SIZE = 7;
	defparam lut_568.mask = 128'h55ff55ff55ff55ff0fff0f0f7fff0f0f;

	lut_sub lut_574 ({sk[112], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x746x);
	defparam lut_574.LUT_SIZE = 7;
	defparam lut_574.mask = 128'h55ff55ff55ff55ff0010000000000000;

	lut_sub lut_576 ({sk[113], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x1525x);
	defparam lut_576.LUT_SIZE = 7;
	defparam lut_576.mask = 128'h55ff55ff55ff55ff0000000010100000;

	lut_sub lut_579 ({sk[114], x18214x, n_n3033, n_n3393}, n_n3027);
	defparam lut_579.LUT_SIZE = 4;
	defparam lut_579.mask = 16'h557f;

	lut_sub lut_583 ({sk[115], i_7_, i_8_, i_6_, x740x, x157x}, n_n4308);
	defparam lut_583.LUT_SIZE = 6;
	defparam lut_583.mask = 64'h11ffffff00000100;

	lut_sub lut_585 ({sk[116], i_8_, x740x, x3607x, n_n18, x17554x, x1823x}, n_n3085);
	defparam lut_585.LUT_SIZE = 7;
	defparam lut_585.mask = 128'h55ff55ff55ff55ff33ff37ff33ff33ff;

	lut_sub lut_589 ({sk[117], i_7_, i_8_, i_6_, n_n170, x285x}, n_n6268);
	defparam lut_589.LUT_SIZE = 6;
	defparam lut_589.mask = 64'h11ffffff01000000;

	lut_sub lut_591 ({sk[118], i_7_, i_8_, i_6_, n_n156, x740x, x725x}, x512x);
	defparam lut_591.LUT_SIZE = 7;
	defparam lut_591.mask = 128'h55ff55ff55ff55ff0000000000010000;

	lut_sub lut_593 ({sk[119], n_n5144, n_n124, x435x, n_n177, x285x, x18221x}, x18223x);
	defparam lut_593.LUT_SIZE = 7;
	defparam lut_593.mask = 128'h55ff55ff55ff55ff55ff57ffffffffff;

	lut_sub lut_598 ({sk[120], x18184x, x18185x, x18187x, x18211x, x21373x}, x18214x);
	defparam lut_598.LUT_SIZE = 6;
	defparam lut_598.mask = 64'h11ffffffbfffffff;

	lut_sub lut_604 ({sk[121], n_n5144, n_n3031, n_n3042, n_n3029, x18266x, x21369x}, x18292x);
	defparam lut_604.LUT_SIZE = 7;
	defparam lut_604.mask = 128'h55ff55ff55ff55ffbfffffffffffffff;

	lut_sub lut_611 ({sk[122], x18170x, x18171x, x18175x, x18176x, x18180x}, n_n3033);
	defparam lut_611.LUT_SIZE = 6;
	defparam lut_611.mask = 64'h11ffffff7fffffff;

	lut_sub lut_617 ({sk[123], x18192x, x18193x, x18200x, x18201x, x18203x, x18204x}, n_n3393);
	defparam lut_617.LUT_SIZE = 7;
	defparam lut_617.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_624 ({sk[124], n_n41, x245x, n_n5055, n_n132, x150x, x4902x}, x18295x);
	defparam lut_624.LUT_SIZE = 7;
	defparam lut_624.mask = 128'h55ff55ff55ff55ff55ff55ff7fffffff;

	lut_sub lut_630 ({sk[125], n_n51, n_n41, n_n40, n_n5056, x608x, x1815x}, x18296x);
	defparam lut_630.LUT_SIZE = 7;
	defparam lut_630.mask = 128'h55ff55ff55ff55ff3f7f3f7f3f7fffff;

	lut_sub lut_635 ({sk[126], i_9_, i_10_, i_11_, x729x}, n_n65);
	defparam lut_635.LUT_SIZE = 5;
	defparam lut_635.mask = 32'h1f1f0400;

	lut_sub lut_637 ({sk[127], i_14_, i_13_, i_12_, i_15_, n_n149}, x77x);
	defparam lut_637.LUT_SIZE = 6;
	defparam lut_637.mask = 64'h11ffffff10004000;

	lut_sub lut_640 ({sk[128], i_7_, i_8_, i_6_, n_n162, n_n159}, n_n10);
	defparam lut_640.LUT_SIZE = 6;
	defparam lut_640.mask = 64'h11ffffff00000100;

	lut_sub lut_642 ({sk[129], i_9_, i_10_, i_11_, x725x, n_n7294, x751x}, x525x);
	defparam lut_642.LUT_SIZE = 7;
	defparam lut_642.mask = 128'h55ff55ff55ff55ff3333373333333333;

	lut_sub lut_645 ({sk[130], i_14_, i_13_, i_12_, i_15_, n_n191}, x270x);
	defparam lut_645.LUT_SIZE = 6;
	defparam lut_645.mask = 64'h11ffffff10404000;

	lut_sub lut_649 ({sk[131], n_n33, x127x, x1850x, x3442x, x18309x, x18310x}, x18313x);
	defparam lut_649.LUT_SIZE = 7;
	defparam lut_649.mask = 128'h55ff55ff55ff55ff7f7f7f7f7fffffff;

	lut_sub lut_655 ({sk[132], i_7_, i_8_, i_6_, x734x}, n_n33);
	defparam lut_655.LUT_SIZE = 5;
	defparam lut_655.mask = 32'h1f1f0040;

	lut_sub lut_657 ({sk[133], n_n33, n_n32, x130x, x48x, x1883x, n_n2733}, x18304x);
	defparam lut_657.LUT_SIZE = 7;
	defparam lut_657.mask = 128'h55ff55ff55ff55ff555577ff5f5f7fff;

	lut_sub lut_662 ({sk[134], i_14_, i_13_, i_12_, i_15_, n_n191}, x52x);
	defparam lut_662.LUT_SIZE = 6;
	defparam lut_662.mask = 64'h11ffffff11010000;

	lut_sub lut_666 ({sk[135], i_14_, i_13_, i_12_, i_15_, n_n191}, x63x);
	defparam lut_666.LUT_SIZE = 6;
	defparam lut_666.mask = 64'h11ffffff00004044;

	lut_sub lut_670 ({sk[136], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1887x);
	defparam lut_670.LUT_SIZE = 7;
	defparam lut_670.mask = 128'h55ff55ff55ff55ff5030353000500000;

	lut_sub lut_677 ({sk[137], i_14_, i_13_, i_12_, i_15_}, x725x);
	defparam lut_677.LUT_SIZE = 5;
	defparam lut_677.mask = 32'h1f1f8000;

	lut_sub lut_679 ({sk[138], i_7_, i_8_, i_6_, n_n159, n_n48}, n_n6);
	defparam lut_679.LUT_SIZE = 6;
	defparam lut_679.mask = 64'h11ffffff10000000;

	lut_sub lut_681 ({sk[139], i_9_, i_10_, i_11_}, n_n184);
	defparam lut_681.LUT_SIZE = 4;
	defparam lut_681.mask = 16'h5580;

	lut_sub lut_683 ({sk[140], i_7_, i_8_, i_6_, n_n159, n_n111}, x267x);
	defparam lut_683.LUT_SIZE = 6;
	defparam lut_683.mask = 64'h11ffffff00110000;

	lut_sub lut_686 ({sk[141], i_9_, i_10_, i_11_, x729x, x717x, x730x}, x768x);
	defparam lut_686.LUT_SIZE = 7;
	defparam lut_686.mask = 128'h55ff55ff55ff55ff00007f007f007f00;

	lut_sub lut_696 ({sk[142], n_n9, n_n3389, n_n3378, x388x, n_n151, x370x}, x18330x);
	defparam lut_696.LUT_SIZE = 7;
	defparam lut_696.mask = 128'h55ff55ff55ff55ff0fffffff7fffffff;

	lut_sub lut_702 ({sk[143], n_n65, n_n4, x77x, n_n259, x87x, x18322x}, x530x);
	defparam lut_702.LUT_SIZE = 7;
	defparam lut_702.mask = 128'h55ff55ff55ff55ff5f5f7fff5f5fffff;

	lut_sub lut_708 ({sk[144], i_7_, i_8_, i_6_, n_n159, n_n111}, n_n5);
	defparam lut_708.LUT_SIZE = 6;
	defparam lut_708.mask = 64'h11ffffff01000000;

	lut_sub lut_710 ({sk[145], i_14_, i_13_, i_12_, i_15_, n_n156}, x370x);
	defparam lut_710.LUT_SIZE = 6;
	defparam lut_710.mask = 64'h11ffffff00404000;

	lut_sub lut_713 ({sk[146], i_14_, i_13_, i_12_, i_15_, n_n156, n_n191}, x404x);
	defparam lut_713.LUT_SIZE = 7;
	defparam lut_713.mask = 128'h55ff55ff55ff55ff0300500050000000;

	lut_sub lut_717 ({sk[147], n_n5144, n_n9, n_n144, n_n7259, n_n10, x145x}, x18327x);
	defparam lut_717.LUT_SIZE = 7;
	defparam lut_717.mask = 128'h55ff55ff55ff55ff1f1f1fffffffffff;

	lut_sub lut_722 ({sk[148], i_7_, i_8_, i_6_, n_n159, n_n48}, n_n14);
	defparam lut_722.LUT_SIZE = 6;
	defparam lut_722.mask = 64'h11ffffff00000100;

	lut_sub lut_724 ({sk[149], i_14_, i_13_, i_12_, i_15_, n_n149}, x185x);
	defparam lut_724.LUT_SIZE = 6;
	defparam lut_724.mask = 64'h11ffffff10404000;

	lut_sub lut_728 ({sk[150], n_n112, x63x, n_n113, x1113x, x1112x, x18353x}, x18355x);
	defparam lut_728.LUT_SIZE = 7;
	defparam lut_728.mask = 128'h55ff55ff55ff55ff555f555f777fffff;

	lut_sub lut_733 ({sk[151], n_n59, n_n112, x613x, x222x, x628x, x697x}, x18344x);
	defparam lut_733.LUT_SIZE = 7;
	defparam lut_733.mask = 128'h55ff55ff55ff55ff77ff7fff77ffffff;

	lut_sub lut_739 ({sk[152], x734x, x725x, n_n161, n_n184, n_n1566, x217x}, x18347x);
	defparam lut_739.LUT_SIZE = 7;
	defparam lut_739.mask = 128'h55ff55ff55ff55ff333333333377337f;

	lut_sub lut_743 ({sk[153], n_n138, n_n42, x172x, n_n43, x216x, x526x}, x18348x);
	defparam lut_743.LUT_SIZE = 7;
	defparam lut_743.mask = 128'h55ff55ff55ff55ff575f575f575fffff;

	lut_sub lut_748 ({sk[154], n_n42, n_n43, n_n190, x1781x, x1786x, x1785x}, x21368x);
	defparam lut_748.LUT_SIZE = 7;
	defparam lut_748.mask = 128'h55ff55ff55ff55ffffffc0c0aa008000;

	lut_sub lut_753 ({sk[155], x608x, x18361x, n_n3177, n_n3176, x18360x, x18376x}, n_n3166);
	defparam lut_753.LUT_SIZE = 7;
	defparam lut_753.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_760 ({sk[156], n_n3173, n_n3175, x18436x, n_n3170, n_n3172, x18488x}, x421x);
	defparam lut_760.LUT_SIZE = 7;
	defparam lut_760.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_767 ({sk[157], x729x, n_n149, n_n2, n_n191, x87x, x18511x}, x18512x);
	defparam lut_767.LUT_SIZE = 7;
	defparam lut_767.mask = 128'h55ff55ff55ff55ff55775577557f55ff;

	lut_sub lut_772 ({sk[158], x729x, n_n9, x77x, n_n10, x238x, n_n191}, n_n2927);
	defparam lut_772.LUT_SIZE = 7;
	defparam lut_772.mask = 128'h55ff55ff55ff55ff030f333f030f777f;

	lut_sub lut_777 ({sk[159], n_n89, x77x, n_n14, x238x, n_n12, x18494x}, x18495x);
	defparam lut_777.LUT_SIZE = 7;
	defparam lut_777.mask = 128'h55ff55ff55ff55ff575f77ff77ff77ff;

	lut_sub lut_785 ({sk[160], x729x, n_n6, n_n5, x238x, n_n191, x3244x}, x18498x);
	defparam lut_785.LUT_SIZE = 7;
	defparam lut_785.mask = 128'h55ff55ff55ff55ff555f5f5f557f7f7f;

	lut_sub lut_791 ({sk[161], x729x, n_n149, n_n4, x77x, x270x, x18497x}, x18499x);
	defparam lut_791.LUT_SIZE = 7;
	defparam lut_791.mask = 128'h55ff55ff55ff55ff557f557f557f55ff;

	lut_sub lut_796 ({sk[162], x569x, n_n7255, n_n7254, n_n231, x18503x, x18504x}, x18507x);
	defparam lut_796.LUT_SIZE = 7;
	defparam lut_796.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_803 ({sk[163], n_n124, x46x, x735x, n_n126, x147x, x958x}, x18526x);
	defparam lut_803.LUT_SIZE = 7;
	defparam lut_803.mask = 128'h55ff55ff55ff55ff00070007007700ff;

	lut_sub lut_809 ({sk[164], n_n123, x18547x, x3220x, x18533x, x18541x, x1396x}, n_n2803);
	defparam lut_809.LUT_SIZE = 7;
	defparam lut_809.mask = 128'h55ff55ff55ff55ff3fffffff7fffffff;

	lut_sub lut_815 ({sk[165], n_n123, n_n2813, n_n125, x1696x, x1695x, x18561x}, n_n2805);
	defparam lut_815.LUT_SIZE = 7;
	defparam lut_815.mask = 128'h55ff55ff55ff55ff555fffff777fffff;

	lut_sub lut_820 ({sk[166], n_n124, x735x, n_n126, x52x, x1531x, x1530x}, n_n2812);
	defparam lut_820.LUT_SIZE = 7;
	defparam lut_820.mask = 128'h55ff55ff55ff55ff0000003300005f7f;

	lut_sub lut_824 ({sk[167], n_n5144, n_n123, n_n125, x1466x, x1465x, x21438x}, x21454x);
	defparam lut_824.LUT_SIZE = 7;
	defparam lut_824.mask = 128'h55ff55ff55ff55ffaa88a08000000000;

	lut_sub lut_829 ({sk[168], i_7_, i_5_, i_6_, i_3_, i_4_, n_n159}, x18572x);
	defparam lut_829.LUT_SIZE = 7;
	defparam lut_829.mask = 128'h55ff55ff55ff55ff0000010050410000;

	lut_sub lut_835 ({sk[169], i_7_, i_5_, i_6_, i_3_, i_4_, n_n159}, n_n7346);
	defparam lut_835.LUT_SIZE = 7;
	defparam lut_835.mask = 128'h55ff55ff55ff55ff0000000000100000;

	lut_sub lut_837 ({sk[170], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x748x);
	defparam lut_837.LUT_SIZE = 7;
	defparam lut_837.mask = 128'h55ff55ff55ff55ff0000000000000008;

	lut_sub lut_839 ({sk[171], n_n4441, x575x, x18577x, x18578x, x18621x}, x18622x);
	defparam lut_839.LUT_SIZE = 6;
	defparam lut_839.mask = 64'h11ffffff7fffffff;

	lut_sub lut_845 ({sk[172], x18584x, x18585x, x18589x, x18590x, x18591x, x18592x}, n_n2747);
	defparam lut_845.LUT_SIZE = 7;
	defparam lut_845.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_852 ({sk[173], i_8_, n_n17, x735x, n_n2760, x1654x, x3143x}, x18615x);
	defparam lut_852.LUT_SIZE = 7;
	defparam lut_852.mask = 128'h55ff55ff55ff55ff5f5f5f7f5f5f5f5f;

	lut_sub lut_856 ({sk[174], x18602x, x18603x, x18607x, x18608x}, x18616x);
	defparam lut_856.LUT_SIZE = 5;
	defparam lut_856.mask = 32'h1f1f7fff;

	lut_sub lut_861 ({sk[175], n_n108, x1024x, x18638x, n_n4762, x18680x, x18681x}, x18684x);
	defparam lut_861.LUT_SIZE = 7;
	defparam lut_861.mask = 128'h55ff55ff55ff55ff7fff7fff7fffffff;

	lut_sub lut_867 ({sk[176], x734x, n_n126, n_n148, x234x, x18652x, x21434x}, x18655x);
	defparam lut_867.LUT_SIZE = 7;
	defparam lut_867.mask = 128'h55ff55ff55ff55ffbbbbbbbbbbbbbfff;

	lut_sub lut_872 ({sk[177], x18641x, x18642x, x3111x, x18650x}, x18656x);
	defparam lut_872.LUT_SIZE = 5;
	defparam lut_872.mask = 32'h1f1f7fff;

	lut_sub lut_877 ({sk[178], n_n101, n_n4903, x544x, x1019x, n_n4763, x18668x}, n_n4753);
	defparam lut_877.LUT_SIZE = 7;
	defparam lut_877.mask = 128'h55ff55ff55ff55ff77ffffff7fffffff;

	lut_sub lut_883 ({sk[179], n_n42, n_n4774, x172x, n_n43, x1879x, x18691x}, x18693x);
	defparam lut_883.LUT_SIZE = 7;
	defparam lut_883.mask = 128'h55ff55ff55ff55ff5757ffff57ffffff;

	lut_sub lut_888 ({sk[180], x18627x, x18628x, x18631x, x18632x}, x18694x);
	defparam lut_888.LUT_SIZE = 5;
	defparam lut_888.mask = 32'h1f1f7fff;

	lut_sub lut_893 ({sk[181], x608x, n_n3034, x18712x, x18711x, x18716x, x18717x}, n_n3028);
	defparam lut_893.LUT_SIZE = 7;
	defparam lut_893.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_900 ({sk[182], x18684x, n_n4849, n_n4850, x18655x, x18656x, n_n4753}, x18795x);
	defparam lut_900.LUT_SIZE = 7;
	defparam lut_900.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_907 ({sk[183], n_n31, n_n30, x1021x, x1020x, x18776x, x18788x}, x18790x);
	defparam lut_907.LUT_SIZE = 7;
	defparam lut_907.mask = 128'h55ff55ff55ff55ff777777ff7f7f7fff;

	lut_sub lut_912 ({sk[184], n_n30, x646x, x2977x, x18783x, x18786x, x1096x}, x18791x);
	defparam lut_912.LUT_SIZE = 7;
	defparam lut_912.mask = 128'h55ff55ff55ff55ff3fffffff7fffffff;

	lut_sub lut_918 ({sk[185], n_n5144, n_n31, n_n4855, n_n4857, x794x, x18735x}, x18792x);
	defparam lut_918.LUT_SIZE = 7;
	defparam lut_918.mask = 128'h55ff55ff55ff55ff5fff7fffffffffff;

	lut_sub lut_924 ({sk[186], i_5_, i_3_, i_4_}, n_n162);
	defparam lut_924.LUT_SIZE = 4;
	defparam lut_924.mask = 16'h5508;

	lut_sub lut_926 ({sk[187], i_7_, i_6_}, n_n18);
	defparam lut_926.LUT_SIZE = 3;
	defparam lut_926.mask = 8'h51;

	lut_sub lut_928 ({sk[188], i_1_, i_2_, i_0_}, n_n163);
	defparam lut_928.LUT_SIZE = 4;
	defparam lut_928.mask = 16'h5504;

	lut_sub lut_930 ({sk[189], i_9_, i_10_, i_8_, i_11_, n_n17, x285x}, x18802x);
	defparam lut_930.LUT_SIZE = 7;
	defparam lut_930.mask = 128'h55ff55ff55ff55ff0001001001001000;

	lut_sub lut_935 ({sk[190], i_9_, i_10_, i_8_, i_11_, n_n16, x285x}, x18803x);
	defparam lut_935.LUT_SIZE = 7;
	defparam lut_935.mask = 128'h55ff55ff55ff55ff0001100001000010;

	lut_sub lut_940 ({sk[191], n_n5144, n_n149, n_n6266, n_n6268, n_n200, x285x}, x18804x);
	defparam lut_940.LUT_SIZE = 7;
	defparam lut_940.mask = 128'h55ff55ff55ff55ff0fff1fffffffffff;

	lut_sub lut_945 ({sk[192], x435x, n_n200, x419x, x445x, n_n170, x285x}, x18805x);
	defparam lut_945.LUT_SIZE = 7;
	defparam lut_945.mask = 128'h55ff55ff55ff55ff0fff1fffffffffff;

	lut_sub lut_950 ({sk[193], x608x, x18814x, x18815x, x18361x, x18360x, x18816x}, x18818x);
	defparam lut_950.LUT_SIZE = 7;
	defparam lut_950.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_957 ({sk[194], x708x, n_n1797, n_n1855, x19032x, x19034x}, x19036x);
	defparam lut_957.LUT_SIZE = 6;
	defparam lut_957.mask = 64'h11ffffff7fffffff;

	lut_sub lut_963 ({sk[195], n_n1807, x18929x, x18930x, x18950x, x18951x, n_n1803}, x19029x);
	defparam lut_963.LUT_SIZE = 7;
	defparam lut_963.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_970 ({sk[196], n_n1802, n_n1829, n_n1830, x19004x}, x19027x);
	defparam lut_970.LUT_SIZE = 5;
	defparam lut_970.mask = 32'h1f1f7fff;

	lut_sub lut_975 ({sk[197], x18874x, x18875x, x18900x, x18901x, x19022x, x19023x}, x19028x);
	defparam lut_975.LUT_SIZE = 7;
	defparam lut_975.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_982 ({sk[198], x19126x, n_n1150, x19097x, x19098x}, n_n1139);
	defparam lut_982.LUT_SIZE = 5;
	defparam lut_982.mask = 32'h1f1f7fff;

	lut_sub lut_987 ({sk[199], n_n1155, x19325x, x19326x, n_n1153}, x19348x);
	defparam lut_987.LUT_SIZE = 5;
	defparam lut_987.mask = 32'h1f1f7fff;

	lut_sub lut_992 ({sk[200], n_n1158, n_n1156, x19211x, x19278x, x19275x, x19276x}, x19349x);
	defparam lut_992.LUT_SIZE = 7;
	defparam lut_992.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_999 ({sk[201], n_n5144, n_n1146, n_n1145, n_n1148}, x19457x);
	defparam lut_999.LUT_SIZE = 5;
	defparam lut_999.mask = 32'h1f1f7fff;

	lut_sub lut_1004 ({sk[202], n_n1144, n_n1147, x19430x, x19431x, n_n1143}, x19458x);
	defparam lut_1004.LUT_SIZE = 6;
	defparam lut_1004.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1010 ({sk[203], n_n31, n_n30, x111x, n_n799, x1810x, x1809x}, x19503x);
	defparam lut_1010.LUT_SIZE = 7;
	defparam lut_1010.mask = 128'h55ff55ff55ff55ff0f0f3fff5f5f7fff;

	lut_sub lut_1015 ({sk[204], n_n34, x1711x, x19491x, x19498x, x19499x}, x19504x);
	defparam lut_1015.LUT_SIZE = 6;
	defparam lut_1015.mask = 64'h11ffffff7f7f7fff;

	lut_sub lut_1020 ({sk[205], x19559x, x19560x, n_n746, n_n747, n_n748}, x19682x);
	defparam lut_1020.LUT_SIZE = 6;
	defparam lut_1020.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1026 ({sk[206], n_n752, x19541x, n_n750, n_n751, x21343x}, x19683x);
	defparam lut_1026.LUT_SIZE = 6;
	defparam lut_1026.mask = 64'h11ffffffbfffffff;

	lut_sub lut_1032 ({sk[207], n_n31, x19478x, x1302x, x19466x, n_n756, x19688x}, x19689x);
	defparam lut_1032.LUT_SIZE = 7;
	defparam lut_1032.mask = 128'h55ff55ff55ff55ff7f7fffff7fffffff;

	lut_sub lut_1038 ({sk[208], x19893x, n_n296, n_n360, n_n362, x19890x, x19912x}, x19914x);
	defparam lut_1038.LUT_SIZE = 7;
	defparam lut_1038.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_1045 ({sk[209], x19738x, x19739x, x19757x, x19758x, x19868x}, x19870x);
	defparam lut_1045.LUT_SIZE = 6;
	defparam lut_1045.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1051 ({sk[210], n_n306, n_n301, n_n304, n_n305, n_n303, n_n302}, x19871x);
	defparam lut_1051.LUT_SIZE = 7;
	defparam lut_1051.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_1058 ({sk[211], i_7_, i_6_}, n_n16);
	defparam lut_1058.LUT_SIZE = 3;
	defparam lut_1058.mask = 8'h54;

	lut_sub lut_1060 ({sk[212], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x288x);
	defparam lut_1060.LUT_SIZE = 7;
	defparam lut_1060.mask = 128'h55ff55ff55ff55ff0800000000000000;

	lut_sub lut_1062 ({sk[213], i_9_, i_10_, i_11_, x729x, x717x, x730x}, x780x);
	defparam lut_1062.LUT_SIZE = 7;
	defparam lut_1062.mask = 128'h55ff55ff55ff55ff00000f007f007f00;

	lut_sub lut_1070 ({sk[214], i_7_, i_6_, n_n5144, n_n219, n_n162, n_n19}, x19920x);
	defparam lut_1070.LUT_SIZE = 7;
	defparam lut_1070.mask = 128'h55ff55ff55ff55ff13ff13ff13ff13ff;

	lut_sub lut_1080 ({sk[215], n_n135, n_n51, x288x, n_n126, n_n59, x454x}, x19921x);
	defparam lut_1080.LUT_SIZE = 7;
	defparam lut_1080.mask = 128'h55ff55ff55ff55ff5557555f555f555f;

	lut_sub lut_1085 ({sk[216], i_7_, i_6_, i_1_, i_2_, i_0_, n_n111}, n_n7259);
	defparam lut_1085.LUT_SIZE = 7;
	defparam lut_1085.mask = 128'h55ff55ff55ff55ff1000000000000000;

	lut_sub lut_1087 ({sk[217], i_7_, i_6_, i_1_, i_2_, i_0_, n_n111}, n_n3389);
	defparam lut_1087.LUT_SIZE = 7;
	defparam lut_1087.mask = 128'h55ff55ff55ff55ff0000100010001000;

	lut_sub lut_1091 ({sk[218], i_7_, i_8_, i_6_, x725x, x288x, n_n184}, x468x);
	defparam lut_1091.LUT_SIZE = 7;
	defparam lut_1091.mask = 128'h55ff55ff55ff55ff0000010100000000;

	lut_sub lut_1094 ({sk[219], i_8_, n_n16, x288x, x370x, x404x, x19925x}, x19927x);
	defparam lut_1094.LUT_SIZE = 7;
	defparam lut_1094.mask = 128'h55ff55ff55ff55ff5555557f55555555;

	lut_sub lut_1098 ({sk[220], x729x, x372x, n_n2, n_n191, x87x, x19945x}, x19946x);
	defparam lut_1098.LUT_SIZE = 7;
	defparam lut_1098.mask = 128'h55ff55ff55ff55ff557755ff557f55ff;

	lut_sub lut_1103 ({sk[221], i_8_, i_5_, i_3_, i_4_, n_n159, n_n16}, n_n3);
	defparam lut_1103.LUT_SIZE = 7;
	defparam lut_1103.mask = 128'h55ff55ff55ff55ff0100000000000000;

	lut_sub lut_1105 ({sk[222], i_7_, i_6_, n_n219, x744x, x525x, n_n48}, n_n275);
	defparam lut_1105.LUT_SIZE = 7;
	defparam lut_1105.mask = 128'h55ff55ff55ff55ff3f7f3f7f3f7f3f3f;

	lut_sub lut_1114 ({sk[223], i_9_, i_10_, i_11_, x729x, x717x, x730x}, x936x);
	defparam lut_1114.LUT_SIZE = 7;
	defparam lut_1114.mask = 128'h55ff55ff55ff55ff00000f007f007f00;

	lut_sub lut_1122 ({sk[224], x725x, n_n191, n_n7242, x462x, x751x, x19940x}, x19941x);
	defparam lut_1122.LUT_SIZE = 7;
	defparam lut_1122.mask = 128'h55ff55ff55ff55ff5fff5fff5fff7fff;

	lut_sub lut_1127 ({sk[225], x453x, n_n3389, x388x, n_n7252, x567x, n_n7262}, x16870x);
	defparam lut_1127.LUT_SIZE = 7;
	defparam lut_1127.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_1134 ({sk[226], i_3_, i_1_, i_2_, i_0_}, x386x);
	defparam lut_1134.LUT_SIZE = 5;
	defparam lut_1134.mask = 32'h1f1f0040;

	lut_sub lut_1136 ({sk[227], i_7_, i_6_, i_1_, i_2_, i_0_, n_n48}, x463x);
	defparam lut_1136.LUT_SIZE = 7;
	defparam lut_1136.mask = 128'h55ff55ff55ff55ff0000000010001000;

	lut_sub lut_1139 ({sk[228], i_5_, i_3_, i_4_, x725x, n_n184, x717x}, x1369x);
	defparam lut_1139.LUT_SIZE = 7;
	defparam lut_1139.mask = 128'h55ff55ff55ff55ff0300000000110000;

	lut_sub lut_1142 ({sk[229], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x16862x);
	defparam lut_1142.LUT_SIZE = 7;
	defparam lut_1142.mask = 128'h55ff55ff55ff55ff2000000000000000;

	lut_sub lut_1144 ({sk[230], i_7_, i_5_, i_6_, i_3_, i_4_, n_n19}, n_n231);
	defparam lut_1144.LUT_SIZE = 7;
	defparam lut_1144.mask = 128'h55ff55ff55ff55ff4040404040404050;

	lut_sub lut_1154 ({sk[231], i_3_, i_1_, i_2_, i_0_, x423x}, x16886x);
	defparam lut_1154.LUT_SIZE = 6;
	defparam lut_1154.mask = 64'h11ffffff55557755;

	lut_sub lut_1158 ({sk[232], i_3_, n_n219, x711x, x569x, n_n19, x567x}, x16895x);
	defparam lut_1158.LUT_SIZE = 7;
	defparam lut_1158.mask = 128'h55ff55ff55ff55ff5fff5fff7fffffff;

	lut_sub lut_1164 ({sk[233], i_7_, i_5_, i_6_, i_3_, i_4_, n_n219}, x16896x);
	defparam lut_1164.LUT_SIZE = 7;
	defparam lut_1164.mask = 128'h55ff55ff55ff55ff0000405050405050;

	lut_sub lut_1175 ({sk[234], i_9_, i_10_, i_11_, x729x}, n_n71);
	defparam lut_1175.LUT_SIZE = 5;
	defparam lut_1175.mask = 32'h1f1f0004;

	lut_sub lut_1177 ({sk[235], i_9_, i_10_, i_11_, x729x}, n_n89);
	defparam lut_1177.LUT_SIZE = 5;
	defparam lut_1177.mask = 32'h1f1f0040;

	lut_sub lut_1179 ({sk[236], i_7_, i_8_, i_6_, n_n159, n_n48}, n_n12);
	defparam lut_1179.LUT_SIZE = 6;
	defparam lut_1179.mask = 64'h11ffffff01000000;

	lut_sub lut_1181 ({sk[237], i_7_, i_8_, i_6_, n_n162, n_n159, n_n48}, x1042x);
	defparam lut_1181.LUT_SIZE = 7;
	defparam lut_1181.mask = 128'h55ff55ff55ff55ff0013000000130000;

	lut_sub lut_1186 ({sk[238], i_9_, i_10_, i_11_, n_n5144, x729x, n_n9}, x16910x);
	defparam lut_1186.LUT_SIZE = 7;
	defparam lut_1186.mask = 128'h55ff55ff55ff55ff0f0f0f0f0f0f1f0f;

	lut_sub lut_1189 ({sk[239], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x740x);
	defparam lut_1189.LUT_SIZE = 7;
	defparam lut_1189.mask = 128'h55ff55ff55ff55ff0000000000800000;

	lut_sub lut_1191 ({sk[240], i_14_, i_13_, i_12_, i_15_, n_n156}, x244x);
	defparam lut_1191.LUT_SIZE = 6;
	defparam lut_1191.mask = 64'h11ffffff00000144;

	lut_sub lut_1195 ({sk[241], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1595x);
	defparam lut_1195.LUT_SIZE = 7;
	defparam lut_1195.mask = 128'h55ff55ff55ff55ff0000007707070770;

	lut_sub lut_1208 ({sk[242], x132x, n_n36, x126x, n_n4569, x4970x, x16960x}, x16961x);
	defparam lut_1208.LUT_SIZE = 7;
	defparam lut_1208.mask = 128'h55ff55ff55ff55ff7f7f7fff7f7fffff;

	lut_sub lut_1214 ({sk[243], n_n36, n_n4169, x942x, x16950x, x16955x, x16956x}, x16962x);
	defparam lut_1214.LUT_SIZE = 7;
	defparam lut_1214.mask = 128'h55ff55ff55ff55ff7f7fffff7fffffff;

	lut_sub lut_1220 ({sk[244], x16975x, n_n4154, x16967x, x4961x, x16974x}, n_n4400);
	defparam lut_1220.LUT_SIZE = 6;
	defparam lut_1220.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1226 ({sk[245], x16943x, x599x, n_n33, x1783x, x17169x, x17170x}, x17173x);
	defparam lut_1226.LUT_SIZE = 7;
	defparam lut_1226.mask = 128'h55ff55ff55ff55ff777fffffffffffff;

	lut_sub lut_1232 ({sk[246], n_n40, x714x, x17002x, x984x, x983x, x17345x}, x17347x);
	defparam lut_1232.LUT_SIZE = 7;
	defparam lut_1232.mask = 128'h55ff55ff55ff55ff5555555f7777777f;

	lut_sub lut_1236 ({sk[247], x17342x, x4531x, x17331x, x17333x, x21403x}, x17348x);
	defparam lut_1236.LUT_SIZE = 6;
	defparam lut_1236.mask = 64'h11ffffffbfffffff;

	lut_sub lut_1242 ({sk[248], x17355x, x17358x, x17359x, x17363x, x21401x}, n_n2231);
	defparam lut_1242.LUT_SIZE = 6;
	defparam lut_1242.mask = 64'h11ffffffbfffffff;

	lut_sub lut_1248 ({sk[249], x17379x, x17369x, x17370x, x4482x, x17375x}, n_n2234);
	defparam lut_1248.LUT_SIZE = 6;
	defparam lut_1248.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1254 ({sk[250], x17389x, x17390x, x17393x, x17394x, x17397x, x17398x}, n_n2233);
	defparam lut_1254.LUT_SIZE = 7;
	defparam lut_1254.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_1261 ({sk[251], n_n4119, n_n4154, x17430x, x17431x, x17433x}, n_n4105);
	defparam lut_1261.LUT_SIZE = 6;
	defparam lut_1261.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1267 ({sk[252], n_n36, n_n4169, x950x, x17451x}, x17453x);
	defparam lut_1267.LUT_SIZE = 5;
	defparam lut_1267.mask = 32'h1f1f5f7f;

	lut_sub lut_1271 ({sk[253], x17438x, x17439x, x17445x, x17446x}, x17454x);
	defparam lut_1271.LUT_SIZE = 5;
	defparam lut_1271.mask = 32'h1f1f7fff;

	lut_sub lut_1276 ({sk[254], n_n5144, x599x, x17412x, x17420x, x21387x}, x17584x);
	defparam lut_1276.LUT_SIZE = 6;
	defparam lut_1276.mask = 64'h11ffffffbfffffff;

	lut_sub lut_1282 ({sk[255], i_9_, i_10_, i_11_, x725x}, n_n135);
	defparam lut_1282.LUT_SIZE = 5;
	defparam lut_1282.mask = 32'h1f1f4000;

	lut_sub lut_1284 ({sk[256], i_7_, i_8_, i_6_, n_n159, n_n111}, n_n4);
	defparam lut_1284.LUT_SIZE = 6;
	defparam lut_1284.mask = 64'h11ffffff10000000;

	lut_sub lut_1286 ({sk[257], i_9_, i_10_, i_11_, x725x}, n_n59);
	defparam lut_1286.LUT_SIZE = 5;
	defparam lut_1286.mask = 32'h1f1f0040;

	lut_sub lut_1288 ({sk[258], i_9_, i_10_, i_11_, x729x, x717x, x730x}, x1495x);
	defparam lut_1288.LUT_SIZE = 7;
	defparam lut_1288.mask = 128'h55ff55ff55ff55ff00000f007f007700;

	lut_sub lut_1295 ({sk[259], n_n3467, x17932x, x17933x, x17934x}, n_n3454);
	defparam lut_1295.LUT_SIZE = 5;
	defparam lut_1295.mask = 32'h1f1f7fff;

	lut_sub lut_1300 ({sk[260], x3810x, x3811x, x17948x, x17949x, x17951x, x17952x}, n_n3455);
	defparam lut_1300.LUT_SIZE = 7;
	defparam lut_1300.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_1307 ({sk[261], x17958x, x17959x, x17961x, x17962x, x17966x, x17967x}, n_n3456);
	defparam lut_1307.LUT_SIZE = 7;
	defparam lut_1307.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_1314 ({sk[262], n_n5144, n_n31, x172x, x125x, x17922x, x17923x}, x18145x);
	defparam lut_1314.LUT_SIZE = 7;
	defparam lut_1314.mask = 128'h55ff55ff55ff55ff00007fffffffffff;

	lut_sub lut_1320 ({sk[263], n_n156, n_n4, n_n5, x717x, n_n3, n_n2}, x3622x);
	defparam lut_1320.LUT_SIZE = 7;
	defparam lut_1320.mask = 128'h55ff55ff55ff55ff00000000070f0f0f;

	lut_sub lut_1325 ({sk[264], i_9_, i_10_, i_11_, x717x}, x253x);
	defparam lut_1325.LUT_SIZE = 5;
	defparam lut_1325.mask = 32'h1f1f0440;

	lut_sub lut_1328 ({sk[265], i_7_, i_8_, i_6_, n_n159, n_n111}, x1550x);
	defparam lut_1328.LUT_SIZE = 6;
	defparam lut_1328.mask = 64'h11ffffff11000000;

	lut_sub lut_1331 ({sk[266], i_7_, i_6_, x741x, x744x, n_n7255, x18164x}, x18165x);
	defparam lut_1331.LUT_SIZE = 7;
	defparam lut_1331.mask = 128'h55ff55ff55ff55ff7f7f77777fff7777;

	lut_sub lut_1337 ({sk[267], i_14_, i_13_, i_12_, i_15_, n_n149}, x127x);
	defparam lut_1337.LUT_SIZE = 6;
	defparam lut_1337.mask = 64'h11ffffff00004044;

	lut_sub lut_1341 ({sk[268], i_14_, i_13_, i_12_, i_15_, n_n149, n_n170}, x1850x);
	defparam lut_1341.LUT_SIZE = 7;
	defparam lut_1341.mask = 128'h55ff55ff55ff55ff0050505003030300;

	lut_sub lut_1348 ({sk[269], x734x, n_n200, x172x, x133x, x158x, x147x}, x3442x);
	defparam lut_1348.LUT_SIZE = 7;
	defparam lut_1348.mask = 128'h55ff55ff55ff55ff0000000000007fff;

	lut_sub lut_1353 ({sk[270], i_15_, n_n32, x1417x, x18300x, n_n184, n_n201}, x18309x);
	defparam lut_1353.LUT_SIZE = 7;
	defparam lut_1353.mask = 128'h55ff55ff55ff55ff0f0f0fff0f0f1fff;

	lut_sub lut_1357 ({sk[271], n_n5144, n_n33, n_n32, x124x, x1858x, n_n138}, x18310x);
	defparam lut_1357.LUT_SIZE = 7;
	defparam lut_1357.mask = 128'h55ff55ff55ff55ff000f777fffffffff;

	lut_sub lut_1362 ({sk[272], i_7_, i_8_, i_6_, n_n162, n_n159}, n_n9);
	defparam lut_1362.LUT_SIZE = 6;
	defparam lut_1362.mask = 64'h11ffffff01000000;

	lut_sub lut_1364 ({sk[273], n_n9, n_n144, n_n186, n_n10, x145x, x170x}, n_n3378);
	defparam lut_1364.LUT_SIZE = 7;
	defparam lut_1364.mask = 128'h55ff55ff55ff55ff050f0f0f77ff7fff;

	lut_sub lut_1371 ({sk[274], i_7_, i_6_, i_1_, i_2_, i_0_, n_n162}, x388x);
	defparam lut_1371.LUT_SIZE = 7;
	defparam lut_1371.mask = 128'h55ff55ff55ff55ff1000100010000000;

	lut_sub lut_1375 ({sk[275], i_9_, i_10_, i_11_, x717x}, n_n151);
	defparam lut_1375.LUT_SIZE = 5;
	defparam lut_1375.mask = 32'h1f1f0004;

	lut_sub lut_1377 ({sk[276], x740x, n_n200, x714x, x17002x, x122x, x1865x}, x608x);
	defparam lut_1377.LUT_SIZE = 7;
	defparam lut_1377.mask = 128'h55ff55ff55ff55ff0003000300035557;

	lut_sub lut_1380 ({sk[277], n_n5056, n_n5060, x461x, x4906x, x4902x, x4903x}, x18361x);
	defparam lut_1380.LUT_SIZE = 7;
	defparam lut_1380.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_1387 ({sk[278], i_7_, i_8_, i_6_, x750x, x1429x, x18364x}, n_n3177);
	defparam lut_1387.LUT_SIZE = 7;
	defparam lut_1387.mask = 128'h55ff55ff55ff55ff5757555555555555;

	lut_sub lut_1391 ({sk[279], n_n65, x77x, n_n7346, n_n3, n_n5319, x18368x}, n_n3176);
	defparam lut_1391.LUT_SIZE = 7;
	defparam lut_1391.mask = 128'h55ff55ff55ff55ff77ff7fff7fff7fff;

	lut_sub lut_1397 ({sk[280], x245x, n_n5055, x714x, x17002x, x150x}, x18360x);
	defparam lut_1397.LUT_SIZE = 6;
	defparam lut_1397.mask = 64'h11ffffff01ff03ff;

	lut_sub lut_1401 ({sk[281], x428x, n_n14, x387x, x270x, x423x, x18373x}, x18376x);
	defparam lut_1401.LUT_SIZE = 7;
	defparam lut_1401.mask = 128'h55ff55ff55ff55ff77ff7fffffffffff;

	lut_sub lut_1407 ({sk[282], x18393x, x18397x, x18398x, x18401x, x21367x}, n_n3173);
	defparam lut_1407.LUT_SIZE = 6;
	defparam lut_1407.mask = 64'h11ffffffbfffffff;

	lut_sub lut_1413 ({sk[283], n_n3195, n_n3257, x18413x, x18414x, x18420x}, n_n3175);
	defparam lut_1413.LUT_SIZE = 6;
	defparam lut_1413.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1419 ({sk[284], x714x, x17051x, n_n3194, n_n3192, x1221x, x18433x}, x18436x);
	defparam lut_1419.LUT_SIZE = 7;
	defparam lut_1419.mask = 128'h55ff55ff55ff55ff5fff5fff5fff7fff;

	lut_sub lut_1424 ({sk[285], x18455x, x18456x, x18461x, x18462x, x18469x}, n_n3170);
	defparam lut_1424.LUT_SIZE = 6;
	defparam lut_1424.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1430 ({sk[286], x18475x, x18476x, n_n3186, x18486x}, n_n3172);
	defparam lut_1430.LUT_SIZE = 5;
	defparam lut_1430.mask = 32'h1f1f7fff;

	lut_sub lut_1435 ({sk[287], i_3_, i_1_, i_2_, i_0_, n_n3184, x21366x}, x18488x);
	defparam lut_1435.LUT_SIZE = 7;
	defparam lut_1435.mask = 128'h55ff55ff55ff55ffbbfbbbfbfbfbbbfb;

	lut_sub lut_1440 ({sk[288], i_8_, i_5_, i_3_, i_4_, n_n159, n_n157}, n_n2);
	defparam lut_1440.LUT_SIZE = 7;
	defparam lut_1440.mask = 128'h55ff55ff55ff55ff0100000000000000;

	lut_sub lut_1442 ({sk[289], i_9_, i_10_, i_11_}, n_n191);
	defparam lut_1442.LUT_SIZE = 4;
	defparam lut_1442.mask = 16'h5508;

	lut_sub lut_1444 ({sk[290], i_14_, i_13_, i_12_, i_15_, n_n191}, x87x);
	defparam lut_1444.LUT_SIZE = 6;
	defparam lut_1444.mask = 64'h11ffffff10004000;

	lut_sub lut_1447 ({sk[291], n_n5144, n_n149, x717x, n_n7346, n_n3, x708x}, x18511x);
	defparam lut_1447.LUT_SIZE = 7;
	defparam lut_1447.mask = 128'h55ff55ff55ff55ff5f5f5f7fffffffff;

	lut_sub lut_1452 ({sk[292], x181x, n_n197, n_n212, x151x, x1572x, x1224x}, n_n4441);
	defparam lut_1452.LUT_SIZE = 7;
	defparam lut_1452.mask = 128'h55ff55ff55ff55ff003f557f00ff55ff;

	lut_sub lut_1457 ({sk[293], n_n197, n_n212, x168x, x47x, x1855x, x1854x}, x575x);
	defparam lut_1457.LUT_SIZE = 7;
	defparam lut_1457.mask = 128'h55ff55ff55ff55ff000055ff3f3f7fff;

	lut_sub lut_1462 ({sk[294], x181x, x735x, n_n200, n_n212, x48x, x1732x}, x18577x);
	defparam lut_1462.LUT_SIZE = 7;
	defparam lut_1462.mask = 128'h55ff55ff55ff55ff07070707070707ff;

	lut_sub lut_1466 ({sk[295], x735x, n_n200, n_n212, x63x, x1857x, x1602x}, x18578x);
	defparam lut_1466.LUT_SIZE = 7;
	defparam lut_1466.mask = 128'h55ff55ff55ff55ff003f003f003f557f;

	lut_sub lut_1470 ({sk[296], i_7_, i_8_, i_6_, x735x, x774x, x18620x}, x18621x);
	defparam lut_1470.LUT_SIZE = 7;
	defparam lut_1470.mask = 128'h55ff55ff55ff55ff5555555557555555;

	lut_sub lut_1473 ({sk[297], n_n74, n_n92, n_n3, n_n2, x815x, x3067x}, n_n3034);
	defparam lut_1473.LUT_SIZE = 7;
	defparam lut_1473.mask = 128'h55ff55ff55ff55ff55557fff7fff7fff;

	lut_sub lut_1481 ({sk[298], n_n41, x245x, n_n5055, n_n5056, n_n18, x732x}, x18712x);
	defparam lut_1481.LUT_SIZE = 7;
	defparam lut_1481.mask = 128'h55ff55ff55ff55ff1fff1fff1fffffff;

	lut_sub lut_1486 ({sk[299], x387x, n_n132, x714x, x17002x, x150x, x4902x}, x18711x);
	defparam lut_1486.LUT_SIZE = 7;
	defparam lut_1486.mask = 128'h55ff55ff55ff55ff5557555fffffffff;

	lut_sub lut_1491 ({sk[300], n_n9, n_n74, n_n68, n_n10, n_n92, x18715x}, x18716x);
	defparam lut_1491.LUT_SIZE = 7;
	defparam lut_1491.mask = 128'h55ff55ff55ff55ff575f575f77ffffff;

	lut_sub lut_1498 ({sk[301], x18701x, x18702x, n_n3054}, x18717x);
	defparam lut_1498.LUT_SIZE = 4;
	defparam lut_1498.mask = 16'h557f;

	lut_sub lut_1502 ({sk[302], n_n31, x18749x, x865x, x18755x, x21365x}, n_n4849);
	defparam lut_1502.LUT_SIZE = 6;
	defparam lut_1502.mask = 64'h11ffffffbbffbfff;

	lut_sub lut_1507 ({sk[303], x18761x, x18762x, x18766x, x18767x, x18768x}, n_n4850);
	defparam lut_1507.LUT_SIZE = 6;
	defparam lut_1507.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1513 ({sk[304], x729x, n_n156, x387x, n_n3, n_n2, n_n12}, x18814x);
	defparam lut_1513.LUT_SIZE = 7;
	defparam lut_1513.mask = 128'h55ff55ff55ff55ff00ff00ff00ff7fff;

	lut_sub lut_1518 ({sk[305], n_n71, n_n4, n_n5319, x95x, x786x, x21364x}, x18815x);
	defparam lut_1518.LUT_SIZE = 7;
	defparam lut_1518.mask = 128'h55ff55ff55ff55ff0aff0aff3bffffff;

	lut_sub lut_1523 ({sk[306], i_7_, i_5_, i_6_, x286x, n_n2, x95x}, x18816x);
	defparam lut_1523.LUT_SIZE = 7;
	defparam lut_1523.mask = 128'h55ff55ff55ff55ff11111f1111111111;

	lut_sub lut_1526 ({sk[307], n_n30, n_n356, x1916x, x19878x, x1567x, x1908x}, x19893x);
	defparam lut_1526.LUT_SIZE = 7;
	defparam lut_1526.mask = 128'h55ff55ff55ff55ff5fffffff7fffffff;

	lut_sub lut_1532 ({sk[308], n_n31, x516x, x19898x, n_n310, x1592x, x19907x}, n_n296);
	defparam lut_1532.LUT_SIZE = 7;
	defparam lut_1532.mask = 128'h55ff55ff55ff55ff5fffffff7fffffff;

	lut_sub lut_1538 ({sk[309], i_9_, i_10_, i_11_, n_n36, n_n34, x728x}, n_n360);
	defparam lut_1538.LUT_SIZE = 7;
	defparam lut_1538.mask = 128'h55ff55ff55ff55ff1511001515050011;

	lut_sub lut_1548 ({sk[310], n_n149, n_n36, n_n34, x720x, x127x, x1780x}, n_n362);
	defparam lut_1548.LUT_SIZE = 7;
	defparam lut_1548.mask = 128'h55ff55ff55ff55ff0077337700773f7f;

	lut_sub lut_1553 ({sk[311], n_n149, n_n36, x726x, x718x, n_n64, x19889x}, x19890x);
	defparam lut_1553.LUT_SIZE = 7;
	defparam lut_1553.mask = 128'h55ff55ff55ff55ff5555777755557fff;

	lut_sub lut_1558 ({sk[312], n_n5144, x185x, n_n7346, n_n3, x19697x, x19698x}, x19912x);
	defparam lut_1558.LUT_SIZE = 7;
	defparam lut_1558.mask = 128'h55ff55ff55ff55ff77ff7fffffffffff;

	lut_sub lut_1564 ({sk[313], n_n149, n_n5, x717x, n_n191, x18317x, x170x}, n_n259);
	defparam lut_1564.LUT_SIZE = 7;
	defparam lut_1564.mask = 128'h55ff55ff55ff55ff3333777f333377ff;

	lut_sub lut_1569 ({sk[314], i_7_, i_6_, x733x, x288x, n_n7252, x732x}, x18322x);
	defparam lut_1569.LUT_SIZE = 7;
	defparam lut_1569.mask = 128'h55ff55ff55ff55ff77ff77ff7fff77ff;

	lut_sub lut_1580 ({sk[315], i_14_, i_13_, i_12_, i_15_, n_n156}, x372x);
	defparam lut_1580.LUT_SIZE = 6;
	defparam lut_1580.mask = 64'h11ffffff10404000;

	lut_sub lut_1584 ({sk[316], n_n5144, x77x, n_n7346, n_n3, x707x}, x19945x);
	defparam lut_1584.LUT_SIZE = 6;
	defparam lut_1584.mask = 64'h11ffffff5f7fffff;

	lut_sub lut_1589 ({sk[317], i_7_, i_6_, i_1_, i_2_, i_0_, n_n162}, n_n7252);
	defparam lut_1589.LUT_SIZE = 7;
	defparam lut_1589.mask = 128'h55ff55ff55ff55ff0000000000001000;

	lut_sub lut_1591 ({sk[318], i_7_, i_5_, i_6_, i_3_, i_4_, n_n219}, x567x);
	defparam lut_1591.LUT_SIZE = 7;
	defparam lut_1591.mask = 128'h55ff55ff55ff55ff0000100000100000;

	lut_sub lut_1594 ({sk[319], i_7_, i_6_, i_1_, i_2_, i_0_, n_n48}, n_n7262);
	defparam lut_1594.LUT_SIZE = 7;
	defparam lut_1594.mask = 128'h55ff55ff55ff55ff0000100000000000;

	lut_sub lut_1596 ({sk[320], i_1_, i_2_, i_0_}, n_n219);
	defparam lut_1596.LUT_SIZE = 4;
	defparam lut_1596.mask = 16'h5540;

	lut_sub lut_1598 ({sk[321], i_7_, i_5_, i_6_, i_3_, i_4_, n_n219}, x711x);
	defparam lut_1598.LUT_SIZE = 7;
	defparam lut_1598.mask = 128'h55ff55ff55ff55ff1010000000000000;

	lut_sub lut_1601 ({sk[322], i_9_, i_10_, i_11_}, n_n156);
	defparam lut_1601.LUT_SIZE = 4;
	defparam lut_1601.mask = 16'h5502;

	lut_sub lut_1603 ({sk[323], i_5_, i_3_, i_4_}, n_n111);
	defparam lut_1603.LUT_SIZE = 4;
	defparam lut_1603.mask = 16'h5580;

	lut_sub lut_1605 ({sk[324], i_5_, i_3_, i_4_}, n_n48);
	defparam lut_1605.LUT_SIZE = 4;
	defparam lut_1605.mask = 16'h5504;

	lut_sub lut_1607 ({sk[325], i_7_, i_8_, i_6_}, n_n124);
	defparam lut_1607.LUT_SIZE = 4;
	defparam lut_1607.mask = 16'h5540;

	lut_sub lut_1609 ({sk[326], i_7_, i_8_, i_6_, x740x}, n_n38);
	defparam lut_1609.LUT_SIZE = 5;
	defparam lut_1609.mask = 32'h1f1f1000;

	lut_sub lut_1611 ({sk[327], i_7_, i_8_, i_6_, x740x}, n_n39);
	defparam lut_1611.LUT_SIZE = 5;
	defparam lut_1611.mask = 32'h1f1f0100;

	lut_sub lut_1613 ({sk[328], i_14_, i_13_, i_12_}, n_n209);
	defparam lut_1613.LUT_SIZE = 4;
	defparam lut_1613.mask = 16'h5501;

	lut_sub lut_1615 ({sk[329], i_9_, i_10_, i_11_, i_15_, n_n209}, n_n134);
	defparam lut_1615.LUT_SIZE = 6;
	defparam lut_1615.mask = 64'h11ffffff00000100;

	lut_sub lut_1617 ({sk[330], i_7_, i_8_, i_6_}, n_n126);
	defparam lut_1617.LUT_SIZE = 4;
	defparam lut_1617.mask = 16'h5510;

	lut_sub lut_1619 ({sk[331], i_9_, i_10_, i_11_}, n_n177);
	defparam lut_1619.LUT_SIZE = 4;
	defparam lut_1619.mask = 16'h5504;

	lut_sub lut_1621 ({sk[332], i_15_, x740x, n_n126, n_n177, n_n209}, n_n6642);
	defparam lut_1621.LUT_SIZE = 6;
	defparam lut_1621.mask = 64'h11ffffff00000001;

	lut_sub lut_1623 ({sk[333], i_14_, i_13_, i_12_, i_15_, n_n149}, x235x);
	defparam lut_1623.LUT_SIZE = 6;
	defparam lut_1623.mask = 64'h11ffffff05004000;

	lut_sub lut_1627 ({sk[334], i_14_, i_13_, i_12_, i_15_, n_n149}, x236x);
	defparam lut_1627.LUT_SIZE = 6;
	defparam lut_1627.mask = 64'h11ffffff00000144;

	lut_sub lut_1631 ({sk[335], i_14_, i_13_, i_12_, i_15_, n_n156}, x140x);
	defparam lut_1631.LUT_SIZE = 6;
	defparam lut_1631.mask = 64'h11ffffff05004000;

	lut_sub lut_1635 ({sk[336], i_14_, i_13_, i_12_, i_15_, n_n170}, n_n132);
	defparam lut_1635.LUT_SIZE = 6;
	defparam lut_1635.mask = 64'h11ffffff00000001;

	lut_sub lut_1637 ({sk[337], i_7_, i_8_, i_6_, x740x, n_n6642, n_n132}, n_n969);
	defparam lut_1637.LUT_SIZE = 7;
	defparam lut_1637.mask = 128'h55ff55ff55ff55ff3337333733333333;

	lut_sub lut_1641 ({sk[338], i_14_, i_13_, i_12_, i_15_}, x728x);
	defparam lut_1641.LUT_SIZE = 5;
	defparam lut_1641.mask = 32'h1f1f0020;

	lut_sub lut_1643 ({sk[339], i_9_, i_10_, i_11_, x740x, n_n126, x728x}, n_n6646);
	defparam lut_1643.LUT_SIZE = 7;
	defparam lut_1643.mask = 128'h55ff55ff55ff55ff0000000000000100;

	lut_sub lut_1645 ({sk[340], i_9_, i_10_, i_11_, x728x}, n_n52);
	defparam lut_1645.LUT_SIZE = 5;
	defparam lut_1645.mask = 32'h1f1f0400;

	lut_sub lut_1647 ({sk[341], i_7_, i_8_, i_6_, x740x, n_n6646, n_n52}, n_n519);
	defparam lut_1647.LUT_SIZE = 7;
	defparam lut_1647.mask = 128'h55ff55ff55ff55ff3337333733333333;

	lut_sub lut_1651 ({sk[342], i_14_, i_13_, i_12_, i_15_}, x719x);
	defparam lut_1651.LUT_SIZE = 5;
	defparam lut_1651.mask = 32'h1f1f0001;

	lut_sub lut_1653 ({sk[343], i_7_, i_8_, i_6_, x740x, n_n177, x719x}, x393x);
	defparam lut_1653.LUT_SIZE = 7;
	defparam lut_1653.mask = 128'h55ff55ff55ff55ff0001000000000000;

	lut_sub lut_1655 ({sk[344], i_7_, i_8_, i_6_, x740x, n_n134, n_n132}, n_n4597);
	defparam lut_1655.LUT_SIZE = 7;
	defparam lut_1655.mask = 128'h55ff55ff55ff55ff0007000500000000;

	lut_sub lut_1659 ({sk[345], i_14_, i_13_, i_12_, i_15_}, x730x);
	defparam lut_1659.LUT_SIZE = 5;
	defparam lut_1659.mask = 32'h1f1f0080;

	lut_sub lut_1661 ({sk[346], i_9_, i_10_, i_11_, x730x}, n_n74);
	defparam lut_1661.LUT_SIZE = 5;
	defparam lut_1661.mask = 32'h1f1f0004;

	lut_sub lut_1663 ({sk[347], i_7_, i_8_, i_6_, x740x, n_n6646, n_n52}, x390x);
	defparam lut_1663.LUT_SIZE = 7;
	defparam lut_1663.mask = 128'h55ff55ff55ff55ff3337333333333333;

	lut_sub lut_1666 ({sk[348], i_7_, i_8_, i_6_, n_n156, x740x, x728x}, x392x);
	defparam lut_1666.LUT_SIZE = 7;
	defparam lut_1666.mask = 128'h55ff55ff55ff55ff0001000000000000;

	lut_sub lut_1668 ({sk[349], n_n149, n_n156, n_n124, x740x, n_n126, x728x}, x712x);
	defparam lut_1668.LUT_SIZE = 7;
	defparam lut_1668.mask = 128'h55ff55ff55ff55ff0000000501010105;

	lut_sub lut_1671 ({sk[350], i_8_, i_1_, i_2_, i_0_}, x714x);
	defparam lut_1671.LUT_SIZE = 5;
	defparam lut_1671.mask = 32'h1f1f0080;

	lut_sub lut_1673 ({sk[351], i_7_, i_5_, i_6_, i_3_, i_4_, x714x}, n_n31);
	defparam lut_1673.LUT_SIZE = 7;
	defparam lut_1673.mask = 128'h55ff55ff55ff55ff0000400000000000;

	lut_sub lut_1675 ({sk[352], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x734x);
	defparam lut_1675.LUT_SIZE = 7;
	defparam lut_1675.mask = 128'h55ff55ff55ff55ff0000000080000000;

	lut_sub lut_1677 ({sk[353], i_7_, i_8_, i_6_, x734x}, n_n30);
	defparam lut_1677.LUT_SIZE = 5;
	defparam lut_1677.mask = 32'h1f1f4000;

	lut_sub lut_1679 ({sk[354], i_9_, i_10_, i_11_}, n_n216);
	defparam lut_1679.LUT_SIZE = 4;
	defparam lut_1679.mask = 16'h5501;

	lut_sub lut_1681 ({sk[355], i_14_, i_13_, i_12_, i_15_, n_n216}, x1449x);
	defparam lut_1681.LUT_SIZE = 6;
	defparam lut_1681.mask = 64'h11ffffff11015154;

	lut_sub lut_1691 ({sk[356], i_14_, i_13_, i_12_, i_15_, n_n216}, x181x);
	defparam lut_1691.LUT_SIZE = 6;
	defparam lut_1691.mask = 64'h11ffffff04440000;

	lut_sub lut_1695 ({sk[357], i_7_, i_8_, i_6_, x735x}, n_n34);
	defparam lut_1695.LUT_SIZE = 5;
	defparam lut_1695.mask = 32'h1f1f4000;

	lut_sub lut_1697 ({sk[358], i_14_, i_13_, i_12_, i_15_, n_n177}, x78x);
	defparam lut_1697.LUT_SIZE = 6;
	defparam lut_1697.mask = 64'h11ffffff40100000;

	lut_sub lut_1700 ({sk[359], i_14_, i_13_, i_12_, i_15_, n_n216}, x143x);
	defparam lut_1700.LUT_SIZE = 6;
	defparam lut_1700.mask = 64'h11ffffff11010000;

	lut_sub lut_1704 ({sk[360], i_14_, i_13_, i_12_, i_15_, n_n216}, x1825x);
	defparam lut_1704.LUT_SIZE = 6;
	defparam lut_1704.mask = 64'h11ffffff00005154;

	lut_sub lut_1711 ({sk[361], i_7_, i_8_, i_6_, x734x, x719x, n_n170}, x753x);
	defparam lut_1711.LUT_SIZE = 7;
	defparam lut_1711.mask = 128'h55ff55ff55ff55ff0000000001000000;

	lut_sub lut_1713 ({sk[362], n_n31, n_n34, x78x, x143x, x1825x, x753x}, x16943x);
	defparam lut_1713.LUT_SIZE = 7;
	defparam lut_1713.mask = 128'h55ff55ff55ff55ff555555ff7f7f7fff;

	lut_sub lut_1718 ({sk[363], i_14_, i_13_, i_12_, i_15_, n_n170}, x132x);
	defparam lut_1718.LUT_SIZE = 6;
	defparam lut_1718.mask = 64'h11ffffff00001110;

	lut_sub lut_1722 ({sk[364], i_7_, i_5_, i_6_, i_3_, i_4_, x714x}, n_n36);
	defparam lut_1722.LUT_SIZE = 7;
	defparam lut_1722.mask = 128'h55ff55ff55ff55ff1000000000000000;

	lut_sub lut_1724 ({sk[365], i_14_, i_13_, i_12_, i_15_, n_n170}, x126x);
	defparam lut_1724.LUT_SIZE = 6;
	defparam lut_1724.mask = 64'h11ffffff00004044;

	lut_sub lut_1728 ({sk[366], i_7_, i_8_, i_6_, x137x, x735x}, n_n4569);
	defparam lut_1728.LUT_SIZE = 6;
	defparam lut_1728.mask = 64'h11ffffff10000000;

	lut_sub lut_1730 ({sk[367], i_7_, i_8_, i_6_, x46x, x735x}, x4970x);
	defparam lut_1730.LUT_SIZE = 6;
	defparam lut_1730.mask = 64'h11ffffff10000000;

	lut_sub lut_1732 ({sk[368], n_n36, x125x, x149x, x147x, n_n4568, x4968x}, x16960x);
	defparam lut_1732.LUT_SIZE = 7;
	defparam lut_1732.mask = 128'h55ff55ff55ff55ff777777777fffffff;

	lut_sub lut_1738 ({sk[369], n_n36, n_n34, n_n140, x247x, x709x, x153x}, n_n4169);
	defparam lut_1738.LUT_SIZE = 7;
	defparam lut_1738.mask = 128'h55ff55ff55ff55ff333377773fff7fff;

	lut_sub lut_1743 ({sk[370], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x942x);
	defparam lut_1743.LUT_SIZE = 7;
	defparam lut_1743.mask = 128'h55ff55ff55ff55ff7000070000700007;

	lut_sub lut_1752 ({sk[371], x725x, n_n34, x125x, n_n216, x941x}, x16950x);
	defparam lut_1752.LUT_SIZE = 6;
	defparam lut_1752.mask = 64'h11ffffff005f007f;

	lut_sub lut_1756 ({sk[372], x181x, x132x, n_n34, x149x, x147x}, x16955x);
	defparam lut_1756.LUT_SIZE = 6;
	defparam lut_1756.mask = 64'h11ffffff070f0f0f;

	lut_sub lut_1761 ({sk[373], x137x, x46x, n_n36, n_n34, x126x, x1877x}, x16956x);
	defparam lut_1761.LUT_SIZE = 7;
	defparam lut_1761.mask = 128'h55ff55ff55ff55ff035703ff03ff03ff;

	lut_sub lut_1766 ({sk[374], i_14_, i_13_, i_12_, i_15_, n_n177}, x137x);
	defparam lut_1766.LUT_SIZE = 6;
	defparam lut_1766.mask = 64'h11ffffff00004044;

	lut_sub lut_1770 ({sk[375], i_14_, i_13_, i_12_, i_15_, n_n177}, x46x);
	defparam lut_1770.LUT_SIZE = 6;
	defparam lut_1770.mask = 64'h11ffffff00001110;

	lut_sub lut_1774 ({sk[376], i_14_, i_13_, i_12_, i_15_, n_n170}, x149x);
	defparam lut_1774.LUT_SIZE = 6;
	defparam lut_1774.mask = 64'h11ffffff04440000;

	lut_sub lut_1778 ({sk[377], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1806x);
	defparam lut_1778.LUT_SIZE = 7;
	defparam lut_1778.mask = 128'h55ff55ff55ff55ff7555575550705053;

	lut_sub lut_1795 ({sk[378], n_n31, n_n30, x137x, x46x, x149x, x1806x}, x16975x);
	defparam lut_1795.LUT_SIZE = 7;
	defparam lut_1795.mask = 128'h55ff55ff55ff55ff00005fff33337fff;

	lut_sub lut_1800 ({sk[379], n_n31, n_n30, n_n63, x135x, x153x, x1371x}, n_n4154);
	defparam lut_1800.LUT_SIZE = 7;
	defparam lut_1800.mask = 128'h55ff55ff55ff55ff00003f3f55ff7fff;

	lut_sub lut_1805 ({sk[380], n_n31, n_n30, x125x, x80x, x78x, x131x}, x16967x);
	defparam lut_1805.LUT_SIZE = 7;
	defparam lut_1805.mask = 128'h55ff55ff55ff55ff000055553fff7fff;

	lut_sub lut_1810 ({sk[381], n_n30, x719x, n_n63, x125x, x146x, n_n170}, x4961x);
	defparam lut_1810.LUT_SIZE = 7;
	defparam lut_1810.mask = 128'h55ff55ff55ff55ff000000003fff7fff;

	lut_sub lut_1815 ({sk[382], i_14_, i_13_, i_12_, i_15_, n_n31, n_n170}, x16974x);
	defparam lut_1815.LUT_SIZE = 7;
	defparam lut_1815.mask = 128'h55ff55ff55ff55ff1101010111111111;

	lut_sub lut_1829 ({sk[383], n_n46, x70x, n_n47, n_n214, x1841x, x1840x}, x543x);
	defparam lut_1829.LUT_SIZE = 7;
	defparam lut_1829.mask = 128'h55ff55ff55ff55ff005500ff3f7f3fff;

	lut_sub lut_1834 ({sk[384], x16993x, x16994x, x16997x, x16998x, x16999x}, n_n4408);
	defparam lut_1834.LUT_SIZE = 6;
	defparam lut_1834.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1840 ({sk[385], n_n46, n_n47, x180x, x142x, n_n169, x57x}, x17093x);
	defparam lut_1840.LUT_SIZE = 7;
	defparam lut_1840.mask = 128'h55ff55ff55ff55ff000055553fff7fff;

	lut_sub lut_1845 ({sk[386], n_n101, n_n108, x618x, x225x, x148x, x17153x}, x17155x);
	defparam lut_1845.LUT_SIZE = 7;
	defparam lut_1845.mask = 128'h55ff55ff55ff55ff55ff5fff7fff7fff;

	lut_sub lut_1851 ({sk[387], n_n4206, x17070x, x17071x, x17077x, x17078x}, x17156x);
	defparam lut_1851.LUT_SIZE = 6;
	defparam lut_1851.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1857 ({sk[388], n_n46, n_n47, x1031x, x1030x, x1170x, x1169x}, x21405x);
	defparam lut_1857.LUT_SIZE = 7;
	defparam lut_1857.mask = 128'h55ff55ff55ff55ffffffc0c0aa008000;

	lut_sub lut_1862 ({sk[389], i_9_, i_10_, i_11_}, n_n170);
	defparam lut_1862.LUT_SIZE = 4;
	defparam lut_1862.mask = 16'h5540;

	lut_sub lut_1864 ({sk[390], i_14_, i_13_, i_12_, i_15_, n_n170}, x53x);
	defparam lut_1864.LUT_SIZE = 6;
	defparam lut_1864.mask = 64'h11ffffff00000110;

	lut_sub lut_1867 ({sk[391], i_14_, i_13_, i_12_}, n_n211);
	defparam lut_1867.LUT_SIZE = 4;
	defparam lut_1867.mask = 16'h5508;

	lut_sub lut_1869 ({sk[392], i_9_, i_10_, i_11_, i_15_, n_n211}, n_n168);
	defparam lut_1869.LUT_SIZE = 6;
	defparam lut_1869.mask = 64'h11ffffff01000000;

	lut_sub lut_1871 ({sk[393], i_14_, i_13_, i_12_, i_15_, n_n199}, x151x);
	defparam lut_1871.LUT_SIZE = 6;
	defparam lut_1871.mask = 64'h11ffffff00001110;

	lut_sub lut_1875 ({sk[394], i_14_, i_13_, i_12_, i_15_, n_n199}, x1108x);
	defparam lut_1875.LUT_SIZE = 6;
	defparam lut_1875.mask = 64'h11ffffff15454044;

	lut_sub lut_1885 ({sk[395], i_14_, i_13_, i_12_, i_15_, n_n199}, x1864x);
	defparam lut_1885.LUT_SIZE = 6;
	defparam lut_1885.mask = 64'h11ffffff15455154;

	lut_sub lut_1898 ({sk[396], n_n31, n_n30, x181x, x151x, x1108x, x1864x}, x599x);
	defparam lut_1898.LUT_SIZE = 7;
	defparam lut_1898.mask = 128'h55ff55ff55ff55ff000055553fff7fff;

	lut_sub lut_1903 ({sk[397], i_14_, i_13_, i_12_, i_15_, n_n177}, x1899x);
	defparam lut_1903.LUT_SIZE = 6;
	defparam lut_1903.mask = 64'h11ffffff15450000;

	lut_sub lut_1910 ({sk[398], i_7_, i_6_}, n_n17);
	defparam lut_1910.LUT_SIZE = 3;
	defparam lut_1910.mask = 8'h52;

	lut_sub lut_1912 ({sk[399], i_3_, i_4_, i_1_, i_2_, i_0_}, x286x);
	defparam lut_1912.LUT_SIZE = 6;
	defparam lut_1912.mask = 64'h11ffffff00000008;

	lut_sub lut_1914 ({sk[400], i_7_, i_8_, i_6_, x740x}, n_n46);
	defparam lut_1914.LUT_SIZE = 5;
	defparam lut_1914.mask = 32'h1f1f0010;

	lut_sub lut_1916 ({sk[401], i_14_, i_13_, i_12_, i_15_, n_n199}, x168x);
	defparam lut_1916.LUT_SIZE = 6;
	defparam lut_1916.mask = 64'h11ffffff04440000;

	lut_sub lut_1920 ({sk[402], i_8_, i_1_, i_2_, i_0_, x17051x}, n_n47);
	defparam lut_1920.LUT_SIZE = 6;
	defparam lut_1920.mask = 64'h11ffffff00004000;

	lut_sub lut_1922 ({sk[403], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x830x);
	defparam lut_1922.LUT_SIZE = 7;
	defparam lut_1922.mask = 128'h55ff55ff55ff55ff0700000077000000;

	lut_sub lut_1929 ({sk[404], i_9_, i_10_, i_11_, x725x, n_n101, n_n108}, x17187x);
	defparam lut_1929.LUT_SIZE = 7;
	defparam lut_1929.mask = 128'h55ff55ff55ff55ff0000070000000300;

	lut_sub lut_1933 ({sk[405], x181x, n_n46, x168x, n_n47, x830x, x17187x}, x17192x);
	defparam lut_1933.LUT_SIZE = 7;
	defparam lut_1933.mask = 128'h55ff55ff55ff55ff575f77ff5f5fffff;

	lut_sub lut_1941 ({sk[406], x729x, n_n42, n_n43, n_n191, x93x, x967x}, n_n2312);
	defparam lut_1941.LUT_SIZE = 7;
	defparam lut_1941.mask = 128'h55ff55ff55ff55ff00335577003f557f;

	lut_sub lut_1945 ({sk[407], n_n51, n_n43, n_n55, x189x, x611x, x895x}, x17205x);
	defparam lut_1945.LUT_SIZE = 7;
	defparam lut_1945.mask = 128'h55ff55ff55ff55ff333f777f3f3f7f7f;

	lut_sub lut_1950 ({sk[408], x512x, n_n42, n_n43, n_n117, x609x, x301x}, x17204x);
	defparam lut_1950.LUT_SIZE = 7;
	defparam lut_1950.mask = 128'h55ff55ff55ff55ff337f7f7fffffffff;

	lut_sub lut_1957 ({sk[409], x740x, n_n161, n_n47, x176x, x149x, x131x}, x17210x);
	defparam lut_1957.LUT_SIZE = 7;
	defparam lut_1957.mask = 128'h55ff55ff55ff55ff003f003f003f557f;

	lut_sub lut_1961 ({sk[410], n_n46, n_n47, x149x, x200x, x201x, x17208x}, x17211x);
	defparam lut_1961.LUT_SIZE = 7;
	defparam lut_1961.mask = 128'h55ff55ff55ff55ff000077773fff7fff;

	lut_sub lut_1967 ({sk[411], n_n2312, x17205x, x17204x, x17210x, x17211x}, x17213x);
	defparam lut_1967.LUT_SIZE = 6;
	defparam lut_1967.mask = 64'h11ffffff7fffffff;

	lut_sub lut_1973 ({sk[412], n_n135, n_n31, x181x, n_n33, n_n32, x969x}, x17218x);
	defparam lut_1973.LUT_SIZE = 7;
	defparam lut_1973.mask = 128'h55ff55ff55ff55ff050505ff373737ff;

	lut_sub lut_1977 ({sk[413], x729x, n_n32, n_n184, x726x, x202x, x21398x}, x17228x);
	defparam lut_1977.LUT_SIZE = 7;
	defparam lut_1977.mask = 128'h55ff55ff55ff55ffaaaabbbfaaaabbff;

	lut_sub lut_1982 ({sk[414], n_n33, x60x, x307x, x1054x, x17225x, x4656x}, x17229x);
	defparam lut_1982.LUT_SIZE = 7;
	defparam lut_1982.mask = 128'h55ff55ff55ff55ff555555557fffffff;

	lut_sub lut_1988 ({sk[415], n_n31, n_n30, x181x, x129x, x900x, x970x}, x21397x);
	defparam lut_1988.LUT_SIZE = 7;
	defparam lut_1988.mask = 128'h55ff55ff55ff55ff00007fff7f7f7fff;

	lut_sub lut_2005 ({sk[416], n_n135, n_n30, n_n63, x176x, x299x, x17237x}, x4639x);
	defparam lut_2005.LUT_SIZE = 7;
	defparam lut_2005.mask = 128'h55ff55ff55ff55ff00007fff0000ffff;

	lut_sub lut_2011 ({sk[417], n_n31, n_n63, x158x, x299x, x17235x, x4640x}, x17241x);
	defparam lut_2011.LUT_SIZE = 7;
	defparam lut_2011.mask = 128'h55ff55ff55ff55ff555555557fffffff;

	lut_sub lut_2017 ({sk[418], i_9_, i_10_, i_11_, n_n31, n_n30, x725x}, n_n2235);
	defparam lut_2017.LUT_SIZE = 7;
	defparam lut_2017.mask = 128'h55ff55ff55ff55ff0515150011151500;

	lut_sub lut_2028 ({sk[419], i_8_, n_n157, n_n31, x734x, x149x, x131x}, x17245x);
	defparam lut_2028.LUT_SIZE = 7;
	defparam lut_2028.mask = 128'h55ff55ff55ff55ff0033053700330033;

	lut_sub lut_2031 ({sk[420], n_n31, n_n30, x149x, x200x, x201x, x17244x}, x17247x);
	defparam lut_2031.LUT_SIZE = 7;
	defparam lut_2031.mask = 128'h55ff55ff55ff55ff00003fff7f7f7fff;

	lut_sub lut_2038 ({sk[421], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x735x);
	defparam lut_2038.LUT_SIZE = 7;
	defparam lut_2038.mask = 128'h55ff55ff55ff55ff0080000000000000;

	lut_sub lut_2040 ({sk[422], i_9_, i_10_, i_11_, x729x}, n_n77);
	defparam lut_2040.LUT_SIZE = 5;
	defparam lut_2040.mask = 32'h1f1f1000;

	lut_sub lut_2042 ({sk[423], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x974x);
	defparam lut_2042.LUT_SIZE = 7;
	defparam lut_2042.mask = 128'h55ff55ff55ff55ff0550005077000000;

	lut_sub lut_2050 ({sk[424], n_n123, n_n125, n_n83, x975x, x1234x, x120x}, x17276x);
	defparam lut_2050.LUT_SIZE = 7;
	defparam lut_2050.mask = 128'h55ff55ff55ff55ff00003f3f55ff7fff;

	lut_sub lut_2055 ({sk[425], i_8_, n_n16, x735x, n_n77, x974x, x17276x}, x17277x);
	defparam lut_2055.LUT_SIZE = 7;
	defparam lut_2055.mask = 128'h55ff55ff55ff55ff5555557f55555555;

	lut_sub lut_2059 ({sk[426], x735x, n_n161, x62x, n_n113, x885x, x202x}, n_n2339);
	defparam lut_2059.LUT_SIZE = 7;
	defparam lut_2059.mask = 128'h55ff55ff55ff55ff050f050f050f373f;

	lut_sub lut_2063 ({sk[427], x729x, n_n156, x735x, n_n126, x972x}, x17256x);
	defparam lut_2063.LUT_SIZE = 6;
	defparam lut_2063.mask = 64'h11ffffff01010103;

	lut_sub lut_2066 ({sk[428], n_n135, n_n71, n_n123, n_n125, x971x, x1177x}, x17257x);
	defparam lut_2066.LUT_SIZE = 7;
	defparam lut_2066.mask = 128'h55ff55ff55ff55ff057705ff0fff0fff;

	lut_sub lut_2073 ({sk[429], x725x, n_n170, n_n113, x255x, n_n182, x21394x}, n_n2340);
	defparam lut_2073.LUT_SIZE = 7;
	defparam lut_2073.mask = 128'h55ff55ff55ff55ff5577557755775f7f;

	lut_sub lut_2077 ({sk[430], x734x, n_n126, n_n210, x21392x, x21456x}, x17268x);
	defparam lut_2077.LUT_SIZE = 6;
	defparam lut_2077.mask = 64'h11ffffffeeeeeeef;

	lut_sub lut_2081 ({sk[431], n_n2339, x17256x, x17257x, n_n2340, x17268x}, x17278x);
	defparam lut_2081.LUT_SIZE = 6;
	defparam lut_2081.mask = 64'h11ffffff7fffffff;

	lut_sub lut_2087 ({sk[432], i_9_, i_10_, i_11_, x730x}, n_n92);
	defparam lut_2087.LUT_SIZE = 5;
	defparam lut_2087.mask = 32'h1f1f0040;

	lut_sub lut_2089 ({sk[433], i_9_, i_10_, i_11_, i_15_, n_n211}, n_n189);
	defparam lut_2089.LUT_SIZE = 6;
	defparam lut_2089.mask = 64'h11ffffff00001000;

	lut_sub lut_2091 ({sk[434], i_14_, i_13_, i_12_, i_15_, n_n199}, x360x);
	defparam lut_2091.LUT_SIZE = 6;
	defparam lut_2091.mask = 64'h11ffffff00005000;

	lut_sub lut_2094 ({sk[435], x729x, n_n36, n_n34, n_n199, x977x, x243x}, x17302x);
	defparam lut_2094.LUT_SIZE = 7;
	defparam lut_2094.mask = 128'h55ff55ff55ff55ff00775577007f5f7f;

	lut_sub lut_2100 ({sk[436], n_n36, n_n34, n_n102, x360x, x495x, x1275x}, x21430x);
	defparam lut_2100.LUT_SIZE = 7;
	defparam lut_2100.mask = 128'h55ff55ff55ff55ffccccc00088008000;

	lut_sub lut_2105 ({sk[437], n_n36, n_n92, n_n189, x360x, x17302x, x21430x}, x17304x);
	defparam lut_2105.LUT_SIZE = 7;
	defparam lut_2105.mask = 128'h55ff55ff55ff55ffbbbbbbbbbfffffff;

	lut_sub lut_2111 ({sk[438], n_n149, x725x, x190x, x17288x, x21390x, x21391x}, x17290x);
	defparam lut_2111.LUT_SIZE = 7;
	defparam lut_2111.mask = 128'h55ff55ff55ff55ffefefefefefefefff;

	lut_sub lut_2116 ({sk[439], n_n40, x714x, x17002x, n_n61, x351x, x17293x}, x17297x);
	defparam lut_2116.LUT_SIZE = 7;
	defparam lut_2116.mask = 128'h55ff55ff55ff55ff0000007f0f0f0f7f;

	lut_sub lut_2121 ({sk[440], n_n41, n_n40, x377x, x363x, x17296x, x21389x}, x17298x);
	defparam lut_2121.LUT_SIZE = 7;
	defparam lut_2121.mask = 128'h55ff55ff55ff55ff0f0fbfbf0fffbfff;

	lut_sub lut_2126 ({sk[441], i_9_, i_10_, i_11_, x725x, n_n41, n_n40}, n_n2298);
	defparam lut_2126.LUT_SIZE = 7;
	defparam lut_2126.mask = 128'h55ff55ff55ff55ff0707000007070300;

	lut_sub lut_2136 ({sk[442], n_n38, n_n74, n_n68, n_n84, n_n143, n_n175}, x4581x);
	defparam lut_2136.LUT_SIZE = 7;
	defparam lut_2136.mask = 128'h55ff55ff55ff55ff000000007fffffff;

	lut_sub lut_2142 ({sk[443], x17290x, x17297x, x17298x, n_n2298, x4581x}, x17305x);
	defparam lut_2142.LUT_SIZE = 6;
	defparam lut_2142.mask = 64'h11ffffff7fffffff;

	lut_sub lut_2148 ({sk[444], n_n135, n_n36, n_n34, x820x, n_n55, x17307x}, n_n2284);
	defparam lut_2148.LUT_SIZE = 7;
	defparam lut_2148.mask = 128'h55ff55ff55ff55ff55777f7f55ffffff;

	lut_sub lut_2155 ({sk[445], i_9_, i_10_, i_11_, x725x, n_n36, x821x}, x17314x);
	defparam lut_2155.LUT_SIZE = 7;
	defparam lut_2155.mask = 128'h55ff55ff55ff55ff1111111111111113;

	lut_sub lut_2158 ({sk[446], x729x, n_n36, n_n34, n_n184, x93x, x17318x}, x17321x);
	defparam lut_2158.LUT_SIZE = 7;
	defparam lut_2158.mask = 128'h55ff55ff55ff55ff0077007700770f7f;

	lut_sub lut_2162 ({sk[447], n_n89, n_n36, n_n34, x93x, x1235x, x1238x}, x17322x);
	defparam lut_2162.LUT_SIZE = 7;
	defparam lut_2162.mask = 128'h55ff55ff55ff55ff00335f7f0033ffff;

	lut_sub lut_2167 ({sk[448], x729x, n_n149, n_n156, n_n34, x17313x, x115x}, x4554x);
	defparam lut_2167.LUT_SIZE = 7;
	defparam lut_2167.mask = 128'h55ff55ff55ff55ff07070707070f0f0f;

	lut_sub lut_2172 ({sk[449], n_n2284, x17314x, x17321x, x17322x, x4554x}, x17328x);
	defparam lut_2172.LUT_SIZE = 6;
	defparam lut_2172.mask = 64'h11ffffff7fffffff;

	lut_sub lut_2178 ({sk[450], i_7_, i_8_, i_6_, x740x}, n_n40);
	defparam lut_2178.LUT_SIZE = 5;
	defparam lut_2178.mask = 32'h1f1f0040;

	lut_sub lut_2180 ({sk[451], i_7_, i_5_, i_6_, i_3_, i_4_}, x17002x);
	defparam lut_2180.LUT_SIZE = 6;
	defparam lut_2180.mask = 64'h11ffffff00000040;

	lut_sub lut_2182 ({sk[452], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x984x);
	defparam lut_2182.LUT_SIZE = 7;
	defparam lut_2182.mask = 128'h55ff55ff55ff55ff0700007077000000;

	lut_sub lut_2191 ({sk[453], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x983x);
	defparam lut_2191.LUT_SIZE = 7;
	defparam lut_2191.mask = 128'h55ff55ff55ff55ff0570705055000000;

	lut_sub lut_2200 ({sk[454], n_n41, n_n40, n_n154, x69x, x397x, x1337x}, x17345x);
	defparam lut_2200.LUT_SIZE = 7;
	defparam lut_2200.mask = 128'h55ff55ff55ff55ff333377773fff7fff;

	lut_sub lut_2205 ({sk[455], n_n41, n_n40, x263x, x361x, x1733x, x1794x}, x17342x);
	defparam lut_2205.LUT_SIZE = 7;
	defparam lut_2205.mask = 128'h55ff55ff55ff55ff0f0f5fff3f3f7fff;

	lut_sub lut_2210 ({sk[456], i_8_, x734x, x725x, n_n184, n_n18, x93x}, x4531x);
	defparam lut_2210.LUT_SIZE = 7;
	defparam lut_2210.mask = 128'h55ff55ff55ff55ff0000111300000000;

	lut_sub lut_2213 ({sk[457], n_n135, n_n89, n_n42, n_n59, n_n43, x632x}, x17331x);
	defparam lut_2213.LUT_SIZE = 7;
	defparam lut_2213.mask = 128'h55ff55ff55ff55ff575f57ff777f77ff;

	lut_sub lut_2219 ({sk[458], x729x, x714x, x17002x, n_n199, n_n216, x726x}, x17333x);
	defparam lut_2219.LUT_SIZE = 7;
	defparam lut_2219.mask = 128'h55ff55ff55ff55ff000000150000003f;

	lut_sub lut_2224 ({sk[459], n_n41, n_n40, x51x, x1052x, x1051x, x1795x}, x21403x);
	defparam lut_2224.LUT_SIZE = 7;
	defparam lut_2224.mask = 128'h55ff55ff55ff55fffffff0f088008000;

	lut_sub lut_2229 ({sk[460], n_n101, n_n108, x62x, x202x, x17351x, x21402x}, x17355x);
	defparam lut_2229.LUT_SIZE = 7;
	defparam lut_2229.mask = 128'h55ff55ff55ff55ff00000fffbbbbbfff;

	lut_sub lut_2234 ({sk[461], n_n124, x734x, n_n126, x964x, x963x, x57x}, x17358x);
	defparam lut_2234.LUT_SIZE = 7;
	defparam lut_2234.mask = 128'h55ff55ff55ff55ff0000000f0000777f;

	lut_sub lut_2238 ({sk[462], i_7_, i_8_, i_6_, x734x, x1061x, x1060x}, x17359x);
	defparam lut_2238.LUT_SIZE = 7;
	defparam lut_2238.mask = 128'h55ff55ff55ff55ff0005000300000000;

	lut_sub lut_2241 ({sk[463], n_n101, n_n108, x86x, x263x, x1063x, x1787x}, x17363x);
	defparam lut_2241.LUT_SIZE = 7;
	defparam lut_2241.mask = 128'h55ff55ff55ff55ff000055553fff7fff;

	lut_sub lut_2246 ({sk[464], x734x, n_n126, x51x, x57x, x17354x, x1064x}, x21401x);
	defparam lut_2246.LUT_SIZE = 7;
	defparam lut_2246.mask = 128'h55ff55ff55ff55ffffffffffffff8000;

	lut_sub lut_2250 ({sk[465], i_7_, i_8_, i_6_, x735x}, n_n197);
	defparam lut_2250.LUT_SIZE = 5;
	defparam lut_2250.mask = 32'h1f1f0040;

	lut_sub lut_2252 ({sk[466], i_7_, i_5_, i_6_, i_3_, i_4_, x714x}, n_n212);
	defparam lut_2252.LUT_SIZE = 7;
	defparam lut_2252.mask = 128'h55ff55ff55ff55ff0000000010000000;

	lut_sub lut_2254 ({sk[467], i_14_, i_13_, i_12_, i_15_, n_n191}, x306x);
	defparam lut_2254.LUT_SIZE = 6;
	defparam lut_2254.mask = 64'h11ffffff10005000;

	lut_sub lut_2258 ({sk[468], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1123x);
	defparam lut_2258.LUT_SIZE = 7;
	defparam lut_2258.mask = 128'h55ff55ff55ff55ff0700000077000000;

	lut_sub lut_2265 ({sk[469], x181x, n_n197, n_n212, x168x, x306x, x1123x}, x17379x);
	defparam lut_2265.LUT_SIZE = 7;
	defparam lut_2265.mask = 128'h55ff55ff55ff55ff007f5f7f00ffffff;

	lut_sub lut_2273 ({sk[470], x735x, n_n200, n_n212, x176x, x149x, x965x}, x17369x);
	defparam lut_2273.LUT_SIZE = 7;
	defparam lut_2273.mask = 128'h55ff55ff55ff55ff005f005f005f337f;

	lut_sub lut_2277 ({sk[471], x735x, n_n200, n_n212, x149x, x131x, x966x}, x17370x);
	defparam lut_2277.LUT_SIZE = 7;
	defparam lut_2277.mask = 128'h55ff55ff55ff55ff000f000f000f777f;

	lut_sub lut_2281 ({sk[472], n_n212, x129x, x131x, x17373x}, x4482x);
	defparam lut_2281.LUT_SIZE = 5;
	defparam lut_2281.mask = 32'h1f1f007f;

	lut_sub lut_2285 ({sk[473], n_n197, n_n212, x129x, x130x, x306x, x17371x}, x17375x);
	defparam lut_2285.LUT_SIZE = 7;
	defparam lut_2285.mask = 128'h55ff55ff55ff55ff00000f0f77ff7fff;

	lut_sub lut_2290 ({sk[474], n_n197, n_n212, n_n59, x158x, x299x, x417x}, x17389x);
	defparam lut_2290.LUT_SIZE = 7;
	defparam lut_2290.mask = 128'h55ff55ff55ff55ff00007fff0f0f7fff;

	lut_sub lut_2296 ({sk[475], i_8_, n_n17, x735x, x308x, x21400x, x21422x}, x17390x);
	defparam lut_2296.LUT_SIZE = 7;
	defparam lut_2296.mask = 128'h55ff55ff55ff55ffdddddddfdddddddd;

	lut_sub lut_2300 ({sk[476], n_n123, n_n125, n_n117, n_n102, x94x, x1274x}, x17393x);
	defparam lut_2300.LUT_SIZE = 7;
	defparam lut_2300.mask = 128'h55ff55ff55ff55ff000055ff3fff7fff;

	lut_sub lut_2306 ({sk[477], n_n124, x735x, n_n126, x362x, x1185x, x1183x}, x17394x);
	defparam lut_2306.LUT_SIZE = 7;
	defparam lut_2306.mask = 128'h55ff55ff55ff55ff0000003f0000557f;

	lut_sub lut_2310 ({sk[478], x729x, x735x, n_n126, n_n216, x1125x}, x17397x);
	defparam lut_2310.LUT_SIZE = 6;
	defparam lut_2310.mask = 64'h11ffffff00050007;

	lut_sub lut_2313 ({sk[479], n_n124, x735x, n_n126, x818x, x1124x, x21399x}, x17398x);
	defparam lut_2313.LUT_SIZE = 7;
	defparam lut_2313.mask = 128'h55ff55ff55ff55ffaaaaaaafaaaabbbf;

	lut_sub lut_2317 ({sk[480], n_n31, n_n30, x158x, x1226x, x1225x}, n_n4119);
	defparam lut_2317.LUT_SIZE = 6;
	defparam lut_2317.mask = 64'h11ffffff00335f7f;

	lut_sub lut_2321 ({sk[481], n_n149, n_n31, n_n30, x719x, x122x, x144x}, x17430x);
	defparam lut_2321.LUT_SIZE = 7;
	defparam lut_2321.mask = 128'h55ff55ff55ff55ff00007777000f777f;

	lut_sub lut_2325 ({sk[482], n_n31, n_n30, x125x, x176x, x123x}, x17431x);
	defparam lut_2325.LUT_SIZE = 6;
	defparam lut_2325.mask = 64'h11ffffff00770f7f;

	lut_sub lut_2329 ({sk[483], n_n30, x725x, n_n216, x122x, x646x, x17429x}, x17433x);
	defparam lut_2329.LUT_SIZE = 7;
	defparam lut_2329.mask = 128'h55ff55ff55ff55ff333333337f7f7fff;

	lut_sub lut_2334 ({sk[484], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x950x);
	defparam lut_2334.LUT_SIZE = 7;
	defparam lut_2334.mask = 128'h55ff55ff55ff55ff7000070000700007;

	lut_sub lut_2343 ({sk[485], x725x, n_n34, x125x, n_n216, x949x}, x17451x);
	defparam lut_2343.LUT_SIZE = 6;
	defparam lut_2343.mask = 64'h11ffffff005f007f;

	lut_sub lut_2347 ({sk[486], n_n36, n_n34, x55x, x158x, x176x, x123x}, x17438x);
	defparam lut_2347.LUT_SIZE = 7;
	defparam lut_2347.mask = 128'h55ff55ff55ff55ff00000fff77777fff;

	lut_sub lut_2352 ({sk[487], x181x, n_n36, n_n34, x133x, x127x, x1828x}, x17439x);
	defparam lut_2352.LUT_SIZE = 7;
	defparam lut_2352.mask = 128'h55ff55ff55ff55ff003f557f00ff55ff;

	lut_sub lut_2357 ({sk[488], n_n36, n_n34, x125x, x133x, x176x, x156x}, x17445x);
	defparam lut_2357.LUT_SIZE = 7;
	defparam lut_2357.mask = 128'h55ff55ff55ff55ff000077770fff7fff;

	lut_sub lut_2362 ({sk[489], n_n36, x55x, x127x, x158x, n_n4268, n_n4266}, x17446x);
	defparam lut_2362.LUT_SIZE = 7;
	defparam lut_2362.mask = 128'h55ff55ff55ff55ff777777777fffffff;

	lut_sub lut_2368 ({sk[490], n_n124, x735x, n_n4225, x17461x, x804x, x17460x}, x17466x);
	defparam lut_2368.LUT_SIZE = 7;
	defparam lut_2368.mask = 128'h55ff55ff55ff55ff5fff5fff5fff7fff;

	lut_sub lut_2373 ({sk[491], n_n123, n_n3912, x17456x, n_n142, x141x, x21420x}, x17467x);
	defparam lut_2373.LUT_SIZE = 7;
	defparam lut_2373.mask = 128'h55ff55ff55ff55ffaaffffffbfffffff;

	lut_sub lut_2379 ({sk[492], n_n4441, x575x, x17519x, x17520x, x17521x}, n_n4116);
	defparam lut_2379.LUT_SIZE = 6;
	defparam lut_2379.mask = 64'h11ffffff7fffffff;

	lut_sub lut_2385 ({sk[493], n_n197, n_n212, x158x, n_n4231, n_n3925, x1849x}, x17578x);
	defparam lut_2385.LUT_SIZE = 7;
	defparam lut_2385.mask = 128'h55ff55ff55ff55ff3f3f3fff7f7f7fff;

	lut_sub lut_2390 ({sk[494], n_n212, n_n3921, x1270x, x17573x, x17114x, x17115x}, x17579x);
	defparam lut_2390.LUT_SIZE = 7;
	defparam lut_2390.mask = 128'h55ff55ff55ff55ff7f7fffff7fffffff;

	lut_sub lut_2396 ({sk[495], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x733x);
	defparam lut_2396.LUT_SIZE = 7;
	defparam lut_2396.mask = 128'h55ff55ff55ff55ff1000000000000000;

	lut_sub lut_2398 ({sk[496], i_7_, i_8_, i_6_}, x747x);
	defparam lut_2398.LUT_SIZE = 4;
	defparam lut_2398.mask = 16'h5520;

	lut_sub lut_2400 ({sk[497], i_14_, i_13_, i_12_, i_15_}, x717x);
	defparam lut_2400.LUT_SIZE = 5;
	defparam lut_2400.mask = 32'h1f1f4000;

	lut_sub lut_2402 ({sk[498], i_9_, i_10_, i_11_, x717x}, n_n144);
	defparam lut_2402.LUT_SIZE = 5;
	defparam lut_2402.mask = 32'h1f1f0400;

	lut_sub lut_2404 ({sk[499], i_9_, i_10_, i_11_, x730x}, n_n68);
	defparam lut_2404.LUT_SIZE = 5;
	defparam lut_2404.mask = 32'h1f1f0400;

	lut_sub lut_2406 ({sk[500], i_7_, i_6_, i_1_, i_2_, i_0_, n_n111}, n_n7257);
	defparam lut_2406.LUT_SIZE = 7;
	defparam lut_2406.mask = 128'h55ff55ff55ff55ff0000000010000000;

	lut_sub lut_2408 ({sk[501], i_7_, i_6_, i_1_, i_2_, i_0_, n_n111}, x568x);
	defparam lut_2408.LUT_SIZE = 7;
	defparam lut_2408.mask = 128'h55ff55ff55ff55ff0000000010001000;

	lut_sub lut_2411 ({sk[502], i_7_, i_6_, i_1_, i_2_, i_0_, n_n111}, n_n7258);
	defparam lut_2411.LUT_SIZE = 7;
	defparam lut_2411.mask = 128'h55ff55ff55ff55ff0000100000000000;

	lut_sub lut_2413 ({sk[503], i_9_, i_10_, i_11_, x725x}, n_n53);
	defparam lut_2413.LUT_SIZE = 5;
	defparam lut_2413.mask = 32'h1f1f0004;

	lut_sub lut_2415 ({sk[504], n_n101, n_n108, x176x, x1892x, x1317x, x1316x}, n_n3822);
	defparam lut_2415.LUT_SIZE = 7;
	defparam lut_2415.mask = 128'h55ff55ff55ff55ff00005fff33337fff;

	lut_sub lut_2420 ({sk[505], n_n124, x734x, n_n126, x1489x, x1319x, x1318x}, n_n3823);
	defparam lut_2420.LUT_SIZE = 7;
	defparam lut_2420.mask = 128'h55ff55ff55ff55ff0000005f0000337f;

	lut_sub lut_2424 ({sk[506], n_n53, x157x, n_n101, x445x, n_n108, x1488x}, n_n3895);
	defparam lut_2424.LUT_SIZE = 7;
	defparam lut_2424.mask = 128'h55ff55ff55ff55ff0f5f3f7f3f7f3f7f;

	lut_sub lut_2429 ({sk[507], n_n134, x725x, n_n101, x721x, n_n216, x17625x}, x4173x);
	defparam lut_2429.LUT_SIZE = 7;
	defparam lut_2429.mask = 128'h55ff55ff55ff55ff0057007700ff00ff;

	lut_sub lut_2434 ({sk[508], n_n124, x734x, n_n126, n_n59, x80x, x1320x}, x17626x);
	defparam lut_2434.LUT_SIZE = 7;
	defparam lut_2434.mask = 128'h55ff55ff55ff55ff0000007700000f7f;

	lut_sub lut_2438 ({sk[509], n_n3822, n_n3823, n_n3895, x4173x, x17626x}, n_n3794);
	defparam lut_2438.LUT_SIZE = 6;
	defparam lut_2438.mask = 64'h11ffffff7fffffff;

	lut_sub lut_2444 ({sk[510], n_n53, n_n6267, n_n6266, x172x, n_n47, x21415x}, x17639x);
	defparam lut_2444.LUT_SIZE = 7;
	defparam lut_2444.mask = 128'h55ff55ff55ff55ff57ffffff77ffffff;

	lut_sub lut_2450 ({sk[511], i_7_, i_8_, i_6_, x740x, x1314x, x21443x}, x17640x);
	defparam lut_2450.LUT_SIZE = 7;
	defparam lut_2450.mask = 128'h55ff55ff55ff55ffaaaaaaaaaaabaaaa;

	lut_sub lut_2453 ({sk[512], n_n46, n_n138, n_n47, x4100x, x176x, x1895x}, x17690x);
	defparam lut_2453.LUT_SIZE = 7;
	defparam lut_2453.mask = 128'h55ff55ff55ff55ff0f0f0fff7f7f7fff;

	lut_sub lut_2458 ({sk[513], x714x, x17051x, x125x, x123x, x21444x}, x17691x);
	defparam lut_2458.LUT_SIZE = 6;
	defparam lut_2458.mask = 64'h11ffffffaaaaaabf;

	lut_sub lut_2462 ({sk[514], i_8_, x734x, n_n18, n_n43, x63x, x48x}, x17693x);
	defparam lut_2462.LUT_SIZE = 7;
	defparam lut_2462.mask = 128'h55ff55ff55ff55ff0707077707070707;

	lut_sub lut_2467 ({sk[515], x734x, n_n161, n_n43, x52x, x129x, x222x}, x17694x);
	defparam lut_2467.LUT_SIZE = 7;
	defparam lut_2467.mask = 128'h55ff55ff55ff55ff007f007f007f3f7f;

	lut_sub lut_2473 ({sk[516], x17639x, x17640x, x17690x, x17691x, x17693x, x17694x}, x17697x);
	defparam lut_2473.LUT_SIZE = 7;
	defparam lut_2473.mask = 128'h55ff55ff55ff55ff7fffffffffffffff;

	lut_sub lut_2480 ({sk[517], i_8_, x734x, n_n18, x1322x, x17657x, x21411x}, x17659x);
	defparam lut_2480.LUT_SIZE = 7;
	defparam lut_2480.mask = 128'h55ff55ff55ff55ffbbbbbbbfbbbbbbbb;

	lut_sub lut_2484 ({sk[518], x17646x, x17647x, x17650x, x17651x}, x17660x);
	defparam lut_2484.LUT_SIZE = 5;
	defparam lut_2484.mask = 32'h1f1f7fff;

	lut_sub lut_2489 ({sk[519], n_n41, n_n40, n_n3866, x1852x, x1323x, x17681x}, x17684x);
	defparam lut_2489.LUT_SIZE = 7;
	defparam lut_2489.mask = 128'h55ff55ff55ff55ff55ff5fff77ff7fff;

	lut_sub lut_2494 ({sk[520], n_n3864, x17671x, x17676x, x17677x, x17670x}, x17685x);
	defparam lut_2494.LUT_SIZE = 6;
	defparam lut_2494.mask = 64'h11ffffff7fffffff;

	lut_sub lut_2500 ({sk[521], x740x, x181x, n_n161, n_n47, x143x, x154x}, x17703x);
	defparam lut_2500.LUT_SIZE = 7;
	defparam lut_2500.mask = 128'h00ff00ffffffffff03030f0f03770f7f;

	lut_sub lut_2505 ({sk[522], x181x, n_n46, n_n47, x47x, x154x, x17700x}, x17704x);
	defparam lut_2505.LUT_SIZE = 7;
	defparam lut_2505.mask = 128'h00ff00ffffffffff557f5f7f557fffff;

	lut_sub lut_2511 ({sk[523], x46x, n_n46, n_n47, x52x, x129x, x131x}, x17708x);
	defparam lut_2511.LUT_SIZE = 7;
	defparam lut_2511.mask = 128'h00ff00ffffffffff00337f7f00ff7fff;

	lut_sub lut_2517 ({sk[524], x714x, x17051x, x52x, x63x, x48x, x1458x}, x17709x);
	defparam lut_2517.LUT_SIZE = 7;
	defparam lut_2517.mask = 128'h00ff00ffffffffff0000000000007fff;

	lut_sub lut_2522 ({sk[525], x46x, n_n46, n_n47, x1845x, x1886x, x1884x}, x17710x);
	defparam lut_2522.LUT_SIZE = 7;
	defparam lut_2522.mask = 128'h00ff00ffffffffff00335f7f0033ffff;

	lut_sub lut_2527 ({sk[526], x17703x, x17704x, x17708x, x17709x, x17710x}, n_n3793);
	defparam lut_2527.LUT_SIZE = 6;
	defparam lut_2527.mask = 64'h0055ffff7fffffff;

	lut_sub lut_2533 ({sk[527], x734x, n_n126, n_n112, x47x, x160x, x21382x}, x17718x);
	defparam lut_2533.LUT_SIZE = 7;
	defparam lut_2533.mask = 128'h00ff00ffffffffffaabbaabbaabbafbf;

	lut_sub lut_2537 ({sk[528], n_n123, n_n125, x80x, n_n57, x78x, x1574x}, n_n3909);
	defparam lut_2537.LUT_SIZE = 7;
	defparam lut_2537.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_2542 ({sk[529], x181x, n_n101, n_n108, x1894x, x1378x, x1454x}, x21380x);
	defparam lut_2542.LUT_SIZE = 7;
	defparam lut_2542.mask = 128'h00ff00ffffffffffffc08880ff000000;

	lut_sub lut_2547 ({sk[530], n_n124, n_n53, x157x, x735x, n_n161, x1455x}, x21381x);
	defparam lut_2547.LUT_SIZE = 7;
	defparam lut_2547.mask = 128'h00ff00fffffffffffefefefefef0f0f0;

	lut_sub lut_2553 ({sk[531], x17718x, n_n3909, x21380x, x21381x}, n_n3795);
	defparam lut_2553.LUT_SIZE = 5;
	defparam lut_2553.mask = 32'h5757efff;

	lut_sub lut_2558 ({sk[532], x137x, x46x, n_n197, n_n212, x63x, x48x}, x17768x);
	defparam lut_2558.LUT_SIZE = 7;
	defparam lut_2558.mask = 128'h00ff00ffffffffff00770f7f0f7f0f7f;

	lut_sub lut_2563 ({sk[533], x735x, n_n200, n_n212, x52x, x129x, x63x}, x17769x);
	defparam lut_2563.LUT_SIZE = 7;
	defparam lut_2563.mask = 128'h00ff00ffffffffff007f007f007f3f7f;

	lut_sub lut_2569 ({sk[534], n_n197, n_n212, x123x, x1878x, x131x, x1230x}, x17771x);
	defparam lut_2569.LUT_SIZE = 7;
	defparam lut_2569.mask = 128'h00ff00ffffffffff00000fff77777fff;

	lut_sub lut_2574 ({sk[535], x181x, n_n197, n_n212, x143x, x48x, x154x}, x17774x);
	defparam lut_2574.LUT_SIZE = 7;
	defparam lut_2574.mask = 128'h00ff00ffffffffff00335f7f0033ffff;

	lut_sub lut_2579 ({sk[536], x181x, n_n212, x1572x, n_n4692, x629x, x1833x}, x21384x);
	defparam lut_2579.LUT_SIZE = 7;
	defparam lut_2579.mask = 128'h00ff00ffffffffffc0c08000c0c00000;

	lut_sub lut_2582 ({sk[537], x17768x, x17769x, x17771x, x17774x, x21384x}, x17778x);
	defparam lut_2582.LUT_SIZE = 6;
	defparam lut_2582.mask = 64'h0055ffffbfffffff;

	lut_sub lut_2588 ({sk[538], n_n3912, n_n3828, x17734x, x17746x, x21383x}, n_n3796);
	defparam lut_2588.LUT_SIZE = 6;
	defparam lut_2588.mask = 64'h0055ffffbfffffff;

	lut_sub lut_2594 ({sk[539], n_n123, n_n125, x86x, x180x, x1422x, x17763x}, x17764x);
	defparam lut_2594.LUT_SIZE = 7;
	defparam lut_2594.mask = 128'h00ff00ffffffffff555577775fff7fff;

	lut_sub lut_2599 ({sk[540], n_n3921, n_n3925, x17752x, x17756x, x17751x, x17755x}, x17765x);
	defparam lut_2599.LUT_SIZE = 7;
	defparam lut_2599.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_2606 ({sk[541], i_9_, i_10_, i_11_, i_15_, n_n209}, n_n138);
	defparam lut_2606.LUT_SIZE = 6;
	defparam lut_2606.mask = 64'h0055ffff00001000;

	lut_sub lut_2608 ({sk[542], i_14_, i_13_, i_12_, i_15_, n_n191}, x172x);
	defparam lut_2608.LUT_SIZE = 6;
	defparam lut_2608.mask = 64'h0055ffff40100400;

	lut_sub lut_2612 ({sk[543], i_14_, i_13_, i_12_, i_15_, n_n177, n_n191}, x1457x);
	defparam lut_2612.LUT_SIZE = 7;
	defparam lut_2612.mask = 128'h00ff00ffffffffff7000070000700007;

	lut_sub lut_2621 ({sk[544], i_14_, i_13_, i_12_, i_15_, n_n216}, x1873x);
	defparam lut_2621.LUT_SIZE = 6;
	defparam lut_2621.mask = 64'h0055ffff40100401;

	lut_sub lut_2626 ({sk[545], n_n31, n_n30, n_n138, x172x, x1457x, x1873x}, x17786x);
	defparam lut_2626.LUT_SIZE = 7;
	defparam lut_2626.mask = 128'h00ff00ffffffffff000077770fff7fff;

	lut_sub lut_2631 ({sk[546], i_14_, i_13_, i_12_, i_15_, n_n177, n_n191}, x1492x);
	defparam lut_2631.LUT_SIZE = 7;
	defparam lut_2631.mask = 128'h00ff00ffffffffff0757505700000000;

	lut_sub lut_2641 ({sk[547], n_n31, n_n30, x137x, x46x, x1899x, x1492x}, x17798x);
	defparam lut_2641.LUT_SIZE = 7;
	defparam lut_2641.mask = 128'h00ff00ffffffffff00005fff3fff7fff;

	lut_sub lut_2648 ({sk[548], i_14_, i_13_, i_12_, i_15_, n_n156}, x1827x);
	defparam lut_2648.LUT_SIZE = 6;
	defparam lut_2648.mask = 64'h0055ffff00005154;

	lut_sub lut_2655 ({sk[549], i_14_, i_13_, i_12_, i_15_, n_n156}, x1876x);
	defparam lut_2655.LUT_SIZE = 6;
	defparam lut_2655.mask = 64'h0055ffff15450000;

	lut_sub lut_2662 ({sk[550], n_n30, x176x, x134x, x123x, x156x, x131x}, x17789x);
	defparam lut_2662.LUT_SIZE = 7;
	defparam lut_2662.mask = 128'h00ff00ffffffffff000000007fffffff;

	lut_sub lut_2668 ({sk[551], n_n31, n_n30, x181x, x129x, x1725x, x1491x}, n_n3802);
	defparam lut_2668.LUT_SIZE = 7;
	defparam lut_2668.mask = 128'h00ff00ffffffffff000055ff3f3f7fff;

	lut_sub lut_2673 ({sk[552], n_n31, x17798x, x1827x, x1876x, x17789x, n_n3802}, n_n3787);
	defparam lut_2673.LUT_SIZE = 7;
	defparam lut_2673.mask = 128'h00ff00ffffffffff7777ffff7fffffff;

	lut_sub lut_2679 ({sk[553], n_n31, n_n30, x181x, n_n33, x47x, x1519x}, x17819x);
	defparam lut_2679.LUT_SIZE = 7;
	defparam lut_2679.mask = 128'h00ff00ffffffffff0505373705ff37ff;

	lut_sub lut_2683 ({sk[554], n_n31, n_n33, n_n138, x143x, x1825x, x17819x}, x17820x);
	defparam lut_2683.LUT_SIZE = 7;
	defparam lut_2683.mask = 128'h00ff00ffffffffff555555ff7f7f7fff;

	lut_sub lut_2688 ({sk[555], x734x, n_n36, n_n200, n_n190, x187x, x1452x}, x17812x);
	defparam lut_2688.LUT_SIZE = 7;
	defparam lut_2688.mask = 128'h00ff00ffffffffff00005555003f557f;

	lut_sub lut_2692 ({sk[556], i_8_, n_n157, n_n36, x735x, x125x, x1315x}, x17803x);
	defparam lut_2692.LUT_SIZE = 7;
	defparam lut_2692.mask = 128'h00ff00ffffffffff0033053700330033;

	lut_sub lut_2695 ({sk[557], n_n36, n_n191, x719x, n_n63, x176x, x123x}, x17804x);
	defparam lut_2695.LUT_SIZE = 7;
	defparam lut_2695.mask = 128'h00ff00ffffffffff000000007f7f7fff;

	lut_sub lut_2700 ({sk[558], n_n53, x157x, n_n36, n_n34, x588x, x174x}, x17811x);
	defparam lut_2700.LUT_SIZE = 7;
	defparam lut_2700.mask = 128'h00ff00ffffffffff373737ff37ff37ff;

	lut_sub lut_2705 ({sk[559], n_n34, x176x, x134x, x123x, x156x, x1453x}, x21379x);
	defparam lut_2705.LUT_SIZE = 7;
	defparam lut_2705.mask = 128'h00ff00ffffffffffffffffff80000000;

	lut_sub lut_2708 ({sk[560], x17812x, x17803x, x17804x, x17811x, x21379x}, x17821x);
	defparam lut_2708.LUT_SIZE = 6;
	defparam lut_2708.mask = 64'h0055ffffbfffffff;

	lut_sub lut_2714 ({sk[561], x181x, n_n36, n_n34, x143x, x154x}, x17829x);
	defparam lut_2714.LUT_SIZE = 6;
	defparam lut_2714.mask = 64'h0055ffff07370f3f;

	lut_sub lut_2719 ({sk[562], i_8_, n_n157, x181x, n_n36, x735x, x47x}, x17827x);
	defparam lut_2719.LUT_SIZE = 7;
	defparam lut_2719.mask = 128'h00ff00ffffffffff000f111f000f000f;

	lut_sub lut_2722 ({sk[563], n_n6646, x393x, x392x, n_n36, x47x, x154x}, x17828x);
	defparam lut_2722.LUT_SIZE = 7;
	defparam lut_2722.mask = 128'h00ff00ffffffffff07ffffffffffffff;

	lut_sub lut_2728 ({sk[564], n_n36, n_n34, x134x, x63x, x156x, x48x}, x17833x);
	defparam lut_2728.LUT_SIZE = 7;
	defparam lut_2728.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_2733 ({sk[565], x137x, x46x, n_n36, n_n34, x63x, x48x}, x17834x);
	defparam lut_2733.LUT_SIZE = 7;
	defparam lut_2733.mask = 128'h00ff00ffffffffff00770f7f0f7f0f7f;

	lut_sub lut_2738 ({sk[566], x17829x, x17827x, x17828x, x17833x, x17834x}, x17839x);
	defparam lut_2738.LUT_SIZE = 6;
	defparam lut_2738.mask = 64'h0055ffff7fffffff;

	lut_sub lut_2744 ({sk[567], i_14_, i_13_, i_12_, i_15_, n_n156}, x83x);
	defparam lut_2744.LUT_SIZE = 6;
	defparam lut_2744.mask = 64'h0055ffff00100400;

	lut_sub lut_2747 ({sk[568], i_14_, i_13_, i_12_, i_15_, n_n156}, x157x);
	defparam lut_2747.LUT_SIZE = 6;
	defparam lut_2747.mask = 64'h0055ffff00100401;

	lut_sub lut_2751 ({sk[569], i_7_, i_8_, i_6_, n_n162, x734x, x714x}, x213x);
	defparam lut_2751.LUT_SIZE = 7;
	defparam lut_2751.mask = 128'h00ff00ffffffffff3700050000000000;

	lut_sub lut_2754 ({sk[570], n_n36, n_n34, x127x, x123x, x146x, x131x}, x17867x);
	defparam lut_2754.LUT_SIZE = 7;
	defparam lut_2754.mask = 128'h00ff00ffffffffff000077ff0f0f7fff;

	lut_sub lut_2759 ({sk[571], x137x, n_n36, n_n34, x55x, x1828x, x176x}, x17868x);
	defparam lut_2759.LUT_SIZE = 7;
	defparam lut_2759.mask = 128'h00ff00ffffffffff000f777f00ff77ff;

	lut_sub lut_2764 ({sk[572], n_n36, n_n34, x130x, x63x, x48x}, x17869x);
	defparam lut_2764.LUT_SIZE = 6;
	defparam lut_2764.mask = 64'h0055ffff00770f7f;

	lut_sub lut_2768 ({sk[573], x137x, x46x, n_n36, n_n3961, x1877x, x3945x}, x17870x);
	defparam lut_2768.LUT_SIZE = 7;
	defparam lut_2768.mask = 128'h00ff00ffffffffff5f7f5fff5fff5fff;

	lut_sub lut_2774 ({sk[574], x132x, n_n36, n_n34, x147x, x126x}, x17874x);
	defparam lut_2774.LUT_SIZE = 6;
	defparam lut_2774.mask = 64'h0055ffff037703ff;

	lut_sub lut_2779 ({sk[575], x46x, n_n36, n_n34, x149x, x126x, x17871x}, x17875x);
	defparam lut_2779.LUT_SIZE = 7;
	defparam lut_2779.mask = 128'h00ff00ffffffffff00770f7f00ff0fff;

	lut_sub lut_2784 ({sk[576], n_n36, n_n34, x168x, x74x, x151x}, n_n4461);
	defparam lut_2784.LUT_SIZE = 6;
	defparam lut_2784.mask = 64'h0055ffff003f557f;

	lut_sub lut_2788 ({sk[577], x181x, n_n36, x143x, x47x, x154x, x21413x}, x597x);
	defparam lut_2788.LUT_SIZE = 7;
	defparam lut_2788.mask = 128'h00ff00ffffffffffaaaabfffaaaaffff;

	lut_sub lut_2794 ({sk[578], n_n36, n_n34, x143x, x866x, x47x, x154x}, x620x);
	defparam lut_2794.LUT_SIZE = 7;
	defparam lut_2794.mask = 128'h00ff00ffffffffff000077ff0f0f7fff;

	lut_sub lut_2799 ({sk[579], n_n36, n_n34, x52x, x129x, x1627x}, x17882x);
	defparam lut_2799.LUT_SIZE = 6;
	defparam lut_2799.mask = 64'h0055ffff00553f7f;

	lut_sub lut_2803 ({sk[580], n_n36, n_n4581, x139x, x63x, x48x, x1882x}, x21378x);
	defparam lut_2803.LUT_SIZE = 7;
	defparam lut_2803.mask = 128'h00ff00ffffffffffffff000080000000;

	lut_sub lut_2806 ({sk[581], n_n34, n_n63, x176x, x4992x, x709x, x153x}, x17893x);
	defparam lut_2806.LUT_SIZE = 7;
	defparam lut_2806.mask = 128'h00ff00ffffffffff3f3f3f3f7fffffff;

	lut_sub lut_2812 ({sk[582], n_n36, n_n34, x125x, x1698x, x1697x}, x17894x);
	defparam lut_2812.LUT_SIZE = 6;
	defparam lut_2812.mask = 64'h0055ffff005f3f7f;

	lut_sub lut_2817 ({sk[583], n_n34, x133x, x134x, x123x, x156x}, x17899x);
	defparam lut_2817.LUT_SIZE = 6;
	defparam lut_2817.mask = 64'h0055ffff00007fff;

	lut_sub lut_2822 ({sk[584], n_n36, n_n34, x55x, x133x, x127x, x158x}, x17900x);
	defparam lut_2822.LUT_SIZE = 7;
	defparam lut_2822.mask = 128'h00ff00ffffffffff000055557fff7fff;

	lut_sub lut_2828 ({sk[585], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x765x);
	defparam lut_2828.LUT_SIZE = 7;
	defparam lut_2828.mask = 128'h00ff00ffffffffff7000070000700007;

	lut_sub lut_2837 ({sk[586], i_9_, i_10_, i_11_, i_15_, n_n209}, n_n128);
	defparam lut_2837.LUT_SIZE = 6;
	defparam lut_2837.mask = 64'h0055ffff00100000;

	lut_sub lut_2839 ({sk[587], i_14_, i_13_, i_12_, i_15_, n_n149}, x152x);
	defparam lut_2839.LUT_SIZE = 6;
	defparam lut_2839.mask = 64'h0055ffff40100400;

	lut_sub lut_2843 ({sk[588], n_n31, x158x, x149x, x1827x, x1876x, x1624x}, n_n3467);
	defparam lut_2843.LUT_SIZE = 7;
	defparam lut_2843.mask = 128'h00ff00ffffffffff000000007fffffff;

	lut_sub lut_2849 ({sk[589], n_n162, n_n157, x46x, x714x, x129x, x1108x}, x17932x);
	defparam lut_2849.LUT_SIZE = 7;
	defparam lut_2849.mask = 128'h00ff00ffffffffff000000000000070f;

	lut_sub lut_2853 ({sk[590], n_n31, x137x, x146x, x131x, x1725x}, x17933x);
	defparam lut_2853.LUT_SIZE = 6;
	defparam lut_2853.mask = 64'h0055ffff00007fff;

	lut_sub lut_2858 ({sk[591], n_n31, x132x, x147x, x126x, x1625x}, x17934x);
	defparam lut_2858.LUT_SIZE = 6;
	defparam lut_2858.mask = 64'h0055ffff00007fff;

	lut_sub lut_2863 ({sk[592], i_14_, i_13_, i_12_, i_15_, n_n32, n_n184}, x3810x);
	defparam lut_2863.LUT_SIZE = 7;
	defparam lut_2863.mask = 128'h00ff00ffffffffff0000000001010110;

	lut_sub lut_2868 ({sk[593], n_n36, n_n132, x78x, x217x, x17941x, x21376x}, x3811x);
	defparam lut_2868.LUT_SIZE = 7;
	defparam lut_2868.mask = 128'h00ff00ffffffffff00000000bfffffff;

	lut_sub lut_2874 ({sk[594], n_n162, n_n157, x714x, x151x, x47x, x154x}, x17948x);
	defparam lut_2874.LUT_SIZE = 7;
	defparam lut_2874.mask = 128'h00ff00ffffffffff000000000000007f;

	lut_sub lut_2878 ({sk[595], n_n31, x181x, n_n32, x143x, x1648x}, x17949x);
	defparam lut_2878.LUT_SIZE = 6;
	defparam lut_2878.mask = 64'h0055ffff050537ff;

	lut_sub lut_2882 ({sk[596], n_n36, n_n138, x176x, x123x, x153x, x356x}, x17951x);
	defparam lut_2882.LUT_SIZE = 7;
	defparam lut_2882.mask = 128'h00ff00ffffffffff000000007fffffff;

	lut_sub lut_2888 ({sk[597], n_n36, x125x, x55x, x133x, x127x, x158x}, x17952x);
	defparam lut_2888.LUT_SIZE = 7;
	defparam lut_2888.mask = 128'h00ff00ffffffffff000000007fffffff;

	lut_sub lut_2894 ({sk[598], i_14_, i_13_, i_12_, i_15_, n_n36, n_n216}, x17958x);
	defparam lut_2894.LUT_SIZE = 7;
	defparam lut_2894.mask = 128'h00ff00ffffffffff0111101111011110;

	lut_sub lut_2907 ({sk[599], n_n39, n_n36, n_n132, x151x, x866x, x434x}, x17959x);
	defparam lut_2907.LUT_SIZE = 7;
	defparam lut_2907.mask = 128'h00ff00ffffffffff55557f7f55ff7fff;

	lut_sub lut_2912 ({sk[600], x132x, n_n36, x134x, x156x, x126x}, x17961x);
	defparam lut_2912.LUT_SIZE = 6;
	defparam lut_2912.mask = 64'h0055ffff007f00ff;

	lut_sub lut_2917 ({sk[601], x137x, n_n36, x149x, x146x, x147x, x131x}, x17962x);
	defparam lut_2917.LUT_SIZE = 7;
	defparam lut_2917.mask = 128'h00ff00ffffffffff00007fff0000ffff;

	lut_sub lut_2923 ({sk[602], i_14_, i_13_, i_12_, i_15_, n_n36, n_n191}, x17966x);
	defparam lut_2923.LUT_SIZE = 7;
	defparam lut_2923.mask = 128'h00ff00ffffffffff0111101111011110;

	lut_sub lut_2936 ({sk[603], x46x, n_n36, x124x, x130x, x139x, x128x}, x17967x);
	defparam lut_2936.LUT_SIZE = 7;
	defparam lut_2936.mask = 128'h00ff00ffffffffff00007fff0000ffff;

	lut_sub lut_2942 ({sk[604], x3676x, x18085x, x3671x, x18091x, x18096x}, n_n3464);
	defparam lut_2942.LUT_SIZE = 6;
	defparam lut_2942.mask = 64'h0055ffff7fffffff;

	lut_sub lut_2948 ({sk[605], n_n3494, x3658x, x18113x, x3653x, x18118x}, n_n3463);
	defparam lut_2948.LUT_SIZE = 6;
	defparam lut_2948.mask = 64'h0055ffff7fffffff;

	lut_sub lut_2954 ({sk[606], n_n3485, x18033x, x18034x, x18037x, x18038x}, n_n3460);
	defparam lut_2954.LUT_SIZE = 6;
	defparam lut_2954.mask = 64'h0055ffff7fffffff;

	lut_sub lut_2960 ({sk[607], n_n3492, n_n3491, x18057x, x18058x}, n_n3462);
	defparam lut_2960.LUT_SIZE = 5;
	defparam lut_2960.mask = 32'h57577fff;

	lut_sub lut_2965 ({sk[608], x445x, n_n3489, x3685x, x21435x}, x18078x);
	defparam lut_2965.LUT_SIZE = 5;
	defparam lut_2965.mask = 32'h5757bfff;

	lut_sub lut_2970 ({sk[609], x18124x, x18127x, x18130x, x18131x, x21374x}, x18134x);
	defparam lut_2970.LUT_SIZE = 6;
	defparam lut_2970.mask = 64'h0055ffffbfffffff;

	lut_sub lut_2976 ({sk[610], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x741x);
	defparam lut_2976.LUT_SIZE = 7;
	defparam lut_2976.mask = 128'h00ff00ffffffffff0000000000400000;

	lut_sub lut_2978 ({sk[611], i_7_, i_6_, i_1_, i_2_, i_0_, n_n48}, n_n7263);
	defparam lut_2978.LUT_SIZE = 7;
	defparam lut_2978.mask = 128'h00ff00ffffffffff1000000000000000;

	lut_sub lut_2980 ({sk[612], i_7_, i_8_, i_6_}, n_n161);
	defparam lut_2980.LUT_SIZE = 4;
	defparam lut_2980.mask = 16'h0f04;

	lut_sub lut_2982 ({sk[613], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x750x);
	defparam lut_2982.LUT_SIZE = 7;
	defparam lut_2982.mask = 128'h00ff00ffffffffff0000000000080000;

	lut_sub lut_2984 ({sk[614], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x744x);
	defparam lut_2984.LUT_SIZE = 7;
	defparam lut_2984.mask = 128'h00ff00ffffffffff0040000000000000;

	lut_sub lut_2986 ({sk[615], i_7_, i_6_, i_1_, i_2_, i_0_, n_n162}, n_n7255);
	defparam lut_2986.LUT_SIZE = 7;
	defparam lut_2986.mask = 128'h00ff00ffffffffff1000000000000000;

	lut_sub lut_2988 ({sk[616], i_7_, i_8_, i_6_, n_n162, n_n159, n_n48}, x1462x);
	defparam lut_2988.LUT_SIZE = 7;
	defparam lut_2988.mask = 128'h00ff00ffffffffff1113000000000000;

	lut_sub lut_2992 ({sk[617], i_9_, i_10_, i_11_, n_n9, x717x}, x18150x);
	defparam lut_2992.LUT_SIZE = 6;
	defparam lut_2992.mask = 64'h0055ffff00101000;

	lut_sub lut_2995 ({sk[618], i_7_, i_6_, i_1_, i_2_, i_0_, n_n162}, n_n7253);
	defparam lut_2995.LUT_SIZE = 7;
	defparam lut_2995.mask = 128'h00ff00ffffffffff0000000010000000;

	lut_sub lut_2997 ({sk[619], i_9_, i_10_, i_11_, x717x}, n_n186);
	defparam lut_2997.LUT_SIZE = 5;
	defparam lut_2997.mask = 32'h57570040;

	lut_sub lut_2999 ({sk[620], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x285x);
	defparam lut_2999.LUT_SIZE = 7;
	defparam lut_2999.mask = 128'h00ff00ffffffffff8000000000000000;

	lut_sub lut_3001 ({sk[621], i_9_, i_10_, i_11_, n_n126, x285x}, n_n6267);
	defparam lut_3001.LUT_SIZE = 6;
	defparam lut_3001.mask = 64'h0055ffff00000010;

	lut_sub lut_3003 ({sk[622], i_14_, i_13_, i_12_, i_15_, n_n149, n_n47}, x3607x);
	defparam lut_3003.LUT_SIZE = 7;
	defparam lut_3003.mask = 128'h00ff00ffffffffff1000010000100000;

	lut_sub lut_3007 ({sk[623], i_15_, n_n149, n_n53, x714x, x17051x, n_n209}, x17554x);
	defparam lut_3007.LUT_SIZE = 7;
	defparam lut_3007.mask = 128'h00ff00ffffffffff0003000300030103;

	lut_sub lut_3010 ({sk[624], i_14_, i_13_, i_12_, i_15_, n_n149}, x1823x);
	defparam lut_3010.LUT_SIZE = 6;
	defparam lut_3010.mask = 64'h0055ffff40100401;

	lut_sub lut_3015 ({sk[625], x740x, n_n161, n_n47, x55x, x127x, x1886x}, x18184x);
	defparam lut_3015.LUT_SIZE = 7;
	defparam lut_3015.mask = 128'h00ff00ffffffffff0055005500553f7f;

	lut_sub lut_3019 ({sk[626], n_n46, n_n47, x176x, x123x, x131x, x1845x}, x18185x);
	defparam lut_3019.LUT_SIZE = 7;
	defparam lut_3019.mask = 128'h00ff00ffffffffff00000fff77777fff;

	lut_sub lut_3024 ({sk[627], x46x, n_n46, n_n47, x52x, x129x, x1458x}, x18187x);
	defparam lut_3024.LUT_SIZE = 7;
	defparam lut_3024.mask = 128'h00ff00ffffffffff00553f7f00ff3fff;

	lut_sub lut_3029 ({sk[628], x740x, x46x, n_n161, n_n47, x149x, x1271x}, x18211x);
	defparam lut_3029.LUT_SIZE = 7;
	defparam lut_3029.mask = 128'h00ff00ffffffffff03030303035703ff;

	lut_sub lut_3033 ({sk[629], n_n46, n_n47, x130x, x147x, x1884x, x1893x}, x21373x);
	defparam lut_3033.LUT_SIZE = 7;
	defparam lut_3033.mask = 128'h00ff00ffffffffffffffa000cccc8000;

	lut_sub lut_3038 ({sk[630], i_7_, i_8_, i_6_, n_n177, x285x}, n_n6266);
	defparam lut_3038.LUT_SIZE = 6;
	defparam lut_3038.mask = 64'h0055ffff00010000;

	lut_sub lut_3040 ({sk[631], i_7_, i_8_, i_6_, n_n149, n_n156, x285x}, x435x);
	defparam lut_3040.LUT_SIZE = 7;
	defparam lut_3040.mask = 128'h00ff00ffffffffff0011000500000000;

	lut_sub lut_3043 ({sk[632], i_8_, i_1_, i_2_, i_0_, x17002x}, n_n41);
	defparam lut_3043.LUT_SIZE = 6;
	defparam lut_3043.mask = 64'h0055ffff00004000;

	lut_sub lut_3045 ({sk[633], i_14_, i_13_, i_12_, i_15_, n_n149}, x245x);
	defparam lut_3045.LUT_SIZE = 6;
	defparam lut_3045.mask = 64'h0055ffff00100401;

	lut_sub lut_3049 ({sk[634], i_7_, i_8_, i_6_}, n_n200);
	defparam lut_3049.LUT_SIZE = 4;
	defparam lut_3049.mask = 16'h0f08;

	lut_sub lut_3051 ({sk[635], i_9_, i_10_, i_11_, x725x}, n_n57);
	defparam lut_3051.LUT_SIZE = 5;
	defparam lut_3051.mask = 32'h57570010;

	lut_sub lut_3053 ({sk[636], i_14_, i_13_, i_12_, i_15_, n_n156}, x144x);
	defparam lut_3053.LUT_SIZE = 6;
	defparam lut_3053.mask = 64'h0055ffff00000401;

	lut_sub lut_3056 ({sk[637], x740x, n_n200, x714x, x17002x, n_n57, x144x}, n_n5055);
	defparam lut_3056.LUT_SIZE = 7;
	defparam lut_3056.mask = 128'h00ff00ffffffffff0005000500053337;

	lut_sub lut_3059 ({sk[638], i_14_, i_13_, i_12_, i_15_, n_n40, n_n177}, n_n5056);
	defparam lut_3059.LUT_SIZE = 7;
	defparam lut_3059.mask = 128'h00ff00ffffffffff0000010000100001;

	lut_sub lut_3063 ({sk[639], i_14_, i_13_, i_12_, i_15_, n_n156}, x1815x);
	defparam lut_3063.LUT_SIZE = 6;
	defparam lut_3063.mask = 64'h0055ffff40100401;

	lut_sub lut_3068 ({sk[640], n_n149, x725x, n_n40, x714x, x17002x, x1815x}, x387x);
	defparam lut_3068.LUT_SIZE = 7;
	defparam lut_3068.mask = 128'h00ff00ffffffffff0055005500550357;

	lut_sub lut_3071 ({sk[641], x18232x, x18237x, x21371x, x21372x}, n_n3031);
	defparam lut_3071.LUT_SIZE = 5;
	defparam lut_3071.mask = 32'h5757efff;

	lut_sub lut_3076 ({sk[642], n_n41, n_n40, n_n117, x98x, x1175x, x1174x}, n_n3042);
	defparam lut_3076.LUT_SIZE = 7;
	defparam lut_3076.mask = 128'h00ff00ffffffffff00003f3f55ff7fff;

	lut_sub lut_3081 ({sk[643], x18273x, x18274x, x3484x, x18283x, x18286x, x18287x}, n_n3029);
	defparam lut_3081.LUT_SIZE = 7;
	defparam lut_3081.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_3088 ({sk[644], i_8_, x740x, n_n17, n_n77, x1331x, x21445x}, x18266x);
	defparam lut_3088.LUT_SIZE = 7;
	defparam lut_3088.mask = 128'h00ff00ffffffffff5555557f55555555;

	lut_sub lut_3092 ({sk[645], n_n89, n_n41, n_n40, x1111x, x1460x, x1459x}, x21369x);
	defparam lut_3092.LUT_SIZE = 7;
	defparam lut_3092.mask = 128'h00ff00ffffffffffffaac080ff00c000;

	lut_sub lut_3097 ({sk[646], i_14_, i_13_, i_12_, i_15_, n_n156}, x122x);
	defparam lut_3097.LUT_SIZE = 6;
	defparam lut_3097.mask = 64'h0055ffff40100000;

	lut_sub lut_3100 ({sk[647], i_14_, i_13_, i_12_, i_15_, n_n149}, x1865x);
	defparam lut_3100.LUT_SIZE = 6;
	defparam lut_3100.mask = 64'h0055ffff40100401;

	lut_sub lut_3105 ({sk[648], i_14_, i_13_, i_12_, i_15_}, x721x);
	defparam lut_3105.LUT_SIZE = 5;
	defparam lut_3105.mask = 32'h57570400;

	lut_sub lut_3107 ({sk[649], x725x, x714x, x17002x, x721x, n_n170, x728x}, x4900x);
	defparam lut_3107.LUT_SIZE = 7;
	defparam lut_3107.mask = 128'h00ff00ffffffffff0000001300000033;

	lut_sub lut_3111 ({sk[650], i_5_, i_3_, i_4_, n_n159, n_n51, x747x}, n_n7294);
	defparam lut_3111.LUT_SIZE = 7;
	defparam lut_3111.mask = 128'h00ff00ffffffffff0001000000000000;

	lut_sub lut_3113 ({sk[651], i_5_, i_3_, i_4_, n_n159, n_n126}, x751x);
	defparam lut_3113.LUT_SIZE = 6;
	defparam lut_3113.mask = 64'h0055ffff01000000;

	lut_sub lut_3115 ({sk[652], i_7_, i_5_, i_6_, i_3_, i_4_, x714x}, n_n32);
	defparam lut_3115.LUT_SIZE = 7;
	defparam lut_3115.mask = 128'h00ff00ffffffffff0000000000004000;

	lut_sub lut_3117 ({sk[653], i_14_, i_13_, i_12_, i_15_, n_n184}, x124x);
	defparam lut_3117.LUT_SIZE = 6;
	defparam lut_3117.mask = 64'h0055ffff00001110;

	lut_sub lut_3121 ({sk[654], i_14_, i_13_, i_12_, i_15_, n_n184}, x1417x);
	defparam lut_3121.LUT_SIZE = 6;
	defparam lut_3121.mask = 64'h0055ffff40000401;

	lut_sub lut_3125 ({sk[655], i_14_, i_13_, i_12_}, n_n201);
	defparam lut_3125.LUT_SIZE = 4;
	defparam lut_3125.mask = 16'h0f20;

	lut_sub lut_3127 ({sk[656], i_9_, i_10_, i_11_, i_15_, n_n32, n_n201}, x3461x);
	defparam lut_3127.LUT_SIZE = 7;
	defparam lut_3127.mask = 128'h00ff00ffffffffff0100000000000000;

	lut_sub lut_3129 ({sk[657], i_7_, i_8_, i_6_, x734x, n_n132, n_n52}, x18300x);
	defparam lut_3129.LUT_SIZE = 7;
	defparam lut_3129.mask = 128'h00ff00ffffffffff0000000007000000;

	lut_sub lut_3132 ({sk[658], i_14_, i_13_, i_12_, i_15_, n_n184}, x130x);
	defparam lut_3132.LUT_SIZE = 6;
	defparam lut_3132.mask = 64'h0055ffff04440000;

	lut_sub lut_3136 ({sk[659], i_14_, i_13_, i_12_, i_15_, n_n191}, x48x);
	defparam lut_3136.LUT_SIZE = 6;
	defparam lut_3136.mask = 64'h0055ffff00001110;

	lut_sub lut_3140 ({sk[660], i_14_, i_13_, i_12_, i_15_, n_n184}, x1883x);
	defparam lut_3140.LUT_SIZE = 6;
	defparam lut_3140.mask = 64'h0055ffff11014044;

	lut_sub lut_3147 ({sk[661], i_14_, i_13_, i_12_, i_15_, n_n149, n_n33}, n_n2733);
	defparam lut_3147.LUT_SIZE = 7;
	defparam lut_3147.mask = 128'h00ff00ffffffffff1000010000000001;

	lut_sub lut_3151 ({sk[662], i_14_, i_13_, i_12_, i_15_, n_n170}, x1858x);
	defparam lut_3151.LUT_SIZE = 6;
	defparam lut_3151.mask = 64'h0055ffff00005154;

	lut_sub lut_3158 ({sk[663], i_14_, i_13_, i_12_, i_15_, n_n191}, x145x);
	defparam lut_3158.LUT_SIZE = 6;
	defparam lut_3158.mask = 64'h0055ffff00404000;

	lut_sub lut_3161 ({sk[664], i_14_, i_13_, i_12_, i_15_, n_n149}, x170x);
	defparam lut_3161.LUT_SIZE = 6;
	defparam lut_3161.mask = 64'h0055ffff00404000;

	lut_sub lut_3164 ({sk[665], n_n71, n_n89, x288x, n_n4, n_n18, x95x}, x18317x);
	defparam lut_3164.LUT_SIZE = 7;
	defparam lut_3164.mask = 128'h00ff00ffffffffff05370f3f0f3f0f3f;

	lut_sub lut_3169 ({sk[666], i_7_, i_8_, i_6_, x735x}, n_n112);
	defparam lut_3169.LUT_SIZE = 5;
	defparam lut_3169.mask = 32'h57570010;

	lut_sub lut_3171 ({sk[667], i_7_, i_5_, i_6_, i_3_, i_4_, x714x}, n_n113);
	defparam lut_3171.LUT_SIZE = 7;
	defparam lut_3171.mask = 128'h00ff00ffffffffff0000000000100000;

	lut_sub lut_3173 ({sk[668], i_14_, i_13_, i_12_, i_15_, n_n184}, x1113x);
	defparam lut_3173.LUT_SIZE = 6;
	defparam lut_3173.mask = 64'h0055ffff55455555;

	lut_sub lut_3189 ({sk[669], i_14_, i_13_, i_12_, i_15_, n_n191}, x1112x);
	defparam lut_3189.LUT_SIZE = 6;
	defparam lut_3189.mask = 64'h0055ffff15451110;

	lut_sub lut_3199 ({sk[670], n_n42, n_n43, x62x, n_n183, x1782x, x1798x}, x18353x);
	defparam lut_3199.LUT_SIZE = 7;
	defparam lut_3199.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_3204 ({sk[671], i_7_, i_5_, i_6_, i_3_, i_4_, n_n159}, x430x);
	defparam lut_3204.LUT_SIZE = 7;
	defparam lut_3204.mask = 128'h00ff00ffffffffff0000000010000000;

	lut_sub lut_3206 ({sk[672], n_n149, x717x, n_n2, x430x, x730x}, x708x);
	defparam lut_3206.LUT_SIZE = 6;
	defparam lut_3206.mask = 64'h0055ffff3333373f;

	lut_sub lut_3210 ({sk[673], i_9_, i_10_, i_11_, x729x, x717x, x730x}, x238x);
	defparam lut_3210.LUT_SIZE = 7;
	defparam lut_3210.mask = 128'h00ff00ffffffffff00000f0077000000;

	lut_sub lut_3214 ({sk[674], i_7_, i_8_, i_6_, x735x}, n_n123);
	defparam lut_3214.LUT_SIZE = 5;
	defparam lut_3214.mask = 32'h57571000;

	lut_sub lut_3216 ({sk[675], i_14_, i_13_, i_12_, i_15_, n_n170}, x147x);
	defparam lut_3216.LUT_SIZE = 6;
	defparam lut_3216.mask = 64'h0055ffff11010000;

	lut_sub lut_3220 ({sk[676], i_14_, i_13_, i_12_, i_15_, n_n170}, x958x);
	defparam lut_3220.LUT_SIZE = 6;
	defparam lut_3220.mask = 64'h0055ffff04445154;

	lut_sub lut_3230 ({sk[677], i_14_, i_13_, i_12_, i_15_, n_n149}, x133x);
	defparam lut_3230.LUT_SIZE = 6;
	defparam lut_3230.mask = 64'h0055ffff11010000;

	lut_sub lut_3234 ({sk[678], i_14_, i_13_, i_12_, i_15_, n_n149}, x960x);
	defparam lut_3234.LUT_SIZE = 6;
	defparam lut_3234.mask = 64'h0055ffff15455154;

	lut_sub lut_3247 ({sk[679], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x959x);
	defparam lut_3247.LUT_SIZE = 7;
	defparam lut_3247.mask = 128'h00ff00ffffffffff0535303555055550;

	lut_sub lut_3260 ({sk[680], n_n124, x735x, n_n126, x133x, x960x, x959x}, x18547x);
	defparam lut_3260.LUT_SIZE = 7;
	defparam lut_3260.mask = 128'h00ff00ffffffffff0000003300005f7f;

	lut_sub lut_3264 ({sk[681], x157x, x735x, n_n126, x186x, x209x, x174x}, x3220x);
	defparam lut_3264.LUT_SIZE = 7;
	defparam lut_3264.mask = 128'h00ff00ffffffffff0000007f000000ff;

	lut_sub lut_3269 ({sk[682], n_n123, n_n125, x1334x, x1333x, x252x, x18530x}, x18533x);
	defparam lut_3269.LUT_SIZE = 7;
	defparam lut_3269.mask = 128'h00ff00ffffffffff000000ff7f7f7fff;

	lut_sub lut_3274 ({sk[683], n_n125, x125x, x247x, x171x, x4055x, x18535x}, x18541x);
	defparam lut_3274.LUT_SIZE = 7;
	defparam lut_3274.mask = 128'h00ff00ffffffffff333333337fffffff;

	lut_sub lut_3280 ({sk[684], n_n116, x125x, x176x, x242x, x135x, x153x}, x1396x);
	defparam lut_3280.LUT_SIZE = 7;
	defparam lut_3280.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_3287 ({sk[685], i_7_, i_8_, i_6_, x735x}, n_n125);
	defparam lut_3287.LUT_SIZE = 5;
	defparam lut_3287.mask = 32'h57570100;

	lut_sub lut_3289 ({sk[686], i_14_, i_13_, i_12_, i_15_, n_n191}, x129x);
	defparam lut_3289.LUT_SIZE = 6;
	defparam lut_3289.mask = 64'h0055ffff04440000;

	lut_sub lut_3293 ({sk[687], i_14_, i_13_, i_12_, i_15_, n_n184}, x1731x);
	defparam lut_3293.LUT_SIZE = 6;
	defparam lut_3293.mask = 64'h0055ffff11015154;

	lut_sub lut_3303 ({sk[688], n_n123, n_n125, x52x, x129x, x130x, x1731x}, n_n2813);
	defparam lut_3303.LUT_SIZE = 7;
	defparam lut_3303.mask = 128'h00ff00ffffffffff00005fff77777fff;

	lut_sub lut_3309 ({sk[689], i_14_, i_13_, i_12_, i_15_, n_n191, n_n199}, x1696x);
	defparam lut_3309.LUT_SIZE = 7;
	defparam lut_3309.mask = 128'h00ff00ffffffffff0555505573037370;

	lut_sub lut_3325 ({sk[690], i_14_, i_13_, i_12_, i_15_, n_n216}, x1695x);
	defparam lut_3325.LUT_SIZE = 6;
	defparam lut_3325.mask = 64'h0055ffff15455154;

	lut_sub lut_3338 ({sk[691], n_n124, x735x, n_n126, x74x, x962x, x961x}, x18561x);
	defparam lut_3338.LUT_SIZE = 7;
	defparam lut_3338.mask = 128'h00ff00ffffffffff0000003300005f7f;

	lut_sub lut_3342 ({sk[692], i_7_, i_5_, i_6_, i_3_, i_4_, n_n159}, n_n5319);
	defparam lut_3342.LUT_SIZE = 7;
	defparam lut_3342.mask = 128'h00ff00ffffffffff0000010000000000;

	lut_sub lut_3344 ({sk[693], x132x, n_n197, n_n212, x149x, x147x, x126x}, x18584x);
	defparam lut_3344.LUT_SIZE = 7;
	defparam lut_3344.mask = 128'h00ff00ffffffffff00770f7f00ff0fff;

	lut_sub lut_3349 ({sk[694], x132x, x46x, n_n197, n_n212, x149x, x1856x}, x18585x);
	defparam lut_3349.LUT_SIZE = 7;
	defparam lut_3349.mask = 128'h00ff00ffffffffff035703ff03ff03ff;

	lut_sub lut_3354 ({sk[695], n_n197, n_n212, x55x, x176x, x63x, x48x}, x18589x);
	defparam lut_3354.LUT_SIZE = 7;
	defparam lut_3354.mask = 128'h00ff00ffffffffff00000f0f77ff7fff;

	lut_sub lut_3359 ({sk[696], x735x, n_n200, n_n212, x52x, x130x, x1833x}, x18590x);
	defparam lut_3359.LUT_SIZE = 7;
	defparam lut_3359.mask = 128'h00ff00ffffffffff0077007700770f7f;

	lut_sub lut_3363 ({sk[697], x137x, x46x, n_n197, n_n212, x127x, x129x}, x18591x);
	defparam lut_3363.LUT_SIZE = 7;
	defparam lut_3363.mask = 128'h00ff00ffffffffff00770f7f0f7f0f7f;

	lut_sub lut_3368 ({sk[698], n_n197, n_n212, x123x, x1878x, x131x, x1230x}, x18592x);
	defparam lut_3368.LUT_SIZE = 7;
	defparam lut_3368.mask = 128'h00ff00ffffffffff00000fff77777fff;

	lut_sub lut_3373 ({sk[699], n_n134, x157x, n_n197, n_n212, x186x, x174x}, n_n2760);
	defparam lut_3373.LUT_SIZE = 7;
	defparam lut_3373.mask = 128'h00ff00ffffffffff03570f5f03ff0fff;

	lut_sub lut_3378 ({sk[700], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1654x);
	defparam lut_3378.LUT_SIZE = 7;
	defparam lut_3378.mask = 128'h00ff00ffffffffff7000070000700007;

	lut_sub lut_3387 ({sk[701], n_n135, n_n134, n_n212, x209x, x217x, x174x}, x3143x);
	defparam lut_3387.LUT_SIZE = 7;
	defparam lut_3387.mask = 128'h00ff00ffffffffff007f00ff00ff00ff;

	lut_sub lut_3393 ({sk[702], n_n197, n_n63, x125x, x4792x, x704x, x153x}, x18602x);
	defparam lut_3393.LUT_SIZE = 7;
	defparam lut_3393.mask = 128'h00ff00ffffffffff3f3f3f3f7fffffff;

	lut_sub lut_3399 ({sk[703], n_n197, n_n212, x125x, x176x, x1653x, x1652x}, x18603x);
	defparam lut_3399.LUT_SIZE = 7;
	defparam lut_3399.mask = 128'h00ff00ffffffffff000033ff5f5f7fff;

	lut_sub lut_3404 ({sk[704], x735x, n_n200, n_n212, x55x, x158x, x1849x}, x18607x);
	defparam lut_3404.LUT_SIZE = 7;
	defparam lut_3404.mask = 128'h00ff00ffffffffff003f003f003f557f;

	lut_sub lut_3408 ({sk[705], n_n197, n_n212, x133x, x127x, x158x, x123x}, x18608x);
	defparam lut_3408.LUT_SIZE = 7;
	defparam lut_3408.mask = 128'h00ff00ffffffffff00000fff77ff7fff;

	lut_sub lut_3414 ({sk[706], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x774x);
	defparam lut_3414.LUT_SIZE = 7;
	defparam lut_3414.mask = 128'h00ff00ffffffffff7000070000700007;

	lut_sub lut_3423 ({sk[707], i_7_, i_8_, i_6_, x734x}, n_n101);
	defparam lut_3423.LUT_SIZE = 5;
	defparam lut_3423.mask = 32'h57571000;

	lut_sub lut_3425 ({sk[708], i_7_, i_8_, i_6_, x734x}, n_n42);
	defparam lut_3425.LUT_SIZE = 5;
	defparam lut_3425.mask = 32'h57570010;

	lut_sub lut_3427 ({sk[709], i_7_, i_5_, i_6_, i_3_, i_4_, x714x}, n_n43);
	defparam lut_3427.LUT_SIZE = 7;
	defparam lut_3427.mask = 128'h00ff00ffffffffff0000000000000040;

	lut_sub lut_3429 ({sk[710], i_14_, i_13_, i_12_, i_15_, n_n184}, x139x);
	defparam lut_3429.LUT_SIZE = 6;
	defparam lut_3429.mask = 64'h0055ffff11010000;

	lut_sub lut_3433 ({sk[711], i_9_, i_10_, i_11_, i_15_, n_n211}, n_n182);
	defparam lut_3433.LUT_SIZE = 6;
	defparam lut_3433.mask = 64'h0055ffff10000000;

	lut_sub lut_3435 ({sk[712], i_14_, i_13_, i_12_, i_15_, n_n184}, x54x);
	defparam lut_3435.LUT_SIZE = 6;
	defparam lut_3435.mask = 64'h0055ffff00000110;

	lut_sub lut_3438 ({sk[713], n_n42, n_n43, x130x, x139x, n_n182, x54x}, x18627x);
	defparam lut_3438.LUT_SIZE = 7;
	defparam lut_3438.mask = 128'h00ff00ffffffffff00000f0f7fff7fff;

	lut_sub lut_3444 ({sk[714], i_14_, i_13_, i_12_, i_15_, n_n184}, x128x);
	defparam lut_3444.LUT_SIZE = 6;
	defparam lut_3444.mask = 64'h0055ffff00004044;

	lut_sub lut_3448 ({sk[715], x124x, n_n42, n_n43, x52x, x129x, x128x}, x18628x);
	defparam lut_3448.LUT_SIZE = 7;
	defparam lut_3448.mask = 128'h00ff00ffffffffff007f557f00ff55ff;

	lut_sub lut_3454 ({sk[716], i_9_, i_10_, i_11_, x725x, n_n43}, x524x);
	defparam lut_3454.LUT_SIZE = 6;
	defparam lut_3454.mask = 64'h0055ffff00001000;

	lut_sub lut_3456 ({sk[717], i_14_, i_13_, i_12_, i_15_, n_n184}, x256x);
	defparam lut_3456.LUT_SIZE = 6;
	defparam lut_3456.mask = 64'h0055ffff40100000;

	lut_sub lut_3459 ({sk[718], i_14_, i_13_, i_12_, i_15_, n_n184}, x216x);
	defparam lut_3459.LUT_SIZE = 6;
	defparam lut_3459.mask = 64'h0055ffff00000401;

	lut_sub lut_3462 ({sk[719], n_n42, x63x, x48x, x524x, x256x, x216x}, x18631x);
	defparam lut_3462.LUT_SIZE = 7;
	defparam lut_3462.mask = 128'h00ff00ffffffffff0f0f0f0f7fffffff;

	lut_sub lut_3468 ({sk[720], i_14_, i_13_, i_12_, i_15_, n_n184}, x940x);
	defparam lut_3468.LUT_SIZE = 6;
	defparam lut_3468.mask = 64'h0055ffff44540401;

	lut_sub lut_3476 ({sk[721], i_14_, i_13_, i_12_, i_15_, n_n191}, x222x);
	defparam lut_3476.LUT_SIZE = 6;
	defparam lut_3476.mask = 64'h0055ffff00100401;

	lut_sub lut_3480 ({sk[722], n_n42, n_n43, x52x, x129x, x940x, x222x}, x18632x);
	defparam lut_3480.LUT_SIZE = 7;
	defparam lut_3480.mask = 128'h00ff00ffffffffff000077770fff7fff;

	lut_sub lut_3485 ({sk[723], i_7_, i_8_, i_6_, x734x}, n_n108);
	defparam lut_3485.LUT_SIZE = 5;
	defparam lut_3485.mask = 32'h57570100;

	lut_sub lut_3487 ({sk[724], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1024x);
	defparam lut_3487.LUT_SIZE = 7;
	defparam lut_3487.mask = 128'h00ff00ffffffffff0707007333033330;

	lut_sub lut_3501 ({sk[725], n_n124, x734x, x250x, x224x, x57x, x618x}, x18638x);
	defparam lut_3501.LUT_SIZE = 7;
	defparam lut_3501.mask = 128'h00ff00ffffffffff5555555555557fff;

	lut_sub lut_3506 ({sk[726], n_n101, n_n108, x62x, n_n190, x1690x, x1689x}, n_n4762);
	defparam lut_3506.LUT_SIZE = 7;
	defparam lut_3506.mask = 128'h00ff00ffffffffff000033ff5f5f7fff;

	lut_sub lut_3511 ({sk[727], n_n101, n_n108, n_n169, x69x, x250x, x1860x}, x18680x);
	defparam lut_3511.LUT_SIZE = 7;
	defparam lut_3511.mask = 128'h00ff00ffffffffff000077ff0f0f7fff;

	lut_sub lut_3516 ({sk[728], n_n101, n_n108, n_n169, x208x, x1859x, x1861x}, x18681x);
	defparam lut_3516.LUT_SIZE = 7;
	defparam lut_3516.mask = 128'h00ff00ffffffffff000055553fff7fff;

	lut_sub lut_3521 ({sk[729], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1267x);
	defparam lut_3521.LUT_SIZE = 7;
	defparam lut_3521.mask = 128'h00ff00ffffffffff7000030000300003;

	lut_sub lut_3527 ({sk[730], i_14_, i_13_, i_12_, i_15_, n_n177}, x1266x);
	defparam lut_3527.LUT_SIZE = 6;
	defparam lut_3527.mask = 64'h0055ffff40100401;

	lut_sub lut_3532 ({sk[731], i_7_, i_8_, i_6_, x734x, x1267x, x1266x}, n_n4774);
	defparam lut_3532.LUT_SIZE = 7;
	defparam lut_3532.mask = 128'h00ff00ffffffffff0005000300000000;

	lut_sub lut_3535 ({sk[732], i_14_, i_13_, i_12_, i_15_, n_n191}, x65x);
	defparam lut_3535.LUT_SIZE = 6;
	defparam lut_3535.mask = 64'h0055ffff00100400;

	lut_sub lut_3538 ({sk[733], i_14_, i_13_, i_12_, i_15_, n_n156}, x381x);
	defparam lut_3538.LUT_SIZE = 6;
	defparam lut_3538.mask = 64'h0055ffff40100400;

	lut_sub lut_3542 ({sk[734], i_14_, i_13_, i_12_, i_15_, n_n191}, x1879x);
	defparam lut_3542.LUT_SIZE = 6;
	defparam lut_3542.mask = 64'h0055ffff00005154;

	lut_sub lut_3549 ({sk[735], n_n33, x3461x, x18300x, n_n59, x3011x, x3012x}, x18749x);
	defparam lut_3549.LUT_SIZE = 7;
	defparam lut_3549.mask = 128'h00ff00ffffffffff77ffffff7fffffff;

	lut_sub lut_3555 ({sk[736], i_14_, i_13_, i_12_, i_15_, n_n199}, x865x);
	defparam lut_3555.LUT_SIZE = 6;
	defparam lut_3555.mask = 64'h0055ffff15455154;

	lut_sub lut_3568 ({sk[737], n_n31, n_n30, x788x, n_n102, x98x, x864x}, x18755x);
	defparam lut_3568.LUT_SIZE = 7;
	defparam lut_3568.mask = 128'h00ff00ffffffffff00005fff33337fff;

	lut_sub lut_3573 ({sk[738], n_n31, n_n30, x861x, x860x, x863x, x862x}, x21365x);
	defparam lut_3573.LUT_SIZE = 7;
	defparam lut_3573.mask = 128'h00ff00ffffffffffffffa0a0cc008000;

	lut_sub lut_3578 ({sk[739], x734x, n_n200, n_n32, x1417x, n_n2733, x1887x}, x18761x);
	defparam lut_3578.LUT_SIZE = 7;
	defparam lut_3578.mask = 128'h00ff00ffffffffff333f333f333f777f;

	lut_sub lut_3582 ({sk[740], x734x, n_n200, n_n32, x130x, x48x, x1543x}, x18762x);
	defparam lut_3582.LUT_SIZE = 7;
	defparam lut_3582.mask = 128'h00ff00ffffffffff000f000f000f777f;

	lut_sub lut_3586 ({sk[741], n_n33, n_n32, x124x, n_n101, x381x, x937x}, x18766x);
	defparam lut_3586.LUT_SIZE = 7;
	defparam lut_3586.mask = 128'h00ff00ffffffffff030303ff575757ff;

	lut_sub lut_3590 ({sk[742], n_n124, x734x, n_n126, n_n4774, x1265x, x1264x}, x18767x);
	defparam lut_3590.LUT_SIZE = 7;
	defparam lut_3590.mask = 128'h00ff00ffffffffff0f0f0f5f0f0f3f7f;

	lut_sub lut_3594 ({sk[743], n_n33, n_n32, x1858x, x1848x, x1850x, x1883x}, x18768x);
	defparam lut_3594.LUT_SIZE = 7;
	defparam lut_3594.mask = 128'h00ff00ffffffffff000055553fff7fff;

	lut_sub lut_3599 ({sk[744], i_14_, i_13_, i_12_, i_15_, n_n156, n_n199}, x1021x);
	defparam lut_3599.LUT_SIZE = 7;
	defparam lut_3599.mask = 128'h00ff00ffffffffff5333353330500005;

	lut_sub lut_3611 ({sk[745], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1020x);
	defparam lut_3611.LUT_SIZE = 7;
	defparam lut_3611.mask = 128'h00ff00ffffffffff7000070000700007;

	lut_sub lut_3620 ({sk[746], n_n31, n_n30, x172x, n_n191, x719x, x1873x}, x18776x);
	defparam lut_3620.LUT_SIZE = 7;
	defparam lut_3620.mask = 128'h00ff00ffffffffff0000555503ff57ff;

	lut_sub lut_3624 ({sk[747], n_n65, n_n31, n_n30, x115x, x1095x, x1161x}, x18788x);
	defparam lut_3624.LUT_SIZE = 7;
	defparam lut_3624.mask = 128'h00ff00ffffffffff00553f7f0055ffff;

	lut_sub lut_3629 ({sk[748], n_n156, n_n31, n_n30, x719x, x728x, x1872x}, x646x);
	defparam lut_3629.LUT_SIZE = 7;
	defparam lut_3629.mask = 128'h00ff00ffffffffff00005555003f557f;

	lut_sub lut_3633 ({sk[749], n_n30, x725x, n_n138, n_n184, x18782x, x186x}, x2977x);
	defparam lut_3633.LUT_SIZE = 7;
	defparam lut_3633.mask = 128'h00ff00ffffffffff0000000077ff7fff;

	lut_sub lut_3638 ({sk[750], n_n31, n_n30, x172x, x1022x, x209x, x1263x}, x18783x);
	defparam lut_3638.LUT_SIZE = 7;
	defparam lut_3638.mask = 128'h00ff00ffffffffff000033ff5f5f7fff;

	lut_sub lut_3643 ({sk[751], n_n31, n_n30, n_n128, x122x, x144x, x1163x}, x18786x);
	defparam lut_3643.LUT_SIZE = 7;
	defparam lut_3643.mask = 128'h00ff00ffffffffff000055ff3f3f7fff;

	lut_sub lut_3648 ({sk[752], i_14_, i_13_, i_12_, i_15_, n_n149}, x1096x);
	defparam lut_3648.LUT_SIZE = 6;
	defparam lut_3648.mask = 64'h0055ffff15455044;

	lut_sub lut_3659 ({sk[753], i_7_, i_8_, i_6_, n_n156, x285x}, x419x);
	defparam lut_3659.LUT_SIZE = 6;
	defparam lut_3659.mask = 64'h0055ffff00000010;

	lut_sub lut_3661 ({sk[754], i_7_, i_8_, i_6_, n_n177, x285x}, x445x);
	defparam lut_3661.LUT_SIZE = 6;
	defparam lut_3661.mask = 64'h0055ffff00000010;

	lut_sub lut_3663 ({sk[755], i_7_, i_8_, i_6_, n_n170, x285x}, x446x);
	defparam lut_3663.LUT_SIZE = 6;
	defparam lut_3663.mask = 64'h0055ffff00001000;

	lut_sub lut_3665 ({sk[756], i_9_, i_10_, i_8_, i_11_, n_n17, x285x}, x448x);
	defparam lut_3665.LUT_SIZE = 7;
	defparam lut_3665.mask = 128'h00ff00ffffffffff0001000001000000;

	lut_sub lut_3668 ({sk[757], i_9_, i_10_, i_8_, i_11_, n_n17, x285x}, x450x);
	defparam lut_3668.LUT_SIZE = 7;
	defparam lut_3668.mask = 128'h00ff00ffffffffff0000001000001000;

	lut_sub lut_3671 ({sk[758], i_7_, i_8_, i_6_, n_n177, n_n170, x285x}, x602x);
	defparam lut_3671.LUT_SIZE = 7;
	defparam lut_3671.mask = 128'h00ff00ffffffffff0005001100000000;

	lut_sub lut_3674 ({sk[759], i_7_, i_8_, i_6_, n_n149, n_n156, x285x}, x603x);
	defparam lut_3674.LUT_SIZE = 7;
	defparam lut_3674.mask = 128'h00ff00ffffffffff0005001100000000;

	lut_sub lut_3677 ({sk[760], i_14_, i_13_, i_12_, i_15_, n_n156}, x95x);
	defparam lut_3677.LUT_SIZE = 6;
	defparam lut_3677.mask = 64'h0055ffff10004000;

	lut_sub lut_3680 ({sk[761], i_7_, i_8_, i_6_, n_n9, x288x, x750x}, x786x);
	defparam lut_3680.LUT_SIZE = 7;
	defparam lut_3680.mask = 128'h00ff00ffffffffff5f3f0f0f0f0f0f0f;

	lut_sub lut_3684 ({sk[762], n_n124, x288x, n_n4, x750x, n_n3, x787x}, x21364x);
	defparam lut_3684.LUT_SIZE = 7;
	defparam lut_3684.mask = 128'h00ff00ffffffffff8800880080000000;

	lut_sub lut_3687 ({sk[763], i_14_, i_13_, i_12_, i_15_, n_n41, n_n177}, n_n5060);
	defparam lut_3687.LUT_SIZE = 7;
	defparam lut_3687.mask = 128'h00ff00ffffffffff0000010000100001;

	lut_sub lut_3691 ({sk[764], i_9_, i_10_, i_11_, x725x, x714x, x17002x}, x461x);
	defparam lut_3691.LUT_SIZE = 7;
	defparam lut_3691.mask = 128'h00ff00ffffffffff0000000000010000;

	lut_sub lut_3693 ({sk[765], i_7_, i_8_, i_6_, x740x, x209x}, x4906x);
	defparam lut_3693.LUT_SIZE = 6;
	defparam lut_3693.mask = 64'h0055ffff00001000;

	lut_sub lut_3695 ({sk[766], i_7_, i_8_, i_6_, x740x, x186x}, x4902x);
	defparam lut_3695.LUT_SIZE = 6;
	defparam lut_3695.mask = 64'h0055ffff00001000;

	lut_sub lut_3697 ({sk[767], i_15_, x714x, x17002x, n_n170, n_n209}, x4903x);
	defparam lut_3697.LUT_SIZE = 6;
	defparam lut_3697.mask = 64'h0055ffff00000001;

	lut_sub lut_3699 ({sk[768], x18832x, n_n1843, x18841x, x18845x, x21363x}, n_n1797);
	defparam lut_3699.LUT_SIZE = 6;
	defparam lut_3699.mask = 64'h0055ffffbfffffff;

	lut_sub lut_3705 ({sk[769], n_n31, n_n33, n_n137, x2918x, x197x, x1467x}, n_n1855);
	defparam lut_3705.LUT_SIZE = 7;
	defparam lut_3705.mask = 128'h00ff00ffffffffff0f0f5fff3f3f7fff;

	lut_sub lut_3710 ({sk[770], n_n31, n_n30, n_n102, x56x, x1487x, x1485x}, x19032x);
	defparam lut_3710.LUT_SIZE = 7;
	defparam lut_3710.mask = 128'h00ff00ffffffffff000055553fff7fff;

	lut_sub lut_3715 ({sk[771], n_n33, x318x, n_n1811, n_n1857, x18825x, x18827x}, x19034x);
	defparam lut_3715.LUT_SIZE = 7;
	defparam lut_3715.mask = 128'h00ff00ffffffffff5fff5fff7fffffff;

	lut_sub lut_3721 ({sk[772], n_n71, n_n34, x155x, x19042x, x49x, x92x}, x2700x);
	defparam lut_3721.LUT_SIZE = 7;
	defparam lut_3721.mask = 128'h00ff00ffffffffff00007fff0000ffff;

	lut_sub lut_3727 ({sk[773], n_n34, x133x, x127x, x2697x, x614x, x847x}, x19050x);
	defparam lut_3727.LUT_SIZE = 7;
	defparam lut_3727.mask = 128'h00ff00ffffffffff3f3f3f3f7fffffff;

	lut_sub lut_3733 ({sk[774], i_14_, i_13_, i_12_, i_15_, n_n149, n_n170}, x851x);
	defparam lut_3733.LUT_SIZE = 7;
	defparam lut_3733.mask = 128'h00ff00ffffffffff0555500550075750;

	lut_sub lut_3746 ({sk[775], n_n36, n_n127, x2690x, n_n52, x1208x, x2684x}, x19055x);
	defparam lut_3746.LUT_SIZE = 7;
	defparam lut_3746.mask = 128'h00ff00ffffffffff55ff55ff7fffffff;

	lut_sub lut_3752 ({sk[776], n_n36, x2702x, x845x, x848x, x1144x}, x21349x);
	defparam lut_3752.LUT_SIZE = 6;
	defparam lut_3752.mask = 64'h0055ffffff008000;

	lut_sub lut_3755 ({sk[777], n_n33, x2700x, x19050x, x851x, x19055x, x21349x}, n_n1146);
	defparam lut_3755.LUT_SIZE = 7;
	defparam lut_3755.mask = 128'h00ff00ffffffffffbbffffffbfffffff;

	lut_sub lut_3761 ({sk[778], n_n46, n_n43, n_n137, x72x, x378x, x1501x}, x19108x);
	defparam lut_3761.LUT_SIZE = 7;
	defparam lut_3761.mask = 128'h00ff00ffffffffff000055553fff7fff;

	lut_sub lut_3766 ({sk[779], n_n6267, x2643x, x2638x, x2642x, x19106x}, x19109x);
	defparam lut_3766.LUT_SIZE = 6;
	defparam lut_3766.mask = 64'h0055ffff7fffffff;

	lut_sub lut_3772 ({sk[780], x740x, n_n161, n_n155, x1554x, x2630x, x21439x}, x19118x);
	defparam lut_3772.LUT_SIZE = 7;
	defparam lut_3772.mask = 128'h00ff00ffffffffffbbbbbbbbbbbbbfff;

	lut_sub lut_3777 ({sk[781], x729x, n_n149, n_n46, n_n47, x118x, x1888x}, x19122x);
	defparam lut_3777.LUT_SIZE = 7;
	defparam lut_3777.mask = 128'h00ff00ffffffffff07070707070707ff;

	lut_sub lut_3781 ({sk[782], n_n46, n_n47, x1436x, x852x, x19115x, x19116x}, x21354x);
	defparam lut_3781.LUT_SIZE = 7;
	defparam lut_3781.mask = 128'h00ff00ffffffffffffffff0080808000;

	lut_sub lut_3786 ({sk[783], x19108x, x19109x, x19118x, x19122x, x21354x}, x19126x);
	defparam lut_3786.LUT_SIZE = 6;
	defparam lut_3786.mask = 64'h0055ffffbfffffff;

	lut_sub lut_3792 ({sk[784], x19062x, x19069x, x19074x, x21353x}, n_n1150);
	defparam lut_3792.LUT_SIZE = 5;
	defparam lut_3792.mask = 32'h57577fff;

	lut_sub lut_3797 ({sk[785], n_n41, n_n40, n_n4620, n_n6384, x1158x, x1157x}, x19097x);
	defparam lut_3797.LUT_SIZE = 7;
	defparam lut_3797.mask = 128'h00ff00ffffffffff0fff3fff5fff7fff;

	lut_sub lut_3802 ({sk[786], x19083x, x19089x, x19090x, n_n1294, x19082x}, x19098x);
	defparam lut_3802.LUT_SIZE = 6;
	defparam lut_3802.mask = 64'h0055ffff7fffffff;

	lut_sub lut_3808 ({sk[787], i_9_, i_10_, i_11_, x729x}, n_n102);
	defparam lut_3808.LUT_SIZE = 5;
	defparam lut_3808.mask = 32'h57570001;

	lut_sub lut_3810 ({sk[788], i_14_, i_13_, i_12_, i_15_, n_n191}, x98x);
	defparam lut_3810.LUT_SIZE = 6;
	defparam lut_3810.mask = 64'h0055ffff00000110;

	lut_sub lut_3813 ({sk[789], i_14_, i_13_, i_12_, i_15_, n_n191, n_n199}, x926x);
	defparam lut_3813.LUT_SIZE = 7;
	defparam lut_3813.mask = 128'h00ff00ffffffffff0555500570057570;

	lut_sub lut_3827 ({sk[790], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x925x);
	defparam lut_3827.LUT_SIZE = 7;
	defparam lut_3827.mask = 128'h00ff00ffffffffff0575300550055550;

	lut_sub lut_3839 ({sk[791], n_n31, n_n30, n_n102, x98x, x926x, x925x}, x19146x);
	defparam lut_3839.LUT_SIZE = 7;
	defparam lut_3839.mask = 128'h00ff00ffffffffff000055ff3f3f7fff;

	lut_sub lut_3844 ({sk[792], n_n33, n_n52, n_n137, x2918x, x1288x, x2619x}, n_n1240);
	defparam lut_3844.LUT_SIZE = 7;
	defparam lut_3844.mask = 128'h00ff00ffffffffff5f5f5f5f7fffffff;

	lut_sub lut_3850 ({sk[793], i_14_, i_13_, i_12_, i_15_, n_n216}, x922x);
	defparam lut_3850.LUT_SIZE = 6;
	defparam lut_3850.mask = 64'h0055ffff15014154;

	lut_sub lut_3860 ({sk[794], n_n31, n_n30, x74x, n_n102, x68x, x81x}, x19133x);
	defparam lut_3860.LUT_SIZE = 7;
	defparam lut_3860.mask = 128'h00ff00ffffffffff000077ff0f0f7fff;

	lut_sub lut_3865 ({sk[795], n_n33, n_n32, x60x, x1848x, x924x, x923x}, n_n1170);
	defparam lut_3865.LUT_SIZE = 7;
	defparam lut_3865.mask = 128'h00ff00ffffffffff000033335fff7fff;

	lut_sub lut_3870 ({sk[796], n_n31, x19146x, n_n1240, x922x, x19133x, n_n1170}, n_n1145);
	defparam lut_3870.LUT_SIZE = 7;
	defparam lut_3870.mask = 128'h00ff00ffffffffff77ffffff7fffffff;

	lut_sub lut_3876 ({sk[797], n_n101, n_n1199, x997x, x19294x, x19299x, x19300x}, n_n1155);
	defparam lut_3876.LUT_SIZE = 7;
	defparam lut_3876.mask = 128'h00ff00ffffffffff7f7fffff7fffffff;

	lut_sub lut_3882 ({sk[798], n_n46, x70x, n_n47, n_n214, x1897x, x19324x}, x19325x);
	defparam lut_3882.LUT_SIZE = 7;
	defparam lut_3882.mask = 128'h00ff00ffffffffff557755ff5f7f5fff;

	lut_sub lut_3887 ({sk[799], x19309x, x19316x, x19317x, n_n1320, x19308x}, x19326x);
	defparam lut_3887.LUT_SIZE = 6;
	defparam lut_3887.mask = 64'h0055ffff7fffffff;

	lut_sub lut_3893 ({sk[800], n_n46, x19332x, n_n1194, x1507x, x19343x, x19344x}, n_n1153);
	defparam lut_3893.LUT_SIZE = 7;
	defparam lut_3893.mask = 128'h00ff00ffffffffff77ffffff7fffffff;

	lut_sub lut_3899 ({sk[801], n_n125, x19163x, x19164x, n_n1209, x920x, x19176x}, n_n1158);
	defparam lut_3899.LUT_SIZE = 7;
	defparam lut_3899.mask = 128'h00ff00ffffffffff5fffffff7fffffff;

	lut_sub lut_3905 ({sk[802], n_n108, n_n1201, x19192x, x19193x, x1075x, x19200x}, n_n1156);
	defparam lut_3905.LUT_SIZE = 7;
	defparam lut_3905.mask = 128'h00ff00ffffffffff5fffffff7fffffff;

	lut_sub lut_3911 ({sk[803], x19153x, x19158x, x19207x, x19208x, x21350x}, x19211x);
	defparam lut_3911.LUT_SIZE = 6;
	defparam lut_3911.mask = 64'h0055ffffbfffffff;

	lut_sub lut_3917 ({sk[804], x19233x, x19269x, n_n1217, n_n1216, n_n1214, n_n1213}, x19278x);
	defparam lut_3917.LUT_SIZE = 7;
	defparam lut_3917.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_3924 ({sk[805], n_n123, x74x, x68x, x81x, n_n1366, x19273x}, x19275x);
	defparam lut_3924.LUT_SIZE = 7;
	defparam lut_3924.mask = 128'h00ff00ffffffffff777777777fffffff;

	lut_sub lut_3930 ({sk[806], n_n212, x19240x, x19241x, x19249x, x1256x, x2519x}, x19276x);
	defparam lut_3930.LUT_SIZE = 7;
	defparam lut_3930.mask = 128'h00ff00ffffffffff5fffffff7fffffff;

	lut_sub lut_3936 ({sk[807], x392x, n_n34, x68x, n_n1514, x17542x, x495x}, x19354x);
	defparam lut_3936.LUT_SIZE = 7;
	defparam lut_3936.mask = 128'h00ff00ffffffffff7f7f7fffffffffff;

	lut_sub lut_3942 ({sk[808], n_n36, n_n34, n_n102, x81x, n_n4279, x1001x}, x19355x);
	defparam lut_3942.LUT_SIZE = 7;
	defparam lut_3942.mask = 128'h00ff00ffffffffff33333f3f77ff7fff;

	lut_sub lut_3947 ({sk[809], n_n39, x248x, n_n143, x249x, x647x, x457x}, x19362x);
	defparam lut_3947.LUT_SIZE = 7;
	defparam lut_3947.mask = 128'h00ff00ffffffffff777777777fffffff;

	lut_sub lut_3953 ({sk[810], n_n124, x740x, x207x, x572x, x1002x, x21431x}, x19363x);
	defparam lut_3953.LUT_SIZE = 7;
	defparam lut_3953.mask = 128'h00ff00ffffffffffafafafafafafbfff;

	lut_sub lut_3958 ({sk[811], n_n36, n_n34, x70x, x74x, n_n198, x233x}, x19367x);
	defparam lut_3958.LUT_SIZE = 7;
	defparam lut_3958.mask = 128'h00ff00ffffffffff00005fff33337fff;

	lut_sub lut_3963 ({sk[812], n_n36, n_n34, n_n102, x98x, x1005x, x1066x}, x19368x);
	defparam lut_3963.LUT_SIZE = 7;
	defparam lut_3963.mask = 128'h00ff00ffffffffff000055ff3f3f7fff;

	lut_sub lut_3968 ({sk[813], x19354x, x19355x, x19362x, x19363x, x19367x, x19368x}, n_n1148);
	defparam lut_3968.LUT_SIZE = 7;
	defparam lut_3968.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_3975 ({sk[814], i_9_, i_10_, i_11_, x729x, n_n30}, x3025x);
	defparam lut_3975.LUT_SIZE = 6;
	defparam lut_3975.mask = 64'h0055ffff01000000;

	lut_sub lut_3977 ({sk[815], n_n31, n_n30, n_n117, x98x, x914x, x913x}, n_n1167);
	defparam lut_3977.LUT_SIZE = 7;
	defparam lut_3977.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_3982 ({sk[816], i_14_, i_13_, i_12_, i_15_, n_n170}, x1869x);
	defparam lut_3982.LUT_SIZE = 6;
	defparam lut_3982.mask = 64'h0055ffff11014044;

	lut_sub lut_3989 ({sk[817], n_n31, n_n30, x1007x, x1006x, x1069x, x1068x}, x21348x);
	defparam lut_3989.LUT_SIZE = 7;
	defparam lut_3989.mask = 128'h00ff00ffffffffffffffcc00a0a08000;

	lut_sub lut_3994 ({sk[818], n_n31, x53x, x3025x, n_n1167, x1869x, x21348x}, n_n1144);
	defparam lut_3994.LUT_SIZE = 7;
	defparam lut_3994.mask = 128'h00ff00ffffffffffafffafffbfffffff;

	lut_sub lut_4000 ({sk[819], n_n36, n_n34, x52x, n_n117, x63x, n_n176}, x19395x);
	defparam lut_4000.LUT_SIZE = 7;
	defparam lut_4000.mask = 128'h00ff00ffffffffff000033ff5f5f7fff;

	lut_sub lut_4005 ({sk[820], n_n36, n_n34, n_n184, x720x, x52x, x63x}, x19401x);
	defparam lut_4005.LUT_SIZE = 7;
	defparam lut_4005.mask = 128'h00ff00ffffffffff0000000f7777777f;

	lut_sub lut_4009 ({sk[821], n_n36, n_n34, x147x, n_n176, n_n77, x1080x}, x19406x);
	defparam lut_4009.LUT_SIZE = 7;
	defparam lut_4009.mask = 128'h00ff00ffffffffff00007f7f00ff7fff;

	lut_sub lut_4014 ({sk[822], n_n36, n_n34, x126x, x227x, x1067x, x1081x}, x19407x);
	defparam lut_4014.LUT_SIZE = 7;
	defparam lut_4014.mask = 128'h00ff00ffffffffff000033335fff7fff;

	lut_sub lut_4019 ({sk[823], n_n36, n_n34, x1077x, x1076x, x1079x, x1078x}, x21347x);
	defparam lut_4019.LUT_SIZE = 7;
	defparam lut_4019.mask = 128'h00ff00ffffffffffffffaa00c0c08000;

	lut_sub lut_4024 ({sk[824], x19395x, x19401x, x19406x, x19407x, x21347x}, n_n1147);
	defparam lut_4024.LUT_SIZE = 6;
	defparam lut_4024.mask = 64'h0055ffffbfffffff;

	lut_sub lut_4030 ({sk[825], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1083x);
	defparam lut_4030.LUT_SIZE = 7;
	defparam lut_4030.mask = 128'h00ff00ffffffffff0000000300070330;

	lut_sub lut_4036 ({sk[826], i_14_, i_13_, i_12_, i_15_, n_n170}, x1082x);
	defparam lut_4036.LUT_SIZE = 6;
	defparam lut_4036.mask = 64'h0055ffff00010114;

	lut_sub lut_4041 ({sk[827], x740x, n_n200, x2373x, x2371x, x1403x, x1555x}, x19429x);
	defparam lut_4041.LUT_SIZE = 7;
	defparam lut_4041.mask = 128'h00ff00ffffffffff0fff0fff0fff7fff;

	lut_sub lut_4046 ({sk[828], n_n124, x740x, n_n126, x1083x, x1082x, x19429x}, x19430x);
	defparam lut_4046.LUT_SIZE = 7;
	defparam lut_4046.mask = 128'h00ff00ffffffffff5555555f5555777f;

	lut_sub lut_4050 ({sk[829], x740x, n_n200, x92x, x232x, x19413x, x19414x}, x2380x);
	defparam lut_4050.LUT_SIZE = 7;
	defparam lut_4050.mask = 128'h00ff00ffffffffff0000000000007fff;

	lut_sub lut_4055 ({sk[830], n_n41, n_n40, x155x, x227x, x1210x, x315x}, x19417x);
	defparam lut_4055.LUT_SIZE = 7;
	defparam lut_4055.mask = 128'h00ff00ffffffffff00000fff77777fff;

	lut_sub lut_4060 ({sk[831], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1213x);
	defparam lut_4060.LUT_SIZE = 7;
	defparam lut_4060.mask = 128'h00ff00ffffffffff0507000770057770;

	lut_sub lut_4075 ({sk[832], x729x, n_n156, n_n41, n_n40, x118x, x726x}, x19421x);
	defparam lut_4075.LUT_SIZE = 7;
	defparam lut_4075.mask = 128'h00ff00ffffffffff03030357030303ff;

	lut_sub lut_4079 ({sk[833], n_n41, n_n40, n_n148, x133x, x127x, x60x}, x19422x);
	defparam lut_4079.LUT_SIZE = 7;
	defparam lut_4079.mask = 128'h00ff00ffffffffff00007f7f00ff7fff;

	lut_sub lut_4084 ({sk[834], n_n41, x2380x, x19417x, x1213x, x19421x, x19422x}, x19431x);
	defparam lut_4084.LUT_SIZE = 7;
	defparam lut_4084.mask = 128'h00ff00ffffffffff77ffffff7fffffff;

	lut_sub lut_4090 ({sk[835], n_n71, n_n31, n_n30, x118x, x1505x, x1504x}, n_n1164);
	defparam lut_4090.LUT_SIZE = 7;
	defparam lut_4090.mask = 128'h00ff00ffffffffff005f337f005fffff;

	lut_sub lut_4095 ({sk[836], i_8_, n_n157, x734x, x232x, x19444x, x19443x}, x2357x);
	defparam lut_4095.LUT_SIZE = 7;
	defparam lut_4095.mask = 128'h00ff00ffffffffff0000007f00000000;

	lut_sub lut_4099 ({sk[837], n_n31, n_n30, x1537x, x1536x, x1538x}, x19446x);
	defparam lut_4099.LUT_SIZE = 6;
	defparam lut_4099.mask = 64'h0055ffff00335f7f;

	lut_sub lut_4103 ({sk[838], i_8_, n_n157, n_n31, x734x, x1585x, x1584x}, x19451x);
	defparam lut_4103.LUT_SIZE = 7;
	defparam lut_4103.mask = 128'h00ff00ffffffffff0033053700330033;

	lut_sub lut_4106 ({sk[839], n_n1164, x2357x, x19446x, x19451x}, n_n1143);
	defparam lut_4106.LUT_SIZE = 5;
	defparam lut_4106.mask = 32'h57577fff;

	lut_sub lut_4111 ({sk[840], i_14_, i_13_, i_12_, i_15_, n_n177}, x1300x);
	defparam lut_4111.LUT_SIZE = 6;
	defparam lut_4111.mask = 64'h0055ffff00051114;

	lut_sub lut_4118 ({sk[841], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1299x);
	defparam lut_4118.LUT_SIZE = 7;
	defparam lut_4118.mask = 128'h00ff00ffffffffff0000005000030300;

	lut_sub lut_4122 ({sk[842], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1308x);
	defparam lut_4122.LUT_SIZE = 7;
	defparam lut_4122.mask = 128'h00ff00ffffffffff0000003707070770;

	lut_sub lut_4134 ({sk[843], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1307x);
	defparam lut_4134.LUT_SIZE = 7;
	defparam lut_4134.mask = 128'h00ff00ffffffffff0000007505050550;

	lut_sub lut_4142 ({sk[844], n_n31, n_n30, x1300x, x1299x, x1308x, x1307x}, x19478x);
	defparam lut_4142.LUT_SIZE = 7;
	defparam lut_4142.mask = 128'h00ff00ffffffffff000055ff3f3f7fff;

	lut_sub lut_4147 ({sk[845], i_14_, i_13_, i_12_, i_15_, n_n216}, x111x);
	defparam lut_4147.LUT_SIZE = 6;
	defparam lut_4147.mask = 64'h0055ffff00000110;

	lut_sub lut_4150 ({sk[846], n_n32, n_n184, x719x, x753x, x19480x, x21346x}, n_n799);
	defparam lut_4150.LUT_SIZE = 7;
	defparam lut_4150.mask = 128'h00ff00ffffffffffbfbfbfbfbfbfbfff;

	lut_sub lut_4155 ({sk[847], i_14_, i_13_, i_12_, i_15_, n_n199}, x1810x);
	defparam lut_4155.LUT_SIZE = 6;
	defparam lut_4155.mask = 64'h0055ffff00051114;

	lut_sub lut_4162 ({sk[848], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1809x);
	defparam lut_4162.LUT_SIZE = 7;
	defparam lut_4162.mask = 128'h00ff00ffffffffff0000007707030370;

	lut_sub lut_4173 ({sk[849], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1711x);
	defparam lut_4173.LUT_SIZE = 7;
	defparam lut_4173.mask = 128'h00ff00ffffffffff0000007707050770;

	lut_sub lut_4185 ({sk[850], n_n36, n_n34, x1709x, x1708x, x1707x, x1710x}, x19491x);
	defparam lut_4185.LUT_SIZE = 7;
	defparam lut_4185.mask = 128'h00ff00ffffffffff000033ff7f7f7fff;

	lut_sub lut_4191 ({sk[851], n_n32, n_n182, x54x, x19494x, x21449x}, x19498x);
	defparam lut_4191.LUT_SIZE = 6;
	defparam lut_4191.mask = 64'h0055ffffbbbbbfff;

	lut_sub lut_4196 ({sk[852], x734x, n_n200, n_n32, x165x, x1739x, x2317x}, x19499x);
	defparam lut_4196.LUT_SIZE = 7;
	defparam lut_4196.mask = 128'h00ff00ffffffffff555f555f555f777f;

	lut_sub lut_4200 ({sk[853], n_n817, x19556x, x19557x}, x19559x);
	defparam lut_4200.LUT_SIZE = 4;
	defparam lut_4200.mask = 16'h0f7f;

	lut_sub lut_4204 ({sk[854], x740x, n_n200, n_n138, x19549x, x21412x, x21414x}, x19560x);
	defparam lut_4204.LUT_SIZE = 7;
	defparam lut_4204.mask = 128'h00ff00ffffffffffefefefefefefefff;

	lut_sub lut_4209 ({sk[855], n_n832, n_n767, x19570x, x19574x, x19569x}, n_n746);
	defparam lut_4209.LUT_SIZE = 6;
	defparam lut_4209.mask = 64'h0055ffff7fffffff;

	lut_sub lut_4215 ({sk[856], x19582x, x19583x, n_n834, x19591x, x19596x, x19590x}, n_n747);
	defparam lut_4215.LUT_SIZE = 7;
	defparam lut_4215.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_4222 ({sk[857], n_n772, n_n849, x19611x, x19618x, x2190x}, n_n748);
	defparam lut_4222.LUT_SIZE = 6;
	defparam lut_4222.mask = 64'h0055ffff7fffffff;

	lut_sub lut_4228 ({sk[858], n_n785, x19510x, x19511x, x19516x}, n_n752);
	defparam lut_4228.LUT_SIZE = 5;
	defparam lut_4228.mask = 32'h57577fff;

	lut_sub lut_4233 ({sk[859], n_n34, x1604x, x19527x, x19533x, x21453x}, x19541x);
	defparam lut_4233.LUT_SIZE = 6;
	defparam lut_4233.mask = 64'h0055ffffbfbfbfff;

	lut_sub lut_4238 ({sk[860], x19645x, x19646x, n_n860, x19652x, x19657x, x19651x}, n_n750);
	defparam lut_4238.LUT_SIZE = 7;
	defparam lut_4238.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_4245 ({sk[861], n_n123, n_n781, x19670x, x19671x, x1775x, x19674x}, n_n751);
	defparam lut_4245.LUT_SIZE = 7;
	defparam lut_4245.mask = 128'h00ff00ffffffffff5fffffff7fffffff;

	lut_sub lut_4251 ({sk[862], n_n812, n_n777, n_n813, n_n776, x19637x, x19538x}, x21343x);
	defparam lut_4251.LUT_SIZE = 7;
	defparam lut_4251.mask = 128'h00ff00ffffffffff8000000000000000;

	lut_sub lut_4253 ({sk[863], i_9_, i_10_, i_11_, i_15_, n_n209}, x777x);
	defparam lut_4253.LUT_SIZE = 6;
	defparam lut_4253.mask = 64'h0055ffff00100110;

	lut_sub lut_4257 ({sk[864], i_9_, i_10_, i_11_, i_15_, n_n209}, x406x);
	defparam lut_4257.LUT_SIZE = 6;
	defparam lut_4257.mask = 64'h0055ffff00100100;

	lut_sub lut_4260 ({sk[865], i_9_, i_10_, i_11_, i_15_, n_n209}, x776x);
	defparam lut_4260.LUT_SIZE = 6;
	defparam lut_4260.mask = 64'h0055ffff00101110;

	lut_sub lut_4265 ({sk[866], i_9_, i_10_, i_11_, i_15_, n_n209}, n_n116);
	defparam lut_4265.LUT_SIZE = 6;
	defparam lut_4265.mask = 64'h0055ffff10000000;

	lut_sub lut_4267 ({sk[867], i_9_, i_10_, i_11_, i_15_, n_n209}, x775x);
	defparam lut_4267.LUT_SIZE = 6;
	defparam lut_4267.mask = 64'h0055ffff11000000;

	lut_sub lut_4270 ({sk[868], i_14_, i_13_, i_12_, i_15_, n_n156, n_n191}, x1368x);
	defparam lut_4270.LUT_SIZE = 7;
	defparam lut_4270.mask = 128'h00ff00ffffffffff0700700070000000;

	lut_sub lut_4277 ({sk[869], i_9_, i_10_, i_11_, x725x, x751x}, x2098x);
	defparam lut_4277.LUT_SIZE = 6;
	defparam lut_4277.mask = 64'h0055ffff00101000;

	lut_sub lut_4280 ({sk[870], n_n149, n_n31, n_n3, x728x, x1368x, x2098x}, x19697x);
	defparam lut_4280.LUT_SIZE = 7;
	defparam lut_4280.mask = 128'h00ff00ffffffffff5577557755775f7f;

	lut_sub lut_4284 ({sk[871], i_9_, i_10_, i_11_, x728x}, n_n136);
	defparam lut_4284.LUT_SIZE = 5;
	defparam lut_4284.mask = 32'h57574000;

	lut_sub lut_4286 ({sk[872], i_9_, i_10_, i_11_, x728x}, n_n56);
	defparam lut_4286.LUT_SIZE = 5;
	defparam lut_4286.mask = 32'h57571000;

	lut_sub lut_4288 ({sk[873], i_9_, i_10_, i_11_, n_n31, x728x}, x2109x);
	defparam lut_4288.LUT_SIZE = 6;
	defparam lut_4288.mask = 64'h0055ffff00000110;

	lut_sub lut_4291 ({sk[874], i_7_, i_6_, i_1_, i_2_, i_0_, n_n48}, x19694x);
	defparam lut_4291.LUT_SIZE = 7;
	defparam lut_4291.mask = 128'h00ff00ffffffffff1100110011001000;

	lut_sub lut_4299 ({sk[875], i_9_, i_10_, i_11_, n_n30, n_n7242, x728x}, x21337x);
	defparam lut_4299.LUT_SIZE = 7;
	defparam lut_4299.mask = 128'h00ff00ffffffffffccccc8ccc8c8c8cc;

	lut_sub lut_4305 ({sk[876], x213x, n_n136, n_n56, x2109x, x19694x, x21337x}, x19698x);
	defparam lut_4305.LUT_SIZE = 7;
	defparam lut_4305.mask = 128'h00ff00ffffffffffbfbfbfbfbfffffff;

	lut_sub lut_4311 ({sk[877], x2084x, x19712x, n_n371, x19736x}, x19738x);
	defparam lut_4311.LUT_SIZE = 5;
	defparam lut_4311.mask = 32'h57577fff;

	lut_sub lut_4316 ({sk[878], n_n367, x19721x, x19732x, x19733x, x19720x}, x19739x);
	defparam lut_4316.LUT_SIZE = 6;
	defparam lut_4316.mask = 64'h0055ffff7fffffff;

	lut_sub lut_4322 ({sk[879], n_n40, n_n6384, x2051x, x1619x, x19755x, x1684x}, x19757x);
	defparam lut_4322.LUT_SIZE = 7;
	defparam lut_4322.mask = 128'h00ff00ffffffffff00ffffff7fffffff;

	lut_sub lut_4328 ({sk[880], n_n41, n_n171, x19751x, x1617x, n_n388, x19750x}, x19758x);
	defparam lut_4328.LUT_SIZE = 7;
	defparam lut_4328.mask = 128'h00ff00ffffffffff77ff77ff7fffffff;

	lut_sub lut_4334 ({sk[881], n_n373, n_n374, n_n319, x19709x, x19710x, x19864x}, x19868x);
	defparam lut_4334.LUT_SIZE = 7;
	defparam lut_4334.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_4341 ({sk[882], n_n197, n_n212, x166x, n_n339, n_n338, x1366x}, n_n306);
	defparam lut_4341.LUT_SIZE = 7;
	defparam lut_4341.mask = 128'h00ff00ffffffffff3f3f7fff7f7f7fff;

	lut_sub lut_4347 ({sk[883], n_n390, x2017x, x19799x, x19807x, x19806x, x19811x}, n_n301);
	defparam lut_4347.LUT_SIZE = 7;
	defparam lut_4347.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_4354 ({sk[884], x19859x, x19846x, x19847x, x19854x, x19855x}, n_n304);
	defparam lut_4354.LUT_SIZE = 6;
	defparam lut_4354.mask = 64'h0055ffff7fffffff;

	lut_sub lut_4360 ({sk[885], x19829x, x1968x, x19834x, x19837x, x21331x}, n_n305);
	defparam lut_4360.LUT_SIZE = 6;
	defparam lut_4360.mask = 64'h0055ffffbfffffff;

	lut_sub lut_4366 ({sk[886], n_n330, n_n331, x19776x}, n_n303);
	defparam lut_4366.LUT_SIZE = 4;
	defparam lut_4366.mask = 16'h0f7f;

	lut_sub lut_4370 ({sk[887], n_n406, x19786x, x2026x, x21329x}, n_n302);
	defparam lut_4370.LUT_SIZE = 5;
	defparam lut_4370.mask = 32'h5757bfff;

	lut_sub lut_4375 ({sk[888], n_n33, n_n32, n_n52, n_n136, x1219x, x1911x}, n_n356);
	defparam lut_4375.LUT_SIZE = 7;
	defparam lut_4375.mask = 128'h00ff00ffffffffff55555f5f77ff7fff;

	lut_sub lut_4380 ({sk[889], n_n33, x166x, x235x, x236x, x282x, x283x}, x1916x);
	defparam lut_4380.LUT_SIZE = 7;
	defparam lut_4380.mask = 128'h00ff00ffffffffff000000007fffffff;

	lut_sub lut_4386 ({sk[890], n_n36, n_n32, n_n56, x269x, x275x, x21341x}, x19878x);
	defparam lut_4386.LUT_SIZE = 7;
	defparam lut_4386.mask = 128'h00ff00ffffffffff55557f7f55ff7fff;

	lut_sub lut_4391 ({sk[891], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1567x);
	defparam lut_4391.LUT_SIZE = 7;
	defparam lut_4391.mask = 128'h00ff00ffffffffff0033000030073070;

	lut_sub lut_4400 ({sk[892], i_7_, i_6_, n_n162, x714x, x1568x}, x1908x);
	defparam lut_4400.LUT_SIZE = 6;
	defparam lut_4400.mask = 64'h0055ffff01000000;

	lut_sub lut_4402 ({sk[893], n_n31, n_n170, x726x, x110x, x1484x}, x516x);
	defparam lut_4402.LUT_SIZE = 6;
	defparam lut_4402.mask = 64'h0055ffff0000777f;

	lut_sub lut_4406 ({sk[894], n_n31, n_n30, x161x, x329x, x1484x, x21339x}, x19898x);
	defparam lut_4406.LUT_SIZE = 7;
	defparam lut_4406.mask = 128'h00ff00ffffffffff0000bbbb0fffbfff;

	lut_sub lut_4411 ({sk[895], n_n31, n_n30, x1590x, x1589x, x1722x, x1721x}, n_n310);
	defparam lut_4411.LUT_SIZE = 7;
	defparam lut_4411.mask = 128'h00ff00ffffffffff000055ff3f3f7fff;

	lut_sub lut_4416 ({sk[896], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1592x);
	defparam lut_4416.LUT_SIZE = 7;
	defparam lut_4416.mask = 128'h00ff00ffffffffff0077000070037030;

	lut_sub lut_4427 ({sk[897], n_n31, n_n30, x248x, n_n64, x416x, x21338x}, x19907x);
	defparam lut_4427.LUT_SIZE = 7;
	defparam lut_4427.mask = 128'h00ff00ffffffffff0000aaff3f3fbfff;

	lut_sub lut_4432 ({sk[898], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x732x);
	defparam lut_4432.LUT_SIZE = 7;
	defparam lut_4432.mask = 128'h00ff00ffffffffff0000000010000000;

	lut_sub lut_4434 ({sk[899], i_7_, i_8_, i_6_, n_n159, x77x, n_n111}, x454x);
	defparam lut_4434.LUT_SIZE = 7;
	defparam lut_4434.mask = 128'h00ff00ffffffffff0001000000050005;

	lut_sub lut_4437 ({sk[900], i_7_, i_6_, i_1_, i_2_, i_0_, n_n162}, n_n7254);
	defparam lut_4437.LUT_SIZE = 7;
	defparam lut_4437.mask = 128'h00ff00ffffffffff0000100000000000;

	lut_sub lut_4439 ({sk[901], x729x, n_n149, x717x, n_n2, x430x, x730x}, x707x);
	defparam lut_4439.LUT_SIZE = 7;
	defparam lut_4439.mask = 128'h00ff00ffffffffff3333373f33333f3f;

	lut_sub lut_4444 ({sk[902], i_9_, i_10_, i_11_}, n_n199);
	defparam lut_4444.LUT_SIZE = 4;
	defparam lut_4444.mask = 16'h0f10;

	lut_sub lut_4446 ({sk[903], i_14_, i_13_, i_12_, i_15_, n_n199}, x70x);
	defparam lut_4446.LUT_SIZE = 6;
	defparam lut_4446.mask = 64'h0055ffff04400000;

	lut_sub lut_4449 ({sk[904], i_7_, i_8_, i_6_, x740x, x168x}, n_n5118);
	defparam lut_4449.LUT_SIZE = 6;
	defparam lut_4449.mask = 64'h0055ffff00000100;

	lut_sub lut_4451 ({sk[905], i_7_, i_5_, i_6_, i_3_, i_4_}, x17051x);
	defparam lut_4451.LUT_SIZE = 6;
	defparam lut_4451.mask = 64'h0055ffff00000004;

	lut_sub lut_4453 ({sk[906], i_14_, i_13_, i_12_, i_15_, n_n216}, n_n141);
	defparam lut_4453.LUT_SIZE = 6;
	defparam lut_4453.mask = 64'h0055ffff00100000;

	lut_sub lut_4455 ({sk[907], i_9_, i_10_, i_11_, x725x}, n_n63);
	defparam lut_4455.LUT_SIZE = 5;
	defparam lut_4455.mask = 32'h57570001;

	lut_sub lut_4457 ({sk[908], i_14_, i_13_, i_12_, i_15_, n_n46, n_n216}, x4100x);
	defparam lut_4457.LUT_SIZE = 7;
	defparam lut_4457.mask = 128'h00ff00ffffffffff1000010000000000;

	lut_sub lut_4460 ({sk[909], i_14_, i_13_, i_12_, i_15_, n_n149}, x82x);
	defparam lut_4460.LUT_SIZE = 6;
	defparam lut_4460.mask = 64'h0055ffff00100400;

	lut_sub lut_4463 ({sk[910], i_7_, i_8_, i_6_, n_n162, n_n159, n_n48}, x787x);
	defparam lut_4463.LUT_SIZE = 7;
	defparam lut_4463.mask = 128'h00ff00ffffffffff1103000000000000;

	lut_sub lut_4466 ({sk[911], i_14_, i_13_, i_12_, i_15_}, x720x);
	defparam lut_4466.LUT_SIZE = 5;
	defparam lut_4466.mask = 32'h57570010;

	lut_sub lut_4468 ({sk[912], i_9_, i_10_, i_11_, x720x}, n_n148);
	defparam lut_4468.LUT_SIZE = 5;
	defparam lut_4468.mask = 32'h57570400;

	lut_sub lut_4470 ({sk[913], i_14_, i_13_, i_12_, i_15_}, x726x);
	defparam lut_4470.LUT_SIZE = 5;
	defparam lut_4470.mask = 32'h57572000;

	lut_sub lut_4472 ({sk[914], i_9_, i_10_, i_11_, x726x}, n_n150);
	defparam lut_4472.LUT_SIZE = 5;
	defparam lut_4472.mask = 32'h57570004;

	lut_sub lut_4474 ({sk[915], i_14_, i_13_, i_12_, i_15_, n_n156}, x90x);
	defparam lut_4474.LUT_SIZE = 6;
	defparam lut_4474.mask = 64'h0055ffff04400000;

	lut_sub lut_4477 ({sk[916], x729x, n_n156, x734x, n_n126, x726x}, x4331x);
	defparam lut_4477.LUT_SIZE = 6;
	defparam lut_4477.mask = 64'h0055ffff00010003;

	lut_sub lut_4480 ({sk[917], i_7_, i_8_, i_6_, n_n149, x734x, x720x}, x4332x);
	defparam lut_4480.LUT_SIZE = 7;
	defparam lut_4480.mask = 128'h00ff00ffffffffff0001000000000000;

	lut_sub lut_4482 ({sk[918], i_14_, i_13_, i_12_, i_15_, n_n216}, x788x);
	defparam lut_4482.LUT_SIZE = 6;
	defparam lut_4482.mask = 64'h0055ffff15054000;

	lut_sub lut_4489 ({sk[919], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x790x);
	defparam lut_4489.LUT_SIZE = 7;
	defparam lut_4489.mask = 128'h00ff00ffffffffff0333503333033330;

	lut_sub lut_4502 ({sk[920], i_14_, i_13_, i_12_, i_15_, n_n177}, x789x);
	defparam lut_4502.LUT_SIZE = 6;
	defparam lut_4502.mask = 64'h0055ffff15455154;

	lut_sub lut_4515 ({sk[921], i_14_, i_13_, i_12_, i_15_, n_n149}, x118x);
	defparam lut_4515.LUT_SIZE = 6;
	defparam lut_4515.mask = 64'h0055ffff00000110;

	lut_sub lut_4518 ({sk[922], n_n71, n_n31, n_n30, x790x, x789x, x118x}, n_n4855);
	defparam lut_4518.LUT_SIZE = 7;
	defparam lut_4518.mask = 128'h00ff00ffffffffff00770f7f0077ffff;

	lut_sub lut_4523 ({sk[923], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x792x);
	defparam lut_4523.LUT_SIZE = 7;
	defparam lut_4523.mask = 128'h00ff00ffffffffff0337003775055550;

	lut_sub lut_4538 ({sk[924], i_14_, i_13_, i_12_, i_15_, n_n191}, x791x);
	defparam lut_4538.LUT_SIZE = 6;
	defparam lut_4538.mask = 64'h0055ffff15455044;

	lut_sub lut_4549 ({sk[925], i_9_, i_10_, i_11_, x729x}, n_n117);
	defparam lut_4549.LUT_SIZE = 5;
	defparam lut_4549.mask = 32'h57574000;

	lut_sub lut_4551 ({sk[926], n_n31, n_n30, x792x, x791x, n_n117, x98x}, n_n4857);
	defparam lut_4551.LUT_SIZE = 7;
	defparam lut_4551.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_4556 ({sk[927], i_14_, i_13_, i_12_, i_15_, n_n170}, x795x);
	defparam lut_4556.LUT_SIZE = 6;
	defparam lut_4556.mask = 64'h0055ffff15055044;

	lut_sub lut_4566 ({sk[928], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x794x);
	defparam lut_4566.LUT_SIZE = 7;
	defparam lut_4566.mask = 128'h00ff00ffffffffff0775307555005050;

	lut_sub lut_4580 ({sk[929], i_14_, i_13_, i_12_, i_15_, n_n216}, x1818x);
	defparam lut_4580.LUT_SIZE = 6;
	defparam lut_4580.mask = 64'h0055ffff00015054;

	lut_sub lut_4587 ({sk[930], i_14_, i_13_, i_12_, i_15_, n_n216}, x125x);
	defparam lut_4587.LUT_SIZE = 6;
	defparam lut_4587.mask = 64'h0055ffff00100401;

	lut_sub lut_4591 ({sk[931], i_9_, i_10_, i_11_, x720x}, n_n214);
	defparam lut_4591.LUT_SIZE = 5;
	defparam lut_4591.mask = 32'h57570001;

	lut_sub lut_4593 ({sk[932], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x797x);
	defparam lut_4593.LUT_SIZE = 7;
	defparam lut_4593.mask = 128'h00ff00ffffffffff7000070000700007;

	lut_sub lut_4602 ({sk[933], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x796x);
	defparam lut_4602.LUT_SIZE = 7;
	defparam lut_4602.mask = 128'h00ff00ffffffffff7000070000700007;

	lut_sub lut_4611 ({sk[934], n_n197, n_n63, n_n125, x1818x, x125x, n_n214}, x17108x);
	defparam lut_4611.LUT_SIZE = 7;
	defparam lut_4611.mask = 128'h00ff00ffffffffff005f005f337fffff;

	lut_sub lut_4616 ({sk[935], i_8_, n_n17, x735x, n_n212, x797x, x796x}, x17109x);
	defparam lut_4616.LUT_SIZE = 7;
	defparam lut_4616.mask = 128'h00ff00ffffffffff0505053705050505;

	lut_sub lut_4619 ({sk[936], i_14_, i_13_, i_12_, i_15_, n_n149}, x55x);
	defparam lut_4619.LUT_SIZE = 6;
	defparam lut_4619.mask = 64'h0055ffff00001110;

	lut_sub lut_4623 ({sk[937], i_9_, i_10_, i_11_, i_15_, n_n209}, n_n69);
	defparam lut_4623.LUT_SIZE = 6;
	defparam lut_4623.mask = 64'h0055ffff00400000;

	lut_sub lut_4625 ({sk[938], i_14_, i_13_, i_12_, i_15_, n_n149}, x207x);
	defparam lut_4625.LUT_SIZE = 6;
	defparam lut_4625.mask = 64'h0055ffff00000104;

	lut_sub lut_4628 ({sk[939], i_7_, i_8_, i_6_, x740x, x207x}, x4283x);
	defparam lut_4628.LUT_SIZE = 6;
	defparam lut_4628.mask = 64'h0055ffff01000000;

	lut_sub lut_4630 ({sk[940], i_14_, i_13_, i_12_, i_15_, n_n156}, x800x);
	defparam lut_4630.LUT_SIZE = 6;
	defparam lut_4630.mask = 64'h0055ffff15455154;

	lut_sub lut_4643 ({sk[941], i_14_, i_13_, i_12_, i_15_, n_n149, n_n216}, x799x);
	defparam lut_4643.LUT_SIZE = 7;
	defparam lut_4643.mask = 128'h00ff00ffffffffff0050500333033330;

	lut_sub lut_4653 ({sk[942], i_14_, i_13_, i_12_, i_15_, n_n216}, x180x);
	defparam lut_4653.LUT_SIZE = 6;
	defparam lut_4653.mask = 64'h0055ffff11040000;

	lut_sub lut_4657 ({sk[943], i_14_, i_13_, i_12_, i_15_, n_n216}, x142x);
	defparam lut_4657.LUT_SIZE = 6;
	defparam lut_4657.mask = 64'h0055ffff00014040;

	lut_sub lut_4661 ({sk[944], n_n46, n_n47, x800x, x799x, x180x, x142x}, n_n4136);
	defparam lut_4661.LUT_SIZE = 7;
	defparam lut_4661.mask = 128'h00ff00ffffffffff000000ff7f7f7fff;

	lut_sub lut_4666 ({sk[945], i_7_, i_8_, i_6_, x181x, x735x}, n_n4581);
	defparam lut_4666.LUT_SIZE = 6;
	defparam lut_4666.mask = 64'h0055ffff10000000;

	lut_sub lut_4668 ({sk[946], i_14_, i_13_, i_12_, i_15_, n_n156}, x1828x);
	defparam lut_4668.LUT_SIZE = 6;
	defparam lut_4668.mask = 64'h0055ffff00005154;

	lut_sub lut_4675 ({sk[947], i_14_, i_13_, i_12_, i_15_, n_n149}, x158x);
	defparam lut_4675.LUT_SIZE = 6;
	defparam lut_4675.mask = 64'h0055ffff04440000;

	lut_sub lut_4679 ({sk[948], i_14_, i_13_, i_12_, i_15_, n_n156}, x176x);
	defparam lut_4679.LUT_SIZE = 6;
	defparam lut_4679.mask = 64'h0055ffff04440000;

	lut_sub lut_4683 ({sk[949], i_14_, i_13_, i_12_, i_15_, n_n156}, x123x);
	defparam lut_4683.LUT_SIZE = 6;
	defparam lut_4683.mask = 64'h0055ffff11010000;

	lut_sub lut_4687 ({sk[950], i_15_, x735x, n_n126, n_n216, n_n209}, x601x);
	defparam lut_4687.LUT_SIZE = 6;
	defparam lut_4687.mask = 64'h0055ffff00000001;

	lut_sub lut_4689 ({sk[951], i_14_, i_13_, i_12_, i_15_, n_n216}, n_n142);
	defparam lut_4689.LUT_SIZE = 6;
	defparam lut_4689.mask = 64'h0055ffff00000001;

	lut_sub lut_4691 ({sk[952], i_14_, i_13_, i_12_, i_15_, n_n156}, x1172x);
	defparam lut_4691.LUT_SIZE = 6;
	defparam lut_4691.mask = 64'h0055ffff15454040;

	lut_sub lut_4700 ({sk[953], i_7_, i_8_, i_6_, x735x, n_n142, x1172x}, n_n3912);
	defparam lut_4700.LUT_SIZE = 7;
	defparam lut_4700.mask = 128'h00ff00ffffffffff0005000300000000;

	lut_sub lut_4703 ({sk[954], i_14_, i_13_, i_12_, i_15_, n_n216}, x141x);
	defparam lut_4703.LUT_SIZE = 6;
	defparam lut_4703.mask = 64'h0055ffff40100400;

	lut_sub lut_4707 ({sk[955], i_14_, i_13_, i_12_, i_15_, n_n199}, x135x);
	defparam lut_4707.LUT_SIZE = 6;
	defparam lut_4707.mask = 64'h0055ffff00000401;

	lut_sub lut_4710 ({sk[956], i_14_, i_13_, i_12_, i_15_, n_n199}, x1171x);
	defparam lut_4710.LUT_SIZE = 6;
	defparam lut_4710.mask = 64'h0055ffff40100401;

	lut_sub lut_4715 ({sk[957], x157x, n_n123, n_n125, x141x, x135x, x1171x}, x17456x);
	defparam lut_4715.LUT_SIZE = 7;
	defparam lut_4715.mask = 128'h00ff00ffffffffff003f557f00ff55ff;

	lut_sub lut_4720 ({sk[958], i_14_, i_13_, i_12_, i_15_, n_n156}, x155x);
	defparam lut_4720.LUT_SIZE = 6;
	defparam lut_4720.mask = 64'h0055ffff00014040;

	lut_sub lut_4724 ({sk[959], i_14_, i_13_, i_12_, i_15_, n_n216}, x85x);
	defparam lut_4724.LUT_SIZE = 6;
	defparam lut_4724.mask = 64'h0055ffff00001014;

	lut_sub lut_4728 ({sk[960], n_n123, x70x, n_n125, n_n214, x85x, x142x}, n_n4225);
	defparam lut_4728.LUT_SIZE = 7;
	defparam lut_4728.mask = 128'h00ff00ffffffffff000000ff7f7f7fff;

	lut_sub lut_4733 ({sk[961], i_14_, i_13_, i_12_, i_15_, n_n216}, x86x);
	defparam lut_4733.LUT_SIZE = 6;
	defparam lut_4733.mask = 64'h0055ffff04400000;

	lut_sub lut_4736 ({sk[962], i_14_, i_13_, i_12_, i_15_, n_n156}, x1851x);
	defparam lut_4736.LUT_SIZE = 6;
	defparam lut_4736.mask = 64'h0055ffff15440000;

	lut_sub lut_4742 ({sk[963], i_9_, i_10_, i_11_, x720x}, n_n155);
	defparam lut_4742.LUT_SIZE = 5;
	defparam lut_4742.mask = 32'h57570004;

	lut_sub lut_4744 ({sk[964], i_14_, i_13_, i_12_, i_15_, n_n156}, x215x);
	defparam lut_4744.LUT_SIZE = 6;
	defparam lut_4744.mask = 64'h0055ffff00001014;

	lut_sub lut_4748 ({sk[965], n_n123, n_n125, x155x, x180x, n_n155, x215x}, x17461x);
	defparam lut_4748.LUT_SIZE = 7;
	defparam lut_4748.mask = 128'h00ff00ffffffffff000077ff0f0f7fff;

	lut_sub lut_4753 ({sk[966], i_14_, i_13_, i_12_, i_15_, n_n149}, x805x);
	defparam lut_4753.LUT_SIZE = 6;
	defparam lut_4753.mask = 64'h0055ffff11055054;

	lut_sub lut_4763 ({sk[967], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x804x);
	defparam lut_4763.LUT_SIZE = 7;
	defparam lut_4763.mask = 128'h00ff00ffffffffff0303003337053770;

	lut_sub lut_4777 ({sk[968], i_14_, i_13_, i_12_, i_15_, n_n149}, x60x);
	defparam lut_4777.LUT_SIZE = 6;
	defparam lut_4777.mask = 64'h0055ffff04400000;

	lut_sub lut_4780 ({sk[969], n_n124, x735x, n_n126, n_n148, x86x, x1851x}, x17460x);
	defparam lut_4780.LUT_SIZE = 7;
	defparam lut_4780.mask = 128'h00ff00ffffffffff0000005500003f7f;

	lut_sub lut_4784 ({sk[970], n_n123, n_n148, n_n125, x805x, x60x, x153x}, x21420x);
	defparam lut_4784.LUT_SIZE = 7;
	defparam lut_4784.mask = 128'h00ff00ffffffffffff80ff00cc80cc00;

	lut_sub lut_4788 ({sk[971], i_14_, i_13_, i_12_, i_15_, n_n149}, x234x);
	defparam lut_4788.LUT_SIZE = 6;
	defparam lut_4788.mask = 64'h0055ffff00014040;

	lut_sub lut_4792 ({sk[972], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x946x);
	defparam lut_4792.LUT_SIZE = 7;
	defparam lut_4792.mask = 128'h00ff00ffffffffff0303003775007550;

	lut_sub lut_4805 ({sk[973], n_n101, n_n108, n_n148, x60x, x234x, x946x}, x17479x);
	defparam lut_4805.LUT_SIZE = 7;
	defparam lut_4805.mask = 128'h00ff00ffffffffff000033ff5f5f7fff;

	lut_sub lut_4810 ({sk[974], i_9_, i_10_, i_11_, x720x}, n_n198);
	defparam lut_4810.LUT_SIZE = 5;
	defparam lut_4810.mask = 32'h57570100;

	lut_sub lut_4812 ({sk[975], i_14_, i_13_, i_12_, i_15_, n_n216}, x1448x);
	defparam lut_4812.LUT_SIZE = 6;
	defparam lut_4812.mask = 64'h0055ffff15454040;

	lut_sub lut_4821 ({sk[976], i_8_, x740x, n_n18, n_n47, n_n198, x1448x}, n_n4206);
	defparam lut_4821.LUT_SIZE = 7;
	defparam lut_4821.mask = 128'h00ff00ffffffffff0505053705050505;

	lut_sub lut_4824 ({sk[977], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x807x);
	defparam lut_4824.LUT_SIZE = 7;
	defparam lut_4824.mask = 128'h00ff00ffffffffff7000070000500005;

	lut_sub lut_4831 ({sk[978], i_14_, i_13_, i_12_, i_15_, n_n149}, x806x);
	defparam lut_4831.LUT_SIZE = 6;
	defparam lut_4831.mask = 64'h0055ffff40100401;

	lut_sub lut_4836 ({sk[979], i_8_, x734x, n_n16, x450x, x807x, x21432x}, x17484x);
	defparam lut_4836.LUT_SIZE = 7;
	defparam lut_4836.mask = 128'h00ff00ffffffffffafafafbfafafafaf;

	lut_sub lut_4840 ({sk[980], n_n47, n_n108, n_n4206, x85x, x806x, x17484x}, x17486x);
	defparam lut_4840.LUT_SIZE = 7;
	defparam lut_4840.mask = 128'h00ff00ffffffffff55ff77ff5fff7fff;

	lut_sub lut_4845 ({sk[981], n_n101, n_n108, x90x, n_n142, x141x, x598x}, x17472x);
	defparam lut_4845.LUT_SIZE = 7;
	defparam lut_4845.mask = 128'h00ff00ffffffffff55557f7f55ff7fff;

	lut_sub lut_4850 ({sk[982], n_n53, n_n101, n_n108, x218x, x141x, x944x}, x21410x);
	defparam lut_4850.LUT_SIZE = 7;
	defparam lut_4850.mask = 128'h00ff00ffffffffffffff8080ff008000;

	lut_sub lut_4855 ({sk[983], x157x, n_n108, x60x, x4362x, x84x, x220x}, x21436x);
	defparam lut_4855.LUT_SIZE = 7;
	defparam lut_4855.mask = 128'h00ff00fffffffffff0f08000f0f00000;

	lut_sub lut_4858 ({sk[984], x17479x, x17472x, x21410x, x21436x}, x17487x);
	defparam lut_4858.LUT_SIZE = 5;
	defparam lut_4858.mask = 32'h5757efff;

	lut_sub lut_4863 ({sk[985], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1841x);
	defparam lut_4863.LUT_SIZE = 7;
	defparam lut_4863.mask = 128'h00ff00ffffffffff0333303337003770;

	lut_sub lut_4878 ({sk[986], i_14_, i_13_, i_12_, i_15_, n_n199}, x1840x);
	defparam lut_4878.LUT_SIZE = 6;
	defparam lut_4878.mask = 64'h0055ffff11055154;

	lut_sub lut_4889 ({sk[987], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x809x);
	defparam lut_4889.LUT_SIZE = 7;
	defparam lut_4889.mask = 128'h00ff00ffffffffff0737307555005550;

	lut_sub lut_4904 ({sk[988], i_14_, i_13_, i_12_, i_15_, n_n149}, x808x);
	defparam lut_4904.LUT_SIZE = 6;
	defparam lut_4904.mask = 64'h0055ffff11055154;

	lut_sub lut_4915 ({sk[989], i_14_, i_13_, i_12_, i_15_, n_n149}, x84x);
	defparam lut_4915.LUT_SIZE = 6;
	defparam lut_4915.mask = 64'h0055ffff00001014;

	lut_sub lut_4919 ({sk[990], n_n124, x734x, n_n148, x4331x, x86x, x84x}, x17504x);
	defparam lut_4919.LUT_SIZE = 7;
	defparam lut_4919.mask = 128'h00ff00ffffffffff0f0f0f0f0f0f7fff;

	lut_sub lut_4924 ({sk[991], i_14_, i_13_, i_12_, i_15_, n_n216}, x1019x);
	defparam lut_4924.LUT_SIZE = 6;
	defparam lut_4924.mask = 64'h0055ffff11055054;

	lut_sub lut_4934 ({sk[992], i_14_, i_13_, i_12_, i_15_, n_n156}, x867x);
	defparam lut_4934.LUT_SIZE = 6;
	defparam lut_4934.mask = 64'h0055ffff11055154;

	lut_sub lut_4945 ({sk[993], i_7_, i_8_, i_6_, x734x, x1019x, x867x}, x17505x);
	defparam lut_4945.LUT_SIZE = 7;
	defparam lut_4945.mask = 128'h00ff00ffffffffff0003000500000000;

	lut_sub lut_4948 ({sk[994], i_14_, i_13_, i_12_, i_15_, n_n216}, x1104x);
	defparam lut_4948.LUT_SIZE = 6;
	defparam lut_4948.mask = 64'h0055ffff11055054;

	lut_sub lut_4958 ({sk[995], i_9_, i_10_, i_8_, i_11_, n_n18, x285x}, x17506x);
	defparam lut_4958.LUT_SIZE = 7;
	defparam lut_4958.mask = 128'h00ff00ffffffffff0000001000001000;

	lut_sub lut_4961 ({sk[996], i_14_, i_13_, i_12_, i_15_, n_n199}, x219x);
	defparam lut_4961.LUT_SIZE = 6;
	defparam lut_4961.mask = 64'h0055ffff00001014;

	lut_sub lut_4965 ({sk[997], i_14_, i_13_, i_12_, i_15_, n_n199}, x108x);
	defparam lut_4965.LUT_SIZE = 6;
	defparam lut_4965.mask = 64'h0055ffff00014040;

	lut_sub lut_4969 ({sk[998], n_n101, n_n108, x86x, n_n198, x219x, x108x}, n_n4903);
	defparam lut_4969.LUT_SIZE = 7;
	defparam lut_4969.mask = 128'h00ff00ffffffffff000000ff7f7f7fff;

	lut_sub lut_4974 ({sk[999], i_14_, i_13_, i_12_, i_15_, n_n199}, x1844x);
	defparam lut_4974.LUT_SIZE = 6;
	defparam lut_4974.mask = 64'h0055ffff15455154;

	lut_sub lut_4987 ({sk[1000], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1843x);
	defparam lut_4987.LUT_SIZE = 7;
	defparam lut_4987.mask = 128'h00ff00ffffffffff0333303000050000;

	lut_sub lut_4994 ({sk[1001], i_7_, i_8_, i_6_, x734x, x1844x, x1843x}, x544x);
	defparam lut_4994.LUT_SIZE = 7;
	defparam lut_4994.mask = 128'h00ff00ffffffffff0005000300000000;

	lut_sub lut_4997 ({sk[1002], i_7_, i_8_, i_6_, n_n216, x285x}, n_n5739);
	defparam lut_4997.LUT_SIZE = 6;
	defparam lut_4997.mask = 64'h0055ffff00000100;

	lut_sub lut_4999 ({sk[1003], x734x, n_n126, x720x, x17506x, n_n216, x21437x}, x17509x);
	defparam lut_4999.LUT_SIZE = 7;
	defparam lut_4999.mask = 128'h00ff00ffffffffff5f5f5f5f5f5f5f7f;

	lut_sub lut_5003 ({sk[1004], n_n123, n_n108, n_n125, x1104x, x1106x, x1105x}, x17510x);
	defparam lut_5003.LUT_SIZE = 7;
	defparam lut_5003.mask = 128'h00ff00ffffffffff00330f3f55775f7f;

	lut_sub lut_5007 ({sk[1005], x17504x, x17505x, n_n4903, x544x, x17509x, x17510x}, x17514x);
	defparam lut_5007.LUT_SIZE = 7;
	defparam lut_5007.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_5014 ({sk[1006], n_n46, n_n47, n_n155, x60x, x809x, x808x}, x17500x);
	defparam lut_5014.LUT_SIZE = 7;
	defparam lut_5014.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_5019 ({sk[1007], i_14_, i_13_, i_12_}, n_n207);
	defparam lut_5019.LUT_SIZE = 4;
	defparam lut_5019.mask = 16'h0f10;

	lut_sub lut_5021 ({sk[1008], i_9_, i_10_, i_11_, i_15_, n_n207}, n_n72);
	defparam lut_5021.LUT_SIZE = 6;
	defparam lut_5021.mask = 64'h0055ffff00000040;

	lut_sub lut_5023 ({sk[1009], i_14_, i_13_, i_12_, i_15_, n_n191}, x51x);
	defparam lut_5023.LUT_SIZE = 6;
	defparam lut_5023.mask = 64'h0055ffff04400000;

	lut_sub lut_5026 ({sk[1010], i_9_, i_10_, i_11_, i_15_, n_n201}, n_n133);
	defparam lut_5026.LUT_SIZE = 6;
	defparam lut_5026.mask = 64'h0055ffff00000100;

	lut_sub lut_5028 ({sk[1011], i_14_, i_13_, i_12_, i_15_, n_n177}, x80x);
	defparam lut_5028.LUT_SIZE = 6;
	defparam lut_5028.mask = 64'h0055ffff00000401;

	lut_sub lut_5031 ({sk[1012], i_15_, n_n156, x714x, x17002x, n_n57, n_n209}, x17661x);
	defparam lut_5031.LUT_SIZE = 7;
	defparam lut_5031.mask = 128'h00ff00ffffffffff0003000300030007;

	lut_sub lut_5034 ({sk[1013], x740x, n_n200, x80x, n_n5060, x78x, x17661x}, n_n3866);
	defparam lut_5034.LUT_SIZE = 7;
	defparam lut_5034.mask = 128'h00ff00ffffffffff5f5f5f5f5f5f7fff;

	lut_sub lut_5039 ({sk[1014], i_9_, i_10_, i_11_, i_15_, n_n211}, n_n154);
	defparam lut_5039.LUT_SIZE = 6;
	defparam lut_5039.mask = 64'h0055ffff00000010;

	lut_sub lut_5041 ({sk[1015], i_14_, i_13_, i_12_, i_15_, n_n156}, x59x);
	defparam lut_5041.LUT_SIZE = 6;
	defparam lut_5041.mask = 64'h0055ffff00000110;

	lut_sub lut_5044 ({sk[1016], i_14_, i_13_, i_12_, i_15_, n_n156}, x134x);
	defparam lut_5044.LUT_SIZE = 6;
	defparam lut_5044.mask = 64'h0055ffff00001110;

	lut_sub lut_5048 ({sk[1017], i_7_, i_8_, i_6_, x735x, x134x}, n_n4268);
	defparam lut_5048.LUT_SIZE = 6;
	defparam lut_5048.mask = 64'h0055ffff10000000;

	lut_sub lut_5050 ({sk[1018], i_1_, i_2_, i_0_}, n_n19);
	defparam lut_5050.LUT_SIZE = 4;
	defparam lut_5050.mask = 16'h0f10;

	lut_sub lut_5052 ({sk[1019], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x731x);
	defparam lut_5052.LUT_SIZE = 7;
	defparam lut_5052.mask = 128'h00ff00ffffffffff0000000000100000;

	lut_sub lut_5054 ({sk[1020], i_14_, i_13_, i_12_}, n_n213);
	defparam lut_5054.LUT_SIZE = 4;
	defparam lut_5054.mask = 16'h0f02;

	lut_sub lut_5056 ({sk[1021], i_9_, i_10_, i_11_, i_15_, n_n213}, n_n82);
	defparam lut_5056.LUT_SIZE = 6;
	defparam lut_5056.mask = 64'h0055ffff01000000;

	lut_sub lut_5058 ({sk[1022], i_9_, i_10_, i_11_, x720x}, n_n169);
	defparam lut_5058.LUT_SIZE = 5;
	defparam lut_5058.mask = 32'h57571000;

	lut_sub lut_5060 ({sk[1023], i_14_, i_13_, i_12_, i_15_, n_n170}, x812x);
	defparam lut_5060.LUT_SIZE = 6;
	defparam lut_5060.mask = 64'h0055ffff15454000;

	lut_sub lut_5068 ({sk[1024], i_9_, i_10_, i_11_, x729x}, n_n83);
	defparam lut_5068.LUT_SIZE = 5;
	defparam lut_5068.mask = 32'h57570010;

	lut_sub lut_5070 ({sk[1025], i_7_, i_6_, i_1_, i_2_, i_0_, n_n48}, n_n7242);
	defparam lut_5070.LUT_SIZE = 7;
	defparam lut_5070.mask = 128'h00ff00ffffffffff0000000000000100;

	lut_sub lut_5072 ({sk[1026], i_7_, i_8_, i_6_, n_n159, n_n111}, x815x);
	defparam lut_5072.LUT_SIZE = 6;
	defparam lut_5072.mask = 64'h0055ffff11000000;

	lut_sub lut_5075 ({sk[1027], n_n149, n_n6, n_n3, n_n2, x730x, x815x}, x3067x);
	defparam lut_5075.LUT_SIZE = 7;
	defparam lut_5075.mask = 128'h00ff00ffffffffff0000000013333333;

	lut_sub lut_5080 ({sk[1028], i_7_, i_5_, i_6_, i_3_, i_4_, n_n219}, x21407x);
	defparam lut_5080.LUT_SIZE = 7;
	defparam lut_5080.mask = 128'h00ff00ffffffffffffffffffefefafef;

	lut_sub lut_5086 ({sk[1029], i_7_, i_6_}, x231x);
	defparam lut_5086.LUT_SIZE = 3;
	defparam lut_5086.mask = 8'h36;

	lut_sub lut_5089 ({sk[1030], i_5_, i_3_, i_4_, n_n159, n_n124, n_n2}, x1044x);
	defparam lut_5089.LUT_SIZE = 7;
	defparam lut_5089.mask = 128'h00ff00ffffffffff5557555555555555;

	lut_sub lut_5092 ({sk[1031], i_7_, i_5_, i_6_, i_3_, i_4_, n_n19}, x462x);
	defparam lut_5092.LUT_SIZE = 7;
	defparam lut_5092.mask = 128'h00ff00ffffffffff0000000010100000;

	lut_sub lut_5095 ({sk[1032], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x816x);
	defparam lut_5095.LUT_SIZE = 7;
	defparam lut_5095.mask = 128'h00ff00ffffffffff1000000000000008;

	lut_sub lut_5098 ({sk[1033], i_9_, i_10_, i_11_, i_15_, n_n207}, n_n78);
	defparam lut_5098.LUT_SIZE = 6;
	defparam lut_5098.mask = 64'h0055ffff04000000;

	lut_sub lut_5100 ({sk[1034], i_14_, i_13_, i_12_, i_15_, n_n170}, x69x);
	defparam lut_5100.LUT_SIZE = 6;
	defparam lut_5100.mask = 64'h0055ffff04400000;

	lut_sub lut_5103 ({sk[1035], i_14_, i_13_, i_12_, i_15_, n_n184}, x62x);
	defparam lut_5103.LUT_SIZE = 6;
	defparam lut_5103.mask = 64'h0055ffff04400000;

	lut_sub lut_5106 ({sk[1036], i_7_, i_8_, i_6_, x735x, n_n212}, x188x);
	defparam lut_5106.LUT_SIZE = 6;
	defparam lut_5106.mask = 64'h0055ffff55557555;

	lut_sub lut_5109 ({sk[1037], i_14_, i_13_, i_12_, i_15_, n_n216}, x818x);
	defparam lut_5109.LUT_SIZE = 6;
	defparam lut_5109.mask = 64'h0055ffff14045000;

	lut_sub lut_5115 ({sk[1038], i_14_, i_13_, i_12_}, n_n204);
	defparam lut_5115.LUT_SIZE = 4;
	defparam lut_5115.mask = 16'h0f80;

	lut_sub lut_5117 ({sk[1039], i_9_, i_10_, i_11_, i_15_, x725x, n_n204}, x820x);
	defparam lut_5117.LUT_SIZE = 7;
	defparam lut_5117.mask = 128'h00ff00ffffffffff0000005033330000;

	lut_sub lut_5121 ({sk[1040], i_9_, i_10_, i_11_, x725x}, n_n55);
	defparam lut_5121.LUT_SIZE = 5;
	defparam lut_5121.mask = 32'h57571000;

	lut_sub lut_5123 ({sk[1041], i_9_, i_10_, i_11_, x725x, n_n34}, x17307x);
	defparam lut_5123.LUT_SIZE = 6;
	defparam lut_5123.mask = 64'h0055ffff00001001;

	lut_sub lut_5126 ({sk[1042], i_14_, i_13_, i_12_, i_15_, n_n156, n_n199}, x17313x);
	defparam lut_5126.LUT_SIZE = 7;
	defparam lut_5126.mask = 128'h00ff00ffffffffff5330003033000000;

	lut_sub lut_5133 ({sk[1043], i_14_, i_13_, i_12_, i_15_, n_n149}, x115x);
	defparam lut_5133.LUT_SIZE = 6;
	defparam lut_5133.mask = 64'h0055ffff14040000;

	lut_sub lut_5137 ({sk[1044], i_14_, i_13_, i_12_, i_15_, n_n149}, x821x);
	defparam lut_5137.LUT_SIZE = 6;
	defparam lut_5137.mask = 64'h0055ffff14445000;

	lut_sub lut_5144 ({sk[1045], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x825x);
	defparam lut_5144.LUT_SIZE = 7;
	defparam lut_5144.mask = 128'h00ff00ffffffffff0700000077000000;

	lut_sub lut_5151 ({sk[1046], i_14_, i_13_, i_12_, i_15_, n_n177}, x200x);
	defparam lut_5151.LUT_SIZE = 6;
	defparam lut_5151.mask = 64'h0055ffff10005000;

	lut_sub lut_5155 ({sk[1047], n_n46, n_n47, x129x, x130x, x825x, x200x}, n_n2253);
	defparam lut_5155.LUT_SIZE = 7;
	defparam lut_5155.mask = 128'h00ff00ffffffffff00007fff3fff7fff;

	lut_sub lut_5163 ({sk[1048], i_9_, i_10_, i_11_, i_15_, n_n204}, n_n61);
	defparam lut_5163.LUT_SIZE = 6;
	defparam lut_5163.mask = 64'h0055ffff00040000;

	lut_sub lut_5165 ({sk[1049], i_14_, i_13_, i_12_, i_15_, n_n149}, x17183x);
	defparam lut_5165.LUT_SIZE = 6;
	defparam lut_5165.mask = 64'h0055ffff10045000;

	lut_sub lut_5170 ({sk[1050], i_14_, i_13_, i_12_, i_15_, n_n156}, x17182x);
	defparam lut_5170.LUT_SIZE = 6;
	defparam lut_5170.mask = 64'h0055ffff10045000;

	lut_sub lut_5175 ({sk[1051], i_9_, i_10_, i_11_, x725x, n_n101, n_n108}, x21395x);
	defparam lut_5175.LUT_SIZE = 7;
	defparam lut_5175.mask = 128'h00ff00fffffffffffff8fffff8f8faff;

	lut_sub lut_5182 ({sk[1052], n_n135, n_n101, n_n108, x90x, n_n61, x21395x}, x17185x);
	defparam lut_5182.LUT_SIZE = 7;
	defparam lut_5182.mask = 128'h00ff00ffffffffffaabbbfbfaaffffff;

	lut_sub lut_5189 ({sk[1053], n_n101, n_n63, n_n108, x60x, x17183x, x17182x}, x17186x);
	defparam lut_5189.LUT_SIZE = 7;
	defparam lut_5189.mask = 128'h00ff00ffffffffff003f00ff5f7fffff;

	lut_sub lut_5196 ({sk[1054], i_14_, i_13_, i_12_, i_15_, n_n156}, x175x);
	defparam lut_5196.LUT_SIZE = 6;
	defparam lut_5196.mask = 64'h0055ffff00000050;

	lut_sub lut_5199 ({sk[1055], i_14_, i_13_, i_12_, i_15_, n_n156}, x832x);
	defparam lut_5199.LUT_SIZE = 6;
	defparam lut_5199.mask = 64'h0055ffff11010050;

	lut_sub lut_5205 ({sk[1056], i_14_, i_13_, i_12_, i_15_, n_n177}, x146x);
	defparam lut_5205.LUT_SIZE = 6;
	defparam lut_5205.mask = 64'h0055ffff11010000;

	lut_sub lut_5209 ({sk[1057], i_14_, i_13_, i_12_, i_15_, n_n177}, x831x);
	defparam lut_5209.LUT_SIZE = 6;
	defparam lut_5209.mask = 64'h0055ffff11410000;

	lut_sub lut_5214 ({sk[1058], i_14_, i_13_, i_12_, i_15_, n_n191}, x257x);
	defparam lut_5214.LUT_SIZE = 6;
	defparam lut_5214.mask = 64'h0055ffff00000050;

	lut_sub lut_5217 ({sk[1059], i_9_, i_10_, i_11_, i_15_, n_n213}, n_n122);
	defparam lut_5217.LUT_SIZE = 6;
	defparam lut_5217.mask = 64'h0055ffff10000000;

	lut_sub lut_5219 ({sk[1060], i_14_, i_13_, i_12_, i_15_, n_n184}, x313x);
	defparam lut_5219.LUT_SIZE = 6;
	defparam lut_5219.mask = 64'h0055ffff00000050;

	lut_sub lut_5222 ({sk[1061], n_n42, n_n43, x139x, n_n117, x257x, x313x}, n_n1886);
	defparam lut_5222.LUT_SIZE = 7;
	defparam lut_5222.mask = 128'h00ff00ffffffffff00005fff3f3f7fff;

	lut_sub lut_5228 ({sk[1062], i_14_, i_13_, i_12_, i_15_, n_n149}, x835x);
	defparam lut_5228.LUT_SIZE = 6;
	defparam lut_5228.mask = 64'h0055ffff11410050;

	lut_sub lut_5235 ({sk[1063], i_9_, i_10_, i_11_, i_15_, n_n201}, n_n129);
	defparam lut_5235.LUT_SIZE = 6;
	defparam lut_5235.mask = 64'h0055ffff00000010;

	lut_sub lut_5237 ({sk[1064], i_9_, i_10_, i_11_, i_15_, n_n207}, n_n166);
	defparam lut_5237.LUT_SIZE = 6;
	defparam lut_5237.mask = 64'h0055ffff01000000;

	lut_sub lut_5239 ({sk[1065], i_9_, i_10_, i_11_, i_15_, n_n201}, n_n127);
	defparam lut_5239.LUT_SIZE = 6;
	defparam lut_5239.mask = 64'h0055ffff00100000;

	lut_sub lut_5241 ({sk[1066], i_9_, i_10_, i_11_, n_n41, n_n40, x721x}, n_n1873);
	defparam lut_5241.LUT_SIZE = 7;
	defparam lut_5241.mask = 128'h00ff00ffffffffff1515000015150500;

	lut_sub lut_5251 ({sk[1067], i_9_, i_10_, i_11_, i_15_, n_n213}, n_n88);
	defparam lut_5251.LUT_SIZE = 6;
	defparam lut_5251.mask = 64'h0055ffff00000100;

	lut_sub lut_5253 ({sk[1068], i_9_, i_10_, i_11_, i_15_, n_n207}, n_n173);
	defparam lut_5253.LUT_SIZE = 6;
	defparam lut_5253.mask = 64'h0055ffff00000100;

	lut_sub lut_5255 ({sk[1069], i_9_, i_10_, i_11_, x718x}, n_n73);
	defparam lut_5255.LUT_SIZE = 5;
	defparam lut_5255.mask = 32'h57570004;

	lut_sub lut_5257 ({sk[1070], i_9_, i_10_, i_11_, x723x, x718x}, x1128x);
	defparam lut_5257.LUT_SIZE = 6;
	defparam lut_5257.mask = 64'h0055ffff00700030;

	lut_sub lut_5261 ({sk[1071], n_n38, n_n39, n_n88, n_n173, n_n73, x1128x}, n_n1871);
	defparam lut_5261.LUT_SIZE = 7;
	defparam lut_5261.mask = 128'h00ff00ffffffffff000077775fff7fff;

	lut_sub lut_5267 ({sk[1072], i_7_, i_8_, i_6_, x740x, x714x, x17002x}, x190x);
	defparam lut_5267.LUT_SIZE = 7;
	defparam lut_5267.mask = 128'h00ff00ffffffffff111111111f111111;

	lut_sub lut_5270 ({sk[1073], i_15_, n_n149, n_n40, x714x, x17002x, n_n201}, x2904x);
	defparam lut_5270.LUT_SIZE = 7;
	defparam lut_5270.mask = 128'h00ff00ffffffffff0000000000000155;

	lut_sub lut_5273 ({sk[1074], n_n38, n_n39, n_n82, n_n166, n_n88, n_n173}, x21358x);
	defparam lut_5273.LUT_SIZE = 7;
	defparam lut_5273.mask = 128'h00ff00ffffffffffffff8000f0f08000;

	lut_sub lut_5277 ({sk[1075], n_n38, n_n40, n_n82, n_n129, x2904x, x21358x}, x18857x);
	defparam lut_5277.LUT_SIZE = 7;
	defparam lut_5277.mask = 128'h00ff00ffffffffffbbbbbfbfbbffbfff;

	lut_sub lut_5282 ({sk[1076], i_9_, i_10_, i_11_, i_15_, n_n201}, n_n139);
	defparam lut_5282.LUT_SIZE = 6;
	defparam lut_5282.mask = 64'h0055ffff00010000;

	lut_sub lut_5284 ({sk[1077], i_14_, i_13_, i_12_, i_15_, n_n156, n_n216}, x838x);
	defparam lut_5284.LUT_SIZE = 7;
	defparam lut_5284.mask = 128'h00ff00ffffffffff0303350300003000;

	lut_sub lut_5291 ({sk[1078], i_15_, n_n41, n_n40, n_n199, x838x, n_n201}, x18863x);
	defparam lut_5291.LUT_SIZE = 7;
	defparam lut_5291.mask = 128'h00ff00ffffffffff0000333300053737;

	lut_sub lut_5295 ({sk[1079], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x21357x);
	defparam lut_5295.LUT_SIZE = 7;
	defparam lut_5295.mask = 128'h00ff00fffffffffffcfccffcffffc8ff;

	lut_sub lut_5306 ({sk[1080], n_n40, x714x, x17002x, x835x, x838x, x21357x}, x18864x);
	defparam lut_5306.LUT_SIZE = 7;
	defparam lut_5306.mask = 128'h00ff00ffffffffff0000000fbbbbbbbf;

	lut_sub lut_5310 ({sk[1081], i_14_, i_13_, i_12_, i_15_}, x718x);
	defparam lut_5310.LUT_SIZE = 5;
	defparam lut_5310.mask = 32'h57571000;

	lut_sub lut_5312 ({sk[1082], n_n156, n_n38, n_n36, x143x, n_n102, x718x}, x18867x);
	defparam lut_5312.LUT_SIZE = 7;
	defparam lut_5312.mask = 128'h00ff00ffffffffff003f003f003f557f;

	lut_sub lut_5316 ({sk[1083], i_14_, i_13_, i_12_, i_15_, n_n199}, x74x);
	defparam lut_5316.LUT_SIZE = 6;
	defparam lut_5316.mask = 64'h0055ffff11010000;

	lut_sub lut_5320 ({sk[1084], i_14_, i_13_, i_12_, i_15_, n_n191, n_n199}, x840x);
	defparam lut_5320.LUT_SIZE = 7;
	defparam lut_5320.mask = 128'h00ff00ffffffffff0505500500007700;

	lut_sub lut_5329 ({sk[1085], i_9_, i_10_, i_11_, x729x}, n_n95);
	defparam lut_5329.LUT_SIZE = 5;
	defparam lut_5329.mask = 32'h57570100;

	lut_sub lut_5331 ({sk[1086], i_14_, i_13_, i_12_, i_15_, n_n216}, x364x);
	defparam lut_5331.LUT_SIZE = 6;
	defparam lut_5331.mask = 64'h0055ffff00000050;

	lut_sub lut_5334 ({sk[1087], i_7_, i_8_, i_6_, x735x, x136x}, x2892x);
	defparam lut_5334.LUT_SIZE = 6;
	defparam lut_5334.mask = 64'h0055ffff10000000;

	lut_sub lut_5336 ({sk[1088], n_n34, x143x, x74x, n_n102, n_n95, x364x}, x18872x);
	defparam lut_5336.LUT_SIZE = 7;
	defparam lut_5336.mask = 128'h00ff00ffffffffff000000007fffffff;

	lut_sub lut_5342 ({sk[1089], n_n36, x18867x, x840x, x364x, x2892x, x18872x}, x18874x);
	defparam lut_5342.LUT_SIZE = 7;
	defparam lut_5342.mask = 128'h00ff00ffffffffff7777ffff7fffffff;

	lut_sub lut_5348 ({sk[1090], n_n1873, n_n1871, x18857x, x18863x, x18864x}, x18875x);
	defparam lut_5348.LUT_SIZE = 6;
	defparam lut_5348.mask = 64'h0055ffff7fffffff;

	lut_sub lut_5354 ({sk[1091], i_14_, i_13_, i_12_, i_15_, n_n199}, x68x);
	defparam lut_5354.LUT_SIZE = 6;
	defparam lut_5354.mask = 64'h0055ffff00004044;

	lut_sub lut_5358 ({sk[1092], i_9_, i_10_, i_11_, x720x}, n_n190);
	defparam lut_5358.LUT_SIZE = 5;
	defparam lut_5358.mask = 32'h57570040;

	lut_sub lut_5360 ({sk[1093], i_14_, i_13_, i_12_, i_15_, n_n184}, x842x);
	defparam lut_5360.LUT_SIZE = 6;
	defparam lut_5360.mask = 64'h0055ffff15414440;

	lut_sub lut_5369 ({sk[1094], i_14_, i_13_, i_12_, i_15_, n_n191}, x841x);
	defparam lut_5369.LUT_SIZE = 6;
	defparam lut_5369.mask = 64'h0055ffff15410110;

	lut_sub lut_5377 ({sk[1095], i_14_, i_13_, i_12_, i_15_, n_n184}, x276x);
	defparam lut_5377.LUT_SIZE = 6;
	defparam lut_5377.mask = 64'h0055ffff00000114;

	lut_sub lut_5381 ({sk[1096], i_9_, i_10_, i_11_, n_n123, x721x, x728x}, x2602x);
	defparam lut_5381.LUT_SIZE = 7;
	defparam lut_5381.mask = 128'h00ff00ffffffffff0000070000000700;

	lut_sub lut_5386 ({sk[1097], i_14_, i_13_, i_12_, i_15_, n_n149, n_n125}, x2603x);
	defparam lut_5386.LUT_SIZE = 7;
	defparam lut_5386.mask = 128'h00ff00ffffffffff0000010000100000;

	lut_sub lut_5389 ({sk[1098], n_n113, x842x, x276x, x2602x, x2603x}, x19153x);
	defparam lut_5389.LUT_SIZE = 6;
	defparam lut_5389.mask = 64'h0055ffff77777fff;

	lut_sub lut_5394 ({sk[1099], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x844x);
	defparam lut_5394.LUT_SIZE = 7;
	defparam lut_5394.mask = 128'h00ff00ffffffffff0555000570057570;

	lut_sub lut_5407 ({sk[1100], i_14_, i_13_, i_12_, i_15_, n_n149}, x843x);
	defparam lut_5407.LUT_SIZE = 6;
	defparam lut_5407.mask = 64'h0055ffff15414054;

	lut_sub lut_5417 ({sk[1101], n_n123, n_n148, n_n125, x133x, x60x, x843x}, x19158x);
	defparam lut_5417.LUT_SIZE = 7;
	defparam lut_5417.mask = 128'h00ff00ffffffffff005500ff3f7f3fff;

	lut_sub lut_5422 ({sk[1102], i_9_, i_10_, i_11_, n_n34, x721x, x728x}, x2702x);
	defparam lut_5422.LUT_SIZE = 7;
	defparam lut_5422.mask = 128'h00ff00ffffffffff0700000007000000;

	lut_sub lut_5427 ({sk[1103], i_14_, i_13_, i_12_, i_15_, n_n156}, x19042x);
	defparam lut_5427.LUT_SIZE = 6;
	defparam lut_5427.mask = 64'h0055ffff15000114;

	lut_sub lut_5434 ({sk[1104], i_14_, i_13_, i_12_, i_15_, n_n216}, x49x);
	defparam lut_5434.LUT_SIZE = 6;
	defparam lut_5434.mask = 64'h0055ffff00100400;

	lut_sub lut_5437 ({sk[1105], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x845x);
	defparam lut_5437.LUT_SIZE = 7;
	defparam lut_5437.mask = 128'h00ff00ffffffffff0000005700000057;

	lut_sub lut_5442 ({sk[1106], i_14_, i_13_, i_12_, i_15_, n_n199}, x92x);
	defparam lut_5442.LUT_SIZE = 6;
	defparam lut_5442.mask = 64'h0055ffff00100400;

	lut_sub lut_5445 ({sk[1107], i_9_, i_10_, i_11_, n_n36, x720x}, x2697x);
	defparam lut_5445.LUT_SIZE = 6;
	defparam lut_5445.mask = 64'h0055ffff00100000;

	lut_sub lut_5447 ({sk[1108], i_9_, i_10_, i_11_, x729x, n_n36}, x614x);
	defparam lut_5447.LUT_SIZE = 6;
	defparam lut_5447.mask = 64'h0055ffff00000010;

	lut_sub lut_5449 ({sk[1109], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x848x);
	defparam lut_5449.LUT_SIZE = 7;
	defparam lut_5449.mask = 128'h00ff00ffffffffff0777300770007330;

	lut_sub lut_5465 ({sk[1110], i_14_, i_13_, i_12_, i_15_, n_n149}, x847x);
	defparam lut_5465.LUT_SIZE = 6;
	defparam lut_5465.mask = 64'h0055ffff04400110;

	lut_sub lut_5470 ({sk[1111], i_9_, i_10_, i_11_, n_n34, x721x, x728x}, x2690x);
	defparam lut_5470.LUT_SIZE = 7;
	defparam lut_5470.mask = 128'h00ff00ffffffffff0007000000070000;

	lut_sub lut_5475 ({sk[1112], n_n40, x51x, x98x, x397x, x3523x, x4157x}, x19062x);
	defparam lut_5475.LUT_SIZE = 7;
	defparam lut_5475.mask = 128'h00ff00ffffffffff7f7f7f7f7fffffff;

	lut_sub lut_5481 ({sk[1113], n_n41, n_n40, x51x, n_n102, x98x, x1153x}, x19069x);
	defparam lut_5481.LUT_SIZE = 7;
	defparam lut_5481.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_5486 ({sk[1114], x53x, n_n41, x69x, x4898x, x3518x, x1155x}, x19074x);
	defparam lut_5486.LUT_SIZE = 7;
	defparam lut_5486.mask = 128'h00ff00ffffffffff3f3f7fff3f3fffff;

	lut_sub lut_5492 ({sk[1115], n_n41, n_n40, x1152x, x1151x, x1154x, x1156x}, x21353x);
	defparam lut_5492.LUT_SIZE = 7;
	defparam lut_5492.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_5503 ({sk[1116], x740x, n_n200, x70x, x714x, x17002x, n_n198}, n_n4620);
	defparam lut_5503.LUT_SIZE = 7;
	defparam lut_5503.mask = 128'h00ff00ffffffffff01010101010101ff;

	lut_sub lut_5506 ({sk[1117], i_7_, i_8_, i_6_, x740x, n_n216, x726x}, n_n6384);
	defparam lut_5506.LUT_SIZE = 7;
	defparam lut_5506.mask = 128'h00ff00ffffffffff0000000001000000;

	lut_sub lut_5508 ({sk[1118], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1158x);
	defparam lut_5508.LUT_SIZE = 7;
	defparam lut_5508.mask = 128'h00ff00ffffffffff0707000770057570;

	lut_sub lut_5523 ({sk[1119], i_14_, i_13_, i_12_, i_15_, n_n199}, x1157x);
	defparam lut_5523.LUT_SIZE = 6;
	defparam lut_5523.mask = 64'h0055ffff15414054;

	lut_sub lut_5533 ({sk[1120], x740x, n_n200, x81x, x3543x, n_n1566, x21457x}, x19083x);
	defparam lut_5533.LUT_SIZE = 7;
	defparam lut_5533.mask = 128'h00ff00ffffffffffbfbfbfbfbfbfbfff;

	lut_sub lut_5538 ({sk[1121], x729x, n_n42, n_n43, n_n191, x139x, x1296x}, x19089x);
	defparam lut_5538.LUT_SIZE = 7;
	defparam lut_5538.mask = 128'h00ff00ffffffffff00007777000f777f;

	lut_sub lut_5542 ({sk[1122], n_n42, n_n43, x62x, n_n183, x128x, x1297x}, x19090x);
	defparam lut_5542.LUT_SIZE = 7;
	defparam lut_5542.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_5547 ({sk[1123], x729x, n_n42, x65x, n_n43, n_n191, x1402x}, n_n1294);
	defparam lut_5547.LUT_SIZE = 7;
	defparam lut_5547.mask = 128'h00ff00ffffffffff000f555f000f777f;

	lut_sub lut_5551 ({sk[1124], n_n42, n_n43, n_n136, n_n6348, x391x, x88x}, x19082x);
	defparam lut_5551.LUT_SIZE = 7;
	defparam lut_5551.mask = 128'h00ff00ffffffffff3f3f3fff7f7f7fff;

	lut_sub lut_5556 ({sk[1125], i_14_, i_13_, i_12_, i_15_, n_n156}, x1436x);
	defparam lut_5556.LUT_SIZE = 6;
	defparam lut_5556.mask = 64'h0055ffff15414054;

	lut_sub lut_5566 ({sk[1126], i_9_, i_10_, i_11_, i_15_, n_n201}, n_n137);
	defparam lut_5566.LUT_SIZE = 6;
	defparam lut_5566.mask = 64'h0055ffff00001000;

	lut_sub lut_5568 ({sk[1127], i_14_, i_13_, i_12_, i_15_, n_n170}, x72x);
	defparam lut_5568.LUT_SIZE = 6;
	defparam lut_5568.mask = 64'h0055ffff00100400;

	lut_sub lut_5571 ({sk[1128], i_14_, i_13_, i_12_, i_15_, n_n177}, x378x);
	defparam lut_5571.LUT_SIZE = 6;
	defparam lut_5571.mask = 64'h0055ffff00100400;

	lut_sub lut_5574 ({sk[1129], i_14_, i_13_, i_12_, i_15_, n_n191}, x1501x);
	defparam lut_5574.LUT_SIZE = 6;
	defparam lut_5574.mask = 64'h0055ffff00014154;

	lut_sub lut_5581 ({sk[1130], i_9_, i_10_, i_11_, n_n46, x721x, x728x}, x2643x);
	defparam lut_5581.LUT_SIZE = 7;
	defparam lut_5581.mask = 128'h00ff00ffffffffff0000070000000700;

	lut_sub lut_5586 ({sk[1131], i_9_, i_10_, i_11_, n_n47, x721x, x728x}, x2638x);
	defparam lut_5586.LUT_SIZE = 7;
	defparam lut_5586.mask = 128'h00ff00ffffffffff0007000000070000;

	lut_sub lut_5591 ({sk[1132], i_9_, i_10_, i_11_, n_n47, x721x, x728x}, x2642x);
	defparam lut_5591.LUT_SIZE = 7;
	defparam lut_5591.mask = 128'h00ff00ffffffffff0000070000000700;

	lut_sub lut_5596 ({sk[1133], i_7_, i_8_, i_6_, n_n149, n_n156, x285x}, x19106x);
	defparam lut_5596.LUT_SIZE = 7;
	defparam lut_5596.mask = 128'h00ff00ffffffffff0015000500000000;

	lut_sub lut_5600 ({sk[1134], i_14_, i_13_, i_12_, i_15_, n_n156, n_n199}, x1554x);
	defparam lut_5600.LUT_SIZE = 7;
	defparam lut_5600.mask = 128'h00ff00ffffffffff0330350000500000;

	lut_sub lut_5606 ({sk[1135], i_9_, i_10_, i_11_, n_n47, x721x, x728x}, x2630x);
	defparam lut_5606.LUT_SIZE = 7;
	defparam lut_5606.mask = 128'h00ff00ffffffffff0700000007000000;

	lut_sub lut_5611 ({sk[1136], n_n47, x60x, n_n199, x721x, n_n216, x728x}, x21439x);
	defparam lut_5611.LUT_SIZE = 7;
	defparam lut_5611.mask = 128'h00ff00ffffffffffffffffffeca00000;

	lut_sub lut_5615 ({sk[1137], i_14_, i_13_, i_12_, i_15_, n_n149}, x1888x);
	defparam lut_5615.LUT_SIZE = 6;
	defparam lut_5615.mask = 64'h0055ffff11014044;

	lut_sub lut_5622 ({sk[1138], i_14_, i_13_, i_12_, i_15_, n_n149}, x852x);
	defparam lut_5622.LUT_SIZE = 6;
	defparam lut_5622.mask = 64'h0055ffff15014154;

	lut_sub lut_5632 ({sk[1139], i_14_, i_13_, i_12_, i_15_, n_n199}, n_n140);
	defparam lut_5632.LUT_SIZE = 6;
	defparam lut_5632.mask = 64'h0055ffff00000001;

	lut_sub lut_5634 ({sk[1140], i_14_, i_13_, i_12_, i_15_, n_n156}, x194x);
	defparam lut_5634.LUT_SIZE = 6;
	defparam lut_5634.mask = 64'h0055ffff00050004;

	lut_sub lut_5638 ({sk[1141], i_14_, i_13_, i_12_, i_15_, n_n156}, x853x);
	defparam lut_5638.LUT_SIZE = 6;
	defparam lut_5638.mask = 64'h0055ffff00051114;

	lut_sub lut_5645 ({sk[1142], i_14_, i_13_, i_12_, i_15_, n_n216}, x855x);
	defparam lut_5645.LUT_SIZE = 6;
	defparam lut_5645.mask = 64'h0055ffff00051114;

	lut_sub lut_5652 ({sk[1143], i_9_, i_10_, i_11_, i_15_, n_n207}, x425x);
	defparam lut_5652.LUT_SIZE = 6;
	defparam lut_5652.mask = 64'h0055ffff00050000;

	lut_sub lut_5655 ({sk[1144], n_n36, n_n34, n_n191, x720x, x855x, x425x}, n_n812);
	defparam lut_5655.LUT_SIZE = 7;
	defparam lut_5655.mask = 128'h00ff00ffffffffff00003333555f777f;

	lut_sub lut_5659 ({sk[1145], i_14_, i_13_, i_12_, i_15_, n_n149}, x199x);
	defparam lut_5659.LUT_SIZE = 6;
	defparam lut_5659.mask = 64'h0055ffff00011004;

	lut_sub lut_5663 ({sk[1146], i_14_, i_13_, i_12_, i_15_, n_n149}, x857x);
	defparam lut_5663.LUT_SIZE = 6;
	defparam lut_5663.mask = 64'h0055ffff00051004;

	lut_sub lut_5668 ({sk[1147], i_14_, i_13_, i_12_, i_15_, n_n156}, x290x);
	defparam lut_5668.LUT_SIZE = 6;
	defparam lut_5668.mask = 64'h0055ffff00011004;

	lut_sub lut_5672 ({sk[1148], i_14_, i_13_, i_12_, i_15_, n_n156}, x856x);
	defparam lut_5672.LUT_SIZE = 6;
	defparam lut_5672.mask = 64'h0055ffff00011114;

	lut_sub lut_5678 ({sk[1149], i_7_, i_8_, i_6_, x735x}, x255x);
	defparam lut_5678.LUT_SIZE = 5;
	defparam lut_5678.mask = 32'h57571100;

	lut_sub lut_5681 ({sk[1150], i_9_, i_10_, i_11_, i_15_, n_n207, n_n209}, x19642x);
	defparam lut_5681.LUT_SIZE = 7;
	defparam lut_5681.mask = 128'h00ff00ffffffffff0000000505003005;

	lut_sub lut_5686 ({sk[1151], i_14_, i_13_, i_12_, i_15_, n_n149}, x19643x);
	defparam lut_5686.LUT_SIZE = 6;
	defparam lut_5686.mask = 64'h0055ffff00051114;

	lut_sub lut_5693 ({sk[1152], i_9_, i_10_, i_11_, i_15_, n_n209}, x401x);
	defparam lut_5693.LUT_SIZE = 6;
	defparam lut_5693.mask = 64'h0055ffff00011000;

	lut_sub lut_5696 ({sk[1153], i_8_, n_n16, x735x, n_n184, x719x, x601x}, x19644x);
	defparam lut_5696.LUT_SIZE = 7;
	defparam lut_5696.mask = 128'h00ff00ffffffffff5555555755555557;

	lut_sub lut_5700 ({sk[1154], x735x, n_n126, x118x, n_n72, x401x, x19644x}, x19645x);
	defparam lut_5700.LUT_SIZE = 7;
	defparam lut_5700.mask = 128'h00ff00ffffffffff5555555555557fff;

	lut_sub lut_5705 ({sk[1155], n_n123, n_n125, x857x, x856x, x19642x, x19643x}, x19646x);
	defparam lut_5705.LUT_SIZE = 7;
	defparam lut_5705.mask = 128'h00ff00ffffffffff000000ff7f7f7fff;

	lut_sub lut_5710 ({sk[1156], i_14_, i_13_, i_12_, i_15_}, x723x);
	defparam lut_5710.LUT_SIZE = 5;
	defparam lut_5710.mask = 32'h57570008;

	lut_sub lut_5712 ({sk[1157], i_9_, i_10_, i_11_, i_15_, n_n207}, n_n103);
	defparam lut_5712.LUT_SIZE = 6;
	defparam lut_5712.mask = 64'h0055ffff00000004;

	lut_sub lut_5714 ({sk[1158], i_9_, i_10_, i_11_, i_15_, n_n201}, n_n115);
	defparam lut_5714.LUT_SIZE = 6;
	defparam lut_5714.mask = 64'h0055ffff10000000;

	lut_sub lut_5716 ({sk[1159], i_9_, i_10_, i_11_, x728x}, n_n54);
	defparam lut_5716.LUT_SIZE = 5;
	defparam lut_5716.mask = 32'h57570004;

	lut_sub lut_5718 ({sk[1160], i_14_, i_13_, i_12_, i_15_}, x727x);
	defparam lut_5718.LUT_SIZE = 5;
	defparam lut_5718.mask = 32'h57570002;

	lut_sub lut_5720 ({sk[1161], i_9_, i_10_, i_11_, x726x}, n_n178);
	defparam lut_5720.LUT_SIZE = 5;
	defparam lut_5720.mask = 32'h57574000;

	lut_sub lut_5722 ({sk[1162], i_9_, i_10_, i_11_, x720x}, n_n183);
	defparam lut_5722.LUT_SIZE = 5;
	defparam lut_5722.mask = 32'h57574000;

	lut_sub lut_5724 ({sk[1163], i_9_, i_10_, i_11_, x728x}, n_n62);
	defparam lut_5724.LUT_SIZE = 5;
	defparam lut_5724.mask = 32'h57570100;

	lut_sub lut_5726 ({sk[1164], i_9_, i_10_, i_11_, i_15_, n_n207}, n_n84);
	defparam lut_5726.LUT_SIZE = 6;
	defparam lut_5726.mask = 64'h0055ffff00000400;

	lut_sub lut_5728 ({sk[1165], i_9_, i_10_, i_11_, i_15_, n_n211}, n_n210);
	defparam lut_5728.LUT_SIZE = 6;
	defparam lut_5728.mask = 64'h0055ffff00000001;

	lut_sub lut_5730 ({sk[1166], i_9_, i_10_, i_11_, x720x}, n_n176);
	defparam lut_5730.LUT_SIZE = 5;
	defparam lut_5730.mask = 32'h57570010;

	lut_sub lut_5732 ({sk[1167], i_9_, i_10_, i_11_, x728x}, n_n60);
	defparam lut_5732.LUT_SIZE = 5;
	defparam lut_5732.mask = 32'h57570040;

	lut_sub lut_5734 ({sk[1168], i_14_, i_13_, i_12_, i_15_, n_n199}, x81x);
	defparam lut_5734.LUT_SIZE = 6;
	defparam lut_5734.mask = 64'h0055ffff00000110;

	lut_sub lut_5737 ({sk[1169], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x861x);
	defparam lut_5737.LUT_SIZE = 7;
	defparam lut_5737.mask = 128'h00ff00ffffffffff0555505557037370;

	lut_sub lut_5753 ({sk[1170], i_14_, i_13_, i_12_, i_15_, n_n184}, x860x);
	defparam lut_5753.LUT_SIZE = 6;
	defparam lut_5753.mask = 64'h0055ffff15455154;

	lut_sub lut_5766 ({sk[1171], i_7_, i_8_, i_6_, x734x, x81x}, x3011x);
	defparam lut_5766.LUT_SIZE = 6;
	defparam lut_5766.mask = 64'h0055ffff10000000;

	lut_sub lut_5768 ({sk[1172], i_9_, i_10_, i_11_, x729x, n_n31}, x3012x);
	defparam lut_5768.LUT_SIZE = 6;
	defparam lut_5768.mask = 64'h0055ffff00000001;

	lut_sub lut_5770 ({sk[1173], i_14_, i_13_, i_12_, i_15_, n_n216}, x863x);
	defparam lut_5770.LUT_SIZE = 6;
	defparam lut_5770.mask = 64'h0055ffff15055154;

	lut_sub lut_5782 ({sk[1174], i_14_, i_13_, i_12_, i_15_, n_n199}, x862x);
	defparam lut_5782.LUT_SIZE = 6;
	defparam lut_5782.mask = 64'h0055ffff15055044;

	lut_sub lut_5792 ({sk[1175], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x864x);
	defparam lut_5792.LUT_SIZE = 7;
	defparam lut_5792.mask = 128'h00ff00ffffffffff0000300005055550;

	lut_sub lut_5799 ({sk[1176], i_14_, i_13_, i_12_, i_15_, n_n212, n_n199}, x4792x);
	defparam lut_5799.LUT_SIZE = 7;
	defparam lut_5799.mask = 128'h00ff00ffffffffff0000000000000001;

	lut_sub lut_5801 ({sk[1177], i_14_, i_13_, i_12_, i_15_, n_n199}, x247x);
	defparam lut_5801.LUT_SIZE = 6;
	defparam lut_5801.mask = 64'h0055ffff40100400;

	lut_sub lut_5805 ({sk[1178], n_n197, n_n212, x719x, n_n63, n_n199, x728x}, x704x);
	defparam lut_5805.LUT_SIZE = 7;
	defparam lut_5805.mask = 128'h00ff00ffffffffff00000f0f11331f3f;

	lut_sub lut_5809 ({sk[1179], i_14_, i_13_, i_12_, i_15_, n_n199}, x153x);
	defparam lut_5809.LUT_SIZE = 6;
	defparam lut_5809.mask = 64'h0055ffff40100000;

	lut_sub lut_5812 ({sk[1180], n_n197, n_n212, n_n140, x247x, x704x, x153x}, n_n4231);
	defparam lut_5812.LUT_SIZE = 7;
	defparam lut_5812.mask = 128'h00ff00ffffffffff33333fff77777fff;

	lut_sub lut_5817 ({sk[1181], i_14_, i_13_, i_12_, i_15_, n_n199}, x218x);
	defparam lut_5817.LUT_SIZE = 6;
	defparam lut_5817.mask = 64'h0055ffff00100401;

	lut_sub lut_5821 ({sk[1182], i_14_, i_13_, i_12_, i_15_, n_n216}, x56x);
	defparam lut_5821.LUT_SIZE = 6;
	defparam lut_5821.mask = 64'h0055ffff11000000;

	lut_sub lut_5824 ({sk[1183], i_14_, i_13_, i_12_, i_15_, n_n156}, x248x);
	defparam lut_5824.LUT_SIZE = 6;
	defparam lut_5824.mask = 64'h0055ffff01004040;

	lut_sub lut_5828 ({sk[1184], i_14_, i_13_, i_12_, i_15_, n_n199}, x866x);
	defparam lut_5828.LUT_SIZE = 6;
	defparam lut_5828.mask = 64'h0055ffff15454044;

	lut_sub lut_5838 ({sk[1185], i_7_, i_8_, i_6_, x734x, x84x}, x4329x);
	defparam lut_5838.LUT_SIZE = 6;
	defparam lut_5838.mask = 64'h0055ffff01000000;

	lut_sub lut_5840 ({sk[1186], i_14_, i_13_, i_12_, i_15_, n_n216}, x1572x);
	defparam lut_5840.LUT_SIZE = 6;
	defparam lut_5840.mask = 64'h0055ffff11015154;

	lut_sub lut_5850 ({sk[1187], i_14_, i_13_, i_12_, i_15_, n_n199}, x1224x);
	defparam lut_5850.LUT_SIZE = 6;
	defparam lut_5850.mask = 64'h0055ffff15455154;

	lut_sub lut_5863 ({sk[1188], i_14_, i_13_, i_12_, i_15_, n_n216}, x47x);
	defparam lut_5863.LUT_SIZE = 6;
	defparam lut_5863.mask = 64'h0055ffff00001110;

	lut_sub lut_5867 ({sk[1189], i_14_, i_13_, i_12_, i_15_, n_n216}, x1855x);
	defparam lut_5867.LUT_SIZE = 6;
	defparam lut_5867.mask = 64'h0055ffff11014044;

	lut_sub lut_5874 ({sk[1190], i_14_, i_13_, i_12_, i_15_, n_n199}, x1854x);
	defparam lut_5874.LUT_SIZE = 6;
	defparam lut_5874.mask = 64'h0055ffff11014044;

	lut_sub lut_5881 ({sk[1191], i_14_, i_13_, i_12_, i_15_, n_n156}, x1878x);
	defparam lut_5881.LUT_SIZE = 6;
	defparam lut_5881.mask = 64'h0055ffff00005154;

	lut_sub lut_5888 ({sk[1192], n_n197, n_n212, x55x, x133x, x127x, x176x}, x17519x);
	defparam lut_5888.LUT_SIZE = 7;
	defparam lut_5888.mask = 128'h00ff00ffffffffff00007f7f00ff7fff;

	lut_sub lut_5893 ({sk[1193], x181x, x735x, n_n200, n_n212, x55x, x1878x}, x17520x);
	defparam lut_5893.LUT_SIZE = 7;
	defparam lut_5893.mask = 128'h00ff00ffffffffff07070707070707ff;

	lut_sub lut_5897 ({sk[1194], n_n197, n_n212, x133x, x127x, x158x, x123x}, x17521x);
	defparam lut_5897.LUT_SIZE = 7;
	defparam lut_5897.mask = 128'h00ff00ffffffffff000055553fff7fff;

	lut_sub lut_5902 ({sk[1195], i_7_, i_8_, i_6_, x740x, x172x}, n_n5061);
	defparam lut_5902.LUT_SIZE = 6;
	defparam lut_5902.mask = 64'h0055ffff00001000;

	lut_sub lut_5904 ({sk[1196], i_7_, i_8_, i_6_, x735x, x123x}, n_n4266);
	defparam lut_5904.LUT_SIZE = 6;
	defparam lut_5904.mask = 64'h0055ffff10000000;

	lut_sub lut_5906 ({sk[1197], i_14_, i_13_, i_12_, i_15_, n_n156}, x156x);
	defparam lut_5906.LUT_SIZE = 6;
	defparam lut_5906.mask = 64'h0055ffff00004044;

	lut_sub lut_5910 ({sk[1198], i_14_, i_13_, i_12_, i_15_, n_n177}, x104x);
	defparam lut_5910.LUT_SIZE = 6;
	defparam lut_5910.mask = 64'h0055ffff00000110;

	lut_sub lut_5913 ({sk[1199], i_7_, i_8_, i_6_, x729x, x740x, n_n191}, x3352x);
	defparam lut_5913.LUT_SIZE = 7;
	defparam lut_5913.mask = 128'h00ff00ffffffffff0000000000010000;

	lut_sub lut_5915 ({sk[1200], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x869x);
	defparam lut_5915.LUT_SIZE = 7;
	defparam lut_5915.mask = 128'h00ff00ffffffffff0337303775005050;

	lut_sub lut_5929 ({sk[1201], i_14_, i_13_, i_12_, i_15_, n_n191}, x868x);
	defparam lut_5929.LUT_SIZE = 6;
	defparam lut_5929.mask = 64'h0055ffff15055154;

	lut_sub lut_5941 ({sk[1202], n_n89, n_n46, n_n47, x104x, x869x, x868x}, n_n3194);
	defparam lut_5941.LUT_SIZE = 7;
	defparam lut_5941.mask = 128'h00ff00ffffffffff003f557f003fffff;

	lut_sub lut_5946 ({sk[1203], i_7_, i_6_, n_n111, n_n7252, n_n19, x746x}, x18701x);
	defparam lut_5946.LUT_SIZE = 7;
	defparam lut_5946.mask = 128'h00ff00ffffffffff0f0f0f3f0f0f5f7f;

	lut_sub lut_5951 ({sk[1204], i_7_, i_6_, x732x, n_n7254, x731x, x746x}, x18702x);
	defparam lut_5951.LUT_SIZE = 7;
	defparam lut_5951.mask = 128'h00ff00ffffffffff0f0f7fff0f0f3f3f;

	lut_sub lut_5957 ({sk[1205], i_14_, i_13_, i_12_, i_15_, n_n216}, x154x);
	defparam lut_5957.LUT_SIZE = 6;
	defparam lut_5957.mask = 64'h0055ffff00004044;

	lut_sub lut_5961 ({sk[1206], x181x, n_n46, n_n47, x143x, x48x, x154x}, x18170x);
	defparam lut_5961.LUT_SIZE = 7;
	defparam lut_5961.mask = 128'h00ff00ffffffffff00335f7f0033ffff;

	lut_sub lut_5966 ({sk[1207], i_14_, i_13_, i_12_, i_15_, n_n199}, x1897x);
	defparam lut_5966.LUT_SIZE = 6;
	defparam lut_5966.mask = 64'h0055ffff11014044;

	lut_sub lut_5973 ({sk[1208], n_n46, x168x, n_n47, x63x, x47x, x1897x}, x18171x);
	defparam lut_5973.LUT_SIZE = 7;
	defparam lut_5973.mask = 128'h00ff00ffffffffff005f00ff337f33ff;

	lut_sub lut_5978 ({sk[1209], i_7_, i_8_, i_6_, x740x, x151x}, n_n5121);
	defparam lut_5978.LUT_SIZE = 6;
	defparam lut_5978.mask = 64'h0055ffff00000100;

	lut_sub lut_5980 ({sk[1210], x181x, n_n46, x168x, n_n47, x74x, x68x}, x18175x);
	defparam lut_5980.LUT_SIZE = 7;
	defparam lut_5980.mask = 128'h00ff00ffffffffff000077ff0f0f7fff;

	lut_sub lut_5985 ({sk[1211], n_n46, n_n47, x143x, x151x, x47x, x154x}, x18176x);
	defparam lut_5985.LUT_SIZE = 7;
	defparam lut_5985.mask = 128'h00ff00ffffffffff00007fff0f0f7fff;

	lut_sub lut_5991 ({sk[1212], i_14_, i_13_, i_12_, i_15_, n_n184}, x875x);
	defparam lut_5991.LUT_SIZE = 6;
	defparam lut_5991.mask = 64'h0055ffff15455154;

	lut_sub lut_6004 ({sk[1213], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x874x);
	defparam lut_6004.LUT_SIZE = 7;
	defparam lut_6004.mask = 128'h00ff00ffffffffff0707000730003030;

	lut_sub lut_6014 ({sk[1214], n_n46, x124x, n_n47, x129x, x875x, x874x}, x18180x);
	defparam lut_6014.LUT_SIZE = 7;
	defparam lut_6014.mask = 128'h00ff00ffffffffff005f00ff337f33ff;

	lut_sub lut_6019 ({sk[1215], i_7_, i_6_, n_n89, x741x, x744x, n_n10}, x18494x);
	defparam lut_6019.LUT_SIZE = 7;
	defparam lut_6019.mask = 128'h00ff00ffffffffff3f7f337733773377;

	lut_sub lut_6026 ({sk[1216], x729x, n_n149, x717x, n_n3, n_n191, x730x}, x3244x);
	defparam lut_6026.LUT_SIZE = 7;
	defparam lut_6026.mask = 128'h00ff00ffffffffff0103050703030f0f;

	lut_sub lut_6032 ({sk[1217], n_n9, n_n17, x288x, x77x, n_n6, x454x}, x18497x);
	defparam lut_6032.LUT_SIZE = 7;
	defparam lut_6032.mask = 128'h00ff00ffffffffff575757ff5f5f5fff;

	lut_sub lut_6037 ({sk[1218], i_7_, i_5_, i_6_, i_3_, i_4_, n_n19}, x423x);
	defparam lut_6037.LUT_SIZE = 7;
	defparam lut_6037.mask = 128'h00ff00ffffffffff1010101010101000;

	lut_sub lut_6045 ({sk[1219], i_14_, i_13_, i_12_, i_15_, n_n191}, x307x);
	defparam lut_6045.LUT_SIZE = 6;
	defparam lut_6045.mask = 64'h0055ffff10044000;

	lut_sub lut_6049 ({sk[1220], i_14_, i_13_, i_12_, i_15_, n_n191}, x885x);
	defparam lut_6049.LUT_SIZE = 6;
	defparam lut_6049.mask = 64'h0055ffff10045000;

	lut_sub lut_6054 ({sk[1221], i_14_, i_13_, i_12_, i_15_, n_n184}, x202x);
	defparam lut_6054.LUT_SIZE = 6;
	defparam lut_6054.mask = 64'h0055ffff10044000;

	lut_sub lut_6058 ({sk[1222], i_9_, i_10_, i_11_, i_15_, x95x, n_n211}, x308x);
	defparam lut_6058.LUT_SIZE = 7;
	defparam lut_6058.mask = 128'h00ff00ffffffffff3333333333333733;

	lut_sub lut_6061 ({sk[1223], i_14_, i_13_, i_12_, i_15_, n_n149}, x299x);
	defparam lut_6061.LUT_SIZE = 6;
	defparam lut_6061.mask = 64'h0055ffff10005000;

	lut_sub lut_6065 ({sk[1224], i_9_, i_10_, i_11_, x725x}, x417x);
	defparam lut_6065.LUT_SIZE = 5;
	defparam lut_6065.mask = 32'h57574010;

	lut_sub lut_6068 ({sk[1225], i_9_, i_10_, i_11_, x725x, n_n197, n_n212}, x21400x);
	defparam lut_6068.LUT_SIZE = 7;
	defparam lut_6068.mask = 128'h00ff00fffffffffffcf8fffffcfcfffc;

	lut_sub lut_6076 ({sk[1226], x735x, n_n200, n_n212, n_n63, x176x, n_n61}, x21422x);
	defparam lut_6076.LUT_SIZE = 7;
	defparam lut_6076.mask = 128'h00ff00ffffffffff005f005f005f777f;

	lut_sub lut_6088 ({sk[1227], i_7_, i_8_, i_6_, x740x, x714x, x17051x}, x189x);
	defparam lut_6088.LUT_SIZE = 7;
	defparam lut_6088.mask = 128'h00ff00ffffffffff11111111111f1111;

	lut_sub lut_6091 ({sk[1228], i_14_, i_13_, i_12_, i_15_, n_n149, n_n191}, x890x);
	defparam lut_6091.LUT_SIZE = 7;
	defparam lut_6091.mask = 128'h00ff00ffffffffff5330303033000000;

	lut_sub lut_6099 ({sk[1229], i_9_, i_10_, i_11_, i_15_, n_n204, x308x}, x17195x);
	defparam lut_6099.LUT_SIZE = 7;
	defparam lut_6099.mask = 128'h00ff00ffffffffff7555555555555575;

	lut_sub lut_6103 ({sk[1230], i_14_, i_13_, i_12_, i_15_, n_n156}, x116x);
	defparam lut_6103.LUT_SIZE = 6;
	defparam lut_6103.mask = 64'h0055ffff14040000;

	lut_sub lut_6107 ({sk[1231], i_14_, i_13_, i_12_, i_15_, n_n156}, x892x);
	defparam lut_6107.LUT_SIZE = 6;
	defparam lut_6107.mask = 64'h0055ffff14045000;

	lut_sub lut_6113 ({sk[1232], i_14_, i_13_, i_12_, i_15_, n_n149}, x369x);
	defparam lut_6113.LUT_SIZE = 6;
	defparam lut_6113.mask = 64'h0055ffff00005000;

	lut_sub lut_6116 ({sk[1233], i_9_, i_10_, i_11_, x729x, x369x}, x891x);
	defparam lut_6116.LUT_SIZE = 6;
	defparam lut_6116.mask = 64'h0055ffff55555755;

	lut_sub lut_6119 ({sk[1234], i_14_, i_13_, i_12_, i_15_, n_n191}, x93x);
	defparam lut_6119.LUT_SIZE = 6;
	defparam lut_6119.mask = 64'h0055ffff14040000;

	lut_sub lut_6123 ({sk[1235], i_14_, i_13_, i_12_, i_15_, n_n184}, x967x);
	defparam lut_6123.LUT_SIZE = 6;
	defparam lut_6123.mask = 64'h0055ffff14045000;

	lut_sub lut_6129 ({sk[1236], i_9_, i_10_, i_11_, x725x, x714x, x17051x}, x609x);
	defparam lut_6129.LUT_SIZE = 7;
	defparam lut_6129.mask = 128'h00ff00ffffffffff0000000000000100;

	lut_sub lut_6131 ({sk[1237], i_7_, i_8_, i_6_, x740x, x725x, n_n177}, x611x);
	defparam lut_6131.LUT_SIZE = 7;
	defparam lut_6131.mask = 128'h00ff00ffffffffff0000000000010000;

	lut_sub lut_6133 ({sk[1238], i_14_, i_13_, i_12_, i_15_, n_n184}, x94x);
	defparam lut_6133.LUT_SIZE = 6;
	defparam lut_6133.mask = 64'h0055ffff14040000;

	lut_sub lut_6137 ({sk[1239], i_14_, i_13_, i_12_, i_15_, n_n184}, x895x);
	defparam lut_6137.LUT_SIZE = 6;
	defparam lut_6137.mask = 64'h0055ffff14045000;

	lut_sub lut_6143 ({sk[1240], i_14_, i_13_, i_12_, i_15_, n_n191}, x301x);
	defparam lut_6143.LUT_SIZE = 6;
	defparam lut_6143.mask = 64'h0055ffff00005000;

	lut_sub lut_6146 ({sk[1241], i_14_, i_13_, i_12_, i_15_, n_n177}, x131x);
	defparam lut_6146.LUT_SIZE = 6;
	defparam lut_6146.mask = 64'h0055ffff04440000;

	lut_sub lut_6150 ({sk[1242], i_14_, i_13_, i_12_, i_15_, n_n170}, x201x);
	defparam lut_6150.LUT_SIZE = 6;
	defparam lut_6150.mask = 64'h0055ffff10005000;

	lut_sub lut_6154 ({sk[1243], i_14_, i_13_, i_12_, i_15_, n_n156, n_n177}, x17208x);
	defparam lut_6154.LUT_SIZE = 7;
	defparam lut_6154.mask = 128'h00ff00ffffffffff0350505033000000;

	lut_sub lut_6161 ({sk[1244], i_9_, i_10_, i_11_, x729x, x725x, x726x}, x969x);
	defparam lut_6161.LUT_SIZE = 7;
	defparam lut_6161.mask = 128'h00ff00ffffffffff003333007f000000;

	lut_sub lut_6167 ({sk[1245], i_9_, i_10_, i_11_, x725x, n_n36, n_n34}, x21398x);
	defparam lut_6167.LUT_SIZE = 7;
	defparam lut_6167.mask = 128'h00ff00fffffffffffffff8fffffaf8ff;

	lut_sub lut_6176 ({sk[1246], i_14_, i_13_, i_12_, i_15_, n_n149, n_n170}, x1054x);
	defparam lut_6176.LUT_SIZE = 7;
	defparam lut_6176.mask = 128'h00ff00ffffffffff0350503033000000;

	lut_sub lut_6183 ({sk[1247], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x17225x);
	defparam lut_6183.LUT_SIZE = 7;
	defparam lut_6183.mask = 128'h00ff00ffffffffff0500005057000000;

	lut_sub lut_6189 ({sk[1248], i_9_, i_10_, i_11_, i_15_, n_n32, n_n211}, x4656x);
	defparam lut_6189.LUT_SIZE = 7;
	defparam lut_6189.mask = 128'h00ff00ffffffffff0100000000000000;

	lut_sub lut_6191 ({sk[1249], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x900x);
	defparam lut_6191.LUT_SIZE = 7;
	defparam lut_6191.mask = 128'h00ff00ffffffffff0730303077000000;

	lut_sub lut_6201 ({sk[1250], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x17237x);
	defparam lut_6201.LUT_SIZE = 7;
	defparam lut_6201.mask = 128'h00ff00ffffffffff0530303055000000;

	lut_sub lut_6208 ({sk[1251], i_9_, i_10_, i_11_, x725x, x176x}, x17235x);
	defparam lut_6208.LUT_SIZE = 6;
	defparam lut_6208.mask = 64'h0055ffff55557555;

	lut_sub lut_6211 ({sk[1252], i_7_, i_8_, i_6_, n_n31, x734x, n_n61}, x4640x);
	defparam lut_6211.LUT_SIZE = 7;
	defparam lut_6211.mask = 128'h00ff00ffffffffff1505050505050505;

	lut_sub lut_6214 ({sk[1253], i_14_, i_13_, i_12_, i_15_, n_n156, n_n177}, x17244x);
	defparam lut_6214.LUT_SIZE = 7;
	defparam lut_6214.mask = 128'h00ff00ffffffffff0350505033000000;

	lut_sub lut_6221 ({sk[1254], i_14_, i_13_, i_12_, i_15_, n_n149}, x376x);
	defparam lut_6221.LUT_SIZE = 6;
	defparam lut_6221.mask = 64'h0055ffff00000050;

	lut_sub lut_6224 ({sk[1255], n_n65, n_n71, n_n123, n_n125, x133x, x376x}, n_n1918);
	defparam lut_6224.LUT_SIZE = 7;
	defparam lut_6224.mask = 128'h00ff00ffffffffff05770f7f05ff0fff;

	lut_sub lut_6230 ({sk[1256], i_14_, i_13_, i_12_, i_15_, n_n184}, x310x);
	defparam lut_6230.LUT_SIZE = 6;
	defparam lut_6230.mask = 64'h0055ffff01010040;

	lut_sub lut_6234 ({sk[1257], i_14_, i_13_, i_12_, i_15_, n_n184}, x906x);
	defparam lut_6234.LUT_SIZE = 6;
	defparam lut_6234.mask = 64'h0055ffff11410050;

	lut_sub lut_6241 ({sk[1258], i_14_, i_13_, i_12_, i_15_, n_n191}, x293x);
	defparam lut_6241.LUT_SIZE = 6;
	defparam lut_6241.mask = 64'h0055ffff10400000;

	lut_sub lut_6244 ({sk[1259], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x905x);
	defparam lut_6244.LUT_SIZE = 7;
	defparam lut_6244.mask = 128'h00ff00ffffffffff0500500000000300;

	lut_sub lut_6248 ({sk[1260], i_9_, i_10_, i_11_, n_n36, n_n34, x721x}, n_n1859);
	defparam lut_6248.LUT_SIZE = 7;
	defparam lut_6248.mask = 128'h00ff00ffffffffff1515000515050011;

	lut_sub lut_6258 ({sk[1261], i_9_, i_10_, i_11_, i_15_, x175x, n_n201}, x908x);
	defparam lut_6258.LUT_SIZE = 7;
	defparam lut_6258.mask = 128'h00ff00ffffffffff3333733733337333;

	lut_sub lut_6263 ({sk[1262], i_8_, n_n157, x735x, x133x, x123x, x908x}, x18883x);
	defparam lut_6263.LUT_SIZE = 7;
	defparam lut_6263.mask = 128'h00ff00ffffffffff0000007f00000000;

	lut_sub lut_6267 ({sk[1263], i_7_, i_8_, i_6_, x735x, x52x}, n_n3961);
	defparam lut_6267.LUT_SIZE = 6;
	defparam lut_6267.mask = 64'h0055ffff10000000;

	lut_sub lut_6269 ({sk[1264], x729x, n_n36, n_n34, n_n184, x139x, x257x}, x18886x);
	defparam lut_6269.LUT_SIZE = 7;
	defparam lut_6269.mask = 128'h00ff00ffffffffff00553377005f337f;

	lut_sub lut_6273 ({sk[1265], i_14_, i_13_, i_12_, i_15_, n_n177, n_n191}, x910x);
	defparam lut_6273.LUT_SIZE = 7;
	defparam lut_6273.mask = 128'h00ff00ffffffffff0303500300003300;

	lut_sub lut_6280 ({sk[1266], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x909x);
	defparam lut_6280.LUT_SIZE = 7;
	defparam lut_6280.mask = 128'h00ff00ffffffffff0303500300003300;

	lut_sub lut_6287 ({sk[1267], i_8_, n_n157, n_n36, x735x, x910x, x909x}, x18890x);
	defparam lut_6287.LUT_SIZE = 7;
	defparam lut_6287.mask = 128'h00ff00ffffffffff0033053700330033;

	lut_sub lut_6290 ({sk[1268], i_7_, i_8_, i_6_, x735x, x146x}, n_n4568);
	defparam lut_6290.LUT_SIZE = 6;
	defparam lut_6290.mask = 64'h0055ffff10000000;

	lut_sub lut_6292 ({sk[1269], x729x, n_n36, n_n34, n_n177, x123x, x376x}, x18893x);
	defparam lut_6292.LUT_SIZE = 7;
	defparam lut_6292.mask = 128'h00ff00ffffffffff00553377005f337f;

	lut_sub lut_6296 ({sk[1270], i_14_, i_13_, i_12_, i_15_, n_n170}, x183x);
	defparam lut_6296.LUT_SIZE = 6;
	defparam lut_6296.mask = 64'h0055ffff00000050;

	lut_sub lut_6299 ({sk[1271], i_14_, i_13_, i_12_, i_15_, n_n177}, x383x);
	defparam lut_6299.LUT_SIZE = 6;
	defparam lut_6299.mask = 64'h0055ffff00000050;

	lut_sub lut_6302 ({sk[1272], n_n36, n_n34, n_n83, n_n77, x183x, x383x}, x18897x);
	defparam lut_6302.LUT_SIZE = 7;
	defparam lut_6302.mask = 128'h00ff00ffffffffff000077773fff7fff;

	lut_sub lut_6308 ({sk[1273], x729x, n_n36, n_n34, x146x, n_n170, x147x}, x18898x);
	defparam lut_6308.LUT_SIZE = 7;
	defparam lut_6308.mask = 128'h00ff00ffffffffff005f555f007f557f;

	lut_sub lut_6313 ({sk[1274], n_n71, n_n36, x175x, x18893x, x18897x, x18898x}, x18900x);
	defparam lut_6313.LUT_SIZE = 7;
	defparam lut_6313.mask = 128'h00ff00ffffffffff7f7f7fff7f7fffff;

	lut_sub lut_6319 ({sk[1275], x729x, n_n149, n_n36, n_n141, x133x, x376x}, x18882x);
	defparam lut_6319.LUT_SIZE = 7;
	defparam lut_6319.mask = 128'h00ff00ffffffffff007f007f007f00ff;

	lut_sub lut_6324 ({sk[1276], n_n36, n_n34, x52x, n_n117, x313x, x18886x}, x21356x);
	defparam lut_6324.LUT_SIZE = 7;
	defparam lut_6324.mask = 128'h00ff00ffffffffffaaaaaa0080008000;

	lut_sub lut_6328 ({sk[1277], n_n1859, x18883x, x18890x, x18882x, x21356x}, x18901x);
	defparam lut_6328.LUT_SIZE = 6;
	defparam lut_6328.mask = 64'h0055ffffbfffffff;

	lut_sub lut_6334 ({sk[1278], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x914x);
	defparam lut_6334.LUT_SIZE = 7;
	defparam lut_6334.mask = 128'h00ff00ffffffffff0777500730033330;

	lut_sub lut_6349 ({sk[1279], i_14_, i_13_, i_12_, i_15_, n_n184}, x913x);
	defparam lut_6349.LUT_SIZE = 6;
	defparam lut_6349.mask = 64'h0055ffff15414154;

	lut_sub lut_6360 ({sk[1280], i_7_, i_8_, i_6_, x735x, n_n177, x720x}, x4757x);
	defparam lut_6360.LUT_SIZE = 7;
	defparam lut_6360.mask = 128'h00ff00ffffffffff0001000000000000;

	lut_sub lut_6362 ({sk[1281], i_14_, i_13_, i_12_, i_15_, n_n149, n_n177}, x916x);
	defparam lut_6362.LUT_SIZE = 7;
	defparam lut_6362.mask = 128'h00ff00ffffffffff0555500550035750;

	lut_sub lut_6374 ({sk[1282], i_14_, i_13_, i_12_, i_15_, n_n156}, x227x);
	defparam lut_6374.LUT_SIZE = 6;
	defparam lut_6374.mask = 64'h0055ffff00000114;

	lut_sub lut_6378 ({sk[1283], i_14_, i_13_, i_12_, i_15_, n_n156}, x232x);
	defparam lut_6378.LUT_SIZE = 6;
	defparam lut_6378.mask = 64'h0055ffff15000000;

	lut_sub lut_6382 ({sk[1284], i_14_, i_13_, i_12_, i_15_, n_n156, n_n125}, x19163x);
	defparam lut_6382.LUT_SIZE = 7;
	defparam lut_6382.mask = 128'h00ff00ffffffffff0111100110011110;

	lut_sub lut_6393 ({sk[1285], n_n123, n_n125, x69x, x147x, n_n176, x916x}, x19164x);
	defparam lut_6393.LUT_SIZE = 7;
	defparam lut_6393.mask = 128'h00ff00ffffffffff00000fff77777fff;

	lut_sub lut_6398 ({sk[1286], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x918x);
	defparam lut_6398.LUT_SIZE = 7;
	defparam lut_6398.mask = 128'h00ff00ffffffffff0333300370057770;

	lut_sub lut_6413 ({sk[1287], i_14_, i_13_, i_12_, i_15_, n_n184}, x917x);
	defparam lut_6413.LUT_SIZE = 6;
	defparam lut_6413.mask = 64'h0055ffff15014154;

	lut_sub lut_6423 ({sk[1288], n_n123, n_n125, x52x, n_n117, x918x, x917x}, n_n1209);
	defparam lut_6423.LUT_SIZE = 7;
	defparam lut_6423.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_6428 ({sk[1289], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x920x);
	defparam lut_6428.LUT_SIZE = 7;
	defparam lut_6428.mask = 128'h00ff00ffffffffff0333300370057770;

	lut_sub lut_6443 ({sk[1290], i_14_, i_13_, i_12_, i_15_, n_n170}, x919x);
	defparam lut_6443.LUT_SIZE = 6;
	defparam lut_6443.mask = 64'h0055ffff15014154;

	lut_sub lut_6453 ({sk[1291], n_n123, n_n125, x51x, n_n176, n_n77, x919x}, x19176x);
	defparam lut_6453.LUT_SIZE = 7;
	defparam lut_6453.mask = 128'h00ff00ffffffffff00000f0f77ff7fff;

	lut_sub lut_6458 ({sk[1292], i_9_, i_10_, i_11_, i_15_, n_n32, n_n201}, x2918x);
	defparam lut_6458.LUT_SIZE = 7;
	defparam lut_6458.mask = 128'h00ff00ffffffffff0100000000000000;

	lut_sub lut_6460 ({sk[1293], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1288x);
	defparam lut_6460.LUT_SIZE = 7;
	defparam lut_6460.mask = 128'h00ff00ffffffffff0057030075000000;

	lut_sub lut_6466 ({sk[1294], i_9_, i_10_, i_11_, n_n32, x728x}, x2619x);
	defparam lut_6466.LUT_SIZE = 6;
	defparam lut_6466.mask = 64'h0055ffff10000000;

	lut_sub lut_6468 ({sk[1295], i_14_, i_13_, i_12_, i_15_, n_n216}, x251x);
	defparam lut_6468.LUT_SIZE = 6;
	defparam lut_6468.mask = 64'h0055ffff15000000;

	lut_sub lut_6472 ({sk[1296], i_14_, i_13_, i_12_, i_15_, n_n149}, x1848x);
	defparam lut_6472.LUT_SIZE = 6;
	defparam lut_6472.mask = 64'h0055ffff11014044;

	lut_sub lut_6479 ({sk[1297], i_14_, i_13_, i_12_, i_15_, n_n184}, x924x);
	defparam lut_6479.LUT_SIZE = 6;
	defparam lut_6479.mask = 64'h0055ffff15414154;

	lut_sub lut_6490 ({sk[1298], i_14_, i_13_, i_12_, i_15_, n_n191}, x923x);
	defparam lut_6490.LUT_SIZE = 6;
	defparam lut_6490.mask = 64'h0055ffff15014154;

	lut_sub lut_6500 ({sk[1299], n_n101, n_n108, x62x, n_n190, x1071x, x1070x}, n_n1201);
	defparam lut_6500.LUT_SIZE = 7;
	defparam lut_6500.mask = 128'h00ff00ffffffffff000055ff3f3f7fff;

	lut_sub lut_6505 ({sk[1300], n_n108, n_n112, n_n60, n_n137, x1894x, x19188x}, x19192x);
	defparam lut_6505.LUT_SIZE = 7;
	defparam lut_6505.mask = 128'h00ff00ffffffffff55555fff77777fff;

	lut_sub lut_6510 ({sk[1301], n_n124, x734x, n_n198, x613x, x1073x, x21409x}, x19193x);
	defparam lut_6510.LUT_SIZE = 7;
	defparam lut_6510.mask = 128'h00ff00ffffffffffafafafafafafbfff;

	lut_sub lut_6515 ({sk[1302], i_14_, i_13_, i_12_, i_15_, n_n199}, x1075x);
	defparam lut_6515.LUT_SIZE = 6;
	defparam lut_6515.mask = 64'h0055ffff15414154;

	lut_sub lut_6526 ({sk[1303], n_n101, n_n108, x86x, n_n190, x1074x, x1535x}, x19200x);
	defparam lut_6526.LUT_SIZE = 7;
	defparam lut_6526.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_6531 ({sk[1304], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1253x);
	defparam lut_6531.LUT_SIZE = 7;
	defparam lut_6531.mask = 128'h00ff00ffffffffff0057000000030000;

	lut_sub lut_6535 ({sk[1305], i_8_, n_n16, x735x, n_n177, x728x, x1253x}, x2558x);
	defparam lut_6535.LUT_SIZE = 7;
	defparam lut_6535.mask = 128'h00ff00ffffffffff0000005700000000;

	lut_sub lut_6538 ({sk[1306], i_9_, i_10_, i_11_, n_n123, x721x, x728x}, x2556x);
	defparam lut_6538.LUT_SIZE = 7;
	defparam lut_6538.mask = 128'h00ff00ffffffffff0700000007000000;

	lut_sub lut_6543 ({sk[1307], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x927x);
	defparam lut_6543.LUT_SIZE = 7;
	defparam lut_6543.mask = 128'h00ff00ffffffffff0000005700003057;

	lut_sub lut_6549 ({sk[1308], i_7_, i_8_, i_6_, x735x, x927x, x2549x}, x19207x);
	defparam lut_6549.LUT_SIZE = 7;
	defparam lut_6549.mask = 128'h00ff00ffffffffff5557555555555555;

	lut_sub lut_6552 ({sk[1309], x735x, n_n126, x2558x, x2556x, x1252x, x1563x}, x19208x);
	defparam lut_6552.LUT_SIZE = 7;
	defparam lut_6552.mask = 128'h00ff00ffffffffff0fff0fff0fff7fff;

	lut_sub lut_6557 ({sk[1310], n_n124, x735x, n_n161, x63x, x841x, x844x}, x21350x);
	defparam lut_6557.LUT_SIZE = 7;
	defparam lut_6557.mask = 128'h00ff00ffffffffffffffffc0ffffaa80;

	lut_sub lut_6563 ({sk[1311], i_14_, i_13_, i_12_, i_15_, n_n216}, x1141x);
	defparam lut_6563.LUT_SIZE = 6;
	defparam lut_6563.mask = 64'h0055ffff00014154;

	lut_sub lut_6570 ({sk[1312], x83x, n_n197, n_n212, n_n125, n_n127, x1141x}, n_n1366);
	defparam lut_6570.LUT_SIZE = 7;
	defparam lut_6570.mask = 128'h00ff00ffffffffff053705370537ffff;

	lut_sub lut_6574 ({sk[1313], i_14_, i_13_, i_12_, i_15_, n_n216}, x1150x);
	defparam lut_6574.LUT_SIZE = 6;
	defparam lut_6574.mask = 64'h0055ffff15414154;

	lut_sub lut_6585 ({sk[1314], i_14_, i_13_, i_12_, i_15_, n_n199}, x1149x);
	defparam lut_6585.LUT_SIZE = 6;
	defparam lut_6585.mask = 64'h0055ffff11014154;

	lut_sub lut_6594 ({sk[1315], i_14_, i_13_, i_12_, i_15_, n_n199}, x1340x);
	defparam lut_6594.LUT_SIZE = 6;
	defparam lut_6594.mask = 64'h0055ffff01014154;

	lut_sub lut_6602 ({sk[1316], n_n197, n_n212, x70x, x1150x, x1149x, x1340x}, x19233x);
	defparam lut_6602.LUT_SIZE = 7;
	defparam lut_6602.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_6607 ({sk[1317], n_n123, n_n125, x52x, x51x, x142x, n_n102}, x19240x);
	defparam lut_6607.LUT_SIZE = 7;
	defparam lut_6607.mask = 128'h00ff00ffffffffff00000fff77777fff;

	lut_sub lut_6612 ({sk[1318], i_14_, i_13_, i_12_, i_15_, n_n191, n_n199}, x1255x);
	defparam lut_6612.LUT_SIZE = 7;
	defparam lut_6612.mask = 128'h00ff00ffffffffff0555500570033330;

	lut_sub lut_6624 ({sk[1319], i_14_, i_13_, i_12_, i_15_, n_n184, n_n216}, x19235x);
	defparam lut_6624.LUT_SIZE = 7;
	defparam lut_6624.mask = 128'h00ff00ffffffffff0000000000070550;

	lut_sub lut_6629 ({sk[1320], n_n124, x735x, n_n126, x251x, x1255x, x19235x}, x19241x);
	defparam lut_6629.LUT_SIZE = 7;
	defparam lut_6629.mask = 128'h00ff00ffffffffff0000003300005f7f;

	lut_sub lut_6633 ({sk[1321], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1559x);
	defparam lut_6633.LUT_SIZE = 7;
	defparam lut_6633.mask = 128'h00ff00ffffffffff0357000057000000;

	lut_sub lut_6639 ({sk[1322], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1558x);
	defparam lut_6639.LUT_SIZE = 7;
	defparam lut_6639.mask = 128'h00ff00ffffffffff5700000000570000;

	lut_sub lut_6644 ({sk[1323], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1561x);
	defparam lut_6644.LUT_SIZE = 7;
	defparam lut_6644.mask = 128'h00ff00ffffffffff5500005700000057;

	lut_sub lut_6650 ({sk[1324], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1560x);
	defparam lut_6650.LUT_SIZE = 7;
	defparam lut_6650.mask = 128'h00ff00ffffffffff0000005757000000;

	lut_sub lut_6655 ({sk[1325], n_n197, n_n212, x1559x, x1558x, x1561x, x1560x}, x19249x);
	defparam lut_6655.LUT_SIZE = 7;
	defparam lut_6655.mask = 128'h00ff00ffffffffff00005f5f33ff7fff;

	lut_sub lut_6660 ({sk[1326], i_14_, i_13_, i_12_, i_15_, n_n170}, x1847x);
	defparam lut_6660.LUT_SIZE = 6;
	defparam lut_6660.mask = 64'h0055ffff11014044;

	lut_sub lut_6667 ({sk[1327], i_14_, i_13_, i_12_, i_15_, n_n170}, x1294x);
	defparam lut_6667.LUT_SIZE = 6;
	defparam lut_6667.mask = 64'h0055ffff15414154;

	lut_sub lut_6678 ({sk[1328], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1293x);
	defparam lut_6678.LUT_SIZE = 7;
	defparam lut_6678.mask = 128'h00ff00ffffffffff0333300330053730;

	lut_sub lut_6690 ({sk[1329], x735x, n_n200, n_n212, x1847x, x1294x, x1293x}, x19269x);
	defparam lut_6690.LUT_SIZE = 7;
	defparam lut_6690.mask = 128'h00ff00ffffffffff005f005f005f337f;

	lut_sub lut_6694 ({sk[1330], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x930x);
	defparam lut_6694.LUT_SIZE = 7;
	defparam lut_6694.mask = 128'h00ff00ffffffffff0555000000003330;

	lut_sub lut_6701 ({sk[1331], x735x, n_n200, n_n212, x63x, x1146x, x1145x}, n_n1217);
	defparam lut_6701.LUT_SIZE = 7;
	defparam lut_6701.mask = 128'h00ff00ffffffffff005f005f005f337f;

	lut_sub lut_6705 ({sk[1332], x735x, n_n200, n_n212, x52x, x1148x, x1147x}, n_n1216);
	defparam lut_6705.LUT_SIZE = 7;
	defparam lut_6705.mask = 128'h00ff00ffffffffff0055005500553f7f;

	lut_sub lut_6709 ({sk[1333], x735x, n_n200, n_n212, x127x, x1290x, x1289x}, n_n1214);
	defparam lut_6709.LUT_SIZE = 7;
	defparam lut_6709.mask = 128'h00ff00ffffffffff0055005500553f7f;

	lut_sub lut_6713 ({sk[1334], x735x, n_n200, n_n212, x133x, x1292x, x1291x}, n_n1213);
	defparam lut_6713.LUT_SIZE = 7;
	defparam lut_6713.mask = 128'h00ff00ffffffffff0055005500553f7f;

	lut_sub lut_6717 ({sk[1335], n_n101, n_n108, x250x, x1892x, x996x, x995x}, n_n1199);
	defparam lut_6717.LUT_SIZE = 7;
	defparam lut_6717.mask = 128'h00ff00ffffffffff00003f3f55ff7fff;

	lut_sub lut_6722 ({sk[1336], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x997x);
	defparam lut_6722.LUT_SIZE = 7;
	defparam lut_6722.mask = 128'h00ff00ffffffffff0333300370057770;

	lut_sub lut_6737 ({sk[1337], x734x, n_n126, x4331x, x4332x, x234x, x998x}, x19294x);
	defparam lut_6737.LUT_SIZE = 7;
	defparam lut_6737.mask = 128'h00ff00ffffffffff0fff0fff0fff7fff;

	lut_sub lut_6742 ({sk[1338], n_n101, n_n108, n_n169, x69x, x250x, x1000x}, x19299x);
	defparam lut_6742.LUT_SIZE = 7;
	defparam lut_6742.mask = 128'h00ff00ffffffffff000077ff0f0f7fff;

	lut_sub lut_6747 ({sk[1339], i_8_, x734x, n_n16, x2488x, x999x, x1142x}, x19300x);
	defparam lut_6747.LUT_SIZE = 7;
	defparam lut_6747.mask = 128'h00ff00ffffffffff0f0f0f7f0f0f0f0f;

	lut_sub lut_6751 ({sk[1340], n_n46, n_n47, x81x, x1214x, x108x, x19319x}, x19324x);
	defparam lut_6751.LUT_SIZE = 7;
	defparam lut_6751.mask = 128'h00ff00ffffffffff000000ff7f7f7fff;

	lut_sub lut_6756 ({sk[1341], n_n101, n_n47, n_n108, n_n129, x378x, x1344x}, x19309x);
	defparam lut_6756.LUT_SIZE = 7;
	defparam lut_6756.mask = 128'h00ff00ffffffffff000f555f333f777f;

	lut_sub lut_6760 ({sk[1342], i_7_, i_8_, i_6_, x734x, x90x, x1408x}, x19316x);
	defparam lut_6760.LUT_SIZE = 7;
	defparam lut_6760.mask = 128'h00ff00ffffffffff0003000500000000;

	lut_sub lut_6763 ({sk[1343], n_n124, x734x, n_n126, x1406x, x19314x, x21351x}, x19317x);
	defparam lut_6763.LUT_SIZE = 7;
	defparam lut_6763.mask = 128'h00ff00ffffffffff0000000f0000bbbf;

	lut_sub lut_6767 ({sk[1344], n_n124, x734x, x450x, n_n129, x19303x, x21433x}, n_n1320);
	defparam lut_6767.LUT_SIZE = 7;
	defparam lut_6767.mask = 128'h00ff00ffffffffffbbffbbffbbffbfff;

	lut_sub lut_6772 ({sk[1345], n_n156, n_n101, x82x, n_n108, x728x, x2470x}, x19308x);
	defparam lut_6772.LUT_SIZE = 7;
	defparam lut_6772.mask = 128'h00ff00ffffffffff555f55ff575f77ff;

	lut_sub lut_6778 ({sk[1346], n_n47, x104x, x3352x, x57x, x4817x, x1506x}, x19332x);
	defparam lut_6778.LUT_SIZE = 7;
	defparam lut_6778.mask = 128'h00ff00ffffffffff33ff33ff7fffffff;

	lut_sub lut_6784 ({sk[1347], n_n89, n_n46, n_n47, x54x, x1509x, x1508x}, n_n1194);
	defparam lut_6784.LUT_SIZE = 7;
	defparam lut_6784.mask = 128'h00ff00ffffffffff00335f7f00ff5fff;

	lut_sub lut_6789 ({sk[1348], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1507x);
	defparam lut_6789.LUT_SIZE = 7;
	defparam lut_6789.mask = 128'h00ff00ffffffffff0333000330037770;

	lut_sub lut_6802 ({sk[1349], x740x, n_n161, n_n47, n_n77, x104x, x1845x}, x19343x);
	defparam lut_6802.LUT_SIZE = 7;
	defparam lut_6802.mask = 128'h00ff00ffffffffff000f000f000f777f;

	lut_sub lut_6806 ({sk[1350], i_8_, x740x, n_n18, n_n47, x1216x, x1215x}, x19344x);
	defparam lut_6806.LUT_SIZE = 7;
	defparam lut_6806.mask = 128'h00ff00ffffffffff0303035703030303;

	lut_sub lut_6809 ({sk[1351], i_15_, x740x, n_n126, x720x, n_n170, n_n213}, x4885x);
	defparam lut_6809.LUT_SIZE = 7;
	defparam lut_6809.mask = 128'h00ff00ffffffffff0000000300000013;

	lut_sub lut_6812 ({sk[1352], i_7_, i_8_, i_6_, x740x, n_n78}, x4886x);
	defparam lut_6812.LUT_SIZE = 6;
	defparam lut_6812.mask = 64'h0055ffff01000000;

	lut_sub lut_6814 ({sk[1353], i_14_, i_13_, i_12_, i_15_, n_n177}, x279x);
	defparam lut_6814.LUT_SIZE = 6;
	defparam lut_6814.mask = 64'h0055ffff00011004;

	lut_sub lut_6818 ({sk[1354], i_9_, i_10_, i_11_, x726x}, n_n171);
	defparam lut_6818.LUT_SIZE = 5;
	defparam lut_6818.mask = 32'h57570010;

	lut_sub lut_6820 ({sk[1355], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x934x);
	defparam lut_6820.LUT_SIZE = 7;
	defparam lut_6820.mask = 128'h00ff00ffffffffff0033000000050000;

	lut_sub lut_6824 ({sk[1356], i_5_, i_3_, i_4_, n_n159, x747x, n_n59}, x527x);
	defparam lut_6824.LUT_SIZE = 7;
	defparam lut_6824.mask = 128'h00ff00ffffffffff0001000000000000;

	lut_sub lut_6826 ({sk[1357], i_7_, i_5_, i_6_, i_3_, i_4_, n_n19}, x551x);
	defparam lut_6826.LUT_SIZE = 7;
	defparam lut_6826.mask = 128'h00ff00ffffffffff1010000000000000;

	lut_sub lut_6829 ({sk[1358], i_14_, i_13_, i_12_, i_15_, n_n170}, n_n131);
	defparam lut_6829.LUT_SIZE = 6;
	defparam lut_6829.mask = 64'h0055ffff00100000;

	lut_sub lut_6831 ({sk[1359], i_9_, i_10_, i_11_, x726x}, n_n143);
	defparam lut_6831.LUT_SIZE = 5;
	defparam lut_6831.mask = 32'h57570400;

	lut_sub lut_6833 ({sk[1360], i_9_, i_10_, i_11_, x728x}, n_n64);
	defparam lut_6833.LUT_SIZE = 5;
	defparam lut_6833.mask = 32'h57570001;

	lut_sub lut_6835 ({sk[1361], i_9_, i_10_, i_11_, i_15_, n_n211}, n_n175);
	defparam lut_6835.LUT_SIZE = 6;
	defparam lut_6835.mask = 64'h0055ffff00000100;

	lut_sub lut_6837 ({sk[1362], i_14_, i_13_, i_12_, i_15_, n_n191}, x1543x);
	defparam lut_6837.LUT_SIZE = 6;
	defparam lut_6837.mask = 64'h0055ffff11114445;

	lut_sub lut_6847 ({sk[1363], i_14_, i_13_, i_12_, i_15_, n_n149, n_n170}, x937x);
	defparam lut_6847.LUT_SIZE = 7;
	defparam lut_6847.mask = 128'h00ff00ffffffffff0535303500000000;

	lut_sub lut_6854 ({sk[1364], i_14_, i_13_, i_12_, i_15_, n_n184}, x242x);
	defparam lut_6854.LUT_SIZE = 6;
	defparam lut_6854.mask = 64'h0055ffff40100400;

	lut_sub lut_6858 ({sk[1365], i_14_, i_13_, i_12_, i_15_, n_n36, n_n199}, x4992x);
	defparam lut_6858.LUT_SIZE = 7;
	defparam lut_6858.mask = 128'h00ff00ffffffffff0000000000000001;

	lut_sub lut_6860 ({sk[1366], n_n36, n_n34, x719x, n_n63, n_n199, x728x}, x709x);
	defparam lut_6860.LUT_SIZE = 7;
	defparam lut_6860.mask = 128'h00ff00ffffffffff000011330f0f1f3f;

	lut_sub lut_6864 ({sk[1367], i_14_, i_13_, i_12_, i_15_, n_n170}, x150x);
	defparam lut_6864.LUT_SIZE = 6;
	defparam lut_6864.mask = 64'h0055ffff40100400;

	lut_sub lut_6868 ({sk[1368], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x941x);
	defparam lut_6868.LUT_SIZE = 7;
	defparam lut_6868.mask = 128'h00ff00ffffffffff5000050000700007;

	lut_sub lut_6875 ({sk[1369], i_9_, i_10_, i_11_, x714x, x17002x, x726x}, n_n6348);
	defparam lut_6875.LUT_SIZE = 7;
	defparam lut_6875.mask = 128'h00ff00ffffffffff0000000000000001;

	lut_sub lut_6877 ({sk[1370], x729x, x714x, x17002x, n_n216, x726x}, x359x);
	defparam lut_6877.LUT_SIZE = 6;
	defparam lut_6877.mask = 64'h0055ffff00010003;

	lut_sub lut_6880 ({sk[1371], n_n41, n_n40, x180x, n_n198, x359x, x219x}, n_n4191);
	defparam lut_6880.LUT_SIZE = 7;
	defparam lut_6880.mask = 128'h00ff00ffffffffff33337f7f33ff7fff;

	lut_sub lut_6885 ({sk[1372], i_7_, i_8_, i_6_, x740x, x392x, n_n52}, n_n1514);
	defparam lut_6885.LUT_SIZE = 7;
	defparam lut_6885.mask = 128'h00ff00ffffffffff3337333733333333;

	lut_sub lut_6889 ({sk[1373], i_7_, i_8_, i_6_, x735x, x68x, x151x}, x21413x);
	defparam lut_6889.LUT_SIZE = 7;
	defparam lut_6889.mask = 128'h00ff00fffffffffff8ffffffffffffff;

	lut_sub lut_6895 ({sk[1374], i_8_, n_n156, x740x, n_n16, x726x, x728x}, x17541x);
	defparam lut_6895.LUT_SIZE = 7;
	defparam lut_6895.mask = 128'h00ff00ffffffffff0000000700000000;

	lut_sub lut_6898 ({sk[1375], i_7_, i_8_, i_6_, x740x, n_n6646, n_n52}, x17542x);
	defparam lut_6898.LUT_SIZE = 7;
	defparam lut_6898.mask = 128'h00ff00ffffffffff3337333733333333;

	lut_sub lut_6902 ({sk[1376], i_7_, i_8_, i_6_, x734x, n_n61, n_n142}, x4838x);
	defparam lut_6902.LUT_SIZE = 7;
	defparam lut_6902.mask = 128'h00ff00ffffffffff0007000000000000;

	lut_sub lut_6905 ({sk[1377], i_14_, i_13_, i_12_, i_15_, n_n199}, x1863x);
	defparam lut_6905.LUT_SIZE = 6;
	defparam lut_6905.mask = 64'h0055ffff40100401;

	lut_sub lut_6910 ({sk[1378], i_7_, i_8_, i_6_, x734x, x4838x, x1863x}, x598x);
	defparam lut_6910.LUT_SIZE = 7;
	defparam lut_6910.mask = 128'h00ff00ffffffffff3333333733333333;

	lut_sub lut_6913 ({sk[1379], i_14_, i_13_, i_12_, i_15_, n_n149}, x204x);
	defparam lut_6913.LUT_SIZE = 6;
	defparam lut_6913.mask = 64'h0055ffff00000401;

	lut_sub lut_6916 ({sk[1380], i_14_, i_13_, i_12_, i_15_, n_n156}, x205x);
	defparam lut_6916.LUT_SIZE = 6;
	defparam lut_6916.mask = 64'h0055ffff11040000;

	lut_sub lut_6920 ({sk[1381], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x944x);
	defparam lut_6920.LUT_SIZE = 7;
	defparam lut_6920.mask = 128'h00ff00ffffffffff0505005000300003;

	lut_sub lut_6926 ({sk[1382], i_7_, i_8_, i_6_, n_n156, x734x, x720x}, x4362x);
	defparam lut_6926.LUT_SIZE = 7;
	defparam lut_6926.mask = 128'h00ff00ffffffffff0001000000000000;

	lut_sub lut_6928 ({sk[1383], i_14_, i_13_, i_12_, i_15_, n_n149}, x220x);
	defparam lut_6928.LUT_SIZE = 6;
	defparam lut_6928.mask = 64'h0055ffff11040000;

	lut_sub lut_6932 ({sk[1384], i_8_, n_n157, x734x, x1449x, x181x, x55x}, x17412x);
	defparam lut_6932.LUT_SIZE = 7;
	defparam lut_6932.mask = 128'h00ff00ffffffffff0000007f00000000;

	lut_sub lut_6936 ({sk[1385], i_14_, i_13_, i_12_, i_15_, n_n149}, x947x);
	defparam lut_6936.LUT_SIZE = 6;
	defparam lut_6936.mask = 64'h0055ffff51155554;

	lut_sub lut_6950 ({sk[1386], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1226x);
	defparam lut_6950.LUT_SIZE = 7;
	defparam lut_6950.mask = 128'h00ff00ffffffffff0333303375057570;

	lut_sub lut_6966 ({sk[1387], i_14_, i_13_, i_12_, i_15_, n_n149}, x1225x);
	defparam lut_6966.LUT_SIZE = 6;
	defparam lut_6966.mask = 64'h0055ffff11015154;

	lut_sub lut_6976 ({sk[1388], i_14_, i_13_, i_12_, i_15_, n_n199}, x1371x);
	defparam lut_6976.LUT_SIZE = 6;
	defparam lut_6976.mask = 64'h0055ffff40100401;

	lut_sub lut_6981 ({sk[1389], i_14_, i_13_, i_12_, i_15_, n_n149}, x1872x);
	defparam lut_6981.LUT_SIZE = 6;
	defparam lut_6981.mask = 64'h0055ffff40100401;

	lut_sub lut_6986 ({sk[1390], i_14_, i_13_, i_12_, i_15_, n_n149, n_n216}, x17429x);
	defparam lut_6986.LUT_SIZE = 7;
	defparam lut_6986.mask = 128'h00ff00ffffffffff3000070000700005;

	lut_sub lut_6993 ({sk[1391], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x949x);
	defparam lut_6993.LUT_SIZE = 7;
	defparam lut_6993.mask = 128'h00ff00ffffffffff3000030000700007;

	lut_sub lut_7000 ({sk[1392], n_n124, x740x, n_n126, n_n84, x104x, x279x}, n_n3864);
	defparam lut_7000.LUT_SIZE = 7;
	defparam lut_7000.mask = 128'h00ff00ffffffffff0000005f0000777f;

	lut_sub lut_7005 ({sk[1393], i_9_, i_10_, i_11_, x729x, x714x, x17002x}, x3506x);
	defparam lut_7005.LUT_SIZE = 7;
	defparam lut_7005.mask = 128'h00ff00ffffffffff0000010000000000;

	lut_sub lut_7007 ({sk[1394], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x952x);
	defparam lut_7007.LUT_SIZE = 7;
	defparam lut_7007.mask = 128'h00ff00ffffffffff0555005557037370;

	lut_sub lut_7022 ({sk[1395], i_14_, i_13_, i_12_, i_15_, n_n184}, x951x);
	defparam lut_7022.LUT_SIZE = 6;
	defparam lut_7022.mask = 64'h0055ffff15455044;

	lut_sub lut_7033 ({sk[1396], n_n89, n_n46, n_n47, x952x, x951x, x54x}, n_n3195);
	defparam lut_7033.LUT_SIZE = 7;
	defparam lut_7033.mask = 128'h00ff00ffffffffff000f777f00ff77ff;

	lut_sub lut_7038 ({sk[1397], i_14_, i_13_, i_12_, i_15_, n_n177}, x1845x);
	defparam lut_7038.LUT_SIZE = 6;
	defparam lut_7038.mask = 64'h0055ffff11014044;

	lut_sub lut_7045 ({sk[1398], i_14_, i_13_, i_12_, i_15_, n_n156}, x1886x);
	defparam lut_7045.LUT_SIZE = 6;
	defparam lut_7045.mask = 64'h0055ffff00005154;

	lut_sub lut_7052 ({sk[1399], i_14_, i_13_, i_12_, i_15_, n_n177}, x1458x);
	defparam lut_7052.LUT_SIZE = 6;
	defparam lut_7052.mask = 64'h0055ffff15454044;

	lut_sub lut_7062 ({sk[1400], i_14_, i_13_, i_12_, i_15_, n_n191}, x1884x);
	defparam lut_7062.LUT_SIZE = 6;
	defparam lut_7062.mask = 64'h0055ffff00005154;

	lut_sub lut_7069 ({sk[1401], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x1531x);
	defparam lut_7069.LUT_SIZE = 7;
	defparam lut_7069.mask = 128'h00ff00ffffffffff0575707555055550;

	lut_sub lut_7085 ({sk[1402], i_14_, i_13_, i_12_, i_15_, n_n191}, x1530x);
	defparam lut_7085.LUT_SIZE = 6;
	defparam lut_7085.mask = 64'h0055ffff04445154;

	lut_sub lut_7095 ({sk[1403], i_14_, i_13_, i_12_, i_15_, n_n170}, x186x);
	defparam lut_7095.LUT_SIZE = 6;
	defparam lut_7095.mask = 64'h0055ffff40100000;

	lut_sub lut_7098 ({sk[1404], i_14_, i_13_, i_12_, i_15_, n_n170}, x209x);
	defparam lut_7098.LUT_SIZE = 6;
	defparam lut_7098.mask = 64'h0055ffff00000401;

	lut_sub lut_7101 ({sk[1405], i_14_, i_13_, i_12_, i_15_, n_n177}, x174x);
	defparam lut_7101.LUT_SIZE = 6;
	defparam lut_7101.mask = 64'h0055ffff40100400;

	lut_sub lut_7105 ({sk[1406], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x1334x);
	defparam lut_7105.LUT_SIZE = 7;
	defparam lut_7105.mask = 128'h00ff00ffffffffff3000030000300007;

	lut_sub lut_7111 ({sk[1407], i_14_, i_13_, i_12_, i_15_, n_n191}, x1333x);
	defparam lut_7111.LUT_SIZE = 6;
	defparam lut_7111.mask = 64'h0055ffff40100401;

	lut_sub lut_7116 ({sk[1408], i_14_, i_13_, i_12_, i_15_, n_n170}, x252x);
	defparam lut_7116.LUT_SIZE = 6;
	defparam lut_7116.mask = 64'h0055ffff00100401;

	lut_sub lut_7120 ({sk[1409], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x18530x);
	defparam lut_7120.LUT_SIZE = 7;
	defparam lut_7120.mask = 128'h00ff00ffffffffff7000030000300003;

	lut_sub lut_7126 ({sk[1410], i_14_, i_13_, i_12_, i_15_, n_n191}, x171x);
	defparam lut_7126.LUT_SIZE = 6;
	defparam lut_7126.mask = 64'h0055ffff00000401;

	lut_sub lut_7129 ({sk[1411], i_7_, i_8_, i_6_, x725x, x735x, n_n216}, x4055x);
	defparam lut_7129.LUT_SIZE = 7;
	defparam lut_7129.mask = 128'h00ff00ffffffffff0001000000000000;

	lut_sub lut_7131 ({sk[1412], i_9_, i_10_, i_11_, x725x, x719x, x721x}, x18535x);
	defparam lut_7131.LUT_SIZE = 7;
	defparam lut_7131.mask = 128'h00ff00ffffffffff000000335f00000f;

	lut_sub lut_7136 ({sk[1413], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x962x);
	defparam lut_7136.LUT_SIZE = 7;
	defparam lut_7136.mask = 128'h00ff00ffffffffff0555505557075750;

	lut_sub lut_7152 ({sk[1414], i_14_, i_13_, i_12_, i_15_, n_n199}, x961x);
	defparam lut_7152.LUT_SIZE = 6;
	defparam lut_7152.mask = 64'h0055ffff04445154;

	lut_sub lut_7162 ({sk[1415], i_14_, i_13_, i_12_, i_15_, n_n156}, x377x);
	defparam lut_7162.LUT_SIZE = 6;
	defparam lut_7162.mask = 64'h0055ffff10044000;

	lut_sub lut_7166 ({sk[1416], i_14_, i_13_, i_12_, i_15_, n_n156}, x964x);
	defparam lut_7166.LUT_SIZE = 6;
	defparam lut_7166.mask = 64'h0055ffff14444000;

	lut_sub lut_7172 ({sk[1417], i_14_, i_13_, i_12_, i_15_, n_n149}, x351x);
	defparam lut_7172.LUT_SIZE = 6;
	defparam lut_7172.mask = 64'h0055ffff10044000;

	lut_sub lut_7176 ({sk[1418], i_14_, i_13_, i_12_, i_15_, n_n149}, x963x);
	defparam lut_7176.LUT_SIZE = 6;
	defparam lut_7176.mask = 64'h0055ffff10045000;

	lut_sub lut_7181 ({sk[1419], i_9_, i_10_, i_11_, i_15_, x717x, n_n211}, x966x);
	defparam lut_7181.LUT_SIZE = 7;
	defparam lut_7181.mask = 128'h00ff00ffffffffff0077770000770000;

	lut_sub lut_7191 ({sk[1420], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x965x);
	defparam lut_7191.LUT_SIZE = 7;
	defparam lut_7191.mask = 128'h00ff00ffffffffff0700000077000000;

	lut_sub lut_7198 ({sk[1421], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x970x);
	defparam lut_7198.LUT_SIZE = 7;
	defparam lut_7198.mask = 128'h00ff00ffffffffff0730303077000000;

	lut_sub lut_7208 ({sk[1422], i_14_, i_13_, i_12_, i_15_, n_n149}, x972x);
	defparam lut_7208.LUT_SIZE = 6;
	defparam lut_7208.mask = 64'h0055ffff14445000;

	lut_sub lut_7215 ({sk[1423], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x971x);
	defparam lut_7215.LUT_SIZE = 7;
	defparam lut_7215.mask = 128'h00ff00ffffffffff0770307077000000;

	lut_sub lut_7227 ({sk[1424], i_9_, i_10_, i_11_, i_15_, x725x, n_n204}, x1177x);
	defparam lut_7227.LUT_SIZE = 7;
	defparam lut_7227.mask = 128'h00ff00ffffffffff0000005033000033;

	lut_sub lut_7231 ({sk[1425], i_9_, i_10_, i_11_, x725x, n_n123, n_n125}, x21394x);
	defparam lut_7231.LUT_SIZE = 7;
	defparam lut_7231.mask = 128'h00ff00ffffffffff0000070000070700;

	lut_sub lut_7240 ({sk[1426], x725x, n_n184, n_n191, x51x, n_n112, n_n113}, x21392x);
	defparam lut_7240.LUT_SIZE = 7;
	defparam lut_7240.mask = 128'h00ff00fffffffffffcfcfcfcfccca888;

	lut_sub lut_7247 ({sk[1427], i_9_, i_8_, n_n18, x285x}, x21456x);
	defparam lut_7247.LUT_SIZE = 5;
	defparam lut_7247.mask = 32'h5757ffef;

	lut_sub lut_7252 ({sk[1428], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x975x);
	defparam lut_7252.LUT_SIZE = 7;
	defparam lut_7252.mask = 128'h00ff00ffffffffff0770707055000000;

	lut_sub lut_7263 ({sk[1429], i_9_, i_10_, i_11_, n_n39, x730x, x726x}, x17288x);
	defparam lut_7263.LUT_SIZE = 7;
	defparam lut_7263.mask = 128'h00ff00ffffffffff0000070000000700;

	lut_sub lut_7268 ({sk[1430], n_n38, n_n39, n_n168, n_n78, n_n84, n_n175}, x21390x);
	defparam lut_7268.LUT_SIZE = 7;
	defparam lut_7268.mask = 128'h00ff00ffffffffffffff8000f0f08000;

	lut_sub lut_7272 ({sk[1431], i_7_, i_8_, i_6_, x740x, n_n168, n_n53}, x21391x);
	defparam lut_7272.LUT_SIZE = 7;
	defparam lut_7272.mask = 128'h00ff00fffffffffffffcfffffaffffff;

	lut_sub lut_7282 ({sk[1432], i_14_, i_13_, i_12_, i_15_, n_n149, n_n216}, x17293x);
	defparam lut_7282.LUT_SIZE = 7;
	defparam lut_7282.mask = 128'h00ff00ffffffffff5030300003000000;

	lut_sub lut_7287 ({sk[1433], x729x, n_n156, x714x, x17002x, x726x}, x363x);
	defparam lut_7287.LUT_SIZE = 6;
	defparam lut_7287.mask = 64'h0055ffff00010003;

	lut_sub lut_7290 ({sk[1434], i_14_, i_13_, i_12_, i_15_, n_n156, n_n216}, x17296x);
	defparam lut_7290.LUT_SIZE = 7;
	defparam lut_7290.mask = 128'h00ff00ffffffffff5300003033000000;

	lut_sub lut_7296 ({sk[1435], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x21389x);
	defparam lut_7296.LUT_SIZE = 7;
	defparam lut_7296.mask = 128'h00ff00fffffffffffc8f8fcfccffffff;

	lut_sub lut_7307 ({sk[1436], i_14_, i_13_, i_12_, i_15_, n_n216}, x977x);
	defparam lut_7307.LUT_SIZE = 6;
	defparam lut_7307.mask = 64'h0055ffff14045000;

	lut_sub lut_7313 ({sk[1437], i_14_, i_13_, i_12_, i_15_, n_n199}, x243x);
	defparam lut_7313.LUT_SIZE = 6;
	defparam lut_7313.mask = 64'h0055ffff14040000;

	lut_sub lut_7317 ({sk[1438], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x17318x);
	defparam lut_7317.LUT_SIZE = 7;
	defparam lut_7317.mask = 128'h00ff00ffffffffff0000700055000000;

	lut_sub lut_7322 ({sk[1439], i_14_, i_13_, i_12_, i_15_, n_n184}, x1235x);
	defparam lut_7322.LUT_SIZE = 6;
	defparam lut_7322.mask = 64'h0055ffff14045000;

	lut_sub lut_7328 ({sk[1440], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x1238x);
	defparam lut_7328.LUT_SIZE = 7;
	defparam lut_7328.mask = 128'h00ff00ffffffffff0770007077000000;

	lut_sub lut_7339 ({sk[1441], i_14_, i_13_, i_12_, i_15_, n_n170}, x982x);
	defparam lut_7339.LUT_SIZE = 6;
	defparam lut_7339.mask = 64'h0055ffff14045000;

	lut_sub lut_7345 ({sk[1442], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x980x);
	defparam lut_7345.LUT_SIZE = 7;
	defparam lut_7345.mask = 128'h00ff00ffffffffff0770007077000000;

	lut_sub lut_7356 ({sk[1443], i_14_, i_13_, i_12_, i_15_, n_n216}, x263x);
	defparam lut_7356.LUT_SIZE = 6;
	defparam lut_7356.mask = 64'h0055ffff10044000;

	lut_sub lut_7360 ({sk[1444], i_8_, x729x, x740x, n_n17, n_n216, x726x}, x361x);
	defparam lut_7360.LUT_SIZE = 7;
	defparam lut_7360.mask = 128'h00ff00ffffffffff0001000300000000;

	lut_sub lut_7363 ({sk[1445], i_14_, i_13_, i_12_, i_15_, n_n191}, x1733x);
	defparam lut_7363.LUT_SIZE = 6;
	defparam lut_7363.mask = 64'h0055ffff10045000;

	lut_sub lut_7368 ({sk[1446], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1794x);
	defparam lut_7368.LUT_SIZE = 7;
	defparam lut_7368.mask = 128'h00ff00ffffffffff0730307077000000;

	lut_sub lut_7379 ({sk[1447], x729x, n_n177, x714x, x17002x, x726x}, x397x);
	defparam lut_7379.LUT_SIZE = 6;
	defparam lut_7379.mask = 64'h0055ffff00010003;

	lut_sub lut_7382 ({sk[1448], n_n65, n_n123, n_n125, x133x, x123x, x175x}, n_n1917);
	defparam lut_7382.LUT_SIZE = 7;
	defparam lut_7382.mask = 128'h00ff00ffffffffff000f777f00ff77ff;

	lut_sub lut_7387 ({sk[1449], i_14_, i_13_, i_12_, i_15_, n_n177}, x991x);
	defparam lut_7387.LUT_SIZE = 6;
	defparam lut_7387.mask = 64'h0055ffff11010050;

	lut_sub lut_7393 ({sk[1450], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x990x);
	defparam lut_7393.LUT_SIZE = 7;
	defparam lut_7393.mask = 128'h00ff00ffffffffff0300300000000500;

	lut_sub lut_7397 ({sk[1451], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x994x);
	defparam lut_7397.LUT_SIZE = 7;
	defparam lut_7397.mask = 128'h00ff00ffffffffff0707700300003300;

	lut_sub lut_7407 ({sk[1452], i_14_, i_13_, i_12_, i_15_, n_n156}, x321x);
	defparam lut_7407.LUT_SIZE = 6;
	defparam lut_7407.mask = 64'h0055ffff00010050;

	lut_sub lut_7411 ({sk[1453], i_9_, i_10_, i_11_, i_15_, n_n201}, x410x);
	defparam lut_7411.LUT_SIZE = 6;
	defparam lut_7411.mask = 64'h0055ffff10000001;

	lut_sub lut_7414 ({sk[1454], i_15_, n_n31, n_n30, n_n199, n_n201}, x2937x);
	defparam lut_7414.LUT_SIZE = 6;
	defparam lut_7414.mask = 64'h0055ffff00000111;

	lut_sub lut_7417 ({sk[1455], n_n30, x994x, x321x, x410x, x2937x}, x18832x);
	defparam lut_7417.LUT_SIZE = 6;
	defparam lut_7417.mask = 64'h0055ffff55557fff;

	lut_sub lut_7422 ({sk[1456], i_14_, i_13_, i_12_, i_15_, n_n177}, x250x);
	defparam lut_7422.LUT_SIZE = 6;
	defparam lut_7422.mask = 64'h0055ffff00014040;

	lut_sub lut_7426 ({sk[1457], i_14_, i_13_, i_12_, i_15_, n_n156}, x1892x);
	defparam lut_7426.LUT_SIZE = 6;
	defparam lut_7426.mask = 64'h0055ffff11014044;

	lut_sub lut_7433 ({sk[1458], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x996x);
	defparam lut_7433.LUT_SIZE = 7;
	defparam lut_7433.mask = 128'h00ff00ffffffffff0555500550035750;

	lut_sub lut_7445 ({sk[1459], i_14_, i_13_, i_12_, i_15_, n_n177}, x995x);
	defparam lut_7445.LUT_SIZE = 6;
	defparam lut_7445.mask = 64'h0055ffff15400114;

	lut_sub lut_7453 ({sk[1460], i_14_, i_13_, i_12_, i_15_, n_n149}, x998x);
	defparam lut_7453.LUT_SIZE = 6;
	defparam lut_7453.mask = 64'h0055ffff15400114;

	lut_sub lut_7461 ({sk[1461], i_14_, i_13_, i_12_, i_15_, n_n177, n_n108}, x2488x);
	defparam lut_7461.LUT_SIZE = 7;
	defparam lut_7461.mask = 128'h00ff00ffffffffff0000000000010110;

	lut_sub lut_7465 ({sk[1462], i_14_, i_13_, i_12_, i_15_, n_n177}, x1000x);
	defparam lut_7465.LUT_SIZE = 6;
	defparam lut_7465.mask = 64'h0055ffff15400000;

	lut_sub lut_7470 ({sk[1463], i_14_, i_13_, i_12_, i_15_, n_n170}, x999x);
	defparam lut_7470.LUT_SIZE = 6;
	defparam lut_7470.mask = 64'h0055ffff11014154;

	lut_sub lut_7479 ({sk[1464], i_7_, i_8_, i_6_, x740x, x248x}, n_n4279);
	defparam lut_7479.LUT_SIZE = 6;
	defparam lut_7479.mask = 64'h0055ffff01000000;

	lut_sub lut_7481 ({sk[1465], i_14_, i_13_, i_12_, i_15_, n_n216}, x1001x);
	defparam lut_7481.LUT_SIZE = 6;
	defparam lut_7481.mask = 64'h0055ffff15014154;

	lut_sub lut_7491 ({sk[1466], i_7_, i_8_, i_6_, n_n156, x740x, x726x}, x495x);
	defparam lut_7491.LUT_SIZE = 7;
	defparam lut_7491.mask = 128'h00ff00ffffffffff0001000000000000;

	lut_sub lut_7493 ({sk[1467], i_14_, i_13_, i_12_, i_15_, n_n149}, x249x);
	defparam lut_7493.LUT_SIZE = 6;
	defparam lut_7493.mask = 64'h0055ffff01004040;

	lut_sub lut_7497 ({sk[1468], i_14_, i_13_, i_12_, i_15_, n_n156}, x110x);
	defparam lut_7497.LUT_SIZE = 6;
	defparam lut_7497.mask = 64'h0055ffff00000104;

	lut_sub lut_7500 ({sk[1469], i_7_, i_8_, i_6_, x740x, x110x}, x647x);
	defparam lut_7500.LUT_SIZE = 6;
	defparam lut_7500.mask = 64'h0055ffff01000000;

	lut_sub lut_7502 ({sk[1470], i_7_, i_8_, i_6_, x740x, x207x, n_n143}, x457x);
	defparam lut_7502.LUT_SIZE = 7;
	defparam lut_7502.mask = 128'h00ff00ffffffffff0005000300000000;

	lut_sub lut_7505 ({sk[1471], i_7_, i_8_, i_6_, x740x, x110x}, x572x);
	defparam lut_7505.LUT_SIZE = 6;
	defparam lut_7505.mask = 64'h0055ffff00010000;

	lut_sub lut_7507 ({sk[1472], i_14_, i_13_, i_12_, i_15_, n_n149, n_n177}, x1002x);
	defparam lut_7507.LUT_SIZE = 7;
	defparam lut_7507.mask = 128'h00ff00ffffffffff0003000530053550;

	lut_sub lut_7515 ({sk[1473], n_n39, n_n150, n_n82, n_n170, n_n166, x727x}, x21431x);
	defparam lut_7515.LUT_SIZE = 7;
	defparam lut_7515.mask = 128'h00ff00ffffffffffffffffffc8000000;

	lut_sub lut_7519 ({sk[1474], i_14_, i_13_, i_12_, i_15_, n_n199}, x1005x);
	defparam lut_7519.LUT_SIZE = 6;
	defparam lut_7519.mask = 64'h0055ffff15414054;

	lut_sub lut_7529 ({sk[1475], i_14_, i_13_, i_12_, i_15_, n_n216}, x233x);
	defparam lut_7529.LUT_SIZE = 6;
	defparam lut_7529.mask = 64'h0055ffff00000114;

	lut_sub lut_7533 ({sk[1476], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1007x);
	defparam lut_7533.LUT_SIZE = 7;
	defparam lut_7533.mask = 128'h00ff00ffffffffff0777300770057570;

	lut_sub lut_7551 ({sk[1477], i_14_, i_13_, i_12_, i_15_, n_n177}, x1006x);
	defparam lut_7551.LUT_SIZE = 6;
	defparam lut_7551.mask = 64'h0055ffff15414154;

	lut_sub lut_7562 ({sk[1478], i_14_, i_13_, i_12_, i_15_, n_n216}, x1009x);
	defparam lut_7562.LUT_SIZE = 6;
	defparam lut_7562.mask = 64'h0055ffff00011114;

	lut_sub lut_7568 ({sk[1479], i_9_, i_10_, i_11_, i_15_, n_n207}, x340x);
	defparam lut_7568.LUT_SIZE = 6;
	defparam lut_7568.mask = 64'h0055ffff50000000;

	lut_sub lut_7571 ({sk[1480], i_14_, i_13_, i_12_, i_15_, n_n191}, x187x);
	defparam lut_7571.LUT_SIZE = 6;
	defparam lut_7571.mask = 64'h0055ffff00001014;

	lut_sub lut_7575 ({sk[1481], i_14_, i_13_, i_12_, i_15_, n_n191}, x1010x);
	defparam lut_7575.LUT_SIZE = 6;
	defparam lut_7575.mask = 64'h0055ffff00051014;

	lut_sub lut_7581 ({sk[1482], n_n138, n_n42, n_n43, n_n190, x340x, x1010x}, n_n832);
	defparam lut_7581.LUT_SIZE = 7;
	defparam lut_7581.mask = 128'h00ff00ffffffffff00335f7f00ff5fff;

	lut_sub lut_7586 ({sk[1483], i_14_, i_13_, i_12_, i_15_, n_n191}, x1015x);
	defparam lut_7586.LUT_SIZE = 6;
	defparam lut_7586.mask = 64'h0055ffff00051114;

	lut_sub lut_7593 ({sk[1484], i_14_, i_13_, i_12_, i_15_, n_n184, n_n216}, x1014x);
	defparam lut_7593.LUT_SIZE = 7;
	defparam lut_7593.mask = 128'h00ff00ffffffffff0000005000030300;

	lut_sub lut_7597 ({sk[1485], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1017x);
	defparam lut_7597.LUT_SIZE = 7;
	defparam lut_7597.mask = 128'h00ff00ffffffffff0000003707070770;

	lut_sub lut_7609 ({sk[1486], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1016x);
	defparam lut_7609.LUT_SIZE = 7;
	defparam lut_7609.mask = 128'h00ff00ffffffffff0000007303030330;

	lut_sub lut_7617 ({sk[1487], n_n101, n_n108, x1015x, x1014x, x1017x, x1016x}, n_n777);
	defparam lut_7617.LUT_SIZE = 7;
	defparam lut_7617.mask = 128'h00ff00ffffffffff000055ff3f3f7fff;

	lut_sub lut_7622 ({sk[1488], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x18782x);
	defparam lut_7622.LUT_SIZE = 7;
	defparam lut_7622.mask = 128'h00ff00ffffffffff0000070000700007;

	lut_sub lut_7629 ({sk[1489], i_14_, i_13_, i_12_, i_15_, n_n184, n_n170}, x1022x);
	defparam lut_7629.LUT_SIZE = 7;
	defparam lut_7629.mask = 128'h00ff00ffffffffff7000070000700007;

	lut_sub lut_7638 ({sk[1490], i_14_, i_13_, i_12_, i_15_, n_n177}, x1263x);
	defparam lut_7638.LUT_SIZE = 6;
	defparam lut_7638.mask = 64'h0055ffff40100401;

	lut_sub lut_7643 ({sk[1491], i_14_, i_13_, i_12_, i_15_, n_n177}, x224x);
	defparam lut_7643.LUT_SIZE = 6;
	defparam lut_7643.mask = 64'h0055ffff11040000;

	lut_sub lut_7647 ({sk[1492], i_14_, i_13_, i_12_, i_15_, n_n177}, x57x);
	defparam lut_7647.LUT_SIZE = 6;
	defparam lut_7647.mask = 64'h0055ffff04400000;

	lut_sub lut_7650 ({sk[1493], i_7_, i_8_, i_6_, x734x, n_n83, n_n171}, x617x);
	defparam lut_7650.LUT_SIZE = 7;
	defparam lut_7650.mask = 128'h00ff00ffffffffff0007000000000000;

	lut_sub lut_7653 ({sk[1494], i_14_, i_13_, i_12_, i_15_, n_n177}, x100x);
	defparam lut_7653.LUT_SIZE = 6;
	defparam lut_7653.mask = 64'h0055ffff00001014;

	lut_sub lut_7657 ({sk[1495], n_n124, x734x, n_n126, x69x, n_n176, x100x}, x618x);
	defparam lut_7657.LUT_SIZE = 7;
	defparam lut_7657.mask = 128'h00ff00ffffffffff0000000f0000777f;

	lut_sub lut_7661 ({sk[1496], i_14_, i_13_, i_12_, i_15_, n_n156}, x1025x);
	defparam lut_7661.LUT_SIZE = 6;
	defparam lut_7661.mask = 64'h0055ffff11055054;

	lut_sub lut_7671 ({sk[1497], n_n101, n_n108, x90x, n_n142, x141x, x598x}, x18641x);
	defparam lut_7671.LUT_SIZE = 7;
	defparam lut_7671.mask = 128'h00ff00ffffffffff55557f7f55ff7fff;

	lut_sub lut_7676 ({sk[1498], i_8_, x734x, n_n16, x218x, x141x, x1025x}, x18642x);
	defparam lut_7676.LUT_SIZE = 7;
	defparam lut_7676.mask = 128'h00ff00ffffffffff0000007f00000000;

	lut_sub lut_7680 ({sk[1499], i_7_, i_8_, i_6_, x734x, x80x}, x4190x);
	defparam lut_7680.LUT_SIZE = 6;
	defparam lut_7680.mask = 64'h0055ffff00010000;

	lut_sub lut_7682 ({sk[1500], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x18648x);
	defparam lut_7682.LUT_SIZE = 7;
	defparam lut_7682.mask = 128'h00ff00ffffffffff3000070000700005;

	lut_sub lut_7689 ({sk[1501], i_14_, i_13_, i_12_, i_15_, n_n184, n_n170}, x18644x);
	defparam lut_7689.LUT_SIZE = 7;
	defparam lut_7689.mask = 128'h00ff00ffffffffff5000050000700003;

	lut_sub lut_7695 ({sk[1502], n_n59, n_n116, n_n108, x78x, x18648x, x252x}, x3111x);
	defparam lut_7695.LUT_SIZE = 7;
	defparam lut_7695.mask = 128'h00ff00ffffffffff007f00ff00ff00ff;

	lut_sub lut_7701 ({sk[1503], i_14_, i_13_, i_12_, i_15_, n_n184, n_n170}, x18643x);
	defparam lut_7701.LUT_SIZE = 7;
	defparam lut_7701.mask = 128'h00ff00ffffffffff3000030000000005;

	lut_sub lut_7705 ({sk[1504], n_n101, n_n59, x4190x, x18644x, x222x, x18643x}, x18650x);
	defparam lut_7705.LUT_SIZE = 7;
	defparam lut_7705.mask = 128'h00ff00ffffffffff00ff00ff7fffffff;

	lut_sub lut_7711 ({sk[1505], i_14_, i_13_, i_12_, i_15_, n_n149}, x1028x);
	defparam lut_7711.LUT_SIZE = 6;
	defparam lut_7711.mask = 64'h0055ffff11054040;

	lut_sub lut_7718 ({sk[1506], n_n108, x4331x, x4332x, x60x, x4329x, x4362x}, x18652x);
	defparam lut_7718.LUT_SIZE = 7;
	defparam lut_7718.mask = 128'h00ff00ffffffffff77ffffff7fffffff;

	lut_sub lut_7724 ({sk[1507], n_n101, n_n108, x60x, x84x, x220x, x1028x}, x21434x);
	defparam lut_7724.LUT_SIZE = 7;
	defparam lut_7724.mask = 128'h00ff00ffffffffffffffc0c0aa008000;

	lut_sub lut_7729 ({sk[1508], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1031x);
	defparam lut_7729.LUT_SIZE = 7;
	defparam lut_7729.mask = 128'h00ff00ffffffffff0757507333033330;

	lut_sub lut_7745 ({sk[1509], i_14_, i_13_, i_12_, i_15_, n_n170}, x1030x);
	defparam lut_7745.LUT_SIZE = 6;
	defparam lut_7745.mask = 64'h0055ffff15455154;

	lut_sub lut_7758 ({sk[1510], i_14_, i_13_, i_12_, i_15_, n_n149}, x1173x);
	defparam lut_7758.LUT_SIZE = 6;
	defparam lut_7758.mask = 64'h0055ffff11055154;

	lut_sub lut_7769 ({sk[1511], x740x, n_n200, x180x, x361x, x363x, x1173x}, x17530x);
	defparam lut_7769.LUT_SIZE = 7;
	defparam lut_7769.mask = 128'h00ff00ffffffffff3f3f3f3f3f3f7fff;

	lut_sub lut_7774 ({sk[1512], n_n41, n_n40, n_n155, x215x, x60x, x220x}, x17533x);
	defparam lut_7774.LUT_SIZE = 7;
	defparam lut_7774.mask = 128'h00ff00ffffffffff00000fff77777fff;

	lut_sub lut_7779 ({sk[1513], i_15_, x714x, x17002x, n_n199, n_n201, n_n204}, x4905x);
	defparam lut_7779.LUT_SIZE = 7;
	defparam lut_7779.mask = 128'h00ff00ffffffffff0000000500000003;

	lut_sub lut_7782 ({sk[1514], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1034x);
	defparam lut_7782.LUT_SIZE = 7;
	defparam lut_7782.mask = 128'h00ff00ffffffffff7000070000700007;

	lut_sub lut_7791 ({sk[1515], i_14_, i_13_, i_12_, i_15_, n_n149}, x173x);
	defparam lut_7791.LUT_SIZE = 6;
	defparam lut_7791.mask = 64'h0055ffff40100000;

	lut_sub lut_7794 ({sk[1516], i_14_, i_13_, i_12_, i_15_, n_n216}, x1867x);
	defparam lut_7794.LUT_SIZE = 6;
	defparam lut_7794.mask = 64'h0055ffff40100401;

	lut_sub lut_7799 ({sk[1517], n_n40, x204x, x173x, n_n4604, x1103x, x4909x}, x17537x);
	defparam lut_7799.LUT_SIZE = 7;
	defparam lut_7799.mask = 128'h00ff00ffffffffff5f5f5f5f7fffffff;

	lut_sub lut_7805 ({sk[1518], n_n41, n_n40, x1034x, x153x, x1867x, x17537x}, x17539x);
	defparam lut_7805.LUT_SIZE = 7;
	defparam lut_7805.mask = 128'h00ff00ffffffffff555577775fff7fff;

	lut_sub lut_7810 ({sk[1519], n_n41, n_n40, n_n148, x90x, x60x, n_n142}, x17531x);
	defparam lut_7810.LUT_SIZE = 7;
	defparam lut_7810.mask = 128'h00ff00ffffffffff00003f3f55ff7fff;

	lut_sub lut_7815 ({sk[1520], n_n41, n_n40, x155x, x205x, x1819x, x1880x}, x21386x);
	defparam lut_7815.LUT_SIZE = 7;
	defparam lut_7815.mask = 128'h00ff00fffffffffffffff00080008000;

	lut_sub lut_7819 ({sk[1521], x17530x, x17533x, x17531x, x21386x}, x17540x);
	defparam lut_7819.LUT_SIZE = 5;
	defparam lut_7819.mask = 32'h5757bfff;

	lut_sub lut_7824 ({sk[1522], i_14_, i_13_, i_12_, i_15_, n_n156}, x1852x);
	defparam lut_7824.LUT_SIZE = 6;
	defparam lut_7824.mask = 64'h0055ffff40100401;

	lut_sub lut_7829 ({sk[1523], n_n124, x740x, n_n4461, x249x, x457x, x620x}, x17552x);
	defparam lut_7829.LUT_SIZE = 7;
	defparam lut_7829.mask = 128'h00ff00ffffffffff77ff77ff77ff7fff;

	lut_sub lut_7834 ({sk[1524], n_n39, n_n40, n_n150, x4283x, x110x, x1852x}, x17548x);
	defparam lut_7834.LUT_SIZE = 7;
	defparam lut_7834.mask = 128'h00ff00ffffffffff0f0f5f5f3fff7fff;

	lut_sub lut_7839 ({sk[1525], n_n38, n_n39, x248x, n_n143, x249x, x110x}, x17549x);
	defparam lut_7839.LUT_SIZE = 7;
	defparam lut_7839.mask = 128'h00ff00ffffffffff00003fff55ff7fff;

	lut_sub lut_7845 ({sk[1526], n_n1514, x597x, x17541x, x17542x, x17548x, x17549x}, x17553x);
	defparam lut_7845.LUT_SIZE = 7;
	defparam lut_7845.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_7852 ({sk[1527], n_n46, n_n47, x218x, x141x, x17554x, x1823x}, x17557x);
	defparam lut_7852.LUT_SIZE = 7;
	defparam lut_7852.mask = 128'h00ff00ffffffffff33333f3f77ff7fff;

	lut_sub lut_7857 ({sk[1528], x714x, x17002x, x720x, x85x, x142x, n_n216}, x549x);
	defparam lut_7857.LUT_SIZE = 7;
	defparam lut_7857.mask = 128'h00ff00ffffffffff0000000000003f7f;

	lut_sub lut_7861 ({sk[1529], n_n41, n_n40, x70x, x85x, x142x, n_n198}, x17008x);
	defparam lut_7861.LUT_SIZE = 7;
	defparam lut_7861.mask = 128'h00ff00ffffffffff00003fff55ff7fff;

	lut_sub lut_7867 ({sk[1530], i_14_, i_13_, i_12_, i_15_, n_n199}, x1107x);
	defparam lut_7867.LUT_SIZE = 6;
	defparam lut_7867.mask = 64'h0055ffff11055054;

	lut_sub lut_7877 ({sk[1531], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1868x);
	defparam lut_7877.LUT_SIZE = 7;
	defparam lut_7877.mask = 128'h00ff00ffffffffff0303003330053000;

	lut_sub lut_7885 ({sk[1532], x740x, n_n200, x714x, x17002x, x1107x, x1868x}, x17009x);
	defparam lut_7885.LUT_SIZE = 7;
	defparam lut_7885.mask = 128'h00ff00ffffffffff0003000300035557;

	lut_sub lut_7888 ({sk[1533], n_n41, n_n214, x85x, x142x, n_n4191, x17562x}, x17564x);
	defparam lut_7888.LUT_SIZE = 7;
	defparam lut_7888.mask = 128'h00ff00ffffffffff777777777fffffff;

	lut_sub lut_7894 ({sk[1534], x17557x, x17008x, x17009x, n_n4195, x17556x}, x17565x);
	defparam lut_7894.LUT_SIZE = 6;
	defparam lut_7894.mask = 64'h0055ffff7fffffff;

	lut_sub lut_7900 ({sk[1535], i_14_, i_13_, i_12_, i_15_, n_n216}, x1035x);
	defparam lut_7900.LUT_SIZE = 6;
	defparam lut_7900.mask = 64'h0055ffff15454000;

	lut_sub lut_7908 ({sk[1536], i_8_, x740x, n_n18, n_n47, x98x, x1035x}, n_n3257);
	defparam lut_7908.LUT_SIZE = 7;
	defparam lut_7908.mask = 128'h00ff00ffffffffff0303035703030303;

	lut_sub lut_7911 ({sk[1537], i_9_, i_10_, i_11_, x729x, x714x, x17002x}, x3523x);
	defparam lut_7911.LUT_SIZE = 7;
	defparam lut_7911.mask = 128'h00ff00ffffffffff0100000000000000;

	lut_sub lut_7913 ({sk[1538], i_14_, i_13_, i_12_, i_15_, n_n184, n_n216}, x1037x);
	defparam lut_7913.LUT_SIZE = 7;
	defparam lut_7913.mask = 128'h00ff00ffffffffff0507005773033330;

	lut_sub lut_7927 ({sk[1539], i_14_, i_13_, i_12_, i_15_, n_n191}, x1036x);
	defparam lut_7927.LUT_SIZE = 6;
	defparam lut_7927.mask = 64'h0055ffff15455044;

	lut_sub lut_7938 ({sk[1540], n_n41, n_n40, n_n102, x98x, n_n6384, x1036x}, x18232x);
	defparam lut_7938.LUT_SIZE = 7;
	defparam lut_7938.mask = 128'h00ff00ffffffffff333333ff7f7f7fff;

	lut_sub lut_7943 ({sk[1541], i_7_, i_8_, i_6_, x740x, x81x}, x3542x);
	defparam lut_7943.LUT_SIZE = 6;
	defparam lut_7943.mask = 64'h0055ffff00001000;

	lut_sub lut_7945 ({sk[1542], i_9_, i_10_, i_11_, x729x, x714x, x17002x}, x3543x);
	defparam lut_7945.LUT_SIZE = 7;
	defparam lut_7945.mask = 128'h00ff00ffffffffff0000000000000001;

	lut_sub lut_7947 ({sk[1543], i_15_, x714x, x17002x, x720x, n_n216, n_n213}, x391x);
	defparam lut_7947.LUT_SIZE = 7;
	defparam lut_7947.mask = 128'h00ff00ffffffffff0000000300000013;

	lut_sub lut_7950 ({sk[1544], i_14_, i_13_, i_12_, i_15_, n_n216}, x1038x);
	defparam lut_7950.LUT_SIZE = 6;
	defparam lut_7950.mask = 64'h0055ffff11055044;

	lut_sub lut_7959 ({sk[1545], n_n4308, x512x, n_n6348, x3542x, x3543x, x391x}, x18237x);
	defparam lut_7959.LUT_SIZE = 7;
	defparam lut_7959.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_7966 ({sk[1546], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1040x);
	defparam lut_7966.LUT_SIZE = 7;
	defparam lut_7966.mask = 128'h00ff00ffffffffff0333003337057570;

	lut_sub lut_7981 ({sk[1547], i_14_, i_13_, i_12_, i_15_, n_n199}, x1039x);
	defparam lut_7981.LUT_SIZE = 6;
	defparam lut_7981.mask = 64'h0055ffff14440000;

	lut_sub lut_7986 ({sk[1548], n_n3085, n_n40, x714x, x17002x, x1037x, x1038x}, x21371x);
	defparam lut_7986.LUT_SIZE = 7;
	defparam lut_7986.mask = 128'h00ff00fffffffffffffaccc800000000;

	lut_sub lut_7993 ({sk[1549], n_n41, n_n40, n_n95, x1040x, x1039x, x1272x}, x21372x);
	defparam lut_7993.LUT_SIZE = 7;
	defparam lut_7993.mask = 128'h00ff00fffffffffffffff00088888000;

	lut_sub lut_7998 ({sk[1550], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x17373x);
	defparam lut_7998.LUT_SIZE = 7;
	defparam lut_7998.mask = 128'h00ff00ffffffffff0700000077000000;

	lut_sub lut_8005 ({sk[1551], i_14_, i_13_, i_12_, i_15_, n_n184}, x17371x);
	defparam lut_8005.LUT_SIZE = 6;
	defparam lut_8005.mask = 64'h0055ffff14445000;

	lut_sub lut_8012 ({sk[1552], i_9_, i_10_, i_11_, x725x, n_n42, n_n43}, x526x);
	defparam lut_8012.LUT_SIZE = 7;
	defparam lut_8012.mask = 128'h00ff00ffffffffff0500000003000000;

	lut_sub lut_8015 ({sk[1553], i_15_, x714x, x17002x, n_n216, n_n211}, x632x);
	defparam lut_8015.LUT_SIZE = 6;
	defparam lut_8015.mask = 64'h0055ffff00000001;

	lut_sub lut_8017 ({sk[1554], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1052x);
	defparam lut_8017.LUT_SIZE = 7;
	defparam lut_8017.mask = 128'h00ff00ffffffffff0330303037000000;

	lut_sub lut_8025 ({sk[1555], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1051x);
	defparam lut_8025.LUT_SIZE = 7;
	defparam lut_8025.mask = 128'h00ff00ffffffffff0700007073000000;

	lut_sub lut_8033 ({sk[1556], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x17354x);
	defparam lut_8033.LUT_SIZE = 7;
	defparam lut_8033.mask = 128'h00ff00ffffffffff0500005057000000;

	lut_sub lut_8039 ({sk[1557], i_14_, i_13_, i_12_, i_15_, n_n184, n_n170}, x17351x);
	defparam lut_8039.LUT_SIZE = 7;
	defparam lut_8039.mask = 128'h00ff00ffffffffff0300003037000000;

	lut_sub lut_8045 ({sk[1558], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x21402x);
	defparam lut_8045.LUT_SIZE = 7;
	defparam lut_8045.mask = 128'h00ff00fffffffffffa8f8fafaaffffff;

	lut_sub lut_8056 ({sk[1559], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1061x);
	defparam lut_8056.LUT_SIZE = 7;
	defparam lut_8056.mask = 128'h00ff00ffffffffff0550505057000000;

	lut_sub lut_8064 ({sk[1560], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1060x);
	defparam lut_8064.LUT_SIZE = 7;
	defparam lut_8064.mask = 128'h00ff00ffffffffff0750507073000000;

	lut_sub lut_8074 ({sk[1561], i_14_, i_13_, i_12_, i_15_, n_n199}, x1065x);
	defparam lut_8074.LUT_SIZE = 6;
	defparam lut_8074.mask = 64'h0055ffff14445000;

	lut_sub lut_8081 ({sk[1562], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1064x);
	defparam lut_8081.LUT_SIZE = 7;
	defparam lut_8081.mask = 128'h00ff00ffffffffff0770707073000000;

	lut_sub lut_8093 ({sk[1563], i_9_, i_10_, i_11_, i_15_, n_n211, x1065x}, x1063x);
	defparam lut_8093.LUT_SIZE = 7;
	defparam lut_8093.mask = 128'h00ff00ffffffffff5555555555555557;

	lut_sub lut_8096 ({sk[1564], i_14_, i_13_, i_12_, i_15_, n_n216}, x1066x);
	defparam lut_8096.LUT_SIZE = 6;
	defparam lut_8096.mask = 64'h0055ffff15014040;

	lut_sub lut_8103 ({sk[1565], i_14_, i_13_, i_12_, i_15_, n_n177}, x1067x);
	defparam lut_8103.LUT_SIZE = 6;
	defparam lut_8103.mask = 64'h0055ffff15414000;

	lut_sub lut_8110 ({sk[1566], i_14_, i_13_, i_12_, i_15_, n_n177}, x1069x);
	defparam lut_8110.LUT_SIZE = 6;
	defparam lut_8110.mask = 64'h0055ffff15414154;

	lut_sub lut_8121 ({sk[1567], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1068x);
	defparam lut_8121.LUT_SIZE = 7;
	defparam lut_8121.mask = 128'h00ff00ffffffffff0050500330033330;

	lut_sub lut_8130 ({sk[1568], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1071x);
	defparam lut_8130.LUT_SIZE = 7;
	defparam lut_8130.mask = 128'h00ff00ffffffffff0333300330037770;

	lut_sub lut_8144 ({sk[1569], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1070x);
	defparam lut_8144.LUT_SIZE = 7;
	defparam lut_8144.mask = 128'h00ff00ffffffffff0753500330033330;

	lut_sub lut_8156 ({sk[1570], i_7_, i_8_, i_6_, x285x}, n_n109);
	defparam lut_8156.LUT_SIZE = 5;
	defparam lut_8156.mask = 32'h57570001;

	lut_sub lut_8158 ({sk[1571], i_9_, i_10_, i_11_, i_15_, n_n113, n_n201}, x613x);
	defparam lut_8158.LUT_SIZE = 7;
	defparam lut_8158.mask = 128'h00ff00ffffffffff0100000000000000;

	lut_sub lut_8160 ({sk[1572], i_14_, i_13_, i_12_, i_15_, n_n216}, x1894x);
	defparam lut_8160.LUT_SIZE = 6;
	defparam lut_8160.mask = 64'h0055ffff11014044;

	lut_sub lut_8167 ({sk[1573], i_9_, i_10_, i_8_, i_11_, n_n18, x285x}, x760x);
	defparam lut_8167.LUT_SIZE = 7;
	defparam lut_8167.mask = 128'h00ff00ffffffffff0010000100000000;

	lut_sub lut_8170 ({sk[1574], i_14_, i_13_, i_12_, i_15_, n_n199}, x1073x);
	defparam lut_8170.LUT_SIZE = 6;
	defparam lut_8170.mask = 64'h0055ffff15414054;

	lut_sub lut_8180 ({sk[1575], i_9_, i_10_, i_8_, i_11_, n_n18, x285x}, x19188x);
	defparam lut_8180.LUT_SIZE = 7;
	defparam lut_8180.mask = 128'h00ff00ffffffffff0011001100000000;

	lut_sub lut_8185 ({sk[1576], i_7_, i_8_, i_6_, x734x, x86x, x111x}, x21409x);
	defparam lut_8185.LUT_SIZE = 7;
	defparam lut_8185.mask = 128'h00ff00fffffffffffffffff8ffffffff;

	lut_sub lut_8191 ({sk[1577], i_14_, i_13_, i_12_, i_15_, n_n216}, x1074x);
	defparam lut_8191.LUT_SIZE = 6;
	defparam lut_8191.mask = 64'h0055ffff11014154;

	lut_sub lut_8200 ({sk[1578], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1077x);
	defparam lut_8200.LUT_SIZE = 7;
	defparam lut_8200.mask = 128'h00ff00ffffffffff0030300550075750;

	lut_sub lut_8211 ({sk[1579], i_14_, i_13_, i_12_, i_15_, n_n177}, x1076x);
	defparam lut_8211.LUT_SIZE = 6;
	defparam lut_8211.mask = 64'h0055ffff15414054;

	lut_sub lut_8221 ({sk[1580], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1079x);
	defparam lut_8221.LUT_SIZE = 7;
	defparam lut_8221.mask = 128'h00ff00ffffffffff0373500330033330;

	lut_sub lut_8233 ({sk[1581], i_14_, i_13_, i_12_, i_15_, n_n184}, x1078x);
	defparam lut_8233.LUT_SIZE = 6;
	defparam lut_8233.mask = 64'h0055ffff15414054;

	lut_sub lut_8243 ({sk[1582], i_14_, i_13_, i_12_, i_15_, n_n170}, x1081x);
	defparam lut_8243.LUT_SIZE = 6;
	defparam lut_8243.mask = 64'h0055ffff04400110;

	lut_sub lut_8248 ({sk[1583], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1080x);
	defparam lut_8248.LUT_SIZE = 7;
	defparam lut_8248.mask = 128'h00ff00ffffffffff0555000000003330;

	lut_sub lut_8255 ({sk[1584], i_9_, i_10_, i_11_, i_15_, n_n201}, x19413x);
	defparam lut_8255.LUT_SIZE = 6;
	defparam lut_8255.mask = 64'h0055ffff10000040;

	lut_sub lut_8258 ({sk[1585], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x19414x);
	defparam lut_8258.LUT_SIZE = 7;
	defparam lut_8258.mask = 128'h00ff00ffffffffff5500000000000057;

	lut_sub lut_8262 ({sk[1586], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1210x);
	defparam lut_8262.LUT_SIZE = 7;
	defparam lut_8262.mask = 128'h00ff00ffffffffff5700005757000057;

	lut_sub lut_8271 ({sk[1587], i_14_, i_13_, i_12_, i_15_, n_n149}, x315x);
	defparam lut_8271.LUT_SIZE = 6;
	defparam lut_8271.mask = 64'h0055ffff14400000;

	lut_sub lut_8275 ({sk[1588], i_9_, i_10_, i_11_, n_n41, x721x, x728x}, x2373x);
	defparam lut_8275.LUT_SIZE = 7;
	defparam lut_8275.mask = 128'h00ff00ffffffffff0000070000000700;

	lut_sub lut_8280 ({sk[1589], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1557x);
	defparam lut_8280.LUT_SIZE = 7;
	defparam lut_8280.mask = 128'h00ff00ffffffffff0057000000550000;

	lut_sub lut_8284 ({sk[1590], i_15_, n_n177, x714x, x17002x, n_n201, x1557x}, x2371x);
	defparam lut_8284.LUT_SIZE = 7;
	defparam lut_8284.mask = 128'h00ff00ffffffffff0005000500050007;

	lut_sub lut_8287 ({sk[1591], i_14_, i_13_, i_12_, i_15_, n_n216}, x1085x);
	defparam lut_8287.LUT_SIZE = 6;
	defparam lut_8287.mask = 64'h0055ffff00011114;

	lut_sub lut_8293 ({sk[1592], i_14_, i_13_, i_12_, i_15_, n_n191, n_n112}, x2152x);
	defparam lut_8293.LUT_SIZE = 7;
	defparam lut_8293.mask = 128'h00ff00ffffffffff0000001100000001;

	lut_sub lut_8297 ({sk[1593], n_n184, x719x, n_n108, n_n113, x1085x, x2152x}, n_n860);
	defparam lut_8297.LUT_SIZE = 7;
	defparam lut_8297.mask = 128'h00ff00ffffffffff5577557755775f7f;

	lut_sub lut_8301 ({sk[1594], i_14_, i_13_, i_12_, i_15_, n_n184}, x107x);
	defparam lut_8301.LUT_SIZE = 6;
	defparam lut_8301.mask = 64'h0055ffff00001014;

	lut_sub lut_8305 ({sk[1595], i_14_, i_13_, i_12_, i_15_, n_n184}, x1088x);
	defparam lut_8305.LUT_SIZE = 6;
	defparam lut_8305.mask = 64'h0055ffff00051114;

	lut_sub lut_8312 ({sk[1596], i_9_, i_10_, i_11_, i_15_, n_n123, n_n209}, x2147x);
	defparam lut_8312.LUT_SIZE = 7;
	defparam lut_8312.mask = 128'h00ff00ffffffffff0000010000010100;

	lut_sub lut_8316 ({sk[1597], x719x, n_n170, n_n113, x255x, x1088x, x2147x}, x19652x);
	defparam lut_8316.LUT_SIZE = 7;
	defparam lut_8316.mask = 128'h00ff00ffffffffff5577557755775f7f;

	lut_sub lut_8320 ({sk[1598], i_9_, i_10_, i_11_, x728x}, x416x);
	defparam lut_8320.LUT_SIZE = 5;
	defparam lut_8320.mask = 32'h57570140;

	lut_sub lut_8323 ({sk[1599], i_7_, i_8_, i_6_, x740x, x186x}, x4861x);
	defparam lut_8323.LUT_SIZE = 6;
	defparam lut_8323.mask = 64'h0055ffff00000100;

	lut_sub lut_8325 ({sk[1600], i_14_, i_13_, i_12_, i_15_, n_n216}, x212x);
	defparam lut_8325.LUT_SIZE = 6;
	defparam lut_8325.mask = 64'h0055ffff00000401;

	lut_sub lut_8328 ({sk[1601], i_7_, i_8_, i_6_, x740x, x212x}, x3501x);
	defparam lut_8328.LUT_SIZE = 6;
	defparam lut_8328.mask = 64'h0055ffff00001000;

	lut_sub lut_8330 ({sk[1602], i_15_, x714x, x17002x, n_n199, n_n204}, x3502x);
	defparam lut_8330.LUT_SIZE = 6;
	defparam lut_8330.mask = 64'h0055ffff00010000;

	lut_sub lut_8332 ({sk[1603], i_9_, i_10_, i_11_, x725x, x152x, x721x}, x1163x);
	defparam lut_8332.LUT_SIZE = 7;
	defparam lut_8332.mask = 128'h00ff00ffffffffff33333333333f7f33;

	lut_sub lut_8337 ({sk[1604], i_14_, i_13_, i_12_, i_15_, n_n149}, x1095x);
	defparam lut_8337.LUT_SIZE = 6;
	defparam lut_8337.mask = 64'h0055ffff01015154;

	lut_sub lut_8346 ({sk[1605], n_n101, n_n108, x86x, n_n190, x1724x, x1723x}, n_n4763);
	defparam lut_8346.LUT_SIZE = 7;
	defparam lut_8346.mask = 128'h00ff00ffffffffff00003f3f55ff7fff;

	lut_sub lut_8351 ({sk[1606], x734x, n_n126, n_n214, x1104x, x17506x, x18666x}, x18668x);
	defparam lut_8351.LUT_SIZE = 7;
	defparam lut_8351.mask = 128'h00ff00ffffffffff7777777777777fff;

	lut_sub lut_8356 ({sk[1607], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x1690x);
	defparam lut_8356.LUT_SIZE = 7;
	defparam lut_8356.mask = 128'h00ff00ffffffffff0303003337053770;

	lut_sub lut_8370 ({sk[1608], i_14_, i_13_, i_12_, i_15_, n_n191}, x1689x);
	defparam lut_8370.LUT_SIZE = 6;
	defparam lut_8370.mask = 64'h0055ffff15455054;

	lut_sub lut_8382 ({sk[1609], i_14_, i_13_, i_12_, i_15_, n_n170}, x208x);
	defparam lut_8382.LUT_SIZE = 6;
	defparam lut_8382.mask = 64'h0055ffff00001014;

	lut_sub lut_8386 ({sk[1610], i_14_, i_13_, i_12_, i_15_, n_n170}, x1859x);
	defparam lut_8386.LUT_SIZE = 6;
	defparam lut_8386.mask = 64'h0055ffff11054040;

	lut_sub lut_8393 ({sk[1611], i_14_, i_13_, i_12_, i_15_, n_n170}, x1860x);
	defparam lut_8393.LUT_SIZE = 6;
	defparam lut_8393.mask = 64'h0055ffff00015054;

	lut_sub lut_8400 ({sk[1612], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1099x);
	defparam lut_8400.LUT_SIZE = 7;
	defparam lut_8400.mask = 128'h00ff00ffffffffff7000070000700007;

	lut_sub lut_8409 ({sk[1613], i_14_, i_13_, i_12_, i_15_, n_n170}, x1098x);
	defparam lut_8409.LUT_SIZE = 6;
	defparam lut_8409.mask = 64'h0055ffff40100401;

	lut_sub lut_8414 ({sk[1614], i_9_, i_10_, i_8_, i_11_, n_n18, x285x}, x16991x);
	defparam lut_8414.LUT_SIZE = 7;
	defparam lut_8414.mask = 128'h00ff00ffffffffff0001000101000100;

	lut_sub lut_8419 ({sk[1615], n_n108, n_n125, n_n214, n_n57, x1098x, x16991x}, x16993x);
	defparam lut_8419.LUT_SIZE = 7;
	defparam lut_8419.mask = 128'h00ff00ffffffffff55557f7f55ff7fff;

	lut_sub lut_8424 ({sk[1616], i_8_, n_n16, x735x, n_n108, x1104x, x1099x}, x16994x);
	defparam lut_8424.LUT_SIZE = 7;
	defparam lut_8424.mask = 128'h00ff00ffffffffff0303035703030303;

	lut_sub lut_8427 ({sk[1617], n_n124, x734x, n_n126, x86x, n_n4903, x250x}, x16997x);
	defparam lut_8427.LUT_SIZE = 7;
	defparam lut_8427.mask = 128'h00ff00ffffffffff3333337733333f7f;

	lut_sub lut_8431 ({sk[1618], n_n124, x734x, n_n126, n_n169, x1019x, x1861x}, x16998x);
	defparam lut_8431.LUT_SIZE = 7;
	defparam lut_8431.mask = 128'h00ff00ffffffffff0000005500003f7f;

	lut_sub lut_8435 ({sk[1619], n_n101, n_n108, x544x, n_n176, x208x, x100x}, x16999x);
	defparam lut_8435.LUT_SIZE = 7;
	defparam lut_8435.mask = 128'h00ff00ffffffffff00ff5fff33ff7fff;

	lut_sub lut_8440 ({sk[1620], i_14_, i_13_, i_12_, i_15_, n_n177}, x1900x);
	defparam lut_8440.LUT_SIZE = 6;
	defparam lut_8440.mask = 64'h0055ffff11054040;

	lut_sub lut_8447 ({sk[1621], n_n177, x714x, x17002x, x720x, x100x, x1900x}, x17014x);
	defparam lut_8447.LUT_SIZE = 7;
	defparam lut_8447.mask = 128'h00ff00ffffffffff000000770000007f;

	lut_sub lut_8451 ({sk[1622], i_14_, i_13_, i_12_, i_15_, n_n170}, x1789x);
	defparam lut_8451.LUT_SIZE = 6;
	defparam lut_8451.mask = 64'h0055ffff11055154;

	lut_sub lut_8462 ({sk[1623], x740x, n_n200, x180x, x397x, x361x, x1789x}, x17015x);
	defparam lut_8462.LUT_SIZE = 7;
	defparam lut_8462.mask = 128'h00ff00ffffffffff3f3f3f3f3f3f7fff;

	lut_sub lut_8467 ({sk[1624], x4900x, n_n5060, x461x, x4906x, x4902x, x4903x}, x17018x);
	defparam lut_8467.LUT_SIZE = 7;
	defparam lut_8467.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_8474 ({sk[1625], i_8_, i_1_, i_2_, i_0_, x17002x, x141x}, n_n4604);
	defparam lut_8474.LUT_SIZE = 7;
	defparam lut_8474.mask = 128'h00ff00ffffffffff0000000010000000;

	lut_sub lut_8476 ({sk[1626], i_14_, i_13_, i_12_, i_15_, n_n199}, x1103x);
	defparam lut_8476.LUT_SIZE = 6;
	defparam lut_8476.mask = 64'h0055ffff40100401;

	lut_sub lut_8481 ({sk[1627], i_15_, x714x, x17002x, n_n199, n_n209, x728x}, x4909x);
	defparam lut_8481.LUT_SIZE = 7;
	defparam lut_8481.mask = 128'h00ff00ffffffffff0000000500000007;

	lut_sub lut_8484 ({sk[1628], n_n40, x4905x, n_n4604, x1103x, x1867x, x4909x}, x17019x);
	defparam lut_8484.LUT_SIZE = 7;
	defparam lut_8484.mask = 128'h00ff00ffffffffff55ffffff7fffffff;

	lut_sub lut_8490 ({sk[1629], i_7_, i_8_, i_6_, x740x, n_n177, x720x}, x4898x);
	defparam lut_8490.LUT_SIZE = 7;
	defparam lut_8490.mask = 128'h00ff00ffffffffff0000000001000000;

	lut_sub lut_8492 ({sk[1630], i_14_, i_13_, i_12_, i_15_, n_n170}, x1898x);
	defparam lut_8492.LUT_SIZE = 6;
	defparam lut_8492.mask = 64'h0055ffff00015054;

	lut_sub lut_8499 ({sk[1631], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1102x);
	defparam lut_8499.LUT_SIZE = 7;
	defparam lut_8499.mask = 128'h00ff00ffffffffff0050500333003330;

	lut_sub lut_8508 ({sk[1632], i_14_, i_13_, i_12_, i_15_, n_n170}, x225x);
	defparam lut_8508.LUT_SIZE = 6;
	defparam lut_8508.mask = 64'h0055ffff11040000;

	lut_sub lut_8512 ({sk[1633], n_n41, n_n169, x69x, n_n142, x4898x, x225x}, x17023x);
	defparam lut_8512.LUT_SIZE = 7;
	defparam lut_8512.mask = 128'h00ff00ffffffffff333333337fffffff;

	lut_sub lut_8518 ({sk[1634], n_n41, n_n40, x224x, x57x, x1898x, x1102x}, x17024x);
	defparam lut_8518.LUT_SIZE = 7;
	defparam lut_8518.mask = 128'h00ff00ffffffffff00005fff33337fff;

	lut_sub lut_8523 ({sk[1635], x17014x, x17015x, x17018x, x17019x, x17023x, x17024x}, n_n4404);
	defparam lut_8523.LUT_SIZE = 7;
	defparam lut_8523.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_8530 ({sk[1636], i_8_, x740x, n_n16, n_n177, x719x, x635x}, x17039x);
	defparam lut_8530.LUT_SIZE = 7;
	defparam lut_8530.mask = 128'h00ff00ffffffffff5555555755555557;

	lut_sub lut_8534 ({sk[1637], n_n38, n_n39, n_n134, n_n132, n_n84, x17039x}, x17041x);
	defparam lut_8534.LUT_SIZE = 7;
	defparam lut_8534.mask = 128'h00ff00ffffffffff55555f5f7fff7fff;

	lut_sub lut_8540 ({sk[1638], i_7_, i_8_, i_6_, x740x, x104x}, x503x);
	defparam lut_8540.LUT_SIZE = 6;
	defparam lut_8540.mask = 64'h0055ffff00010000;

	lut_sub lut_8542 ({sk[1639], n_n40, n_n5056, n_n57, x4885x, x4886x, x503x}, x17045x);
	defparam lut_8542.LUT_SIZE = 7;
	defparam lut_8542.mask = 128'h00ff00ffffffffff7f7fffff7fffffff;

	lut_sub lut_8548 ({sk[1640], i_7_, i_8_, i_6_, x740x, n_n4461, x279x}, x17046x);
	defparam lut_8548.LUT_SIZE = 7;
	defparam lut_8548.mask = 128'h00ff00ffffffffff3337333733333333;

	lut_sub lut_8552 ({sk[1641], n_n38, n_n39, n_n84, x104x, x1822x, x1881x}, x17047x);
	defparam lut_8552.LUT_SIZE = 7;
	defparam lut_8552.mask = 128'h00ff00ffffffffff000033ff5f5f7fff;

	lut_sub lut_8557 ({sk[1642], x597x, x620x, x17041x, x17045x, x17046x, x17047x}, n_n4403);
	defparam lut_8557.LUT_SIZE = 7;
	defparam lut_8557.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_8564 ({sk[1643], n_n46, n_n132, n_n47, x218x, x141x, x57x}, x21418x);
	defparam lut_8564.LUT_SIZE = 7;
	defparam lut_8564.mask = 128'h00ff00ffffffffffffccff00a080a000;

	lut_sub lut_8569 ({sk[1644], x714x, x17051x, x719x, n_n216, x4861x, x21418x}, x17055x);
	defparam lut_8569.LUT_SIZE = 7;
	defparam lut_8569.mask = 128'h00ff00ffffffffffbbbbbbbbbbbbbbbf;

	lut_sub lut_8573 ({sk[1645], i_8_, x740x, n_n18, n_n47, x1223x, x1222x}, n_n4195);
	defparam lut_8573.LUT_SIZE = 7;
	defparam lut_8573.mask = 128'h00ff00ffffffffff0505053705050505;

	lut_sub lut_8576 ({sk[1646], i_14_, i_13_, i_12_, i_15_, n_n177}, x1846x);
	defparam lut_8576.LUT_SIZE = 6;
	defparam lut_8576.mask = 64'h0055ffff40100401;

	lut_sub lut_8581 ({sk[1647], x740x, n_n161, n_n47, x209x, n_n4195, x1846x}, x17056x);
	defparam lut_8581.LUT_SIZE = 7;
	defparam lut_8581.mask = 128'h00ff00ffffffffff3377337733773f7f;

	lut_sub lut_8585 ({sk[1648], i_14_, i_13_, i_12_, i_15_, n_n46, n_n177}, x4840x);
	defparam lut_8585.LUT_SIZE = 7;
	defparam lut_8585.mask = 128'h00ff00ffffffffff0000010000100001;

	lut_sub lut_8589 ({sk[1649], x725x, x714x, x17051x, x721x, n_n170, x728x}, x4841x);
	defparam lut_8589.LUT_SIZE = 7;
	defparam lut_8589.mask = 128'h00ff00ffffffffff0000001300000033;

	lut_sub lut_8593 ({sk[1650], n_n6266, n_n6268, x602x, x611x, x4840x, x4841x}, x17060x);
	defparam lut_8593.LUT_SIZE = 7;
	defparam lut_8593.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_8600 ({sk[1651], x17008x, x17009x, x17055x, x17056x}, x17063x);
	defparam lut_8600.LUT_SIZE = 5;
	defparam lut_8600.mask = 32'h57577fff;

	lut_sub lut_8605 ({sk[1652], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1106x);
	defparam lut_8605.LUT_SIZE = 7;
	defparam lut_8605.mask = 128'h00ff00ffffffffff7000030000300003;

	lut_sub lut_8611 ({sk[1653], i_14_, i_13_, i_12_, i_15_, n_n149}, x1105x);
	defparam lut_8611.LUT_SIZE = 6;
	defparam lut_8611.mask = 64'h0055ffff40100401;

	lut_sub lut_8616 ({sk[1654], i_14_, i_13_, i_12_, i_15_, n_n199}, x258x);
	defparam lut_8616.LUT_SIZE = 6;
	defparam lut_8616.mask = 64'h0055ffff11040000;

	lut_sub lut_8620 ({sk[1655], i_9_, i_10_, i_11_, x714x, x17002x, x720x}, x4157x);
	defparam lut_8620.LUT_SIZE = 7;
	defparam lut_8620.mask = 128'h00ff00ffffffffff0000000000010000;

	lut_sub lut_8622 ({sk[1656], i_14_, i_13_, i_12_, i_15_, n_n216}, x1109x);
	defparam lut_8622.LUT_SIZE = 6;
	defparam lut_8622.mask = 64'h0055ffff11014044;

	lut_sub lut_8629 ({sk[1657], x181x, n_n46, n_n47, x143x, x74x, x68x}, x18413x);
	defparam lut_8629.LUT_SIZE = 7;
	defparam lut_8629.mask = 128'h00ff00ffffffffff000f777f00ff77ff;

	lut_sub lut_8634 ({sk[1658], n_n5319, n_n5118, n_n47, x47x, x154x, n_n5121}, x18414x);
	defparam lut_8634.LUT_SIZE = 7;
	defparam lut_8634.mask = 128'h00ff00ffffffffff557fffffffffffff;

	lut_sub lut_8640 ({sk[1659], i_14_, i_13_, i_12_, i_15_, n_n177}, x1111x);
	defparam lut_8640.LUT_SIZE = 6;
	defparam lut_8640.mask = 64'h0055ffff01015154;

	lut_sub lut_8649 ({sk[1660], i_14_, i_13_, i_12_, i_15_, n_n184}, x1274x);
	defparam lut_8649.LUT_SIZE = 6;
	defparam lut_8649.mask = 64'h0055ffff14045000;

	lut_sub lut_8655 ({sk[1661], i_14_, i_13_, i_12_, i_15_, n_n177}, x362x);
	defparam lut_8655.LUT_SIZE = 6;
	defparam lut_8655.mask = 64'h0055ffff00005000;

	lut_sub lut_8658 ({sk[1662], i_14_, i_13_, i_12_, i_15_, n_n191}, x1185x);
	defparam lut_8658.LUT_SIZE = 6;
	defparam lut_8658.mask = 64'h0055ffff14445000;

	lut_sub lut_8665 ({sk[1663], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1183x);
	defparam lut_8665.LUT_SIZE = 7;
	defparam lut_8665.mask = 128'h00ff00ffffffffff0550505077000000;

	lut_sub lut_8674 ({sk[1664], i_14_, i_13_, i_12_, i_15_, n_n199}, x1125x);
	defparam lut_8674.LUT_SIZE = 6;
	defparam lut_8674.mask = 64'h0055ffff14445000;

	lut_sub lut_8681 ({sk[1665], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1124x);
	defparam lut_8681.LUT_SIZE = 7;
	defparam lut_8681.mask = 128'h00ff00ffffffffff0770307077000000;

	lut_sub lut_8693 ({sk[1666], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1131x);
	defparam lut_8693.LUT_SIZE = 7;
	defparam lut_8693.mask = 128'h00ff00ffffffffff0707700300003300;

	lut_sub lut_8703 ({sk[1667], i_14_, i_13_, i_12_, i_15_, n_n191}, x319x);
	defparam lut_8703.LUT_SIZE = 6;
	defparam lut_8703.mask = 64'h0055ffff00010050;

	lut_sub lut_8707 ({sk[1668], i_14_, i_13_, i_12_, i_15_, n_n177}, x331x);
	defparam lut_8707.LUT_SIZE = 6;
	defparam lut_8707.mask = 64'h0055ffff00010050;

	lut_sub lut_8711 ({sk[1669], i_14_, i_13_, i_12_, i_15_, n_n177}, x312x);
	defparam lut_8711.LUT_SIZE = 6;
	defparam lut_8711.mask = 64'h0055ffff11400000;

	lut_sub lut_8715 ({sk[1670], n_n197, n_n212, x1131x, x319x, x331x, x312x}, n_n1839);
	defparam lut_8715.LUT_SIZE = 7;
	defparam lut_8715.mask = 128'h00ff00ffffffffff000077ff0fff7fff;

	lut_sub lut_8721 ({sk[1671], i_14_, i_13_, i_12_, i_15_, n_n170}, x18907x);
	defparam lut_8721.LUT_SIZE = 6;
	defparam lut_8721.mask = 64'h0055ffff11410050;

	lut_sub lut_8728 ({sk[1672], i_14_, i_13_, i_12_, i_15_, n_n149, n_n177}, x18908x);
	defparam lut_8728.LUT_SIZE = 7;
	defparam lut_8728.mask = 128'h00ff00ffffffffff0505500700007700;

	lut_sub lut_8738 ({sk[1673], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1132x);
	defparam lut_8738.LUT_SIZE = 7;
	defparam lut_8738.mask = 128'h00ff00ffffffffff0707700700007700;

	lut_sub lut_8751 ({sk[1674], x735x, n_n200, n_n212, x18907x, x18908x, x1132x}, n_n1838);
	defparam lut_8751.LUT_SIZE = 7;
	defparam lut_8751.mask = 128'h00ff00ffffffffff0055005500553f7f;

	lut_sub lut_8755 ({sk[1675], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1135x);
	defparam lut_8755.LUT_SIZE = 7;
	defparam lut_8755.mask = 128'h00ff00ffffffffff0707700700007700;

	lut_sub lut_8768 ({sk[1676], n_n197, n_n212, x319x, n_n1839, n_n1838, x1135x}, n_n1807);
	defparam lut_8768.LUT_SIZE = 7;
	defparam lut_8768.mask = 128'h00ff00ffffffffff3f3f7fff7f7f7fff;

	lut_sub lut_8774 ({sk[1677], i_8_, n_n16, x735x, x52x, x313x, n_n102}, x21452x);
	defparam lut_8774.LUT_SIZE = 7;
	defparam lut_8774.mask = 128'h00ff00ffffffffff0000007f00000000;

	lut_sub lut_8780 ({sk[1678], x729x, x735x, n_n126, n_n184, x383x, x21452x}, x18917x);
	defparam lut_8780.LUT_SIZE = 7;
	defparam lut_8780.mask = 128'h00ff00ffffffffff555555775555557f;

	lut_sub lut_8784 ({sk[1679], i_14_, i_13_, i_12_, i_15_, n_n191}, x1279x);
	defparam lut_8784.LUT_SIZE = 6;
	defparam lut_8784.mask = 64'h0055ffff00400050;

	lut_sub lut_8788 ({sk[1680], i_14_, i_13_, i_12_, i_15_, n_n184}, x1398x);
	defparam lut_8788.LUT_SIZE = 6;
	defparam lut_8788.mask = 64'h0055ffff11010050;

	lut_sub lut_8794 ({sk[1681], i_14_, i_13_, i_12_, i_15_, n_n184}, x1397x);
	defparam lut_8794.LUT_SIZE = 6;
	defparam lut_8794.mask = 64'h0055ffff11410000;

	lut_sub lut_8799 ({sk[1682], n_n123, n_n125, x52x, x1279x, x1398x, x1397x}, x18918x);
	defparam lut_8799.LUT_SIZE = 7;
	defparam lut_8799.mask = 128'h00ff00ffffffffff00003fff5f5f7fff;

	lut_sub lut_8805 ({sk[1683], i_14_, i_13_, i_12_, i_15_, n_n156}, x1468x);
	defparam lut_8805.LUT_SIZE = 6;
	defparam lut_8805.mask = 64'h0055ffff11410050;

	lut_sub lut_8812 ({sk[1684], n_n197, n_n212, n_n141, n_n139, n_n131, x1468x}, x18922x);
	defparam lut_8812.LUT_SIZE = 7;
	defparam lut_8812.mask = 128'h00ff00ffffffffff00003fff7f7f7fff;

	lut_sub lut_8819 ({sk[1685], i_9_, i_10_, i_11_, i_15_, n_n201}, x403x);
	defparam lut_8819.LUT_SIZE = 6;
	defparam lut_8819.mask = 64'h0055ffff10000100;

	lut_sub lut_8822 ({sk[1686], i_14_, i_13_, i_12_, i_15_, n_n149, n_n191}, x1283x);
	defparam lut_8822.LUT_SIZE = 7;
	defparam lut_8822.mask = 128'h00ff00ffffffffff0303350000000000;

	lut_sub lut_8827 ({sk[1687], i_9_, i_10_, i_11_, i_15_, n_n201}, x18921x);
	defparam lut_8827.LUT_SIZE = 6;
	defparam lut_8827.mask = 64'h0055ffff10000101;

	lut_sub lut_8831 ({sk[1688], i_14_, i_13_, i_12_, i_15_, n_n149}, x316x);
	defparam lut_8831.LUT_SIZE = 6;
	defparam lut_8831.mask = 64'h0055ffff00010050;

	lut_sub lut_8835 ({sk[1689], n_n197, n_n212, x403x, x1283x, x18921x, x316x}, x18923x);
	defparam lut_8835.LUT_SIZE = 7;
	defparam lut_8835.mask = 128'h00ff00ffffffffff00005fff3f3f7fff;

	lut_sub lut_8841 ({sk[1690], i_7_, i_8_, i_6_, x735x, n_n212, n_n129}, x2824x);
	defparam lut_8841.LUT_SIZE = 7;
	defparam lut_8841.mask = 128'h00ff00ffffffffff1111111115111111;

	lut_sub lut_8844 ({sk[1691], n_n125, x188x, n_n127, x143x, x364x, x2824x}, n_n1927);
	defparam lut_8844.LUT_SIZE = 7;
	defparam lut_8844.mask = 128'h00ff00ffffffffff555555ff7f7f7fff;

	lut_sub lut_8849 ({sk[1692], i_14_, i_13_, i_12_, i_15_, n_n199}, x136x);
	defparam lut_8849.LUT_SIZE = 6;
	defparam lut_8849.mask = 64'h0055ffff00000050;

	lut_sub lut_8852 ({sk[1693], n_n124, x735x, n_n126, x74x, n_n95, x136x}, x18926x);
	defparam lut_8852.LUT_SIZE = 7;
	defparam lut_8852.mask = 128'h00ff00ffffffffff0000007f0000777f;

	lut_sub lut_8858 ({sk[1694], n_n123, n_n125, x143x, x74x, n_n102, x364x}, x18927x);
	defparam lut_8858.LUT_SIZE = 7;
	defparam lut_8858.mask = 128'h00ff00ffffffffff000033335fff7fff;

	lut_sub lut_8863 ({sk[1695], n_n1927, x18926x, x18927x}, x18929x);
	defparam lut_8863.LUT_SIZE = 4;
	defparam lut_8863.mask = 16'h0f7f;

	lut_sub lut_8867 ({sk[1696], x18917x, x18918x, x18922x, x18923x}, x18930x);
	defparam lut_8867.LUT_SIZE = 5;
	defparam lut_8867.mask = 32'h57577fff;

	lut_sub lut_8872 ({sk[1697], i_9_, i_10_, i_11_, i_15_, n_n201}, x1242x);
	defparam lut_8872.LUT_SIZE = 6;
	defparam lut_8872.mask = 64'h0055ffff00011001;

	lut_sub lut_8876 ({sk[1698], i_9_, i_10_, i_11_, i_15_, x729x, n_n201}, x1241x);
	defparam lut_8876.LUT_SIZE = 7;
	defparam lut_8876.mask = 128'h00ff00ffffffffff0000000505003305;

	lut_sub lut_8881 ({sk[1699], n_n124, x735x, n_n126, n_n115, x1242x, x1241x}, x18935x);
	defparam lut_8881.LUT_SIZE = 7;
	defparam lut_8881.mask = 128'h00ff00ffffffffff0000003f00005f7f;

	lut_sub lut_8886 ({sk[1700], n_n112, x293x, n_n137, n_n109, x760x, x412x}, x21362x);
	defparam lut_8886.LUT_SIZE = 7;
	defparam lut_8886.mask = 128'h00ff00ffffffffffc8c8c8c8c8000000;

	lut_sub lut_8891 ({sk[1701], i_15_, n_n108, n_n216, n_n213, x613x, x21362x}, n_n1913);
	defparam lut_8891.LUT_SIZE = 7;
	defparam lut_8891.mask = 128'h00ff00ffffffffffbbbbbbbbbbbbbbbf;

	lut_sub lut_8895 ({sk[1702], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x18946x);
	defparam lut_8895.LUT_SIZE = 7;
	defparam lut_8895.mask = 128'h00ff00ffffffffff0000700000005500;

	lut_sub lut_8900 ({sk[1703], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1139x);
	defparam lut_8900.LUT_SIZE = 7;
	defparam lut_8900.mask = 128'h00ff00ffffffffff0505000500007700;

	lut_sub lut_8908 ({sk[1704], n_n123, n_n125, x832x, x831x, x147x, n_n77}, x18949x);
	defparam lut_8908.LUT_SIZE = 7;
	defparam lut_8908.mask = 128'h00ff00ffffffffff000033ff5f5f7fff;

	lut_sub lut_8913 ({sk[1705], n_n123, n_n125, x146x, x18946x, x1139x, x18949x}, x18950x);
	defparam lut_8913.LUT_SIZE = 7;
	defparam lut_8913.mask = 128'h00ff00ffffffffff55555fff77777fff;

	lut_sub lut_8918 ({sk[1706], x735x, n_n161, n_n113, x310x, x1192x, x305x}, n_n1914);
	defparam lut_8918.LUT_SIZE = 7;
	defparam lut_8918.mask = 128'h00ff00ffffffffff005f005f005f337f;

	lut_sub lut_8922 ({sk[1707], n_n123, n_n125, n_n122, n_n113, n_n131, x21361x}, x18942x);
	defparam lut_8922.LUT_SIZE = 7;
	defparam lut_8922.mask = 128'h00ff00ffffffffffaaafbbbfbbbfbbbf;

	lut_sub lut_8927 ({sk[1708], n_n1918, n_n1917, x18935x, n_n1913, n_n1914, x18942x}, x18951x);
	defparam lut_8927.LUT_SIZE = 7;
	defparam lut_8927.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_8934 ({sk[1709], i_14_, i_13_, i_12_, i_15_, n_n191}, x1142x);
	defparam lut_8934.LUT_SIZE = 6;
	defparam lut_8934.mask = 64'h0055ffff15414000;

	lut_sub lut_8941 ({sk[1710], i_14_, i_13_, i_12_, i_15_, n_n184}, x88x);
	defparam lut_8941.LUT_SIZE = 6;
	defparam lut_8941.mask = 64'h0055ffff00100400;

	lut_sub lut_8944 ({sk[1711], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1144x);
	defparam lut_8944.LUT_SIZE = 7;
	defparam lut_8944.mask = 128'h00ff00ffffffffff5700000057550000;

	lut_sub lut_8950 ({sk[1712], i_14_, i_13_, i_12_, i_15_, n_n184, n_n216}, x1146x);
	defparam lut_8950.LUT_SIZE = 7;
	defparam lut_8950.mask = 128'h00ff00ffffffffff0555500550077770;

	lut_sub lut_8965 ({sk[1713], i_14_, i_13_, i_12_, i_15_, n_n191, n_n199}, x1145x);
	defparam lut_8965.LUT_SIZE = 7;
	defparam lut_8965.mask = 128'h00ff00ffffffffff0773700300030300;

	lut_sub lut_8976 ({sk[1714], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1148x);
	defparam lut_8976.LUT_SIZE = 7;
	defparam lut_8976.mask = 128'h00ff00ffffffffff0373700370055550;

	lut_sub lut_8990 ({sk[1715], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x1147x);
	defparam lut_8990.LUT_SIZE = 7;
	defparam lut_8990.mask = 128'h00ff00ffffffffff0333300330073330;

	lut_sub lut_9002 ({sk[1716], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x1152x);
	defparam lut_9002.LUT_SIZE = 7;
	defparam lut_9002.mask = 128'h00ff00ffffffffff0737000550005550;

	lut_sub lut_9013 ({sk[1717], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1151x);
	defparam lut_9013.LUT_SIZE = 7;
	defparam lut_9013.mask = 128'h00ff00ffffffffff0303000330053570;

	lut_sub lut_9023 ({sk[1718], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1154x);
	defparam lut_9023.LUT_SIZE = 7;
	defparam lut_9023.mask = 128'h00ff00ffffffffff0505000770037370;

	lut_sub lut_9036 ({sk[1719], i_14_, i_13_, i_12_, i_15_, n_n184}, x1153x);
	defparam lut_9036.LUT_SIZE = 6;
	defparam lut_9036.mask = 64'h0055ffff15414154;

	lut_sub lut_9047 ({sk[1720], i_7_, i_8_, i_6_, x729x, x740x, n_n170}, x3518x);
	defparam lut_9047.LUT_SIZE = 7;
	defparam lut_9047.mask = 128'h00ff00ffffffffff0000000001000000;

	lut_sub lut_9049 ({sk[1721], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1156x);
	defparam lut_9049.LUT_SIZE = 7;
	defparam lut_9049.mask = 128'h00ff00ffffffffff0777300770007330;

	lut_sub lut_9065 ({sk[1722], i_14_, i_13_, i_12_, i_15_, n_n170}, x1155x);
	defparam lut_9065.LUT_SIZE = 6;
	defparam lut_9065.mask = 64'h0055ffff11014044;

	lut_sub lut_9072 ({sk[1723], n_n184, n_n42, n_n43, n_n191, x721x, x728x}, n_n1566);
	defparam lut_9072.LUT_SIZE = 7;
	defparam lut_9072.mask = 128'h00ff00ffffffffff0000070700330737;

	lut_sub lut_9076 ({sk[1724], i_14_, i_13_, i_12_, i_15_, n_n41, n_n216}, x21457x);
	defparam lut_9076.LUT_SIZE = 7;
	defparam lut_9076.mask = 128'h00ff00fffffffffffefefffeefffefef;

	lut_sub lut_9085 ({sk[1725], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1296x);
	defparam lut_9085.LUT_SIZE = 7;
	defparam lut_9085.mask = 128'h00ff00ffffffffff0000000000070750;

	lut_sub lut_9091 ({sk[1726], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1297x);
	defparam lut_9091.LUT_SIZE = 7;
	defparam lut_9091.mask = 128'h00ff00ffffffffff0777300330003330;

	lut_sub lut_9104 ({sk[1727], i_9_, i_10_, i_11_, n_n41, n_n40, x719x}, x19543x);
	defparam lut_9104.LUT_SIZE = 7;
	defparam lut_9104.mask = 128'h00ff00ffffffffff0015150000111100;

	lut_sub lut_9111 ({sk[1728], i_14_, i_13_, i_12_, i_15_, n_n156}, x1161x);
	defparam lut_9111.LUT_SIZE = 6;
	defparam lut_9111.mask = 64'h0055ffff00001154;

	lut_sub lut_9117 ({sk[1729], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1724x);
	defparam lut_9117.LUT_SIZE = 7;
	defparam lut_9117.mask = 128'h00ff00ffffffffff0555505555035550;

	lut_sub lut_9130 ({sk[1730], i_14_, i_13_, i_12_, i_15_, n_n184}, x1723x);
	defparam lut_9130.LUT_SIZE = 6;
	defparam lut_9130.mask = 64'h0055ffff15455154;

	lut_sub lut_9143 ({sk[1731], i_14_, i_13_, i_12_, i_15_, n_n177, n_n216}, x1165x);
	defparam lut_9143.LUT_SIZE = 7;
	defparam lut_9143.mask = 128'h00ff00ffffffffff7000070000700003;

	lut_sub lut_9151 ({sk[1732], n_n124, x734x, x218x, x141x, x224x, x209x}, x17070x);
	defparam lut_9151.LUT_SIZE = 7;
	defparam lut_9151.mask = 128'h00ff00ffffffffff0000000000007fff;

	lut_sub lut_9156 ({sk[1733], n_n108, n_n142, x4838x, x617x, x1165x, x1863x}, x17071x);
	defparam lut_9156.LUT_SIZE = 7;
	defparam lut_9156.mask = 128'h00ff00ffffffffff0fff0fff7fffffff;

	lut_sub lut_9162 ({sk[1734], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1168x);
	defparam lut_9162.LUT_SIZE = 7;
	defparam lut_9162.mask = 128'h00ff00ffffffffff7000070000300003;

	lut_sub lut_9169 ({sk[1735], i_7_, i_8_, i_6_, x740x, x720x, n_n170}, x4817x);
	defparam lut_9169.LUT_SIZE = 7;
	defparam lut_9169.mask = 128'h00ff00ffffffffff0000000000010000;

	lut_sub lut_9171 ({sk[1736], i_14_, i_13_, i_12_, i_15_, n_n177}, x1170x);
	defparam lut_9171.LUT_SIZE = 6;
	defparam lut_9171.mask = 64'h0055ffff11055154;

	lut_sub lut_9182 ({sk[1737], i_14_, i_13_, i_12_, i_15_, n_n170}, x148x);
	defparam lut_9182.LUT_SIZE = 6;
	defparam lut_9182.mask = 64'h0055ffff00014040;

	lut_sub lut_9186 ({sk[1738], i_14_, i_13_, i_12_, i_15_, n_n170, n_n216}, x1169x);
	defparam lut_9186.LUT_SIZE = 7;
	defparam lut_9186.mask = 128'h00ff00ffffffffff0050500333003330;

	lut_sub lut_9195 ({sk[1739], i_7_, i_8_, i_6_, x735x, x141x}, n_n4658);
	defparam lut_9195.LUT_SIZE = 6;
	defparam lut_9195.mask = 64'h0055ffff00010000;

	lut_sub lut_9197 ({sk[1740], i_14_, i_13_, i_12_, i_15_, n_n156}, x1819x);
	defparam lut_9197.LUT_SIZE = 6;
	defparam lut_9197.mask = 64'h0055ffff00001114;

	lut_sub lut_9202 ({sk[1741], i_14_, i_13_, i_12_, i_15_, n_n156}, x1824x);
	defparam lut_9202.LUT_SIZE = 6;
	defparam lut_9202.mask = 64'h0055ffff11054040;

	lut_sub lut_9209 ({sk[1742], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1175x);
	defparam lut_9209.LUT_SIZE = 7;
	defparam lut_9209.mask = 128'h00ff00ffffffffff0775307555005050;

	lut_sub lut_9223 ({sk[1743], i_14_, i_13_, i_12_, i_15_, n_n184}, x1174x);
	defparam lut_9223.LUT_SIZE = 6;
	defparam lut_9223.mask = 64'h0055ffff15055154;

	lut_sub lut_9235 ({sk[1744], i_14_, i_13_, i_12_, i_15_, n_n191}, x318x);
	defparam lut_9235.LUT_SIZE = 6;
	defparam lut_9235.mask = 64'h0055ffff01010040;

	lut_sub lut_9239 ({sk[1745], i_14_, i_13_, i_12_, i_15_, n_n191}, x1192x);
	defparam lut_9239.LUT_SIZE = 6;
	defparam lut_9239.mask = 64'h0055ffff01010050;

	lut_sub lut_9244 ({sk[1746], i_14_, i_13_, i_12_, i_15_, n_n184}, x305x);
	defparam lut_9244.LUT_SIZE = 6;
	defparam lut_9244.mask = 64'h0055ffff10400000;

	lut_sub lut_9247 ({sk[1747], i_14_, i_13_, i_12_, i_15_, n_n177}, x1194x);
	defparam lut_9247.LUT_SIZE = 6;
	defparam lut_9247.mask = 64'h0055ffff11410050;

	lut_sub lut_9254 ({sk[1748], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1193x);
	defparam lut_9254.LUT_SIZE = 7;
	defparam lut_9254.mask = 128'h00ff00ffffffffff0500500000000300;

	lut_sub lut_9258 ({sk[1749], i_9_, i_10_, i_11_, n_n31, n_n30, x721x}, n_n1843);
	defparam lut_9258.LUT_SIZE = 7;
	defparam lut_9258.mask = 128'h00ff00ffffffffff0515150011150500;

	lut_sub lut_9268 ({sk[1750], i_9_, i_10_, i_11_, x729x, x717x, x730x}, x1198x);
	defparam lut_9268.LUT_SIZE = 7;
	defparam lut_9268.mask = 128'h00ff00ffffffffff00000f007f007f00;

	lut_sub lut_9276 ({sk[1751], i_9_, i_10_, i_11_, i_15_, n_n201}, x1470x);
	defparam lut_9276.LUT_SIZE = 6;
	defparam lut_9276.mask = 64'h0055ffff01001100;

	lut_sub lut_9280 ({sk[1752], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x18959x);
	defparam lut_9280.LUT_SIZE = 7;
	defparam lut_9280.mask = 128'h00ff00ffffffffff0700700000000000;

	lut_sub lut_9285 ({sk[1753], i_14_, i_13_, i_12_, i_15_, n_n156, n_n216}, x18960x);
	defparam lut_9285.LUT_SIZE = 7;
	defparam lut_9285.mask = 128'h00ff00ffffffffff0003050300003300;

	lut_sub lut_9291 ({sk[1754], i_9_, i_10_, i_11_, n_n101, n_n108, x721x}, x21360x);
	defparam lut_9291.LUT_SIZE = 7;
	defparam lut_9291.mask = 128'h00ff00ffffffffffeaeeffffeeeeeeff;

	lut_sub lut_9299 ({sk[1755], n_n124, x734x, x1470x, x18959x, x18960x, x21360x}, x18962x);
	defparam lut_9299.LUT_SIZE = 7;
	defparam lut_9299.mask = 128'h00ff00ffffffffffaaaaaaaaaaaabfff;

	lut_sub lut_9304 ({sk[1756], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1200x);
	defparam lut_9304.LUT_SIZE = 7;
	defparam lut_9304.mask = 128'h00ff00ffffffffff0707700700007700;

	lut_sub lut_9317 ({sk[1757], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1401x);
	defparam lut_9317.LUT_SIZE = 7;
	defparam lut_9317.mask = 128'h00ff00ffffffffff0707700700007700;

	lut_sub lut_9330 ({sk[1758], i_8_, n_n149, n_n156, x734x, n_n16, x721x}, x18965x);
	defparam lut_9330.LUT_SIZE = 7;
	defparam lut_9330.mask = 128'h00ff00ffffffffff0001010100000101;

	lut_sub lut_9334 ({sk[1759], n_n46, n_n47, x1200x, x331x, x1401x, x18965x}, x18967x);
	defparam lut_9334.LUT_SIZE = 7;
	defparam lut_9334.mask = 128'h00ff00ffffffffff55557fff77ff7fff;

	lut_sub lut_9341 ({sk[1760], i_14_, i_13_, i_12_, i_15_, n_n149, n_n216}, x1471x);
	defparam lut_9341.LUT_SIZE = 7;
	defparam lut_9341.mask = 128'h00ff00ffffffffff0303350300003300;

	lut_sub lut_9349 ({sk[1761], n_n101, n_n108, n_n139, x18962x, x18967x, x1471x}, n_n1803);
	defparam lut_9349.LUT_SIZE = 7;
	defparam lut_9349.mask = 128'h00ff00ffffffffff3f3f7fff3fff7fff;

	lut_sub lut_9355 ({sk[1762], n_n42, n_n43, x52x, x139x, x257x, x313x}, x18975x);
	defparam lut_9355.LUT_SIZE = 7;
	defparam lut_9355.mask = 128'h00ff00ffffffffff000033ff5f5f7fff;

	lut_sub lut_9360 ({sk[1763], i_14_, i_13_, i_12_, i_15_, n_n156}, x303x);
	defparam lut_9360.LUT_SIZE = 6;
	defparam lut_9360.mask = 64'h0055ffff11400000;

	lut_sub lut_9364 ({sk[1764], i_14_, i_13_, i_12_, i_15_, n_n149, n_n191}, x1768x);
	defparam lut_9364.LUT_SIZE = 7;
	defparam lut_9364.mask = 128'h00ff00ffffffffff0303350300003300;

	lut_sub lut_9372 ({sk[1765], x740x, n_n161, x321x, x303x, x1768x, x410x}, x2755x);
	defparam lut_9372.LUT_SIZE = 7;
	defparam lut_9372.mask = 128'h00ff00ffffffffff0000000000007fff;

	lut_sub lut_9377 ({sk[1766], i_15_, x740x, n_n161, n_n47, n_n199, n_n201}, x2756x);
	defparam lut_9377.LUT_SIZE = 7;
	defparam lut_9377.mask = 128'h00ff00ffffffffff0000000001010111;

	lut_sub lut_9380 ({sk[1767], x714x, x17051x, n_n141, x403x, x1768x, x2756x}, x18981x);
	defparam lut_9380.LUT_SIZE = 7;
	defparam lut_9380.mask = 128'h00ff00ffffffffff5555555555557fff;

	lut_sub lut_9385 ({sk[1768], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1203x);
	defparam lut_9385.LUT_SIZE = 7;
	defparam lut_9385.mask = 128'h00ff00ffffffffff0707700500005500;

	lut_sub lut_9395 ({sk[1769], x729x, n_n43, n_n47, n_n191, n_n129, x18971x}, x18974x);
	defparam lut_9395.LUT_SIZE = 7;
	defparam lut_9395.mask = 128'h00ff00ffffffffff5577557755775f7f;

	lut_sub lut_9399 ({sk[1770], n_n46, n_n47, x1203x, x331x, x321x, x303x}, x18984x);
	defparam lut_9399.LUT_SIZE = 7;
	defparam lut_9399.mask = 128'h00ff00ffffffffff000077ff0fff7fff;

	lut_sub lut_9405 ({sk[1771], n_n1886, x18975x, x2755x, x18981x, x18974x, x18984x}, n_n1802);
	defparam lut_9405.LUT_SIZE = 7;
	defparam lut_9405.mask = 128'h00ff00ffffffffff7fffffffffffffff;

	lut_sub lut_9412 ({sk[1772], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1498x);
	defparam lut_9412.LUT_SIZE = 7;
	defparam lut_9412.mask = 128'h00ff00ffffffffff0307300700007500;

	lut_sub lut_9422 ({sk[1773], i_14_, i_13_, i_12_, i_15_, n_n149, n_n170}, x1497x);
	defparam lut_9422.LUT_SIZE = 7;
	defparam lut_9422.mask = 128'h00ff00ffffffffff0507500700007300;

	lut_sub lut_9432 ({sk[1774], n_n101, n_n108, x1194x, x1193x, x1498x, x1497x}, n_n1829);
	defparam lut_9432.LUT_SIZE = 7;
	defparam lut_9432.mask = 128'h00ff00ffffffffff00003f3f55ff7fff;

	lut_sub lut_9437 ({sk[1775], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x1533x);
	defparam lut_9437.LUT_SIZE = 7;
	defparam lut_9437.mask = 128'h00ff00ffffffffff0707700700007500;

	lut_sub lut_9449 ({sk[1776], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1532x);
	defparam lut_9449.LUT_SIZE = 7;
	defparam lut_9449.mask = 128'h00ff00ffffffffff0303300300003700;

	lut_sub lut_9457 ({sk[1777], n_n101, n_n108, x906x, x905x, x1533x, x1532x}, n_n1830);
	defparam lut_9457.LUT_SIZE = 7;
	defparam lut_9457.mask = 128'h00ff00ffffffffff00003f3f55ff7fff;

	lut_sub lut_9462 ({sk[1778], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1205x);
	defparam lut_9462.LUT_SIZE = 7;
	defparam lut_9462.mask = 128'h00ff00ffffffffff0707700700007300;

	lut_sub lut_9474 ({sk[1779], i_14_, i_13_, i_12_, i_15_, n_n191}, x1552x);
	defparam lut_9474.LUT_SIZE = 6;
	defparam lut_9474.mask = 64'h0055ffff01010050;

	lut_sub lut_9479 ({sk[1780], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x21359x);
	defparam lut_9479.LUT_SIZE = 7;
	defparam lut_9479.mask = 128'h00ff00fffffffffff8f88ff8ffff88ff;

	lut_sub lut_9492 ({sk[1781], n_n124, x734x, n_n126, x1205x, x1552x, x21359x}, x19004x);
	defparam lut_9492.LUT_SIZE = 7;
	defparam lut_9492.mask = 128'h00ff00ffffffffff0000003f0000aabf;

	lut_sub lut_9496 ({sk[1782], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1208x);
	defparam lut_9496.LUT_SIZE = 7;
	defparam lut_9496.mask = 128'h00ff00ffffffffff0057000000035700;

	lut_sub lut_9502 ({sk[1783], i_14_, i_13_, i_12_, i_15_, n_n216}, x1344x);
	defparam lut_9502.LUT_SIZE = 6;
	defparam lut_9502.mask = 64'h0055ffff15414000;

	lut_sub lut_9509 ({sk[1784], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1408x);
	defparam lut_9509.LUT_SIZE = 7;
	defparam lut_9509.mask = 128'h00ff00ffffffffff5500005757000057;

	lut_sub lut_9517 ({sk[1785], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1406x);
	defparam lut_9517.LUT_SIZE = 7;
	defparam lut_9517.mask = 128'h00ff00ffffffffff0357000000570000;

	lut_sub lut_9523 ({sk[1786], i_14_, i_13_, i_12_, i_15_, n_n156, n_n184}, x19314x);
	defparam lut_9523.LUT_SIZE = 7;
	defparam lut_9523.mask = 128'h00ff00ffffffffff0303050300500000;

	lut_sub lut_9529 ({sk[1787], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x21351x);
	defparam lut_9529.LUT_SIZE = 7;
	defparam lut_9529.mask = 128'h00ff00ffffffffffffa8ffa8a8ffffa8;

	lut_sub lut_9535 ({sk[1788], i_14_, i_13_, i_12_, i_15_, n_n216}, x1214x);
	defparam lut_9535.LUT_SIZE = 6;
	defparam lut_9535.mask = 64'h0055ffff15414054;

	lut_sub lut_9545 ({sk[1789], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x1506x);
	defparam lut_9545.LUT_SIZE = 7;
	defparam lut_9545.mask = 128'h00ff00ffffffffff0735300550005050;

	lut_sub lut_9555 ({sk[1790], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1509x);
	defparam lut_9555.LUT_SIZE = 7;
	defparam lut_9555.mask = 128'h00ff00ffffffffff0557000770077770;

	lut_sub lut_9572 ({sk[1791], i_14_, i_13_, i_12_, i_15_, n_n184}, x1508x);
	defparam lut_9572.LUT_SIZE = 6;
	defparam lut_9572.mask = 64'h0055ffff15414044;

	lut_sub lut_9581 ({sk[1792], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1216x);
	defparam lut_9581.LUT_SIZE = 7;
	defparam lut_9581.mask = 128'h00ff00ffffffffff0555000550075550;

	lut_sub lut_9592 ({sk[1793], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1215x);
	defparam lut_9592.LUT_SIZE = 7;
	defparam lut_9592.mask = 128'h00ff00ffffffffff0575700550000000;

	lut_sub lut_9601 ({sk[1794], i_14_, i_13_, i_12_, i_15_, n_n199}, x385x);
	defparam lut_9601.LUT_SIZE = 6;
	defparam lut_9601.mask = 64'h0055ffff05000000;

	lut_sub lut_9604 ({sk[1795], i_14_, i_13_, i_12_, i_15_, n_n34, n_n216}, x2084x);
	defparam lut_9604.LUT_SIZE = 7;
	defparam lut_9604.mask = 128'h00ff00ffffffffff0011000000010000;

	lut_sub lut_9608 ({sk[1796], n_n36, n_n34, n_n191, x720x, x154x, x385x}, x19712x);
	defparam lut_9608.LUT_SIZE = 7;
	defparam lut_9608.mask = 128'h00ff00ffffffffff00003333555f777f;

	lut_sub lut_9612 ({sk[1797], i_14_, i_13_, i_12_, i_15_, n_n216}, x335x);
	defparam lut_9612.LUT_SIZE = 6;
	defparam lut_9612.mask = 64'h0055ffff00000104;

	lut_sub lut_9615 ({sk[1798], i_14_, i_13_, i_12_, i_15_, n_n191}, x278x);
	defparam lut_9615.LUT_SIZE = 6;
	defparam lut_9615.mask = 64'h0055ffff05004000;

	lut_sub lut_9619 ({sk[1799], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1219x);
	defparam lut_9619.LUT_SIZE = 7;
	defparam lut_9619.mask = 128'h00ff00ffffffffff0033000030700000;

	lut_sub lut_9625 ({sk[1800], i_14_, i_13_, i_12_, i_15_, n_n31, n_n216}, x1911x);
	defparam lut_9625.LUT_SIZE = 7;
	defparam lut_9625.mask = 128'h00ff00ffffffffff0000000000010010;

	lut_sub lut_9628 ({sk[1801], x172x, n_n47, n_n191, x719x, x4100x, x1324x}, x18393x);
	defparam lut_9628.LUT_SIZE = 7;
	defparam lut_9628.mask = 128'h00ff00ffffffffff3333777f3333ffff;

	lut_sub lut_9633 ({sk[1802], n_n132, n_n47, x150x, x4861x, x4840x, x1379x}, x18397x);
	defparam lut_9633.LUT_SIZE = 7;
	defparam lut_9633.mask = 128'h00ff00ffffffffff3f3f7fff3f3fffff;

	lut_sub lut_9639 ({sk[1803], n_n46, n_n47, x209x, x217x, x18395x, x1846x}, x18398x);
	defparam lut_9639.LUT_SIZE = 7;
	defparam lut_9639.mask = 128'h00ff00ffffffffff000055553fff7fff;

	lut_sub lut_9644 ({sk[1804], x729x, n_n149, n_n46, n_n47, x118x, x1328x}, x18401x);
	defparam lut_9644.LUT_SIZE = 7;
	defparam lut_9644.mask = 128'h00ff00ffffffffff0707070707070fff;

	lut_sub lut_9649 ({sk[1805], n_n46, x247x, x116x, x1327x, x198x, x18389x}, x21367x);
	defparam lut_9649.LUT_SIZE = 7;
	defparam lut_9649.mask = 128'h00ff00ffffffffffffffffff80000000;

	lut_sub lut_9652 ({sk[1806], n_n46, n_n5319, n_n47, x151x, x1330x, x1329x}, x18420x);
	defparam lut_9652.LUT_SIZE = 7;
	defparam lut_9652.mask = 128'h00ff00ffffffffff003fffff557fffff;

	lut_sub lut_9657 ({sk[1807], i_14_, i_13_, i_12_, i_15_, n_n156}, x1576x);
	defparam lut_9657.LUT_SIZE = 6;
	defparam lut_9657.mask = 64'h0055ffff15455154;

	lut_sub lut_9670 ({sk[1808], i_14_, i_13_, i_12_, i_15_, n_n149, n_n177}, x1575x);
	defparam lut_9670.LUT_SIZE = 7;
	defparam lut_9670.mask = 128'h00ff00ffffffffff0555505555035350;

	lut_sub lut_9683 ({sk[1809], n_n46, n_n47, n_n77, x104x, x1576x, x1575x}, n_n3192);
	defparam lut_9683.LUT_SIZE = 7;
	defparam lut_9683.mask = 128'h00ff00ffffffffff000033ff5f5f7fff;

	lut_sub lut_9688 ({sk[1810], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1221x);
	defparam lut_9688.LUT_SIZE = 7;
	defparam lut_9688.mask = 128'h00ff00ffffffffff0775307555005050;

	lut_sub lut_9702 ({sk[1811], i_14_, i_13_, i_12_, i_15_, n_n170}, x1220x);
	defparam lut_9702.LUT_SIZE = 6;
	defparam lut_9702.mask = 64'h0055ffff00001154;

	lut_sub lut_9708 ({sk[1812], n_n46, n_n47, n_n82, n_n169, x812x, x1220x}, x18433x);
	defparam lut_9708.LUT_SIZE = 7;
	defparam lut_9708.mask = 128'h00ff00ffffffffff00000fff77777fff;

	lut_sub lut_9713 ({sk[1813], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1223x);
	defparam lut_9713.LUT_SIZE = 7;
	defparam lut_9713.mask = 128'h00ff00ffffffffff7000050000500005;

	lut_sub lut_9719 ({sk[1814], i_14_, i_13_, i_12_, i_15_, n_n199}, x1222x);
	defparam lut_9719.LUT_SIZE = 6;
	defparam lut_9719.mask = 64'h0055ffff40100401;

	lut_sub lut_9724 ({sk[1815], i_14_, i_13_, i_12_, i_15_, n_n184, n_n216}, x1228x);
	defparam lut_9724.LUT_SIZE = 7;
	defparam lut_9724.mask = 128'h00ff00ffffffffff7000030000300003;

	lut_sub lut_9730 ({sk[1816], i_14_, i_13_, i_12_, i_15_, n_n191}, x160x);
	defparam lut_9730.LUT_SIZE = 6;
	defparam lut_9730.mask = 64'h0055ffff40100000;

	lut_sub lut_9733 ({sk[1817], i_14_, i_13_, i_12_, i_15_, n_n191}, x1227x);
	defparam lut_9733.LUT_SIZE = 6;
	defparam lut_9733.mask = 64'h0055ffff40100401;

	lut_sub lut_9738 ({sk[1818], i_7_, i_5_, i_6_, i_3_, i_4_, n_n219}, x18707x);
	defparam lut_9738.LUT_SIZE = 7;
	defparam lut_9738.mask = 128'h00ff00ffffffffff0010001000100010;

	lut_sub lut_9743 ({sk[1819], n_n219, n_n14, n_n92, n_n18, n_n111, n_n12}, x21406x);
	defparam lut_9743.LUT_SIZE = 7;
	defparam lut_9743.mask = 128'h00ff00ffffffffffffaaff00fca8fc00;

	lut_sub lut_9750 ({sk[1820], n_n149, n_n7258, n_n14, x730x, x18707x, x21406x}, n_n3054);
	defparam lut_9750.LUT_SIZE = 7;
	defparam lut_9750.mask = 128'h00ff00ffffffffffbbbbffffbbbfffff;

	lut_sub lut_9755 ({sk[1821], i_14_, i_13_, i_12_, i_15_, n_n177}, x1230x);
	defparam lut_9755.LUT_SIZE = 6;
	defparam lut_9755.mask = 64'h0055ffff11014044;

	lut_sub lut_9762 ({sk[1822], i_14_, i_13_, i_12_, i_15_, n_n156}, x1234x);
	defparam lut_9762.LUT_SIZE = 6;
	defparam lut_9762.mask = 64'h5757ffff14045000;

	lut_sub lut_9768 ({sk[1823], i_14_, i_13_, i_12_, i_15_, n_n177}, x120x);
	defparam lut_9768.LUT_SIZE = 6;
	defparam lut_9768.mask = 64'h3f3f3fff14040000;

	lut_sub lut_9772 ({sk[1824], i_9_, i_10_, i_11_}, x412x);
	defparam lut_9772.LUT_SIZE = 4;
	defparam lut_9772.mask = 16'h5560;

	lut_sub lut_9775 ({sk[1825], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1246x);
	defparam lut_9775.LUT_SIZE = 7;
	defparam lut_9775.mask = 128'h3fff3fff3fff3fff0707700700007700;

	lut_sub lut_9788 ({sk[1826], x729x, n_n31, n_n30, n_n216, x56x, x1246x}, n_n1811);
	defparam lut_9788.LUT_SIZE = 7;
	defparam lut_9788.mask = 128'h3fff3fff3fff3fff00775577007f557f;

	lut_sub lut_9793 ({sk[1827], i_14_, i_13_, i_12_, i_15_, n_n149, n_n170}, x1399x);
	defparam lut_9793.LUT_SIZE = 7;
	defparam lut_9793.mask = 128'h3fff3fff3fff3fff0703700300003300;

	lut_sub lut_9802 ({sk[1828], i_8_, x734x, n_n17, n_n32, n_n122, x1399x}, n_n1857);
	defparam lut_9802.LUT_SIZE = 7;
	defparam lut_9802.mask = 128'h3fff3fff3fff3fff0303035703030303;

	lut_sub lut_9805 ({sk[1829], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x18825x);
	defparam lut_9805.LUT_SIZE = 7;
	defparam lut_9805.mask = 128'h3fff3fff3fff3fff0005000500005700;

	lut_sub lut_9811 ({sk[1830], i_14_, i_13_, i_12_, i_15_, n_n184}, x1248x);
	defparam lut_9811.LUT_SIZE = 6;
	defparam lut_9811.mask = 64'h1f5f1f5f11410040;

	lut_sub lut_9817 ({sk[1831], i_9_, i_10_, i_11_, i_15_, n_n201}, x1247x);
	defparam lut_9817.LUT_SIZE = 6;
	defparam lut_9817.mask = 64'h1f5f1f5f00100010;

	lut_sub lut_9820 ({sk[1832], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1252x);
	defparam lut_9820.LUT_SIZE = 7;
	defparam lut_9820.mask = 128'h3fff3fff3fff3fff0057000000035700;

	lut_sub lut_9826 ({sk[1833], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1256x);
	defparam lut_9826.LUT_SIZE = 7;
	defparam lut_9826.mask = 128'h3fff3fff3fff3fff0057550000005700;

	lut_sub lut_9832 ({sk[1834], i_14_, i_13_, i_12_, i_15_, n_n170}, x1822x);
	defparam lut_9832.LUT_SIZE = 6;
	defparam lut_9832.mask = 64'h1f5f1f5f00051004;

	lut_sub lut_9837 ({sk[1835], n_n38, n_n39, x53x, n_n78, x104x, x1822x}, n_n817);
	defparam lut_9837.LUT_SIZE = 7;
	defparam lut_9837.mask = 128'h3fff3fff3fff3fff000055ff3f3f7fff;

	lut_sub lut_9842 ({sk[1836], i_14_, i_13_, i_12_, i_15_, n_n191}, x167x);
	defparam lut_9842.LUT_SIZE = 6;
	defparam lut_9842.mask = 64'h1f5f1f5f00050004;

	lut_sub lut_9846 ({sk[1837], i_9_, i_10_, i_11_, i_15_, n_n33, n_n209}, x19480x);
	defparam lut_9846.LUT_SIZE = 7;
	defparam lut_9846.mask = 128'h3fff3fff3fff3fff0000010001000000;

	lut_sub lut_9849 ({sk[1838], i_8_, n_n31, x734x, n_n17, x111x, x167x}, x21346x);
	defparam lut_9849.LUT_SIZE = 7;
	defparam lut_9849.mask = 128'h3fff3fff3fff3ffffffaccc8ffffcccc;

	lut_sub lut_9858 ({sk[1839], i_14_, i_13_, i_12_, i_15_, n_n191}, x1259x);
	defparam lut_9858.LUT_SIZE = 6;
	defparam lut_9858.mask = 64'h1f5f1f5f00051114;

	lut_sub lut_9865 ({sk[1840], i_14_, i_13_, i_12_, i_15_, n_n184, n_n216}, x1258x);
	defparam lut_9865.LUT_SIZE = 7;
	defparam lut_9865.mask = 128'h0fff0fff7fff7fff0000005000030300;

	lut_sub lut_9869 ({sk[1841], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1261x);
	defparam lut_9869.LUT_SIZE = 7;
	defparam lut_9869.mask = 128'h0fff0fff7fff7fff0000007707050570;

	lut_sub lut_9880 ({sk[1842], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x1260x);
	defparam lut_9880.LUT_SIZE = 7;
	defparam lut_9880.mask = 128'h0fff0fff7fff7fff0000003303070730;

	lut_sub lut_9889 ({sk[1843], n_n123, n_n125, x1259x, x1258x, x1261x, x1260x}, n_n781);
	defparam lut_9889.LUT_SIZE = 7;
	defparam lut_9889.mask = 128'h0fff0fff7fff7fff000055ff3f3f7fff;

	lut_sub lut_9894 ({sk[1844], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1265x);
	defparam lut_9894.LUT_SIZE = 7;
	defparam lut_9894.mask = 128'h0fff0fff7fff7fff3000030000300007;

	lut_sub lut_9900 ({sk[1845], i_14_, i_13_, i_12_, i_15_, n_n149}, x1264x);
	defparam lut_9900.LUT_SIZE = 6;
	defparam lut_9900.mask = 64'h7777777740100401;

	lut_sub lut_9905 ({sk[1846], i_14_, i_13_, i_12_, i_15_, n_n156, n_n197}, x4238x);
	defparam lut_9905.LUT_SIZE = 7;
	defparam lut_9905.mask = 128'h0fff0fff7fff7fff1000010000000000;

	lut_sub lut_9908 ({sk[1847], x735x, n_n126, x720x, x1818x, n_n216, x4238x}, n_n3921);
	defparam lut_9908.LUT_SIZE = 7;
	defparam lut_9908.mask = 128'h0fff0fff7fff7fff5555555555555f7f;

	lut_sub lut_9912 ({sk[1848], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1270x);
	defparam lut_9912.LUT_SIZE = 7;
	defparam lut_9912.mask = 128'h0fff0fff7fff7fff7000070000700007;

	lut_sub lut_9921 ({sk[1849], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1269x);
	defparam lut_9921.LUT_SIZE = 7;
	defparam lut_9921.mask = 128'h0fff0fff7fff7fff3000030000700007;

	lut_sub lut_9928 ({sk[1850], i_8_, n_n17, x735x, n_n63, x125x, x1269x}, x17573x);
	defparam lut_9928.LUT_SIZE = 7;
	defparam lut_9928.mask = 128'h0fff0fff7fff7fff0000007f00000000;

	lut_sub lut_9932 ({sk[1851], x740x, n_n161, n_n47, n_n63, x176x, x1388x}, x18192x);
	defparam lut_9932.LUT_SIZE = 7;
	defparam lut_9932.mask = 128'h0fff0fff7fff7fff000f000f000f777f;

	lut_sub lut_9936 ({sk[1852], n_n46, n_n47, x125x, x1228x, x1227x, x1387x}, x18193x);
	defparam lut_9936.LUT_SIZE = 7;
	defparam lut_9936.mask = 128'h0fff0fff7fff7fff000077ff0f0f7fff;

	lut_sub lut_9941 ({sk[1853], x157x, n_n46, n_n177, n_n47, x719x, x174x}, x18200x);
	defparam lut_9941.LUT_SIZE = 7;
	defparam lut_9941.mask = 128'h0fff0fff7fff7fff000055770f0f5f7f;

	lut_sub lut_9945 ({sk[1854], x740x, n_n161, n_n47, x18198x, x18199x, x1546x}, x18201x);
	defparam lut_9945.LUT_SIZE = 7;
	defparam lut_9945.mask = 128'h0fff0fff7fff7fff003f003f003f557f;

	lut_sub lut_9949 ({sk[1855], i_8_, x740x, n_n18, x133x, x158x, x1895x}, x18203x);
	defparam lut_9949.LUT_SIZE = 7;
	defparam lut_9949.mask = 128'h0fff0fff7fff7fff0000007f00000000;

	lut_sub lut_9953 ({sk[1856], n_n46, n_n47, x55x, x158x, x134x, x1888x}, x18204x);
	defparam lut_9953.LUT_SIZE = 7;
	defparam lut_9953.mask = 128'h0fff0fff7fff7fff00005fff33337fff;

	lut_sub lut_9958 ({sk[1857], i_14_, i_13_, i_12_, i_15_, n_n170}, x1893x);
	defparam lut_9958.LUT_SIZE = 6;
	defparam lut_9958.mask = 64'h7777777700005154;

	lut_sub lut_9965 ({sk[1858], i_14_, i_13_, i_12_, i_15_, n_n170}, x1271x);
	defparam lut_9965.LUT_SIZE = 6;
	defparam lut_9965.mask = 64'h7777777715455154;

	lut_sub lut_9978 ({sk[1859], i_14_, i_13_, i_12_, i_15_, n_n199}, x1272x);
	defparam lut_9978.LUT_SIZE = 6;
	defparam lut_9978.mask = 64'h7777777701015154;

	lut_sub lut_9987 ({sk[1860], i_7_, i_8_, i_6_, x46x, x735x}, n_n4692);
	defparam lut_9987.LUT_SIZE = 6;
	defparam lut_9987.mask = 64'h7777777700001000;

	lut_sub lut_9989 ({sk[1861], i_14_, i_13_, i_12_, i_15_, n_n216}, x1275x);
	defparam lut_9989.LUT_SIZE = 6;
	defparam lut_9989.mask = 64'h7777777714045000;

	lut_sub lut_9995 ({sk[1862], i_15_, n_n89, n_n41, n_n42, n_n216, n_n213}, x21421x);
	defparam lut_9995.LUT_SIZE = 7;
	defparam lut_9995.mask = 128'h0fff0fff7fff7ffffffff0f0ffeef0e0;

	lut_sub lut_10004 ({sk[1863], n_n42, n_n43, x52x, n_n115, n_n137, x21421x}, n_n1885);
	defparam lut_10004.LUT_SIZE = 7;
	defparam lut_10004.mask = 128'h0fff0fff7fff7fffaaaabfbfbfffbfff;

	lut_sub lut_10011 ({sk[1864], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1285x);
	defparam lut_10011.LUT_SIZE = 7;
	defparam lut_10011.mask = 128'h0fff0fff7fff7fff0707700700007700;

	lut_sub lut_10024 ({sk[1865], n_n30, n_n7294, n_n129, x527x, x551x, x18839x}, x18841x);
	defparam lut_10024.LUT_SIZE = 7;
	defparam lut_10024.mask = 128'h0fff0fff7fff7fff7f7fffff7fffffff;

	lut_sub lut_10030 ({sk[1866], i_8_, n_n157, n_n31, x734x, x1285x, x321x}, x18845x);
	defparam lut_10030.LUT_SIZE = 7;
	defparam lut_10030.mask = 128'h0fff0fff7fff7fff0077037700770077;

	lut_sub lut_10034 ({sk[1867], n_n31, n_n2, n_n141, n_n137, x994x, x1198x}, x21363x);
	defparam lut_10034.LUT_SIZE = 7;
	defparam lut_10034.mask = 128'h0fff0fff7fff7fffffffaaaac0008000;

	lut_sub lut_10039 ({sk[1868], i_14_, i_13_, i_12_, i_15_, n_n149, n_n177}, x1290x);
	defparam lut_10039.LUT_SIZE = 7;
	defparam lut_10039.mask = 128'h0fff0fff7fff7fff0555500550075750;

	lut_sub lut_10052 ({sk[1869], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1289x);
	defparam lut_10052.LUT_SIZE = 7;
	defparam lut_10052.mask = 128'h0fff0fff7fff7fff0373700330033330;

	lut_sub lut_10065 ({sk[1870], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1292x);
	defparam lut_10065.LUT_SIZE = 7;
	defparam lut_10065.mask = 128'h0fff0fff7fff7fff0575700550055550;

	lut_sub lut_10078 ({sk[1871], i_14_, i_13_, i_12_, i_15_, n_n149, n_n216}, x1291x);
	defparam lut_10078.LUT_SIZE = 7;
	defparam lut_10078.mask = 128'h0fff0fff7fff7fff0333350330533330;

	lut_sub lut_10091 ({sk[1872], i_14_, i_13_, i_12_, i_15_, n_n191}, x1402x);
	defparam lut_10091.LUT_SIZE = 6;
	defparam lut_10091.mask = 64'h7777777715014040;

	lut_sub lut_10098 ({sk[1873], i_14_, i_13_, i_12_, i_15_, n_n191}, x1298x);
	defparam lut_10098.LUT_SIZE = 6;
	defparam lut_10098.mask = 64'h7777777700051014;

	lut_sub lut_10104 ({sk[1874], i_14_, i_13_, i_12_, i_15_, n_n149}, x1303x);
	defparam lut_10104.LUT_SIZE = 6;
	defparam lut_10104.mask = 64'h7777777700051114;

	lut_sub lut_10111 ({sk[1875], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1302x);
	defparam lut_10111.LUT_SIZE = 7;
	defparam lut_10111.mask = 128'h0fff0fff7fff7fff0000007707030370;

	lut_sub lut_10122 ({sk[1876], i_15_, x59x, n_n216, n_n209, x1303x, x402x}, x21342x);
	defparam lut_10122.LUT_SIZE = 7;
	defparam lut_10122.mask = 128'h0fff0fff7fff7fff8888000088800000;

	lut_sub lut_10126 ({sk[1877], n_n31, n_n30, n_n142, x290x, x401x, x21342x}, x19466x);
	defparam lut_10126.LUT_SIZE = 7;
	defparam lut_10126.mask = 128'h0fff0fff7fff7fff0000afaf33ffbfff;

	lut_sub lut_10131 ({sk[1878], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1305x);
	defparam lut_10131.LUT_SIZE = 7;
	defparam lut_10131.mask = 128'h0fff0fff7fff7fff0000003707070770;

	lut_sub lut_10143 ({sk[1879], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1304x);
	defparam lut_10143.LUT_SIZE = 7;
	defparam lut_10143.mask = 128'h0fff0fff7fff7fff0000007303030330;

	lut_sub lut_10151 ({sk[1880], i_14_, i_13_, i_12_, i_15_, n_n191}, x1672x);
	defparam lut_10151.LUT_SIZE = 6;
	defparam lut_10151.mask = 64'h7777777700011114;

	lut_sub lut_10157 ({sk[1881], i_14_, i_13_, i_12_, i_15_, n_n216}, x1671x);
	defparam lut_10157.LUT_SIZE = 6;
	defparam lut_10157.mask = 64'h7777777700051004;

	lut_sub lut_10162 ({sk[1882], n_n31, n_n30, x1305x, x1304x, x1672x, x1671x}, n_n756);
	defparam lut_10162.LUT_SIZE = 7;
	defparam lut_10162.mask = 128'h0fff0fff7fff7fff000055ff3f3f7fff;

	lut_sub lut_10167 ({sk[1883], i_14_, i_13_, i_12_, i_15_, n_n170}, x237x);
	defparam lut_10167.LUT_SIZE = 6;
	defparam lut_10167.mask = 64'h7777777700011004;

	lut_sub lut_10171 ({sk[1884], i_14_, i_13_, i_12_, i_15_, n_n184}, x1310x);
	defparam lut_10171.LUT_SIZE = 6;
	defparam lut_10171.mask = 64'h7777777705004144;

	lut_sub lut_10178 ({sk[1885], i_14_, i_13_, i_12_, i_15_, n_n184}, x346x);
	defparam lut_10178.LUT_SIZE = 6;
	defparam lut_10178.mask = 64'h7777777705000000;

	lut_sub lut_10181 ({sk[1886], n_n36, n_n34, n_n191, x720x, x1310x, x346x}, n_n367);
	defparam lut_10181.LUT_SIZE = 7;
	defparam lut_10181.mask = 128'h0fff0fff7fff7fff0000555f3333777f;

	lut_sub lut_10185 ({sk[1887], i_14_, i_13_, i_12_, i_15_, n_n170}, x161x);
	defparam lut_10185.LUT_SIZE = 6;
	defparam lut_10185.mask = 64'h7777777700000104;

	lut_sub lut_10188 ({sk[1888], i_14_, i_13_, i_12_, i_15_, n_n170}, x329x);
	defparam lut_10188.LUT_SIZE = 6;
	defparam lut_10188.mask = 64'h7777777701004040;

	lut_sub lut_10192 ({sk[1889], i_14_, i_13_, i_12_, i_15_, n_n177, n_n125}, n_n4657);
	defparam lut_10192.LUT_SIZE = 7;
	defparam lut_10192.mask = 128'h0fff0fff7fff7fff0000010000100001;

	lut_sub lut_10196 ({sk[1890], i_14_, i_13_, i_12_, i_15_, n_n191, n_n216}, x1313x);
	defparam lut_10196.LUT_SIZE = 7;
	defparam lut_10196.mask = 128'h0fff0fff7fff7fff3000070000700007;

	lut_sub lut_10204 ({sk[1891], i_14_, i_13_, i_12_, i_15_, n_n156, n_n191}, x1314x);
	defparam lut_10204.LUT_SIZE = 7;
	defparam lut_10204.mask = 128'h0fff0fff7fff7fff7000070000700007;

	lut_sub lut_10213 ({sk[1892], n_n156, n_n124, n_n177, n_n47, x80x, x285x}, x21415x);
	defparam lut_10213.LUT_SIZE = 7;
	defparam lut_10213.mask = 128'h0fff0fff7fff7fff0303035703035757;

	lut_sub lut_10222 ({sk[1893], n_n134, x157x, n_n46, n_n47, x78x, x174x}, x21443x);
	defparam lut_10222.LUT_SIZE = 7;
	defparam lut_10222.mask = 128'h0fff0fff7fff7ffffca8f0a0fc00f000;

	lut_sub lut_10227 ({sk[1894], i_14_, i_13_, i_12_, i_15_, n_n216}, x1315x);
	defparam lut_10227.LUT_SIZE = 6;
	defparam lut_10227.mask = 64'h7777777740100401;

	lut_sub lut_10232 ({sk[1895], i_14_, i_13_, i_12_, i_15_, n_n156, n_n216}, x1317x);
	defparam lut_10232.LUT_SIZE = 7;
	defparam lut_10232.mask = 128'h0fff0fff7fff7fff0333303333533335;

	lut_sub lut_10247 ({sk[1896], i_14_, i_13_, i_12_, i_15_, n_n216}, x1316x);
	defparam lut_10247.LUT_SIZE = 6;
	defparam lut_10247.mask = 64'h7777777740100401;

	lut_sub lut_10252 ({sk[1897], i_14_, i_13_, i_12_, i_15_, n_n177}, x1489x);
	defparam lut_10252.LUT_SIZE = 6;
	defparam lut_10252.mask = 64'h7777777711015154;

	lut_sub lut_10262 ({sk[1898], i_14_, i_13_, i_12_, i_15_, n_n177}, x1319x);
	defparam lut_10262.LUT_SIZE = 6;
	defparam lut_10262.mask = 64'h7777777715455154;

	lut_sub lut_10275 ({sk[1899], i_14_, i_13_, i_12_, i_15_, n_n156, n_n177}, x1318x);
	defparam lut_10275.LUT_SIZE = 7;
	defparam lut_10275.mask = 128'h0fff0fff7fff7fff0050505003030300;

	lut_sub lut_10282 ({sk[1900], i_14_, i_13_, i_12_, i_15_, n_n156}, x1488x);
	defparam lut_10282.LUT_SIZE = 6;
	defparam lut_10282.mask = 64'h7777777740100401;

	lut_sub lut_10287 ({sk[1901], i_14_, i_13_, i_12_, i_15_, n_n177, n_n191}, x17625x);
	defparam lut_10287.LUT_SIZE = 7;
	defparam lut_10287.mask = 128'h0fff0fff7fff7fff3000070000700005;

	lut_sub lut_10294 ({sk[1902], i_14_, i_13_, i_12_, i_15_, n_n177, n_n191}, x1320x);
	defparam lut_10294.LUT_SIZE = 7;
	defparam lut_10294.mask = 128'h0fff0fff7fff7fff7000070000500005;

	lut_sub lut_10301 ({sk[1903], i_14_, i_13_, i_12_, i_15_, n_n191}, x240x);
	defparam lut_10301.LUT_SIZE = 6;
	defparam lut_10301.mask = 64'h7777777711040000;

	lut_sub lut_10305 ({sk[1904], n_n41, n_n40, x51x, n_n176, x361x, x240x}, x17646x);
	defparam lut_10305.LUT_SIZE = 7;
	defparam lut_10305.mask = 128'h0fff0fff7fff7fff333333ff7fff7fff;

	lut_sub lut_10311 ({sk[1905], i_14_, i_13_, i_12_, i_15_, n_n191}, x1832x);
	defparam lut_10311.LUT_SIZE = 6;
	defparam lut_10311.mask = 64'h7777777700015154;

	lut_sub lut_10319 ({sk[1906], i_14_, i_13_, i_12_, i_15_, n_n191}, x1450x);
	defparam lut_10319.LUT_SIZE = 6;
	defparam lut_10319.mask = 64'h7777777711055154;

	lut_sub lut_10330 ({sk[1907], x740x, n_n200, x714x, x17002x, x1832x, x1450x}, x17647x);
	defparam lut_10330.LUT_SIZE = 7;
	defparam lut_10330.mask = 128'h0fff0fff7fff7fff0003000300035557;

	lut_sub lut_10333 ({sk[1908], x714x, x17002x, n_n155, x215x, x100x, x1900x}, x17650x);
	defparam lut_10333.LUT_SIZE = 7;
	defparam lut_10333.mask = 128'h0fff0fff7fff7fff0000000000007fff;

	lut_sub lut_10338 ({sk[1909], i_14_, i_13_, i_12_, i_15_, n_n177}, x1691x);
	defparam lut_10338.LUT_SIZE = 6;
	defparam lut_10338.mask = 64'h7777777700015154;

	lut_sub lut_10346 ({sk[1910], n_n41, n_n40, n_n83, n_n171, x224x, x1691x}, x17651x);
	defparam lut_10346.LUT_SIZE = 7;
	defparam lut_10346.mask = 128'h0fff0fff7fff7fff00007fff0fff7fff;

	lut_sub lut_10353 ({sk[1911], i_14_, i_13_, i_12_, i_15_, n_n191}, x1322x);
	defparam lut_10353.LUT_SIZE = 6;
	defparam lut_10353.mask = 64'h7777777740100401;

	lut_sub lut_10358 ({sk[1912], n_n40, x714x, x17002x, n_n214, x180x, x142x}, x17657x);
	defparam lut_10358.LUT_SIZE = 7;
	defparam lut_10358.mask = 128'h0fff0fff7fff7fff0000007f3f3f3f7f;

	lut_sub lut_10364 ({sk[1913], n_n41, n_n40, x85x, x142x, x524x, x359x}, x21411x);
	defparam lut_10364.LUT_SIZE = 7;
	defparam lut_10364.mask = 128'h0fff0fff7fff7fff8888800088008000;

	lut_sub lut_10368 ({sk[1914], i_8_, n_n156, x740x, n_n16, x726x, x728x}, x17668x);
	defparam lut_10368.LUT_SIZE = 7;
	defparam lut_10368.mask = 128'h0fff0fff7fff7fff0000000700000007;

	lut_sub lut_10373 ({sk[1915], i_7_, i_8_, i_6_, x740x, x248x, x17668x}, x17671x);
	defparam lut_10373.LUT_SIZE = 7;
	defparam lut_10373.mask = 128'h0fff0fff7fff7fff5557555755555555;

	lut_sub lut_10377 ({sk[1916], i_14_, i_13_, i_12_, i_15_, n_n156}, x1871x);
	defparam lut_10377.LUT_SIZE = 6;
	defparam lut_10377.mask = 64'h7777777711054040;

	lut_sub lut_10384 ({sk[1917], i_8_, x740x, n_n17, n_n4604, x363x, x1871x}, x17676x);
	defparam lut_10384.LUT_SIZE = 7;
	defparam lut_10384.mask = 128'h0fff0fff7fff7fff3f3f3f7f3f3f3f3f;

	lut_sub lut_10388 ({sk[1918], i_14_, i_13_, i_12_, i_15_, n_n156, n_n216}, x1692x);
	defparam lut_10388.LUT_SIZE = 7;
	defparam lut_10388.mask = 128'h0fff0fff7fff7fff0000050003530335;

	lut_sub lut_10396 ({sk[1919], n_n41, n_n40, x90x, n_n142, x1824x, x1692x}, x17677x);
	defparam lut_10396.LUT_SIZE = 7;
	defparam lut_10396.mask = 128'h0fff0fff7fff7fff000055ff3f3f7fff;

	lut_sub lut_10401 ({sk[1920], i_14_, i_13_, i_12_, i_15_, n_n156, n_n191}, x1323x);
	defparam lut_10401.LUT_SIZE = 7;
	defparam lut_10401.mask = 128'h0fff0fff7fff7fff7000070000700005;

	lut_sub lut_10409 ({sk[1921], x740x, n_n200, n_n138, x172x, n_n63, x503x}, x17681x);
	defparam lut_10409.LUT_SIZE = 7;
	defparam lut_10409.mask = 128'h0fff0fff7fff7fff5555555555557fff;

	lut_sub lut_10414 ({sk[1922], n_n38, n_n39, n_n177, x719x, n_n84, x110x}, x17670x);
	defparam lut_10414.LUT_SIZE = 7;
	defparam lut_10414.mask = 128'h0fff0fff7fff7fff0000555f777f777f;

	lut_sub lut_10420 ({sk[1923], i_14_, i_13_, i_12_, i_15_, n_n156}, x1895x);
	defparam lut_10420.LUT_SIZE = 6;
	defparam lut_10420.mask = 64'h7777777711014044;

	lut_sub lut_10427 ({sk[1924], n_n46, n_n47, n_n63, x176x, x134x, x212x}, x21444x);
	defparam lut_10427.LUT_SIZE = 7;
	defparam lut_10427.mask = 128'h0fff0fff7fff7ffffffff00088888000;

	lut_sub lut_10432 ({sk[1925], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1324x);
	defparam lut_10432.LUT_SIZE = 7;
	defparam lut_10432.mask = 128'h0fff0fff7fff7fff7000070000700007;

	lut_sub lut_10441 ({sk[1926], i_14_, i_13_, i_12_, i_15_, n_n184}, x1379x);
	defparam lut_10441.LUT_SIZE = 6;
	defparam lut_10441.mask = 64'h7777777740100401;

	lut_sub lut_10446 ({sk[1927], i_14_, i_13_, i_12_, i_15_, n_n184}, x217x);
	defparam lut_10446.LUT_SIZE = 6;
	defparam lut_10446.mask = 64'h7777777700100401;

	lut_sub lut_10450 ({sk[1928], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x18395x);
	defparam lut_10450.LUT_SIZE = 7;
	defparam lut_10450.mask = 128'h0fff0fff7fff7fff7000050000500005;

	lut_sub lut_10456 ({sk[1929], i_14_, i_13_, i_12_, i_15_, n_n149}, x1328x);
	defparam lut_10456.LUT_SIZE = 6;
	defparam lut_10456.mask = 64'h7777777715055044;

	lut_sub lut_10466 ({sk[1930], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1327x);
	defparam lut_10466.LUT_SIZE = 7;
	defparam lut_10466.mask = 128'h0fff0fff7fff7fff0333003337057570;

	lut_sub lut_10481 ({sk[1931], i_14_, i_13_, i_12_, i_15_, n_n199}, x1330x);
	defparam lut_10481.LUT_SIZE = 6;
	defparam lut_10481.mask = 64'h7777777715454044;

	lut_sub lut_10491 ({sk[1932], i_14_, i_13_, i_12_, i_15_, n_n216}, x1329x);
	defparam lut_10491.LUT_SIZE = 6;
	defparam lut_10491.mask = 64'h7777777700001154;

	lut_sub lut_10497 ({sk[1933], i_14_, i_13_, i_12_, i_15_, n_n41, n_n216}, x3503x);
	defparam lut_10497.LUT_SIZE = 7;
	defparam lut_10497.mask = 128'h0fff0fff7fff7fff1000010000000000;

	lut_sub lut_10500 ({sk[1934], i_14_, i_13_, i_12_, i_15_, n_n40, n_n216}, x3497x);
	defparam lut_10500.LUT_SIZE = 7;
	defparam lut_10500.mask = 128'h0fff0fff7fff7fff1000010000000000;

	lut_sub lut_10503 ({sk[1935], n_n5060, x461x, n_n5061, x3501x, x3502x, x4906x}, x18273x);
	defparam lut_10503.LUT_SIZE = 7;
	defparam lut_10503.mask = 128'h0fff0fff7fff7fff7fffffffffffffff;

	lut_sub lut_10510 ({sk[1936], i_14_, i_13_, i_12_, i_15_, n_n184}, x1820x);
	defparam lut_10510.LUT_SIZE = 6;
	defparam lut_10510.mask = 64'h7777777740100401;

	lut_sub lut_10515 ({sk[1937], x725x, n_n40, n_n184, n_n191, x719x, x88x}, x21447x);
	defparam lut_10515.LUT_SIZE = 7;
	defparam lut_10515.mask = 128'h0fff0fff7fff7fffffffa888ffffa800;

	lut_sub lut_10520 ({sk[1938], n_n41, n_n138, x172x, x3497x, x1820x, x21447x}, x18274x);
	defparam lut_10520.LUT_SIZE = 7;
	defparam lut_10520.mask = 128'h0fff0fff7fff7fffafafafafbfffffff;

	lut_sub lut_10526 ({sk[1939], i_14_, i_13_, i_12_, i_15_, n_n177}, x469x);
	defparam lut_10526.LUT_SIZE = 6;
	defparam lut_10526.mask = 64'h7777777710040000;

	lut_sub lut_10529 ({sk[1940], i_14_, i_13_, i_12_, i_15_, n_n170}, x1331x);
	defparam lut_10529.LUT_SIZE = 6;
	defparam lut_10529.mask = 64'h7777777715055154;

	lut_sub lut_10541 ({sk[1941], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1433x);
	defparam lut_10541.LUT_SIZE = 7;
	defparam lut_10541.mask = 128'h0fff0fff7fff7fff0507005773033330;

	lut_sub lut_10555 ({sk[1942], i_8_, i_1_, i_2_, i_0_, x17002x, x1433x}, x3484x);
	defparam lut_10555.LUT_SIZE = 7;
	defparam lut_10555.mask = 128'h0fff0fff7fff7fff0000000010000000;

	lut_sub lut_10557 ({sk[1943], i_14_, i_13_, i_12_, i_15_, n_n149}, x1432x);
	defparam lut_10557.LUT_SIZE = 6;
	defparam lut_10557.mask = 64'h7777777715455044;

	lut_sub lut_10568 ({sk[1944], n_n71, n_n41, n_n40, n_n150, x118x, x1432x}, x18283x);
	defparam lut_10568.LUT_SIZE = 7;
	defparam lut_10568.mask = 128'h0fff0fff7fff7fff00770f7f0077ffff;

	lut_sub lut_10573 ({sk[1945], i_8_, i_1_, i_2_, i_0_, x17002x, x218x}, x3482x);
	defparam lut_10573.LUT_SIZE = 7;
	defparam lut_10573.mask = 128'h0fff0fff7fff7fff0000000010000000;

	lut_sub lut_10575 ({sk[1946], i_15_, x714x, x17002x, n_n216, n_n209, x728x}, x3480x);
	defparam lut_10575.LUT_SIZE = 7;
	defparam lut_10575.mask = 128'h0fff0fff7fff7fff0000000500000007;

	lut_sub lut_10578 ({sk[1947], i_14_, i_13_, i_12_, i_15_, n_n156}, x198x);
	defparam lut_10578.LUT_SIZE = 6;
	defparam lut_10578.mask = 64'h7777777701014000;

	lut_sub lut_10582 ({sk[1948], i_14_, i_13_, i_12_, i_15_, n_n156}, x1332x);
	defparam lut_10582.LUT_SIZE = 6;
	defparam lut_10582.mask = 64'h7777777701015044;

	lut_sub lut_10589 ({sk[1949], n_n40, x59x, n_n140, x3506x, x3503x, x1332x}, x18286x);
	defparam lut_10589.LUT_SIZE = 7;
	defparam lut_10589.mask = 128'h0fff0fff7fff7fff3f3f3f3f7fffffff;

	lut_sub lut_10595 ({sk[1950], n_n41, n_n40, x218x, x212x, x1889x, x21448x}, x18287x);
	defparam lut_10595.LUT_SIZE = 7;
	defparam lut_10595.mask = 128'h0fff0fff7fff7fffaaaabbbbafffbfff;

	lut_sub lut_10600 ({sk[1951], i_14_, i_13_, i_12_, i_15_, n_n177}, x1337x);
	defparam lut_10600.LUT_SIZE = 6;
	defparam lut_10600.mask = 64'h7777777714445000;

	lut_sub lut_10607 ({sk[1952], i_9_, i_10_, i_8_, i_11_, n_n17, x285x}, x19303x);
	defparam lut_10607.LUT_SIZE = 7;
	defparam lut_10607.mask = 128'h0fff0fff7fff7fff0000100000000010;

	lut_sub lut_10610 ({sk[1953], i_14_, i_13_, i_12_, i_15_, n_n47, n_n216}, x21433x);
	defparam lut_10610.LUT_SIZE = 7;
	defparam lut_10610.mask = 128'h0fff0fff7fff7ffffffffffffffeeeef;

	lut_sub lut_10617 ({sk[1954], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1348x);
	defparam lut_10617.LUT_SIZE = 7;
	defparam lut_10617.mask = 128'h0fff0fff7fff7fff0000007703030370;

	lut_sub lut_10627 ({sk[1955], i_14_, i_13_, i_12_, i_15_, n_n177}, x280x);
	defparam lut_10627.LUT_SIZE = 6;
	defparam lut_10627.mask = 64'h7777777700050004;

	lut_sub lut_10631 ({sk[1956], x46x, n_n197, n_n212, x48x, x1348x, x280x}, n_n785);
	defparam lut_10631.LUT_SIZE = 7;
	defparam lut_10631.mask = 128'h0fff0fff7fff7fff00773f7f00ff3fff;

	lut_sub lut_10637 ({sk[1957], i_14_, i_13_, i_12_, i_15_, n_n149, n_n170}, x19508x);
	defparam lut_10637.LUT_SIZE = 7;
	defparam lut_10637.mask = 128'h0fff0fff7fff7fff0000005503030350;

	lut_sub lut_10644 ({sk[1958], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1349x);
	defparam lut_10644.LUT_SIZE = 7;
	defparam lut_10644.mask = 128'h0fff0fff7fff7fff0000007703030370;

	lut_sub lut_10654 ({sk[1959], i_8_, x132x, x46x, n_n17, x735x, n_n212}, x19510x);
	defparam lut_10654.LUT_SIZE = 7;
	defparam lut_10654.mask = 128'h0fff0fff7fff7fff0003575700005555;

	lut_sub lut_10658 ({sk[1960], x735x, n_n200, n_n212, x280x, x19508x, x1349x}, x19511x);
	defparam lut_10658.LUT_SIZE = 7;
	defparam lut_10658.mask = 128'h0fff0fff7fff7fff0055005500553f7f;

	lut_sub lut_10662 ({sk[1961], i_7_, i_8_, i_6_, x735x, x47x}, x629x);
	defparam lut_10662.LUT_SIZE = 6;
	defparam lut_10662.mask = 64'h7777777700001000;

	lut_sub lut_10664 ({sk[1962], i_9_, i_10_, i_11_, i_15_, n_n207, n_n209}, x1353x);
	defparam lut_10664.LUT_SIZE = 7;
	defparam lut_10664.mask = 128'h0fff0fff7fff7fff0000007300000073;

	lut_sub lut_10671 ({sk[1963], n_n197, n_n212, x151x, x48x, x47x, x1353x}, x19516x);
	defparam lut_10671.LUT_SIZE = 7;
	defparam lut_10671.mask = 128'h0fff0fff7fff7fff00007fff77ff7fff;

	lut_sub lut_10679 ({sk[1964], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1356x);
	defparam lut_10679.LUT_SIZE = 7;
	defparam lut_10679.mask = 128'h0fff0fff7fff7fff0077000070033030;

	lut_sub lut_10689 ({sk[1965], i_14_, i_13_, i_12_, i_15_, n_n191}, x166x);
	defparam lut_10689.LUT_SIZE = 6;
	defparam lut_10689.mask = 64'h7777777700000144;

	lut_sub lut_10693 ({sk[1966], i_14_, i_13_, i_12_, i_15_, n_n177}, x325x);
	defparam lut_10693.LUT_SIZE = 6;
	defparam lut_10693.mask = 64'h7777777700000144;

	lut_sub lut_10697 ({sk[1967], i_14_, i_13_, i_12_, i_15_, n_n177}, x354x);
	defparam lut_10697.LUT_SIZE = 6;
	defparam lut_10697.mask = 64'h7777777705004000;

	lut_sub lut_10701 ({sk[1968], n_n197, n_n212, x1356x, x166x, x325x, x354x}, n_n339);
	defparam lut_10701.LUT_SIZE = 7;
	defparam lut_10701.mask = 128'h0fff0fff7fff7fff000077ff0fff7fff;

	lut_sub lut_10707 ({sk[1969], i_9_, i_10_, i_11_, x726x, x728x}, x1358x);
	defparam lut_10707.LUT_SIZE = 6;
	defparam lut_10707.mask = 64'h7777777700055035;

	lut_sub lut_10712 ({sk[1970], i_9_, i_10_, i_11_, x734x, n_n126, x728x}, x2031x);
	defparam lut_10712.LUT_SIZE = 7;
	defparam lut_10712.mask = 128'h0fff0fff7fff7fff0000000101000001;

	lut_sub lut_10716 ({sk[1971], n_n124, x734x, n_n126, n_n136, x1358x, x2031x}, n_n406);
	defparam lut_10716.LUT_SIZE = 7;
	defparam lut_10716.mask = 128'h0fff0fff7fff7fff5555555f55557f7f;

	lut_sub lut_10721 ({sk[1972], i_9_, i_10_, i_11_, x726x, x728x}, x19784x);
	defparam lut_10721.LUT_SIZE = 6;
	defparam lut_10721.mask = 64'h7777777700700550;

	lut_sub lut_10726 ({sk[1973], n_n101, x419x, n_n108, x249x, n_n56, x19784x}, x19786x);
	defparam lut_10726.LUT_SIZE = 7;
	defparam lut_10726.mask = 128'h0fff0fff7fff7fff007fffff337fffff;

	lut_sub lut_10732 ({sk[1974], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1363x);
	defparam lut_10732.LUT_SIZE = 7;
	defparam lut_10732.mask = 128'h0fff0fff7fff7fff0077000070077070;

	lut_sub lut_10745 ({sk[1975], n_n170, x723x, x161x, x236x, x325x, x282x}, x21335x);
	defparam lut_10745.LUT_SIZE = 7;
	defparam lut_10745.mask = 128'h0fff0fff7fff7fff8000800080000000;

	lut_sub lut_10748 ({sk[1976], x735x, n_n200, n_n212, x1363x, x354x, x21335x}, n_n338);
	defparam lut_10748.LUT_SIZE = 7;
	defparam lut_10748.mask = 128'h0fff0fff7fff7fff000f000f000fbbbf;

	lut_sub lut_10752 ({sk[1977], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1366x);
	defparam lut_10752.LUT_SIZE = 7;
	defparam lut_10752.mask = 128'h0fff0fff7fff7fff0077000070077070;

	lut_sub lut_10765 ({sk[1978], x735x, n_n200, n_n212, x125x, x176x, x123x}, n_n3925);
	defparam lut_10765.LUT_SIZE = 7;
	defparam lut_10765.mask = 128'h0fff0fff7fff7fff000f000f000f777f;

	lut_sub lut_10769 ({sk[1979], i_14_, i_13_, i_12_, i_15_, n_n156, n_n177}, x1373x);
	defparam lut_10769.LUT_SIZE = 7;
	defparam lut_10769.mask = 128'h0fff0fff7fff7fff0555505557035770;

	lut_sub lut_10785 ({sk[1980], i_14_, i_13_, i_12_, i_15_, n_n156}, x1830x);
	defparam lut_10785.LUT_SIZE = 6;
	defparam lut_10785.mask = 64'h7777777700001114;

	lut_sub lut_10790 ({sk[1981], n_n123, n_n125, x155x, x1851x, x1373x, x1830x}, n_n3828);
	defparam lut_10790.LUT_SIZE = 7;
	defparam lut_10790.mask = 128'h0fff0fff7fff7fff00005fff33337fff;

	lut_sub lut_10795 ({sk[1982], i_14_, i_13_, i_12_, i_15_, n_n177}, x1877x);
	defparam lut_10795.LUT_SIZE = 6;
	defparam lut_10795.mask = 64'h7777777715450000;

	lut_sub lut_10802 ({sk[1983], i_9_, i_10_, i_8_, i_11_, n_n17, x285x}, x17700x);
	defparam lut_10802.LUT_SIZE = 7;
	defparam lut_10802.mask = 128'h0fff0fff7fff7fff0000000001001010;

	lut_sub lut_10806 ({sk[1984], i_9_, i_8_, n_n18, x285x}, x21382x);
	defparam lut_10806.LUT_SIZE = 5;
	defparam lut_10806.mask = 32'h33ffffef;

	lut_sub lut_10811 ({sk[1985], i_14_, i_13_, i_12_, i_15_, n_n191}, x1378x);
	defparam lut_10811.LUT_SIZE = 6;
	defparam lut_10811.mask = 64'h7777777715455154;

	lut_sub lut_10824 ({sk[1986], n_n40, x172x, x247x, x212x, x3502x, x3482x}, x18455x);
	defparam lut_10824.LUT_SIZE = 7;
	defparam lut_10824.mask = 128'h0fff0fff7fff7fff777777777fffffff;

	lut_sub lut_10830 ({sk[1987], x725x, n_n40, n_n184, n_n191, x719x, x88x}, x21446x);
	defparam lut_10830.LUT_SIZE = 7;
	defparam lut_10830.mask = 128'h0fff0fff7fff7fffffffa888ffffa800;

	lut_sub lut_10835 ({sk[1988], n_n41, n_n138, x172x, x3497x, x1820x, x21446x}, x18456x);
	defparam lut_10835.LUT_SIZE = 7;
	defparam lut_10835.mask = 128'h0fff0fff7fff7fffafafafafbfffffff;

	lut_sub lut_10841 ({sk[1989], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1545x);
	defparam lut_10841.LUT_SIZE = 7;
	defparam lut_10841.mask = 128'h0fff0fff7fff7fff0737303755055550;

	lut_sub lut_10857 ({sk[1990], i_14_, i_13_, i_12_, i_15_, n_n177}, x1544x);
	defparam lut_10857.LUT_SIZE = 6;
	defparam lut_10857.mask = 64'h7777777711055154;

	lut_sub lut_10868 ({sk[1991], n_n40, x714x, x17002x, x397x, x1545x, x1544x}, n_n3184);
	defparam lut_10868.LUT_SIZE = 7;
	defparam lut_10868.mask = 128'h0fff0fff7fff7fff0f0f0f5f3f3f3f7f;

	lut_sub lut_10872 ({sk[1992], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1382x);
	defparam lut_10872.LUT_SIZE = 7;
	defparam lut_10872.mask = 128'h0fff0fff7fff7fff0373707333033330;

	lut_sub lut_10888 ({sk[1993], i_14_, i_13_, i_12_, i_15_, n_n170}, x1381x);
	defparam lut_10888.LUT_SIZE = 6;
	defparam lut_10888.mask = 64'h7777777715455154;

	lut_sub lut_10901 ({sk[1994], i_14_, i_13_, i_12_, i_15_, n_n156}, x1889x);
	defparam lut_10901.LUT_SIZE = 6;
	defparam lut_10901.mask = 64'h7777777714440000;

	lut_sub lut_10906 ({sk[1995], n_n40, n_n5319, x59x, x3506x, x3480x, x1889x}, x18461x);
	defparam lut_10906.LUT_SIZE = 7;
	defparam lut_10906.mask = 128'h0fff0fff7fff7fff3f3fffff7fffffff;

	lut_sub lut_10912 ({sk[1996], i_14_, i_13_, i_12_, i_15_, n_n149}, x1431x);
	defparam lut_10912.LUT_SIZE = 6;
	defparam lut_10912.mask = 64'h7777777715054044;

	lut_sub lut_10921 ({sk[1997], i_14_, i_13_, i_12_, i_15_, n_n156}, x1430x);
	defparam lut_10921.LUT_SIZE = 6;
	defparam lut_10921.mask = 64'h7777777701015044;

	lut_sub lut_10928 ({sk[1998], n_n41, n_n40, n_n140, x3503x, x1431x, x1430x}, x18462x);
	defparam lut_10928.LUT_SIZE = 7;
	defparam lut_10928.mask = 128'h0fff0fff7fff7fff0f0f5fff3f3f7fff;

	lut_sub lut_10933 ({sk[1999], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1384x);
	defparam lut_10933.LUT_SIZE = 7;
	defparam lut_10933.mask = 128'h0fff0fff7fff7fff0505005557075750;

	lut_sub lut_10947 ({sk[2000], i_14_, i_13_, i_12_, i_15_, n_n149}, x1383x);
	defparam lut_10947.LUT_SIZE = 6;
	defparam lut_10947.mask = 64'h7777777715455154;

	lut_sub lut_10960 ({sk[2001], n_n40, x714x, x17002x, x363x, x1384x, x1383x}, x18469x);
	defparam lut_10960.LUT_SIZE = 7;
	defparam lut_10960.mask = 128'h0fff0fff7fff7fff0f0f0f3f5f5f5f7f;

	lut_sub lut_10964 ({sk[2002], n_n41, n_n5319, n_n210, x611x, x391x, x1109x}, x18475x);
	defparam lut_10964.LUT_SIZE = 7;
	defparam lut_10964.mask = 128'h0fff0fff7fff7fff3f3fffff7fffffff;

	lut_sub lut_10970 ({sk[2003], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1425x);
	defparam lut_10970.LUT_SIZE = 7;
	defparam lut_10970.mask = 128'h0fff0fff7fff7fff7000070000700007;

	lut_sub lut_10979 ({sk[2004], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1424x);
	defparam lut_10979.LUT_SIZE = 7;
	defparam lut_10979.mask = 128'h0fff0fff7fff7fff7000070000700007;

	lut_sub lut_10988 ({sk[2005], i_8_, x740x, n_n18, n_n47, x1425x, x1424x}, x18476x);
	defparam lut_10988.LUT_SIZE = 7;
	defparam lut_10988.mask = 128'h0fff0fff7fff7fff0303035703030303;

	lut_sub lut_10991 ({sk[2006], i_14_, i_13_, i_12_, i_15_, n_n184, n_n216}, x1494x);
	defparam lut_10991.LUT_SIZE = 7;
	defparam lut_10991.mask = 128'h0fff0fff7fff7fff0505005557075750;

	lut_sub lut_11005 ({sk[2007], i_14_, i_13_, i_12_, i_15_, n_n191}, x1493x);
	defparam lut_11005.LUT_SIZE = 6;
	defparam lut_11005.mask = 64'h7777777715455154;

	lut_sub lut_11018 ({sk[2008], n_n40, x714x, x17002x, x361x, x1494x, x1493x}, n_n3186);
	defparam lut_11018.LUT_SIZE = 7;
	defparam lut_11018.mask = 128'h0fff0fff7fff7fff0f0f0f5f3f3f3f7f;

	lut_sub lut_11022 ({sk[2009], i_14_, i_13_, i_12_, i_15_, n_n199}, x1386x);
	defparam lut_11022.LUT_SIZE = 6;
	defparam lut_11022.mask = 64'h7777777715455154;

	lut_sub lut_11035 ({sk[2010], n_n40, x714x, x17002x, n_n103, x359x, x1386x}, x18486x);
	defparam lut_11035.LUT_SIZE = 7;
	defparam lut_11035.mask = 128'h0fff0fff7fff7fff3333337f7777777f;

	lut_sub lut_11040 ({sk[2011], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1388x);
	defparam lut_11040.LUT_SIZE = 7;
	defparam lut_11040.mask = 128'h0fff0fff7fff7fff3000070000700007;

	lut_sub lut_11048 ({sk[2012], i_14_, i_13_, i_12_, i_15_, n_n199}, x1387x);
	defparam lut_11048.LUT_SIZE = 6;
	defparam lut_11048.mask = 64'h7777777740100401;

	lut_sub lut_11053 ({sk[2013], n_n9, n_n144, n_n14, n_n10, n_n12, x170x}, n_n2954);
	defparam lut_11053.LUT_SIZE = 7;
	defparam lut_11053.mask = 128'h0fff0fff7fff7fff15153fff55557fff;

	lut_sub lut_11060 ({sk[2014], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1403x);
	defparam lut_11060.LUT_SIZE = 7;
	defparam lut_11060.mask = 128'h0fff0fff7fff7fff0000570000035700;

	lut_sub lut_11066 ({sk[2015], n_n36, n_n34, x720x, n_n199, x425x, x219x}, n_n813);
	defparam lut_11066.LUT_SIZE = 7;
	defparam lut_11066.mask = 128'h0fff0fff7fff7fff00007777555f777f;

	lut_sub lut_11071 ({sk[2016], i_14_, i_13_, i_12_, i_15_, n_n149}, x1412x);
	defparam lut_11071.LUT_SIZE = 6;
	defparam lut_11071.mask = 64'h7777777705004144;

	lut_sub lut_11078 ({sk[2017], i_9_, i_10_, i_11_, x720x, x726x, x727x}, x1411x);
	defparam lut_11078.LUT_SIZE = 7;
	defparam lut_11078.mask = 128'h0fff0fff7fff7fff00005f0000003300;

	lut_sub lut_11082 ({sk[2018], i_14_, i_13_, i_12_, i_15_, n_n216}, x1413x);
	defparam lut_11082.LUT_SIZE = 6;
	defparam lut_11082.mask = 64'h7777777705004144;

	lut_sub lut_11089 ({sk[2019], x712x, n_n36, n_n34, x720x, n_n199, x1413x}, n_n371);
	defparam lut_11089.LUT_SIZE = 7;
	defparam lut_11089.mask = 128'h0fff0fff7fff7fff00035557ffffffff;

	lut_sub lut_11093 ({sk[2020], i_9_, i_10_, i_11_, x728x}, x409x);
	defparam lut_11093.LUT_SIZE = 5;
	defparam lut_11093.mask = 32'h33ff0410;

	lut_sub lut_11096 ({sk[2021], i_14_, i_13_, i_12_, i_15_, n_n149}, x1880x);
	defparam lut_11096.LUT_SIZE = 6;
	defparam lut_11096.mask = 64'h7777777700015054;

	lut_sub lut_11103 ({sk[2022], i_14_, i_13_, i_12_, i_15_, n_n177}, x1817x);
	defparam lut_11103.LUT_SIZE = 6;
	defparam lut_11103.mask = 64'h7777777715454040;

	lut_sub lut_11112 ({sk[2023], i_14_, i_13_, i_12_, i_15_, n_n177, n_n191}, x1420x);
	defparam lut_11112.LUT_SIZE = 7;
	defparam lut_11112.mask = 128'h0fff0fff7fff7fff0505005555075550;

	lut_sub lut_11124 ({sk[2024], n_n125, x141x, x160x, x171x, x4055x, n_n4657}, x17734x);
	defparam lut_11124.LUT_SIZE = 7;
	defparam lut_11124.mask = 128'h0fff0fff7fff7fff777777777fffffff;

	lut_sub lut_11130 ({sk[2025], i_7_, i_8_, i_6_, x735x, x1817x, x1420x}, x17746x);
	defparam lut_11130.LUT_SIZE = 7;
	defparam lut_11130.mask = 128'h0fff0fff7fff7fff0005000300000000;

	lut_sub lut_11133 ({sk[2026], n_n123, n_n125, x51x, n_n176, x100x, x1313x}, x21383x);
	defparam lut_11133.LUT_SIZE = 7;
	defparam lut_11133.mask = 128'h0fff0fff7fff7fffffffc000aa008000;

	lut_sub lut_11138 ({sk[2027], i_14_, i_13_, i_12_, i_15_, n_n156, n_n191}, x1516x);
	defparam lut_11138.LUT_SIZE = 7;
	defparam lut_11138.mask = 128'h0fff0fff7fff7fff5000050000700007;

	lut_sub lut_11145 ({sk[2028], x157x, x735x, n_n200, n_n212, x174x, x1516x}, x17752x);
	defparam lut_11145.LUT_SIZE = 7;
	defparam lut_11145.mask = 128'h0fff0fff7fff7fff000000770f0f0f7f;

	lut_sub lut_11149 ({sk[2029], n_n212, x172x, n_n191, x719x, n_n63, x176x}, x17756x);
	defparam lut_11149.LUT_SIZE = 7;
	defparam lut_11149.mask = 128'h0fff0fff7fff7fff00000000777fffff;

	lut_sub lut_11154 ({sk[2030], i_14_, i_13_, i_12_, i_15_, n_n191}, x1596x);
	defparam lut_11154.LUT_SIZE = 6;
	defparam lut_11154.mask = 64'h7777777711055054;

	lut_sub lut_11164 ({sk[2031], i_14_, i_13_, i_12_, i_15_, n_n191, n_n216}, x1422x);
	defparam lut_11164.LUT_SIZE = 7;
	defparam lut_11164.mask = 128'h0fff0fff7fff7fff0555505000030000;

	lut_sub lut_11171 ({sk[2032], n_n123, n_n125, n_n214, x85x, x142x, x1596x}, x17763x);
	defparam lut_11171.LUT_SIZE = 7;
	defparam lut_11171.mask = 128'h0fff0fff7fff7fff000055553fff7fff;

	lut_sub lut_11176 ({sk[2033], n_n134, n_n53, n_n197, n_n212, x80x, x78x}, x17751x);
	defparam lut_11176.LUT_SIZE = 7;
	defparam lut_11176.mask = 128'h0fff0fff7fff7fff07070f0f07ff0fff;

	lut_sub lut_11181 ({sk[2034], i_7_, i_8_, i_6_, x735x, x1849x, x1518x}, x17755x);
	defparam lut_11181.LUT_SIZE = 7;
	defparam lut_11181.mask = 128'h0fff0fff7fff7fff0000000007000000;

	lut_sub lut_11184 ({sk[2035], i_9_, i_10_, i_11_, x729x, x717x, x730x}, x1429x);
	defparam lut_11184.LUT_SIZE = 7;
	defparam lut_11184.mask = 128'h0fff0fff7fff7fff00007f007f007f00;

	lut_sub lut_11194 ({sk[2036], n_n89, n_n14, x185x, x372x, n_n3, x87x}, x18364x);
	defparam lut_11194.LUT_SIZE = 7;
	defparam lut_11194.mask = 128'h0fff0fff7fff7fff131313ff333333ff;

	lut_sub lut_11199 ({sk[2037], i_14_, i_13_, i_12_, i_15_, n_n184}, x165x);
	defparam lut_11199.LUT_SIZE = 6;
	defparam lut_11199.mask = 64'h7777777700050004;

	lut_sub lut_11203 ({sk[2038], i_9_, i_10_, i_11_, i_15_, n_n207, n_n209}, x1438x);
	defparam lut_11203.LUT_SIZE = 7;
	defparam lut_11203.mask = 128'h0fff0fff7fff7fff7300000073000000;

	lut_sub lut_11210 ({sk[2039], x46x, n_n46, x124x, n_n47, x48x, x1438x}, n_n772);
	defparam lut_11210.LUT_SIZE = 7;
	defparam lut_11210.mask = 128'h0fff0fff7fff7fff070f77ff0f0f7fff;

	lut_sub lut_11218 ({sk[2040], x140x, n_n197, n_n212, n_n62, n_n64, x244x}, n_n433);
	defparam lut_11218.LUT_SIZE = 7;
	defparam lut_11218.mask = 128'h0fff0fff7fff7fff003f5f7f003fffff;

	lut_sub lut_11224 ({sk[2041], i_9_, i_10_, i_11_, x728x, x235x}, x1442x);
	defparam lut_11224.LUT_SIZE = 6;
	defparam lut_11224.mask = 64'h7777777755557555;

	lut_sub lut_11227 ({sk[2042], i_9_, i_10_, i_11_, x728x}, x19827x);
	defparam lut_11227.LUT_SIZE = 5;
	defparam lut_11227.mask = 32'h33ff4011;

	lut_sub lut_11231 ({sk[2043], i_9_, i_10_, i_11_, x728x}, x413x);
	defparam lut_11231.LUT_SIZE = 5;
	defparam lut_11231.mask = 32'h33ff4010;

	lut_sub lut_11234 ({sk[2044], n_n197, n_n212, x236x, x1442x, x19827x, x413x}, x19829x);
	defparam lut_11234.LUT_SIZE = 7;
	defparam lut_11234.mask = 128'h0fff0fff7fff7fff00005fff3f3f7fff;

	lut_sub lut_11240 ({sk[2045], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1444x);
	defparam lut_11240.LUT_SIZE = 7;
	defparam lut_11240.mask = 128'h0fff0fff7fff7fff0077000070077070;

	lut_sub lut_11253 ({sk[2046], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1447x);
	defparam lut_11253.LUT_SIZE = 7;
	defparam lut_11253.mask = 128'h0fff0fff7fff7fff0033000030077070;

	lut_sub lut_11263 ({sk[2047], i_14_, i_13_, i_12_, i_15_, n_n156}, x19701x);
	defparam lut_11263.LUT_SIZE = 6;
	defparam lut_11263.mask = 64'h7777777701004000;

	lut_sub lut_11266 ({sk[2048], i_14_, i_13_, i_12_, i_15_, n_n156, n_n177}, x19700x);
	defparam lut_11266.LUT_SIZE = 7;
	defparam lut_11266.mask = 128'h0fff0fff7fff7fff0077000070000000;

	lut_sub lut_11273 ({sk[2049], n_n41, n_n40, n_n150, x1447x, x19701x, x19700x}, n_n319);
	defparam lut_11273.LUT_SIZE = 7;
	defparam lut_11273.mask = 128'h0fff0fff7fff7fff00005f5f3fff7fff;

	lut_sub lut_11279 ({sk[2050], i_9_, i_10_, i_11_, i_15_, n_n34, n_n209}, x588x);
	defparam lut_11279.LUT_SIZE = 7;
	defparam lut_11279.mask = 128'h0fff0fff7fff7fff0000000000010000;

	lut_sub lut_11281 ({sk[2051], i_14_, i_13_, i_12_, i_15_, n_n156, n_n191}, x1453x);
	defparam lut_11281.LUT_SIZE = 7;
	defparam lut_11281.mask = 128'h0fff0fff7fff7fff7000070000700007;

	lut_sub lut_11290 ({sk[2052], i_14_, i_13_, i_12_, i_15_, n_n177, n_n191}, x1452x);
	defparam lut_11290.LUT_SIZE = 7;
	defparam lut_11290.mask = 128'h0fff0fff7fff7fff7000070000700003;

	lut_sub lut_11298 ({sk[2053], i_14_, i_13_, i_12_, i_15_, n_n216}, x1454x);
	defparam lut_11298.LUT_SIZE = 6;
	defparam lut_11298.mask = 64'h7777777711015154;

	lut_sub lut_11308 ({sk[2054], i_14_, i_13_, i_12_, i_15_, n_n156}, x1574x);
	defparam lut_11308.LUT_SIZE = 6;
	defparam lut_11308.mask = 64'h7777777740100401;

	lut_sub lut_11313 ({sk[2055], i_14_, i_13_, i_12_, i_15_, n_n191}, x1455x);
	defparam lut_11313.LUT_SIZE = 6;
	defparam lut_11313.mask = 64'h7777777715455555;

	lut_sub lut_11328 ({sk[2056], i_14_, i_13_, i_12_, i_15_, n_n156, n_n177}, x1456x);
	defparam lut_11328.LUT_SIZE = 7;
	defparam lut_11328.mask = 128'h0fff0fff7fff7fff5000070000700007;

	lut_sub lut_11336 ({sk[2057], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1460x);
	defparam lut_11336.LUT_SIZE = 7;
	defparam lut_11336.mask = 128'h0fff0fff7fff7fff0555505557037370;

	lut_sub lut_11352 ({sk[2058], i_14_, i_13_, i_12_, i_15_, n_n177}, x1459x);
	defparam lut_11352.LUT_SIZE = 6;
	defparam lut_11352.mask = 64'h7777777715455154;

	lut_sub lut_11365 ({sk[2059], i_7_, i_5_, i_6_, i_3_, i_4_, n_n19}, x17590x);
	defparam lut_11365.LUT_SIZE = 7;
	defparam lut_11365.mask = 128'h0fff0fff7fff7fff4040505000000000;

	lut_sub lut_11372 ({sk[2060], i_14_, i_13_, i_12_, i_15_, n_n149, n_n177}, x1466x);
	defparam lut_11372.LUT_SIZE = 7;
	defparam lut_11372.mask = 128'h0fff0fff7fff7fff0555505573037370;

	lut_sub lut_11388 ({sk[2061], i_14_, i_13_, i_12_, i_15_, n_n156}, x1465x);
	defparam lut_11388.LUT_SIZE = 6;
	defparam lut_11388.mask = 64'h7777777715455154;

	lut_sub lut_11401 ({sk[2062], i_14_, i_13_, i_12_, i_15_, n_n216}, x197x);
	defparam lut_11401.LUT_SIZE = 6;
	defparam lut_11401.mask = 64'h7777777700010050;

	lut_sub lut_11405 ({sk[2063], i_9_, i_10_, i_11_, x729x, x717x, x721x}, x1467x);
	defparam lut_11405.LUT_SIZE = 7;
	defparam lut_11405.mask = 128'h0fff0fff7fff7fff005555003f000000;

	lut_sub lut_11410 ({sk[2064], i_9_, i_10_, i_11_, i_15_, n_n207, n_n209}, x402x);
	defparam lut_11410.LUT_SIZE = 7;
	defparam lut_11410.mask = 128'h0fff0fff7fff7fff0000000500003000;

	lut_sub lut_11413 ({sk[2065], i_9_, i_10_, i_11_, i_15_, n_n207, n_n209}, x1473x);
	defparam lut_11413.LUT_SIZE = 7;
	defparam lut_11413.mask = 128'h0fff0fff7fff7fff0000000505003005;

	lut_sub lut_11418 ({sk[2066], n_n101, n_n116, n_n108, n_n142, x401x, x1473x}, n_n849);
	defparam lut_11418.LUT_SIZE = 7;
	defparam lut_11418.mask = 128'h0fff0fff7fff7fff003f00ff557fffff;

	lut_sub lut_11424 ({sk[2067], i_14_, i_13_, i_12_, i_15_, n_n216}, x333x);
	defparam lut_11424.LUT_SIZE = 6;
	defparam lut_11424.mask = 64'h7777777701004040;

	lut_sub lut_11428 ({sk[2068], i_14_, i_13_, i_12_, i_15_, n_n216}, x1474x);
	defparam lut_11428.LUT_SIZE = 6;
	defparam lut_11428.mask = 64'h7777777701004144;

	lut_sub lut_11434 ({sk[2069], i_9_, i_10_, i_11_, x728x}, x414x);
	defparam lut_11434.LUT_SIZE = 5;
	defparam lut_11434.mask = 32'h33ff4001;

	lut_sub lut_11437 ({sk[2070], i_9_, i_10_, i_11_, x714x, x17002x, x728x}, x2093x);
	defparam lut_11437.LUT_SIZE = 7;
	defparam lut_11437.mask = 128'h0fff0fff7fff7fff0100000001010001;

	lut_sub lut_11442 ({sk[2071], i_9_, i_10_, i_11_, i_15_, x720x, n_n209}, x19706x);
	defparam lut_11442.LUT_SIZE = 7;
	defparam lut_11442.mask = 128'h0fff0fff7fff7fff0073000000730000;

	lut_sub lut_11447 ({sk[2072], i_14_, i_13_, i_12_, i_15_, n_n177}, x259x);
	defparam lut_11447.LUT_SIZE = 6;
	defparam lut_11447.mask = 64'h7777777700000104;

	lut_sub lut_11450 ({sk[2073], i_9_, i_10_, i_11_, x728x}, x1478x);
	defparam lut_11450.LUT_SIZE = 5;
	defparam lut_11450.mask = 32'h33ff1400;

	lut_sub lut_11453 ({sk[2074], i_7_, i_8_, i_6_, x740x, n_n177, x728x}, x2090x);
	defparam lut_11453.LUT_SIZE = 7;
	defparam lut_11453.mask = 128'h0fff0fff7fff7fff0000000001000000;

	lut_sub lut_11455 ({sk[2075], n_n39, x190x, x244x, x19706x, x1478x, x2090x}, x19709x);
	defparam lut_11455.LUT_SIZE = 7;
	defparam lut_11455.mask = 128'h0fff0fff7fff7fff555577775fff7fff;

	lut_sub lut_11460 ({sk[2076], i_9_, i_10_, i_11_, x740x, n_n200, x728x}, x2092x);
	defparam lut_11460.LUT_SIZE = 7;
	defparam lut_11460.mask = 128'h0fff0fff7fff7fff0100000001000001;

	lut_sub lut_11464 ({sk[2077], n_n38, n_n41, n_n40, n_n54, x161x, x259x}, x21336x);
	defparam lut_11464.LUT_SIZE = 7;
	defparam lut_11464.mask = 128'h0fff0fff7fff7ffffff0f0f088808080;

	lut_sub lut_11469 ({sk[2078], n_n199, x190x, x728x, x2093x, x2092x, x21336x}, x19710x);
	defparam lut_11469.LUT_SIZE = 7;
	defparam lut_11469.mask = 128'h0fff0fff7fff7fffbfbfbfbfbfbfbfff;

	lut_sub lut_11474 ({sk[2079], i_14_, i_13_, i_12_, i_15_, n_n177}, x1484x);
	defparam lut_11474.LUT_SIZE = 6;
	defparam lut_11474.mask = 64'h7777777705004144;

	lut_sub lut_11481 ({sk[2080], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x21339x);
	defparam lut_11481.LUT_SIZE = 7;
	defparam lut_11481.mask = 128'h0fff0fff7fff7fffff8affffaffaafaf;

	lut_sub lut_11492 ({sk[2081], i_14_, i_13_, i_12_, i_15_, n_n199}, x1487x);
	defparam lut_11492.LUT_SIZE = 6;
	defparam lut_11492.mask = 64'h7777777711410050;

	lut_sub lut_11499 ({sk[2082], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1485x);
	defparam lut_11499.LUT_SIZE = 7;
	defparam lut_11499.mask = 128'h0fff0fff7fff7fff0303300700007700;

	lut_sub lut_11509 ({sk[2083], i_14_, i_13_, i_12_, i_15_, n_n156}, x1849x);
	defparam lut_11509.LUT_SIZE = 6;
	defparam lut_11509.mask = 64'h7777777700005154;

	lut_sub lut_11516 ({sk[2084], x735x, n_n126, x86x, x180x, x258x, x108x}, x17114x);
	defparam lut_11516.LUT_SIZE = 7;
	defparam lut_11516.mask = 128'h0fff0fff7fff7fff0000000000007fff;

	lut_sub lut_11521 ({sk[2085], i_14_, i_13_, i_12_, i_15_, n_n199}, x1853x);
	defparam lut_11521.LUT_SIZE = 6;
	defparam lut_11521.mask = 64'h7777777711055154;

	lut_sub lut_11532 ({sk[2086], n_n123, x70x, n_n125, n_n198, x219x, x1853x}, x17115x);
	defparam lut_11532.LUT_SIZE = 7;
	defparam lut_11532.mask = 128'h0fff0fff7fff7fff003f003f557fffff;

	lut_sub lut_11537 ({sk[2087], i_14_, i_13_, i_12_, i_15_, n_n191}, x1857x);
	defparam lut_11537.LUT_SIZE = 6;
	defparam lut_11537.mask = 64'h7777777715450000;

	lut_sub lut_11544 ({sk[2088], i_14_, i_13_, i_12_, i_15_, n_n177}, x1833x);
	defparam lut_11544.LUT_SIZE = 6;
	defparam lut_11544.mask = 64'h7777777715450000;

	lut_sub lut_11551 ({sk[2089], i_14_, i_13_, i_12_, i_15_, n_n191}, x1725x);
	defparam lut_11551.LUT_SIZE = 6;
	defparam lut_11551.mask = 64'h7777777711015154;

	lut_sub lut_11561 ({sk[2090], i_14_, i_13_, i_12_, i_15_, n_n191, n_n216}, x1491x);
	defparam lut_11561.LUT_SIZE = 7;
	defparam lut_11561.mask = 128'h0fff0fff7fff7fff0505000573037370;

	lut_sub lut_11574 ({sk[2091], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1505x);
	defparam lut_11574.LUT_SIZE = 7;
	defparam lut_11574.mask = 128'h0fff0fff7fff7fff0777300330033330;

	lut_sub lut_11588 ({sk[2092], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1504x);
	defparam lut_11588.LUT_SIZE = 7;
	defparam lut_11588.mask = 128'h0fff0fff7fff7fff0333300330053570;

	lut_sub lut_11600 ({sk[2093], i_14_, i_13_, i_12_, i_15_, n_n184}, x314x);
	defparam lut_11600.LUT_SIZE = 6;
	defparam lut_11600.mask = 64'h7777777701004040;

	lut_sub lut_11604 ({sk[2094], i_14_, i_13_, i_12_, i_15_, n_n184}, x338x);
	defparam lut_11604.LUT_SIZE = 6;
	defparam lut_11604.mask = 64'h7777777700000104;

	lut_sub lut_11607 ({sk[2095], i_14_, i_13_, i_12_, i_15_, n_n191}, x1514x);
	defparam lut_11607.LUT_SIZE = 6;
	defparam lut_11607.mask = 64'h7777777705004144;

	lut_sub lut_11614 ({sk[2096], x735x, n_n126, n_n184, x726x, x259x, x1514x}, x1968x);
	defparam lut_11614.LUT_SIZE = 7;
	defparam lut_11614.mask = 128'h0fff0fff7fff7fff000000000000777f;

	lut_sub lut_11618 ({sk[2097], i_14_, i_13_, i_12_, i_15_, n_n184, n_n216}, x21332x);
	defparam lut_11618.LUT_SIZE = 7;
	defparam lut_11618.mask = 128'h0fff0fff7fff7fffff8cffffcffccfcf;

	lut_sub lut_11629 ({sk[2098], n_n123, n_n125, x314x, x338x, x1514x, x21332x}, x19834x);
	defparam lut_11629.LUT_SIZE = 7;
	defparam lut_11629.mask = 128'h0fff0fff7fff7fff00000fffbbbbbfff;

	lut_sub lut_11634 ({sk[2099], i_14_, i_13_, i_12_, i_15_, n_n216}, x1518x);
	defparam lut_11634.LUT_SIZE = 6;
	defparam lut_11634.mask = 64'h7777777740100401;

	lut_sub lut_11639 ({sk[2100], i_14_, i_13_, i_12_, i_15_, n_n191}, x1519x);
	defparam lut_11639.LUT_SIZE = 6;
	defparam lut_11639.mask = 64'h7777777755554440;

	lut_sub lut_11651 ({sk[2101], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1521x);
	defparam lut_11651.LUT_SIZE = 7;
	defparam lut_11651.mask = 128'h0fff0fff7fff7fff0333303375057570;

	lut_sub lut_11667 ({sk[2102], i_14_, i_13_, i_12_, i_15_, n_n184}, x1520x);
	defparam lut_11667.LUT_SIZE = 6;
	defparam lut_11667.mask = 64'h7777777715455154;

	lut_sub lut_11680 ({sk[2103], x370x, x404x, x717x, n_n2, x707x, n_n191}, x18368x);
	defparam lut_11680.LUT_SIZE = 7;
	defparam lut_11680.mask = 128'h0fff0fff7fff7fff33373f3f3f3f3f3f;

	lut_sub lut_11685 ({sk[2104], i_14_, i_13_, i_12_, i_15_, n_n191}, x1535x);
	defparam lut_11685.LUT_SIZE = 6;
	defparam lut_11685.mask = 64'h7777777701014054;

	lut_sub lut_11692 ({sk[2105], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1537x);
	defparam lut_11692.LUT_SIZE = 7;
	defparam lut_11692.mask = 128'h0fff0fff7fff7fff5700000000570000;

	lut_sub lut_11697 ({sk[2106], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1536x);
	defparam lut_11697.LUT_SIZE = 7;
	defparam lut_11697.mask = 128'h0fff0fff7fff7fff0357000057000000;

	lut_sub lut_11703 ({sk[2107], i_14_, i_13_, i_12_, i_15_, n_n156, n_n184}, x19444x);
	defparam lut_11703.LUT_SIZE = 7;
	defparam lut_11703.mask = 128'h0fff0fff7fff7fff0000300330503000;

	lut_sub lut_11709 ({sk[2108], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1538x);
	defparam lut_11709.LUT_SIZE = 7;
	defparam lut_11709.mask = 128'h0fff0fff7fff7fff0000005757000057;

	lut_sub lut_11716 ({sk[2109], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x19443x);
	defparam lut_11716.LUT_SIZE = 7;
	defparam lut_11716.mask = 128'h0fff0fff7fff7fff0000005700000057;

	lut_sub lut_11721 ({sk[2110], i_14_, i_13_, i_12_, i_15_, n_n191}, x348x);
	defparam lut_11721.LUT_SIZE = 6;
	defparam lut_11721.mask = 64'h7777777705000000;

	lut_sub lut_11724 ({sk[2111], x137x, n_n36, n_n34, x63x, x348x}, x19721x);
	defparam lut_11724.LUT_SIZE = 6;
	defparam lut_11724.mask = 64'h77777777037703ff;

	lut_sub lut_11729 ({sk[2112], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1542x);
	defparam lut_11729.LUT_SIZE = 7;
	defparam lut_11729.mask = 128'h0fff0fff7fff7fff0077000030033030;

	lut_sub lut_11738 ({sk[2113], i_14_, i_13_, i_12_, i_15_, n_n149, n_n177}, x1541x);
	defparam lut_11738.LUT_SIZE = 7;
	defparam lut_11738.mask = 128'h0fff0fff7fff7fff0055000000030000;

	lut_sub lut_11742 ({sk[2114], x137x, n_n36, n_n34, n_n176, x126x, x1541x}, x19732x);
	defparam lut_11742.LUT_SIZE = 7;
	defparam lut_11742.mask = 128'h0fff0fff7fff7fff005f337f00ff33ff;

	lut_sub lut_11747 ({sk[2115], i_14_, i_13_, i_12_, i_15_, n_n34, n_n170}, x21408x);
	defparam lut_11747.LUT_SIZE = 7;
	defparam lut_11747.mask = 128'h0fff0fff7fff7fffffeeffffeffeefef;

	lut_sub lut_11755 ({sk[2116], n_n36, x934x, x1542x, x21408x}, x19733x);
	defparam lut_11755.LUT_SIZE = 5;
	defparam lut_11755.mask = 32'h33ffaabf;

	lut_sub lut_11759 ({sk[2117], n_n36, n_n34, x720x, n_n199, x68x, x385x}, x19736x);
	defparam lut_11759.LUT_SIZE = 7;
	defparam lut_11759.mask = 128'h0fff0fff7fff7fff00007777333f777f;

	lut_sub lut_11764 ({sk[2118], n_n36, n_n34, n_n183, n_n176, x128x, x348x}, x19720x);
	defparam lut_11764.LUT_SIZE = 7;
	defparam lut_11764.mask = 128'h0fff0fff7fff7fff000077ff0f0f7fff;

	lut_sub lut_11769 ({sk[2119], x714x, x17002x, x278x, x275x, x332x, x19742x}, x2051x);
	defparam lut_11769.LUT_SIZE = 7;
	defparam lut_11769.mask = 128'h0fff0fff7fff7fff0000000000007fff;

	lut_sub lut_11774 ({sk[2120], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1619x);
	defparam lut_11774.LUT_SIZE = 7;
	defparam lut_11774.mask = 128'h0fff0fff7fff7fff0055000050077070;

	lut_sub lut_11784 ({sk[2121], i_14_, i_13_, i_12_, i_15_, n_n191}, x19755x);
	defparam lut_11784.LUT_SIZE = 6;
	defparam lut_11784.mask = 64'h7777777705004144;

	lut_sub lut_11791 ({sk[2122], i_14_, i_13_, i_12_, i_15_, n_n184, n_n216}, x1684x);
	defparam lut_11791.LUT_SIZE = 7;
	defparam lut_11791.mask = 128'h0fff0fff7fff7fff0037000070077070;

	lut_sub lut_11803 ({sk[2123], i_8_, x734x, n_n18, x63x, x348x, x19749x}, x19751x);
	defparam lut_11803.LUT_SIZE = 7;
	defparam lut_11803.mask = 128'h0fff0fff7fff7fff5555557f55555555;

	lut_sub lut_11807 ({sk[2124], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1617x);
	defparam lut_11807.LUT_SIZE = 7;
	defparam lut_11807.mask = 128'h0fff0fff7fff7fff0057000070077070;

	lut_sub lut_11819 ({sk[2125], n_n184, n_n42, n_n43, n_n191, x728x, x19748x}, n_n388);
	defparam lut_11819.LUT_SIZE = 7;
	defparam lut_11819.mask = 128'h0fff0fff7fff7fff5555575755777777;

	lut_sub lut_11824 ({sk[2126], x740x, n_n200, x714x, x17002x, x296x, x332x}, x19750x);
	defparam lut_11824.LUT_SIZE = 7;
	defparam lut_11824.mask = 128'h0fff0fff7fff7fff0003000300037777;

	lut_sub lut_11828 ({sk[2127], x734x, n_n161, n_n43, n_n183, x128x, x346x}, n_n390);
	defparam lut_11828.LUT_SIZE = 7;
	defparam lut_11828.mask = 128'h0fff0fff7fff7fff003f003f003f777f;

	lut_sub lut_11833 ({sk[2128], x740x, x140x, n_n161, x244x, x414x, x1638x}, x2017x);
	defparam lut_11833.LUT_SIZE = 7;
	defparam lut_11833.mask = 128'h0fff0fff7fff7fff00000000007f00ff;

	lut_sub lut_11838 ({sk[2129], n_n46, n_n47, n_n199, x728x, x1638x, x19796x}, x19799x);
	defparam lut_11838.LUT_SIZE = 7;
	defparam lut_11838.mask = 128'h0fff0fff7fff7fff0000777f000f777f;

	lut_sub lut_11843 ({sk[2130], n_n162, n_n18, x714x, x63x, x348x, x19805x}, x19807x);
	defparam lut_11843.LUT_SIZE = 7;
	defparam lut_11843.mask = 128'h0fff0fff7fff7fff555555555555557f;

	lut_sub lut_11847 ({sk[2131], x435x, x603x, n_n52, x189x, n_n56, x697x}, x19806x);
	defparam lut_11847.LUT_SIZE = 7;
	defparam lut_11847.mask = 128'h0fff0fff7fff7fff575fffffffffffff;

	lut_sub lut_11853 ({sk[2132], n_n46, n_n47, x325x, x19810x, x354x, x19809x}, x19811x);
	defparam lut_11853.LUT_SIZE = 7;
	defparam lut_11853.mask = 128'h0fff0fff7fff7fff00007f7f77ff7fff;

	lut_sub lut_11860 ({sk[2133], n_n123, n_n125, x1665x, x1664x, x1761x, x1760x}, x19859x);
	defparam lut_11860.LUT_SIZE = 7;
	defparam lut_11860.mask = 128'h0fff0fff7fff7fff000033ff5f5f7fff;

	lut_sub lut_11865 ({sk[2134], x734x, n_n126, n_n113, x335x, x333x, x1719x}, x19846x);
	defparam lut_11865.LUT_SIZE = 7;
	defparam lut_11865.mask = 128'h0fff0fff7fff7fff0055005500553f7f;

	lut_sub lut_11869 ({sk[2135], n_n184, x720x, n_n113, x1957x, x21334x, x21450x}, x19847x);
	defparam lut_11869.LUT_SIZE = 7;
	defparam lut_11869.mask = 128'h0fff0fff7fff7fffefefefefefefefff;

	lut_sub lut_11874 ({sk[2136], n_n123, n_n125, x207x, n_n136, x416x, x19848x}, x19854x);
	defparam lut_11874.LUT_SIZE = 7;
	defparam lut_11874.mask = 128'h0fff0fff7fff7fff00007fff0f0f7fff;

	lut_sub lut_11880 ({sk[2137], n_n123, n_n125, n_n143, x249x, x19853x, x21333x}, x19855x);
	defparam lut_11880.LUT_SIZE = 7;
	defparam lut_11880.mask = 128'h0fff0fff7fff7fff00000fffbbbbbfff;

	lut_sub lut_11885 ({sk[2138], i_7_, i_8_, i_6_, x735x, x129x}, x3945x);
	defparam lut_11885.LUT_SIZE = 6;
	defparam lut_11885.mask = 64'h7777777710000000;

	lut_sub lut_11887 ({sk[2139], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x18198x);
	defparam lut_11887.LUT_SIZE = 7;
	defparam lut_11887.mask = 128'h0fff0fff7fff7fff3000030000300007;

	lut_sub lut_11893 ({sk[2140], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x18199x);
	defparam lut_11893.LUT_SIZE = 7;
	defparam lut_11893.mask = 128'h0fff0fff7fff7fff7000070000700005;

	lut_sub lut_11901 ({sk[2141], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1546x);
	defparam lut_11901.LUT_SIZE = 7;
	defparam lut_11901.mask = 128'h0fff0fff7fff7fff7000070000700007;

	lut_sub lut_11910 ({sk[2142], i_14_, i_13_, i_12_, i_15_, n_n216}, x261x);
	defparam lut_11910.LUT_SIZE = 6;
	defparam lut_11910.mask = 64'h7777777701010040;

	lut_sub lut_11914 ({sk[2143], i_14_, i_13_, i_12_, i_15_, n_n216}, x375x);
	defparam lut_11914.LUT_SIZE = 6;
	defparam lut_11914.mask = 64'h7777777710400000;

	lut_sub lut_11917 ({sk[2144], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1555x);
	defparam lut_11917.LUT_SIZE = 7;
	defparam lut_11917.mask = 128'h0fff0fff7fff7fff0057000057550000;

	lut_sub lut_11923 ({sk[2145], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1563x);
	defparam lut_11923.LUT_SIZE = 7;
	defparam lut_11923.mask = 128'h0fff0fff7fff7fff5700000057550000;

	lut_sub lut_11929 ({sk[2146], i_14_, i_13_, i_12_, i_15_, n_n184}, x269x);
	defparam lut_11929.LUT_SIZE = 6;
	defparam lut_11929.mask = 64'h7777777700000144;

	lut_sub lut_11933 ({sk[2147], i_14_, i_13_, i_12_, i_15_, n_n184}, x275x);
	defparam lut_11933.LUT_SIZE = 6;
	defparam lut_11933.mask = 64'h7777777705004000;

	lut_sub lut_11937 ({sk[2148], i_14_, i_13_, i_12_, i_15_, n_n170}, x282x);
	defparam lut_11937.LUT_SIZE = 6;
	defparam lut_11937.mask = 64'h7777777705004000;

	lut_sub lut_11941 ({sk[2149], i_14_, i_13_, i_12_, i_15_, n_n170}, x283x);
	defparam lut_11941.LUT_SIZE = 6;
	defparam lut_11941.mask = 64'h7777777700000144;

	lut_sub lut_11945 ({sk[2150], i_9_, i_10_, i_11_, n_n36, n_n34, x728x}, x21341x);
	defparam lut_11945.LUT_SIZE = 7;
	defparam lut_11945.mask = 128'h0fff0fff7fff7fff0000150000111500;

	lut_sub lut_11951 ({sk[2151], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1568x);
	defparam lut_11951.LUT_SIZE = 7;
	defparam lut_11951.mask = 128'h0fff0fff7fff7fff0077000070037030;

	lut_sub lut_11962 ({sk[2152], i_14_, i_13_, i_12_, i_15_, n_n149}, x1780x);
	defparam lut_11962.LUT_SIZE = 6;
	defparam lut_11962.mask = 64'h7777777705000000;

	lut_sub lut_11965 ({sk[2153], i_14_, i_13_, i_12_, i_15_, n_n199}, x19319x);
	defparam lut_11965.LUT_SIZE = 6;
	defparam lut_11965.mask = 64'h7777777715400000;

	lut_sub lut_11970 ({sk[2154], i_9_, i_10_, i_11_, x721x, x728x, x727x}, x19115x);
	defparam lut_11970.LUT_SIZE = 7;
	defparam lut_11970.mask = 128'h0fff0fff7fff7fff000000003300553f;

	lut_sub lut_11975 ({sk[2155], i_14_, i_13_, i_12_, i_15_, n_n156, n_n184}, x19116x);
	defparam lut_11975.LUT_SIZE = 7;
	defparam lut_11975.mask = 128'h0fff0fff7fff7fff0003050330503300;

	lut_sub lut_11983 ({sk[2156], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1585x);
	defparam lut_11983.LUT_SIZE = 7;
	defparam lut_11983.mask = 128'h0fff0fff7fff7fff0057570000005700;

	lut_sub lut_11990 ({sk[2157], i_9_, i_10_, i_11_, i_15_, n_n201, x728x}, x1584x);
	defparam lut_11990.LUT_SIZE = 7;
	defparam lut_11990.mask = 128'h0fff0fff7fff7fff0000570000575700;

	lut_sub lut_11997 ({sk[2158], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1587x);
	defparam lut_11997.LUT_SIZE = 7;
	defparam lut_11997.mask = 128'h0fff0fff7fff7fff0037000070077070;

	lut_sub lut_12009 ({sk[2159], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1586x);
	defparam lut_12009.LUT_SIZE = 7;
	defparam lut_12009.mask = 128'h0fff0fff7fff7fff0073000030033030;

	lut_sub lut_12017 ({sk[2160], n_n125, x188x, n_n52, x1474x, x1586x, x1973x}, x19837x);
	defparam lut_12017.LUT_SIZE = 7;
	defparam lut_12017.mask = 128'h0fff0fff7fff7fff555555ff7f7f7fff;

	lut_sub lut_12022 ({sk[2161], n_n124, x735x, x188x, n_n56, n_n433, x1587x}, x21331x);
	defparam lut_12022.LUT_SIZE = 7;
	defparam lut_12022.mask = 128'h0fff0fff7fff7fffccc0ccc0ccc08880;

	lut_sub lut_12029 ({sk[2162], i_14_, i_13_, i_12_, i_15_, n_n184, n_n216}, x1590x);
	defparam lut_12029.LUT_SIZE = 7;
	defparam lut_12029.mask = 128'h0fff0fff7fff7fff0077000070037030;

	lut_sub lut_12040 ({sk[2163], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1589x);
	defparam lut_12040.LUT_SIZE = 7;
	defparam lut_12040.mask = 128'h0fff0fff7fff7fff0055000050075070;

	lut_sub lut_12049 ({sk[2164], i_14_, i_13_, i_12_, i_15_, n_n184}, x1722x);
	defparam lut_12049.LUT_SIZE = 6;
	defparam lut_12049.mask = 64'h7777777705004040;

	lut_sub lut_12054 ({sk[2165], i_14_, i_13_, i_12_, i_15_, n_n191}, x1721x);
	defparam lut_12054.LUT_SIZE = 6;
	defparam lut_12054.mask = 64'h7777777701004144;

	lut_sub lut_12060 ({sk[2166], i_14_, i_13_, i_12_, i_15_, n_n149}, x1593x);
	defparam lut_12060.LUT_SIZE = 6;
	defparam lut_12060.mask = 64'h7777777705004144;

	lut_sub lut_12067 ({sk[2167], i_9_, i_10_, i_11_, x740x, n_n126, x728x}, x434x);
	defparam lut_12067.LUT_SIZE = 7;
	defparam lut_12067.mask = 128'h0fff0fff7fff7fff0000010000000100;

	lut_sub lut_12070 ({sk[2168], i_15_, x740x, n_n126, n_n170, n_n209}, x522x);
	defparam lut_12070.LUT_SIZE = 6;
	defparam lut_12070.mask = 64'h7777777700000001;

	lut_sub lut_12072 ({sk[2169], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x18083x);
	defparam lut_12072.LUT_SIZE = 7;
	defparam lut_12072.mask = 128'h0fff0fff7fff7fff7000070000700007;

	lut_sub lut_12081 ({sk[2170], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x353x);
	defparam lut_12081.LUT_SIZE = 7;
	defparam lut_12081.mask = 128'h0fff0fff7fff7fff3000030000000005;

	lut_sub lut_12085 ({sk[2171], i_9_, i_10_, i_11_, x725x, x719x, x728x}, x355x);
	defparam lut_12085.LUT_SIZE = 7;
	defparam lut_12085.mask = 128'h0fff0fff7fff7fff0f00000000770000;

	lut_sub lut_12089 ({sk[2172], n_n212, x150x, x217x, x18083x, x353x, x355x}, x3676x);
	defparam lut_12089.LUT_SIZE = 7;
	defparam lut_12089.mask = 128'h0fff0fff7fff7fff000000007fffffff;

	lut_sub lut_12095 ({sk[2173], x735x, n_n126, x720x, x1818x, n_n216}, x18085x);
	defparam lut_12095.LUT_SIZE = 6;
	defparam lut_12095.mask = 64'h7777777700000037;

	lut_sub lut_12098 ({sk[2174], i_14_, i_13_, i_12_, i_15_, n_n191, n_n199}, x350x);
	defparam lut_12098.LUT_SIZE = 7;
	defparam lut_12098.mask = 128'h0fff0fff7fff7fff5000050000000003;

	lut_sub lut_12102 ({sk[2175], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x356x);
	defparam lut_12102.LUT_SIZE = 7;
	defparam lut_12102.mask = 128'h0fff0fff7fff7fff5000000000300003;

	lut_sub lut_12106 ({sk[2176], n_n212, x172x, x133x, x127x, x350x, x356x}, x3671x);
	defparam lut_12106.LUT_SIZE = 7;
	defparam lut_12106.mask = 128'h0fff0fff7fff7fff000000007fffffff;

	lut_sub lut_12112 ({sk[2177], n_n212, x125x, x55x, x158x, x176x}, x18091x);
	defparam lut_12112.LUT_SIZE = 6;
	defparam lut_12112.mask = 64'h7777777700007fff;

	lut_sub lut_12117 ({sk[2178], i_14_, i_13_, i_12_, i_15_, n_n199}, x1837x);
	defparam lut_12117.LUT_SIZE = 6;
	defparam lut_12117.mask = 64'h7777777711054040;

	lut_sub lut_12124 ({sk[2179], i_14_, i_13_, i_12_, i_15_, n_n216}, x1838x);
	defparam lut_12124.LUT_SIZE = 6;
	defparam lut_12124.mask = 64'h7777777715440000;

	lut_sub lut_12130 ({sk[2180], i_14_, i_13_, i_12_, i_15_, n_n191, n_n199}, x18093x);
	defparam lut_12130.LUT_SIZE = 7;
	defparam lut_12130.mask = 128'h0fff0fff7fff7fff0050500000070000;

	lut_sub lut_12135 ({sk[2181], n_n125, x219x, x1596x, x1837x, x1838x, x18093x}, x18096x);
	defparam lut_12135.LUT_SIZE = 7;
	defparam lut_12135.mask = 128'h0fff0fff7fff7fff000000007fffffff;

	lut_sub lut_12141 ({sk[2182], i_14_, i_13_, i_12_, i_15_, n_n149, n_n170}, x17918x);
	defparam lut_12141.LUT_SIZE = 7;
	defparam lut_12141.mask = 128'h0fff0fff7fff7fff7000070000700000;

	lut_sub lut_12148 ({sk[2183], i_15_, n_n191, n_n209, x153x, x217x, x17918x}, x17922x);
	defparam lut_12148.LUT_SIZE = 7;
	defparam lut_12148.mask = 128'h0fff0fff7fff7fff7f7f7f7f7f7f7fff;

	lut_sub lut_12153 ({sk[2184], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x17917x);
	defparam lut_12153.LUT_SIZE = 7;
	defparam lut_12153.mask = 128'h0fff0fff7fff7fff5000050000500007;

	lut_sub lut_12159 ({sk[2185], x719x, x78x, n_n170, x356x, x355x, x17917x}, x17923x);
	defparam lut_12159.LUT_SIZE = 7;
	defparam lut_12159.mask = 128'h0fff0fff7fff7fff7f7fffff7fffffff;

	lut_sub lut_12165 ({sk[2186], i_14_, i_13_, i_12_, i_15_, n_n184}, x1732x);
	defparam lut_12165.LUT_SIZE = 6;
	defparam lut_12165.mask = 64'h7777777711015154;

	lut_sub lut_12175 ({sk[2187], i_14_, i_13_, i_12_, i_15_, n_n184}, x1602x);
	defparam lut_12175.LUT_SIZE = 6;
	defparam lut_12175.mask = 64'h7777777715455154;

	lut_sub lut_12188 ({sk[2188], i_7_, i_8_, i_6_, x735x, x131x}, x4968x);
	defparam lut_12188.LUT_SIZE = 6;
	defparam lut_12188.mask = 64'h7777777710000000;

	lut_sub lut_12190 ({sk[2189], i_14_, i_13_, i_12_, i_15_, n_n170}, x17871x);
	defparam lut_12190.LUT_SIZE = 6;
	defparam lut_12190.mask = 64'h7777777704441110;

	lut_sub lut_12197 ({sk[2190], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1605x);
	defparam lut_12197.LUT_SIZE = 7;
	defparam lut_12197.mask = 128'h0fff0fff7fff7fff0000007707030770;

	lut_sub lut_12209 ({sk[2191], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1604x);
	defparam lut_12209.LUT_SIZE = 7;
	defparam lut_12209.mask = 128'h0fff0fff7fff7fff0000003303050330;

	lut_sub lut_12216 ({sk[2192], n_n36, n_n34, n_n176, x100x, x1298x, x1605x}, x19527x);
	defparam lut_12216.LUT_SIZE = 7;
	defparam lut_12216.mask = 128'h0fff0fff7fff7fff000033335fff7fff;

	lut_sub lut_12221 ({sk[2193], i_14_, i_13_, i_12_, i_15_, n_n170}, x1608x);
	defparam lut_12221.LUT_SIZE = 6;
	defparam lut_12221.mask = 64'h7777777700051114;

	lut_sub lut_12228 ({sk[2194], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1607x);
	defparam lut_12228.LUT_SIZE = 7;
	defparam lut_12228.mask = 128'h0fff0fff7fff7fff0000007705050550;

	lut_sub lut_12237 ({sk[2195], n_n36, n_n34, x100x, x1608x, x1607x}, x19533x);
	defparam lut_12237.LUT_SIZE = 6;
	defparam lut_12237.mask = 64'h77777777003f557f;

	lut_sub lut_12241 ({sk[2196], i_14_, i_13_, i_12_, i_15_, n_n216}, x1609x);
	defparam lut_12241.LUT_SIZE = 6;
	defparam lut_12241.mask = 64'h7777777700051114;

	lut_sub lut_12248 ({sk[2197], n_n36, n_n34, n_n183, n_n176, x1770x, x1769x}, x21453x);
	defparam lut_12248.LUT_SIZE = 7;
	defparam lut_12248.mask = 128'h0fff0fff7fff7fffffffa000cccc8000;

	lut_sub lut_12253 ({sk[2198], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1611x);
	defparam lut_12253.LUT_SIZE = 7;
	defparam lut_12253.mask = 128'h0fff0fff7fff7fff0037000070077070;

	lut_sub lut_12265 ({sk[2199], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x21330x);
	defparam lut_12265.LUT_SIZE = 7;
	defparam lut_12265.mask = 128'h0fff0fff7fff7fffff88ffff8ff88f8f;

	lut_sub lut_12272 ({sk[2200], n_n101, n_n108, n_n178, x314x, x1611x, x21330x}, n_n330);
	defparam lut_12272.LUT_SIZE = 7;
	defparam lut_12272.mask = 128'h0fff0fff7fff7fff0000aaaa3fffbfff;

	lut_sub lut_12277 ({sk[2201], i_14_, i_13_, i_12_, i_15_, n_n199}, x1614x);
	defparam lut_12277.LUT_SIZE = 6;
	defparam lut_12277.mask = 64'h7777777705004144;

	lut_sub lut_12284 ({sk[2202], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1613x);
	defparam lut_12284.LUT_SIZE = 7;
	defparam lut_12284.mask = 128'h0fff0fff7fff7fff0037000070077070;

	lut_sub lut_12296 ({sk[2203], i_9_, i_10_, i_11_, x726x, x1614x}, x1612x);
	defparam lut_12296.LUT_SIZE = 6;
	defparam lut_12296.mask = 64'h7777777755555557;

	lut_sub lut_12299 ({sk[2204], i_14_, i_13_, i_12_, i_15_, n_n191}, x1681x);
	defparam lut_12299.LUT_SIZE = 6;
	defparam lut_12299.mask = 64'h7777777705004144;

	lut_sub lut_12306 ({sk[2205], i_9_, i_10_, i_11_, x720x, x726x, x727x}, x1680x);
	defparam lut_12306.LUT_SIZE = 7;
	defparam lut_12306.mask = 128'h0fff0fff7fff7fff5f00000000000033;

	lut_sub lut_12310 ({sk[2206], n_n101, n_n108, x1613x, x1612x, x1681x, x1680x}, n_n331);
	defparam lut_12310.LUT_SIZE = 7;
	defparam lut_12310.mask = 128'h0fff0fff7fff7fff00003f3f55ff7fff;

	lut_sub lut_12315 ({sk[2207], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1616x);
	defparam lut_12315.LUT_SIZE = 7;
	defparam lut_12315.mask = 128'h0fff0fff7fff7fff0057000070077070;

	lut_sub lut_12327 ({sk[2208], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1615x);
	defparam lut_12327.LUT_SIZE = 7;
	defparam lut_12327.mask = 128'h0fff0fff7fff7fff0073000030033030;

	lut_sub lut_12335 ({sk[2209], n_n101, n_n108, x1412x, x1411x, x1616x, x1615x}, x19776x);
	defparam lut_12335.LUT_SIZE = 7;
	defparam lut_12335.mask = 128'h0fff0fff7fff7fff00003f3f55ff7fff;

	lut_sub lut_12340 ({sk[2210], i_14_, i_13_, i_12_, i_15_, n_n199}, x332x);
	defparam lut_12340.LUT_SIZE = 6;
	defparam lut_12340.mask = 64'h7777777705004000;

	lut_sub lut_12344 ({sk[2211], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x19742x);
	defparam lut_12344.LUT_SIZE = 7;
	defparam lut_12344.mask = 128'h0fff0fff7fff7fff0000000000077070;

	lut_sub lut_12351 ({sk[2212], n_n42, n_n43, n_n191, x720x, x728x, x346x}, x19749x);
	defparam lut_12351.LUT_SIZE = 7;
	defparam lut_12351.mask = 128'h0fff0fff7fff7fff00005577000f557f;

	lut_sub lut_12355 ({sk[2213], n_n47, x149x, x147x, x1886x, x1458x, x1893x}, n_n3485);
	defparam lut_12355.LUT_SIZE = 7;
	defparam lut_12355.mask = 128'h0fff0fff7fff7fff000000007fffffff;

	lut_sub lut_12361 ({sk[2214], n_n39, n_n150, x207x, n_n78, x248x, x110x}, n_n3532);
	defparam lut_12361.LUT_SIZE = 7;
	defparam lut_12361.mask = 128'h0fff0fff7fff7fff000000007fffffff;

	lut_sub lut_12367 ({sk[2215], i_14_, i_13_, i_12_, i_15_, n_n149, n_n184}, x18105x);
	defparam lut_12367.LUT_SIZE = 7;
	defparam lut_12367.mask = 128'h0fff0fff7fff7fff5333353330503005;

	lut_sub lut_12380 ({sk[2216], i_14_, i_13_, i_12_, i_15_, n_n191}, x18100x);
	defparam lut_12380.LUT_SIZE = 6;
	defparam lut_12380.mask = 64'h7777777740100401;

	lut_sub lut_12385 ({sk[2217], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x18101x);
	defparam lut_12385.LUT_SIZE = 7;
	defparam lut_12385.mask = 128'h0fff0fff7fff7fff3000030000300007;

	lut_sub lut_12391 ({sk[2218], n_n125, x141x, n_n4657, x18105x, x18100x, x18101x}, n_n3494);
	defparam lut_12391.LUT_SIZE = 7;
	defparam lut_12391.mask = 128'h0fff0fff7fff7fff00ff00ff7fffffff;

	lut_sub lut_12397 ({sk[2219], i_14_, i_13_, i_12_, i_15_, n_n184}, x18110x);
	defparam lut_12397.LUT_SIZE = 6;
	defparam lut_12397.mask = 64'h7777777711054040;

	lut_sub lut_12404 ({sk[2220], i_9_, i_10_, i_11_, x720x, x107x}, x18109x);
	defparam lut_12404.LUT_SIZE = 6;
	defparam lut_12404.mask = 64'h7777777777555555;

	lut_sub lut_12408 ({sk[2221], x735x, n_n126, x62x, n_n176, x18110x, x18109x}, x3658x);
	defparam lut_12408.LUT_SIZE = 7;
	defparam lut_12408.mask = 128'h0fff0fff7fff7fff0000000000007fff;

	lut_sub lut_12413 ({sk[2222], x735x, n_n126, x51x, x100x, x1817x}, x18113x);
	defparam lut_12413.LUT_SIZE = 6;
	defparam lut_12413.mask = 64'h777777770000007f;

	lut_sub lut_12417 ({sk[2223], i_14_, i_13_, i_12_, i_15_, n_n170}, x1901x);
	defparam lut_12417.LUT_SIZE = 6;
	defparam lut_12417.mask = 64'h7777777700015054;

	lut_sub lut_12424 ({sk[2224], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x18116x);
	defparam lut_12424.LUT_SIZE = 7;
	defparam lut_12424.mask = 128'h0fff0fff7fff7fff0505005003000330;

	lut_sub lut_12431 ({sk[2225], n_n148, x90x, n_n125, x69x, x225x, x18116x}, x3653x);
	defparam lut_12431.LUT_SIZE = 7;
	defparam lut_12431.mask = 128'h0fff0fff7fff7fff007f00ff00ff00ff;

	lut_sub lut_12437 ({sk[2226], x735x, n_n126, x155x, x208x, x148x, x1830x}, x18118x);
	defparam lut_12437.LUT_SIZE = 7;
	defparam lut_12437.mask = 128'h0fff0fff7fff7fff0000000000007fff;

	lut_sub lut_12442 ({sk[2227], i_14_, i_13_, i_12_, i_15_, n_n149}, x1624x);
	defparam lut_12442.LUT_SIZE = 6;
	defparam lut_12442.mask = 64'h7777777711015154;

	lut_sub lut_12452 ({sk[2228], i_14_, i_13_, i_12_, i_15_, n_n184}, x1625x);
	defparam lut_12452.LUT_SIZE = 6;
	defparam lut_12452.mask = 64'h7777777715455154;

	lut_sub lut_12465 ({sk[2229], i_14_, i_13_, i_12_, i_15_, n_n170}, x1856x);
	defparam lut_12465.LUT_SIZE = 6;
	defparam lut_12465.mask = 64'h7777777711014044;

	lut_sub lut_12472 ({sk[2230], i_14_, i_13_, i_12_, i_15_, n_n184}, x1882x);
	defparam lut_12472.LUT_SIZE = 6;
	defparam lut_12472.mask = 64'h7777777700005154;

	lut_sub lut_12479 ({sk[2231], i_14_, i_13_, i_12_, i_15_, n_n184}, x1627x);
	defparam lut_12479.LUT_SIZE = 6;
	defparam lut_12479.mask = 64'h7777777715455154;

	lut_sub lut_12492 ({sk[2232], i_14_, i_13_, i_12_, i_15_, n_n191, n_n199}, x19565x);
	defparam lut_12492.LUT_SIZE = 7;
	defparam lut_12492.mask = 128'h0fff0fff7fff7fff0000007703030370;

	lut_sub lut_12502 ({sk[2233], i_14_, i_13_, i_12_, i_15_, n_n184, n_n216}, x1628x);
	defparam lut_12502.LUT_SIZE = 7;
	defparam lut_12502.mask = 128'h0fff0fff7fff7fff0000007707070770;

	lut_sub lut_12515 ({sk[2234], n_n41, n_n40, x124x, x165x, x19565x, x1628x}, n_n767);
	defparam lut_12515.LUT_SIZE = 7;
	defparam lut_12515.mask = 128'h0fff0fff7fff7fff000055553fff7fff;

	lut_sub lut_12520 ({sk[2235], i_14_, i_13_, i_12_, i_15_, n_n170}, x1881x);
	defparam lut_12520.LUT_SIZE = 6;
	defparam lut_12520.mask = 64'h7777777700011114;

	lut_sub lut_12526 ({sk[2236], i_9_, i_10_, i_11_, i_15_, n_n41, n_n209}, x2257x);
	defparam lut_12526.LUT_SIZE = 7;
	defparam lut_12526.mask = 128'h0fff0fff7fff7fff0100000001010000;

	lut_sub lut_12530 ({sk[2237], i_9_, i_10_, i_11_, n_n41, n_n40, x719x}, x21345x);
	defparam lut_12530.LUT_SIZE = 7;
	defparam lut_12530.mask = 128'h0fff0fff7fff7fffeeffffeaffffffee;

	lut_sub lut_12540 ({sk[2238], n_n38, n_n39, n_n84, x1881x, x2257x, x21345x}, x19549x);
	defparam lut_12540.LUT_SIZE = 7;
	defparam lut_12540.mask = 128'h0fff0fff7fff7fffbbbbbbffbfbfbfff;

	lut_sub lut_12545 ({sk[2239], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1632x);
	defparam lut_12545.LUT_SIZE = 7;
	defparam lut_12545.mask = 128'h0fff0fff7fff7fff0000007707070770;

	lut_sub lut_12558 ({sk[2240], i_7_, i_8_, i_6_, x740x, n_n6642, n_n132}, x635x);
	defparam lut_12558.LUT_SIZE = 7;
	defparam lut_12558.mask = 128'h0fff0fff7fff7fff3337333333333333;

	lut_sub lut_12561 ({sk[2241], n_n39, x393x, n_n148, n_n69, x647x, x635x}, x19556x);
	defparam lut_12561.LUT_SIZE = 7;
	defparam lut_12561.mask = 128'h0fff0fff7fff7fff7777ffff7fffffff;

	lut_sub lut_12567 ({sk[2242], n_n38, n_n969, x207x, n_n84, x279x, x572x}, x19557x);
	defparam lut_12567.LUT_SIZE = 7;
	defparam lut_12567.mask = 128'h0fff0fff7fff7fff5555ffff7fffffff;

	lut_sub lut_12573 ({sk[2243], n_n156, n_n41, x719x, n_n216, x503x, x19543x}, x21412x);
	defparam lut_12573.LUT_SIZE = 7;
	defparam lut_12573.mask = 128'h0fff0fff7fff7fff8888888088888800;

	lut_sub lut_12577 ({sk[2244], n_n39, n_n41, n_n40, x279x, x280x, x1632x}, x21414x);
	defparam lut_12577.LUT_SIZE = 7;
	defparam lut_12577.mask = 128'h0fff0fff7fff7fffff88aa88f080a080;

	lut_sub lut_12584 ({sk[2245], i_14_, i_13_, i_12_, i_15_, n_n149, n_n191}, x1638x);
	defparam lut_12584.LUT_SIZE = 7;
	defparam lut_12584.mask = 128'h0fff0fff7fff7fff0033000030533030;

	lut_sub lut_12592 ({sk[2246], i_9_, i_10_, i_11_, x728x}, x19796x);
	defparam lut_12592.LUT_SIZE = 5;
	defparam lut_12592.mask = 32'h33ff4011;

	lut_sub lut_12596 ({sk[2247], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1640x);
	defparam lut_12596.LUT_SIZE = 7;
	defparam lut_12596.mask = 128'h0fff0fff7fff7fff0077000070077070;

	lut_sub lut_12609 ({sk[2248], n_n124, x734x, n_n54, x248x, x110x, x409x}, x2026x);
	defparam lut_12609.LUT_SIZE = 7;
	defparam lut_12609.mask = 128'h0fff0fff7fff7fff0000000000007fff;

	lut_sub lut_12614 ({sk[2249], n_n46, n_n47, x1444x, x325x, x1640x, x19792x}, x21329x);
	defparam lut_12614.LUT_SIZE = 7;
	defparam lut_12614.mask = 128'h0fff0fff7fff7fffaaaa800088008000;

	lut_sub lut_12618 ({sk[2250], n_n156, n_n46, n_n177, n_n47, x728x, x628x}, x19805x);
	defparam lut_12618.LUT_SIZE = 7;
	defparam lut_12618.mask = 128'h0fff0fff7fff7fff5555557757577777;

	lut_sub lut_12623 ({sk[2251], i_14_, i_13_, i_12_, i_15_, n_n156}, x19810x);
	defparam lut_12623.LUT_SIZE = 6;
	defparam lut_12623.mask = 64'h7777777705004144;

	lut_sub lut_12630 ({sk[2252], i_14_, i_13_, i_12_, i_15_, n_n149}, x1645x);
	defparam lut_12630.LUT_SIZE = 6;
	defparam lut_12630.mask = 64'h7777777740100401;

	lut_sub lut_12635 ({sk[2253], i_14_, i_13_, i_12_, i_15_, n_n184}, x268x);
	defparam lut_12635.LUT_SIZE = 6;
	defparam lut_12635.mask = 64'h7777777700001044;

	lut_sub lut_12639 ({sk[2254], i_9_, i_10_, i_11_, x725x, x719x, x728x}, x17941x);
	defparam lut_12639.LUT_SIZE = 7;
	defparam lut_12639.mask = 128'h0fff0fff7fff7fff0f00770000770f00;

	lut_sub lut_12646 ({sk[2255], x725x, x157x, x172x, n_n170, x173x, x72x}, x21376x);
	defparam lut_12646.LUT_SIZE = 7;
	defparam lut_12646.mask = 128'h0fff0fff7fff7fff8800000080000000;

	lut_sub lut_12649 ({sk[2256], i_14_, i_13_, i_12_, i_15_, n_n184}, x1648x);
	defparam lut_12649.LUT_SIZE = 6;
	defparam lut_12649.mask = 64'h7777777755554441;

	lut_sub lut_12662 ({sk[2257], i_14_, i_13_, i_12_, i_15_, n_n191, n_n199}, x1653x);
	defparam lut_12662.LUT_SIZE = 7;
	defparam lut_12662.mask = 128'h0fff0fff7fff7fff7000070000700003;

	lut_sub lut_12670 ({sk[2258], i_14_, i_13_, i_12_, i_15_, n_n184}, x1652x);
	defparam lut_12670.LUT_SIZE = 6;
	defparam lut_12670.mask = 64'h7777777740100401;

	lut_sub lut_12675 ({sk[2259], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1657x);
	defparam lut_12675.LUT_SIZE = 7;
	defparam lut_12675.mask = 128'h0fff0fff7fff7fff0000005503030350;

	lut_sub lut_12682 ({sk[2260], i_14_, i_13_, i_12_, i_15_, n_n199}, x1656x);
	defparam lut_12682.LUT_SIZE = 6;
	defparam lut_12682.mask = 64'h7777777700051114;

	lut_sub lut_12689 ({sk[2261], x740x, n_n200, x714x, x17002x, x1657x, x1656x}, x19570x);
	defparam lut_12689.LUT_SIZE = 7;
	defparam lut_12689.mask = 128'h0fff0fff7fff7fff0003000300035557;

	lut_sub lut_12692 ({sk[2262], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1661x);
	defparam lut_12692.LUT_SIZE = 7;
	defparam lut_12692.mask = 128'h0fff0fff7fff7fff0000005507070750;

	lut_sub lut_12702 ({sk[2263], n_n41, n_n40, x48x, x167x, x280x, x1661x}, x19574x);
	defparam lut_12702.LUT_SIZE = 7;
	defparam lut_12702.mask = 128'h0fff0fff7fff7fff00005fff77777fff;

	lut_sub lut_12708 ({sk[2264], n_n138, n_n42, n_n43, n_n116, x391x, x632x}, x19569x);
	defparam lut_12708.LUT_SIZE = 7;
	defparam lut_12708.mask = 128'h0fff0fff7fff7fff777f7f7f777fffff;

	lut_sub lut_12714 ({sk[2265], i_14_, i_13_, i_12_, i_15_, n_n156}, x1665x);
	defparam lut_12714.LUT_SIZE = 6;
	defparam lut_12714.mask = 64'h7777777701004144;

	lut_sub lut_12720 ({sk[2266], i_14_, i_13_, i_12_, i_15_, n_n177}, x1664x);
	defparam lut_12720.LUT_SIZE = 6;
	defparam lut_12720.mask = 64'h7777777705004040;

	lut_sub lut_12725 ({sk[2267], i_7_, i_8_, i_6_, x734x, n_n184, x720x}, x628x);
	defparam lut_12725.LUT_SIZE = 7;
	defparam lut_12725.mask = 128'h0fff0fff7fff7fff0000000000010000;

	lut_sub lut_12727 ({sk[2268], i_9_, i_10_, i_11_, n_n43, x720x}, x697x);
	defparam lut_12727.LUT_SIZE = 6;
	defparam lut_12727.mask = 64'h7777777700001000;

	lut_sub lut_12729 ({sk[2269], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1761x);
	defparam lut_12729.LUT_SIZE = 7;
	defparam lut_12729.mask = 128'h0fff0fff7fff7fff0077000070057050;

	lut_sub lut_12740 ({sk[2270], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1760x);
	defparam lut_12740.LUT_SIZE = 7;
	defparam lut_12740.mask = 128'h0fff0fff7fff7fff0055000050075070;

	lut_sub lut_12749 ({sk[2271], i_9_, i_10_, i_11_, x725x, x719x, x728x}, x17972x);
	defparam lut_12749.LUT_SIZE = 7;
	defparam lut_12749.mask = 128'h0fff0fff7fff7fff0f00770000770f00;

	lut_sub lut_12756 ({sk[2272], i_14_, i_13_, i_12_, i_15_, n_n149, n_n170}, x17970x);
	defparam lut_12756.LUT_SIZE = 7;
	defparam lut_12756.mask = 128'h0fff0fff7fff7fff7000070000500000;

	lut_sub lut_12762 ({sk[2273], x714x, x17051x, x217x, x17972x, x353x, x17970x}, x3773x);
	defparam lut_12762.LUT_SIZE = 7;
	defparam lut_12762.mask = 128'h0fff0fff7fff7fff0000000000007fff;

	lut_sub lut_12767 ({sk[2274], i_9_, i_10_, i_11_, n_n126, x285x}, x17976x);
	defparam lut_12767.LUT_SIZE = 6;
	defparam lut_12767.mask = 64'h7777777701100110;

	lut_sub lut_12772 ({sk[2275], x157x, x172x, x714x, x17051x, x17976x}, x17978x);
	defparam lut_12772.LUT_SIZE = 6;
	defparam lut_12772.mask = 64'h7777777755575757;

	lut_sub lut_12776 ({sk[2276], n_n212, x130x, x63x, x1732x}, x18124x);
	defparam lut_12776.LUT_SIZE = 5;
	defparam lut_12776.mask = 32'h33ff007f;

	lut_sub lut_12780 ({sk[2277], x132x, n_n212, x134x, x123x, x149x, x156x}, x18127x);
	defparam lut_12780.LUT_SIZE = 7;
	defparam lut_12780.mask = 128'h0fff0fff7fff7fff00007fff0000ffff;

	lut_sub lut_12786 ({sk[2278], x157x, n_n36, n_n34, x186x, x588x, x174x}, n_n2635);
	defparam lut_12786.LUT_SIZE = 7;
	defparam lut_12786.mask = 128'h0fff0fff7fff7fff33773f7f3377ffff;

	lut_sub lut_12791 ({sk[2279], i_9_, i_10_, i_11_, i_15_, n_n207, n_n209}, x163x);
	defparam lut_12791.LUT_SIZE = 7;
	defparam lut_12791.mask = 128'h0fff0fff7fff7fff0000730000000000;

	lut_sub lut_12795 ({sk[2280], i_14_, i_13_, i_12_, i_15_, n_n149, x163x}, x19578x);
	defparam lut_12795.LUT_SIZE = 7;
	defparam lut_12795.mask = 128'h0fff0fff7fff7fff5555555557575755;

	lut_sub lut_12800 ({sk[2281], i_9_, i_10_, i_11_, i_15_, x194x, n_n209}, x19579x);
	defparam lut_12800.LUT_SIZE = 7;
	defparam lut_12800.mask = 128'h0fff0fff7fff7fff3733333337333337;

	lut_sub lut_12805 ({sk[2282], i_9_, i_10_, i_11_, i_15_, n_n207, n_n209}, x1673x);
	defparam lut_12805.LUT_SIZE = 7;
	defparam lut_12805.mask = 128'h0fff0fff7fff7fff0500730005050000;

	lut_sub lut_12812 ({sk[2283], n_n46, n_n47, x719x, n_n199, n_n216, x1673x}, x19582x);
	defparam lut_12812.LUT_SIZE = 7;
	defparam lut_12812.mask = 128'h0fff0fff7fff7fff0000557f000f557f;

	lut_sub lut_12817 ({sk[2284], n_n46, n_n47, x55x, x134x, x19578x, x19579x}, x19583x);
	defparam lut_12817.LUT_SIZE = 7;
	defparam lut_12817.mask = 128'h0fff0fff7fff7fff000000ff7f7f7fff;

	lut_sub lut_12822 ({sk[2285], i_14_, i_13_, i_12_, i_15_, n_n191}, x1737x);
	defparam lut_12822.LUT_SIZE = 6;
	defparam lut_12822.mask = 64'h7777777700051014;

	lut_sub lut_12828 ({sk[2286], n_n42, n_n43, x602x, n_n190, n_n183, x1737x}, n_n834);
	defparam lut_12828.LUT_SIZE = 7;
	defparam lut_12828.mask = 128'h0fff0fff7fff7fff00ff5fff33ff7fff;

	lut_sub lut_12833 ({sk[2287], n_n6266, n_n6268, n_n42, n_n43, x340x, x107x}, x19591x);
	defparam lut_12833.LUT_SIZE = 7;
	defparam lut_12833.mask = 128'h77777f7fffffffff0577ffffffffffff;

	lut_sub lut_12839 ({sk[2288], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1679x);
	defparam lut_12839.LUT_SIZE = 7;
	defparam lut_12839.mask = 128'h77777f7fffffffff0000007705050570;

	lut_sub lut_12849 ({sk[2289], x46x, n_n46, n_n47, x134x, x194x, x1679x}, x19596x);
	defparam lut_12849.LUT_SIZE = 7;
	defparam lut_12849.mask = 128'h77777f7fffffffff007f557f007fffff;

	lut_sub lut_12855 ({sk[2290], n_n46, n_n43, n_n177, x719x, n_n183, x19588x}, x19590x);
	defparam lut_12855.LUT_SIZE = 7;
	defparam lut_12855.mask = 128'h77777f7fffffffff55557777555f777f;

	lut_sub lut_12859 ({sk[2291], i_14_, i_13_, i_12_, i_15_, n_n41, n_n216}, x19748x);
	defparam lut_12859.LUT_SIZE = 7;
	defparam lut_12859.mask = 128'h77777f7fffffffff0011000010011010;

	lut_sub lut_12866 ({sk[2292], i_14_, i_13_, i_12_, i_15_, n_n199}, x296x);
	defparam lut_12866.LUT_SIZE = 6;
	defparam lut_12866.mask = 64'h55ffffff00000144;

	lut_sub lut_12870 ({sk[2293], n_n43, x130x, n_n182, x128x, x54x, x222x}, x17981x);
	defparam lut_12870.LUT_SIZE = 7;
	defparam lut_12870.mask = 128'h77777f7fffffffff000000007fffffff;

	lut_sub lut_12876 ({sk[2294], n_n43, x52x, x129x, x139x, x63x, x48x}, x17982x);
	defparam lut_12876.LUT_SIZE = 7;
	defparam lut_12876.mask = 128'h77777f7fffffffff000000007fffffff;

	lut_sub lut_12882 ({sk[2295], i_14_, i_13_, i_12_, i_15_, n_n47, n_n216}, x18033x);
	defparam lut_12882.LUT_SIZE = 7;
	defparam lut_12882.mask = 128'h77777f7fffffffff0111101111011110;

	lut_sub lut_12895 ({sk[2296], i_9_, i_10_, i_8_, i_11_, n_n17, x285x}, x18031x);
	defparam lut_12895.LUT_SIZE = 7;
	defparam lut_12895.mask = 128'h33ffffff33ffffff0001001000000010;

	lut_sub lut_12899 ({sk[2297], x168x, x714x, x17051x, x151x, x1897x, x18031x}, x18034x);
	defparam lut_12899.LUT_SIZE = 7;
	defparam lut_12899.mask = 128'h33ffffff33ffffff5555557f555555ff;

	lut_sub lut_12904 ({sk[2298], x714x, x17051x, x129x, x130x, x139x, x128x}, x18037x);
	defparam lut_12904.LUT_SIZE = 7;
	defparam lut_12904.mask = 128'h33ffffff33ffffff0000000000007fff;

	lut_sub lut_12909 ({sk[2299], x46x, x124x, n_n47, x52x, x63x, x48x}, x18038x);
	defparam lut_12909.LUT_SIZE = 7;
	defparam lut_12909.mask = 128'h33ffffff33ffffff007f00ff00ff00ff;

	lut_sub lut_12915 ({sk[2300], i_14_, i_13_, i_12_, i_15_, n_n191, n_n199}, x1698x);
	defparam lut_12915.LUT_SIZE = 7;
	defparam lut_12915.mask = 128'h33ffffff33ffffff7000070000700003;

	lut_sub lut_12923 ({sk[2301], i_14_, i_13_, i_12_, i_15_, n_n184}, x1697x);
	defparam lut_12923.LUT_SIZE = 6;
	defparam lut_12923.mask = 64'h00ffffff40100401;

	lut_sub lut_12928 ({sk[2302], i_14_, i_13_, i_12_, i_15_, n_n184}, x1700x);
	defparam lut_12928.LUT_SIZE = 6;
	defparam lut_12928.mask = 64'h00ffffff11410050;

	lut_sub lut_12935 ({sk[2303], i_14_, i_13_, i_12_, i_15_, n_n184}, x1703x);
	defparam lut_12935.LUT_SIZE = 6;
	defparam lut_12935.mask = 64'h00ffffff11410040;

	lut_sub lut_12941 ({sk[2304], i_14_, i_13_, i_12_, i_15_, n_n191}, x1701x);
	defparam lut_12941.LUT_SIZE = 6;
	defparam lut_12941.mask = 64'h00ffffff01010050;

	lut_sub lut_12946 ({sk[2305], n_n41, n_n40, n_n122, x293x, x1700x, x1703x}, x19010x);
	defparam lut_12946.LUT_SIZE = 7;
	defparam lut_12946.mask = 128'h33ffffff33ffffff000033335fff7fff;

	lut_sub lut_12951 ({sk[2306], i_14_, i_13_, i_12_, i_15_, n_n191}, x1706x);
	defparam lut_12951.LUT_SIZE = 6;
	defparam lut_12951.mask = 64'h00ffffff00051114;

	lut_sub lut_12958 ({sk[2307], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x1705x);
	defparam lut_12958.LUT_SIZE = 7;
	defparam lut_12958.mask = 128'h33ffffff33ffffff0000003000050500;

	lut_sub lut_12962 ({sk[2308], i_9_, i_10_, i_11_, i_15_, n_n209}, x1709x);
	defparam lut_12962.LUT_SIZE = 6;
	defparam lut_12962.mask = 64'h00ffffff01001001;

	lut_sub lut_12966 ({sk[2309], i_9_, i_10_, i_11_, i_15_, n_n209}, x1708x);
	defparam lut_12966.LUT_SIZE = 6;
	defparam lut_12966.mask = 64'h3f3f3f3f00001100;

	lut_sub lut_12969 ({sk[2310], i_9_, i_10_, i_11_, i_15_, n_n209}, x1707x);
	defparam lut_12969.LUT_SIZE = 6;
	defparam lut_12969.mask = 64'h3f3f3f3f10010000;

	lut_sub lut_12972 ({sk[2311], i_14_, i_13_, i_12_, i_15_, n_n149, n_n216}, x1710x);
	defparam lut_12972.LUT_SIZE = 7;
	defparam lut_12972.mask = 128'h3f3f3f3f3f3f3f7f0000003303030335;

	lut_sub lut_12980 ({sk[2312], i_9_, i_10_, i_11_, i_15_, n_n207, n_n209}, x19609x);
	defparam lut_12980.LUT_SIZE = 7;
	defparam lut_12980.mask = 128'h3f3f3f3f3f3f3f7f0000350000050500;

	lut_sub lut_12985 ({sk[2313], n_n101, x445x, n_n132, n_n108, x199x, x19609x}, x19611x);
	defparam lut_12985.LUT_SIZE = 7;
	defparam lut_12985.mask = 128'h3f3f3f3f3f3f3f7f070fffff07ffffff;

	lut_sub lut_12991 ({sk[2314], i_9_, i_10_, i_11_, i_15_, n_n207, n_n209}, x1715x);
	defparam lut_12991.LUT_SIZE = 7;
	defparam lut_12991.mask = 128'h3f3f3f3f3f3f3f7f0000007300000073;

	lut_sub lut_12998 ({sk[2315], i_9_, i_10_, i_8_, i_11_, n_n17, x285x}, x19613x);
	defparam lut_12998.LUT_SIZE = 7;
	defparam lut_12998.mask = 128'h3f3f3f3f3f3f3f7f0101000001000000;

	lut_sub lut_13002 ({sk[2316], n_n46, n_n47, x151x, x47x, x1715x, x19613x}, x19618x);
	defparam lut_13002.LUT_SIZE = 7;
	defparam lut_13002.mask = 128'h3f3f3f3f3f3f3f7f55557fff7fff7fff;

	lut_sub lut_13010 ({sk[2317], n_n156, n_n101, x406x, x719x, x59x, x290x}, x2190x);
	defparam lut_13010.LUT_SIZE = 7;
	defparam lut_13010.mask = 128'h3f3f3f3f3f3f3f7f000077ff00007fff;

	lut_sub lut_13015 ({sk[2318], i_14_, i_13_, i_12_, i_15_, n_n184}, x1719x);
	defparam lut_13015.LUT_SIZE = 6;
	defparam lut_13015.mask = 64'h3f3f3f3f05004444;

	lut_sub lut_13022 ({sk[2319], i_9_, i_10_, i_11_, x735x, n_n126, x728x}, x1957x);
	defparam lut_13022.LUT_SIZE = 7;
	defparam lut_13022.mask = 128'h3f3f3f3f3f3f3f7f0000010000010100;

	lut_sub lut_13026 ({sk[2320], n_n190, n_n112, x255x, n_n60, n_n56, x348x}, x21334x);
	defparam lut_13026.LUT_SIZE = 7;
	defparam lut_13026.mask = 128'h3f3f3f3f3f3f3f7fffcca080ffcc0000;

	lut_sub lut_13031 ({sk[2321], n_n156, n_n123, n_n112, x63x, x728x, x409x}, x21450x);
	defparam lut_13031.LUT_SIZE = 7;
	defparam lut_13031.mask = 128'h3f3f3f3f3f3f3f7ffff0aaa0fff08880;

	lut_sub lut_13038 ({sk[2322], i_14_, i_13_, i_12_, i_15_, n_n184}, x1726x);
	defparam lut_13038.LUT_SIZE = 6;
	defparam lut_13038.mask = 64'h3f3f3f3f40100401;

	lut_sub lut_13043 ({sk[2323], n_n41, n_n214, x180x, x85x, x142x, n_n198}, x17987x);
	defparam lut_13043.LUT_SIZE = 7;
	defparam lut_13043.mask = 128'h3f3f3f3f3f3f3f7f000000007fffffff;

	lut_sub lut_13049 ({sk[2324], n_n41, n_n59, n_n43, x359x, x1107x, x1726x}, x17988x);
	defparam lut_13049.LUT_SIZE = 7;
	defparam lut_13049.mask = 128'h3f3f3f3f3f3f3f7f0f5f0fff3f7f3fff;

	lut_sub lut_13054 ({sk[2325], i_14_, i_13_, i_12_, i_15_, n_n184}, x17992x);
	defparam lut_13054.LUT_SIZE = 6;
	defparam lut_13054.mask = 64'h3f3f3f3f11054040;

	lut_sub lut_13061 ({sk[2326], i_9_, i_10_, i_11_, x729x, x720x, x726x}, x17990x);
	defparam lut_13061.LUT_SIZE = 7;
	defparam lut_13061.mask = 128'h3f3f3f3f3f3f3f7f7f00000000330000;

	lut_sub lut_13066 ({sk[2327], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x17991x);
	defparam lut_13066.LUT_SIZE = 7;
	defparam lut_13066.mask = 128'h3f3f3f3f3f3f3f7f0505005003000330;

	lut_sub lut_13073 ({sk[2328], x729x, x714x, n_n191, x17002x, n_n199, x726x}, x17994x);
	defparam lut_13073.LUT_SIZE = 7;
	defparam lut_13073.mask = 128'h3f3f3f3f3f3f3f7f000001050000030f;

	lut_sub lut_13078 ({sk[2329], n_n41, x1832x, x17992x, x17990x, x17991x, x17994x}, n_n3480);
	defparam lut_13078.LUT_SIZE = 7;
	defparam lut_13078.mask = 128'h3f3f3f3f3f3f3f7f555555557fffffff;

	lut_sub lut_13084 ({sk[2330], x714x, x17002x, x720x, n_n170, x225x, x1819x}, x17998x);
	defparam lut_13084.LUT_SIZE = 7;
	defparam lut_13084.mask = 128'h3f3f3f3f3f3f3f7f000000000000777f;

	lut_sub lut_13088 ({sk[2331], n_n41, x69x, x397x, x100x, x1898x, x1900x}, x17999x);
	defparam lut_13088.LUT_SIZE = 7;
	defparam lut_13088.mask = 128'h3f3f3f3f3f3f3f7f00ff00ff7fffffff;

	lut_sub lut_13094 ({sk[2332], x245x, x714x, x17002x, n_n5060, n_n57, x503x}, x18012x);
	defparam lut_13094.LUT_SIZE = 7;
	defparam lut_13094.mask = 128'h3f3f3f3f3f3f3f7f5f5f5f7f5f5f5fff;

	lut_sub lut_13099 ({sk[2333], i_14_, i_13_, i_12_, i_15_, n_n191}, x18005x);
	defparam lut_13099.LUT_SIZE = 6;
	defparam lut_13099.mask = 64'h3f3f3f3f40100401;

	lut_sub lut_13104 ({sk[2334], i_14_, i_13_, i_12_, i_15_, n_n184, n_n199}, x18006x);
	defparam lut_13104.LUT_SIZE = 7;
	defparam lut_13104.mask = 128'h3f3f3f3f3f3f3f7f7000030000300003;

	lut_sub lut_13110 ({sk[2335], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x18009x);
	defparam lut_13110.LUT_SIZE = 7;
	defparam lut_13110.mask = 128'h3f3f3f3f3f3f3f7f7000050000500005;

	lut_sub lut_13116 ({sk[2336], n_n41, x186x, x209x, x18005x, x18006x, x18009x}, x18013x);
	defparam lut_13116.LUT_SIZE = 7;
	defparam lut_13116.mask = 128'h3f3f3f3f3f3f3f7f000000007fffffff;

	lut_sub lut_13122 ({sk[2337], i_14_, i_13_, i_12_, i_15_, n_n149, n_n216}, x18015x);
	defparam lut_13122.LUT_SIZE = 7;
	defparam lut_13122.mask = 128'h3f3f3f3f3f3f3f7f0030300000030005;

	lut_sub lut_13127 ({sk[2338], i_14_, i_13_, i_12_, i_15_, n_n149, n_n199}, x18016x);
	defparam lut_13127.LUT_SIZE = 7;
	defparam lut_13127.mask = 128'h3f3f3f3f3f3f3f7f0303053000500005;

	lut_sub lut_13134 ({sk[2339], x714x, x17002x, x141x, x363x, x18015x, x18016x}, x18019x);
	defparam lut_13134.LUT_SIZE = 7;
	defparam lut_13134.mask = 128'h3f3f3f3f3f3f3f7f0f0f0f0f0f0f7fff;

	lut_sub lut_13139 ({sk[2340], i_14_, i_13_, i_12_, i_15_, n_n149, n_n170}, x18020x);
	defparam lut_13139.LUT_SIZE = 7;
	defparam lut_13139.mask = 128'h3f3f3f3f3f3f3f7f0030000000050500;

	lut_sub lut_13143 ({sk[2341], n_n39, n_n84, x279x, x249x, x237x, x18020x}, x21440x);
	defparam lut_13143.LUT_SIZE = 7;
	defparam lut_13143.mask = 128'h3f3f3f3f3f3f3f7fffffffff80000000;

	lut_sub lut_13146 ({sk[2342], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1735x);
	defparam lut_13146.LUT_SIZE = 7;
	defparam lut_13146.mask = 128'h3f3f3f3f3f3f3f7f0707700700007300;

	lut_sub lut_13158 ({sk[2343], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1734x);
	defparam lut_13158.LUT_SIZE = 7;
	defparam lut_13158.mask = 128'h3f3f3f3f3f3f3f7f0303300300003700;

	lut_sub lut_13166 ({sk[2344], i_14_, i_13_, i_12_, i_15_, n_n149, n_n170}, x1739x);
	defparam lut_13166.LUT_SIZE = 7;
	defparam lut_13166.mask = 128'h3f3f3f3f3f3f3f7f0000007707070770;

	lut_sub lut_13179 ({sk[2345], i_9_, i_10_, i_11_, i_15_, n_n34, n_n209}, x19494x);
	defparam lut_13179.LUT_SIZE = 7;
	defparam lut_13179.mask = 128'h3f3f3f3f3f3f3f7f0000000000010100;

	lut_sub lut_13182 ({sk[2346], n_n156, n_n36, n_n33, x719x, n_n170, x48x}, x21449x);
	defparam lut_13182.LUT_SIZE = 7;
	defparam lut_13182.mask = 128'h3f3f3f3f3f3f3f7fffaafca8ffaaf0a0;

	lut_sub lut_13189 ({sk[2347], i_15_, n_n149, n_n36, n_n34, n_n209}, x2317x);
	defparam lut_13189.LUT_SIZE = 6;
	defparam lut_13189.mask = 64'h3f3f3f3f00000015;

	lut_sub lut_13192 ({sk[2348], i_14_, i_13_, i_12_, i_15_, n_n184, n_n177}, x1741x);
	defparam lut_13192.LUT_SIZE = 7;
	defparam lut_13192.mask = 128'h3f3f3f3f3f3f3f7f0000005707030370;

	lut_sub lut_13202 ({sk[2349], i_14_, i_13_, i_12_, i_15_, n_n184, n_n170}, x1740x);
	defparam lut_13202.LUT_SIZE = 7;
	defparam lut_13202.mask = 128'h3f3f3f3f3f3f3f7f0000003707050570;

	lut_sub lut_13212 ({sk[2350], n_n101, n_n108, x1706x, x1705x, x1741x, x1740x}, n_n776);
	defparam lut_13212.LUT_SIZE = 7;
	defparam lut_13212.mask = 128'h3f3f3f3f3f3f3f7f00003f3f55ff7fff;

	lut_sub lut_13217 ({sk[2351], i_14_, i_13_, i_12_, i_15_, n_n149, n_n177}, x1743x);
	defparam lut_13217.LUT_SIZE = 7;
	defparam lut_13217.mask = 128'h3f3f3f3f3f3f3f7f0000007707030370;

	lut_sub lut_13228 ({sk[2352], i_14_, i_13_, i_12_, i_15_, n_n149, n_n156}, x1742x);
	defparam lut_13228.LUT_SIZE = 7;
	defparam lut_13228.mask = 128'h3f3f3f3f3f3f3f7f0000005505070750;

	lut_sub lut_13237 ({sk[2353], i_14_, i_13_, i_12_, i_15_, n_n170}, x1756x);
	defparam lut_13237.LUT_SIZE = 6;
	defparam lut_13237.mask = 64'h3f3f3f3f00051114;

	lut_sub lut_13244 ({sk[2354], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1755x);
	defparam lut_13244.LUT_SIZE = 7;
	defparam lut_13244.mask = 128'h33ff33ff33ff33ff0000005000030300;

	lut_sub lut_13248 ({sk[2355], n_n101, n_n108, x1743x, x1742x, x1756x, x1755x}, x19637x);
	defparam lut_13248.LUT_SIZE = 7;
	defparam lut_13248.mask = 128'h33ff33ff33ff33ff00003f3f55ff7fff;

	lut_sub lut_13253 ({sk[2356], i_14_, i_13_, i_12_, i_15_, n_n149, n_n216}, x19853x);
	defparam lut_13253.LUT_SIZE = 7;
	defparam lut_13253.mask = 128'h33ff33ff33ff33ff0003000030533030;

	lut_sub lut_13260 ({sk[2357], i_9_, i_10_, i_11_, x726x, x728x}, x19848x);
	defparam lut_13260.LUT_SIZE = 6;
	defparam lut_13260.mask = 64'h3f3fffff00000035;

	lut_sub lut_13263 ({sk[2358], n_n150, n_n62, n_n60, x248x, n_n143, x110x}, x21333x);
	defparam lut_13263.LUT_SIZE = 7;
	defparam lut_13263.mask = 128'h0000ffffffffffff8000000000000000;

	lut_sub lut_13265 ({sk[2359], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1748x);
	defparam lut_13265.LUT_SIZE = 7;
	defparam lut_13265.mask = 128'h0000ffffffffffff0303000337073730;

	lut_sub lut_13278 ({sk[2360], i_9_, n_n113, x256x, n_n109}, x21375x);
	defparam lut_13278.LUT_SIZE = 5;
	defparam lut_13278.mask = 32'h7777a8fc;

	lut_sub lut_13283 ({sk[2361], x734x, x181x, n_n126, x1894x, x1748x, x21375x}, n_n3492);
	defparam lut_13283.LUT_SIZE = 7;
	defparam lut_13283.mask = 128'h0000ffffffffffffaaaaaaaaaabfaaff;

	lut_sub lut_13288 ({sk[2362], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x18051x);
	defparam lut_13288.LUT_SIZE = 7;
	defparam lut_13288.mask = 128'h0000ffffffffffff0373707350005050;

	lut_sub lut_13301 ({sk[2363], i_14_, i_13_, i_12_, i_15_, n_n191, n_n199}, x18046x);
	defparam lut_13301.LUT_SIZE = 7;
	defparam lut_13301.mask = 128'h0000ffffffffffff0353505300000000;

	lut_sub lut_13308 ({sk[2364], x124x, n_n108, x48x, x128x, x18051x, x18046x}, n_n3491);
	defparam lut_13308.LUT_SIZE = 7;
	defparam lut_13308.mask = 128'h0000ffffffffffff00007fff0000ffff;

	lut_sub lut_13314 ({sk[2365], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1751x);
	defparam lut_13314.LUT_SIZE = 7;
	defparam lut_13314.mask = 128'h0f1f1f1f0f1f1f1f7000070000700007;

	lut_sub lut_13323 ({sk[2366], i_14_, i_13_, i_12_, i_15_, n_n184}, x1750x);
	defparam lut_13323.LUT_SIZE = 6;
	defparam lut_13323.mask = 64'h1f1f1fff15454401;

	lut_sub lut_13333 ({sk[2367], n_n125, n_n57, n_n113, x54x, x1645x, x268x}, x18057x);
	defparam lut_13333.LUT_SIZE = 7;
	defparam lut_13333.mask = 128'h0f1f1f1f0f1f1f1f005f005f337fffff;

	lut_sub lut_13338 ({sk[2368], x735x, n_n126, n_n113, x1751x, x1750x}, x18058x);
	defparam lut_13338.LUT_SIZE = 6;
	defparam lut_13338.mask = 64'h1f1f1fff05050537;

	lut_sub lut_13341 ({sk[2369], i_14_, i_13_, i_12_, i_15_, n_n149}, x18064x);
	defparam lut_13341.LUT_SIZE = 6;
	defparam lut_13341.mask = 64'h1f1f1fff15455154;

	lut_sub lut_13354 ({sk[2370], n_n108, x125x, x176x, x1892x, x356x, x18064x}, n_n3489);
	defparam lut_13354.LUT_SIZE = 7;
	defparam lut_13354.mask = 128'h0f1f1f1f0f1f1f1f000000007fffffff;

	lut_sub lut_13360 ({sk[2371], i_14_, i_13_, i_12_, i_15_, n_n149, n_n191}, x18065x);
	defparam lut_13360.LUT_SIZE = 7;
	defparam lut_13360.mask = 128'h0f1f1f1f0f1f1f1f7000070000500000;

	lut_sub lut_13366 ({sk[2372], i_9_, i_10_, i_11_, x725x, x719x, x721x}, x18067x);
	defparam lut_13366.LUT_SIZE = 7;
	defparam lut_13366.mask = 128'h0fff0fffffffffff0033005f335f0000;

	lut_sub lut_13373 ({sk[2373], i_9_, i_10_, i_11_, x725x, x719x, x728x}, x18068x);
	defparam lut_13373.LUT_SIZE = 7;
	defparam lut_13373.mask = 128'h0fff0fffffffffff0f00770000770f00;

	lut_sub lut_13380 ({sk[2374], n_n108, x150x, x217x, x18065x, x18067x, x18068x}, x3685x);
	defparam lut_13380.LUT_SIZE = 7;
	defparam lut_13380.mask = 128'h0fff0fffffffffff000000007fffffff;

	lut_sub lut_13386 ({sk[2375], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x18075x);
	defparam lut_13386.LUT_SIZE = 7;
	defparam lut_13386.mask = 128'h0fff0fffffffffff0555505507070700;

	lut_sub lut_13399 ({sk[2376], x157x, n_n108, x131x, x126x, x1489x, x18075x}, x21435x);
	defparam lut_13399.LUT_SIZE = 7;
	defparam lut_13399.mask = 128'h0fff0fffffffffffffff8000ffff0000;

	lut_sub lut_13402 ({sk[2377], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1758x);
	defparam lut_13402.LUT_SIZE = 7;
	defparam lut_13402.mask = 128'h0fff0fffffffffff0000007707050570;

	lut_sub lut_13413 ({sk[2378], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x21344x);
	defparam lut_13413.LUT_SIZE = 7;
	defparam lut_13413.mask = 128'h0fff0fffffffffffffffff88f8f8f88f;

	lut_sub lut_13422 ({sk[2379], n_n123, n_n125, x59x, x290x, x1758x, x21344x}, x19657x);
	defparam lut_13422.LUT_SIZE = 7;
	defparam lut_13422.mask = 128'h77ff77ff77ff77ff00003fffaaaabfff;

	lut_sub lut_13427 ({sk[2380], x735x, n_n161, n_n191, x720x, x187x, x2149x}, x19651x);
	defparam lut_13427.LUT_SIZE = 7;
	defparam lut_13427.mask = 128'h77ff77ff77ff77ff555555555555777f;

	lut_sub lut_13431 ({sk[2381], i_14_, i_13_, i_12_, i_15_, n_n212, n_n199}, x18130x);
	defparam lut_13431.LUT_SIZE = 7;
	defparam lut_13431.mask = 128'h77ff77ff77ff77ff0111101111011110;

	lut_sub lut_13444 ({sk[2382], x181x, n_n212, x48x, x1572x}, x18131x);
	defparam lut_13444.LUT_SIZE = 5;
	defparam lut_13444.mask = 32'h33ff070f;

	lut_sub lut_13448 ({sk[2383], x137x, x46x, n_n212, x1847x, x1857x, x1833x}, x21374x);
	defparam lut_13448.LUT_SIZE = 7;
	defparam lut_13448.mask = 128'h77ff77ff77ff77ffff80ff00ff00ff00;

	lut_sub lut_13451 ({sk[2384], i_14_, i_13_, i_12_, i_15_, n_n156}, x1770x);
	defparam lut_13451.LUT_SIZE = 6;
	defparam lut_13451.mask = 64'h3fff3fff00051114;

	lut_sub lut_13458 ({sk[2385], i_9_, i_10_, i_11_, i_15_, x720x, n_n207}, x1769x);
	defparam lut_13458.LUT_SIZE = 7;
	defparam lut_13458.mask = 128'h77ff77ff77ff77ff0000330000550000;

	lut_sub lut_13462 ({sk[2386], i_9_, i_10_, i_11_, i_15_, n_n207, n_n209}, x1772x);
	defparam lut_13462.LUT_SIZE = 7;
	defparam lut_13462.mask = 128'h77ff77ff77ff77ff0500730005000005;

	lut_sub lut_13469 ({sk[2387], i_9_, i_10_, i_11_, i_15_, n_n207, n_n209}, x1771x);
	defparam lut_13469.LUT_SIZE = 7;
	defparam lut_13469.mask = 128'h77ff77ff77ff77ff0500730005050000;

	lut_sub lut_13476 ({sk[2388], n_n197, n_n212, n_n140, n_n142, x853x, x1771x}, x19670x);
	defparam lut_13476.LUT_SIZE = 7;
	defparam lut_13476.mask = 128'h77ff77ff77ff77ff00005fff33ff7fff;

	lut_sub lut_13482 ({sk[2389], n_n134, n_n197, n_n212, n_n132, x55x, x1772x}, x19671x);
	defparam lut_13482.LUT_SIZE = 7;
	defparam lut_13482.mask = 128'h77ff77ff77ff77ff003f5f7f003fffff;

	lut_sub lut_13488 ({sk[2390], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1775x);
	defparam lut_13488.LUT_SIZE = 7;
	defparam lut_13488.mask = 128'h77ff77ff77ff77ff0000003707070770;

	lut_sub lut_13500 ({sk[2391], i_14_, i_13_, i_12_, i_15_, n_n199, n_n216}, x1774x);
	defparam lut_13500.LUT_SIZE = 7;
	defparam lut_13500.mask = 128'h77ff77ff77ff77ff0000007303030330;

	lut_sub lut_13508 ({sk[2392], n_n128, n_n125, x188x, x1009x, x1774x, x2138x}, x19674x);
	defparam lut_13508.LUT_SIZE = 7;
	defparam lut_13508.mask = 128'h77ff77ff77ff77ff55557f7f55ff7fff;

	lut_sub lut_13513 ({sk[2393], i_14_, i_13_, i_12_, i_15_, n_n191}, x1782x);
	defparam lut_13513.LUT_SIZE = 6;
	defparam lut_13513.mask = 64'h3fff3fff15455054;

	lut_sub lut_13525 ({sk[2394], i_14_, i_13_, i_12_, i_15_, n_n184, n_n191}, x1781x);
	defparam lut_13525.LUT_SIZE = 7;
	defparam lut_13525.mask = 128'h77ff77ff77ff77ff0333303000000005;

	lut_sub lut_13532 ({sk[2395], i_14_, i_13_, i_12_, i_15_, n_n170}, x1783x);
	defparam lut_13532.LUT_SIZE = 6;
	defparam lut_13532.mask = 64'h3fff3fff55555554;

	lut_sub lut_13548 ({sk[2396], i_14_, i_13_, i_12_, i_15_, n_n191}, x1786x);
	defparam lut_13548.LUT_SIZE = 6;
	defparam lut_13548.mask = 64'h3fff3fff15455054;

	lut_sub lut_13560 ({sk[2397], i_14_, i_13_, i_12_, i_15_, n_n184}, x1785x);
	defparam lut_13560.LUT_SIZE = 6;
	defparam lut_13560.mask = 64'h3fff3fff11055054;

	lut_sub lut_13570 ({sk[2398], i_14_, i_13_, i_12_, i_15_, n_n191}, x1787x);
	defparam lut_13570.LUT_SIZE = 6;
	defparam lut_13570.mask = 64'h3fff3fff10045000;

	lut_sub lut_13575 ({sk[2399], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1800x);
	defparam lut_13575.LUT_SIZE = 7;
	defparam lut_13575.mask = 128'h77ff77ff77ff77ff0707700700007300;

	lut_sub lut_13587 ({sk[2400], n_n41, n_n40, n_n83, x991x, x990x, x1799x}, x19021x);
	defparam lut_13587.LUT_SIZE = 7;
	defparam lut_13587.mask = 128'h77ff77ff77ff77ff000033335fff7fff;

	lut_sub lut_13592 ({sk[2401], i_7_, i_8_, i_6_, x740x, x1800x, x19021x}, x19022x);
	defparam lut_13592.LUT_SIZE = 7;
	defparam lut_13592.mask = 128'h77ff77ff77ff77ff5555555557555555;

	lut_sub lut_13595 ({sk[2402], n_n41, n_n40, x261x, x375x, x1701x, x1735x}, x21355x);
	defparam lut_13595.LUT_SIZE = 7;
	defparam lut_13595.mask = 128'h77ff77ff77ff77ffffffc00088888000;

	lut_sub lut_13600 ({sk[2403], x740x, n_n200, n_n1885, x19010x, x1734x, x21355x}, x19023x);
	defparam lut_13600.LUT_SIZE = 7;
	defparam lut_13600.mask = 128'h77ff77ff77ff77ffafffafffafffbfff;

	lut_sub lut_13605 ({sk[2404], i_14_, i_13_, i_12_, i_15_, n_n184}, x1795x);
	defparam lut_13605.LUT_SIZE = 6;
	defparam lut_13605.mask = 64'h3fff3fff14445000;

	lut_sub lut_13612 ({sk[2405], i_7_, i_8_, i_6_, x735x, n_n4225, x1817x}, x17129x);
	defparam lut_13612.LUT_SIZE = 7;
	defparam lut_13612.mask = 128'h77ff77ff77ff77ff3333333733333333;

	lut_sub lut_13615 ({sk[2406], x137x, n_n197, n_n212, x149x, x146x, x131x}, x17118x);
	defparam lut_13615.LUT_SIZE = 7;
	defparam lut_13615.mask = 128'h77ff77ff77ff77ff000f777f000fffff;

	lut_sub lut_13620 ({sk[2407], x46x, n_n197, n_n212, x125x, n_n4231, x17118x}, x17120x);
	defparam lut_13620.LUT_SIZE = 7;
	defparam lut_13620.mask = 128'h77ff77ff77ff77ff777f777f777fffff;

	lut_sub lut_13625 ({sk[2408], n_n125, x17108x, x17109x, x17115x, x1837x, x1838x}, x17121x);
	defparam lut_13625.LUT_SIZE = 7;
	defparam lut_13625.mask = 128'h77ff77ff77ff77ff0fffffff7fffffff;

	lut_sub lut_13631 ({sk[2409], n_n125, n_n169, x69x, x4757x, x225x, x1901x}, x17134x);
	defparam lut_13631.LUT_SIZE = 7;
	defparam lut_13631.mask = 128'h77ff77ff77ff77ff0f0f0f0f7fffffff;

	lut_sub lut_13637 ({sk[2410], i_14_, i_13_, i_12_, i_15_, n_n177}, x1797x);
	defparam lut_13637.LUT_SIZE = 6;
	defparam lut_13637.mask = 64'h3fff3fff15454040;

	lut_sub lut_13646 ({sk[2411], n_n123, x601x, n_n4658, x1171x, n_n4657, x4769x}, x17137x);
	defparam lut_13646.LUT_SIZE = 7;
	defparam lut_13646.mask = 128'h77ff77ff77ff77ff77ffffff7fffffff;

	lut_sub lut_13652 ({sk[2412], n_n123, n_n125, n_n142, x141x, x153x, x1797x}, x17138x);
	defparam lut_13652.LUT_SIZE = 7;
	defparam lut_13652.mask = 128'h77ff77ff77ff77ff000033335fff7fff;

	lut_sub lut_13657 ({sk[2413], n_n124, x735x, x86x, x180x, x1802x, x21458x}, x21404x);
	defparam lut_13657.LUT_SIZE = 7;
	defparam lut_13657.mask = 128'h77ff77ff77ff77ff5555555555554000;

	lut_sub lut_13661 ({sk[2414], x17129x, x17134x, x17137x, x17138x, x21404x}, n_n4409);
	defparam lut_13661.LUT_SIZE = 6;
	defparam lut_13661.mask = 64'h3fff3fffbfffffff;

	lut_sub lut_13667 ({sk[2415], x137x, x46x, n_n212, x147x, x126x}, x17143x);
	defparam lut_13667.LUT_SIZE = 6;
	defparam lut_13667.mask = 64'h3fff3fff070f0f0f;

	lut_sub lut_13672 ({sk[2416], i_8_, n_n17, x735x, n_n212, x1833x, x1856x}, x17144x);
	defparam lut_13672.LUT_SIZE = 7;
	defparam lut_13672.mask = 128'h77ff77ff77ff77ff0303035703030303;

	lut_sub lut_13675 ({sk[2417], x181x, x132x, x735x, n_n200, n_n212, x149x}, x17145x);
	defparam lut_13675.LUT_SIZE = 7;
	defparam lut_13675.mask = 128'h77ff77ff77ff77ff0005333f000f333f;

	lut_sub lut_13680 ({sk[2418], n_n4441, x575x, x17143x, x17144x, x17145x}, x17149x);
	defparam lut_13680.LUT_SIZE = 6;
	defparam lut_13680.mask = 64'h3fff3fff7fffffff;

	lut_sub lut_13686 ({sk[2419], i_14_, i_13_, i_12_, i_15_, n_n184}, x1798x);
	defparam lut_13686.LUT_SIZE = 6;
	defparam lut_13686.mask = 64'h3fff3fff00015054;

	lut_sub lut_13693 ({sk[2420], i_14_, i_13_, i_12_, i_15_, n_n156, n_n170}, x1799x);
	defparam lut_13693.LUT_SIZE = 7;
	defparam lut_13693.mask = 128'h77ff77ff77ff77ff0505500500005700;

	lut_sub lut_13701 ({sk[2421], i_14_, i_13_, i_12_, i_15_, n_n177, n_n170}, x1802x);
	defparam lut_13701.LUT_SIZE = 7;
	defparam lut_13701.mask = 128'h77ff77ff77ff77ff0555505557005770;

	lut_sub lut_13716 ({sk[2422], i_14_, i_13_, i_12_, i_15_, n_n191, n_n170}, x1813x);
	defparam lut_13716.LUT_SIZE = 7;
	defparam lut_13716.mask = 128'h77ff77ff77ff77ff7000070000700007;

	lut_sub lut_13725 ({sk[2423], i_14_, i_13_, i_12_, i_15_, n_n177}, x1861x);
	defparam lut_13725.LUT_SIZE = 6;
	defparam lut_13725.mask = 64'h3fff3fff15440000;

	lut_sub lut_13731 ({sk[2424], i_14_, i_13_, i_12_, i_15_, n_n170}, x19809x);
	defparam lut_13731.LUT_SIZE = 6;
	defparam lut_13731.mask = 64'h3fff3fff05004144;

	lut_sub lut_13738 ({sk[2425], i_7_, i_8_, i_6_, x735x, n_n212, n_n54}, x1973x);
	defparam lut_13738.LUT_SIZE = 7;
	defparam lut_13738.mask = 128'h77ff77ff77ff77ff1111111115111111;

	lut_sub lut_13741 ({sk[2426], i_15_, n_n156, x735x, n_n200, n_n212, n_n209}, x2138x);
	defparam lut_13741.LUT_SIZE = 7;
	defparam lut_13741.mask = 128'h77ff77ff77ff77ff0000000000001115;

	lut_sub lut_13744 ({sk[2427], i_9_, i_10_, i_11_, i_15_, n_n125, n_n209}, x2149x);
	defparam lut_13744.LUT_SIZE = 7;
	defparam lut_13744.mask = 128'h77ff77ff77ff77ff0000010000010100;

	lut_sub lut_13748 ({sk[2428], i_14_, i_13_, i_12_, i_15_, n_n46, n_n199}, x2470x);
	defparam lut_13748.LUT_SIZE = 7;
	defparam lut_13748.mask = 128'h77ff77ff77ff77ff0000000000010110;

	lut_sub lut_13752 ({sk[2429], i_9_, i_10_, i_11_, n_n197, x721x, x728x}, x2519x);
	defparam lut_13752.LUT_SIZE = 7;
	defparam lut_13752.mask = 128'h77ff77ff77ff77ff0000070000070000;

	lut_sub lut_13757 ({sk[2430], i_9_, i_10_, i_11_, n_n125, x721x, x728x}, x2549x);
	defparam lut_13757.LUT_SIZE = 7;
	defparam lut_13757.mask = 128'h77ff77ff77ff77ff0000000700000007;

	lut_sub lut_13762 ({sk[2431], i_9_, i_10_, i_11_, n_n34, x721x, x728x}, x2684x);
	defparam lut_13762.LUT_SIZE = 7;
	defparam lut_13762.mask = 128'h77ff77ff77ff77ff0000070000000700;

	lut_sub lut_13767 ({sk[2432], n_n135, n_n134, n_n36, x209x, x217x, x174x}, x3836x);
	defparam lut_13767.LUT_SIZE = 7;
	defparam lut_13767.mask = 128'h77ff77ff77ff77ff007f00ff00ff00ff;

	lut_sub lut_13773 ({sk[2433], i_7_, i_8_, i_6_, x735x, x135x}, x4769x);
	defparam lut_13773.LUT_SIZE = 6;
	defparam lut_13773.mask = 64'h3fff3fff00010000;

	lut_sub lut_13775 ({sk[2434], x445x, x446x, x448x, n_n47, n_n214, x85x}, x17077x);
	defparam lut_13775.LUT_SIZE = 7;
	defparam lut_13775.mask = 128'h77ff77ff77ff77ff07ffffffffffffff;

	lut_sub lut_13781 ({sk[2435], n_n124, x734x, n_n126, n_n132, x150x, x1168x}, x17078x);
	defparam lut_13781.LUT_SIZE = 7;
	defparam lut_13781.mask = 128'h77ff77ff77ff77ff0000003f0000557f;

	lut_sub lut_13785 ({sk[2436], n_n101, n_n108, n_n169, x69x, x250x, x1860x}, x17153x);
	defparam lut_13785.LUT_SIZE = 7;
	defparam lut_13785.mask = 128'h77ff77ff77ff77ff000055ff3f3f7fff;

	lut_sub lut_13790 ({sk[2437], n_n5144, n_n31, n_n30, x181x, x137x, x46x}, x17169x);
	defparam lut_13790.LUT_SIZE = 7;
	defparam lut_13790.mask = 128'h77ff77ff77ff77ff000f777fffffffff;

	lut_sub lut_13795 ({sk[2438], n_n31, n_n30, x1449x, x132x, x146x, x131x}, x17170x);
	defparam lut_13795.LUT_SIZE = 7;
	defparam lut_13795.mask = 128'h77ff77ff77ff77ff00000fff77777fff;

	lut_sub lut_13800 ({sk[2439], n_n71, n_n36, n_n34, n_n77, x892x, x891x}, x17325x);
	defparam lut_13800.LUT_SIZE = 7;
	defparam lut_13800.mask = 128'h77ff77ff77ff77ff005f337f005fffff;

	lut_sub lut_13805 ({sk[2440], n_n36, n_n34, n_n83, n_n77, x982x, x980x}, x17326x);
	defparam lut_13805.LUT_SIZE = 7;
	defparam lut_13805.mask = 128'h77ff77ff77ff77ff000055553fff7fff;

	lut_sub lut_13810 ({sk[2441], i_10_, i_11_, x725x, n_n197, n_n212}, x21399x);
	defparam lut_13810.LUT_SIZE = 6;
	defparam lut_13810.mask = 64'h3fff3ffffffff8ff;

	lut_sub lut_13815 ({sk[2442], n_n46, n_n47, x890x, x17195x, x417x, x21429x}, x21455x);
	defparam lut_13815.LUT_SIZE = 7;
	defparam lut_13815.mask = 128'h77ff77ff77ff77ffaaaa8800a0008000;

	lut_sub lut_13820 ({sk[2443], i_14_, i_13_, i_12_, i_15_, n_n149, n_n33}, x17417x);
	defparam lut_13820.LUT_SIZE = 7;
	defparam lut_13820.mask = 128'h77ff77ff77ff77ff0010100000000001;

	lut_sub lut_13824 ({sk[2444], n_n31, n_n34, x143x, x122x, x1825x, x17417x}, x17420x);
	defparam lut_13824.LUT_SIZE = 7;
	defparam lut_13824.mask = 128'h77ff77ff77ff77ff55555f5f77ff7fff;

	lut_sub lut_13829 ({sk[2445], n_n149, n_n200, x419x, n_n47, n_n214, x285x}, x21432x);
	defparam lut_13829.LUT_SIZE = 7;
	defparam lut_13829.mask = 128'h77ff77ff77ff77fffc00fc00fc00a800;

	lut_sub lut_13836 ({sk[2446], n_n53, x157x, n_n123, n_n5739, n_n199, n_n109}, x21437x);
	defparam lut_13836.LUT_SIZE = 7;
	defparam lut_13836.mask = 128'h77ff77ff77ff77ff1f1f1fff1fff1fff;

	lut_sub lut_13847 ({sk[2447], x740x, x157x, n_n161, n_n47, x90x, n_n142}, x17556x);
	defparam lut_13847.LUT_SIZE = 7;
	defparam lut_13847.mask = 128'h77ff77ff77ff77ff05050f0f05370f3f;

	lut_sub lut_13851 ({sk[2448], x152x, n_n4308, x435x, x512x, x603x, n_n47}, x17562x);
	defparam lut_13851.LUT_SIZE = 7;
	defparam lut_13851.mask = 128'h77ff77ff77ff77ff3fffffff7fffffff;

	lut_sub lut_13857 ({sk[2449], n_n31, x734x, n_n200, x947x, x1827x, x1876x}, x21387x);
	defparam lut_13857.LUT_SIZE = 7;
	defparam lut_13857.mask = 128'h77ff77ff77ff77fffffffff088888880;

	lut_sub lut_13864 ({sk[2450], i_7_, i_5_, i_6_, x286x, x741x, x744x}, x17598x);
	defparam lut_13864.LUT_SIZE = 7;
	defparam lut_13864.mask = 128'h77ff77ff77ff77ff55775577000f0000;

	lut_sub lut_13869 ({sk[2451], n_n36, n_n34, x52x, x129x, x146x, x131x}, x17835x);
	defparam lut_13869.LUT_SIZE = 7;
	defparam lut_13869.mask = 128'h77ff77ff77ff77ff000077770fff7fff;

	lut_sub lut_13874 ({sk[2452], x137x, x46x, n_n36, n_n3961, x1877x, x3945x}, x17836x);
	defparam lut_13874.LUT_SIZE = 7;
	defparam lut_13874.mask = 128'h77ff77ff77ff77ff5f7f5fff5fff5fff;

	lut_sub lut_13880 ({sk[2453], n_n5144, n_n156, n_n31, n_n30, x725x, x157x}, x17841x);
	defparam lut_13880.LUT_SIZE = 7;
	defparam lut_13880.mask = 128'h77ff77ff77ff77ff05050737ffffffff;

	lut_sub lut_13885 ({sk[2454], n_n31, x17786x, n_n63, x125x, x1456x, x17841x}, x17842x);
	defparam lut_13885.LUT_SIZE = 7;
	defparam lut_13885.mask = 128'h77ff77ff77ff77ff5555ffff7fffffff;

	lut_sub lut_13891 ({sk[2455], i_7_, i_5_, i_6_, i_3_, i_4_, n_n19}, x17857x);
	defparam lut_13891.LUT_SIZE = 7;
	defparam lut_13891.mask = 128'h77ff77ff77ff77ff0000000050101000;

	lut_sub lut_13896 ({sk[2456], i_7_, i_6_, n_n219, n_n162, n_n19, n_n48}, x17858x);
	defparam lut_13896.LUT_SIZE = 7;
	defparam lut_13896.mask = 128'h77ff77ff77ff77ff000000000303131f;

	lut_sub lut_13901 ({sk[2457], n_n5144, n_n156, x725x, n_n36, n_n128, x152x}, x17912x);
	defparam lut_13901.LUT_SIZE = 7;
	defparam lut_13901.mask = 128'h77ff77ff77ff77ff0707070fffffffff;

	lut_sub lut_13906 ({sk[2458], x714x, x17051x, x176x, x123x, x350x, x356x}, x18137x);
	defparam lut_13906.LUT_SIZE = 7;
	defparam lut_13906.mask = 128'h77ff77ff77ff77ff0000000000007fff;

	lut_sub lut_13911 ({sk[2459], x714x, x17051x, x125x, x55x, x158x, x1888x}, x18138x);
	defparam lut_13911.LUT_SIZE = 7;
	defparam lut_13911.mask = 128'h77ff77ff77ff77ff0000000000007fff;

	lut_sub lut_13916 ({sk[2460], n_n5144, n_n7257, n_n7259, n_n7263, n_n14, x253x}, x18164x);
	defparam lut_13916.LUT_SIZE = 7;
	defparam lut_13916.mask = 128'h77ff77ff77ff77ff1fffffffffffffff;

	lut_sub lut_13922 ({sk[2461], i_9_, i_10_, i_8_, i_11_, n_n16, x285x}, x18221x);
	defparam lut_13922.LUT_SIZE = 7;
	defparam lut_13922.mask = 128'h77ff77ff77ff77ff0001100000010010;

	lut_sub lut_13927 ({sk[2462], x729x, x53x, n_n41, n_n177, x726x, x469x}, x21445x);
	defparam lut_13927.LUT_SIZE = 7;
	defparam lut_13927.mask = 128'h77ff77ff77ff77ff005700ff005f00ff;

	lut_sub lut_13936 ({sk[2463], x740x, n_n200, x714x, x17002x, x115x, x247x}, x21448x);
	defparam lut_13936.LUT_SIZE = 7;
	defparam lut_13936.mask = 128'h77ff77ff77ff77fffffcfffcfffcaaa8;

	lut_sub lut_13946 ({sk[2464], i_7_, i_6_, x741x, x744x, x748x, x731x}, x18373x);
	defparam lut_13946.LUT_SIZE = 7;
	defparam lut_13946.mask = 128'h77ff77ff77ff77ff33ff00ff00ff5fff;

	lut_sub lut_13954 ({sk[2465], i_9_, i_10_, i_11_, x729x, x719x, x728x}, x18389x);
	defparam lut_13954.LUT_SIZE = 7;
	defparam lut_13954.mask = 128'h77ff77ff77ff77ff0000003300000f77;

	lut_sub lut_13959 ({sk[2466], n_n41, n_n40, x1382x, x1381x, x1521x, x1520x}, x21366x);
	defparam lut_13959.LUT_SIZE = 7;
	defparam lut_13959.mask = 128'h77ff77ff77ff77ffffffcc00a0a08000;

	lut_sub lut_13964 ({sk[2467], i_7_, i_5_, i_6_, i_3_, i_4_, n_n219}, x18503x);
	defparam lut_13964.LUT_SIZE = 7;
	defparam lut_13964.mask = 128'h77ff77ff77ff77ff0000000040404040;

	lut_sub lut_13969 ({sk[2468], i_7_, i_6_, n_n219, n_n19, n_n48, x746x}, x18504x);
	defparam lut_13969.LUT_SIZE = 7;
	defparam lut_13969.mask = 128'h77ff77ff77ff77ff5757577757775577;

	lut_sub lut_13980 ({sk[2469], n_n5144, n_n156, x725x, n_n128, x152x, n_n212}, x18620x);
	defparam lut_13980.LUT_SIZE = 7;
	defparam lut_13980.mask = 128'h77ff77ff77ff77ff15151555ffffffff;

	lut_sub lut_13985 ({sk[2470], i_9_, i_10_, i_8_, i_11_, n_n18, x285x}, x18666x);
	defparam lut_13985.LUT_SIZE = 7;
	defparam lut_13985.mask = 128'h77ff77ff77ff77ff0011000111000100;

	lut_sub lut_13992 ({sk[2471], n_n138, n_n101, n_n42, n_n108, x1265x, x1264x}, x21451x);
	defparam lut_13992.LUT_SIZE = 7;
	defparam lut_13992.mask = 128'h77ff77ff77ff77fffafac8c8fa00c800;

	lut_sub lut_14001 ({sk[2472], i_8_, n_n5144, x734x, n_n16, x381x, x21451x}, x18691x);
	defparam lut_14001.LUT_SIZE = 7;
	defparam lut_14001.mask = 128'h77ff77ff77ff77ffaaabffffaaaaffff;

	lut_sub lut_14005 ({sk[2473], i_9_, i_10_, i_11_, n_n6, n_n12, x730x}, x18715x);
	defparam lut_14005.LUT_SIZE = 7;
	defparam lut_14005.mask = 128'h77ff77ff77ff77ff0000110005001500;

	lut_sub lut_14010 ({sk[2474], n_n31, n_n30, x795x, n_n82, n_n169, n_n77}, x18735x);
	defparam lut_14010.LUT_SIZE = 7;
	defparam lut_14010.mask = 128'h77ff77ff77ff77ff00007fff3f3f7fff;

	lut_sub lut_14017 ({sk[2475], n_n36, n_n34, n_n32, n_n133, x1248x, x1247x}, x18827x);
	defparam lut_14017.LUT_SIZE = 7;
	defparam lut_14017.mask = 128'h77ff77ff77ff77ff00335f7f55775f7f;

	lut_sub lut_14022 ({sk[2476], i_7_, i_6_, x744x, x746x}, x18839x);
	defparam lut_14022.LUT_SIZE = 5;
	defparam lut_14022.mask = 32'h33ff3377;

	lut_sub lut_14029 ({sk[2477], i_9_, i_10_, i_11_, n_n123, n_n125, x721x}, x21361x);
	defparam lut_14029.LUT_SIZE = 7;
	defparam lut_14029.mask = 128'h77ff77ff77ff77ffffffeaffffeaeaff;

	lut_sub lut_14048 ({sk[2478], i_9_, i_10_, i_11_, n_n46, n_n47, x721x}, x18971x);
	defparam lut_14048.LUT_SIZE = 7;
	defparam lut_14048.mask = 128'h77ff77ff77ff77ff0015150000050500;

	lut_sub lut_14055 ({sk[2479], n_n123, x70x, n_n125, n_n102, n_n198, x930x}, x19273x);
	defparam lut_14055.LUT_SIZE = 7;
	defparam lut_14055.mask = 128'h77ff77ff77ff77ff007f007f007fffff;

	lut_sub lut_14060 ({sk[2480], x393x, n_n36, n_n34, n_n198, x522x, x1609x}, x19538x);
	defparam lut_14060.LUT_SIZE = 7;
	defparam lut_14060.mask = 128'h77ff77ff77ff77ff333f777fffffffff;

	lut_sub lut_14065 ({sk[2481], i_9_, i_10_, i_11_, n_n46, n_n47, x719x}, x19588x);
	defparam lut_14065.LUT_SIZE = 7;
	defparam lut_14065.mask = 128'h77ff77ff77ff77ff0015150000001500;

	lut_sub lut_14072 ({sk[2482], n_n5144, n_n31, n_n30, x777x, x776x, x775x}, x19688x);
	defparam lut_14072.LUT_SIZE = 7;
	defparam lut_14072.mask = 128'h77ff77ff77ff77ff00775f7fffffffff;

	lut_sub lut_14078 ({sk[2483], i_9_, i_10_, i_8_, i_11_, n_n17, x285x}, x19792x);
	defparam lut_14078.LUT_SIZE = 7;
	defparam lut_14078.mask = 128'h77ff77ff77ff77ff0000101000001000;

	lut_sub lut_14082 ({sk[2484], n_n149, n_n156, n_n38, n_n39, x140x, x728x}, x19864x);
	defparam lut_14082.LUT_SIZE = 7;
	defparam lut_14082.mask = 128'h77ff77ff77ff77ff0033057705770577;

	lut_sub lut_14088 ({sk[2485], i_14_, i_13_, i_12_, i_15_, n_n156, n_n34}, x19889x);
	defparam lut_14088.LUT_SIZE = 7;
	defparam lut_14088.mask = 128'h77ff77ff77ff77ff0011000010011010;

	lut_sub lut_14095 ({sk[2486], n_n150, n_n199, n_n216, x728x, x110x, x1593x}, x21338x);
	defparam lut_14095.LUT_SIZE = 7;
	defparam lut_14095.mask = 128'h77ff77ff77ff77ff8880808000000000;

	lut_sub lut_14098 ({sk[2487], i_9_, i_10_, i_11_, x725x, x267x, x388x}, x19925x);
	defparam lut_14098.LUT_SIZE = 7;
	defparam lut_14098.mask = 128'h77ff77ff77ff77ff5555575557555555;

	lut_sub lut_14102 ({sk[2488], i_7_, i_6_, x741x, x731x, x746x, x527x}, x19940x);
	defparam lut_14102.LUT_SIZE = 7;
	defparam lut_14102.mask = 128'h77ff77ff77ff77ff7f7f7f7f5f5f55ff;

	lut_sub lut_14110 ({sk[2489], n_n124, x735x, n_n126, n_n169, n_n176, x100x}, x21458x);
	defparam lut_14110.LUT_SIZE = 7;
	defparam lut_14110.mask = 128'h77ff77ff77ff77ffffffff88fffff080;

	lut_sub lut_14116 ({sk[2490], x740x, n_n161, n_n47, n_n63, x176x, n_n61}, x21429x);
	defparam lut_14116.LUT_SIZE = 7;
	defparam lut_14116.mask = 128'h77ff77ff77ff77ff005f005f005f777f;

	lut_sub lut_14127 ({sk[2491], n_n53, x157x, n_n123, n_n125, x1106x, x1105x}, x21438x);
	defparam lut_14127.LUT_SIZE = 7;
	defparam lut_14127.mask = 128'h77ff77ff77ff77ff035703ff03ff03ff;


endmodule