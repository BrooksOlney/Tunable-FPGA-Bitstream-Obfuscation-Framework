module misex3_qmap_map (sk, b, e, f, g, n, m, k, j, l, h, i, d, c, a, r2, s2, t2, u2, n2, o2, p2, q2, h2, i2, j2, k2, m2, l2);

	input b;
	input e;
	input f;
	input g;
	input n;
	input m;
	input k;
	input j;
	input l;
	input h;
	input i;
	input d;
	input c;
	input a;
	output r2;
	output s2;
	output t2;
	output u2;
	output n2;
	output o2;
	output p2;
	output q2;
	output h2;
	output i2;
	output j2;
	output k2;
	output m2;
	output l2;



	wire g53, g103, g129, g173, g217, g235, g252, g274, g295, g328, g339, g345, g351, g1, g2, g3, g4, g5, g6, g7, g8;
	wire g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29;
	wire g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50;
	wire g51, g455, g52, g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71;
	wire g72, g73, g74, g75, g76, g77, g78, g79, g80, g81, g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92;
	wire g93, g94, g95, g96, g97, g98, g99, g100, g101, g539, g102, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113;
	wire g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g130, g131, g132, g532, g133, g134;
	wire g135, g136, g137, g138, g139, g140, g141, g142, g525, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154;
	wire g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g511, g170, g171, g172, g518, g174;
	wire g175, g176, g504, g177, g178, g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194;
	wire g195, g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207, g208, g497, g209, g210, g211, g212, g213, g214;
	wire g215, g216, g218, g219, g220, g221, g222, g223, g224, g225, g226, g227, g228, g229, g230, g231, g232, g233, g234, g236, g237;
	wire g238, g239, g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250, g251, g253, g254, g255, g256, g257, g258, g259;
	wire g260, g261, g262, g263, g264, g265, g266, g267, g268, g269, g270, g271, g479, g272, g273, g486, g275, g276, g277, g278, g279;
	wire g280, g281, g282, g283, g284, g285, g286, g287, g472, g288, g289, g290, g291, g292, g293, g294, g296, g297, g298, g299, g300;
	wire g301, g302, g303, g304, g305, g306, g307, g308, g309, g310, g311, g312, g313, g314, g315, g316, g317, g318, g319, g320, g321;
	wire g322, g323, g324, g325, g326, g327, g329, g330, g331, g332, g333, g334, g335, g336, g337, g338, g340, g341, g342, g343, g344;
	wire g346, g347, g348, g349, g350, g352, g353, g354, g355, g356, g357, g358, g359, g360, g361, g362, g363, g364, g365, g366, g367;
	wire g368, g369, g370, g371, g372, g373, g374, g375, g376, g377, g378, g379, g380, g381, g462, g382, g383, g384, g385, g386, g387;
	wire g388, g389, g390, g391, g392, g393, g394, g395, g396, g397, g398, g399, g400, g401, g402, g403, g404, g405, g406, g407, g408;
	wire g409, g410, g411, g412, g413, g414, g415, g416, g417, g418, g419, g420, g421, g422, g423, g424, g425, g426, g427, g428, g429;
	wire g430, g431, g432, g433, g434, g435, g436, g437, g438, g439, g440, g441, g442, g443, g444, g445, g446, g456, g447, g448, g449;
	wire g450, g451, g453, g454, g457, g458, g459, g460, g461, g463, g464, g465, g468, g466, g467, g469, g470, g471, g473, g474, g475;
	wire g476, g477, g478, g480, g481, g482, g483, g484, g485, g487, g488, g489, g492, g490, g491, g494, g495, g493, g496, g498, g499;
	wire g500, g501, g502, g503, g505, g506, g507, g508, g509, g510, g512, g513, g514, g515, g516, g517, g519, g520, g521, g522, g523;
	wire g524, g526, g527, g528, g529, g530, g531, g533, g534, g535, g536, g537, g538, g540, g541, g542, g545, g543, g544, g547, g548;
	wire g546, g549;

	lut_sub lut_19 ({g53}, r2);
	defparam lut_19.LUT_SIZE = 1;
	defparam lut_19.mask = 2'b10;

	lut_sub lut_23 ({g103}, s2);
	defparam lut_23.LUT_SIZE = 1;
	defparam lut_23.mask = 2'b10;

	lut_sub lut_27 ({g129}, t2);
	defparam lut_27.LUT_SIZE = 1;
	defparam lut_27.mask = 2'b10;

	lut_sub lut_31 ({g173}, u2);
	defparam lut_31.LUT_SIZE = 1;
	defparam lut_31.mask = 2'b10;

	lut_sub lut_35 ({g217}, n2);
	defparam lut_35.LUT_SIZE = 1;
	defparam lut_35.mask = 2'b10;

	lut_sub lut_39 ({g235}, o2);
	defparam lut_39.LUT_SIZE = 1;
	defparam lut_39.mask = 2'b10;

	lut_sub lut_43 ({g252}, p2);
	defparam lut_43.LUT_SIZE = 1;
	defparam lut_43.mask = 2'b10;

	lut_sub lut_47 ({g274}, q2);
	defparam lut_47.LUT_SIZE = 1;
	defparam lut_47.mask = 2'b10;

	lut_sub lut_51 ({g295}, h2);
	defparam lut_51.LUT_SIZE = 1;
	defparam lut_51.mask = 2'b10;

	lut_sub lut_55 ({g328}, i2);
	defparam lut_55.LUT_SIZE = 1;
	defparam lut_55.mask = 2'b10;

	lut_sub lut_59 ({g339}, j2);
	defparam lut_59.LUT_SIZE = 1;
	defparam lut_59.mask = 2'b10;

	lut_sub lut_63 ({g345}, k2);
	defparam lut_63.LUT_SIZE = 1;
	defparam lut_63.mask = 2'b10;

	lut_sub lut_67 ({g351}, m2);
	defparam lut_67.LUT_SIZE = 1;
	defparam lut_67.mask = 2'b10;

	lut_sub lut_71 ({n, m}, g1);
	defparam lut_71.LUT_SIZE = 2;
	defparam lut_71.mask = 4'b0010;

	lut_sub lut_75 ({n, m, j, l}, g2);
	defparam lut_75.LUT_SIZE = 4;
	defparam lut_75.mask = 16'h0040;

	lut_sub lut_81 ({k, g1, g2}, g3);
	defparam lut_81.LUT_SIZE = 3;
	defparam lut_81.mask = 8'ha8;

	lut_sub lut_88 ({k, g1}, g4);
	defparam lut_88.LUT_SIZE = 2;
	defparam lut_88.mask = 4'b0001;

	lut_sub lut_93 ({h, g, j, i, g4}, g5);
	defparam lut_93.LUT_SIZE = 5;
	defparam lut_93.mask = 32'h33005400;

	lut_sub lut_103 ({h, j, k, l}, g6);
	defparam lut_103.LUT_SIZE = 4;
	defparam lut_103.mask = 16'h002e;

	lut_sub lut_114 ({g, g1, g3, g5, g6}, g7);
	defparam lut_114.LUT_SIZE = 5;
	defparam lut_114.mask = 32'h30753030;

	lut_sub lut_129 ({e, f, g7}, g8);
	defparam lut_129.LUT_SIZE = 3;
	defparam lut_129.mask = 8'h10;

	lut_sub lut_133 ({n, m}, g9);
	defparam lut_133.LUT_SIZE = 2;
	defparam lut_133.mask = 4'b1000;

	lut_sub lut_137 ({h, i}, g10);
	defparam lut_137.LUT_SIZE = 2;
	defparam lut_137.mask = 4'b0100;

	lut_sub lut_141 ({h, j, k, i, l}, g11);
	defparam lut_141.LUT_SIZE = 5;
	defparam lut_141.mask = 32'h03030ffe;

	lut_sub lut_162 ({j, l, g9, g10, g11}, g12);
	defparam lut_162.LUT_SIZE = 5;
	defparam lut_162.mask = 32'h05070505;

	lut_sub lut_175 ({d, e, f, g12, c}, g13);
	defparam lut_175.LUT_SIZE = 5;
	defparam lut_175.mask = 32'h01010100;

	lut_sub lut_181 ({h, j, k, l}, g14);
	defparam lut_181.LUT_SIZE = 4;
	defparam lut_181.mask = 16'h0073;

	lut_sub lut_189 ({n, m}, g15);
	defparam lut_189.LUT_SIZE = 2;
	defparam lut_189.mask = 4'b0100;

	lut_sub lut_193 ({b, d, a}, g16);
	defparam lut_193.LUT_SIZE = 3;
	defparam lut_193.mask = 8'h01;

	lut_sub lut_197 ({h, j, k, i, l}, g17);
	defparam lut_197.LUT_SIZE = 5;
	defparam lut_197.mask = 32'he4a8b101;

	lut_sub lut_213 ({j, k, i, g17}, g18);
	defparam lut_213.LUT_SIZE = 4;
	defparam lut_213.mask = 16'h5415;

	lut_sub lut_226 ({e, g, g14, g15, g16, g18}, g19);
	defparam lut_226.LUT_SIZE = 6;
	defparam lut_226.mask = 64'h0003020200000000;

	lut_sub lut_233 ({d, e, c}, g20);
	defparam lut_233.LUT_SIZE = 3;
	defparam lut_233.mask = 8'h01;

	lut_sub lut_237 ({n, m, j, k, l}, g21);
	defparam lut_237.LUT_SIZE = 5;
	defparam lut_237.mask = 32'h73000000;

	lut_sub lut_247 ({f, g10, g21}, g22);
	defparam lut_247.LUT_SIZE = 3;
	defparam lut_247.mask = 8'h10;

	lut_sub lut_251 ({f, h}, g23);
	defparam lut_251.LUT_SIZE = 2;
	defparam lut_251.mask = 4'b0100;

	lut_sub lut_257 ({j, k, i, l, g9, g23}, g24);
	defparam lut_257.LUT_SIZE = 6;
	defparam lut_257.mask = 64'h0000111111111110;

	lut_sub lut_272 ({b, h, i, g1}, g25);
	defparam lut_272.LUT_SIZE = 4;
	defparam lut_272.mask = 16'h0015;

	lut_sub lut_278 ({h, j, k, i, l}, g26);
	defparam lut_278.LUT_SIZE = 5;
	defparam lut_278.mask = 32'ha0f0f001;

	lut_sub lut_294 ({e, f, c, g25, g26}, g27);
	defparam lut_294.LUT_SIZE = 5;
	defparam lut_294.mask = 32'h00000200;

	lut_sub lut_303 ({g19, g20, g22, g24, g27}, g28);
	defparam lut_303.LUT_SIZE = 5;
	defparam lut_303.mask = 32'haa800000;

	lut_sub lut_311 ({j, k, i}, g29);
	defparam lut_311.LUT_SIZE = 3;
	defparam lut_311.mask = 8'h18;

	lut_sub lut_316 ({b, d, e, c, a}, g30);
	defparam lut_316.LUT_SIZE = 5;
	defparam lut_316.mask = 32'h00000e0a;

	lut_sub lut_324 ({n, m, j, k, i, l}, g31);
	defparam lut_324.LUT_SIZE = 6;
	defparam lut_324.mask = 64'h000000000ffe0000;

	lut_sub lut_338 ({n, m, j, k, i, l}, g32);
	defparam lut_338.LUT_SIZE = 6;
	defparam lut_338.mask = 64'h0000000013030000;

	lut_sub lut_348 ({h, g31, g32}, g33);
	defparam lut_348.LUT_SIZE = 3;
	defparam lut_348.mask = 8'hac;

	lut_sub lut_355 ({e, g}, g34);
	defparam lut_355.LUT_SIZE = 2;
	defparam lut_355.mask = 4'b0100;

	lut_sub lut_359 ({b, c}, g35);
	defparam lut_359.LUT_SIZE = 2;
	defparam lut_359.mask = 4'b0001;

	lut_sub lut_364 ({d, g35}, g36);
	defparam lut_364.LUT_SIZE = 2;
	defparam lut_364.mask = 4'b0100;

	lut_sub lut_368 ({b, d, c}, g37);
	defparam lut_368.LUT_SIZE = 3;
	defparam lut_368.mask = 8'h02;

	lut_sub lut_376 ({f, g33, g34, g36, g37}, g38);
	defparam lut_376.LUT_SIZE = 5;
	defparam lut_376.mask = 32'h03005700;

	lut_sub lut_386 ({b, d, e}, g39);
	defparam lut_386.LUT_SIZE = 3;
	defparam lut_386.mask = 8'hfb;

	lut_sub lut_396 ({f, h, g}, g40);
	defparam lut_396.LUT_SIZE = 3;
	defparam lut_396.mask = 8'h01;

	lut_sub lut_400 ({f, h, g}, g41);
	defparam lut_400.LUT_SIZE = 3;
	defparam lut_400.mask = 8'h04;

	lut_sub lut_408 ({g40, g31, g41, g32}, g42);
	defparam lut_408.LUT_SIZE = 4;
	defparam lut_408.mask = 16'h111f;

	lut_sub lut_418 ({b, d, e}, g43);
	defparam lut_418.LUT_SIZE = 3;
	defparam lut_418.mask = 8'h02;

	lut_sub lut_422 ({f, h}, g44);
	defparam lut_422.LUT_SIZE = 2;
	defparam lut_422.mask = 4'b0001;

	lut_sub lut_428 ({g44, j, k, i, l, g1}, g45);
	defparam lut_428.LUT_SIZE = 6;
	defparam lut_428.mask = 64'h0000000000555554;

	lut_sub lut_447 ({f, g10, g4, g2, g43, g45}, g46);
	defparam lut_447.LUT_SIZE = 6;
	defparam lut_447.mask = 64'h1111111111111333;

	lut_sub lut_471 ({g14, g15}, g47);
	defparam lut_471.LUT_SIZE = 2;
	defparam lut_471.mask = 4'b0001;

	lut_sub lut_478 ({g15, g29, g17}, g48);
	defparam lut_478.LUT_SIZE = 3;
	defparam lut_478.mask = 8'h0b;

	lut_sub lut_485 ({d, a, g35}, g49);
	defparam lut_485.LUT_SIZE = 3;
	defparam lut_485.mask = 8'h10;

	lut_sub lut_492 ({e, g, g47, g48, g49}, g50);
	defparam lut_492.LUT_SIZE = 5;
	defparam lut_492.mask = 32'h00000511;

	lut_sub lut_503 ({g39, g42, g46, g50}, g51);
	defparam lut_503.LUT_SIZE = 4;
	defparam lut_503.mask = 16'h8088;

	lut_sub lut_513 ({g455, g30, g38, g51}, g52);
	defparam lut_513.LUT_SIZE = 4;
	defparam lut_513.mask = 16'h4044;

	lut_sub lut_523 ({b, g8, g13, g28, g52}, g53);
	defparam lut_523.LUT_SIZE = 5;
	defparam lut_523.mask = 32'h10101000;

	lut_sub lut_529 ({n, m, k}, g54);
	defparam lut_529.LUT_SIZE = 3;
	defparam lut_529.mask = 8'h10;

	lut_sub lut_534 ({h, g, g54}, g55);
	defparam lut_534.LUT_SIZE = 3;
	defparam lut_534.mask = 8'h04;

	lut_sub lut_539 ({e, g55}, g56);
	defparam lut_539.LUT_SIZE = 2;
	defparam lut_539.mask = 4'b0100;

	lut_sub lut_543 ({f, g}, g57);
	defparam lut_543.LUT_SIZE = 2;
	defparam lut_543.mask = 4'b0001;

	lut_sub lut_547 ({j, i}, g58);
	defparam lut_547.LUT_SIZE = 2;
	defparam lut_547.mask = 4'b0010;

	lut_sub lut_552 ({m, k, l, g58}, g59);
	defparam lut_552.LUT_SIZE = 4;
	defparam lut_552.mask = 16'h0008;

	lut_sub lut_556 ({m, j, k, i, l}, g60);
	defparam lut_556.LUT_SIZE = 5;
	defparam lut_556.mask = 32'h000000c4;

	lut_sub lut_562 ({m, k, l}, g61);
	defparam lut_562.LUT_SIZE = 3;
	defparam lut_562.mask = 8'h04;

	lut_sub lut_566 ({m, l}, g62);
	defparam lut_566.LUT_SIZE = 2;
	defparam lut_566.mask = 4'b0001;

	lut_sub lut_571 ({h, j, k, i, g62}, g63);
	defparam lut_571.LUT_SIZE = 5;
	defparam lut_571.mask = 32'h11510051;

	lut_sub lut_582 ({m, j, l}, g64);
	defparam lut_582.LUT_SIZE = 3;
	defparam lut_582.mask = 8'h04;

	lut_sub lut_586 ({m, j, i, l}, g65);
	defparam lut_586.LUT_SIZE = 4;
	defparam lut_586.mask = 16'h004e;

	lut_sub lut_597 ({g44, g, g54, g64, g65}, g66);
	defparam lut_597.LUT_SIZE = 5;
	defparam lut_597.mask = 32'h00003f55;

	lut_sub lut_614 ({h, g57, g61, g63, g66}, g67);
	defparam lut_614.LUT_SIZE = 5;
	defparam lut_614.mask = 32'haa88aaa8;

	lut_sub lut_634 ({n, g57, g59, g60, g67}, g68);
	defparam lut_634.LUT_SIZE = 5;
	defparam lut_634.mask = 32'haabf0000;

	lut_sub lut_649 ({j, g61}, g69);
	defparam lut_649.LUT_SIZE = 2;
	defparam lut_649.mask = 4'b0001;

	lut_sub lut_657 ({h, g34, g65, g60, g69}, g70);
	defparam lut_657.LUT_SIZE = 5;
	defparam lut_657.mask = 32'h0077007f;

	lut_sub lut_673 ({n, m, k, l}, g71);
	defparam lut_673.LUT_SIZE = 4;
	defparam lut_673.mask = 16'h0200;

	lut_sub lut_678 ({e, h, g, j, i, g62}, g72);
	defparam lut_678.LUT_SIZE = 6;
	defparam lut_678.mask = 64'h0011500000000000;

	lut_sub lut_690 ({n, g58, g34, g70, g71, g72}, g73);
	defparam lut_690.LUT_SIZE = 6;
	defparam lut_690.mask = 64'h5f7f5f5f00000000;

	lut_sub lut_722 ({f, g12, a, g56, g68, g73}, g74);
	defparam lut_722.LUT_SIZE = 6;
	defparam lut_722.mask = 64'hff80ff80ff800000;

	lut_sub lut_752 ({e, h, g}, g75);
	defparam lut_752.LUT_SIZE = 3;
	defparam lut_752.mask = 8'h02;

	lut_sub lut_756 ({e, g}, g76);
	defparam lut_756.LUT_SIZE = 2;
	defparam lut_756.mask = 4'b0001;

	lut_sub lut_760 ({m, j, k}, g77);
	defparam lut_760.LUT_SIZE = 3;
	defparam lut_760.mask = 8'h04;

	lut_sub lut_767 ({h, i, g76, g62, g77}, g78);
	defparam lut_767.LUT_SIZE = 5;
	defparam lut_767.mask = 32'h00070005;

	lut_sub lut_780 ({h, g76, g59, g65, g60, g69}, g79);
	defparam lut_780.LUT_SIZE = 6;
	defparam lut_780.mask = 64'h000077ff00007fff;

	lut_sub lut_817 ({n, g54, g75, g64, g78, g79}, g80);
	defparam lut_817.LUT_SIZE = 6;
	defparam lut_817.mask = 64'h777f77ff00000000;

	lut_sub lut_847 ({b, c, a}, g81);
	defparam lut_847.LUT_SIZE = 3;
	defparam lut_847.mask = 8'hef;

	lut_sub lut_857 ({d, e, f}, g82);
	defparam lut_857.LUT_SIZE = 3;
	defparam lut_857.mask = 8'h01;

	lut_sub lut_864 ({g81, g82, g455}, g83);
	defparam lut_864.LUT_SIZE = 3;
	defparam lut_864.mask = 8'h20;

	lut_sub lut_868 ({b, d, a}, g84);
	defparam lut_868.LUT_SIZE = 3;
	defparam lut_868.mask = 8'h02;

	lut_sub lut_874 ({e, f, g, g47, g48}, g85);
	defparam lut_874.LUT_SIZE = 5;
	defparam lut_874.mask = 32'h00350000;

	lut_sub lut_881 ({j, i}, g86);
	defparam lut_881.LUT_SIZE = 2;
	defparam lut_881.mask = 4'b0100;

	lut_sub lut_886 ({n, m, k, g86}, g87);
	defparam lut_886.LUT_SIZE = 4;
	defparam lut_886.mask = 16'h0100;

	lut_sub lut_890 ({d, c, a}, g88);
	defparam lut_890.LUT_SIZE = 3;
	defparam lut_890.mask = 8'hfb;

	lut_sub lut_904 ({g57, g34, g87, g88}, g89);
	defparam lut_904.LUT_SIZE = 4;
	defparam lut_904.mask = 16'h0222;

	lut_sub lut_910 ({b, d, c}, g90);
	defparam lut_910.LUT_SIZE = 3;
	defparam lut_910.mask = 8'h01;

	lut_sub lut_917 ({e, g44, g31, g90}, g91);
	defparam lut_917.LUT_SIZE = 4;
	defparam lut_917.mask = 16'h0100;

	lut_sub lut_923 ({e, f, h, g32, g90}, g92);
	defparam lut_923.LUT_SIZE = 5;
	defparam lut_923.mask = 32'h00100000;

	lut_sub lut_927 ({b, f, c}, g93);
	defparam lut_927.LUT_SIZE = 3;
	defparam lut_927.mask = 8'h10;

	lut_sub lut_934 ({j, l, g1, g10, g11}, g94);
	defparam lut_934.LUT_SIZE = 5;
	defparam lut_934.mask = 32'h05070505;

	lut_sub lut_950 ({f, g34, g36, g93, g94}, g95);
	defparam lut_950.LUT_SIZE = 5;
	defparam lut_950.mask = 32'h11111115;

	lut_sub lut_968 ({g81, g85, g89, g91, g92, g95}, g96);
	defparam lut_968.LUT_SIZE = 6;
	defparam lut_968.mask = 64'h8000000080008000;

	lut_sub lut_974 ({d, c}, g97);
	defparam lut_974.LUT_SIZE = 2;
	defparam lut_974.mask = 4'b0001;

	lut_sub lut_980 ({g9, g6}, g98);
	defparam lut_980.LUT_SIZE = 2;
	defparam lut_980.mask = 4'b0001;

	lut_sub lut_984 ({j, i}, g99);
	defparam lut_984.LUT_SIZE = 2;
	defparam lut_984.mask = 4'b0001;

	lut_sub lut_991 ({g44, k, g9, g99}, g100);
	defparam lut_991.LUT_SIZE = 4;
	defparam lut_991.mask = 16'h0002;

	lut_sub lut_999 ({f, g10, g21, g98, g100}, g101);
	defparam lut_999.LUT_SIZE = 5;
	defparam lut_999.mask = 32'haaaa8880;

	lut_sub lut_1019 ({g80, g83, g28, g84, g96, g539}, g102);
	defparam lut_1019.LUT_SIZE = 6;
	defparam lut_1019.mask = 64'h0011000000100000;

	lut_sub lut_1028 ({d, c, g8, g74, g102}, g103);
	defparam lut_1028.LUT_SIZE = 5;
	defparam lut_1028.mask = 32'h55501150;

	lut_sub lut_1044 ({f, g10, g3, g45}, g104);
	defparam lut_1044.LUT_SIZE = 4;
	defparam lut_1044.mask = 16'haaa2;

	lut_sub lut_1056 ({f, h, g, g31, g32}, g105);
	defparam lut_1056.LUT_SIZE = 5;
	defparam lut_1056.mask = 32'h05030000;

	lut_sub lut_1066 ({e, f, g37, g94, g105}, g106);
	defparam lut_1066.LUT_SIZE = 5;
	defparam lut_1066.mask = 32'h05050507;

	lut_sub lut_1078 ({b, e, c}, g107);
	defparam lut_1078.LUT_SIZE = 3;
	defparam lut_1078.mask = 8'h10;

	lut_sub lut_1083 ({e, f, g12, c}, g108);
	defparam lut_1083.LUT_SIZE = 4;
	defparam lut_1083.mask = 16'h0010;

	lut_sub lut_1089 ({g57, g87}, g109);
	defparam lut_1089.LUT_SIZE = 2;
	defparam lut_1089.mask = 4'b0001;

	lut_sub lut_1094 ({b, d, e, a, g109}, g110);
	defparam lut_1094.LUT_SIZE = 5;
	defparam lut_1094.mask = 32'h00104410;

	lut_sub lut_1101 ({b, d, f, a}, g111);
	defparam lut_1101.LUT_SIZE = 4;
	defparam lut_1101.mask = 16'h0100;

	lut_sub lut_1108 ({f, g, g47, g48, g111}, g112);
	defparam lut_1108.LUT_SIZE = 5;
	defparam lut_1108.mask = 32'h05010511;

	lut_sub lut_1118 ({b, c, a}, g113);
	defparam lut_1118.LUT_SIZE = 3;
	defparam lut_1118.mask = 8'h04;

	lut_sub lut_1122 ({d, c, a}, g114);
	defparam lut_1122.LUT_SIZE = 3;
	defparam lut_1122.mask = 8'h10;

	lut_sub lut_1130 ({g, g14, g15, g29, g17}, g115);
	defparam lut_1130.LUT_SIZE = 5;
	defparam lut_1130.mask = 32'h000f0b0b;

	lut_sub lut_1146 ({d, e, f, g113, g114, g115}, g116);
	defparam lut_1146.LUT_SIZE = 6;
	defparam lut_1146.mask = 64'h0005001500000011;

	lut_sub lut_1161 ({g108, g110, g27, g112, g116}, g117);
	defparam lut_1161.LUT_SIZE = 5;
	defparam lut_1161.mask = 32'h80000000;

	lut_sub lut_1166 ({g, g10}, g118);
	defparam lut_1166.LUT_SIZE = 2;
	defparam lut_1166.mask = 4'b0001;

	lut_sub lut_1170 ({h, g, j}, g119);
	defparam lut_1170.LUT_SIZE = 3;
	defparam lut_1170.mask = 8'h01;

	lut_sub lut_1176 ({k, g1, g119}, g120);
	defparam lut_1176.LUT_SIZE = 3;
	defparam lut_1176.mask = 8'h10;

	lut_sub lut_1182 ({h, g, k, g1, g99}, g121);
	defparam lut_1182.LUT_SIZE = 5;
	defparam lut_1182.mask = 32'h00000002;

	lut_sub lut_1187 ({h, g, k, l, g1}, g122);
	defparam lut_1187.LUT_SIZE = 5;
	defparam lut_1187.mask = 32'h00000004;

	lut_sub lut_1196 ({g3, g118, g120, g121, g122}, g123);
	defparam lut_1196.LUT_SIZE = 5;
	defparam lut_1196.mask = 32'h80008080;

	lut_sub lut_1204 ({j, k, i, l, g1, g23}, g124);
	defparam lut_1204.LUT_SIZE = 6;
	defparam lut_1204.mask = 64'h0000111111111110;

	lut_sub lut_1221 ({f, g10, g3, g124}, g125);
	defparam lut_1221.LUT_SIZE = 4;
	defparam lut_1221.mask = 16'ha2aa;

	lut_sub lut_1232 ({d, e, c, g101}, g126);
	defparam lut_1232.LUT_SIZE = 4;
	defparam lut_1232.mask = 16'h0208;

	lut_sub lut_1241 ({g39, g123, g125, g126}, g127);
	defparam lut_1241.LUT_SIZE = 4;
	defparam lut_1241.mask = 16'h02aa;

	lut_sub lut_1251 ({b, d, e, a, g68, g109}, g128);
	defparam lut_1251.LUT_SIZE = 6;
	defparam lut_1251.mask = 64'h0000030030700370;

	lut_sub lut_1272 ({g104, g106, g107, g117, g127, g128}, g129);
	defparam lut_1272.LUT_SIZE = 6;
	defparam lut_1272.mask = 64'h0200000002020000;

	lut_sub lut_1280 ({g75, g114}, g130);
	defparam lut_1280.LUT_SIZE = 2;
	defparam lut_1280.mask = 4'b0001;

	lut_sub lut_1284 ({b, d, e, c, a}, g131);
	defparam lut_1284.LUT_SIZE = 5;
	defparam lut_1284.mask = 32'hfafefaaa;

	lut_sub lut_1310 ({b, d, e, c, a}, g132);
	defparam lut_1310.LUT_SIZE = 5;
	defparam lut_1310.mask = 32'heeaa11ab;

	lut_sub lut_1332 ({g130, g532}, g133);
	defparam lut_1332.LUT_SIZE = 2;
	defparam lut_1332.mask = 4'b0100;

	lut_sub lut_1336 ({b, e, f, a}, g134);
	defparam lut_1336.LUT_SIZE = 4;
	defparam lut_1336.mask = 16'hfff1;

	lut_sub lut_1352 ({h, g, i}, g135);
	defparam lut_1352.LUT_SIZE = 3;
	defparam lut_1352.mask = 8'h04;

	lut_sub lut_1356 ({h, g, i}, g136);
	defparam lut_1356.LUT_SIZE = 3;
	defparam lut_1356.mask = 8'h01;

	lut_sub lut_1362 ({m, j, l, g135, g136}, g137);
	defparam lut_1362.LUT_SIZE = 5;
	defparam lut_1362.mask = 32'h00000350;

	lut_sub lut_1373 ({g, g99, g61, g134, g137}, g138);
	defparam lut_1373.LUT_SIZE = 5;
	defparam lut_1373.mask = 32'h4444444c;

	lut_sub lut_1385 ({m, j, k, i, l}, g139);
	defparam lut_1385.LUT_SIZE = 5;
	defparam lut_1385.mask = 32'h0ffe0000;

	lut_sub lut_1399 ({d, e, c}, g140);
	defparam lut_1399.LUT_SIZE = 3;
	defparam lut_1399.mask = 8'h10;

	lut_sub lut_1404 ({m, k, i, g41}, g141);
	defparam lut_1404.LUT_SIZE = 4;
	defparam lut_1404.mask = 16'h0100;

	lut_sub lut_1412 ({g40, g139, g140, g141}, g142);
	defparam lut_1412.LUT_SIZE = 4;
	defparam lut_1412.mask = 16'h1113;

	lut_sub lut_1424 ({i, g62, g138, g525, g142}, g143);
	defparam lut_1424.LUT_SIZE = 5;
	defparam lut_1424.mask = 32'ha0a0a020;

	lut_sub lut_1436 ({m, k, i, g133, g143}, g144);
	defparam lut_1436.LUT_SIZE = 5;
	defparam lut_1436.mask = 32'h55555551;

	lut_sub lut_1454 ({j, k}, g145);
	defparam lut_1454.LUT_SIZE = 2;
	defparam lut_1454.mask = 4'b0010;

	lut_sub lut_1458 ({f, h, g}, g146);
	defparam lut_1458.LUT_SIZE = 3;
	defparam lut_1458.mask = 8'h10;

	lut_sub lut_1462 ({d, e, g, c, a}, g147);
	defparam lut_1462.LUT_SIZE = 5;
	defparam lut_1462.mask = 32'h00010000;

	lut_sub lut_1471 ({h, g40, g34, g88, g147, g132}, g148);
	defparam lut_1471.LUT_SIZE = 6;
	defparam lut_1471.mask = 64'h0000aaaa33f3bbfb;

	lut_sub lut_1508 ({g146, g131, g148}, g149);
	defparam lut_1508.LUT_SIZE = 3;
	defparam lut_1508.mask = 8'ha2;

	lut_sub lut_1516 ({g34, g88}, g150);
	defparam lut_1516.LUT_SIZE = 2;
	defparam lut_1516.mask = 4'b0010;

	lut_sub lut_1523 ({f, g, i, g150, g131, g132}, g151);
	defparam lut_1523.LUT_SIZE = 6;
	defparam lut_1523.mask = 64'hffffff30ffffff50;

	lut_sub lut_1579 ({g, g134}, g152);
	defparam lut_1579.LUT_SIZE = 2;
	defparam lut_1579.mask = 4'b0010;

	lut_sub lut_1585 ({g86, g152}, g153);
	defparam lut_1585.LUT_SIZE = 2;
	defparam lut_1585.mask = 4'b0001;

	lut_sub lut_1591 ({g54, g153}, g154);
	defparam lut_1591.LUT_SIZE = 2;
	defparam lut_1591.mask = 4'b0001;

	lut_sub lut_1595 ({e, c, a}, g155);
	defparam lut_1595.LUT_SIZE = 3;
	defparam lut_1595.mask = 8'h01;

	lut_sub lut_1602 ({f, g, g81, g87, g155}, g156);
	defparam lut_1602.LUT_SIZE = 5;
	defparam lut_1602.mask = 32'h00110030;

	lut_sub lut_1612 ({f, g, g113, g16, g87}, g157);
	defparam lut_1612.LUT_SIZE = 5;
	defparam lut_1612.mask = 32'h00110005;

	lut_sub lut_1620 ({d, e, f, g, a, g87}, g158);
	defparam lut_1620.LUT_SIZE = 6;
	defparam lut_1620.mask = 64'h0000010000000000;

	lut_sub lut_1627 ({g87, g158, g147}, g159);
	defparam lut_1627.LUT_SIZE = 3;
	defparam lut_1627.mask = 8'hc8;

	lut_sub lut_1639 ({g89, g110, g154, g156, g157, g159}, g160);
	defparam lut_1639.LUT_SIZE = 6;
	defparam lut_1639.mask = 64'h4000000000000000;

	lut_sub lut_1648 ({g33, g34, g36, g71, g151}, g161);
	defparam lut_1648.LUT_SIZE = 5;
	defparam lut_1648.mask = 32'h222f2222;

	lut_sub lut_1664 ({l, g86, g15}, g162);
	defparam lut_1664.LUT_SIZE = 3;
	defparam lut_1664.mask = 8'h01;

	lut_sub lut_1670 ({h, g, k, g9, g99}, g163);
	defparam lut_1670.LUT_SIZE = 5;
	defparam lut_1670.mask = 32'h00000002;

	lut_sub lut_1678 ({g, g10, g21, g98, g163}, g164);
	defparam lut_1678.LUT_SIZE = 5;
	defparam lut_1678.mask = 32'haaaa8880;

	lut_sub lut_1693 ({d, e, f, c, g164}, g165);
	defparam lut_1693.LUT_SIZE = 5;
	defparam lut_1693.mask = 32'h02208a28;

	lut_sub lut_1706 ({h, n, i, g62, g71, g147}, g166);
	defparam lut_1706.LUT_SIZE = 6;
	defparam lut_1706.mask = 64'h0015001100110011;

	lut_sub lut_1722 ({l, g41, g86, g9, g140}, g167);
	defparam lut_1722.LUT_SIZE = 5;
	defparam lut_1722.mask = 32'h00000001;

	lut_sub lut_1730 ({g54, g134, g135, g167}, g168);
	defparam lut_1730.LUT_SIZE = 4;
	defparam lut_1730.mask = 16'haa8a;

	lut_sub lut_1742 ({b, c, g76, g33}, g169);
	defparam lut_1742.LUT_SIZE = 4;
	defparam lut_1742.mask = 16'h0020;

	lut_sub lut_1752 ({g42, g43, g166, g511, g168, g169}, g170);
	defparam lut_1752.LUT_SIZE = 6;
	defparam lut_1752.mask = 64'h0200020002000000;

	lut_sub lut_1759 ({b, e, f, c, g123}, g171);
	defparam lut_1759.LUT_SIZE = 5;
	defparam lut_1759.mask = 32'h220200a0;

	lut_sub lut_1773 ({g133, g161, g162, g165, g170, g171}, g172);
	defparam lut_1773.LUT_SIZE = 6;
	defparam lut_1773.mask = 64'h2000000020200000;

	lut_sub lut_1783 ({n, m, g144, g518, g160, g172}, g173);
	defparam lut_1783.LUT_SIZE = 6;
	defparam lut_1783.mask = 64'h0011000111111111;

	lut_sub lut_1800 ({h, i, g15, g147, g525}, g174);
	defparam lut_1800.LUT_SIZE = 5;
	defparam lut_1800.mask = 32'h000b000a;

	lut_sub lut_1809 ({k, g174}, g175);
	defparam lut_1809.LUT_SIZE = 2;
	defparam lut_1809.mask = 4'b0001;

	lut_sub lut_1813 ({b, d, e, f, c}, g176);
	defparam lut_1813.LUT_SIZE = 5;
	defparam lut_1813.mask = 32'hffffcac8;

	lut_sub lut_1841 ({g4, g504}, g177);
	defparam lut_1841.LUT_SIZE = 2;
	defparam lut_1841.mask = 4'b0010;

	lut_sub lut_1845 ({d, e, c}, g178);
	defparam lut_1845.LUT_SIZE = 3;
	defparam lut_1845.mask = 8'hf7;

	lut_sub lut_1858 ({n, m, g145, g136, g178}, g179);
	defparam lut_1858.LUT_SIZE = 5;
	defparam lut_1858.mask = 32'h02000000;

	lut_sub lut_1862 ({d, e, f, g, c}, g180);
	defparam lut_1862.LUT_SIZE = 5;
	defparam lut_1862.mask = 32'h05550f5e;

	lut_sub lut_1883 ({h, k, g9, g99, g180}, g181);
	defparam lut_1883.LUT_SIZE = 5;
	defparam lut_1883.mask = 32'h00000100;

	lut_sub lut_1887 ({h, j, i}, g182);
	defparam lut_1887.LUT_SIZE = 3;
	defparam lut_1887.mask = 8'h01;

	lut_sub lut_1894 ({k, g1, g93, g182}, g183);
	defparam lut_1894.LUT_SIZE = 4;
	defparam lut_1894.mask = 16'h0100;

	lut_sub lut_1901 ({g15, g16, g146}, g184);
	defparam lut_1901.LUT_SIZE = 3;
	defparam lut_1901.mask = 8'h01;

	lut_sub lut_1907 ({d, e, g40, c, a, g146}, g185);
	defparam lut_1907.LUT_SIZE = 6;
	defparam lut_1907.mask = 64'h0000111100330101;

	lut_sub lut_1924 ({h, g40, g34, g88, g147}, g186);
	defparam lut_1924.LUT_SIZE = 5;
	defparam lut_1924.mask = 32'h00cc5ddd;

	lut_sub lut_1945 ({h, g, g184, g185, g186}, g187);
	defparam lut_1945.LUT_SIZE = 5;
	defparam lut_1945.mask = 32'ha0a0a080;

	lut_sub lut_1956 ({b, d, g40, c, a}, g188);
	defparam lut_1956.LUT_SIZE = 5;
	defparam lut_1956.mask = 32'h01010e04;

	lut_sub lut_1967 ({b, e, k, a, g15, g119}, g189);
	defparam lut_1967.LUT_SIZE = 6;
	defparam lut_1967.mask = 64'h0000000000001000;

	lut_sub lut_1976 ({g145, g15, g187, g188, g189}, g190);
	defparam lut_1976.LUT_SIZE = 5;
	defparam lut_1976.mask = 32'haaaaaa08;

	lut_sub lut_1992 ({b, d, e, f, c}, g191);
	defparam lut_1992.LUT_SIZE = 5;
	defparam lut_1992.mask = 32'hafafa051;

	lut_sub lut_2013 ({h, g, g191}, g192);
	defparam lut_2013.LUT_SIZE = 3;
	defparam lut_2013.mask = 8'h02;

	lut_sub lut_2018 ({m, g145, i}, g193);
	defparam lut_2018.LUT_SIZE = 3;
	defparam lut_2018.mask = 8'h10;

	lut_sub lut_2022 ({b, d, e, f, h}, g194);
	defparam lut_2022.LUT_SIZE = 5;
	defparam lut_2022.mask = 32'h00000410;

	lut_sub lut_2032 ({n, g135, g176, g192, g193, g194}, g195);
	defparam lut_2032.LUT_SIZE = 6;
	defparam lut_2032.mask = 64'h0000000013133313;

	lut_sub lut_2053 ({g179, g181, g183, g190, g195}, g196);
	defparam lut_2053.LUT_SIZE = 5;
	defparam lut_2053.mask = 32'h20000000;

	lut_sub lut_2059 ({n, m, k, g178, g191}, g197);
	defparam lut_2059.LUT_SIZE = 5;
	defparam lut_2059.mask = 32'h0c000a00;

	lut_sub lut_2068 ({h, g, g99, g197}, g198);
	defparam lut_2068.LUT_SIZE = 4;
	defparam lut_2068.mask = 16'h0004;

	lut_sub lut_2074 ({n, m, g93, g180}, g199);
	defparam lut_2074.LUT_SIZE = 4;
	defparam lut_2074.mask = 16'h5030;

	lut_sub lut_2083 ({h, k, g99, g199}, g200);
	defparam lut_2083.LUT_SIZE = 4;
	defparam lut_2083.mask = 16'h0004;

	lut_sub lut_2090 ({f, g, i, g150, g131, g132}, g201);
	defparam lut_2090.LUT_SIZE = 6;
	defparam lut_2090.mask = 64'h0f00cf000f00af00;

	lut_sub lut_2113 ({j, k, l}, g202);
	defparam lut_2113.LUT_SIZE = 3;
	defparam lut_2113.mask = 8'hfe;

	lut_sub lut_2125 ({g15, g202}, g203);
	defparam lut_2125.LUT_SIZE = 2;
	defparam lut_2125.mask = 4'b0010;

	lut_sub lut_2131 ({j, k, l, g15, g152}, g204);
	defparam lut_2131.LUT_SIZE = 5;
	defparam lut_2131.mask = 32'h00100000;

	lut_sub lut_2136 ({n, m, k, g134}, g205);
	defparam lut_2136.LUT_SIZE = 4;
	defparam lut_2136.mask = 16'h0200;

	lut_sub lut_2142 ({g, l, g10, g58}, g206);
	defparam lut_2142.LUT_SIZE = 4;
	defparam lut_2142.mask = 16'h0007;

	lut_sub lut_2152 ({j, g71, g147, g205, g206}, g207);
	defparam lut_2152.LUT_SIZE = 5;
	defparam lut_2152.mask = 32'h111f1111;

	lut_sub lut_2171 ({i, g147, g201, g203, g204, g207}, g208);
	defparam lut_2171.LUT_SIZE = 6;
	defparam lut_2171.mask = 64'h8880808088808880;

	lut_sub lut_2190 ({g4, g198, g497, g200, g208}, g209);
	defparam lut_2190.LUT_SIZE = 5;
	defparam lut_2190.mask = 32'h44000400;

	lut_sub lut_2199 ({f, g, g150, g131, g132}, g210);
	defparam lut_2199.LUT_SIZE = 5;
	defparam lut_2199.mask = 32'hf030f050;

	lut_sub lut_2214 ({h, g, i}, g211);
	defparam lut_2214.LUT_SIZE = 3;
	defparam lut_2214.mask = 8'hfd;

	lut_sub lut_2224 ({j, i, l}, g212);
	defparam lut_2224.LUT_SIZE = 3;
	defparam lut_2224.mask = 8'h40;

	lut_sub lut_2229 ({d, e, c, a, g146}, g213);
	defparam lut_2229.LUT_SIZE = 5;
	defparam lut_2229.mask = 32'h00110001;

	lut_sub lut_2240 ({g15, g148, g184, g212, g213}, g214);
	defparam lut_2240.LUT_SIZE = 5;
	defparam lut_2240.mask = 32'h03031333;

	lut_sub lut_2258 ({n, g211, g64, g134, g214}, g215);
	defparam lut_2258.LUT_SIZE = 5;
	defparam lut_2258.mask = 32'ha2aaaaaa;

	lut_sub lut_2281 ({j, g71, g118, g134, g210, g215}, g216);
	defparam lut_2281.LUT_SIZE = 6;
	defparam lut_2281.mask = 64'h5555110155555505;

	lut_sub lut_2315 ({g175, g177, g160, g196, g209, g216}, g217);
	defparam lut_2315.LUT_SIZE = 6;
	defparam lut_2315.mask = 64'h0001000000000000;

	lut_sub lut_2319 ({m, j, k}, g218);
	defparam lut_2319.LUT_SIZE = 3;
	defparam lut_2319.mask = 8'h40;

	lut_sub lut_2324 ({n, g218, i}, g219);
	defparam lut_2324.LUT_SIZE = 3;
	defparam lut_2324.mask = 8'h01;

	lut_sub lut_2332 ({k, g10, g199, g194, g219}, g220);
	defparam lut_2332.LUT_SIZE = 5;
	defparam lut_2332.mask = 32'h1111111f;

	lut_sub lut_2349 ({g44, j, g71, g132}, g221);
	defparam lut_2349.LUT_SIZE = 4;
	defparam lut_2349.mask = 16'h0020;

	lut_sub lut_2357 ({n, g218, g135, g176, g221}, g222);
	defparam lut_2357.LUT_SIZE = 5;
	defparam lut_2357.mask = 32'haaaaaaa2;

	lut_sub lut_2376 ({k, l, g15}, g223);
	defparam lut_2376.LUT_SIZE = 3;
	defparam lut_2376.mask = 8'h01;

	lut_sub lut_2381 ({j, i, g223}, g224);
	defparam lut_2381.LUT_SIZE = 3;
	defparam lut_2381.mask = 8'h40;

	lut_sub lut_2388 ({g39, f, g, g10, g176}, g225);
	defparam lut_2388.LUT_SIZE = 5;
	defparam lut_2388.mask = 32'h33202020;

	lut_sub lut_2401 ({f, g10, g43, g225}, g226);
	defparam lut_2401.LUT_SIZE = 4;
	defparam lut_2401.mask = 16'haaa8;

	lut_sub lut_2413 ({n, g178, g191}, g227);
	defparam lut_2413.LUT_SIZE = 3;
	defparam lut_2413.mask = 8'h35;

	lut_sub lut_2425 ({g218, g4, g136, g226, g227}, g228);
	defparam lut_2425.LUT_SIZE = 5;
	defparam lut_2425.mask = 32'h00cc0ace;

	lut_sub lut_2441 ({n, m, k, g93, g180}, g229);
	defparam lut_2441.LUT_SIZE = 5;
	defparam lut_2441.mask = 32'h05000300;

	lut_sub lut_2451 ({f, a, g140, g131, g178}, g230);
	defparam lut_2451.LUT_SIZE = 5;
	defparam lut_2451.mask = 32'h3310ff50;

	lut_sub lut_2472 ({h, j, i, g71, g229, g230}, g231);
	defparam lut_2472.LUT_SIZE = 6;
	defparam lut_2472.mask = 64'h000000000a3b0000;

	lut_sub lut_2488 ({g15, g29, g149, g224, g228, g231}, g232);
	defparam lut_2488.LUT_SIZE = 6;
	defparam lut_2488.mask = 64'h8088808880880088;

	lut_sub lut_2503 ({h, g, j, g205}, g233);
	defparam lut_2503.LUT_SIZE = 4;
	defparam lut_2503.mask = 16'h0054;

	lut_sub lut_2514 ({g54, g118, g133, g197, g233}, g234);
	defparam lut_2514.LUT_SIZE = 5;
	defparam lut_2514.mask = 32'haa880a08;

	lut_sub lut_2531 ({g196, g220, g222, g232, g234}, g235);
	defparam lut_2531.LUT_SIZE = 5;
	defparam lut_2531.mask = 32'h00000100;

	lut_sub lut_2536 ({j, k, l, g174}, g236);
	defparam lut_2536.LUT_SIZE = 4;
	defparam lut_2536.mask = 16'h1015;

	lut_sub lut_2544 ({n, m, g133}, g237);
	defparam lut_2544.LUT_SIZE = 3;
	defparam lut_2544.mask = 8'h13;

	lut_sub lut_2553 ({n, g118, g226, g227}, g238);
	defparam lut_2553.LUT_SIZE = 4;
	defparam lut_2553.mask = 16'h0ace;

	lut_sub lut_2565 ({m, g211, g227}, g239);
	defparam lut_2565.LUT_SIZE = 3;
	defparam lut_2565.mask = 8'h70;

	lut_sub lut_2574 ({n, j, k, g497, g238, g239}, g240);
	defparam lut_2574.LUT_SIZE = 6;
	defparam lut_2574.mask = 64'h000000bb000000fb;

	lut_sub lut_2592 ({j, k, l, g15, g118}, g241);
	defparam lut_2592.LUT_SIZE = 5;
	defparam lut_2592.mask = 32'h01000111;

	lut_sub lut_2601 ({g, k, l, g15, g58}, g242);
	defparam lut_2601.LUT_SIZE = 5;
	defparam lut_2601.mask = 32'h00001101;

	lut_sub lut_2611 ({j, g55, g134, g241, g242}, g243);
	defparam lut_2611.LUT_SIZE = 5;
	defparam lut_2611.mask = 32'h707070f0;

	lut_sub lut_2627 ({n, m, j, k, l}, g244);
	defparam lut_2627.LUT_SIZE = 5;
	defparam lut_2627.mask = 32'h000d0000;

	lut_sub lut_2635 ({n, g60, g147}, g245);
	defparam lut_2635.LUT_SIZE = 3;
	defparam lut_2635.mask = 8'h10;

	lut_sub lut_2642 ({h, g145, g199, g245}, g246);
	defparam lut_2642.LUT_SIZE = 4;
	defparam lut_2642.mask = 16'haaa8;

	lut_sub lut_2654 ({h, g, j, g176, g194}, g247);
	defparam lut_2654.LUT_SIZE = 5;
	defparam lut_2654.mask = 32'h05050d05;

	lut_sub lut_2667 ({h, j, i, g229}, g248);
	defparam lut_2667.LUT_SIZE = 4;
	defparam lut_2667.mask = 16'h0104;

	lut_sub lut_2675 ({n, m, k, g119, g178, g191}, g249);
	defparam lut_2675.LUT_SIZE = 6;
	defparam lut_2675.mask = 64'h0c0000000a000000;

	lut_sub lut_2686 ({k, g1, g247, g248, g249}, g250);
	defparam lut_2686.LUT_SIZE = 5;
	defparam lut_2686.mask = 32'h88808888;

	lut_sub lut_2701 ({g201, g243, g244, g246, g250}, g251);
	defparam lut_2701.LUT_SIZE = 5;
	defparam lut_2701.mask = 32'h11001000;

	lut_sub lut_2712 ({g236, g237, g190, g240, g251}, g252);
	defparam lut_2712.LUT_SIZE = 5;
	defparam lut_2712.mask = 32'h04050000;

	lut_sub lut_2720 ({h, g147, g525}, g253);
	defparam lut_2720.LUT_SIZE = 3;
	defparam lut_2720.mask = 8'h45;

	lut_sub lut_2727 ({h, g, j, k, g134}, g254);
	defparam lut_2727.LUT_SIZE = 5;
	defparam lut_2727.mask = 32'h0008a208;

	lut_sub lut_2738 ({j, l, g15, g253, g254}, g255);
	defparam lut_2738.LUT_SIZE = 5;
	defparam lut_2738.mask = 32'h0005000d;

	lut_sub lut_2746 ({m, k, l}, g256);
	defparam lut_2746.LUT_SIZE = 3;
	defparam lut_2746.mask = 8'h01;

	lut_sub lut_2753 ({j, k, g62, g532, g210}, g257);
	defparam lut_2753.LUT_SIZE = 5;
	defparam lut_2753.mask = 32'h0c0c0a00;

	lut_sub lut_2762 ({m, k, l}, g258);
	defparam lut_2762.LUT_SIZE = 3;
	defparam lut_2762.mask = 8'h10;

	lut_sub lut_2768 ({h, g, j, g62, g134}, g259);
	defparam lut_2768.LUT_SIZE = 5;
	defparam lut_2768.mask = 32'h00020000;

	lut_sub lut_2776 ({h, n, g58, g180, g258, g259}, g260);
	defparam lut_2776.LUT_SIZE = 6;
	defparam lut_2776.mask = 64'haaaa0000aaa80000;

	lut_sub lut_2799 ({g153, g133, g256, g257, g260}, g261);
	defparam lut_2799.LUT_SIZE = 5;
	defparam lut_2799.mask = 32'h40444040;

	lut_sub lut_2807 ({m, k, l}, g262);
	defparam lut_2807.LUT_SIZE = 3;
	defparam lut_2807.mask = 8'h40;

	lut_sub lut_2814 ({h, g58, g93, g504}, g263);
	defparam lut_2814.LUT_SIZE = 4;
	defparam lut_2814.mask = 16'h5554;

	lut_sub lut_2825 ({n, m, j, l, g225}, g264);
	defparam lut_2825.LUT_SIZE = 5;
	defparam lut_2825.mask = 32'h0000efff;

	lut_sub lut_2848 ({g247, g258, g262, g263, g264}, g265);
	defparam lut_2848.LUT_SIZE = 5;
	defparam lut_2848.mask = 32'h55115010;

	lut_sub lut_2863 ({j, i, g147, g151, g223}, g266);
	defparam lut_2863.LUT_SIZE = 5;
	defparam lut_2863.mask = 32'h44450000;

	lut_sub lut_2875 ({n, g64, g69, g147, g130}, g267);
	defparam lut_2875.LUT_SIZE = 5;
	defparam lut_2875.mask = 32'h03570000;

	lut_sub lut_2885 ({h, j, k, i}, g268);
	defparam lut_2885.LUT_SIZE = 4;
	defparam lut_2885.mask = 16'h513c;

	lut_sub lut_2898 ({n, m, l, g93, g180, g268}, g269);
	defparam lut_2898.LUT_SIZE = 6;
	defparam lut_2898.mask = 64'h0011000000050000;

	lut_sub lut_2908 ({f, g10, g2, g43}, g270);
	defparam lut_2908.LUT_SIZE = 4;
	defparam lut_2908.mask = 16'h0001;

	lut_sub lut_2916 ({g119, g270, g227, g262}, g271);
	defparam lut_2916.LUT_SIZE = 4;
	defparam lut_2916.mask = 16'hf0b0;

	lut_sub lut_2931 ({g227, g479, g267, g269, g271}, g272);
	defparam lut_2931.LUT_SIZE = 5;
	defparam lut_2931.mask = 32'h00404040;

	lut_sub lut_2942 ({g238, g258, g266, g215, g272}, g273);
	defparam lut_2942.LUT_SIZE = 5;
	defparam lut_2942.mask = 32'h10101000;

	lut_sub lut_2953 ({g255, g261, g265, g486, g273}, g274);
	defparam lut_2953.LUT_SIZE = 5;
	defparam lut_2953.mask = 32'h01110000;

	lut_sub lut_2961 ({g, g23, g54}, g275);
	defparam lut_2961.LUT_SIZE = 3;
	defparam lut_2961.mask = 8'h10;

	lut_sub lut_2967 ({f, h, g, g61, g63}, g276);
	defparam lut_2967.LUT_SIZE = 5;
	defparam lut_2967.mask = 32'h05010000;

	lut_sub lut_2976 ({f, h, g, g59, g64, g60}, g277);
	defparam lut_2976.LUT_SIZE = 6;
	defparam lut_2976.mask = 64'h005f335f00000000;

	lut_sub lut_2999 ({n, g65, g146, g276, g277}, g278);
	defparam lut_2999.LUT_SIZE = 5;
	defparam lut_2999.mask = 32'h777f0000;

	lut_sub lut_3017 ({g275, g278}, g279);
	defparam lut_3017.LUT_SIZE = 2;
	defparam lut_3017.mask = 4'b1000;

	lut_sub lut_3024 ({g54, g75, g114}, g280);
	defparam lut_3024.LUT_SIZE = 3;
	defparam lut_3024.mask = 8'h01;

	lut_sub lut_3028 ({d, c}, g281);
	defparam lut_3028.LUT_SIZE = 2;
	defparam lut_3028.mask = 4'b1000;

	lut_sub lut_3034 ({e, l, g9, g281}, g282);
	defparam lut_3034.LUT_SIZE = 4;
	defparam lut_3034.mask = 16'h0001;

	lut_sub lut_3041 ({g40, k, g86, g282}, g283);
	defparam lut_3041.LUT_SIZE = 4;
	defparam lut_3041.mask = 16'h0010;

	lut_sub lut_3048 ({h, n, g65, g87, g147}, g284);
	defparam lut_3048.LUT_SIZE = 5;
	defparam lut_3048.mask = 32'h11111511;

	lut_sub lut_3064 ({j, g71, g147, g166, g284}, g285);
	defparam lut_3064.LUT_SIZE = 5;
	defparam lut_3064.mask = 32'h88808888;

	lut_sub lut_3079 ({g245, g267, g280, g283, g285}, g286);
	defparam lut_3079.LUT_SIZE = 5;
	defparam lut_3079.mask = 32'h40000000;

	lut_sub lut_3086 ({d, f, a, g35, g80, g115}, g287);
	defparam lut_3086.LUT_SIZE = 6;
	defparam lut_3086.mask = 64'h0300070003000300;

	lut_sub lut_3102 ({g81, g68, g156, g472}, g288);
	defparam lut_3102.LUT_SIZE = 4;
	defparam lut_3102.mask = 16'h4044;

	lut_sub lut_3109 ({h, g, i, g9}, g289);
	defparam lut_3109.LUT_SIZE = 4;
	defparam lut_3109.mask = 16'h4000;

	lut_sub lut_3115 ({g135, g202}, g290);
	defparam lut_3115.LUT_SIZE = 2;
	defparam lut_3115.mask = 4'b0010;

	lut_sub lut_3122 ({k, l, g9, g289, g290}, g291);
	defparam lut_3122.LUT_SIZE = 5;
	defparam lut_3122.mask = 32'h37050505;

	lut_sub lut_3138 ({f, g281, g291}, g292);
	defparam lut_3138.LUT_SIZE = 3;
	defparam lut_3138.mask = 8'h10;

	lut_sub lut_3145 ({k, g41, g58, g282}, g293);
	defparam lut_3145.LUT_SIZE = 4;
	defparam lut_3145.mask = 16'h0001;

	lut_sub lut_3153 ({a, g97, g85, g292, g293}, g294);
	defparam lut_3153.LUT_SIZE = 5;
	defparam lut_3153.mask = 32'h88888880;

	lut_sub lut_3169 ({g155, g279, g286, g287, g288, g294}, g295);
	defparam lut_3169.LUT_SIZE = 6;
	defparam lut_3169.mask = 64'h0010001000000010;

	lut_sub lut_3177 ({d, e, a, g275, g278}, g296);
	defparam lut_3177.LUT_SIZE = 5;
	defparam lut_3177.mask = 32'h00070000;

	lut_sub lut_3184 ({h, g, i, g1, c}, g297);
	defparam lut_3184.LUT_SIZE = 5;
	defparam lut_3184.mask = 32'h01000000;

	lut_sub lut_3190 ({j, k, l, g105, g297}, g298);
	defparam lut_3190.LUT_SIZE = 5;
	defparam lut_3190.mask = 32'hc888cc88;

	lut_sub lut_3207 ({f, g, g47, g48, g81}, g299);
	defparam lut_3207.LUT_SIZE = 5;
	defparam lut_3207.mask = 32'h0a220000;

	lut_sub lut_3216 ({b, d, e, g298, g299}, g300);
	defparam lut_3216.LUT_SIZE = 5;
	defparam lut_3216.mask = 32'h0505050d;

	lut_sub lut_3229 ({b, d, f, g7}, g301);
	defparam lut_3229.LUT_SIZE = 4;
	defparam lut_3229.mask = 16'h0001;

	lut_sub lut_3237 ({b, g33, g34, g97, g104}, g302);
	defparam lut_3237.LUT_SIZE = 5;
	defparam lut_3237.mask = 32'h23220000;

	lut_sub lut_3247 ({e, l, g9, g97}, g303);
	defparam lut_3247.LUT_SIZE = 4;
	defparam lut_3247.mask = 16'h0100;

	lut_sub lut_3252 ({f, h, g, k, g58}, g304);
	defparam lut_3252.LUT_SIZE = 5;
	defparam lut_3252.mask = 32'h01000000;

	lut_sub lut_3259 ({h, g58, g34, g258}, g305);
	defparam lut_3259.LUT_SIZE = 4;
	defparam lut_3259.mask = 16'h0100;

	lut_sub lut_3267 ({f, g90, g303, g304, g305}, g306);
	defparam lut_3267.LUT_SIZE = 5;
	defparam lut_3267.mask = 32'h03570303;

	lut_sub lut_3282 ({d, e, l, g9, c}, g307);
	defparam lut_3282.LUT_SIZE = 5;
	defparam lut_3282.mask = 32'h00000002;

	lut_sub lut_3288 ({b, f, n, g76, g97}, g308);
	defparam lut_3288.LUT_SIZE = 5;
	defparam lut_3288.mask = 32'h01000000;

	lut_sub lut_3297 ({h, g58, g258, g304, g307, g308}, g309);
	defparam lut_3297.LUT_SIZE = 6;
	defparam lut_3297.mask = 64'h0303035703030303;

	lut_sub lut_3321 ({k, g86, g146}, g310);
	defparam lut_3321.LUT_SIZE = 3;
	defparam lut_3321.mask = 8'h10;

	lut_sub lut_3327 ({h, g86, g262}, g311);
	defparam lut_3327.LUT_SIZE = 3;
	defparam lut_3327.mask = 8'h01;

	lut_sub lut_3336 ({f, g34, g90, g303, g310, g311}, g312);
	defparam lut_3336.LUT_SIZE = 6;
	defparam lut_3336.mask = 64'h0303035703030303;

	lut_sub lut_3360 ({i, g9, g281}, g313);
	defparam lut_3360.LUT_SIZE = 3;
	defparam lut_3360.mask = 8'h10;

	lut_sub lut_3364 ({e, f, h, g}, g314);
	defparam lut_3364.LUT_SIZE = 4;
	defparam lut_3364.mask = 16'h8000;

	lut_sub lut_3370 ({k, l, g313, g314}, g315);
	defparam lut_3370.LUT_SIZE = 4;
	defparam lut_3370.mask = 16'h1000;

	lut_sub lut_3379 ({g46, g19, g158, g312, g315}, g316);
	defparam lut_3379.LUT_SIZE = 5;
	defparam lut_3379.mask = 32'h80000000;

	lut_sub lut_3385 ({k, l, g9, g99}, g317);
	defparam lut_3385.LUT_SIZE = 4;
	defparam lut_3385.mask = 16'h0001;

	lut_sub lut_3392 ({g, g23, g281, g317}, g318);
	defparam lut_3392.LUT_SIZE = 4;
	defparam lut_3392.mask = 16'h0100;

	lut_sub lut_3398 ({f, g76, g90}, g319);
	defparam lut_3398.LUT_SIZE = 3;
	defparam lut_3398.mask = 8'h01;

	lut_sub lut_3405 ({k, l, g41, g58, g20}, g320);
	defparam lut_3405.LUT_SIZE = 5;
	defparam lut_3405.mask = 32'h01000000;

	lut_sub lut_3410 ({h, k, l, g58}, g321);
	defparam lut_3410.LUT_SIZE = 4;
	defparam lut_3410.mask = 16'h4000;

	lut_sub lut_3417 ({n, m, g319, g320, g321}, g322);
	defparam lut_3417.LUT_SIZE = 5;
	defparam lut_3417.mask = 32'h37000500;

	lut_sub lut_3430 ({g31, g90, g75}, g323);
	defparam lut_3430.LUT_SIZE = 3;
	defparam lut_3430.mask = 8'h01;

	lut_sub lut_3434 ({b, d, c, a}, g324);
	defparam lut_3434.LUT_SIZE = 4;
	defparam lut_3434.mask = 16'h1504;

	lut_sub lut_3444 ({d, e, f, g113, g115, g324}, g325);
	defparam lut_3444.LUT_SIZE = 6;
	defparam lut_3444.mask = 64'h0003001300000011;

	lut_sub lut_3458 ({e, g318, g322, g323, g325}, g326);
	defparam lut_3458.LUT_SIZE = 5;
	defparam lut_3458.mask = 32'h80008080;

	lut_sub lut_3470 ({g37, g123, g306, g309, g316, g326}, g327);
	defparam lut_3470.LUT_SIZE = 6;
	defparam lut_3470.mask = 64'h1000100000001000;

	lut_sub lut_3482 ({g296, g300, g286, g301, g302, g327}, g328);
	defparam lut_3482.LUT_SIZE = 6;
	defparam lut_3482.mask = 64'h0040000000000000;

	lut_sub lut_3490 ({g310, g311, g307, g308}, g329);
	defparam lut_3490.LUT_SIZE = 4;
	defparam lut_3490.mask = 16'h0537;

	lut_sub lut_3500 ({j, k}, g330);
	defparam lut_3500.LUT_SIZE = 2;
	defparam lut_3500.mask = 4'b1000;

	lut_sub lut_3505 ({d, e, f, a, g35}, g331);
	defparam lut_3505.LUT_SIZE = 5;
	defparam lut_3505.mask = 32'h00000400;

	lut_sub lut_3514 ({l, g15, g330, g136, g293, g331}, g332);
	defparam lut_3514.LUT_SIZE = 6;
	defparam lut_3514.mask = 64'hccccccccccccccc8;

	lut_sub lut_3551 ({j, g10, g262, g308}, g333);
	defparam lut_3551.LUT_SIZE = 4;
	defparam lut_3551.mask = 16'h0001;

	lut_sub lut_3556 ({f, h, g, k, g99}, g334);
	defparam lut_3556.LUT_SIZE = 5;
	defparam lut_3556.mask = 32'h04000000;

	lut_sub lut_3564 ({g145, l, g15, g135, g331}, g335);
	defparam lut_3564.LUT_SIZE = 5;
	defparam lut_3564.mask = 32'h00000001;

	lut_sub lut_3573 ({g306, g307, g333, g334, g335}, g336);
	defparam lut_3573.LUT_SIZE = 5;
	defparam lut_3573.mask = 32'ha0800000;

	lut_sub lut_3581 ({f, l, g330, g281}, g337);
	defparam lut_3581.LUT_SIZE = 4;
	defparam lut_3581.mask = 16'h1000;

	lut_sub lut_3588 ({e, g289, g318, g337}, g338);
	defparam lut_3588.LUT_SIZE = 4;
	defparam lut_3588.mask = 16'h3705;

	lut_sub lut_3603 ({g312, g329, g332, g336, g338}, g339);
	defparam lut_3603.LUT_SIZE = 5;
	defparam lut_3603.mask = 32'h02000000;

	lut_sub lut_3609 ({a, g35, g82}, g340);
	defparam lut_3609.LUT_SIZE = 3;
	defparam lut_3609.mask = 8'h01;

	lut_sub lut_3616 ({g136, g203, g340}, g341);
	defparam lut_3616.LUT_SIZE = 3;
	defparam lut_3616.mask = 8'h01;

	lut_sub lut_3623 ({g182, g258, g319}, g342);
	defparam lut_3623.LUT_SIZE = 3;
	defparam lut_3623.mask = 8'h01;

	lut_sub lut_3632 ({g40, g20, g317, g309, g342}, g343);
	defparam lut_3632.LUT_SIZE = 5;
	defparam lut_3632.mask = 32'h88888880;

	lut_sub lut_3647 ({g312, g329, g332, g341, g343}, g344);
	defparam lut_3647.LUT_SIZE = 5;
	defparam lut_3647.mask = 32'h04000000;

	lut_sub lut_3654 ({e, g318, g315, g344}, g345);
	defparam lut_3654.LUT_SIZE = 4;
	defparam lut_3654.mask = 16'h4440;

	lut_sub lut_3662 ({h, g, a, g36, g223}, g346);
	defparam lut_3662.LUT_SIZE = 5;
	defparam lut_3662.mask = 32'h00ef00ff;

	lut_sub lut_3681 ({b, h, n, k, g97}, g347);
	defparam lut_3681.LUT_SIZE = 5;
	defparam lut_3681.mask = 32'h00440040;

	lut_sub lut_3688 ({g, m, l, g347}, g348);
	defparam lut_3688.LUT_SIZE = 4;
	defparam lut_3688.mask = 16'hef00;

	lut_sub lut_3698 ({e, f, j, i}, g349);
	defparam lut_3698.LUT_SIZE = 4;
	defparam lut_3698.mask = 16'h8000;

	lut_sub lut_3707 ({g322, g346, g348, g283, g349}, g350);
	defparam lut_3707.LUT_SIZE = 5;
	defparam lut_3707.mask = 32'h8ccc0000;

	lut_sub lut_3721 ({g292, g336, g344, g350}, g351);
	defparam lut_3721.LUT_SIZE = 4;
	defparam lut_3721.mask = 16'h0100;

	lut_sub lut_3727 ({h, k, l, g9, g99}, g352);
	defparam lut_3727.LUT_SIZE = 5;
	defparam lut_3727.mask = 32'h11000001;

	lut_sub lut_3733 ({h, j, k, i}, g353);
	defparam lut_3733.LUT_SIZE = 4;
	defparam lut_3733.mask = 16'h0040;

	lut_sub lut_3739 ({g15, g353}, g354);
	defparam lut_3739.LUT_SIZE = 2;
	defparam lut_3739.mask = 4'b0001;

	lut_sub lut_3745 ({e, g, g1, g281}, g355);
	defparam lut_3745.LUT_SIZE = 4;
	defparam lut_3745.mask = 16'h0e0f;

	lut_sub lut_3755 ({e, h, m, i, c}, g356);
	defparam lut_3755.LUT_SIZE = 5;
	defparam lut_3755.mask = 32'h80000000;

	lut_sub lut_3760 ({b, e, h, i, g1}, g357);
	defparam lut_3760.LUT_SIZE = 5;
	defparam lut_3760.mask = 32'h40000000;

	lut_sub lut_3769 ({g35, g182, g223, g356, g357}, g358);
	defparam lut_3769.LUT_SIZE = 5;
	defparam lut_3769.mask = 32'h88808888;

	lut_sub lut_3782 ({f, g313, g355, g358}, g359);
	defparam lut_3782.LUT_SIZE = 4;
	defparam lut_3782.mask = 16'h1011;

	lut_sub lut_3792 ({d, a, g35, g352, g354, g359}, g360);
	defparam lut_3792.LUT_SIZE = 6;
	defparam lut_3792.mask = 64'h4040404044554444;

	lut_sub lut_3809 ({e, f, c}, g361);
	defparam lut_3809.LUT_SIZE = 3;
	defparam lut_3809.mask = 8'h40;

	lut_sub lut_3816 ({e, f, g145, a, g15, g90}, g362);
	defparam lut_3816.LUT_SIZE = 6;
	defparam lut_3816.mask = 64'h0033002300330033;

	lut_sub lut_3835 ({g9, c}, g363);
	defparam lut_3835.LUT_SIZE = 2;
	defparam lut_3835.mask = 4'b0001;

	lut_sub lut_3842 ({h, i, g281, g317, g363}, g364);
	defparam lut_3842.LUT_SIZE = 5;
	defparam lut_3842.mask = 32'h55003030;

	lut_sub lut_3856 ({h, g, g54, g362, g364}, g365);
	defparam lut_3856.LUT_SIZE = 5;
	defparam lut_3856.mask = 32'h80008800;

	lut_sub lut_3866 ({i, g9, g330, g361, g365}, g366);
	defparam lut_3866.LUT_SIZE = 5;
	defparam lut_3866.mask = 32'h55455544;

	lut_sub lut_3883 ({b, d, e, l, c, g330}, g367);
	defparam lut_3883.LUT_SIZE = 6;
	defparam lut_3883.mask = 64'h0105010100ff0033;

	lut_sub lut_3904 ({e, c, g90}, g368);
	defparam lut_3904.LUT_SIZE = 3;
	defparam lut_3904.mask = 8'h10;

	lut_sub lut_3909 ({b, h, j, k, i, g368}, g369);
	defparam lut_3909.LUT_SIZE = 6;
	defparam lut_3909.mask = 64'h5511055555310555;

	lut_sub lut_3940 ({g, g1, g367, g369}, g370);
	defparam lut_3940.LUT_SIZE = 4;
	defparam lut_3940.mask = 16'h0d05;

	lut_sub lut_3950 ({d, a, g15, g212}, g371);
	defparam lut_3950.LUT_SIZE = 4;
	defparam lut_3950.mask = 16'h0111;

	lut_sub lut_3958 ({i, l, g1, g371}, g372);
	defparam lut_3958.LUT_SIZE = 4;
	defparam lut_3958.mask = 16'h8aaa;

	lut_sub lut_3968 ({b, h, k, i}, g373);
	defparam lut_3968.LUT_SIZE = 4;
	defparam lut_3968.mask = 16'h88a0;

	lut_sub lut_3978 ({e, g1, c, g352, g373}, g374);
	defparam lut_3978.LUT_SIZE = 5;
	defparam lut_3978.mask = 32'h03030357;

	lut_sub lut_3995 ({f, h, g370, g372, g374}, g375);
	defparam lut_3995.LUT_SIZE = 5;
	defparam lut_3995.mask = 32'hdf5f0000;

	lut_sub lut_4012 ({b, k, l, g1}, g376);
	defparam lut_4012.LUT_SIZE = 4;
	defparam lut_4012.mask = 16'h5515;

	lut_sub lut_4024 ({h, n, i, g64, g376}, g377);
	defparam lut_4024.LUT_SIZE = 5;
	defparam lut_4024.mask = 32'h70500000;

	lut_sub lut_4034 ({e, g, n, m, g281, g353}, g378);
	defparam lut_4034.LUT_SIZE = 6;
	defparam lut_4034.mask = 64'h7000400070304000;

	lut_sub lut_4047 ({d, e, h, k, a}, g379);
	defparam lut_4047.LUT_SIZE = 5;
	defparam lut_4047.mask = 32'h0000a200;

	lut_sub lut_4054 ({d, e, i, a, g35}, g380);
	defparam lut_4054.LUT_SIZE = 5;
	defparam lut_4054.mask = 32'h1100c000;

	lut_sub lut_4065 ({b, g15, g281, g379, g380}, g381);
	defparam lut_4065.LUT_SIZE = 5;
	defparam lut_4065.mask = 32'h007f0077;

	lut_sub lut_4084 ({k, l, g182, g462, g381}, g382);
	defparam lut_4084.LUT_SIZE = 5;
	defparam lut_4084.mask = 32'haaaaaaa8;

	lut_sub lut_4104 ({h, k, g34, g99}, g383);
	defparam lut_4104.LUT_SIZE = 4;
	defparam lut_4104.mask = 16'h1000;

	lut_sub lut_4110 ({g57, g20}, g384);
	defparam lut_4110.LUT_SIZE = 2;
	defparam lut_4110.mask = 4'b0001;

	lut_sub lut_4115 ({j, k, i, l, g384}, g385);
	defparam lut_4115.LUT_SIZE = 5;
	defparam lut_4115.mask = 32'h15551454;

	lut_sub lut_4133 ({g, l, g211, g281, g361}, g386);
	defparam lut_4133.LUT_SIZE = 5;
	defparam lut_4133.mask = 32'h55507750;

	lut_sub lut_4150 ({h, g, j, k, i}, g387);
	defparam lut_4150.LUT_SIZE = 5;
	defparam lut_4150.mask = 32'h5051001f;

	lut_sub lut_4163 ({e, f, g, j, l, c}, g388);
	defparam lut_4163.LUT_SIZE = 6;
	defparam lut_4163.mask = 64'h00f8ffff00f800f8;

	lut_sub lut_4200 ({h, g40, i, g20, g388}, g389);
	defparam lut_4200.LUT_SIZE = 5;
	defparam lut_4200.mask = 32'h50700030;

	lut_sub lut_4212 ({e, f, c, g387, g389}, g390);
	defparam lut_4212.LUT_SIZE = 5;
	defparam lut_4212.mask = 32'ha8aa8aaa;

	lut_sub lut_4234 ({g9, g383, g385, g386, g390}, g391);
	defparam lut_4234.LUT_SIZE = 5;
	defparam lut_4234.mask = 32'h0000bfff;

	lut_sub lut_4256 ({f, g377, g378, g382, g391}, g392);
	defparam lut_4256.LUT_SIZE = 5;
	defparam lut_4256.mask = 32'haaaa2000;

	lut_sub lut_4270 ({f, m, g145, g10}, g393);
	defparam lut_4270.LUT_SIZE = 4;
	defparam lut_4270.mask = 16'h0010;

	lut_sub lut_4274 ({g, m, j, i, l}, g394);
	defparam lut_4274.LUT_SIZE = 5;
	defparam lut_4274.mask = 32'h3000e000;

	lut_sub lut_4284 ({h, k, g393, g394}, g395);
	defparam lut_4284.LUT_SIZE = 4;
	defparam lut_4284.mask = 16'hcc8c;

	lut_sub lut_4296 ({d, e, l, g57, g182}, g396);
	defparam lut_4296.LUT_SIZE = 5;
	defparam lut_4296.mask = 32'h01010100;

	lut_sub lut_4304 ({m, j, k, g340, g396}, g397);
	defparam lut_4304.LUT_SIZE = 5;
	defparam lut_4304.mask = 32'h00000705;

	lut_sub lut_4312 ({d, f, h, g, k, c}, g398);
	defparam lut_4312.LUT_SIZE = 6;
	defparam lut_4312.mask = 64'h0c080808ac00aa00;

	lut_sub lut_4328 ({e, f, h, g, c}, g399);
	defparam lut_4328.LUT_SIZE = 5;
	defparam lut_4328.mask = 32'h08005a00;

	lut_sub lut_4338 ({m, i, g398, g399}, g400);
	defparam lut_4338.LUT_SIZE = 4;
	defparam lut_4338.mask = 16'h7000;

	lut_sub lut_4346 ({g44, g, m, g330}, g401);
	defparam lut_4346.LUT_SIZE = 4;
	defparam lut_4346.mask = 16'h0040;

	lut_sub lut_4350 ({h, j, k, i, l}, g402);
	defparam lut_4350.LUT_SIZE = 5;
	defparam lut_4350.mask = 32'h808080b3;

	lut_sub lut_4362 ({f, g, m, c, g402}, g403);
	defparam lut_4362.LUT_SIZE = 5;
	defparam lut_4362.mask = 32'h80000000;

	lut_sub lut_4368 ({f, m, g86, g281}, g404);
	defparam lut_4368.LUT_SIZE = 4;
	defparam lut_4368.mask = 16'h1000;

	lut_sub lut_4377 ({g193, g384, g401, g403, g404}, g405);
	defparam lut_4377.LUT_SIZE = 5;
	defparam lut_4377.mask = 32'h80808000;

	lut_sub lut_4384 ({d, e, f, a, g35}, g406);
	defparam lut_4384.LUT_SIZE = 5;
	defparam lut_4384.mask = 32'hf000cc01;

	lut_sub lut_4398 ({g, m, g145, g406}, g407);
	defparam lut_4398.LUT_SIZE = 4;
	defparam lut_4398.mask = 16'h0400;

	lut_sub lut_4407 ({g395, g397, g400, g405, g407}, g408);
	defparam lut_4407.LUT_SIZE = 5;
	defparam lut_4407.mask = 32'h00002000;

	lut_sub lut_4411 ({d, e, f, a}, g409);
	defparam lut_4411.LUT_SIZE = 4;
	defparam lut_4411.mask = 16'hc080;

	lut_sub lut_4417 ({b, e, f}, g410);
	defparam lut_4417.LUT_SIZE = 3;
	defparam lut_4417.mask = 8'h20;

	lut_sub lut_4423 ({g1, g410}, g411);
	defparam lut_4423.LUT_SIZE = 2;
	defparam lut_4423.mask = 4'b0001;

	lut_sub lut_4429 ({b, e, j, k, g1, g97}, g412);
	defparam lut_4429.LUT_SIZE = 6;
	defparam lut_4429.mask = 64'h2000200020003000;

	lut_sub lut_4441 ({j, g15, g409, g411, g412}, g413);
	defparam lut_4441.LUT_SIZE = 5;
	defparam lut_4441.mask = 32'haaa08880;

	lut_sub lut_4453 ({d, e, f}, g414);
	defparam lut_4453.LUT_SIZE = 3;
	defparam lut_4453.mask = 8'h0d;

	lut_sub lut_4459 ({b, e, n, i, c}, g415);
	defparam lut_4459.LUT_SIZE = 5;
	defparam lut_4459.mask = 32'h23002000;

	lut_sub lut_4470 ({m, g330, g414, g363, g415}, g416);
	defparam lut_4470.LUT_SIZE = 5;
	defparam lut_4470.mask = 32'h00750030;

	lut_sub lut_4482 ({n, m, j, i, g97, g61}, g417);
	defparam lut_4482.LUT_SIZE = 6;
	defparam lut_4482.mask = 64'h50005000c0c00000;

	lut_sub lut_4493 ({h, n, k, i, l}, g418);
	defparam lut_4493.LUT_SIZE = 5;
	defparam lut_4493.mask = 32'hdfff0000;

	lut_sub lut_4512 ({d, j, i, g9, c}, g419);
	defparam lut_4512.LUT_SIZE = 5;
	defparam lut_4512.mask = 32'h12100000;

	lut_sub lut_4522 ({j, g411, g417, g418, g419}, g420);
	defparam lut_4522.LUT_SIZE = 5;
	defparam lut_4522.mask = 32'h20002020;

	lut_sub lut_4529 ({b, e, f, g, g145}, g421);
	defparam lut_4529.LUT_SIZE = 5;
	defparam lut_4529.mask = 32'hd1c01100;

	lut_sub lut_4543 ({g, k, l, g1, g58, g421}, g422);
	defparam lut_4543.LUT_SIZE = 6;
	defparam lut_4543.mask = 64'h0f0505050d050505;

	lut_sub lut_4570 ({h, g313, g413, g416, g420, g422}, g423);
	defparam lut_4570.LUT_SIZE = 6;
	defparam lut_4570.mask = 64'h2222222222f22222;

	lut_sub lut_4593 ({b, d, c, g410}, g424);
	defparam lut_4593.LUT_SIZE = 4;
	defparam lut_4593.mask = 16'hdc50;

	lut_sub lut_4607 ({j, g1, g290, g319, g424}, g425);
	defparam lut_4607.LUT_SIZE = 5;
	defparam lut_4607.mask = 32'h007f005f;

	lut_sub lut_4625 ({g44, j, k, g1}, g426);
	defparam lut_4625.LUT_SIZE = 4;
	defparam lut_4625.mask = 16'h0040;

	lut_sub lut_4629 ({b, e, f, c, a}, g427);
	defparam lut_4629.LUT_SIZE = 5;
	defparam lut_4629.mask = 32'hb0008000;

	lut_sub lut_4640 ({h, k, g15, g340, g426, g427}, g428);
	defparam lut_4640.LUT_SIZE = 6;
	defparam lut_4640.mask = 64'hcc80cc80cc80cc88;

	lut_sub lut_4665 ({d, e, g, g145}, g429);
	defparam lut_4665.LUT_SIZE = 4;
	defparam lut_4665.mask = 16'h0010;

	lut_sub lut_4672 ({i, a, g35, g82, g429}, g430);
	defparam lut_4672.LUT_SIZE = 5;
	defparam lut_4672.mask = 32'h55035500;

	lut_sub lut_4686 ({f, h, g, g409}, g431);
	defparam lut_4686.LUT_SIZE = 4;
	defparam lut_4686.mask = 16'h2aaa;

	lut_sub lut_4698 ({j, l, g406, g431}, g432);
	defparam lut_4698.LUT_SIZE = 4;
	defparam lut_4698.mask = 16'h30ba;

	lut_sub lut_4708 ({f, h, g}, g433);
	defparam lut_4708.LUT_SIZE = 3;
	defparam lut_4708.mask = 8'h08;

	lut_sub lut_4713 ({b, l, a, g330}, g434);
	defparam lut_4713.LUT_SIZE = 4;
	defparam lut_4713.mask = 16'hdc50;

	lut_sub lut_4725 ({e, f, h, g, g212, g353}, g435);
	defparam lut_4725.LUT_SIZE = 6;
	defparam lut_4725.mask = 64'h0000000037050505;

	lut_sub lut_4743 ({d, c, g433, g410, g434, g435}, g436);
	defparam lut_4743.LUT_SIZE = 6;
	defparam lut_4743.mask = 64'h8800880080008800;

	lut_sub lut_4756 ({g99, g146, g223}, g437);
	defparam lut_4756.LUT_SIZE = 3;
	defparam lut_4756.mask = 8'h01;

	lut_sub lut_4764 ({h, g58, g34, g71, g317}, g438);
	defparam lut_4764.LUT_SIZE = 5;
	defparam lut_4764.mask = 32'h00330505;

	lut_sub lut_4781 ({g15, g430, g432, g436, g437, g438}, g439);
	defparam lut_4781.LUT_SIZE = 6;
	defparam lut_4781.mask = 64'h8888888808000000;

	lut_sub lut_4798 ({n, g408, g423, g425, g428, g439}, g440);
	defparam lut_4798.LUT_SIZE = 6;
	defparam lut_4798.mask = 64'h0000001000100010;

	lut_sub lut_4806 ({g, j, g281, g361}, g441);
	defparam lut_4806.LUT_SIZE = 4;
	defparam lut_4806.mask = 16'h0507;

	lut_sub lut_4818 ({g41, g9, g20, g441}, g442);
	defparam lut_4818.LUT_SIZE = 4;
	defparam lut_4818.mask = 16'h0507;

	lut_sub lut_4828 ({k, l, g1, g319}, g443);
	defparam lut_4828.LUT_SIZE = 4;
	defparam lut_4828.mask = 16'h1110;

	lut_sub lut_4837 ({h, g1, c, g82, g202}, g444);
	defparam lut_4837.LUT_SIZE = 5;
	defparam lut_4837.mask = 32'h000000a8;

	lut_sub lut_4844 ({f, g, k, g9, c}, g445);
	defparam lut_4844.LUT_SIZE = 5;
	defparam lut_4844.mask = 32'h20000000;

	lut_sub lut_4850 ({n, g218, g281}, g446);
	defparam lut_4850.LUT_SIZE = 3;
	defparam lut_4850.mask = 8'h10;

	lut_sub lut_4859 ({g443, g444, g445, g446, g456}, g447);
	defparam lut_4859.LUT_SIZE = 5;
	defparam lut_4859.mask = 32'h40000000;

	lut_sub lut_4863 ({h, k, i, l}, g448);
	defparam lut_4863.LUT_SIZE = 4;
	defparam lut_4863.mask = 16'h8033;

	lut_sub lut_4873 ({m, k, g58, g410}, g449);
	defparam lut_4873.LUT_SIZE = 4;
	defparam lut_4873.mask = 16'h0400;

	lut_sub lut_4881 ({m, g319, g395, g448, g449}, g450);
	defparam lut_4881.LUT_SIZE = 5;
	defparam lut_4881.mask = 32'h0a020a0a;

	lut_sub lut_4894 ({n, i, g442, g447, g450}, g451);
	defparam lut_4894.LUT_SIZE = 5;
	defparam lut_4894.mask = 32'hff305510;

	lut_sub lut_4918 ({g360, g366, g375, g392, g440, g451}, l2);
	defparam lut_4918.LUT_SIZE = 6;
	defparam lut_4918.mask = 64'hfffffefffefffeff;

	lut_sub lut_4983 ({h, k, j, g15, l}, g453);
	defparam lut_4983.LUT_SIZE = 5;
	defparam lut_4983.mask = 32'h00001033;

	lut_sub lut_4992 ({h, i, k, j, g15, l}, g454);
	defparam lut_4992.LUT_SIZE = 6;
	defparam lut_4992.mask = 64'h0321113313330332;

	lut_sub lut_5019 ({g453, g454, g}, g455);
	defparam lut_5019.LUT_SIZE = 3;
	defparam lut_5019.mask = 8'he4;

	lut_sub lut_5027 ({n, g457}, g456);
	defparam lut_5027.LUT_SIZE = 2;
	defparam lut_5027.mask = 4'b1000;

	lut_sub lut_5032 ({n, g458}, g457);
	defparam lut_5032.LUT_SIZE = 2;
	defparam lut_5032.mask = 4'b0100;

	lut_sub lut_5038 ({g459, g460}, g458);
	defparam lut_5038.LUT_SIZE = 2;
	defparam lut_5038.mask = 4'b1000;

	lut_sub lut_5043 ({m, g461}, g459);
	defparam lut_5043.LUT_SIZE = 2;
	defparam lut_5043.mask = 4'b0100;

	lut_sub lut_5048 ({m, g431}, g460);
	defparam lut_5048.LUT_SIZE = 2;
	defparam lut_5048.mask = 4'b0001;

	lut_sub lut_5053 ({g34, c, l, f}, g461);
	defparam lut_5053.LUT_SIZE = 4;
	defparam lut_5053.mask = 16'h7fff;

	lut_sub lut_5073 ({g463, g464}, g462);
	defparam lut_5073.LUT_SIZE = 2;
	defparam lut_5073.mask = 4'b1000;

	lut_sub lut_5078 ({a, g465}, g463);
	defparam lut_5078.LUT_SIZE = 2;
	defparam lut_5078.mask = 4'b0100;

	lut_sub lut_5083 ({a, g468}, g464);
	defparam lut_5083.LUT_SIZE = 2;
	defparam lut_5083.mask = 4'b0001;

	lut_sub lut_5089 ({g466, g467}, g465);
	defparam lut_5089.LUT_SIZE = 2;
	defparam lut_5089.mask = 4'b1000;

	lut_sub lut_5094 ({m, g469}, g466);
	defparam lut_5094.LUT_SIZE = 2;
	defparam lut_5094.mask = 4'b0100;

	lut_sub lut_5099 ({m, g470}, g467);
	defparam lut_5099.LUT_SIZE = 2;
	defparam lut_5099.mask = 4'b0001;

	lut_sub lut_5104 ({m, g471}, g468);
	defparam lut_5104.LUT_SIZE = 2;
	defparam lut_5104.mask = 4'b0100;

	lut_sub lut_5108 ({c, l, b, n}, g469);
	defparam lut_5108.LUT_SIZE = 4;
	defparam lut_5108.mask = 16'hce44;

	lut_sub lut_5118 ({g, n}, g470);
	defparam lut_5118.LUT_SIZE = 2;
	defparam lut_5118.mask = 4'b0010;

	lut_sub lut_5122 ({c, l, b, n}, g471);
	defparam lut_5122.LUT_SIZE = 4;
	defparam lut_5122.mask = 16'hce44;

	lut_sub lut_5133 ({f, g473}, g472);
	defparam lut_5133.LUT_SIZE = 2;
	defparam lut_5133.mask = 4'b1000;

	lut_sub lut_5138 ({f, g474}, g473);
	defparam lut_5138.LUT_SIZE = 2;
	defparam lut_5138.mask = 4'b0100;

	lut_sub lut_5144 ({g475, g476}, g474);
	defparam lut_5144.LUT_SIZE = 2;
	defparam lut_5144.mask = 4'b1000;

	lut_sub lut_5149 ({g, g477}, g475);
	defparam lut_5149.LUT_SIZE = 2;
	defparam lut_5149.mask = 4'b0100;

	lut_sub lut_5154 ({g, g478}, g476);
	defparam lut_5154.LUT_SIZE = 2;
	defparam lut_5154.mask = 4'b0001;

	lut_sub lut_5160 ({g35, a, g47, d}, g477);
	defparam lut_5160.LUT_SIZE = 4;
	defparam lut_5160.mask = 16'hfffe;

	lut_sub lut_5180 ({g35, a, g48, d}, g478);
	defparam lut_5180.LUT_SIZE = 4;
	defparam lut_5180.mask = 16'hfffe;

	lut_sub lut_5199 ({m, g480}, g479);
	defparam lut_5199.LUT_SIZE = 2;
	defparam lut_5199.mask = 4'b1000;

	lut_sub lut_5204 ({m, g481}, g480);
	defparam lut_5204.LUT_SIZE = 2;
	defparam lut_5204.mask = 4'b0100;

	lut_sub lut_5210 ({g482, g483}, g481);
	defparam lut_5210.LUT_SIZE = 2;
	defparam lut_5210.mask = 4'b1000;

	lut_sub lut_5215 ({h, g484}, g482);
	defparam lut_5215.LUT_SIZE = 2;
	defparam lut_5215.mask = 4'b0100;

	lut_sub lut_5220 ({h, g485}, g483);
	defparam lut_5220.LUT_SIZE = 2;
	defparam lut_5220.mask = 4'b0001;

	lut_sub lut_5224 ({g, l, i, j}, g484);
	defparam lut_5224.LUT_SIZE = 4;
	defparam lut_5224.mask = 16'hfffd;

	lut_sub lut_5242 ({g, l, k, j}, g485);
	defparam lut_5242.LUT_SIZE = 4;
	defparam lut_5242.mask = 16'hfffd;

	lut_sub lut_5262 ({g487, g488}, g486);
	defparam lut_5262.LUT_SIZE = 2;
	defparam lut_5262.mask = 4'b1000;

	lut_sub lut_5268 ({g211, g489}, g487);
	defparam lut_5268.LUT_SIZE = 2;
	defparam lut_5268.mask = 4'b0100;

	lut_sub lut_5274 ({g211, g492}, g488);
	defparam lut_5274.LUT_SIZE = 2;
	defparam lut_5274.mask = 4'b0001;

	lut_sub lut_5280 ({g490, g491}, g489);
	defparam lut_5280.LUT_SIZE = 2;
	defparam lut_5280.mask = 4'b1000;

	lut_sub lut_5285 ({n, g494}, g490);
	defparam lut_5285.LUT_SIZE = 2;
	defparam lut_5285.mask = 4'b0100;

	lut_sub lut_5290 ({n, g495}, g491);
	defparam lut_5290.LUT_SIZE = 2;
	defparam lut_5290.mask = 4'b0001;

	lut_sub lut_5295 ({n, g493}, g492);
	defparam lut_5295.LUT_SIZE = 2;
	defparam lut_5295.mask = 4'b0010;

	lut_sub lut_5300 ({n, g496}, g493);
	defparam lut_5300.LUT_SIZE = 2;
	defparam lut_5300.mask = 4'b0001;

	lut_sub lut_5306 ({m, g202, g178}, g494);
	defparam lut_5306.LUT_SIZE = 3;
	defparam lut_5306.mask = 8'h7f;

	lut_sub lut_5319 ({m, g202, g497, g191}, g495);
	defparam lut_5319.LUT_SIZE = 4;
	defparam lut_5319.mask = 16'h1fff;

	lut_sub lut_5337 ({m, g202, g497}, g496);
	defparam lut_5337.LUT_SIZE = 3;
	defparam lut_5337.mask = 8'h7f;

	lut_sub lut_5348 ({h, g498}, g497);
	defparam lut_5348.LUT_SIZE = 2;
	defparam lut_5348.mask = 4'b0010;

	lut_sub lut_5353 ({h, g499}, g498);
	defparam lut_5353.LUT_SIZE = 2;
	defparam lut_5353.mask = 4'b0001;

	lut_sub lut_5359 ({g500, g501}, g499);
	defparam lut_5359.LUT_SIZE = 2;
	defparam lut_5359.mask = 4'b1000;

	lut_sub lut_5364 ({f, g502}, g500);
	defparam lut_5364.LUT_SIZE = 2;
	defparam lut_5364.mask = 4'b0100;

	lut_sub lut_5369 ({f, g503}, g501);
	defparam lut_5369.LUT_SIZE = 2;
	defparam lut_5369.mask = 4'b0001;

	lut_sub lut_5375 ({g176, g, g39, i}, g502);
	defparam lut_5375.LUT_SIZE = 4;
	defparam lut_5375.mask = 16'h5777;

	lut_sub lut_5391 ({g176, g, g43, i}, g503);
	defparam lut_5391.LUT_SIZE = 4;
	defparam lut_5391.mask = 16'h5ddd;

	lut_sub lut_5406 ({h, g505}, g504);
	defparam lut_5406.LUT_SIZE = 2;
	defparam lut_5406.mask = 4'b0010;

	lut_sub lut_5411 ({h, g506}, g505);
	defparam lut_5411.LUT_SIZE = 2;
	defparam lut_5411.mask = 4'b0001;

	lut_sub lut_5417 ({g507, g508}, g506);
	defparam lut_5417.LUT_SIZE = 2;
	defparam lut_5417.mask = 4'b1000;

	lut_sub lut_5422 ({f, g509}, g507);
	defparam lut_5422.LUT_SIZE = 2;
	defparam lut_5422.mask = 4'b0100;

	lut_sub lut_5427 ({f, g510}, g508);
	defparam lut_5427.LUT_SIZE = 2;
	defparam lut_5427.mask = 4'b0001;

	lut_sub lut_5433 ({g176, j, g39, g}, g509);
	defparam lut_5433.LUT_SIZE = 4;
	defparam lut_5433.mask = 16'h1f3f;

	lut_sub lut_5449 ({g176, j, g43, g}, g510);
	defparam lut_5449.LUT_SIZE = 4;
	defparam lut_5449.mask = 16'h4fcf;

	lut_sub lut_5465 ({g15, g512}, g511);
	defparam lut_5465.LUT_SIZE = 2;
	defparam lut_5465.mask = 4'b0010;

	lut_sub lut_5471 ({g15, g513}, g512);
	defparam lut_5471.LUT_SIZE = 2;
	defparam lut_5471.mask = 4'b0001;

	lut_sub lut_5477 ({g514, g515}, g513);
	defparam lut_5477.LUT_SIZE = 2;
	defparam lut_5477.mask = 4'b1000;

	lut_sub lut_5482 ({l, g516}, g514);
	defparam lut_5482.LUT_SIZE = 2;
	defparam lut_5482.mask = 4'b0100;

	lut_sub lut_5487 ({l, g517}, g515);
	defparam lut_5487.LUT_SIZE = 2;
	defparam lut_5487.mask = 4'b0001;

	lut_sub lut_5492 ({i, g134, k, g}, g516);
	defparam lut_5492.LUT_SIZE = 4;
	defparam lut_5492.mask = 16'hffef;

	lut_sub lut_5511 ({i, g134, h, g}, g517);
	defparam lut_5511.LUT_SIZE = 4;
	defparam lut_5511.mask = 16'hffbf;

	lut_sub lut_5530 ({j, g519}, g518);
	defparam lut_5530.LUT_SIZE = 2;
	defparam lut_5530.mask = 4'b0010;

	lut_sub lut_5535 ({j, g520}, g519);
	defparam lut_5535.LUT_SIZE = 2;
	defparam lut_5535.mask = 4'b0001;

	lut_sub lut_5541 ({g521, g522}, g520);
	defparam lut_5541.LUT_SIZE = 2;
	defparam lut_5541.mask = 4'b1000;

	lut_sub lut_5546 ({l, g523}, g521);
	defparam lut_5546.LUT_SIZE = 2;
	defparam lut_5546.mask = 4'b0100;

	lut_sub lut_5551 ({l, g524}, g522);
	defparam lut_5551.LUT_SIZE = 2;
	defparam lut_5551.mask = 4'b0001;

	lut_sub lut_5556 ({i, g149}, g523);
	defparam lut_5556.LUT_SIZE = 2;
	defparam lut_5556.mask = 4'b1101;

	lut_sub lut_5564 ({g147, i, g151, k}, g524);
	defparam lut_5564.LUT_SIZE = 4;
	defparam lut_5564.mask = 16'h7775;

	lut_sub lut_5579 ({h, g526}, g525);
	defparam lut_5579.LUT_SIZE = 2;
	defparam lut_5579.mask = 4'b1000;

	lut_sub lut_5584 ({h, g527}, g526);
	defparam lut_5584.LUT_SIZE = 2;
	defparam lut_5584.mask = 4'b0100;

	lut_sub lut_5590 ({g528, g529}, g527);
	defparam lut_5590.LUT_SIZE = 2;
	defparam lut_5590.mask = 4'b1000;

	lut_sub lut_5595 ({f, g530}, g528);
	defparam lut_5595.LUT_SIZE = 2;
	defparam lut_5595.mask = 4'b0100;

	lut_sub lut_5600 ({f, g531}, g529);
	defparam lut_5600.LUT_SIZE = 2;
	defparam lut_5600.mask = 4'b0001;

	lut_sub lut_5606 ({g, e, g131, g88}, g530);
	defparam lut_5606.LUT_SIZE = 4;
	defparam lut_5606.mask = 16'hff13;

	lut_sub lut_5622 ({g, e, g132, g88}, g531);
	defparam lut_5622.LUT_SIZE = 4;
	defparam lut_5622.mask = 16'hff13;

	lut_sub lut_5637 ({h, g533}, g532);
	defparam lut_5637.LUT_SIZE = 2;
	defparam lut_5637.mask = 4'b0010;

	lut_sub lut_5642 ({h, g534}, g533);
	defparam lut_5642.LUT_SIZE = 2;
	defparam lut_5642.mask = 4'b0001;

	lut_sub lut_5648 ({g535, g536}, g534);
	defparam lut_5648.LUT_SIZE = 2;
	defparam lut_5648.mask = 4'b1000;

	lut_sub lut_5653 ({f, g537}, g535);
	defparam lut_5653.LUT_SIZE = 2;
	defparam lut_5653.mask = 4'b0100;

	lut_sub lut_5658 ({f, g538}, g536);
	defparam lut_5658.LUT_SIZE = 2;
	defparam lut_5658.mask = 4'b0001;

	lut_sub lut_5664 ({g88, e, g131, g}, g537);
	defparam lut_5664.LUT_SIZE = 4;
	defparam lut_5664.mask = 16'h5777;

	lut_sub lut_5680 ({g88, e, g132, g}, g538);
	defparam lut_5680.LUT_SIZE = 4;
	defparam lut_5680.mask = 16'h5777;

	lut_sub lut_5696 ({g540, g541}, g539);
	defparam lut_5696.LUT_SIZE = 2;
	defparam lut_5696.mask = 4'b1000;

	lut_sub lut_5702 ({g101, g542}, g540);
	defparam lut_5702.LUT_SIZE = 2;
	defparam lut_5702.mask = 4'b0100;

	lut_sub lut_5708 ({g101, g545}, g541);
	defparam lut_5708.LUT_SIZE = 2;
	defparam lut_5708.mask = 4'b0001;

	lut_sub lut_5714 ({g543, g544}, g542);
	defparam lut_5714.LUT_SIZE = 2;
	defparam lut_5714.mask = 4'b1000;

	lut_sub lut_5719 ({e, g547}, g543);
	defparam lut_5719.LUT_SIZE = 2;
	defparam lut_5719.mask = 4'b0100;

	lut_sub lut_5724 ({e, g548}, g544);
	defparam lut_5724.LUT_SIZE = 2;
	defparam lut_5724.mask = 4'b0001;

	lut_sub lut_5729 ({e, g546}, g545);
	defparam lut_5729.LUT_SIZE = 2;
	defparam lut_5729.mask = 4'b0010;

	lut_sub lut_5734 ({e, g549}, g546);
	defparam lut_5734.LUT_SIZE = 2;
	defparam lut_5734.mask = 4'b0001;

	lut_sub lut_5738 ({c, d}, g547);
	defparam lut_5738.LUT_SIZE = 2;
	defparam lut_5738.mask = 4'b1110;

	lut_sub lut_5746 ({g81, f, g455, d}, g548);
	defparam lut_5746.LUT_SIZE = 4;
	defparam lut_5746.mask = 16'hbfff;

	lut_sub lut_5766 ({g81, f, g455, d}, g549);
	defparam lut_5766.LUT_SIZE = 4;
	defparam lut_5766.mask = 16'hbfff;


endmodule