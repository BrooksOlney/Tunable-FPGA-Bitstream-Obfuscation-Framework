`timescale 10ns/1ns
module alu4_orig (/* input clk, */ input n, input j, input k, input l, input i, input a, input e, input m, input b, input f, input c, input g, input d, input houtput wire o, output wire p, output wire q, output wire r, output wire s, output wire t, output wire u, output wire v);

//reg [13:0] inputs;
//reg [7:0] outputs;
//always @(posedge clk) inputs = {n, j, k, l, i, a, e, m, b, f, c, g, d, h};
//always @(posedge clk) outputs = {o, p, q, r, s, t, u, v};

	wire g163, g121, g179, g182, g1, g8, g11, g9, g10, g12, g7;
	wire g13, g15, g17, g14, g16, g18, g19, g20, g22, g23, g27;
	wire g28, g26, g29, g21, g24, g25, g30, g33, g34, g35, g32;
	wire g36, g2, g3, g4, g41, g42, g38, g39, g40, g43, g44;
	wire g45, g46, g47, g50, g51, g54, g55, g48, g49, g52, g206;
	wire g62, g63, g64, g65, g67, g68, g69, g60, g61, g66, g70;
	wire g71, g58, g59, g72, g76, g74, g75, g77, g31, g73, g78;
	wire g81, g83, g84, g85, g86, g82, g87, g88, g89, g90, g53;
	wire g57, g92, g93, g95, g96, g91, g94, g97, g99, g100, g102;
	wire g103, g104, g106, g111, g108, g109, g110, g112, g98, g101, g105;
	wire g107, g113, g114, g118, g122, g123, g125, g126, g129, g130, g127;
	wire g128, g131, g124, g132, g133, g134, g120, g135, g136, g138, g139;
	wire g141, g147, g148, g149, g144, g145, g146, g150, g152, g153, g154;
	wire g137, g140, g142, g143, g151, g155, g159, g157, g158, g160, g80;
	wire g115, g156, g161, g168, g171, g183, g173, g169, g170, g172, g174;
	wire g165, g166, g167, g175, g164, g176, g178, g180, g181, g184, g185;
	wire g186, g189, g187, g188, g190, g191, g192, g194, g195, g196, g199;
	wire g197, g198, g202, g203, g200, g201, g204, g205, g119, g116, g117;
	wire g207, g208, g209, g212, g210, g211, g215, g216, g213, g214, g217;
	wire g218, g56, g220, g221, g222, g225, g223, g224, g228, g229, g226;
	wire g227, g230, g231, g37, g5, g6;


	assign s = (((!g163)));
	assign t = (((g121)));
	assign v = (((!g179)));
	assign g1 = (((k) & (!l)));
	assign g2 = (((!k) & (!l) & (n) & (!i) & (j)) + ((!k) & (l) & (n) & (!i) & (j)) + ((k) & (!l) & (!n) & (i) & (j)) + ((k) & (!l) & (n) & (i) & (j)) + ((k) & (l) & (!n) & (i) & (!j)) + ((k) & (l) & (n) & (!i) & (j)));
	assign g3 = (((!k) & (!l) & (!n) & (!i) & (!j)) + ((!k) & (!l) & (!n) & (!i) & (j)) + ((!k) & (l) & (!n) & (!i) & (!j)));
	assign g4 = (((!k) & (!l) & (!n) & (i) & (!j)) + ((k) & (!l) & (n) & (i) & (!j)) + ((k) & (l) & (n) & (i) & (!j)));
	assign g5 = (((!k) & (!l) & (!i) & (!a) & (!e) & (g182)) + ((!k) & (!l) & (!i) & (!a) & (e) & (g182)) + ((!k) & (!l) & (!i) & (a) & (!e) & (g182)) + ((!k) & (!l) & (!i) & (a) & (e) & (g182)) + ((!k) & (!l) & (i) & (!a) & (!e) & (!g182)) + ((!k) & (!l) & (i) & (!a) & (e) & (!g182)) + ((!k) & (!l) & (i) & (a) & (!e) & (!g182)) + ((!k) & (!l) & (i) & (a) & (e) & (!g182)) + ((!k) & (l) & (!i) & (!a) & (!e) & (g182)) + ((!k) & (l) & (!i) & (!a) & (e) & (g182)) + ((!k) & (l) & (!i) & (a) & (!e) & (!g182)) + ((!k) & (l) & (!i) & (a) & (!e) & (g182)) + ((!k) & (l) & (!i) & (a) & (e) & (g182)) + ((!k) & (l) & (i) & (!a) & (e) & (!g182)) + ((!k) & (l) & (i) & (!a) & (e) & (g182)) + ((!k) & (l) & (i) & (a) & (!e) & (!g182)) + ((!k) & (l) & (i) & (a) & (!e) & (g182)) + ((k) & (!l) & (!i) & (!a) & (!e) & (!g182)) + ((k) & (!l) & (!i) & (!a) & (e) & (!g182)) + ((k) & (!l) & (!i) & (a) & (!e) & (!g182)) + ((k) & (!l) & (!i) & (a) & (e) & (!g182)) + ((k) & (!l) & (i) & (!a) & (!e) & (!g182)) + ((k) & (!l) & (i) & (!a) & (!e) & (g182)) + ((k) & (!l) & (i) & (a) & (!e) & (!g182)) + ((k) & (!l) & (i) & (a) & (!e) & (g182)) + ((k) & (l) & (!i) & (!a) & (!e) & (!g182)) + ((k) & (l) & (!i) & (!a) & (!e) & (g182)) + ((k) & (l) & (!i) & (!a) & (e) & (!g182)) + ((k) & (l) & (!i) & (!a) & (e) & (g182)) + ((k) & (l) & (!i) & (a) & (!e) & (!g182)) + ((k) & (l) & (!i) & (a) & (!e) & (g182)) + ((k) & (l) & (!i) & (a) & (e) & (!g182)) + ((k) & (l) & (!i) & (a) & (e) & (g182)) + ((k) & (l) & (i) & (!a) & (!e) & (g182)) + ((k) & (l) & (i) & (!a) & (e) & (g182)) + ((k) & (l) & (i) & (a) & (!e) & (!g182)) + ((k) & (l) & (i) & (a) & (!e) & (g182)) + ((k) & (l) & (i) & (a) & (e) & (g182)));
	assign g6 = (((!k) & (l) & (!i) & (!a) & (e) & (!g182)) + ((!k) & (l) & (!i) & (!a) & (e) & (g182)) + ((!k) & (l) & (!i) & (a) & (e) & (!g182)) + ((!k) & (l) & (!i) & (a) & (e) & (g182)) + ((k) & (!l) & (!i) & (!a) & (!e) & (!g182)) + ((k) & (!l) & (!i) & (!a) & (!e) & (g182)) + ((k) & (!l) & (i) & (a) & (!e) & (g182)) + ((k) & (!l) & (i) & (a) & (e) & (g182)) + ((k) & (l) & (!i) & (!a) & (e) & (!g182)) + ((k) & (l) & (!i) & (!a) & (e) & (g182)) + ((k) & (l) & (!i) & (a) & (e) & (!g182)) + ((k) & (l) & (!i) & (a) & (e) & (g182)) + ((k) & (l) & (i) & (a) & (!e) & (g182)) + ((k) & (l) & (i) & (a) & (e) & (g182)));
	assign g7 = (((n) & (i) & (!j) & (g1)));
	assign g8 = (((i) & (j)));
	assign g9 = (((n) & (g8) & (g1)));
	assign g10 = (((n) & (!i) & (!j) & (g1)));
	assign g11 = (((n) & (!i) & (j)));
	assign g12 = (((l) & (g11)));
	assign g13 = (((!a) & (!g182) & (!g9) & (!g10) & (!g12)) + ((!a) & (!g182) & (!g9) & (!g10) & (g12)) + ((!a) & (!g182) & (g9) & (!g10) & (!g12)) + ((!a) & (!g182) & (g9) & (!g10) & (g12)) + ((!a) & (g182) & (!g9) & (!g10) & (!g12)) + ((!a) & (g182) & (!g9) & (g10) & (!g12)) + ((!a) & (g182) & (g9) & (!g10) & (!g12)) + ((!a) & (g182) & (g9) & (g10) & (!g12)) + ((a) & (!g182) & (!g9) & (!g10) & (!g12)) + ((a) & (!g182) & (g9) & (!g10) & (!g12)) + ((a) & (g182) & (!g9) & (!g10) & (!g12)) + ((a) & (g182) & (!g9) & (g10) & (!g12)));
	assign g14 = (((!a) & (!e) & (!g7) & (g13)) + ((!a) & (!e) & (g7) & (g13)) + ((!a) & (e) & (!g7) & (g13)) + ((!a) & (e) & (g7) & (g13)) + ((a) & (!e) & (!g7) & (g13)) + ((a) & (!e) & (g7) & (g13)) + ((a) & (e) & (!g7) & (g13)));
	assign g15 = (((!k) & (g12)));
	assign g16 = (((!a) & (!e) & (g7) & (g13) & (!g15)) + ((!a) & (!e) & (g7) & (g13) & (g15)) + ((!a) & (e) & (g7) & (g13) & (!g15)) + ((!a) & (e) & (g7) & (g13) & (g15)) + ((a) & (!e) & (g7) & (g13) & (!g15)) + ((a) & (!e) & (g7) & (g13) & (g15)) + ((a) & (e) & (!g7) & (!g13) & (g15)) + ((a) & (e) & (!g7) & (g13) & (g15)) + ((a) & (e) & (g7) & (!g13) & (g15)) + ((a) & (e) & (g7) & (g13) & (g15)));
	assign g17 = (((!k) & (!i) & (j)));
	assign g18 = (((l) & (g17)));
	assign g19 = (((!l) & (!i) & (!j) & (a) & (!e) & (!g182)) + ((!l) & (!i) & (!j) & (a) & (!e) & (g182)) + ((!l) & (!i) & (!j) & (a) & (e) & (!g182)) + ((!l) & (!i) & (!j) & (a) & (e) & (g182)) + ((!l) & (!i) & (j) & (!a) & (!e) & (g182)) + ((!l) & (!i) & (j) & (!a) & (e) & (g182)) + ((!l) & (!i) & (j) & (a) & (!e) & (!g182)) + ((!l) & (!i) & (j) & (a) & (!e) & (g182)) + ((!l) & (!i) & (j) & (a) & (e) & (!g182)) + ((!l) & (!i) & (j) & (a) & (e) & (g182)) + ((!l) & (i) & (!j) & (!a) & (e) & (!g182)) + ((!l) & (i) & (!j) & (!a) & (e) & (g182)) + ((!l) & (i) & (!j) & (a) & (!e) & (!g182)) + ((!l) & (i) & (!j) & (a) & (!e) & (g182)) + ((l) & (!i) & (!j) & (a) & (!e) & (!g182)) + ((l) & (!i) & (!j) & (a) & (e) & (!g182)) + ((l) & (i) & (!j) & (!a) & (e) & (!g182)) + ((l) & (i) & (!j) & (!a) & (e) & (g182)) + ((l) & (i) & (!j) & (a) & (!e) & (!g182)) + ((l) & (i) & (!j) & (a) & (!e) & (g182)));
	assign g20 = (((!k) & (l) & (!i) & (!j) & (!a) & (g182)) + ((k) & (l) & (!i) & (!j) & (!a) & (g182)) + ((k) & (l) & (!i) & (!j) & (a) & (!g182)) + ((k) & (l) & (!i) & (j) & (!a) & (g182)) + ((k) & (l) & (!i) & (j) & (a) & (!g182)) + ((k) & (l) & (i) & (!j) & (!a) & (g182)) + ((k) & (l) & (i) & (!j) & (a) & (!g182)) + ((k) & (l) & (i) & (j) & (!a) & (g182)));
	assign g21 = (((!k) & (!g14) & (!g16) & (!g18) & (!g19) & (!g20)) + ((!k) & (!g14) & (g16) & (!g18) & (!g19) & (!g20)) + ((!k) & (!g14) & (g16) & (g18) & (!g19) & (!g20)) + ((!k) & (g14) & (!g16) & (!g18) & (!g19) & (!g20)) + ((!k) & (g14) & (!g16) & (g18) & (!g19) & (!g20)) + ((!k) & (g14) & (g16) & (!g18) & (!g19) & (!g20)) + ((k) & (!g14) & (!g16) & (!g18) & (!g19) & (!g20)) + ((k) & (!g14) & (!g16) & (!g18) & (g19) & (!g20)) + ((k) & (!g14) & (g16) & (!g18) & (!g19) & (!g20)) + ((k) & (!g14) & (g16) & (!g18) & (g19) & (!g20)) + ((k) & (!g14) & (g16) & (g18) & (!g19) & (!g20)) + ((k) & (!g14) & (g16) & (g18) & (g19) & (!g20)) + ((k) & (g14) & (!g16) & (!g18) & (!g19) & (!g20)) + ((k) & (g14) & (!g16) & (!g18) & (g19) & (!g20)) + ((k) & (g14) & (!g16) & (g18) & (!g19) & (!g20)) + ((k) & (g14) & (!g16) & (g18) & (g19) & (!g20)) + ((k) & (g14) & (g16) & (!g18) & (!g19) & (!g20)) + ((k) & (g14) & (g16) & (!g18) & (g19) & (!g20)));
	assign g22 = (((!l) & (n) & (!j)));
	assign g23 = (((k) & (i) & (g22)));
	assign g24 = (((!g182) & (g16) & (g23)) + ((g182) & (!g16) & (g23)));
	assign g25 = (((k) & (!l) & (n) & (g8) & (!a) & (g14)) + ((k) & (!l) & (n) & (g8) & (a) & (g14)) + ((k) & (l) & (n) & (g8) & (!a) & (!g14)) + ((k) & (l) & (n) & (g8) & (!a) & (g14)));
	assign g26 = (((!i) & (g22)));
	assign g27 = (((!k) & (l) & (n) & (i) & (j)) + ((k) & (!l) & (n) & (!i) & (j)));
	assign g28 = (((i) & (g22)));
	assign g29 = (((!k) & (!e) & (!g182) & (g27) & (!g28)) + ((!k) & (!e) & (!g182) & (g27) & (g28)) + ((!k) & (e) & (!g182) & (!g27) & (g28)) + ((!k) & (e) & (!g182) & (g27) & (!g28)) + ((!k) & (e) & (!g182) & (g27) & (g28)) + ((!k) & (e) & (g182) & (!g27) & (g28)) + ((!k) & (e) & (g182) & (g27) & (g28)) + ((k) & (!e) & (!g182) & (g27) & (!g28)) + ((k) & (!e) & (!g182) & (g27) & (g28)) + ((k) & (e) & (!g182) & (g27) & (!g28)) + ((k) & (e) & (!g182) & (g27) & (g28)));
	assign g30 = (((!k) & (!a) & (!g14) & (!g26) & (!g29)) + ((!k) & (!a) & (!g14) & (g26) & (!g29)) + ((!k) & (!a) & (g14) & (!g26) & (!g29)) + ((!k) & (!a) & (g14) & (g26) & (!g29)) + ((!k) & (a) & (!g14) & (!g26) & (!g29)) + ((!k) & (a) & (!g14) & (g26) & (!g29)) + ((!k) & (a) & (g14) & (!g26) & (!g29)) + ((k) & (!a) & (!g14) & (!g26) & (!g29)) + ((k) & (!a) & (g14) & (!g26) & (!g29)) + ((k) & (!a) & (g14) & (g26) & (!g29)) + ((k) & (a) & (!g14) & (!g26) & (!g29)) + ((k) & (a) & (!g14) & (g26) & (!g29)) + ((k) & (a) & (g14) & (!g26) & (!g29)));
	assign g31 = (((!n) & (!g21) & (!g24) & (!g25) & (!g30)) + ((!n) & (!g21) & (!g24) & (g25) & (!g30)) + ((!n) & (!g21) & (!g24) & (g25) & (g30)) + ((!n) & (!g21) & (g24) & (!g25) & (!g30)) + ((!n) & (!g21) & (g24) & (!g25) & (g30)) + ((!n) & (!g21) & (g24) & (g25) & (!g30)) + ((!n) & (!g21) & (g24) & (g25) & (g30)) + ((!n) & (g21) & (!g24) & (!g25) & (!g30)) + ((!n) & (g21) & (!g24) & (g25) & (!g30)) + ((!n) & (g21) & (!g24) & (g25) & (g30)) + ((!n) & (g21) & (g24) & (!g25) & (!g30)) + ((!n) & (g21) & (g24) & (!g25) & (g30)) + ((!n) & (g21) & (g24) & (g25) & (!g30)) + ((!n) & (g21) & (g24) & (g25) & (g30)) + ((n) & (!g21) & (!g24) & (!g25) & (!g30)) + ((n) & (!g21) & (!g24) & (!g25) & (g30)) + ((n) & (!g21) & (!g24) & (g25) & (!g30)) + ((n) & (!g21) & (!g24) & (g25) & (g30)) + ((n) & (!g21) & (g24) & (!g25) & (!g30)) + ((n) & (!g21) & (g24) & (!g25) & (g30)) + ((n) & (!g21) & (g24) & (g25) & (!g30)) + ((n) & (!g21) & (g24) & (g25) & (g30)) + ((n) & (g21) & (!g24) & (!g25) & (!g30)) + ((n) & (g21) & (!g24) & (g25) & (!g30)) + ((n) & (g21) & (!g24) & (g25) & (g30)) + ((n) & (g21) & (g24) & (!g25) & (!g30)) + ((n) & (g21) & (g24) & (!g25) & (g30)) + ((n) & (g21) & (g24) & (g25) & (!g30)) + ((n) & (g21) & (g24) & (g25) & (g30)));
	assign g32 = (((!k) & (!n) & (!i)));
	assign g33 = (((!k) & (!l) & (n) & (i) & (j)) + ((k) & (l) & (!n) & (!i) & (!j)));
	assign g34 = (((!k) & (l) & (!n) & (!i) & (j)) + ((!k) & (l) & (!n) & (i) & (j)) + ((k) & (!l) & (!n) & (!i) & (j)) + ((k) & (l) & (!n) & (!i) & (j)) + ((k) & (l) & (!n) & (i) & (j)));
	assign g35 = (((!k) & (l) & (!n) & (!i) & (!j)) + ((k) & (l) & (!n) & (!i) & (!j)) + ((k) & (l) & (!n) & (!i) & (j)) + ((k) & (l) & (!n) & (i) & (!j)) + ((k) & (l) & (!n) & (i) & (j)));
	assign g36 = (((!g33) & (!a) & (!e) & (!g34) & (!g35)) + ((!g33) & (!a) & (!e) & (!g34) & (g35)) + ((!g33) & (!a) & (!e) & (g34) & (!g35)) + ((!g33) & (!a) & (!e) & (g34) & (g35)) + ((!g33) & (!a) & (e) & (!g34) & (!g35)) + ((!g33) & (!a) & (e) & (!g34) & (g35)) + ((!g33) & (!a) & (e) & (g34) & (!g35)) + ((!g33) & (!a) & (e) & (g34) & (g35)) + ((!g33) & (a) & (!e) & (!g34) & (!g35)) + ((!g33) & (a) & (!e) & (g34) & (!g35)) + ((!g33) & (a) & (e) & (!g34) & (!g35)));
	assign g37 = (((!e) & (!g32) & (!g182) & (!g36)) + ((!e) & (!g32) & (g182) & (!g36)) + ((!e) & (g32) & (!g182) & (!g36)) + ((!e) & (g32) & (g182) & (!g36)) + ((e) & (!g32) & (!g182) & (!g36)) + ((e) & (!g32) & (g182) & (!g36)) + ((e) & (g32) & (!g182) & (!g36)) + ((e) & (g32) & (g182) & (!g36)) + ((e) & (g32) & (g182) & (g36)));
	assign g38 = (((k) & (l) & (n) & (!i) & (!j)));
	assign g39 = (((!a) & (!e) & (!g1) & (!f) & (b)) + ((!a) & (!e) & (g1) & (!f) & (b)) + ((!a) & (!e) & (g1) & (f) & (!b)) + ((!a) & (e) & (!g1) & (!f) & (!b)) + ((!a) & (e) & (g1) & (!f) & (!b)) + ((a) & (!e) & (!g1) & (!f) & (b)) + ((a) & (!e) & (g1) & (!f) & (b)) + ((a) & (!e) & (g1) & (f) & (!b)) + ((a) & (e) & (!g1) & (!f) & (b)) + ((a) & (e) & (g1) & (!f) & (b)) + ((a) & (e) & (g1) & (f) & (!b)));
	assign g40 = (((!g2) & (g3) & (!f) & (!b)) + ((!g2) & (g3) & (f) & (!b)) + ((g2) & (!g3) & (!f) & (!b)) + ((g2) & (!g3) & (!f) & (b)) + ((g2) & (g3) & (!f) & (!b)) + ((g2) & (g3) & (!f) & (b)) + ((g2) & (g3) & (f) & (!b)));
	assign g41 = (((!k) & (l) & (n) & (!i) & (!j)) + ((!k) & (l) & (n) & (i) & (j)) + ((k) & (!l) & (!n) & (!i) & (!j)) + ((k) & (!l) & (n) & (!i) & (!j)) + ((k) & (!l) & (n) & (i) & (!j)));
	assign g42 = (((n) & (!i) & (!a) & (e) & (g1)));
	assign g43 = (((!g4) & (f) & (b) & (!g41) & (g42)) + ((!g4) & (f) & (b) & (g41) & (!g42)) + ((!g4) & (f) & (b) & (g41) & (g42)) + ((g4) & (!f) & (b) & (!g41) & (!g42)) + ((g4) & (!f) & (b) & (!g41) & (g42)) + ((g4) & (!f) & (b) & (g41) & (!g42)) + ((g4) & (!f) & (b) & (g41) & (g42)) + ((g4) & (f) & (!b) & (!g41) & (!g42)) + ((g4) & (f) & (!b) & (!g41) & (g42)) + ((g4) & (f) & (!b) & (g41) & (!g42)) + ((g4) & (f) & (!b) & (g41) & (g42)) + ((g4) & (f) & (b) & (!g41) & (!g42)) + ((g4) & (f) & (b) & (!g41) & (g42)) + ((g4) & (f) & (b) & (g41) & (!g42)) + ((g4) & (f) & (b) & (g41) & (g42)));
	assign g44 = (((!a) & (!g11) & (!g38) & (!g39) & (!g40) & (g43)) + ((!a) & (!g11) & (!g38) & (!g39) & (g40) & (!g43)) + ((!a) & (!g11) & (!g38) & (!g39) & (g40) & (g43)) + ((!a) & (!g11) & (!g38) & (g39) & (!g40) & (g43)) + ((!a) & (!g11) & (!g38) & (g39) & (g40) & (!g43)) + ((!a) & (!g11) & (!g38) & (g39) & (g40) & (g43)) + ((!a) & (!g11) & (g38) & (!g39) & (!g40) & (g43)) + ((!a) & (!g11) & (g38) & (!g39) & (g40) & (!g43)) + ((!a) & (!g11) & (g38) & (!g39) & (g40) & (g43)) + ((!a) & (!g11) & (g38) & (g39) & (!g40) & (g43)) + ((!a) & (!g11) & (g38) & (g39) & (g40) & (!g43)) + ((!a) & (!g11) & (g38) & (g39) & (g40) & (g43)) + ((!a) & (g11) & (!g38) & (!g39) & (!g40) & (g43)) + ((!a) & (g11) & (!g38) & (!g39) & (g40) & (!g43)) + ((!a) & (g11) & (!g38) & (!g39) & (g40) & (g43)) + ((!a) & (g11) & (!g38) & (g39) & (!g40) & (!g43)) + ((!a) & (g11) & (!g38) & (g39) & (!g40) & (g43)) + ((!a) & (g11) & (!g38) & (g39) & (g40) & (!g43)) + ((!a) & (g11) & (!g38) & (g39) & (g40) & (g43)) + ((!a) & (g11) & (g38) & (!g39) & (!g40) & (g43)) + ((!a) & (g11) & (g38) & (!g39) & (g40) & (!g43)) + ((!a) & (g11) & (g38) & (!g39) & (g40) & (g43)) + ((!a) & (g11) & (g38) & (g39) & (!g40) & (!g43)) + ((!a) & (g11) & (g38) & (g39) & (!g40) & (g43)) + ((!a) & (g11) & (g38) & (g39) & (g40) & (!g43)) + ((!a) & (g11) & (g38) & (g39) & (g40) & (g43)) + ((a) & (!g11) & (!g38) & (!g39) & (!g40) & (g43)) + ((a) & (!g11) & (!g38) & (!g39) & (g40) & (!g43)) + ((a) & (!g11) & (!g38) & (!g39) & (g40) & (g43)) + ((a) & (!g11) & (!g38) & (g39) & (!g40) & (g43)) + ((a) & (!g11) & (!g38) & (g39) & (g40) & (!g43)) + ((a) & (!g11) & (!g38) & (g39) & (g40) & (g43)) + ((a) & (!g11) & (g38) & (!g39) & (!g40) & (!g43)) + ((a) & (!g11) & (g38) & (!g39) & (!g40) & (g43)) + ((a) & (!g11) & (g38) & (!g39) & (g40) & (!g43)) + ((a) & (!g11) & (g38) & (!g39) & (g40) & (g43)) + ((a) & (!g11) & (g38) & (g39) & (!g40) & (!g43)) + ((a) & (!g11) & (g38) & (g39) & (!g40) & (g43)) + ((a) & (!g11) & (g38) & (g39) & (g40) & (!g43)) + ((a) & (!g11) & (g38) & (g39) & (g40) & (g43)) + ((a) & (g11) & (!g38) & (!g39) & (!g40) & (g43)) + ((a) & (g11) & (!g38) & (!g39) & (g40) & (!g43)) + ((a) & (g11) & (!g38) & (!g39) & (g40) & (g43)) + ((a) & (g11) & (!g38) & (g39) & (!g40) & (!g43)) + ((a) & (g11) & (!g38) & (g39) & (!g40) & (g43)) + ((a) & (g11) & (!g38) & (g39) & (g40) & (!g43)) + ((a) & (g11) & (!g38) & (g39) & (g40) & (g43)) + ((a) & (g11) & (g38) & (!g39) & (!g40) & (!g43)) + ((a) & (g11) & (g38) & (!g39) & (!g40) & (g43)) + ((a) & (g11) & (g38) & (!g39) & (g40) & (!g43)) + ((a) & (g11) & (g38) & (!g39) & (g40) & (g43)) + ((a) & (g11) & (g38) & (g39) & (!g40) & (!g43)) + ((a) & (g11) & (g38) & (g39) & (!g40) & (g43)) + ((a) & (g11) & (g38) & (g39) & (g40) & (!g43)) + ((a) & (g11) & (g38) & (g39) & (g40) & (g43)));
	assign g45 = (((g7) & (f)));
	assign g46 = (((!g9) & (!g10) & (!g12) & (!b) & (!g44) & (!g45)) + ((!g9) & (!g10) & (!g12) & (!b) & (!g44) & (g45)) + ((!g9) & (!g10) & (!g12) & (!b) & (g44) & (!g45)) + ((!g9) & (!g10) & (!g12) & (!b) & (g44) & (g45)) + ((!g9) & (!g10) & (!g12) & (b) & (!g44) & (!g45)) + ((!g9) & (!g10) & (!g12) & (b) & (g44) & (!g45)) + ((!g9) & (!g10) & (g12) & (!b) & (!g44) & (!g45)) + ((!g9) & (!g10) & (g12) & (!b) & (!g44) & (g45)) + ((!g9) & (g10) & (!g12) & (!b) & (g44) & (!g45)) + ((!g9) & (g10) & (!g12) & (!b) & (g44) & (g45)) + ((!g9) & (g10) & (!g12) & (b) & (g44) & (!g45)) + ((g9) & (!g10) & (!g12) & (!b) & (!g44) & (!g45)) + ((g9) & (!g10) & (!g12) & (!b) & (!g44) & (g45)) + ((g9) & (!g10) & (!g12) & (!b) & (g44) & (!g45)) + ((g9) & (!g10) & (!g12) & (!b) & (g44) & (g45)) + ((g9) & (!g10) & (!g12) & (b) & (!g44) & (!g45)) + ((g9) & (!g10) & (g12) & (!b) & (!g44) & (!g45)) + ((g9) & (!g10) & (g12) & (!b) & (!g44) & (g45)) + ((g9) & (g10) & (!g12) & (!b) & (g44) & (!g45)) + ((g9) & (g10) & (!g12) & (!b) & (g44) & (g45)));
	assign g47 = (((g15) & (f) & (b)));
	assign g48 = (((!g7) & (!g46) & (!g47)) + ((!g7) & (g46) & (!g47)) + ((g7) & (!g46) & (!g47)));
	assign g49 = (((!k) & (l) & (!i) & (j) & (a) & (e)));
	assign g50 = (((a) & (g182)));
	assign g51 = (((!k) & (l) & (!i) & (!j)) + ((k) & (l) & (!i) & (!j)) + ((k) & (l) & (!i) & (j)) + ((k) & (l) & (i) & (!j)));
	assign g52 = (((g50) & (!b) & (!g44) & (g51)));
	assign g53 = (((!k) & (!l) & (!i) & (!j)) + ((!k) & (l) & (!i) & (!j)) + ((k) & (l) & (!i) & (!j)) + ((k) & (l) & (!i) & (j)) + ((k) & (l) & (i) & (!j)));
	assign g54 = (((!l) & (g17)));
	assign g55 = (((!k) & (!l) & (!i) & (j)) + ((!k) & (l) & (i) & (j)) + ((k) & (!l) & (!i) & (j)));
	assign g56 = (((!g182) & (g54) & (!g55)) + ((!g182) & (g54) & (g55)) + ((g182) & (!g54) & (g55)) + ((g182) & (g54) & (!g55)) + ((g182) & (g54) & (g55)));
	assign g57 = (((!k) & (!l) & (!g8)));
	assign g58 = (((n) & (!g46) & (!g48) & (!g49) & (!g52) & (g206)) + ((n) & (!g46) & (!g48) & (!g49) & (g52) & (!g206)) + ((n) & (!g46) & (!g48) & (!g49) & (g52) & (g206)) + ((n) & (!g46) & (!g48) & (g49) & (!g52) & (g206)) + ((n) & (!g46) & (!g48) & (g49) & (g52) & (!g206)) + ((n) & (!g46) & (!g48) & (g49) & (g52) & (g206)) + ((n) & (!g46) & (g48) & (!g49) & (!g52) & (g206)) + ((n) & (!g46) & (g48) & (!g49) & (g52) & (!g206)) + ((n) & (!g46) & (g48) & (!g49) & (g52) & (g206)) + ((n) & (!g46) & (g48) & (g49) & (!g52) & (g206)) + ((n) & (!g46) & (g48) & (g49) & (g52) & (!g206)) + ((n) & (!g46) & (g48) & (g49) & (g52) & (g206)) + ((n) & (g46) & (!g48) & (!g49) & (!g52) & (g206)) + ((n) & (g46) & (!g48) & (!g49) & (g52) & (!g206)) + ((n) & (g46) & (!g48) & (!g49) & (g52) & (g206)) + ((n) & (g46) & (!g48) & (g49) & (!g52) & (g206)) + ((n) & (g46) & (!g48) & (g49) & (g52) & (!g206)) + ((n) & (g46) & (!g48) & (g49) & (g52) & (g206)) + ((n) & (g46) & (g48) & (!g49) & (!g52) & (g206)) + ((n) & (g46) & (g48) & (!g49) & (g52) & (!g206)) + ((n) & (g46) & (g48) & (!g49) & (g52) & (g206)) + ((n) & (g46) & (g48) & (g49) & (!g52) & (!g206)) + ((n) & (g46) & (g48) & (g49) & (!g52) & (g206)) + ((n) & (g46) & (g48) & (g49) & (g52) & (!g206)) + ((n) & (g46) & (g48) & (g49) & (g52) & (g206)));
	assign g59 = (((!g182) & (!g16) & (g23) & (!g44) & (!g48)) + ((!g182) & (!g16) & (g23) & (g44) & (g48)) + ((!g182) & (g16) & (g23) & (!g44) & (!g48)) + ((!g182) & (g16) & (g23) & (g44) & (g48)) + ((g182) & (!g16) & (g23) & (!g44) & (!g48)) + ((g182) & (!g16) & (g23) & (g44) & (g48)) + ((g182) & (g16) & (g23) & (!g44) & (g48)) + ((g182) & (g16) & (g23) & (g44) & (!g48)));
	assign g60 = (((k) & (n) & (g8)));
	assign g61 = (((!l) & (!a) & (!g14) & (!b) & (!g46)) + ((!l) & (!a) & (!g14) & (b) & (!g46)) + ((!l) & (!a) & (g14) & (!b) & (g46)) + ((!l) & (!a) & (g14) & (b) & (g46)) + ((!l) & (a) & (!g14) & (!b) & (!g46)) + ((!l) & (a) & (!g14) & (b) & (!g46)) + ((!l) & (a) & (g14) & (!b) & (g46)) + ((!l) & (a) & (g14) & (b) & (g46)) + ((l) & (!a) & (!g14) & (!b) & (!g46)) + ((l) & (!a) & (!g14) & (!b) & (g46)) + ((l) & (!a) & (g14) & (!b) & (!g46)) + ((l) & (!a) & (g14) & (!b) & (g46)) + ((l) & (a) & (!g14) & (b) & (!g46)) + ((l) & (a) & (!g14) & (b) & (g46)) + ((l) & (a) & (g14) & (b) & (!g46)) + ((l) & (a) & (g14) & (b) & (g46)));
	assign g62 = (((!g182) & (!g44)));
	assign g63 = (((!k) & (i) & (g22) & (f)));
	assign g64 = (((!l) & (!a) & (!e) & (!f) & (b)) + ((!l) & (!a) & (!e) & (f) & (!b)) + ((!l) & (!a) & (e) & (!f) & (b)) + ((!l) & (!a) & (e) & (f) & (!b)) + ((!l) & (a) & (!e) & (!f) & (b)) + ((!l) & (a) & (!e) & (f) & (!b)) + ((!l) & (a) & (e) & (f) & (b)) + ((l) & (!a) & (!e) & (!f) & (b)) + ((l) & (!a) & (!e) & (f) & (!b)) + ((l) & (!a) & (e) & (!f) & (b)) + ((l) & (!a) & (e) & (f) & (!b)) + ((l) & (a) & (!e) & (!f) & (b)) + ((l) & (a) & (!e) & (f) & (!b)) + ((l) & (a) & (e) & (!f) & (!b)) + ((l) & (a) & (e) & (f) & (b)));
	assign g65 = (((!k) & (n) & (i) & (!j)));
	assign g66 = (((!g27) & (!g62) & (!g63) & (!g64) & (!g65)) + ((!g27) & (!g62) & (!g63) & (!g64) & (g65)) + ((!g27) & (!g62) & (!g63) & (g64) & (!g65)) + ((!g27) & (g62) & (!g63) & (!g64) & (!g65)) + ((!g27) & (g62) & (!g63) & (!g64) & (g65)) + ((!g27) & (g62) & (!g63) & (g64) & (!g65)) + ((g27) & (!g62) & (!g63) & (!g64) & (!g65)) + ((g27) & (!g62) & (!g63) & (!g64) & (g65)) + ((g27) & (!g62) & (!g63) & (g64) & (!g65)));
	assign g67 = (((a) & (e) & (g15)));
	assign g68 = (((!k) & (l) & (g11)));
	assign g69 = (((l) & (!i) & (a) & (e)));
	assign g70 = (((!g7) & (!g67) & (!g46) & (!g47) & (g68) & (!g69)) + ((!g7) & (!g67) & (!g46) & (!g47) & (g68) & (g69)) + ((!g7) & (!g67) & (!g46) & (g47) & (!g68) & (g69)) + ((!g7) & (!g67) & (!g46) & (g47) & (g68) & (g69)) + ((!g7) & (!g67) & (g46) & (g47) & (g68) & (!g69)) + ((!g7) & (!g67) & (g46) & (g47) & (g68) & (g69)) + ((!g7) & (g67) & (!g46) & (g47) & (!g68) & (g69)) + ((!g7) & (g67) & (!g46) & (g47) & (g68) & (g69)) + ((g7) & (!g67) & (!g46) & (!g47) & (g68) & (!g69)) + ((g7) & (!g67) & (!g46) & (!g47) & (g68) & (g69)) + ((g7) & (!g67) & (!g46) & (g47) & (!g68) & (g69)) + ((g7) & (!g67) & (!g46) & (g47) & (g68) & (g69)) + ((g7) & (!g67) & (g46) & (!g47) & (g68) & (!g69)) + ((g7) & (!g67) & (g46) & (!g47) & (g68) & (g69)) + ((g7) & (!g67) & (g46) & (g47) & (g68) & (!g69)) + ((g7) & (!g67) & (g46) & (g47) & (g68) & (g69)) + ((g7) & (g67) & (!g46) & (g47) & (!g68) & (g69)) + ((g7) & (g67) & (!g46) & (g47) & (g68) & (g69)));
	assign g71 = (((!k) & (!a) & (!g14) & (g26) & (b) & (g46)) + ((!k) & (!a) & (g14) & (g26) & (b) & (g46)) + ((!k) & (a) & (!g14) & (g26) & (b) & (!g46)) + ((!k) & (a) & (g14) & (g26) & (b) & (g46)) + ((k) & (!a) & (!g14) & (g26) & (!b) & (!g46)) + ((k) & (!a) & (!g14) & (g26) & (b) & (g46)) + ((k) & (!a) & (g14) & (g26) & (!b) & (!g46)) + ((k) & (!a) & (g14) & (g26) & (b) & (g46)) + ((k) & (a) & (!g14) & (g26) & (!b) & (g46)) + ((k) & (a) & (!g14) & (g26) & (b) & (!g46)) + ((k) & (a) & (g14) & (g26) & (!b) & (!g46)) + ((k) & (a) & (g14) & (g26) & (b) & (g46)));
	assign g72 = (((!g60) & (!g61) & (g66) & (!g70) & (!g71)) + ((!g60) & (g61) & (g66) & (!g70) & (!g71)) + ((g60) & (!g61) & (g66) & (!g70) & (!g71)));
	assign g73 = (((!g58) & (!g59) & (g72)));
	assign g74 = (((!k) & (!l) & (!i) & (!f) & (!b) & (!g44)) + ((!k) & (!l) & (!i) & (!f) & (b) & (!g44)) + ((!k) & (!l) & (!i) & (f) & (!b) & (!g44)) + ((!k) & (!l) & (!i) & (f) & (b) & (!g44)) + ((!k) & (!l) & (i) & (!f) & (!b) & (g44)) + ((!k) & (!l) & (i) & (!f) & (b) & (g44)) + ((!k) & (!l) & (i) & (f) & (!b) & (g44)) + ((!k) & (!l) & (i) & (f) & (b) & (g44)) + ((!k) & (l) & (!i) & (!f) & (!b) & (!g44)) + ((!k) & (l) & (!i) & (f) & (!b) & (!g44)) + ((!k) & (l) & (!i) & (f) & (b) & (!g44)) + ((!k) & (l) & (i) & (!f) & (!b) & (!g44)) + ((!k) & (l) & (i) & (!f) & (!b) & (g44)) + ((!k) & (l) & (i) & (f) & (b) & (!g44)) + ((!k) & (l) & (i) & (f) & (b) & (g44)) + ((k) & (!l) & (!i) & (!f) & (!b) & (g44)) + ((k) & (!l) & (!i) & (!f) & (b) & (g44)) + ((k) & (!l) & (!i) & (f) & (!b) & (g44)) + ((k) & (!l) & (!i) & (f) & (b) & (g44)) + ((k) & (!l) & (i) & (f) & (!b) & (!g44)) + ((k) & (!l) & (i) & (f) & (!b) & (g44)) + ((k) & (!l) & (i) & (f) & (b) & (!g44)) + ((k) & (!l) & (i) & (f) & (b) & (g44)) + ((k) & (l) & (i) & (!f) & (!b) & (!g44)) + ((k) & (l) & (i) & (f) & (!b) & (!g44)) + ((k) & (l) & (i) & (f) & (b) & (!g44)));
	assign g75 = (((!k) & (l) & (!i) & (f) & (!b) & (!g44)) + ((!k) & (l) & (!i) & (f) & (!b) & (g44)) + ((!k) & (l) & (!i) & (f) & (b) & (!g44)) + ((!k) & (l) & (!i) & (f) & (b) & (g44)) + ((k) & (!l) & (!i) & (!f) & (!b) & (!g44)) + ((k) & (!l) & (!i) & (!f) & (!b) & (g44)) + ((k) & (!l) & (i) & (!f) & (b) & (g44)) + ((k) & (!l) & (i) & (f) & (b) & (g44)) + ((k) & (l) & (!i) & (f) & (!b) & (!g44)) + ((k) & (l) & (!i) & (f) & (!b) & (g44)) + ((k) & (l) & (!i) & (f) & (b) & (!g44)) + ((k) & (l) & (!i) & (f) & (b) & (g44)) + ((k) & (l) & (i) & (!f) & (b) & (g44)) + ((k) & (l) & (i) & (f) & (b) & (g44)));
	assign g76 = (((!g34) & (g35) & (!f) & (b)) + ((!g34) & (g35) & (f) & (b)) + ((g34) & (!g35) & (f) & (b)) + ((g34) & (g35) & (!f) & (b)) + ((g34) & (g35) & (f) & (b)));
	assign g77 = (((!g33) & (!g32) & (!f) & (!g44) & (!g76)) + ((!g33) & (!g32) & (!f) & (g44) & (!g76)) + ((!g33) & (!g32) & (f) & (!g44) & (!g76)) + ((!g33) & (!g32) & (f) & (g44) & (!g76)) + ((!g33) & (g32) & (!f) & (!g44) & (!g76)) + ((!g33) & (g32) & (!f) & (g44) & (!g76)) + ((!g33) & (g32) & (f) & (!g44) & (!g76)));
	assign g78 = (((!n) & (!j) & (g74) & (!g75) & (g77)) + ((!n) & (!j) & (g74) & (g75) & (g77)) + ((!n) & (j) & (!g74) & (!g75) & (g77)) + ((!n) & (j) & (g74) & (!g75) & (g77)) + ((n) & (!j) & (!g74) & (!g75) & (g77)) + ((n) & (!j) & (!g74) & (g75) & (g77)) + ((n) & (!j) & (g74) & (!g75) & (g77)) + ((n) & (!j) & (g74) & (g75) & (g77)) + ((n) & (j) & (!g74) & (!g75) & (g77)) + ((n) & (j) & (!g74) & (g75) & (g77)) + ((n) & (j) & (g74) & (!g75) & (g77)) + ((n) & (j) & (g74) & (g75) & (g77)));
	assign p = (((!n) & (!m) & (!g31) & (!g73) & (!g78)) + ((!n) & (!m) & (!g31) & (g73) & (!g78)) + ((!n) & (!m) & (g31) & (!g73) & (!g78)) + ((!n) & (!m) & (g31) & (g73) & (!g78)) + ((!n) & (m) & (!g31) & (!g73) & (!g78)) + ((!n) & (m) & (!g31) & (g73) & (!g78)) + ((!n) & (m) & (g31) & (!g73) & (!g78)) + ((!n) & (m) & (g31) & (g73) & (!g78)) + ((n) & (!m) & (!g31) & (!g73) & (!g78)) + ((n) & (!m) & (!g31) & (!g73) & (g78)) + ((n) & (!m) & (!g31) & (g73) & (!g78)) + ((n) & (!m) & (g31) & (!g73) & (!g78)) + ((n) & (!m) & (g31) & (g73) & (!g78)) + ((n) & (!m) & (g31) & (g73) & (g78)) + ((n) & (m) & (!g31) & (!g73) & (!g78)) + ((n) & (m) & (!g31) & (!g73) & (g78)) + ((n) & (m) & (!g31) & (g73) & (!g78)) + ((n) & (m) & (g31) & (!g73) & (!g78)) + ((n) & (m) & (g31) & (!g73) & (g78)) + ((n) & (m) & (g31) & (g73) & (!g78)));
	assign g80 = (((!m) & (!g31) & (!g58) & (!g59) & (!g72)) + ((!m) & (!g31) & (!g58) & (!g59) & (g72)) + ((!m) & (!g31) & (!g58) & (g59) & (!g72)) + ((!m) & (!g31) & (!g58) & (g59) & (g72)) + ((!m) & (!g31) & (g58) & (!g59) & (!g72)) + ((!m) & (!g31) & (g58) & (!g59) & (g72)) + ((!m) & (!g31) & (g58) & (g59) & (!g72)) + ((!m) & (!g31) & (g58) & (g59) & (g72)) + ((!m) & (g31) & (!g58) & (!g59) & (g72)) + ((m) & (!g31) & (!g58) & (!g59) & (!g72)) + ((m) & (!g31) & (!g58) & (!g59) & (g72)) + ((m) & (!g31) & (!g58) & (g59) & (!g72)) + ((m) & (!g31) & (!g58) & (g59) & (g72)) + ((m) & (!g31) & (g58) & (!g59) & (!g72)) + ((m) & (!g31) & (g58) & (!g59) & (g72)) + ((m) & (!g31) & (g58) & (g59) & (!g72)) + ((m) & (!g31) & (g58) & (g59) & (g72)) + ((m) & (g31) & (!g58) & (!g59) & (!g72)) + ((m) & (g31) & (!g58) & (!g59) & (g72)) + ((m) & (g31) & (!g58) & (g59) & (!g72)) + ((m) & (g31) & (!g58) & (g59) & (g72)) + ((m) & (g31) & (g58) & (!g59) & (!g72)) + ((m) & (g31) & (g58) & (!g59) & (g72)) + ((m) & (g31) & (g58) & (g59) & (!g72)) + ((m) & (g31) & (g58) & (g59) & (g72)));
	assign g81 = (((!a) & (!e) & (f) & (!b)) + ((!a) & (e) & (!f) & (!b)) + ((!a) & (e) & (f) & (!b)) + ((!a) & (e) & (f) & (b)) + ((a) & (!e) & (f) & (!b)) + ((a) & (e) & (f) & (!b)));
	assign g82 = (((!g1) & (g11) & (c) & (!g) & (!g81)) + ((g1) & (g11) & (!c) & (g) & (!g81)) + ((g1) & (g11) & (c) & (!g) & (!g81)));
	assign g83 = (((!j) & (g1) & (c) & (g)) + ((j) & (!g1) & (!c) & (!g)) + ((j) & (g1) & (!c) & (!g)) + ((j) & (g1) & (c) & (g)));
	assign g84 = (((n) & (!i) & (g81) & (g83)));
	assign g85 = (((!g2) & (g3) & (!c) & (!g)) + ((!g2) & (g3) & (!c) & (g)) + ((g2) & (!g3) & (!c) & (!g)) + ((g2) & (!g3) & (c) & (!g)) + ((g2) & (g3) & (!c) & (!g)) + ((g2) & (g3) & (!c) & (g)) + ((g2) & (g3) & (c) & (!g)));
	assign g86 = (((!g4) & (g41) & (c) & (g)) + ((g4) & (!g41) & (!c) & (g)) + ((g4) & (!g41) & (c) & (!g)) + ((g4) & (!g41) & (c) & (g)) + ((g4) & (g41) & (!c) & (g)) + ((g4) & (g41) & (c) & (!g)) + ((g4) & (g41) & (c) & (g)));
	assign g87 = (((!b) & (!g38) & (!g84) & (!g85) & (!g86)) + ((!b) & (g38) & (!g84) & (!g85) & (!g86)) + ((b) & (!g38) & (!g84) & (!g85) & (!g86)));
	assign g88 = (((!g9) & (!g12) & (!c)) + ((!g9) & (!g12) & (c)) + ((g9) & (!g12) & (!c)));
	assign g89 = (((!g7) & (g12) & (c) & (!g)) + ((!g7) & (g12) & (c) & (g)) + ((g7) & (!g12) & (c) & (g)) + ((g7) & (g12) & (c) & (!g)) + ((g7) & (g12) & (c) & (g)));
	assign g90 = (((!g10) & (!g82) & (!g87) & (g88) & (!g89)) + ((!g10) & (!g82) & (g87) & (!g88) & (!g89)) + ((!g10) & (!g82) & (g87) & (g88) & (!g89)) + ((!g10) & (g82) & (!g87) & (g88) & (!g89)) + ((!g10) & (g82) & (g87) & (g88) & (!g89)) + ((g10) & (!g82) & (!g87) & (g88) & (!g89)) + ((g10) & (g82) & (!g87) & (g88) & (!g89)) + ((g10) & (g82) & (g87) & (g88) & (!g89)));
	assign g91 = (((!a) & (!g14) & (!b) & (!g46) & (!g90)) + ((!a) & (!g14) & (!b) & (g46) & (!g90)) + ((!a) & (!g14) & (b) & (!g46) & (g90)) + ((!a) & (!g14) & (b) & (g46) & (!g90)) + ((!a) & (g14) & (!b) & (!g46) & (!g90)) + ((!a) & (g14) & (!b) & (g46) & (!g90)) + ((!a) & (g14) & (b) & (!g46) & (g90)) + ((!a) & (g14) & (b) & (g46) & (!g90)) + ((a) & (!g14) & (!b) & (!g46) & (g90)) + ((a) & (!g14) & (!b) & (g46) & (!g90)) + ((a) & (!g14) & (b) & (!g46) & (g90)) + ((a) & (!g14) & (b) & (g46) & (g90)) + ((a) & (g14) & (!b) & (!g46) & (!g90)) + ((a) & (g14) & (!b) & (g46) & (!g90)) + ((a) & (g14) & (b) & (!g46) & (g90)) + ((a) & (g14) & (b) & (g46) & (!g90)));
	assign g92 = (((!g50) & (b) & (g44)) + ((g50) & (!b) & (g44)) + ((g50) & (b) & (!g44)) + ((g50) & (b) & (g44)));
	assign g93 = (((!g82) & (g87)));
	assign g94 = (((n) & (!g53) & (g57) & (!g92) & (!g93)) + ((n) & (!g53) & (g57) & (!g92) & (g93)) + ((n) & (!g53) & (g57) & (g92) & (!g93)) + ((n) & (!g53) & (g57) & (g92) & (g93)) + ((n) & (g53) & (!g57) & (!g92) & (g93)) + ((n) & (g53) & (g57) & (!g92) & (!g93)) + ((n) & (g53) & (g57) & (!g92) & (g93)) + ((n) & (g53) & (g57) & (g92) & (!g93)) + ((n) & (g53) & (g57) & (g92) & (g93)));
	assign g95 = (((l) & (!a) & (b) & (g60)) + ((l) & (a) & (!b) & (g60)) + ((l) & (a) & (b) & (g60)));
	assign g96 = (((!a) & (!e) & (f) & (b)) + ((!a) & (e) & (f) & (b)) + ((a) & (!e) & (f) & (b)) + ((a) & (e) & (!f) & (b)) + ((a) & (e) & (f) & (!b)) + ((a) & (e) & (f) & (b)));
	assign g97 = (((!g65) & (!g) & (!g95) & (!g96)) + ((!g65) & (!g) & (!g95) & (g96)) + ((!g65) & (g) & (!g95) & (!g96)) + ((!g65) & (g) & (!g95) & (g96)) + ((g65) & (!g) & (!g95) & (g96)) + ((g65) & (g) & (!g95) & (!g96)));
	assign g98 = (((!g26) & (c) & (!g91) & (!g94) & (!g97)) + ((!g26) & (c) & (!g91) & (g94) & (!g97)) + ((!g26) & (c) & (!g91) & (g94) & (g97)) + ((!g26) & (c) & (g91) & (!g94) & (!g97)) + ((!g26) & (c) & (g91) & (g94) & (!g97)) + ((!g26) & (c) & (g91) & (g94) & (g97)) + ((g26) & (c) & (!g91) & (!g94) & (!g97)) + ((g26) & (c) & (!g91) & (!g94) & (g97)) + ((g26) & (c) & (!g91) & (g94) & (!g97)) + ((g26) & (c) & (!g91) & (g94) & (g97)) + ((g26) & (c) & (g91) & (!g94) & (!g97)) + ((g26) & (c) & (g91) & (g94) & (!g97)) + ((g26) & (c) & (g91) & (g94) & (g97)));
	assign g99 = (((!l) & (g65) & (g) & (!g96)) + ((l) & (g65) & (!g) & (g96)) + ((l) & (g65) & (g) & (!g96)));
	assign g100 = (((!n) & (!g51) & (!g92) & (!g93) & (!g99)) + ((!n) & (!g51) & (!g92) & (g93) & (!g99)) + ((!n) & (!g51) & (g92) & (!g93) & (!g99)) + ((!n) & (!g51) & (g92) & (g93) & (!g99)) + ((!n) & (g51) & (!g92) & (!g93) & (!g99)) + ((!n) & (g51) & (!g92) & (g93) & (!g99)) + ((!n) & (g51) & (g92) & (!g93) & (!g99)) + ((!n) & (g51) & (g92) & (g93) & (!g99)) + ((n) & (!g51) & (!g92) & (!g93) & (!g99)) + ((n) & (!g51) & (!g92) & (g93) & (!g99)) + ((n) & (!g51) & (g92) & (!g93) & (!g99)) + ((n) & (!g51) & (g92) & (g93) & (!g99)) + ((n) & (g51) & (!g92) & (!g93) & (!g99)) + ((n) & (g51) & (!g92) & (g93) & (!g99)) + ((n) & (g51) & (g92) & (!g93) & (!g99)));
	assign g101 = (((!k) & (!g26) & (!c) & (!g91) & (!g100)) + ((!k) & (!g26) & (!c) & (g91) & (!g100)) + ((!k) & (g26) & (!c) & (!g91) & (!g100)) + ((!k) & (g26) & (!c) & (g91) & (!g100)) + ((k) & (!g26) & (!c) & (!g91) & (!g100)) + ((k) & (!g26) & (!c) & (g91) & (!g100)) + ((k) & (g26) & (!c) & (!g91) & (!g100)) + ((k) & (g26) & (!c) & (g91) & (!g100)) + ((k) & (g26) & (!c) & (g91) & (g100)));
	assign g102 = (((g15) & (c) & (g)));
	assign g103 = (((!g7) & (!g90) & (!g102)) + ((!g7) & (g90) & (!g102)) + ((g7) & (!g90) & (!g102)));
	assign g104 = (((!g182) & (!g7) & (!g16) & (g44) & (!g46) & (g47)) + ((!g182) & (!g7) & (!g16) & (g44) & (g46) & (g47)) + ((!g182) & (!g7) & (g16) & (g44) & (!g46) & (g47)) + ((!g182) & (!g7) & (g16) & (g44) & (g46) & (g47)) + ((!g182) & (g7) & (!g16) & (g44) & (!g46) & (g47)) + ((!g182) & (g7) & (!g16) & (g44) & (g46) & (!g47)) + ((!g182) & (g7) & (!g16) & (g44) & (g46) & (g47)) + ((!g182) & (g7) & (g16) & (g44) & (!g46) & (g47)) + ((!g182) & (g7) & (g16) & (g44) & (g46) & (!g47)) + ((!g182) & (g7) & (g16) & (g44) & (g46) & (g47)) + ((g182) & (!g7) & (!g16) & (g44) & (!g46) & (g47)) + ((g182) & (!g7) & (!g16) & (g44) & (g46) & (g47)) + ((g182) & (!g7) & (g16) & (!g44) & (!g46) & (g47)) + ((g182) & (!g7) & (g16) & (!g44) & (g46) & (g47)) + ((g182) & (!g7) & (g16) & (g44) & (!g46) & (!g47)) + ((g182) & (!g7) & (g16) & (g44) & (!g46) & (g47)) + ((g182) & (!g7) & (g16) & (g44) & (g46) & (!g47)) + ((g182) & (!g7) & (g16) & (g44) & (g46) & (g47)) + ((g182) & (g7) & (!g16) & (g44) & (!g46) & (g47)) + ((g182) & (g7) & (!g16) & (g44) & (g46) & (!g47)) + ((g182) & (g7) & (!g16) & (g44) & (g46) & (g47)) + ((g182) & (g7) & (g16) & (!g44) & (!g46) & (g47)) + ((g182) & (g7) & (g16) & (!g44) & (g46) & (!g47)) + ((g182) & (g7) & (g16) & (!g44) & (g46) & (g47)) + ((g182) & (g7) & (g16) & (g44) & (!g46) & (!g47)) + ((g182) & (g7) & (g16) & (g44) & (!g46) & (g47)) + ((g182) & (g7) & (g16) & (g44) & (g46) & (!g47)) + ((g182) & (g7) & (g16) & (g44) & (g46) & (g47)));
	assign g105 = (((!k) & (g28) & (g) & (!g93) & (!g103) & (!g104)) + ((!k) & (g28) & (g) & (!g93) & (!g103) & (g104)) + ((!k) & (g28) & (g) & (!g93) & (g103) & (!g104)) + ((!k) & (g28) & (g) & (!g93) & (g103) & (g104)) + ((!k) & (g28) & (g) & (g93) & (!g103) & (!g104)) + ((!k) & (g28) & (g) & (g93) & (!g103) & (g104)) + ((!k) & (g28) & (g) & (g93) & (g103) & (!g104)) + ((!k) & (g28) & (g) & (g93) & (g103) & (g104)) + ((k) & (g28) & (!g) & (!g93) & (!g103) & (g104)) + ((k) & (g28) & (!g) & (!g93) & (g103) & (!g104)) + ((k) & (g28) & (!g) & (g93) & (!g103) & (!g104)) + ((k) & (g28) & (!g) & (g93) & (g103) & (g104)) + ((k) & (g28) & (g) & (!g93) & (!g103) & (g104)) + ((k) & (g28) & (g) & (!g93) & (g103) & (!g104)) + ((k) & (g28) & (g) & (g93) & (!g103) & (!g104)) + ((k) & (g28) & (g) & (g93) & (g103) & (g104)));
	assign g106 = (((!g7) & (!g67) & (!g46) & (!g47)) + ((!g7) & (!g67) & (g46) & (!g47)) + ((!g7) & (!g67) & (g46) & (g47)) + ((!g7) & (g67) & (g46) & (!g47)) + ((g7) & (!g67) & (!g46) & (!g47)) + ((g7) & (!g67) & (g46) & (!g47)) + ((g7) & (!g67) & (g46) & (g47)));
	assign g107 = (((g68) & (!g90) & (!g103) & (!g106)) + ((g68) & (g90) & (!g103) & (g106)));
	assign g108 = (((l) & (!a) & (!b) & (g60) & (!c)));
	assign g109 = (((g27) & (g62) & (g93)));
	assign g110 = (((!l) & (!g14) & (!g46) & (g60) & (!g90)) + ((!l) & (!g14) & (g46) & (g60) & (!g90)) + ((!l) & (g14) & (!g46) & (g60) & (!g90)) + ((!l) & (g14) & (g46) & (g60) & (g90)));
	assign g111 = (((!g182) & (!g44) & (!g54) & (!g55)) + ((!g182) & (!g44) & (!g54) & (g55)) + ((!g182) & (g44) & (!g54) & (!g55)) + ((g182) & (!g44) & (!g54) & (!g55)) + ((g182) & (g44) & (!g54) & (!g55)));
	assign g112 = (((!g51) & (!g53) & (!c) & (!g92) & (g111)) + ((!g51) & (!g53) & (!c) & (g92) & (g111)) + ((!g51) & (!g53) & (c) & (!g92) & (g111)) + ((!g51) & (!g53) & (c) & (g92) & (g111)) + ((!g51) & (g53) & (!c) & (!g92) & (g111)) + ((!g51) & (g53) & (!c) & (g92) & (g111)) + ((!g51) & (g53) & (c) & (!g92) & (g111)) + ((g51) & (!g53) & (!c) & (g92) & (g111)) + ((g51) & (!g53) & (c) & (!g92) & (g111)) + ((g51) & (!g53) & (c) & (g92) & (g111)) + ((g51) & (g53) & (!c) & (g92) & (g111)) + ((g51) & (g53) & (c) & (!g92) & (g111)));
	assign g113 = (((!n) & (!g93) & (!g108) & (!g109) & (!g110) & (!g112)) + ((!n) & (!g93) & (!g108) & (!g109) & (!g110) & (g112)) + ((!n) & (g93) & (!g108) & (!g109) & (!g110) & (!g112)) + ((!n) & (g93) & (!g108) & (!g109) & (!g110) & (g112)) + ((n) & (!g93) & (!g108) & (!g109) & (!g110) & (g112)) + ((n) & (g93) & (!g108) & (!g109) & (!g110) & (!g112)) + ((n) & (g93) & (!g108) & (!g109) & (!g110) & (g112)));
	assign g114 = (((g68) & (!g90) & (g103) & (g106)) + ((g68) & (g90) & (g103) & (!g106)));
	assign g115 = (((!g98) & (!g101) & (!g105) & (!g107) & (!g113) & (!g114)) + ((!g98) & (!g101) & (!g105) & (!g107) & (!g113) & (g114)) + ((!g98) & (!g101) & (!g105) & (!g107) & (g113) & (g114)) + ((!g98) & (!g101) & (!g105) & (g107) & (!g113) & (!g114)) + ((!g98) & (!g101) & (!g105) & (g107) & (!g113) & (g114)) + ((!g98) & (!g101) & (!g105) & (g107) & (g113) & (!g114)) + ((!g98) & (!g101) & (!g105) & (g107) & (g113) & (g114)) + ((!g98) & (!g101) & (g105) & (!g107) & (!g113) & (!g114)) + ((!g98) & (!g101) & (g105) & (!g107) & (!g113) & (g114)) + ((!g98) & (!g101) & (g105) & (!g107) & (g113) & (!g114)) + ((!g98) & (!g101) & (g105) & (!g107) & (g113) & (g114)) + ((!g98) & (!g101) & (g105) & (g107) & (!g113) & (!g114)) + ((!g98) & (!g101) & (g105) & (g107) & (!g113) & (g114)) + ((!g98) & (!g101) & (g105) & (g107) & (g113) & (!g114)) + ((!g98) & (!g101) & (g105) & (g107) & (g113) & (g114)) + ((!g98) & (g101) & (!g105) & (!g107) & (!g113) & (!g114)) + ((!g98) & (g101) & (!g105) & (!g107) & (!g113) & (g114)) + ((!g98) & (g101) & (!g105) & (!g107) & (g113) & (!g114)) + ((!g98) & (g101) & (!g105) & (!g107) & (g113) & (g114)) + ((!g98) & (g101) & (!g105) & (g107) & (!g113) & (!g114)) + ((!g98) & (g101) & (!g105) & (g107) & (!g113) & (g114)) + ((!g98) & (g101) & (!g105) & (g107) & (g113) & (!g114)) + ((!g98) & (g101) & (!g105) & (g107) & (g113) & (g114)) + ((!g98) & (g101) & (g105) & (!g107) & (!g113) & (!g114)) + ((!g98) & (g101) & (g105) & (!g107) & (!g113) & (g114)) + ((!g98) & (g101) & (g105) & (!g107) & (g113) & (!g114)) + ((!g98) & (g101) & (g105) & (!g107) & (g113) & (g114)) + ((!g98) & (g101) & (g105) & (g107) & (!g113) & (!g114)) + ((!g98) & (g101) & (g105) & (g107) & (!g113) & (g114)) + ((!g98) & (g101) & (g105) & (g107) & (g113) & (!g114)) + ((!g98) & (g101) & (g105) & (g107) & (g113) & (g114)) + ((g98) & (!g101) & (!g105) & (!g107) & (!g113) & (!g114)) + ((g98) & (!g101) & (!g105) & (!g107) & (!g113) & (g114)) + ((g98) & (!g101) & (!g105) & (!g107) & (g113) & (!g114)) + ((g98) & (!g101) & (!g105) & (!g107) & (g113) & (g114)) + ((g98) & (!g101) & (!g105) & (g107) & (!g113) & (!g114)) + ((g98) & (!g101) & (!g105) & (g107) & (!g113) & (g114)) + ((g98) & (!g101) & (!g105) & (g107) & (g113) & (!g114)) + ((g98) & (!g101) & (!g105) & (g107) & (g113) & (g114)) + ((g98) & (!g101) & (g105) & (!g107) & (!g113) & (!g114)) + ((g98) & (!g101) & (g105) & (!g107) & (!g113) & (g114)) + ((g98) & (!g101) & (g105) & (!g107) & (g113) & (!g114)) + ((g98) & (!g101) & (g105) & (!g107) & (g113) & (g114)) + ((g98) & (!g101) & (g105) & (g107) & (!g113) & (!g114)) + ((g98) & (!g101) & (g105) & (g107) & (!g113) & (g114)) + ((g98) & (!g101) & (g105) & (g107) & (g113) & (!g114)) + ((g98) & (!g101) & (g105) & (g107) & (g113) & (g114)) + ((g98) & (g101) & (!g105) & (!g107) & (!g113) & (!g114)) + ((g98) & (g101) & (!g105) & (!g107) & (!g113) & (g114)) + ((g98) & (g101) & (!g105) & (!g107) & (g113) & (!g114)) + ((g98) & (g101) & (!g105) & (!g107) & (g113) & (g114)) + ((g98) & (g101) & (!g105) & (g107) & (!g113) & (!g114)) + ((g98) & (g101) & (!g105) & (g107) & (!g113) & (g114)) + ((g98) & (g101) & (!g105) & (g107) & (g113) & (!g114)) + ((g98) & (g101) & (!g105) & (g107) & (g113) & (g114)) + ((g98) & (g101) & (g105) & (!g107) & (!g113) & (!g114)) + ((g98) & (g101) & (g105) & (!g107) & (!g113) & (g114)) + ((g98) & (g101) & (g105) & (!g107) & (g113) & (!g114)) + ((g98) & (g101) & (g105) & (!g107) & (g113) & (g114)) + ((g98) & (g101) & (g105) & (g107) & (!g113) & (!g114)) + ((g98) & (g101) & (g105) & (g107) & (!g113) & (g114)) + ((g98) & (g101) & (g105) & (g107) & (g113) & (!g114)) + ((g98) & (g101) & (g105) & (g107) & (g113) & (g114)));
	assign g116 = (((!k) & (!l) & (!i) & (!c) & (!g) & (!g93)) + ((!k) & (!l) & (!i) & (!c) & (g) & (!g93)) + ((!k) & (!l) & (!i) & (c) & (!g) & (!g93)) + ((!k) & (!l) & (!i) & (c) & (g) & (!g93)) + ((!k) & (!l) & (i) & (!c) & (!g) & (g93)) + ((!k) & (!l) & (i) & (!c) & (g) & (g93)) + ((!k) & (!l) & (i) & (c) & (!g) & (g93)) + ((!k) & (!l) & (i) & (c) & (g) & (g93)) + ((!k) & (l) & (!i) & (!c) & (!g) & (!g93)) + ((!k) & (l) & (!i) & (!c) & (g) & (!g93)) + ((!k) & (l) & (!i) & (c) & (!g) & (!g93)) + ((!k) & (l) & (!i) & (c) & (!g) & (g93)) + ((!k) & (l) & (!i) & (c) & (g) & (!g93)) + ((!k) & (l) & (i) & (!c) & (g) & (!g93)) + ((!k) & (l) & (i) & (!c) & (g) & (g93)) + ((!k) & (l) & (i) & (c) & (!g) & (!g93)) + ((!k) & (l) & (i) & (c) & (!g) & (g93)) + ((k) & (!l) & (!i) & (!c) & (!g) & (g93)) + ((k) & (!l) & (!i) & (!c) & (g) & (g93)) + ((k) & (!l) & (!i) & (c) & (!g) & (g93)) + ((k) & (!l) & (!i) & (c) & (g) & (g93)) + ((k) & (!l) & (i) & (!c) & (!g) & (!g93)) + ((k) & (!l) & (i) & (!c) & (!g) & (g93)) + ((k) & (!l) & (i) & (c) & (!g) & (!g93)) + ((k) & (!l) & (i) & (c) & (!g) & (g93)) + ((k) & (l) & (!i) & (!c) & (!g) & (!g93)) + ((k) & (l) & (!i) & (!c) & (!g) & (g93)) + ((k) & (l) & (!i) & (!c) & (g) & (!g93)) + ((k) & (l) & (!i) & (!c) & (g) & (g93)) + ((k) & (l) & (!i) & (c) & (!g) & (!g93)) + ((k) & (l) & (!i) & (c) & (!g) & (g93)) + ((k) & (l) & (!i) & (c) & (g) & (!g93)) + ((k) & (l) & (!i) & (c) & (g) & (g93)) + ((k) & (l) & (i) & (!c) & (!g) & (!g93)) + ((k) & (l) & (i) & (!c) & (g) & (!g93)) + ((k) & (l) & (i) & (c) & (!g) & (!g93)) + ((k) & (l) & (i) & (c) & (!g) & (g93)) + ((k) & (l) & (i) & (c) & (g) & (!g93)));
	assign g117 = (((!k) & (l) & (!i) & (!c) & (g) & (!g93)) + ((!k) & (l) & (!i) & (!c) & (g) & (g93)) + ((!k) & (l) & (!i) & (c) & (g) & (!g93)) + ((!k) & (l) & (!i) & (c) & (g) & (g93)) + ((k) & (!l) & (!i) & (!c) & (!g) & (!g93)) + ((k) & (!l) & (!i) & (!c) & (!g) & (g93)) + ((k) & (!l) & (i) & (c) & (!g) & (!g93)) + ((k) & (!l) & (i) & (c) & (g) & (!g93)) + ((k) & (l) & (!i) & (!c) & (g) & (!g93)) + ((k) & (l) & (!i) & (!c) & (g) & (g93)) + ((k) & (l) & (!i) & (c) & (g) & (!g93)) + ((k) & (l) & (!i) & (c) & (g) & (g93)) + ((k) & (l) & (i) & (c) & (!g) & (!g93)) + ((k) & (l) & (i) & (c) & (g) & (!g93)));
	assign g118 = (((!g34) & (g32) & (!c) & (!g93)) + ((!g34) & (g32) & (c) & (!g93)) + ((g34) & (!g32) & (c) & (!g93)) + ((g34) & (!g32) & (c) & (g93)) + ((g34) & (g32) & (!c) & (!g93)) + ((g34) & (g32) & (c) & (!g93)) + ((g34) & (g32) & (c) & (g93)));
	assign g119 = (((!g33) & (!g35) & (!c) & (g) & (g118)) + ((!g33) & (!g35) & (c) & (g) & (g118)) + ((!g33) & (g35) & (!c) & (g) & (g118)) + ((!g33) & (g35) & (c) & (!g) & (!g118)) + ((!g33) & (g35) & (c) & (!g) & (g118)) + ((!g33) & (g35) & (c) & (g) & (!g118)) + ((!g33) & (g35) & (c) & (g) & (g118)) + ((g33) & (!g35) & (!c) & (!g) & (!g118)) + ((g33) & (!g35) & (!c) & (!g) & (g118)) + ((g33) & (!g35) & (!c) & (g) & (!g118)) + ((g33) & (!g35) & (!c) & (g) & (g118)) + ((g33) & (!g35) & (c) & (!g) & (!g118)) + ((g33) & (!g35) & (c) & (!g) & (g118)) + ((g33) & (!g35) & (c) & (g) & (!g118)) + ((g33) & (!g35) & (c) & (g) & (g118)) + ((g33) & (g35) & (!c) & (!g) & (!g118)) + ((g33) & (g35) & (!c) & (!g) & (g118)) + ((g33) & (g35) & (!c) & (g) & (!g118)) + ((g33) & (g35) & (!c) & (g) & (g118)) + ((g33) & (g35) & (c) & (!g) & (!g118)) + ((g33) & (g35) & (c) & (!g) & (g118)) + ((g33) & (g35) & (c) & (g) & (!g118)) + ((g33) & (g35) & (c) & (g) & (g118)));
	assign g120 = (((g14) & (g46) & (g90)));
	assign g121 = (((d) & (h)));
	assign g122 = (((!c) & (!g) & (g81)) + ((!c) & (g) & (!g81)) + ((!c) & (g) & (g81)) + ((c) & (g) & (g81)));
	assign g123 = (((!k) & (l) & (!i) & (!j) & (!g122)) + ((!k) & (l) & (!i) & (!j) & (g122)) + ((!k) & (l) & (i) & (j) & (!g122)) + ((!k) & (l) & (i) & (j) & (g122)) + ((k) & (!l) & (!i) & (!j) & (!g122)) + ((k) & (!l) & (!i) & (!j) & (g122)) + ((k) & (!l) & (!i) & (j) & (g122)) + ((k) & (!l) & (i) & (!j) & (!g122)) + ((k) & (!l) & (i) & (!j) & (g122)));
	assign g124 = (((n) & (g121) & (g123)));
	assign g125 = (((n) & (j) & (!h)));
	assign g126 = (((!k) & (!l) & (!n) & (!j)) + ((!k) & (!l) & (!n) & (j)) + ((!k) & (l) & (!n) & (!j)));
	assign g127 = (((!i) & (!d) & (!g122) & (!g125) & (g126)) + ((!i) & (!d) & (!g122) & (g125) & (g126)) + ((!i) & (!d) & (g122) & (!g125) & (g126)) + ((!i) & (!d) & (g122) & (g125) & (!g126)) + ((!i) & (!d) & (g122) & (g125) & (g126)));
	assign g128 = (((!g1) & (d) & (!h)) + ((g1) & (!d) & (h)) + ((g1) & (d) & (!h)));
	assign g129 = (((k) & (!l) & (!n) & (!c) & (g121)) + ((k) & (!l) & (!n) & (c) & (g121)) + ((k) & (!l) & (n) & (!c) & (g121)) + ((k) & (!l) & (n) & (c) & (g121)) + ((k) & (l) & (n) & (c) & (!g121)) + ((k) & (l) & (n) & (c) & (g121)));
	assign g130 = (((!g2) & (!g4) & (!d) & (!h)) + ((!g2) & (!g4) & (!d) & (h)) + ((!g2) & (!g4) & (d) & (!h)) + ((!g2) & (!g4) & (d) & (h)) + ((!g2) & (g4) & (!d) & (!h)) + ((g2) & (!g4) & (!d) & (h)) + ((g2) & (!g4) & (d) & (h)));
	assign g131 = (((!i) & (!j) & (!g129) & (g130)) + ((!i) & (j) & (!g129) & (g130)) + ((!i) & (j) & (g129) & (g130)) + ((i) & (!j) & (!g129) & (g130)) + ((i) & (!j) & (g129) & (g130)) + ((i) & (j) & (!g129) & (g130)) + ((i) & (j) & (g129) & (g130)));
	assign g132 = (((!g11) & (!g122) & (!g127) & (!g128) & (g131)) + ((!g11) & (!g122) & (!g127) & (g128) & (g131)) + ((!g11) & (g122) & (!g127) & (!g128) & (g131)) + ((!g11) & (g122) & (!g127) & (g128) & (g131)) + ((g11) & (!g122) & (!g127) & (!g128) & (g131)) + ((g11) & (g122) & (!g127) & (!g128) & (g131)) + ((g11) & (g122) & (!g127) & (g128) & (g131)));
	assign g133 = (((!g9) & (!g12) & (!d)) + ((!g9) & (!g12) & (d)) + ((g9) & (!g12) & (!d)));
	assign g134 = (((!g7) & (g12) & (d) & (!h)) + ((!g7) & (g12) & (d) & (h)) + ((g7) & (!g12) & (d) & (h)) + ((g7) & (g12) & (d) & (!h)) + ((g7) & (g12) & (d) & (h)));
	assign g135 = (((!g10) & (!g124) & (!g132) & (g133) & (!g134)) + ((!g10) & (!g124) & (g132) & (!g133) & (!g134)) + ((!g10) & (!g124) & (g132) & (g133) & (!g134)) + ((!g10) & (g124) & (!g132) & (g133) & (!g134)) + ((!g10) & (g124) & (g132) & (g133) & (!g134)) + ((g10) & (!g124) & (!g132) & (g133) & (!g134)) + ((g10) & (g124) & (!g132) & (g133) & (!g134)) + ((g10) & (g124) & (g132) & (g133) & (!g134)));
	assign g136 = (((!a) & (!b) & (!c) & (!d)) + ((!a) & (!b) & (c) & (d)) + ((!a) & (b) & (!c) & (d)) + ((!a) & (b) & (c) & (d)) + ((a) & (!b) & (!c) & (d)) + ((a) & (!b) & (c) & (d)) + ((a) & (b) & (!c) & (d)) + ((a) & (b) & (c) & (d)));
	assign g137 = (((!l) & (g60) & (!g120) & (!g135) & (!g136)) + ((!l) & (g60) & (!g120) & (!g135) & (g136)) + ((!l) & (g60) & (g120) & (g135) & (!g136)) + ((!l) & (g60) & (g120) & (g135) & (g136)) + ((l) & (g60) & (!g120) & (!g135) & (g136)) + ((l) & (g60) & (!g120) & (g135) & (g136)) + ((l) & (g60) & (g120) & (!g135) & (g136)) + ((l) & (g60) & (g120) & (g135) & (g136)));
	assign g138 = (((!g7) & (g15) & (g121) & (!g135)) + ((!g7) & (g15) & (g121) & (g135)) + ((g7) & (!g15) & (!g121) & (g135)) + ((g7) & (!g15) & (g121) & (g135)) + ((g7) & (g15) & (!g121) & (g135)) + ((g7) & (g15) & (g121) & (!g135)) + ((g7) & (g15) & (g121) & (g135)));
	assign g139 = (((!g7) & (!g67) & (!g46) & (!g47) & (!g90) & (!g102)) + ((!g7) & (!g67) & (!g46) & (!g47) & (g90) & (!g102)) + ((!g7) & (!g67) & (!g46) & (!g47) & (g90) & (g102)) + ((!g7) & (!g67) & (!g46) & (g47) & (g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (!g47) & (!g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (!g47) & (g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (!g47) & (g90) & (g102)) + ((!g7) & (!g67) & (g46) & (g47) & (!g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (g47) & (g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (g47) & (g90) & (g102)) + ((!g7) & (g67) & (!g46) & (!g47) & (g90) & (!g102)) + ((!g7) & (g67) & (!g46) & (g47) & (g90) & (!g102)) + ((!g7) & (g67) & (g46) & (!g47) & (!g90) & (!g102)) + ((!g7) & (g67) & (g46) & (!g47) & (g90) & (!g102)) + ((!g7) & (g67) & (g46) & (!g47) & (g90) & (g102)) + ((!g7) & (g67) & (g46) & (g47) & (g90) & (!g102)) + ((g7) & (!g67) & (!g46) & (!g47) & (!g90) & (!g102)) + ((g7) & (!g67) & (!g46) & (!g47) & (g90) & (!g102)) + ((g7) & (!g67) & (!g46) & (!g47) & (g90) & (g102)) + ((g7) & (!g67) & (g46) & (!g47) & (!g90) & (!g102)) + ((g7) & (!g67) & (g46) & (!g47) & (g90) & (!g102)) + ((g7) & (!g67) & (g46) & (!g47) & (g90) & (g102)) + ((g7) & (!g67) & (g46) & (g47) & (!g90) & (!g102)) + ((g7) & (!g67) & (g46) & (g47) & (g90) & (!g102)) + ((g7) & (!g67) & (g46) & (g47) & (g90) & (g102)));
	assign g140 = (((n) & (g18) & (!g135) & (!g138) & (g139)) + ((n) & (g18) & (!g135) & (g138) & (!g139)) + ((n) & (g18) & (g135) & (!g138) & (!g139)) + ((n) & (g18) & (g135) & (g138) & (g139)));
	assign g141 = (((!g124) & (g132)));
	assign g142 = (((g7) & (!g93) & (g103) & (!g104) & (!g141) & (!g138)) + ((g7) & (!g93) & (g103) & (!g104) & (g141) & (g138)) + ((g7) & (g93) & (!g103) & (!g104) & (!g141) & (!g138)) + ((g7) & (g93) & (!g103) & (!g104) & (g141) & (g138)) + ((g7) & (g93) & (g103) & (!g104) & (!g141) & (!g138)) + ((g7) & (g93) & (g103) & (!g104) & (g141) & (g138)) + ((g7) & (g93) & (g103) & (g104) & (!g141) & (!g138)) + ((g7) & (g93) & (g103) & (g104) & (g141) & (g138)));
	assign g143 = (((g7) & (!g93) & (!g103) & (!g104) & (!g141) & (g138)) + ((g7) & (!g93) & (!g103) & (!g104) & (g141) & (!g138)) + ((g7) & (!g93) & (!g103) & (g104) & (!g141) & (g138)) + ((g7) & (!g93) & (!g103) & (g104) & (g141) & (!g138)) + ((g7) & (!g93) & (g103) & (g104) & (!g141) & (g138)) + ((g7) & (!g93) & (g103) & (g104) & (g141) & (!g138)) + ((g7) & (g93) & (!g103) & (g104) & (!g141) & (g138)) + ((g7) & (g93) & (!g103) & (g104) & (g141) & (!g138)));
	assign g144 = (((!g53) & (!g57) & (!c) & (!g92) & (!g93) & (!g141)) + ((!g53) & (!g57) & (!c) & (!g92) & (!g93) & (g141)) + ((!g53) & (!g57) & (!c) & (!g92) & (g93) & (!g141)) + ((!g53) & (!g57) & (!c) & (!g92) & (g93) & (g141)) + ((!g53) & (!g57) & (!c) & (g92) & (!g93) & (!g141)) + ((!g53) & (!g57) & (!c) & (g92) & (!g93) & (g141)) + ((!g53) & (!g57) & (!c) & (g92) & (g93) & (!g141)) + ((!g53) & (!g57) & (!c) & (g92) & (g93) & (g141)) + ((!g53) & (!g57) & (c) & (!g92) & (!g93) & (!g141)) + ((!g53) & (!g57) & (c) & (!g92) & (!g93) & (g141)) + ((!g53) & (!g57) & (c) & (!g92) & (g93) & (!g141)) + ((!g53) & (!g57) & (c) & (!g92) & (g93) & (g141)) + ((!g53) & (!g57) & (c) & (g92) & (!g93) & (!g141)) + ((!g53) & (!g57) & (c) & (g92) & (!g93) & (g141)) + ((!g53) & (!g57) & (c) & (g92) & (g93) & (!g141)) + ((!g53) & (!g57) & (c) & (g92) & (g93) & (g141)) + ((g53) & (!g57) & (!c) & (!g92) & (!g93) & (!g141)) + ((g53) & (!g57) & (!c) & (!g92) & (g93) & (!g141)) + ((g53) & (!g57) & (!c) & (g92) & (!g93) & (g141)) + ((g53) & (!g57) & (!c) & (g92) & (g93) & (!g141)) + ((g53) & (!g57) & (c) & (!g92) & (!g93) & (g141)) + ((g53) & (!g57) & (c) & (!g92) & (g93) & (!g141)) + ((g53) & (!g57) & (c) & (g92) & (!g93) & (g141)) + ((g53) & (!g57) & (c) & (g92) & (g93) & (g141)));
	assign g145 = (((n) & (d)));
	assign g146 = (((n) & (!g62) & (!g54) & (g55) & (!g93) & (!g141)) + ((n) & (!g62) & (!g54) & (g55) & (g93) & (!g141)) + ((n) & (!g62) & (g54) & (!g55) & (!g93) & (!g141)) + ((n) & (!g62) & (g54) & (!g55) & (g93) & (!g141)) + ((n) & (!g62) & (g54) & (g55) & (!g93) & (!g141)) + ((n) & (!g62) & (g54) & (g55) & (g93) & (!g141)) + ((n) & (g62) & (!g54) & (g55) & (!g93) & (!g141)) + ((n) & (g62) & (g54) & (!g55) & (!g93) & (!g141)) + ((n) & (g62) & (g54) & (!g55) & (g93) & (!g141)) + ((n) & (g62) & (g54) & (g55) & (!g93) & (!g141)) + ((n) & (g62) & (g54) & (g55) & (g93) & (!g141)));
	assign g147 = (((!c) & (g) & (g96)) + ((c) & (!g) & (g96)) + ((c) & (g) & (!g96)) + ((c) & (g) & (g96)));
	assign g148 = (((!l) & (g65) & (!d) & (h) & (!g147)) + ((!l) & (g65) & (!d) & (h) & (g147)) + ((!l) & (g65) & (d) & (!h) & (!g147)) + ((!l) & (g65) & (d) & (h) & (!g147)) + ((!l) & (g65) & (d) & (h) & (g147)) + ((l) & (g65) & (!d) & (!h) & (g147)) + ((l) & (g65) & (!d) & (h) & (!g147)) + ((l) & (g65) & (d) & (!h) & (!g147)) + ((l) & (g65) & (d) & (h) & (g147)));
	assign g149 = (((n) & (g51) & (!d)));
	assign g150 = (((!c) & (!g92) & (!g93) & (!g141) & (!g148) & (!g149)) + ((!c) & (!g92) & (!g93) & (g141) & (!g148) & (!g149)) + ((!c) & (!g92) & (!g93) & (g141) & (!g148) & (g149)) + ((!c) & (!g92) & (g93) & (!g141) & (!g148) & (!g149)) + ((!c) & (!g92) & (g93) & (g141) & (!g148) & (!g149)) + ((!c) & (!g92) & (g93) & (g141) & (!g148) & (g149)) + ((!c) & (g92) & (!g93) & (!g141) & (!g148) & (!g149)) + ((!c) & (g92) & (!g93) & (!g141) & (!g148) & (g149)) + ((!c) & (g92) & (!g93) & (g141) & (!g148) & (!g149)) + ((!c) & (g92) & (g93) & (!g141) & (!g148) & (!g149)) + ((!c) & (g92) & (g93) & (g141) & (!g148) & (!g149)) + ((!c) & (g92) & (g93) & (g141) & (!g148) & (g149)) + ((c) & (!g92) & (!g93) & (!g141) & (!g148) & (!g149)) + ((c) & (!g92) & (!g93) & (!g141) & (!g148) & (g149)) + ((c) & (!g92) & (!g93) & (g141) & (!g148) & (!g149)) + ((c) & (!g92) & (g93) & (!g141) & (!g148) & (!g149)) + ((c) & (!g92) & (g93) & (g141) & (!g148) & (!g149)) + ((c) & (!g92) & (g93) & (g141) & (!g148) & (g149)) + ((c) & (g92) & (!g93) & (!g141) & (!g148) & (!g149)) + ((c) & (g92) & (!g93) & (!g141) & (!g148) & (g149)) + ((c) & (g92) & (!g93) & (g141) & (!g148) & (!g149)) + ((c) & (g92) & (g93) & (!g141) & (!g148) & (!g149)) + ((c) & (g92) & (g93) & (!g141) & (!g148) & (g149)) + ((c) & (g92) & (g93) & (g141) & (!g148) & (!g149)));
	assign g151 = (((!g109) & (!g141) & (!g144) & (!g145) & (!g146) & (g150)) + ((!g109) & (!g141) & (g144) & (!g145) & (!g146) & (g150)) + ((!g109) & (!g141) & (g144) & (g145) & (!g146) & (g150)) + ((!g109) & (g141) & (!g144) & (!g145) & (!g146) & (g150)) + ((!g109) & (g141) & (g144) & (!g145) & (!g146) & (g150)) + ((!g109) & (g141) & (g144) & (g145) & (!g146) & (g150)) + ((g109) & (!g141) & (!g144) & (!g145) & (!g146) & (g150)) + ((g109) & (!g141) & (g144) & (!g145) & (!g146) & (g150)) + ((g109) & (!g141) & (g144) & (g145) & (!g146) & (g150)));
	assign g152 = (((!a) & (!g14) & (!b) & (!g46) & (c) & (!g90)) + ((!a) & (!g14) & (!b) & (g46) & (c) & (!g90)) + ((!a) & (!g14) & (b) & (!g46) & (!c) & (!g90)) + ((!a) & (!g14) & (b) & (!g46) & (c) & (!g90)) + ((!a) & (!g14) & (b) & (!g46) & (c) & (g90)) + ((!a) & (!g14) & (b) & (g46) & (c) & (!g90)) + ((!a) & (g14) & (!b) & (!g46) & (c) & (!g90)) + ((!a) & (g14) & (!b) & (g46) & (c) & (!g90)) + ((!a) & (g14) & (b) & (!g46) & (!c) & (!g90)) + ((!a) & (g14) & (b) & (!g46) & (c) & (!g90)) + ((!a) & (g14) & (b) & (!g46) & (c) & (g90)) + ((!a) & (g14) & (b) & (g46) & (c) & (!g90)) + ((a) & (!g14) & (!b) & (!g46) & (!c) & (!g90)) + ((a) & (!g14) & (!b) & (!g46) & (c) & (!g90)) + ((a) & (!g14) & (!b) & (!g46) & (c) & (g90)) + ((a) & (!g14) & (!b) & (g46) & (c) & (!g90)) + ((a) & (!g14) & (b) & (!g46) & (!c) & (!g90)) + ((a) & (!g14) & (b) & (!g46) & (c) & (!g90)) + ((a) & (!g14) & (b) & (!g46) & (c) & (g90)) + ((a) & (!g14) & (b) & (g46) & (!c) & (!g90)) + ((a) & (!g14) & (b) & (g46) & (c) & (!g90)) + ((a) & (!g14) & (b) & (g46) & (c) & (g90)) + ((a) & (g14) & (!b) & (!g46) & (c) & (!g90)) + ((a) & (g14) & (!b) & (g46) & (c) & (!g90)) + ((a) & (g14) & (b) & (!g46) & (!c) & (!g90)) + ((a) & (g14) & (b) & (!g46) & (c) & (!g90)) + ((a) & (g14) & (b) & (!g46) & (c) & (g90)) + ((a) & (g14) & (b) & (g46) & (c) & (!g90)));
	assign g153 = (((!l) & (!i) & (!j) & (d)));
	assign g154 = (((!i) & (!j) & (g1) & (!d)));
	assign g155 = (((n) & (!g135) & (!g152) & (!g153) & (g154)) + ((n) & (!g135) & (!g152) & (g153) & (g154)) + ((n) & (!g135) & (g152) & (g153) & (!g154)) + ((n) & (!g135) & (g152) & (g153) & (g154)) + ((n) & (g135) & (!g152) & (g153) & (!g154)) + ((n) & (g135) & (!g152) & (g153) & (g154)) + ((n) & (g135) & (g152) & (!g153) & (g154)) + ((n) & (g135) & (g152) & (g153) & (g154)));
	assign g156 = (((!g137) & (!g140) & (!g142) & (!g143) & (g151) & (!g155)));
	assign g157 = (((!k) & (!l) & (!i) & (!d) & (!h) & (g141)) + ((!k) & (!l) & (!i) & (!d) & (h) & (g141)) + ((!k) & (!l) & (!i) & (d) & (!h) & (g141)) + ((!k) & (!l) & (!i) & (d) & (h) & (g141)) + ((!k) & (!l) & (i) & (!d) & (!h) & (!g141)) + ((!k) & (!l) & (i) & (!d) & (h) & (!g141)) + ((!k) & (!l) & (i) & (d) & (!h) & (!g141)) + ((!k) & (!l) & (i) & (d) & (h) & (!g141)) + ((!k) & (l) & (!i) & (!d) & (!h) & (g141)) + ((!k) & (l) & (!i) & (!d) & (h) & (g141)) + ((!k) & (l) & (!i) & (d) & (h) & (g141)) + ((!k) & (l) & (i) & (!d) & (!h) & (!g141)) + ((!k) & (l) & (i) & (!d) & (!h) & (g141)) + ((!k) & (l) & (i) & (d) & (h) & (!g141)) + ((!k) & (l) & (i) & (d) & (h) & (g141)) + ((k) & (!l) & (!i) & (!d) & (!h) & (!g141)) + ((k) & (!l) & (!i) & (!d) & (h) & (!g141)) + ((k) & (!l) & (!i) & (d) & (!h) & (!g141)) + ((k) & (!l) & (!i) & (d) & (h) & (!g141)) + ((k) & (!l) & (i) & (!d) & (h) & (!g141)) + ((k) & (!l) & (i) & (!d) & (h) & (g141)) + ((k) & (!l) & (i) & (d) & (h) & (!g141)) + ((k) & (!l) & (i) & (d) & (h) & (g141)) + ((k) & (l) & (i) & (!d) & (!h) & (g141)) + ((k) & (l) & (i) & (!d) & (h) & (g141)) + ((k) & (l) & (i) & (d) & (h) & (g141)));
	assign g158 = (((!k) & (l) & (!i) & (!d) & (h) & (!g141)) + ((!k) & (l) & (!i) & (!d) & (h) & (g141)) + ((!k) & (l) & (!i) & (d) & (h) & (!g141)) + ((!k) & (l) & (!i) & (d) & (h) & (g141)) + ((k) & (!l) & (!i) & (!d) & (!h) & (!g141)) + ((k) & (!l) & (!i) & (!d) & (!h) & (g141)) + ((k) & (!l) & (i) & (d) & (!h) & (!g141)) + ((k) & (!l) & (i) & (d) & (h) & (!g141)) + ((k) & (l) & (!i) & (!d) & (h) & (!g141)) + ((k) & (l) & (!i) & (!d) & (h) & (g141)) + ((k) & (l) & (!i) & (d) & (h) & (!g141)) + ((k) & (l) & (!i) & (d) & (h) & (g141)) + ((k) & (l) & (i) & (d) & (!h) & (!g141)) + ((k) & (l) & (i) & (d) & (h) & (!g141)));
	assign g159 = (((!g33) & (!g34) & (!g35) & (!d) & (!h)) + ((!g33) & (!g34) & (!g35) & (!d) & (h)) + ((!g33) & (!g34) & (!g35) & (d) & (!h)) + ((!g33) & (!g34) & (!g35) & (d) & (h)) + ((!g33) & (!g34) & (g35) & (!d) & (!h)) + ((!g33) & (!g34) & (g35) & (!d) & (h)) + ((!g33) & (g34) & (!g35) & (!d) & (!h)) + ((!g33) & (g34) & (!g35) & (!d) & (h)) + ((!g33) & (g34) & (!g35) & (d) & (!h)) + ((!g33) & (g34) & (g35) & (!d) & (!h)) + ((!g33) & (g34) & (g35) & (!d) & (h)));
	assign g160 = (((!g32) & (!h) & (!g141) & (g159)) + ((!g32) & (!h) & (g141) & (g159)) + ((!g32) & (h) & (!g141) & (g159)) + ((!g32) & (h) & (g141) & (g159)) + ((g32) & (!h) & (!g141) & (g159)) + ((g32) & (!h) & (g141) & (g159)) + ((g32) & (h) & (g141) & (g159)));
	assign g161 = (((!n) & (!j) & (g157) & (!g158) & (g160)) + ((!n) & (!j) & (g157) & (g158) & (g160)) + ((!n) & (j) & (!g157) & (!g158) & (g160)) + ((!n) & (j) & (g157) & (!g158) & (g160)) + ((n) & (!j) & (!g157) & (!g158) & (g160)) + ((n) & (!j) & (!g157) & (g158) & (g160)) + ((n) & (!j) & (g157) & (!g158) & (g160)) + ((n) & (!j) & (g157) & (g158) & (g160)) + ((n) & (j) & (!g157) & (!g158) & (g160)) + ((n) & (j) & (!g157) & (g158) & (g160)) + ((n) & (j) & (g157) & (!g158) & (g160)) + ((n) & (j) & (g157) & (g158) & (g160)));
	assign r = (((!n) & (!g80) & (!g115) & (!g156) & (!g161)) + ((!n) & (!g80) & (!g115) & (g156) & (!g161)) + ((!n) & (!g80) & (g115) & (!g156) & (!g161)) + ((!n) & (!g80) & (g115) & (g156) & (!g161)) + ((!n) & (g80) & (!g115) & (!g156) & (!g161)) + ((!n) & (g80) & (!g115) & (g156) & (!g161)) + ((!n) & (g80) & (g115) & (!g156) & (!g161)) + ((!n) & (g80) & (g115) & (g156) & (!g161)) + ((n) & (!g80) & (!g115) & (!g156) & (!g161)) + ((n) & (!g80) & (!g115) & (!g156) & (g161)) + ((n) & (!g80) & (!g115) & (g156) & (!g161)) + ((n) & (!g80) & (g115) & (!g156) & (!g161)) + ((n) & (!g80) & (g115) & (g156) & (!g161)) + ((n) & (!g80) & (g115) & (g156) & (g161)) + ((n) & (g80) & (!g115) & (!g156) & (!g161)) + ((n) & (g80) & (!g115) & (!g156) & (g161)) + ((n) & (g80) & (!g115) & (g156) & (!g161)) + ((n) & (g80) & (g115) & (!g156) & (!g161)) + ((n) & (g80) & (g115) & (!g156) & (g161)) + ((n) & (g80) & (g115) & (g156) & (!g161)));
	assign g163 = (((!d) & (h)) + ((d) & (!h)));
	assign g164 = (((!k) & (!l) & (g8) & (!g120) & (!g135)) + ((!k) & (!l) & (g8) & (!g120) & (g135)) + ((!k) & (!l) & (g8) & (g120) & (!g135)) + ((!k) & (!l) & (g8) & (g120) & (g135)) + ((k) & (!l) & (g8) & (g120) & (g135)));
	assign g165 = (((!i) & (d) & (!g135) & (!g152)) + ((!i) & (d) & (!g135) & (g152)) + ((!i) & (d) & (g135) & (g152)));
	assign g166 = (((i) & (!g93) & (!g103) & (!g104) & (!g141) & (!g138)) + ((i) & (!g93) & (!g103) & (!g104) & (!g141) & (g138)) + ((i) & (!g93) & (!g103) & (!g104) & (g141) & (g138)) + ((i) & (!g93) & (!g103) & (g104) & (!g141) & (!g138)) + ((i) & (!g93) & (!g103) & (g104) & (!g141) & (g138)) + ((i) & (!g93) & (!g103) & (g104) & (g141) & (g138)) + ((i) & (!g93) & (g103) & (g104) & (!g141) & (!g138)) + ((i) & (!g93) & (g103) & (g104) & (!g141) & (g138)) + ((i) & (!g93) & (g103) & (g104) & (g141) & (g138)) + ((i) & (g93) & (!g103) & (g104) & (!g141) & (!g138)) + ((i) & (g93) & (!g103) & (g104) & (!g141) & (g138)) + ((i) & (g93) & (!g103) & (g104) & (g141) & (g138)));
	assign g167 = (((!i) & (!g141) & (!g135) & (!g138) & (g152)) + ((!i) & (!g141) & (!g135) & (g138) & (g152)) + ((!i) & (g141) & (!g135) & (!g138) & (g152)) + ((!i) & (g141) & (!g135) & (g138) & (g152)) + ((i) & (!g141) & (!g135) & (g138) & (!g152)) + ((i) & (!g141) & (!g135) & (g138) & (g152)) + ((i) & (!g141) & (g135) & (g138) & (!g152)) + ((i) & (!g141) & (g135) & (g138) & (g152)));
	assign g168 = (((!k) & (!i) & (!j)) + ((k) & (!i) & (!j)) + ((k) & (!i) & (j)) + ((k) & (i) & (!j)));
	assign g169 = (((!c) & (!g92) & (!g93) & (d) & (!g141) & (g168)) + ((!c) & (!g92) & (g93) & (d) & (!g141) & (g168)) + ((!c) & (g92) & (!g93) & (!d) & (!g141) & (g168)) + ((!c) & (g92) & (!g93) & (d) & (!g141) & (g168)) + ((!c) & (g92) & (!g93) & (d) & (g141) & (g168)) + ((!c) & (g92) & (g93) & (d) & (!g141) & (g168)) + ((c) & (!g92) & (!g93) & (!d) & (!g141) & (g168)) + ((c) & (!g92) & (!g93) & (d) & (!g141) & (g168)) + ((c) & (!g92) & (!g93) & (d) & (g141) & (g168)) + ((c) & (!g92) & (g93) & (d) & (!g141) & (g168)) + ((c) & (g92) & (!g93) & (!d) & (!g141) & (g168)) + ((c) & (g92) & (!g93) & (d) & (!g141) & (g168)) + ((c) & (g92) & (!g93) & (d) & (g141) & (g168)) + ((c) & (g92) & (g93) & (!d) & (!g141) & (g168)) + ((c) & (g92) & (g93) & (d) & (!g141) & (g168)) + ((c) & (g92) & (g93) & (d) & (g141) & (g168)));
	assign g170 = (((!g7) & (!g15) & (g17) & (!g121) & (!g135)) + ((!g7) & (!g15) & (g17) & (g121) & (!g135)) + ((!g7) & (g15) & (g17) & (!g121) & (!g135)) + ((!g7) & (g15) & (g17) & (g121) & (!g135)) + ((!g7) & (g15) & (g17) & (g121) & (g135)) + ((g7) & (!g15) & (g17) & (!g121) & (!g135)) + ((g7) & (!g15) & (g17) & (!g121) & (g135)) + ((g7) & (!g15) & (g17) & (g121) & (!g135)) + ((g7) & (!g15) & (g17) & (g121) & (g135)) + ((g7) & (g15) & (g17) & (!g121) & (!g135)) + ((g7) & (g15) & (g17) & (!g121) & (g135)) + ((g7) & (g15) & (g17) & (g121) & (!g135)) + ((g7) & (g15) & (g17) & (g121) & (g135)));
	assign g171 = (((!a) & (!b) & (!c) & (!d)));
	assign g172 = (((!k) & (!g8) & (!g171) & (g183)) + ((!k) & (!g8) & (g171) & (g183)) + ((!k) & (g8) & (!g171) & (g183)) + ((!k) & (g8) & (g171) & (g183)) + ((k) & (g8) & (g171) & (!g183)) + ((k) & (g8) & (g171) & (g183)));
	assign g173 = (((!k) & (!l) & (i) & (j)) + ((!k) & (l) & (i) & (j)) + ((k) & (!l) & (!i) & (j)));
	assign g174 = (((g62) & (g93) & (g141) & (g173)));
	assign g175 = (((!l) & (!g139) & (!g169) & (!g170) & (!g172) & (!g174)) + ((!l) & (!g139) & (!g169) & (!g170) & (g172) & (!g174)) + ((!l) & (!g139) & (!g169) & (g170) & (!g172) & (!g174)) + ((!l) & (!g139) & (!g169) & (g170) & (g172) & (!g174)) + ((!l) & (!g139) & (g169) & (!g170) & (!g172) & (!g174)) + ((!l) & (!g139) & (g169) & (!g170) & (g172) & (!g174)) + ((!l) & (!g139) & (g169) & (g170) & (!g172) & (!g174)) + ((!l) & (!g139) & (g169) & (g170) & (g172) & (!g174)) + ((!l) & (g139) & (!g169) & (!g170) & (!g172) & (!g174)) + ((!l) & (g139) & (!g169) & (!g170) & (g172) & (!g174)) + ((!l) & (g139) & (!g169) & (g170) & (!g172) & (!g174)) + ((!l) & (g139) & (!g169) & (g170) & (g172) & (!g174)) + ((!l) & (g139) & (g169) & (!g170) & (!g172) & (!g174)) + ((!l) & (g139) & (g169) & (!g170) & (g172) & (!g174)) + ((!l) & (g139) & (g169) & (g170) & (!g172) & (!g174)) + ((!l) & (g139) & (g169) & (g170) & (g172) & (!g174)) + ((l) & (!g139) & (!g169) & (!g170) & (!g172) & (!g174)) + ((l) & (g139) & (!g169) & (!g170) & (!g172) & (!g174)) + ((l) & (g139) & (!g169) & (g170) & (!g172) & (!g174)));
	assign g176 = (((!j) & (!g1) & (!g165) & (!g166) & (!g167) & (g175)) + ((!j) & (!g1) & (!g165) & (!g166) & (g167) & (g175)) + ((!j) & (!g1) & (!g165) & (g166) & (!g167) & (g175)) + ((!j) & (!g1) & (!g165) & (g166) & (g167) & (g175)) + ((!j) & (!g1) & (g165) & (!g166) & (!g167) & (g175)) + ((!j) & (!g1) & (g165) & (!g166) & (g167) & (g175)) + ((!j) & (!g1) & (g165) & (g166) & (!g167) & (g175)) + ((!j) & (!g1) & (g165) & (g166) & (g167) & (g175)) + ((!j) & (g1) & (!g165) & (!g166) & (!g167) & (g175)) + ((j) & (!g1) & (!g165) & (!g166) & (!g167) & (g175)) + ((j) & (!g1) & (!g165) & (!g166) & (g167) & (g175)) + ((j) & (!g1) & (!g165) & (g166) & (!g167) & (g175)) + ((j) & (!g1) & (!g165) & (g166) & (g167) & (g175)) + ((j) & (!g1) & (g165) & (!g166) & (!g167) & (g175)) + ((j) & (!g1) & (g165) & (!g166) & (g167) & (g175)) + ((j) & (!g1) & (g165) & (g166) & (!g167) & (g175)) + ((j) & (!g1) & (g165) & (g166) & (g167) & (g175)) + ((j) & (g1) & (!g165) & (!g166) & (!g167) & (g175)) + ((j) & (g1) & (!g165) & (!g166) & (g167) & (g175)) + ((j) & (g1) & (!g165) & (g166) & (!g167) & (g175)) + ((j) & (g1) & (!g165) & (g166) & (g167) & (g175)) + ((j) & (g1) & (g165) & (!g166) & (!g167) & (g175)) + ((j) & (g1) & (g165) & (!g166) & (g167) & (g175)) + ((j) & (g1) & (g165) & (g166) & (!g167) & (g175)) + ((j) & (g1) & (g165) & (g166) & (g167) & (g175)));
	assign u = (((n) & (!g80) & (!g115) & (!g156) & (!g164) & (!g176)) + ((n) & (!g80) & (!g115) & (!g156) & (g164) & (!g176)) + ((n) & (!g80) & (!g115) & (!g156) & (g164) & (g176)) + ((n) & (!g80) & (!g115) & (g156) & (!g164) & (!g176)) + ((n) & (!g80) & (!g115) & (g156) & (g164) & (!g176)) + ((n) & (!g80) & (!g115) & (g156) & (g164) & (g176)) + ((n) & (!g80) & (g115) & (!g156) & (!g164) & (!g176)) + ((n) & (!g80) & (g115) & (!g156) & (!g164) & (g176)) + ((n) & (!g80) & (g115) & (!g156) & (g164) & (!g176)) + ((n) & (!g80) & (g115) & (!g156) & (g164) & (g176)) + ((n) & (!g80) & (g115) & (g156) & (!g164) & (!g176)) + ((n) & (!g80) & (g115) & (g156) & (g164) & (!g176)) + ((n) & (!g80) & (g115) & (g156) & (g164) & (g176)) + ((n) & (g80) & (!g115) & (!g156) & (!g164) & (!g176)) + ((n) & (g80) & (!g115) & (!g156) & (g164) & (!g176)) + ((n) & (g80) & (!g115) & (!g156) & (g164) & (g176)) + ((n) & (g80) & (!g115) & (g156) & (!g164) & (!g176)) + ((n) & (g80) & (!g115) & (g156) & (g164) & (!g176)) + ((n) & (g80) & (!g115) & (g156) & (g164) & (g176)) + ((n) & (g80) & (g115) & (!g156) & (!g164) & (!g176)) + ((n) & (g80) & (g115) & (!g156) & (g164) & (!g176)) + ((n) & (g80) & (g115) & (!g156) & (g164) & (g176)) + ((n) & (g80) & (g115) & (g156) & (!g164) & (!g176)) + ((n) & (g80) & (g115) & (g156) & (g164) & (!g176)) + ((n) & (g80) & (g115) & (g156) & (g164) & (g176)));
	assign g178 = (((!a) & (!e) & (!g163)) + ((a) & (e) & (!g163)));
	assign g179 = (((!f) & (!b) & (!c) & (!g) & (!g178)) + ((!f) & (!b) & (!c) & (g) & (!g178)) + ((!f) & (!b) & (!c) & (g) & (g178)) + ((!f) & (!b) & (c) & (!g) & (!g178)) + ((!f) & (!b) & (c) & (!g) & (g178)) + ((!f) & (!b) & (c) & (g) & (!g178)) + ((!f) & (b) & (!c) & (!g) & (!g178)) + ((!f) & (b) & (!c) & (!g) & (g178)) + ((!f) & (b) & (!c) & (g) & (!g178)) + ((!f) & (b) & (!c) & (g) & (g178)) + ((!f) & (b) & (c) & (!g) & (!g178)) + ((!f) & (b) & (c) & (!g) & (g178)) + ((!f) & (b) & (c) & (g) & (!g178)) + ((!f) & (b) & (c) & (g) & (g178)) + ((f) & (!b) & (!c) & (!g) & (!g178)) + ((f) & (!b) & (!c) & (!g) & (g178)) + ((f) & (!b) & (!c) & (g) & (!g178)) + ((f) & (!b) & (!c) & (g) & (g178)) + ((f) & (!b) & (c) & (!g) & (!g178)) + ((f) & (!b) & (c) & (!g) & (g178)) + ((f) & (!b) & (c) & (g) & (!g178)) + ((f) & (!b) & (c) & (g) & (g178)) + ((f) & (b) & (!c) & (!g) & (!g178)) + ((f) & (b) & (!c) & (g) & (!g178)) + ((f) & (b) & (!c) & (g) & (g178)) + ((f) & (b) & (c) & (!g) & (!g178)) + ((f) & (b) & (c) & (!g) & (g178)) + ((f) & (b) & (c) & (g) & (!g178)));
	assign g180 = (((!l) & (!k) & (!e) & (!a) & (!j) & (!n)) + ((!l) & (!k) & (!e) & (!a) & (j) & (!n)) + ((!l) & (!k) & (!e) & (!a) & (j) & (n)) + ((!l) & (!k) & (!e) & (a) & (j) & (n)) + ((!l) & (!k) & (e) & (!a) & (!j) & (!n)) + ((!l) & (!k) & (e) & (!a) & (j) & (!n)) + ((!l) & (k) & (!e) & (a) & (j) & (n)) + ((!l) & (k) & (e) & (!a) & (j) & (n)) + ((!l) & (k) & (e) & (a) & (!j) & (!n)) + ((!l) & (k) & (e) & (a) & (!j) & (n)) + ((l) & (!k) & (!e) & (!a) & (!j) & (!n)) + ((l) & (!k) & (!e) & (!a) & (j) & (n)) + ((l) & (!k) & (!e) & (a) & (j) & (n)) + ((l) & (!k) & (e) & (!a) & (!j) & (!n)) + ((l) & (!k) & (e) & (a) & (!j) & (n)) + ((l) & (k) & (!e) & (!a) & (j) & (n)) + ((l) & (k) & (!e) & (a) & (j) & (n)));
	assign g181 = (((!l) & (!k) & (!e) & (a) & (!j) & (!n)) + ((!l) & (!k) & (e) & (!a) & (!j) & (!n)) + ((!l) & (!k) & (e) & (a) & (!j) & (!n)) + ((!l) & (k) & (!e) & (!a) & (j) & (!n)) + ((!l) & (k) & (!e) & (!a) & (j) & (n)) + ((!l) & (k) & (!e) & (a) & (!j) & (n)) + ((!l) & (k) & (!e) & (a) & (j) & (!n)) + ((!l) & (k) & (!e) & (a) & (j) & (n)) + ((!l) & (k) & (e) & (!a) & (!j) & (n)) + ((!l) & (k) & (e) & (a) & (!j) & (n)) + ((l) & (!k) & (e) & (a) & (j) & (n)) + ((l) & (k) & (!e) & (!a) & (!j) & (!n)) + ((l) & (k) & (!e) & (a) & (!j) & (!n)) + ((l) & (k) & (!e) & (a) & (!j) & (n)) + ((l) & (k) & (e) & (!a) & (!j) & (n)) + ((l) & (k) & (e) & (a) & (!j) & (n)));
	assign g182 = (((!g180) & (g181) & (i)) + ((g180) & (!g181) & (!i)) + ((g180) & (g181) & (!i)) + ((g180) & (g181) & (i)));
	assign g183 = (((!g184) & (!g185)));
	assign g184 = (((!k) & (g186)));
	assign g185 = (((k) & (g189)));
	assign g186 = (((!g187) & (!g188)));
	assign g187 = (((!j) & (g190)));
	assign g188 = (((j) & (g191)));
	assign g189 = (((!j) & (g192)));
	assign g190 = (((!h) & (d) & (g147) & (i)) + ((h) & (!d) & (g147) & (i)) + ((h) & (d) & (!g147) & (i)) + ((h) & (d) & (g147) & (i)));
	assign g191 = (((h) & (d) & (g12) & (!i)));
	assign g192 = (((!h) & (d) & (g147) & (i)) + ((h) & (!d) & (g147) & (i)) + ((h) & (d) & (!g147) & (i)) + ((h) & (d) & (g147) & (i)));
	assign q = (((!g194) & (!g195)));
	assign g194 = (((!n) & (g196)));
	assign g195 = (((n) & (g199)));
	assign g196 = (((!g197) & (!g198)));
	assign g197 = (((!j) & (g202)));
	assign g198 = (((j) & (g203)));
	assign g199 = (((!g200) & (!g201)));
	assign g200 = (((!j) & (g204)));
	assign g201 = (((j) & (g205)));
	assign g202 = (((!g119) & (g116)) + ((g119) & (!g116)) + ((g119) & (g116)));
	assign g203 = (((!g119) & (g117)) + ((g119) & (!g117)) + ((g119) & (g117)));
	assign g204 = (((!g119) & (!g115) & (!g80)) + ((!g119) & (g115) & (g80)) + ((g119) & (!g115) & (!g80)) + ((g119) & (!g115) & (g80)) + ((g119) & (g115) & (!g80)) + ((g119) & (g115) & (g80)));
	assign g205 = (((!g119) & (!g115) & (!g80)) + ((!g119) & (g115) & (g80)) + ((g119) & (!g115) & (!g80)) + ((g119) & (!g115) & (g80)) + ((g119) & (g115) & (!g80)) + ((g119) & (g115) & (g80)));
	assign g206 = (((!g207) & (!g208)));
	assign g207 = (((!g50) & (g209)));
	assign g208 = (((g50) & (g212)));
	assign g209 = (((!g210) & (!g211)));
	assign g210 = (((!b) & (g215)));
	assign g211 = (((b) & (g216)));
	assign g212 = (((!g213) & (!g214)));
	assign g213 = (((!b) & (g217)));
	assign g214 = (((b) & (g218)));
	assign g215 = (((!g56) & (g51) & (g44)) + ((g56) & (!g51) & (g44)) + ((g56) & (g51) & (g44)));
	assign g216 = (((!g56) & (!g57) & (g53) & (!g44)) + ((!g56) & (g57) & (!g53) & (!g44)) + ((!g56) & (g57) & (!g53) & (g44)) + ((!g56) & (g57) & (g53) & (!g44)) + ((!g56) & (g57) & (g53) & (g44)) + ((g56) & (!g57) & (!g53) & (g44)) + ((g56) & (!g57) & (g53) & (!g44)) + ((g56) & (!g57) & (g53) & (g44)) + ((g56) & (g57) & (!g53) & (!g44)) + ((g56) & (g57) & (!g53) & (g44)) + ((g56) & (g57) & (g53) & (!g44)) + ((g56) & (g57) & (g53) & (g44)));
	assign g217 = (((g56) & (g44)));
	assign g218 = (((!g56) & (!g57) & (g53) & (g44)) + ((!g56) & (g57) & (!g53) & (!g44)) + ((!g56) & (g57) & (!g53) & (g44)) + ((!g56) & (g57) & (g53) & (!g44)) + ((!g56) & (g57) & (g53) & (g44)) + ((g56) & (!g57) & (!g53) & (g44)) + ((g56) & (!g57) & (g53) & (g44)) + ((g56) & (g57) & (!g53) & (!g44)) + ((g56) & (g57) & (!g53) & (g44)) + ((g56) & (g57) & (g53) & (!g44)) + ((g56) & (g57) & (g53) & (g44)));
	assign o = (((!g220) & (!g221)));
	assign g220 = (((!n) & (g222)));
	assign g221 = (((n) & (g225)));
	assign g222 = (((!g223) & (!g224)));
	assign g223 = (((!j) & (g228)));
	assign g224 = (((j) & (g229)));
	assign g225 = (((!g226) & (!g227)));
	assign g226 = (((!j) & (g230)));
	assign g227 = (((j) & (g231)));
	assign g228 = (((!g37) & (g5)) + ((g37) & (!g5)) + ((g37) & (g5)));
	assign g229 = (((!g37) & (g6)) + ((g37) & (!g6)) + ((g37) & (g6)));
	assign g230 = (((!g37) & (!g31) & (!m)) + ((!g37) & (g31) & (m)) + ((g37) & (!g31) & (!m)) + ((g37) & (!g31) & (m)) + ((g37) & (g31) & (!m)) + ((g37) & (g31) & (m)));
	assign g231 = (((!g37) & (!g31) & (!m)) + ((!g37) & (g31) & (m)) + ((g37) & (!g31) & (!m)) + ((g37) & (!g31) & (m)) + ((g37) & (g31) & (!m)) + ((g37) & (g31) & (m)));
endmodule
