module sqrt_qmap_o (input [127:0] a, output [63:0] asqrt);




	wire g3496, g3400, g3395, g3187, g3178, g2980, g3030, g2779, g2825, g2585, g2627;
	wire g2398, g2436, g2218, g2252, g2045, g2075, g1879, g1905, g1720, g1742, g1568;
	wire g1586, g1423, g1437, g1285, g1295, g1154, g1160, g1030, g1032, g914, g851;
	wire g803, g744, g700, g645, g604, g553, g515, g468, g433, g390, g358;
	wire g319, g290, g255, g229, g198, g174, g147, g127, g104, g87, g68;
	wire g54, g39, g27, g18, g8, g2, g4, g1, g3, g5, g6;
	wire g7, g9, g10, g11, g12, g13, g14, g15, g16, g17, g19;
	wire g20, g21, g22, g23, g24, g25, g26, g28, g29, g30, g31;
	wire g32, g33, g34, g35, g36, g37, g38, g40, g41, g42, g43;
	wire g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g55;
	wire g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66;
	wire g67, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78;
	wire g79, g80, g81, g82, g83, g84, g85, g86, g88, g89, g90;
	wire g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101;
	wire g102, g103, g105, g106, g107, g108, g109, g110, g111, g112, g113;
	wire g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124;
	wire g125, g126, g128, g129, g130, g131, g132, g133, g134, g135, g136;
	wire g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g148;
	wire g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159;
	wire g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g170;
	wire g171, g172, g173, g175, g176, g177, g178, g179, g180, g181, g182;
	wire g183, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193;
	wire g194, g195, g196, g197, g199, g200, g201, g202, g203, g204, g205;
	wire g206, g207, g208, g209, g210, g211, g212, g213, g214, g215, g216;
	wire g217, g218, g219, g220, g221, g222, g223, g224, g225, g226, g227;
	wire g228, g230, g231, g232, g233, g234, g235, g236, g237, g238, g239;
	wire g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250;
	wire g251, g252, g253, g254, g256, g257, g258, g259, g260, g261, g262;
	wire g263, g264, g265, g266, g267, g268, g269, g270, g271, g272, g273;
	wire g274, g275, g276, g277, g278, g279, g280, g281, g282, g283, g284;
	wire g285, g286, g287, g288, g289, g291, g292, g293, g294, g295, g296;
	wire g297, g298, g299, g300, g301, g302, g303, g304, g305, g306, g307;
	wire g308, g309, g310, g311, g312, g313, g314, g315, g316, g317, g318;
	wire g320, g321, g322, g323, g324, g325, g326, g327, g328, g329, g330;
	wire g331, g332, g333, g334, g335, g336, g337, g338, g339, g340, g341;
	wire g342, g343, g344, g345, g346, g347, g348, g349, g350, g351, g352;
	wire g353, g354, g355, g356, g357, g359, g360, g361, g362, g363, g364;
	wire g365, g366, g367, g368, g369, g370, g371, g372, g373, g374, g375;
	wire g376, g377, g378, g379, g380, g381, g382, g383, g384, g385, g386;
	wire g387, g388, g389, g391, g392, g393, g394, g395, g396, g397, g398;
	wire g399, g400, g401, g402, g403, g404, g405, g406, g407, g408, g409;
	wire g410, g411, g412, g413, g414, g415, g416, g417, g418, g419, g420;
	wire g421, g422, g423, g424, g425, g426, g427, g428, g429, g430, g431;
	wire g432, g434, g435, g436, g437, g438, g439, g440, g441, g442, g443;
	wire g444, g445, g446, g447, g448, g449, g450, g451, g452, g453, g454;
	wire g455, g456, g457, g458, g459, g460, g461, g462, g463, g464, g465;
	wire g466, g467, g469, g470, g471, g472, g473, g474, g475, g476, g477;
	wire g478, g479, g480, g481, g482, g483, g484, g485, g486, g487, g488;
	wire g489, g490, g491, g492, g493, g494, g495, g496, g497, g498, g499;
	wire g500, g501, g502, g503, g504, g505, g506, g507, g508, g509, g510;
	wire g511, g512, g513, g514, g516, g517, g518, g519, g520, g521, g522;
	wire g523, g524, g525, g526, g527, g528, g529, g530, g531, g532, g533;
	wire g534, g535, g536, g537, g538, g539, g540, g541, g542, g543, g544;
	wire g545, g546, g547, g548, g549, g550, g551, g552, g554, g555, g556;
	wire g557, g558, g559, g560, g561, g562, g563, g564, g565, g566, g567;
	wire g568, g569, g570, g571, g572, g573, g574, g575, g576, g577, g578;
	wire g579, g580, g581, g582, g583, g584, g585, g586, g587, g588, g589;
	wire g590, g591, g592, g593, g594, g595, g596, g597, g598, g599, g600;
	wire g601, g602, g603, g605, g606, g607, g608, g609, g610, g611, g612;
	wire g613, g614, g615, g616, g617, g618, g619, g620, g621, g622, g623;
	wire g624, g625, g626, g627, g628, g629, g630, g631, g632, g633, g634;
	wire g635, g636, g637, g638, g639, g640, g641, g642, g643, g644, g646;
	wire g647, g648, g649, g650, g651, g652, g653, g654, g655, g656, g657;
	wire g658, g659, g660, g661, g662, g663, g664, g665, g666, g667, g668;
	wire g669, g670, g671, g672, g673, g674, g675, g676, g677, g678, g679;
	wire g680, g681, g682, g683, g684, g685, g686, g687, g688, g689, g690;
	wire g691, g692, g693, g694, g695, g696, g697, g698, g699, g701, g702;
	wire g703, g704, g705, g706, g707, g708, g709, g710, g711, g712, g713;
	wire g714, g715, g716, g717, g718, g719, g720, g721, g722, g723, g724;
	wire g725, g726, g727, g728, g729, g730, g731, g732, g733, g734, g735;
	wire g736, g737, g738, g739, g740, g741, g742, g743, g745, g746, g747;
	wire g748, g749, g750, g751, g752, g753, g754, g755, g756, g757, g758;
	wire g759, g760, g761, g762, g763, g764, g765, g766, g767, g768, g769;
	wire g770, g771, g772, g773, g774, g775, g776, g777, g778, g779, g780;
	wire g781, g782, g783, g784, g785, g786, g787, g788, g789, g790, g791;
	wire g792, g793, g794, g795, g796, g797, g798, g799, g800, g801, g802;
	wire g804, g805, g806, g807, g808, g809, g810, g811, g812, g813, g814;
	wire g815, g816, g817, g818, g819, g820, g821, g822, g823, g824, g825;
	wire g826, g827, g828, g829, g830, g831, g832, g833, g834, g835, g836;
	wire g837, g838, g839, g840, g841, g842, g843, g844, g845, g846, g847;
	wire g848, g849, g850, g852, g853, g854, g855, g856, g857, g858, g859;
	wire g860, g861, g862, g863, g864, g865, g866, g867, g868, g869, g870;
	wire g871, g872, g873, g874, g875, g876, g877, g878, g879, g880, g881;
	wire g882, g883, g884, g885, g886, g887, g888, g889, g890, g891, g892;
	wire g893, g894, g895, g896, g897, g898, g899, g900, g901, g902, g903;
	wire g904, g905, g906, g907, g908, g909, g910, g911, g912, g913, g915;
	wire g916, g917, g918, g919, g920, g921, g922, g923, g924, g925, g926;
	wire g927, g928, g929, g930, g931, g932, g933, g934, g935, g936, g937;
	wire g938, g939, g940, g941, g942, g943, g944, g945, g946, g947, g948;
	wire g949, g950, g951, g952, g953, g954, g955, g956, g957, g958, g959;
	wire g960, g961, g962, g963, g964, g965, g966, g967, g968, g969, g970;
	wire g971, g972, g973, g974, g975, g976, g977, g978, g979, g980, g981;
	wire g982, g983, g984, g985, g986, g987, g988, g989, g990, g991, g992;
	wire g993, g994, g995, g996, g997, g998, g999, g1000, g1001, g1002, g1003;
	wire g1004, g1005, g1006, g1007, g1008, g1009, g1010, g1011, g1012, g1013, g1014;
	wire g1015, g1016, g1017, g1018, g1019, g1020, g1021, g1022, g1023, g1024, g1025;
	wire g1026, g1027, g1028, g1029, g1031, g1033, g1034, g1035, g1036, g1037, g1038;
	wire g1039, g1040, g1041, g1042, g1043, g1044, g1045, g1046, g1047, g1048, g1049;
	wire g1050, g1051, g1052, g1053, g1054, g1055, g1056, g1057, g1058, g1059, g1060;
	wire g1061, g1062, g1063, g1064, g1065, g1066, g1067, g1068, g1069, g1070, g1071;
	wire g1072, g1073, g1074, g1075, g1076, g1077, g1078, g1079, g1080, g1081, g1082;
	wire g1083, g1084, g1085, g1086, g1087, g1088, g1089, g1090, g1091, g1092, g1093;
	wire g1094, g1095, g1096, g1097, g1098, g1099, g1100, g1101, g1102, g1103, g1104;
	wire g1105, g1106, g1107, g1108, g1109, g1110, g1111, g1112, g1113, g1114, g1115;
	wire g1116, g1117, g1118, g1119, g1120, g1121, g1122, g1123, g1124, g1125, g1126;
	wire g1127, g1128, g1129, g1130, g1131, g1132, g1133, g1134, g1135, g1136, g1137;
	wire g1138, g1139, g1140, g1141, g1142, g1143, g1144, g1145, g1146, g1147, g1148;
	wire g1149, g1150, g1151, g1152, g1153, g1155, g1156, g1157, g1158, g1159, g1161;
	wire g1162, g1163, g1164, g1165, g1166, g1167, g1168, g1169, g1170, g1171, g1172;
	wire g1173, g1174, g1175, g1176, g1177, g1178, g1179, g1180, g1181, g1182, g1183;
	wire g1184, g1185, g1186, g1187, g1188, g1189, g1190, g1191, g1192, g1193, g1194;
	wire g1195, g1196, g1197, g1198, g1199, g1200, g1201, g1202, g1203, g1204, g1205;
	wire g1206, g1207, g1208, g1209, g1210, g1211, g1212, g1213, g1214, g1215, g1216;
	wire g1217, g1218, g1219, g1220, g1221, g1222, g1223, g1224, g1225, g1226, g1227;
	wire g1228, g1229, g1230, g1231, g1232, g1233, g1234, g1235, g1236, g1237, g1238;
	wire g1239, g1240, g1241, g1242, g1243, g1244, g1245, g1246, g1247, g1248, g1249;
	wire g1250, g1251, g1252, g1253, g1254, g1255, g1256, g1257, g1258, g1259, g1260;
	wire g1261, g1262, g1263, g1264, g1265, g1266, g1267, g1268, g1269, g1270, g1271;
	wire g1272, g1273, g1274, g1275, g1276, g1277, g1278, g1279, g1280, g1281, g1282;
	wire g1283, g1284, g1286, g1287, g1288, g1289, g1290, g1291, g1292, g1293, g1294;
	wire g1296, g1297, g1298, g1299, g1300, g1301, g1302, g1303, g1304, g1305, g1306;
	wire g1307, g1308, g1309, g1310, g1311, g1312, g1313, g1314, g1315, g1316, g1317;
	wire g1318, g1319, g1320, g1321, g1322, g1323, g1324, g1325, g1326, g1327, g1328;
	wire g1329, g1330, g1331, g1332, g1333, g1334, g1335, g1336, g1337, g1338, g1339;
	wire g1340, g1341, g1342, g1343, g1344, g1345, g1346, g1347, g1348, g1349, g1350;
	wire g1351, g1352, g1353, g1354, g1355, g1356, g1357, g1358, g1359, g1360, g1361;
	wire g1362, g1363, g1364, g1365, g1366, g1367, g1368, g1369, g1370, g1371, g1372;
	wire g1373, g1374, g1375, g1376, g1377, g1378, g1379, g1380, g1381, g1382, g1383;
	wire g1384, g1385, g1386, g1387, g1388, g1389, g1390, g1391, g1392, g1393, g1394;
	wire g1395, g1396, g1397, g1398, g1399, g1400, g1401, g1402, g1403, g1404, g1405;
	wire g1406, g1407, g1408, g1409, g1410, g1411, g1412, g1413, g1414, g1415, g1416;
	wire g1417, g1418, g1419, g1420, g1421, g1422, g1424, g1425, g1426, g1427, g1428;
	wire g1429, g1430, g1431, g1432, g1433, g1434, g1435, g1436, g1438, g1439, g1440;
	wire g1441, g1442, g1443, g1444, g1445, g1446, g1447, g1448, g1449, g1450, g1451;
	wire g1452, g1453, g1454, g1455, g1456, g1457, g1458, g1459, g1460, g1461, g1462;
	wire g1463, g1464, g1465, g1466, g1467, g1468, g1469, g1470, g1471, g1472, g1473;
	wire g1474, g1475, g1476, g1477, g1478, g1479, g1480, g1481, g1482, g1483, g1484;
	wire g1485, g1486, g1487, g1488, g1489, g1490, g1491, g1492, g1493, g1494, g1495;
	wire g1496, g1497, g1498, g1499, g1500, g1501, g1502, g1503, g1504, g1505, g1506;
	wire g1507, g1508, g1509, g1510, g1511, g1512, g1513, g1514, g1515, g1516, g1517;
	wire g1518, g1519, g1520, g1521, g1522, g1523, g1524, g1525, g1526, g1527, g1528;
	wire g1529, g1530, g1531, g1532, g1533, g1534, g1535, g1536, g1537, g1538, g1539;
	wire g1540, g1541, g1542, g1543, g1544, g1545, g1546, g1547, g1548, g1549, g1550;
	wire g1551, g1552, g1553, g1554, g1555, g1556, g1557, g1558, g1559, g1560, g1561;
	wire g1562, g1563, g1564, g1565, g1566, g1567, g1569, g1570, g1571, g1572, g1573;
	wire g1574, g1575, g1576, g1577, g1578, g1579, g1580, g1581, g1582, g1583, g1584;
	wire g1585, g1587, g1588, g1589, g1590, g1591, g1592, g1593, g1594, g1595, g1596;
	wire g1597, g1598, g1599, g1600, g1601, g1602, g1603, g1604, g1605, g1606, g1607;
	wire g1608, g1609, g1610, g1611, g1612, g1613, g1614, g1615, g1616, g1617, g1618;
	wire g1619, g1620, g1621, g1622, g1623, g1624, g1625, g1626, g1627, g1628, g1629;
	wire g1630, g1631, g1632, g1633, g1634, g1635, g1636, g1637, g1638, g1639, g1640;
	wire g1641, g1642, g1643, g1644, g1645, g1646, g1647, g1648, g1649, g1650, g1651;
	wire g1652, g1653, g1654, g1655, g1656, g1657, g1658, g1659, g1660, g1661, g1662;
	wire g1663, g1664, g1665, g1666, g1667, g1668, g1669, g1670, g1671, g1672, g1673;
	wire g1674, g1675, g1676, g1677, g1678, g1679, g1680, g1681, g1682, g1683, g1684;
	wire g1685, g1686, g1687, g1688, g1689, g1690, g1691, g1692, g1693, g1694, g1695;
	wire g1696, g1697, g1698, g1699, g1700, g1701, g1702, g1703, g1704, g1705, g1706;
	wire g1707, g1708, g1709, g1710, g1711, g1712, g1713, g1714, g1715, g1716, g1717;
	wire g1718, g1719, g1721, g1722, g1723, g1724, g1725, g1726, g1727, g1728, g1729;
	wire g1730, g1731, g1732, g1733, g1734, g1735, g1736, g1737, g1738, g1739, g1740;
	wire g1741, g1743, g1744, g1745, g1746, g1747, g1748, g1749, g1750, g1751, g1752;
	wire g1753, g1754, g1755, g1756, g1757, g1758, g1759, g1760, g1761, g1762, g1763;
	wire g1764, g1765, g1766, g1767, g1768, g1769, g1770, g1771, g1772, g1773, g1774;
	wire g1775, g1776, g1777, g1778, g1779, g1780, g1781, g1782, g1783, g1784, g1785;
	wire g1786, g1787, g1788, g1789, g1790, g1791, g1792, g1793, g1794, g1795, g1796;
	wire g1797, g1798, g1799, g1800, g1801, g1802, g1803, g1804, g1805, g1806, g1807;
	wire g1808, g1809, g1810, g1811, g1812, g1813, g1814, g1815, g1816, g1817, g1818;
	wire g1819, g1820, g1821, g1822, g1823, g1824, g1825, g1826, g1827, g1828, g1829;
	wire g1830, g1831, g1832, g1833, g1834, g1835, g1836, g1837, g1838, g1839, g1840;
	wire g1841, g1842, g1843, g1844, g1845, g1846, g1847, g1848, g1849, g1850, g1851;
	wire g1852, g1853, g1854, g1855, g1856, g1857, g1858, g1859, g1860, g1861, g1862;
	wire g1863, g1864, g1865, g1866, g1867, g1868, g1869, g1870, g1871, g1872, g1873;
	wire g1874, g1875, g1876, g1877, g1878, g1880, g1881, g1882, g1883, g1884, g1885;
	wire g1886, g1887, g1888, g1889, g1890, g1891, g1892, g1893, g1894, g1895, g1896;
	wire g1897, g1898, g1899, g1900, g1901, g1902, g1903, g1904, g1906, g1907, g1908;
	wire g1909, g1910, g1911, g1912, g1913, g1914, g1915, g1916, g1917, g1918, g1919;
	wire g1920, g1921, g1922, g1923, g1924, g1925, g1926, g1927, g1928, g1929, g1930;
	wire g1931, g1932, g1933, g1934, g1935, g1936, g1937, g1938, g1939, g1940, g1941;
	wire g1942, g1943, g1944, g1945, g1946, g1947, g1948, g1949, g1950, g1951, g1952;
	wire g1953, g1954, g1955, g1956, g1957, g1958, g1959, g1960, g1961, g1962, g1963;
	wire g1964, g1965, g1966, g1967, g1968, g1969, g1970, g1971, g1972, g1973, g1974;
	wire g1975, g1976, g1977, g1978, g1979, g1980, g1981, g1982, g1983, g1984, g1985;
	wire g1986, g1987, g1988, g1989, g1990, g1991, g1992, g1993, g1994, g1995, g1996;
	wire g1997, g1998, g1999, g2000, g2001, g2002, g2003, g2004, g2005, g2006, g2007;
	wire g2008, g2009, g2010, g2011, g2012, g2013, g2014, g2015, g2016, g2017, g2018;
	wire g2019, g2020, g2021, g2022, g2023, g2024, g2025, g2026, g2027, g2028, g2029;
	wire g2030, g2031, g2032, g2033, g2034, g2035, g2036, g2037, g2038, g2039, g2040;
	wire g2041, g2042, g2043, g2044, g2046, g2047, g2048, g2049, g2050, g2051, g2052;
	wire g2053, g2054, g2055, g2056, g2057, g2058, g2059, g2060, g2061, g2062, g2063;
	wire g2064, g2065, g2066, g2067, g2068, g2069, g2070, g2071, g2072, g2073, g2074;
	wire g2076, g2077, g2078, g2079, g2080, g2081, g2082, g2083, g2084, g2085, g2086;
	wire g2087, g2088, g2089, g2090, g2091, g2092, g2093, g2094, g2095, g2096, g2097;
	wire g2098, g2099, g2100, g2101, g2102, g2103, g2104, g2105, g2106, g2107, g2108;
	wire g2109, g2110, g2111, g2112, g2113, g2114, g2115, g2116, g2117, g2118, g2119;
	wire g2120, g2121, g2122, g2123, g2124, g2125, g2126, g2127, g2128, g2129, g2130;
	wire g2131, g2132, g2133, g2134, g2135, g2136, g2137, g2138, g2139, g2140, g2141;
	wire g2142, g2143, g2144, g2145, g2146, g2147, g2148, g2149, g2150, g2151, g2152;
	wire g2153, g2154, g2155, g2156, g2157, g2158, g2159, g2160, g2161, g2162, g2163;
	wire g2164, g2165, g2166, g2167, g2168, g2169, g2170, g2171, g2172, g2173, g2174;
	wire g2175, g2176, g2177, g2178, g2179, g2180, g2181, g2182, g2183, g2184, g2185;
	wire g2186, g2187, g2188, g2189, g2190, g2191, g2192, g2193, g2194, g2195, g2196;
	wire g2197, g2198, g2199, g2200, g2201, g2202, g2203, g2204, g2205, g2206, g2207;
	wire g2208, g2209, g2210, g2211, g2212, g2213, g2214, g2215, g2216, g2217, g2219;
	wire g2220, g2221, g2222, g2223, g2224, g2225, g2226, g2227, g2228, g2229, g2230;
	wire g2231, g2232, g2233, g2234, g2235, g2236, g2237, g2238, g2239, g2240, g2241;
	wire g2242, g2243, g2244, g2245, g2246, g2247, g2248, g2249, g2250, g2251, g2253;
	wire g2254, g2255, g2256, g2257, g2258, g2259, g2260, g2261, g2262, g2263, g2264;
	wire g2265, g2266, g2267, g2268, g2269, g2270, g2271, g2272, g2273, g2274, g2275;
	wire g2276, g2277, g2278, g2279, g2280, g2281, g2282, g2283, g2284, g2285, g2286;
	wire g2287, g2288, g2289, g2290, g2291, g2292, g2293, g2294, g2295, g2296, g2297;
	wire g2298, g2299, g2300, g2301, g2302, g2303, g2304, g2305, g2306, g2307, g2308;
	wire g2309, g2310, g2311, g2312, g2313, g2314, g2315, g2316, g2317, g2318, g2319;
	wire g2320, g2321, g2322, g2323, g2324, g2325, g2326, g2327, g2328, g2329, g2330;
	wire g2331, g2332, g2333, g2334, g2335, g2336, g2337, g2338, g2339, g2340, g2341;
	wire g2342, g2343, g2344, g2345, g2346, g2347, g2348, g2349, g2350, g2351, g2352;
	wire g2353, g2354, g2355, g2356, g2357, g2358, g2359, g2360, g2361, g2362, g2363;
	wire g2364, g2365, g2366, g2367, g2368, g2369, g2370, g2371, g2372, g2373, g2374;
	wire g2375, g2376, g2377, g2378, g2379, g2380, g2381, g2382, g2383, g2384, g2385;
	wire g2386, g2387, g2388, g2389, g2390, g2391, g2392, g2393, g2394, g2395, g2396;
	wire g2397, g2399, g2400, g2401, g2402, g2403, g2404, g2405, g2406, g2407, g2408;
	wire g2409, g2410, g2411, g2412, g2413, g2414, g2415, g2416, g2417, g2418, g2419;
	wire g2420, g2421, g2422, g2423, g2424, g2425, g2426, g2427, g2428, g2429, g2430;
	wire g2431, g2432, g2433, g2434, g2435, g2437, g2438, g2439, g2440, g2441, g2442;
	wire g2443, g2444, g2445, g2446, g2447, g2448, g2449, g2450, g2451, g2452, g2453;
	wire g2454, g2455, g2456, g2457, g2458, g2459, g2460, g2461, g2462, g2463, g2464;
	wire g2465, g2466, g2467, g2468, g2469, g2470, g2471, g2472, g2473, g2474, g2475;
	wire g2476, g2477, g2478, g2479, g2480, g2481, g2482, g2483, g2484, g2485, g2486;
	wire g2487, g2488, g2489, g2490, g2491, g2492, g2493, g2494, g2495, g2496, g2497;
	wire g2498, g2499, g2500, g2501, g2502, g2503, g2504, g2505, g2506, g2507, g2508;
	wire g2509, g2510, g2511, g2512, g2513, g2514, g2515, g2516, g2517, g2518, g2519;
	wire g2520, g2521, g2522, g2523, g2524, g2525, g2526, g2527, g2528, g2529, g2530;
	wire g2531, g2532, g2533, g2534, g2535, g2536, g2537, g2538, g2539, g2540, g2541;
	wire g2542, g2543, g2544, g2545, g2546, g2547, g2548, g2549, g2550, g2551, g2552;
	wire g2553, g2554, g2555, g2556, g2557, g2558, g2559, g2560, g2561, g2562, g2563;
	wire g2564, g2565, g2566, g2567, g2568, g2569, g2570, g2571, g2572, g2573, g2574;
	wire g2575, g2576, g2577, g2578, g2579, g2580, g2581, g2582, g2583, g2584, g2586;
	wire g2587, g2588, g2589, g2590, g2591, g2592, g2593, g2594, g2595, g2596, g2597;
	wire g2598, g2599, g2600, g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608;
	wire g2609, g2610, g2611, g2612, g2613, g2614, g2615, g2616, g2617, g2618, g2619;
	wire g2620, g2621, g2622, g2623, g2624, g2625, g2626, g2628, g2629, g2630, g2631;
	wire g2632, g2633, g2634, g2635, g2636, g2637, g2638, g2639, g2640, g2641, g2642;
	wire g2643, g2644, g2645, g2646, g2647, g2648, g2649, g2650, g2651, g2652, g2653;
	wire g2654, g2655, g2656, g2657, g2658, g2659, g2660, g2661, g2662, g2663, g2664;
	wire g2665, g2666, g2667, g2668, g2669, g2670, g2671, g2672, g2673, g2674, g2675;
	wire g2676, g2677, g2678, g2679, g2680, g2681, g2682, g2683, g2684, g2685, g2686;
	wire g2687, g2688, g2689, g2690, g2691, g2692, g2693, g2694, g2695, g2696, g2697;
	wire g2698, g2699, g2700, g2701, g2702, g2703, g2704, g2705, g2706, g2707, g2708;
	wire g2709, g2710, g2711, g2712, g2713, g2714, g2715, g2716, g2717, g2718, g2719;
	wire g2720, g2721, g2722, g2723, g2724, g2725, g2726, g2727, g2728, g2729, g2730;
	wire g2731, g2732, g2733, g2734, g2735, g2736, g2737, g2738, g2739, g2740, g2741;
	wire g2742, g2743, g2744, g2745, g2746, g2747, g2748, g2749, g2750, g2751, g2752;
	wire g2753, g2754, g2755, g2756, g2757, g2758, g2759, g2760, g2761, g2762, g2763;
	wire g2764, g2765, g2766, g2767, g2768, g2769, g2770, g2771, g2772, g2773, g2774;
	wire g2775, g2776, g2777, g2778, g2780, g2781, g2782, g2783, g2784, g2785, g2786;
	wire g2787, g2788, g2789, g2790, g2791, g2792, g2793, g2794, g2795, g2796, g2797;
	wire g2798, g2799, g2800, g2801, g2802, g2803, g2804, g2805, g2806, g2807, g2808;
	wire g2809, g2810, g2811, g2812, g2813, g2814, g2815, g2816, g2817, g2818, g2819;
	wire g2820, g2821, g2822, g2823, g2824, g2826, g2827, g2828, g2829, g2830, g2831;
	wire g2832, g2833, g2834, g2835, g2836, g2837, g2838, g2839, g2840, g2841, g2842;
	wire g2843, g2844, g2845, g2846, g2847, g2848, g2849, g2850, g2851, g2852, g2853;
	wire g2854, g2855, g2856, g2857, g2858, g2859, g2860, g2861, g2862, g2863, g2864;
	wire g2865, g2866, g2867, g2868, g2869, g2870, g2871, g2872, g2873, g2874, g2875;
	wire g2876, g2877, g2878, g2879, g2880, g2881, g2882, g2883, g2884, g2885, g2886;
	wire g2887, g2888, g2889, g2890, g2891, g2892, g2893, g2894, g2895, g2896, g2897;
	wire g2898, g2899, g2900, g2901, g2902, g2903, g2904, g2905, g2906, g2907, g2908;
	wire g2909, g2910, g2911, g2912, g2913, g2914, g2915, g2916, g2917, g2918, g2919;
	wire g2920, g2921, g2922, g2923, g2924, g2925, g2926, g2927, g2928, g2929, g2930;
	wire g2931, g2932, g2933, g2934, g2935, g2936, g2937, g2938, g2939, g2940, g2941;
	wire g2942, g2943, g2944, g2945, g2946, g2947, g2948, g2949, g2950, g2951, g2952;
	wire g2953, g2954, g2955, g2956, g2957, g2958, g2959, g2960, g2961, g2962, g2963;
	wire g2964, g2965, g2966, g2967, g2968, g2969, g2970, g2971, g2972, g2973, g2974;
	wire g2975, g2976, g2977, g2978, g2979, g2981, g2982, g2983, g2984, g2985, g2986;
	wire g2987, g2988, g2989, g2990, g2991, g2992, g2993, g2994, g2995, g2996, g2997;
	wire g2998, g2999, g3000, g3001, g3002, g3003, g3004, g3005, g3006, g3007, g3008;
	wire g3009, g3010, g3011, g3012, g3013, g3014, g3015, g3016, g3017, g3018, g3019;
	wire g3020, g3021, g3022, g3023, g3024, g3025, g3026, g3027, g3028, g3029, g3031;
	wire g3032, g3033, g3034, g3035, g3036, g3037, g3038, g3039, g3040, g3041, g3042;
	wire g3043, g3044, g3045, g3046, g3047, g3048, g3049, g3050, g3051, g3052, g3053;
	wire g3054, g3055, g3056, g3057, g3058, g3059, g3060, g3061, g3062, g3063, g3064;
	wire g3065, g3066, g3067, g3068, g3069, g3070, g3071, g3072, g3073, g3074, g3075;
	wire g3076, g3077, g3078, g3079, g3080, g3081, g3082, g3083, g3084, g3085, g3086;
	wire g3087, g3088, g3089, g3090, g3091, g3092, g3093, g3094, g3095, g3096, g3097;
	wire g3098, g3099, g3100, g3101, g3102, g3103, g3104, g3105, g3106, g3107, g3108;
	wire g3109, g3110, g3111, g3112, g3113, g3114, g3115, g3116, g3117, g3118, g3119;
	wire g3120, g3121, g3122, g3123, g3124, g3125, g3126, g3127, g3128, g3129, g3130;
	wire g3131, g3132, g3133, g3134, g3135, g3136, g3137, g3138, g3139, g3140, g3141;
	wire g3142, g3143, g3144, g3145, g3146, g3147, g3148, g3149, g3150, g3151, g3152;
	wire g3153, g3154, g3155, g3156, g3157, g3158, g3159, g3160, g3161, g3162, g3163;
	wire g3164, g3165, g3166, g3167, g3168, g3169, g3170, g3171, g3172, g3173, g3174;
	wire g3175, g3176, g3177, g3179, g3180, g3181, g3182, g3183, g3184, g3185, g3186;
	wire g3188, g3189, g3190, g3191, g3192, g3193, g3194, g3195, g3196, g3197, g3198;
	wire g3199, g3200, g3201, g3202, g3203, g3204, g3205, g3206, g3207, g3208, g3209;
	wire g3210, g3211, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220;
	wire g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231;
	wire g3232, g3233, g3234, g3235, g3236, g3237, g3238, g3239, g3240, g3241, g3242;
	wire g3243, g3244, g3245, g3246, g3247, g3248, g3249, g3250, g3251, g3252, g3253;
	wire g3254, g3255, g3256, g3257, g3258, g3259, g3260, g3261, g3262, g3263, g3264;
	wire g3265, g3266, g3267, g3268, g3269, g3270, g3271, g3272, g3273, g3274, g3275;
	wire g3276, g3277, g3278, g3279, g3280, g3281, g3282, g3283, g3284, g3285, g3286;
	wire g3287, g3288, g3289, g3290, g3291, g3292, g3293, g3294, g3295, g3296, g3297;
	wire g3298, g3299, g3300, g3301, g3302, g3303, g3304, g3305, g3306, g3307, g3308;
	wire g3309, g3310, g3311, g3312, g3313, g3314, g3315, g3316, g3317, g3318, g3319;
	wire g3320, g3321, g3322, g3323, g3324, g3325, g3326, g3327, g3328, g3329, g3330;
	wire g3331, g3332, g3333, g3334, g3335, g3336, g3337, g3338, g3339, g3340, g3341;
	wire g3342, g3343, g3344, g3345, g3346, g3347, g3348, g3349, g3350, g3351, g3352;
	wire g3353, g3354, g3355, g3356, g3357, g3358, g3359, g3360, g3361, g3362, g3363;
	wire g3364, g3365, g3366, g3367, g3368, g3369, g3370, g3371, g3372, g3373, g3374;
	wire g3375, g3376, g3377, g3378, g3379, g3380, g3381, g3382, g3383, g3384, g3385;
	wire g3386, g3387, g3388, g3389, g3390, g3391, g3392,