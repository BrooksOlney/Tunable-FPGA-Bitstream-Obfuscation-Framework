module pdc_qmap_map (sk, i_5_, i_3_, i_4_, i_1_, i_0_, i_2_, i_8_, i_7_, i_6_, i_9_, i_10_, i_11_, i_15_, i_14_, i_12_, i_13_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_);

	input i_5_;
	input i_3_;
	input i_4_;
	input i_1_;
	input i_0_;
	input i_2_;
	input i_8_;
	input i_7_;
	input i_6_;
	input i_9_;
	input i_10_;
	input i_11_;
	input i_15_;
	input i_14_;
	input i_12_;
	input i_13_;
	output o_0_;
	output o_1_;
	output o_2_;
	output o_3_;
	output o_4_;
	output o_5_;
	output o_6_;
	output o_7_;
	output o_8_;
	output o_9_;
	output o_10_;
	output o_11_;
	output o_12_;
	output o_13_;
	output o_14_;
	output o_15_;
	output o_16_;
	output o_17_;
	output o_18_;
	output o_19_;
	output o_20_;
	output o_21_;
	output o_22_;
	output o_23_;
	output o_24_;
	output o_25_;
	output o_26_;
	output o_27_;
	output o_28_;
	output o_29_;
	output o_30_;
	output o_31_;
	output o_32_;
	output o_33_;
	output o_34_;
	output o_35_;
	output o_36_;
	output o_37_;
	output o_38_;
	output o_39_;



	wire g854, g68, g874, g1029, g1640, g1094, g1137, g29, g1138, g1437, g1467, g1469, g1476, g1477, g1491, g1503, g1506, g1509, g1530, g1, g2;
	wire g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23;
	wire g24, g25, g26, g27, g28, g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44, g45;
	wire g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66;
	wire g67, g69, g70, g71, g72, g73, g75, g76, g77, g78, g79, g80, g81, g82, g1544, g83, g85, g87, g88, g89, g90;
	wire g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111;
	wire g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g132;
	wire g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153;
	wire g154, g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g1775, g168, g1782, g169, g170, g171, g172;
	wire g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193;
	wire g194, g195, g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207, g208, g209, g210, g211, g212, g213, g214;
	wire g215, g216, g217, g218, g219, g220, g221, g222, g223, g224, g225, g226, g227, g228, g229, g230, g231, g232, g233, g234, g1543;
	wire g235, g236, g237, g238, g239, g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250, g251, g252, g253, g254, g255;
	wire g256, g257, g258, g259, g260, g261, g262, g263, g264, g265, g266, g267, g268, g269, g270, g271, g272, g273, g274, g275, g276;
	wire g277, g278, g279, g280, g281, g282, g283, g284, g285, g286, g287, g288, g289, g290, g291, g292, g293, g294, g295, g296, g297;
	wire g298, g299, g300, g301, g302, g303, g304, g305, g306, g307, g308, g309, g310, g311, g312, g313, g314, g315, g316, g317, g318;
	wire g319, g320, g321, g1768, g322, g323, g324, g325, g326, g327, g328, g329, g330, g331, g332, g333, g334, g1761, g335, g336, g337;
	wire g338, g339, g340, g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351, g352, g353, g354, g355, g356, g357, g358;
	wire g359, g360, g361, g362, g363, g364, g365, g366, g367, g368, g369, g370, g371, g372, g373, g1754, g374, g375, g376, g377, g378;
	wire g379, g380, g381, g382, g383, g384, g385, g386, g387, g388, g389, g390, g391, g392, g393, g394, g395, g396, g397, g398, g399;
	wire g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410, g1747, g411, g412, g413, g414, g415, g416, g417, g418, g419;
	wire g420, g421, g422, g423, g424, g425, g426, g427, g428, g429, g430, g431, g432, g433, g434, g435, g436, g437, g438, g439, g440;
	wire g441, g442, g443, g444, g445, g446, g447, g448, g449, g450, g451, g452, g453, g454, g455, g456, g457, g458, g460, g461, g462;
	wire g463, g464, g465, g466, g467, g468, g469, g470, g471, g472, g473, g474, g475, g476, g477, g478, g479, g480, g481, g482, g483;
	wire g484, g485, g486, g487, g488, g489, g490, g491, g492, g493, g494, g495, g496, g497, g498, g499, g500, g501, g502, g503, g504;
	wire g505, g506, g507, g508, g509, g510, g511, g512, g513, g514, g515, g516, g517, g518, g519, g520, g1737, g1728, g521, g522, g523;
	wire g524, g525, g526, g527, g528, g529, g530, g531, g532, g533, g534, g535, g536, g537, g538, g539, g540, g541, g542, g1721, g543;
	wire g544, g545, g546, g547, g548, g549, g550, g551, g552, g553, g554, g555, g556, g557, g558, g559, g560, g561, g562, g563, g564;
	wire g565, g566, g567, g1708, g568, g569, g570, g571, g572, g573, g574, g575, g576, g577, g578, g579, g580, g581, g582, g583, g584;
	wire g585, g586, g587, g588, g589, g590, g591, g592, g593, g594, g595, g596, g597, g598, g599, g600, g601, g602, g603, g604, g605;
	wire g606, g1695, g607, g608, g609, g610, g611, g612, g613, g614, g615, g616, g617, g618, g619, g620, g621, g622, g623, g624, g625;
	wire g626, g627, g628, g629, g630, g631, g632, g1686, g633, g634, g635, g636, g637, g638, g639, g640, g641, g642, g643, g644, g645;
	wire g646, g647, g648, g649, g650, g651, g652, g653, g654, g655, g656, g657, g658, g659, g660, g661, g662, g663, g664, g666, g667;
	wire g668, g669, g670, g671, g672, g673, g674, g675, g676, g677, g678, g679, g680, g681, g682, g683, g684, g685, g686, g687, g688;
	wire g689, g690, g691, g692, g693, g694, g695, g696, g697, g698, g699, g700, g701, g702, g703, g704, g705, g706, g707, g708, g709;
	wire g710, g711, g712, g713, g714, g715, g716, g717, g718, g719, g720, g721, g722, g723, g724, g725, g726, g727, g728, g729, g730;
	wire g731, g732, g733, g734, g735, g736, g737, g738, g739, g740, g741, g742, g743, g744, g745, g746, g747, g748, g749, g750, g751;
	wire g752, g753, g754, g755, g756, g757, g758, g759, g760, g761, g762, g763, g764, g765, g766, g767, g768, g769, g770, g771, g772;
	wire g773, g774, g775, g776, g777, g778, g779, g780, g781, g782, g783, g784, g785, g786, g787, g788, g789, g790, g791, g792, g793;
	wire g794, g795, g796, g797, g798, g799, g800, g801, g802, g803, g804, g805, g806, g807, g808, g809, g810, g811, g812, g813, g814;
	wire g815, g1673, g1666, g816, g817, g818, g819, g820, g821, g822, g823, g824, g825, g826, g827, g828, g829, g830, g831, g832, g833;
	wire g834, g835, g836, g837, g838, g839, g840, g1653, g841, g842, g843, g844, g845, g846, g847, g848, g849, g850, g851, g852, g853;
	wire g855, g857, g858, g859, g860, g861, g862, g863, g864, g865, g866, g867, g868, g869, g870, g871, g872, g873, g875, g876, g877;
	wire g878, g879, g880, g881, g882, g883, g884, g885, g886, g887, g888, g889, g890, g891, g892, g893, g894, g895, g896, g897, g898;
	wire g899, g900, g901, g902, g903, g904, g905, g906, g907, g908, g909, g910, g911, g912, g913, g914, g915, g916, g917, g918, g919;
	wire g920, g921, g922, g923, g924, g925, g926, g927, g928, g929, g930, g931, g932, g933, g934, g935, g936, g937, g938, g939, g940;
	wire g941, g942, g943, g944, g945, g946, g947, g948, g949, g950, g951, g952, g953, g954, g955, g956, g957, g958, g959, g960, g961;
	wire g962, g963, g964, g965, g966, g967, g968, g970, g971, g972, g973, g974, g975, g976, g977, g978, g979, g980, g981, g982, g983;
	wire g984, g985, g986, g987, g988, g989, g990, g991, g992, g993, g994, g995, g996, g997, g998, g999, g1000, g1001, g1002, g1003, g1004;
	wire g1005, g1006, g1007, g1008, g1009, g1010, g1011, g1012, g1013, g1014, g1015, g1016, g1017, g1018, g1019, g1020, g1021, g1022, g1023, g1024, g1025;
	wire g1026, g1027, g1542, g1028, g1030, g1031, g1032, g1033, g1034, g1035, g1036, g1037, g1038, g1039, g1040, g1041, g1042, g1043, g1044, g1045, g1046;
	wire g1047, g1048, g1049, g1050, g1051, g1052, g1053, g1054, g1055, g1056, g1057, g1058, g1059, g1060, g1061, g1062, g1063, g1064, g1065, g1066, g1067;
	wire g1068, g1069, g1070, g1071, g1072, g1073, g1074, g1075, g1076, g1077, g1078, g1079, g1080, g1081, g1082, g1083, g1084, g1085, g1086, g1087, g1088;
	wire g1089, g1090, g1091, g1092, g1093, g1095, g1096, g1097, g1098, g1099, g1100, g1541, g1101, g1102, g1103, g1104, g1628, g1622, g1105, g1106, g1107;
	wire g1108, g1109, g1110, g1111, g1112, g1113, g1114, g1115, g1116, g1117, g1118, g1616, g1119, g1120, g1121, g1122, g1123, g1124, g1125, g1126, g1127;
	wire g1128, g1129, g1130, g1131, g1132, g1133, g1134, g1135, g1136, g1139, g1140, g1141, g1142, g1143, g1144, g1145, g1146, g1147, g1148, g1149, g1150;
	wire g1151, g1152, g1153, g1154, g1155, g1156, g1157, g1158, g1159, g1160, g1161, g1162, g1163, g1164, g1165, g1166, g1167, g1168, g1169, g1170, g1171;
	wire g1172, g1173, g1174, g1175, g1176, g1177, g1178, g1179, g1180, g1181, g1182, g1183, g1184, g1185, g1186, g1187, g1188, g1189, g1191, g1192, g1193;
	wire g1194, g1195, g1196, g1197, g1198, g1199, g1200, g1201, g1202, g1203, g1204, g1205, g1206, g1207, g1208, g1209, g1210, g1211, g1212, g1213, g1214;
	wire g1215, g1216, g1607, g1217, g1218, g1219, g1220, g1221, g1222, g1223, g1224, g1225, g1226, g1227, g1228, g1229, g1230, g1231, g1232, g1233, g1234;
	wire g1235, g1236, g1237, g1238, g1239, g1240, g1241, g1242, g1243, g1244, g1245, g1246, g1247, g1248, g1249, g1250, g1251, g1252, g1253, g1254, g1255;
	wire g1256, g1257, g1258, g1259, g1260, g1261, g1262, g1263, g1264, g1265, g1266, g1267, g1268, g1269, g1270, g1271, g1272, g1273, g1274, g1275, g1276;
	wire g1277, g1278, g1279, g1280, g1281, g1282, g1283, g1284, g1285, g1286, g1287, g1288, g1289, g1290, g1291, g1292, g1293, g1294, g1295, g1296, g1297;
	wire g1298, g1299, g1596, g1300, g1301, g1303, g1304, g1305, g1306, g1307, g1308, g1309, g1310, g1311, g1312, g1313, g1314, g1315, g1316, g1317, g1318;
	wire g1319, g1320, g1321, g1322, g1323, g1324, g1325, g1326, g1327, g1328, g1329, g1589, g1330, g1331, g1332, g1333, g1334, g1335, g1336, g1337, g1338;
	wire g1339, g1340, g1341, g1342, g1343, g1344, g1345, g1346, g1347, g1348, g1349, g1350, g1351, g1352, g1353, g1354, g1355, g1356, g1357, g1358, g1359;
	wire g1360, g1361, g1362, g1363, g1364, g1365, g1366, g1367, g1368, g1369, g1370, g1371, g1372, g1580, g1373, g1374, g1375, g1376, g1377, g1378, g1379;
	wire g1380, g1381, g1382, g1384, g1385, g1386, g1387, g1388, g1389, g1390, g1391, g1538, g1392, g1393, g1394, g1395, g1396, g1397, g1398, g1399, g1400;
	wire g1401, g1402, g1403, g1404, g1405, g1406, g1407, g1408, g1409, g1410, g1411, g1558, g1412, g1413, g1568, g1415, g1416, g1417, g1418, g1419, g1420;
	wire g1421, g1422, g1423, g1424, g1425, g1426, g1427, g1428, g1429, g1430, g1431, g1432, g1433, g1434, g1435, g1438, g1439, g1441, g1442, g1443, g1444;
	wire g1445, g1446, g1447, g1448, g1449, g1450, g1451, g1545, g1452, g1453, g1454, g1455, g1456, g1457, g1458, g1459, g1460, g1461, g1462, g1463, g1464;
	wire g1465, g1466, g1468, g1470, g1471, g1472, g1473, g1474, g1475, g1479, g1480, g1481, g1482, g1483, g1484, g1485, g1486, g1487, g1488, g1489, g1490;
	wire g1492, g1493, g1494, g1495, g1496, g1497, g1498, g1499, g1501, g1502, g1504, g1507, g1508, g1510, g1511, g1512, g1513, g1514, g1515, g1516, g1517;
	wire g1518, g1519, g1520, g1521, g1522, g1524, g1526, g1527, g1528, g1529, g1531, g1532, g1536, g1537, g1539, g1540, g1546, g1547, g1548, g1551, g1549;
	wire g1550, g1554, g1555, g1552, g1553, g1556, g1557, g1559, g1560, g1561, g1564, g1562, g1563, g1566, g1565, g1567, g1569, g1570, g1571, g1574, g1572;
	wire g1573, g1577, g1578, g1575, g1576, g1579, g1581, g1582, g1583, g1585, g1584, g1587, g1586, g1588, g1590, g1591, g1592, g1593, g1594, g1595, g1597;
	wire g1598, g1599, g1601, g1600, g1604, g1602, g1603, g1605, g1606, g1608, g1609, g1610, g1613, g1611, g1612, g1614, g1615, g1617, g1618, g1619, g1620;
	wire g1621, g1623, g1624, g1625, g1626, g1627, g1629, g1630, g1631, g1634, g1632, g1633, g1637, g1635, g1636, g1638, g1639, g1641, g1642, g1643, g1646;
	wire g1644, g1645, g1649, g1650, g1647, g1648, g1651, g1652, g1654, g1655, g1656, g1659, g1657, g1658, g1662, g1663, g1660, g1661, g1664, g1665, g1667;
	wire g1668, g1669, g1670, g1671, g1672, g1674, g1675, g1676, g1679, g1677, g1678, g1682, g1683, g1680, g1681, g1684, g1685, g1687, g1688, g1689, g1691;
	wire g1690, g1693, g1692, g1694, g1696, g1697, g1698, g1701, g1699, g1700, g1704, g1705, g1702, g1703, g1706, g1707, g1709, g1710, g1711, g1714, g1712;
	wire g1713, g1717, g1718, g1715, g1716, g1719, g1720, g1722, g1723, g1724, g1725, g1726, g1727, g1729, g1730, g1731, g1732, g1733, g1734, g1735, g1736;
	wire g1738, g1739, g1740, g1741, g1744, g1742, g1743, g1745, g1746, g1748, g1749, g1750, g1751, g1752, g1753, g1755, g1756, g1757, g1758, g1759, g1760;
	wire g1762, g1763, g1764, g1765, g1766, g1767, g1769, g1770, g1771, g1772, g1773, g1774, g1776, g1777, g1778, g1779, g1780, g1781, g1783, g1784, g1785;
	wire g1786, g1789, g1787, g1788, g1790, g1791;

	lut_sub lut_5 ({g854}, o_5_);
	defparam lut_5.LUT_SIZE = 1;
	defparam lut_5.mask = 2'b10;

	lut_sub lut_9 ({g68}, o_6_);
	defparam lut_9.LUT_SIZE = 1;
	defparam lut_9.mask = 2'b10;

	lut_sub lut_13 ({g874}, o_8_);
	defparam lut_13.LUT_SIZE = 1;
	defparam lut_13.mask = 2'b10;

	lut_sub lut_17 ({g1029}, o_10_);
	defparam lut_17.LUT_SIZE = 1;
	defparam lut_17.mask = 2'b10;

	lut_sub lut_21 ({g1640}, o_11_);
	defparam lut_21.LUT_SIZE = 1;
	defparam lut_21.mask = 2'b10;

	lut_sub lut_25 ({g1094}, o_12_);
	defparam lut_25.LUT_SIZE = 1;
	defparam lut_25.mask = 2'b10;

	lut_sub lut_29 ({g1137}, o_13_);
	defparam lut_29.LUT_SIZE = 1;
	defparam lut_29.mask = 2'b10;

	lut_sub lut_33 ({g29}, o_14_);
	defparam lut_33.LUT_SIZE = 1;
	defparam lut_33.mask = 2'b01;

	lut_sub lut_37 ({g1138}, o_15_);
	defparam lut_37.LUT_SIZE = 1;
	defparam lut_37.mask = 2'b10;

	lut_sub lut_41 ({g1437}, o_21_);
	defparam lut_41.LUT_SIZE = 1;
	defparam lut_41.mask = 2'b10;

	lut_sub lut_45 ({g1467}, o_23_);
	defparam lut_45.LUT_SIZE = 1;
	defparam lut_45.mask = 2'b10;

	lut_sub lut_49 ({g1469}, o_24_);
	defparam lut_49.LUT_SIZE = 1;
	defparam lut_49.mask = 2'b10;

	lut_sub lut_53 ({g1476}, o_25_);
	defparam lut_53.LUT_SIZE = 1;
	defparam lut_53.mask = 2'b10;

	lut_sub lut_57 ({g1477}, o_26_);
	defparam lut_57.LUT_SIZE = 1;
	defparam lut_57.mask = 2'b10;

	lut_sub lut_61 ({g1491}, o_28_);
	defparam lut_61.LUT_SIZE = 1;
	defparam lut_61.mask = 2'b10;

	lut_sub lut_65 ({g1503}, o_30_);
	defparam lut_65.LUT_SIZE = 1;
	defparam lut_65.mask = 2'b10;

	lut_sub lut_69 ({g1506}, o_32_);
	defparam lut_69.LUT_SIZE = 1;
	defparam lut_69.mask = 2'b10;

	lut_sub lut_73 ({g1509}, o_33_);
	defparam lut_73.LUT_SIZE = 1;
	defparam lut_73.mask = 2'b10;

	lut_sub lut_77 ({g1530}, o_36_);
	defparam lut_77.LUT_SIZE = 1;
	defparam lut_77.mask = 2'b10;

	lut_sub lut_81 ({i_1_, i_0_, i_2_}, g1);
	defparam lut_81.LUT_SIZE = 3;
	defparam lut_81.mask = 8'h08;

	lut_sub lut_86 ({i_5_, i_3_, i_4_, g1}, g2);
	defparam lut_86.LUT_SIZE = 4;
	defparam lut_86.mask = 16'h4000;

	lut_sub lut_91 ({g2, i_8_, i_7_}, g3);
	defparam lut_91.LUT_SIZE = 3;
	defparam lut_91.mask = 8'h02;

	lut_sub lut_95 ({i_6_, i_7_}, g4);
	defparam lut_95.LUT_SIZE = 2;
	defparam lut_95.mask = 4'b0001;

	lut_sub lut_99 ({i_9_, i_10_}, g5);
	defparam lut_99.LUT_SIZE = 2;
	defparam lut_99.mask = 4'b1000;

	lut_sub lut_103 ({i_11_, i_9_, i_10_}, g6);
	defparam lut_103.LUT_SIZE = 3;
	defparam lut_103.mask = 8'h20;

	lut_sub lut_107 ({i_14_, i_12_, i_13_}, g7);
	defparam lut_107.LUT_SIZE = 3;
	defparam lut_107.mask = 8'h80;

	lut_sub lut_113 ({g6, i_15_, g7}, g8);
	defparam lut_113.LUT_SIZE = 3;
	defparam lut_113.mask = 8'hfe;

	lut_sub lut_123 ({i_14_, i_12_, i_13_}, g9);
	defparam lut_123.LUT_SIZE = 3;
	defparam lut_123.mask = 8'h40;

	lut_sub lut_129 ({g6, i_15_, g9}, g10);
	defparam lut_129.LUT_SIZE = 3;
	defparam lut_129.mask = 8'h04;

	lut_sub lut_133 ({i_11_, i_9_, i_10_, i_15_}, g11);
	defparam lut_133.LUT_SIZE = 4;
	defparam lut_133.mask = 16'h0200;

	lut_sub lut_139 ({g11, g9}, g12);
	defparam lut_139.LUT_SIZE = 2;
	defparam lut_139.mask = 4'b0001;

	lut_sub lut_143 ({i_14_, i_12_, i_13_}, g13);
	defparam lut_143.LUT_SIZE = 3;
	defparam lut_143.mask = 8'h08;

	lut_sub lut_149 ({g6, i_15_, g13}, g14);
	defparam lut_149.LUT_SIZE = 3;
	defparam lut_149.mask = 8'h04;

	lut_sub lut_153 ({i_11_, i_9_, i_10_, i_15_}, g15);
	defparam lut_153.LUT_SIZE = 4;
	defparam lut_153.mask = 16'hdfff;

	lut_sub lut_173 ({g15, g9}, g16);
	defparam lut_173.LUT_SIZE = 2;
	defparam lut_173.mask = 4'b1011;

	lut_sub lut_182 ({g12, g14, g16}, g17);
	defparam lut_182.LUT_SIZE = 3;
	defparam lut_182.mask = 8'h40;

	lut_sub lut_186 ({i_11_, i_9_, i_10_, i_15_}, g18);
	defparam lut_186.LUT_SIZE = 4;
	defparam lut_186.mask = 16'hefff;

	lut_sub lut_206 ({g7, g18}, g19);
	defparam lut_206.LUT_SIZE = 2;
	defparam lut_206.mask = 4'b0010;

	lut_sub lut_212 ({g15, g13}, g20);
	defparam lut_212.LUT_SIZE = 2;
	defparam lut_212.mask = 4'b1011;

	lut_sub lut_220 ({g13, g11}, g21);
	defparam lut_220.LUT_SIZE = 2;
	defparam lut_220.mask = 4'b0001;

	lut_sub lut_224 ({i_11_, i_9_, i_10_, i_15_}, g22);
	defparam lut_224.LUT_SIZE = 4;
	defparam lut_224.mask = 16'h0100;

	lut_sub lut_230 ({g7, g22}, g23);
	defparam lut_230.LUT_SIZE = 2;
	defparam lut_230.mask = 4'b0001;

	lut_sub lut_238 ({g19, g20, g21, g23}, g24);
	defparam lut_238.LUT_SIZE = 4;
	defparam lut_238.mask = 16'h0800;

	lut_sub lut_246 ({g8, g10, g17, g24}, g25);
	defparam lut_246.LUT_SIZE = 4;
	defparam lut_246.mask = 16'h0010;

	lut_sub lut_252 ({g5, g25}, g26);
	defparam lut_252.LUT_SIZE = 2;
	defparam lut_252.mask = 4'b0100;

	lut_sub lut_256 ({i_8_, i_6_, i_7_}, g27);
	defparam lut_256.LUT_SIZE = 3;
	defparam lut_256.mask = 8'h20;

	lut_sub lut_264 ({g2, g4, g26, g27}, g28);
	defparam lut_264.LUT_SIZE = 4;
	defparam lut_264.mask = 16'h004f;

	lut_sub lut_272 ({i_1_, i_0_}, g29);
	defparam lut_272.LUT_SIZE = 2;
	defparam lut_272.mask = 4'b0100;

	lut_sub lut_276 ({i_6_, i_7_}, g30);
	defparam lut_276.LUT_SIZE = 2;
	defparam lut_276.mask = 4'b1000;

	lut_sub lut_281 ({i_8_, g30}, g31);
	defparam lut_281.LUT_SIZE = 2;
	defparam lut_281.mask = 4'b0100;

	lut_sub lut_287 ({g2, g31}, g32);
	defparam lut_287.LUT_SIZE = 2;
	defparam lut_287.mask = 4'b0001;

	lut_sub lut_295 ({g10, g23, g17, g5}, g33);
	defparam lut_295.LUT_SIZE = 4;
	defparam lut_295.mask = 16'h2000;

	lut_sub lut_299 ({i_6_, i_7_}, g34);
	defparam lut_299.LUT_SIZE = 2;
	defparam lut_299.mask = 4'b0100;

	lut_sub lut_308 ({g8, g2, g31, g19, g34}, g35);
	defparam lut_308.LUT_SIZE = 5;
	defparam lut_308.mask = 32'h005f0057;

	lut_sub lut_327 ({g32, g20, g21, g33, g35}, g36);
	defparam lut_327.LUT_SIZE = 5;
	defparam lut_327.mask = 32'haaaa0020;

	lut_sub lut_342 ({i_3_, i_4_, g28, g29, g36}, g37);
	defparam lut_342.LUT_SIZE = 5;
	defparam lut_342.mask = 32'h40505050;

	lut_sub lut_353 ({i_8_, g4}, g38);
	defparam lut_353.LUT_SIZE = 2;
	defparam lut_353.mask = 4'b0100;

	lut_sub lut_357 ({i_5_, i_3_, i_4_}, g39);
	defparam lut_357.LUT_SIZE = 3;
	defparam lut_357.mask = 8'h40;

	lut_sub lut_363 ({g1, g39}, g40);
	defparam lut_363.LUT_SIZE = 2;
	defparam lut_363.mask = 4'b0001;

	lut_sub lut_368 ({i_8_, i_7_, g40}, g41);
	defparam lut_368.LUT_SIZE = 3;
	defparam lut_368.mask = 8'h40;

	lut_sub lut_373 ({i_5_, i_3_, g1}, g42);
	defparam lut_373.LUT_SIZE = 3;
	defparam lut_373.mask = 8'h04;

	lut_sub lut_379 ({g7, g15}, g43);
	defparam lut_379.LUT_SIZE = 2;
	defparam lut_379.mask = 4'b0010;

	lut_sub lut_385 ({g18, g9}, g44);
	defparam lut_385.LUT_SIZE = 2;
	defparam lut_385.mask = 4'b0100;

	lut_sub lut_391 ({g6, i_15_, g13}, g45);
	defparam lut_391.LUT_SIZE = 3;
	defparam lut_391.mask = 8'h01;

	lut_sub lut_397 ({g6, i_15_, g9}, g46);
	defparam lut_397.LUT_SIZE = 3;
	defparam lut_397.mask = 8'h01;

	lut_sub lut_403 ({g18, g13}, g47);
	defparam lut_403.LUT_SIZE = 2;
	defparam lut_403.mask = 4'b0100;

	lut_sub lut_407 ({i_14_, i_12_, i_13_}, g48);
	defparam lut_407.LUT_SIZE = 3;
	defparam lut_407.mask = 8'hfb;

	lut_sub lut_418 ({i_11_, i_9_, i_10_, i_12_, g48}, g49);
	defparam lut_418.LUT_SIZE = 5;
	defparam lut_418.mask = 32'h0bb00ff0;

	lut_sub lut_440 ({g44, g45, g46, g47, g49}, g50);
	defparam lut_440.LUT_SIZE = 5;
	defparam lut_440.mask = 32'h80000000;

	lut_sub lut_449 ({g38, g41, g42, g43, g50}, g51);
	defparam lut_449.LUT_SIZE = 5;
	defparam lut_449.mask = 32'h00bb0bbb;

	lut_sub lut_467 ({i_5_, i_3_, i_4_}, g52);
	defparam lut_467.LUT_SIZE = 3;
	defparam lut_467.mask = 8'h08;

	lut_sub lut_471 ({i_11_, i_15_}, g53);
	defparam lut_471.LUT_SIZE = 2;
	defparam lut_471.mask = 4'b1000;

	lut_sub lut_477 ({i_9_, i_10_, g7, i_4_, g53}, g54);
	defparam lut_477.LUT_SIZE = 5;
	defparam lut_477.mask = 32'h04050500;

	lut_sub lut_485 ({i_5_, i_3_, i_8_, i_7_}, g55);
	defparam lut_485.LUT_SIZE = 4;
	defparam lut_485.mask = 16'h2000;

	lut_sub lut_492 ({i_0_, g52, g54, g55}, g56);
	defparam lut_492.LUT_SIZE = 4;
	defparam lut_492.mask = 16'h44f4;

	lut_sub lut_502 ({i_1_, i_0_, i_2_}, g57);
	defparam lut_502.LUT_SIZE = 3;
	defparam lut_502.mask = 8'h80;

	lut_sub lut_507 ({i_5_, i_3_, i_4_, g57}, g58);
	defparam lut_507.LUT_SIZE = 4;
	defparam lut_507.mask = 16'h4000;

	lut_sub lut_513 ({g58, g38}, g59);
	defparam lut_513.LUT_SIZE = 2;
	defparam lut_513.mask = 4'b0001;

	lut_sub lut_519 ({i_11_, i_12_, g59, g41}, g60);
	defparam lut_519.LUT_SIZE = 4;
	defparam lut_519.mask = 16'hc8cc;

	lut_sub lut_530 ({i_5_, i_3_, i_4_, g1}, g61);
	defparam lut_530.LUT_SIZE = 4;
	defparam lut_530.mask = 16'h0100;

	lut_sub lut_535 ({i_5_, i_3_, i_4_, g1}, g62);
	defparam lut_535.LUT_SIZE = 4;
	defparam lut_535.mask = 16'h0400;

	lut_sub lut_542 ({g31, g61, g62}, g63);
	defparam lut_542.LUT_SIZE = 3;
	defparam lut_542.mask = 8'h07;

	lut_sub lut_549 ({i_5_, i_3_, i_4_, g1}, g64);
	defparam lut_549.LUT_SIZE = 4;
	defparam lut_549.mask = 16'h0010;

	lut_sub lut_555 ({g1, g52}, g65);
	defparam lut_555.LUT_SIZE = 2;
	defparam lut_555.mask = 4'b0001;

	lut_sub lut_561 ({g6, i_15_, g7}, g66);
	defparam lut_561.LUT_SIZE = 3;
	defparam lut_561.mask = 8'h04;

	lut_sub lut_566 ({i_9_, i_10_, g66}, g67);
	defparam lut_566.LUT_SIZE = 3;
	defparam lut_566.mask = 8'h28;

	lut_sub lut_571 ({i_3_, i_1_, i_0_}, g68);
	defparam lut_571.LUT_SIZE = 3;
	defparam lut_571.mask = 8'hf7;

	lut_sub lut_584 ({i_8_, i_6_, g64, g65, g68}, g69);
	defparam lut_584.LUT_SIZE = 5;
	defparam lut_584.mask = 32'h55555540;

	lut_sub lut_602 ({i_11_, i_9_, i_10_, g59, g69}, g70);
	defparam lut_602.LUT_SIZE = 5;
	defparam lut_602.mask = 32'h55555545;

	lut_sub lut_625 ({g38, g64, g65, g67, g70}, g71);
	defparam lut_625.LUT_SIZE = 5;
	defparam lut_625.mask = 32'h55555111;

	lut_sub lut_644 ({i_9_, i_10_, g60, g63, g71}, g72);
	defparam lut_644.LUT_SIZE = 5;
	defparam lut_644.mask = 32'h44555504;

	lut_sub lut_661 ({i_1_, i_2_, g51, g56, g72}, g73);
	defparam lut_661.LUT_SIZE = 5;
	defparam lut_661.mask = 32'h50504050;

	lut_sub lut_674 ({g3, g37, g73}, o_0_);
	defparam lut_674.LUT_SIZE = 3;
	defparam lut_674.mask = 8'h45;

	lut_sub lut_682 ({g27, g40}, g75);
	defparam lut_682.LUT_SIZE = 2;
	defparam lut_682.mask = 4'b0001;

	lut_sub lut_691 ({g21, g23, g4, g27, g40}, g76);
	defparam lut_691.LUT_SIZE = 5;
	defparam lut_691.mask = 32'h05151515;

	lut_sub lut_706 ({i_5_, i_3_, i_4_, g29}, g77);
	defparam lut_706.LUT_SIZE = 4;
	defparam lut_706.mask = 16'h0010;

	lut_sub lut_712 ({g31, g40}, g78);
	defparam lut_712.LUT_SIZE = 2;
	defparam lut_712.mask = 4'b0001;

	lut_sub lut_720 ({g21, g10, g23, g12}, g79);
	defparam lut_720.LUT_SIZE = 4;
	defparam lut_720.mask = 16'h8000;

	lut_sub lut_727 ({i_8_, i_6_, i_7_, g19, g20, g40}, g80);
	defparam lut_727.LUT_SIZE = 6;
	defparam lut_727.mask = 64'h4555000000550000;

	lut_sub lut_746 ({g8, g14, g16, g78, g80}, g81);
	defparam lut_746.LUT_SIZE = 5;
	defparam lut_746.mask = 32'h88888a88;

	lut_sub lut_763 ({g29, g39, g78, g79, g81}, g82);
	defparam lut_763.LUT_SIZE = 5;
	defparam lut_763.mask = 32'h51515100;

	lut_sub lut_780 ({g17, g75, g76, g1544, g82}, g83);
	defparam lut_780.LUT_SIZE = 5;
	defparam lut_780.mask = 32'h10001010;

	lut_sub lut_790 ({i_8_, i_7_, g5, g40, g73, g83}, o_1_);
	defparam lut_790.LUT_SIZE = 6;
	defparam lut_790.mask = 64'h2223222223232222;

	lut_sub lut_813 ({g2, i_8_, i_6_, i_7_}, g85);
	defparam lut_813.LUT_SIZE = 4;
	defparam lut_813.mask = 16'h0002;

	lut_sub lut_822 ({g28, g52, g29, g73, g85}, o_2_);
	defparam lut_822.LUT_SIZE = 5;
	defparam lut_822.mask = 32'h11133333;

	lut_sub lut_840 ({g57, g39}, g87);
	defparam lut_840.LUT_SIZE = 2;
	defparam lut_840.mask = 4'b0001;

	lut_sub lut_846 ({g34, g87}, g88);
	defparam lut_846.LUT_SIZE = 2;
	defparam lut_846.mask = 4'b0001;

	lut_sub lut_851 ({i_8_, g88}, g89);
	defparam lut_851.LUT_SIZE = 2;
	defparam lut_851.mask = 4'b1011;

	lut_sub lut_859 ({g6, i_15_, g48}, g90);
	defparam lut_859.LUT_SIZE = 3;
	defparam lut_859.mask = 8'hf7;

	lut_sub lut_869 ({i_14_, i_12_, i_13_}, g91);
	defparam lut_869.LUT_SIZE = 3;
	defparam lut_869.mask = 8'hdf;

	lut_sub lut_881 ({g6, i_15_, g91}, g92);
	defparam lut_881.LUT_SIZE = 3;
	defparam lut_881.mask = 8'hfd;

	lut_sub lut_891 ({i_11_, i_9_, i_10_, i_15_}, g93);
	defparam lut_891.LUT_SIZE = 4;
	defparam lut_891.mask = 16'hffbf;

	lut_sub lut_911 ({g91, g93}, g94);
	defparam lut_911.LUT_SIZE = 2;
	defparam lut_911.mask = 4'b1000;

	lut_sub lut_915 ({i_11_, i_9_, i_10_, i_15_}, g95);
	defparam lut_915.LUT_SIZE = 4;
	defparam lut_915.mask = 16'h0080;

	lut_sub lut_921 ({g48, g95}, g96);
	defparam lut_921.LUT_SIZE = 2;
	defparam lut_921.mask = 4'b1011;

	lut_sub lut_930 ({g89, g94, g96}, g97);
	defparam lut_930.LUT_SIZE = 3;
	defparam lut_930.mask = 8'hb0;

	lut_sub lut_937 ({i_5_, i_3_, i_4_, g57}, g98);
	defparam lut_937.LUT_SIZE = 4;
	defparam lut_937.mask = 16'h0010;

	lut_sub lut_943 ({g38, g98}, g99);
	defparam lut_943.LUT_SIZE = 2;
	defparam lut_943.mask = 4'b0001;

	lut_sub lut_949 ({g4, g98}, g100);
	defparam lut_949.LUT_SIZE = 2;
	defparam lut_949.mask = 4'b0001;

	lut_sub lut_954 ({i_8_, g100}, g101);
	defparam lut_954.LUT_SIZE = 2;
	defparam lut_954.mask = 4'b0001;

	lut_sub lut_958 ({i_11_, i_9_, i_10_, i_15_}, g102);
	defparam lut_958.LUT_SIZE = 4;
	defparam lut_958.mask = 16'hffdf;

	lut_sub lut_978 ({g48, g102}, g103);
	defparam lut_978.LUT_SIZE = 2;
	defparam lut_978.mask = 4'b0111;

	lut_sub lut_984 ({i_11_, i_9_, i_10_, i_15_}, g104);
	defparam lut_984.LUT_SIZE = 4;
	defparam lut_984.mask = 16'h0002;

	lut_sub lut_990 ({g48, g104}, g105);
	defparam lut_990.LUT_SIZE = 2;
	defparam lut_990.mask = 4'b0100;

	lut_sub lut_999 ({g99, g101, g103, g90, g105}, g106);
	defparam lut_999.LUT_SIZE = 5;
	defparam lut_999.mask = 32'hff220a02;

	lut_sub lut_1020 ({g89, g90, g92, g97, g106}, g107);
	defparam lut_1020.LUT_SIZE = 5;
	defparam lut_1020.mask = 32'h00044444;

	lut_sub lut_1030 ({g34, g98}, g108);
	defparam lut_1030.LUT_SIZE = 2;
	defparam lut_1030.mask = 4'b0001;

	lut_sub lut_1035 ({i_8_, g108}, g109);
	defparam lut_1035.LUT_SIZE = 2;
	defparam lut_1035.mask = 4'b0100;

	lut_sub lut_1041 ({g52, g57}, g110);
	defparam lut_1041.LUT_SIZE = 2;
	defparam lut_1041.mask = 4'b0001;

	lut_sub lut_1046 ({i_8_, g30}, g111);
	defparam lut_1046.LUT_SIZE = 2;
	defparam lut_1046.mask = 4'b0001;

	lut_sub lut_1052 ({g110, g111}, g112);
	defparam lut_1052.LUT_SIZE = 2;
	defparam lut_1052.mask = 4'b0001;

	lut_sub lut_1056 ({i_9_, i_10_}, g113);
	defparam lut_1056.LUT_SIZE = 2;
	defparam lut_1056.mask = 4'b0001;

	lut_sub lut_1063 ({g53, g113, g48}, g114);
	defparam lut_1063.LUT_SIZE = 3;
	defparam lut_1063.mask = 8'h02;

	lut_sub lut_1067 ({i_11_, i_9_, i_10_, i_15_}, g115);
	defparam lut_1067.LUT_SIZE = 4;
	defparam lut_1067.mask = 16'hffef;

	lut_sub lut_1087 ({g91, g115}, g116);
	defparam lut_1087.LUT_SIZE = 2;
	defparam lut_1087.mask = 4'b1000;

	lut_sub lut_1093 ({g18, g91}, g117);
	defparam lut_1093.LUT_SIZE = 2;
	defparam lut_1093.mask = 4'b1000;

	lut_sub lut_1099 ({g31, g110}, g118);
	defparam lut_1099.LUT_SIZE = 2;
	defparam lut_1099.mask = 4'b0001;

	lut_sub lut_1103 ({i_11_, i_9_, i_10_, i_15_}, g119);
	defparam lut_1103.LUT_SIZE = 4;
	defparam lut_1103.mask = 16'h0008;

	lut_sub lut_1109 ({g48, g119}, g120);
	defparam lut_1109.LUT_SIZE = 2;
	defparam lut_1109.mask = 4'b1011;

	lut_sub lut_1118 ({g118, g120, g90}, g121);
	defparam lut_1118.LUT_SIZE = 3;
	defparam lut_1118.mask = 8'h0e;

	lut_sub lut_1124 ({i_11_, i_9_, i_10_, i_15_}, g122);
	defparam lut_1124.LUT_SIZE = 4;
	defparam lut_1124.mask = 16'hfffb;

	lut_sub lut_1144 ({g91, g122}, g123);
	defparam lut_1144.LUT_SIZE = 2;
	defparam lut_1144.mask = 4'b1000;

	lut_sub lut_1148 ({i_11_, i_9_, i_10_, i_15_}, g124);
	defparam lut_1148.LUT_SIZE = 4;
	defparam lut_1148.mask = 16'h0001;

	lut_sub lut_1154 ({g91, g124}, g125);
	defparam lut_1154.LUT_SIZE = 2;
	defparam lut_1154.mask = 4'b0100;

	lut_sub lut_1162 ({g118, g112, g123, g125}, g126);
	defparam lut_1162.LUT_SIZE = 4;
	defparam lut_1162.mask = 16'hf8a8;

	lut_sub lut_1175 ({g22, g91}, g127);
	defparam lut_1175.LUT_SIZE = 2;
	defparam lut_1175.mask = 4'b1101;

	lut_sub lut_1184 ({g88, g127, g125}, g128);
	defparam lut_1184.LUT_SIZE = 3;
	defparam lut_1184.mask = 8'h0d;

	lut_sub lut_1196 ({g89, g116, g117, g121, g126, g128}, g129);
	defparam lut_1196.LUT_SIZE = 6;
	defparam lut_1196.mask = 64'h2000000020202020;

	lut_sub lut_1210 ({g99, g101, g109, g112, g114, g129}, g130);
	defparam lut_1210.LUT_SIZE = 6;
	defparam lut_1210.mask = 64'h5444444444444444;

	lut_sub lut_1232 ({g53, g5}, g131);
	defparam lut_1232.LUT_SIZE = 2;
	defparam lut_1232.mask = 4'b0001;

	lut_sub lut_1238 ({g48, g131}, g132);
	defparam lut_1238.LUT_SIZE = 2;
	defparam lut_1238.mask = 4'b1011;

	lut_sub lut_1246 ({i_11_, i_9_, i_10_, i_15_, g91, g109}, g133);
	defparam lut_1246.LUT_SIZE = 6;
	defparam lut_1246.mask = 64'hfbfffbfbfbfbfbff;

	lut_sub lut_1309 ({g27, g58}, g134);
	defparam lut_1309.LUT_SIZE = 2;
	defparam lut_1309.mask = 4'b0001;

	lut_sub lut_1314 ({i_6_, i_7_, g58}, g135);
	defparam lut_1314.LUT_SIZE = 3;
	defparam lut_1314.mask = 8'h04;

	lut_sub lut_1319 ({i_8_, g135}, g136);
	defparam lut_1319.LUT_SIZE = 2;
	defparam lut_1319.mask = 4'b0001;

	lut_sub lut_1329 ({g134, g136, g120, g103, g116, g123}, g137);
	defparam lut_1329.LUT_SIZE = 6;
	defparam lut_1329.mask = 64'hffff000caaaa0008;

	lut_sub lut_1363 ({g118, g94, g92, g116}, g138);
	defparam lut_1363.LUT_SIZE = 4;
	defparam lut_1363.mask = 16'h00df;

	lut_sub lut_1377 ({g134, g103, g96, g105}, g139);
	defparam lut_1377.LUT_SIZE = 4;
	defparam lut_1377.mask = 16'h00fd;

	lut_sub lut_1391 ({g134, g94, g116, g125}, g140);
	defparam lut_1391.LUT_SIZE = 4;
	defparam lut_1391.mask = 16'h007f;

	lut_sub lut_1401 ({i_9_, i_10_}, g141);
	defparam lut_1401.LUT_SIZE = 2;
	defparam lut_1401.mask = 4'b0100;

	lut_sub lut_1407 ({i_11_, i_15_, g141, g48}, g142);
	defparam lut_1407.LUT_SIZE = 4;
	defparam lut_1407.mask = 16'h2000;

	lut_sub lut_1416 ({g59, g134, g99, g142, g90}, g143);
	defparam lut_1416.LUT_SIZE = 5;
	defparam lut_1416.mask = 32'hf5444444;

	lut_sub lut_1435 ({g138, g139, g140, g143}, g144);
	defparam lut_1435.LUT_SIZE = 4;
	defparam lut_1435.mask = 16'h4000;

	lut_sub lut_1440 ({i_8_, g108}, g145);
	defparam lut_1440.LUT_SIZE = 2;
	defparam lut_1440.mask = 4'b0001;

	lut_sub lut_1446 ({i_8_, g88, g112}, g146);
	defparam lut_1446.LUT_SIZE = 3;
	defparam lut_1446.mask = 8'ha8;

	lut_sub lut_1458 ({g145, g146, g127, g125, g114, g105}, g147);
	defparam lut_1458.LUT_SIZE = 6;
	defparam lut_1458.mask = 64'haaaaffff00800080;

	lut_sub lut_1493 ({g118, g127, g117, g137, g144, g147}, g148);
	defparam lut_1493.LUT_SIZE = 6;
	defparam lut_1493.mask = 64'h0101010100000100;

	lut_sub lut_1503 ({g27, g98}, g149);
	defparam lut_1503.LUT_SIZE = 2;
	defparam lut_1503.mask = 4'b0001;

	lut_sub lut_1510 ({g149, g127, g114}, g150);
	defparam lut_1510.LUT_SIZE = 3;
	defparam lut_1510.mask = 8'h0d;

	lut_sub lut_1517 ({i_8_, g88}, g151);
	defparam lut_1517.LUT_SIZE = 2;
	defparam lut_1517.mask = 4'b0001;

	lut_sub lut_1524 ({g99, g142, g117}, g152);
	defparam lut_1524.LUT_SIZE = 3;
	defparam lut_1524.mask = 8'h07;

	lut_sub lut_1533 ({g134, g127, g114}, g153);
	defparam lut_1533.LUT_SIZE = 3;
	defparam lut_1533.mask = 8'h0d;

	lut_sub lut_1544 ({g136, g151, g114, g152, g153}, g154);
	defparam lut_1544.LUT_SIZE = 5;
	defparam lut_1544.mask = 32'h88808080;

	lut_sub lut_1556 ({i_8_, g100, g108, g142, g117}, g155);
	defparam lut_1556.LUT_SIZE = 5;
	defparam lut_1556.mask = 32'h07070033;

	lut_sub lut_1574 ({g109, g136, g125, g105, g155}, g156);
	defparam lut_1574.LUT_SIZE = 5;
	defparam lut_1574.mask = 32'haa888080;

	lut_sub lut_1590 ({g136, g125, g150, g154, g156}, g157);
	defparam lut_1590.LUT_SIZE = 5;
	defparam lut_1590.mask = 32'h10101000;

	lut_sub lut_1596 ({i_11_, i_9_, i_10_, i_15_}, g158);
	defparam lut_1596.LUT_SIZE = 4;
	defparam lut_1596.mask = 16'h4000;

	lut_sub lut_1602 ({g91, g158}, g159);
	defparam lut_1602.LUT_SIZE = 2;
	defparam lut_1602.mask = 4'b0100;

	lut_sub lut_1612 ({g134, g118, g145, g151, g159, g96}, g160);
	defparam lut_1612.LUT_SIZE = 6;
	defparam lut_1612.mask = 64'hf5c45544c4c44444;

	lut_sub lut_1643 ({i_8_, g135, g92, g123}, g161);
	defparam lut_1643.LUT_SIZE = 4;
	defparam lut_1643.mask = 16'h0c0d;

	lut_sub lut_1652 ({i_11_, i_9_, i_10_, i_15_, g48}, g162);
	defparam lut_1652.LUT_SIZE = 5;
	defparam lut_1652.mask = 32'h80000080;

	lut_sub lut_1660 ({i_8_, g88, g108, g90}, g163);
	defparam lut_1660.LUT_SIZE = 4;
	defparam lut_1660.mask = 16'h222a;

	lut_sub lut_1669 ({i_15_, g141}, g164);
	defparam lut_1669.LUT_SIZE = 2;
	defparam lut_1669.mask = 4'b0001;

	lut_sub lut_1675 ({g91, g164}, g165);
	defparam lut_1675.LUT_SIZE = 2;
	defparam lut_1675.mask = 4'b0100;

	lut_sub lut_1683 ({g100, g112, g127, g165}, g166);
	defparam lut_1683.LUT_SIZE = 4;
	defparam lut_1683.mask = 16'hf232;

	lut_sub lut_1699 ({g134, g117, g162, g163, g166}, g167);
	defparam lut_1699.LUT_SIZE = 5;
	defparam lut_1699.mask = 32'h44444000;

	lut_sub lut_1711 ({g160, g1775, g161, g167}, g168);
	defparam lut_1711.LUT_SIZE = 4;
	defparam lut_1711.mask = 16'h0004;

	lut_sub lut_1721 ({g107, g130, g1782, g148, g157, g168}, g169);
	defparam lut_1721.LUT_SIZE = 6;
	defparam lut_1721.mask = 64'h0000000000000001;

	lut_sub lut_1727 ({i_14_, i_12_, i_13_, g102, g119}, g170);
	defparam lut_1727.LUT_SIZE = 5;
	defparam lut_1727.mask = 32'h0000dd05;

	lut_sub lut_1738 ({i_14_, i_12_, i_13_}, g171);
	defparam lut_1738.LUT_SIZE = 3;
	defparam lut_1738.mask = 8'hfe;

	lut_sub lut_1750 ({g15, g171}, g172);
	defparam lut_1750.LUT_SIZE = 2;
	defparam lut_1750.mask = 4'b1000;

	lut_sub lut_1756 ({g102, g171}, g173);
	defparam lut_1756.LUT_SIZE = 2;
	defparam lut_1756.mask = 4'b1000;

	lut_sub lut_1764 ({g20, g172, g142, g173}, g174);
	defparam lut_1764.LUT_SIZE = 4;
	defparam lut_1764.mask = 16'h0080;

	lut_sub lut_1770 ({i_14_, i_12_, i_13_, g119, g131}, g175);
	defparam lut_1770.LUT_SIZE = 5;
	defparam lut_1770.mask = 32'h00007707;

	lut_sub lut_1786 ({i_8_, g88, g170, g174, g175}, g176);
	defparam lut_1786.LUT_SIZE = 5;
	defparam lut_1786.mask = 32'h005500cf;

	lut_sub lut_1801 ({g11, g171}, g177);
	defparam lut_1801.LUT_SIZE = 2;
	defparam lut_1801.mask = 4'b0010;

	lut_sub lut_1805 ({i_11_, i_9_, i_10_}, g178);
	defparam lut_1805.LUT_SIZE = 3;
	defparam lut_1805.mask = 8'h28;

	lut_sub lut_1812 ({i_15_, g171, g178}, g179);
	defparam lut_1812.LUT_SIZE = 3;
	defparam lut_1812.mask = 8'h40;

	lut_sub lut_1818 ({i_14_, i_12_, i_13_, g59, g95}, g180);
	defparam lut_1818.LUT_SIZE = 5;
	defparam lut_1818.mask = 32'h00001101;

	lut_sub lut_1826 ({g91, g119}, g181);
	defparam lut_1826.LUT_SIZE = 2;
	defparam lut_1826.mask = 4'b0100;

	lut_sub lut_1830 ({i_14_, i_12_, i_13_}, g182);
	defparam lut_1830.LUT_SIZE = 3;
	defparam lut_1830.mask = 8'h02;

	lut_sub lut_1836 ({g119, g182}, g183);
	defparam lut_1836.LUT_SIZE = 2;
	defparam lut_1836.mask = 4'b0001;

	lut_sub lut_1844 ({g181, g118, g112, g183}, g184);
	defparam lut_1844.LUT_SIZE = 4;
	defparam lut_1844.mask = 16'h0537;

	lut_sub lut_1856 ({g104, g91}, g185);
	defparam lut_1856.LUT_SIZE = 2;
	defparam lut_1856.mask = 4'b1101;

	lut_sub lut_1865 ({g31, g34, g87}, g186);
	defparam lut_1865.LUT_SIZE = 3;
	defparam lut_1865.mask = 8'h15;

	lut_sub lut_1873 ({g104, g182}, g187);
	defparam lut_1873.LUT_SIZE = 2;
	defparam lut_1873.mask = 4'b0001;

	lut_sub lut_1882 ({g134, g118, g185, g186, g187}, g188);
	defparam lut_1882.LUT_SIZE = 5;
	defparam lut_1882.mask = 32'heeaa0e0a;

	lut_sub lut_1906 ({g151, g177, g179, g180, g184, g188}, g189);
	defparam lut_1906.LUT_SIZE = 6;
	defparam lut_1906.mask = 64'h4040404040000000;

	lut_sub lut_1916 ({i_14_, g99, g131}, g190);
	defparam lut_1916.LUT_SIZE = 3;
	defparam lut_1916.mask = 8'h01;

	lut_sub lut_1922 ({g15, g182}, g191);
	defparam lut_1922.LUT_SIZE = 2;
	defparam lut_1922.mask = 4'b0100;

	lut_sub lut_1929 ({i_8_, i_6_, i_7_, g58, g98, g191}, g192);
	defparam lut_1929.LUT_SIZE = 6;
	defparam lut_1929.mask = 64'h0011111500110000;

	lut_sub lut_1943 ({g102, g182}, g193);
	defparam lut_1943.LUT_SIZE = 2;
	defparam lut_1943.mask = 4'b0100;

	lut_sub lut_1950 ({i_8_, g108, g183, g193}, g194);
	defparam lut_1950.LUT_SIZE = 4;
	defparam lut_1950.mask = 16'h0507;

	lut_sub lut_1960 ({g104, g171}, g195);
	defparam lut_1960.LUT_SIZE = 2;
	defparam lut_1960.mask = 4'b0010;

	lut_sub lut_1968 ({i_8_, g108, g185, g195, g187}, g196);
	defparam lut_1968.LUT_SIZE = 5;
	defparam lut_1968.mask = 32'h00f70033;

	lut_sub lut_1984 ({g6, i_15_, g171}, g197);
	defparam lut_1984.LUT_SIZE = 3;
	defparam lut_1984.mask = 8'h08;

	lut_sub lut_1991 ({i_8_, g108, g197, g177}, g198);
	defparam lut_1991.LUT_SIZE = 4;
	defparam lut_1991.mask = 16'h0507;

	lut_sub lut_2001 ({g119, g171}, g199);
	defparam lut_2001.LUT_SIZE = 2;
	defparam lut_2001.mask = 4'b0010;

	lut_sub lut_2008 ({i_8_, g181, g135, g199}, g200);
	defparam lut_2008.LUT_SIZE = 4;
	defparam lut_2008.mask = 16'h0013;

	lut_sub lut_2016 ({g11, g182}, g201);
	defparam lut_2016.LUT_SIZE = 2;
	defparam lut_2016.mask = 4'b1110;

	lut_sub lut_2024 ({i_8_, i_6_, i_7_, g98, g201}, g202);
	defparam lut_2024.LUT_SIZE = 5;
	defparam lut_2024.mask = 32'h00220200;

	lut_sub lut_2032 ({g182, g93}, g203);
	defparam lut_2032.LUT_SIZE = 2;
	defparam lut_2032.mask = 4'b0010;

	lut_sub lut_2038 ({g182, g158}, g204);
	defparam lut_2038.LUT_SIZE = 2;
	defparam lut_2038.mask = 4'b1110;

	lut_sub lut_2047 ({i_8_, g100, g203, g204}, g205);
	defparam lut_2047.LUT_SIZE = 4;
	defparam lut_2047.mask = 16'h000b;

	lut_sub lut_2055 ({g11, g91}, g206);
	defparam lut_2055.LUT_SIZE = 2;
	defparam lut_2055.mask = 4'b1101;

	lut_sub lut_2063 ({g91, g131}, g207);
	defparam lut_2063.LUT_SIZE = 2;
	defparam lut_2063.mask = 4'b0100;

	lut_sub lut_2071 ({i_8_, g4, g206, g98, g207}, g208);
	defparam lut_2071.LUT_SIZE = 5;
	defparam lut_2071.mask = 32'h00300031;

	lut_sub lut_2081 ({g6, i_15_, g182}, g209);
	defparam lut_2081.LUT_SIZE = 3;
	defparam lut_2081.mask = 8'h04;

	lut_sub lut_2088 ({i_8_, g100, g183, g209}, g210);
	defparam lut_2088.LUT_SIZE = 4;
	defparam lut_2088.mask = 16'h0007;

	lut_sub lut_2100 ({g198, g200, g202, g205, g208, g210}, g211);
	defparam lut_2100.LUT_SIZE = 6;
	defparam lut_2100.mask = 64'h8000000000000000;

	lut_sub lut_2108 ({i_8_, g59, g108, g112, g135}, g212);
	defparam lut_2108.LUT_SIZE = 5;
	defparam lut_2108.mask = 32'h80008800;

	lut_sub lut_2116 ({g95, g182}, g213);
	defparam lut_2116.LUT_SIZE = 2;
	defparam lut_2116.mask = 4'b0001;

	lut_sub lut_2121 ({i_8_, i_6_, g87}, g214);
	defparam lut_2121.LUT_SIZE = 3;
	defparam lut_2121.mask = 8'h40;

	lut_sub lut_2127 ({g118, g214}, g215);
	defparam lut_2127.LUT_SIZE = 2;
	defparam lut_2127.mask = 4'b1000;

	lut_sub lut_2133 ({g13, g119}, g216);
	defparam lut_2133.LUT_SIZE = 2;
	defparam lut_2133.mask = 4'b0001;

	lut_sub lut_2141 ({g112, g216, g199, g120}, g217);
	defparam lut_2141.LUT_SIZE = 4;
	defparam lut_2141.mask = 16'h00bf;

	lut_sub lut_2155 ({g212, g213, g215, g217}, g218);
	defparam lut_2155.LUT_SIZE = 4;
	defparam lut_2155.mask = 16'ha0a2;

	lut_sub lut_2167 ({g134, g183, g187, g193}, g219);
	defparam lut_2167.LUT_SIZE = 4;
	defparam lut_2167.mask = 16'h007f;

	lut_sub lut_2179 ({g91, g102}, g220);
	defparam lut_2179.LUT_SIZE = 2;
	defparam lut_2179.mask = 4'b1000;

	lut_sub lut_2185 ({g6, i_15_, g91}, g221);
	defparam lut_2185.LUT_SIZE = 3;
	defparam lut_2185.mask = 8'hf7;

	lut_sub lut_2197 ({g15, g91}, g222);
	defparam lut_2197.LUT_SIZE = 2;
	defparam lut_2197.mask = 4'b1000;

	lut_sub lut_2205 ({g99, g220, g221, g222}, g223);
	defparam lut_2205.LUT_SIZE = 4;
	defparam lut_2205.mask = 16'h00df;

	lut_sub lut_2217 ({g6, i_15_, g182}, g224);
	defparam lut_2217.LUT_SIZE = 3;
	defparam lut_2217.mask = 8'h01;

	lut_sub lut_2225 ({g99, g183, g224, g213}, g225);
	defparam lut_2225.LUT_SIZE = 4;
	defparam lut_2225.mask = 16'h007f;

	lut_sub lut_2237 ({g22, g182}, g226);
	defparam lut_2237.LUT_SIZE = 2;
	defparam lut_2237.mask = 4'b1110;

	lut_sub lut_2245 ({g38, g87}, g227);
	defparam lut_2245.LUT_SIZE = 2;
	defparam lut_2245.mask = 4'b0001;

	lut_sub lut_2249 ({i_11_, i_9_, i_10_, i_15_}, g228);
	defparam lut_2249.LUT_SIZE = 4;
	defparam lut_2249.mask = 16'h0140;

	lut_sub lut_2258 ({i_3_, i_4_, g57, g38, g182, g228}, g229);
	defparam lut_2258.LUT_SIZE = 6;
	defparam lut_2258.mask = 64'h0000000100000000;

	lut_sub lut_2267 ({g99, g226, g203, g227, g229}, g230);
	defparam lut_2267.LUT_SIZE = 5;
	defparam lut_2267.mask = 32'h15001515;

	lut_sub lut_2281 ({g182, g124}, g231);
	defparam lut_2281.LUT_SIZE = 2;
	defparam lut_2281.mask = 4'b1110;

	lut_sub lut_2289 ({g182, g115}, g232);
	defparam lut_2289.LUT_SIZE = 2;
	defparam lut_2289.mask = 4'b0010;

	lut_sub lut_2297 ({g99, g193, g231, g232}, g233);
	defparam lut_2297.LUT_SIZE = 4;
	defparam lut_2297.mask = 16'h00df;

	lut_sub lut_2312 ({g219, g223, g225, g230, g233}, g234);
	defparam lut_2312.LUT_SIZE = 5;
	defparam lut_2312.mask = 32'h80000000;

	lut_sub lut_2322 ({g176, g189, g1543, g211, g218, g234}, g235);
	defparam lut_2322.LUT_SIZE = 6;
	defparam lut_2322.mask = 64'h0000000100000000;

	lut_sub lut_2328 ({i_8_, g34, g110}, g236);
	defparam lut_2328.LUT_SIZE = 3;
	defparam lut_2328.mask = 8'h10;

	lut_sub lut_2334 ({g6, g236}, g237);
	defparam lut_2334.LUT_SIZE = 2;
	defparam lut_2334.mask = 4'b0001;

	lut_sub lut_2340 ({g31, g98}, g238);
	defparam lut_2340.LUT_SIZE = 2;
	defparam lut_2340.mask = 4'b0001;

	lut_sub lut_2346 ({g227, g224}, g239);
	defparam lut_2346.LUT_SIZE = 2;
	defparam lut_2346.mask = 4'b0001;

	lut_sub lut_2353 ({g99, g187, g209}, g240);
	defparam lut_2353.LUT_SIZE = 3;
	defparam lut_2353.mask = 8'h07;

	lut_sub lut_2362 ({i_8_, g108, g183, g201}, g241);
	defparam lut_2362.LUT_SIZE = 4;
	defparam lut_2362.mask = 16'h0b00;

	lut_sub lut_2374 ({g14, g237, g238, g239, g240, g241}, g242);
	defparam lut_2374.LUT_SIZE = 6;
	defparam lut_2374.mask = 64'h8080000080000000;

	lut_sub lut_2382 ({g30, g87}, g243);
	defparam lut_2382.LUT_SIZE = 2;
	defparam lut_2382.mask = 4'b0001;

	lut_sub lut_2387 ({i_15_, g91}, g244);
	defparam lut_2387.LUT_SIZE = 2;
	defparam lut_2387.mask = 4'b1000;

	lut_sub lut_2392 ({i_11_, i_9_, i_10_, g244}, g245);
	defparam lut_2392.LUT_SIZE = 4;
	defparam lut_2392.mask = 16'h0104;

	lut_sub lut_2398 ({i_14_, i_12_, i_13_, g131}, g246);
	defparam lut_2398.LUT_SIZE = 4;
	defparam lut_2398.mask = 16'h0051;

	lut_sub lut_2408 ({g221, g183, g199, g197}, g247);
	defparam lut_2408.LUT_SIZE = 4;
	defparam lut_2408.mask = 16'h0080;

	lut_sub lut_2417 ({g245, g185, g246, g120, g247}, g248);
	defparam lut_2417.LUT_SIZE = 5;
	defparam lut_2417.mask = 32'h00100000;

	lut_sub lut_2423 ({i_14_, i_12_, i_13_, g100, g108}, g249);
	defparam lut_2423.LUT_SIZE = 5;
	defparam lut_2423.mask = 32'h00300005;

	lut_sub lut_2434 ({g119, g243, g248, g249}, g250);
	defparam lut_2434.LUT_SIZE = 4;
	defparam lut_2434.mask = 16'h0c5d;

	lut_sub lut_2447 ({i_8_, g88, g118, g243}, g251);
	defparam lut_2447.LUT_SIZE = 4;
	defparam lut_2447.mask = 16'h7f77;

	lut_sub lut_2464 ({i_11_, i_9_, i_10_, i_15_, g171}, g252);
	defparam lut_2464.LUT_SIZE = 5;
	defparam lut_2464.mask = 32'h00008008;

	lut_sub lut_2471 ({g131, g182}, g253);
	defparam lut_2471.LUT_SIZE = 2;
	defparam lut_2471.mask = 4'b0001;

	lut_sub lut_2477 ({i_15_, g141, g171}, g254);
	defparam lut_2477.LUT_SIZE = 3;
	defparam lut_2477.mask = 8'h20;

	lut_sub lut_2483 ({g141, g244}, g255);
	defparam lut_2483.LUT_SIZE = 2;
	defparam lut_2483.mask = 4'b0001;

	lut_sub lut_2492 ({g193, g177, g253, g254, g255}, g256);
	defparam lut_2492.LUT_SIZE = 5;
	defparam lut_2492.mask = 32'h80000000;

	lut_sub lut_2497 ({g6, i_15_, i_14_, i_12_}, g257);
	defparam lut_2497.LUT_SIZE = 4;
	defparam lut_2497.mask = 16'h0010;

	lut_sub lut_2506 ({g212, g251, g252, g256, g257}, g258);
	defparam lut_2506.LUT_SIZE = 5;
	defparam lut_2506.mask = 32'haa20ff30;

	lut_sub lut_2526 ({g207, g204}, g259);
	defparam lut_2526.LUT_SIZE = 2;
	defparam lut_2526.mask = 4'b0100;

	lut_sub lut_2532 ({i_11_, g113, g236}, g260);
	defparam lut_2532.LUT_SIZE = 3;
	defparam lut_2532.mask = 8'h10;

	lut_sub lut_2538 ({i_8_, g88, g231}, g261);
	defparam lut_2538.LUT_SIZE = 3;
	defparam lut_2538.mask = 8'h02;

	lut_sub lut_2546 ({i_8_, g30, g20, g21, g98}, g262);
	defparam lut_2546.LUT_SIZE = 5;
	defparam lut_2546.mask = 32'h00110050;

	lut_sub lut_2559 ({g99, g251, g259, g260, g261, g262}, g263);
	defparam lut_2559.LUT_SIZE = 6;
	defparam lut_2559.mask = 64'h8080008000800080;

	lut_sub lut_2569 ({g13, g102}, g264);
	defparam lut_2569.LUT_SIZE = 2;
	defparam lut_2569.mask = 4'b0010;

	lut_sub lut_2577 ({g185, g216, g120, g173}, g265);
	defparam lut_2577.LUT_SIZE = 4;
	defparam lut_2577.mask = 16'h0020;

	lut_sub lut_2585 ({i_8_, g4, g98, g221, g185}, g266);
	defparam lut_2585.LUT_SIZE = 5;
	defparam lut_2585.mask = 32'h000a000c;

	lut_sub lut_2598 ({g264, g101, g199, g265, g103, g266}, g267);
	defparam lut_2598.LUT_SIZE = 6;
	defparam lut_2598.mask = 64'haaaa0200aaaa0000;

	lut_sub lut_2620 ({g95, g171}, g268);
	defparam lut_2620.LUT_SIZE = 2;
	defparam lut_2620.mask = 4'b0010;

	lut_sub lut_2625 ({i_14_, i_12_, i_13_, g102}, g269);
	defparam lut_2625.LUT_SIZE = 4;
	defparam lut_2625.mask = 16'h00a2;

	lut_sub lut_2633 ({g91, g95}, g270);
	defparam lut_2633.LUT_SIZE = 2;
	defparam lut_2633.mask = 4'b1011;

	lut_sub lut_2643 ({i_8_, g4, g98, g270, g255}, g271);
	defparam lut_2643.LUT_SIZE = 5;
	defparam lut_2643.mask = 32'h000c000d;

	lut_sub lut_2656 ({g134, g118, g201, g209, g246}, g272);
	defparam lut_2656.LUT_SIZE = 5;
	defparam lut_2656.mask = 32'hff080f08;

	lut_sub lut_2679 ({g145, g268, g172, g269, g271, g272}, g273);
	defparam lut_2679.LUT_SIZE = 6;
	defparam lut_2679.mask = 64'h4444444440000000;

	lut_sub lut_2697 ({g242, g250, g258, g263, g267, g273}, g274);
	defparam lut_2697.LUT_SIZE = 6;
	defparam lut_2697.mask = 64'h0000000000010000;

	lut_sub lut_2703 ({g235, g274}, g275);
	defparam lut_2703.LUT_SIZE = 2;
	defparam lut_2703.mask = 4'b0001;

	lut_sub lut_2711 ({g17, g75, g76, g1544}, g276);
	defparam lut_2711.LUT_SIZE = 4;
	defparam lut_2711.mask = 16'h4044;

	lut_sub lut_2719 ({g134, g118}, g277);
	defparam lut_2719.LUT_SIZE = 2;
	defparam lut_2719.mask = 4'b1000;

	lut_sub lut_2726 ({g191, g277, g214}, g278);
	defparam lut_2726.LUT_SIZE = 3;
	defparam lut_2726.mask = 8'h0d;

	lut_sub lut_2734 ({g131, g171}, g279);
	defparam lut_2734.LUT_SIZE = 2;
	defparam lut_2734.mask = 4'b0010;

	lut_sub lut_2740 ({i_9_, g53, g182}, g280);
	defparam lut_2740.LUT_SIZE = 3;
	defparam lut_2740.mask = 8'h01;

	lut_sub lut_2748 ({g142, g103, g114, g105}, g281);
	defparam lut_2748.LUT_SIZE = 4;
	defparam lut_2748.mask = 16'h0800;

	lut_sub lut_2757 ({i_8_, g88, g118, g216, g243, g281}, g282);
	defparam lut_2757.LUT_SIZE = 6;
	defparam lut_2757.mask = 64'hdd505550dd50dd50;

	lut_sub lut_2795 ({g145, g279, g214, g280, g282}, g283);
	defparam lut_2795.LUT_SIZE = 5;
	defparam lut_2795.mask = 32'h54545400;

	lut_sub lut_2809 ({i_8_, g4, g58}, g284);
	defparam lut_2809.LUT_SIZE = 3;
	defparam lut_2809.mask = 8'h01;

	lut_sub lut_2815 ({i_8_, g134, g108}, g285);
	defparam lut_2815.LUT_SIZE = 3;
	defparam lut_2815.mask = 8'h8c;

	lut_sub lut_2827 ({g100, g251, g253, g284, g159, g285}, g286);
	defparam lut_2827.LUT_SIZE = 6;
	defparam lut_2827.mask = 64'hfc54cc44cc44cc44;

	lut_sub lut_2860 ({g99, g94, g116}, g287);
	defparam lut_2860.LUT_SIZE = 3;
	defparam lut_2860.mask = 8'h07;

	lut_sub lut_2868 ({i_8_, i_6_, i_7_, g5, g40}, g288);
	defparam lut_2868.LUT_SIZE = 5;
	defparam lut_2868.mask = 32'h00100050;

	lut_sub lut_2876 ({i_11_, i_9_, i_10_, i_15_, g91, g100}, g289);
	defparam lut_2876.LUT_SIZE = 6;
	defparam lut_2876.mask = 64'h0000000000000c04;

	lut_sub lut_2886 ({i_8_, g4, g98, g92, g165}, g290);
	defparam lut_2886.LUT_SIZE = 5;
	defparam lut_2886.mask = 32'h000c000d;

	lut_sub lut_2900 ({g100, g251, g287, g288, g289, g290}, g291);
	defparam lut_2900.LUT_SIZE = 6;
	defparam lut_2900.mask = 64'ha000800080008000;

	lut_sub lut_2912 ({g127, g90, g116, g125}, g292);
	defparam lut_2912.LUT_SIZE = 4;
	defparam lut_2912.mask = 16'h0008;

	lut_sub lut_2920 ({i_8_, g48, g91, g95, g216}, g293);
	defparam lut_2920.LUT_SIZE = 5;
	defparam lut_2920.mask = 32'h888aaaaa;

	lut_sub lut_2937 ({i_11_, i_9_, i_10_, i_15_, g91}, g294);
	defparam lut_2937.LUT_SIZE = 5;
	defparam lut_2937.mask = 32'h02202000;

	lut_sub lut_2948 ({g59, g243, g292, g293, g294}, g295);
	defparam lut_2948.LUT_SIZE = 5;
	defparam lut_2948.mask = 32'hff02aa02;

	lut_sub lut_2971 ({g134, g252, g283, g286, g291, g295}, g296);
	defparam lut_2971.LUT_SIZE = 6;
	defparam lut_2971.mask = 64'h0001000100010000;

	lut_sub lut_2979 ({g13, g104}, g297);
	defparam lut_2979.LUT_SIZE = 2;
	defparam lut_2979.mask = 4'b0001;

	lut_sub lut_2985 ({i_11_, i_9_, i_10_, g59, g244}, g298);
	defparam lut_2985.LUT_SIZE = 5;
	defparam lut_2985.mask = 32'h01001000;

	lut_sub lut_2994 ({i_8_, g20, g4, g98, g216}, g299);
	defparam lut_2994.LUT_SIZE = 5;
	defparam lut_2994.mask = 32'h01010300;

	lut_sub lut_3006 ({g14, g4, g98, g118, g299}, g300);
	defparam lut_3006.LUT_SIZE = 5;
	defparam lut_3006.mask = 32'haaaa8880;

	lut_sub lut_3026 ({g297, g89, g245, g136, g298, g300}, g301);
	defparam lut_3026.LUT_SIZE = 6;
	defparam lut_3026.mask = 64'h4400444440004040;

	lut_sub lut_3041 ({i_8_, g220, g264, g135}, g302);
	defparam lut_3041.LUT_SIZE = 4;
	defparam lut_3041.mask = 16'h0015;

	lut_sub lut_3050 ({i_8_, g297, g264, g108}, g303);
	defparam lut_3050.LUT_SIZE = 4;
	defparam lut_3050.mask = 16'h1505;

	lut_sub lut_3060 ({g13, g95}, g304);
	defparam lut_3060.LUT_SIZE = 2;
	defparam lut_3060.mask = 4'b0001;

	lut_sub lut_3069 ({i_8_, g59, g221, g88, g304, g270}, g305);
	defparam lut_3069.LUT_SIZE = 6;
	defparam lut_3069.mask = 64'h0f0bff0b0000ff00;

	lut_sub lut_3103 ({g89, g185, g302, g303, g305}, g306);
	defparam lut_3103.LUT_SIZE = 5;
	defparam lut_3103.mask = 32'h00808080;

	lut_sub lut_3113 ({g206, g118, g112, g185}, g307);
	defparam lut_3113.LUT_SIZE = 4;
	defparam lut_3113.mask = 16'hc0d5;

	lut_sub lut_3126 ({g21, g149, g108}, g308);
	defparam lut_3126.LUT_SIZE = 3;
	defparam lut_3126.mask = 8'h07;

	lut_sub lut_3136 ({g221, g181, g118, g270}, g309);
	defparam lut_3136.LUT_SIZE = 4;
	defparam lut_3136.mask = 16'h3323;

	lut_sub lut_3150 ({g20, g99, g304, g264}, g310);
	defparam lut_3150.LUT_SIZE = 4;
	defparam lut_3150.mask = 16'h0f07;

	lut_sub lut_3164 ({g21, g297, g134, g304}, g311);
	defparam lut_3164.LUT_SIZE = 4;
	defparam lut_3164.mask = 16'h1333;

	lut_sub lut_3178 ({g134, g220, g221, g181}, g312);
	defparam lut_3178.LUT_SIZE = 4;
	defparam lut_3178.mask = 16'h00df;

	lut_sub lut_3194 ({g307, g308, g309, g310, g311, g312}, g313);
	defparam lut_3194.LUT_SIZE = 6;
	defparam lut_3194.mask = 64'h0000000080000000;

	lut_sub lut_3201 ({i_8_, g20, g108, g222}, g314);
	defparam lut_3201.LUT_SIZE = 4;
	defparam lut_3201.mask = 16'h3100;

	lut_sub lut_3210 ({i_8_, g304, g108, g270}, g315);
	defparam lut_3210.LUT_SIZE = 4;
	defparam lut_3210.mask = 16'h2300;

	lut_sub lut_3218 ({g13, g131}, g316);
	defparam lut_3218.LUT_SIZE = 2;
	defparam lut_3218.mask = 4'b0001;

	lut_sub lut_3225 ({i_8_, g108, g316, g216}, g317);
	defparam lut_3225.LUT_SIZE = 4;
	defparam lut_3225.mask = 16'h0700;

	lut_sub lut_3234 ({i_8_, g206, g181, g108}, g318);
	defparam lut_3234.LUT_SIZE = 4;
	defparam lut_3234.mask = 16'h5100;

	lut_sub lut_3243 ({i_8_, g220, g221, g108}, g319);
	defparam lut_3243.LUT_SIZE = 4;
	defparam lut_3243.mask = 16'h4500;

	lut_sub lut_3253 ({g134, g206, g149, g222}, g320);
	defparam lut_3253.LUT_SIZE = 4;
	defparam lut_3253.mask = 16'hcf0a;

	lut_sub lut_3270 ({g314, g315, g317, g318, g319, g320}, g321);
	defparam lut_3270.LUT_SIZE = 6;
	defparam lut_3270.mask = 64'h4000000000000000;

	lut_sub lut_3279 ({g301, g1768, g306, g313, g321}, g322);
	defparam lut_3279.LUT_SIZE = 5;
	defparam lut_3279.mask = 32'h00000001;

	lut_sub lut_3285 ({g87, g111}, g323);
	defparam lut_3285.LUT_SIZE = 2;
	defparam lut_3285.mask = 4'b0001;

	lut_sub lut_3292 ({i_8_, g297, g100, g316}, g324);
	defparam lut_3292.LUT_SIZE = 4;
	defparam lut_3292.mask = 16'h0313;

	lut_sub lut_3306 ({g14, g145, g323, g186, g212, g324}, g325);
	defparam lut_3306.LUT_SIZE = 6;
	defparam lut_3306.mask = 64'haaaaaaaa20000000;

	lut_sub lut_3327 ({i_15_, g13}, g326);
	defparam lut_3327.LUT_SIZE = 2;
	defparam lut_3327.mask = 4'b0100;

	lut_sub lut_3333 ({i_10_, g326, g251}, g327);
	defparam lut_3333.LUT_SIZE = 3;
	defparam lut_3333.mask = 8'h01;

	lut_sub lut_3341 ({g270, g316, g216, g207}, g328);
	defparam lut_3341.LUT_SIZE = 4;
	defparam lut_3341.mask = 16'h0080;

	lut_sub lut_3350 ({g297, g134, g264, g328, g146}, g329);
	defparam lut_3350.LUT_SIZE = 5;
	defparam lut_3350.mask = 32'hff305510;

	lut_sub lut_3371 ({g59, g112, g135}, g330);
	defparam lut_3371.LUT_SIZE = 3;
	defparam lut_3371.mask = 8'h80;

	lut_sub lut_3379 ({i_9_, i_10_, g53, g13, g145, g330}, g331);
	defparam lut_3379.LUT_SIZE = 6;
	defparam lut_3379.mask = 64'h0003000a00000000;

	lut_sub lut_3390 ({g21, g304, g118, g112}, g332);
	defparam lut_3390.LUT_SIZE = 4;
	defparam lut_3390.mask = 16'h0357;

	lut_sub lut_3405 ({i_8_, g21, g4, g98, g135, g216}, g333);
	defparam lut_3405.LUT_SIZE = 6;
	defparam lut_3405.mask = 64'h0000000f1111333f;

	lut_sub lut_3431 ({g304, g136, g151, g243, g333}, g334);
	defparam lut_3431.LUT_SIZE = 5;
	defparam lut_3431.mask = 32'haaaa8000;

	lut_sub lut_3449 ({g327, g329, g331, g1761, g332, g334}, g335);
	defparam lut_3449.LUT_SIZE = 6;
	defparam lut_3449.mask = 64'h0000040000000000;

	lut_sub lut_3459 ({g276, g278, g296, g322, g325, g335}, g336);
	defparam lut_3459.LUT_SIZE = 6;
	defparam lut_3459.mask = 64'h0000000000010000;

	lut_sub lut_3466 ({g136, g204, g279}, g337);
	defparam lut_3466.LUT_SIZE = 3;
	defparam lut_3466.mask = 8'h0d;

	lut_sub lut_3473 ({i_8_, i_6_, i_7_, g98}, g338);
	defparam lut_3473.LUT_SIZE = 4;
	defparam lut_3473.mask = 16'hfffb;

	lut_sub lut_3493 ({g18, g182}, g339);
	defparam lut_3493.LUT_SIZE = 2;
	defparam lut_3493.mask = 4'b0100;

	lut_sub lut_3500 ({g172, g338, g339}, g340);
	defparam lut_3500.LUT_SIZE = 3;
	defparam lut_3500.mask = 8'h4c;

	lut_sub lut_3509 ({g203, g268, g338}, g341);
	defparam lut_3509.LUT_SIZE = 3;
	defparam lut_3509.mask = 8'h2a;

	lut_sub lut_3519 ({g112, g203, g224, g254}, g342);
	defparam lut_3519.LUT_SIZE = 4;
	defparam lut_3519.mask = 16'h007f;

	lut_sub lut_3533 ({g112, g323, g226, g231}, g343);
	defparam lut_3533.LUT_SIZE = 4;
	defparam lut_3533.mask = 16'hf311;

	lut_sub lut_3549 ({i_8_, g100, g226, g268, g279, g339}, g344);
	defparam lut_3549.LUT_SIZE = 6;
	defparam lut_3549.mask = 64'h000000000000ff7f;

	lut_sub lut_3572 ({g340, g341, g342, g343, g344}, g345);
	defparam lut_3572.LUT_SIZE = 5;
	defparam lut_3572.mask = 32'h20000000;

	lut_sub lut_3579 ({i_8_, g88, g224, g232}, g346);
	defparam lut_3579.LUT_SIZE = 4;
	defparam lut_3579.mask = 16'h0007;

	lut_sub lut_3591 ({g112, g151, g204, g279, g284, g346}, g347);
	defparam lut_3591.LUT_SIZE = 6;
	defparam lut_3591.mask = 64'h88a800a000a000a0;

	lut_sub lut_3609 ({g323, g224, g232, g339}, g348);
	defparam lut_3609.LUT_SIZE = 4;
	defparam lut_3609.mask = 16'h007f;

	lut_sub lut_3621 ({g182, g122}, g349);
	defparam lut_3621.LUT_SIZE = 2;
	defparam lut_3621.mask = 4'b0010;

	lut_sub lut_3629 ({g112, g232, g349, g339}, g350);
	defparam lut_3629.LUT_SIZE = 4;
	defparam lut_3629.mask = 16'h007f;

	lut_sub lut_3642 ({i_8_, g135, g231, g349}, g351);
	defparam lut_3642.LUT_SIZE = 4;
	defparam lut_3642.mask = 16'h000d;

	lut_sub lut_3653 ({i_8_, g135, g226, g224, g232, g339}, g352);
	defparam lut_3653.LUT_SIZE = 6;
	defparam lut_3653.mask = 64'h000000000000ff7f;

	lut_sub lut_3677 ({g136, g203, g348, g350, g351, g352}, g353);
	defparam lut_3677.LUT_SIZE = 6;
	defparam lut_3677.mask = 64'h8000800080000000;

	lut_sub lut_3686 ({g151, g226, g339}, g354);
	defparam lut_3686.LUT_SIZE = 3;
	defparam lut_3686.mask = 8'h0d;

	lut_sub lut_3695 ({i_8_, g108, g203, g204}, g355);
	defparam lut_3695.LUT_SIZE = 4;
	defparam lut_3695.mask = 16'h000b;

	lut_sub lut_3706 ({i_8_, g108, g226, g224, g231, g232}, g356);
	defparam lut_3706.LUT_SIZE = 6;
	defparam lut_3706.mask = 64'h000000000000ffdf;

	lut_sub lut_3730 ({g323, g151, g203, g349, g355, g356}, g357);
	defparam lut_3730.LUT_SIZE = 6;
	defparam lut_3730.mask = 64'h8888800080008000;

	lut_sub lut_3746 ({g337, g345, g347, g353, g354, g357}, g358);
	defparam lut_3746.LUT_SIZE = 6;
	defparam lut_3746.mask = 64'h0000000400000000;

	lut_sub lut_3755 ({g244, g112, g136, g222, g178}, g359);
	defparam lut_3755.LUT_SIZE = 5;
	defparam lut_3755.mask = 32'h03330377;

	lut_sub lut_3778 ({g145, g112, g136, g222, g151, g284}, g360);
	defparam lut_3778.LUT_SIZE = 6;
	defparam lut_3778.mask = 64'h8880000000000000;

	lut_sub lut_3786 ({i_14_, i_12_, i_13_, g15, g338}, g361);
	defparam lut_3786.LUT_SIZE = 5;
	defparam lut_3786.mask = 32'h00808000;

	lut_sub lut_3794 ({g220, g145, g361}, g362);
	defparam lut_3794.LUT_SIZE = 3;
	defparam lut_3794.mask = 8'ha8;

	lut_sub lut_3803 ({i_8_, g20, g108, g222}, g363);
	defparam lut_3803.LUT_SIZE = 4;
	defparam lut_3803.mask = 16'h0031;

	lut_sub lut_3812 ({i_8_, g221, g88, g270}, g364);
	defparam lut_3812.LUT_SIZE = 4;
	defparam lut_3812.mask = 16'h0032;

	lut_sub lut_3821 ({i_8_, g206, g88, g181}, g365);
	defparam lut_3821.LUT_SIZE = 4;
	defparam lut_3821.mask = 16'h0031;

	lut_sub lut_3830 ({i_8_, g206, g108, g185}, g366);
	defparam lut_3830.LUT_SIZE = 4;
	defparam lut_3830.mask = 16'h0032;

	lut_sub lut_3840 ({i_8_, g304, g108, g270, g216}, g367);
	defparam lut_3840.LUT_SIZE = 5;
	defparam lut_3840.mask = 32'h00000d0f;

	lut_sub lut_3855 ({g363, g364, g365, g366, g367}, g368);
	defparam lut_3855.LUT_SIZE = 5;
	defparam lut_3855.mask = 32'h80000000;

	lut_sub lut_3861 ({i_8_, g304, g100}, g369);
	defparam lut_3861.LUT_SIZE = 3;
	defparam lut_3861.mask = 8'h01;

	lut_sub lut_3868 ({i_8_, g206, g221, g135}, g370);
	defparam lut_3868.LUT_SIZE = 4;
	defparam lut_3868.mask = 16'h0054;

	lut_sub lut_3877 ({g220, g112, g316}, g371);
	defparam lut_3877.LUT_SIZE = 3;
	defparam lut_3877.mask = 8'h13;

	lut_sub lut_3887 ({i_8_, g88, g135, g316, g284}, g372);
	defparam lut_3887.LUT_SIZE = 5;
	defparam lut_3887.mask = 32'h11111333;

	lut_sub lut_3907 ({g270, g136, g369, g370, g371, g372}, g373);
	defparam lut_3907.LUT_SIZE = 6;
	defparam lut_3907.mask = 64'h8000000080008000;

	lut_sub lut_3919 ({g359, g1754, g360, g362, g368, g373}, g374);
	defparam lut_3919.LUT_SIZE = 6;
	defparam lut_3919.mask = 64'h0001010100010001;

	lut_sub lut_3930 ({i_8_, g4, g87, g182}, g375);
	defparam lut_3930.LUT_SIZE = 4;
	defparam lut_3930.mask = 16'h0001;

	lut_sub lut_3935 ({i_11_, i_9_, i_15_, g375}, g376);
	defparam lut_3935.LUT_SIZE = 4;
	defparam lut_3935.mask = 16'h1000;

	lut_sub lut_3941 ({i_8_, g34, g110}, g377);
	defparam lut_3941.LUT_SIZE = 3;
	defparam lut_3941.mask = 8'h01;

	lut_sub lut_3947 ({i_11_, g141, g377}, g378);
	defparam lut_3947.LUT_SIZE = 3;
	defparam lut_3947.mask = 8'h10;

	lut_sub lut_3955 ({g112, g323, g191, g201}, g379);
	defparam lut_3955.LUT_SIZE = 4;
	defparam lut_3955.mask = 16'h03ab;

	lut_sub lut_3971 ({g145, g151, g213, g209, g378, g379}, g380);
	defparam lut_3971.LUT_SIZE = 6;
	defparam lut_3971.mask = 64'h8888880080808000;

	lut_sub lut_3987 ({i_11_, g5, g112, g253, g377}, g381);
	defparam lut_3987.LUT_SIZE = 5;
	defparam lut_3987.mask = 32'h03570303;

	lut_sub lut_4003 ({i_5_, i_3_, g57, g111}, g382);
	defparam lut_4003.LUT_SIZE = 4;
	defparam lut_4003.mask = 16'h0010;

	lut_sub lut_4013 ({g98, g112, g316, g268, g381, g382}, g383);
	defparam lut_4013.LUT_SIZE = 6;
	defparam lut_4013.mask = 64'hccc8c8c8cc88c888;

	lut_sub lut_4043 ({i_9_, i_10_, g53, g323, g182}, g384);
	defparam lut_4043.LUT_SIZE = 5;
	defparam lut_4043.mask = 32'h05000100;

	lut_sub lut_4054 ({g323, g151, g209, g284, g384}, g385);
	defparam lut_4054.LUT_SIZE = 5;
	defparam lut_4054.mask = 32'h11551555;

	lut_sub lut_4073 ({i_8_, g100, g191, g201}, g386);
	defparam lut_4073.LUT_SIZE = 4;
	defparam lut_4073.mask = 16'h000b;

	lut_sub lut_4082 ({i_8_, g100, g193, g232}, g387);
	defparam lut_4082.LUT_SIZE = 4;
	defparam lut_4082.mask = 16'h0007;

	lut_sub lut_4091 ({i_8_, g135, g187, g193}, g388);
	defparam lut_4091.LUT_SIZE = 4;
	defparam lut_4091.mask = 16'h0007;

	lut_sub lut_4101 ({g112, g183, g187, g193}, g389);
	defparam lut_4101.LUT_SIZE = 4;
	defparam lut_4101.mask = 16'h007f;

	lut_sub lut_4116 ({i_8_, g108, g323, g187, g201, g213}, g390);
	defparam lut_4116.LUT_SIZE = 6;
	defparam lut_4116.mask = 64'hff20ff20ff20a020;

	lut_sub lut_4154 ({g386, g387, g388, g389, g390}, g391);
	defparam lut_4154.LUT_SIZE = 5;
	defparam lut_4154.mask = 32'h40000000;

	lut_sub lut_4161 ({i_8_, g88, g193, g255}, g392);
	defparam lut_4161.LUT_SIZE = 4;
	defparam lut_4161.mask = 16'h0007;

	lut_sub lut_4170 ({i_8_, g100, g213, g253}, g393);
	defparam lut_4170.LUT_SIZE = 4;
	defparam lut_4170.mask = 16'h0007;

	lut_sub lut_4179 ({i_8_, g100, g187, g231}, g394);
	defparam lut_4179.LUT_SIZE = 4;
	defparam lut_4179.mask = 16'h000b;

	lut_sub lut_4188 ({i_8_, g100, g224, g349}, g395);
	defparam lut_4188.LUT_SIZE = 4;
	defparam lut_4188.mask = 16'h0007;

	lut_sub lut_4199 ({i_8_, g135, g183, g191, g201, g338}, g396);
	defparam lut_4199.LUT_SIZE = 6;
	defparam lut_4199.mask = 64'h8a8a8a8a8a8aceff;

	lut_sub lut_4238 ({g392, g393, g394, g395, g396}, g397);
	defparam lut_4238.LUT_SIZE = 5;
	defparam lut_4238.mask = 32'h80000000;

	lut_sub lut_4248 ({g376, g380, g383, g385, g391, g397}, g398);
	defparam lut_4248.LUT_SIZE = 6;
	defparam lut_4248.mask = 64'h0000001000000000;

	lut_sub lut_4254 ({g142, g117}, g399);
	defparam lut_4254.LUT_SIZE = 2;
	defparam lut_4254.mask = 4'b1000;

	lut_sub lut_4259 ({i_6_, g58}, g400);
	defparam lut_4259.LUT_SIZE = 2;
	defparam lut_4259.mask = 4'b0001;

	lut_sub lut_4268 ({i_8_, g88, g132, g94, g165, g400}, g401);
	defparam lut_4268.LUT_SIZE = 6;
	defparam lut_4268.mask = 64'h000000005500ff3f;

	lut_sub lut_4292 ({g136, g399, g401}, g402);
	defparam lut_4292.LUT_SIZE = 3;
	defparam lut_4292.mask = 8'ha2;

	lut_sub lut_4303 ({i_8_, g88, g135, g159, g92, g96}, g403);
	defparam lut_4303.LUT_SIZE = 6;
	defparam lut_4303.mask = 64'h0000000000afcfef;

	lut_sub lut_4330 ({g101, g112, g103, g96, g403}, g404);
	defparam lut_4330.LUT_SIZE = 5;
	defparam lut_4330.mask = 32'haa0a2202;

	lut_sub lut_4345 ({g112, g132, g159}, g405);
	defparam lut_4345.LUT_SIZE = 3;
	defparam lut_4345.mask = 8'h0d;

	lut_sub lut_4354 ({i_8_, g108, g94, g116}, g406);
	defparam lut_4354.LUT_SIZE = 4;
	defparam lut_4354.mask = 16'h0007;

	lut_sub lut_4363 ({i_8_, g100, g108, g132}, g407);
	defparam lut_4363.LUT_SIZE = 4;
	defparam lut_4363.mask = 16'h002a;

	lut_sub lut_4372 ({g112, g94, g92}, g408);
	defparam lut_4372.LUT_SIZE = 3;
	defparam lut_4372.mask = 8'h0b;

	lut_sub lut_4382 ({i_8_, g112, g135, g142, g90}, g409);
	defparam lut_4382.LUT_SIZE = 5;
	defparam lut_4382.mask = 32'h00bb0abb;

	lut_sub lut_4404 ({g405, g406, g407, g408, g409}, g410);
	defparam lut_4404.LUT_SIZE = 5;
	defparam lut_4404.mask = 32'h80000000;

	lut_sub lut_4414 ({g338, g399, g402, g404, g410, g1747}, g411);
	defparam lut_4414.LUT_SIZE = 6;
	defparam lut_4414.mask = 64'h0000000100010001;

	lut_sub lut_4425 ({g15, g91, g131, g182, g268}, g412);
	defparam lut_4425.LUT_SIZE = 5;
	defparam lut_4425.mask = 32'h8088a0a8;

	lut_sub lut_4438 ({i_8_, g135, g172}, g413);
	defparam lut_4438.LUT_SIZE = 3;
	defparam lut_4438.mask = 8'h01;

	lut_sub lut_4445 ({i_8_, g108, g349, g339}, g414);
	defparam lut_4445.LUT_SIZE = 4;
	defparam lut_4445.mask = 16'h0007;

	lut_sub lut_4454 ({i_14_, i_12_, i_13_, g95, g112, g323}, g415);
	defparam lut_4454.LUT_SIZE = 6;
	defparam lut_4454.mask = 64'h0000050003070000;

	lut_sub lut_4468 ({i_8_, g100, g135, g94, g127}, g416);
	defparam lut_4468.LUT_SIZE = 5;
	defparam lut_4468.mask = 32'h00000a3b;

	lut_sub lut_4484 ({g151, g280, g413, g414, g415, g416}, g417);
	defparam lut_4484.LUT_SIZE = 6;
	defparam lut_4484.mask = 64'h8000800080000000;

	lut_sub lut_4494 ({i_9_, i_10_, g53, g145, g146, g182}, g418);
	defparam lut_4494.LUT_SIZE = 6;
	defparam lut_4494.mask = 64'h0005004400000000;

	lut_sub lut_4505 ({g136, g412, g417, g418}, g419);
	defparam lut_4505.LUT_SIZE = 4;
	defparam lut_4505.mask = 16'h2202;

	lut_sub lut_4516 ({g358, g374, g398, g411, g419}, g420);
	defparam lut_4516.LUT_SIZE = 5;
	defparam lut_4516.mask = 32'h00000001;

	lut_sub lut_4525 ({g203, g199, g224, g177, g339}, g421);
	defparam lut_4525.LUT_SIZE = 5;
	defparam lut_4525.mask = 32'h80000000;

	lut_sub lut_4534 ({g134, g109, g172, g349, g421}, g422);
	defparam lut_4534.LUT_SIZE = 5;
	defparam lut_4534.mask = 32'hffcc5040;

	lut_sub lut_4554 ({g31, g87}, g423);
	defparam lut_4554.LUT_SIZE = 2;
	defparam lut_4554.mask = 4'b0001;

	lut_sub lut_4560 ({i_15_, g113, g182}, g424);
	defparam lut_4560.LUT_SIZE = 3;
	defparam lut_4560.mask = 8'h01;

	lut_sub lut_4566 ({g423, g424}, g425);
	defparam lut_4566.LUT_SIZE = 2;
	defparam lut_4566.mask = 4'b0001;

	lut_sub lut_4573 ({g204, g279, g285}, g426);
	defparam lut_4573.LUT_SIZE = 3;
	defparam lut_4573.mask = 8'ha2;

	lut_sub lut_4581 ({g203, g214}, g427);
	defparam lut_4581.LUT_SIZE = 2;
	defparam lut_4581.mask = 4'b0001;

	lut_sub lut_4586 ({i_5_, i_3_, i_4_, g57}, g428);
	defparam lut_4586.LUT_SIZE = 4;
	defparam lut_4586.mask = 16'h1040;

	lut_sub lut_4593 ({g31, g428}, g429);
	defparam lut_4593.LUT_SIZE = 2;
	defparam lut_4593.mask = 4'b0001;

	lut_sub lut_4600 ({g110, g111, g177}, g430);
	defparam lut_4600.LUT_SIZE = 3;
	defparam lut_4600.mask = 8'h01;

	lut_sub lut_4607 ({g31, g110, g199}, g431);
	defparam lut_4607.LUT_SIZE = 3;
	defparam lut_4607.mask = 8'h01;

	lut_sub lut_4617 ({g59, g99, g172, g339, g430, g431}, g432);
	defparam lut_4617.LUT_SIZE = 6;
	defparam lut_4617.mask = 64'h8888800080008000;

	lut_sub lut_4633 ({g277, g232, g339, g427, g429, g432}, g433);
	defparam lut_4633.LUT_SIZE = 6;
	defparam lut_4633.mask = 64'h5040000050405040;

	lut_sub lut_4648 ({g134, g118, g231}, g434);
	defparam lut_4648.LUT_SIZE = 3;
	defparam lut_4648.mask = 8'h2a;

	lut_sub lut_4657 ({g118, g224, g197}, g435);
	defparam lut_4657.LUT_SIZE = 3;
	defparam lut_4657.mask = 8'h07;

	lut_sub lut_4667 ({i_8_, g134, g135, g177, g173}, g436);
	defparam lut_4667.LUT_SIZE = 5;
	defparam lut_4667.mask = 32'h00550757;

	lut_sub lut_4685 ({i_8_, g100, g177, g172}, g437);
	defparam lut_4685.LUT_SIZE = 4;
	defparam lut_4685.mask = 16'h0007;

	lut_sub lut_4695 ({i_8_, g108, g226, g224, g231}, g438);
	defparam lut_4695.LUT_SIZE = 5;
	defparam lut_4695.mask = 32'h00fb0000;

	lut_sub lut_4710 ({g434, g435, g436, g437, g438}, g439);
	defparam lut_4710.LUT_SIZE = 5;
	defparam lut_4710.mask = 32'h80000000;

	lut_sub lut_4719 ({i_8_, g4, g98, g195, g197, g173}, g440);
	defparam lut_4719.LUT_SIZE = 6;
	defparam lut_4719.mask = 64'h0000005f0000003f;

	lut_sub lut_4740 ({g109, g146, g195, g232, g173, g440}, g441);
	defparam lut_4740.LUT_SIZE = 6;
	defparam lut_4740.mask = 64'haa00aaaa80008080;

	lut_sub lut_4761 ({i_8_, g88, g224, g197}, g442);
	defparam lut_4761.LUT_SIZE = 4;
	defparam lut_4761.mask = 16'h0700;

	lut_sub lut_4773 ({g109, g203, g268, g172, g339, g442}, g443);
	defparam lut_4773.LUT_SIZE = 6;
	defparam lut_4773.mask = 64'haaaaaaaa80000000;

	lut_sub lut_4796 ({i_8_, g88, g323, g231}, g444);
	defparam lut_4796.LUT_SIZE = 4;
	defparam lut_4796.mask = 16'h2a22;

	lut_sub lut_4807 ({i_8_, g88, g232, g339}, g445);
	defparam lut_4807.LUT_SIZE = 4;
	defparam lut_4807.mask = 16'h0700;

	lut_sub lut_4816 ({i_8_, g88, g226, g349}, g446);
	defparam lut_4816.LUT_SIZE = 4;
	defparam lut_4816.mask = 16'h0d00;

	lut_sub lut_4825 ({g134, g226, g349}, g447);
	defparam lut_4825.LUT_SIZE = 3;
	defparam lut_4825.mask = 8'h0d;

	lut_sub lut_4835 ({g224, g232, g349, g423}, g448);
	defparam lut_4835.LUT_SIZE = 4;
	defparam lut_4835.mask = 16'h1555;

	lut_sub lut_4849 ({g118, g226, g203, g349}, g449);
	defparam lut_4849.LUT_SIZE = 4;
	defparam lut_4849.mask = 16'h00f7;

	lut_sub lut_4865 ({g444, g445, g446, g447, g448, g449}, g450);
	defparam lut_4865.LUT_SIZE = 6;
	defparam lut_4865.mask = 64'h8000000000000000;

	lut_sub lut_4872 ({g99, g226, g177}, g451);
	defparam lut_4872.LUT_SIZE = 3;
	defparam lut_4872.mask = 8'h0d;

	lut_sub lut_4881 ({g149, g226, g177}, g452);
	defparam lut_4881.LUT_SIZE = 3;
	defparam lut_4881.mask = 8'hf2;

	lut_sub lut_4892 ({g59, g203, g224}, g453);
	defparam lut_4892.LUT_SIZE = 3;
	defparam lut_4892.mask = 8'h07;

	lut_sub lut_4901 ({g149, g199, g349}, g454);
	defparam lut_4901.LUT_SIZE = 3;
	defparam lut_4901.mask = 8'h07;

	lut_sub lut_4912 ({g99, g199, g197, g268, g349}, g455);
	defparam lut_4912.LUT_SIZE = 5;
	defparam lut_4912.mask = 32'h00007fff;

	lut_sub lut_4935 ({g451, g452, g453, g454, g455}, g456);
	defparam lut_4935.LUT_SIZE = 5;
	defparam lut_4935.mask = 32'h00800000;

	lut_sub lut_4945 ({g433, g439, g441, g443, g450, g456}, g457);
	defparam lut_4945.LUT_SIZE = 6;
	defparam lut_4945.mask = 64'h0000000000000001;

	lut_sub lut_4955 ({g136, g195, g422, g425, g426, g457}, g458);
	defparam lut_4955.LUT_SIZE = 6;
	defparam lut_4955.mask = 64'h0040004000400000;

	lut_sub lut_4967 ({g73, g169, g275, g336, g420, g458}, o_3_);
	defparam lut_4967.LUT_SIZE = 6;
	defparam lut_4967.mask = 64'h00000000fffffffe;

	lut_sub lut_5003 ({g48, g158}, g460);
	defparam lut_5003.LUT_SIZE = 2;
	defparam lut_5003.mask = 4'b0100;

	lut_sub lut_5007 ({i_14_, i_12_, i_13_}, g461);
	defparam lut_5007.LUT_SIZE = 3;
	defparam lut_5007.mask = 8'h10;

	lut_sub lut_5013 ({g18, g461}, g462);
	defparam lut_5013.LUT_SIZE = 2;
	defparam lut_5013.mask = 4'b1011;

	lut_sub lut_5022 ({g151, g460, g462}, g463);
	defparam lut_5022.LUT_SIZE = 3;
	defparam lut_5022.mask = 8'h0b;

	lut_sub lut_5030 ({i_11_, i_15_, g113, g48}, g464);
	defparam lut_5030.LUT_SIZE = 4;
	defparam lut_5030.mask = 16'hfdff;

	lut_sub lut_5050 ({i_11_, i_15_, g141, g48}, g465);
	defparam lut_5050.LUT_SIZE = 4;
	defparam lut_5050.mask = 16'hfdff;

	lut_sub lut_5070 ({g284, g460}, g466);
	defparam lut_5070.LUT_SIZE = 2;
	defparam lut_5070.mask = 4'b0001;

	lut_sub lut_5076 ({g6, i_15_, g48}, g467);
	defparam lut_5076.LUT_SIZE = 3;
	defparam lut_5076.mask = 8'hfd;

	lut_sub lut_5088 ({g6, i_15_, g461}, g468);
	defparam lut_5088.LUT_SIZE = 3;
	defparam lut_5088.mask = 8'hfe;

	lut_sub lut_5101 ({g112, g467, g468}, g469);
	defparam lut_5101.LUT_SIZE = 3;
	defparam lut_5101.mask = 8'h0e;

	lut_sub lut_5109 ({g158, g461}, g470);
	defparam lut_5109.LUT_SIZE = 2;
	defparam lut_5109.mask = 4'b0001;

	lut_sub lut_5117 ({g87, g110, g111, g465}, g471);
	defparam lut_5117.LUT_SIZE = 4;
	defparam lut_5117.mask = 16'h0222;

	lut_sub lut_5128 ({i_8_, g135, g323, g467, g470, g471}, g472);
	defparam lut_5128.LUT_SIZE = 6;
	defparam lut_5128.mask = 64'haa0aaa0aaa0a8808;

	lut_sub lut_5158 ({g101, g464, g465, g466, g469, g472}, g473);
	defparam lut_5158.LUT_SIZE = 6;
	defparam lut_5158.mask = 64'h4040404000000040;

	lut_sub lut_5168 ({g48, g93}, g474);
	defparam lut_5168.LUT_SIZE = 2;
	defparam lut_5168.mask = 4'b1000;

	lut_sub lut_5174 ({g93, g461}, g475);
	defparam lut_5174.LUT_SIZE = 2;
	defparam lut_5174.mask = 4'b1011;

	lut_sub lut_5183 ({g338, g474, g475}, g476);
	defparam lut_5183.LUT_SIZE = 3;
	defparam lut_5183.mask = 8'hb0;

	lut_sub lut_5191 ({g48, g115}, g477);
	defparam lut_5191.LUT_SIZE = 2;
	defparam lut_5191.mask = 4'b0111;

	lut_sub lut_5199 ({g48, g124}, g478);
	defparam lut_5199.LUT_SIZE = 2;
	defparam lut_5199.mask = 4'b0100;

	lut_sub lut_5207 ({g112, g323, g477, g478}, g479);
	defparam lut_5207.LUT_SIZE = 4;
	defparam lut_5207.mask = 16'hf322;

	lut_sub lut_5221 ({g112, g323, g464}, g480);
	defparam lut_5221.LUT_SIZE = 3;
	defparam lut_5221.mask = 8'h2a;

	lut_sub lut_5229 ({g48, g122}, g481);
	defparam lut_5229.LUT_SIZE = 2;
	defparam lut_5229.mask = 4'b0111;

	lut_sub lut_5238 ({g323, g481, g474}, g482);
	defparam lut_5238.LUT_SIZE = 3;
	defparam lut_5238.mask = 8'h0d;

	lut_sub lut_5249 ({i_8_, g88, g112, g460, g470, g475}, g483);
	defparam lut_5249.LUT_SIZE = 6;
	defparam lut_5249.mask = 64'hff40ff40ff40cc40;

	lut_sub lut_5289 ({g476, g479, g480, g482, g483}, g484);
	defparam lut_5289.LUT_SIZE = 5;
	defparam lut_5289.mask = 32'h00400000;

	lut_sub lut_5295 ({g122, g461}, g485);
	defparam lut_5295.LUT_SIZE = 2;
	defparam lut_5295.mask = 4'b0100;

	lut_sub lut_5302 ({g145, g485, g475}, g486);
	defparam lut_5302.LUT_SIZE = 3;
	defparam lut_5302.mask = 8'h0b;

	lut_sub lut_5310 ({g115, g461}, g487);
	defparam lut_5310.LUT_SIZE = 2;
	defparam lut_5310.mask = 4'b0100;

	lut_sub lut_5317 ({g145, g487, g462}, g488);
	defparam lut_5317.LUT_SIZE = 3;
	defparam lut_5317.mask = 8'h0b;

	lut_sub lut_5325 ({i_11_, i_9_, i_10_, i_15_, g48, g136}, g489);
	defparam lut_5325.LUT_SIZE = 6;
	defparam lut_5325.mask = 64'h0004040404040004;

	lut_sub lut_5340 ({g463, g473, g484, g486, g488, g489}, g490);
	defparam lut_5340.LUT_SIZE = 6;
	defparam lut_5340.mask = 64'h0000008000000000;

	lut_sub lut_5346 ({g112, g485}, g491);
	defparam lut_5346.LUT_SIZE = 2;
	defparam lut_5346.mask = 4'b1110;

	lut_sub lut_5356 ({g59, g135, g474, g460}, g492);
	defparam lut_5356.LUT_SIZE = 4;
	defparam lut_5356.mask = 16'hfac8;

	lut_sub lut_5373 ({g99, g118, g464, g467, g468}, g493);
	defparam lut_5373.LUT_SIZE = 5;
	defparam lut_5373.mask = 32'hff010f01;

	lut_sub lut_5394 ({g59, g429, g465, g493}, g494);
	defparam lut_5394.LUT_SIZE = 4;
	defparam lut_5394.mask = 16'h5111;

	lut_sub lut_5404 ({g30, g110}, g495);
	defparam lut_5404.LUT_SIZE = 2;
	defparam lut_5404.mask = 4'b0001;

	lut_sub lut_5412 ({g124, g461, g474, g495}, g496);
	defparam lut_5412.LUT_SIZE = 4;
	defparam lut_5412.mask = 16'h1115;

	lut_sub lut_5423 ({g109, g465, g462}, g497);
	defparam lut_5423.LUT_SIZE = 3;
	defparam lut_5423.mask = 8'h0e;

	lut_sub lut_5432 ({i_8_, i_7_, g400, g467, g487}, g498);
	defparam lut_5432.LUT_SIZE = 5;
	defparam lut_5432.mask = 32'h050c0000;

	lut_sub lut_5444 ({g323, g478, g496, g497, g498}, g499);
	defparam lut_5444.LUT_SIZE = 5;
	defparam lut_5444.mask = 32'h80808000;

	lut_sub lut_5453 ({g118, g478, g487}, g500);
	defparam lut_5453.LUT_SIZE = 3;
	defparam lut_5453.mask = 8'h07;

	lut_sub lut_5463 ({g18, g118, g228, g461}, g501);
	defparam lut_5463.LUT_SIZE = 4;
	defparam lut_5463.mask = 16'h0501;

	lut_sub lut_5473 ({g22, g88, g124, g461}, g502);
	defparam lut_5473.LUT_SIZE = 4;
	defparam lut_5473.mask = 16'h0105;

	lut_sub lut_5484 ({g22, g134, g93, g124, g461}, g503);
	defparam lut_5484.LUT_SIZE = 5;
	defparam lut_5484.mask = 32'h00510055;

	lut_sub lut_5500 ({g134, g149, g99, g423, g481, g467}, g504);
	defparam lut_5500.LUT_SIZE = 6;
	defparam lut_5500.mask = 64'hf131313131313131;

	lut_sub lut_5534 ({g500, g501, g502, g503, g504}, g505);
	defparam lut_5534.LUT_SIZE = 5;
	defparam lut_5534.mask = 32'h40000000;

	lut_sub lut_5540 ({g22, g461}, g506);
	defparam lut_5540.LUT_SIZE = 2;
	defparam lut_5540.mask = 4'b0001;

	lut_sub lut_5547 ({i_8_, g108, g506, g470}, g507);
	defparam lut_5547.LUT_SIZE = 4;
	defparam lut_5547.mask = 16'h0703;

	lut_sub lut_5559 ({g136, g124, g115, g461}, g508);
	defparam lut_5559.LUT_SIZE = 4;
	defparam lut_5559.mask = 16'h0045;

	lut_sub lut_5569 ({i_8_, g108, g124, g115, g461}, g509);
	defparam lut_5569.LUT_SIZE = 5;
	defparam lut_5569.mask = 32'h00450005;

	lut_sub lut_5580 ({i_8_, g108, g474, g475}, g510);
	defparam lut_5580.LUT_SIZE = 4;
	defparam lut_5580.mask = 16'h0b00;

	lut_sub lut_5591 ({g149, g109, g477, g485, g510}, g511);
	defparam lut_5591.LUT_SIZE = 5;
	defparam lut_5591.mask = 32'haa088808;

	lut_sub lut_5607 ({g505, g507, g508, g509, g511}, g512);
	defparam lut_5607.LUT_SIZE = 5;
	defparam lut_5607.mask = 32'h00004000;

	lut_sub lut_5616 ({g110, g111, g428, g487, g506}, g513);
	defparam lut_5616.LUT_SIZE = 5;
	defparam lut_5616.mask = 32'h00030057;

	lut_sub lut_5629 ({i_8_, g88, g108, g468}, g514);
	defparam lut_5629.LUT_SIZE = 4;
	defparam lut_5629.mask = 16'h222a;

	lut_sub lut_5642 ({i_8_, g135, g485, g506, g468, g475}, g515);
	defparam lut_5642.LUT_SIZE = 6;
	defparam lut_5642.mask = 64'h0000cccc0000efff;

	lut_sub lut_5673 ({g100, g506, g513, g514, g515}, g516);
	defparam lut_5673.LUT_SIZE = 5;
	defparam lut_5673.mask = 32'h80808000;

	lut_sub lut_5684 ({g464, g467, g474, g465, g485}, g517);
	defparam lut_5684.LUT_SIZE = 5;
	defparam lut_5684.mask = 32'h00000020;

	lut_sub lut_5689 ({i_11_, i_10_, i_15_, g461}, g518);
	defparam lut_5689.LUT_SIZE = 4;
	defparam lut_5689.mask = 16'h0010;

	lut_sub lut_5699 ({g134, g145, g151, g470, g517, g518}, g519);
	defparam lut_5699.LUT_SIZE = 6;
	defparam lut_5699.mask = 64'hffaaf0a030203020;

	lut_sub lut_5730 ({g109, g460, g516, g519}, g520);
	defparam lut_5730.LUT_SIZE = 4;
	defparam lut_5730.mask = 16'h1110;

	lut_sub lut_5742 ({g490, g1737, g499, g1728, g512, g520}, g521);
	defparam lut_5742.LUT_SIZE = 6;
	defparam lut_5742.mask = 64'h0000000000000001;

	lut_sub lut_5748 ({g93, g171}, g522);
	defparam lut_5748.LUT_SIZE = 2;
	defparam lut_5748.mask = 4'b1000;

	lut_sub lut_5756 ({g100, g212, g251, g522}, g523);
	defparam lut_5756.LUT_SIZE = 4;
	defparam lut_5756.mask = 16'h5155;

	lut_sub lut_5767 ({i_11_, i_9_, i_15_, g375}, g524);
	defparam lut_5767.LUT_SIZE = 4;
	defparam lut_5767.mask = 16'h0010;

	lut_sub lut_5774 ({i_11_, i_9_, g326, g98, g111}, g525);
	defparam lut_5774.LUT_SIZE = 5;
	defparam lut_5774.mask = 32'h00000100;

	lut_sub lut_5784 ({g297, g216, g227, g231, g238, g349}, g526);
	defparam lut_5784.LUT_SIZE = 6;
	defparam lut_5784.mask = 64'hff0acc08cc08cc08;

	lut_sub lut_5817 ({g261, g523, g524, g525, g526}, g527);
	defparam lut_5817.LUT_SIZE = 5;
	defparam lut_5817.mask = 32'h40000000;

	lut_sub lut_5823 ({g45, g197}, g528);
	defparam lut_5823.LUT_SIZE = 2;
	defparam lut_5823.mask = 4'b1000;

	lut_sub lut_5829 ({g467, g528}, g529);
	defparam lut_5829.LUT_SIZE = 2;
	defparam lut_5829.mask = 4'b0001;

	lut_sub lut_5835 ({g22, g171}, g530);
	defparam lut_5835.LUT_SIZE = 2;
	defparam lut_5835.mask = 4'b0010;

	lut_sub lut_5841 ({g6, i_15_, g171}, g531);
	defparam lut_5841.LUT_SIZE = 3;
	defparam lut_5841.mask = 8'h02;

	lut_sub lut_5847 ({g13, g124}, g532);
	defparam lut_5847.LUT_SIZE = 2;
	defparam lut_5847.mask = 4'b0001;

	lut_sub lut_5855 ({g134, g195, g532, g478}, g533);
	defparam lut_5855.LUT_SIZE = 4;
	defparam lut_5855.mask = 16'h007f;

	lut_sub lut_5867 ({g171, g124}, g534);
	defparam lut_5867.LUT_SIZE = 2;
	defparam lut_5867.mask = 4'b0100;

	lut_sub lut_5874 ({g45, g224, g467}, g535);
	defparam lut_5874.LUT_SIZE = 3;
	defparam lut_5874.mask = 8'h40;

	lut_sub lut_5883 ({g99, g534, g530, g531, g535}, g536);
	defparam lut_5883.LUT_SIZE = 5;
	defparam lut_5883.mask = 32'h0000bfff;

	lut_sub lut_5906 ({g423, g464, g478, g533, g536}, g537);
	defparam lut_5906.LUT_SIZE = 5;
	defparam lut_5906.mask = 32'h88880080;

	lut_sub lut_5916 ({i_8_, i_6_, i_7_, g98, g87}, g538);
	defparam lut_5916.LUT_SIZE = 5;
	defparam lut_5916.mask = 32'h57330700;

	lut_sub lut_5937 ({g99, g251, g277, g158, g285, g538}, g539);
	defparam lut_5937.LUT_SIZE = 6;
	defparam lut_5937.mask = 64'h00a200a000a000a0;

	lut_sub lut_5951 ({g171, g122}, g540);
	defparam lut_5951.LUT_SIZE = 2;
	defparam lut_5951.mask = 4'b1000;

	lut_sub lut_5956 ({i_11_, i_9_, i_10_, i_15_, g171}, g541);
	defparam lut_5956.LUT_SIZE = 5;
	defparam lut_5956.mask = 32'h20000020;

	lut_sub lut_5966 ({g99, g251, g285, g540, g541}, g542);
	defparam lut_5966.LUT_SIZE = 5;
	defparam lut_5966.mask = 32'h51555555;

	lut_sub lut_5990 ({g109, g529, g1721, g537, g539, g542}, g543);
	defparam lut_5990.LUT_SIZE = 6;
	defparam lut_5990.mask = 64'h000b000b0000000b;

	lut_sub lut_6004 ({g6, i_15_, g461}, g544);
	defparam lut_6004.LUT_SIZE = 3;
	defparam lut_6004.mask = 8'hfb;

	lut_sub lut_6017 ({g45, g118, g544}, g545);
	defparam lut_6017.LUT_SIZE = 3;
	defparam lut_6017.mask = 8'h23;

	lut_sub lut_6025 ({g13, g115}, g546);
	defparam lut_6025.LUT_SIZE = 2;
	defparam lut_6025.mask = 4'b0010;

	lut_sub lut_6031 ({g13, g122}, g547);
	defparam lut_6031.LUT_SIZE = 2;
	defparam lut_6031.mask = 4'b1101;

	lut_sub lut_6039 ({g119, g461}, g548);
	defparam lut_6039.LUT_SIZE = 2;
	defparam lut_6039.mask = 4'b0001;

	lut_sub lut_6045 ({g547, g548}, g549);
	defparam lut_6045.LUT_SIZE = 2;
	defparam lut_6045.mask = 4'b0010;

	lut_sub lut_6051 ({g102, g461}, g550);
	defparam lut_6051.LUT_SIZE = 2;
	defparam lut_6051.mask = 4'b0100;

	lut_sub lut_6057 ({g104, g461}, g551);
	defparam lut_6057.LUT_SIZE = 2;
	defparam lut_6057.mask = 4'b0001;

	lut_sub lut_6066 ({i_8_, g108, g135, g550, g546, g551}, g552);
	defparam lut_6066.LUT_SIZE = 6;
	defparam lut_6066.mask = 64'h00000f0f007f557f;

	lut_sub lut_6100 ({g149, g151, g549, g532, g552}, g553);
	defparam lut_6100.LUT_SIZE = 5;
	defparam lut_6100.mask = 32'haa880a08;

	lut_sub lut_6114 ({g95, g461}, g554);
	defparam lut_6114.LUT_SIZE = 2;
	defparam lut_6114.mask = 4'b0001;

	lut_sub lut_6120 ({g13, g93}, g555);
	defparam lut_6120.LUT_SIZE = 2;
	defparam lut_6120.mask = 4'b0010;

	lut_sub lut_6126 ({g554, g555}, g556);
	defparam lut_6126.LUT_SIZE = 2;
	defparam lut_6126.mask = 4'b1000;

	lut_sub lut_6134 ({g18, g15, g13, g461}, g557);
	defparam lut_6134.LUT_SIZE = 4;
	defparam lut_6134.mask = 16'h7350;

	lut_sub lut_6147 ({g45, g556, g557}, g558);
	defparam lut_6147.LUT_SIZE = 3;
	defparam lut_6147.mask = 8'h20;

	lut_sub lut_6156 ({g109, g186, g330, g544, g558}, g559);
	defparam lut_6156.LUT_SIZE = 5;
	defparam lut_6156.mask = 32'h1f131313;

	lut_sub lut_6175 ({g13, g22}, g560);
	defparam lut_6175.LUT_SIZE = 2;
	defparam lut_6175.mask = 4'b0001;

	lut_sub lut_6181 ({g11, g461}, g561);
	defparam lut_6181.LUT_SIZE = 2;
	defparam lut_6181.mask = 4'b0001;

	lut_sub lut_6188 ({g112, g560, g561}, g562);
	defparam lut_6188.LUT_SIZE = 3;
	defparam lut_6188.mask = 8'h07;

	lut_sub lut_6198 ({i_8_, g15, g11, g108, g461}, g563);
	defparam lut_6198.LUT_SIZE = 5;
	defparam lut_6198.mask = 32'h11010101;

	lut_sub lut_6209 ({i_8_, g108, g548, g554}, g564);
	defparam lut_6209.LUT_SIZE = 4;
	defparam lut_6209.mask = 16'h0700;

	lut_sub lut_6221 ({g100, g136, g560, g562, g563, g564}, g565);
	defparam lut_6221.LUT_SIZE = 6;
	defparam lut_6221.mask = 64'h8080800080008000;

	lut_sub lut_6231 ({g13, g158}, g566);
	defparam lut_6231.LUT_SIZE = 2;
	defparam lut_6231.mask = 4'b0001;

	lut_sub lut_6240 ({g131, g251, g461, g566, g556}, g567);
	defparam lut_6240.LUT_SIZE = 5;
	defparam lut_6240.mask = 32'h00bb00bf;

	lut_sub lut_6262 ({g545, g1708, g553, g559, g565, g567}, g568);
	defparam lut_6262.LUT_SIZE = 6;
	defparam lut_6262.mask = 64'h0000000200000000;

	lut_sub lut_6268 ({g112, g566}, g569);
	defparam lut_6268.LUT_SIZE = 2;
	defparam lut_6268.mask = 4'b0001;

	lut_sub lut_6275 ({i_14_, i_12_, i_13_, g99, g101, g115}, g570);
	defparam lut_6275.LUT_SIZE = 6;
	defparam lut_6275.mask = 64'h000000000a2a2a00;

	lut_sub lut_6290 ({g45, g547, g546, g532}, g571);
	defparam lut_6290.LUT_SIZE = 4;
	defparam lut_6290.mask = 16'h0800;

	lut_sub lut_6294 ({i_14_, i_12_, i_13_}, g572);
	defparam lut_6294.LUT_SIZE = 3;
	defparam lut_6294.mask = 8'h06;

	lut_sub lut_6304 ({g13, g99, g100, g124, g572}, g573);
	defparam lut_6304.LUT_SIZE = 5;
	defparam lut_6304.mask = 32'h01010133;

	lut_sub lut_6316 ({g122, g572}, g574);
	defparam lut_6316.LUT_SIZE = 2;
	defparam lut_6316.mask = 4'b0100;

	lut_sub lut_6326 ({g101, g224, g467, g571, g573, g574}, g575);
	defparam lut_6326.LUT_SIZE = 6;
	defparam lut_6326.mask = 64'hcccccccc00080000;

	lut_sub lut_6349 ({g131, g461, g566}, g576);
	defparam lut_6349.LUT_SIZE = 3;
	defparam lut_6349.mask = 8'ha8;

	lut_sub lut_6358 ({i_8_, g88, g284, g576}, g577);
	defparam lut_6358.LUT_SIZE = 4;
	defparam lut_6358.mask = 16'h222a;

	lut_sub lut_6370 ({i_8_, g15, g119, g108, g461}, g578);
	defparam lut_6370.LUT_SIZE = 5;
	defparam lut_6370.mask = 32'h00001101;

	lut_sub lut_6379 ({i_8_, g108, g554, g550}, g579);
	defparam lut_6379.LUT_SIZE = 4;
	defparam lut_6379.mask = 16'h0007;

	lut_sub lut_6390 ({g338, g577, g556, g578, g579}, g580);
	defparam lut_6390.LUT_SIZE = 5;
	defparam lut_6390.mask = 32'h08008800;

	lut_sub lut_6401 ({g102, g112, g131, g461, g546}, g581);
	defparam lut_6401.LUT_SIZE = 5;
	defparam lut_6401.mask = 32'h00770057;

	lut_sub lut_6418 ({g151, g554, g581}, g582);
	defparam lut_6418.LUT_SIZE = 3;
	defparam lut_6418.mask = 8'ha8;

	lut_sub lut_6428 ({g45, g195, g532, g478}, g583);
	defparam lut_6428.LUT_SIZE = 4;
	defparam lut_6428.mask = 16'h8000;

	lut_sub lut_6434 ({i_11_, i_9_, g48, g214}, g584);
	defparam lut_6434.LUT_SIZE = 4;
	defparam lut_6434.mask = 16'h0040;

	lut_sub lut_6441 ({g141, g99, g171}, g585);
	defparam lut_6441.LUT_SIZE = 3;
	defparam lut_6441.mask = 8'h02;

	lut_sub lut_6449 ({i_15_, g89, g583, g584, g585}, g586);
	defparam lut_6449.LUT_SIZE = 5;
	defparam lut_6449.mask = 32'h0fff0888;

	lut_sub lut_6473 ({g569, g570, g575, g580, g582, g586}, g587);
	defparam lut_6473.LUT_SIZE = 6;
	defparam lut_6473.mask = 64'h0001000000000000;

	lut_sub lut_6479 ({i_12_, i_13_, g18, g179}, g588);
	defparam lut_6479.LUT_SIZE = 4;
	defparam lut_6479.mask = 16'haaa2;

	lut_sub lut_6495 ({g109, g330, g413, g414, g531, g588}, g589);
	defparam lut_6495.LUT_SIZE = 6;
	defparam lut_6495.mask = 64'h4000f0004000c000;

	lut_sub lut_6507 ({i_11_, i_9_, i_10_, i_15_, g461}, g590);
	defparam lut_6507.LUT_SIZE = 5;
	defparam lut_6507.mask = 32'hfbfbfbab;

	lut_sub lut_6537 ({i_11_, i_9_, i_10_, i_15_, g171}, g591);
	defparam lut_6537.LUT_SIZE = 5;
	defparam lut_6537.mask = 32'h0a028a02;

	lut_sub lut_6552 ({g204, g279, g460, g470, g591}, g592);
	defparam lut_6552.LUT_SIZE = 5;
	defparam lut_6552.mask = 32'hffff7fff;

	lut_sub lut_6589 ({g177, g560, g561}, g593);
	defparam lut_6589.LUT_SIZE = 3;
	defparam lut_6589.mask = 8'h80;

	lut_sub lut_6595 ({g464, g593}, g594);
	defparam lut_6595.LUT_SIZE = 2;
	defparam lut_6595.mask = 4'b0001;

	lut_sub lut_6605 ({g112, g136, g151, g548, g478, g594}, g595);
	defparam lut_6605.LUT_SIZE = 6;
	defparam lut_6605.mask = 64'hff40f040f040f040;

	lut_sub lut_6636 ({i_8_, g108, g177, g560, g464}, g596);
	defparam lut_6636.LUT_SIZE = 5;
	defparam lut_6636.mask = 32'h000000bf;

	lut_sub lut_6651 ({g145, g195, g532, g596, g478}, g597);
	defparam lut_6651.LUT_SIZE = 5;
	defparam lut_6651.mask = 32'hcccc8000;

	lut_sub lut_6667 ({g99, g203, g555, g474}, g598);
	defparam lut_6667.LUT_SIZE = 4;
	defparam lut_6667.mask = 16'h007f;

	lut_sub lut_6680 ({g100, g284, g470}, g599);
	defparam lut_6680.LUT_SIZE = 3;
	defparam lut_6680.mask = 8'h15;

	lut_sub lut_6690 ({i_8_, g4, g98, g279, g173}, g600);
	defparam lut_6690.LUT_SIZE = 5;
	defparam lut_6690.mask = 32'h00030005;

	lut_sub lut_6698 ({i_11_, i_9_, g236}, g601);
	defparam lut_6698.LUT_SIZE = 3;
	defparam lut_6698.mask = 8'h01;

	lut_sub lut_6706 ({g134, g149, g534, g522}, g602);
	defparam lut_6706.LUT_SIZE = 4;
	defparam lut_6706.mask = 16'h0537;

	lut_sub lut_6719 ({i_8_, g100, g199, g531}, g603);
	defparam lut_6719.LUT_SIZE = 4;
	defparam lut_6719.mask = 16'h0007;

	lut_sub lut_6731 ({g598, g599, g600, g601, g602, g603}, g604);
	defparam lut_6731.LUT_SIZE = 6;
	defparam lut_6731.mask = 64'h8000000000000000;

	lut_sub lut_6739 ({i_8_, g108, g177, g560, g464}, g605);
	defparam lut_6739.LUT_SIZE = 5;
	defparam lut_6739.mask = 32'h00bf0000;

	lut_sub lut_6754 ({g109, g195, g605, g532, g478}, g606);
	defparam lut_6754.LUT_SIZE = 5;
	defparam lut_6754.mask = 32'hf0f08000;

	lut_sub lut_6772 ({g589, g1695, g595, g597, g604, g606}, g607);
	defparam lut_6772.LUT_SIZE = 6;
	defparam lut_6772.mask = 64'h0000000000010000;

	lut_sub lut_6780 ({g136, g199, g547, g481}, g608);
	defparam lut_6780.LUT_SIZE = 4;
	defparam lut_6780.mask = 16'h00ef;

	lut_sub lut_6794 ({i_8_, g108, g135, g561, g544}, g609);
	defparam lut_6794.LUT_SIZE = 5;
	defparam lut_6794.mask = 32'h000003ab;

	lut_sub lut_6806 ({i_11_, i_15_, g141, g461}, g610);
	defparam lut_6806.LUT_SIZE = 4;
	defparam lut_6806.mask = 16'h5051;

	lut_sub lut_6818 ({g6, i_15_, g323, g186, g610}, g611);
	defparam lut_6818.LUT_SIZE = 5;
	defparam lut_6818.mask = 32'h00110511;

	lut_sub lut_6832 ({g136, g532, g495, g609, g611}, g612);
	defparam lut_6832.LUT_SIZE = 5;
	defparam lut_6832.mask = 32'h88808800;

	lut_sub lut_6842 ({g199, g547}, g613);
	defparam lut_6842.LUT_SIZE = 2;
	defparam lut_6842.mask = 4'b0100;

	lut_sub lut_6851 ({g18, g13, g195, g124, g461}, g614);
	defparam lut_6851.LUT_SIZE = 5;
	defparam lut_6851.mask = 32'ha080e0c0;

	lut_sub lut_6867 ({g177, g560, g613, g506, g614}, g615);
	defparam lut_6867.LUT_SIZE = 5;
	defparam lut_6867.mask = 32'h04000000;

	lut_sub lut_6872 ({i_11_, i_9_, i_10_, i_15_, g461}, g616);
	defparam lut_6872.LUT_SIZE = 5;
	defparam lut_6872.mask = 32'hbfafaefe;

	lut_sub lut_6901 ({i_11_, i_9_, i_10_, i_15_, g13}, g617);
	defparam lut_6901.LUT_SIZE = 5;
	defparam lut_6901.mask = 32'h00010010;

	lut_sub lut_6908 ({i_14_, i_12_, i_13_, g99, g158}, g618);
	defparam lut_6908.LUT_SIZE = 5;
	defparam lut_6908.mask = 32'h00001110;

	lut_sub lut_6916 ({i_15_, g178, g461}, g619);
	defparam lut_6916.LUT_SIZE = 3;
	defparam lut_6916.mask = 8'h01;

	lut_sub lut_6923 ({g59, g243, g619}, g620);
	defparam lut_6923.LUT_SIZE = 3;
	defparam lut_6923.mask = 8'h15;

	lut_sub lut_6931 ({g135, g576}, g621);
	defparam lut_6931.LUT_SIZE = 2;
	defparam lut_6931.mask = 4'b0010;

	lut_sub lut_6938 ({i_15_, g113, g118, g171}, g622);
	defparam lut_6938.LUT_SIZE = 4;
	defparam lut_6938.mask = 16'h0200;

	lut_sub lut_6948 ({g277, g617, g618, g620, g621, g622}, g623);
	defparam lut_6948.LUT_SIZE = 6;
	defparam lut_6948.mask = 64'h8000000080008000;

	lut_sub lut_6959 ({g108, g131, g171, g164, g461}, g624);
	defparam lut_6959.LUT_SIZE = 5;
	defparam lut_6959.mask = 32'h00003075;

	lut_sub lut_6973 ({g47, g566, g546, g555}, g625);
	defparam lut_6973.LUT_SIZE = 4;
	defparam lut_6973.mask = 16'h8000;

	lut_sub lut_6980 ({g199, g547, g481}, g626);
	defparam lut_6980.LUT_SIZE = 3;
	defparam lut_6980.mask = 8'h10;

	lut_sub lut_6987 ({g177, g560, g464}, g627);
	defparam lut_6987.LUT_SIZE = 3;
	defparam lut_6987.mask = 8'h40;

	lut_sub lut_6995 ({i_8_, g88, g108, g626, g627}, g628);
	defparam lut_6995.LUT_SIZE = 5;
	defparam lut_6995.mask = 32'h0cee0000;

	lut_sub lut_7011 ({g109, g534, g624, g625, g628}, g629);
	defparam lut_7011.LUT_SIZE = 5;
	defparam lut_7011.mask = 32'ha0a02000;

	lut_sub lut_7021 ({g171, g115}, g630);
	defparam lut_7021.LUT_SIZE = 2;
	defparam lut_7021.mask = 4'b1000;

	lut_sub lut_7029 ({g548, g550, g561, g630}, g631);
	defparam lut_7029.LUT_SIZE = 4;
	defparam lut_7029.mask = 16'h8000;

	lut_sub lut_7038 ({g134, g109, g146, g551, g631}, g632);
	defparam lut_7038.LUT_SIZE = 5;
	defparam lut_7038.mask = 32'hcfcc4444;

	lut_sub lut_7061 ({g608, g612, g1686, g623, g629, g632}, g633);
	defparam lut_7061.LUT_SIZE = 6;
	defparam lut_7061.mask = 64'h0000000100000000;

	lut_sub lut_7071 ({g527, g543, g568, g587, g607, g633}, g634);
	defparam lut_7071.LUT_SIZE = 6;
	defparam lut_7071.mask = 64'h0000000000000001;

	lut_sub lut_7079 ({g145, g268, g555, g474}, g635);
	defparam lut_7079.LUT_SIZE = 4;
	defparam lut_7079.mask = 16'h007f;

	lut_sub lut_7092 ({g47, g172, g465}, g636);
	defparam lut_7092.LUT_SIZE = 3;
	defparam lut_7092.mask = 8'h40;

	lut_sub lut_7100 ({g101, g151, g530, g636}, g637);
	defparam lut_7100.LUT_SIZE = 4;
	defparam lut_7100.mask = 16'h0a3b;

	lut_sub lut_7113 ({g279, g566, g460}, g638);
	defparam lut_7113.LUT_SIZE = 3;
	defparam lut_7113.mask = 8'h80;

	lut_sub lut_7123 ({g101, g145, g203, g555, g474, g638}, g639);
	defparam lut_7123.LUT_SIZE = 6;
	defparam lut_7123.mask = 64'hffff5555c0004000;

	lut_sub lut_7156 ({g173, g546, g477}, g640);
	defparam lut_7156.LUT_SIZE = 3;
	defparam lut_7156.mask = 8'h40;

	lut_sub lut_7162 ({g18, g171}, g641);
	defparam lut_7162.LUT_SIZE = 2;
	defparam lut_7162.mask = 4'b1000;

	lut_sub lut_7169 ({g530, g641, g531}, g642);
	defparam lut_7169.LUT_SIZE = 3;
	defparam lut_7169.mask = 8'h80;

	lut_sub lut_7177 ({g15, g102, g461, g642}, g643);
	defparam lut_7177.LUT_SIZE = 4;
	defparam lut_7177.mask = 16'h4445;

	lut_sub lut_7190 ({g145, g151, g640, g529, g643}, g644);
	defparam lut_7190.LUT_SIZE = 5;
	defparam lut_7190.mask = 32'hff010f01;

	lut_sub lut_7212 ({g151, g268, g555, g474, g644}, g645);
	defparam lut_7212.LUT_SIZE = 5;
	defparam lut_7212.mask = 32'h55554000;

	lut_sub lut_7229 ({i_8_, g88, g108, g112, g135, g284}, g646);
	defparam lut_7229.LUT_SIZE = 6;
	defparam lut_7229.mask = 64'ha0a0a0a080000000;

	lut_sub lut_7244 ({g171, g158, g646}, g647);
	defparam lut_7244.LUT_SIZE = 3;
	defparam lut_7244.mask = 8'h20;

	lut_sub lut_7250 ({i_14_, g101, g158}, g648);
	defparam lut_7250.LUT_SIZE = 3;
	defparam lut_7250.mask = 8'h01;

	lut_sub lut_7257 ({g101, g641, g630}, g649);
	defparam lut_7257.LUT_SIZE = 3;
	defparam lut_7257.mask = 8'h07;

	lut_sub lut_7266 ({i_8_, g88, g108, g534}, g650);
	defparam lut_7266.LUT_SIZE = 4;
	defparam lut_7266.mask = 16'h0015;

	lut_sub lut_7276 ({g112, g534, g530, g540}, g651);
	defparam lut_7276.LUT_SIZE = 4;
	defparam lut_7276.mask = 16'h007f;

	lut_sub lut_7291 ({i_8_, g135, g534, g530, g630, g540}, g652);
	defparam lut_7291.LUT_SIZE = 6;
	defparam lut_7291.mask = 64'h0000000000007fff;

	lut_sub lut_7314 ({g145, g530, g531, g651, g652}, g653);
	defparam lut_7314.LUT_SIZE = 5;
	defparam lut_7314.mask = 32'h88888000;

	lut_sub lut_7328 ({g45, g145, g197, g626, g467, g636}, g654);
	defparam lut_7328.LUT_SIZE = 6;
	defparam lut_7328.mask = 64'h0000feff0000ffff;

	lut_sub lut_7368 ({g647, g648, g649, g650, g653, g654}, g655);
	defparam lut_7368.LUT_SIZE = 6;
	defparam lut_7368.mask = 64'h2000000000000000;

	lut_sub lut_7376 ({i_8_, g100, g323, g338, g540}, g656);
	defparam lut_7376.LUT_SIZE = 5;
	defparam lut_7376.mask = 32'h45454555;

	lut_sub lut_7397 ({g101, g151, g534, g626, g656}, g657);
	defparam lut_7397.LUT_SIZE = 5;
	defparam lut_7397.mask = 32'haa22a020;

	lut_sub lut_7411 ({i_11_, g141, g377}, g658);
	defparam lut_7411.LUT_SIZE = 3;
	defparam lut_7411.mask = 8'h01;

	lut_sub lut_7417 ({i_11_, g5, g377}, g659);
	defparam lut_7417.LUT_SIZE = 3;
	defparam lut_7417.mask = 8'h01;

	lut_sub lut_7423 ({i_3_, i_4_, i_8_, g34, g57}, g660);
	defparam lut_7423.LUT_SIZE = 5;
	defparam lut_7423.mask = 32'h00010000;

	lut_sub lut_7430 ({i_14_, i_12_, g112, g199, g122}, g661);
	defparam lut_7430.LUT_SIZE = 5;
	defparam lut_7430.mask = 32'h03030b03;

	lut_sub lut_7448 ({g338, g658, g659, g522, g660, g661}, g662);
	defparam lut_7448.LUT_SIZE = 6;
	defparam lut_7448.mask = 64'ha0000000a8000000;

	lut_sub lut_7460 ({g146, g630, g657, g662}, g663);
	defparam lut_7460.LUT_SIZE = 4;
	defparam lut_7460.mask = 16'h1011;

	lut_sub lut_7472 ({g635, g637, g639, g645, g655, g663}, g664);
	defparam lut_7472.LUT_SIZE = 6;
	defparam lut_7472.mask = 64'h0001000000000000;

	lut_sub lut_7482 ({g73, g358, g458, g521, g634, g664}, o_4_);
	defparam lut_7482.LUT_SIZE = 6;
	defparam lut_7482.mask = 64'h00000000fffffffe;

	lut_sub lut_7521 ({g107, g130, g1782, g148, g157}, g666);
	defparam lut_7521.LUT_SIZE = 5;
	defparam lut_7521.mask = 32'h00000001;

	lut_sub lut_7530 ({g490, g1737, g499, g1728, g512}, g667);
	defparam lut_7530.LUT_SIZE = 5;
	defparam lut_7530.mask = 32'h00000001;

	lut_sub lut_7537 ({g19, g16, g145}, g668);
	defparam lut_7537.LUT_SIZE = 3;
	defparam lut_7537.mask = 8'h45;

	lut_sub lut_7545 ({g7, g93}, g669);
	defparam lut_7545.LUT_SIZE = 2;
	defparam lut_7545.mask = 4'b1101;

	lut_sub lut_7553 ({g9, g119}, g670);
	defparam lut_7553.LUT_SIZE = 2;
	defparam lut_7553.mask = 4'b0001;

	lut_sub lut_7559 ({g7, g122}, g671);
	defparam lut_7559.LUT_SIZE = 2;
	defparam lut_7559.mask = 4'b0010;

	lut_sub lut_7565 ({g9, g102}, g672);
	defparam lut_7565.LUT_SIZE = 2;
	defparam lut_7565.mask = 4'b0010;

	lut_sub lut_7572 ({i_8_, g16, g100, g672}, g673);
	defparam lut_7572.LUT_SIZE = 4;
	defparam lut_7572.mask = 16'h0031;

	lut_sub lut_7584 ({g101, g145, g669, g670, g671, g673}, g674);
	defparam lut_7584.LUT_SIZE = 6;
	defparam lut_7584.mask = 64'haaaa0080a0a00080;

	lut_sub lut_7603 ({g7, g115}, g675);
	defparam lut_7603.LUT_SIZE = 2;
	defparam lut_7603.mask = 4'b0010;

	lut_sub lut_7609 ({g7, g158}, g676);
	defparam lut_7609.LUT_SIZE = 2;
	defparam lut_7609.mask = 4'b0001;

	lut_sub lut_7615 ({g9, g131}, g677);
	defparam lut_7615.LUT_SIZE = 2;
	defparam lut_7615.mask = 4'b0001;

	lut_sub lut_7621 ({g9, g95}, g678);
	defparam lut_7621.LUT_SIZE = 2;
	defparam lut_7621.mask = 4'b1110;

	lut_sub lut_7631 ({g323, g284, g678, g677}, g679);
	defparam lut_7631.LUT_SIZE = 4;
	defparam lut_7631.mask = 16'hfa22;

	lut_sub lut_7648 ({g145, g675, g672, g676, g677, g679}, g680);
	defparam lut_7648.LUT_SIZE = 6;
	defparam lut_7648.mask = 64'h5555555540000000;

	lut_sub lut_7671 ({g19, g16, g112}, g681);
	defparam lut_7671.LUT_SIZE = 3;
	defparam lut_7671.mask = 8'h45;

	lut_sub lut_7680 ({g112, g678, g669}, g682);
	defparam lut_7680.LUT_SIZE = 3;
	defparam lut_7680.mask = 8'h0e;

	lut_sub lut_7689 ({g112, g676, g677}, g683);
	defparam lut_7689.LUT_SIZE = 3;
	defparam lut_7689.mask = 8'h07;

	lut_sub lut_7698 ({g112, g675, g672}, g684);
	defparam lut_7698.LUT_SIZE = 3;
	defparam lut_7698.mask = 8'h07;

	lut_sub lut_7707 ({i_8_, g100, g678, g677}, g685);
	defparam lut_7707.LUT_SIZE = 4;
	defparam lut_7707.mask = 16'h000d;

	lut_sub lut_7717 ({g12, g112, g323, g670}, g686);
	defparam lut_7717.LUT_SIZE = 4;
	defparam lut_7717.mask = 16'hfac0;

	lut_sub lut_7734 ({g681, g682, g683, g684, g685, g686}, g687);
	defparam lut_7734.LUT_SIZE = 6;
	defparam lut_7734.mask = 64'h4000000000000000;

	lut_sub lut_7744 ({g19, g16, g136, g151, g678, g669}, g688);
	defparam lut_7744.LUT_SIZE = 6;
	defparam lut_7744.mask = 64'hf000f1f1f000f000;

	lut_sub lut_7772 ({i_8_, g12, g135, g672}, g689);
	defparam lut_7772.LUT_SIZE = 4;
	defparam lut_7772.mask = 16'h0013;

	lut_sub lut_7781 ({i_8_, g135, g669, g676}, g690);
	defparam lut_7781.LUT_SIZE = 4;
	defparam lut_7781.mask = 16'h000d;

	lut_sub lut_7790 ({i_8_, g135, g678, g670}, g691);
	defparam lut_7790.LUT_SIZE = 4;
	defparam lut_7790.mask = 16'h000d;

	lut_sub lut_7801 ({i_8_, g12, g88, g108, g675, g676}, g692);
	defparam lut_7801.LUT_SIZE = 6;
	defparam lut_7801.mask = 64'h0000000000770fff;

	lut_sub lut_7828 ({g151, g670, g689, g690, g691, g692}, g693);
	defparam lut_7828.LUT_SIZE = 6;
	defparam lut_7828.mask = 64'h8000800080000000;

	lut_sub lut_7840 ({g668, g674, g680, g687, g688, g693}, g694);
	defparam lut_7840.LUT_SIZE = 6;
	defparam lut_7840.mask = 64'h0000000100000000;

	lut_sub lut_7846 ({g8, g145}, g695);
	defparam lut_7846.LUT_SIZE = 2;
	defparam lut_7846.mask = 4'b0100;

	lut_sub lut_7852 ({g9, g104}, g696);
	defparam lut_7852.LUT_SIZE = 2;
	defparam lut_7852.mask = 4'b1110;

	lut_sub lut_7862 ({g112, g136, g151, g696}, g697);
	defparam lut_7862.LUT_SIZE = 4;
	defparam lut_7862.mask = 16'h2aaa;

	lut_sub lut_7878 ({g8, g10, g112, g323, g696, g670}, g698);
	defparam lut_7878.LUT_SIZE = 6;
	defparam lut_7878.mask = 64'hf200f000f2f2f000;

	lut_sub lut_7910 ({g10, g12, g101, g145, g696, g698}, g699);
	defparam lut_7910.LUT_SIZE = 6;
	defparam lut_7910.mask = 64'h5111510051005100;

	lut_sub lut_7932 ({g8, g10, g23, g136, g151}, g700);
	defparam lut_7932.LUT_SIZE = 5;
	defparam lut_7932.mask = 32'h8888fc88;

	lut_sub lut_7951 ({g695, g697, g699, g700}, g701);
	defparam lut_7951.LUT_SIZE = 4;
	defparam lut_7951.mask = 16'h1000;

	lut_sub lut_7957 ({g9, g124}, g702);
	defparam lut_7957.LUT_SIZE = 2;
	defparam lut_7957.mask = 4'b0001;

	lut_sub lut_7963 ({g9, g22}, g703);
	defparam lut_7963.LUT_SIZE = 2;
	defparam lut_7963.mask = 4'b0001;

	lut_sub lut_7969 ({g9, g122}, g704);
	defparam lut_7969.LUT_SIZE = 2;
	defparam lut_7969.mask = 4'b0010;

	lut_sub lut_7977 ({g46, g118, g702, g704}, g705);
	defparam lut_7977.LUT_SIZE = 4;
	defparam lut_7977.mask = 16'h070f;

	lut_sub lut_7989 ({g9, g115}, g706);
	defparam lut_7989.LUT_SIZE = 2;
	defparam lut_7989.mask = 4'b0010;

	lut_sub lut_7995 ({g477, g703}, g707);
	defparam lut_7995.LUT_SIZE = 2;
	defparam lut_7995.mask = 4'b0010;

	lut_sub lut_8004 ({i_8_, g108, g464, g696, g706, g707}, g708);
	defparam lut_8004.LUT_SIZE = 6;
	defparam lut_8004.mask = 64'h0000fff30000ffbb;

	lut_sub lut_8040 ({g109, g702, g703, g705, g708}, g709);
	defparam lut_8040.LUT_SIZE = 5;
	defparam lut_8040.mask = 32'h88888000;

	lut_sub lut_8050 ({g9, g158}, g710);
	defparam lut_8050.LUT_SIZE = 2;
	defparam lut_8050.mask = 4'b0001;

	lut_sub lut_8054 ({i_14_, i_12_}, g711);
	defparam lut_8054.LUT_SIZE = 2;
	defparam lut_8054.mask = 4'b0100;

	lut_sub lut_8062 ({g7, i_8_, g115, g122, g711}, g712);
	defparam lut_8062.LUT_SIZE = 5;
	defparam lut_8062.mask = 32'h0054f0fc;

	lut_sub lut_8081 ({g6, i_15_, g7, g461}, g713);
	defparam lut_8081.LUT_SIZE = 4;
	defparam lut_8081.mask = 16'h0007;

	lut_sub lut_8092 ({g4, g98, g92, g712, g713}, g714);
	defparam lut_8092.LUT_SIZE = 5;
	defparam lut_8092.mask = 32'h000000f7;

	lut_sub lut_8106 ({g251, g281, g710, g714}, g715);
	defparam lut_8106.LUT_SIZE = 4;
	defparam lut_8106.mask = 16'haa08;

	lut_sub lut_8117 ({i_8_, g99, g108, g467}, g716);
	defparam lut_8117.LUT_SIZE = 4;
	defparam lut_8117.mask = 16'h0a2a;

	lut_sub lut_8129 ({g19, g99, g115, g711}, g717);
	defparam lut_8129.LUT_SIZE = 4;
	defparam lut_8129.mask = 16'h040f;

	lut_sub lut_8140 ({i_8_, g46, g88, g704}, g718);
	defparam lut_8140.LUT_SIZE = 4;
	defparam lut_8140.mask = 16'h1300;

	lut_sub lut_8149 ({i_8_, g100, g474, g460}, g719);
	defparam lut_8149.LUT_SIZE = 4;
	defparam lut_8149.mask = 16'h0007;

	lut_sub lut_8161 ({g112, g186, g120, g477, g474, g671}, g720);
	defparam lut_8161.LUT_SIZE = 6;
	defparam lut_8161.mask = 64'hffff0c0c00aa0008;

	lut_sub lut_8194 ({g716, g717, g718, g719, g720}, g721);
	defparam lut_8194.LUT_SIZE = 5;
	defparam lut_8194.mask = 32'h40000000;

	lut_sub lut_8201 ({g44, g118, g186}, g722);
	defparam lut_8201.LUT_SIZE = 3;
	defparam lut_8201.mask = 8'h07;

	lut_sub lut_8210 ({g44, g108, g710}, g723);
	defparam lut_8210.LUT_SIZE = 3;
	defparam lut_8210.mask = 8'h13;

	lut_sub lut_8219 ({g7, g158, g711}, g724);
	defparam lut_8219.LUT_SIZE = 3;
	defparam lut_8219.mask = 8'h13;

	lut_sub lut_8229 ({g99, g724, g677, g710}, g725);
	defparam lut_8229.LUT_SIZE = 4;
	defparam lut_8229.mask = 16'h007f;

	lut_sub lut_8241 ({g7, g711}, g726);
	defparam lut_8241.LUT_SIZE = 2;
	defparam lut_8241.mask = 4'b1000;

	lut_sub lut_8246 ({g6, i_15_, i_14_, i_12_, i_13_}, g727);
	defparam lut_8246.LUT_SIZE = 5;
	defparam lut_8246.mask = 32'h000000b0;

	lut_sub lut_8256 ({g18, g59, g726, g727}, g728);
	defparam lut_8256.LUT_SIZE = 4;
	defparam lut_8256.mask = 16'h0d05;

	lut_sub lut_8267 ({i_14_, i_12_, i_13_, g59, g99, g93}, g729);
	defparam lut_8267.LUT_SIZE = 6;
	defparam lut_8267.mask = 64'h2a222a2a00000000;

	lut_sub lut_8286 ({g722, g723, g725, g728, g729}, g730);
	defparam lut_8286.LUT_SIZE = 5;
	defparam lut_8286.mask = 32'h80000000;

	lut_sub lut_8294 ({g44, g46, g99, g678}, g731);
	defparam lut_8294.LUT_SIZE = 4;
	defparam lut_8294.mask = 16'h2333;

	lut_sub lut_8308 ({g99, g477, g474, g460}, g732);
	defparam lut_8308.LUT_SIZE = 4;
	defparam lut_8308.mask = 16'h00f7;

	lut_sub lut_8322 ({g99, g702, g706, g703}, g733);
	defparam lut_8322.LUT_SIZE = 4;
	defparam lut_8322.mask = 16'h007f;

	lut_sub lut_8334 ({g7, g124}, g734);
	defparam lut_8334.LUT_SIZE = 2;
	defparam lut_8334.mask = 4'b0001;

	lut_sub lut_8342 ({g134, g478, g734, g702}, g735);
	defparam lut_8342.LUT_SIZE = 4;
	defparam lut_8342.mask = 16'h007f;

	lut_sub lut_8355 ({i_8_, i_6_, i_7_, g98, g478, g704}, g736);
	defparam lut_8355.LUT_SIZE = 6;
	defparam lut_8355.mask = 64'h0007000700030005;

	lut_sub lut_8373 ({g731, g732, g733, g735, g736}, g737);
	defparam lut_8373.LUT_SIZE = 5;
	defparam lut_8373.mask = 32'h80000000;

	lut_sub lut_8378 ({i_11_, i_9_, i_10_, i_15_, g7}, g738);
	defparam lut_8378.LUT_SIZE = 5;
	defparam lut_8378.mask = 32'h01100100;

	lut_sub lut_8389 ({g23, g96, g734, g669, g738}, g739);
	defparam lut_8389.LUT_SIZE = 5;
	defparam lut_8389.mask = 32'h00200000;

	lut_sub lut_8397 ({g46, g90, g704, g739}, g740);
	defparam lut_8397.LUT_SIZE = 4;
	defparam lut_8397.mask = 16'h0400;

	lut_sub lut_8406 ({g243, g251, g460, g724, g740}, g741);
	defparam lut_8406.LUT_SIZE = 5;
	defparam lut_8406.mask = 32'hffc05540;

	lut_sub lut_8429 ({g715, g721, g730, g737, g741}, g742);
	defparam lut_8429.LUT_SIZE = 5;
	defparam lut_8429.mask = 32'h00000001;

	lut_sub lut_8438 ({g7, g9, g22, g100, g277}, g743);
	defparam lut_8438.LUT_SIZE = 5;
	defparam lut_8438.mask = 32'h000a030b;

	lut_sub lut_8451 ({i_14_, i_12_, i_13_, g101, g145, g93}, g744);
	defparam lut_8451.LUT_SIZE = 6;
	defparam lut_8451.mask = 64'h0a000a0a00220000;

	lut_sub lut_8467 ({i_8_, g18, g4, g98, g122, g726}, g745);
	defparam lut_8467.LUT_SIZE = 6;
	defparam lut_8467.mask = 64'h00080008000a0000;

	lut_sub lut_8475 ({i_6_, g87}, g746);
	defparam lut_8475.LUT_SIZE = 2;
	defparam lut_8475.mask = 4'b0100;

	lut_sub lut_8484 ({i_8_, g134, g135, g746, g671, g704}, g747);
	defparam lut_8484.LUT_SIZE = 6;
	defparam lut_8484.mask = 64'h0303575703335777;

	lut_sub lut_8524 ({g145, g135, g460, g710, g745, g747}, g748);
	defparam lut_8524.LUT_SIZE = 6;
	defparam lut_8524.mask = 64'h8888808088008000;

	lut_sub lut_8538 ({i_11_, i_9_, i_10_, i_15_, g9, g660}, g749);
	defparam lut_8538.LUT_SIZE = 6;
	defparam lut_8538.mask = 64'h0000000000030100;

	lut_sub lut_8549 ({g134, g251, g660, g704, g749}, g750);
	defparam lut_8549.LUT_SIZE = 5;
	defparam lut_8549.mask = 32'h01555555;

	lut_sub lut_8569 ({i_8_, g10, g4, g46, g98}, g751);
	defparam lut_8569.LUT_SIZE = 5;
	defparam lut_8569.mask = 32'h00050101;

	lut_sub lut_8580 ({g186, g423, g702, g703}, g752);
	defparam lut_8580.LUT_SIZE = 4;
	defparam lut_8580.mask = 16'h0357;

	lut_sub lut_8592 ({g481, g702}, g753);
	defparam lut_8592.LUT_SIZE = 2;
	defparam lut_8592.mask = 4'b0010;

	lut_sub lut_8601 ({i_8_, g88, g108, g467, g465, g753}, g754);
	defparam lut_8601.LUT_SIZE = 6;
	defparam lut_8601.mask = 64'h00f0aafa0000fefe;

	lut_sub lut_8637 ({g186, g677, g751, g752, g754}, g755);
	defparam lut_8637.LUT_SIZE = 5;
	defparam lut_8637.mask = 32'h80808000;

	lut_sub lut_8645 ({g9, g93}, g756);
	defparam lut_8645.LUT_SIZE = 2;
	defparam lut_8645.mask = 4'b0010;

	lut_sub lut_8655 ({g44, g46, g109, g330, g215, g756}, g757);
	defparam lut_8655.LUT_SIZE = 6;
	defparam lut_8655.mask = 64'habaa0b000b0a0b00;

	lut_sub lut_8684 ({g743, g744, g748, g750, g755, g757}, g758);
	defparam lut_8684.LUT_SIZE = 6;
	defparam lut_8684.mask = 64'h0010000000000000;

	lut_sub lut_8694 ({g411, g694, g701, g709, g742, g758}, g759);
	defparam lut_8694.LUT_SIZE = 6;
	defparam lut_8694.mask = 64'h0000000000000001;

	lut_sub lut_8701 ({i_8_, g135, g481, g704}, g760);
	defparam lut_8701.LUT_SIZE = 4;
	defparam lut_8701.mask = 16'h000d;

	lut_sub lut_8710 ({i_8_, g108, g702, g756}, g761);
	defparam lut_8710.LUT_SIZE = 4;
	defparam lut_8710.mask = 16'h0007;

	lut_sub lut_8719 ({i_8_, g135, g706, g703}, g762);
	defparam lut_8719.LUT_SIZE = 4;
	defparam lut_8719.mask = 16'h0007;

	lut_sub lut_8729 ({i_8_, g100, g481, g467, g478}, g763);
	defparam lut_8729.LUT_SIZE = 5;
	defparam lut_8729.mask = 32'h000000fd;

	lut_sub lut_8745 ({g284, g724, g760, g761, g762, g763}, g764);
	defparam lut_8745.LUT_SIZE = 6;
	defparam lut_8745.mask = 64'h8000800080000000;

	lut_sub lut_8757 ({g46, g151, g284, g706, g756, g710}, g765);
	defparam lut_8757.LUT_SIZE = 6;
	defparam lut_8757.mask = 64'hffaa8080ffaa0000;

	lut_sub lut_8792 ({g46, g101, g145, g136, g323, g702}, g766);
	defparam lut_8792.LUT_SIZE = 6;
	defparam lut_8792.mask = 64'heaeaaaaaea00aa00;

	lut_sub lut_8825 ({i_8_, g100, g477, g706}, g767);
	defparam lut_8825.LUT_SIZE = 4;
	defparam lut_8825.mask = 16'h000d;

	lut_sub lut_8835 ({g112, g702, g706, g703}, g768);
	defparam lut_8835.LUT_SIZE = 4;
	defparam lut_8835.mask = 16'h007f;

	lut_sub lut_8849 ({g112, g481, g704, g710}, g769);
	defparam lut_8849.LUT_SIZE = 4;
	defparam lut_8849.mask = 16'h00f7;

	lut_sub lut_8862 ({i_8_, g100, g703, g710}, g770);
	defparam lut_8862.LUT_SIZE = 4;
	defparam lut_8862.mask = 16'h0007;

	lut_sub lut_8873 ({i_8_, g44, g100, g323, g703, g756}, g771);
	defparam lut_8873.LUT_SIZE = 6;
	defparam lut_8873.mask = 64'hf8f8f0f0f8a8f000;

	lut_sub lut_8911 ({g767, g768, g769, g770, g771}, g772);
	defparam lut_8911.LUT_SIZE = 5;
	defparam lut_8911.mask = 32'h40000000;

	lut_sub lut_8919 ({g764, g765, g766, g772}, g773);
	defparam lut_8919.LUT_SIZE = 4;
	defparam lut_8919.mask = 16'h0001;

	lut_sub lut_8926 ({g8, g10, g118}, g774);
	defparam lut_8926.LUT_SIZE = 3;
	defparam lut_8926.mask = 8'h51;

	lut_sub lut_8935 ({i_8_, g19, g23, g108}, g775);
	defparam lut_8935.LUT_SIZE = 4;
	defparam lut_8935.mask = 16'h0511;

	lut_sub lut_8946 ({i_9_, g53, g9, g119, g214}, g776);
	defparam lut_8946.LUT_SIZE = 5;
	defparam lut_8946.mask = 32'h01010105;

	lut_sub lut_8957 ({i_8_, g88, g423, g696}, g777);
	defparam lut_8957.LUT_SIZE = 4;
	defparam lut_8957.mask = 16'h2a22;

	lut_sub lut_8971 ({g429, g678, g774, g775, g776, g777}, g778);
	defparam lut_8971.LUT_SIZE = 6;
	defparam lut_8971.mask = 64'h8000800000008000;

	lut_sub lut_8981 ({g134, g696, g675, g672}, g779);
	defparam lut_8981.LUT_SIZE = 4;
	defparam lut_8981.mask = 16'h00f7;

	lut_sub lut_8997 ({g19, g16, g89, g678, g669, g779}, g780);
	defparam lut_8997.LUT_SIZE = 6;
	defparam lut_8997.mask = 64'h00aa02aa00aa00aa;

	lut_sub lut_9020 ({g19, g16, g134}, g781);
	defparam lut_9020.LUT_SIZE = 3;
	defparam lut_9020.mask = 8'h45;

	lut_sub lut_9029 ({g118, g670, g671}, g782);
	defparam lut_9029.LUT_SIZE = 3;
	defparam lut_9029.mask = 8'h07;

	lut_sub lut_9038 ({g134, g670, g671}, g783);
	defparam lut_9038.LUT_SIZE = 3;
	defparam lut_9038.mask = 8'h07;

	lut_sub lut_9047 ({g8, i_8_, g88, g675}, g784);
	defparam lut_9047.LUT_SIZE = 4;
	defparam lut_9047.mask = 16'h3010;

	lut_sub lut_9058 ({g8, i_8_, g108, g678, g670, g671}, g785);
	defparam lut_9058.LUT_SIZE = 6;
	defparam lut_9058.mask = 64'h00ff000000f70000;

	lut_sub lut_9081 ({g781, g782, g783, g784, g785}, g786);
	defparam lut_9081.LUT_SIZE = 5;
	defparam lut_9081.mask = 32'h80000000;

	lut_sub lut_9088 ({g10, g12, g134}, g787);
	defparam lut_9088.LUT_SIZE = 3;
	defparam lut_9088.mask = 8'h15;

	lut_sub lut_9097 ({g12, g16, g99}, g788);
	defparam lut_9097.LUT_SIZE = 3;
	defparam lut_9097.mask = 8'h45;

	lut_sub lut_9106 ({g23, g88, g734}, g789);
	defparam lut_9106.LUT_SIZE = 3;
	defparam lut_9106.mask = 8'h13;

	lut_sub lut_9115 ({g23, g112, g734}, g790);
	defparam lut_9115.LUT_SIZE = 3;
	defparam lut_9115.mask = 8'h13;

	lut_sub lut_9124 ({i_8_, g108, g734, g669}, g791);
	defparam lut_9124.LUT_SIZE = 4;
	defparam lut_9124.mask = 16'h0b03;

	lut_sub lut_9135 ({i_8_, g135, g734, g675}, g792);
	defparam lut_9135.LUT_SIZE = 4;
	defparam lut_9135.mask = 16'h0007;

	lut_sub lut_9147 ({g787, g788, g789, g790, g791, g792}, g793);
	defparam lut_9147.LUT_SIZE = 6;
	defparam lut_9147.mask = 64'h8000000000000000;

	lut_sub lut_9155 ({g99, g696, g670, g672}, g794);
	defparam lut_9155.LUT_SIZE = 4;
	defparam lut_9155.mask = 16'h00f7;

	lut_sub lut_9169 ({g10, g16, g59, g678}, g795);
	defparam lut_9169.LUT_SIZE = 4;
	defparam lut_9169.mask = 16'h3233;

	lut_sub lut_9183 ({g8, g23, g134, g669}, g796);
	defparam lut_9183.LUT_SIZE = 4;
	defparam lut_9183.mask = 16'h3323;

	lut_sub lut_9195 ({i_9_, g53, g9}, g797);
	defparam lut_9195.LUT_SIZE = 3;
	defparam lut_9195.mask = 8'h10;

	lut_sub lut_9203 ({g12, g118, g696, g797}, g798);
	defparam lut_9203.LUT_SIZE = 4;
	defparam lut_9203.mask = 16'h0d0f;

	lut_sub lut_9215 ({i_11_, i_9_, i_10_, i_15_, g7, g118}, g799);
	defparam lut_9215.LUT_SIZE = 6;
	defparam lut_9215.mask = 64'h0001000101010001;

	lut_sub lut_9228 ({g794, g795, g796, g798, g799}, g800);
	defparam lut_9228.LUT_SIZE = 5;
	defparam lut_9228.mask = 32'h80000000;

	lut_sub lut_9234 ({g676, g677}, g801);
	defparam lut_9234.LUT_SIZE = 2;
	defparam lut_9234.mask = 4'b1000;

	lut_sub lut_9244 ({g23, g12, g109, g675, g672, g801}, g802);
	defparam lut_9244.LUT_SIZE = 6;
	defparam lut_9244.mask = 64'h00bf00ff00ff00ff;

	lut_sub lut_9284 ({g778, g780, g786, g793, g800, g802}, g803);
	defparam lut_9284.LUT_SIZE = 6;
	defparam lut_9284.mask = 64'h0000000000000002;

	lut_sub lut_9292 ({g21, g112, g127, g506}, g804);
	defparam lut_9292.LUT_SIZE = 4;
	defparam lut_9292.mask = 16'h0d0f;

	lut_sub lut_9304 ({g20, g59}, g805);
	defparam lut_9304.LUT_SIZE = 2;
	defparam lut_9304.mask = 4'b0100;

	lut_sub lut_9310 ({g18, g711}, g806);
	defparam lut_9310.LUT_SIZE = 2;
	defparam lut_9310.mask = 4'b0100;

	lut_sub lut_9316 ({g20, g806}, g807);
	defparam lut_9316.LUT_SIZE = 2;
	defparam lut_9316.mask = 4'b0010;

	lut_sub lut_9323 ({i_8_, g20, g21, g135}, g808);
	defparam lut_9323.LUT_SIZE = 4;
	defparam lut_9323.mask = 16'h5051;

	lut_sub lut_9335 ({g20, g16, g118, g423}, g809);
	defparam lut_9335.LUT_SIZE = 4;
	defparam lut_9335.mask = 16'h7350;

	lut_sub lut_9350 ({g136, g127, g506, g808, g809}, g810);
	defparam lut_9350.LUT_SIZE = 5;
	defparam lut_9350.mask = 32'h88880080;

	lut_sub lut_9359 ({g6, i_15_, i_14_, i_12_, i_13_}, g811);
	defparam lut_9359.LUT_SIZE = 5;
	defparam lut_9359.mask = 32'h00000c10;

	lut_sub lut_9369 ({g186, g122, g280, g711}, g812);
	defparam lut_9369.LUT_SIZE = 4;
	defparam lut_9369.mask = 16'h0073;

	lut_sub lut_9378 ({i_14_, i_12_, g95}, g813);
	defparam lut_9378.LUT_SIZE = 3;
	defparam lut_9378.mask = 8'h04;

	lut_sub lut_9387 ({g297, g270, g243, g813, g495}, g814);
	defparam lut_9387.LUT_SIZE = 5;
	defparam lut_9387.mask = 32'he0eea0aa;

	lut_sub lut_9411 ({g101, g109, g811, g676, g812, g814}, g815);
	defparam lut_9411.LUT_SIZE = 6;
	defparam lut_9411.mask = 64'h4444440040404000;

	lut_sub lut_9429 ({g804, g805, g1673, g810, g1666, g815}, g816);
	defparam lut_9429.LUT_SIZE = 6;
	defparam lut_9429.mask = 64'h0001000000000000;

	lut_sub lut_9434 ({g6, i_15_, i_14_, i_12_, i_13_}, g817);
	defparam lut_9434.LUT_SIZE = 5;
	defparam lut_9434.mask = 32'h00000830;

	lut_sub lut_9443 ({g304, g94, g475}, g818);
	defparam lut_9443.LUT_SIZE = 3;
	defparam lut_9443.mask = 8'h40;

	lut_sub lut_9451 ({i_8_, g10, g108, g158, g572}, g819);
	defparam lut_9451.LUT_SIZE = 5;
	defparam lut_9451.mask = 32'h0101000f;

	lut_sub lut_9465 ({g216, g423, g817, g818, g819}, g820);
	defparam lut_9465.LUT_SIZE = 5;
	defparam lut_9465.mask = 32'haa20aa00;

	lut_sub lut_9483 ({g301, g1768, g306, g313, g321, g820}, g821);
	defparam lut_9483.LUT_SIZE = 6;
	defparam lut_9483.mask = 64'h0000000000000001;

	lut_sub lut_9489 ({i_14_, i_12_, g18, g119}, g822);
	defparam lut_9489.LUT_SIZE = 4;
	defparam lut_9489.mask = 16'h0c50;

	lut_sub lut_9501 ({g270, g204, g817, g724, g822}, g823);
	defparam lut_9501.LUT_SIZE = 5;
	defparam lut_9501.mask = 32'h00000080;

	lut_sub lut_9510 ({g246, g421, g517, g678, g823}, g824);
	defparam lut_9510.LUT_SIZE = 5;
	defparam lut_9510.mask = 32'h00010000;

	lut_sub lut_9516 ({g134, g824}, g825);
	defparam lut_9516.LUT_SIZE = 2;
	defparam lut_9516.mask = 4'b0010;

	lut_sub lut_9523 ({g464, g478, g487}, g826);
	defparam lut_9523.LUT_SIZE = 3;
	defparam lut_9523.mask = 8'h08;

	lut_sub lut_9530 ({g264, g115, g711}, g827);
	defparam lut_9530.LUT_SIZE = 3;
	defparam lut_9530.mask = 8'hb0;

	lut_sub lut_9539 ({i_8_, g124, g572, g672}, g828);
	defparam lut_9539.LUT_SIZE = 4;
	defparam lut_9539.mask = 16'h0355;

	lut_sub lut_9552 ({g243, g423, g827, g828}, g829);
	defparam lut_9552.LUT_SIZE = 4;
	defparam lut_9552.mask = 16'h0c5d;

	lut_sub lut_9567 ({g113, g326, g88, g826, g829}, g830);
	defparam lut_9567.LUT_SIZE = 5;
	defparam lut_9567.mask = 32'ha2a2a2a0;

	lut_sub lut_9585 ({g135, g195, g412, g677}, g831);
	defparam lut_9585.LUT_SIZE = 4;
	defparam lut_9585.mask = 16'h00df;

	lut_sub lut_9601 ({g6, g141, g326, g59, g89, g831}, g832);
	defparam lut_9601.LUT_SIZE = 6;
	defparam lut_9601.mask = 64'haaaaaa22aa20aa20;

	lut_sub lut_9633 ({i_8_, g10, g16, g108, g574, g678}, g833);
	defparam lut_9633.LUT_SIZE = 6;
	defparam lut_9633.mask = 64'h0f030f0f0b0b0b0b;

	lut_sub lut_9666 ({g145, g339, g465, g833}, g834);
	defparam lut_9666.LUT_SIZE = 4;
	defparam lut_9666.mask = 16'haa20;

	lut_sub lut_9677 ({g216, g122, g711}, g835);
	defparam lut_9677.LUT_SIZE = 3;
	defparam lut_9677.mask = 8'hb0;

	lut_sub lut_9687 ({i_14_, i_12_, g100, g108, g131, g734}, g836);
	defparam lut_9687.LUT_SIZE = 6;
	defparam lut_9687.mask = 64'h0055005500550357;

	lut_sub lut_9712 ({g297, g124, g711}, g837);
	defparam lut_9712.LUT_SIZE = 3;
	defparam lut_9712.mask = 8'he0;

	lut_sub lut_9721 ({g21, g22, g711}, g838);
	defparam lut_9721.LUT_SIZE = 3;
	defparam lut_9721.mask = 8'he0;

	lut_sub lut_9732 ({g99, g323, g423, g837, g838}, g839);
	defparam lut_9732.LUT_SIZE = 5;
	defparam lut_9732.mask = 32'hf1111111;

	lut_sub lut_9751 ({g21, g118, g835, g836, g839}, g840);
	defparam lut_9751.LUT_SIZE = 5;
	defparam lut_9751.mask = 32'h44044400;

	lut_sub lut_9765 ({g825, g1653, g830, g832, g834, g840}, g841);
	defparam lut_9765.LUT_SIZE = 6;
	defparam lut_9765.mask = 64'h0000000100000000;

	lut_sub lut_9775 ({g457, g773, g803, g816, g821, g841}, g842);
	defparam lut_9775.LUT_SIZE = 6;
	defparam lut_9775.mask = 64'h0000000000000001;

	lut_sub lut_9783 ({g136, g462, g817, g818}, g843);
	defparam lut_9783.LUT_SIZE = 4;
	defparam lut_9783.mask = 16'h00fb;

	lut_sub lut_9798 ({i_8_, g21, g22, g100, g711, g837}, g844);
	defparam lut_9798.LUT_SIZE = 6;
	defparam lut_9798.mask = 64'h5544554455445040;

	lut_sub lut_9828 ({g101, g136, g216, g123, g485, g844}, g845);
	defparam lut_9828.LUT_SIZE = 6;
	defparam lut_9828.mask = 64'hffffc00055554000;

	lut_sub lut_9864 ({g14, g112, g323, g835, g807, g827}, g846);
	defparam lut_9864.LUT_SIZE = 6;
	defparam lut_9864.mask = 64'hff011101ff010000;

	lut_sub lut_9892 ({g145, g151, g811, g846}, g847);
	defparam lut_9892.LUT_SIZE = 4;
	defparam lut_9892.mask = 16'h5444;

	lut_sub lut_9903 ({g316, g158, g711}, g848);
	defparam lut_9903.LUT_SIZE = 3;
	defparam lut_9903.mask = 8'he0;

	lut_sub lut_9912 ({i_8_, g88, g813, g475}, g849);
	defparam lut_9912.LUT_SIZE = 4;
	defparam lut_9912.mask = 16'h000b;

	lut_sub lut_9921 ({g323, g817, g818}, g850);
	defparam lut_9921.LUT_SIZE = 3;
	defparam lut_9921.mask = 8'h0b;

	lut_sub lut_9932 ({g101, g145, g848, g849, g850}, g851);
	defparam lut_9932.LUT_SIZE = 5;
	defparam lut_9932.mask = 32'h88080808;

	lut_sub lut_9944 ({g843, g845, g847, g851}, g852);
	defparam lut_9944.LUT_SIZE = 4;
	defparam lut_9944.mask = 16'h0100;

	lut_sub lut_9954 ({g235, g274, g358, g374, g398, g852}, g853);
	defparam lut_9954.LUT_SIZE = 6;
	defparam lut_9954.mask = 64'h0000000000000001;

	lut_sub lut_9964 ({g73, g666, g667, g759, g842, g853}, g854);
	defparam lut_9964.LUT_SIZE = 6;
	defparam lut_9964.mask = 64'hffffffff00000001;

	lut_sub lut_10001 ({i_5_, i_3_, i_4_, g29}, g855);
	defparam lut_10001.LUT_SIZE = 4;
	defparam lut_10001.mask = 16'h4000;

	lut_sub lut_10010 ({g2, g36, g73, g111, g855}, o_7_);
	defparam lut_10010.LUT_SIZE = 5;
	defparam lut_10010.mask = 32'h0f050f07;

	lut_sub lut_10032 ({g10, g16, g134, g109, g678, g801}, g857);
	defparam lut_10032.LUT_SIZE = 6;
	defparam lut_10032.mask = 64'hf010ff11f010f010;

	lut_sub lut_10064 ({g251, g672, g803, g857}, g858);
	defparam lut_10064.LUT_SIZE = 4;
	defparam lut_10064.mask = 16'h1110;

	lut_sub lut_10074 ({g145, g151, g142, g103}, g859);
	defparam lut_10074.LUT_SIZE = 4;
	defparam lut_10074.mask = 16'hf454;

	lut_sub lut_10090 ({g764, g765, g766, g772, g859}, g860);
	defparam lut_10090.LUT_SIZE = 5;
	defparam lut_10090.mask = 32'h00000001;

	lut_sub lut_10098 ({i_8_, g88, g108, g678, g672}, g861);
	defparam lut_10098.LUT_SIZE = 5;
	defparam lut_10098.mask = 32'h00000c5d;

	lut_sub lut_10113 ({g136, g186, g677, g826, g861}, g862);
	defparam lut_10113.LUT_SIZE = 5;
	defparam lut_10113.mask = 32'haa22a020;

	lut_sub lut_10128 ({i_8_, g108, g481, g465}, g863);
	defparam lut_10128.LUT_SIZE = 4;
	defparam lut_10128.mask = 16'h0c0e;

	lut_sub lut_10140 ({i_8_, g100, g124, g158, g726}, g864);
	defparam lut_10140.LUT_SIZE = 5;
	defparam lut_10140.mask = 32'h000a002a;

	lut_sub lut_10153 ({g10, g145, g136, g127, g864}, g865);
	defparam lut_10153.LUT_SIZE = 5;
	defparam lut_10153.mask = 32'ha2a2a200;

	lut_sub lut_10168 ({i_8_, g30, g5, g40}, g866);
	defparam lut_10168.LUT_SIZE = 4;
	defparam lut_10168.mask = 16'h0105;

	lut_sub lut_10179 ({i_8_, g100, g120, g746, g103, g866}, g867);
	defparam lut_10179.LUT_SIZE = 6;
	defparam lut_10179.mask = 64'ha0aaa0aaa0aa0022;

	lut_sub lut_10208 ({g59, g112, g135, g96, g462, g867}, g868);
	defparam lut_10208.LUT_SIZE = 6;
	defparam lut_10208.mask = 64'h5511010105010101;

	lut_sub lut_10226 ({i_11_, i_9_, i_10_, i_15_, g91, g711}, g869);
	defparam lut_10226.LUT_SIZE = 6;
	defparam lut_10226.mask = 64'h00050c050c0c0005;

	lut_sub lut_10245 ({g16, g243, g619, g869}, g870);
	defparam lut_10245.LUT_SIZE = 4;
	defparam lut_10245.mask = 16'h0f07;

	lut_sub lut_10260 ({g251, g132, g122, g711, g870}, g871);
	defparam lut_10260.LUT_SIZE = 5;
	defparam lut_10260.mask = 32'haaaa008a;

	lut_sub lut_10280 ({g99, g132, g863, g865, g868, g871}, g872);
	defparam lut_10280.LUT_SIZE = 6;
	defparam lut_10280.mask = 64'h0100010000000100;

	lut_sub lut_10290 ({g82, g860, g862, g872}, g873);
	defparam lut_10290.LUT_SIZE = 4;
	defparam lut_10290.mask = 16'h0001;

	lut_sub lut_10300 ({g73, g169, g521, g759, g858, g873}, g874);
	defparam lut_10300.LUT_SIZE = 6;
	defparam lut_10300.mask = 64'hffffffff00000001;

	lut_sub lut_10337 ({i_15_, g7}, g875);
	defparam lut_10337.LUT_SIZE = 2;
	defparam lut_10337.mask = 4'b0100;

	lut_sub lut_10342 ({i_11_, i_9_, i_10_, g875}, g876);
	defparam lut_10342.LUT_SIZE = 4;
	defparam lut_10342.mask = 16'h1440;

	lut_sub lut_10349 ({i_11_, i_9_, i_10_, g875}, g877);
	defparam lut_10349.LUT_SIZE = 4;
	defparam lut_10349.mask = 16'h4010;

	lut_sub lut_10358 ({g99, g251, g285, g877}, g878);
	defparam lut_10358.LUT_SIZE = 4;
	defparam lut_10358.mask = 16'h4555;

	lut_sub lut_10372 ({g212, g568, g876, g878}, g879);
	defparam lut_10372.LUT_SIZE = 4;
	defparam lut_10372.mask = 16'h080a;

	lut_sub lut_10381 ({g569, g580, g582}, g880);
	defparam lut_10381.LUT_SIZE = 3;
	defparam lut_10381.mask = 8'h10;

	lut_sub lut_10387 ({g7, g104}, g881);
	defparam lut_10387.LUT_SIZE = 2;
	defparam lut_10387.mask = 4'b0001;

	lut_sub lut_10393 ({g551, g734}, g882);
	defparam lut_10393.LUT_SIZE = 2;
	defparam lut_10393.mask = 4'b1000;

	lut_sub lut_10401 ({i_8_, g23, g206, g100, g561}, g883);
	defparam lut_10401.LUT_SIZE = 5;
	defparam lut_10401.mask = 32'haa008a00;

	lut_sub lut_10416 ({g101, g185, g881, g882, g883}, g884);
	defparam lut_10416.LUT_SIZE = 5;
	defparam lut_10416.mask = 32'h0000ffef;

	lut_sub lut_10436 ({i_11_, i_9_, i_10_, g323, g875}, g885);
	defparam lut_10436.LUT_SIZE = 5;
	defparam lut_10436.mask = 32'h00100001;

	lut_sub lut_10445 ({i_8_, g10, g66, g100, g108}, g886);
	defparam lut_10445.LUT_SIZE = 5;
	defparam lut_10445.mask = 32'h00000757;

	lut_sub lut_10459 ({g181, g548, g671}, g887);
	defparam lut_10459.LUT_SIZE = 3;
	defparam lut_10459.mask = 8'h80;

	lut_sub lut_10468 ({g8, g221, g323, g544, g887}, g888);
	defparam lut_10468.LUT_SIZE = 5;
	defparam lut_10468.mask = 32'h0f0f0f0e;

	lut_sub lut_10492 ({g136, g609, g881, g885, g886, g888}, g889);
	defparam lut_10492.LUT_SIZE = 6;
	defparam lut_10492.mask = 64'h8080000080000000;

	lut_sub lut_10504 ({g695, g697, g699, g700, g884, g889}, g890);
	defparam lut_10504.LUT_SIZE = 6;
	defparam lut_10504.mask = 64'h0004000000000000;

	lut_sub lut_10511 ({g270, g554, g669}, g891);
	defparam lut_10511.LUT_SIZE = 3;
	defparam lut_10511.mask = 8'h04;

	lut_sub lut_10516 ({i_8_, i_7_, g98}, g892);
	defparam lut_10516.LUT_SIZE = 3;
	defparam lut_10516.mask = 8'h01;

	lut_sub lut_10524 ({i_6_, g43, g131, g461, g892}, g893);
	defparam lut_10524.LUT_SIZE = 5;
	defparam lut_10524.mask = 32'h01010055;

	lut_sub lut_10538 ({g101, g136, g576, g891, g893}, g894);
	defparam lut_10538.LUT_SIZE = 5;
	defparam lut_10538.mask = 32'haa0a2202;

	lut_sub lut_10552 ({g7, g119}, g895);
	defparam lut_10552.LUT_SIZE = 2;
	defparam lut_10552.mask = 4'b0001;

	lut_sub lut_10557 ({i_11_, i_9_, i_10_, g875}, g896);
	defparam lut_10557.LUT_SIZE = 4;
	defparam lut_10557.mask = 16'h1040;

	lut_sub lut_10566 ({i_5_, g141, g326, g660, g896}, g897);
	defparam lut_10566.LUT_SIZE = 5;
	defparam lut_10566.mask = 32'h11131111;

	lut_sub lut_10580 ({g15, g711}, g898);
	defparam lut_10580.LUT_SIZE = 2;
	defparam lut_10580.mask = 4'b0100;

	lut_sub lut_10586 ({g19, g898}, g899);
	defparam lut_10586.LUT_SIZE = 2;
	defparam lut_10586.mask = 4'b1000;

	lut_sub lut_10592 ({i_8_, g100, g899}, g900);
	defparam lut_10592.LUT_SIZE = 3;
	defparam lut_10592.mask = 8'h02;

	lut_sub lut_10601 ({i_8_, g181, g135, g548, g671, g895}, g901);
	defparam lut_10601.LUT_SIZE = 6;
	defparam lut_10601.mask = 64'h00000000007f00ff;

	lut_sub lut_10624 ({g151, g895, g897, g900, g901}, g902);
	defparam lut_10624.LUT_SIZE = 5;
	defparam lut_10624.mask = 32'h80808000;

	lut_sub lut_10634 ({i_8_, g91, g100, g131, g461}, g903);
	defparam lut_10634.LUT_SIZE = 5;
	defparam lut_10634.mask = 32'h11111311;

	lut_sub lut_10652 ({g101, g136, g676, g677, g861, g903}, g904);
	defparam lut_10652.LUT_SIZE = 6;
	defparam lut_10652.mask = 64'hccccc0c088008000;

	lut_sub lut_10675 ({g7, g102, g131, g146, g646}, g905);
	defparam lut_10675.LUT_SIZE = 5;
	defparam lut_10675.mask = 32'h0000ce0a;

	lut_sub lut_10689 ({g7, i_8_, g95, g100, g131}, g906);
	defparam lut_10689.LUT_SIZE = 5;
	defparam lut_10689.mask = 32'h00000013;

	lut_sub lut_10697 ({g7, g102}, g907);
	defparam lut_10697.LUT_SIZE = 2;
	defparam lut_10697.mask = 4'b0010;

	lut_sub lut_10703 ({g7, g11}, g908);
	defparam lut_10703.LUT_SIZE = 2;
	defparam lut_10703.mask = 4'b0001;

	lut_sub lut_10710 ({i_8_, g100, g907, g908}, g909);
	defparam lut_10710.LUT_SIZE = 4;
	defparam lut_10710.mask = 16'h0007;

	lut_sub lut_10719 ({i_8_, g135, g907, g908}, g910);
	defparam lut_10719.LUT_SIZE = 4;
	defparam lut_10719.mask = 16'h0007;

	lut_sub lut_10729 ({g112, g895, g908, g881}, g911);
	defparam lut_10729.LUT_SIZE = 4;
	defparam lut_10729.mask = 16'h007f;

	lut_sub lut_10744 ({i_8_, g264, g108, g895, g907, g881}, g912);
	defparam lut_10744.LUT_SIZE = 6;
	defparam lut_10744.mask = 64'h00000000007f00ff;

	lut_sub lut_10767 ({g906, g909, g910, g911, g912}, g913);
	defparam lut_10767.LUT_SIZE = 5;
	defparam lut_10767.mask = 32'h80000000;

	lut_sub lut_10774 ({g102, g711, g675}, g914);
	defparam lut_10774.LUT_SIZE = 3;
	defparam lut_10774.mask = 8'h8a;

	lut_sub lut_10784 ({i_8_, g100, g112, g887, g914}, g915);
	defparam lut_10784.LUT_SIZE = 5;
	defparam lut_10784.mask = 32'h0c0c0cee;

	lut_sub lut_10804 ({g323, g914, g908, g899, g915}, g916);
	defparam lut_10804.LUT_SIZE = 5;
	defparam lut_10804.mask = 32'haaaa0020;

	lut_sub lut_10822 ({g894, g902, g904, g905, g913, g916}, g917);
	defparam lut_10822.LUT_SIZE = 6;
	defparam lut_10822.mask = 64'h0000000000000010;

	lut_sub lut_10830 ({g880, g694, g890, g917}, g918);
	defparam lut_10830.LUT_SIZE = 4;
	defparam lut_10830.mask = 16'h0001;

	lut_sub lut_10838 ({g316, g216, g207, g895}, g919);
	defparam lut_10838.LUT_SIZE = 4;
	defparam lut_10838.mask = 16'h8000;

	lut_sub lut_10846 ({g547, g532, g676, g896}, g920);
	defparam lut_10846.LUT_SIZE = 4;
	defparam lut_10846.mask = 16'h0080;

	lut_sub lut_10853 ({g185, g551, g734}, g921);
	defparam lut_10853.LUT_SIZE = 3;
	defparam lut_10853.mask = 8'h08;

	lut_sub lut_10860 ({g134, g881, g921}, g922);
	defparam lut_10860.LUT_SIZE = 3;
	defparam lut_10860.mask = 8'h0b;

	lut_sub lut_10870 ({g251, g919, g920, g922}, g923);
	defparam lut_10870.LUT_SIZE = 4;
	defparam lut_10870.mask = 16'haa02;

	lut_sub lut_10883 ({g19, g15, g91, g99, g461}, g924);
	defparam lut_10883.LUT_SIZE = 5;
	defparam lut_10883.mask = 32'h31003333;

	lut_sub lut_10901 ({g316, g669, g676, g896}, g925);
	defparam lut_10901.LUT_SIZE = 4;
	defparam lut_10901.mask = 16'h0800;

	lut_sub lut_10909 ({g99, g887, g924, g925}, g926);
	defparam lut_10909.LUT_SIZE = 4;
	defparam lut_10909.mask = 16'hcc04;

	lut_sub lut_10921 ({g47, g108, g560, g926}, g927);
	defparam lut_10921.LUT_SIZE = 4;
	defparam lut_10921.mask = 16'h5450;

	lut_sub lut_10933 ({g23, g206, g99, g561}, g928);
	defparam lut_10933.LUT_SIZE = 4;
	defparam lut_10933.mask = 16'h3133;

	lut_sub lut_10947 ({g99, g220, g550, g675}, g929);
	defparam lut_10947.LUT_SIZE = 4;
	defparam lut_10947.mask = 16'h007f;

	lut_sub lut_10961 ({g45, g746, g928, g929}, g930);
	defparam lut_10961.LUT_SIZE = 4;
	defparam lut_10961.mask = 16'h8880;

	lut_sub lut_10970 ({g99, g185, g882}, g931);
	defparam lut_10970.LUT_SIZE = 3;
	defparam lut_10970.mask = 8'h0e;

	lut_sub lut_10981 ({g8, g10, g99, g221, g544}, g932);
	defparam lut_10981.LUT_SIZE = 5;
	defparam lut_10981.mask = 32'h0f0f0e0f;

	lut_sub lut_11003 ({g264, g101, g931, g932}, g933);
	defparam lut_11003.LUT_SIZE = 4;
	defparam lut_11003.mask = 16'h8880;

	lut_sub lut_11011 ({g108, g908}, g934);
	defparam lut_11011.LUT_SIZE = 2;
	defparam lut_11011.mask = 4'b0001;

	lut_sub lut_11019 ({g23, g206, g423, g561}, g935);
	defparam lut_11019.LUT_SIZE = 4;
	defparam lut_11019.mask = 16'h3133;

	lut_sub lut_11031 ({i_14_, i_12_, i_13_, g99, g131}, g936);
	defparam lut_11031.LUT_SIZE = 5;
	defparam lut_11031.mask = 32'h01110000;

	lut_sub lut_11039 ({i_14_, i_12_, i_13_, g99, g95}, g937);
	defparam lut_11039.LUT_SIZE = 5;
	defparam lut_11039.mask = 32'h01110000;

	lut_sub lut_11050 ({g99, g908, g935, g936, g937}, g938);
	defparam lut_11050.LUT_SIZE = 5;
	defparam lut_11050.mask = 32'h80808000;

	lut_sub lut_11061 ({g112, g135, g547, g934, g938}, g939);
	defparam lut_11061.LUT_SIZE = 5;
	defparam lut_11061.mask = 32'h44040404;

	lut_sub lut_11074 ({g100, g108, g566, g555, g571}, g940);
	defparam lut_11074.LUT_SIZE = 5;
	defparam lut_11074.mask = 32'hff404040;

	lut_sub lut_11093 ({g8, g221, g101, g544, g940}, g941);
	defparam lut_11093.LUT_SIZE = 5;
	defparam lut_11093.mask = 32'h50505051;

	lut_sub lut_11111 ({g923, g927, g930, g933, g939, g941}, g942);
	defparam lut_11111.LUT_SIZE = 6;
	defparam lut_11111.mask = 64'h0000000000000001;

	lut_sub lut_11117 ({g220, g898}, g943);
	defparam lut_11117.LUT_SIZE = 2;
	defparam lut_11117.mask = 4'b1000;

	lut_sub lut_11127 ({g186, g548, g550, g671, g677, g943}, g944);
	defparam lut_11127.LUT_SIZE = 6;
	defparam lut_11127.mask = 64'h00000000bfffffff;

	lut_sub lut_11167 ({g99, g109, g423, g429, g881, g921}, g945);
	defparam lut_11167.LUT_SIZE = 6;
	defparam lut_11167.mask = 64'hfc54cc44cc44cc44;

	lut_sub lut_11200 ({i_11_, i_9_, i_10_, g99, g186, g875}, g946);
	defparam lut_11200.LUT_SIZE = 6;
	defparam lut_11200.mask = 64'h0000151100000000;

	lut_sub lut_11212 ({g16, g270, g243, g669}, g947);
	defparam lut_11212.LUT_SIZE = 4;
	defparam lut_11212.mask = 16'h3332;

	lut_sub lut_11227 ({g101, g216, g146, g946, g947}, g948);
	defparam lut_11227.LUT_SIZE = 5;
	defparam lut_11227.mask = 32'h88088800;

	lut_sub lut_11239 ({g47, g546, g555, g617}, g949);
	defparam lut_11239.LUT_SIZE = 4;
	defparam lut_11239.mask = 16'h8000;

	lut_sub lut_11246 ({g221, g181, g738}, g950);
	defparam lut_11246.LUT_SIZE = 3;
	defparam lut_11246.mask = 8'h08;

	lut_sub lut_11253 ({i_8_, i_6_, i_7_, g87, g949, g950}, g951);
	defparam lut_11253.LUT_SIZE = 6;
	defparam lut_11253.mask = 64'h0a000000000c0000;

	lut_sub lut_11264 ({g88, g551, g561, g881}, g952);
	defparam lut_11264.LUT_SIZE = 4;
	defparam lut_11264.mask = 16'h007f;

	lut_sub lut_11277 ({i_8_, g100, g108, g895}, g953);
	defparam lut_11277.LUT_SIZE = 4;
	defparam lut_11277.mask = 16'h1505;

	lut_sub lut_11286 ({i_11_, i_9_, i_10_, i_15_, g7}, g954);
	defparam lut_11286.LUT_SIZE = 5;
	defparam lut_11286.mask = 32'h01101000;

	lut_sub lut_11297 ({g59, g66, g118, g943, g954}, g955);
	defparam lut_11297.LUT_SIZE = 5;
	defparam lut_11297.mask = 32'hf3f0a2a0;

	lut_sub lut_11320 ({g284, g676, g952, g953, g955}, g956);
	defparam lut_11320.LUT_SIZE = 5;
	defparam lut_11320.mask = 32'h40404000;

	lut_sub lut_11326 ({i_11_, i_9_, i_10_, i_15_}, g957);
	defparam lut_11326.LUT_SIZE = 4;
	defparam lut_11326.mask = 16'h0180;

	lut_sub lut_11335 ({i_15_, g13, g59, g112, g957}, g958);
	defparam lut_11335.LUT_SIZE = 5;
	defparam lut_11335.mask = 32'h00150055;

	lut_sub lut_11350 ({i_15_, g134, g251, g576, g895, g958}, g959);
	defparam lut_11350.LUT_SIZE = 6;
	defparam lut_11350.mask = 64'haaaa0808ffaa0808;

	lut_sub lut_11383 ({g944, g945, g948, g951, g956, g959}, g960);
	defparam lut_11383.LUT_SIZE = 6;
	defparam lut_11383.mask = 64'h0000001000000000;

	lut_sub lut_11388 ({i_14_, i_12_, i_13_, g104}, g961);
	defparam lut_11388.LUT_SIZE = 4;
	defparam lut_11388.mask = 16'h1500;

	lut_sub lut_11399 ({g23, g206, g323, g561, g921}, g962);
	defparam lut_11399.LUT_SIZE = 5;
	defparam lut_11399.mask = 32'h0f0b0f0f;

	lut_sub lut_11421 ({g112, g135, g532, g962}, g963);
	defparam lut_11421.LUT_SIZE = 4;
	defparam lut_11421.mask = 16'ha888;

	lut_sub lut_11431 ({i_12_, i_13_, i_8_, g108, g135}, g964);
	defparam lut_11431.LUT_SIZE = 5;
	defparam lut_11431.mask = 32'h00000530;

	lut_sub lut_11442 ({g548, g550, g561, g908}, g965);
	defparam lut_11442.LUT_SIZE = 4;
	defparam lut_11442.mask = 16'h8000;

	lut_sub lut_11450 ({i_14_, g131, g277, g964, g965}, g966);
	defparam lut_11450.LUT_SIZE = 5;
	defparam lut_11450.mask = 32'ha0b3a0a0;

	lut_sub lut_11470 ({g109, g551, g495, g961, g963, g966}, g967);
	defparam lut_11470.LUT_SIZE = 6;
	defparam lut_11470.mask = 64'h2222220020202000;

	lut_sub lut_11488 ({g322, g325, g335, g374, g960, g967}, g968);
	defparam lut_11488.LUT_SIZE = 6;
	defparam lut_11488.mask = 64'h0000000000000001;

	lut_sub lut_11498 ({g73, g858, g879, g918, g942, g968}, o_9_);
	defparam lut_11498.LUT_SIZE = 6;
	defparam lut_11498.mask = 64'h00000000fffffffe;

	lut_sub lut_11535 ({g20, g101, g806}, g970);
	defparam lut_11535.LUT_SIZE = 3;
	defparam lut_11535.mask = 8'h31;

	lut_sub lut_11545 ({g101, g339, g465, g924}, g971);
	defparam lut_11545.LUT_SIZE = 4;
	defparam lut_11545.mask = 16'haa20;

	lut_sub lut_11557 ({i_8_, g21, g22, g100, g711}, g972);
	defparam lut_11557.LUT_SIZE = 5;
	defparam lut_11557.mask = 32'h00000133;

	lut_sub lut_11568 ({i_14_, i_12_, i_13_, g18, g15, g99}, g973);
	defparam lut_11568.LUT_SIZE = 6;
	defparam lut_11568.mask = 64'h0044000054005044;

	lut_sub lut_11586 ({g99, g152, g465, g462, g972, g973}, g974);
	defparam lut_11586.LUT_SIZE = 6;
	defparam lut_11586.mask = 64'h8888000000080000;

	lut_sub lut_11599 ({g47, g101, g172, g142, g883}, g975);
	defparam lut_11599.LUT_SIZE = 5;
	defparam lut_11599.mask = 32'h00bf00ff;

	lut_sub lut_11623 ({g12, g101, g970, g971, g974, g975}, g976);
	defparam lut_11623.LUT_SIZE = 6;
	defparam lut_11623.mask = 64'h0200020002000000;

	lut_sub lut_11634 ({g99, g114, g560, g464, g838}, g977);
	defparam lut_11634.LUT_SIZE = 5;
	defparam lut_11634.mask = 32'h0000efff;

	lut_sub lut_11655 ({g451, g928, g977}, g978);
	defparam lut_11655.LUT_SIZE = 3;
	defparam lut_11655.mask = 8'h80;

	lut_sub lut_11661 ({g630, g907}, g979);
	defparam lut_11661.LUT_SIZE = 2;
	defparam lut_11661.mask = 4'b1000;

	lut_sub lut_11667 ({g193, g706}, g980);
	defparam lut_11667.LUT_SIZE = 2;
	defparam lut_11667.mask = 4'b1000;

	lut_sub lut_11674 ({g99, g979, g980}, g981);
	defparam lut_11674.LUT_SIZE = 3;
	defparam lut_11674.mask = 8'h0e;

	lut_sub lut_11682 ({g702, g881}, g982);
	defparam lut_11682.LUT_SIZE = 2;
	defparam lut_11682.mask = 4'b1000;

	lut_sub lut_11692 ({g101, g193, g630, g706, g981, g982}, g983);
	defparam lut_11692.LUT_SIZE = 6;
	defparam lut_11692.mask = 64'hcccccccc40000000;

	lut_sub lut_11717 ({g12, g16, g99, g101, g187}, g984);
	defparam lut_11717.LUT_SIZE = 5;
	defparam lut_11717.mask = 32'hcceec0e0;

	lut_sub lut_11741 ({g101, g534, g899, g978, g983, g984}, g985);
	defparam lut_11741.LUT_SIZE = 6;
	defparam lut_11741.mask = 64'h0101010100010000;

	lut_sub lut_11751 ({g7, g95}, g986);
	defparam lut_11751.LUT_SIZE = 2;
	defparam lut_11751.mask = 4'b0001;

	lut_sub lut_11758 ({i_8_, g100, g522, g986}, g987);
	defparam lut_11758.LUT_SIZE = 4;
	defparam lut_11758.mask = 16'h0703;

	lut_sub lut_11769 ({g99, g835, g887}, g988);
	defparam lut_11769.LUT_SIZE = 3;
	defparam lut_11769.mask = 8'h0e;

	lut_sub lut_11780 ({g46, g66, g99, g209, g531}, g989);
	defparam lut_11780.LUT_SIZE = 5;
	defparam lut_11780.mask = 32'h070f0f0f;

	lut_sub lut_11804 ({g7, g101, g131, g540, g710, g989}, g990);
	defparam lut_11804.LUT_SIZE = 6;
	defparam lut_11804.mask = 64'haaaa8080aaaa8000;

	lut_sub lut_11830 ({i_8_, g4, g98, g213, g986}, g991);
	defparam lut_11830.LUT_SIZE = 5;
	defparam lut_11830.mask = 32'h00030007;

	lut_sub lut_11842 ({g99, g101, g756, g991}, g992);
	defparam lut_11842.LUT_SIZE = 4;
	defparam lut_11842.mask = 16'ha888;

	lut_sub lut_11854 ({g101, g183, g704, g895}, g993);
	defparam lut_11854.LUT_SIZE = 4;
	defparam lut_11854.mask = 16'h007f;

	lut_sub lut_11869 ({g987, g988, g990, g992, g993}, g994);
	defparam lut_11869.LUT_SIZE = 5;
	defparam lut_11869.mask = 32'h02000000;

	lut_sub lut_11878 ({i_8_, g4, g44, g98, g530, g641}, g995);
	defparam lut_11878.LUT_SIZE = 6;
	defparam lut_11878.mask = 64'h0000070f0000050f;

	lut_sub lut_11899 ({g4, g43, g98, g191, g995}, g996);
	defparam lut_11899.LUT_SIZE = 5;
	defparam lut_11899.mask = 32'haaaaa8a0;

	lut_sub lut_11920 ({g99, g101, g187, g534, g907}, g997);
	defparam lut_11920.LUT_SIZE = 5;
	defparam lut_11920.mask = 32'hffaac080;

	lut_sub lut_11942 ({g99, g201, g702, g881}, g998);
	defparam lut_11942.LUT_SIZE = 4;
	defparam lut_11942.mask = 16'h00f7;

	lut_sub lut_11955 ({g996, g997, g998}, g999);
	defparam lut_11955.LUT_SIZE = 3;
	defparam lut_11955.mask = 8'h02;

	lut_sub lut_11963 ({g976, g985, g994, g999}, g1000);
	defparam lut_11963.LUT_SIZE = 4;
	defparam lut_11963.mask = 16'h0001;

	lut_sub lut_11970 ({g46, g209, g531}, g1001);
	defparam lut_11970.LUT_SIZE = 3;
	defparam lut_11970.mask = 8'h80;

	lut_sub lut_11977 ({i_14_, i_12_, i_13_, g99, g95, g93}, g1002);
	defparam lut_11977.LUT_SIZE = 6;
	defparam lut_11977.mask = 64'h000303030a0a0a00;

	lut_sub lut_11997 ({g99, g268, g96, g669, g818}, g1003);
	defparam lut_11997.LUT_SIZE = 5;
	defparam lut_11997.mask = 32'h0000feff;

	lut_sub lut_12018 ({i_14_, i_12_, i_13_, g95, g101, g93}, g1004);
	defparam lut_12018.LUT_SIZE = 6;
	defparam lut_12018.mask = 64'h0000000023232203;

	lut_sub lut_12036 ({g101, g94, g475, g678, g891}, g1005);
	defparam lut_12036.LUT_SIZE = 5;
	defparam lut_12036.mask = 32'h0000feff;

	lut_sub lut_12058 ({g1002, g1003, g1004, g1005}, g1006);
	defparam lut_12058.LUT_SIZE = 4;
	defparam lut_12058.mask = 16'h8000;

	lut_sub lut_12065 ({i_9_, i_8_, g30, g326, g98}, g1007);
	defparam lut_12065.LUT_SIZE = 5;
	defparam lut_12065.mask = 32'h00010100;

	lut_sub lut_12074 ({g101, g1001, g1006, g1007}, g1008);
	defparam lut_12074.LUT_SIZE = 4;
	defparam lut_12074.mask = 16'h2202;

	lut_sub lut_12085 ({g99, g264, g115, g711, g672}, g1009);
	defparam lut_12085.LUT_SIZE = 5;
	defparam lut_12085.mask = 32'h000075ff;

	lut_sub lut_12105 ({g101, g696, g672, g1009}, g1010);
	defparam lut_12105.LUT_SIZE = 4;
	defparam lut_12105.mask = 16'haa08;

	lut_sub lut_12117 ({g99, g101, g696, g670}, g1011);
	defparam lut_12117.LUT_SIZE = 4;
	defparam lut_12117.mask = 16'h05cd;

	lut_sub lut_12133 ({g10, g99, g220, g221, g550, g544}, g1012);
	defparam lut_12133.LUT_SIZE = 6;
	defparam lut_12133.mask = 64'h0000fbff0000ffff;

	lut_sub lut_12173 ({g10, g14, g101, g677, g903, g1012}, g1013);
	defparam lut_12173.LUT_SIZE = 6;
	defparam lut_12173.mask = 64'haa80aa00aa00aa00;

	lut_sub lut_12197 ({g102, g119, g544, g711}, g1014);
	defparam lut_12197.LUT_SIZE = 4;
	defparam lut_12197.mask = 16'h2232;

	lut_sub lut_12208 ({i_8_, g100, g551, g1014}, g1015);
	defparam lut_12208.LUT_SIZE = 4;
	defparam lut_12208.mask = 16'h030b;

	lut_sub lut_12220 ({g324, g440, g864, g1015}, g1016);
	defparam lut_12220.LUT_SIZE = 4;
	defparam lut_12220.mask = 16'h8000;

	lut_sub lut_12229 ({g267, g714, g1011, g1013, g1016}, g1017);
	defparam lut_12229.LUT_SIZE = 5;
	defparam lut_12229.mask = 32'h00001000;

	lut_sub lut_12238 ({g106, g570, g575, g1010, g1017}, g1018);
	defparam lut_12238.LUT_SIZE = 5;
	defparam lut_12238.mask = 32'h00000100;

	lut_sub lut_12246 ({i_8_, g100, g177, g114, g560}, g1019);
	defparam lut_12246.LUT_SIZE = 5;
	defparam lut_12246.mask = 32'haaaaaa80;

	lut_sub lut_12264 ({g101, g1019}, g1020);
	defparam lut_12264.LUT_SIZE = 2;
	defparam lut_12264.mask = 4'b0010;

	lut_sub lut_12274 ({g99, g101, g226, g464, g703, g908}, g1021);
	defparam lut_12274.LUT_SIZE = 6;
	defparam lut_12274.mask = 64'hffff000888880008;

	lut_sub lut_12302 ({i_14_, i_12_, i_13_, g99, g119, g122}, g1022);
	defparam lut_12302.LUT_SIZE = 6;
	defparam lut_12302.mask = 64'h000b00000a0b0b0b;

	lut_sub lut_12322 ({g99, g535, g1022}, g1023);
	defparam lut_12322.LUT_SIZE = 3;
	defparam lut_12322.mask = 8'ha2;

	lut_sub lut_12333 ({g14, g99, g197, g90, g895}, g1024);
	defparam lut_12333.LUT_SIZE = 5;
	defparam lut_12333.mask = 32'h00df00ff;

	lut_sub lut_12355 ({g101, g201, g530, g1024}, g1025);
	defparam lut_12355.LUT_SIZE = 4;
	defparam lut_12355.mask = 16'haa08;

	lut_sub lut_12367 ({g7, g131, g171, g158}, g1026);
	defparam lut_12367.LUT_SIZE = 4;
	defparam lut_12367.mask = 16'h444f;

	lut_sub lut_12382 ({i_8_, g66, g100, g253, g132, g279}, g1027);
	defparam lut_12382.LUT_SIZE = 6;
	defparam lut_12382.mask = 64'h0000000000df00ff;

	lut_sub lut_12406 ({g648, g1020, g1021, g1023, g1025, g1542}, g1028);
	defparam lut_12406.LUT_SIZE = 6;
	defparam lut_12406.mask = 64'h0001000000000000;

	lut_sub lut_12415 ({g73, g1000, g1008, g1018, g1028}, g1029);
	defparam lut_12415.LUT_SIZE = 5;
	defparam lut_12415.mask = 32'hffff0001;

	lut_sub lut_12439 ({g213, g557, g522, g756}, g1030);
	defparam lut_12439.LUT_SIZE = 4;
	defparam lut_12439.mask = 16'h8000;

	lut_sub lut_12449 ({g44, g556, g544, g641, g876, g1030}, g1031);
	defparam lut_12449.LUT_SIZE = 6;
	defparam lut_12449.mask = 64'h0000004000000000;

	lut_sub lut_12455 ({i_14_, i_12_, i_13_, g131, g158}, g1032);
	defparam lut_12455.LUT_SIZE = 5;
	defparam lut_12455.mask = 32'hc8ccafca;

	lut_sub lut_12477 ({g6, i_15_, i_14_, i_12_, i_13_, g59}, g1033);
	defparam lut_12477.LUT_SIZE = 6;
	defparam lut_12477.mask = 64'h0000000014555555;

	lut_sub lut_12499 ({g18, g59, g142, g465, g726}, g1034);
	defparam lut_12499.LUT_SIZE = 5;
	defparam lut_12499.mask = 32'h00ef00cf;

	lut_sub lut_12518 ({i_14_, i_12_, i_13_, g18, g15, g59}, g1035);
	defparam lut_12518.LUT_SIZE = 6;
	defparam lut_12518.mask = 64'h0044440000005444;

	lut_sub lut_12533 ({i_14_, i_12_, i_13_, g59, g95, g93}, g1036);
	defparam lut_12533.LUT_SIZE = 6;
	defparam lut_12533.mask = 64'h0a030b0a030b0a03;

	lut_sub lut_12557 ({i_14_, i_12_, i_13_, g131, g158, g284}, g1037);
	defparam lut_12557.LUT_SIZE = 6;
	defparam lut_12557.mask = 64'h1100111105151105;

	lut_sub lut_12580 ({g1033, g1034, g1035, g1036, g1037}, g1038);
	defparam lut_12580.LUT_SIZE = 5;
	defparam lut_12580.mask = 32'h80000000;

	lut_sub lut_12585 ({i_11_, i_15_, i_14_, i_12_, i_13_, g113}, g1039);
	defparam lut_12585.LUT_SIZE = 6;
	defparam lut_12585.mask = 64'h0551454000000000;

	lut_sub lut_12599 ({g323, g1039}, g1040);
	defparam lut_12599.LUT_SIZE = 2;
	defparam lut_12599.mask = 4'b0001;

	lut_sub lut_12607 ({g12, g177, g114, g560}, g1041);
	defparam lut_12607.LUT_SIZE = 4;
	defparam lut_12607.mask = 16'h8000;

	lut_sub lut_12614 ({g323, g187, g534}, g1042);
	defparam lut_12614.LUT_SIZE = 3;
	defparam lut_12614.mask = 8'h07;

	lut_sub lut_12625 ({g12, g323, g201, g703, g908}, g1043);
	defparam lut_12625.LUT_SIZE = 5;
	defparam lut_12625.mask = 32'h00f700ff;

	lut_sub lut_12648 ({g423, g838, g935, g1042, g1043}, g1044);
	defparam lut_12648.LUT_SIZE = 5;
	defparam lut_12648.mask = 32'h80800080;

	lut_sub lut_12658 ({g423, g1040, g1041, g1044}, g1045);
	defparam lut_12658.LUT_SIZE = 4;
	defparam lut_12658.mask = 16'h5010;

	lut_sub lut_12667 ({g323, g226, g464}, g1046);
	defparam lut_12667.LUT_SIZE = 3;
	defparam lut_12667.mask = 8'h0e;

	lut_sub lut_12679 ({g323, g224, g423, g467, g817, g1046}, g1047);
	defparam lut_12679.LUT_SIZE = 6;
	defparam lut_12679.mask = 64'haa08aa0008080000;

	lut_sub lut_12695 ({i_14_, i_12_, i_13_, g119, g122}, g1048);
	defparam lut_12695.LUT_SIZE = 5;
	defparam lut_12695.mask = 32'ha3bb3000;

	lut_sub lut_12712 ({i_14_, i_12_, i_13_, g104, g124}, g1049);
	defparam lut_12712.LUT_SIZE = 5;
	defparam lut_12712.mask = 32'h00557303;

	lut_sub lut_12731 ({g323, g90, g528, g921, g1049}, g1050);
	defparam lut_12731.LUT_SIZE = 5;
	defparam lut_12731.mask = 32'h0000fffd;

	lut_sub lut_12752 ({g423, g1048, g1050}, g1051);
	defparam lut_12752.LUT_SIZE = 3;
	defparam lut_12752.mask = 8'ha8;

	lut_sub lut_12760 ({i_14_, i_12_, i_13_, g95, g93}, g1052);
	defparam lut_12760.LUT_SIZE = 5;
	defparam lut_12760.mask = 32'h5c44445c;

	lut_sub lut_12780 ({g120, g349, g423, g613, g481}, g1053);
	defparam lut_12780.LUT_SIZE = 5;
	defparam lut_12780.mask = 32'h0f0f0e0f;

	lut_sub lut_12801 ({g323, g835, g1053}, g1054);
	defparam lut_12801.LUT_SIZE = 3;
	defparam lut_12801.mask = 8'ha2;

	lut_sub lut_12809 ({i_14_, i_12_, i_13_, g95, g93}, g1055);
	defparam lut_12809.LUT_SIZE = 5;
	defparam lut_12809.mask = 32'ha033a303;

	lut_sub lut_12828 ({g323, g678, g670, g756}, g1056);
	defparam lut_12828.LUT_SIZE = 4;
	defparam lut_12828.mask = 16'h00f7;

	lut_sub lut_12842 ({g323, g203, g213, g474}, g1057);
	defparam lut_12842.LUT_SIZE = 4;
	defparam lut_12842.mask = 16'h007f;

	lut_sub lut_12858 ({g323, g818, g887, g1055, g1056, g1057}, g1058);
	defparam lut_12858.LUT_SIZE = 6;
	defparam lut_12858.mask = 64'h8888888800000080;

	lut_sub lut_12874 ({g423, g1052, g1054, g1058}, g1059);
	defparam lut_12874.LUT_SIZE = 4;
	defparam lut_12874.mask = 16'h1101;

	lut_sub lut_12883 ({g6, i_15_, g7, g182}, g1060);
	defparam lut_12883.LUT_SIZE = 4;
	defparam lut_12883.mask = 16'h0070;

	lut_sub lut_12891 ({i_14_, i_12_, i_13_, g131, g158}, g1061);
	defparam lut_12891.LUT_SIZE = 5;
	defparam lut_12891.mask = 32'h35000575;

	lut_sub lut_12910 ({g46, g642, g522, g896, g1061}, g1062);
	defparam lut_12910.LUT_SIZE = 5;
	defparam lut_12910.mask = 32'h00800000;

	lut_sub lut_12918 ({i_11_, g113, g9, g423, g1049}, g1063);
	defparam lut_12918.LUT_SIZE = 5;
	defparam lut_12918.mask = 32'h11111113;

	lut_sub lut_12933 ({g183, g704, g895}, g1064);
	defparam lut_12933.LUT_SIZE = 3;
	defparam lut_12933.mask = 8'h80;

	lut_sub lut_12941 ({g323, g120, g613, g1064}, g1065);
	defparam lut_12941.LUT_SIZE = 4;
	defparam lut_12941.mask = 16'h00fe;

	lut_sub lut_12955 ({g47, g323, g172, g142}, g1066);
	defparam lut_12955.LUT_SIZE = 4;
	defparam lut_12955.mask = 16'h070f;

	lut_sub lut_12970 ({g44, g323, g191, g339, g807}, g1067);
	defparam lut_12970.LUT_SIZE = 5;
	defparam lut_12970.mask = 32'h00bf00ff;

	lut_sub lut_12993 ({g323, g465, g899, g1066, g1067}, g1068);
	defparam lut_12993.LUT_SIZE = 5;
	defparam lut_12993.mask = 32'h88880008;

	lut_sub lut_13005 ({g323, g349, g481, g540}, g1069);
	defparam lut_13005.LUT_SIZE = 4;
	defparam lut_13005.mask = 16'h00df;

	lut_sub lut_13021 ({g10, g323, g423, g677, g921, g1069}, g1070);
	defparam lut_13021.LUT_SIZE = 6;
	defparam lut_13021.mask = 64'haa22a020aa220000;

	lut_sub lut_13044 ({g207, g323, g246, g576, g724}, g1071);
	defparam lut_13044.LUT_SIZE = 5;
	defparam lut_13044.mask = 32'h00df00ff;

	lut_sub lut_13067 ({g8, g221, g323, g544, g1071}, g1072);
	defparam lut_13067.LUT_SIZE = 5;
	defparam lut_13067.mask = 32'ha0a0a0a2;

	lut_sub lut_13084 ({g1063, g1065, g1068, g1070, g1072}, g1073);
	defparam lut_13084.LUT_SIZE = 5;
	defparam lut_13084.mask = 32'h01000000;

	lut_sub lut_13093 ({g243, g1673, g1060, g1062, g1073}, g1074);
	defparam lut_13093.LUT_SIZE = 5;
	defparam lut_13093.mask = 32'h00550010;

	lut_sub lut_13105 ({g142, g540, g724, g895}, g1075);
	defparam lut_13105.LUT_SIZE = 4;
	defparam lut_13105.mask = 16'h8000;

	lut_sub lut_13110 ({i_14_, i_12_, i_13_, g102}, g1076);
	defparam lut_13110.LUT_SIZE = 4;
	defparam lut_13110.mask = 16'h2a00;

	lut_sub lut_13117 ({g6, i_15_, i_14_, i_12_, i_13_}, g1077);
	defparam lut_13117.LUT_SIZE = 5;
	defparam lut_13117.mask = 32'h00006588;

	lut_sub lut_13130 ({g232, g103, g1076, g1077}, g1078);
	defparam lut_13130.LUT_SIZE = 4;
	defparam lut_13130.mask = 16'h0800;

	lut_sub lut_13139 ({g44, g183, g191, g704, g756}, g1079);
	defparam lut_13139.LUT_SIZE = 5;
	defparam lut_13139.mask = 32'h80000000;

	lut_sub lut_13148 ({g316, g172, g173, g339, g1079}, g1080);
	defparam lut_13148.LUT_SIZE = 5;
	defparam lut_13148.mask = 32'h40000000;

	lut_sub lut_13157 ({g222, g908, g1075, g1078, g1080}, g1081);
	defparam lut_13157.LUT_SIZE = 5;
	defparam lut_13157.mask = 32'h01000000;

	lut_sub lut_13162 ({i_14_, i_12_, g115}, g1082);
	defparam lut_13162.LUT_SIZE = 3;
	defparam lut_13162.mask = 8'h08;

	lut_sub lut_13172 ({g19, g201, g675, g797, g703, g1082}, g1083);
	defparam lut_13172.LUT_SIZE = 6;
	defparam lut_13172.mask = 64'h0000800000000000;

	lut_sub lut_13181 ({g132, g576, g557, g465, g1083}, g1084);
	defparam lut_13181.LUT_SIZE = 5;
	defparam lut_13181.mask = 32'h00000010;

	lut_sub lut_13190 ({g207, g213, g279, g544, g881}, g1085);
	defparam lut_13190.LUT_SIZE = 5;
	defparam lut_13190.mask = 32'h20000000;

	lut_sub lut_13197 ({g243, g630, g980}, g1086);
	defparam lut_13197.LUT_SIZE = 3;
	defparam lut_13197.mask = 8'h0b;

	lut_sub lut_13207 ({g323, g173, g103, g546}, g1087);
	defparam lut_13207.LUT_SIZE = 4;
	defparam lut_13207.mask = 16'h00df;

	lut_sub lut_13222 ({g187, g423, g534, g907, g1087}, g1088);
	defparam lut_13222.LUT_SIZE = 5;
	defparam lut_13222.mask = 32'haa80aa00;

	lut_sub lut_13236 ({i_11_, i_10_, g323, g875}, g1089);
	defparam lut_13236.LUT_SIZE = 4;
	defparam lut_13236.mask = 16'h0001;

	lut_sub lut_13245 ({g48, g323, g182, g124, g115}, g1090);
	defparam lut_13245.LUT_SIZE = 5;
	defparam lut_13245.mask = 32'h00bb000b;

	lut_sub lut_13263 ({g323, g696, g702, g827, g914, g1090}, g1091);
	defparam lut_13263.LUT_SIZE = 6;
	defparam lut_13263.mask = 64'haaaaaaaa00000200;

	lut_sub lut_13288 ({g829, g1086, g1088, g1089, g1091}, g1092);
	defparam lut_13288.LUT_SIZE = 5;
	defparam lut_13288.mask = 32'h04000000;

	lut_sub lut_13297 ({g423, g1081, g1084, g1085, g1092}, g1093);
	defparam lut_13297.LUT_SIZE = 5;
	defparam lut_13297.mask = 32'h55550001;

	lut_sub lut_13315 ({g1045, g1047, g1051, g1059, g1074, g1093}, g1094);
	defparam lut_13315.LUT_SIZE = 6;
	defparam lut_13315.mask = 64'h0000000000000001;

	lut_sub lut_13321 ({g89, g627}, g1095);
	defparam lut_13321.LUT_SIZE = 2;
	defparam lut_13321.mask = 4'b1000;

	lut_sub lut_13327 ({g21, g114}, g1096);
	defparam lut_13327.LUT_SIZE = 2;
	defparam lut_13327.mask = 4'b1000;

	lut_sub lut_13332 ({i_14_, i_13_, g22}, g1097);
	defparam lut_13332.LUT_SIZE = 3;
	defparam lut_13332.mask = 8'h40;

	lut_sub lut_13341 ({g151, g506, g594, g1096, g1097}, g1098);
	defparam lut_13341.LUT_SIZE = 5;
	defparam lut_13341.mask = 32'h0000fdff;

	lut_sub lut_13361 ({g187, g982}, g1099);
	defparam lut_13361.LUT_SIZE = 2;
	defparam lut_13361.mask = 4'b0100;

	lut_sub lut_13368 ({g151, g534, g1099}, g1100);
	defparam lut_13368.LUT_SIZE = 3;
	defparam lut_13368.mask = 8'h0b;

	lut_sub lut_13378 ({g1095, g1098, g1100, g1541}, g1101);
	defparam lut_13378.LUT_SIZE = 4;
	defparam lut_13378.mask = 16'h4000;

	lut_sub lut_13386 ({i_8_, g46, g88, g224, g811}, g1102);
	defparam lut_13386.LUT_SIZE = 5;
	defparam lut_13386.mask = 32'hfffff8f0;

	lut_sub lut_13416 ({i_14_, i_12_, i_13_, g104, g124}, g1103);
	defparam lut_13416.LUT_SIZE = 5;
	defparam lut_13416.mask = 32'hafa888ac;

	lut_sub lut_13439 ({g14, g46, g89, g442, g1103}, g1104);
	defparam lut_13439.LUT_SIZE = 5;
	defparam lut_13439.mask = 32'h4c0c0c0c;

	lut_sub lut_13454 ({g1628, g1622, g1104}, g1105);
	defparam lut_13454.LUT_SIZE = 3;
	defparam lut_13454.mask = 8'h01;

	lut_sub lut_13461 ({i_14_, i_12_, i_13_, g95, g151, g93}, g1106);
	defparam lut_13461.LUT_SIZE = 6;
	defparam lut_13461.mask = 64'h2323220022220023;

	lut_sub lut_13482 ({i_8_, g88, g203, g475}, g1107);
	defparam lut_13482.LUT_SIZE = 4;
	defparam lut_13482.mask = 16'h0a03;

	lut_sub lut_13493 ({i_8_, g88, g304, g270, g213}, g1108);
	defparam lut_13493.LUT_SIZE = 5;
	defparam lut_13493.mask = 32'h00cf00dd;

	lut_sub lut_13514 ({g89, g93, g572, g849, g1107, g1108}, g1109);
	defparam lut_13514.LUT_SIZE = 6;
	defparam lut_13514.mask = 64'h8000808080808080;

	lut_sub lut_13530 ({g89, g97, g678, g669, g1106, g1109}, g1110);
	defparam lut_13530.LUT_SIZE = 6;
	defparam lut_13530.mask = 64'h0004000044440000;

	lut_sub lut_13543 ({g268, g172, g556, g986, g1030}, g1111);
	defparam lut_13543.LUT_SIZE = 5;
	defparam lut_13543.mask = 32'h04000000;

	lut_sub lut_13551 ({g20, g460, g1032, g1111}, g1112);
	defparam lut_13551.LUT_SIZE = 4;
	defparam lut_13551.mask = 16'h0010;

	lut_sub lut_13560 ({g204, g548, g881, g1096, g1075}, g1113);
	defparam lut_13560.LUT_SIZE = 5;
	defparam lut_13560.mask = 32'h00001000;

	lut_sub lut_13569 ({g181, g123, g670, g671, g702}, g1114);
	defparam lut_13569.LUT_SIZE = 5;
	defparam lut_13569.mask = 32'h80000000;

	lut_sub lut_13578 ({g10, g45, g221, g187, g1114}, g1115);
	defparam lut_13578.LUT_SIZE = 5;
	defparam lut_13578.mask = 32'h04000000;

	lut_sub lut_13586 ({i_8_, g88, g534, g979, g980}, g1116);
	defparam lut_13586.LUT_SIZE = 5;
	defparam lut_13586.mask = 32'hff10ff11;

	lut_sub lut_13610 ({i_14_, i_12_, i_13_, g102, g115}, g1117);
	defparam lut_13610.LUT_SIZE = 5;
	defparam lut_13610.mask = 32'h000aee0c;

	lut_sub lut_13627 ({i_8_, g88, g232, g116, g675}, g1118);
	defparam lut_13627.LUT_SIZE = 5;
	defparam lut_13627.mask = 32'hff80fff0;

	lut_sub lut_13656 ({g89, g1112, g1113, g1115, g1616}, g1119);
	defparam lut_13656.LUT_SIZE = 5;
	defparam lut_13656.mask = 32'h00015555;

	lut_sub lut_13672 ({g115, g554, g460, g711}, g1120);
	defparam lut_13672.LUT_SIZE = 4;
	defparam lut_13672.mask = 16'h80c0;

	lut_sub lut_13682 ({g253, g710, g1026, g1120}, g1121);
	defparam lut_13682.LUT_SIZE = 4;
	defparam lut_13682.mask = 16'h4000;

	lut_sub lut_13689 ({g44, g191, g641}, g1122);
	defparam lut_13689.LUT_SIZE = 3;
	defparam lut_13689.mask = 8'h80;

	lut_sub lut_13695 ({g6, i_15_, i_14_, i_12_, i_13_, g122}, g1123);
	defparam lut_13695.LUT_SIZE = 6;
	defparam lut_13695.mask = 64'h02a002a003ac02a3;

	lut_sub lut_13718 ({i_9_, i_10_, g7, g53, g91}, g1124);
	defparam lut_13718.LUT_SIZE = 5;
	defparam lut_13718.mask = 32'h00230303;

	lut_sub lut_13732 ({g1076, g1122, g1123, g1124}, g1125);
	defparam lut_13732.LUT_SIZE = 4;
	defparam lut_13732.mask = 16'h0800;

	lut_sub lut_13740 ({i_8_, g88, g1084, g1121, g1125}, g1126);
	defparam lut_13740.LUT_SIZE = 5;
	defparam lut_13740.mask = 32'h00aa00fe;

	lut_sub lut_13756 ({i_14_, i_12_, i_13_, g119, g122}, g1127);
	defparam lut_13756.LUT_SIZE = 5;
	defparam lut_13756.mask = 32'haaa3003a;

	lut_sub lut_13776 ({i_8_, g88, g349, g670, g704, g895}, g1128);
	defparam lut_13776.LUT_SIZE = 6;
	defparam lut_13776.mask = 64'h000033ff00005fff;

	lut_sub lut_13810 ({i_8_, g88, g181, g183, g1127, g1128}, g1129);
	defparam lut_13810.LUT_SIZE = 6;
	defparam lut_13810.mask = 64'haaaaa0a0aaaa8800;

	lut_sub lut_13839 ({i_8_, g88, g339, g117, g806}, g1130);
	defparam lut_13839.LUT_SIZE = 5;
	defparam lut_13839.mask = 32'h003f005f;

	lut_sub lut_13860 ({g19, g16, g89, g465, g462, g1130}, g1131);
	defparam lut_13860.LUT_SIZE = 6;
	defparam lut_13860.mask = 64'h00aa02aa00aa00aa;

	lut_sub lut_13882 ({i_14_, i_12_, i_13_, g104, g124}, g1132);
	defparam lut_13882.LUT_SIZE = 5;
	defparam lut_13882.mask = 32'h50577703;

	lut_sub lut_13904 ({i_8_, g88, g185, g696, g1132}, g1133);
	defparam lut_13904.LUT_SIZE = 5;
	defparam lut_13904.mask = 32'h00fc0055;

	lut_sub lut_13920 ({i_14_, i_12_, i_13_, g131, g151, g158}, g1134);
	defparam lut_13920.LUT_SIZE = 6;
	defparam lut_13920.mask = 64'h1100131103001103;

	lut_sub lut_13941 ({g8, g10, g151, g1133, g1134}, g1135);
	defparam lut_13941.LUT_SIZE = 5;
	defparam lut_13941.mask = 32'h80808880;

	lut_sub lut_13954 ({g176, g1126, g1129, g1131, g1135}, g1136);
	defparam lut_13954.LUT_SIZE = 5;
	defparam lut_13954.mask = 32'h01000000;

	lut_sub lut_13963 ({g1101, g1105, g1110, g1119, g1136}, g1137);
	defparam lut_13963.LUT_SIZE = 5;
	defparam lut_13963.mask = 32'h00000001;

	lut_sub lut_13967 ({i_1_, i_0_, i_2_}, g1138);
	defparam lut_13967.LUT_SIZE = 3;
	defparam lut_13967.mask = 8'h9b;

	lut_sub lut_13978 ({g20, g460, g710}, g1139);
	defparam lut_13978.LUT_SIZE = 3;
	defparam lut_13978.mask = 8'h08;

	lut_sub lut_13984 ({g528, g1031}, g1140);
	defparam lut_13984.LUT_SIZE = 2;
	defparam lut_13984.mask = 4'b0001;

	lut_sub lut_13991 ({i_8_, g23, g108, g506}, g1141);
	defparam lut_13991.LUT_SIZE = 4;
	defparam lut_13991.mask = 16'h0013;

	lut_sub lut_14000 ({i_8_, g21, g108, g561}, g1142);
	defparam lut_14000.LUT_SIZE = 4;
	defparam lut_14000.mask = 16'h0013;

	lut_sub lut_14012 ({g145, g127, g114, g596, g1141, g1142}, g1143);
	defparam lut_14012.LUT_SIZE = 6;
	defparam lut_14012.mask = 64'h8080808000008000;

	lut_sub lut_14026 ({g112, g136, g474, g1139, g1140, g1143}, g1144);
	defparam lut_14026.LUT_SIZE = 6;
	defparam lut_14026.mask = 64'h5555010111000100;

	lut_sub lut_14048 ({g880, g694, g860, g890, g917, g1144}, g1145);
	defparam lut_14048.LUT_SIZE = 6;
	defparam lut_14048.mask = 64'h0000000000000001;

	lut_sub lut_14054 ({i_11_, i_9_, i_10_, i_15_, g7, g9}, g1146);
	defparam lut_14054.LUT_SIZE = 6;
	defparam lut_14054.mask = 64'h5005303500000000;

	lut_sub lut_14071 ({g151, g544, g487, g1146}, g1147);
	defparam lut_14071.LUT_SIZE = 4;
	defparam lut_14071.mask = 16'h00f7;

	lut_sub lut_14084 ({g112, g114, g464}, g1148);
	defparam lut_14084.LUT_SIZE = 3;
	defparam lut_14084.mask = 8'h0b;

	lut_sub lut_14093 ({i_14_, i_12_, i_13_, g11, g22, g112}, g1149);
	defparam lut_14093.LUT_SIZE = 6;
	defparam lut_14093.mask = 64'h1105050000001105;

	lut_sub lut_14111 ({g112, g183, g123, g670, g887}, g1150);
	defparam lut_14111.LUT_SIZE = 5;
	defparam lut_14111.mask = 32'h0000bfff;

	lut_sub lut_14134 ({g562, g804, g1148, g1149, g1150}, g1151);
	defparam lut_14134.LUT_SIZE = 5;
	defparam lut_14134.mask = 32'h80000000;

	lut_sub lut_14141 ({i_14_, i_12_, i_13_, g104, g136, g124}, g1152);
	defparam lut_14141.LUT_SIZE = 6;
	defparam lut_14141.mask = 64'h1100131313030003;

	lut_sub lut_14162 ({i_14_, i_12_, i_13_, g104, g112, g124}, g1153);
	defparam lut_14162.LUT_SIZE = 6;
	defparam lut_14162.mask = 64'h1100131313030003;

	lut_sub lut_14185 ({g101, g323, g231, g478, g1001}, g1154);
	defparam lut_14185.LUT_SIZE = 5;
	defparam lut_14185.mask = 32'hff0c5504;

	lut_sub lut_14206 ({i_14_, i_12_, i_13_, g104, g145, g124}, g1155);
	defparam lut_14206.LUT_SIZE = 6;
	defparam lut_14206.mask = 64'h1100111313130003;

	lut_sub lut_14229 ({g1151, g1152, g1153, g1154, g1155}, g1156);
	defparam lut_14229.LUT_SIZE = 5;
	defparam lut_14229.mask = 32'h00002000;

	lut_sub lut_14237 ({i_8_, g108, g183, g540, g704}, g1157);
	defparam lut_14237.LUT_SIZE = 5;
	defparam lut_14237.mask = 32'h88888880;

	lut_sub lut_14249 ({g145, g1157}, g1158);
	defparam lut_14249.LUT_SIZE = 2;
	defparam lut_14249.mask = 4'b0010;

	lut_sub lut_14258 ({g268, g556, g669, g672, g979}, g1159);
	defparam lut_14258.LUT_SIZE = 5;
	defparam lut_14258.mask = 32'h00040000;

	lut_sub lut_14268 ({g16, g323, g534, g980, g1062, g1159}, g1160);
	defparam lut_14268.LUT_SIZE = 6;
	defparam lut_14268.mask = 64'h0000ffff0000feff;

	lut_sub lut_14304 ({i_14_, i_12_, g119, g485}, g1161);
	defparam lut_14304.LUT_SIZE = 4;
	defparam lut_14304.mask = 16'haa8a;

	lut_sub lut_14317 ({g112, g199, g547}, g1162);
	defparam lut_14317.LUT_SIZE = 3;
	defparam lut_14317.mask = 8'h0b;

	lut_sub lut_14328 ({g101, g151, g1064, g1161, g1162}, g1163);
	defparam lut_14328.LUT_SIZE = 5;
	defparam lut_14328.mask = 32'haa220a02;

	lut_sub lut_14342 ({g6, i_15_, i_14_, i_12_, i_13_, g101}, g1164);
	defparam lut_14342.LUT_SIZE = 6;
	defparam lut_14342.mask = 64'h0000000005514540;

	lut_sub lut_14358 ({i_8_, g108, g201, g703, g908}, g1165);
	defparam lut_14358.LUT_SIZE = 5;
	defparam lut_14358.mask = 32'h000000f7;

	lut_sub lut_14373 ({g101, g199, g120, g547, g1165}, g1166);
	defparam lut_14373.LUT_SIZE = 5;
	defparam lut_14373.mask = 32'haaaa0200;

	lut_sub lut_14391 ({g1065, g1158, g1160, g1163, g1164, g1166}, g1167);
	defparam lut_14391.LUT_SIZE = 6;
	defparam lut_14391.mask = 64'h0400000000000000;

	lut_sub lut_14396 ({i_12_, i_13_, g93}, g1168);
	defparam lut_14396.LUT_SIZE = 3;
	defparam lut_14396.mask = 8'h02;

	lut_sub lut_14403 ({g13, g115, g711}, g1169);
	defparam lut_14403.LUT_SIZE = 3;
	defparam lut_14403.mask = 8'h4c;

	lut_sub lut_14413 ({i_8_, g264, g100, g103, g1169}, g1170);
	defparam lut_14413.LUT_SIZE = 5;
	defparam lut_14413.mask = 32'haaaaa2a0;

	lut_sub lut_14435 ({g20, g101, g173, g806, g1168, g1170}, g1171);
	defparam lut_14435.LUT_SIZE = 6;
	defparam lut_14435.mask = 64'h0000ffff0000bfff;

	lut_sub lut_14475 ({g145, g261, g524, g525, g710, g1122}, g1172);
	defparam lut_14475.LUT_SIZE = 6;
	defparam lut_14475.mask = 64'hf000000040000000;

	lut_sub lut_14489 ({g843, g845, g847, g851, g1171, g1172}, g1173);
	defparam lut_14489.LUT_SIZE = 6;
	defparam lut_14489.mask = 64'h0000000400000000;

	lut_sub lut_14497 ({g112, g216, g120, g485}, g1174);
	defparam lut_14497.LUT_SIZE = 4;
	defparam lut_14497.mask = 16'h00df;

	lut_sub lut_14512 ({g136, g226, g506, g670, g1001}, g1175);
	defparam lut_14512.LUT_SIZE = 5;
	defparam lut_14512.mask = 32'h0000ffbf;

	lut_sub lut_14534 ({i_8_, g135, g114, g560, g464}, g1176);
	defparam lut_14534.LUT_SIZE = 5;
	defparam lut_14534.mask = 32'h000000bf;

	lut_sub lut_14549 ({g21, g136, g177, g120, g1176}, g1177);
	defparam lut_14549.LUT_SIZE = 5;
	defparam lut_14549.mask = 32'haa20aa00;

	lut_sub lut_14565 ({g608, g1174, g1175, g1177}, g1178);
	defparam lut_14565.LUT_SIZE = 4;
	defparam lut_14565.mask = 16'h4000;

	lut_sub lut_14572 ({i_8_, g108, g630, g980}, g1179);
	defparam lut_14572.LUT_SIZE = 4;
	defparam lut_14572.mask = 16'h000b;

	lut_sub lut_14583 ({g47, g101, g172, g142, g1179}, g1180);
	defparam lut_14583.LUT_SIZE = 5;
	defparam lut_14583.mask = 32'haa80aa00;

	lut_sub lut_14598 ({i_14_, i_12_, i_13_, g102, g136, g115}, g1181);
	defparam lut_14598.LUT_SIZE = 6;
	defparam lut_14598.mask = 64'h2200323232300030;

	lut_sub lut_14620 ({g1050, g1071, g1040, g1066}, g1182);
	defparam lut_14620.LUT_SIZE = 4;
	defparam lut_14620.mask = 16'h8000;

	lut_sub lut_14628 ({g151, g1127, g1099, g1132}, g1183);
	defparam lut_14628.LUT_SIZE = 4;
	defparam lut_14628.mask = 16'h00df;

	lut_sub lut_14642 ({i_8_, g100, g195, g105, g532}, g1184);
	defparam lut_14642.LUT_SIZE = 5;
	defparam lut_14642.mask = 32'ha0a0a080;

	lut_sub lut_14655 ({g20, g98, g111}, g1185);
	defparam lut_14655.LUT_SIZE = 3;
	defparam lut_14655.mask = 8'h10;

	lut_sub lut_14664 ({i_8_, g100, g112, g1185, g835, g1001}, g1186);
	defparam lut_14664.LUT_SIZE = 6;
	defparam lut_14664.mask = 64'hf050f050f0503010;

	lut_sub lut_14693 ({g101, g1019, g1087, g1184, g1186}, g1187);
	defparam lut_14693.LUT_SIZE = 5;
	defparam lut_14693.mask = 32'h50500010;

	lut_sub lut_14707 ({g1098, g1180, g1181, g1182, g1183, g1187}, g1188);
	defparam lut_14707.LUT_SIZE = 6;
	defparam lut_14707.mask = 64'h0000040000000000;

	lut_sub lut_14717 ({g1147, g1156, g1167, g1173, g1178, g1188}, g1189);
	defparam lut_14717.LUT_SIZE = 6;
	defparam lut_14717.mask = 64'h0000000100000000;

	lut_sub lut_14727 ({g73, g420, g490, g664, g1145, g1189}, o_16_);
	defparam lut_14727.LUT_SIZE = 6;
	defparam lut_14727.mask = 64'h00000000fffffffe;

	lut_sub lut_14764 ({i_14_, i_12_, i_13_, g104, g109, g124}, g1191);
	defparam lut_14764.LUT_SIZE = 6;
	defparam lut_14764.mask = 64'h1103131313131103;

	lut_sub lut_14789 ({g6, i_15_, i_14_, i_12_, i_13_, g145}, g1192);
	defparam lut_14789.LUT_SIZE = 6;
	defparam lut_14789.mask = 64'h0000000004510554;

	lut_sub lut_14806 ({g10, g99, g109, g92, g468}, g1193);
	defparam lut_14806.LUT_SIZE = 5;
	defparam lut_14806.mask = 32'hff11f010;

	lut_sub lut_14830 ({g101, g224, g467, g574, g1192, g1193}, g1194);
	defparam lut_14830.LUT_SIZE = 6;
	defparam lut_14830.mask = 64'h4444444400400000;

	lut_sub lut_14848 ({g932, g978, g1164, g1166, g1191, g1194}, g1195);
	defparam lut_14848.LUT_SIZE = 6;
	defparam lut_14848.mask = 64'h0000040000000000;

	lut_sub lut_14854 ({g1020, g1021}, g1196);
	defparam lut_14854.LUT_SIZE = 2;
	defparam lut_14854.mask = 4'b0100;

	lut_sub lut_14862 ({g21, g12, g134, g136}, g1197);
	defparam lut_14862.LUT_SIZE = 4;
	defparam lut_14862.mask = 16'hf8c8;

	lut_sub lut_14876 ({i_14_, i_12_, i_13_, g11, g22, g136}, g1198);
	defparam lut_14876.LUT_SIZE = 6;
	defparam lut_14876.mask = 64'h0511000500000511;

	lut_sub lut_14891 ({i_14_, i_12_, i_13_, g11, g22}, g1199);
	defparam lut_14891.LUT_SIZE = 5;
	defparam lut_14891.mask = 32'h75300070;

	lut_sub lut_14909 ({g112, g201, g530, g703, g908}, g1200);
	defparam lut_14909.LUT_SIZE = 5;
	defparam lut_14909.mask = 32'h0000ff7f;

	lut_sub lut_14930 ({g134, g1199, g1200}, g1201);
	defparam lut_14930.LUT_SIZE = 3;
	defparam lut_14930.mask = 8'ha8;

	lut_sub lut_14942 ({g134, g153, g506, g1197, g1198, g1201}, g1202);
	defparam lut_14942.LUT_SIZE = 6;
	defparam lut_14942.mask = 64'h0404000004000000;

	lut_sub lut_14953 ({g21, g109, g114, g605, g908}, g1203);
	defparam lut_14953.LUT_SIZE = 5;
	defparam lut_14953.mask = 32'hcc80cc00;

	lut_sub lut_14968 ({i_8_, g108, g530, g703}, g1204);
	defparam lut_14968.LUT_SIZE = 4;
	defparam lut_14968.mask = 16'h0503;

	lut_sub lut_14980 ({i_8_, g12, g206, g108, g226, g506}, g1205);
	defparam lut_14980.LUT_SIZE = 6;
	defparam lut_14980.mask = 64'h0d0d0d0d0f0c0f0f;

	lut_sub lut_15013 ({g1143, g1203, g1204, g1205}, g1206);
	defparam lut_15013.LUT_SIZE = 4;
	defparam lut_15013.mask = 16'h0008;

	lut_sub lut_15021 ({g562, g804, g1148, g1149}, g1207);
	defparam lut_15021.LUT_SIZE = 4;
	defparam lut_15021.mask = 16'h8000;

	lut_sub lut_15028 ({g136, g177, g1176}, g1208);
	defparam lut_15028.LUT_SIZE = 3;
	defparam lut_15028.mask = 8'ha8;

	lut_sub lut_15037 ({i_8_, i_6_, i_7_, g87, g424, g530}, g1209);
	defparam lut_15037.LUT_SIZE = 6;
	defparam lut_15037.mask = 64'h0500000305000000;

	lut_sub lut_15051 ({g151, g201, g423, g703, g1209}, g1210);
	defparam lut_15051.LUT_SIZE = 5;
	defparam lut_15051.mask = 32'ha0a80088;

	lut_sub lut_15066 ({g134, g89, g118, g593, g1096}, g1211);
	defparam lut_15066.LUT_SIZE = 5;
	defparam lut_15066.mask = 32'h51f11131;

	lut_sub lut_15084 ({g99, g201}, g1212);
	defparam lut_15084.LUT_SIZE = 2;
	defparam lut_15084.mask = 4'b0010;

	lut_sub lut_15090 ({g118, g506}, g1213);
	defparam lut_15090.LUT_SIZE = 2;
	defparam lut_15090.mask = 4'b0001;

	lut_sub lut_15096 ({g134, g464}, g1214);
	defparam lut_15096.LUT_SIZE = 2;
	defparam lut_15096.mask = 4'b0010;

	lut_sub lut_15104 ({i_8_, g23, g206, g135, g226}, g1215);
	defparam lut_15104.LUT_SIZE = 5;
	defparam lut_15104.mask = 32'h00003233;

	lut_sub lut_15120 ({g297, g1212, g238, g1213, g1214, g1215}, g1216);
	defparam lut_15120.LUT_SIZE = 6;
	defparam lut_15120.mask = 64'h8080000080000000;

	lut_sub lut_15132 ({g1207, g1208, g1210, g1607, g1211, g1216}, g1217);
	defparam lut_15132.LUT_SIZE = 6;
	defparam lut_15132.mask = 64'h0000000000000001;

	lut_sub lut_15139 ({i_14_, i_12_, i_13_, g11, g22, g118}, g1218);
	defparam lut_15139.LUT_SIZE = 6;
	defparam lut_15139.mask = 64'h0515110000001511;

	lut_sub lut_15160 ({g23, g206, g118, g260, g464, g1218}, g1219);
	defparam lut_15160.LUT_SIZE = 6;
	defparam lut_15160.mask = 64'ha000a020a000a000;

	lut_sub lut_15177 ({g1095, g1098, g1100, g1541, g1219}, g1220);
	defparam lut_15177.LUT_SIZE = 5;
	defparam lut_15177.mask = 32'h10000000;

	lut_sub lut_15187 ({g1196, g1045, g1202, g1206, g1217, g1220}, g1221);
	defparam lut_15187.LUT_SIZE = 6;
	defparam lut_15187.mask = 64'h0000000000000001;

	lut_sub lut_15193 ({i_8_, g135, g224}, g1222);
	defparam lut_15193.LUT_SIZE = 3;
	defparam lut_15193.mask = 8'h01;

	lut_sub lut_15199 ({g10, g134}, g1223);
	defparam lut_15199.LUT_SIZE = 2;
	defparam lut_15199.mask = 4'b0001;

	lut_sub lut_15205 ({g66, g118}, g1224);
	defparam lut_15205.LUT_SIZE = 2;
	defparam lut_15205.mask = 4'b0001;

	lut_sub lut_15213 ({i_8_, g134, g221, g135, g127}, g1225);
	defparam lut_15213.LUT_SIZE = 5;
	defparam lut_15213.mask = 32'h00f022f2;

	lut_sub lut_15231 ({i_8_, g134, g135, g90, g467}, g1226);
	defparam lut_15231.LUT_SIZE = 5;
	defparam lut_15231.mask = 32'h00cc0ece;

	lut_sub lut_15252 ({g370, g1222, g1223, g1224, g1225, g1226}, g1227);
	defparam lut_15252.LUT_SIZE = 6;
	defparam lut_15252.mask = 64'h8000000000000000;

	lut_sub lut_15261 ({g8, i_8_, g135, g528, g817, g1001}, g1228);
	defparam lut_15261.LUT_SIZE = 6;
	defparam lut_15261.mask = 64'h00ff00f300fa00f3;

	lut_sub lut_15296 ({g608, g1174, g1175, g1177, g1227, g1228}, g1229);
	defparam lut_15296.LUT_SIZE = 6;
	defparam lut_15296.mask = 64'h0200000000000000;

	lut_sub lut_15305 ({g145, g187, g534, g702, g881}, g1230);
	defparam lut_15305.LUT_SIZE = 5;
	defparam lut_15305.mask = 32'h00007fff;

	lut_sub lut_15325 ({g6, i_15_, i_14_, i_12_, i_13_, g109}, g1231);
	defparam lut_15325.LUT_SIZE = 6;
	defparam lut_15325.mask = 64'h0000000004504504;

	lut_sub lut_15339 ({i_8_, g46, g209, g531, g1060}, g1232);
	defparam lut_15339.LUT_SIZE = 5;
	defparam lut_15339.mask = 32'haa00c0c0;

	lut_sub lut_15354 ({i_8_, g206, g108, g127, g561}, g1233);
	defparam lut_15354.LUT_SIZE = 5;
	defparam lut_15354.mask = 32'h0f0d0000;

	lut_sub lut_15369 ({i_8_, g23, g12, g108, g1232, g1233}, g1234);
	defparam lut_15369.LUT_SIZE = 6;
	defparam lut_15369.mask = 64'ha2a0a0a0a2a2a2a2;

	lut_sub lut_15399 ({g1628, g1622, g1104, g1230, g1231, g1234}, g1235);
	defparam lut_15399.LUT_SIZE = 6;
	defparam lut_15399.mask = 64'h0000000000000040;

	lut_sub lut_15405 ({g6, i_15_, i_14_, i_12_, i_13_, g112}, g1236);
	defparam lut_15405.LUT_SIZE = 6;
	defparam lut_15405.mask = 64'h0000000004551555;

	lut_sub lut_15422 ({g6, i_15_, i_14_, i_12_, i_13_, g118}, g1237);
	defparam lut_15422.LUT_SIZE = 6;
	defparam lut_15422.mask = 64'h0000000015555554;

	lut_sub lut_15441 ({g1236, g1237}, g1238);
	defparam lut_15441.LUT_SIZE = 2;
	defparam lut_15441.mask = 4'b1000;

	lut_sub lut_15450 ({g109, g529, g1721, g537, g1238}, g1239);
	defparam lut_15450.LUT_SIZE = 5;
	defparam lut_15450.mask = 32'h01010001;

	lut_sub lut_15458 ({g46, g243}, g1240);
	defparam lut_15458.LUT_SIZE = 2;
	defparam lut_15458.mask = 4'b0001;

	lut_sub lut_15468 ({g185, g151, g187, g429, g1033, g1240}, g1241);
	defparam lut_15468.LUT_SIZE = 6;
	defparam lut_15468.mask = 64'h8880000088808880;

	lut_sub lut_15484 ({g8, g197, g90, g424}, g1242);
	defparam lut_15484.LUT_SIZE = 4;
	defparam lut_15484.mask = 16'h0020;

	lut_sub lut_15491 ({i_8_, g108, g185, g231}, g1243);
	defparam lut_15491.LUT_SIZE = 4;
	defparam lut_15491.mask = 16'h000e;

	lut_sub lut_15502 ({g66, g330, g423, g1242, g1243}, g1244);
	defparam lut_15502.LUT_SIZE = 5;
	defparam lut_15502.mask = 32'ha2a200a2;

	lut_sub lut_15517 ({i_8_, g88, g108, g531}, g1245);
	defparam lut_15517.LUT_SIZE = 4;
	defparam lut_15517.mask = 16'h1105;

	lut_sub lut_15528 ({g227, g209, g746, g349}, g1246);
	defparam lut_15528.LUT_SIZE = 4;
	defparam lut_15528.mask = 16'h0357;

	lut_sub lut_15541 ({g12, g46, g99}, g1247);
	defparam lut_15541.LUT_SIZE = 3;
	defparam lut_15541.mask = 8'h15;

	lut_sub lut_15552 ({g134, g118, g231, g534, g478}, g1248);
	defparam lut_15552.LUT_SIZE = 5;
	defparam lut_15552.mask = 32'hff080f08;

	lut_sub lut_15574 ({g972, g1245, g1246, g1247, g1248}, g1249);
	defparam lut_15574.LUT_SIZE = 5;
	defparam lut_15574.mask = 32'h40000000;

	lut_sub lut_15584 ({g766, g1025, g1054, g1241, g1244, g1249}, g1250);
	defparam lut_15584.LUT_SIZE = 6;
	defparam lut_15584.mask = 64'h0000000000000001;

	lut_sub lut_15592 ({g10, g45, g221, g534}, g1251);
	defparam lut_15592.LUT_SIZE = 4;
	defparam lut_15592.mask = 16'h2000;

	lut_sub lut_15600 ({g134, g224, g467, g817}, g1252);
	defparam lut_15600.LUT_SIZE = 4;
	defparam lut_15600.mask = 16'h00df;

	lut_sub lut_15614 ({g214, g946, g1251, g1252}, g1253);
	defparam lut_15614.LUT_SIZE = 4;
	defparam lut_15614.mask = 16'ha020;

	lut_sub lut_15622 ({i_11_, i_9_, i_10_, g326, g238}, g1254);
	defparam lut_15622.LUT_SIZE = 5;
	defparam lut_15622.mask = 32'h00010010;

	lut_sub lut_15628 ({i_14_, i_12_, i_13_, g122}, g1255);
	defparam lut_15628.LUT_SIZE = 4;
	defparam lut_15628.mask = 16'h2002;

	lut_sub lut_15638 ({g109, g186, g330, g544, g1255}, g1256);
	defparam lut_15638.LUT_SIZE = 5;
	defparam lut_15638.mask = 32'h3f332222;

	lut_sub lut_15661 ({g242, g1253, g1047, g1051, g1254, g1256}, g1257);
	defparam lut_15661.LUT_SIZE = 6;
	defparam lut_15661.mask = 64'h0000000000000004;

	lut_sub lut_15671 ({g890, g1229, g1235, g1239, g1250, g1257}, g1258);
	defparam lut_15671.LUT_SIZE = 6;
	defparam lut_15671.mask = 64'h0000000000000001;

	lut_sub lut_15678 ({g1065, g1158, g1163}, g1259);
	defparam lut_15678.LUT_SIZE = 3;
	defparam lut_15678.mask = 8'h40;

	lut_sub lut_15685 ({g187, g534, g702}, g1260);
	defparam lut_15685.LUT_SIZE = 3;
	defparam lut_15685.mask = 8'h80;

	lut_sub lut_15693 ({g89, g109, g1099, g1260}, g1261);
	defparam lut_15693.LUT_SIZE = 4;
	defparam lut_15693.mask = 16'hce0a;

	lut_sub lut_15708 ({i_8_, g134, g135, g187, g534, g702}, g1262);
	defparam lut_15708.LUT_SIZE = 6;
	defparam lut_15708.mask = 64'hffff8080ffc08080;

	lut_sub lut_15746 ({g136, g231, g478, g922, g1262}, g1263);
	defparam lut_15746.LUT_SIZE = 5;
	defparam lut_15746.mask = 32'h44440040;

	lut_sub lut_15760 ({g134, g99, g105, g837, g696, g702}, g1264);
	defparam lut_15760.LUT_SIZE = 6;
	defparam lut_15760.mask = 64'hffffaaaa03000200;

	lut_sub lut_15796 ({g945, g1063, g1261, g1263, g1133, g1264}, g1265);
	defparam lut_15796.LUT_SIZE = 6;
	defparam lut_15796.mask = 64'h0000000004000000;

	lut_sub lut_15802 ({g101, g1184}, g1266);
	defparam lut_15802.LUT_SIZE = 2;
	defparam lut_15802.mask = 4'b0010;

	lut_sub lut_15810 ({g99, g195, g105, g696}, g1267);
	defparam lut_15810.LUT_SIZE = 4;
	defparam lut_15810.mask = 16'h00bf;

	lut_sub lut_15825 ({g99, g101, g573, g837, g1267}, g1268);
	defparam lut_15825.LUT_SIZE = 5;
	defparam lut_15825.mask = 32'ha0202020;

	lut_sub lut_15836 ({i_14_, i_12_, i_13_, g104, g112, g124}, g1269);
	defparam lut_15836.LUT_SIZE = 6;
	defparam lut_15836.mask = 64'hfca0f0a0a0f0fff0;

	lut_sub lut_15874 ({i_8_, g495, g982, g1269}, g1270);
	defparam lut_15874.LUT_SIZE = 4;
	defparam lut_15874.mask = 16'h0a08;

	lut_sub lut_15883 ({i_14_, i_12_, i_13_, g118, g112, g124}, g1271);
	defparam lut_15883.LUT_SIZE = 6;
	defparam lut_15883.mask = 64'h0500050000111111;

	lut_sub lut_15901 ({i_11_, g113, g112, g187, g236, g1271}, g1272);
	defparam lut_15901.LUT_SIZE = 6;
	defparam lut_15901.mask = 64'haaa0aaa0aaa08880;

	lut_sub lut_15930 ({g931, g1266, g1268, g1270, g1272}, g1273);
	defparam lut_15930.LUT_SIZE = 5;
	defparam lut_15930.mask = 32'h04000000;

	lut_sub lut_15937 ({i_14_, i_12_, i_13_, g119, g118, g122}, g1274);
	defparam lut_15937.LUT_SIZE = 6;
	defparam lut_15937.mask = 64'h2223232203232300;

	lut_sub lut_15960 ({i_11_, i_9_, i_10_, g236, g1274}, g1275);
	defparam lut_15960.LUT_SIZE = 5;
	defparam lut_15960.mask = 32'haaaaaa8a;

	lut_sub lut_15981 ({i_8_, g108, g216, g548}, g1276);
	defparam lut_15981.LUT_SIZE = 4;
	defparam lut_15981.mask = 16'h0507;

	lut_sub lut_15993 ({i_8_, g181, g108, g123, g485}, g1277);
	defparam lut_15993.LUT_SIZE = 5;
	defparam lut_15993.mask = 32'h070f050f;

	lut_sub lut_16014 ({i_8_, g108, g670, g671, g1276, g1277}, g1278);
	defparam lut_16014.LUT_SIZE = 6;
	defparam lut_16014.mask = 64'h8888808088888000;

	lut_sub lut_16033 ({i_8_, g108, g216, g120, g123, g670}, g1279);
	defparam lut_16033.LUT_SIZE = 6;
	defparam lut_16033.mask = 64'h0000f5ff0000f3f3;

	lut_sub lut_16064 ({g108, g349}, g1280);
	defparam lut_16064.LUT_SIZE = 2;
	defparam lut_16064.mask = 4'b0001;

	lut_sub lut_16073 ({g101, g835, g670, g887, g1280}, g1281);
	defparam lut_16073.LUT_SIZE = 5;
	defparam lut_16073.mask = 32'haaaa0020;

	lut_sub lut_16088 ({i_8_, g108, g626, g895}, g1282);
	defparam lut_16088.LUT_SIZE = 4;
	defparam lut_16088.mask = 16'h0d0c;

	lut_sub lut_16102 ({g657, g1275, g1278, g1279, g1281, g1282}, g1283);
	defparam lut_16102.LUT_SIZE = 6;
	defparam lut_16102.mask = 64'h0000000000000020;

	lut_sub lut_16110 ({i_8_, g88, g120, g626, g1048}, g1284);
	defparam lut_16110.LUT_SIZE = 5;
	defparam lut_16110.mask = 32'h00fd0000;

	lut_sub lut_16125 ({g101, g136, g187, g670, g1284}, g1285);
	defparam lut_16125.LUT_SIZE = 5;
	defparam lut_16125.mask = 32'haa88a080;

	lut_sub lut_16140 ({i_14_, i_12_, i_13_, g149, g119, g122}, g1286);
	defparam lut_16140.LUT_SIZE = 6;
	defparam lut_16140.mask = 64'h0000000b0a0a0a0b;

	lut_sub lut_16161 ({g277, g214, g613, g540, g895, g1286}, g1287);
	defparam lut_16161.LUT_SIZE = 6;
	defparam lut_16161.mask = 64'h00800080aaaa8080;

	lut_sub lut_16178 ({g988, g1022}, g1288);
	defparam lut_16178.LUT_SIZE = 2;
	defparam lut_16178.mask = 4'b1000;

	lut_sub lut_16184 ({i_8_, g108, g895}, g1289);
	defparam lut_16184.LUT_SIZE = 3;
	defparam lut_16184.mask = 8'h01;

	lut_sub lut_16190 ({g134, g1161}, g1290);
	defparam lut_16190.LUT_SIZE = 2;
	defparam lut_16190.mask = 4'b0010;

	lut_sub lut_16197 ({g183, g423, g704}, g1291);
	defparam lut_16197.LUT_SIZE = 3;
	defparam lut_16197.mask = 8'h13;

	lut_sub lut_16206 ({g134, g118, g548}, g1292);
	defparam lut_16206.LUT_SIZE = 3;
	defparam lut_16206.mask = 8'h15;

	lut_sub lut_16216 ({g112, g323, g349, g481}, g1293);
	defparam lut_16216.LUT_SIZE = 4;
	defparam lut_16216.mask = 16'hf454;

	lut_sub lut_16233 ({g491, g1289, g1290, g1291, g1292, g1293}, g1294);
	defparam lut_16233.LUT_SIZE = 6;
	defparam lut_16233.mask = 64'h0000000040000000;

	lut_sub lut_16243 ({g1150, g1129, g1285, g1287, g1288, g1294}, g1295);
	defparam lut_16243.LUT_SIZE = 6;
	defparam lut_16243.mask = 64'h0000000100000000;

	lut_sub lut_16252 ({g112, g349, g540, g704, g895}, g1296);
	defparam lut_16252.LUT_SIZE = 5;
	defparam lut_16252.mask = 32'h00007fff;

	lut_sub lut_16275 ({g134, g136, g120, g123, g1296}, g1297);
	defparam lut_16275.LUT_SIZE = 5;
	defparam lut_16275.mask = 32'haa0a8808;

	lut_sub lut_16290 ({g136, g349, g540}, g1298);
	defparam lut_16290.LUT_SIZE = 3;
	defparam lut_16290.mask = 8'h07;

	lut_sub lut_16299 ({i_14_, i_12_, i_13_, g119, g136, g122}, g1299);
	defparam lut_16299.LUT_SIZE = 6;
	defparam lut_16299.mask = 64'h2300232323000003;

	lut_sub lut_16321 ({g760, g1297, g1298, g1596, g1299}, g1300);
	defparam lut_16321.LUT_SIZE = 5;
	defparam lut_16321.mask = 32'h00200000;

	lut_sub lut_16331 ({g1259, g1265, g1273, g1283, g1295, g1300}, g1301);
	defparam lut_16331.LUT_SIZE = 6;
	defparam lut_16331.mask = 64'h0000000000000001;

	lut_sub lut_16341 ({g73, g1156, g1195, g1221, g1258, g1301}, o_17_);
	defparam lut_16341.LUT_SIZE = 6;
	defparam lut_16341.mask = 64'h00000000fffffffe;

	lut_sub lut_16377 ({g1265, g1273}, g1303);
	defparam lut_16377.LUT_SIZE = 2;
	defparam lut_16377.mask = 4'b0001;

	lut_sub lut_16383 ({i_14_, i_12_, i_13_, g102, g115}, g1304);
	defparam lut_16383.LUT_SIZE = 5;
	defparam lut_16383.mask = 32'h0ceccea0;

	lut_sub lut_16405 ({g118, g187, g534, g980, g1304}, g1305);
	defparam lut_16405.LUT_SIZE = 5;
	defparam lut_16405.mask = 32'h0000dfff;

	lut_sub lut_16427 ({g546, g477, g706, g979}, g1306);
	defparam lut_16427.LUT_SIZE = 4;
	defparam lut_16427.mask = 16'h0400;

	lut_sub lut_16435 ({g109, g1179, g1243, g1306}, g1307);
	defparam lut_16435.LUT_SIZE = 4;
	defparam lut_16435.mask = 16'hc040;

	lut_sub lut_16446 ({i_8_, g108, g193, g232, g173, g103}, g1308);
	defparam lut_16446.LUT_SIZE = 6;
	defparam lut_16446.mask = 64'h0000bfff00000000;

	lut_sub lut_16469 ({i_8_, g264, g108, g696, g907, g1308}, g1309);
	defparam lut_16469.LUT_SIZE = 6;
	defparam lut_16469.mask = 64'haaaaaa00aa08aa08;

	lut_sub lut_16497 ({g220, g112, g827}, g1310);
	defparam lut_16497.LUT_SIZE = 3;
	defparam lut_16497.mask = 8'h23;

	lut_sub lut_16508 ({g48, g102, g112, g182, g115}, g1311);
	defparam lut_16508.LUT_SIZE = 5;
	defparam lut_16508.mask = 32'h0f0a0302;

	lut_sub lut_16524 ({g112, g675, g672, g706}, g1312);
	defparam lut_16524.LUT_SIZE = 4;
	defparam lut_16524.mask = 16'h007f;

	lut_sub lut_16539 ({g118, g231, g478, g487, g675}, g1313);
	defparam lut_16539.LUT_SIZE = 5;
	defparam lut_16539.mask = 32'h0000ff7f;

	lut_sub lut_16562 ({g658, g1310, g1311, g1312, g1313}, g1314);
	defparam lut_16562.LUT_SIZE = 5;
	defparam lut_16562.mask = 32'h80000000;

	lut_sub lut_16569 ({g173, g546, g907}, g1315);
	defparam lut_16569.LUT_SIZE = 3;
	defparam lut_16569.mask = 8'h80;

	lut_sub lut_16576 ({g550, g630, g696}, g1316);
	defparam lut_16576.LUT_SIZE = 3;
	defparam lut_16576.mask = 8'h40;

	lut_sub lut_16585 ({g112, g495, g1153, g1315, g1316}, g1317);
	defparam lut_16585.LUT_SIZE = 5;
	defparam lut_16585.mask = 32'hf0305010;

	lut_sub lut_16603 ({g1155, g1305, g1307, g1309, g1314, g1317}, g1318);
	defparam lut_16603.LUT_SIZE = 6;
	defparam lut_16603.mask = 64'h0001000000000000;

	lut_sub lut_16613 ({g101, g185, g173, g914, g882, g1170}, g1319);
	defparam lut_16613.LUT_SIZE = 6;
	defparam lut_16613.mask = 64'h00000000fffffeff;

	lut_sub lut_16651 ({g99, g173, g103, g929}, g1320);
	defparam lut_16651.LUT_SIZE = 4;
	defparam lut_16651.mask = 16'haa20;

	lut_sub lut_16663 ({g570, g1010, g1319, g1320}, g1321);
	defparam lut_16663.LUT_SIZE = 4;
	defparam lut_16663.mask = 16'h0400;

	lut_sub lut_16672 ({g136, g193, g696, g672, g702}, g1322);
	defparam lut_16672.LUT_SIZE = 5;
	defparam lut_16672.mask = 32'h0000f7ff;

	lut_sub lut_16692 ({i_14_, i_12_, i_13_, g102, g115}, g1323);
	defparam lut_16692.LUT_SIZE = 5;
	defparam lut_16692.mask = 32'h35511511;

	lut_sub lut_16711 ({g134, g533, g779, g1323}, g1324);
	defparam lut_16711.LUT_SIZE = 4;
	defparam lut_16711.mask = 16'hc040;

	lut_sub lut_16721 ({g134, g136, g231, g232}, g1325);
	defparam lut_16721.LUT_SIZE = 4;
	defparam lut_16721.mask = 16'h05cd;

	lut_sub lut_16734 ({i_8_, g135, g907, g881}, g1326);
	defparam lut_16734.LUT_SIZE = 4;
	defparam lut_16734.mask = 16'h0007;

	lut_sub lut_16745 ({g134, g220, g103, g105, g837}, g1327);
	defparam lut_16745.LUT_SIZE = 5;
	defparam lut_16745.mask = 32'h0000fbff;

	lut_sub lut_16769 ({g136, g477, g630, g706, g1326, g1327}, g1328);
	defparam lut_16769.LUT_SIZE = 6;
	defparam lut_16769.mask = 64'h8888888800008000;

	lut_sub lut_16787 ({g1152, g1181, g1322, g1324, g1325, g1328}, g1329);
	defparam lut_16787.LUT_SIZE = 6;
	defparam lut_16787.mask = 64'h0400000000000000;

	lut_sub lut_16796 ({g145, g269, g1082, g1191, g1589}, g1330);
	defparam lut_16796.LUT_SIZE = 5;
	defparam lut_16796.mask = 32'h44444000;

	lut_sub lut_16806 ({g89, g1103}, g1331);
	defparam lut_16806.LUT_SIZE = 2;
	defparam lut_16806.mask = 4'b1000;

	lut_sub lut_16815 ({g323, g195, g105, g532, g921}, g1332);
	defparam lut_16815.LUT_SIZE = 5;
	defparam lut_16815.mask = 32'h0000bfff;

	lut_sub lut_16836 ({i_8_, g88, g115, g711}, g1333);
	defparam lut_16836.LUT_SIZE = 4;
	defparam lut_16836.mask = 16'h0004;

	lut_sub lut_16844 ({g118, g232, g423, g630}, g1334);
	defparam lut_16844.LUT_SIZE = 4;
	defparam lut_16844.mask = 16'h0357;

	lut_sub lut_16858 ({g88, g103, g423, g1076}, g1335);
	defparam lut_16858.LUT_SIZE = 4;
	defparam lut_16858.mask = 16'hce8a;

	lut_sub lut_16874 ({i_8_, g88, g264, g103, g423, g675}, g1336);
	defparam lut_16874.LUT_SIZE = 6;
	defparam lut_16874.mask = 64'h111111111111f5ff;

	lut_sub lut_16909 ({g323, g837, g1333, g1334, g1335, g1336}, g1337);
	defparam lut_16909.LUT_SIZE = 6;
	defparam lut_16909.mask = 64'h2000200000002000;

	lut_sub lut_16918 ({i_8_, g88, g423, g640}, g1338);
	defparam lut_16918.LUT_SIZE = 4;
	defparam lut_16918.mask = 16'h222a;

	lut_sub lut_16932 ({g145, g187, g534, g702, g881, g1338}, g1339);
	defparam lut_16932.LUT_SIZE = 6;
	defparam lut_16932.mask = 64'haaaaaaaa80000000;

	lut_sub lut_16958 ({g997, g1331, g1616, g1332, g1337, g1339}, g1340);
	defparam lut_16958.LUT_SIZE = 6;
	defparam lut_16958.mask = 64'h0000000000100000;

	lut_sub lut_16968 ({g1092, g1318, g1321, g1329, g1330, g1340}, g1341);
	defparam lut_16968.LUT_SIZE = 6;
	defparam lut_16968.mask = 64'h0000000000000001;

	lut_sub lut_16976 ({g44, g43, g191, g530}, g1342);
	defparam lut_16976.LUT_SIZE = 4;
	defparam lut_16976.mask = 16'h8000;

	lut_sub lut_16984 ({i_8_, g108, g142, g117, g1342}, g1343);
	defparam lut_16984.LUT_SIZE = 5;
	defparam lut_16984.mask = 32'h00bf003f;

	lut_sub lut_17003 ({i_8_, g19, g108, g462}, g1344);
	defparam lut_17003.LUT_SIZE = 4;
	defparam lut_17003.mask = 16'h0322;

	lut_sub lut_17012 ({i_14_, i_12_, i_13_, i_8_, g15, g108}, g1345);
	defparam lut_17012.LUT_SIZE = 6;
	defparam lut_17012.mask = 64'h0400444444000000;

	lut_sub lut_17028 ({g109, g201, g172, g339, g1344, g1345}, g1346);
	defparam lut_17028.LUT_SIZE = 6;
	defparam lut_17028.mask = 64'h8888888800008000;

	lut_sub lut_17046 ({g145, g497, g668, g1122, g1343, g1346}, g1347);
	defparam lut_17046.LUT_SIZE = 6;
	defparam lut_17046.mask = 64'h4400000004000000;

	lut_sub lut_17056 ({g134, g136, g142, g465}, g1348);
	defparam lut_17056.LUT_SIZE = 4;
	defparam lut_17056.mask = 16'h0a3b;

	lut_sub lut_17069 ({g134, g222, g530}, g1349);
	defparam lut_17069.LUT_SIZE = 3;
	defparam lut_17069.mask = 8'h07;

	lut_sub lut_17080 ({g43, g135, g781, g1122, g1349}, g1350);
	defparam lut_17080.LUT_SIZE = 5;
	defparam lut_17080.mask = 32'ha020a000;

	lut_sub lut_17093 ({g19, g16, g136, g222, g399}, g1351);
	defparam lut_17093.LUT_SIZE = 5;
	defparam lut_17093.mask = 32'h0f0b0f0f;

	lut_sub lut_17116 ({g136, g339, g1348, g1350, g1351}, g1352);
	defparam lut_17116.LUT_SIZE = 5;
	defparam lut_17116.mask = 32'h20202000;

	lut_sub lut_17128 ({g149, g191, g338, g340, g399, g361}, g1353);
	defparam lut_17128.LUT_SIZE = 6;
	defparam lut_17128.mask = 64'h20a000a020a00000;

	lut_sub lut_17145 ({g804, g805, g1673, g810, g1666, g1353}, g1354);
	defparam lut_17145.LUT_SIZE = 6;
	defparam lut_17145.mask = 64'h0001000000000000;

	lut_sub lut_17153 ({g19, g118, g117, g462}, g1355);
	defparam lut_17153.LUT_SIZE = 4;
	defparam lut_17153.mask = 16'h0b0f;

	lut_sub lut_17166 ({g112, g222, g807}, g1356);
	defparam lut_17166.LUT_SIZE = 3;
	defparam lut_17166.mask = 8'h0b;

	lut_sub lut_17178 ({g19, g16, g112, g142, g339, g465}, g1357);
	defparam lut_17178.LUT_SIZE = 6;
	defparam lut_17178.mask = 64'h00ff00bf00ff00ff;

	lut_sub lut_17218 ({g16, g118, g378, g1355, g1356, g1357}, g1358);
	defparam lut_17218.LUT_SIZE = 6;
	defparam lut_17218.mask = 64'h8000000080008000;

	lut_sub lut_17229 ({i_8_, g108, g201, g641, g703, g908}, g1359);
	defparam lut_17229.LUT_SIZE = 6;
	defparam lut_17229.mask = 64'h00000f0f0000ff77;

	lut_sub lut_17256 ({g996, g1359}, g1360);
	defparam lut_17256.LUT_SIZE = 2;
	defparam lut_17256.mask = 4'b0010;

	lut_sub lut_17262 ({g43, g641}, g1361);
	defparam lut_17262.LUT_SIZE = 2;
	defparam lut_17262.mask = 4'b1000;

	lut_sub lut_17270 ({g118, g186, g142, g898}, g1362);
	defparam lut_17270.LUT_SIZE = 4;
	defparam lut_17270.mask = 16'hf888;

	lut_sub lut_17284 ({g59, g44, g186, g495}, g1363);
	defparam lut_17284.LUT_SIZE = 4;
	defparam lut_17284.mask = 16'h070f;

	lut_sub lut_17300 ({g59, g146, g251, g1361, g1362, g1363}, g1364);
	defparam lut_17300.LUT_SIZE = 6;
	defparam lut_17300.mask = 64'h0202220202020202;

	lut_sub lut_17314 ({i_8_, g100, g201}, g1365);
	defparam lut_17314.LUT_SIZE = 3;
	defparam lut_17314.mask = 8'h02;

	lut_sub lut_17320 ({g134, g117}, g1366);
	defparam lut_17320.LUT_SIZE = 2;
	defparam lut_17320.mask = 4'b0001;

	lut_sub lut_17326 ({g20, g88}, g1367);
	defparam lut_17326.LUT_SIZE = 2;
	defparam lut_17326.mask = 4'b0100;

	lut_sub lut_17332 ({g186, g908}, g1368);
	defparam lut_17332.LUT_SIZE = 2;
	defparam lut_17332.mask = 4'b0001;

	lut_sub lut_17339 ({g98, g264, g111}, g1369);
	defparam lut_17339.LUT_SIZE = 3;
	defparam lut_17339.mask = 8'h01;

	lut_sub lut_17349 ({g1365, g1366, g1046, g1367, g1368, g1369}, g1370);
	defparam lut_17349.LUT_SIZE = 6;
	defparam lut_17349.mask = 64'h8000000000000000;

	lut_sub lut_17358 ({g15, g59, g112, g135, g461}, g1371);
	defparam lut_17358.LUT_SIZE = 5;
	defparam lut_17358.mask = 32'h15550000;

	lut_sub lut_17373 ({g375, g164, g1371, g1034, g1035}, g1372);
	defparam lut_17373.LUT_SIZE = 5;
	defparam lut_17373.mask = 32'h80808000;

	lut_sub lut_17385 ({g1358, g1360, g1580, g1364, g1370, g1372}, g1373);
	defparam lut_17385.LUT_SIZE = 6;
	defparam lut_17385.mask = 64'h0000000000000001;

	lut_sub lut_17393 ({g23, g12, g109, g1233}, g1374);
	defparam lut_17393.LUT_SIZE = 4;
	defparam lut_17393.mask = 16'ha888;

	lut_sub lut_17406 ({g31, g19, g87, g339, g465}, g1375);
	defparam lut_17406.LUT_SIZE = 5;
	defparam lut_17406.mask = 32'h00000b0f;

	lut_sub lut_17420 ({g172, g214, g495, g1375}, g1376);
	defparam lut_17420.LUT_SIZE = 4;
	defparam lut_17420.mask = 16'haa80;

	lut_sub lut_17432 ({g277, g339, g465, g1376}, g1377);
	defparam lut_17432.LUT_SIZE = 4;
	defparam lut_17432.mask = 16'h1055;

	lut_sub lut_17445 ({i_8_, g19, g16, g88, g231, g262}, g1378);
	defparam lut_17445.LUT_SIZE = 6;
	defparam lut_17445.mask = 64'haaaaaaaaa0a2a0a0;

	lut_sub lut_17478 ({g101, g151, g530, g636, g1378}, g1379);
	defparam lut_17478.LUT_SIZE = 5;
	defparam lut_17478.mask = 32'h55115010;

	lut_sub lut_17494 ({i_8_, g16, g108, g339, g636}, g1380);
	defparam lut_17494.LUT_SIZE = 5;
	defparam lut_17494.mask = 32'h0f000b0b;

	lut_sub lut_17513 ({g1374, g1377, g1379, g1380, g1068, g1131}, g1381);
	defparam lut_17513.LUT_SIZE = 6;
	defparam lut_17513.mask = 64'h0000000000000010;

	lut_sub lut_17523 ({g976, g1347, g1352, g1354, g1373, g1381}, g1382);
	defparam lut_17523.LUT_SIZE = 6;
	defparam lut_17523.mask = 64'h0000000000000001;

	lut_sub lut_17533 ({g73, g985, g1221, g1303, g1341, g1382}, o_18_);
	defparam lut_17533.LUT_SIZE = 6;
	defparam lut_17533.mask = 64'h00000000fffffffe;

	lut_sub lut_17571 ({g203, g678, g669, g818}, g1384);
	defparam lut_17571.LUT_SIZE = 4;
	defparam lut_17571.mask = 16'h0100;

	lut_sub lut_17579 ({g134, g304, g270, g136}, g1385);
	defparam lut_17579.LUT_SIZE = 4;
	defparam lut_17579.mask = 16'h444f;

	lut_sub lut_17592 ({g134, g94, g475}, g1386);
	defparam lut_17592.LUT_SIZE = 3;
	defparam lut_17592.mask = 8'h0b;

	lut_sub lut_17603 ({g136, g96, g474, g1385, g1386}, g1387);
	defparam lut_17603.LUT_SIZE = 5;
	defparam lut_17603.mask = 32'h88880080;

	lut_sub lut_17615 ({g109, g94, g96, g678}, g1388);
	defparam lut_17615.LUT_SIZE = 4;
	defparam lut_17615.mask = 16'h00ef;

	lut_sub lut_17628 ({i_8_, g108, g96, g986}, g1389);
	defparam lut_17628.LUT_SIZE = 4;
	defparam lut_17628.mask = 16'h050d;

	lut_sub lut_17642 ({g109, g203, g183, g268, g1255, g1389}, g1390);
	defparam lut_17642.LUT_SIZE = 6;
	defparam lut_17642.mask = 64'haaaaaaaa80000000;

	lut_sub lut_17664 ({i_14_, i_12_, i_13_, i_8_, g108, g93}, g1391);
	defparam lut_17664.LUT_SIZE = 6;
	defparam lut_17664.mask = 64'h0020000000000002;

	lut_sub lut_17674 ({g510, g1388, g1390, g1538, g1391}, g1392);
	defparam lut_17674.LUT_SIZE = 5;
	defparam lut_17674.mask = 32'h02000000;

	lut_sub lut_17682 ({g89, g135, g268, g495}, g1393);
	defparam lut_17682.LUT_SIZE = 4;
	defparam lut_17682.mask = 16'h3313;

	lut_sub lut_17694 ({g474, g495}, g1394);
	defparam lut_17694.LUT_SIZE = 2;
	defparam lut_17694.mask = 4'b0001;

	lut_sub lut_17701 ({i_8_, g270, g475, g495}, g1395);
	defparam lut_17701.LUT_SIZE = 4;
	defparam lut_17701.mask = 16'h4450;

	lut_sub lut_17712 ({g118, g270, g813, g495}, g1396);
	defparam lut_17712.LUT_SIZE = 4;
	defparam lut_17712.mask = 16'h11f1;

	lut_sub lut_17725 ({i_14_, i_12_, i_13_, g118, g112, g93}, g1397);
	defparam lut_17725.LUT_SIZE = 6;
	defparam lut_17725.mask = 64'h0a002a2200002a00;

	lut_sub lut_17744 ({g659, g682, g1394, g1395, g1396, g1397}, g1398);
	defparam lut_17744.LUT_SIZE = 6;
	defparam lut_17744.mask = 64'h8000000000000000;

	lut_sub lut_17753 ({g118, g423, g429, g556, g1048}, g1399);
	defparam lut_17753.LUT_SIZE = 5;
	defparam lut_17753.mask = 32'h04050c0d;

	lut_sub lut_17768 ({g983, g1393, g1398, g1399}, g1400);
	defparam lut_17768.LUT_SIZE = 4;
	defparam lut_17768.mask = 16'h0020;

	lut_sub lut_17777 ({g145, g268, g555, g474, g678}, g1401);
	defparam lut_17777.LUT_SIZE = 5;
	defparam lut_17777.mask = 32'h0000bfff;

	lut_sub lut_17800 ({g1002, g1003, g1004, g1005, g1401}, g1402);
	defparam lut_17800.LUT_SIZE = 5;
	defparam lut_17800.mask = 32'h80000000;

	lut_sub lut_17807 ({g118, g214, g756}, g1403);
	defparam lut_17807.LUT_SIZE = 3;
	defparam lut_17807.mask = 8'h15;

	lut_sub lut_17817 ({g7, g95, g461, g756}, g1404);
	defparam lut_17817.LUT_SIZE = 4;
	defparam lut_17817.mask = 16'ha8a0;

	lut_sub lut_17831 ({g99, g330, g251, g986, g1403, g1404}, g1405);
	defparam lut_17831.LUT_SIZE = 6;
	defparam lut_17831.mask = 64'h5550ddd05050d0d0;

	lut_sub lut_17864 ({g212, g213, g215, g217, g1036}, g1406);
	defparam lut_17864.LUT_SIZE = 5;
	defparam lut_17864.mask = 32'h88008808;

	lut_sub lut_17877 ({i_8_, g88, g212, g534, g555, g1099}, g1407);
	defparam lut_17877.LUT_SIZE = 6;
	defparam lut_17877.mask = 64'h330033333300bfaf;

	lut_sub lut_17913 ({g99, g88, g554, g895}, g1408);
	defparam lut_17913.LUT_SIZE = 4;
	defparam lut_17913.mask = 16'h0357;

	lut_sub lut_17929 ({g99, g101, g756, g991, g1042, g1408}, g1409);
	defparam lut_17929.LUT_SIZE = 6;
	defparam lut_17929.mask = 64'h8080800080008000;

	lut_sub lut_17943 ({g149, g338, g341, g556, g522, g476}, g1410);
	defparam lut_17943.LUT_SIZE = 6;
	defparam lut_17943.mask = 64'h0800aa0008008800;

	lut_sub lut_17959 ({i_8_, g100, g199, g120, g547, g574}, g1411);
	defparam lut_17959.LUT_SIZE = 6;
	defparam lut_17959.mask = 64'h000000000000fdff;

	lut_sub lut_17983 ({g1405, g1406, g1407, g1409, g1410, g1558}, g1412);
	defparam lut_17983.LUT_SIZE = 6;
	defparam lut_17983.mask = 64'h0000000000000200;

	lut_sub lut_17993 ({g527, g1110, g1059, g1400, g1402, g1412}, g1413);
	defparam lut_17993.LUT_SIZE = 6;
	defparam lut_17993.mask = 64'h0000000000000001;

	lut_sub lut_18003 ({g73, g1301, g1341, g1568, g1392, g1413}, o_19_);
	defparam lut_18003.LUT_SIZE = 6;
	defparam lut_18003.mask = 64'h00000000fffffffe;

	lut_sub lut_18040 ({g1305, g1314, g1317}, g1415);
	defparam lut_18040.LUT_SIZE = 3;
	defparam lut_18040.mask = 8'h10;

	lut_sub lut_18047 ({i_8_, g222, g531, g630}, g1416);
	defparam lut_18047.LUT_SIZE = 4;
	defparam lut_18047.mask = 16'h8000;

	lut_sub lut_18055 ({g246, g593, g678, g1416}, g1417);
	defparam lut_18055.LUT_SIZE = 4;
	defparam lut_18055.mask = 16'h0100;

	lut_sub lut_18064 ({g339, g613, g465, g506, g1417}, g1418);
	defparam lut_18064.LUT_SIZE = 5;
	defparam lut_18064.mask = 32'h00040000;

	lut_sub lut_18071 ({g6, i_15_, g7, g461}, g1419);
	defparam lut_18071.LUT_SIZE = 4;
	defparam lut_18071.mask = 16'h0070;

	lut_sub lut_18081 ({i_8_, g495, g1026, g1111, g1419}, g1420);
	defparam lut_18081.LUT_SIZE = 5;
	defparam lut_18081.mask = 32'h00ff00df;

	lut_sub lut_18103 ({g1112, g1113, g1418, g1420}, g1421);
	defparam lut_18103.LUT_SIZE = 4;
	defparam lut_18103.mask = 16'h5554;

	lut_sub lut_18116 ({g1238, g1270, g1272}, g1422);
	defparam lut_18116.LUT_SIZE = 3;
	defparam lut_18116.mask = 8'h04;

	lut_sub lut_18124 ({g237, g661, g1224, g1200}, g1423);
	defparam lut_18124.LUT_SIZE = 4;
	defparam lut_18124.mask = 16'h8000;

	lut_sub lut_18132 ({g43, g495, g1122, g1296}, g1424);
	defparam lut_18132.LUT_SIZE = 4;
	defparam lut_18132.mask = 16'ha2a0;

	lut_sub lut_18143 ({i_14_, i_12_, i_13_, g112, g131, g158}, g1425);
	defparam lut_18143.LUT_SIZE = 6;
	defparam lut_18143.mask = 64'h0507070707070503;

	lut_sub lut_18172 ({g8, g10, g112, g1174, g1425}, g1426);
	defparam lut_18172.LUT_SIZE = 5;
	defparam lut_18172.mask = 32'h80808880;

	lut_sub lut_18185 ({g381, g1275, g1423, g1424, g1426}, g1427);
	defparam lut_18185.LUT_SIZE = 5;
	defparam lut_18185.mask = 32'h00010000;

	lut_sub lut_18192 ({g1151, g1358, g1398}, g1428);
	defparam lut_18192.LUT_SIZE = 3;
	defparam lut_18192.mask = 8'h01;

	lut_sub lut_18202 ({g1219, g1415, g1421, g1422, g1427, g1428}, g1429);
	defparam lut_18202.LUT_SIZE = 6;
	defparam lut_18202.mask = 64'h0000000000000100;

	lut_sub lut_18211 ({g560, g561, g549, g540, g895}, g1430);
	defparam lut_18211.LUT_SIZE = 5;
	defparam lut_18211.mask = 32'h08000000;

	lut_sub lut_18219 ({g134, g824, g1300, g1430}, g1431);
	defparam lut_18219.LUT_SIZE = 4;
	defparam lut_18219.mask = 16'h3301;

	lut_sub lut_18233 ({g8, g10, g23, g136, g132, g462}, g1432);
	defparam lut_18233.LUT_SIZE = 6;
	defparam lut_18233.mask = 64'h0f0f0f0f0e0f0f0f;

	lut_sub lut_18270 ({i_14_, i_12_, i_13_, g136, g131, g158}, g1433);
	defparam lut_18270.LUT_SIZE = 6;
	defparam lut_18270.mask = 64'h0500050503000503;

	lut_sub lut_18291 ({g135, g1112, g1263, g1419, g1432, g1433}, g1434);
	defparam lut_18291.LUT_SIZE = 6;
	defparam lut_18291.mask = 64'h0088008800000080;

	lut_sub lut_18304 ({g1202, g1229, g1352, g1434, g1640}, g1435);
	defparam lut_18304.LUT_SIZE = 5;
	defparam lut_18304.mask = 32'h00000001;

	lut_sub lut_18314 ({g73, g1329, g1568, g1429, g1431, g1435}, o_20_);
	defparam lut_18314.LUT_SIZE = 6;
	defparam lut_18314.mask = 64'h00000000fffffffe;

	lut_sub lut_18350 ({g73, g1429}, g1437);
	defparam lut_18350.LUT_SIZE = 2;
	defparam lut_18350.mask = 4'b1101;

	lut_sub lut_18356 ({i_11_, i_9_, i_10_, i_8_}, g1438);
	defparam lut_18356.LUT_SIZE = 4;
	defparam lut_18356.mask = 16'h5a52;

	lut_sub lut_18370 ({i_15_, g4, g87, g182, g1438}, g1439);
	defparam lut_18370.LUT_SIZE = 5;
	defparam lut_18370.mask = 32'h00000001;

	lut_sub lut_18378 ({g227, g349, g1007, g1439}, o_22_);
	defparam lut_18378.LUT_SIZE = 4;
	defparam lut_18378.mask = 16'h777f;

	lut_sub lut_18395 ({i_5_, i_3_, i_4_, g1}, g1441);
	defparam lut_18395.LUT_SIZE = 4;
	defparam lut_18395.mask = 16'h0001;

	lut_sub lut_18401 ({g30, g1441}, g1442);
	defparam lut_18401.LUT_SIZE = 2;
	defparam lut_18401.mask = 4'b0001;

	lut_sub lut_18411 ({g1155, g1230, g1231, g1234, g1307, g1309}, g1443);
	defparam lut_18411.LUT_SIZE = 6;
	defparam lut_18411.mask = 64'h0100000000000000;

	lut_sub lut_18420 ({g132, g159, g566, g531, g522}, g1444);
	defparam lut_18420.LUT_SIZE = 5;
	defparam lut_18420.mask = 32'h00008000;

	lut_sub lut_18429 ({i_8_, g66, g108, g207, g1085, g1444}, g1445);
	defparam lut_18429.LUT_SIZE = 6;
	defparam lut_18429.mask = 64'h00ee00ee000e00ff;

	lut_sub lut_18457 ({i_14_, i_12_, i_13_, g131, g158}, g1446);
	defparam lut_18457.LUT_SIZE = 5;
	defparam lut_18457.mask = 32'h35030035;

	lut_sub lut_18475 ({g46, g101, g108, g209, g1446}, g1447);
	defparam lut_18475.LUT_SIZE = 5;
	defparam lut_18475.mask = 32'hfac8fa00;

	lut_sub lut_18498 ({g109, g529, g801, g819, g1260}, g1448);
	defparam lut_18498.LUT_SIZE = 5;
	defparam lut_18498.mask = 32'hcccc0004;

	lut_sub lut_18513 ({i_8_, g108, g316, g132}, g1449);
	defparam lut_18513.LUT_SIZE = 4;
	defparam lut_18513.mask = 16'h030a;

	lut_sub lut_18524 ({g8, i_8_, g46, g108, g895}, g1450);
	defparam lut_18524.LUT_SIZE = 5;
	defparam lut_18524.mask = 32'hffccffec;

	lut_sub lut_18557 ({g145, g638, g676, g677, g1157}, g1451);
	defparam lut_18557.LUT_SIZE = 5;
	defparam lut_18557.mask = 32'h0000ffbf;

	lut_sub lut_18581 ({g1445, g1447, g1448, g1449, g1545, g1451}, g1452);
	defparam lut_18581.LUT_SIZE = 6;
	defparam lut_18581.mask = 64'h0000002000000000;

	lut_sub lut_18591 ({g1028, g1206, g1347, g1392, g1443, g1452}, g1453);
	defparam lut_18591.LUT_SIZE = 6;
	defparam lut_18591.mask = 64'h0000000000000001;

	lut_sub lut_18597 ({g613, g555}, g1454);
	defparam lut_18597.LUT_SIZE = 2;
	defparam lut_18597.mask = 4'b0010;

	lut_sub lut_18606 ({i_8_, g108, g268, g172, g895, g1454}, g1455);
	defparam lut_18606.LUT_SIZE = 6;
	defparam lut_18606.mask = 64'h0000bbbb0000afff;

	lut_sub lut_18639 ({i_8_, g100, g270, g554, g678}, g1456);
	defparam lut_18639.LUT_SIZE = 5;
	defparam lut_18639.mask = 32'h000000fb;

	lut_sub lut_18654 ({g47, g108, g598, g937, g1456}, g1457);
	defparam lut_18654.LUT_SIZE = 5;
	defparam lut_18654.mask = 32'h80808000;

	lut_sub lut_18666 ({g744, g834, g1192, g1359, g1455, g1457}, g1458);
	defparam lut_18666.LUT_SIZE = 6;
	defparam lut_18666.mask = 64'h0000400000000000;

	lut_sub lut_18676 ({g1003, g1004, g1278, g1279, g1330, g1458}, g1459);
	defparam lut_18676.LUT_SIZE = 6;
	defparam lut_18676.mask = 64'h0010000000000000;

	lut_sub lut_18685 ({g101, g531, g996, g997, g998}, g1460);
	defparam lut_18685.LUT_SIZE = 5;
	defparam lut_18685.mask = 32'h02020200;

	lut_sub lut_18692 ({i_3_, i_4_, g1, i_8_, i_6_, i_7_}, g1461);
	defparam lut_18692.LUT_SIZE = 6;
	defparam lut_18692.mask = 64'h002000a000000000;

	lut_sub lut_18702 ({g32, g21, g900, g1461}, g1462);
	defparam lut_18702.LUT_SIZE = 4;
	defparam lut_18702.mask = 16'hc8c0;

	lut_sub lut_18715 ({g101, g534, g983, g984, g1462}, g1463);
	defparam lut_18715.LUT_SIZE = 5;
	defparam lut_18715.mask = 32'h01010100;

	lut_sub lut_18723 ({g32, g1461}, g1464);
	defparam lut_18723.LUT_SIZE = 2;
	defparam lut_18723.mask = 4'b1000;

	lut_sub lut_18731 ({g23, g12, g978, g1464}, g1465);
	defparam lut_18731.LUT_SIZE = 4;
	defparam lut_18731.mask = 16'h3111;

	lut_sub lut_18744 ({g976, g994, g1460, g1463, g1465}, g1466);
	defparam lut_18744.LUT_SIZE = 5;
	defparam lut_18744.mask = 32'h00000001;

	lut_sub lut_18754 ({g73, g1018, g1442, g1453, g1459, g1466}, g1467);
	defparam lut_18754.LUT_SIZE = 6;
	defparam lut_18754.mask = 64'hffffffff00000100;

	lut_sub lut_18792 ({g31, g64}, g1468);
	defparam lut_18792.LUT_SIZE = 2;
	defparam lut_18792.mask = 4'b0001;

	lut_sub lut_18801 ({g7, g25, g3, g131, g1468}, g1469);
	defparam lut_18801.LUT_SIZE = 5;
	defparam lut_18801.mask = 32'haaffa8fc;

	lut_sub lut_18830 ({g12, g101, g971, g974, g975}, g1470);
	defparam lut_18830.LUT_SIZE = 5;
	defparam lut_18830.mask = 32'h02020200;

	lut_sub lut_18841 ({g101, g534, g978, g983, g984}, g1471);
	defparam lut_18841.LUT_SIZE = 5;
	defparam lut_18841.mask = 32'h01010100;

	lut_sub lut_18850 ({g987, g990, g992}, g1472);
	defparam lut_18850.LUT_SIZE = 3;
	defparam lut_18850.mask = 8'h10;

	lut_sub lut_18857 ({g99, g119, g711}, g1473);
	defparam lut_18857.LUT_SIZE = 3;
	defparam lut_18857.mask = 8'h01;

	lut_sub lut_18867 ({g101, g299, g745, g898, g1064, g1473}, g1474);
	defparam lut_18867.LUT_SIZE = 6;
	defparam lut_18867.mask = 64'haa00000020000000;

	lut_sub lut_18880 ({g1470, g1471, g1472, g1460, g1474}, g1475);
	defparam lut_18880.LUT_SIZE = 5;
	defparam lut_18880.mask = 32'h00000001;

	lut_sub lut_18889 ({g73, g1018, g1453, g1459, g1475}, g1476);
	defparam lut_18889.LUT_SIZE = 5;
	defparam lut_18889.mask = 32'hffff0001;

	lut_sub lut_18915 ({g338, g540, g1286, g1607, g1353, g1410}, g1477);
	defparam lut_18915.LUT_SIZE = 6;
	defparam lut_18915.mask = 64'h0100000001000100;

	lut_sub lut_18923 ({i_1_, i_0_, i_2_, g4, g73}, o_27_);
	defparam lut_18923.LUT_SIZE = 5;
	defparam lut_18923.mask = 32'h00000010;

	lut_sub lut_18929 ({g2, i_8_, i_6_, i_7_, g42}, g1479);
	defparam lut_18929.LUT_SIZE = 5;
	defparam lut_18929.mask = 32'h05000d00;

	lut_sub lut_18941 ({g32, g75, g1468, g1479}, g1480);
	defparam lut_18941.LUT_SIZE = 4;
	defparam lut_18941.mask = 16'h8000;

	lut_sub lut_18946 ({i_3_, i_4_, i_6_, i_7_, g29}, g1481);
	defparam lut_18946.LUT_SIZE = 5;
	defparam lut_18946.mask = 32'h00040000;

	lut_sub lut_18955 ({g32, g20, g75, g1468, g1481}, g1482);
	defparam lut_18955.LUT_SIZE = 5;
	defparam lut_18955.mask = 32'h80aa00aa;

	lut_sub lut_18969 ({i_3_, i_4_, g30, g29}, g1483);
	defparam lut_18969.LUT_SIZE = 4;
	defparam lut_18969.mask = 16'h0100;

	lut_sub lut_18978 ({g32, g19, g75, g1468, g1483}, g1484);
	defparam lut_18978.LUT_SIZE = 5;
	defparam lut_18978.mask = 32'haa80aa00;

	lut_sub lut_18994 ({g19, g20, g1479, g1484}, g1485);
	defparam lut_18994.LUT_SIZE = 4;
	defparam lut_18994.mask = 16'h4544;

	lut_sub lut_19006 ({g16, g1480, g1482, g1485}, g1486);
	defparam lut_19006.LUT_SIZE = 4;
	defparam lut_19006.mask = 16'h0111;

	lut_sub lut_19013 ({i_3_, i_4_, g29}, g1487);
	defparam lut_19013.LUT_SIZE = 3;
	defparam lut_19013.mask = 8'h40;

	lut_sub lut_19021 ({g5, g61, g62, g111}, g1488);
	defparam lut_19021.LUT_SIZE = 4;
	defparam lut_19021.mask = 16'h0015;

	lut_sub lut_19031 ({i_7_, g141, g1487, g63, g1488}, g1489);
	defparam lut_19031.LUT_SIZE = 5;
	defparam lut_19031.mask = 32'ha080aa88;

	lut_sub lut_19048 ({g19, g20, g16, g78, g1489}, g1490);
	defparam lut_19048.LUT_SIZE = 5;
	defparam lut_19048.mask = 32'h44454444;

	lut_sub lut_19065 ({g30, g61, g73, g1486, g1490}, g1491);
	defparam lut_19065.LUT_SIZE = 5;
	defparam lut_19065.mask = 32'hf1f0f1f1;

	lut_sub lut_19092 ({g14, g4, g29, g39, g1480}, g1492);
	defparam lut_19092.LUT_SIZE = 5;
	defparam lut_19092.mask = 32'h0003aaab;

	lut_sub lut_19111 ({g8, g32, g75, g1468, g1479}, g1493);
	defparam lut_19111.LUT_SIZE = 5;
	defparam lut_19111.mask = 32'h7fff0000;

	lut_sub lut_19132 ({i_3_, i_4_, g34, g29, g1493}, g1494);
	defparam lut_19132.LUT_SIZE = 5;
	defparam lut_19132.mask = 32'haaa8aaaa;

	lut_sub lut_19155 ({g10, g78, g1480, g1492, g1494}, g1495);
	defparam lut_19155.LUT_SIZE = 5;
	defparam lut_19155.mask = 32'h44440400;

	lut_sub lut_19164 ({i_5_, i_3_, i_4_, g29}, g1496);
	defparam lut_19164.LUT_SIZE = 4;
	defparam lut_19164.mask = 16'h4050;

	lut_sub lut_19174 ({g14, g4, g78, g1496}, g1497);
	defparam lut_19174.LUT_SIZE = 4;
	defparam lut_19174.mask = 16'h0537;

	lut_sub lut_19188 ({g8, g34, g1487, g78}, g1498);
	defparam lut_19188.LUT_SIZE = 4;
	defparam lut_19188.mask = 16'h5703;

	lut_sub lut_19203 ({g30, g1441, g1488, g1497, g1498}, g1499);
	defparam lut_19203.LUT_SIZE = 5;
	defparam lut_19203.mask = 32'h80008080;

	lut_sub lut_19213 ({i_9_, i_10_, g63, g73, g1495, g1499}, o_29_);
	defparam lut_19213.LUT_SIZE = 6;
	defparam lut_19213.mask = 64'h0e0e0e0e0e0f0e0e;

	lut_sub lut_19244 ({g2, i_6_, i_7_, g40, g77}, g1501);
	defparam lut_19244.LUT_SIZE = 5;
	defparam lut_19244.mask = 32'h00070f0f;

	lut_sub lut_19260 ({i_3_, i_4_, g29, g1501}, g1502);
	defparam lut_19260.LUT_SIZE = 4;
	defparam lut_19260.mask = 16'h8aaa;

	lut_sub lut_19275 ({g73, g81, g1486, g1495, g1502}, g1503);
	defparam lut_19275.LUT_SIZE = 5;
	defparam lut_19275.mask = 32'hffff0001;

	lut_sub lut_19298 ({i_3_, i_4_, g1, g32, g27}, g1504);
	defparam lut_19298.LUT_SIZE = 5;
	defparam lut_19298.mask = 32'hc8cccccc;

	lut_sub lut_19319 ({i_9_, i_10_, g63, g1488, g1504}, o_31_);
	defparam lut_19319.LUT_SIZE = 5;
	defparam lut_19319.mask = 32'hbb3f3f33;

	lut_sub lut_19345 ({i_5_, i_3_, i_4_, g1, i_6_, i_7_}, g1506);
	defparam lut_19345.LUT_SIZE = 6;
	defparam lut_19345.mask = 64'hfafafffefffffff6;

	lut_sub lut_19410 ({g19, g5, g41, g78, g1479}, g1507);
	defparam lut_19410.LUT_SIZE = 5;
	defparam lut_19410.mask = 32'h000f770f;

	lut_sub lut_19432 ({g30, g23, g1487, g1464, g1498}, g1508);
	defparam lut_19432.LUT_SIZE = 5;
	defparam lut_19432.mask = 32'haa22a020;

	lut_sub lut_19449 ({g73, g1484, g1494, g1507, g1508}, g1509);
	defparam lut_19449.LUT_SIZE = 5;
	defparam lut_19449.mask = 32'hffff0004;

	lut_sub lut_19473 ({g976, g994, g1460, g1463}, g1510);
	defparam lut_19473.LUT_SIZE = 4;
	defparam lut_19473.mask = 16'h0001;

	lut_sub lut_19480 ({g931, g1266, g1268}, g1511);
	defparam lut_19480.LUT_SIZE = 3;
	defparam lut_19480.mask = 8'h40;

	lut_sub lut_19489 ({g1278, g1279, g1281, g1282, g1492}, g1512);
	defparam lut_19489.LUT_SIZE = 5;
	defparam lut_19489.mask = 32'h00000800;

	lut_sub lut_19494 ({i_11_, i_9_, i_10_, i_15_, g13}, g1513);
	defparam lut_19494.LUT_SIZE = 5;
	defparam lut_19494.mask = 32'h01001000;

	lut_sub lut_19505 ({g101, g109, g641, g676, g903, g1513}, g1514);
	defparam lut_19505.LUT_SIZE = 6;
	defparam lut_19505.mask = 64'hffffaa00c0c08000;

	lut_sub lut_19535 ({i_14_, i_12_, i_8_, g102, g108}, g1515);
	defparam lut_19535.LUT_SIZE = 5;
	defparam lut_19535.mask = 32'h00000400;

	lut_sub lut_19544 ({g20, g78, g1479, g1482, g1515}, g1516);
	defparam lut_19544.LUT_SIZE = 5;
	defparam lut_19544.mask = 32'h20002222;

	lut_sub lut_19555 ({i_3_, i_4_, g1, g5, g27}, g1517);
	defparam lut_19555.LUT_SIZE = 5;
	defparam lut_19555.mask = 32'h00010000;

	lut_sub lut_19561 ({i_6_, i_7_, g1487, g1517}, g1518);
	defparam lut_19561.LUT_SIZE = 4;
	defparam lut_19561.mask = 16'haa8a;

	lut_sub lut_19576 ({i_8_, g10, g100, g108, g640, g677}, g1519);
	defparam lut_19576.LUT_SIZE = 6;
	defparam lut_19576.mask = 64'h000000000c5d0cff;

	lut_sub lut_19601 ({g101, g848, g1497, g1518, g1519}, g1520);
	defparam lut_19601.LUT_SIZE = 5;
	defparam lut_19601.mask = 32'h20200020;

	lut_sub lut_19612 ({g1589, g1380, g1514, g1516, g1520}, g1521);
	defparam lut_19612.LUT_SIZE = 5;
	defparam lut_19612.mask = 32'h00000100;

	lut_sub lut_19621 ({g1511, g1321, g1402, g1512, g1521}, g1522);
	defparam lut_19621.LUT_SIZE = 5;
	defparam lut_19621.mask = 32'h00000001;

	lut_sub lut_19630 ({g73, g1195, g1453, g1510, g1522}, o_34_);
	defparam lut_19630.LUT_SIZE = 5;
	defparam lut_19630.mask = 32'h0000fffe;

	lut_sub lut_19653 ({g10, g16, g5, g78, g1480}, g1524);
	defparam lut_19653.LUT_SIZE = 5;
	defparam lut_19653.mask = 32'h44fc4444;

	lut_sub lut_19672 ({g12, g73, g1464, g1524}, o_35_);
	defparam lut_19672.LUT_SIZE = 4;
	defparam lut_19672.mask = 16'h0a0e;

	lut_sub lut_19683 ({i_8_, g30, g5, g61}, g1526);
	defparam lut_19683.LUT_SIZE = 4;
	defparam lut_19683.mask = 16'h0501;

	lut_sub lut_19694 ({g38, g64, g101, g531, g1526}, g1527);
	defparam lut_19694.LUT_SIZE = 5;
	defparam lut_19694.mask = 32'ha8a8a800;

	lut_sub lut_19711 ({g31, g25, g27, g64, g1527}, g1528);
	defparam lut_19711.LUT_SIZE = 5;
	defparam lut_19711.mask = 32'h54554455;

	lut_sub lut_19733 ({g83, g976, g985, g994, g999, g1528}, g1529);
	defparam lut_19733.LUT_SIZE = 6;
	defparam lut_19733.mask = 64'h0000000000000001;

	lut_sub lut_19743 ({g73, g1018, g1442, g1453, g1459, g1529}, g1530);
	defparam lut_19743.LUT_SIZE = 6;
	defparam lut_19743.mask = 64'hffffffff00000100;

	lut_sub lut_19782 ({g26, g27, g38}, g1531);
	defparam lut_19782.LUT_SIZE = 3;
	defparam lut_19782.mask = 8'h8a;

	lut_sub lut_19791 ({i_8_, g30, g5, g62}, g1532);
	defparam lut_19791.LUT_SIZE = 4;
	defparam lut_19791.mask = 16'h0501;

	lut_sub lut_19802 ({g37, g65, g73, g1531, g1532}, o_37_);
	defparam lut_19802.LUT_SIZE = 5;
	defparam lut_19802.mask = 32'h0f0f050d;

	lut_sub lut_19820 ({i_3_, i_4_, g1, g34}, o_38_);
	defparam lut_19820.LUT_SIZE = 4;
	defparam lut_19820.mask = 16'h0001;

	lut_sub lut_19825 ({i_3_, i_4_, g1, i_6_, i_7_}, o_39_);
	defparam lut_19825.LUT_SIZE = 5;
	defparam lut_19825.mask = 32'h00000002;

	lut_sub lut_19832 ({g95, i_13_, i_12_, i_14_, g93, g108}, g1536);
	defparam lut_19832.LUT_SIZE = 6;
	defparam lut_19832.mask = 64'h4000000045500050;

	lut_sub lut_19846 ({g95, i_13_, i_12_, i_14_, g93, g108}, g1537);
	defparam lut_19846.LUT_SIZE = 6;
	defparam lut_19846.mask = 64'h4044404045554050;

	lut_sub lut_19866 ({g1536, g1537, i_8_}, g1538);
	defparam lut_19866.LUT_SIZE = 3;
	defparam lut_19866.mask = 8'he4;

	lut_sub lut_19876 ({g22, i_13_, i_12_, i_14_, g11, g88}, g1539);
	defparam lut_19876.LUT_SIZE = 6;
	defparam lut_19876.mask = 64'h0011101050555055;

	lut_sub lut_19898 ({g22, i_13_, i_12_, i_14_, g11, g88}, g1540);
	defparam lut_19898.LUT_SIZE = 6;
	defparam lut_19898.mask = 64'h0010100000151005;

	lut_sub lut_19911 ({g1539, g1540, i_8_}, g1541);
	defparam lut_19911.LUT_SIZE = 3;
	defparam lut_19911.mask = 8'he4;

	lut_sub lut_19922 ({g158, g131, g1027, g99}, g1542);
	defparam lut_19922.LUT_SIZE = 4;
	defparam lut_19922.mask = 16'hc888;

	lut_sub lut_19936 ({g183, g88, g196, g194, g192, g190}, g1543);
	defparam lut_19936.LUT_SIZE = 6;
	defparam lut_19936.mask = 64'h8000800080000000;

	lut_sub lut_19948 ({g10, g20, g19, g77, g75, g8}, g1544);
	defparam lut_19948.LUT_SIZE = 6;
	defparam lut_19948.mask = 64'hc0c0d0c0c0c0c0c0;

	lut_sub lut_19970 ({g1546, g1547}, g1545);
	defparam lut_19970.LUT_SIZE = 2;
	defparam lut_19970.mask = 4'b1000;

	lut_sub lut_19976 ({g544, g1548}, g1546);
	defparam lut_19976.LUT_SIZE = 2;
	defparam lut_19976.mask = 4'b0100;

	lut_sub lut_19982 ({g544, g1551}, g1547);
	defparam lut_19982.LUT_SIZE = 2;
	defparam lut_19982.mask = 4'b0001;

	lut_sub lut_19988 ({g1549, g1550}, g1548);
	defparam lut_19988.LUT_SIZE = 2;
	defparam lut_19988.mask = 4'b1000;

	lut_sub lut_19993 ({i_8_, g1554}, g1549);
	defparam lut_19993.LUT_SIZE = 2;
	defparam lut_19993.mask = 4'b0100;

	lut_sub lut_19998 ({i_8_, g1555}, g1550);
	defparam lut_19998.LUT_SIZE = 2;
	defparam lut_19998.mask = 4'b0001;

	lut_sub lut_20004 ({g1552, g1553}, g1551);
	defparam lut_20004.LUT_SIZE = 2;
	defparam lut_20004.mask = 4'b1000;

	lut_sub lut_20009 ({i_8_, g1556}, g1552);
	defparam lut_20009.LUT_SIZE = 2;
	defparam lut_20009.mask = 4'b0100;

	lut_sub lut_20014 ({i_8_, g1557}, g1553);
	defparam lut_20014.LUT_SIZE = 2;
	defparam lut_20014.mask = 4'b0001;

	lut_sub lut_20021 ({g108, g1450, g470}, g1554);
	defparam lut_20021.LUT_SIZE = 3;
	defparam lut_20021.mask = 8'h32;

	lut_sub lut_20029 ({g108, g1450}, g1555);
	defparam lut_20029.LUT_SIZE = 2;
	defparam lut_20029.mask = 4'b0100;

	lut_sub lut_20036 ({g108, g1450, g470}, g1556);
	defparam lut_20036.LUT_SIZE = 3;
	defparam lut_20036.mask = 8'h32;

	lut_sub lut_20046 ({g108, g1450, g204, g848}, g1557);
	defparam lut_20046.LUT_SIZE = 4;
	defparam lut_20046.mask = 16'h0f01;

	lut_sub lut_20056 ({g1559, g1560}, g1558);
	defparam lut_20056.LUT_SIZE = 2;
	defparam lut_20056.mask = 4'b1000;

	lut_sub lut_20062 ({g134, g1561}, g1559);
	defparam lut_20062.LUT_SIZE = 2;
	defparam lut_20062.mask = 4'b0100;

	lut_sub lut_20068 ({g134, g1564}, g1560);
	defparam lut_20068.LUT_SIZE = 2;
	defparam lut_20068.mask = 4'b0001;

	lut_sub lut_20074 ({g1562, g1563}, g1561);
	defparam lut_20074.LUT_SIZE = 2;
	defparam lut_20074.mask = 4'b1000;

	lut_sub lut_20080 ({g678, g1566}, g1562);
	defparam lut_20080.LUT_SIZE = 2;
	defparam lut_20080.mask = 4'b0100;

	lut_sub lut_20086 ({g678, g1411}, g1563);
	defparam lut_20086.LUT_SIZE = 2;
	defparam lut_20086.mask = 4'b0001;

	lut_sub lut_20092 ({g678, g1565}, g1564);
	defparam lut_20092.LUT_SIZE = 2;
	defparam lut_20092.mask = 4'b0010;

	lut_sub lut_20098 ({g678, g1567}, g1565);
	defparam lut_20098.LUT_SIZE = 2;
	defparam lut_20098.mask = 4'b0001;

	lut_sub lut_20104 ({g118, g1411}, g1566);
	defparam lut_20104.LUT_SIZE = 2;
	defparam lut_20104.mask = 4'b0111;

	lut_sub lut_20114 ({g572, g93, g270, g1411}, g1567);
	defparam lut_20114.LUT_SIZE = 4;
	defparam lut_20114.mask = 16'hddfd;

	lut_sub lut_20132 ({g1569, g1570}, g1568);
	defparam lut_20132.LUT_SIZE = 2;
	defparam lut_20132.mask = 4'b1000;

	lut_sub lut_20138 ({g96, g1571}, g1569);
	defparam lut_20138.LUT_SIZE = 2;
	defparam lut_20138.mask = 4'b0100;

	lut_sub lut_20144 ({g96, g1574}, g1570);
	defparam lut_20144.LUT_SIZE = 2;
	defparam lut_20144.mask = 4'b0001;

	lut_sub lut_20150 ({g1572, g1573}, g1571);
	defparam lut_20150.LUT_SIZE = 2;
	defparam lut_20150.mask = 4'b1000;

	lut_sub lut_20156 ({g1384, g1577}, g1572);
	defparam lut_20156.LUT_SIZE = 2;
	defparam lut_20156.mask = 4'b0100;

	lut_sub lut_20162 ({g1384, g1578}, g1573);
	defparam lut_20162.LUT_SIZE = 2;
	defparam lut_20162.mask = 4'b0001;

	lut_sub lut_20168 ({g1575, g1576}, g1574);
	defparam lut_20168.LUT_SIZE = 2;
	defparam lut_20168.mask = 4'b1000;

	lut_sub lut_20174 ({g1384, g1579}, g1575);
	defparam lut_20174.LUT_SIZE = 2;
	defparam lut_20174.mask = 4'b0100;

	lut_sub lut_20180 ({g1384, g1387}, g1576);
	defparam lut_20180.LUT_SIZE = 2;
	defparam lut_20180.mask = 4'b0001;

	lut_sub lut_20186 ({g135, g1387}, g1577);
	defparam lut_20186.LUT_SIZE = 2;
	defparam lut_20186.mask = 4'b0100;

	lut_sub lut_20193 ({g135, g1387, g134}, g1578);
	defparam lut_20193.LUT_SIZE = 3;
	defparam lut_20193.mask = 8'h32;

	lut_sub lut_20202 ({g135, g1387, i_8_, g669}, g1579);
	defparam lut_20202.LUT_SIZE = 4;
	defparam lut_20202.mask = 16'h0f04;

	lut_sub lut_20212 ({g1581, g1582}, g1580);
	defparam lut_20212.LUT_SIZE = 2;
	defparam lut_20212.mask = 4'b1000;

	lut_sub lut_20217 ({i_14_, g1583}, g1581);
	defparam lut_20217.LUT_SIZE = 2;
	defparam lut_20217.mask = 4'b0100;

	lut_sub lut_20222 ({i_14_, g1585}, g1582);
	defparam lut_20222.LUT_SIZE = 2;
	defparam lut_20222.mask = 4'b0001;

	lut_sub lut_20227 ({i_13_, g1584}, g1583);
	defparam lut_20227.LUT_SIZE = 2;
	defparam lut_20227.mask = 4'b0010;

	lut_sub lut_20232 ({i_13_, g1587}, g1584);
	defparam lut_20232.LUT_SIZE = 2;
	defparam lut_20232.mask = 4'b0001;

	lut_sub lut_20237 ({i_13_, g1586}, g1585);
	defparam lut_20237.LUT_SIZE = 2;
	defparam lut_20237.mask = 4'b1000;

	lut_sub lut_20242 ({i_13_, g1588}, g1586);
	defparam lut_20242.LUT_SIZE = 2;
	defparam lut_20242.mask = 4'b0100;

	lut_sub lut_20248 ({g18, i_12_, g135}, g1587);
	defparam lut_20248.LUT_SIZE = 3;
	defparam lut_20248.mask = 8'hef;

	lut_sub lut_20261 ({g18, i_12_, g212, g215}, g1588);
	defparam lut_20261.LUT_SIZE = 4;
	defparam lut_20261.mask = 16'h1fff;

	lut_sub lut_20279 ({g108, g1590}, g1589);
	defparam lut_20279.LUT_SIZE = 2;
	defparam lut_20279.mask = 4'b0010;

	lut_sub lut_20285 ({g108, g1591}, g1590);
	defparam lut_20285.LUT_SIZE = 2;
	defparam lut_20285.mask = 4'b0001;

	lut_sub lut_20291 ({g1592, g1593}, g1591);
	defparam lut_20291.LUT_SIZE = 2;
	defparam lut_20291.mask = 4'b1000;

	lut_sub lut_20296 ({i_14_, g1594}, g1592);
	defparam lut_20296.LUT_SIZE = 2;
	defparam lut_20296.mask = 4'b0100;

	lut_sub lut_20301 ({i_14_, g1595}, g1593);
	defparam lut_20301.LUT_SIZE = 2;
	defparam lut_20301.mask = 4'b0001;

	lut_sub lut_20307 ({i_13_, i_12_, g102, g115}, g1594);
	defparam lut_20307.LUT_SIZE = 4;
	defparam lut_20307.mask = 16'h5131;

	lut_sub lut_20317 ({i_13_, i_12_, i_8_, g115}, g1595);
	defparam lut_20317.LUT_SIZE = 4;
	defparam lut_20317.mask = 16'hfdff;

	lut_sub lut_20337 ({g1597, g1598}, g1596);
	defparam lut_20337.LUT_SIZE = 2;
	defparam lut_20337.mask = 4'b1000;

	lut_sub lut_20343 ({g119, g1599}, g1597);
	defparam lut_20343.LUT_SIZE = 2;
	defparam lut_20343.mask = 4'b0100;

	lut_sub lut_20349 ({g119, g1601}, g1598);
	defparam lut_20349.LUT_SIZE = 2;
	defparam lut_20349.mask = 4'b0001;

	lut_sub lut_20355 ({g134, g1600}, g1599);
	defparam lut_20355.LUT_SIZE = 2;
	defparam lut_20355.mask = 4'b0010;

	lut_sub lut_20361 ({g134, g1604}, g1600);
	defparam lut_20361.LUT_SIZE = 2;
	defparam lut_20361.mask = 4'b0001;

	lut_sub lut_20367 ({g1602, g1603}, g1601);
	defparam lut_20367.LUT_SIZE = 2;
	defparam lut_20367.mask = 4'b1000;

	lut_sub lut_20373 ({g134, g1605}, g1602);
	defparam lut_20373.LUT_SIZE = 2;
	defparam lut_20373.mask = 4'b0100;

	lut_sub lut_20379 ({g134, g1606}, g1603);
	defparam lut_20379.LUT_SIZE = 2;
	defparam lut_20379.mask = 4'b0001;

	lut_sub lut_20384 ({i_13_, i_12_, g122, i_14_}, g1604);
	defparam lut_20384.LUT_SIZE = 4;
	defparam lut_20384.mask = 16'h7b3f;

	lut_sub lut_20400 ({i_13_, i_12_, g136, i_14_}, g1605);
	defparam lut_20400.LUT_SIZE = 4;
	defparam lut_20400.mask = 16'hfeff;

	lut_sub lut_20419 ({i_13_, i_12_, g122, i_14_}, g1606);
	defparam lut_20419.LUT_SIZE = 4;
	defparam lut_20419.mask = 16'h701f;

	lut_sub lut_20432 ({g1608, g1609}, g1607);
	defparam lut_20432.LUT_SIZE = 2;
	defparam lut_20432.mask = 4'b1000;

	lut_sub lut_20438 ({g149, g1610}, g1608);
	defparam lut_20438.LUT_SIZE = 2;
	defparam lut_20438.mask = 4'b0100;

	lut_sub lut_20444 ({g149, g1613}, g1609);
	defparam lut_20444.LUT_SIZE = 2;
	defparam lut_20444.mask = 4'b0001;

	lut_sub lut_20450 ({g1611, g1612}, g1610);
	defparam lut_20450.LUT_SIZE = 2;
	defparam lut_20450.mask = 4'b1000;

	lut_sub lut_20456 ({g201, g1614}, g1611);
	defparam lut_20456.LUT_SIZE = 2;
	defparam lut_20456.mask = 4'b0100;

	lut_sub lut_20462 ({g201, g452}, g1612);
	defparam lut_20462.LUT_SIZE = 2;
	defparam lut_20462.mask = 4'b0001;

	lut_sub lut_20468 ({g201, g1615}, g1613);
	defparam lut_20468.LUT_SIZE = 2;
	defparam lut_20468.mask = 4'b0001;

	lut_sub lut_20474 ({g452, g338}, g1614);
	defparam lut_20474.LUT_SIZE = 2;
	defparam lut_20474.mask = 4'b0001;

	lut_sub lut_20482 ({g1096, g452, g206, g127}, g1615);
	defparam lut_20482.LUT_SIZE = 4;
	defparam lut_20482.mask = 16'h0001;

	lut_sub lut_20488 ({g1116, g1617}, g1616);
	defparam lut_20488.LUT_SIZE = 2;
	defparam lut_20488.mask = 4'b0001;

	lut_sub lut_20494 ({g1618, g1619}, g1617);
	defparam lut_20494.LUT_SIZE = 2;
	defparam lut_20494.mask = 4'b1000;

	lut_sub lut_20499 ({i_8_, g1620}, g1618);
	defparam lut_20499.LUT_SIZE = 2;
	defparam lut_20499.mask = 4'b0100;

	lut_sub lut_20504 ({i_8_, g1621}, g1619);
	defparam lut_20504.LUT_SIZE = 2;
	defparam lut_20504.mask = 4'b0001;

	lut_sub lut_20511 ({g88, g1117, g1118}, g1620);
	defparam lut_20511.LUT_SIZE = 3;
	defparam lut_20511.mask = 8'h54;

	lut_sub lut_20521 ({g696, g88, g185, g1118}, g1621);
	defparam lut_20521.LUT_SIZE = 4;
	defparam lut_20521.mask = 16'h5051;

	lut_sub lut_20531 ({g1102, g1623}, g1622);
	defparam lut_20531.LUT_SIZE = 2;
	defparam lut_20531.mask = 4'b0001;

	lut_sub lut_20537 ({g1624, g1625}, g1623);
	defparam lut_20537.LUT_SIZE = 2;
	defparam lut_20537.mask = 4'b1000;

	lut_sub lut_20542 ({i_8_, g1626}, g1624);
	defparam lut_20542.LUT_SIZE = 2;
	defparam lut_20542.mask = 4'b0100;

	lut_sub lut_20547 ({i_8_, g1627}, g1625);
	defparam lut_20547.LUT_SIZE = 2;
	defparam lut_20547.mask = 4'b0001;

	lut_sub lut_20553 ({g8, g88}, g1626);
	defparam lut_20553.LUT_SIZE = 2;
	defparam lut_20553.mask = 4'b1011;

	lut_sub lut_20563 ({g92, g221, g231, g88}, g1627);
	defparam lut_20563.LUT_SIZE = 4;
	defparam lut_20563.mask = 16'haaab;

	lut_sub lut_20577 ({g1629, g1630}, g1628);
	defparam lut_20577.LUT_SIZE = 2;
	defparam lut_20577.mask = 4'b1000;

	lut_sub lut_20583 ({g90, g1631}, g1629);
	defparam lut_20583.LUT_SIZE = 2;
	defparam lut_20583.mask = 4'b0100;

	lut_sub lut_20589 ({g90, g1634}, g1630);
	defparam lut_20589.LUT_SIZE = 2;
	defparam lut_20589.mask = 4'b0001;

	lut_sub lut_20595 ({g1632, g1633}, g1631);
	defparam lut_20595.LUT_SIZE = 2;
	defparam lut_20595.mask = 4'b1000;

	lut_sub lut_20600 ({i_8_, g88}, g1632);
	defparam lut_20600.LUT_SIZE = 2;
	defparam lut_20600.mask = 4'b1000;

	lut_sub lut_20605 ({i_8_, g1637}, g1633);
	defparam lut_20605.LUT_SIZE = 2;
	defparam lut_20605.mask = 4'b0001;

	lut_sub lut_20611 ({g1635, g1636}, g1634);
	defparam lut_20611.LUT_SIZE = 2;
	defparam lut_20611.mask = 4'b1000;

	lut_sub lut_20616 ({i_8_, g1638}, g1635);
	defparam lut_20616.LUT_SIZE = 2;
	defparam lut_20616.mask = 4'b0100;

	lut_sub lut_20621 ({i_8_, g1639}, g1636);
	defparam lut_20621.LUT_SIZE = 2;
	defparam lut_20621.mask = 4'b0001;

	lut_sub lut_20628 ({g467, g528, g88}, g1637);
	defparam lut_20628.LUT_SIZE = 3;
	defparam lut_20628.mask = 8'hab;

	lut_sub lut_20640 ({g468, g467, g92, g88}, g1638);
	defparam lut_20640.LUT_SIZE = 4;
	defparam lut_20640.mask = 16'haaab;

	lut_sub lut_20655 ({g467, g528, g88}, g1639);
	defparam lut_20655.LUT_SIZE = 3;
	defparam lut_20655.mask = 8'hab;

	lut_sub lut_20665 ({g1641, g1642}, g1640);
	defparam lut_20665.LUT_SIZE = 2;
	defparam lut_20665.mask = 4'b1000;

	lut_sub lut_20671 ({g1031, g1643}, g1641);
	defparam lut_20671.LUT_SIZE = 2;
	defparam lut_20671.mask = 4'b0100;

	lut_sub lut_20677 ({g1031, g1646}, g1642);
	defparam lut_20677.LUT_SIZE = 2;
	defparam lut_20677.mask = 4'b0001;

	lut_sub lut_20683 ({g1644, g1645}, g1643);
	defparam lut_20683.LUT_SIZE = 2;
	defparam lut_20683.mask = 4'b1000;

	lut_sub lut_20688 ({i_8_, g1649}, g1644);
	defparam lut_20688.LUT_SIZE = 2;
	defparam lut_20688.mask = 4'b0100;

	lut_sub lut_20693 ({i_8_, g1650}, g1645);
	defparam lut_20693.LUT_SIZE = 2;
	defparam lut_20693.mask = 4'b0001;

	lut_sub lut_20699 ({g1647, g1648}, g1646);
	defparam lut_20699.LUT_SIZE = 2;
	defparam lut_20699.mask = 4'b1000;

	lut_sub lut_20704 ({i_8_, g1651}, g1647);
	defparam lut_20704.LUT_SIZE = 2;
	defparam lut_20704.mask = 4'b0100;

	lut_sub lut_20709 ({i_8_, g1652}, g1648);
	defparam lut_20709.LUT_SIZE = 2;
	defparam lut_20709.mask = 4'b0001;

	lut_sub lut_20715 ({g400, i_7_, g1038}, g1649);
	defparam lut_20715.LUT_SIZE = 3;
	defparam lut_20715.mask = 8'h54;

	lut_sub lut_20724 ({g400, i_7_, g1032, g1038}, g1650);
	defparam lut_20724.LUT_SIZE = 4;
	defparam lut_20724.mask = 16'h5551;

	lut_sub lut_20737 ({g400, i_7_, g20, g1038}, g1651);
	defparam lut_20737.LUT_SIZE = 4;
	defparam lut_20737.mask = 16'h5551;

	lut_sub lut_20750 ({g400, i_7_, g1032, g1038}, g1652);
	defparam lut_20750.LUT_SIZE = 4;
	defparam lut_20750.mask = 16'h5551;

	lut_sub lut_20762 ({g1654, g1655}, g1653);
	defparam lut_20762.LUT_SIZE = 2;
	defparam lut_20762.mask = 4'b1000;

	lut_sub lut_20768 ({g118, g1656}, g1654);
	defparam lut_20768.LUT_SIZE = 2;
	defparam lut_20768.mask = 4'b0100;

	lut_sub lut_20774 ({g118, g1659}, g1655);
	defparam lut_20774.LUT_SIZE = 2;
	defparam lut_20774.mask = 4'b0001;

	lut_sub lut_20780 ({g1657, g1658}, g1656);
	defparam lut_20780.LUT_SIZE = 2;
	defparam lut_20780.mask = 4'b1000;

	lut_sub lut_20785 ({i_13_, g1662}, g1657);
	defparam lut_20785.LUT_SIZE = 2;
	defparam lut_20785.mask = 4'b0100;

	lut_sub lut_20790 ({i_13_, g1663}, g1658);
	defparam lut_20790.LUT_SIZE = 2;
	defparam lut_20790.mask = 4'b0001;

	lut_sub lut_20796 ({g1660, g1661}, g1659);
	defparam lut_20796.LUT_SIZE = 2;
	defparam lut_20796.mask = 4'b1000;

	lut_sub lut_20801 ({i_13_, g1664}, g1660);
	defparam lut_20801.LUT_SIZE = 2;
	defparam lut_20801.mask = 4'b0100;

	lut_sub lut_20806 ({i_13_, g1665}, g1661);
	defparam lut_20806.LUT_SIZE = 2;
	defparam lut_20806.mask = 4'b0001;

	lut_sub lut_20812 ({i_12_, i_14_, g134, g102}, g1662);
	defparam lut_20812.LUT_SIZE = 4;
	defparam lut_20812.mask = 16'hfdff;

	lut_sub lut_20832 ({i_12_, i_14_, g186, g102}, g1663);
	defparam lut_20832.LUT_SIZE = 4;
	defparam lut_20832.mask = 16'hdfff;

	lut_sub lut_20851 ({i_12_, i_14_, g102}, g1664);
	defparam lut_20851.LUT_SIZE = 3;
	defparam lut_20851.mask = 8'hdf;

	lut_sub lut_20862 ({i_12_, i_14_, g102}, g1665);
	defparam lut_20862.LUT_SIZE = 3;
	defparam lut_20862.mask = 8'h7f;

	lut_sub lut_20873 ({i_14_, g1667}, g1666);
	defparam lut_20873.LUT_SIZE = 2;
	defparam lut_20873.mask = 4'b0010;

	lut_sub lut_20878 ({i_14_, g1668}, g1667);
	defparam lut_20878.LUT_SIZE = 2;
	defparam lut_20878.mask = 4'b0001;

	lut_sub lut_20884 ({g1669, g1670}, g1668);
	defparam lut_20884.LUT_SIZE = 2;
	defparam lut_20884.mask = 4'b1000;

	lut_sub lut_20889 ({i_13_, g1671}, g1669);
	defparam lut_20889.LUT_SIZE = 2;
	defparam lut_20889.mask = 4'b0100;

	lut_sub lut_20894 ({i_13_, g1672}, g1670);
	defparam lut_20894.LUT_SIZE = 2;
	defparam lut_20894.mask = 4'b0001;

	lut_sub lut_20901 ({g495, i_12_, g186, g15}, g1671);
	defparam lut_20901.LUT_SIZE = 4;
	defparam lut_20901.mask = 16'hfdf5;

	lut_sub lut_20919 ({i_12_, g135, g15}, g1672);
	defparam lut_20919.LUT_SIZE = 3;
	defparam lut_20919.mask = 8'hfd;

	lut_sub lut_20931 ({g1674, g1675}, g1673);
	defparam lut_20931.LUT_SIZE = 2;
	defparam lut_20931.mask = 4'b1000;

	lut_sub lut_20937 ({g807, g1676}, g1674);
	defparam lut_20937.LUT_SIZE = 2;
	defparam lut_20937.mask = 4'b0100;

	lut_sub lut_20943 ({g807, g1679}, g1675);
	defparam lut_20943.LUT_SIZE = 2;
	defparam lut_20943.mask = 4'b0001;

	lut_sub lut_20949 ({g1677, g1678}, g1676);
	defparam lut_20949.LUT_SIZE = 2;
	defparam lut_20949.mask = 4'b1000;

	lut_sub lut_20954 ({i_8_, g1682}, g1677);
	defparam lut_20954.LUT_SIZE = 2;
	defparam lut_20954.mask = 4'b0100;

	lut_sub lut_20959 ({i_8_, g1683}, g1678);
	defparam lut_20959.LUT_SIZE = 2;
	defparam lut_20959.mask = 4'b0001;

	lut_sub lut_20965 ({g1680, g1681}, g1679);
	defparam lut_20965.LUT_SIZE = 2;
	defparam lut_20965.mask = 4'b1000;

	lut_sub lut_20970 ({i_8_, g1684}, g1680);
	defparam lut_20970.LUT_SIZE = 2;
	defparam lut_20970.mask = 4'b0100;

	lut_sub lut_20975 ({i_8_, g1685}, g1681);
	defparam lut_20975.LUT_SIZE = 2;
	defparam lut_20975.mask = 4'b0001;

	lut_sub lut_20981 ({g30, g87}, g1682);
	defparam lut_20981.LUT_SIZE = 2;
	defparam lut_20981.mask = 4'b1110;

	lut_sub lut_20990 ({g30, g16, g87}, g1683);
	defparam lut_20990.LUT_SIZE = 3;
	defparam lut_20990.mask = 8'hfb;

	lut_sub lut_21004 ({g30, g464, g226, g87}, g1684);
	defparam lut_21004.LUT_SIZE = 4;
	defparam lut_21004.mask = 16'hffab;

	lut_sub lut_21023 ({g30, g16, g87}, g1685);
	defparam lut_21023.LUT_SIZE = 3;
	defparam lut_21023.mask = 8'hfb;

	lut_sub lut_21035 ({g1687, g1688}, g1686);
	defparam lut_21035.LUT_SIZE = 2;
	defparam lut_21035.mask = 4'b1000;

	lut_sub lut_21040 ({i_6_, g1689}, g1687);
	defparam lut_21040.LUT_SIZE = 2;
	defparam lut_21040.mask = 4'b0100;

	lut_sub lut_21045 ({i_6_, g1691}, g1688);
	defparam lut_21045.LUT_SIZE = 2;
	defparam lut_21045.mask = 4'b0001;

	lut_sub lut_21050 ({i_7_, g1690}, g1689);
	defparam lut_21050.LUT_SIZE = 2;
	defparam lut_21050.mask = 4'b1000;

	lut_sub lut_21055 ({i_7_, g1693}, g1690);
	defparam lut_21055.LUT_SIZE = 2;
	defparam lut_21055.mask = 4'b0100;

	lut_sub lut_21060 ({i_7_, g1692}, g1691);
	defparam lut_21060.LUT_SIZE = 2;
	defparam lut_21060.mask = 4'b0010;

	lut_sub lut_21065 ({i_7_, g1694}, g1692);
	defparam lut_21065.LUT_SIZE = 2;
	defparam lut_21065.mask = 4'b0001;

	lut_sub lut_21072 ({g87, g615, g528}, g1693);
	defparam lut_21072.LUT_SIZE = 3;
	defparam lut_21072.mask = 8'hf1;

	lut_sub lut_21082 ({g98, g616}, g1694);
	defparam lut_21082.LUT_SIZE = 2;
	defparam lut_21082.mask = 4'b1101;

	lut_sub lut_21090 ({g1696, g1697}, g1695);
	defparam lut_21090.LUT_SIZE = 2;
	defparam lut_21090.mask = 4'b1000;

	lut_sub lut_21096 ({g100, g1698}, g1696);
	defparam lut_21096.LUT_SIZE = 2;
	defparam lut_21096.mask = 4'b0100;

	lut_sub lut_21102 ({g100, g1701}, g1697);
	defparam lut_21102.LUT_SIZE = 2;
	defparam lut_21102.mask = 4'b0001;

	lut_sub lut_21108 ({g1699, g1700}, g1698);
	defparam lut_21108.LUT_SIZE = 2;
	defparam lut_21108.mask = 4'b1000;

	lut_sub lut_21113 ({i_8_, g1704}, g1699);
	defparam lut_21113.LUT_SIZE = 2;
	defparam lut_21113.mask = 4'b0100;

	lut_sub lut_21118 ({i_8_, g1705}, g1700);
	defparam lut_21118.LUT_SIZE = 2;
	defparam lut_21118.mask = 4'b0001;

	lut_sub lut_21124 ({g1702, g1703}, g1701);
	defparam lut_21124.LUT_SIZE = 2;
	defparam lut_21124.mask = 4'b1000;

	lut_sub lut_21129 ({i_8_, g1706}, g1702);
	defparam lut_21129.LUT_SIZE = 2;
	defparam lut_21129.mask = 4'b0100;

	lut_sub lut_21134 ({i_8_, g1707}, g1703);
	defparam lut_21134.LUT_SIZE = 2;
	defparam lut_21134.mask = 4'b0001;

	lut_sub lut_21141 ({g592, g590, g251}, g1704);
	defparam lut_21141.LUT_SIZE = 3;
	defparam lut_21141.mask = 8'h45;

	lut_sub lut_21150 ({g592, g590, g251}, g1705);
	defparam lut_21150.LUT_SIZE = 3;
	defparam lut_21150.mask = 8'h45;

	lut_sub lut_21160 ({g592, g590, g547, g251}, g1706);
	defparam lut_21160.LUT_SIZE = 4;
	defparam lut_21160.mask = 16'hfcfd;

	lut_sub lut_21180 ({g592, g590, g462, g251}, g1707);
	defparam lut_21180.LUT_SIZE = 4;
	defparam lut_21180.mask = 16'hfcfd;

	lut_sub lut_21198 ({g1709, g1710}, g1708);
	defparam lut_21198.LUT_SIZE = 2;
	defparam lut_21198.mask = 4'b1000;

	lut_sub lut_21204 ({g134, g1711}, g1709);
	defparam lut_21204.LUT_SIZE = 2;
	defparam lut_21204.mask = 4'b0100;

	lut_sub lut_21210 ({g134, g1714}, g1710);
	defparam lut_21210.LUT_SIZE = 2;
	defparam lut_21210.mask = 4'b0001;

	lut_sub lut_21216 ({g1712, g1713}, g1711);
	defparam lut_21216.LUT_SIZE = 2;
	defparam lut_21216.mask = 4'b1000;

	lut_sub lut_21222 ({g100, g1717}, g1712);
	defparam lut_21222.LUT_SIZE = 2;
	defparam lut_21222.mask = 4'b0100;

	lut_sub lut_21228 ({g100, g1718}, g1713);
	defparam lut_21228.LUT_SIZE = 2;
	defparam lut_21228.mask = 4'b0001;

	lut_sub lut_21234 ({g1715, g1716}, g1714);
	defparam lut_21234.LUT_SIZE = 2;
	defparam lut_21234.mask = 4'b1000;

	lut_sub lut_21240 ({g100, g1719}, g1715);
	defparam lut_21240.LUT_SIZE = 2;
	defparam lut_21240.mask = 4'b0100;

	lut_sub lut_21246 ({g100, g1720}, g1716);
	defparam lut_21246.LUT_SIZE = 2;
	defparam lut_21246.mask = 4'b0001;

	lut_sub lut_21253 ({g164, g13, g251}, g1717);
	defparam lut_21253.LUT_SIZE = 3;
	defparam lut_21253.mask = 8'hfe;

	lut_sub lut_21267 ({g164, g13, g18, g251}, g1718);
	defparam lut_21267.LUT_SIZE = 4;
	defparam lut_21267.mask = 16'hfff2;

	lut_sub lut_21287 ({g164, g13, g115, g251}, g1719);
	defparam lut_21287.LUT_SIZE = 4;
	defparam lut_21287.mask = 16'hfff2;

	lut_sub lut_21305 ({g164, g13}, g1720);
	defparam lut_21305.LUT_SIZE = 2;
	defparam lut_21305.mask = 4'b1110;

	lut_sub lut_21313 ({g171, g1722}, g1721);
	defparam lut_21313.LUT_SIZE = 2;
	defparam lut_21313.mask = 4'b1000;

	lut_sub lut_21319 ({g171, g1723}, g1722);
	defparam lut_21319.LUT_SIZE = 2;
	defparam lut_21319.mask = 4'b0100;

	lut_sub lut_21325 ({g1724, g1725}, g1723);
	defparam lut_21325.LUT_SIZE = 2;
	defparam lut_21325.mask = 4'b1000;

	lut_sub lut_21330 ({i_10_, g1726}, g1724);
	defparam lut_21330.LUT_SIZE = 2;
	defparam lut_21330.mask = 4'b0100;

	lut_sub lut_21335 ({i_10_, g1727}, g1725);
	defparam lut_21335.LUT_SIZE = 2;
	defparam lut_21335.mask = 4'b0001;

	lut_sub lut_21340 ({i_9_, i_11_, g251, i_15_}, g1726);
	defparam lut_21340.LUT_SIZE = 4;
	defparam lut_21340.mask = 16'hffef;

	lut_sub lut_21359 ({i_9_, i_11_, g285, i_15_}, g1727);
	defparam lut_21359.LUT_SIZE = 4;
	defparam lut_21359.mask = 16'hffbf;

	lut_sub lut_21379 ({g1729, g1730}, g1728);
	defparam lut_21379.LUT_SIZE = 2;
	defparam lut_21379.mask = 4'b1000;

	lut_sub lut_21385 ({g465, g1731}, g1729);
	defparam lut_21385.LUT_SIZE = 2;
	defparam lut_21385.mask = 4'b0100;

	lut_sub lut_21391 ({g465, g1732}, g1730);
	defparam lut_21391.LUT_SIZE = 2;
	defparam lut_21391.mask = 4'b0001;

	lut_sub lut_21397 ({g89, g99}, g1731);
	defparam lut_21397.LUT_SIZE = 2;
	defparam lut_21397.mask = 4'b0010;

	lut_sub lut_21403 ({g1733, g1734}, g1732);
	defparam lut_21403.LUT_SIZE = 2;
	defparam lut_21403.mask = 4'b1000;

	lut_sub lut_21409 ({g89, g1735}, g1733);
	defparam lut_21409.LUT_SIZE = 2;
	defparam lut_21409.mask = 4'b0100;

	lut_sub lut_21415 ({g89, g1736}, g1734);
	defparam lut_21415.LUT_SIZE = 2;
	defparam lut_21415.mask = 4'b0001;

	lut_sub lut_21423 ({g468, g467, g475, g462}, g1735);
	defparam lut_21423.LUT_SIZE = 4;
	defparam lut_21423.mask = 16'h0001;

	lut_sub lut_21429 ({g99, g462}, g1736);
	defparam lut_21429.LUT_SIZE = 2;
	defparam lut_21429.mask = 4'b1101;

	lut_sub lut_21437 ({g1738, g1739}, g1737);
	defparam lut_21437.LUT_SIZE = 2;
	defparam lut_21437.mask = 4'b1000;

	lut_sub lut_21443 ({g477, g1740}, g1738);
	defparam lut_21443.LUT_SIZE = 2;
	defparam lut_21443.mask = 4'b0100;

	lut_sub lut_21449 ({g477, g1741}, g1739);
	defparam lut_21449.LUT_SIZE = 2;
	defparam lut_21449.mask = 4'b0001;

	lut_sub lut_21455 ({g118, g1744}, g1740);
	defparam lut_21455.LUT_SIZE = 2;
	defparam lut_21455.mask = 4'b0100;

	lut_sub lut_21461 ({g1742, g1743}, g1741);
	defparam lut_21461.LUT_SIZE = 2;
	defparam lut_21461.mask = 4'b1000;

	lut_sub lut_21467 ({g118, g1745}, g1742);
	defparam lut_21467.LUT_SIZE = 2;
	defparam lut_21467.mask = 4'b0100;

	lut_sub lut_21473 ({g118, g1746}, g1743);
	defparam lut_21473.LUT_SIZE = 2;
	defparam lut_21473.mask = 4'b0001;

	lut_sub lut_21481 ({g491, g494, g134, g492}, g1744);
	defparam lut_21481.LUT_SIZE = 4;
	defparam lut_21481.mask = 16'h0004;

	lut_sub lut_21488 ({g491, g494, g492}, g1745);
	defparam lut_21488.LUT_SIZE = 3;
	defparam lut_21488.mask = 8'h01;

	lut_sub lut_21496 ({g491, g494, g481, g492}, g1746);
	defparam lut_21496.LUT_SIZE = 4;
	defparam lut_21496.mask = 16'h0001;

	lut_sub lut_21502 ({g145, g1748}, g1747);
	defparam lut_21502.LUT_SIZE = 2;
	defparam lut_21502.mask = 4'b0010;

	lut_sub lut_21508 ({g145, g1749}, g1748);
	defparam lut_21508.LUT_SIZE = 2;
	defparam lut_21508.mask = 4'b0001;

	lut_sub lut_21514 ({g1750, g1751}, g1749);
	defparam lut_21514.LUT_SIZE = 2;
	defparam lut_21514.mask = 4'b1000;

	lut_sub lut_21519 ({i_15_, g1752}, g1750);
	defparam lut_21519.LUT_SIZE = 2;
	defparam lut_21519.mask = 4'b0100;

	lut_sub lut_21524 ({i_15_, g1753}, g1751);
	defparam lut_21524.LUT_SIZE = 2;
	defparam lut_21524.mask = 4'b0001;

	lut_sub lut_21529 ({i_10_, i_9_, g48, i_11_}, g1752);
	defparam lut_21529.LUT_SIZE = 4;
	defparam lut_21529.mask = 16'hbb7f;

	lut_sub lut_21546 ({i_10_, i_9_, g91, i_11_}, g1753);
	defparam lut_21546.LUT_SIZE = 4;
	defparam lut_21546.mask = 16'hf37f;

	lut_sub lut_21564 ({g91, g1755}, g1754);
	defparam lut_21564.LUT_SIZE = 2;
	defparam lut_21564.mask = 4'b1000;

	lut_sub lut_21570 ({g91, g1756}, g1755);
	defparam lut_21570.LUT_SIZE = 2;
	defparam lut_21570.mask = 4'b0100;

	lut_sub lut_21576 ({g1757, g1758}, g1756);
	defparam lut_21576.LUT_SIZE = 2;
	defparam lut_21576.mask = 4'b1000;

	lut_sub lut_21581 ({i_10_, g1759}, g1757);
	defparam lut_21581.LUT_SIZE = 2;
	defparam lut_21581.mask = 4'b0100;

	lut_sub lut_21586 ({i_10_, g1760}, g1758);
	defparam lut_21586.LUT_SIZE = 2;
	defparam lut_21586.mask = 4'b0001;

	lut_sub lut_21591 ({i_15_, i_11_, g145, i_9_}, g1759);
	defparam lut_21591.LUT_SIZE = 4;
	defparam lut_21591.mask = 16'h4eff;

	lut_sub lut_21607 ({i_15_, i_11_, g151, i_9_}, g1760);
	defparam lut_21607.LUT_SIZE = 4;
	defparam lut_21607.mask = 16'hfeff;

	lut_sub lut_21627 ({g13, g1762}, g1761);
	defparam lut_21627.LUT_SIZE = 2;
	defparam lut_21627.mask = 4'b0010;

	lut_sub lut_21633 ({g13, g1763}, g1762);
	defparam lut_21633.LUT_SIZE = 2;
	defparam lut_21633.mask = 4'b0001;

	lut_sub lut_21639 ({g1764, g1765}, g1763);
	defparam lut_21639.LUT_SIZE = 2;
	defparam lut_21639.mask = 4'b1000;

	lut_sub lut_21644 ({i_9_, g1766}, g1764);
	defparam lut_21644.LUT_SIZE = 2;
	defparam lut_21644.mask = 4'b0100;

	lut_sub lut_21649 ({i_9_, g1767}, g1765);
	defparam lut_21649.LUT_SIZE = 2;
	defparam lut_21649.mask = 4'b0001;

	lut_sub lut_21654 ({i_15_, i_10_, g112, i_11_}, g1766);
	defparam lut_21654.LUT_SIZE = 4;
	defparam lut_21654.mask = 16'hfeff;

	lut_sub lut_21673 ({i_15_, i_10_, g151, i_11_}, g1767);
	defparam lut_21673.LUT_SIZE = 4;
	defparam lut_21673.mask = 16'hfdff;

	lut_sub lut_21693 ({g91, g1769}, g1768);
	defparam lut_21693.LUT_SIZE = 2;
	defparam lut_21693.mask = 4'b1000;

	lut_sub lut_21699 ({g91, g1770}, g1769);
	defparam lut_21699.LUT_SIZE = 2;
	defparam lut_21699.mask = 4'b0100;

	lut_sub lut_21705 ({g1771, g1772}, g1770);
	defparam lut_21705.LUT_SIZE = 2;
	defparam lut_21705.mask = 4'b1000;

	lut_sub lut_21710 ({i_10_, g1773}, g1771);
	defparam lut_21710.LUT_SIZE = 2;
	defparam lut_21710.mask = 4'b0100;

	lut_sub lut_21715 ({i_10_, g1774}, g1772);
	defparam lut_21715.LUT_SIZE = 2;
	defparam lut_21715.mask = 4'b0001;

	lut_sub lut_21720 ({i_15_, i_9_, g109, i_11_}, g1773);
	defparam lut_21720.LUT_SIZE = 4;
	defparam lut_21720.mask = 16'hdfff;

	lut_sub lut_21739 ({i_15_, i_9_, g136, i_11_}, g1774);
	defparam lut_21739.LUT_SIZE = 4;
	defparam lut_21739.mask = 16'hfeff;

	lut_sub lut_21759 ({g91, g1776}, g1775);
	defparam lut_21759.LUT_SIZE = 2;
	defparam lut_21759.mask = 4'b1000;

	lut_sub lut_21765 ({g91, g1777}, g1776);
	defparam lut_21765.LUT_SIZE = 2;
	defparam lut_21765.mask = 4'b0100;

	lut_sub lut_21771 ({g1778, g1779}, g1777);
	defparam lut_21771.LUT_SIZE = 2;
	defparam lut_21771.mask = 4'b1000;

	lut_sub lut_21776 ({i_9_, g1780}, g1778);
	defparam lut_21776.LUT_SIZE = 2;
	defparam lut_21776.mask = 4'b0100;

	lut_sub lut_21781 ({i_9_, g1781}, g1779);
	defparam lut_21781.LUT_SIZE = 2;
	defparam lut_21781.mask = 4'b0001;

	lut_sub lut_21786 ({i_15_, i_10_, g136, i_11_}, g1780);
	defparam lut_21786.LUT_SIZE = 4;
	defparam lut_21786.mask = 16'hffef;

	lut_sub lut_21805 ({i_15_, i_10_, g151, i_11_}, g1781);
	defparam lut_21805.LUT_SIZE = 4;
	defparam lut_21805.mask = 16'hffef;

	lut_sub lut_21825 ({g1783, g1784}, g1782);
	defparam lut_21825.LUT_SIZE = 2;
	defparam lut_21825.mask = 4'b1000;

	lut_sub lut_21831 ({g132, g1785}, g1783);
	defparam lut_21831.LUT_SIZE = 2;
	defparam lut_21831.mask = 4'b0100;

	lut_sub lut_21837 ({g132, g1786}, g1784);
	defparam lut_21837.LUT_SIZE = 2;
	defparam lut_21837.mask = 4'b0001;

	lut_sub lut_21843 ({g109, g1789}, g1785);
	defparam lut_21843.LUT_SIZE = 2;
	defparam lut_21843.mask = 4'b0100;

	lut_sub lut_21849 ({g1787, g1788}, g1786);
	defparam lut_21849.LUT_SIZE = 2;
	defparam lut_21849.mask = 4'b1000;

	lut_sub lut_21855 ({g109, g1790}, g1787);
	defparam lut_21855.LUT_SIZE = 2;
	defparam lut_21855.mask = 4'b0100;

	lut_sub lut_21861 ({g109, g1791}, g1788);
	defparam lut_21861.LUT_SIZE = 2;
	defparam lut_21861.mask = 4'b0001;

	lut_sub lut_21869 ({g96, g133, g99, g120}, g1789);
	defparam lut_21869.LUT_SIZE = 4;
	defparam lut_21869.mask = 16'h0c0d;

	lut_sub lut_21881 ({g96, g133, g99, g120}, g1790);
	defparam lut_21881.LUT_SIZE = 4;
	defparam lut_21881.mask = 16'h0c0d;

	lut_sub lut_21893 ({g96, g133, g103, g120}, g1791);
	defparam lut_21893.LUT_SIZE = 4;
	defparam lut_21893.mask = 16'h0001;


endmodule