module alu4_qmap_map (sk, n, j, k, l, i, a, e, m, b, f, c, g, d, h, o, p, q, r, s, t, u, v);

	input n;
	input j;
	input k;
	input l;
	input i;
	input a;
	input e;
	input m;
	input b;
	input f;
	input c;
	input g;
	input d;
	input h;
	output o;
	output p;
	output q;
	output r;
	output s;
	output t;
	output u;
	output v;



	wire g163, g121, g179, g1, g2, g3, g4, g182, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17;
	wire g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37, g38;
	wire g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57, g206, g58;
	wire g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g80;
	wire g81, g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101;
	wire g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g122, g123;
	wire g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144;
	wire g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159, g160, g161, g164, g165, g166, g167;
	wire g168, g169, g170, g171, g183, g172, g173, g174, g175, g176, g178, g180, g181, g184, g185, g186, g189, g187, g188, g190, g191;
	wire g192, g194, g195, g196, g199, g197, g198, g202, g203, g200, g201, g204, g205, g207, g208, g209, g212, g210, g211, g215, g216;
	wire g213, g214, g217, g218, g220, g221, g222, g225, g223, g224, g228, g229, g226, g227, g230, g231;

	lut_sub lut_5 ({g163}, s);
	defparam lut_5.LUT_SIZE = 1;
	defparam lut_5.mask = 2'b10;

	lut_sub lut_9 ({g121}, t);
	defparam lut_9.LUT_SIZE = 1;
	defparam lut_9.mask = 2'b01;

	lut_sub lut_13 ({g179}, v);
	defparam lut_13.LUT_SIZE = 1;
	defparam lut_13.mask = 2'b10;

	lut_sub lut_17 ({k, l}, g1);
	defparam lut_17.LUT_SIZE = 2;
	defparam lut_17.mask = 4'b0010;

	lut_sub lut_21 ({k, l, n, i, j}, g2);
	defparam lut_21.LUT_SIZE = 5;
	defparam lut_21.mask = 32'h04041124;

	lut_sub lut_30 ({k, l, n, i, j}, g3);
	defparam lut_30.LUT_SIZE = 5;
	defparam lut_30.mask = 32'hc0800000;

	lut_sub lut_36 ({k, l, n, i, j}, g4);
	defparam lut_36.LUT_SIZE = 5;
	defparam lut_36.mask = 32'h20000202;

	lut_sub lut_43 ({k, l, i, a, e, g182}, g5);
	defparam lut_43.LUT_SIZE = 6;
	defparam lut_43.mask = 64'h55aa5d3caaccff5d;

	lut_sub lut_85 ({k, l, i, a, e, g182}, g6);
	defparam lut_85.LUT_SIZE = 6;
	defparam lut_85.mask = 64'h00003300c0053305;

	lut_sub lut_103 ({n, i, j, g1}, g7);
	defparam lut_103.LUT_SIZE = 4;
	defparam lut_103.mask = 16'h0004;

	lut_sub lut_107 ({i, j}, g8);
	defparam lut_107.LUT_SIZE = 2;
	defparam lut_107.mask = 4'b0001;

	lut_sub lut_113 ({n, g8, g1}, g9);
	defparam lut_113.LUT_SIZE = 3;
	defparam lut_113.mask = 8'h01;

	lut_sub lut_118 ({n, i, j, g1}, g10);
	defparam lut_118.LUT_SIZE = 4;
	defparam lut_118.mask = 16'h0040;

	lut_sub lut_122 ({n, i, j}, g11);
	defparam lut_122.LUT_SIZE = 3;
	defparam lut_122.mask = 8'h04;

	lut_sub lut_127 ({l, g11}, g12);
	defparam lut_127.LUT_SIZE = 2;
	defparam lut_127.mask = 4'b0001;

	lut_sub lut_135 ({a, g182, g9, g10, g12}, g13);
	defparam lut_135.LUT_SIZE = 5;
	defparam lut_135.mask = 32'hccaa88a0;

	lut_sub lut_152 ({a, e, g7, g13}, g14);
	defparam lut_152.LUT_SIZE = 4;
	defparam lut_152.mask = 16'h5554;

	lut_sub lut_163 ({k, g12}, g15);
	defparam lut_163.LUT_SIZE = 2;
	defparam lut_163.mask = 4'b0100;

	lut_sub lut_170 ({a, e, g7, g13, g15}, g16);
	defparam lut_170.LUT_SIZE = 5;
	defparam lut_170.mask = 32'h03030355;

	lut_sub lut_183 ({k, i, j}, g17);
	defparam lut_183.LUT_SIZE = 3;
	defparam lut_183.mask = 8'h40;

	lut_sub lut_188 ({l, g17}, g18);
	defparam lut_188.LUT_SIZE = 2;
	defparam lut_188.mask = 4'b0001;

	lut_sub lut_193 ({l, i, j, a, e, g182}, g19);
	defparam lut_193.LUT_SIZE = 6;
	defparam lut_193.mask = 64'h0f5f3c000a003c00;

	lut_sub lut_217 ({k, l, i, j, a, g182}, g20);
	defparam lut_217.LUT_SIZE = 6;
	defparam lut_217.mask = 64'h0000400000006664;

	lut_sub lut_233 ({k, g14, g16, g18, g19, g20}, g21);
	defparam lut_233.LUT_SIZE = 6;
	defparam lut_233.mask = 64'h80888880a0aaaaa0;

	lut_sub lut_254 ({l, n, j}, g22);
	defparam lut_254.LUT_SIZE = 3;
	defparam lut_254.mask = 8'h20;

	lut_sub lut_259 ({k, i, g22}, g23);
	defparam lut_259.LUT_SIZE = 3;
	defparam lut_259.mask = 8'h01;

	lut_sub lut_266 ({g182, g16, g23}, g24);
	defparam lut_266.LUT_SIZE = 3;
	defparam lut_266.mask = 8'h14;

	lut_sub lut_273 ({k, l, n, g8, a, g14}, g25);
	defparam lut_273.LUT_SIZE = 6;
	defparam lut_273.mask = 64'h000000000005000c;

	lut_sub lut_281 ({i, g22}, g26);
	defparam lut_281.LUT_SIZE = 2;
	defparam lut_281.mask = 4'b0100;

	lut_sub lut_285 ({k, l, n, i, j}, g27);
	defparam lut_285.LUT_SIZE = 5;
	defparam lut_285.mask = 32'h00010400;

	lut_sub lut_291 ({i, g22}, g28);
	defparam lut_291.LUT_SIZE = 2;
	defparam lut_291.mask = 4'b0001;

	lut_sub lut_298 ({k, e, g182, g27, g28}, g29);
	defparam lut_298.LUT_SIZE = 5;
	defparam lut_298.mask = 32'h30753030;

	lut_sub lut_315 ({k, a, g14, g26, g29}, g30);
	defparam lut_315.LUT_SIZE = 5;
	defparam lut_315.mask = 32'haaa88aa8;

	lut_sub lut_335 ({n, g21, g24, g25, g30}, g31);
	defparam lut_335.LUT_SIZE = 5;
	defparam lut_335.mask = 32'hbfbfffbf;

	lut_sub lut_367 ({k, n, i}, g32);
	defparam lut_367.LUT_SIZE = 3;
	defparam lut_367.mask = 8'h80;

	lut_sub lut_371 ({k, l, n, i, j}, g33);
	defparam lut_371.LUT_SIZE = 5;
	defparam lut_371.mask = 32'h01000080;

	lut_sub lut_376 ({k, l, n, i, j}, g34);
	defparam lut_376.LUT_SIZE = 5;
	defparam lut_376.mask = 32'h00504050;

	lut_sub lut_384 ({k, l, n, i, j}, g35);
	defparam lut_384.LUT_SIZE = 5;
	defparam lut_384.mask = 32'h008000f0;

	lut_sub lut_395 ({g33, a, e, g34, g35}, g36);
	defparam lut_395.LUT_SIZE = 5;
	defparam lut_395.mask = 32'hffa80000;

	lut_sub lut_412 ({e, g32, g182, g36}, g37);
	defparam lut_412.LUT_SIZE = 4;
	defparam lut_412.mask = 16'haaab;

	lut_sub lut_424 ({k, l, n, i, j}, g38);
	defparam lut_424.LUT_SIZE = 5;
	defparam lut_424.mask = 32'h00000008;

	lut_sub lut_429 ({a, e, g1, f, b}, g39);
	defparam lut_429.LUT_SIZE = 5;
	defparam lut_429.mask = 32'h46884646;

	lut_sub lut_445 ({g2, g3, f, b}, g40);
	defparam lut_445.LUT_SIZE = 4;
	defparam lut_445.mask = 16'h0ace;

	lut_sub lut_455 ({k, l, n, i, j}, g41);
	defparam lut_455.LUT_SIZE = 5;
	defparam lut_455.mask = 32'h00098a00;

	lut_sub lut_464 ({n, i, a, e, g1}, g42);
	defparam lut_464.LUT_SIZE = 5;
	defparam lut_464.mask = 32'h00001000;

	lut_sub lut_471 ({g4, f, b, g41, g42}, g43);
	defparam lut_471.LUT_SIZE = 5;
	defparam lut_471.mask = 32'h00070fff;

	lut_sub lut_494 ({a, g11, g38, g39, g40, g43}, g44);
	defparam lut_494.LUT_SIZE = 6;
	defparam lut_494.mask = 64'h77777f7f77ff7fff;

	lut_sub lut_553 ({g7, f}, g45);
	defparam lut_553.LUT_SIZE = 2;
	defparam lut_553.mask = 4'b0001;

	lut_sub lut_562 ({g9, g10, g12, b, g44, g45}, g46);
	defparam lut_562.LUT_SIZE = 6;
	defparam lut_562.mask = 64'hfac03200f8c03000;

	lut_sub lut_586 ({g15, f, b}, g47);
	defparam lut_586.LUT_SIZE = 3;
	defparam lut_586.mask = 8'h01;

	lut_sub lut_593 ({g7, g46, g47}, g48);
	defparam lut_593.LUT_SIZE = 3;
	defparam lut_593.mask = 8'ha8;

	lut_sub lut_599 ({k, l, i, j, a, e}, g49);
	defparam lut_599.LUT_SIZE = 6;
	defparam lut_599.mask = 64'h0000010000000000;

	lut_sub lut_604 ({a, g182}, g50);
	defparam lut_604.LUT_SIZE = 2;
	defparam lut_604.mask = 4'b0001;

	lut_sub lut_608 ({k, l, i, j}, g51);
	defparam lut_608.LUT_SIZE = 4;
	defparam lut_608.mask = 16'h080e;

	lut_sub lut_618 ({g50, b, g44, g51}, g52);
	defparam lut_618.LUT_SIZE = 4;
	defparam lut_618.mask = 16'h0040;

	lut_sub lut_622 ({k, l, i, j}, g53);
	defparam lut_622.LUT_SIZE = 4;
	defparam lut_622.mask = 16'h880e;

	lut_sub lut_631 ({l, g17}, g54);
	defparam lut_631.LUT_SIZE = 2;
	defparam lut_631.mask = 4'b0100;

	lut_sub lut_635 ({k, l, i, j}, g55);
	defparam lut_635.LUT_SIZE = 4;
	defparam lut_635.mask = 16'h4140;

	lut_sub lut_644 ({g182, g54, g55}, g56);
	defparam lut_644.LUT_SIZE = 3;
	defparam lut_644.mask = 8'h37;

	lut_sub lut_653 ({k, l, g8}, g57);
	defparam lut_653.LUT_SIZE = 3;
	defparam lut_653.mask = 8'h80;

	lut_sub lut_662 ({n, g46, g48, g49, g52, g206}, g58);
	defparam lut_662.LUT_SIZE = 6;
	defparam lut_662.mask = 64'h000000007777777f;

	lut_sub lut_695 ({g182, g16, g23, g44, g48}, g59);
	defparam lut_695.LUT_SIZE = 5;
	defparam lut_695.mask = 32'h09090906;

	lut_sub lut_707 ({k, n, g8}, g60);
	defparam lut_707.LUT_SIZE = 3;
	defparam lut_707.mask = 8'h01;

	lut_sub lut_713 ({l, a, g14, b, g46}, g61);
	defparam lut_713.LUT_SIZE = 5;
	defparam lut_713.mask = 32'ha5a5cc33;

	lut_sub lut_734 ({g182, g44}, g62);
	defparam lut_734.LUT_SIZE = 2;
	defparam lut_734.mask = 4'b1000;

	lut_sub lut_739 ({k, i, g22, f}, g63);
	defparam lut_739.LUT_SIZE = 4;
	defparam lut_739.mask = 16'h0100;

	lut_sub lut_743 ({l, a, e, f, b}, g64);
	defparam lut_743.LUT_SIZE = 5;
	defparam lut_743.mask = 32'h66616669;

	lut_sub lut_761 ({k, n, i, j}, g65);
	defparam lut_761.LUT_SIZE = 4;
	defparam lut_761.mask = 16'h0200;

	lut_sub lut_770 ({g27, g62, g63, g64, g65}, g66);
	defparam lut_770.LUT_SIZE = 5;
	defparam lut_770.mask = 32'he0e0e000;

	lut_sub lut_783 ({a, e, g15}, g67);
	defparam lut_783.LUT_SIZE = 3;
	defparam lut_783.mask = 8'h01;

	lut_sub lut_788 ({k, l, g11}, g68);
	defparam lut_788.LUT_SIZE = 3;
	defparam lut_788.mask = 8'h10;

	lut_sub lut_792 ({l, i, a, e}, g69);
	defparam lut_792.LUT_SIZE = 4;
	defparam lut_792.mask = 16'h0010;

	lut_sub lut_802 ({g7, g67, g46, g47, g68, g69}, g70);
	defparam lut_802.LUT_SIZE = 6;
	defparam lut_802.mask = 64'h3503050035330500;

	lut_sub lut_826 ({k, a, g14, g26, b, g46}, g71);
	defparam lut_826.LUT_SIZE = 6;
	defparam lut_826.mask = 64'h0101020109090609;

	lut_sub lut_846 ({g60, g61, g66, g70, g71}, g72);
	defparam lut_846.LUT_SIZE = 5;
	defparam lut_846.mask = 32'h08080800;

	lut_sub lut_855 ({g58, g59, g72}, g73);
	defparam lut_855.LUT_SIZE = 3;
	defparam lut_855.mask = 8'h40;

	lut_sub lut_860 ({k, l, i, f, b, g44}, g74);
	defparam lut_860.LUT_SIZE = 6;
	defparam lut_860.mask = 64'haa558ac3550f008a;

	lut_sub lut_890 ({k, l, i, f, b, g44}, g75);
	defparam lut_890.LUT_SIZE = 6;
	defparam lut_890.mask = 64'h00000f00c0110f11;

	lut_sub lut_909 ({g34, g35, f, b}, g76);
	defparam lut_909.LUT_SIZE = 4;
	defparam lut_909.mask = 16'h0515;

	lut_sub lut_921 ({g33, g32, f, g44, g76}, g77);
	defparam lut_921.LUT_SIZE = 5;
	defparam lut_921.mask = 32'haaa80000;

	lut_sub lut_934 ({n, j, g74, g75, g77}, g78);
	defparam lut_934.LUT_SIZE = 5;
	defparam lut_934.mask = 32'h05445555;

	lut_sub lut_952 ({n, m, g31, g73, g78}, p);
	defparam lut_952.LUT_SIZE = 5;
	defparam lut_952.mask = 32'haaaaebee;

	lut_sub lut_979 ({m, g31, g58, g59, g72}, g80);
	defparam lut_979.LUT_SIZE = 5;
	defparam lut_979.mask = 32'hff40ffff;

	lut_sub lut_1007 ({a, e, f, b}, g81);
	defparam lut_1007.LUT_SIZE = 4;
	defparam lut_1007.mask = 16'h2b22;

	lut_sub lut_1019 ({g1, g11, c, g, g81}, g82);
	defparam lut_1019.LUT_SIZE = 5;
	defparam lut_1019.mask = 32'h00080028;

	lut_sub lut_1026 ({j, g1, c, g}, g83);
	defparam lut_1026.LUT_SIZE = 4;
	defparam lut_1026.mask = 16'h0189;

	lut_sub lut_1035 ({n, i, g81, g83}, g84);
	defparam lut_1035.LUT_SIZE = 4;
	defparam lut_1035.mask = 16'h0010;

	lut_sub lut_1041 ({g2, g3, c, g}, g85);
	defparam lut_1041.LUT_SIZE = 4;
	defparam lut_1041.mask = 16'h0cae;

	lut_sub lut_1053 ({g4, g41, c, g}, g86);
	defparam lut_1053.LUT_SIZE = 4;
	defparam lut_1053.mask = 16'h0177;

	lut_sub lut_1067 ({b, g38, g84, g85, g86}, g87);
	defparam lut_1067.LUT_SIZE = 5;
	defparam lut_1067.mask = 32'h80808000;

	lut_sub lut_1075 ({g9, g12, c}, g88);
	defparam lut_1075.LUT_SIZE = 3;
	defparam lut_1075.mask = 8'hc8;

	lut_sub lut_1083 ({g7, g12, c, g}, g89);
	defparam lut_1083.LUT_SIZE = 4;
	defparam lut_1083.mask = 16'h0313;

	lut_sub lut_1096 ({g10, g82, g87, g88, g89}, g90);
	defparam lut_1096.LUT_SIZE = 5;
	defparam lut_1096.mask = 32'h2a222022;

	lut_sub lut_1110 ({a, g14, b, g46, g90}, g91);
	defparam lut_1110.LUT_SIZE = 5;
	defparam lut_1110.mask = 32'ha6a665a6;

	lut_sub lut_1131 ({g50, b, g44}, g92);
	defparam lut_1131.LUT_SIZE = 3;
	defparam lut_1131.mask = 8'h17;

	lut_sub lut_1140 ({g82, g87}, g93);
	defparam lut_1140.LUT_SIZE = 2;
	defparam lut_1140.mask = 4'b0100;

	lut_sub lut_1148 ({n, g53, g57, g92, g93}, g94);
	defparam lut_1148.LUT_SIZE = 5;
	defparam lut_1148.mask = 32'h00000f4f;

	lut_sub lut_1161 ({l, a, b, g60}, g95);
	defparam lut_1161.LUT_SIZE = 4;
	defparam lut_1161.mask = 16'h0015;

	lut_sub lut_1167 ({a, e, f, b}, g96);
	defparam lut_1167.LUT_SIZE = 4;
	defparam lut_1167.mask = 16'h1117;

	lut_sub lut_1179 ({g65, g, g95, g96}, g97);
	defparam lut_1179.LUT_SIZE = 4;
	defparam lut_1179.mask = 16'hcc48;

	lut_sub lut_1192 ({g26, c, g91, g94, g97}, g98);
	defparam lut_1192.LUT_SIZE = 5;
	defparam lut_1192.mask = 32'h00bb00fb;

	lut_sub lut_1210 ({l, g65, g, g96}, g99);
	defparam lut_1210.LUT_SIZE = 4;
	defparam lut_1210.mask = 16'h0206;

	lut_sub lut_1220 ({n, g51, g92, g93, g99}, g100);
	defparam lut_1220.LUT_SIZE = 5;
	defparam lut_1220.mask = 32'haaaaaaa8;

	lut_sub lut_1241 ({k, g26, c, g91, g100}, g101);
	defparam lut_1241.LUT_SIZE = 5;
	defparam lut_1241.mask = 32'ha0a0a0b0;

	lut_sub lut_1254 ({g15, c, g}, g102);
	defparam lut_1254.LUT_SIZE = 3;
	defparam lut_1254.mask = 8'h01;

	lut_sub lut_1261 ({g7, g90, g102}, g103);
	defparam lut_1261.LUT_SIZE = 3;
	defparam lut_1261.mask = 8'ha8;

	lut_sub lut_1273 ({g182, g7, g16, g44, g46, g47}, g104);
	defparam lut_1273.LUT_SIZE = 6;
	defparam lut_1273.mask = 64'h05050707055f077f;

	lut_sub lut_1308 ({k, g28, g, g93, g103, g104}, g105);
	defparam lut_1308.LUT_SIZE = 6;
	defparam lut_1308.mask = 64'h000000ff00006969;

	lut_sub lut_1331 ({g7, g67, g46, g47}, g106);
	defparam lut_1331.LUT_SIZE = 4;
	defparam lut_1331.mask = 16'hb2b0;

	lut_sub lut_1345 ({g68, g90, g103, g106}, g107);
	defparam lut_1345.LUT_SIZE = 4;
	defparam lut_1345.mask = 16'h0084;

	lut_sub lut_1351 ({l, a, b, g60, c}, g108);
	defparam lut_1351.LUT_SIZE = 5;
	defparam lut_1351.mask = 32'h00002000;

	lut_sub lut_1358 ({g27, g62, g93}, g109);
	defparam lut_1358.LUT_SIZE = 3;
	defparam lut_1358.mask = 8'h01;

	lut_sub lut_1366 ({l, g14, g46, g60, g90}, g110);
	defparam lut_1366.LUT_SIZE = 5;
	defparam lut_1366.mask = 32'h22210000;

	lut_sub lut_1377 ({g182, g44, g54, g55}, g111);
	defparam lut_1377.LUT_SIZE = 4;
	defparam lut_1377.mask = 16'hc888;

	lut_sub lut_1389 ({g51, g53, c, g92, g111}, g112);
	defparam lut_1389.LUT_SIZE = 5;
	defparam lut_1389.mask = 32'h55541514;

	lut_sub lut_1409 ({n, g93, g108, g109, g110, g112}, g113);
	defparam lut_1409.LUT_SIZE = 6;
	defparam lut_1409.mask = 64'hc000c0004000c000;

	lut_sub lut_1423 ({g68, g90, g103, g106}, g114);
	defparam lut_1423.LUT_SIZE = 4;
	defparam lut_1423.mask = 16'h0012;

	lut_sub lut_1434 ({g98, g101, g105, g107, g113, g114}, g115);
	defparam lut_1434.LUT_SIZE = 6;
	defparam lut_1434.mask = 64'hdfffffffffffffff;

	lut_sub lut_1501 ({k, l, i, c, g, g93}, g116);
	defparam lut_1501.LUT_SIZE = 6;
	defparam lut_1501.mask = 64'haa55ae3c55ccffae;

	lut_sub lut_1543 ({k, l, i, c, g, g93}, g117);
	defparam lut_1543.LUT_SIZE = 6;
	defparam lut_1543.mask = 64'h00003300c00a330a;

	lut_sub lut_1563 ({g34, g32, c, g93}, g118);
	defparam lut_1563.LUT_SIZE = 4;
	defparam lut_1563.mask = 16'h0a3b;

	lut_sub lut_1576 ({g33, g35, c, g, g118}, g119);
	defparam lut_1576.LUT_SIZE = 5;
	defparam lut_1576.mask = 32'h111fffff;

	lut_sub lut_1605 ({g14, g46, g90}, g120);
	defparam lut_1605.LUT_SIZE = 3;
	defparam lut_1605.mask = 8'h01;

	lut_sub lut_1609 ({d, h}, g121);
	defparam lut_1609.LUT_SIZE = 2;
	defparam lut_1609.mask = 4'b0001;

	lut_sub lut_1614 ({c, g, g81}, g122);
	defparam lut_1614.LUT_SIZE = 3;
	defparam lut_1614.mask = 8'h71;

	lut_sub lut_1622 ({k, l, i, j, g122}, g123);
	defparam lut_1622.LUT_SIZE = 5;
	defparam lut_1622.mask = 32'h00c3dc00;

	lut_sub lut_1636 ({n, g121, g123}, g124);
	defparam lut_1636.LUT_SIZE = 3;
	defparam lut_1636.mask = 8'h01;

	lut_sub lut_1640 ({n, j, h}, g125);
	defparam lut_1640.LUT_SIZE = 3;
	defparam lut_1640.mask = 8'h02;

	lut_sub lut_1644 ({k, l, n, j}, g126);
	defparam lut_1644.LUT_SIZE = 4;
	defparam lut_1644.mask = 16'hc800;

	lut_sub lut_1653 ({i, d, g122, g125, g126}, g127);
	defparam lut_1653.LUT_SIZE = 5;
	defparam lut_1653.mask = 32'h57000000;

	lut_sub lut_1662 ({g1, d, h}, g128);
	defparam lut_1662.LUT_SIZE = 3;
	defparam lut_1662.mask = 8'h26;

	lut_sub lut_1669 ({k, l, n, c, g121}, g129);
	defparam lut_1669.LUT_SIZE = 5;
	defparam lut_1669.mask = 32'h00005503;

	lut_sub lut_1680 ({g2, g4, d, h}, g130);
	defparam lut_1680.LUT_SIZE = 4;
	defparam lut_1680.mask = 16'hf850;

	lut_sub lut_1692 ({i, j, g129, g130}, g131);
	defparam lut_1692.LUT_SIZE = 4;
	defparam lut_1692.mask = 16'h4555;

	lut_sub lut_1707 ({g11, g122, g127, g128, g131}, g132);
	defparam lut_1707.LUT_SIZE = 5;
	defparam lut_1707.mask = 32'h50504050;

	lut_sub lut_1719 ({g9, g12, d}, g133);
	defparam lut_1719.LUT_SIZE = 3;
	defparam lut_1719.mask = 8'hc8;

	lut_sub lut_1727 ({g7, g12, d, h}, g134);
	defparam lut_1727.LUT_SIZE = 4;
	defparam lut_1727.mask = 16'h0313;

	lut_sub lut_1740 ({g10, g124, g132, g133, g134}, g135);
	defparam lut_1740.LUT_SIZE = 5;
	defparam lut_1740.mask = 32'h2a222022;

	lut_sub lut_1751 ({a, b, c, d}, g136);
	defparam lut_1751.LUT_SIZE = 4;
	defparam lut_1751.mask = 16'h9555;

	lut_sub lut_1766 ({l, g60, g120, g135, g136}, g137);
	defparam lut_1766.LUT_SIZE = 5;
	defparam lut_1766.mask = 32'h00c30055;

	lut_sub lut_1781 ({g7, g15, g121, g135}, g138);
	defparam lut_1781.LUT_SIZE = 4;
	defparam lut_1781.mask = 16'h0357;

	lut_sub lut_1797 ({g7, g67, g46, g47, g90, g102}, g139);
	defparam lut_1797.LUT_SIZE = 6;
	defparam lut_1797.mask = 64'hb2bb22b2b0bb0000;

	lut_sub lut_1829 ({n, g18, g135, g138, g139}, g140);
	defparam lut_1829.LUT_SIZE = 5;
	defparam lut_1829.mask = 32'h00000069;

	lut_sub lut_1838 ({g124, g132}, g141);
	defparam lut_1838.LUT_SIZE = 2;
	defparam lut_1838.mask = 4'b0100;

	lut_sub lut_1848 ({g7, g93, g103, g104, g141, g138}, g142);
	defparam lut_1848.LUT_SIZE = 6;
	defparam lut_1848.mask = 64'h0000000000909099;

	lut_sub lut_1865 ({g7, g93, g103, g104, g141, g138}, g143);
	defparam lut_1865.LUT_SIZE = 6;
	defparam lut_1865.mask = 64'h0000000066060600;

	lut_sub lut_1881 ({g53, g57, c, g92, g93, g141}, g144);
	defparam lut_1881.LUT_SIZE = 6;
	defparam lut_1881.mask = 64'hffff0000a6650000;

	lut_sub lut_1908 ({n, d}, g145);
	defparam lut_1908.LUT_SIZE = 2;
	defparam lut_1908.mask = 4'b0001;

	lut_sub lut_1917 ({n, g62, g54, g55, g93, g141}, g146);
	defparam lut_1917.LUT_SIZE = 6;
	defparam lut_1917.mask = 64'h000000000aaa08aa;

	lut_sub lut_1932 ({c, g, g96}, g147);
	defparam lut_1932.LUT_SIZE = 3;
	defparam lut_1932.mask = 8'h17;

	lut_sub lut_1941 ({l, g65, d, h, g147}, g148);
	defparam lut_1941.LUT_SIZE = 5;
	defparam lut_1941.mask = 32'h003b0069;

	lut_sub lut_1954 ({n, g51, d}, g149);
	defparam lut_1954.LUT_SIZE = 3;
	defparam lut_1954.mask = 8'h02;

	lut_sub lut_1963 ({c, g92, g93, g141, g148, g149}, g150);
	defparam lut_1963.LUT_SIZE = 6;
	defparam lut_1963.mask = 64'h8c8cc88cc88cc8c8;

	lut_sub lut_1996 ({g109, g141, g144, g145, g146, g150}, g151);
	defparam lut_1996.LUT_SIZE = 6;
	defparam lut_1996.mask = 64'h4044404440440000;

	lut_sub lut_2011 ({a, g14, b, g46, c, g90}, g152);
	defparam lut_2011.LUT_SIZE = 6;
	defparam lut_2011.mask = 64'h22b222b2b2bb22b2;

	lut_sub lut_2042 ({l, i, j, d}, g153);
	defparam lut_2042.LUT_SIZE = 4;
	defparam lut_2042.mask = 16'h4000;

	lut_sub lut_2047 ({i, j, g1, d}, g154);
	defparam lut_2047.LUT_SIZE = 4;
	defparam lut_2047.mask = 16'h2000;

	lut_sub lut_2055 ({n, g135, g152, g153, g154}, g155);
	defparam lut_2055.LUT_SIZE = 5;
	defparam lut_2055.mask = 32'h00005335;

	lut_sub lut_2072 ({g137, g140, g142, g143, g151, g155}, g156);
	defparam lut_2072.LUT_SIZE = 6;
	defparam lut_2072.mask = 64'h2000000000000000;

	lut_sub lut_2077 ({k, l, i, d, h, g141}, g157);
	defparam lut_2077.LUT_SIZE = 6;
	defparam lut_2077.mask = 64'h55aa51c3aa330051;

	lut_sub lut_2107 ({k, l, i, d, h, g141}, g158);
	defparam lut_2107.LUT_SIZE = 6;
	defparam lut_2107.mask = 64'h00003300c00a330a;

	lut_sub lut_2127 ({g33, g34, g35, d, h}, g159);
	defparam lut_2127.LUT_SIZE = 5;
	defparam lut_2127.mask = 32'hfcec0000;

	lut_sub lut_2144 ({g32, h, g141, g159}, g160);
	defparam lut_2144.LUT_SIZE = 4;
	defparam lut_2144.mask = 16'h5551;

	lut_sub lut_2157 ({n, j, g157, g158, g160}, g161);
	defparam lut_2157.LUT_SIZE = 5;
	defparam lut_2157.mask = 32'h05445555;

	lut_sub lut_2176 ({n, g80, g115, g156, g161}, r);
	defparam lut_2176.LUT_SIZE = 5;
	defparam lut_2176.mask = 32'haaaaebee;

	lut_sub lut_2199 ({d, h}, g163);
	defparam lut_2199.LUT_SIZE = 2;
	defparam lut_2199.mask = 4'b0110;

	lut_sub lut_2207 ({k, l, g8, g120, g135}, g164);
	defparam lut_2207.LUT_SIZE = 5;
	defparam lut_2207.mask = 32'h0f000100;

	lut_sub lut_2217 ({i, d, g135, g152}, g165);
	defparam lut_2217.LUT_SIZE = 4;
	defparam lut_2217.mask = 16'h0d00;

	lut_sub lut_2228 ({i, g93, g103, g104, g141, g138}, g166);
	defparam lut_2228.LUT_SIZE = 6;
	defparam lut_2228.mask = 64'h00000000dd0d0d00;

	lut_sub lut_2247 ({i, g141, g135, g138, g152}, g167);
	defparam lut_2247.LUT_SIZE = 5;
	defparam lut_2247.mask = 32'h50503300;

	lut_sub lut_2258 ({k, i, j}, g168);
	defparam lut_2258.LUT_SIZE = 3;
	defparam lut_2258.mask = 8'h8e;

	lut_sub lut_2269 ({c, g92, g93, d, g141, g168}, g169);
	defparam lut_2269.LUT_SIZE = 6;
	defparam lut_2269.mask = 64'h0404450445044545;

	lut_sub lut_2293 ({g7, g15, g17, g121, g135}, g170);
	defparam lut_2293.LUT_SIZE = 5;
	defparam lut_2293.mask = 32'h0a0b0f0f;

	lut_sub lut_2309 ({a, b, c, d}, g171);
	defparam lut_2309.LUT_SIZE = 4;
	defparam lut_2309.mask = 16'h8000;

	lut_sub lut_2316 ({k, g8, g171, g183}, g172);
	defparam lut_2316.LUT_SIZE = 4;
	defparam lut_2316.mask = 16'h5503;

	lut_sub lut_2325 ({k, l, i, j}, g173);
	defparam lut_2325.LUT_SIZE = 4;
	defparam lut_2325.mask = 16'h1140;

	lut_sub lut_2335 ({g62, g93, g141, g173}, g174);
	defparam lut_2335.LUT_SIZE = 4;
	defparam lut_2335.mask = 16'h0001;

	lut_sub lut_2344 ({l, g139, g169, g170, g172, g174}, g175);
	defparam lut_2344.LUT_SIZE = 6;
	defparam lut_2344.mask = 64'haaaaaaaa80008800;

	lut_sub lut_2371 ({j, g1, g165, g166, g167, g175}, g176);
	defparam lut_2371.LUT_SIZE = 6;
	defparam lut_2371.mask = 64'h5555400055555555;

	lut_sub lut_2404 ({n, g80, g115, g156, g164, g176}, u);
	defparam lut_2404.LUT_SIZE = 6;
	defparam lut_2404.mask = 64'h00000000bbfbbbbb;

	lut_sub lut_2433 ({a, e, g163}, g178);
	defparam lut_2433.LUT_SIZE = 3;
	defparam lut_2433.mask = 8'h82;

	lut_sub lut_2439 ({f, b, c, g, g178}, g179);
	defparam lut_2439.LUT_SIZE = 5;
	defparam lut_2439.mask = 32'hbeffffbe;

	lut_sub lut_2470 ({l, k, e, a, j, n}, g180);
	defparam lut_2470.LUT_SIZE = 6;
	defparam lut_2470.mask = 64'hb1a0011c91841100;

	lut_sub lut_2490 ({l, k, e, a, j, n}, g181);
	defparam lut_2490.LUT_SIZE = 6;
	defparam lut_2490.mask = 64'h0888374400018c44;

	lut_sub lut_2511 ({g180, g181, i}, g182);
	defparam lut_2511.LUT_SIZE = 3;
	defparam lut_2511.mask = 8'h1b;

	lut_sub lut_2520 ({g184, g185}, g183);
	defparam lut_2520.LUT_SIZE = 2;
	defparam lut_2520.mask = 4'b1000;

	lut_sub lut_2525 ({k, g186}, g184);
	defparam lut_2525.LUT_SIZE = 2;
	defparam lut_2525.mask = 4'b0100;

	lut_sub lut_2530 ({k, g189}, g185);
	defparam lut_2530.LUT_SIZE = 2;
	defparam lut_2530.mask = 4'b0001;

	lut_sub lut_2536 ({g187, g188}, g186);
	defparam lut_2536.LUT_SIZE = 2;
	defparam lut_2536.mask = 4'b1000;

	lut_sub lut_2541 ({j, g190}, g187);
	defparam lut_2541.LUT_SIZE = 2;
	defparam lut_2541.mask = 4'b0100;

	lut_sub lut_2546 ({j, g191}, g188);
	defparam lut_2546.LUT_SIZE = 2;
	defparam lut_2546.mask = 4'b0001;

	lut_sub lut_2551 ({j, g192}, g189);
	defparam lut_2551.LUT_SIZE = 2;
	defparam lut_2551.mask = 4'b0100;

	lut_sub lut_2556 ({h, d, g147, i}, g190);
	defparam lut_2556.LUT_SIZE = 4;
	defparam lut_2556.mask = 16'h0115;

	lut_sub lut_2564 ({h, d, g12, i}, g191);
	defparam lut_2564.LUT_SIZE = 4;
	defparam lut_2564.mask = 16'h0002;

	lut_sub lut_2569 ({h, d, g147, i}, g192);
	defparam lut_2569.LUT_SIZE = 4;
	defparam lut_2569.mask = 16'h0115;

	lut_sub lut_2578 ({g194, g195}, q);
	defparam lut_2578.LUT_SIZE = 2;
	defparam lut_2578.mask = 4'b1000;

	lut_sub lut_2583 ({n, g196}, g194);
	defparam lut_2583.LUT_SIZE = 2;
	defparam lut_2583.mask = 4'b0100;

	lut_sub lut_2588 ({n, g199}, g195);
	defparam lut_2588.LUT_SIZE = 2;
	defparam lut_2588.mask = 4'b0001;

	lut_sub lut_2594 ({g197, g198}, g196);
	defparam lut_2594.LUT_SIZE = 2;
	defparam lut_2594.mask = 4'b1000;

	lut_sub lut_2599 ({j, g202}, g197);
	defparam lut_2599.LUT_SIZE = 2;
	defparam lut_2599.mask = 4'b0100;

	lut_sub lut_2604 ({j, g203}, g198);
	defparam lut_2604.LUT_SIZE = 2;
	defparam lut_2604.mask = 4'b0001;

	lut_sub lut_2610 ({g200, g201}, g199);
	defparam lut_2610.LUT_SIZE = 2;
	defparam lut_2610.mask = 4'b1000;

	lut_sub lut_2615 ({j, g204}, g200);
	defparam lut_2615.LUT_SIZE = 2;
	defparam lut_2615.mask = 4'b0100;

	lut_sub lut_2620 ({j, g205}, g201);
	defparam lut_2620.LUT_SIZE = 2;
	defparam lut_2620.mask = 4'b0001;

	lut_sub lut_2626 ({g119, g116}, g202);
	defparam lut_2626.LUT_SIZE = 2;
	defparam lut_2626.mask = 4'b0111;

	lut_sub lut_2634 ({g119, g117}, g203);
	defparam lut_2634.LUT_SIZE = 2;
	defparam lut_2634.mask = 4'b0111;

	lut_sub lut_2643 ({g119, g115, g80}, g204);
	defparam lut_2643.LUT_SIZE = 3;
	defparam lut_2643.mask = 8'h9f;

	lut_sub lut_2655 ({g119, g115, g80}, g205);
	defparam lut_2655.LUT_SIZE = 3;
	defparam lut_2655.mask = 8'h9f;

	lut_sub lut_2666 ({g207, g208}, g206);
	defparam lut_2666.LUT_SIZE = 2;
	defparam lut_2666.mask = 4'b1000;

	lut_sub lut_2672 ({g50, g209}, g207);
	defparam lut_2672.LUT_SIZE = 2;
	defparam lut_2672.mask = 4'b0100;

	lut_sub lut_2678 ({g50, g212}, g208);
	defparam lut_2678.LUT_SIZE = 2;
	defparam lut_2678.mask = 4'b0001;

	lut_sub lut_2684 ({g210, g211}, g209);
	defparam lut_2684.LUT_SIZE = 2;
	defparam lut_2684.mask = 4'b1000;

	lut_sub lut_2689 ({b, g215}, g210);
	defparam lut_2689.LUT_SIZE = 2;
	defparam lut_2689.mask = 4'b0100;

	lut_sub lut_2694 ({b, g216}, g211);
	defparam lut_2694.LUT_SIZE = 2;
	defparam lut_2694.mask = 4'b0001;

	lut_sub lut_2700 ({g213, g214}, g212);
	defparam lut_2700.LUT_SIZE = 2;
	defparam lut_2700.mask = 4'b1000;

	lut_sub lut_2705 ({b, g217}, g213);
	defparam lut_2705.LUT_SIZE = 2;
	defparam lut_2705.mask = 4'b0100;

	lut_sub lut_2710 ({b, g218}, g214);
	defparam lut_2710.LUT_SIZE = 2;
	defparam lut_2710.mask = 4'b0001;

	lut_sub lut_2717 ({g56, g51, g44}, g215);
	defparam lut_2717.LUT_SIZE = 3;
	defparam lut_2717.mask = 8'h15;

	lut_sub lut_2727 ({g56, g57, g53, g44}, g216);
	defparam lut_2727.LUT_SIZE = 4;
	defparam lut_2727.mask = 16'h2f7f;

	lut_sub lut_2744 ({g56, g44}, g217);
	defparam lut_2744.LUT_SIZE = 2;
	defparam lut_2744.mask = 4'b0001;

	lut_sub lut_2752 ({g56, g57, g53, g44}, g218);
	defparam lut_2752.LUT_SIZE = 4;
	defparam lut_2752.mask = 16'h1f5f;

	lut_sub lut_2768 ({g220, g221}, o);
	defparam lut_2768.LUT_SIZE = 2;
	defparam lut_2768.mask = 4'b1000;

	lut_sub lut_2773 ({n, g222}, g220);
	defparam lut_2773.LUT_SIZE = 2;
	defparam lut_2773.mask = 4'b0100;

	lut_sub lut_2778 ({n, g225}, g221);
	defparam lut_2778.LUT_SIZE = 2;
	defparam lut_2778.mask = 4'b0001;

	lut_sub lut_2784 ({g223, g224}, g222);
	defparam lut_2784.LUT_SIZE = 2;
	defparam lut_2784.mask = 4'b1000;

	lut_sub lut_2789 ({j, g228}, g223);
	defparam lut_2789.LUT_SIZE = 2;
	defparam lut_2789.mask = 4'b0100;

	lut_sub lut_2794 ({j, g229}, g224);
	defparam lut_2794.LUT_SIZE = 2;
	defparam lut_2794.mask = 4'b0001;

	lut_sub lut_2800 ({g226, g227}, g225);
	defparam lut_2800.LUT_SIZE = 2;
	defparam lut_2800.mask = 4'b1000;

	lut_sub lut_2805 ({j, g230}, g226);
	defparam lut_2805.LUT_SIZE = 2;
	defparam lut_2805.mask = 4'b0100;

	lut_sub lut_2810 ({j, g231}, g227);
	defparam lut_2810.LUT_SIZE = 2;
	defparam lut_2810.mask = 4'b0001;

	lut_sub lut_2816 ({g37, g5}, g228);
	defparam lut_2816.LUT_SIZE = 2;
	defparam lut_2816.mask = 4'b0111;

	lut_sub lut_2824 ({g37, g6}, g229);
	defparam lut_2824.LUT_SIZE = 2;
	defparam lut_2824.mask = 4'b0111;

	lut_sub lut_2832 ({g37, g31, m}, g230);
	defparam lut_2832.LUT_SIZE = 3;
	defparam lut_2832.mask = 8'h9f;

	lut_sub lut_2843 ({g37, g31, m}, g231);
	defparam lut_2843.LUT_SIZE = 3;
	defparam lut_2843.mask = 8'h9f;


endmodule