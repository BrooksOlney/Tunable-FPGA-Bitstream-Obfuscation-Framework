module apex4 (
	i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, 
	i_8_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, 
	o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_);

input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_;

output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_;

wire n4, n5, n6, n7, n8, n9, n3, n11, n12, n13, n14, n15, n16, n17, n10, n19, n18, n20, n22, n23, n24, n25, n26, n27, n28, n21, n30, n31, n32, n33, n34, n35, n36, n29, n38, n39, n40, n41, n42, n43, n37, n45, n46, n47, n44, n49, n50, n51, n52, n53, n54, n55, n56, n48, n57, n59, n60, n61, n62, n63, n64, n65, n66, n58, n68, n69, n70, n71, n72, n73, n74, n75, n67, n77, n78, n79, n80, n81, n82, n83, n84, n76, n85, n87, n88, n91, n92, n86, n94, n95, n96, n97, n98, n99, n93, n103, n104, n101, n102, n100, n106, n107, n108, n109, n110, n111, n112, n113, n105, n117, n118, n115, n116, n114, n120, n121, n122, n119, n124, n125, n123, n128, n129, n126, n127, n130, n131, n132, n134, n135, n136, n133, n140, n141, n138, n139, n137, n142, n143, n144, n145, n146, n147, n149, n150, n151, n148, n153, n154, n152, n157, n156, n155, n159, n160, n158, n162, n163, n164, n161, n168, n166, n167, n165, n170, n169, n171, n172, n173, n174, n175, n176, n177, n178, n181, n182, n179, n180, n184, n186, n183, n188, n189, n187, n192, n190, n191, n196, n197, n194, n195, n193, n202, n199, n200, n201, n198, n204, n205, n203, n209, n208, n206, n212, n210, n214, n213, n216, n220, n226, n227, n228, n229, n230, n231, n225, n233, n234, n235, n232, n236, n237, n238, n239, n240, n241, n242, n248, n247, n250, n251, n249, n253, n254, n255, n256, n257, n258, n252, n260, n261, n262, n263, n264, n265, n266, n259, n268, n269, n270, n271, n272, n273, n267, n275, n276, n277, n274, n279, n280, n278, n282, n283, n284, n285, n286, n281, n288, n287, n289, n291, n292, n293, n290, n295, n294, n297, n296, n298, n299, n300, n301, n302, n303, n304, n306, n305, n310, n315, n314, n317, n316, n319, n318, n322, n323, n321, n327, n325, n326, n324, n328, n329, n330, n331, n332, n333, n335, n334, n337, n336, n338, n339, n340, n341, n342, n343, n344, n346, n345, n348, n347, n350, n349, n352, n351, n354, n353, n358, n355, n359, n364, n363, n366, n367, n368, n369, n370, n371, n365, n374, n375, n373, n372, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n401, n399, n400, n404, n405, n403, n402, n409, n407, n408, n406, n411, n412, n410, n413, n414, n416, n415, n417, n421, n423, n422, n425, n424, n427, n428, n429, n430, n426, n432, n433, n435, n436, n434, n438, n439, n437, n443, n444, n441, n442, n440, n445, n446, n447, n448, n449, n453, n451, n455, n454, n458, n459, n457, n456, n463, n460, n464, n467, n466, n469, n468, n471, n472, n473, n474, n475, n470, n477, n476, n479, n480, n478, n482, n483, n481, n485, n486, n484, n488, n487, n489, n490, n491, n492, n493, n498, n499, n500, n497, n501, n502, n503, n504, n505, n506, n507, n508, n510, n509, n512, n513, n511, n514, n515, n516, n517, n518, n519, n523, n524, n525, n522, n528, n529, n531, n532, n533, n534, n535, n536, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n570, n572, n573, n574, n571, n575, n576, n577, n578, n579, n580, n581, n582, n584, n583, n586, n585, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n599, n600, n598, n602, n603, n604, n605, n601, n607, n608, n609, n610, n611, n612, n613, n615, n616, n617, n614, n618, n619, n621, n622, n620, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n641, n642, n643, n645, n646, n647, n649, n648, n650, n651, n652, n653, n654, n656, n657, n655, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n728, n729, n730, n732, n731, n733, n734, n735, n736, n737, n738, n740, n741, n739, n743, n742, n744, n745, n746, n747, n748, n750, n749, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763;

assign o_0_ =((~ i_0_) & i_0_);
 assign o_1_ = ( (~ n86) ) ;
 assign o_2_ = ( (~ n484) ) ;
 assign o_3_ = ( (~ n85) ) ;
 assign o_4_ = ( (~ n76) ) ;
 assign o_5_ = ( (~ n67) ) ;
 assign o_6_ = ( (~ n58) ) ;
 assign o_7_ = ( (~ n57) ) ;
 assign o_8_ = ( (~ n281) ) ;
 assign o_9_ = ( (~ n48) ) ;
 assign o_10_ = ( (~ n522) ) ;
 assign o_11_ = ( (~ n44) ) ;
 assign o_12_ = ( (~ n37) ) ;
 assign o_13_ = ( (~ n29) ) ;
 assign o_14_ = ( (~ n21) ) ;
 assign o_15_ = ( (~ n20) ) ;
 assign o_16_ = ( (~ n18) ) ;
 assign o_17_ = ( (~ n10) ) ;
 assign o_18_ = ( (~ n3) ) ;
 assign n4 = ( n429 ) | ( n510 ) ;
 assign n5 = ( n542 ) | ( n442 ) ;
 assign n6 = ( n411 ) | ( n543 ) ;
 assign n7 = ( n279 ) | ( n560 ) ;
 assign n8 = ( n650  &  n651  &  n394  &  n622  &  n652  &  n653  &  n648  &  n654 ) ;
 assign n9 = ( n22  &  n513 ) | ( n22  &  n512 ) ;
 assign n3 = ( n4  &  n5  &  n6  &  n7  &  n8  &  n9 ) ;
 assign n11 = ( n649  &  n499  &  n629  &  n625  &  n590 ) ;
 assign n12 = ( n288 ) | ( n595 ) ;
 assign n13 = ( n529 ) | ( n166 ) ;
 assign n14 = ( n411 ) | ( n561 ) ;
 assign n15 = ( n194 ) | ( n580 ) ;
 assign n16 = ( (~ i_6_) ) | ( n533 ) | ( n548 ) ;
 assign n17 = ( n6  &  n756 ) ;
 assign n10 = ( n5  &  n11  &  n12  &  n13  &  n14  &  n15  &  n16  &  n17 ) ;
 assign n19 = ( n658  &  n659  &  n660  &  n661  &  n655  &  n229  &  n609  &  n662 ) ;
 assign n18 = ( n11  &  n19  &  n7  &  n4 ) ;
 assign n20 = ( n8  &  n19  &  n15  &  n13 ) ;
 assign n22 = ( n149 ) | ( n546 ) | ( n512 ) ;
 assign n23 = ( n189 ) | ( n551 ) ;
 assign n24 = ( (~ i_0_) ) | ( n403 ) | ( n432 ) ;
 assign n25 = ( n149 ) | ( n565 ) ;
 assign n26 = ( n663  &  n209  &  n664  &  n626  &  n665  &  n604  &  n666 ) ;
 assign n27 = ( n424  &  n445  &  n509  &  n667  &  n668  &  n511  &  n669  &  n670 ) ;
 assign n28 = ( n501  &  n502  &  n503  &  n504  &  n505  &  n506  &  n507  &  n508 ) ;
 assign n21 = ( n22  &  n23  &  n24  &  n25  &  n26  &  n27  &  n28 ) ;
 assign n30 = ( n234  &  n338  &  n376  &  n423  &  (~ n519)  &  n559  &  n602  &  n672 ) ;
 assign n31 = ( n340  &  n514  &  n384  &  n515  &  n516  &  n517  &  n518 ) ;
 assign n32 = ( n513 ) | ( n205 ) ;
 assign n33 = ( n429 ) | ( n561 ) ;
 assign n34 = ( (~ i_0_) ) | ( n149 ) | ( n212 ) | ( n214 ) ;
 assign n35 = ( n416 ) | ( n403 ) ;
 assign n36 = ( (~ n306) ) | ( n325 ) ;
 assign n29 = ( n30  &  n31  &  n32  &  n27  &  n33  &  n34  &  n35  &  n36 ) ;
 assign n38 = ( n639  &  n598  &  n330  &  n456  &  n87  &  n673  &  n674  &  n675 ) ;
 assign n39 = ( n429 ) | ( n101 ) ;
 assign n40 = ( i_3_ ) | ( n354 ) | ( n403 ) ;
 assign n41 = ( n149 ) | ( n579 ) ;
 assign n42 = ( n323 ) | ( n562 ) ;
 assign n43 = ( n139 ) | ( n579 ) ;
 assign n37 = ( n31  &  n38  &  n39  &  n26  &  n40  &  n41  &  n42  &  n43 ) ;
 assign n45 = ( n563 ) | ( n579 ) ;
 assign n46 = ( (~ i_3_) ) | ( i_5_ ) | ( n429 ) | ( (~ n453) ) ;
 assign n47 = ( (~ i_0_) ) | ( n212 ) | ( n325 ) ;
 assign n44 = ( n45  &  n46  &  n16  &  n47  &  n28  &  n30  &  n38 ) ;
 assign n49 = ( n571  &  n148  &  n158  &  n155  &  n592  &  n593 ) ;
 assign n50 = ( n133  &  n142  &  n137  &  n143  &  n144  &  n145  &  n146  &  n147 ) ;
 assign n51 = ( n93  &  n105  &  n114  &  n119  &  n130  &  n79  &  n131  &  n132 ) ;
 assign n52 = ( n181  &  n182  &  n179 ) | ( n181  &  n182  &  n180 ) ;
 assign n53 = ( n171  &  n172  &  n173  &  n174  &  n175  &  n176  &  n177  &  n178 ) ;
 assign n54 = ( n165  &  n161  &  n587  &  n169  &  n588  &  n589  &  n590  &  n591 ) ;
 assign n55 = ( n80  &  n193  &  n206  &  (~ n216)  &  (~ n220)  &  n583  &  n585 ) ;
 assign n56 = ( n667  &  n693  &  n621  &  n694  &  n695  &  n298  &  n213  &  n692 ) ;
 assign n48 = ( n49  &  n50  &  n51  &  n52  &  n53  &  n54  &  n55  &  n56 ) ;
 assign n57 = ( n59  &  n328  &  n329  &  n324  &  n330  &  n331  &  n332  &  n333 ) ;
 assign n59 = ( n298  &  n299  &  n111  &  n300  &  n301  &  n302  &  n303  &  n304 ) ;
 assign n60 = ( n352  &  i_5_ ) | ( n352  &  n351 ) ;
 assign n61 = ( n350  &  n149 ) | ( n350  &  n179 ) | ( n350  &  n349 ) ;
 assign n62 = ( n635  &  n345  &  n347  &  n108  &  n174  &  n636 ) ;
 assign n63 = ( n110  &  n338  &  n339  &  n340  &  n341  &  n342  &  n343  &  n344 ) ;
 assign n64 = ( n165  &  n236  &  n252  &  (~ n359)  &  n363  &  n583 ) ;
 assign n65 = ( n47  &  n404  &  n724  &  n107  &  n573  &  n725 ) ;
 assign n66 = ( n23  &  n32  &  n43  &  n353  &  (~ n355)  &  n653 ) ;
 assign n58 = ( n59  &  n60  &  n61  &  n62  &  n63  &  n64  &  n65  &  n66 ) ;
 assign n68 = ( n401  &  n399 ) | ( n401  &  n400 ) ;
 assign n69 = ( n180  &  n255  &  n398 ) | ( n255  &  (~ n306)  &  n398 ) ;
 assign n70 = ( n392  &  n36  &  n393  &  n394  &  n6  &  n395  &  n396  &  n397 ) ;
 assign n71 = ( n384  &  n385  &  n386  &  n387  &  n388  &  n389  &  n390  &  n391 ) ;
 assign n72 = ( n376  &  n377  &  n378  &  n379  &  n380  &  n381  &  n382  &  n383 ) ;
 assign n73 = ( n329  &  n406  &  n402  &  n415  &  n51  &  n278 ) ;
 assign n74 = ( n645  &  n663  &  n725  &  n704  &  n14  &  n658 ) ;
 assign n75 = ( n410  &  n413  &  n414  &  n619  &  n43  &  n706 ) ;
 assign n67 = ( n68  &  n69  &  n70  &  n71  &  n72  &  n73  &  n74  &  n75 ) ;
 assign n77 = ( n225  &  n232  &  n236  &  n237  &  n238  &  n239  &  n240  &  n241 ) ;
 assign n78 = ( n287  &  n158  &  n618  &  n619 ) ;
 assign n79 = ( n128  &  n129  &  n126 ) | ( n128  &  n129  &  n127 ) ;
 assign n80 = ( n45  &  n192  &  n190 ) | ( n45  &  n192  &  n191 ) ;
 assign n81 = ( i_0_ ) | ( (~ i_2_) ) | ( n199 ) | ( n399 ) ;
 assign n82 = ( n432 ) | ( n149 ) | ( n433 ) ;
 assign n83 = ( n498  &  n733  &  n734 ) ;
 assign n84 = ( n422  &  n446  &  n426  &  n424  &  n365  &  n68  &  n328  &  n63 ) ;
 assign n76 = ( n77  &  n78  &  n79  &  n80  &  n81  &  n82  &  n83  &  n84 ) ;
 assign n85 = ( n434  &  n445  &  n440  &  n446  &  n72  &  n324  &  n447  &  n448 ) ;
 assign n87 = ( n368  &  n490  &  n102 ) | ( n368  &  n490  &  n315 ) ;
 assign n88 = ( n647  &  n487  &  n489  &  n502  &  n501  &  n624 ) ;
 assign n91 = ( n668  &  n664  &  n491 ) ;
 assign n92 = ( n608  &  n5  &  n25  &  n734  &  n253  &  n145  &  n607  &  n755 ) ;
 assign n86 = ( n54  &  n69  &  n87  &  n88  &  n91  &  n92  &  (~ n492)  &  (~ n493) ) ;
 assign n94 = ( n319 ) | ( n545 ) ;
 assign n95 = ( n429 ) | ( n400 ) ;
 assign n96 = ( n125 ) | ( n544 ) ;
 assign n97 = ( n194 ) | ( n541 ) ;
 assign n98 = ( n429  &  n279 ) | ( n195  &  n279 ) | ( n429  &  n180 ) | ( n195  &  n180 ) ;
 assign n99 = ( n687  &  n275 ) | ( n687  &  n186 ) | ( n687  &  n513 ) ;
 assign n93 = ( n94  &  n95  &  n96  &  n97  &  n98  &  n99 ) ;
 assign n103 = ( n275 ) | ( n335 ) | ( n469 ) ;
 assign n104 = ( n125 ) | ( n322 ) ;
 assign n101 = ( n416 ) | ( n115 ) ;
 assign n102 = ( i_6_ ) | ( i_7_ ) ;
 assign n100 = ( n103  &  n104  &  n101 ) | ( n103  &  n104  &  n102 ) ;
 assign n106 = ( n407 ) | ( n457 ) ;
 assign n107 = ( n126 ) | ( n547 ) ;
 assign n108 = ( n323 ) | ( n348 ) ;
 assign n109 = ( n429 ) | ( n425 ) ;
 assign n110 = ( n125 ) | ( n346 ) ;
 assign n111 = ( (~ i_6_) ) | ( (~ i_8_) ) | ( n441 ) ;
 assign n112 = ( n407 ) | ( n549 ) ;
 assign n113 = ( n100  &  n429 ) | ( n100  &  n190 ) | ( n100  &  n416 ) ;
 assign n105 = ( n106  &  n107  &  n108  &  n109  &  n110  &  n111  &  n112  &  n113 ) ;
 assign n117 = ( n411 ) | ( n438 ) ;
 assign n118 = ( n189 ) | ( n214 ) | ( n186 ) ;
 assign n115 = ( i_5_ ) | ( n535 ) ;
 assign n116 = ( n139 ) | ( (~ n306) ) ;
 assign n114 = ( n117  &  n118  &  n115 ) | ( n117  &  n118  &  n116 ) ;
 assign n120 = ( n531 ) | ( n551 ) ;
 assign n121 = ( n411 ) | ( n549 ) ;
 assign n122 = ( n429  &  n408 ) | ( n536  &  n408 ) | ( n429  &  n442 ) | ( n536  &  n442 ) ;
 assign n119 = ( n120  &  n121  &  n122 ) ;
 assign n124 = ( n139 ) | ( n416 ) ;
 assign n125 = ( i_5_ ) | ( n199 ) ;
 assign n123 = ( n124 ) | ( n125 ) ;
 assign n128 = ( n199 ) | ( n179 ) | ( n166 ) ;
 assign n129 = ( n323 ) | ( n317 ) ;
 assign n126 = ( (~ i_5_) ) | ( n535 ) ;
 assign n127 = ( n411 ) | ( n416 ) ;
 assign n130 = ( n556  &  n557  &  n123  &  n260  &  n558  &  n559 ) ;
 assign n131 = ( n691  &  n472  &  n411 ) | ( n691  &  n472  &  n154 ) ;
 assign n132 = ( n638  &  n477  &  n643  &  n615  &  n689  &  n690  &  n626  &  n688 ) ;
 assign n134 = ( n442 ) | ( n455 ) ;
 assign n135 = ( n194 ) | ( n167 ) ;
 assign n136 = ( n125  &  n115 ) | ( n562  &  n115 ) | ( n125  &  n322 ) | ( n562  &  n322 ) ;
 assign n133 = ( n134  &  n135  &  n136 ) ;
 assign n140 = ( n563 ) | ( n430 ) ;
 assign n141 = ( n533 ) | ( n180 ) ;
 assign n138 = ( n125 ) | ( n279 ) ;
 assign n139 = ( (~ i_6_) ) | ( n531 ) ;
 assign n137 = ( n140  &  n141  &  n138 ) | ( n140  &  n141  &  n139 ) ;
 assign n142 = ( n269  &  n268  &  n566 ) ;
 assign n143 = ( n125 ) | ( n348 ) ;
 assign n144 = ( n531 ) | ( n533 ) | ( n467 ) ;
 assign n145 = ( n184 ) | ( n275 ) | ( (~ n306) ) ;
 assign n146 = ( (~ i_8_)  &  n686 ) | ( n565  &  n686 ) ;
 assign n147 = ( n683  &  n684  &  n238  &  n33  &  n342  &  n629  &  n685  &  n7 ) ;
 assign n149 = ( i_7_ ) | ( i_8_ ) ;
 assign n150 = ( (~ i_6_) ) | ( n546 ) ;
 assign n151 = ( (~ i_0_) ) | ( (~ n463) ) ;
 assign n148 = ( n42  &  n149 ) | ( n42  &  n150 ) | ( n42  &  n151 ) ;
 assign n153 = ( i_6_ ) | ( (~ i_7_) ) ;
 assign n154 = ( n125 ) | ( n179 ) ;
 assign n152 = ( n153 ) | ( n154 ) ;
 assign n157 = ( n400 ) | ( n442 ) ;
 assign n156 = ( n190 ) | ( n179 ) ;
 assign n155 = ( n157  &  n156 ) | ( n157  &  n102 ) ;
 assign n159 = ( n125 ) | ( n570 ) ;
 assign n160 = ( n319 ) | ( n248 ) ;
 assign n158 = ( n159  &  n160  &  n139 ) | ( n159  &  n160  &  n101 ) ;
 assign n162 = ( n125 ) | ( n317 ) ;
 assign n163 = ( n411 ) | ( n167 ) ;
 assign n164 = ( n115  &  n156 ) | ( n191  &  n156 ) | ( n115  &  n442 ) | ( n191  &  n442 ) ;
 assign n161 = ( n162  &  n163  &  n164 ) ;
 assign n168 = ( n102 ) | ( n126 ) | ( (~ n453) ) ;
 assign n166 = ( (~ i_6_) ) | ( n189 ) ;
 assign n167 = ( n200 ) | ( n548 ) ;
 assign n165 = ( n168  &  n166 ) | ( n168  &  n167 ) ;
 assign n170 = ( n179 ) | ( n319 ) ;
 assign n169 = ( n170 ) | ( n166 ) ;
 assign n171 = ( n429 ) | ( n167 ) ;
 assign n172 = ( n115 ) | ( n248 ) ;
 assign n173 = ( n194 ) | ( n576 ) ;
 assign n174 = ( n139 ) | ( n576 ) ;
 assign n175 = ( n399 ) | ( n170 ) ;
 assign n176 = ( n275 ) | ( n150 ) | ( n483 ) ;
 assign n177 = ( n139 ) | ( n170 ) ;
 assign n178 = ( n125  &  n534 ) | ( n577  &  n534 ) | ( n125  &  n102 ) | ( n577  &  n102 ) ;
 assign n181 = ( n533 ) | ( n189 ) | ( n548 ) ;
 assign n182 = ( n16  &  n190 ) | ( n16  &  (~ n306) ) | ( n16  &  n578 ) ;
 assign n179 = ( (~ i_2_) ) | ( n295 ) ;
 assign n180 = ( n411 ) | ( n319 ) ;
 assign n184 = ( i_6_ ) | ( n482 ) ;
 assign n186 = ( (~ i_1_) ) | ( n432 ) ;
 assign n183 = ( (~ i_7_) ) | ( n184 ) | ( n186 ) ;
 assign n188 = ( i_0_ ) | ( n150 ) | ( (~ n463) ) ;
 assign n189 = ( (~ i_7_) ) | ( (~ i_8_) ) ;
 assign n187 = ( n188 ) | ( n189 ) ;
 assign n192 = ( n407 ) | ( n154 ) ;
 assign n190 = ( (~ i_5_) ) | ( n199 ) ;
 assign n191 = ( n139 ) | ( (~ n453) ) ;
 assign n196 = ( n149 ) | ( n513 ) | ( n483 ) ;
 assign n197 = ( n323 ) | ( n351 ) ;
 assign n194 = ( i_6_ ) | ( n531 ) ;
 assign n195 = ( n533 ) | ( n115 ) ;
 assign n193 = ( n196  &  n197  &  n194 ) | ( n196  &  n197  &  n195 ) ;
 assign n202 = ( n295 ) | ( n581 ) ;
 assign n199 = ( (~ i_3_) ) | ( i_4_ ) ;
 assign n200 = ( (~ i_2_) ) | ( n354 ) ;
 assign n201 = ( (~ i_6_) ) | ( i_8_ ) ;
 assign n198 = ( n202  &  n199 ) | ( n202  &  n200 ) | ( n202  &  n201 ) ;
 assign n204 = ( i_6_ ) | ( n297 ) ;
 assign n205 = ( n149 ) | ( (~ n453) ) ;
 assign n203 = ( n204 ) | ( n205 ) ;
 assign n209 = ( n319 ) | ( n577 ) ;
 assign n208 = ( i_3_ ) | ( i_4_ ) | ( i_6_ ) ;
 assign n206 = ( n189  &  n209 ) | ( n209  &  n208 ) | ( n209  &  (~ n306) ) ;
 assign n212 = ( i_2_ ) | ( (~ i_3_) ) ;
 assign n210 = ( (~ i_0_) ) | ( n184 ) | ( n212 ) ;
 assign n214 = ( (~ i_4_) ) | ( i_5_ ) | ( i_6_ ) ;
 assign n213 = ( (~ i_1_) ) | ( (~ i_7_) ) | ( n212 ) | ( n214 ) ;
 assign n216 = ( i_8_  &  (~ n210) ) | ( i_8_  &  (~ n416)  &  (~ n467) ) ;
 assign n220 = ( (~ i_5_)  &  (~ n595) ) | ( (~ i_5_)  &  (~ n407)  &  (~ n564) ) ;
 assign n226 = ( n411 ) | ( n425 ) ;
 assign n227 = ( n364 ) | ( (~ n453) ) ;
 assign n228 = ( n126 ) | ( n348 ) ;
 assign n229 = ( n166 ) | ( n561 ) ;
 assign n230 = ( n125  &  n300 ) | ( n189  &  n300 ) | ( n300  &  (~ n453) ) ;
 assign n231 = ( n275 ) | ( n101 ) ;
 assign n225 = ( n226  &  n227  &  n228  &  n229  &  n230  &  n231 ) ;
 assign n233 = ( n399 ) | ( n541 ) ;
 assign n234 = ( n138 ) | ( n166 ) ;
 assign n235 = ( n582  &  n275 ) | ( n582  &  n200 ) | ( n582  &  n433 ) ;
 assign n232 = ( n35  &  n233  &  n234  &  n235 ) ;
 assign n236 = ( n596  &  n597 ) ;
 assign n237 = ( n193  &  n710  &  n540 ) | ( n193  &  n710  &  n150 ) ;
 assign n238 = ( n319 ) | ( n429 ) | ( (~ n453) ) ;
 assign n239 = ( n323 ) | ( n346 ) ;
 assign n240 = ( n190 ) | ( n200 ) | ( n201 ) ;
 assign n241 = ( n677  &  n709  &  n663  &  n395 ) ;
 assign n242 = ( (~ n195)  &  (~ n399) ) | ( (~ n279)  &  (~ n399)  &  (~ n535) ) ;
 assign n248 = ( n166 ) | ( (~ n306) ) ;
 assign n247 = ( n248 ) | ( n126 ) ;
 assign n250 = ( n433 ) | ( n568 ) ;
 assign n251 = ( (~ i_4_) ) | ( i_5_ ) | ( n346 ) ;
 assign n249 = ( n250  &  n251  &  n184 ) | ( n250  &  n251  &  n205 ) ;
 assign n253 = ( n190 ) | ( n351 ) ;
 assign n254 = ( n531 ) | ( n575 ) ;
 assign n255 = ( n323 ) | ( n116 ) ;
 assign n256 = ( n139 ) | ( n542 ) ;
 assign n257 = ( n701  &  n528 ) | ( n701  &  n547 ) ;
 assign n258 = ( n699  &  n459  &  n700  &  n665  &  n444  &  n656  &  n97  &  n387 ) ;
 assign n252 = ( n253  &  n254  &  n255  &  n256  &  n137  &  n100  &  n257  &  n258 ) ;
 assign n260 = ( n548 ) | ( n248 ) ;
 assign n261 = ( n115 ) | ( n545 ) ;
 assign n262 = ( n534 ) | ( n411 ) ;
 assign n263 = ( n411 ) | ( n441 ) ;
 assign n264 = ( n126 ) | ( n276 ) | ( n416 ) ;
 assign n265 = ( n139 ) | ( n408 ) ;
 assign n266 = ( n534  &  n529 ) | ( n442  &  n529 ) | ( n534  &  n102 ) | ( n442  &  n102 ) ;
 assign n259 = ( n260  &  n95  &  n261  &  n262  &  n263  &  n264  &  n265  &  n266 ) ;
 assign n268 = ( n166 ) | ( n549 ) ;
 assign n269 = ( n429 ) | ( n488 ) ;
 assign n270 = ( n194 ) | ( n567 ) ;
 assign n271 = ( n115 ) | ( n595 ) ;
 assign n272 = ( n115  &  n698 ) | ( n194  &  n698 ) | ( (~ n306)  &  n698 ) ;
 assign n273 = ( n279 ) | ( n189 ) | ( n335 ) ;
 assign n267 = ( n268  &  n269  &  n270  &  n271  &  n272  &  n273 ) ;
 assign n275 = ( (~ i_7_) ) | ( i_8_ ) ;
 assign n276 = ( i_6_ ) | ( (~ i_8_) ) ;
 assign n277 = ( n533 ) | ( n319 ) ;
 assign n274 = ( n275  &  n276 ) | ( n188  &  n276 ) | ( n275  &  n277 ) | ( n188  &  n277 ) ;
 assign n279 = ( i_2_ ) | ( n295 ) ;
 assign n280 = ( i_3_ ) | ( i_5_ ) ;
 assign n278 = ( n202  &  n279 ) | ( n202  &  n194 ) | ( n202  &  n280 ) ;
 assign n282 = ( n607  &  n608  &  n609  &  n516 ) ;
 assign n283 = ( (~ i_1_)  &  n712 ) | ( n139  &  n712 ) | ( n323  &  n712 ) ;
 assign n284 = ( n331  &  n252  &  n77  &  n267  &  n274  &  n259 ) ;
 assign n285 = ( n681  &  n41  &  n647  &  n683  &  n711  &  n24 ) ;
 assign n286 = ( n33  &  n389  &  n177  &  n642  &  n657  &  n36 ) ;
 assign n281 = ( n282  &  n52  &  n278  &  n283  &  n114  &  n284  &  n285  &  n286 ) ;
 assign n288 = ( i_3_ ) | ( n482 ) ;
 assign n287 = ( n116 ) | ( n288 ) ;
 assign n289 = ( n124 ) | ( n190 ) ;
 assign n291 = ( n429 ) | ( n408 ) ;
 assign n292 = ( n149 ) | ( n208 ) | ( (~ n306) ) ;
 assign n293 = ( n194  &  n399 ) | ( n539  &  n399 ) | ( n194  &  n579 ) | ( n539  &  n579 ) ;
 assign n290 = ( n291  &  n292  &  n293 ) ;
 assign n295 = ( i_0_ ) | ( (~ i_1_) ) ;
 assign n294 = ( n150 ) | ( n275 ) | ( n295 ) | ( i_3_ ) ;
 assign n297 = ( i_3_ ) | ( (~ i_5_) ) ;
 assign n296 = ( n166 ) | ( n179 ) | ( n297 ) ;
 assign n298 = ( n540 ) | ( n214 ) ;
 assign n299 = ( n399 ) | ( n457 ) ;
 assign n300 = ( n323 ) | ( n577 ) ;
 assign n301 = ( n718  &  i_0_ ) | ( n718  &  n432 ) | ( n718  &  n403 ) ;
 assign n302 = ( i_3_ ) | ( n570 ) ;
 assign n303 = ( n290  &  n473  &  n267  &  n130  &  n78  &  n614  &  n620 ) ;
 assign n304 = ( n717  &  n176  &  n388  &  n227  &  n109  &  n145  &  n587  &  n716 ) ;
 assign n306 = ( (~ i_2_)  &  (~ n412) ) ;
 assign n305 = ( (~ n126)  &  (~ n191) ) | ( (~ n126)  &  (~ n275)  &  n306 ) ;
 assign n310 = ( (~ n180)  &  (~ n416) ) | ( (~ n288)  &  (~ n416)  &  (~ n531) ) ;
 assign n315 = ( n323 ) | ( n200 ) ;
 assign n314 = ( n315 ) | ( n149 ) ;
 assign n317 = ( (~ n306) ) | ( n407 ) ;
 assign n316 = ( n317 ) | ( n190 ) ;
 assign n319 = ( i_5_ ) | ( n528 ) ;
 assign n318 = ( n201 ) | ( n319 ) | ( (~ n453) ) ;
 assign n322 = ( n399 ) | ( (~ n453) ) ;
 assign n323 = ( (~ i_5_) ) | ( n528 ) ;
 assign n321 = ( n322 ) | ( n323 ) ;
 assign n327 = ( n689  &  n566  &  n713 ) ;
 assign n325 = ( n189 ) | ( n433 ) ;
 assign n326 = ( i_1_ ) | ( (~ n463) ) ;
 assign n324 = ( n198  &  n327  &  n325 ) | ( n198  &  n327  &  n326 ) ;
 assign n328 = ( n626  &  n627  &  n628  &  n629  &  n490  &  n630  &  n631  &  n632 ) ;
 assign n329 = ( n318  &  n321  &  n15  &  n625 ) ;
 assign n330 = ( n623  &  n390  &  n624 ) ;
 assign n331 = ( n610  &  n133  &  n611  &  n612  &  n249  &  n598  &  n601  &  n613 ) ;
 assign n332 = ( n585  &  n148  &  n232 ) ;
 assign n333 = ( n384  &  n228  &  n705  &  n720  &  n503  &  n144  &  n661  &  n719 ) ;
 assign n335 = ( (~ i_6_) ) | ( n482 ) ;
 assign n334 = ( n275 ) | ( n335 ) | ( (~ n453) ) ;
 assign n337 = ( (~ i_4_) ) | ( (~ i_5_) ) ;
 assign n336 = ( n337 ) | ( n124 ) ;
 assign n338 = ( n139 ) | ( n438 ) ;
 assign n339 = ( n200 ) | ( n180 ) ;
 assign n340 = ( n190 ) | ( n139 ) | ( n200 ) ;
 assign n341 = ( n125 ) | ( n116 ) ;
 assign n342 = ( n126 ) | ( n322 ) ;
 assign n343 = ( n4  &  n499  &  n106 ) ;
 assign n344 = ( n393  &  n381  &  n684  &  n157  &  n722  &  n375  &  n723  &  n721 ) ;
 assign n346 = ( n416 ) | ( n166 ) ;
 assign n345 = ( n346 ) | ( n190 ) ;
 assign n348 = ( (~ n306) ) | ( n411 ) ;
 assign n347 = ( n348 ) | ( n115 ) ;
 assign n350 = ( n533 ) | ( n166 ) | ( n550 ) ;
 assign n349 = ( i_6_ ) | ( n550 ) ;
 assign n352 = ( n536 ) | ( n439 ) ;
 assign n351 = ( n411 ) | ( (~ n453) ) ;
 assign n354 = ( (~ i_0_) ) | ( (~ i_1_) ) ;
 assign n353 = ( n354 ) | ( n275 ) | ( n319 ) ;
 assign n358 = ( i_1_  &  (~ i_5_) ) | ( i_1_  &  (~ n412) ) | ( i_5_  &  (~ n412) ) ;
 assign n355 = ( (~ i_4_)  &  n358  &  (~ n442) ) ;
 assign n359 = ( (~ n154)  &  (~ n411) ) | ( (~ n154)  &  (~ n439) ) ;
 assign n364 = ( n190 ) | ( n194 ) ;
 assign n363 = ( (~ n306) ) | ( n364 ) ;
 assign n366 = ( n200 ) | ( n560 ) ;
 assign n367 = ( n408 ) | ( n166 ) ;
 assign n368 = ( n125 ) | ( n594 ) ;
 assign n369 = ( n190 ) | ( n545 ) ;
 assign n370 = ( n126  &  n407 ) | ( n544  &  n407 ) | ( n126  &  n441 ) | ( n544  &  n441 ) ;
 assign n371 = ( (~ i_1_)  &  n730 ) | ( i_2_  &  n730 ) | ( n581  &  n730 ) ;
 assign n365 = ( n366  &  n367  &  n368  &  n369  &  n370  &  n371 ) ;
 assign n374 = ( n407 ) | ( n552 ) ;
 assign n375 = ( n334  &  n336  &  n633  &  n634 ) ;
 assign n373 = ( n531 ) | ( n513 ) ;
 assign n372 = ( n374  &  n375  &  n373 ) | ( n374  &  n375  &  n326 ) ;
 assign n376 = ( n194 ) | ( n552 ) ;
 assign n377 = ( n126 ) | ( n594 ) ;
 assign n378 = ( n399 ) | ( n430 ) ;
 assign n379 = ( n139 ) | ( n567 ) ;
 assign n380 = ( n411 ) | ( n541 ) ;
 assign n381 = ( n166 ) | ( n430 ) ;
 assign n382 = ( n411 ) | ( n430 ) ;
 assign n383 = ( n372  &  n290  &  n365  &  n282  &  n249  &  n731 ) ;
 assign n384 = ( n125 ) | ( n416 ) | ( n442 ) ;
 assign n385 = ( n126 ) | ( n116 ) ;
 assign n386 = ( n288 ) | ( n562 ) ;
 assign n387 = ( n411 ) | ( n567 ) ;
 assign n388 = ( n101 ) | ( n442 ) ;
 assign n389 = ( n288 ) | ( n248 ) ;
 assign n390 = ( n541 ) | ( n166 ) ;
 assign n391 = ( n299  &  n612  &  n256  &  n707  &  n728  &  n729 ) ;
 assign n392 = ( n469 ) | ( n427 ) ;
 assign n393 = ( n288 ) | ( n439 ) | ( (~ n453) ) ;
 assign n394 = ( n439 ) | ( n567 ) ;
 assign n395 = ( n139 ) | ( n457 ) ;
 assign n396 = ( n720  &  n630  &  n540 ) | ( n720  &  n630  &  n208 ) ;
 assign n397 = ( n618  &  n708  &  n722 ) ;
 assign n398 = ( n599  &  n703  &  n47 ) ;
 assign n401 = ( n275 ) | ( n416 ) | ( n214 ) ;
 assign n399 = ( i_6_ ) | ( n275 ) ;
 assign n400 = ( n279 ) | ( n126 ) ;
 assign n404 = ( n399 ) | ( n441 ) ;
 assign n405 = ( n411 ) | ( n580 ) ;
 assign n403 = ( n184 ) | ( n189 ) ;
 assign n402 = ( n404  &  n405  &  n151 ) | ( n404  &  n405  &  n403 ) ;
 assign n409 = ( (~ n306) ) | ( n548 ) | ( n578 ) ;
 assign n407 = ( (~ i_6_) ) | ( n275 ) ;
 assign n408 = ( n125 ) | ( n200 ) ;
 assign n406 = ( n409  &  n407 ) | ( n409  &  n408 ) ;
 assign n411 = ( (~ i_6_) ) | ( n149 ) ;
 assign n412 = ( (~ i_0_) ) | ( i_1_ ) ;
 assign n410 = ( n411 ) | ( n199 ) | ( n412 ) ;
 assign n413 = ( n335 ) | ( i_7_ ) | ( n151 ) ;
 assign n414 = ( n189 ) | ( n200 ) | ( n204 ) ;
 assign n416 = ( i_2_ ) | ( n354 ) ;
 assign n415 = ( n180 ) | ( n416 ) ;
 assign n417 = ( (~ n442)  &  (~ n536) ) | ( (~ n179)  &  (~ n280)  &  (~ n442) ) ;
 assign n421 = ( n351 ) | ( n115 ) ;
 assign n423 = ( n399 ) | ( n549 ) ;
 assign n422 = ( n189  &  n423 ) | ( (~ n306)  &  n423 ) | ( n349  &  n423 ) ;
 assign n425 = ( n179 ) | ( n548 ) ;
 assign n424 = ( n386  &  n194 ) | ( n386  &  n425 ) ;
 assign n427 = ( n189 ) | ( n513 ) ;
 assign n428 = ( (~ i_0_) ) | ( (~ i_2_) ) ;
 assign n429 = ( i_6_ ) | ( n149 ) ;
 assign n430 = ( n179 ) | ( n126 ) ;
 assign n426 = ( n427  &  n429 ) | ( n428  &  n429 ) | ( n427  &  n430 ) | ( n428  &  n430 ) ;
 assign n432 = ( (~ i_2_) ) | ( i_3_ ) ;
 assign n433 = ( i_6_ ) | ( n337 ) ;
 assign n435 = ( n166 ) | ( n488 ) ;
 assign n436 = ( n407  &  n531 ) | ( n579  &  n531 ) | ( n407  &  n430 ) | ( n579  &  n430 ) ;
 assign n434 = ( n435  &  n341  &  n436 ) ;
 assign n438 = ( n416 ) | ( n548 ) ;
 assign n439 = ( (~ i_6_) ) | ( (~ i_7_) ) ;
 assign n437 = ( n438 ) | ( n439 ) ;
 assign n443 = ( n190 ) | ( n348 ) ;
 assign n444 = ( n279 ) | ( n407 ) | ( n535 ) ;
 assign n441 = ( n323 ) | ( n179 ) ;
 assign n442 = ( i_6_ ) | ( n189 ) ;
 assign n440 = ( n443  &  n444  &  n441 ) | ( n443  &  n444  &  n442 ) ;
 assign n445 = ( n642  &  n437  &  n627  &  n584 ) ;
 assign n446 = ( (~ n417)  &  n421  &  n555  &  n556  &  n637  &  n638  &  n639  &  n641 ) ;
 assign n447 = ( n601  &  n206  &  n620 ) ;
 assign n448 = ( n268  &  n271  &  n711  &  n735  &  n161  &  n155  &  n736  &  n105 ) ;
 assign n449 = ( (~ n214)  &  (~ n531) ) ;
 assign n453 = ( i_2_  &  (~ n412) ) ;
 assign n451 = ( n449  &  n453 ) | ( (~ n153)  &  (~ n288)  &  n453 ) ;
 assign n455 = ( n279 ) | ( n319 ) ;
 assign n454 = ( n455 ) | ( n399 ) ;
 assign n458 = ( n139 ) | ( n536 ) ;
 assign n459 = ( n288 ) | ( n346 ) ;
 assign n457 = ( n200 ) | ( n115 ) ;
 assign n456 = ( n458  &  n459  &  n194 ) | ( n458  &  n459  &  n457 ) ;
 assign n463 = ( i_3_  &  i_2_ ) ;
 assign n460 = ( (~ n373)  &  n463 ) | ( (~ n189)  &  (~ n214)  &  n463 ) ;
 assign n464 = ( i_2_  &  (~ n460) ) | ( n280  &  (~ n460) ) | ( n429  &  (~ n460) ) ;
 assign n467 = ( (~ i_6_) ) | ( n528 ) ;
 assign n466 = ( n189  &  i_7_ ) | ( n467  &  i_7_ ) | ( n189  &  n349 ) | ( n467  &  n349 ) ;
 assign n469 = ( i_3_ ) | ( n412 ) ;
 assign n468 = ( n295  &  i_4_ ) | ( n115  &  i_4_ ) | ( n295  &  n469 ) | ( n115  &  n469 ) ;
 assign n471 = ( n107  &  (~ n451)  &  n454  &  n643  &  n645  &  n646 ) ;
 assign n472 = ( n553  &  n554  &  n555 ) ;
 assign n473 = ( n265  &  n294  &  n296 ) ;
 assign n474 = ( (~ i_1_)  &  n746  &  n748 ) | ( n464  &  n746  &  n748 ) ;
 assign n475 = ( n557  &  n711  &  n745  &  n744  &  n381  &  n120  &  n698  &  n739 ) ;
 assign n470 = ( n456  &  n402  &  n471  &  n53  &  n472  &  n473  &  n474  &  n475 ) ;
 assign n477 = ( n429 ) | ( n543 ) ;
 assign n476 = ( n477  &  n156 ) | ( n477  &  n399 ) ;
 assign n479 = ( n276 ) | ( n115 ) ;
 assign n480 = ( n125 ) | ( n194 ) ;
 assign n478 = ( (~ i_5_)  &  n479  &  n480 ) | ( n429  &  n479  &  n480 ) ;
 assign n482 = ( i_4_ ) | ( (~ i_5_) ) ;
 assign n483 = ( (~ i_0_) ) | ( i_2_ ) | ( i_3_ ) ;
 assign n481 = ( n482  &  n354 ) | ( n483  &  n354 ) | ( n482  &  n126 ) | ( n483  &  n126 ) ;
 assign n485 = ( n225  &  n49  &  n614  &  n752  &  n753  &  n751 ) ;
 assign n486 = ( n626  &  n657  &  n651  &  n650  &  n263  &  n121  &  n378  &  n749 ) ;
 assign n484 = ( n476  &  n434  &  n470  &  n71  &  n60  &  n426  &  n485  &  n486 ) ;
 assign n488 = ( n200 ) | ( n288 ) ;
 assign n487 = ( n488 ) | ( n407 ) ;
 assign n489 = ( n167 ) | ( n139 ) ;
 assign n490 = ( n411 ) | ( n488 ) ;
 assign n491 = ( n337 ) | ( n139 ) | ( n326 ) ;
 assign n492 = ( (~ n126)  &  (~ n416)  &  (~ n439) ) | ( (~ n126)  &  (~ n439)  &  n453 ) ;
 assign n493 = ( n306  &  (~ n364) ) | ( n306  &  (~ n480) ) | ( n306  &  (~ n754) ) ;
 assign n498 = ( n102 ) | ( (~ n306) ) | ( n548 ) ;
 assign n499 = ( n533 ) | ( n560 ) ;
 assign n500 = ( n323  &  n439 ) | ( n127  &  n439 ) | ( n323  &  n315 ) | ( n127  &  n315 ) ;
 assign n497 = ( n498  &  n499  &  n500 ) ;
 assign n501 = ( n125 ) | ( n248 ) ;
 assign n502 = ( n115 ) | ( n570 ) ;
 assign n503 = ( n407 ) | ( n580 ) ;
 assign n504 = ( n733  &  n149 ) | ( n733  &  n335 ) | ( n733  &  n564 ) ;
 assign n505 = ( n416 ) | ( n325 ) ;
 assign n506 = ( n471  &  n440  &  n497  &  n259  &  n571  &  n406 ) ;
 assign n507 = ( n617  &  n369  &  n162  &  n171  &  n690  &  n341 ) ;
 assign n508 = ( n291  &  n135  &  n134  &  n650  &  n649  &  n292 ) ;
 assign n510 = ( n125 ) | ( n533 ) ;
 assign n509 = ( n239  &  n411 ) | ( n239  &  n510 ) ;
 assign n512 = ( i_3_ ) | ( n532 ) ;
 assign n513 = ( i_6_ ) | ( n546 ) ;
 assign n511 = ( n512 ) | ( n513 ) ;
 assign n514 = ( n102 ) | ( n579 ) ;
 assign n515 = ( n125 ) | ( n191 ) ;
 assign n516 = ( n126 ) | ( n570 ) ;
 assign n517 = ( n677  &  n374  &  n175  &  n703  &  n159 ) ;
 assign n518 = ( n389  &  n702  &  n339  &  n758  &  n655  &  n648  &  n476  &  n62 ) ;
 assign n519 = ( (~ n190)  &  (~ n547) ) | ( (~ n190)  &  (~ n595) ) ;
 assign n523 = ( n372  &  n61  &  n70  &  n50  &  n93  &  n274 ) ;
 assign n524 = ( n759  &  n760  &  n761  &  n34  &  n367  &  n610 ) ;
 assign n525 = ( n699  &  n240  &  n717  &  n340  &  n4  &  n623 ) ;
 assign n522 = ( n470  &  n422  &  n88  &  n509  &  n497  &  n523  &  n524  &  n525 ) ;
 assign n528 = ( i_3_ ) | ( (~ i_4_) ) ;
 assign n529 = ( n279 ) | ( n323 ) ;
 assign n531 = ( i_7_ ) | ( (~ i_8_) ) ;
 assign n532 = ( i_1_ ) | ( i_0_ ) ;
 assign n533 = ( (~ i_2_) ) | ( n532 ) ;
 assign n534 = ( n323 ) | ( n533 ) ;
 assign n535 = ( (~ i_3_) ) | ( (~ i_4_) ) ;
 assign n536 = ( n126 ) | ( n200 ) ;
 assign n538 = ( i_0_ ) | ( n432 ) | ( n184 ) ;
 assign n539 = ( n319 ) | ( n416 ) ;
 assign n540 = ( n179 ) | ( n189 ) ;
 assign n541 = ( n533 ) | ( n126 ) ;
 assign n542 = ( n279 ) | ( n115 ) ;
 assign n543 = ( n279 ) | ( n288 ) ;
 assign n544 = ( n407 ) | ( n416 ) ;
 assign n545 = ( n166 ) | ( (~ n453) ) ;
 assign n546 = ( i_4_ ) | ( i_5_ ) ;
 assign n547 = ( n399 ) | ( n416 ) ;
 assign n548 = ( i_4_ ) | ( n280 ) ;
 assign n549 = ( n279 ) | ( n548 ) ;
 assign n550 = ( (~ i_3_) ) | ( (~ i_5_) ) ;
 assign n551 = ( n416 ) | ( n349 ) ;
 assign n552 = ( n179 ) | ( n115 ) ;
 assign n553 = ( n190 ) | ( n322 ) ;
 assign n554 = ( n126 ) | ( n351 ) ;
 assign n555 = ( n166 ) | ( n543 ) ;
 assign n556 = ( n139 ) | ( n552 ) ;
 assign n557 = ( n166 ) | ( n455 ) ;
 assign n558 = ( n543 ) | ( n442 ) ;
 assign n559 = ( n411 ) | ( n457 ) ;
 assign n560 = ( n407 ) | ( n319 ) ;
 assign n561 = ( n533 ) | ( n288 ) ;
 assign n562 = ( (~ n306) ) | ( n442 ) ;
 assign n563 = ( (~ i_6_) ) | ( i_7_ ) ;
 assign n564 = ( i_1_ ) | ( n432 ) ;
 assign n565 = ( (~ i_3_) ) | ( n214 ) | ( n412 ) ;
 assign n566 = ( n194 ) | ( n170 ) ;
 assign n567 = ( n279 ) | ( n190 ) ;
 assign n568 = ( n531 ) | ( n469 ) ;
 assign n570 = ( n407 ) | ( (~ n453) ) ;
 assign n572 = ( n194 ) | ( n455 ) ;
 assign n573 = ( n539 ) | ( n563 ) ;
 assign n574 = ( n319 ) | ( n322 ) ;
 assign n571 = ( n572  &  n152  &  n573  &  n574 ) ;
 assign n575 = ( n179 ) | ( n288 ) ;
 assign n576 = ( n200 ) | ( n319 ) ;
 assign n577 = ( (~ n306) ) | ( n399 ) ;
 assign n578 = ( i_6_ ) | ( i_8_ ) ;
 assign n579 = ( (~ n453) ) | ( n548 ) ;
 assign n580 = ( n190 ) | ( n533 ) ;
 assign n581 = ( i_3_ ) | ( n149 ) | ( n433 ) ;
 assign n582 = ( n6  &  n379  &  n409  &  n374  &  n435 ) ;
 assign n584 = ( n429 ) | ( n567 ) ;
 assign n583 = ( n203  &  n582  &  n198  &  n395  &  n584  &  n405 ) ;
 assign n586 = ( (~ n453) ) | ( n480 ) ;
 assign n585 = ( n183  &  n187  &  n443  &  n586 ) ;
 assign n587 = ( n407 ) | ( n430 ) ;
 assign n588 = ( n407 ) | ( n575 ) ;
 assign n589 = ( n139 ) | ( n549 ) ;
 assign n590 = ( n411 ) | ( n400 ) ;
 assign n591 = ( n139 ) | ( n425 ) ;
 assign n592 = ( n680  &  n681  &  n611  &  n682 ) ;
 assign n593 = ( n676  &  n631  &  n677  &  n678  &  n679  &  n261  &  n652  &  n270 ) ;
 assign n594 = ( (~ n306) ) | ( n429 ) ;
 assign n595 = ( n139 ) | ( n533 ) ;
 assign n596 = ( n392  &  n94  &  n702  &  n377  &  n96  &  n703  &  n704  &  n12 ) ;
 assign n597 = ( n705  &  n706  &  n693  &  n695  &  n589  &  n707  &  n708  &  n689 ) ;
 assign n599 = ( n319 ) | ( n562 ) ;
 assign n600 = ( n138 ) | ( n411 ) ;
 assign n598 = ( n405  &  n378  &  n599  &  n600  &  n553 ) ;
 assign n602 = ( (~ n306) ) | ( n560 ) ;
 assign n603 = ( n411 ) | ( n101 ) ;
 assign n604 = ( n429 ) | ( n575 ) ;
 assign n605 = ( n288 ) | ( n544 ) ;
 assign n601 = ( (~ n242)  &  n247  &  n515  &  n602  &  n603  &  n604  &  n605 ) ;
 assign n607 = ( n139 ) | ( n488 ) ;
 assign n608 = ( n190 ) | ( n248 ) ;
 assign n609 = ( n407 ) | ( n561 ) ;
 assign n610 = ( n126 ) | ( n194 ) | ( (~ n453) ) ;
 assign n611 = ( n416 ) | ( n480 ) ;
 assign n612 = ( n166 ) | ( n400 ) ;
 assign n613 = ( n554  &  n694  &  n646  &  n643  &  n679  &  n574  &  n14  &  n660 ) ;
 assign n615 = ( n319 ) | ( n116 ) ;
 assign n616 = ( n407 ) | ( n195 ) ;
 assign n617 = ( n195 ) | ( n442 ) ;
 assign n614 = ( n615  &  n380  &  n289  &  n616  &  n617  &  n376 ) ;
 assign n618 = ( n194 ) | ( n400 ) ;
 assign n619 = ( n542 ) | ( n201 ) ;
 assign n621 = ( n138 ) | ( n276 ) ;
 assign n622 = ( n442 ) | ( n567 ) ;
 assign n620 = ( n621  &  n226  &  n238  &  n196  &  n172  &  n239  &  n7  &  n622 ) ;
 assign n623 = ( n531 ) | ( n538 ) ;
 assign n624 = ( n179 ) | ( n560 ) ;
 assign n625 = ( n534 ) | ( n166 ) ;
 assign n626 = ( n407 ) | ( n541 ) ;
 assign n627 = ( n139 ) | ( n575 ) ;
 assign n628 = ( n138 ) | ( n429 ) ;
 assign n629 = ( n139 ) | ( n455 ) ;
 assign n630 = ( n139 ) | ( n154 ) ;
 assign n631 = ( n568 ) | ( n150 ) ;
 assign n632 = ( n39  &  (~ n305)  &  (~ n310)  &  n314  &  n316  &  n382 ) ;
 assign n633 = ( n411 ) | ( n575 ) ;
 assign n634 = ( n323 ) | ( n248 ) ;
 assign n635 = ( n194 ) | ( n323 ) | ( (~ n453) ) ;
 assign n636 = ( n536 ) | ( n399 ) ;
 assign n637 = ( n190 ) | ( n127 ) ;
 assign n638 = ( n194 ) | ( n542 ) ;
 assign n639 = ( n323 ) | ( n191 ) ;
 assign n641 = ( n214  &  n680 ) | ( (~ n306)  &  n680 ) | ( n531  &  n680 ) ;
 assign n642 = ( n549 ) | ( n442 ) ;
 assign n643 = ( n190 ) | ( n116 ) ;
 assign n645 = ( n139 ) | ( n400 ) ;
 assign n646 = ( n416 ) | ( n560 ) ;
 assign n647 = ( n407 ) | ( n543 ) ;
 assign n649 = ( i_2_ ) | ( n532 ) ;
 assign n648 = ( n387  &  n628  &  n649  &  n379 ) ;
 assign n650 = ( n411 ) | ( n195 ) ;
 assign n651 = ( n195 ) | ( n166 ) ;
 assign n652 = ( n399 ) | ( n567 ) ;
 assign n653 = ( n399 ) | ( n580 ) ;
 assign n654 = ( n97  &  n233  &  n704  &  n616  &  n499  &  n685  &  n271 ) ;
 assign n656 = ( n429 ) | ( n580 ) ;
 assign n657 = ( n429 ) | ( n277 ) ;
 assign n655 = ( n16  &  n14  &  n656  &  n657  &  n591 ) ;
 assign n658 = ( n319 ) | ( n595 ) ;
 assign n659 = ( i_5_ ) | ( n194 ) | ( n512 ) ;
 assign n660 = ( n529 ) | ( n407 ) ;
 assign n661 = ( n277 ) | ( n153 ) ;
 assign n662 = ( n756  &  n12  &  n141 ) ;
 assign n663 = ( n138 ) | ( n442 ) ;
 assign n664 = ( n194 ) | ( n438 ) ;
 assign n665 = ( n156 ) | ( n139 ) ;
 assign n666 = ( n172  &  n197  &  n679  &  n15  &  n659  &  n96 ) ;
 assign n667 = ( n529 ) | ( n411 ) ;
 assign n668 = ( n429 ) | ( n576 ) ;
 assign n669 = ( n740  &  n637  &  n586  &  n192  &  n385  &  n709  &  n588 ) ;
 assign n670 = ( n106  &  n104  &  n651  &  n395  &  n270  &  n160  &  n342  &  n757 ) ;
 assign n672 = ( n658  &  n435  &  n633 ) ;
 assign n673 = ( n678  &  n725  &  n676  &  n638  &  n603  &  n605 ) ;
 assign n674 = ( n141  &  n227  &  n110  &  n6  &  n704  &  n756 ) ;
 assign n675 = ( n388  &  n177  &  n558  &  n377  &  n352  &  n634 ) ;
 assign n676 = ( n399 ) | ( n438 ) ;
 assign n677 = ( n166 ) | ( n552 ) ;
 assign n678 = ( n442 ) | ( n430 ) ;
 assign n679 = ( n429 ) | ( n457 ) ;
 assign n680 = ( n429 ) | ( n154 ) ;
 assign n681 = ( n407 ) | ( n167 ) ;
 assign n682 = ( n194 ) | ( n441 ) ;
 assign n683 = ( n156 ) | ( n411 ) ;
 assign n684 = ( n194 ) | ( n488 ) ;
 assign n685 = ( n429 ) | ( n541 ) ;
 assign n686 = ( n275 ) | ( n564 ) | ( n433 ) ;
 assign n687 = ( n166 ) | ( n277 ) ;
 assign n688 = ( n233  &  n616  &  n13 ) ;
 assign n689 = ( n166 ) | ( n457 ) ;
 assign n690 = ( n542 ) | ( n439 ) ;
 assign n691 = ( (~ i_3_) ) | ( n442 ) | ( (~ n453) ) ;
 assign n692 = ( n665  &  n262  &  n628  &  n660  &  n636  &  n635  &  n600 ) ;
 assign n693 = ( n275 ) | ( n408 ) ;
 assign n694 = ( n275 ) | ( n538 ) ;
 assign n695 = ( n539 ) | ( n189 ) ;
 assign n698 = ( n166 ) | ( n579 ) ;
 assign n699 = ( n407 ) | ( n533 ) | ( n337 ) ;
 assign n700 = ( n200 ) | ( n364 ) ;
 assign n701 = ( n275 ) | ( n200 ) | ( n467 ) ;
 assign n702 = ( n541 ) | ( n442 ) ;
 assign n703 = ( n288 ) | ( n547 ) ;
 assign n704 = ( n429 ) | ( n542 ) ;
 assign n705 = ( n149 ) | ( n551 ) ;
 assign n706 = ( n151 ) | ( n373 ) ;
 assign n707 = ( n166 ) | ( n438 ) ;
 assign n708 = ( n194 ) | ( n315 ) ;
 assign n709 = ( n323 ) | ( n594 ) ;
 assign n710 = ( n112  &  n429 ) | ( n112  &  n179 ) | ( n112  &  n280 ) ;
 assign n711 = ( n429 ) | ( n552 ) ;
 assign n712 = ( (~ i_7_) ) | ( n204 ) | ( n279 ) ;
 assign n713 = ( n528 ) | ( n139 ) | ( n354 ) ;
 assign n716 = ( n645  &  n197  &  n95  &  n685  &  n677  &  n572  &  n175 ) ;
 assign n717 = ( n543 ) | ( n578 ) ;
 assign n718 = ( n411 ) | ( n200 ) | ( n550 ) ;
 assign n719 = ( n119  &  n295 ) | ( n119  &  n399 ) | ( n119  &  n546 ) ;
 assign n720 = ( n138 ) | ( n275 ) ;
 assign n721 = ( (~ i_7_)  &  n682 ) | ( n179  &  n682 ) | ( n208  &  n682 ) ;
 assign n722 = ( n323 ) | ( n544 ) ;
 assign n723 = ( n115 ) | ( n317 ) ;
 assign n724 = ( (~ i_3_) ) | ( i_5_ ) | ( n279 ) | ( n399 ) ;
 assign n725 = ( n407 ) | ( n156 ) ;
 assign n728 = ( n335  &  n724 ) | ( (~ n453)  &  n724 ) | ( n531  &  n724 ) ;
 assign n729 = ( n127 ) | ( n297 ) ;
 assign n730 = ( i_7_ ) | ( n204 ) | ( (~ n453) ) ;
 assign n732 = ( n275 ) | ( n184 ) | ( n186 ) ;
 assign n731 = ( n732  &  n403 ) | ( n732  &  n326 ) ;
 assign n733 = ( n139 ) | ( n441 ) ;
 assign n734 = ( n531 ) | ( n184 ) | ( n483 ) ;
 assign n735 = ( n687  &  n186 ) | ( n687  &  n427 ) ;
 assign n736 = ( n439  &  n179 ) | ( n154  &  n179 ) | ( n439  &  n180 ) | ( n154  &  n180 ) ;
 assign n737 = ( n528  &  n275 ) | ( n153  &  n275 ) | ( n528  &  n190 ) | ( n153  &  n190 ) ;
 assign n738 = ( n531  &  n149 ) | ( n433  &  n149 ) | ( n531  &  n125 ) | ( n433  &  n125 ) ;
 assign n740 = ( n319 ) | ( n191 ) ;
 assign n741 = ( n552 ) | ( n153 ) ;
 assign n739 = ( n514  &  n108  &  n740  &  n741 ) ;
 assign n743 = ( i_8_ ) | ( n214 ) | ( n483 ) ;
 assign n742 = ( n743  &  n199 ) | ( n743  &  n354 ) | ( n743  &  n399 ) ;
 assign n744 = ( i_3_  &  n742 ) | ( n442  &  n742 ) | ( (~ n453)  &  n742 ) ;
 assign n745 = ( n194 ) | ( (~ n306) ) | ( n535 ) ;
 assign n746 = ( n468  &  n466 ) | ( n411  &  n466 ) | ( n468  &  n200 ) | ( n411  &  n200 ) ;
 assign n747 = ( n153  &  n531 ) | ( n510  &  n531 ) | ( n153  &  n543 ) | ( n510  &  n543 ) ;
 assign n748 = ( n747  &  n416 ) | ( n747  &  n738  &  n737 ) ;
 assign n750 = ( (~ i_0_) ) | ( (~ i_2_) ) | ( (~ i_7_) ) | ( n323 ) ;
 assign n749 = ( n254  &  n46  &  n750  &  n366  &  n129  &  n40 ) ;
 assign n751 = ( n190  &  (~ n306) ) | ( n190  &  n478 ) | ( (~ n306)  &  n595 ) | ( n478  &  n595 ) ;
 assign n752 = ( n481 ) | ( n149 ) ;
 assign n753 = ( n354 ) | ( n166 ) | ( n550 ) ;
 assign n754 = ( n535  &  n407 ) | ( n399  &  n407 ) | ( n535  &  n190 ) | ( n399  &  n190 ) ;
 assign n755 = ( n369  &  n269  &  n683 ) ;
 assign n756 = ( i_4_ ) | ( i_6_ ) | ( n512 ) ;
 assign n757 = ( n173  &  n163  &  n700  &  n121  &  n741  &  n228 ) ;
 assign n758 = ( n142  &  n536 ) | ( n142  &  n194 ) ;
 assign n759 = ( (~ i_2_) ) | ( (~ i_5_) ) | ( n762 ) | ( n763 ) ;
 assign n760 = ( i_3_ ) | ( n416 ) | ( n578 ) ;
 assign n761 = ( n482 ) | ( n568 ) ;
 assign n762 = ( i_1_  &  i_4_ ) | ( i_1_  &  n189 ) ;
 assign n763 = ( (~ i_1_)  &  (~ i_4_) ) | ( (~ i_1_)  &  n166 ) ;


endmodule

